module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g18881, g23612, g23652, g73, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29219, g29220, g29221, g30327, g30331,
         g30332, g31656, g31665, g34435, g34839, g36, g44, g53, g54, g56, g57,
         g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6753,
         g84, g90, g91, g92, g99, test_so10, test_so26, test_so35, test_so39,
         test_so42, test_so44, test_so46, test_so80, test_so86, test_so92,
         test_so100, g34783, n2730, n4896, n4895, n4837, n4921, n4920, n5045,
         g559, n4959, g33046, g5057, n5615, g34441, g2771, n5544, g33982,
         g1882, g34007, g2299, Tj_TriggerIN1, g24276, g4040, n5530, g30381,
         g2547, n5782, Tj_TriggerIN2, g30405, g3243, Tj_TriggerIN3, g25604,
         g452, Tj_TriggerIN4, g30416, g3542, Tj_TriggerIN5, g30466, g5232,
         Tj_TriggerIN6, g25736, g5813, Tj_TriggerIN7, g34617, Tj_TriggerIN8,
         g33974, g1744, g30505, g5909, Tj_TriggerIN9, g33554, g1802, n5536,
         g30432, g3554, Tj_TriggerIN10, g33064, g6219, n5385, g34881, g807,
         n5479, g6031, g24216, g847, n5709, g24232, n9367, DFF_24_n1, g34733,
         g4172, n5493, g34882, g4372, g33026, g3512, g31867, n5471, g25668,
         g3490, n5454, g24344, n5432, g4235, g33966, g1600, g33550, g1714,
         n5460, g30393, g3155, n5366, g29248, g2236, g4571, g4555, g24274,
         g3698, g33973, g1736, g30360, g1968, n5664, g34460, g30494, g5607,
         g30384, g2657, n5316, g24340, n5439, g29223, g490, n5708, g26881,
         g311, n5317, g34252, g772, n5334, g30489, g5587, g29301, g6177, n5874,
         g6377, g33022, g3167, n5652, g30496, g5615, g33043, g4567, g29263,
         g30533, g6287, g24256, n5302, g34015, g2563, g34031, g4776, n5707,
         g34452, g4593, n5303, g34646, g6199, n5644, g34001, g2295, g25633,
         g1384, g24259, g1339, n5381, g33049, g5180, n5384, g34609, g2844,
         g31869, g1024, g30490, g30427, g3598, g21894, g4264, g33965, g767,
         n5333, g34645, g5853, n5499, g33571, g2089, g34267, g4933, g26971,
         g4521, n5752, g34644, g5507, n5643, g30534, g6291, g33535, g294,
         n5680, g30498, g25728, g25743, g25684, g3813, g25613, g562, g34438,
         g608, n5475, g24244, g1205, n5547, g30439, g3909, g30541, g6259,
         g30519, g5905, g25621, g921, g34807, g2955, g25599, g203, g24235,
         g34036, g4878, n5283, g30476, g5204, g30429, g3606, g32997, g1926,
         n5510, g33063, g6215, n5651, g30424, g3586, g32977, g291, n5679,
         g34026, g4674, n5440, g30420, g3570, g33560, g29226, g676, n5751,
         g25619, g843, g34455, g4332, n5540, g30457, g4153, g33625, g6336,
         n5592, g34790, g622, n5672, g30414, g3506, n5576, g26966, g4558,
         g25656, g3111, g30390, g25688, g34727, g939, n5415, g278, n5627,
         g26963, g4492, g34034, g4864, n5318, g33541, g1036, g28093, g24236,
         g1178, g30404, g3239, g28051, g718, g29303, g6195, g26917, g1135,
         n5328, g33624, g6395, n5396, g24337, g34911, g554, g33963, g496,
         g34627, g3853, n5641, g29282, g5134, n5807, g25676, g33013, g2485,
         n5509, g32981, g925, n5725, g34976, n9357, DFF_150_n1, g30483, g5555,
         g32994, g1798, n5833, g28070, g34806, g2941, g30453, g3905, g33539,
         g763, n5332, g30526, g6255, g4375, g34035, g4871, n5443, g34636,
         g4722, n5345, g32978, g590, n5472, g30348, g1632, n5836, g24336,
         n5438, g3100, g24250, g29236, g1437, g29298, g6154, n5747, g1579,
         g30499, g5567, g33976, g1752, n5797, g32996, g1917, g30335, g744,
         n5470, g34637, g4737, n5867, g25694, DFF_178_n1, g30528, g6267,
         g24251, g1442, g30521, g26960, g4477, n5849, g24239, g34259, g4643,
         n5382, g30474, g5264, n5703, g33016, g2610, g34643, g5160, n5498,
         g30510, g5933, g29239, g1454, g26897, g753, g34729, g1296, g34625,
         g3151, n5495, g24353, g6727, n5531, g33029, g3530, n5569, g33615,
         g4104, g24253, g1532, g24281, g33997, n9352, g34971, n9351,
         DFF_206_n1, g34263, g4754, n5877, g24237, g1189, n5642, g33584, g2287,
         n5353, g24280, g4273, n5764, g26920, g1389, g33548, g29296, g5835,
         n5663, g30338, g1171, n5363, g21895, g4269, n5763, g33588, g2399,
         n5762, g34041, g4983, n5367, g30495, g5611, g29279, g4572, g25655,
         g3143, n5882, g34795, g2898, g24269, g3343, g30403, g3235, g33042,
         g30419, g3566, g34023, n9348, g28090, g4961, n5770, g34642, g4927,
         n5879, g30370, g2259, n5419, g34448, g2819, n5609, g26946, g5802,
         g34610, g2852, g24209, g417, n5358, g28047, g681, g24206, g437,
         g26891, g30504, g5901, g34798, g2886, g25669, g3494, n5889, g30480,
         g5511, n5575, g33027, g3518, n5645, g33972, g1604, g25697, g5092,
         g28099, g4831, g26947, g4382, n5714, g24350, g6386, g24210, g479,
         g30455, g3965, g28084, g33993, g2008, g736, g30444, g3933, g33537,
         g222, g25650, g3050, n5998, g25625, g1052, g30366, g2122, n5784,
         g33593, g2465, n5523, g30502, g5889, g33036, g4495, g25595, g34462,
         g33024, g3179, n5390, g33552, g1728, n5352, g34014, g2433, g29273,
         g3835, n5662, g25748, g6187, n5453, g34638, g4917, n5408, g30341,
         g1070, g26899, g822, n5422, g30336, g914, n5560, g5339, g26940, g4164,
         g25622, g34447, g2807, n5379, g33613, g4054, n5395, g25749, g6191,
         n5888, g25704, g5077, n5455, g33053, g5523, n5647, g3680, g30555,
         g6637, g25601, g174, n5402, g33971, g1682, g26892, g355, g1087,
         g26915, g1105, n5478, g33008, g30538, g6307, g3802, g25750, g6159,
         g30369, g2255, n5414, g34446, g2815, n5404, g29230, g911, n5559, g43,
         g33975, g1748, g30497, g5551, g30418, g3558, g25721, g5499, n5885,
         g34622, g30438, g3901, g34266, g4888, n5863, g30540, g6251, g32986,
         g1373, g25648, g33960, g157, n5678, g34442, g2783, n5403, g4281,
         g30421, g3574, g33573, g2112, g34730, g1283, n5635, g24205, g4297,
         n5698, g32979, g758, n5331, g4639, n5727, g25763, g6537, n5884,
         g30481, g5543, g30517, g5961, g30539, g6243, g34880, n9340, g24242,
         n5654, g30436, g29265, g3476, n5786, g32990, g1664, g24245, g1246,
         n5756, g30553, g6629, g26907, g246, n6008, g24278, g4049, g26955,
         g24282, g2932, g4575, g31894, g4098, n5350, g33037, g4498, g26894,
         g528, n5327, g34977, n5477, g25654, g3139, n5447, g33962, g34451,
         g4584, n5539, g34250, g142, n5724, g29295, g5831, g26905, g239,
         g25629, g1216, n5442, g34792, g2848, g25703, g5022, g32983, g1030,
         g30402, g3231, g25757, g1430, n9336, g33999, g2241, g24262, g1564,
         g25729, g6148, g30558, g6649, g34781, g110, g26901, g225, n5597,
         g26961, g33039, g4504, g33059, g5873, n5388, g31899, g5037, n5611,
         g33007, g2319, n5375, g25720, g5495, n5446, g21891, g30462, g5208,
         g30487, g5579, g33058, g5869, n5649, g24261, g1589, n5755, g25730,
         g5752, n5996, g30531, g6279, g30506, g34804, g2975, n5750, g25747,
         g6167, n5430, n5701, g33601, g2599, n5524, g26922, g1448, n5343,
         g29250, g2370, g30459, g5164, n5570, g1333, n5616, g33534, g153,
         n5677, g30543, g6549, n5571, g29275, g4087, n5480, g34030, g34980,
         g2984, n5842, g30451, g3961, g25627, g962, n5630, g34657, g101,
         g30552, g6625, g34979, n9332, DFF_420_n1, g30337, g1018, g24254,
         g24277, g4045, g29237, g1467, g30378, g2461, n5840, g33019, n5300,
         g33623, g5990, n5589, g29235, g1256, n5558, g31902, g5029, n5601,
         g29306, g6519, n5806, g25689, g4169, n5729, g33978, g1816, g26970,
         g4369, g4578, g34253, g4459, n5765, g29272, g3831, n5872, g33595,
         g2514, g33610, g3288, n5400, g33589, g34605, g2145, n5307, g30350,
         g1700, n5417, g25611, g513, n5548, g2841, n5963, g33619, g5297, n5588,
         g34022, g2763, g34033, g4793, n5368, g34726, g952, g31870, g1263,
         n5674, g33985, g1950, g29283, g5138, n5871, g34003, g2307, g25677,
         g34463, g4664, g33006, g2223, g29292, g5808, n5749, g30557, g6645,
         g33989, g2016, g33033, g3873, n5387, n5699, g34005, g2315, g26932,
         g2811, g30516, g5957, g33575, g2047, g33032, g30486, g5575, g34974,
         n9327, DFF_477_n1, g25678, g3752, n5994, g30440, g3917, g1585, n5757,
         g26949, g4388, g30530, g6275, g30542, g6311, g25624, g1041, g30383,
         g33597, g2537, g34598, g26957, g4430, g26967, n9325, g28102, g4826,
         g30524, g6239, g26903, g232, g30475, g5268, g34647, g6545, n5497,
         g30377, n9324, g33553, g1772, n5504, g31903, g5052, n5607, g25715,
         g33984, g1890, g33602, g2629, n5521, g28045, g572, n5337, g34603,
         g2130, n5487, g33035, g4108, n5715, g4308, g24208, g475, g990, n5622,
         g31, n5469, g34970, n9322, DFF_514_n1, g33614, g3990, n5594, g33060,
         g30362, g1992, g33023, g3171, n5603, g26898, g812, n5733, g25618,
         g832, g30518, g5897, g4570, n5702, g26959, g4455, g34801, g2902,
         g26884, g333, g25600, g168, n5606, g26933, g28066, g3684, g33612,
         g3639, n5591, g24268, g3338, n5527, g25716, g5406, n5992, g26906,
         g269, g24203, g401, g24346, g6040, g24207, g441, g25701, n5690,
         g29269, g3808, n5745, g9, n5468, g34255, g30450, g3957, g30456, g4093,
         n5340, g32991, g1760, n5602, g24348, n5437, g34249, g160, n5843,
         g30371, g2279, n5778, g29268, g3498, g29224, g586, n5336, g33017,
         g2619, n5508, g30339, g1183, n5599, g33967, g1608, g33559, g1779,
         g29255, g2652, g30368, g2193, n5839, g30375, g2393, n5421, g28052,
         g661, g28089, g4950, n5772, g33055, g5535, n5566, g30392, g2834,
         g30343, g1361, g30523, g6235, g24233, g1146, n5851, g33018, g32976,
         g150, n5676, g30349, g1696, n5628, g33067, g6555, g26900, g33034,
         g3881, n5564, g30551, g6621, g25667, g3470, n5424, g30452, g3897,
         g34719, g518, g538, g33607, g2606, g26923, g1472, n5290, g24211,
         g33050, g5188, n5567, g24341, g5689, n5529, g24201, g405, g30463,
         g5216, g6494, g34464, g4669, g24243, g996, g24335, g4531, g34611,
         g2860, g34262, g4743, g30546, g6593, g25591, g4411, g30347, g1413,
         g30556, g6641, g6, g33562, g1936, n5534, g55, g25610, g504, n5519,
         g33015, g2587, n5372, g31896, g4480, g34004, n9314, g30428, g30485,
         g5571, g30422, g3578, g25714, g29294, g5827, n5809, g30423, g3582,
         g30529, g6271, g34028_Tj_Payload, g4688, n5656, g33587, g2380, g30460,
         g5196, g30401, g3227, g33990, n9312, g29309, g6541, g30411, g3203,
         g33546, g1668, n5598, g28085, g4760, n5775, g26904, g262, g33556,
         g1840, n5451, g25722, g5467, g25605, g460, g33062, g6209, g26893,
         n5704, g28050, g655, g34626, g33583, g2204, n5620, g30472, g5256,
         g34454, g4608, n5274, g34850, g794, n5291, g4423, g24272, g3689,
         n5532, g5685, g24214, g703, n5821, g26909, g862, n5682, g30406, g3247,
         g33569, g2040, n5505, DFF_672_n1, g34628, g4146, n5981, g34458, g4633,
         n5844, g24240, n5304, g34634, g4732, n5296, g25700, n5689, g29293,
         g5817, g33009, g2351, n5511, g33603, g2648, g24355, g6736, g34268,
         g4944, n5875, g25691, g4072, g26890, g29264, g3466, g28072, g4116,
         g31900, g5041, n5605, g26956, g4434, g29271, g3827, n5808, g29304,
         g6500, n5748, g29261, g3133, n5661, g28063, g3333, g979, n5320,
         g34027, g4681, g33961, g298, n5675, g33604, g32995, g1894, n5374,
         g34624, g2988, g30415, g3538, g33536, g301, g26888, n9306, DFF_709_n1,
         g28055, g827, n5728, g24238, g33600, g2555, n5351, g28105, g5011,
         g34721, g199, g29307, g6523, n5870, g30345, g34453, g4601, n5365,
         g32980, g854, g29238, g1484, n5865, g34639, g4922, n5346, g25695,
         g5080, n5893, g33057, g5863, g26969, g4581, n5670, g29253, g2518,
         g34021, g2567, g26895, g568, n5335, g30413, g3263, g30549, g6613,
         g24347, g25758, g6444, n5990, g34808, g2965, g30501, g5857, n5573,
         g33969, n9303, g34440, g890, n5305, g30433, g3562, g21900, g26921,
         g1404, g29270, g3817, n9302, n6010, g33038, g4501, g31865, g26926,
         g2724, n5301, g28083, g4704, n5771, g34797, g22, g2878, g30478, g5220,
         g34724, g617, n5339, g24212, g26883, g316, g32985, g1277, g25761,
         g6513, n5426, g26886, g336, n5824, g34796, g2882, g32982, g33561,
         g1906, n5503, g26880, g305, n5282, g34975, g8, g26931, g2799, g34641,
         g4912, n5297, g34629, g4157, n5983, g33598, g2541, n5461, g33576,
         g2153, n5356, g34720, g550, g26902, g255, g29244, g30468, g5240,
         g26924, g1478, n5289, g33031, g3863, g29245, g1959, g29266, g3480,
         n5868, g30559, g6653, g34794, g2864, n5489, g28087, g4894, n5774,
         g30435, g3857, n5572, g25609, g28057, g1002, g34439, g776, n5330, g28,
         n5324, g1236, g34260, g4646, n5712, g33012, g2476, g32989, g1657,
         n5525, g34006, g2375, g63, g358, g26910, g896, n5431, g28043, g33021,
         g3161, g29251, g2384, n5700, g34456, g4616, n5608, g26968, g4561,
         g33991, g2024, g3451, g26930, g2795, g34599, g613, n5474, g28082,
         g4527, g33557, g1844, g30511, g5937, g33045, g30379, g2523, n5281,
         g24267, n5436, g34020, g2643, g24249, g1489, n5850, g25592, g30382,
         n9295, g29285, g5156, n5526, n9294, DFF_829_n1, g25662, g21896,
         g33563, g1955, g33622, g33582, g2273, n5458, g28086, g4771, n5769,
         g25744, g6098, n5988, g29262, g3147, g24270, g3347, g33581, g2269,
         g191, g24266, g2712, g34849, g626, n5288, g33618, g2729, g5357, n5393,
         g34038, g34032, g4709, n5518, g34803, g2927, g34459, g4340, n5653,
         g30509, g5929, g34640, g4907, n5295, g28069, g4035, g21899, g2946,
         g31868, g918, n5673, g26938, g4082, g25756, g30363, g30334, g577,
         n5294, g33970, g1620, g30391, g2831, g25615, g667, g33540, g930,
         n5731, g30445, g3937, g25617, g817, n5822, g24247, g1249, g24215,
         g837, n5562, g33964, g599, n5550, g25719, g5475, n5425, g29228,
         g30514, g5949, g33627, g6682, n5590, g24231, g904, g34615, g2873,
         n5488, g30356, g1854, n5785, g25696, g5084, n5681, g30493, g5603,
         n5726, g33594, g2495, n5522, g34009, g2437, g30365, g2102, n5666,
         g33004, g2208, g34018, g25685, g4064, n5416, g34040, g4899, n5517,
         g25639, g2719, n5465, g34029, g4785, n5361, g30488, g5583, g34600,
         g781, n5551, g29300, g6173, n5810, g34802, g2917, g25614, g686,
         g28058, g1252, n5554, g29225, g671, g33580, g30532, g6283, g33054,
         g5527, n5389, g26962, g4489, g33564, g1974, n5450, g32984, g1270,
         n5716, g34039, g4966, n5706, g33065, g6227, n5568, g30443, g3929,
         g29291, g5503, g24279, g30508, g5925, g29232, g1124, g34269, g4955,
         n5614, g30464, g5224, g33988, g2012, g30522, g6203, n5574, g25708,
         g5120, g30374, g2389, n5631, g26953, g4438, g34008, g2429, g34444,
         g2787, n5610, g34731, g33606, g2675, n5457, g24334, n5541, g34265,
         g4836, n5713, g30340, g1199, g24257, n5401, g30482, g5547, g34604,
         g2138, n5275, g33591, g2338, g30525, g6247, g26929, g2791, g30448,
         g34602, g1291, n2549, g30513, g5945, g30469, g5244, g33608, g2759,
         g33626, g6741, n5398, g34725, g785, n5293, g30342, g1259, n5553,
         g29267, g3484, n5668, g25593, g209, n5595, g30548, g6609, g33052,
         g5517, g34012, g2449, g34017, n9281, g24263, g2715, n5299, g26912,
         g936, n5557, g30364, g2098, n5280, g34254, g4462, n5671, g34251, g604,
         n5473, g30560, g6589, g33983, n9280, g24204, g429, g33980, g1870,
         g34631, g29243, g1825, g25623, g1008, n5321, g26950, g4392, n5710,
         g30431, g3546, g30467, g5236, g30353, g1768, n5834, g34467, g4854,
         g30442, g3925, g29305, g6509, g25616, g732, n5732, g29252, g2504,
         g4519, g4520, g33003, g2185, n5376, g34613, g37, g4031, g33570, g2070,
         n5535, g34734, g4176, n5494, g24275, n5435, g4405, g872, g29302,
         g6181, n5667, g24349, g34264, g4765, n5613, g30484, g5563, g25634,
         g1395, g33567, g1913, g33585, g2331, n5513, g30527, g6263, g34978,
         n9276, DFF_1012_n1, g30447, g3945, g347, n5860, g34256, g4473, g25630,
         g1266, g29290, g5489, n5660, g29227, g31872, g2748, n5516, g29287,
         g5471, g31897, g4540, g6723, g30562, g6605, g34011, n9274, g33996,
         g2173, g21898, g33014, g2491, g34465, g4849, g33995, g2169, g30372,
         n9273, g30545, g30389, g33590, g2407, n5459, g34616, g2868, g26927,
         g2767, g32992, g1783, n5596, g25631, g1312, n5466, g30477, g5212,
         g34632, g4245, n5640, g28046, g645, g4291, g26896, g25602, g26916,
         g1129, n5329, g33578, g2227, n5538, g33579, g2246, g30354, g1830,
         n5413, g30425, g3590, g24200, g392, g33544, g1592, n5362, g25764,
         g6505, g24246, g1221, g30507, g5921, g26889, g30333, g218, g32998,
         g1932, g32987, g1624, n5370, g25702, g5062, g29286, g5462, n5744,
         g34606, g2689, n5347, g33070, g6573, n5563, g29240, g1677, g32999,
         g2028, n5371, g33605, g2671, g24255, g26945, g33558, g1848, n5464,
         g25699, n5669, g29289, g5485, n5869, g30388, g2741, n5349, n5482,
         g29254, g2638, g28074, g4122, g34450, g4322, n5506, g30512, g5941,
         g33572, g2108, n5452, g25, g33551, g33538, g595, n5476, g33005, g2217,
         n5512, g24248, n9267, DFF_1092_n1, g33002, g2066, n5832, g24234,
         g1152, n5618, g30471, g5252, g34000, g2165, g34016, g2571, g33048,
         g5176, n5650, g25628, g26934, g2827, g34468, g4859, g24202, g424,
         g33542, g1274, n5730, n9265, g34445, g2803, n5545, g33555, g1821,
         g34013, g2509, g28091, g5073, g26919, n5556, g30554, g6633, g29281,
         g5124, g30537, g6303, g28092, g5069, g34732, g2994, n5634, g28049,
         g650, g33545, g1636, n5549, g30441, g3921, g29247, g24354, g6732,
         g25636, g1306, n5796, g26914, g1061, g25670, g3462, g33998, g2181,
         g25626, g956, n5341, g33977, g1756, g29297, g5849, g28071, g4112,
         g30387, n9262, g33577, g2197, n5514, g33592, g26913, g1046, g28044,
         g482, n5820, g26948, g4401, g30344, g1514, n5364, g26885, g329, n5766,
         g33069, g6565, n5386, g34621, g2950, g28059, g1345, g25762, g6533,
         n5445, g34633, g4727, n5312, g24352, g26925, g1536, g30446, g3941,
         g25597, g370, g24342, g5694, g30357, g1858, n5892, g26908, g446,
         g30399, g3219, g29242, g1811, g30547, g6601, g34010, g2441, g33986,
         g1874, g34257, g30544, g6581, g30561, g6597, g5008, n5637, g30430,
         g3610, g34799, g2890, g33565, g1978, g33968, g1612, g34843, g112,
         g34793, g2856, g33566, g1982, n5462, g30465, g28073, g4119, g24351,
         g6390, g30346, g1542, g21893, g4258, g4818, n5636, g31904, g5033,
         g34635, g4717, n5344, g25637, g1554, n5768, g29274, g3849, g30396,
         g3199, g25735, g34037, g4975, n5360, g34791, g790, n5292, g30520,
         g5913, g30358, g1902, n5837, g29299, g6163, g25690, g4125, g28096,
         g4821, g28088, g4939, n5776, g24241, n5392, g30397, g3207, g4483,
         g30409, g29284, g5142, n5658, g30470, g5248, g30367, g2126, g24273,
         g3694, g29288, g5481, n5805, g30359, g1964, n5315, g25698, g5097,
         n5753, g30398, g3215, n9255, g26952, g4427, g26928, g2779, n5694,
         g26954, DFF_1225_n1, g30351, g1720, n5780, g31871, g1367, g5112, g19,
         g26939, g4145, g33994, g2161, g25596, g376, n5633, g33586, g2361,
         n5537, g21901, g31866, g582, n5552, g33000, g2051, g26918, g1193,
         g30373, g2327, n5841, g28056, g907, n5555, g34601, g947, n5286,
         g30355, g1834, n5665, g30426, g3594, g34805, g2999, g34002, g2303,
         g28053, g29229, g723, n5826, g33620, g5703, n5397, g34722, g546,
         n5492, g33599, g2472, n5619, g30515, g5953, g25649, g33979, g1740,
         g30417, g3550, g25683, g3845, n5886, g33574, g2116, n5463, g30410,
         g30454, g3913, g34024, g33547, g1687, g30386, g2681, n5777, g33596,
         g2533, n5761, g26887, g324, n5827, g34607, g2697, n5308, g31895,
         g4417, g33068, g6561, n5646, g29233, g1141, n5691, g24258, n5655,
         g30376, g33549, g1710, g29308, g6527, n5659, g30408, g3255, g29241,
         g1691, g34620, g2936, g33621, g5644, n5593, g25707, g5152, n5883,
         g24339, g5352, g34443, g2775, n5378, g34619, g2922, g29234, g30503,
         g5893, g30550, g6617, g33001, g2060, n5507, g33040, g4512, g30492,
         g5599, g25664, g3401, n5986, g26944, g4366, g34614, n5342, g29260,
         g3129, n5861, g33047, g5170, g24298, g25733, g5821, n5429, g30536,
         g6299, g29246, g2079, g34261, g4698, n5862, g33611, g3703, n5399,
         g25638, g1559, n5441, g34728, n9247, g29222, g411, n5629, g25742,
         g30449, g3953, g34608, g2704, n5377, g24345, g6035, n5528, n9245,
         g25635, g1300, n5483, g25686, g4057, n5711, g30461, g5200, g34466,
         g4843, g31901, g5046, n5578, g29249, g2250, g26882, n5456, g33041,
         g33011, g2453, n5373, g25734, g5841, n5449, n5705, g34618, g2912,
         g33010, g2357, g31864, g164, n5561, g34630, g4253, n5484, g31898,
         g5016, n5369, g25653, g3119, n5423, g25632, g1351, n5322, g32988,
         g33616, g29280, g5115, n5743, g33609, g3352, n5604, g30563, g6657,
         g33044, g4552, g30437, g3893, g30412, g3211, g30491, g5595, g30434,
         g3614, g34612, g29259, g3125, n5781, g25681, g3821, n5428, g25687,
         g4141, n5612, g33617, g30479, g5272, g29256, g2735, n5600, g28054,
         g728, g30535, g6295, g30385, g2661, n5418, g30361, g1988, n5783,
         g25705, g24260, g1548, n5546, g29257, g3106, n5742, g34461, g4659,
         g34258, g4358, n5348, g32993, g1792, n5359, g33992, g2084, g30394,
         g3187, g34449, g4311, n5323, g34019, g2583, g18597, n9240,
         DFF_1381_n1, g29231, g1094, g25682, g21897, g4284, g30395, g3191,
         g21892, g4239, g4180, n5380, g28048, g691, n5520, g34723, g534, n5490,
         g25598, g385, n5632, g33987, g2004, g30380, g2527, n5420, g5456,
         g26965, n6007, g25706, g30458, g4507, n5846, g24338, g5348, g30400,
         g3223, g34623, g2970, g24343, g5698, g30473, g5260, g24252, g1521,
         n5577, g33028, g3522, n5383, g29258, g3115, g30407, g3251, g26958,
         g34457, g33568, g1996, n5355, g25663, g26964, g4515, g34735, g4300,
         n5639, g30352, n9236, g33543, g1379, g24271, n5433, g33981, g1878,
         g30500, g5619, g34649, g71, g29277, g25612, n5287, g28060, n2505,
         n2499, n2668, n3160, n3102, g72, n5960, n4689, n5961, n4708, n3593,
         n3589, n3595, n3574, n3570, n3576, n3517, n3513, n3519, n3628, n3624,
         n3630, n3555, n3551, n3557, n3646, n3642, n3648, n3536, n3532, n3538,
         n3611, n3607, n3613, n3006, n3765, n3505, n3525, n3635, n4888, n3550,
         n2595, n2527, n3524, n3005, n3623, n3549, n3003, n3007, n3569, n3606,
         n3588, n3165, n3799, n3033, n3622, n3587, n3586, n3605, n3604, n3568,
         n3567, n3548, n3512, n3511, n3531, n3530, n3641, n3640, n3131, n3111,
         n4537, n4201, n3745, n3684, n3274, n2982, n2706, n2649, n2556, n2509,
         n2487, n2427, n2423, n2421, n4172, n4173, n4190, n4191, n4388, n4210,
         n3951, n3774, n3842, n3808, n3908, n3984, n3875, n4015, n3914, n3780,
         n3957, n3848, n3990, n3814, n3881, n4022, n4027, n3785, n3962, n3853,
         n3886, n3819, n3995, n3919, n3682, n3272, n2980, n2704, n2647, n2554,
         n2507, n2485, n2425, n2419, n2405, n2760, n2552, n4946, n2404, n3653,
         n4962, n4948, n3195, n2774, n3116, n4945, n4525, n4518, n3281, n3277,
         n3276, n2989, n2991, n3687, n2710, n2707, n3174, n3362, n2644, n3146,
         n3115, n3833, n3023, n3933, n3729, n3664, n3662, n3673, n3671, n3506,
         n2790, n4490, n4178, n4514, n4196, n3736, n3741, n2598, n4519, n2594,
         n3084, n2590, n4722, n3125, n3105, n3145, n3164, n2422, n4037, n4034,
         n4039, n3972, n3969, n3929, n3926, n3863, n3860, n4003, n4002, n4032,
         n4035, n3797, n3792, n3790, n3795, n3891, n3893, n3827, n3826, n3896,
         n4007, n3931, n3793, n3924, n3831, n3829, n3927, n3974, n3898, n3970,
         n4000, n3865, n3861, n3824, n3894, n3967, n3858, n4005, n3395, n4956,
         n5026, n3941, n3733, n4798, n4805, n4175, n4193, n3738, n4721, n4523,
         n4524, n4526, n2573, n2577, n2563, n2567, n4938, n4913, n4714, n4516,
         n4517, n5111, n4819, n3730, n4305, n4283, g34028, n2608, n4447, n4448,
         n4402, n4403, n4425, n4426, n4436, n4437, n4391, n4392, n4379, n4380,
         n4414, n4415, n4458, n4459, n5016, n5014, n3064, n3065, n4535, n5112,
         n3675, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4, Tj_OUT1234, Tj_OUT5,
         test_se_NOT, Tj_Trigger, n5, n26, n43, n45, n47, n52, n54, n57, n73,
         n74, n75, n89, n90, n91, n101, n103, g33959, n176, n183, n184, n190,
         n192, n194, n199, g33533, n266, n324, n353, n408, n420, n422, n430,
         n432, n434, n439, n470, n488, n497, n498, n499, g34788, n513, n536,
         n537, n538, n540, n552, n553, n716, n725, n727, n729, n733, n757,
         n758, n759, n763, n764, n765, n822, n826, n841, n843, n845, n850,
         n869, n905, n955, n956, n957, n959, n999, n1013, g25259, n1037, n1038,
         n1039, n1107, n1108, n1109, n1178, n1179, n1180, g25167, n1205, n1266,
         n1289, n1296, n1426, n1452, n1454, n1456, n1460, n1465, n1577, n1733,
         n1774, n1835, n8330, n8333, n8336, n8337, n8339, n8340, n8355, n8356,
         n8358, n8359, n8363, n8364, n8365, n8368, n8369, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8379, n8381, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8394, n8395, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8421, n8422, n8423, n8425, n8427,
         n8431, n8433, n8435, n8436, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8446, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8460, n8462, n8463, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8479, n8480, n8481, n8484,
         n8485, n8487, n8488, n8490, n8491, n8493, n8494, n8495, n8497, n8500,
         n8502, n8503, n8505, n8507, n8509, n8511, n8512, n8513, n8514, n8547,
         n8549, n8551, n8553, n8555, n8557, n8559, n8560, n8562, n8564, n8566,
         n8568, n8569, n8571, n8573, n8575, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8593, n8598, n8600, n8605, n8608, n8611, n8614, n8617, n8629, n8643,
         n8644, n8645, n8646, n8648, n8649, n8650, n8651, n8655, n8658, n8659,
         n8660, n8662, n8663, n8664, n8665, n8667, n8668, n8669, n8670, n8672,
         n8673, n8674, n8676, n8677, n8678, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8725, n8726, n8727, n8728, n8729, n8732,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8752, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8775, n8776, n8778, n8779, n8781, n8782, n8784,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8837, n8838,
         n8839, n8842, n8843, n8844, n8845, g32975, n8847, n8848, n8849, n8850,
         n8851, n8852, g31860, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9237, n9238, n9239, n9241, n9242,
         n9243, n9244, n9246, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9256, n9257, n9258, n9259, n9260, n9261, n9263, n9264, n9266, n9268,
         n9269, n9270, n9271, n9272, n9275, n9277, n9278, n9279, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9296, n9297, n9298, n9299, n9300, n9301, n9304, n9305, n9307, n9308,
         n9309, n9310, n9311, n9313, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9323, n9326, n9328, n9329, n9330, n9331, n9333, n9334, n9335,
         n9337, n9338, n9339, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9349, n9350, n9353, n9354, n9355, n9356, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, U5116_n1, U5126_n1, U5127_n1, U5128_n1,
         U5129_n1, U5353_n1, U5355_n1, U5961_n1, U5962_n1, U5963_n1, U5964_n1,
         U5965_n1, U5966_n1, U5967_n1, U5968_n1, U6100_n1, U6211_n1, U6212_n1,
         U6213_n1, U6214_n1, U6215_n1, U6216_n1, U6217_n1, U6218_n1, U6279_n1,
         U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1, U6286_n1,
         U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1, U6338_n1,
         U6341_n1, U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1,
         U6348_n1, U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1,
         U6355_n1, U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1,
         U6362_n1, U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1,
         U6369_n1, U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1,
         U6417_n1, U6446_n1, U6465_n1, U6497_n1, U6523_n1, U6542_n1, U6552_n1,
         U6553_n1, U6554_n1, U6555_n1, U6556_n1, U6559_n1, U6560_n1, U6561_n1,
         U6570_n1, U6911_n1, U6912_n1, U6917_n1, U6926_n1, U6927_n1, U6929_n1,
         U6931_n1, U6932_n1, U6933_n1, U6934_n1, U6935_n1, U6936_n1, U6937_n1,
         U6938_n1, U6939_n1, U6940_n1, U6941_n1, U6944_n1, U6950_n1, U6954_n1,
         U6955_n1, U6956_n1, U6957_n1, U7174_n1, U7248_n1, U7249_n1, U7402_n1,
         U7405_n1, U7413_n1, U7416_n1, U7427_n1, U7438_n1, U7449_n1, U7455_n1,
         U7464_n1, U7467_n1, U7482_n1, U7492_n1, U7513_n1, U7516_n1, U7549_n1,
         U7561_n1, U7574_n1, U7577_n1, U7585_n1, U7595_n1, U7614_n1, U7621_n1,
         U7629_n1, U7636_n1, U7639_n1, U7649_n1, U7652_n1, U7668_n1, U7673_n1,
         U7690_n1, U7707_n1, U7712_n1, U7792_n1, U7794_n1, U7895_n1, U7897_n1,
         U7977_n1, U8034_n1, U8036_n1, U8050_n1, U8055_n1, U8060_n1, U8070_n1,
         U8074_n1, U8088_n1, U8112_n1, U8113_n1, U8147_n1, U8165_n1, U8185_n1,
         U8192_n1, U8210_n1, U8223_n1, U8224_n1, U8281_n1, U8307_n1, U8974_n1,
         U8975_n1, U9065_n1, U9070_n1, U9075_n1, U9076_n1, U9080_n1, U9084_n1,
         U9085_n1, U9086_n1, U9090_n1, U9098_n1, U9099_n1, U9101_n1, U9107_n1,
         U9111_n1, U9116_n1, U9120_n1, U9124_n1, U9128_n1, U9132_n1, U9136_n1,
         U9315_n1, U9453_n1, U9825_n1, U9886_n1, U9927_n1, U9953_n1, U9957_n1,
         U9958_n1, U9968_n1, U9972_n1, U9992_n1, U10314_n1, U10318_n1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g34597 = 1'b0;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g29218 = g18881;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g24167 = g73;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20557 = g29213;
  assign g20652 = g29214;
  assign g20901 = g29215;
  assign g21176 = g29216;
  assign g21270 = g29217;
  assign g20654 = g29219;
  assign g21245 = g29220;
  assign g21292 = g29221;
  assign g23002 = g30327;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g31521 = g34435;
  assign g34956 = g34839;
  assign g21698 = g36;
  assign g24185 = g44;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18101 = g6746;
  assign g18097 = g6747;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18100 = g6751;
  assign g18092 = g6753;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g31861 = test_so10;
  assign g25219 = test_so10;
  assign g13881 = test_so26;
  assign g9615 = test_so35;
  assign g8785 = test_so39;
  assign g8291 = test_so42;
  assign g17316 = test_so44;
  assign g8178 = test_so46;
  assign g12470 = test_so80;
  assign g11447 = test_so86;
  assign g9682 = test_so92;
  assign g29210 = test_so100;
  assign g20049 = test_so100;
  assign g24166 = g72;
  assign g28753 = g33959;
  assign g27831 = g33533;
  assign g33894 = g34788;
  assign g31862 = g25259;
  assign g31863 = g25167;
  assign g26801 = g32975;
  assign g25114 = g31860;

  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(n9119), .CLK(n9517), .Q(
        g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(n9088), .CLK(n9532), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(n8930), .CLK(n9611), .Q(
        g1882) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(n8930), .CLK(n9611), .Q(
        g2299), .QN(Tj_TriggerIN1) );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(n9042), .CLK(n9555), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(n9046), .CLK(n9553), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(n9046), .CLK(n9553), .Q(g559), .QN(Tj_TriggerIN2) );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(n9045), .CLK(n9553), .Q(
        g3243), .QN(Tj_TriggerIN3) );
  SDFFX1 DFF_10_Q_reg ( .D(g25604), .SI(g3243), .SE(n9091), .CLK(n9530), .Q(
        g452), .QN(Tj_TriggerIN4) );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(n9091), .CLK(n9530), .Q(
        g3542), .QN(Tj_TriggerIN5) );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(n9110), .CLK(n9521), .Q(
        g5232), .QN(Tj_TriggerIN6) );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(n8942), .CLK(n9605), .Q(
        g5813), .QN(Tj_TriggerIN7) );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(n8941), .CLK(n9606), .Q(
        test_so1), .QN(Tj_TriggerIN8) );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(n9063), .CLK(n9544), 
        .Q(g1744) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(n9018), .CLK(n9567), .Q(
        g5909), .QN(Tj_TriggerIN9) );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(n9048), .CLK(n9552), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(n8928), .CLK(n9612), .Q(
        g3554), .QN(Tj_TriggerIN10) );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(n8927), .CLK(n9613), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(n9031), .CLK(n9561), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(n9031), .CLK(n9561), .Q(
        g6031), .QN(n8683) );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(n9059), .CLK(n9546), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(n8953), .CLK(n9600), .Q(
        n9367), .QN(DFF_24_n1) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(n9080), .CLK(n9536), .Q(
        g4172), .QN(n5493) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(n9084), .CLK(n9534), .Q(
        g4372) );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(n9084), .CLK(n9534), .Q(
        g3512), .QN(n8767) );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(n9033), .CLK(n9560), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(g25668), .SI(test_si3), .SE(n8956), .CLK(n9598), 
        .Q(g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(n8918), .CLK(n9617), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(n8918), .CLK(n9617), .Q(
        g4235), .QN(n8514) );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(n9007), .CLK(n9573), .Q(
        g1600) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(n9065), .CLK(n9543), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(n8970), .CLK(n9591), .Q(
        g14451) );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(n8927), .CLK(n9613), .Q(
        g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(n8918), .CLK(n9617), .Q(
        g2236) );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(n9010), .CLK(n9571), .Q(
        g4555) );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(n9112), .CLK(n9520), .Q(
        g3698), .QN(n8582) );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(n9064), .CLK(n9544), .Q(
        g1736) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(n8984), .CLK(n9584), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(n8983), .CLK(n9584), .Q(
        test_so3), .QN(n8873) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(n9102), .CLK(n9525), 
        .Q(g5607) );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(n9102), .CLK(n9525), .Q(
        g2657), .QN(n5316) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(n8953), .CLK(n9600), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(n8947), .CLK(n9602), .Q(
        g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(n8947), .CLK(n9602), .Q(
        g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(n9032), .CLK(n9560), .Q(
        g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(n9103), .CLK(n9524), .Q(
        g5587) );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(n9099), .CLK(n9526), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(n9009), .CLK(n9571), .Q(
        g6377), .QN(n8703) );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(n9009), .CLK(n9571), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(n9098), .CLK(n9527), .Q(
        g5615) );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(n9021), .CLK(n9565), .Q(
        g4567) );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(n9091), .CLK(n9530), .Q(
        test_so4), .QN(n8891) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(n9016), .CLK(n9568), 
        .Q(g6287) );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(n8973), .CLK(n9589), .Q(
        g7946), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g7946), .SE(n9005), .CLK(n9573), .Q(
        g2563) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(n8975), .CLK(n9589), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(n8998), .CLK(n9577), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(n8998), .CLK(n9577), .Q(
        g6199), .QN(n5644) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(n8997), .CLK(n9577), .Q(
        g2295) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(n9071), .CLK(n9540), .Q(
        g1384), .QN(n8340) );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(n8974), .CLK(n9589), .Q(
        g1339), .QN(n5381) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(n8974), .CLK(n9589), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(n9043), .CLK(n9555), .Q(
        g2844) );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(n9095), .CLK(n9529), .Q(
        g1024), .QN(n8440) );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(n9102), .CLK(n9525), .Q(
        test_so5) );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(n9030), .CLK(n9561), 
        .Q(g3598), .QN(n8488) );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(n9030), .CLK(n9561), .Q(
        g4264) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(n9032), .CLK(n9560), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(n9032), .CLK(n9560), .Q(
        g5853), .QN(n5499) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(n8921), .CLK(n9615), .Q(
        g13865) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(n8991), .CLK(n9580), .Q(
        g2089), .QN(n8385) );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(n9097), .CLK(n9527), .Q(
        g4933) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(n9084), .CLK(n9534), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(n9084), .CLK(n9534), .Q(
        g5507), .QN(n5643) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(n8971), .CLK(n9591), .Q(
        g16656), .QN(n8674) );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(n9015), .CLK(n9568), .Q(
        g6291) );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(n9068), .CLK(n9542), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(n8907), .CLK(n9623), .Q(
        test_so6) );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(n8965), .CLK(n9594), 
        .Q(g9617) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(n9052), .CLK(n9550), .Q(
        g9741), .QN(n8369) );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(n9052), .CLK(n9550), .Q(
        g3813), .QN(n8409) );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(n9052), .CLK(n9550), .Q(
        g562), .QN(n8842) );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(n9050), .CLK(n9551), .Q(
        g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(n9034), .CLK(n9559), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(n9092), .CLK(n9530), .Q(
        g3909), .QN(n8608) );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(n9016), .CLK(n9568), .Q(
        g6259), .QN(n8704) );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(n8988), .CLK(n9582), .Q(
        g5905) );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(n8987), .CLK(n9582), .Q(
        g921), .QN(n8782) );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(n9117), .CLK(n9517), .Q(
        g2955) );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(n8952), .CLK(n9600), .Q(
        g203) );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(n8952), .CLK(n9600), .Q(
        test_so7), .QN(n8865) );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(n8979), .CLK(n9587), 
        .Q(g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(n8978), .CLK(n9587), .Q(
        g5204) );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(n8962), .CLK(n9595), .Q(
        g17604), .QN(n8660) );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(n8927), .CLK(n9612), .Q(
        g3606), .QN(n8673) );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(n8984), .CLK(n9584), .Q(
        g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(n8928), .CLK(n9612), .Q(
        g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(n8928), .CLK(n9612), .Q(
        g3586) );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(n9068), .CLK(n9542), .Q(
        g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(n8979), .CLK(n9586), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(n8945), .CLK(n9604), .Q(
        g3570) );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(n8945), .CLK(n9604), .Q(
        g9048), .QN(n8330) );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(n8944), .CLK(n9604), .Q(
        g17607), .QN(n8551) );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(n8935), .CLK(n9609), .Q(
        test_so8), .QN(n8861) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(n9088), .CLK(n9532), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(n8981), .CLK(n9586), .Q(
        g843), .QN(n8431) );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(n8981), .CLK(n9586), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(n9080), .CLK(n9536), .Q(
        g4153), .QN(n8819) );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(n9077), .CLK(n9537), .Q(
        g17711), .QN(n8568) );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(n9100), .CLK(n9526), .Q(
        g6336), .QN(n5592) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(n9049), .CLK(n9551), .Q(
        g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(n8972), .CLK(n9590), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(n9010), .CLK(n9571), .Q(
        g4558) );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(n9010), .CLK(n9571), .Q(
        g17685), .QN(n8678) );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(n8919), .CLK(n9617), .Q(
        g3111), .QN(n8406) );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(n9004), .CLK(n9574), .Q(
        g29217) );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g29217), .SE(n9004), .CLK(n9574), .Q(
        test_so9) );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(n9060), .CLK(n9546), 
        .Q(g939), .QN(n5415) );
  SDFFX1 DFF_128_Q_reg ( .D(n324), .SI(g939), .SE(n9069), .CLK(n9542), .Q(g278), .QN(n5627) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(n8924), .CLK(n9614), .Q(
        g4492) );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(n8979), .CLK(n9587), .Q(
        g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(n9095), .CLK(n9529), .Q(
        g1036), .QN(n8792) );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(n9029), .CLK(n9562), .Q(
        g29220) );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g29220), .SE(n9028), .CLK(n9562), .Q(
        g1178) );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(n9038), .CLK(n9557), .Q(
        g3239) );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(n8950), .CLK(n9601), .Q(
        g718), .QN(n8829) );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(n8921), .CLK(n9616), .Q(
        g6195) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(n9066), .CLK(n9543), .Q(
        g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(n8933), .CLK(n9609), .Q(
        g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(n8910), .CLK(n9621), .Q(
        test_so10), .QN(n8888) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(n8911), .CLK(n9621), 
        .Q(g554), .QN(n8427) );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(n9107), .CLK(n9522), .Q(
        g496) );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(n9107), .CLK(n9522), .Q(
        g3853), .QN(n5641) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(n9107), .CLK(n9522), .Q(
        g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(n8992), .CLK(n9580), .Q(
        g17404), .QN(n8443) );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(n8917), .CLK(n9618), .Q(
        g8344) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(n9056), .CLK(n9548), .Q(
        g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(n8923), .CLK(n9614), .Q(
        g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(n9117), .CLK(n9518), .Q(
        n9357), .QN(DFF_150_n1) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(n9117), .CLK(n9518), .Q(
        g5555), .QN(n8690) );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(n9057), .CLK(n9548), .Q(
        g14096) );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(n9054), .CLK(n9549), .Q(
        g1798), .QN(n5833) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(n8975), .CLK(n9588), .Q(
        test_so11), .QN(n8878) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(n9093), .CLK(n9529), 
        .Q(g2941), .QN(n8737) );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(n9093), .CLK(n9529), .Q(
        g3905), .QN(n8665) );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(n9033), .CLK(n9560), .Q(
        g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(n9016), .CLK(n9568), .Q(
        g6255), .QN(n8617) );
  SDFFX1 DFF_159_Q_reg ( .D(n1577), .SI(g6255), .SE(n9086), .CLK(n9533), .Q(
        g4375), .QN(n8837) );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(n8979), .CLK(n9587), .Q(
        g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(n8954), .CLK(n9599), .Q(
        g4722), .QN(n5345) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(n9050), .CLK(n9551), .Q(
        g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(n8925), .CLK(n9613), .Q(
        g13099) );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(n9054), .CLK(n9549), .Q(
        g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(n8911), .CLK(n9621), .Q(
        g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(n9064), .CLK(n9544), .Q(
        g3100), .QN(n8799) );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(n8936), .CLK(n9608), .Q(
        test_so12) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(n8936), .CLK(n9608), 
        .Q(g1437) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(n9100), .CLK(n9526), .Q(
        g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(n8974), .CLK(n9589), .Q(
        g1579), .QN(n8436) );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(n9089), .CLK(n9531), .Q(
        g5567), .QN(n8688) );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(n9089), .CLK(n9531), .Q(
        g1752), .QN(n5797) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(n8929), .CLK(n9611), .Q(
        g1917), .QN(n8757) );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(n9033), .CLK(n9559), .Q(
        g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(n8954), .CLK(n9599), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(n8954), .CLK(n9599), .Q(
        g8132), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(n9017), .CLK(n9567), .Q(
        g6267) );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(n8956), .CLK(n9598), .Q(
        g16659), .QN(n8555) );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(n8936), .CLK(n9608), .Q(
        g1442), .QN(n8717) );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(n8912), .CLK(n9620), .Q(
        test_so13) );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(n9022), .CLK(n9565), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(n9022), .CLK(n9565), .Q(
        g10500) );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(n8983), .CLK(n9584), .Q(
        g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(n8945), .CLK(n9603), .Q(
        g5264), .QN(n8649) );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(n8945), .CLK(n9603), .Q(
        g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(n8932), .CLK(n9610), .Q(
        g2610), .QN(n8759) );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(n8932), .CLK(n9610), .Q(
        g5160), .QN(n5498) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(n8989), .CLK(n9581), .Q(
        g5933) );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(n9027), .CLK(n9562), .Q(
        g1454) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(n8942), .CLK(n9605), .Q(
        g753), .QN(n8828) );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(n8941), .CLK(n9605), .Q(
        g1296) );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(n8941), .CLK(n9605), .Q(
        g3151), .QN(n5495) );
  SDFFX1 DFF_197_Q_reg ( .D(n422), .SI(g3151), .SE(n8941), .CLK(n9605), .Q(
        test_so14) );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(n9021), .CLK(n9566), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(n8957), .CLK(n9598), .Q(
        g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(g33615), .SI(g3530), .SE(n9081), .CLK(n9536), .Q(
        g4104), .QN(n8593) );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(n9020), .CLK(n9566), .Q(
        g1532), .QN(n8588) );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(n9020), .CLK(n9566), .Q(
        g9251) );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(n9020), .CLK(n9566), .Q(
        n9352), .QN(n15965) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(n9079), .CLK(n9536), .Q(
        n9351), .QN(DFF_206_n1) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(n9079), .CLK(n9537), .Q(
        g4754), .QN(n5877) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(n8953), .CLK(n9599), .Q(
        g1189), .QN(n5642) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(n8938), .CLK(n9607), .Q(
        g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(n9070), .CLK(n9541), .Q(
        g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(n9071), .CLK(n9540), .Q(
        g1389) );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(n9007), .CLK(n9572), .Q(
        test_so15), .QN(n8899) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(n9078), .CLK(n9537), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(n8954), .CLK(n9599), .Q(
        g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(n8954), .CLK(n9599), .Q(
        g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(g33588), .SI(g4269), .SE(n9026), .CLK(n9563), .Q(
        g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(n9025), .CLK(n9563), .Q(
        g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(n9089), .CLK(n9531), .Q(
        g5611), .QN(n8659) );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(n8971), .CLK(n9591), .Q(
        g16627), .QN(n8559) );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(n9113), .CLK(n9519), .Q(
        g4572), .QN(n8404) );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(n9096), .CLK(n9528), .Q(
        g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(n9096), .CLK(n9528), .Q(
        g2898), .QN(n8740) );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(n9039), .CLK(n9556), .Q(
        g3343), .QN(n8578) );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(n9039), .CLK(n9556), .Q(
        g3235) );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(n9021), .CLK(n9565), .Q(
        test_so16) );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(n8943), .CLK(n9605), 
        .Q(g3566) );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(n8913), .CLK(n9619), .Q(
        n9348), .QN(n15959) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(n9041), .CLK(n9555), .Q(
        g4961), .QN(n5770) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(n8921), .CLK(n9615), .Q(
        g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(n9015), .CLK(n9569), .Q(
        g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(n9073), .CLK(n9540), .Q(
        g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(n8959), .CLK(n9597), .Q(
        g7257) );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(n8958), .CLK(n9597), .Q(
        g5802), .QN(n8800) );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(n9043), .CLK(n9555), .Q(
        g2852) );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(n8952), .CLK(n9600), .Q(
        g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(n8949), .CLK(n9601), .Q(
        g681), .QN(n8441) );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(n9035), .CLK(n9559), .Q(
        g437) );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(n9035), .CLK(n9559), .Q(
        test_so17), .QN(n8886) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(n8987), .CLK(n9583), 
        .Q(g5901), .QN(n8686) );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(n9095), .CLK(n9528), .Q(
        g2886), .QN(n8739) );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(n9090), .CLK(n9531), .Q(
        g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(n9090), .CLK(n9531), .Q(
        g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(n8972), .CLK(n9590), .Q(
        g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(n8946), .CLK(n9603), .Q(
        g1604) );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(n9118), .CLK(n9517), .Q(
        g5092) );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(n8912), .CLK(n9620), .Q(
        g4831) );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(n9086), .CLK(n9533), .Q(
        g4382), .QN(n5714) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(n9053), .CLK(n9550), .Q(
        g6386), .QN(n8580) );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(n8939), .CLK(n9607), .Q(
        g479) );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(n9114), .CLK(n9519), .Q(
        g3965), .QN(n8500) );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(n9077), .CLK(n9538), .Q(
        test_so18), .QN(n8906) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(n8991), .CLK(n9581), 
        .Q(g2008) );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(n8991), .CLK(n9581), .Q(
        g736), .QN(n8791) );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(n8935), .CLK(n9608), .Q(
        g3933) );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(n9068), .CLK(n9542), .Q(
        g222), .QN(n8747) );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(n9064), .CLK(n9544), .Q(
        g3050), .QN(n5998) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(n8963), .CLK(n9595), .Q(
        g1052), .QN(n8779) );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(n8963), .CLK(n9595), .Q(
        g17580), .QN(n8553) );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(n9074), .CLK(n9539), .Q(
        g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(n9074), .CLK(n9539), .Q(
        g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(n8944), .CLK(n9604), .Q(
        g5889) );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(n8966), .CLK(n9593), .Q(
        g4495) );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(n8965), .CLK(n9594), .Q(
        g8719) );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(n8964), .CLK(n9594), .Q(
        test_so19), .QN(n8881) );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(n8919), .CLK(n9616), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(n9047), .CLK(n9552), .Q(
        g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(n8916), .CLK(n9618), .Q(
        g2433) );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(n9074), .CLK(n9539), .Q(
        g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(g25748), .SI(g3835), .SE(n8922), .CLK(n9615), .Q(
        g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(n8922), .CLK(n9615), .Q(
        g4917), .QN(n5408) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(n9028), .CLK(n9562), .Q(
        g1070) );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(n8982), .CLK(n9585), .Q(
        g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(n8981), .CLK(n9585), .Q(
        g17715) );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(n8981), .CLK(n9585), .Q(
        g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(n8930), .CLK(n9611), .Q(
        g5339) );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(n8907), .CLK(n9623), .Q(
        g4164), .QN(n8727) );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(n9094), .CLK(n9529), .Q(
        test_so20), .QN(n8890) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(n9072), .CLK(n9540), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(n8909), .CLK(n9622), .Q(
        g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(n9099), .CLK(n9527), .Q(
        g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(n9099), .CLK(n9527), .Q(
        g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(n9099), .CLK(n9527), .Q(
        g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(n8914), .CLK(n9619), .Q(
        g3680) );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(n9011), .CLK(n9570), .Q(
        g6637) );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(n8952), .CLK(n9600), .Q(
        g174), .QN(n5402) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(n9066), .CLK(n9543), .Q(
        g1682), .QN(n8419) );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(n9035), .CLK(n9559), .Q(
        g355), .QN(n8716) );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(n9034), .CLK(n9559), .Q(
        g1087), .QN(n8723) );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(n8940), .CLK(n9606), .Q(
        g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(n8996), .CLK(n9578), .Q(
        test_so21), .QN(n8869) );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(n9015), .CLK(n9568), 
        .Q(g6307) );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(n9015), .CLK(n9568), .Q(
        g3802), .QN(n8801) );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(n9015), .CLK(n9569), .Q(
        g6159), .QN(n8421) );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(n9015), .CLK(n9569), .Q(
        g2255), .QN(n5414) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(n9072), .CLK(n9540), .Q(
        g2815), .QN(n5404) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(n8987), .CLK(n9583), .Q(
        g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n8843), .SI(g911), .SE(n9109), .CLK(n9521), .Q(g43), .QN(n8776) );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(n8956), .CLK(n9598), .Q(
        g16775), .QN(n8569) );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(n9089), .CLK(n9532), .Q(
        g1748) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(n9103), .CLK(n9525), .Q(
        g5551) );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(n9084), .CLK(n9534), .Q(
        g3558), .QN(n8614) );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(n9076), .CLK(n9538), .Q(
        g5499), .QN(n5885) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(n9076), .CLK(n9538), .Q(
        test_so22), .QN(n8894) );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(n9093), .CLK(n9529), 
        .Q(g3901) );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(n9082), .CLK(n9535), .Q(
        g4888), .QN(n5863) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(n9017), .CLK(n9568), .Q(
        g6251) );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(n8945), .CLK(n9604), .Q(
        g17649), .QN(n8560) );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(n9065), .CLK(n9544), .Q(
        g1373), .QN(n8455) );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(n9064), .CLK(n9544), .Q(
        g8215) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(n9058), .CLK(n9547), .Q(
        g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(n9049), .CLK(n9552), .Q(
        g2783), .QN(n5403) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(n8977), .CLK(n9588), .Q(
        g4281), .QN(n8750) );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(n8927), .CLK(n9612), .Q(
        g3574) );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(n9036), .CLK(n9558), .Q(
        g2112) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(n9036), .CLK(n9558), .Q(
        g1283), .QN(n5635) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(n9036), .CLK(n9558), .Q(
        test_so23) );
  SDFFX1 DFF_325_Q_reg ( .D(g10122), .SI(test_si24), .SE(n9069), .CLK(n9541), 
        .Q(g4297), .QN(n8372) );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(n9069), .CLK(n9541), .Q(
        g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(n9028), .CLK(n9562), .Q(
        g13272), .QN(n8798) );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(n9033), .CLK(n9560), .Q(
        g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(n408), .SI(g758), .SE(n8983), .CLK(n9585), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(n9104), .CLK(n9524), .Q(
        g6537), .QN(n5884) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(n9104), .CLK(n9524), .Q(
        g5543) );
  SDFFX1 DFF_334_Q_reg ( .D(g7946), .SI(g5543), .SE(n8973), .CLK(n9589), .Q(
        g8475), .QN(n8797) );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(n9018), .CLK(n9567), .Q(
        g5961) );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(n9018), .CLK(n9567), .Q(
        g6243) );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(n8908), .CLK(n9622), .Q(
        n9340), .QN(n15963) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(n9061), .CLK(n9546), .Q(
        g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(n8936), .CLK(n9608), .Q(
        test_so24) );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(n9025), .CLK(n9563), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(n9025), .CLK(n9563), .Q(
        g1664) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(n9025), .CLK(n9564), .Q(
        g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(n9013), .CLK(n9569), .Q(
        g6629) );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(n9061), .CLK(n9545), .Q(
        g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(n9042), .CLK(n9555), .Q(
        g4049), .QN(n8586) );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(n9044), .CLK(n9554), .Q(
        g7260) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(n9044), .CLK(n9554), .Q(
        g2932), .QN(n8814) );
  SDFFX1 DFF_350_Q_reg ( .D(n1733), .SI(g2932), .SE(n9110), .CLK(n9521), .Q(
        g4575) );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(n9110), .CLK(n9521), .Q(
        g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(n8966), .CLK(n9593), .Q(
        g4498) );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(n8947), .CLK(n9603), .Q(
        g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(n9117), .CLK(n9517), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(g25654), .SI(test_si26), .SE(n8919), .CLK(n9616), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(n9061), .CLK(n9545), .Q(
        g29215) );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g29215), .SE(n8920), .CLK(n9616), .Q(
        g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(n9068), .CLK(n9542), .Q(
        g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(n8930), .CLK(n9611), .Q(
        g17639), .QN(n8648) );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(n9078), .CLK(n9537), .Q(
        g5831) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(n9027), .CLK(n9563), .Q(
        g239), .QN(n8590) );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(n9000), .CLK(n9576), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(n9116), .CLK(n9518), .Q(
        g2848), .QN(n8821) );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(n8910), .CLK(n9621), .Q(
        g5022), .QN(n8773) );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(n8910), .CLK(n9621), .Q(
        g16955) );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(n9095), .CLK(n9529), .Q(
        g1030), .QN(n8457) );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(n8970), .CLK(n9591), .Q(
        test_so26) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(n9009), .CLK(n9572), 
        .Q(g3231) );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(n8994), .CLK(n9579), .Q(
        g9817), .QN(n8373) );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(n8994), .CLK(n9579), .Q(
        g1430), .QN(n8721) );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(n8994), .CLK(n9579), .Q(
        n9336), .QN(n15961) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(n8969), .CLK(n9592), .Q(
        g2241), .QN(n8418) );
  SDFFX1 DFF_375_Q_reg ( .D(g24262), .SI(g2241), .SE(n8993), .CLK(n9579), .Q(
        g1564), .QN(n8720) );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(n8958), .CLK(n9597), .Q(
        g9680), .QN(n8379) );
  SDFFX1 DFF_377_Q_reg ( .D(test_so92), .SI(g9680), .SE(n8921), .CLK(n9616), 
        .Q(g6148), .QN(n8806) );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(n9012), .CLK(n9570), .Q(
        g6649), .QN(n8668) );
  SDFFX1 DFF_379_Q_reg ( .D(g34781), .SI(g6649), .SE(n9056), .CLK(n9548), .Q(
        g110) );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(n9027), .CLK(n9563), .Q(
        g14147) );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(n8959), .CLK(n9596), .Q(
        g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(n8959), .CLK(n9596), .Q(
        test_so27) );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(n8966), .CLK(n9593), 
        .Q(g4504) );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(n8965), .CLK(n9593), .Q(
        g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(n8965), .CLK(n9593), .Q(
        g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(n8996), .CLK(n9578), .Q(
        g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(g25720), .SI(g2319), .SE(n8924), .CLK(n9614), .Q(
        g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(n9110), .CLK(n9521), .Q(
        g11770) );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(n9110), .CLK(n9521), .Q(
        g5208) );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(n9090), .CLK(n9531), .Q(
        g5579) );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(n8974), .CLK(n9589), .Q(
        g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(n8974), .CLK(n9589), .Q(
        g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(n8958), .CLK(n9597), .Q(
        g5752), .QN(n5996) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(n8990), .CLK(n9581), .Q(
        g6279) );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(n8990), .CLK(n9581), .Q(
        test_so28) );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(n9067), .CLK(n9543), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(n9099), .CLK(n9526), .Q(
        g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(n8956), .CLK(n9598), .Q(
        g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(n8935), .CLK(n9609), .Q(
        g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(n9027), .CLK(n9562), .Q(
        g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(n9027), .CLK(n9563), .Q(
        g14125) );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(n8995), .CLK(n9578), .Q(
        g2370) );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(n8995), .CLK(n9578), .Q(
        g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(n8973), .CLK(n9589), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(n9058), .CLK(n9547), .Q(
        g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(n8972), .CLK(n9590), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(n8975), .CLK(n9588), .Q(
        g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(n8975), .CLK(n9589), .Q(
        test_so29), .QN(n8862) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(n8941), .CLK(n9606), 
        .Q(g2984), .QN(n5842) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(n9114), .CLK(n9519), .Q(
        g3961) );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(n8953), .CLK(n9599), .Q(
        g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(n9106), .CLK(n9523), .Q(
        g101) );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(n9105), .CLK(n9523), .Q(
        g8918), .QN(n15969) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(n9105), .CLK(n9523), .Q(
        g6625) );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(n9095), .CLK(n9528), .Q(
        n9332), .QN(DFF_420_n1) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(n9095), .CLK(n9528), .Q(
        g1018), .QN(n8456) );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(n8992), .CLK(n9580), .Q(
        g17320), .QN(n8444) );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(n9042), .CLK(n9555), .Q(
        g4045), .QN(n8587) );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(n8935), .CLK(n9608), .Q(
        g1467) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(n9073), .CLK(n9539), .Q(
        g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(n9003), .CLK(n9575), .Q(
        test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(n9079), .CLK(n9537), 
        .Q(g5990), .QN(n5589) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(n8939), .CLK(n9606), .Q(
        g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(n9109), .CLK(n9522), .Q(
        g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(g29306), .SI(g5029), .SE(n9082), .CLK(n9535), .Q(
        g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(n9081), .CLK(n9535), .Q(
        g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(n9047), .CLK(n9552), .Q(
        g1816), .QN(n8355) );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(n9023), .CLK(n9565), .Q(
        g4369), .QN(n8591) );
  SDFFX1 DFF_439_Q_reg ( .D(n470), .SI(g4369), .SE(n9023), .CLK(n9565), .Q(
        g4578) );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(n9023), .CLK(n9564), .Q(
        g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(n9075), .CLK(n9539), .Q(
        g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(n9047), .CLK(n9553), .Q(
        g2514), .QN(n8387) );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(n9097), .CLK(n9527), .Q(
        g3288), .QN(n5400) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(n8911), .CLK(n9621), .Q(
        test_so31) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(n9051), .CLK(n9550), 
        .Q(g2145), .QN(n5307) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(n9065), .CLK(n9543), .Q(
        g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(n8950), .CLK(n9601), .Q(
        g513), .QN(n5548) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(n9004), .CLK(n9574), .Q(
        g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(n8985), .CLK(n9584), .Q(
        g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(n8985), .CLK(n9584), .Q(
        g2763), .QN(n8337) );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(n9100), .CLK(n9526), .Q(
        g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(n8953), .CLK(n9599), .Q(
        g952) );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(n8939), .CLK(n9606), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(n8934), .CLK(n9609), .Q(
        g1950), .QN(n8417) );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(n9107), .CLK(n9523), .Q(
        g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(n8997), .CLK(n9578), .Q(
        g2307) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(n8996), .CLK(n9578), .Q(
        test_so32) );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(n9101), .CLK(n9526), 
        .Q(g8398), .QN(n8376) );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(n9100), .CLK(n9526), .Q(
        g4664), .QN(n8377) );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(n8985), .CLK(n9584), .Q(
        g2223) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(n9079), .CLK(n9537), .Q(
        g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(n9013), .CLK(n9569), .Q(
        g6645) );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(n9037), .CLK(n9557), .Q(
        g2016) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(n8971), .CLK(n9590), .Q(
        g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(n8971), .CLK(n9590), .Q(
        g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(n8997), .CLK(n9578), .Q(
        g2315) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(n9019), .CLK(n9567), .Q(
        g2811) );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(n9019), .CLK(n9567), .Q(
        g5957) );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(n8999), .CLK(n9576), .Q(
        g2047) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(n8999), .CLK(n9576), .Q(
        test_so33), .QN(n8868) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(n8945), .CLK(n9603), 
        .Q(g17760), .QN(n8575) );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(n9103), .CLK(n9525), .Q(
        g5575) );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(n9101), .CLK(n9526), .Q(
        n9327), .QN(DFF_477_n1) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(n9101), .CLK(n9526), .Q(
        g3752), .QN(n5994) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(n8935), .CLK(n9608), .Q(
        g3917) );
  SDFFX1 DFF_480_Q_reg ( .D(test_so86), .SI(g3917), .SE(n9006), .CLK(n9573), 
        .Q(g8783), .QN(n15971) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(n9006), .CLK(n9573), .Q(
        g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(n8958), .CLK(n9597), .Q(
        g4388) );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(n9016), .CLK(n9568), .Q(
        g6275) );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(n8912), .CLK(n9620), .Q(
        g6311), .QN(n8490) );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(n8912), .CLK(n9620), .Q(
        g8916) );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(n9094), .CLK(n9529), .Q(
        g1041), .QN(n8339) );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(n8967), .CLK(n9593), .Q(
        test_so34) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(n9046), .CLK(n9553), 
        .Q(g2537) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(n9087), .CLK(n9533), .Q(
        g29221), .QN(g23612) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g29221), .SE(n9086), .CLK(n9533), .Q(
        g4430), .QN(n8405) );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(n8913), .CLK(n9619), .Q(
        n9325) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(n8912), .CLK(n9620), .Q(
        g4826) );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(n9017), .CLK(n9567), .Q(
        g6239), .QN(n8493) );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(n8959), .CLK(n9597), .Q(
        g232), .QN(n8589) );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(n9029), .CLK(n9561), .Q(
        g5268) );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(n9029), .CLK(n9562), .Q(
        g6545), .QN(n5497) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(n9048), .CLK(n9552), .Q(
        n9324) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(n9048), .CLK(n9552), .Q(
        g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(n9108), .CLK(n9522), .Q(
        g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(n9108), .CLK(n9522), .Q(
        test_so35), .QN(n8375) );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(n8967), .CLK(n9592), 
        .Q(g1890) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(n8967), .CLK(n9593), .Q(
        g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(n9052), .CLK(n9550), .Q(
        g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(n9051), .CLK(n9550), .Q(
        g2130), .QN(n5487) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(n9081), .CLK(n9535), .Q(
        g4108), .QN(n5715) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(n9020), .CLK(n9566), .Q(
        g4308) );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(n8963), .CLK(n9594), .Q(
        g475) );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(n8963), .CLK(n9594), .Q(
        g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(n8963), .CLK(n9594), .Q(
        g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(n9115), .CLK(n9518), .Q(
        n9322), .QN(DFF_514_n1) );
  SDFFX1 DFF_515_Q_reg ( .D(n420), .SI(n9322), .SE(n9115), .CLK(n9518), .Q(
        g12184) );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(n9115), .CLK(n9518), .Q(
        g3990), .QN(n5594) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(n8965), .CLK(n9593), .Q(
        test_so36), .QN(n8872) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(n8983), .CLK(n9585), 
        .Q(g1992) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(n8983), .CLK(n9585), .Q(
        g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(n8982), .CLK(n9585), .Q(
        g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(n8920), .CLK(n9616), .Q(
        g832), .QN(n8796) );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(n8989), .CLK(n9581), .Q(
        g5897) );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(n8989), .CLK(n9582), .Q(
        g25689) );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(n9010), .CLK(n9571), .Q(
        g4571) );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(n8961), .CLK(n9595), .Q(
        g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(n8908), .CLK(n9622), .Q(
        g4455) );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(n9076), .CLK(n9538), .Q(
        g2902), .QN(n8823) );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(n9076), .CLK(n9538), .Q(
        g333), .QN(n8715) );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(n8952), .CLK(n9600), .Q(
        g168), .QN(n5606) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(n9073), .CLK(n9540), .Q(
        test_so37) );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(n9083), .CLK(n9535), 
        .Q(g3684) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(n9083), .CLK(n9535), .Q(
        g3639), .QN(n5591) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(n8931), .CLK(n9611), .Q(
        g14597) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(n9040), .CLK(n9556), .Q(
        g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(n9108), .CLK(n9522), .Q(
        g5406), .QN(n5992) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(n9108), .CLK(n9522), .Q(
        g269), .QN(n8472) );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(n9035), .CLK(n9558), .Q(
        g401) );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(n9035), .CLK(n9558), .Q(
        g6040), .QN(n8581) );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(n9035), .CLK(n9558), .Q(
        g441), .QN(n8467) );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(n8910), .CLK(n9621), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(n9115), .CLK(n9519), .Q(
        g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(n9115), .CLK(n9519), .Q(
        g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(n9023), .CLK(n9565), .Q(
        test_so38), .QN(n8864) );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(n9093), .CLK(n9530), 
        .Q(g3957), .QN(n8663) );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(n9081), .CLK(n9535), .Q(
        g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(n9053), .CLK(n9549), .Q(
        g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(n9053), .CLK(n9549), .Q(
        g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(n9058), .CLK(n9547), .Q(
        g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(n9014), .CLK(n9569), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(n8943), .CLK(n9605), .Q(
        g3498) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(n9051), .CLK(n9551), .Q(
        g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(n9057), .CLK(n9547), .Q(
        g14201) );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(n9057), .CLK(n9548), .Q(
        g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(n8954), .CLK(n9599), .Q(
        g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(n9007), .CLK(n9573), .Q(
        g1608) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(n9007), .CLK(n9573), .Q(
        test_so39) );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(n8931), .CLK(n9610), 
        .Q(g17577), .QN(n8650) );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(n8929), .CLK(n9612), .Q(
        g1779) );
  SDFFX1 DFF_568_Q_reg ( .D(g29255), .SI(g1779), .SE(n8916), .CLK(n9618), .Q(
        g2652), .QN(n8513) );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(n9019), .CLK(n9566), .Q(
        g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(n9026), .CLK(n9563), .Q(
        g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(n8950), .CLK(n9601), .Q(
        g661), .QN(n8474) );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(n9112), .CLK(n9520), .Q(
        g4950), .QN(n5772) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(n8924), .CLK(n9614), .Q(
        g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(n9072), .CLK(n9540), .Q(
        g2834), .QN(g23652) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(n9072), .CLK(n9540), .Q(
        g1361), .QN(n8454) );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(n8990), .CLK(n9581), .Q(
        g6235) );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(n8952), .CLK(n9600), .Q(
        g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(n8908), .CLK(n9622), .Q(
        test_so40) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(n9058), .CLK(n9547), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(n9066), .CLK(n9543), .Q(
        g1696), .QN(n5628) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(n8972), .CLK(n9590), .Q(
        g6555), .QN(n8772) );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(n9057), .CLK(n9547), .Q(
        g14189) );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(n8999), .CLK(n9576), .Q(
        g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(n9011), .CLK(n9570), .Q(
        g6621) );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(n9091), .CLK(n9531), .Q(
        g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(n8970), .CLK(n9591), .Q(
        g3897) );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(n9067), .CLK(n9542), .Q(
        g538) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(n8938), .CLK(n9607), .Q(
        g2606) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(n8938), .CLK(n9607), .Q(
        g1472), .QN(n5290) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(n9087), .CLK(n9532), .Q(
        test_so41) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(n9109), .CLK(n9521), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(n8955), .CLK(n9598), .Q(
        g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(n8955), .CLK(n9598), .Q(
        g13259), .QN(n8804) );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(n9059), .CLK(n9547), .Q(
        g405), .QN(n8786) );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(n8994), .CLK(n9579), .Q(
        g5216), .QN(n8600) );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(n8994), .CLK(n9579), .Q(
        g6494), .QN(n8805) );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(n9100), .CLK(n9526), .Q(
        g4669), .QN(n8830) );
  SDFFX1 DFF_606_Q_reg ( .D(g24243), .SI(g4669), .SE(n9022), .CLK(n9565), .Q(
        g996), .QN(n8808) );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(n9085), .CLK(n9534), .Q(
        g4531), .QN(n15958) );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(n9043), .CLK(n9555), .Q(
        g2860), .QN(n8729) );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(n9077), .CLK(n9538), .Q(
        g4743) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(n9013), .CLK(n9570), .Q(
        g6593) );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(n9013), .CLK(n9570), .Q(
        test_so42), .QN(n8903) );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(n8958), .CLK(n9597), 
        .Q(g4411) );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(n9071), .CLK(n9541), .Q(
        g1413) );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(n9022), .CLK(n9565), 
        .Q(g26960) );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(n8931), .CLK(n9611), .Q(
        g13039), .QN(n8629) );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(n9105), .CLK(n9523), .Q(
        g6641), .QN(n8485) );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(n9105), .CLK(n9524), .Q(
        g6), .QN(n8401) );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(n8951), .CLK(n9600), .Q(
        g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n26), .SI(g1936), .SE(n8951), .CLK(n9601), .Q(g55)
         );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(n8950), .CLK(n9601), .Q(
        g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(n8966), .CLK(n9593), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(n8966), .CLK(n9593), .Q(
        g4480) );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(n8997), .CLK(n9578), .Q(
        n9314), .QN(n15964) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(n8928), .CLK(n9612), .Q(
        test_so43) );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(n9104), .CLK(n9524), 
        .Q(g5571) );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(n9083), .CLK(n9534), .Q(
        g3578) );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(n8924), .CLK(n9614), .Q(
        g9555) );
  SDFFX1 DFF_632_Q_reg ( .D(g29294), .SI(g9555), .SE(n9030), .CLK(n9561), .Q(
        g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(n9030), .CLK(n9561), .Q(
        g3582) );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(n9016), .CLK(n9568), .Q(
        g6271) );
  SDFFX1 DFF_635_Q_reg ( .D(g34028_Tj_Payload), .SI(g6271), .SE(n9110), .CLK(
        n9521), .Q(g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(n9026), .CLK(n9563), .Q(
        g2380), .QN(n8386) );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(n8943), .CLK(n9604), .Q(
        g5196) );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(n9038), .CLK(n9557), .Q(
        g3227) );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(n9037), .CLK(n9557), .Q(
        n9312) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(n8960), .CLK(n9596), .Q(
        g14518) );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(n8960), .CLK(n9596), .Q(
        test_so44), .QN(n8895) );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(n9000), .CLK(n9576), 
        .Q(g6541) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(n9039), .CLK(n9557), .Q(
        g3203), .QN(n8646) );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(n9007), .CLK(n9572), .Q(
        g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(n9069), .CLK(n9542), .Q(
        g4760), .QN(n5775) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(n9069), .CLK(n9542), .Q(
        g262), .QN(n8471) );
  SDFFX1 DFF_649_Q_reg ( .D(g33556), .SI(g262), .SE(n9047), .CLK(n9552), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(n9092), .CLK(n9530), .Q(
        g5467), .QN(n8408) );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(n9092), .CLK(n9530), .Q(
        g460) );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(n8928), .CLK(n9612), .Q(
        g6209), .QN(n8768) );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(n9034), .CLK(n9559), .Q(
        g29211) );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g29211), .SE(n9034), .CLK(n9559), .Q(
        g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(n9034), .CLK(n9559), .Q(
        g655), .QN(n8827) );
  SDFFX1 DFF_657_Q_reg ( .D(g34626), .SI(g655), .SE(n9033), .CLK(n9559), .Q(
        test_so45), .QN(n8884) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(n8947), .CLK(n9603), 
        .Q(g2204), .QN(n5620) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(n9041), .CLK(n9556), .Q(
        g5256), .QN(n8495) );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(n8917), .CLK(n9618), .Q(
        g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(n9031), .CLK(n9560), .Q(
        g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(n8909), .CLK(n9621), .Q(
        g13906) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(n9113), .CLK(n9520), .Q(
        g4423) );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(n9113), .CLK(n9520), .Q(
        g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(n8956), .CLK(n9598), .Q(
        g5685), .QN(n8687) );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(n9059), .CLK(n9546), .Q(
        g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(n9061), .CLK(n9545), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(n9009), .CLK(n9572), .Q(
        g3247), .QN(n8477) );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(n9008), .CLK(n9572), .Q(
        g2040), .QN(n5505) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(n9008), .CLK(n9572), .Q(
        test_so46), .QN(DFF_672_n1) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(n9079), .CLK(n9536), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(n8983), .CLK(n9584), .Q(
        g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(n8955), .CLK(n9598), .Q(
        g7916), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g7916), .SE(n8955), .CLK(n9599), .Q(
        g4732), .QN(n5296) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(n9109), .CLK(n9521), .Q(
        g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(n9078), .CLK(n9537), .Q(
        g5817), .QN(n8358) );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(n8996), .CLK(n9578), .Q(
        g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(n8935), .CLK(n9609), .Q(
        g2648), .QN(n8390) );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(n9021), .CLK(n9566), .Q(
        g6736), .QN(n8709) );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(n9112), .CLK(n9520), .Q(
        g4944), .QN(n5875) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(n8976), .CLK(n9588), .Q(
        g4072), .QN(n8820) );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(n9075), .CLK(n9538), .Q(
        g7540) );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(n9075), .CLK(n9538), .Q(
        test_so47) );
  SDFFX1 DFF_688_Q_reg ( .D(g29264), .SI(test_si48), .SE(n9091), .CLK(n9531), 
        .Q(g3466), .QN(n8374) );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(n9080), .CLK(n9536), .Q(
        g4116) );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(n9108), .CLK(n9522), .Q(
        g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(n9075), .CLK(n9539), .Q(
        g4434), .QN(n8403) );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(n9075), .CLK(n9539), .Q(
        g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(n9105), .CLK(n9524), .Q(
        g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(n8961), .CLK(n9596), .Q(
        g17813) );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(n9096), .CLK(n9528), .Q(
        g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(n9045), .CLK(n9554), .Q(
        g3333) );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(n9045), .CLK(n9554), .Q(
        g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(n8979), .CLK(n9586), .Q(
        g4681), .QN(n8713) );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(n9068), .CLK(n9542), .Q(
        g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(n8937), .CLK(n9607), .Q(
        test_so48), .QN(n8897) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(n8946), .CLK(n9603), 
        .Q(g8789), .QN(n8460) );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(n8930), .CLK(n9611), .Q(
        g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(n9044), .CLK(n9554), .Q(
        g2988), .QN(n8762) );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(n8943), .CLK(n9604), .Q(
        g3538) );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(n9058), .CLK(n9547), .Q(
        g301), .QN(n8822) );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(n9058), .CLK(n9547), .Q(
        n9306), .QN(DFF_709_n1) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(n8981), .CLK(n9585), .Q(
        g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(n9055), .CLK(n9549), .Q(
        g17291), .QN(n8433) );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(n8967), .CLK(n9593), .Q(
        g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(n8913), .CLK(n9620), .Q(
        g5011) );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(n8912), .CLK(n9620), .Q(
        g199), .QN(n8746) );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(n9104), .CLK(n9524), .Q(
        g6523), .QN(n5870) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(n8957), .CLK(n9597), .Q(
        test_so49), .QN(n8859) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(n8917), .CLK(n9617), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(n9060), .CLK(n9546), .Q(
        g854) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(n8937), .CLK(n9607), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(n8922), .CLK(n9615), .Q(
        g4922), .QN(n5346) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(n9118), .CLK(n9517), .Q(
        g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(n8973), .CLK(n9590), .Q(
        g5863), .QN(n8770) );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(n9022), .CLK(n9565), .Q(
        g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(g29253), .SI(g4581), .SE(n8916), .CLK(n9618), .Q(
        g2518), .QN(n8512) );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(n9005), .CLK(n9573), .Q(
        g2567) );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(n9052), .CLK(n9550), .Q(
        g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(n9045), .CLK(n9553), .Q(
        g3263), .QN(n8476) );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(n9013), .CLK(n9569), .Q(
        g6613) );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(n9069), .CLK(n9541), .Q(
        test_so50), .QN(n8887) );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(n8994), .CLK(n9579), 
        .Q(g6444), .QN(n5990) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(n9067), .CLK(n9543), .Q(
        g2965), .QN(n8813) );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(n8973), .CLK(n9590), .Q(
        g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(n9055), .CLK(n9549), .Q(
        n9303) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(n9062), .CLK(n9545), .Q(
        g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(n8944), .CLK(n9604), .Q(
        g17646), .QN(n8655) );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(n8927), .CLK(n9613), .Q(
        g3562) );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(n9070), .CLK(n9541), .Q(
        g10122), .QN(n8371) );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122), .SE(n9002), .CLK(n9575), .Q(
        g1404), .QN(n8450) );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(n9115), .CLK(n9519), .Q(
        g3817) );
  SDFFX1 DFF_743_Q_reg ( .D(n8847), .SI(g3817), .SE(n9082), .CLK(n9535), .Q(
        n9302), .QN(n6010) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(n8966), .CLK(n9593), .Q(
        g4501) );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(n8964), .CLK(n9594), .Q(
        test_so51) );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(n9003), .CLK(n9574), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(n9106), .CLK(n9523), .Q(
        g4704), .QN(n5771) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(n9096), .CLK(n9528), .Q(
        g2878), .QN(n8738) );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(n8943), .CLK(n9604), .Q(
        g5220) );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(n9049), .CLK(n9551), .Q(
        g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(n9049), .CLK(n9551), .Q(
        g12368) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(n9001), .CLK(n9575), .Q(
        g316) );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(n8917), .CLK(n9617), .Q(
        g1277), .QN(n8744) );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(n9104), .CLK(n9524), .Q(
        g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(n8916), .CLK(n9618), .Q(
        g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(n9096), .CLK(n9528), .Q(
        g2882), .QN(n8824) );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(n9060), .CLK(n9546), .Q(
        test_so52), .QN(n8748) );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(n8967), .CLK(n9592), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(n8967), .CLK(n9592), .Q(
        g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(g34975), .SI(g305), .SE(n9114), .CLK(n9519), .Q(g8), .QN(n8810) );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(n9019), .CLK(n9566), .Q(
        g2799) );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(n9019), .CLK(n9567), .Q(
        g14167) );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(n8931), .CLK(n9611), .Q(
        g17787) );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(n8921), .CLK(n9615), .Q(
        g4912), .QN(n5297) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(n9079), .CLK(n9536), .Q(
        g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(n9046), .CLK(n9553), .Q(
        g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(n8942), .CLK(n9605), .Q(
        g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(n9087), .CLK(n9533), .Q(
        g550), .QN(n8745) );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(n8959), .CLK(n9597), .Q(
        g255), .QN(n8470) );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(n8929), .CLK(n9611), .Q(
        test_so53), .QN(n8905) );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(n9041), .CLK(n9556), 
        .Q(g5240) );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(n8936), .CLK(n9608), .Q(
        g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(n8936), .CLK(n9608), .Q(
        g3863), .QN(n8771) );
  SDFFX1 DFF_777_Q_reg ( .D(g29245), .SI(g3863), .SE(n8929), .CLK(n9611), .Q(
        g1959), .QN(n8511) );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(n9091), .CLK(n9531), .Q(
        g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(n9011), .CLK(n9570), .Q(
        g6653) );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(n8925), .CLK(n9614), .Q(
        g17764), .QN(n8667) );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(n9114), .CLK(n9519), .Q(
        g2864), .QN(n5489) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(n9082), .CLK(n9535), .Q(
        g4894), .QN(n5774) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(n8961), .CLK(n9596), .Q(
        g17678), .QN(n8658) );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(n8960), .CLK(n9596), .Q(
        g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(n8960), .CLK(n9596), .Q(
        g16693), .QN(n8664) );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(n8950), .CLK(n9601), .Q(
        test_so54) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(n9094), .CLK(n9529), 
        .Q(g1002), .QN(n8449) );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(n9032), .CLK(n9560), .Q(
        g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(n9032), .CLK(n9560), .Q(
        g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(n9022), .CLK(n9565), .Q(
        g1236), .QN(n8435) );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(n8980), .CLK(n9586), .Q(
        g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(n8980), .CLK(n9586), .Q(
        g2476), .QN(n8758) );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(n9025), .CLK(n9564), .Q(
        g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(n9026), .CLK(n9563), .Q(
        g2375), .QN(n8416) );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(n8980), .CLK(n9586), .Q(
        g63) );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(n8980), .CLK(n9586), .Q(
        g17739), .QN(n8566) );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(n8965), .CLK(n9594), .Q(
        g358), .QN(n8473) );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(n8964), .CLK(n9594), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(g28043), .SI(g896), .SE(n8964), .CLK(n9594), .Q(
        test_so55), .QN(n8874) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(n8926), .CLK(n9613), 
        .Q(g3161), .QN(n8752) );
  SDFFX1 DFF_804_Q_reg ( .D(g29251), .SI(g3161), .SE(n8917), .CLK(n9617), .Q(
        g2384), .QN(n8507) );
  SDFFX1 DFF_806_Q_reg ( .D(test_so80), .SI(g2384), .SE(n8998), .CLK(n9577), 
        .Q(g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(n8998), .CLK(n9577), .Q(
        g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(n8915), .CLK(n9619), .Q(
        g4561) );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(n8915), .CLK(n9619), .Q(
        g2024) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(n8914), .CLK(n9619), .Q(
        g3451), .QN(n8807) );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(n9037), .CLK(n9558), .Q(
        g2795) );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(n9050), .CLK(n9551), .Q(
        g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(n8917), .CLK(n9618), .Q(
        g4527), .QN(n8725) );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(n9062), .CLK(n9545), .Q(
        g1844) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(n8988), .CLK(n9582), .Q(
        g5937) );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(n8988), .CLK(n9582), .Q(
        test_so56) );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(n9046), .CLK(n9553), 
        .Q(g2523), .QN(n5281) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(n8962), .CLK(n9595), .Q(
        g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(n8937), .CLK(n9608), .Q(
        g2643), .QN(n8415) );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(n8937), .CLK(n9608), .Q(
        g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(n9068), .CLK(n9542), .Q(
        g8358), .QN(n8452) );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(n9056), .CLK(n9548), .Q(
        n9295) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(n9056), .CLK(n9548), .Q(
        g5156) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(n9056), .CLK(n9548), .Q(
        g30332), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(g34975), .SI(g30332), .SE(n9055), .CLK(n9548), .Q(
        n9294), .QN(DFF_829_n1) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(n8956), .CLK(n9598), .Q(
        g8279) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(n8977), .CLK(n9587), .Q(
        g8839) );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(n8934), .CLK(n9609), .Q(
        g1955), .QN(n8383) );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(n8934), .CLK(n9609), .Q(
        test_so57), .QN(n8866) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(n9014), .CLK(n9569), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(n8925), .CLK(n9614), .Q(
        g14749) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(n9053), .CLK(n9550), .Q(
        g4771), .QN(n5769) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(n9052), .CLK(n9550), .Q(
        g6098), .QN(n5988) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(n8919), .CLK(n9617), .Q(
        g3147) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(n9040), .CLK(n9556), .Q(
        g3347), .QN(n8577) );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(n9014), .CLK(n9569), .Q(
        g2269) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(n9014), .CLK(n9569), .Q(
        g191), .QN(n8453) );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(n9004), .CLK(n9574), .Q(
        g2712), .QN(n8368) );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(n9049), .CLK(n9552), .Q(
        g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(n8985), .CLK(n9583), .Q(
        g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(n8920), .CLK(n9616), .Q(
        test_so58), .QN(n8863) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(n8986), .CLK(n9583), 
        .Q(g17819) );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(n8985), .CLK(n9583), .Q(
        g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(n9094), .CLK(n9529), .Q(
        g2927), .QN(n8815) );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(n9085), .CLK(n9533), .Q(
        g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(n9018), .CLK(n9567), .Q(
        g5929) );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(n8922), .CLK(n9615), .Q(
        g4907), .QN(n5295) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(n8922), .CLK(n9615), .Q(
        g16874) );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(n9113), .CLK(n9519), .Q(
        g4035) );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(n8976), .CLK(n9588), .Q(
        g2946), .QN(n8818) );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(n8976), .CLK(n9588), .Q(
        g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(n8976), .CLK(n9588), .Q(
        g4082), .QN(n8446) );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(n8971), .CLK(n9590), .Q(
        g9743) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(n9037), .CLK(n9557), .Q(
        test_so59) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(n9051), .CLK(n9551), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(n8915), .CLK(n9618), .Q(
        g1620) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(n9088), .CLK(n9532), .Q(
        g2831), .QN(g30331) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(n9088), .CLK(n9532), .Q(
        g667) );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(n9061), .CLK(n9546), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(n8969), .CLK(n9591), .Q(
        g3937) );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(n8982), .CLK(n9585), .Q(
        g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(n8982), .CLK(n9585), .Q(
        g1249) );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(n8981), .CLK(n9586), .Q(
        g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(n8970), .CLK(n9591), .Q(
        g16924) );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(n9050), .CLK(n9551), .Q(
        g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(n9116), .CLK(n9518), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(n9033), .CLK(n9559), .Q(
        test_so60), .QN(n8904) );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(n8989), .CLK(n9581), 
        .Q(g5949) );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(n9082), .CLK(n9535), .Q(
        g6682), .QN(n5590) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(n9061), .CLK(n9546), .Q(
        g904) );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(n9043), .CLK(n9554), .Q(
        g2873), .QN(n5488) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(n9062), .CLK(n9545), .Q(
        g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(n9118), .CLK(n9517), .Q(
        g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(n9103), .CLK(n9524), .Q(
        g5603), .QN(n8481) );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(n9103), .CLK(n9524), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(n9002), .CLK(n9575), .Q(
        g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(n8916), .CLK(n9618), .Q(
        g2437) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(n9036), .CLK(n9558), .Q(
        g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(n8984), .CLK(n9584), .Q(
        g2208), .QN(n8756) );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(n9005), .CLK(n9574), .Q(
        test_so61) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(n8976), .CLK(n9588), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(n8920), .CLK(n9616), .Q(
        g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(n9004), .CLK(n9574), .Q(
        g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(n8975), .CLK(n9589), .Q(
        g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(n9098), .CLK(n9527), .Q(
        g5583) );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(n9032), .CLK(n9560), .Q(
        g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(n9010), .CLK(n9571), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(n9010), .CLK(n9571), .Q(
        g17743), .QN(n8676) );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(n9094), .CLK(n9529), .Q(
        g2917), .QN(n8825) );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(n8949), .CLK(n9602), .Q(
        g686) );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(n8940), .CLK(n9606), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(n9088), .CLK(n9532), .Q(
        g671), .QN(n8364) );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(n8942), .CLK(n9605), .Q(
        test_so62), .QN(n8898) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(n9017), .CLK(n9567), 
        .Q(g6283) );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(n8932), .CLK(n9610), .Q(
        g14705) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(n8931), .CLK(n9610), .Q(
        g17519), .QN(n8549) );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(n8931), .CLK(n9610), .Q(
        g8784), .QN(n15972) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(n8926), .CLK(n9613), .Q(
        g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(n8926), .CLK(n9613), .Q(
        g4489) );
  SDFFX1 DFF_912_Q_reg ( .D(g33564), .SI(g4489), .SE(n8926), .CLK(n9613), .Q(
        g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(n8926), .CLK(n9613), .Q(
        g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(n8923), .CLK(n9615), .Q(
        g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(n8922), .CLK(n9615), .Q(
        g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(n9092), .CLK(n9530), .Q(
        g3929) );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(n9092), .CLK(n9530), .Q(
        g5503) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(n9111), .CLK(n9521), .Q(
        test_so63), .QN(n8741) );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(n8986), .CLK(n9583), 
        .Q(g5925) );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(n8940), .CLK(n9606), .Q(
        g1124) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(n9041), .CLK(n9555), .Q(
        g4955), .QN(n5614) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(n9041), .CLK(n9555), .Q(
        g5224) );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(n8990), .CLK(n9581), .Q(
        g2012) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(n8990), .CLK(n9581), .Q(
        g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(n9055), .CLK(n9548), .Q(
        g5120), .QN(n8407) );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(n9034), .CLK(n9559), .Q(
        g17674), .QN(n8564) );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(n9026), .CLK(n9563), .Q(
        g2389), .QN(n5631) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(n9026), .CLK(n9563), .Q(
        g4438), .QN(n8719) );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(n8916), .CLK(n9618), .Q(
        g2429) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(n9037), .CLK(n9558), .Q(
        g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(n8909), .CLK(n9622), .Q(
        test_so64) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(n9102), .CLK(n9525), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(n9085), .CLK(n9534), .Q(
        g18881), .QN(n5541) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g18881), .SE(n8979), .CLK(n9586), .Q(
        g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(n9028), .CLK(n9562), .Q(
        g1199), .QN(n8763) );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(n9028), .CLK(n9562), .Q(
        g19357), .QN(n5401) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(n9103), .CLK(n9525), .Q(
        g5547) );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(n9051), .CLK(n9550), .Q(
        g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(n8971), .CLK(n9591), .Q(
        g16744), .QN(n8573) );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(n8939), .CLK(n9607), .Q(
        g2338) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(n8939), .CLK(n9607), .Q(
        g8919), .QN(n15970) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(n9017), .CLK(n9568), .Q(
        g6247), .QN(n8706) );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(n8929), .CLK(n9612), .Q(
        g2791) );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(n8929), .CLK(n9612), .Q(
        test_so65), .QN(n8896) );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(n9119), .CLK(n9517), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(n9018), .CLK(n9567), .Q(
        g5945) );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(n8978), .CLK(n9587), .Q(
        g5244) );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(n8978), .CLK(n9587), .Q(
        g2759), .QN(n8336) );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(n9082), .CLK(n9535), .Q(
        g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(n9031), .CLK(n9560), .Q(
        g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(n8939), .CLK(n9606), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(n9090), .CLK(n9531), .Q(
        g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(n9067), .CLK(n9542), .Q(
        g209), .QN(n5595) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(n8944), .CLK(n9604), .Q(
        g6609) );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(n9090), .CLK(n9531), .Q(
        g5517), .QN(n8769) );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(n9074), .CLK(n9539), .Q(
        g2449) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(n8937), .CLK(n9608), .Q(
        test_so66) );
  SDFFX1 DFF_961_Q_reg ( .D(g18881), .SI(test_si67), .SE(n9085), .CLK(n9534), 
        .Q(n9281) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(n9004), .CLK(n9574), .Q(
        g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(n8987), .CLK(n9582), .Q(
        g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(n9024), .CLK(n9564), .Q(
        g2098), .QN(n5280) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(n9024), .CLK(n9564), .Q(
        g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(n9050), .CLK(n9551), .Q(
        g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(n8944), .CLK(n9604), .Q(
        g6589) );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(n8932), .CLK(n9610), .Q(
        n9280) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(n8932), .CLK(n9610), .Q(
        g17845) );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(n8925), .CLK(n9614), .Q(
        g17871) );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(n9036), .CLK(n9558), .Q(
        g429) );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(n8933), .CLK(n9610), .Q(
        g1870) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(n8933), .CLK(n9610), .Q(
        test_so67), .QN(n8902) );
  SDFFX1 DFF_977_Q_reg ( .D(g29243), .SI(test_si68), .SE(n9063), .CLK(n9545), 
        .Q(g1825), .QN(n8505) );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(n9045), .CLK(n9554), .Q(
        g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(n9044), .CLK(n9554), .Q(
        g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(test_so46), .SI(g4392), .SE(n9008), .CLK(n9572), 
        .Q(g8283) );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(n9030), .CLK(n9561), .Q(
        g3546) );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(n9029), .CLK(n9561), .Q(
        g5236) );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(n9089), .CLK(n9532), .Q(
        g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(n8923), .CLK(n9615), .Q(
        g4854), .QN(n8363) );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(n9093), .CLK(n9530), .Q(
        g3925) );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(n9105), .CLK(n9524), .Q(
        g6509), .QN(n8395) );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(n8942), .CLK(n9605), .Q(
        g732), .QN(n5732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(n9002), .CLK(n9575), .Q(
        g2504), .QN(n8761) );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(n9002), .CLK(n9575), .Q(
        test_so68), .QN(n8875) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(n9111), .CLK(n9520), 
        .Q(g4520) );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(n9111), .CLK(n9520), .Q(
        g8917), .QN(n15968) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(n8984), .CLK(n9584), .Q(
        g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(n9042), .CLK(n9555), .Q(
        g37), .QN(g30327) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(n9042), .CLK(n9555), .Q(
        g4031) );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(n8948), .CLK(n9602), .Q(
        g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(n8948), .CLK(n9602), .Q(
        g8235) );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(n9080), .CLK(n9536), .Q(
        g4176), .QN(n5494) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(n8960), .CLK(n9596), .Q(
        g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(n8960), .CLK(n9596), .Q(
        g4405), .QN(n8838) );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(n8959), .CLK(n9596), .Q(
        g872) );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(n9099), .CLK(n9526), .Q(
        g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(n9053), .CLK(n9549), .Q(
        test_so69), .QN(n8889) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(n8908), .CLK(n9622), 
        .Q(g4765), .QN(n5613) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(n9098), .CLK(n9527), .Q(
        g5563), .QN(n8605) );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(n8973), .CLK(n9590), .Q(
        g1395), .QN(n8778) );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(n8968), .CLK(n9592), .Q(
        g1913) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(n8938), .CLK(n9607), .Q(
        g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(n8990), .CLK(n9581), .Q(
        g6263) );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(n9114), .CLK(n9519), .Q(
        n9276), .QN(DFF_1012_n1) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(n9114), .CLK(n9519), .Q(
        g3945) );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(n9075), .CLK(n9538), .Q(
        g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(n9023), .CLK(n9564), .Q(
        g4473), .QN(n8423) );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(n8982), .CLK(n9585), .Q(
        g1266), .QN(n8781) );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(n9076), .CLK(n9538), .Q(
        g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(n9087), .CLK(n9532), .Q(
        test_so70), .QN(n8879) );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(n9003), .CLK(n9575), 
        .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(n9116), .CLK(n9518), .Q(
        g5471), .QN(n8365) );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(n9021), .CLK(n9565), .Q(
        g4540) );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(n9021), .CLK(n9566), .Q(
        g6723) );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(n9012), .CLK(n9570), .Q(
        g6605) );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(n9073), .CLK(n9539), .Q(
        n9274) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(n9019), .CLK(n9566), .Q(
        g2173) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(n8977), .CLK(n9588), .Q(
        g9019) );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(n9056), .CLK(n9548), .Q(
        g2491) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(n8923), .CLK(n9614), .Q(
        g4849), .QN(n8834) );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(n8992), .CLK(n9580), .Q(
        g2169) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(n9014), .CLK(n9569), .Q(
        n9273), .QN(n15967) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(n9014), .CLK(n9569), .Q(
        test_so71) );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(n9048), .CLK(n9552), 
        .Q(g29219) );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g29219), .SE(n9048), .CLK(n9552), 
        .Q(g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(n9043), .CLK(n9554), .Q(
        g2868), .QN(n8728) );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(n9054), .CLK(n9549), .Q(
        g2767) );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(n9054), .CLK(n9549), .Q(
        g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(n8961), .CLK(n9595), .Q(
        g16718), .QN(n8562) );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(n9071), .CLK(n9541), 
        .Q(g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(n8977), .CLK(n9587), .Q(
        g5212), .QN(n8651) );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(n8977), .CLK(n9587), .Q(
        g4245), .QN(n5640) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(n8949), .CLK(n9601), .Q(
        g645) );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(n8949), .CLK(n9601), .Q(
        g4291), .QN(n8749) );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(n8940), .CLK(n9606), .Q(
        g29212) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g29212), .SE(n9059), .CLK(n9547), 
        .Q(test_so72), .QN(n8871) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(n8951), .CLK(n9600), 
        .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(n8946), .CLK(n9603), .Q(
        g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(n8946), .CLK(n9603), .Q(
        g8788) );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(n8969), .CLK(n9592), .Q(
        g2246), .QN(n8389) );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(n9063), .CLK(n9545), .Q(
        g1830), .QN(n5413) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(n8927), .CLK(n9612), .Q(
        g3590) );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(n9059), .CLK(n9546), .Q(
        g392), .QN(n8787) );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(n9007), .CLK(n9572), .Q(
        g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(n9000), .CLK(n9576), .Q(
        g6505), .QN(n8422) );
  SDFFX1 DFF_1057_Q_reg ( .D(g24246), .SI(g6505), .SE(n9000), .CLK(n9576), .Q(
        g1221), .QN(n8722) );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(n8988), .CLK(n9582), .Q(
        g5921) );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(n9057), .CLK(n9547), .Q(
        g29216) );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g29216), .SE(n8907), .CLK(n9622), 
        .Q(test_so73), .QN(n8883) );
  SDFFX1 DFF_1061_Q_reg ( .D(test_so42), .SI(test_si74), .SE(n9012), .CLK(
        n9570), .Q(g218), .QN(n8718) );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(n8984), .CLK(n9584), .Q(
        g1932) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(n8918), .CLK(n9617), .Q(
        g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(n9109), .CLK(n9522), .Q(
        g5062), .QN(n8775) );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(n9117), .CLK(n9518), .Q(
        g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(n9116), .CLK(n9518), .Q(
        g2689), .QN(n5347) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(n8972), .CLK(n9590), .Q(
        g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(n9025), .CLK(n9564), .Q(
        g1677) );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(n9024), .CLK(n9564), .Q(
        g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(n9102), .CLK(n9525), .Q(
        g2671) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(n8974), .CLK(n9589), .Q(
        g10527) );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(n8958), .CLK(n9597), 
        .Q(g7243), .QN(n8839) );
  SDFFX1 DFF_1074_Q_reg ( .D(n26), .SI(g7243), .SE(n8951), .CLK(n9601), .Q(
        test_so74) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(n9062), .CLK(n9545), 
        .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(n9118), .CLK(n9517), .Q(
        g29213), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g29213), .SE(n9117), .CLK(n9517), 
        .Q(g5485), .QN(n5869) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(n9003), .CLK(n9574), .Q(
        g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(n9003), .CLK(n9575), .Q(
        g11678), .QN(n5482) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(n9005), .CLK(n9574), 
        .Q(g2638), .QN(n8789) );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(n9080), .CLK(n9536), .Q(
        g4122) );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(n8980), .CLK(n9586), .Q(
        g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(n8986), .CLK(n9583), .Q(
        g5941) );
  SDFFX1 DFF_1086_Q_reg ( .D(g33572), .SI(g5941), .SE(n8986), .CLK(n9583), .Q(
        g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(n8986), .CLK(n9583), .Q(
        g13068), .QN(n8685) );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(n8986), .CLK(n9583), .Q(
        g25) );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(n9008), .CLK(n9572), .Q(
        test_so75) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(n9050), .CLK(n9551), 
        .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(n8984), .CLK(n9584), .Q(
        g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(n9027), .CLK(n9562), .Q(
        n9267), .QN(DFF_1092_n1) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(n9037), .CLK(n9558), .Q(
        g2066), .QN(n5832) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(n8951), .CLK(n9600), .Q(
        g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(n9029), .CLK(n9561), .Q(
        g5252) );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(n8968), .CLK(n9592), .Q(
        g2165) );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(n9005), .CLK(n9573), .Q(
        g2571) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(n8995), .CLK(n9579), .Q(
        g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(n8995), .CLK(n9579), .Q(
        g8403) );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(n8985), .CLK(n9583), .Q(
        g14673) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(n9000), .CLK(n9576), 
        .Q(test_so76), .QN(n8880) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(n9073), .CLK(n9540), 
        .Q(g2827) );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(n9057), .CLK(n9548), .Q(
        g14217) );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(n8923), .CLK(n9615), 
        .Q(g4859), .QN(n8832) );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(n9060), .CLK(n9546), .Q(
        g424), .QN(n8784) );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(n8993), .CLK(n9580), .Q(
        g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(n8992), .CLK(n9580), .Q(
        g17423), .QN(n8442) );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(n8992), .CLK(n9580), 
        .Q(n9265) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(n9072), .CLK(n9540), .Q(
        g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(n9047), .CLK(n9553), .Q(
        g1821), .QN(n8384) );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(n9047), .CLK(n9553), .Q(
        g2509), .QN(n8414) );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(n9118), .CLK(n9517), .Q(
        g5073), .QN(n8412) );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(n8982), .CLK(n9585), .Q(
        test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(n8948), .CLK(n9602), 
        .Q(g8353) );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(n8948), .CLK(n9602), .Q(
        g13085), .QN(n8705) );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(n9012), .CLK(n9570), 
        .Q(g6633) );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(n9055), .CLK(n9548), .Q(
        g5124), .QN(n8356) );
  SDFFX1 DFF_1122_Q_reg ( .D(test_so44), .SI(g5124), .SE(n9055), .CLK(n9549), 
        .Q(g17400), .QN(n8438) );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(n9016), .CLK(n9568), 
        .Q(g6303), .QN(n8677) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(n9119), .CLK(n9517), .Q(
        g5069), .QN(n8411) );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(n9044), .CLK(n9554), .Q(
        g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(n8949), .CLK(n9602), .Q(
        g650) );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(n9008), .CLK(n9572), .Q(
        g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(n8969), .CLK(n9591), .Q(
        g3921) );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(n9024), .CLK(n9564), .Q(
        test_so78), .QN(n8885) );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(n9020), .CLK(n9566), 
        .Q(g6732), .QN(n8710) );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(n9020), .CLK(n9566), .Q(
        g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(n8953), .CLK(n9600), .Q(
        g1061), .QN(n8451) );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(n8943), .CLK(n9605), .Q(
        g3462), .QN(n8410) );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(n8992), .CLK(n9580), .Q(
        g2181) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(n8991), .CLK(n9580), .Q(
        g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(n9063), .CLK(n9544), .Q(
        g1756) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(n8942), .CLK(n9605), .Q(
        g5849) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(n9081), .CLK(n9536), .Q(
        g4112), .QN(n8708) );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(n9101), .CLK(n9525), .Q(
        n9262), .QN(n15960) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(n8947), .CLK(n9603), .Q(
        g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(n9002), .CLK(n9575), .Q(
        test_so79), .QN(n8860) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(n9094), .CLK(n9529), 
        .Q(g1046), .QN(n8835) );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(n8968), .CLK(n9592), .Q(
        g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(n8957), .CLK(n9597), .Q(
        g4401), .QN(n8402) );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(n8957), .CLK(n9597), .Q(
        g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(n9001), .CLK(n9576), .Q(
        g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(n9001), .CLK(n9576), .Q(
        g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(n8911), .CLK(n9620), .Q(
        g2950), .QN(n8735) );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(n9071), .CLK(n9541), .Q(
        g1345), .QN(n8448) );
  SDFFX1 DFF_1154_Q_reg ( .D(g25762), .SI(g1345), .SE(n9000), .CLK(n9576), .Q(
        g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(n8962), .CLK(n9595), .Q(
        g14421) );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(n8962), .CLK(n9595), 
        .Q(g4727), .QN(n5312) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(n8998), .CLK(n9577), .Q(
        test_so80), .QN(n8882) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(n9070), .CLK(n9541), 
        .Q(g1536), .QN(n8812) );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(n9093), .CLK(n9530), .Q(
        g3941) );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(n8964), .CLK(n9594), .Q(
        g370), .QN(n8816) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(n9077), .CLK(n9537), .Q(
        g5694), .QN(n8585) );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(n9062), .CLK(n9545), .Q(
        g1858), .QN(n5892) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(n9062), .CLK(n9545), .Q(
        g446) );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(n8915), .CLK(n9619), .Q(
        g3219) );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(n9063), .CLK(n9544), .Q(
        g1811) );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(n9012), .CLK(n9570), .Q(
        g6601), .QN(n8611) );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(n9073), .CLK(n9539), .Q(
        g2441) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(n8934), .CLK(n9609), .Q(
        g1874) );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(n8934), .CLK(n9609), .Q(
        test_so81), .QN(n8867) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(n8944), .CLK(n9604), 
        .Q(g6581) );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(n9013), .CLK(n9570), .Q(
        g6597), .QN(n8670) );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(n8995), .CLK(n9579), .Q(
        g5008), .QN(n5637) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(n9083), .CLK(n9534), .Q(
        g3610) );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(n9043), .CLK(n9554), .Q(
        g2890), .QN(n8742) );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(n8926), .CLK(n9613), .Q(
        g1978) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(n9054), .CLK(n9549), .Q(
        g1612) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(n9008), .CLK(n9572), .Q(
        g112), .QN(n8468) );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(n9101), .CLK(n9525), .Q(
        g2856), .QN(n8826) );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(n8925), .CLK(n9613), .Q(
        g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(n8925), .CLK(n9613), .Q(
        g17722), .QN(n8669) );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(n8978), .CLK(n9587), 
        .Q(test_so82) );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(n9080), .CLK(n9536), 
        .Q(g4119) );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(n9053), .CLK(n9550), .Q(
        g6390), .QN(n8579) );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(n9070), .CLK(n9541), .Q(
        g1542), .QN(n8764) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(n9070), .CLK(n9541), .Q(
        g4258) );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(n8948), .CLK(n9602), .Q(
        g4818), .QN(n5636) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(n9109), .CLK(n9522), .Q(
        g5033), .QN(n8795) );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(n8955), .CLK(n9599), .Q(
        g4717), .QN(n5344) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(n8993), .CLK(n9580), .Q(
        g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(n8999), .CLK(n9577), .Q(
        g3849) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(n8998), .CLK(n9577), .Q(
        g17778), .QN(n8571) );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(n9039), .CLK(n9557), 
        .Q(g3199) );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(n8907), .CLK(n9623), .Q(
        test_so83) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(n8920), .CLK(n9616), 
        .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(n9031), .CLK(n9560), .Q(
        g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(n9018), .CLK(n9567), .Q(
        g5913), .QN(n8684) );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(n8930), .CLK(n9611), .Q(
        g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(n9100), .CLK(n9526), .Q(
        g6163) );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(n8989), .CLK(n9582), .Q(
        g4125), .QN(n8707) );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(n9098), .CLK(n9527), .Q(
        g4821) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(n9097), .CLK(n9527), .Q(
        g4939), .QN(n5776) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(n8963), .CLK(n9595), .Q(
        g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(n9038), .CLK(n9557), 
        .Q(g3207), .QN(n8598) );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(n9038), .CLK(n9557), .Q(
        g4483) );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(n9045), .CLK(n9553), .Q(
        test_so84) );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(n9107), .CLK(n9523), 
        .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(n8946), .CLK(n9603), .Q(
        g5248) );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(n8907), .CLK(n9622), .Q(
        g2126) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(n9112), .CLK(n9520), .Q(
        g3694), .QN(n8583) );
  SDFFX1 DFF_1215_Q_reg ( .D(g29288), .SI(g3694), .SE(n9116), .CLK(n9518), .Q(
        g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(n9116), .CLK(n9518), .Q(
        g1964), .QN(n5315) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(n9118), .CLK(n9517), .Q(
        g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(n9009), .CLK(n9572), .Q(
        g3215) );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(n8909), .CLK(n9621), .Q(
        g16748), .QN(n8662) );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(n8909), .CLK(n9621), 
        .Q(n9255) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(n9086), .CLK(n9533), .Q(
        g4427), .QN(n8462) );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(n9086), .CLK(n9533), .Q(
        test_so85), .QN(n8893) );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(n9089), .CLK(n9532), 
        .Q(g2779) );
  SDFFX1 DFF_1224_Q_reg ( .D(test_so39), .SI(g2779), .SE(n9006), .CLK(n9573), 
        .Q(g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(n9006), .CLK(n9573), .Q(
        g7245), .QN(DFF_1225_n1) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(n9065), .CLK(n9544), .Q(
        g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(n9065), .CLK(n9544), .Q(
        g1367), .QN(n8439) );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(n8910), .CLK(n9621), .Q(
        g5112) );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(n8910), .CLK(n9621), .Q(
        g19), .QN(n8809) );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(n9081), .CLK(n9536), .Q(
        g4145), .QN(n8726) );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(n8968), .CLK(n9592), .Q(
        g2161) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(n8968), .CLK(n9592), .Q(
        g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(n8938), .CLK(n9607), .Q(
        g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(n9006), .CLK(n9573), .Q(
        test_so86) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(n9051), .CLK(n9551), 
        .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(n9024), .CLK(n9564), .Q(
        g2051), .QN(n8760) );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(n9028), .CLK(n9562), .Q(
        g1193), .QN(n8811) );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(n8996), .CLK(n9578), .Q(
        g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(n8987), .CLK(n9582), .Q(
        g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(n8987), .CLK(n9583), .Q(
        g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(n9063), .CLK(n9545), .Q(
        g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(n9083), .CLK(n9534), .Q(
        g3594) );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(n9044), .CLK(n9554), .Q(
        g2999) );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(n8997), .CLK(n9577), .Q(
        g2303) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(n8997), .CLK(n9577), .Q(
        g17688), .QN(n8557) );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(n8949), .CLK(n9602), 
        .Q(test_so87) );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(n8920), .CLK(n9616), 
        .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(n8919), .CLK(n9616), .Q(
        g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(n9067), .CLK(n9542), .Q(
        g546), .QN(n5492) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(n9067), .CLK(n9543), .Q(
        g2472), .QN(n5619) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(n8988), .CLK(n9582), .Q(
        g5953) );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(n9064), .CLK(n9544), .Q(
        g8277), .QN(n8381) );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(n9064), .CLK(n9544), .Q(
        g1740) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(n8928), .CLK(n9612), .Q(
        g3550) );
  SDFFX1 DFF_1260_Q_reg ( .D(g25683), .SI(g3550), .SE(n9074), .CLK(n9539), .Q(
        g3845), .QN(n5886) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(n9074), .CLK(n9539), .Q(
        g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(n8961), .CLK(n9596), .Q(
        g14635) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(n8915), .CLK(n9618), 
        .Q(test_so88) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(n9092), .CLK(n9530), 
        .Q(g3913) );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(n9113), .CLK(n9520), .Q(
        g10306) );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(n9066), .CLK(n9543), 
        .Q(g1687), .QN(n8388) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(n9101), .CLK(n9525), .Q(
        g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(g33596), .SI(g2681), .SE(n9002), .CLK(n9575), .Q(
        g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(n9001), .CLK(n9575), .Q(
        g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(n9001), .CLK(n9575), .Q(
        g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(g31895), .SI(g2697), .SE(n9086), .CLK(n9533), .Q(
        g4417), .QN(n8333) );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(n8972), .CLK(n9590), .Q(
        g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(n8932), .CLK(n9610), .Q(
        g1141), .QN(n5691) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(n8993), .CLK(n9580), .Q(
        g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(n9048), .CLK(n9552), 
        .Q(test_so89), .QN(n8892) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(n9065), .CLK(n9543), 
        .Q(g1710) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(n9104), .CLK(n9524), .Q(
        g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(n9038), .CLK(n9557), .Q(
        g3255), .QN(n8644) );
  SDFFX1 DFF_1281_Q_reg ( .D(g29241), .SI(g3255), .SE(n8911), .CLK(n9620), .Q(
        g1691), .QN(n8509) );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(n8911), .CLK(n9620), .Q(
        g2936), .QN(n8736) );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(n9077), .CLK(n9538), .Q(
        g5644), .QN(n5593) );
  SDFFX1 DFF_1284_Q_reg ( .D(g25707), .SI(g5644), .SE(n9107), .CLK(n9523), .Q(
        g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(n9106), .CLK(n9523), .Q(
        g5352), .QN(n8711) );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(n9106), .CLK(n9523), .Q(
        g8915) );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(n9088), .CLK(n9532), .Q(
        g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(n8940), .CLK(n9606), .Q(
        g2922) );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(n8940), .CLK(n9606), .Q(
        test_so90) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(n8989), .CLK(n9582), 
        .Q(g5893) );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(n8961), .CLK(n9595), .Q(
        g16603), .QN(n8547) );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(n9012), .CLK(n9570), 
        .Q(g6617) );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(n9036), .CLK(n9558), .Q(
        g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(n9113), .CLK(n9519), .Q(
        g4512) );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(n9098), .CLK(n9527), .Q(
        g5599) );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(n8914), .CLK(n9619), .Q(
        g3401), .QN(n5986) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(n8914), .CLK(n9619), .Q(
        g4366) );
  SDFFX1 DFF_1300_Q_reg ( .D(test_so26), .SI(g4366), .SE(n8914), .CLK(n9619), 
        .Q(g16722), .QN(n8672) );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(n8914), .CLK(n9619), 
        .Q(g29214), .QN(n5342) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g29214), .SE(n9096), .CLK(n9528), 
        .Q(g3129), .QN(n5861) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(n9040), .CLK(n9556), .Q(
        test_so91) );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(n8995), .CLK(n9578), 
        .Q(g5170), .QN(n8766) );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(n8908), .CLK(n9622), .Q(
        g26959) );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(n9078), .CLK(n9537), 
        .Q(g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(n9017), .CLK(n9568), .Q(
        g6299) );
  SDFFX1 DFF_1308_Q_reg ( .D(g7916), .SI(g6299), .SE(n8955), .CLK(n9599), .Q(
        g8416), .QN(n8803) );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(n9024), .CLK(n9564), .Q(
        g2079), .QN(n8790) );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(n9106), .CLK(n9523), .Q(
        g4698), .QN(n5862) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(n8933), .CLK(n9609), .Q(
        g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(n8993), .CLK(n9579), .Q(
        g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(n9060), .CLK(n9546), .Q(
        n9247), .QN(n15962) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(n9060), .CLK(n9546), .Q(
        g411), .QN(n5629) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(n8921), .CLK(n9616), .Q(
        test_so92) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(n8969), .CLK(n9591), 
        .Q(g3953) );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(n8969), .CLK(n9592), .Q(
        g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(n9031), .CLK(n9561), .Q(
        g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(n9030), .CLK(n9561), .Q(
        n9245) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(n8937), .CLK(n9607), .Q(
        g1300), .QN(n5483) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(n8976), .CLK(n9588), .Q(
        g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(n8978), .CLK(n9587), .Q(
        g5200), .QN(n8497) );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(n8923), .CLK(n9614), .Q(
        g4843), .QN(n8833) );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(n9108), .CLK(n9522), .Q(
        g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(g29249), .SI(g5046), .SE(n8918), .CLK(n9617), .Q(
        g2250), .QN(n8503) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(n9001), .CLK(n9576), .Q(
        g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(n8988), .CLK(n9582), 
        .Q(test_so93) );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(n8980), .CLK(n9586), 
        .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(g25734), .SI(g2453), .SE(n9078), .CLK(n9537), .Q(
        g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(n9078), .CLK(n9537), .Q(
        g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(n8941), .CLK(n9606), 
        .Q(g2912) );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(n8996), .CLK(n9578), .Q(
        g2357) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(n8938), .CLK(n9607), .Q(
        g8920) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(n9059), .CLK(n9547), .Q(
        g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(n9111), .CLK(n9521), .Q(
        g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(n8909), .CLK(n9622), .Q(
        g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(n9097), .CLK(n9528), .Q(
        g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(n9071), .CLK(n9540), .Q(
        g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(n8919), .CLK(n9617), .Q(
        test_so94), .QN(n8870) );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(n9111), .CLK(n9520), 
        .Q(g4519) );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(n9041), .CLK(n9556), .Q(
        g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(n9040), .CLK(n9556), .Q(
        g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(n9011), .CLK(n9571), .Q(
        g6657), .QN(n8484) );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(n9011), .CLK(n9571), .Q(
        g4552) );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(n8970), .CLK(n9591), .Q(
        g3893), .QN(n8502) );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(n9038), .CLK(n9557), .Q(
        g3211) );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(n8962), .CLK(n9595), .Q(
        g13049), .QN(n8689) );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(n8962), .CLK(n9595), 
        .Q(g16624), .QN(n8645) );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(n9090), .CLK(n9531), 
        .Q(g5595) );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(n9083), .CLK(n9535), .Q(
        g3614), .QN(n8487) );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(n9042), .CLK(n9555), .Q(
        test_so95) );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(n9040), .CLK(n9556), 
        .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(n9040), .CLK(n9556), .Q(
        g16686), .QN(n8643) );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(n8999), .CLK(n9577), 
        .Q(g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(n8975), .CLK(n9588), .Q(
        g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(n9011), .CLK(n9571), .Q(
        g4570) );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(n9029), .CLK(n9562), .Q(
        g5272), .QN(n8494) );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(n9003), .CLK(n9574), .Q(
        g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(n8950), .CLK(n9601), .Q(
        g728), .QN(n8475) );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(n8918), .CLK(n9617), .Q(
        g6295), .QN(n8491) );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(n9102), .CLK(n9525), .Q(
        g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(n8924), .CLK(n9614), .Q(
        g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(n8908), .CLK(n9622), .Q(
        test_so96), .QN(n8877) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(n8993), .CLK(n9579), 
        .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(n9097), .CLK(n9528), .Q(
        g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(n8964), .CLK(n9594), .Q(
        g4659), .QN(n8831) );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(n8934), .CLK(n9609), .Q(
        g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(n9054), .CLK(n9549), .Q(
        g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(n8991), .CLK(n9580), .Q(
        g2084), .QN(n8413) );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(n9009), .CLK(n9571), .Q(
        g3187) );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(n8933), .CLK(n9609), .Q(
        g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(n9005), .CLK(n9574), .Q(
        g2583) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(n9066), .CLK(n9543), .Q(
        n9240), .QN(DFF_1381_n1) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(n9066), .CLK(n9543), .Q(
        g1094) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(n8999), .CLK(n9577), .Q(
        test_so97), .QN(n8901) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(n8977), .CLK(n9588), 
        .Q(g4284), .QN(n8788) );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(n8915), .CLK(n9618), .Q(
        g3191), .QN(n8479) );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(n9070), .CLK(n9541), .Q(
        g4239), .QN(n8425) );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(n8946), .CLK(n9603), .Q(
        g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(n9087), .CLK(n9532), .Q(
        g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(n9087), .CLK(n9533), .Q(
        g534), .QN(n5490) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(n8968), .CLK(n9592), .Q(
        g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(n8991), .CLK(n9581), .Q(
        g2004) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(n9046), .CLK(n9553), .Q(
        g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(n8924), .CLK(n9614), .Q(
        g5456), .QN(n8802) );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(n8913), .CLK(n9620), .Q(
        n6007), .QN(n8463) );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(n8913), .CLK(n9620), .Q(
        test_so98), .QN(n8900) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(n9023), .CLK(n9564), 
        .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(n9106), .CLK(n9523), .Q(
        g5348), .QN(n8712) );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(n9039), .CLK(n9557), .Q(
        g3223) );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(n9076), .CLK(n9538), .Q(
        g2970), .QN(n8732) );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(n9077), .CLK(n9537), .Q(
        g5698), .QN(n8584) );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(n8978), .CLK(n9587), .Q(
        g5260) );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(n8957), .CLK(n9598), .Q(
        g1521), .QN(n5577) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(n8957), .CLK(n9598), .Q(
        g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(n9097), .CLK(n9528), .Q(
        g3115), .QN(n8394) );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(n9039), .CLK(n9556), .Q(
        g3251) );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(n9085), .CLK(n9533), .Q(
        g12832) );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(n9085), .CLK(n9533), 
        .Q(test_so99), .QN(n8876) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(n8947), .CLK(n9602), 
        .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(n8913), .CLK(n9619), .Q(
        g8342), .QN(n8359) );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(n9084), .CLK(n9534), .Q(
        g4515), .QN(n8714) );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(n9006), .CLK(n9573), .Q(
        g8787) );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(n9111), .CLK(n9521), .Q(
        g4300), .QN(n5639) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(n8907), .CLK(n9622), .Q(
        n9236), .QN(n15966) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(n9072), .CLK(n9540), .Q(
        g1379), .QN(n8793) );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(n8970), .CLK(n9591), .Q(
        g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(n8933), .CLK(n9610), 
        .Q(g1878) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(n9098), .CLK(n9527), .Q(
        g5619), .QN(n8480) );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(n9112), .CLK(n9520), .Q(
        g71) );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(n9112), .CLK(n9520), .Q(
        test_so100) );
  SDFFX1 DFF_748_Q_reg ( .D(n1465), .SI(g4704), .SE(n8951), .CLK(n9601), .Q(
        g22) );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(n8948), .CLK(n9602), .Q(
        g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(n9049), .CLK(n9552), .Q(
        g2729), .QN(n8469) );
  AND2X1 Trojan1 ( .IN1(Tj_TriggerIN1), .IN2(Tj_TriggerIN2), .Q(Tj_OUT1) );
  AND2X1 Trojan2 ( .IN1(Tj_TriggerIN3), .IN2(Tj_TriggerIN4), .Q(Tj_OUT2) );
  AND2X1 Trojan3 ( .IN1(Tj_TriggerIN5), .IN2(Tj_TriggerIN6), .Q(Tj_OUT3) );
  AND2X1 Trojan4 ( .IN1(Tj_TriggerIN7), .IN2(Tj_TriggerIN8), .Q(Tj_OUT4) );
  NOR4X0 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .QN(Tj_OUT1234) );
  AND2X1 Trojan5 ( .IN1(Tj_TriggerIN9), .IN2(Tj_TriggerIN10), .Q(Tj_OUT5) );
  INVX0 TrojanNOT_test_se ( .INP(n9119), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5), .IN3(test_se_NOT), 
        .Q(Tj_Trigger) );
  OR2X1 Trojan_Payload ( .IN1(Tj_Trigger), .IN2(g34028), .Q(g34028_Tj_Payload)
         );
  NBUFFX2 U8876 ( .INP(n9645), .Z(n9518) );
  NBUFFX2 U8877 ( .INP(n9645), .Z(n9517) );
  NBUFFX2 U8878 ( .INP(n9633), .Z(n9575) );
  NBUFFX2 U8879 ( .INP(n9644), .Z(n9523) );
  NBUFFX2 U8880 ( .INP(n9629), .Z(n9596) );
  NBUFFX2 U8881 ( .INP(n9630), .Z(n9592) );
  NBUFFX2 U8882 ( .INP(n9632), .Z(n9579) );
  NBUFFX2 U8883 ( .INP(n9633), .Z(n9576) );
  NBUFFX2 U8884 ( .INP(n9637), .Z(n9554) );
  NBUFFX2 U8885 ( .INP(n9639), .Z(n9545) );
  NBUFFX2 U8886 ( .INP(n9635), .Z(n9564) );
  NBUFFX2 U8887 ( .INP(n9637), .Z(n9558) );
  NBUFFX2 U8888 ( .INP(n9639), .Z(n9547) );
  NBUFFX2 U8889 ( .INP(n9641), .Z(n9535) );
  NBUFFX2 U8890 ( .INP(n9633), .Z(n9578) );
  NBUFFX2 U8891 ( .INP(n9634), .Z(n9570) );
  NBUFFX2 U8892 ( .INP(n9631), .Z(n9585) );
  NBUFFX2 U8893 ( .INP(n9630), .Z(n9593) );
  NBUFFX2 U8894 ( .INP(n9640), .Z(n9539) );
  NBUFFX2 U8895 ( .INP(n9641), .Z(n9538) );
  NBUFFX2 U8896 ( .INP(n9632), .Z(n9583) );
  NBUFFX2 U8897 ( .INP(n9629), .Z(n9597) );
  NBUFFX2 U8898 ( .INP(n9634), .Z(n9569) );
  NBUFFX2 U8899 ( .INP(n9637), .Z(n9556) );
  NBUFFX2 U8900 ( .INP(n9643), .Z(n9528) );
  NBUFFX2 U8901 ( .INP(n9644), .Z(n9519) );
  NBUFFX2 U8902 ( .INP(n9636), .Z(n9563) );
  NBUFFX2 U8903 ( .INP(n9634), .Z(n9572) );
  NBUFFX2 U8904 ( .INP(n9640), .Z(n9541) );
  NBUFFX2 U8905 ( .INP(n9627), .Z(n9607) );
  NBUFFX2 U8906 ( .INP(n9635), .Z(n9566) );
  NBUFFX2 U8907 ( .INP(n9632), .Z(n9581) );
  NBUFFX2 U8908 ( .INP(n9626), .Z(n9610) );
  NBUFFX2 U8909 ( .INP(n9628), .Z(n9603) );
  NBUFFX2 U8910 ( .INP(n9642), .Z(n9531) );
  NBUFFX2 U8911 ( .INP(n9627), .Z(n9608) );
  NBUFFX2 U8912 ( .INP(n9628), .Z(n9599) );
  NBUFFX2 U8913 ( .INP(n9642), .Z(n9533) );
  NBUFFX2 U8914 ( .INP(n9631), .Z(n9588) );
  NBUFFX2 U8915 ( .INP(n9638), .Z(n9549) );
  NBUFFX2 U8916 ( .INP(n9639), .Z(n9548) );
  NBUFFX2 U8917 ( .INP(n9625), .Z(n9618) );
  NBUFFX2 U8918 ( .INP(n9644), .Z(n9522) );
  NBUFFX2 U8919 ( .INP(n9625), .Z(n9616) );
  NBUFFX2 U8920 ( .INP(n9628), .Z(n9601) );
  NBUFFX2 U8921 ( .INP(n9637), .Z(n9557) );
  NBUFFX2 U8922 ( .INP(n9636), .Z(n9562) );
  NBUFFX2 U8923 ( .INP(n9625), .Z(n9614) );
  NBUFFX2 U8924 ( .INP(n9633), .Z(n9574) );
  NBUFFX2 U8925 ( .INP(n9630), .Z(n9590) );
  NBUFFX2 U8926 ( .INP(n9641), .Z(n9537) );
  NBUFFX2 U8927 ( .INP(n9626), .Z(n9609) );
  NBUFFX2 U8928 ( .INP(n9627), .Z(n9604) );
  NBUFFX2 U8929 ( .INP(n9631), .Z(n9586) );
  NBUFFX2 U8930 ( .INP(n9629), .Z(n9595) );
  NBUFFX2 U8931 ( .INP(n9631), .Z(n9587) );
  NBUFFX2 U8932 ( .INP(n9632), .Z(n9582) );
  NBUFFX2 U8933 ( .INP(n9636), .Z(n9559) );
  NBUFFX2 U8934 ( .INP(n9638), .Z(n9551) );
  NBUFFX2 U8935 ( .INP(n9638), .Z(n9550) );
  NBUFFX2 U8936 ( .INP(n9629), .Z(n9594) );
  NBUFFX2 U8937 ( .INP(n9640), .Z(n9542) );
  NBUFFX2 U8938 ( .INP(n9632), .Z(n9580) );
  NBUFFX2 U8939 ( .INP(n9625), .Z(n9615) );
  NBUFFX2 U8940 ( .INP(n9642), .Z(n9529) );
  NBUFFX2 U8941 ( .INP(n9640), .Z(n9540) );
  NBUFFX2 U8942 ( .INP(n9633), .Z(n9577) );
  NBUFFX2 U8943 ( .INP(n9630), .Z(n9589) );
  NBUFFX2 U8944 ( .INP(n9635), .Z(n9568) );
  NBUFFX2 U8945 ( .INP(n9635), .Z(n9565) );
  NBUFFX2 U8946 ( .INP(n9643), .Z(n9527) );
  NBUFFX2 U8947 ( .INP(n9643), .Z(n9526) );
  NBUFFX2 U8948 ( .INP(n9643), .Z(n9524) );
  NBUFFX2 U8949 ( .INP(n9628), .Z(n9602) );
  NBUFFX2 U8950 ( .INP(n9643), .Z(n9525) );
  NBUFFX2 U8951 ( .INP(n9631), .Z(n9584) );
  NBUFFX2 U8952 ( .INP(n9644), .Z(n9520) );
  NBUFFX2 U8953 ( .INP(n9634), .Z(n9571) );
  NBUFFX2 U8954 ( .INP(n9630), .Z(n9591) );
  NBUFFX2 U8955 ( .INP(n9640), .Z(n9543) );
  NBUFFX2 U8956 ( .INP(n9634), .Z(n9573) );
  NBUFFX2 U8957 ( .INP(n9625), .Z(n9617) );
  NBUFFX2 U8958 ( .INP(n9629), .Z(n9598) );
  NBUFFX2 U8959 ( .INP(n9636), .Z(n9560) );
  NBUFFX2 U8960 ( .INP(n9641), .Z(n9534) );
  NBUFFX2 U8961 ( .INP(n9641), .Z(n9536) );
  NBUFFX2 U8962 ( .INP(n9628), .Z(n9600) );
  NBUFFX2 U8963 ( .INP(n9639), .Z(n9546) );
  NBUFFX2 U8964 ( .INP(n9636), .Z(n9561) );
  NBUFFX2 U8965 ( .INP(n9626), .Z(n9613) );
  NBUFFX2 U8966 ( .INP(n9626), .Z(n9612) );
  NBUFFX2 U8967 ( .INP(n9638), .Z(n9552) );
  NBUFFX2 U8968 ( .INP(n9635), .Z(n9567) );
  NBUFFX2 U8969 ( .INP(n9639), .Z(n9544) );
  NBUFFX2 U8970 ( .INP(n9627), .Z(n9606) );
  NBUFFX2 U8971 ( .INP(n9627), .Z(n9605) );
  NBUFFX2 U8972 ( .INP(n9644), .Z(n9521) );
  NBUFFX2 U8973 ( .INP(n9642), .Z(n9530) );
  NBUFFX2 U8976 ( .INP(n9638), .Z(n9553) );
  NBUFFX2 U8977 ( .INP(n9637), .Z(n9555) );
  NBUFFX2 U8978 ( .INP(n9626), .Z(n9611) );
  NBUFFX2 U8979 ( .INP(n9642), .Z(n9532) );
  INVX0 U8980 ( .INP(n9226), .ZN(n9385) );
  INVX0 U8981 ( .INP(n9237), .ZN(n9411) );
  INVX0 U8982 ( .INP(n9239), .ZN(n9417) );
  INVX0 U8983 ( .INP(n9238), .ZN(n9415) );
  INVX0 U8984 ( .INP(n9239), .ZN(n9419) );
  INVX0 U8985 ( .INP(n9237), .ZN(n9412) );
  INVX0 U8986 ( .INP(n9238), .ZN(n9414) );
  INVX0 U8987 ( .INP(n9241), .ZN(n9420) );
  INVX0 U8988 ( .INP(n9237), .ZN(n9413) );
  INVX0 U8989 ( .INP(n9238), .ZN(n9416) );
  INVX0 U8990 ( .INP(n9239), .ZN(n9418) );
  INVX0 U8991 ( .INP(n9243), .ZN(n9426) );
  INVX0 U8992 ( .INP(n9242), .ZN(n9423) );
  INVX0 U8993 ( .INP(n9243), .ZN(n9428) );
  INVX0 U8994 ( .INP(n9243), .ZN(n9427) );
  INVX0 U8995 ( .INP(n9244), .ZN(n9429) );
  INVX0 U8996 ( .INP(n9242), .ZN(n9424) );
  INVX0 U8997 ( .INP(n9242), .ZN(n9425) );
  INVX0 U8998 ( .INP(n9241), .ZN(n9422) );
  INVX0 U8999 ( .INP(n9244), .ZN(n9430) );
  INVX0 U9000 ( .INP(n9282), .ZN(n9511) );
  INVX0 U9001 ( .INP(n9282), .ZN(n9512) );
  INVX0 U9002 ( .INP(n9283), .ZN(n9514) );
  INVX0 U9003 ( .INP(n9283), .ZN(n9513) );
  INVX0 U9004 ( .INP(n9283), .ZN(n9515) );
  INVX0 U9005 ( .INP(n9235), .ZN(n9408) );
  INVX0 U9006 ( .INP(n9235), .ZN(n9409) );
  INVX0 U9007 ( .INP(n9234), .ZN(n9407) );
  INVX0 U9008 ( .INP(n9235), .ZN(n9410) );
  INVX0 U9009 ( .INP(n9227), .ZN(n9386) );
  INVX0 U9010 ( .INP(n9271), .ZN(n9516) );
  INVX0 U9011 ( .INP(n9241), .ZN(n9421) );
  INVX0 U9012 ( .INP(n9226), .ZN(n9384) );
  INVX0 U9013 ( .INP(n9254), .ZN(n9453) );
  INVX0 U9014 ( .INP(n9250), .ZN(n9441) );
  INVX0 U9015 ( .INP(n9266), .ZN(n9481) );
  INVX0 U9016 ( .INP(n9253), .ZN(n9451) );
  INVX0 U9017 ( .INP(n9275), .ZN(n9499) );
  INVX0 U9018 ( .INP(n9277), .ZN(n9501) );
  INVX0 U9019 ( .INP(n9256), .ZN(n9458) );
  INVX0 U9020 ( .INP(n9258), .ZN(n9462) );
  INVX0 U9021 ( .INP(n9254), .ZN(n9455) );
  INVX0 U9022 ( .INP(n9260), .ZN(n9470) );
  INVX0 U9023 ( .INP(n9264), .ZN(n9479) );
  INVX0 U9024 ( .INP(n9246), .ZN(n9432) );
  INVX0 U9025 ( .INP(n9263), .ZN(n9474) );
  INVX0 U9026 ( .INP(n9258), .ZN(n9464) );
  INVX0 U9027 ( .INP(n9278), .ZN(n9506) );
  INVX0 U9028 ( .INP(n9250), .ZN(n9443) );
  INVX0 U9029 ( .INP(n9253), .ZN(n9452) );
  INVX0 U9030 ( .INP(n9270), .ZN(n9491) );
  INVX0 U9031 ( .INP(n9279), .ZN(n9508) );
  INVX0 U9032 ( .INP(n9275), .ZN(n9500) );
  INVX0 U9033 ( .INP(n9259), .ZN(n9465) );
  INVX0 U9034 ( .INP(n9249), .ZN(n9438) );
  INVX0 U9035 ( .INP(n9258), .ZN(n9463) );
  INVX0 U9036 ( .INP(n9254), .ZN(n9454) );
  INVX0 U9037 ( .INP(n9263), .ZN(n9476) );
  INVX0 U9038 ( .INP(n9261), .ZN(n9471) );
  INVX0 U9039 ( .INP(n9252), .ZN(n9448) );
  INVX0 U9040 ( .INP(n9268), .ZN(n9483) );
  INVX0 U9041 ( .INP(n9249), .ZN(n9440) );
  INVX0 U9042 ( .INP(n9282), .ZN(n9510) );
  INVX0 U9043 ( .INP(n9266), .ZN(n9482) );
  INVX0 U9044 ( .INP(n9272), .ZN(n9496) );
  INVX0 U9045 ( .INP(n9269), .ZN(n9486) );
  INVX0 U9046 ( .INP(n9257), .ZN(n9459) );
  INVX0 U9047 ( .INP(n9278), .ZN(n9505) );
  INVX0 U9048 ( .INP(n9251), .ZN(n9444) );
  INVX0 U9049 ( .INP(n9257), .ZN(n9460) );
  INVX0 U9050 ( .INP(n9256), .ZN(n9456) );
  INVX0 U9051 ( .INP(n9268), .ZN(n9484) );
  INVX0 U9052 ( .INP(n9268), .ZN(n9485) );
  INVX0 U9053 ( .INP(n9259), .ZN(n9466) );
  INVX0 U9054 ( .INP(n9269), .ZN(n9488) );
  INVX0 U9055 ( .INP(n9248), .ZN(n9437) );
  INVX0 U9056 ( .INP(n9277), .ZN(n9502) );
  INVX0 U9057 ( .INP(n9279), .ZN(n9507) );
  INVX0 U9058 ( .INP(n9248), .ZN(n9435) );
  INVX0 U9059 ( .INP(n9270), .ZN(n9490) );
  INVX0 U9060 ( .INP(n9252), .ZN(n9449) );
  INVX0 U9061 ( .INP(n9272), .ZN(n9495) );
  INVX0 U9062 ( .INP(n9275), .ZN(n9498) );
  INVX0 U9063 ( .INP(n9246), .ZN(n9434) );
  INVX0 U9064 ( .INP(n9256), .ZN(n9457) );
  INVX0 U9066 ( .INP(n9248), .ZN(n9436) );
  INVX0 U9067 ( .INP(n9266), .ZN(n9480) );
  INVX0 U9068 ( .INP(n9251), .ZN(n9446) );
  INVX0 U9069 ( .INP(n9253), .ZN(n9450) );
  INVX0 U9071 ( .INP(n9264), .ZN(n9478) );
  INVX0 U9072 ( .INP(n9261), .ZN(n9473) );
  INVX0 U9073 ( .INP(n9251), .ZN(n9445) );
  INVX0 U9074 ( .INP(n9272), .ZN(n9497) );
  INVX0 U9077 ( .INP(n9246), .ZN(n9433) );
  INVX0 U9078 ( .INP(n9271), .ZN(n9493) );
  INVX0 U9079 ( .INP(n9271), .ZN(n9492) );
  INVX0 U9081 ( .INP(n9263), .ZN(n9475) );
  INVX0 U9082 ( .INP(n9257), .ZN(n9461) );
  INVX0 U9083 ( .INP(n9244), .ZN(n9431) );
  INVX0 U9087 ( .INP(n9259), .ZN(n9467) );
  INVX0 U9088 ( .INP(n9279), .ZN(n9509) );
  INVX0 U9089 ( .INP(n9278), .ZN(n9504) );
  INVX0 U9091 ( .INP(n9269), .ZN(n9487) );
  INVX0 U9092 ( .INP(n9271), .ZN(n9494) );
  INVX0 U9093 ( .INP(n9260), .ZN(n9468) );
  INVX0 U9094 ( .INP(n9270), .ZN(n9489) );
  INVX0 U9095 ( .INP(n9249), .ZN(n9439) );
  INVX0 U9096 ( .INP(n9250), .ZN(n9442) );
  INVX0 U9097 ( .INP(n9252), .ZN(n9447) );
  INVX0 U9100 ( .INP(n9261), .ZN(n9472) );
  INVX0 U9102 ( .INP(n9260), .ZN(n9469) );
  INVX0 U9103 ( .INP(n9264), .ZN(n9477) );
  INVX0 U9104 ( .INP(n9277), .ZN(n9503) );
  INVX0 U9105 ( .INP(n9234), .ZN(n9406) );
  INVX0 U9106 ( .INP(n9226), .ZN(n9383) );
  INVX0 U9108 ( .INP(n9227), .ZN(n9387) );
  INVX0 U9109 ( .INP(n9227), .ZN(n9388) );
  INVX0 U9110 ( .INP(n9234), .ZN(n9405) );
  INVX0 U9112 ( .INP(n9228), .ZN(n9390) );
  INVX0 U9113 ( .INP(n9232), .ZN(n9399) );
  INVX0 U9114 ( .INP(n9230), .ZN(n9395) );
  INVX0 U9115 ( .INP(n9231), .ZN(n9398) );
  INVX0 U9117 ( .INP(n9229), .ZN(n9392) );
  INVX0 U9118 ( .INP(n9233), .ZN(n9404) );
  INVX0 U9119 ( .INP(n9232), .ZN(n9401) );
  INVX0 U9121 ( .INP(n9231), .ZN(n9396) );
  INVX0 U9122 ( .INP(n9233), .ZN(n9403) );
  INVX0 U9123 ( .INP(n9229), .ZN(n9394) );
  INVX0 U9125 ( .INP(n9232), .ZN(n9400) );
  INVX0 U9126 ( .INP(n9233), .ZN(n9402) );
  INVX0 U9127 ( .INP(n9228), .ZN(n9389) );
  INVX0 U9129 ( .INP(n9231), .ZN(n9397) );
  INVX0 U9130 ( .INP(n9228), .ZN(n9391) );
  INVX0 U9131 ( .INP(n9229), .ZN(n9393) );
  NBUFFX2 U9133 ( .INP(n9624), .Z(n9622) );
  NBUFFX2 U9134 ( .INP(n9624), .Z(n9619) );
  NBUFFX2 U9135 ( .INP(n9624), .Z(n9620) );
  NBUFFX2 U9137 ( .INP(n9624), .Z(n9621) );
  NBUFFX2 U9138 ( .INP(n9624), .Z(n9623) );
  NBUFFX2 U9139 ( .INP(n9190), .Z(n8907) );
  NBUFFX2 U9140 ( .INP(n9190), .Z(n8908) );
  NBUFFX2 U9141 ( .INP(n9190), .Z(n8909) );
  NBUFFX2 U9142 ( .INP(n9189), .Z(n8910) );
  NBUFFX2 U9143 ( .INP(n9189), .Z(n8911) );
  NBUFFX2 U9144 ( .INP(n9189), .Z(n8912) );
  NBUFFX2 U9145 ( .INP(n9188), .Z(n8913) );
  NBUFFX2 U9146 ( .INP(n9188), .Z(n8914) );
  NBUFFX2 U9147 ( .INP(n9188), .Z(n8915) );
  NBUFFX2 U9148 ( .INP(n9187), .Z(n8916) );
  NBUFFX2 U9149 ( .INP(n9187), .Z(n8917) );
  NBUFFX2 U9150 ( .INP(n9187), .Z(n8918) );
  NBUFFX2 U9151 ( .INP(n9186), .Z(n8919) );
  NBUFFX2 U9152 ( .INP(n9186), .Z(n8920) );
  NBUFFX2 U9153 ( .INP(n9186), .Z(n8921) );
  NBUFFX2 U9154 ( .INP(n9185), .Z(n8922) );
  NBUFFX2 U9155 ( .INP(n9185), .Z(n8923) );
  NBUFFX2 U9156 ( .INP(n9185), .Z(n8924) );
  NBUFFX2 U9157 ( .INP(n9184), .Z(n8925) );
  NBUFFX2 U9158 ( .INP(n9184), .Z(n8926) );
  NBUFFX2 U9159 ( .INP(n9184), .Z(n8927) );
  NBUFFX2 U9160 ( .INP(n9183), .Z(n8928) );
  NBUFFX2 U9161 ( .INP(n9183), .Z(n8929) );
  NBUFFX2 U9162 ( .INP(n9183), .Z(n8930) );
  NBUFFX2 U9163 ( .INP(n9182), .Z(n8931) );
  NBUFFX2 U9164 ( .INP(n9182), .Z(n8932) );
  NBUFFX2 U9165 ( .INP(n9182), .Z(n8933) );
  NBUFFX2 U9166 ( .INP(n9181), .Z(n8934) );
  NBUFFX2 U9167 ( .INP(n9181), .Z(n8935) );
  NBUFFX2 U9168 ( .INP(n9181), .Z(n8936) );
  NBUFFX2 U9169 ( .INP(n9180), .Z(n8937) );
  NBUFFX2 U9170 ( .INP(n9180), .Z(n8938) );
  NBUFFX2 U9171 ( .INP(n9180), .Z(n8939) );
  NBUFFX2 U9172 ( .INP(n9179), .Z(n8940) );
  NBUFFX2 U9173 ( .INP(n9179), .Z(n8941) );
  NBUFFX2 U9174 ( .INP(n9179), .Z(n8942) );
  NBUFFX2 U9175 ( .INP(n9178), .Z(n8943) );
  NBUFFX2 U9176 ( .INP(n9178), .Z(n8944) );
  NBUFFX2 U9177 ( .INP(n9178), .Z(n8945) );
  NBUFFX2 U9178 ( .INP(n9177), .Z(n8946) );
  NBUFFX2 U9179 ( .INP(n9177), .Z(n8947) );
  NBUFFX2 U9180 ( .INP(n9177), .Z(n8948) );
  NBUFFX2 U9181 ( .INP(n9176), .Z(n8949) );
  NBUFFX2 U9182 ( .INP(n9176), .Z(n8950) );
  NBUFFX2 U9183 ( .INP(n9176), .Z(n8951) );
  NBUFFX2 U9184 ( .INP(n9175), .Z(n8952) );
  NBUFFX2 U9185 ( .INP(n9175), .Z(n8953) );
  NBUFFX2 U9186 ( .INP(n9175), .Z(n8954) );
  NBUFFX2 U9187 ( .INP(n9174), .Z(n8955) );
  NBUFFX2 U9188 ( .INP(n9174), .Z(n8956) );
  NBUFFX2 U9189 ( .INP(n9174), .Z(n8957) );
  NBUFFX2 U9190 ( .INP(n9173), .Z(n8958) );
  NBUFFX2 U9191 ( .INP(n9173), .Z(n8959) );
  NBUFFX2 U9192 ( .INP(n9173), .Z(n8960) );
  NBUFFX2 U9193 ( .INP(n9172), .Z(n8961) );
  NBUFFX2 U9194 ( .INP(n9172), .Z(n8962) );
  NBUFFX2 U9195 ( .INP(n9172), .Z(n8963) );
  NBUFFX2 U9196 ( .INP(n9171), .Z(n8964) );
  NBUFFX2 U9197 ( .INP(n9171), .Z(n8965) );
  NBUFFX2 U9198 ( .INP(n9171), .Z(n8966) );
  NBUFFX2 U9199 ( .INP(n9170), .Z(n8967) );
  NBUFFX2 U9200 ( .INP(n9170), .Z(n8968) );
  NBUFFX2 U9201 ( .INP(n9170), .Z(n8969) );
  NBUFFX2 U9202 ( .INP(n9169), .Z(n8970) );
  NBUFFX2 U9203 ( .INP(n9169), .Z(n8971) );
  NBUFFX2 U9204 ( .INP(n9169), .Z(n8972) );
  NBUFFX2 U9205 ( .INP(n9168), .Z(n8973) );
  NBUFFX2 U9206 ( .INP(n9168), .Z(n8974) );
  NBUFFX2 U9207 ( .INP(n9168), .Z(n8975) );
  NBUFFX2 U9208 ( .INP(n9167), .Z(n8976) );
  NBUFFX2 U9209 ( .INP(n9167), .Z(n8977) );
  NBUFFX2 U9210 ( .INP(n9167), .Z(n8978) );
  NBUFFX2 U9211 ( .INP(n9166), .Z(n8979) );
  NBUFFX2 U9212 ( .INP(n9166), .Z(n8980) );
  NBUFFX2 U9213 ( .INP(n9166), .Z(n8981) );
  NBUFFX2 U9214 ( .INP(n9165), .Z(n8982) );
  NBUFFX2 U9215 ( .INP(n9165), .Z(n8983) );
  NBUFFX2 U9216 ( .INP(n9165), .Z(n8984) );
  NBUFFX2 U9217 ( .INP(n9164), .Z(n8985) );
  NBUFFX2 U9218 ( .INP(n9164), .Z(n8986) );
  NBUFFX2 U9219 ( .INP(n9164), .Z(n8987) );
  NBUFFX2 U9220 ( .INP(n9163), .Z(n8988) );
  NBUFFX2 U9221 ( .INP(n9163), .Z(n8989) );
  NBUFFX2 U9222 ( .INP(n9163), .Z(n8990) );
  NBUFFX2 U9223 ( .INP(n9162), .Z(n8991) );
  NBUFFX2 U9224 ( .INP(n9162), .Z(n8992) );
  NBUFFX2 U9225 ( .INP(n9162), .Z(n8993) );
  NBUFFX2 U9226 ( .INP(n9161), .Z(n8994) );
  NBUFFX2 U9227 ( .INP(n9161), .Z(n8995) );
  NBUFFX2 U9228 ( .INP(n9161), .Z(n8996) );
  NBUFFX2 U9229 ( .INP(n9160), .Z(n8997) );
  NBUFFX2 U9230 ( .INP(n9160), .Z(n8998) );
  NBUFFX2 U9231 ( .INP(n9160), .Z(n8999) );
  NBUFFX2 U9232 ( .INP(n9159), .Z(n9000) );
  NBUFFX2 U9233 ( .INP(n9159), .Z(n9001) );
  NBUFFX2 U9234 ( .INP(n9159), .Z(n9002) );
  NBUFFX2 U9235 ( .INP(n9158), .Z(n9003) );
  NBUFFX2 U9236 ( .INP(n9158), .Z(n9004) );
  NBUFFX2 U9237 ( .INP(n9158), .Z(n9005) );
  NBUFFX2 U9238 ( .INP(n9157), .Z(n9006) );
  NBUFFX2 U9239 ( .INP(n9157), .Z(n9007) );
  NBUFFX2 U9240 ( .INP(n9157), .Z(n9008) );
  NBUFFX2 U9241 ( .INP(n9156), .Z(n9009) );
  NBUFFX2 U9242 ( .INP(n9156), .Z(n9010) );
  NBUFFX2 U9243 ( .INP(n9156), .Z(n9011) );
  NBUFFX2 U9244 ( .INP(n9155), .Z(n9012) );
  NBUFFX2 U9245 ( .INP(n9155), .Z(n9013) );
  NBUFFX2 U9246 ( .INP(n9155), .Z(n9014) );
  NBUFFX2 U9247 ( .INP(n9154), .Z(n9015) );
  NBUFFX2 U9248 ( .INP(n9154), .Z(n9016) );
  NBUFFX2 U9249 ( .INP(n9154), .Z(n9017) );
  NBUFFX2 U9250 ( .INP(n9153), .Z(n9018) );
  NBUFFX2 U9251 ( .INP(n9153), .Z(n9019) );
  NBUFFX2 U9252 ( .INP(n9153), .Z(n9020) );
  NBUFFX2 U9253 ( .INP(n9152), .Z(n9021) );
  NBUFFX2 U9254 ( .INP(n9152), .Z(n9022) );
  NBUFFX2 U9255 ( .INP(n9152), .Z(n9023) );
  NBUFFX2 U9256 ( .INP(n9151), .Z(n9024) );
  NBUFFX2 U9257 ( .INP(n9151), .Z(n9025) );
  NBUFFX2 U9258 ( .INP(n9151), .Z(n9026) );
  NBUFFX2 U9259 ( .INP(n9150), .Z(n9027) );
  NBUFFX2 U9260 ( .INP(n9150), .Z(n9028) );
  NBUFFX2 U9261 ( .INP(n9150), .Z(n9029) );
  NBUFFX2 U9262 ( .INP(n9149), .Z(n9030) );
  NBUFFX2 U9263 ( .INP(n9149), .Z(n9031) );
  NBUFFX2 U9264 ( .INP(n9149), .Z(n9032) );
  NBUFFX2 U9265 ( .INP(n9148), .Z(n9033) );
  NBUFFX2 U9266 ( .INP(n9148), .Z(n9034) );
  NBUFFX2 U9267 ( .INP(n9148), .Z(n9035) );
  NBUFFX2 U9268 ( .INP(n9147), .Z(n9036) );
  NBUFFX2 U9269 ( .INP(n9147), .Z(n9037) );
  NBUFFX2 U9270 ( .INP(n9147), .Z(n9038) );
  NBUFFX2 U9271 ( .INP(n9146), .Z(n9039) );
  NBUFFX2 U9272 ( .INP(n9146), .Z(n9040) );
  NBUFFX2 U9273 ( .INP(n9146), .Z(n9041) );
  NBUFFX2 U9274 ( .INP(n9145), .Z(n9042) );
  NBUFFX2 U9275 ( .INP(n9145), .Z(n9043) );
  NBUFFX2 U9276 ( .INP(n9145), .Z(n9044) );
  NBUFFX2 U9277 ( .INP(n9144), .Z(n9045) );
  NBUFFX2 U9278 ( .INP(n9144), .Z(n9046) );
  NBUFFX2 U9279 ( .INP(n9144), .Z(n9047) );
  NBUFFX2 U9280 ( .INP(n9143), .Z(n9048) );
  NBUFFX2 U9281 ( .INP(n9143), .Z(n9049) );
  NBUFFX2 U9282 ( .INP(n9143), .Z(n9050) );
  NBUFFX2 U9283 ( .INP(n9142), .Z(n9051) );
  NBUFFX2 U9284 ( .INP(n9142), .Z(n9052) );
  NBUFFX2 U9285 ( .INP(n9142), .Z(n9053) );
  NBUFFX2 U9286 ( .INP(n9141), .Z(n9054) );
  NBUFFX2 U9287 ( .INP(n9141), .Z(n9055) );
  NBUFFX2 U9288 ( .INP(n9141), .Z(n9056) );
  NBUFFX2 U9289 ( .INP(n9140), .Z(n9057) );
  NBUFFX2 U9290 ( .INP(n9140), .Z(n9058) );
  NBUFFX2 U9291 ( .INP(n9140), .Z(n9059) );
  NBUFFX2 U9292 ( .INP(n9139), .Z(n9060) );
  NBUFFX2 U9293 ( .INP(n9139), .Z(n9061) );
  NBUFFX2 U9294 ( .INP(n9139), .Z(n9062) );
  NBUFFX2 U9295 ( .INP(n9138), .Z(n9063) );
  NBUFFX2 U9296 ( .INP(n9138), .Z(n9064) );
  NBUFFX2 U9297 ( .INP(n9138), .Z(n9065) );
  NBUFFX2 U9298 ( .INP(n9137), .Z(n9066) );
  NBUFFX2 U9299 ( .INP(n9137), .Z(n9067) );
  NBUFFX2 U9300 ( .INP(n9137), .Z(n9068) );
  NBUFFX2 U9301 ( .INP(n9136), .Z(n9069) );
  NBUFFX2 U9302 ( .INP(n9136), .Z(n9070) );
  NBUFFX2 U9303 ( .INP(n9136), .Z(n9071) );
  NBUFFX2 U9304 ( .INP(n9135), .Z(n9072) );
  NBUFFX2 U9305 ( .INP(n9135), .Z(n9073) );
  NBUFFX2 U9306 ( .INP(n9135), .Z(n9074) );
  NBUFFX2 U9307 ( .INP(n9134), .Z(n9075) );
  NBUFFX2 U9308 ( .INP(n9134), .Z(n9076) );
  NBUFFX2 U9309 ( .INP(n9134), .Z(n9077) );
  NBUFFX2 U9310 ( .INP(n9133), .Z(n9078) );
  NBUFFX2 U9311 ( .INP(n9133), .Z(n9079) );
  NBUFFX2 U9312 ( .INP(n9133), .Z(n9080) );
  NBUFFX2 U9313 ( .INP(n9132), .Z(n9081) );
  NBUFFX2 U9314 ( .INP(n9132), .Z(n9082) );
  NBUFFX2 U9316 ( .INP(n9132), .Z(n9083) );
  NBUFFX2 U9317 ( .INP(n9131), .Z(n9084) );
  NBUFFX2 U9318 ( .INP(n9131), .Z(n9085) );
  NBUFFX2 U9319 ( .INP(n9131), .Z(n9086) );
  NBUFFX2 U9320 ( .INP(n9130), .Z(n9087) );
  NBUFFX2 U9321 ( .INP(n9130), .Z(n9088) );
  NBUFFX2 U9322 ( .INP(n9130), .Z(n9089) );
  NBUFFX2 U9323 ( .INP(n9129), .Z(n9090) );
  NBUFFX2 U9324 ( .INP(n9129), .Z(n9091) );
  NBUFFX2 U9325 ( .INP(n9129), .Z(n9092) );
  NBUFFX2 U9326 ( .INP(n9128), .Z(n9093) );
  NBUFFX2 U9327 ( .INP(n9128), .Z(n9094) );
  NBUFFX2 U9328 ( .INP(n9128), .Z(n9095) );
  NBUFFX2 U9329 ( .INP(n9127), .Z(n9096) );
  NBUFFX2 U9330 ( .INP(n9127), .Z(n9097) );
  NBUFFX2 U9331 ( .INP(n9127), .Z(n9098) );
  NBUFFX2 U9332 ( .INP(n9126), .Z(n9099) );
  NBUFFX2 U9333 ( .INP(n9126), .Z(n9100) );
  NBUFFX2 U9334 ( .INP(n9126), .Z(n9101) );
  NBUFFX2 U9335 ( .INP(n9125), .Z(n9102) );
  NBUFFX2 U9336 ( .INP(n9125), .Z(n9103) );
  NBUFFX2 U9337 ( .INP(n9125), .Z(n9104) );
  NBUFFX2 U9338 ( .INP(n9124), .Z(n9105) );
  NBUFFX2 U9339 ( .INP(n9124), .Z(n9106) );
  NBUFFX2 U9340 ( .INP(n9124), .Z(n9107) );
  NBUFFX2 U9341 ( .INP(n9123), .Z(n9108) );
  NBUFFX2 U9342 ( .INP(n9123), .Z(n9109) );
  NBUFFX2 U9343 ( .INP(n9123), .Z(n9110) );
  NBUFFX2 U9344 ( .INP(n9122), .Z(n9111) );
  NBUFFX2 U9345 ( .INP(n9122), .Z(n9112) );
  NBUFFX2 U9346 ( .INP(n9122), .Z(n9113) );
  NBUFFX2 U9347 ( .INP(n9121), .Z(n9114) );
  NBUFFX2 U9348 ( .INP(n9121), .Z(n9115) );
  NBUFFX2 U9349 ( .INP(n9121), .Z(n9116) );
  NBUFFX2 U9350 ( .INP(n9120), .Z(n9117) );
  NBUFFX2 U9351 ( .INP(n9120), .Z(n9118) );
  NBUFFX2 U9352 ( .INP(n9120), .Z(n9119) );
  NBUFFX2 U9353 ( .INP(n9214), .Z(n9120) );
  NBUFFX2 U9354 ( .INP(n9214), .Z(n9121) );
  NBUFFX2 U9355 ( .INP(n9213), .Z(n9122) );
  NBUFFX2 U9356 ( .INP(n9213), .Z(n9123) );
  NBUFFX2 U9357 ( .INP(n9213), .Z(n9124) );
  NBUFFX2 U9358 ( .INP(n9212), .Z(n9125) );
  NBUFFX2 U9359 ( .INP(n9212), .Z(n9126) );
  NBUFFX2 U9360 ( .INP(n9212), .Z(n9127) );
  NBUFFX2 U9361 ( .INP(n9211), .Z(n9128) );
  NBUFFX2 U9362 ( .INP(n9211), .Z(n9129) );
  NBUFFX2 U9363 ( .INP(n9211), .Z(n9130) );
  NBUFFX2 U9364 ( .INP(n9210), .Z(n9131) );
  NBUFFX2 U9365 ( .INP(n9210), .Z(n9132) );
  NBUFFX2 U9366 ( .INP(n9210), .Z(n9133) );
  NBUFFX2 U9367 ( .INP(n9209), .Z(n9134) );
  NBUFFX2 U9368 ( .INP(n9209), .Z(n9135) );
  NBUFFX2 U9369 ( .INP(n9209), .Z(n9136) );
  NBUFFX2 U9370 ( .INP(n9208), .Z(n9137) );
  NBUFFX2 U9371 ( .INP(n9208), .Z(n9138) );
  NBUFFX2 U9372 ( .INP(n9208), .Z(n9139) );
  NBUFFX2 U9373 ( .INP(n9207), .Z(n9140) );
  NBUFFX2 U9374 ( .INP(n9207), .Z(n9141) );
  NBUFFX2 U9375 ( .INP(n9207), .Z(n9142) );
  NBUFFX2 U9376 ( .INP(n9206), .Z(n9143) );
  NBUFFX2 U9377 ( .INP(n9206), .Z(n9144) );
  NBUFFX2 U9378 ( .INP(n9206), .Z(n9145) );
  NBUFFX2 U9379 ( .INP(n9205), .Z(n9146) );
  NBUFFX2 U9380 ( .INP(n9205), .Z(n9147) );
  NBUFFX2 U9381 ( .INP(n9205), .Z(n9148) );
  NBUFFX2 U9382 ( .INP(n9204), .Z(n9149) );
  NBUFFX2 U9383 ( .INP(n9204), .Z(n9150) );
  NBUFFX2 U9384 ( .INP(n9204), .Z(n9151) );
  NBUFFX2 U9385 ( .INP(n9203), .Z(n9152) );
  NBUFFX2 U9386 ( .INP(n9203), .Z(n9153) );
  NBUFFX2 U9387 ( .INP(n9203), .Z(n9154) );
  NBUFFX2 U9388 ( .INP(n9202), .Z(n9155) );
  NBUFFX2 U9389 ( .INP(n9202), .Z(n9156) );
  NBUFFX2 U9390 ( .INP(n9202), .Z(n9157) );
  NBUFFX2 U9391 ( .INP(n9201), .Z(n9158) );
  NBUFFX2 U9392 ( .INP(n9201), .Z(n9159) );
  NBUFFX2 U9393 ( .INP(n9201), .Z(n9160) );
  NBUFFX2 U9394 ( .INP(n9200), .Z(n9161) );
  NBUFFX2 U9395 ( .INP(n9200), .Z(n9162) );
  NBUFFX2 U9396 ( .INP(n9200), .Z(n9163) );
  NBUFFX2 U9397 ( .INP(n9199), .Z(n9164) );
  NBUFFX2 U9398 ( .INP(n9199), .Z(n9165) );
  NBUFFX2 U9399 ( .INP(n9199), .Z(n9166) );
  NBUFFX2 U9400 ( .INP(n9198), .Z(n9167) );
  NBUFFX2 U9401 ( .INP(n9198), .Z(n9168) );
  NBUFFX2 U9402 ( .INP(n9198), .Z(n9169) );
  NBUFFX2 U9403 ( .INP(n9197), .Z(n9170) );
  NBUFFX2 U9404 ( .INP(n9197), .Z(n9171) );
  NBUFFX2 U9405 ( .INP(n9197), .Z(n9172) );
  NBUFFX2 U9406 ( .INP(n9196), .Z(n9173) );
  NBUFFX2 U9407 ( .INP(n9196), .Z(n9174) );
  NBUFFX2 U9408 ( .INP(n9196), .Z(n9175) );
  NBUFFX2 U9409 ( .INP(n9195), .Z(n9176) );
  NBUFFX2 U9410 ( .INP(n9195), .Z(n9177) );
  NBUFFX2 U9411 ( .INP(n9195), .Z(n9178) );
  NBUFFX2 U9412 ( .INP(n9194), .Z(n9179) );
  NBUFFX2 U9413 ( .INP(n9194), .Z(n9180) );
  NBUFFX2 U9414 ( .INP(n9194), .Z(n9181) );
  NBUFFX2 U9415 ( .INP(n9193), .Z(n9182) );
  NBUFFX2 U9416 ( .INP(n9193), .Z(n9183) );
  NBUFFX2 U9417 ( .INP(n9193), .Z(n9184) );
  NBUFFX2 U9418 ( .INP(n9192), .Z(n9185) );
  NBUFFX2 U9419 ( .INP(n9192), .Z(n9186) );
  NBUFFX2 U9420 ( .INP(n9192), .Z(n9187) );
  NBUFFX2 U9421 ( .INP(n9191), .Z(n9188) );
  NBUFFX2 U9422 ( .INP(n9191), .Z(n9189) );
  NBUFFX2 U9423 ( .INP(n9191), .Z(n9190) );
  NBUFFX2 U9424 ( .INP(n9222), .Z(n9191) );
  NBUFFX2 U9425 ( .INP(n9222), .Z(n9192) );
  NBUFFX2 U9426 ( .INP(n9222), .Z(n9193) );
  NBUFFX2 U9427 ( .INP(n9221), .Z(n9194) );
  NBUFFX2 U9428 ( .INP(n9221), .Z(n9195) );
  NBUFFX2 U9429 ( .INP(n9221), .Z(n9196) );
  NBUFFX2 U9430 ( .INP(n9220), .Z(n9197) );
  NBUFFX2 U9431 ( .INP(n9220), .Z(n9198) );
  NBUFFX2 U9432 ( .INP(n9220), .Z(n9199) );
  NBUFFX2 U9433 ( .INP(n9219), .Z(n9200) );
  NBUFFX2 U9434 ( .INP(n9219), .Z(n9201) );
  NBUFFX2 U9435 ( .INP(n9219), .Z(n9202) );
  NBUFFX2 U9436 ( .INP(n9218), .Z(n9203) );
  NBUFFX2 U9437 ( .INP(n9218), .Z(n9204) );
  NBUFFX2 U9438 ( .INP(n9218), .Z(n9205) );
  NBUFFX2 U9439 ( .INP(n9217), .Z(n9206) );
  NBUFFX2 U9440 ( .INP(n9217), .Z(n9207) );
  NBUFFX2 U9441 ( .INP(n9217), .Z(n9208) );
  NBUFFX2 U9442 ( .INP(n9216), .Z(n9209) );
  NBUFFX2 U9443 ( .INP(n9216), .Z(n9210) );
  NBUFFX2 U9444 ( .INP(n9216), .Z(n9211) );
  NBUFFX2 U9445 ( .INP(n9215), .Z(n9212) );
  NBUFFX2 U9446 ( .INP(n9215), .Z(n9213) );
  NBUFFX2 U9447 ( .INP(n9215), .Z(n9214) );
  NBUFFX2 U9448 ( .INP(n9225), .Z(n9215) );
  NBUFFX2 U9449 ( .INP(n9225), .Z(n9216) );
  NBUFFX2 U9450 ( .INP(n9224), .Z(n9217) );
  NBUFFX2 U9451 ( .INP(n9224), .Z(n9218) );
  NBUFFX2 U9452 ( .INP(n9224), .Z(n9219) );
  NBUFFX2 U9454 ( .INP(n9223), .Z(n9220) );
  NBUFFX2 U9455 ( .INP(n9223), .Z(n9221) );
  NBUFFX2 U9456 ( .INP(n9223), .Z(n9222) );
  NBUFFX2 U9457 ( .INP(test_se), .Z(n9223) );
  NBUFFX2 U9458 ( .INP(test_se), .Z(n9224) );
  NBUFFX2 U9459 ( .INP(test_se), .Z(n9225) );
  NBUFFX2 U9460 ( .INP(n9304), .Z(n9226) );
  NBUFFX2 U9461 ( .INP(n9304), .Z(n9227) );
  NBUFFX2 U9462 ( .INP(n9301), .Z(n9228) );
  NBUFFX2 U9463 ( .INP(n9301), .Z(n9229) );
  NBUFFX2 U9464 ( .INP(n9301), .Z(n9230) );
  NBUFFX2 U9465 ( .INP(n9300), .Z(n9231) );
  NBUFFX2 U9466 ( .INP(n9300), .Z(n9232) );
  NBUFFX2 U9467 ( .INP(n9299), .Z(n9233) );
  NBUFFX2 U9468 ( .INP(n9299), .Z(n9234) );
  NBUFFX2 U9469 ( .INP(n9299), .Z(n9235) );
  NBUFFX2 U9470 ( .INP(n9298), .Z(n9237) );
  NBUFFX2 U9471 ( .INP(n9298), .Z(n9238) );
  NBUFFX2 U9472 ( .INP(n9298), .Z(n9239) );
  NBUFFX2 U9473 ( .INP(n9297), .Z(n9241) );
  NBUFFX2 U9474 ( .INP(n9297), .Z(n9242) );
  NBUFFX2 U9475 ( .INP(n9297), .Z(n9243) );
  NBUFFX2 U9476 ( .INP(n9296), .Z(n9244) );
  NBUFFX2 U9477 ( .INP(n9296), .Z(n9246) );
  NBUFFX2 U9478 ( .INP(n9296), .Z(n9248) );
  NBUFFX2 U9479 ( .INP(n9293), .Z(n9249) );
  NBUFFX2 U9480 ( .INP(n9293), .Z(n9250) );
  NBUFFX2 U9481 ( .INP(n9292), .Z(n9251) );
  NBUFFX2 U9482 ( .INP(n9292), .Z(n9252) );
  NBUFFX2 U9483 ( .INP(n9292), .Z(n9253) );
  NBUFFX2 U9484 ( .INP(n9291), .Z(n9254) );
  NBUFFX2 U9485 ( .INP(n9291), .Z(n9256) );
  NBUFFX2 U9486 ( .INP(n9290), .Z(n9257) );
  NBUFFX2 U9487 ( .INP(n9290), .Z(n9258) );
  NBUFFX2 U9488 ( .INP(n9289), .Z(n9259) );
  NBUFFX2 U9489 ( .INP(n9289), .Z(n9260) );
  NBUFFX2 U9490 ( .INP(n9289), .Z(n9261) );
  NBUFFX2 U9491 ( .INP(n9288), .Z(n9263) );
  NBUFFX2 U9492 ( .INP(n9288), .Z(n9264) );
  NBUFFX2 U9493 ( .INP(n9288), .Z(n9266) );
  NBUFFX2 U9494 ( .INP(n9287), .Z(n9268) );
  NBUFFX2 U9495 ( .INP(n9287), .Z(n9269) );
  NBUFFX2 U9496 ( .INP(n9287), .Z(n9270) );
  NBUFFX2 U9497 ( .INP(n9286), .Z(n9271) );
  NBUFFX2 U9498 ( .INP(n9286), .Z(n9272) );
  NBUFFX2 U9499 ( .INP(n9286), .Z(n9275) );
  NBUFFX2 U9500 ( .INP(n9285), .Z(n9277) );
  NBUFFX2 U9501 ( .INP(n9285), .Z(n9278) );
  NBUFFX2 U9502 ( .INP(n9285), .Z(n9279) );
  NBUFFX2 U9503 ( .INP(n9284), .Z(n9282) );
  NBUFFX2 U9504 ( .INP(n9284), .Z(n9283) );
  NBUFFX2 U9505 ( .INP(n9311), .Z(n9284) );
  NBUFFX2 U9506 ( .INP(n9311), .Z(n9285) );
  NBUFFX2 U9507 ( .INP(n9310), .Z(n9286) );
  NBUFFX2 U9508 ( .INP(n9310), .Z(n9287) );
  NBUFFX2 U9509 ( .INP(n9310), .Z(n9288) );
  NBUFFX2 U9510 ( .INP(n9309), .Z(n9289) );
  NBUFFX2 U9511 ( .INP(n9309), .Z(n9290) );
  NBUFFX2 U9512 ( .INP(n9309), .Z(n9291) );
  NBUFFX2 U9513 ( .INP(n9308), .Z(n9292) );
  NBUFFX2 U9514 ( .INP(n9308), .Z(n9293) );
  NBUFFX2 U9515 ( .INP(n9308), .Z(n9296) );
  NBUFFX2 U9516 ( .INP(n9307), .Z(n9297) );
  NBUFFX2 U9517 ( .INP(n9307), .Z(n9298) );
  NBUFFX2 U9518 ( .INP(n9307), .Z(n9299) );
  NBUFFX2 U9519 ( .INP(n9305), .Z(n9300) );
  NBUFFX2 U9520 ( .INP(n9305), .Z(n9301) );
  NBUFFX2 U9521 ( .INP(n9305), .Z(n9304) );
  NBUFFX2 U9522 ( .INP(g35), .Z(n9305) );
  NBUFFX2 U9523 ( .INP(g35), .Z(n9307) );
  NBUFFX2 U9524 ( .INP(g35), .Z(n9308) );
  NBUFFX2 U9525 ( .INP(g35), .Z(n9309) );
  NBUFFX2 U9526 ( .INP(g35), .Z(n9310) );
  NBUFFX2 U9527 ( .INP(g35), .Z(n9311) );
  INVX0 U9528 ( .INP(n9429), .ZN(n9313) );
  INVX0 U9529 ( .INP(n9430), .ZN(n9315) );
  INVX0 U9530 ( .INP(n9430), .ZN(n9316) );
  INVX0 U9531 ( .INP(n9426), .ZN(n9317) );
  INVX0 U9532 ( .INP(n9430), .ZN(n9318) );
  INVX0 U9533 ( .INP(n9430), .ZN(n9319) );
  INVX0 U9534 ( .INP(n9429), .ZN(n9320) );
  INVX0 U9535 ( .INP(n9429), .ZN(n9321) );
  INVX0 U9536 ( .INP(n9429), .ZN(n9323) );
  INVX0 U9537 ( .INP(n9428), .ZN(n9326) );
  INVX0 U9538 ( .INP(n9429), .ZN(n9328) );
  INVX0 U9539 ( .INP(n9428), .ZN(n9329) );
  INVX0 U9540 ( .INP(n9429), .ZN(n9330) );
  INVX0 U9541 ( .INP(n9425), .ZN(n9331) );
  INVX0 U9542 ( .INP(n9428), .ZN(n9333) );
  INVX0 U9543 ( .INP(n9428), .ZN(n9334) );
  INVX0 U9544 ( .INP(n9426), .ZN(n9335) );
  INVX0 U9545 ( .INP(n9427), .ZN(n9337) );
  INVX0 U9546 ( .INP(n9428), .ZN(n9338) );
  INVX0 U9547 ( .INP(n9428), .ZN(n9339) );
  INVX0 U9548 ( .INP(n9427), .ZN(n9341) );
  INVX0 U9549 ( .INP(n9427), .ZN(n9342) );
  INVX0 U9550 ( .INP(n9427), .ZN(n9343) );
  INVX0 U9551 ( .INP(n9427), .ZN(n9344) );
  INVX0 U9552 ( .INP(n9427), .ZN(n9345) );
  INVX0 U9553 ( .INP(n9426), .ZN(n9346) );
  INVX0 U9554 ( .INP(n9426), .ZN(n9347) );
  INVX0 U9555 ( .INP(n9426), .ZN(n9349) );
  INVX0 U9556 ( .INP(n9423), .ZN(n9350) );
  INVX0 U9557 ( .INP(n9425), .ZN(n9353) );
  INVX0 U9558 ( .INP(n9426), .ZN(n9354) );
  INVX0 U9559 ( .INP(n9425), .ZN(n9355) );
  INVX0 U9560 ( .INP(n9425), .ZN(n9356) );
  INVX0 U9561 ( .INP(n9425), .ZN(n9358) );
  INVX0 U9562 ( .INP(n9425), .ZN(n9359) );
  INVX0 U9563 ( .INP(n9423), .ZN(n9360) );
  INVX0 U9564 ( .INP(n9424), .ZN(n9361) );
  INVX0 U9565 ( .INP(n9424), .ZN(n9362) );
  INVX0 U9566 ( .INP(n9424), .ZN(n9363) );
  INVX0 U9567 ( .INP(n9424), .ZN(n9364) );
  INVX0 U9568 ( .INP(n9424), .ZN(n9365) );
  INVX0 U9569 ( .INP(n9424), .ZN(n9366) );
  INVX0 U9570 ( .INP(n9421), .ZN(n9368) );
  INVX0 U9571 ( .INP(n9423), .ZN(n9369) );
  INVX0 U9572 ( .INP(n9423), .ZN(n9370) );
  INVX0 U9573 ( .INP(n9423), .ZN(n9371) );
  INVX0 U9574 ( .INP(n9422), .ZN(n9372) );
  INVX0 U9575 ( .INP(n9423), .ZN(n9373) );
  INVX0 U9576 ( .INP(n9422), .ZN(n9374) );
  INVX0 U9577 ( .INP(n9422), .ZN(n9375) );
  INVX0 U9578 ( .INP(n9422), .ZN(n9376) );
  INVX0 U9579 ( .INP(n9421), .ZN(n9377) );
  INVX0 U9580 ( .INP(n9422), .ZN(n9378) );
  INVX0 U9581 ( .INP(n9422), .ZN(n9379) );
  INVX0 U9582 ( .INP(n9421), .ZN(n9380) );
  INVX0 U9583 ( .INP(n9421), .ZN(n9381) );
  INVX0 U9584 ( .INP(n9421), .ZN(n9382) );
  NBUFFX2 U9585 ( .INP(n9653), .Z(n9624) );
  NBUFFX2 U9586 ( .INP(n9652), .Z(n9625) );
  NBUFFX2 U9587 ( .INP(n9652), .Z(n9626) );
  NBUFFX2 U9588 ( .INP(n9652), .Z(n9627) );
  NBUFFX2 U9589 ( .INP(n9651), .Z(n9628) );
  NBUFFX2 U9590 ( .INP(n9651), .Z(n9629) );
  NBUFFX2 U9591 ( .INP(n9651), .Z(n9630) );
  NBUFFX2 U9592 ( .INP(n9650), .Z(n9631) );
  NBUFFX2 U9593 ( .INP(n9650), .Z(n9632) );
  NBUFFX2 U9594 ( .INP(n9650), .Z(n9633) );
  NBUFFX2 U9595 ( .INP(n9649), .Z(n9634) );
  NBUFFX2 U9596 ( .INP(n9649), .Z(n9635) );
  NBUFFX2 U9597 ( .INP(n9649), .Z(n9636) );
  NBUFFX2 U9598 ( .INP(n9648), .Z(n9637) );
  NBUFFX2 U9599 ( .INP(n9648), .Z(n9638) );
  NBUFFX2 U9600 ( .INP(n9648), .Z(n9639) );
  NBUFFX2 U9601 ( .INP(n9647), .Z(n9640) );
  NBUFFX2 U9602 ( .INP(n9647), .Z(n9641) );
  NBUFFX2 U9603 ( .INP(n9647), .Z(n9642) );
  NBUFFX2 U9604 ( .INP(n9646), .Z(n9643) );
  NBUFFX2 U9605 ( .INP(n9646), .Z(n9644) );
  NBUFFX2 U9606 ( .INP(n9646), .Z(n9645) );
  NBUFFX2 U9607 ( .INP(n9656), .Z(n9646) );
  NBUFFX2 U9608 ( .INP(n9656), .Z(n9647) );
  NBUFFX2 U9609 ( .INP(n9655), .Z(n9648) );
  NBUFFX2 U9610 ( .INP(n9655), .Z(n9649) );
  NBUFFX2 U9611 ( .INP(n9655), .Z(n9650) );
  NBUFFX2 U9612 ( .INP(n9654), .Z(n9651) );
  NBUFFX2 U9613 ( .INP(n9654), .Z(n9652) );
  NBUFFX2 U9614 ( .INP(n9654), .Z(n9653) );
  NBUFFX2 U9615 ( .INP(CK), .Z(n9654) );
  NBUFFX2 U9616 ( .INP(CK), .Z(n9655) );
  NBUFFX2 U9617 ( .INP(CK), .Z(n9656) );
  INVX0 U9618 ( .INP(n9657), .ZN(n959) );
  INVX0 U9619 ( .INP(n9658), .ZN(n91) );
  INVX0 U9620 ( .INP(n9659), .ZN(n89) );
  NOR3X0 U9621 ( .IN1(n9660), .IN2(n9661), .IN3(n9662), .QN(n8843) );
  INVX0 U9622 ( .INP(n9663), .ZN(n869) );
  INVX0 U9623 ( .INP(n9664), .ZN(n822) );
  INVX0 U9624 ( .INP(n9665), .ZN(n765) );
  INVX0 U9625 ( .INP(n9666), .ZN(n763) );
  INVX0 U9626 ( .INP(n9667), .ZN(n759) );
  INVX0 U9627 ( .INP(n9668), .ZN(n757) );
  INVX0 U9628 ( .INP(n9669), .ZN(n74) );
  INVX0 U9629 ( .INP(n9670), .ZN(n73) );
  NAND4X0 U9630 ( .IN1(n9671), .IN2(n9672), .IN3(n9673), .IN4(n9674), .QN(
        n5961) );
  NAND2X0 U9631 ( .IN1(n9675), .IN2(g5348), .QN(n9674) );
  NAND2X0 U9632 ( .IN1(n8712), .IN2(n9676), .QN(n9673) );
  NAND2X0 U9633 ( .IN1(g31860), .IN2(g5352), .QN(n9672) );
  NAND2X0 U9634 ( .IN1(n8711), .IN2(n9677), .QN(n9671) );
  NAND4X0 U9635 ( .IN1(n9678), .IN2(n9679), .IN3(n9680), .IN4(n9681), .QN(
        n5960) );
  NAND2X0 U9636 ( .IN1(n9682), .IN2(g6732), .QN(n9681) );
  NAND2X0 U9637 ( .IN1(n8710), .IN2(n9683), .QN(n9680) );
  NAND2X0 U9638 ( .IN1(n9684), .IN2(g6736), .QN(n9679) );
  NAND2X0 U9639 ( .IN1(n8709), .IN2(n9685), .QN(n9678) );
  INVX0 U9640 ( .INP(n9686), .ZN(n540) );
  INVX0 U9641 ( .INP(n9687), .ZN(n499) );
  INVX0 U9642 ( .INP(n9688), .ZN(n497) );
  INVX0 U9643 ( .INP(n9689), .ZN(n470) );
  NOR2X0 U9644 ( .IN1(n9690), .IN2(g29279), .QN(n9689) );
  NOR2X0 U9645 ( .IN1(n8404), .IN2(n9354), .QN(n9690) );
  NAND2X0 U9646 ( .IN1(n9691), .IN2(g1677), .QN(n4459) );
  NAND2X0 U9647 ( .IN1(n9692), .IN2(g1811), .QN(n4448) );
  NAND2X0 U9648 ( .IN1(test_so53), .IN2(n9693), .QN(n4437) );
  NAND2X0 U9649 ( .IN1(n9694), .IN2(g2079), .QN(n4426) );
  NAND2X0 U9650 ( .IN1(n9695), .IN2(g2236), .QN(n4415) );
  NAND2X0 U9651 ( .IN1(n9696), .IN2(g2370), .QN(n4403) );
  NAND2X0 U9652 ( .IN1(n9697), .IN2(g2504), .QN(n4392) );
  NAND2X0 U9653 ( .IN1(n9698), .IN2(g2638), .QN(n4380) );
  NAND4X0 U9654 ( .IN1(n9699), .IN2(n9700), .IN3(n9701), .IN4(n9702), .QN(
        n4305) );
  NOR2X0 U9655 ( .IN1(n9703), .IN2(n9704), .QN(n9702) );
  NOR2X0 U9656 ( .IN1(n5656), .IN2(g4826), .QN(n9704) );
  NOR2X0 U9657 ( .IN1(n5440), .IN2(g4821), .QN(n9703) );
  NAND2X0 U9658 ( .IN1(g4646), .IN2(g29220), .QN(n9701) );
  NAND4X0 U9659 ( .IN1(n5440), .IN2(n9705), .IN3(n9706), .IN4(n8713), .QN(
        n9700) );
  NOR2X0 U9660 ( .IN1(g4688), .IN2(g4646), .QN(n9706) );
  NAND2X0 U9661 ( .IN1(n9707), .IN2(n9708), .QN(n9705) );
  NAND3X0 U9662 ( .IN1(n9709), .IN2(n9710), .IN3(n9711), .QN(n9707) );
  NAND2X0 U9663 ( .IN1(n9712), .IN2(g4776), .QN(n9711) );
  NAND2X0 U9664 ( .IN1(n5368), .IN2(n9713), .QN(n9712) );
  NAND2X0 U9665 ( .IN1(n9714), .IN2(n9715), .QN(n9713) );
  NAND2X0 U9666 ( .IN1(n9716), .IN2(n9717), .QN(n9715) );
  INVX0 U9667 ( .INP(n9718), .ZN(n9714) );
  NOR2X0 U9668 ( .IN1(n9716), .IN2(n9717), .QN(n9718) );
  NAND4X0 U9669 ( .IN1(n9719), .IN2(n9720), .IN3(n9721), .IN4(n9722), .QN(
        n9716) );
  NAND2X0 U9670 ( .IN1(n9723), .IN2(g4732), .QN(n9722) );
  NAND2X0 U9671 ( .IN1(n9724), .IN2(g4717), .QN(n9721) );
  NAND2X0 U9672 ( .IN1(n9725), .IN2(g4727), .QN(n9720) );
  NAND2X0 U9673 ( .IN1(n9726), .IN2(g4722), .QN(n9719) );
  NAND2X0 U9674 ( .IN1(n9717), .IN2(g4793), .QN(n9710) );
  NAND2X0 U9675 ( .IN1(n5368), .IN2(n9727), .QN(n9709) );
  NAND2X0 U9676 ( .IN1(n8862), .IN2(n9728), .QN(n9727) );
  NAND4X0 U9677 ( .IN1(n5707), .IN2(n9729), .IN3(n9730), .IN4(n9731), .QN(
        n9728) );
  NAND2X0 U9678 ( .IN1(n5867), .IN2(n9725), .QN(n9729) );
  NAND2X0 U9679 ( .IN1(g4831), .IN2(g4681), .QN(n9699) );
  NAND4X0 U9680 ( .IN1(n9732), .IN2(n9733), .IN3(n9734), .IN4(n9735), .QN(
        n4283) );
  NOR2X0 U9681 ( .IN1(n9736), .IN2(n9737), .QN(n9735) );
  NOR2X0 U9682 ( .IN1(n5318), .IN2(g3333), .QN(n9737) );
  NOR2X0 U9683 ( .IN1(n5283), .IN2(g4035), .QN(n9736) );
  NAND2X0 U9684 ( .IN1(g4871), .IN2(g3684), .QN(n9734) );
  NAND4X0 U9685 ( .IN1(n5283), .IN2(n9738), .IN3(n9739), .IN4(n5713), .QN(
        n9733) );
  NOR2X0 U9686 ( .IN1(g4864), .IN2(g4871), .QN(n9739) );
  NAND2X0 U9687 ( .IN1(n9740), .IN2(n9741), .QN(n9738) );
  NAND3X0 U9688 ( .IN1(n9742), .IN2(n9743), .IN3(n9744), .QN(n9740) );
  NAND2X0 U9689 ( .IN1(n9745), .IN2(g4966), .QN(n9744) );
  NAND2X0 U9690 ( .IN1(n5367), .IN2(n9746), .QN(n9745) );
  NAND2X0 U9691 ( .IN1(n9747), .IN2(n9748), .QN(n9746) );
  NAND2X0 U9692 ( .IN1(n9749), .IN2(n9750), .QN(n9748) );
  INVX0 U9693 ( .INP(n9751), .ZN(n9747) );
  NOR2X0 U9694 ( .IN1(n9749), .IN2(n9750), .QN(n9751) );
  NAND4X0 U9695 ( .IN1(n9752), .IN2(n9753), .IN3(n9754), .IN4(n9755), .QN(
        n9749) );
  NAND2X0 U9696 ( .IN1(n9756), .IN2(g4912), .QN(n9755) );
  NAND2X0 U9697 ( .IN1(n9757), .IN2(g4917), .QN(n9754) );
  NAND2X0 U9698 ( .IN1(n9758), .IN2(g4922), .QN(n9753) );
  NAND2X0 U9699 ( .IN1(n9759), .IN2(g4907), .QN(n9752) );
  NAND2X0 U9700 ( .IN1(n9750), .IN2(g4983), .QN(n9743) );
  NAND2X0 U9701 ( .IN1(n5367), .IN2(n9760), .QN(n9742) );
  NAND2X0 U9702 ( .IN1(n8863), .IN2(n9761), .QN(n9760) );
  NAND4X0 U9703 ( .IN1(n5706), .IN2(n9762), .IN3(n9763), .IN4(n9764), .QN(
        n9761) );
  NAND2X0 U9704 ( .IN1(n5879), .IN2(n9757), .QN(n9762) );
  NAND2X0 U9705 ( .IN1(g4836), .IN2(g5011), .QN(n9732) );
  INVX0 U9706 ( .INP(n9765), .ZN(n422) );
  NOR2X0 U9707 ( .IN1(n9766), .IN2(n9767), .QN(n9765) );
  NOR2X0 U9708 ( .IN1(n9358), .IN2(n8739), .QN(n9767) );
  NOR2X0 U9709 ( .IN1(n9768), .IN2(n9410), .QN(n9766) );
  NOR2X0 U9710 ( .IN1(test_so74), .IN2(test_so14), .QN(n9768) );
  INVX0 U9711 ( .INP(n9769), .ZN(n420) );
  NOR2X0 U9712 ( .IN1(n9770), .IN2(g24212), .QN(n9769) );
  NOR2X0 U9713 ( .IN1(n8828), .IN2(n9355), .QN(n9770) );
  NOR3X0 U9714 ( .IN1(g3167), .IN2(g3155), .IN3(g3161), .QN(n4034) );
  NOR3X0 U9715 ( .IN1(g3518), .IN2(g3512), .IN3(g3506), .QN(n4002) );
  NOR3X0 U9716 ( .IN1(g3863), .IN2(test_so33), .IN3(g3857), .QN(n3969) );
  NOR4X0 U9717 ( .IN1(n8776), .IN2(n1835), .IN3(n9662), .IN4(n9660), .QN(n3933) );
  INVX0 U9718 ( .INP(n9771), .ZN(n9660) );
  INVX0 U9719 ( .INP(n9772), .ZN(n9662) );
  NOR3X0 U9720 ( .IN1(g5176), .IN2(g5164), .IN3(g5170), .QN(n3926) );
  NOR3X0 U9721 ( .IN1(g5523), .IN2(g5511), .IN3(g5517), .QN(n3893) );
  NOR3X0 U9722 ( .IN1(g5863), .IN2(g5857), .IN3(g5869), .QN(n3860) );
  NOR3X0 U9723 ( .IN1(g6209), .IN2(g6203), .IN3(g6215), .QN(n3826) );
  NOR3X0 U9724 ( .IN1(g6561), .IN2(g6549), .IN3(g6555), .QN(n3792) );
  INVX0 U9725 ( .INP(n9773), .ZN(n3729) );
  NAND4X0 U9726 ( .IN1(n5520), .IN2(n5358), .IN3(n9774), .IN4(n9775), .QN(
        n3675) );
  NAND2X0 U9727 ( .IN1(n8787), .IN2(n9776), .QN(n9775) );
  NAND3X0 U9728 ( .IN1(n9777), .IN2(n9778), .IN3(n5629), .QN(n9776) );
  NAND2X0 U9729 ( .IN1(test_so72), .IN2(g174), .QN(n9778) );
  NAND2X0 U9730 ( .IN1(n5402), .IN2(n8871), .QN(n9777) );
  NAND2X0 U9731 ( .IN1(n9779), .IN2(g392), .QN(n9774) );
  NAND2X0 U9732 ( .IN1(n8467), .IN2(n9780), .QN(n9779) );
  NAND2X0 U9733 ( .IN1(n9781), .IN2(n9782), .QN(n9780) );
  INVX0 U9734 ( .INP(n9783), .ZN(n9782) );
  NOR2X0 U9735 ( .IN1(n8871), .IN2(g452), .QN(n9783) );
  NAND2X0 U9736 ( .IN1(g452), .IN2(n8871), .QN(n9781) );
  NAND3X0 U9737 ( .IN1(g2741), .IN2(n5300), .IN3(n5516), .QN(n3635) );
  INVX0 U9738 ( .INP(n9784), .ZN(n324) );
  NAND3X0 U9739 ( .IN1(n9785), .IN2(n9313), .IN3(n9786), .QN(n9784) );
  NOR2X0 U9740 ( .IN1(n9787), .IN2(n9788), .QN(n3174) );
  NOR2X0 U9741 ( .IN1(n9789), .IN2(n9790), .QN(n9788) );
  NOR2X0 U9742 ( .IN1(g72), .IN2(g482), .QN(n9790) );
  NOR2X0 U9743 ( .IN1(n5820), .IN2(n9791), .QN(n9789) );
  NOR2X0 U9744 ( .IN1(n9792), .IN2(n9793), .QN(n9787) );
  NOR2X0 U9745 ( .IN1(n5708), .IN2(n9794), .QN(n9793) );
  NOR2X0 U9746 ( .IN1(g73), .IN2(g490), .QN(n9792) );
  NOR2X0 U9747 ( .IN1(n1835), .IN2(n6010), .QN(n3084) );
  NAND3X0 U9748 ( .IN1(n9347), .IN2(g4104), .IN3(n9795), .QN(n3065) );
  NAND2X0 U9749 ( .IN1(n9796), .IN2(g4108), .QN(n9795) );
  NAND2X0 U9750 ( .IN1(n9797), .IN2(n9798), .QN(n2608) );
  NAND2X0 U9751 ( .IN1(n5323), .IN2(n9799), .QN(n9798) );
  NAND2X0 U9752 ( .IN1(n103), .IN2(g4311), .QN(n9797) );
  INVX0 U9753 ( .INP(n9800), .ZN(n199) );
  INVX0 U9754 ( .INP(n9801), .ZN(n176) );
  NAND2X0 U9755 ( .IN1(n9802), .IN2(n9803), .QN(n1733) );
  INVX0 U9756 ( .INP(g29277), .ZN(n9803) );
  NAND2X0 U9757 ( .IN1(n9431), .IN2(test_so100), .QN(n9802) );
  INVX0 U9758 ( .INP(n9804), .ZN(n1577) );
  NOR2X0 U9759 ( .IN1(n9805), .IN2(g26953), .QN(n9804) );
  NOR2X0 U9760 ( .IN1(n8462), .IN2(n9355), .QN(n9805) );
  INVX0 U9761 ( .INP(n9806), .ZN(n1460) );
  INVX0 U9762 ( .INP(n9807), .ZN(n1426) );
  INVX0 U9763 ( .INP(n9808), .ZN(n1289) );
  INVX0 U9764 ( .INP(n9809), .ZN(n1266) );
  INVX0 U9765 ( .INP(n9810), .ZN(n1179) );
  INVX0 U9766 ( .INP(n9811), .ZN(n1178) );
  INVX0 U9767 ( .INP(n9812), .ZN(n1108) );
  INVX0 U9768 ( .INP(n9813), .ZN(n1107) );
  INVX0 U9769 ( .INP(n9814), .ZN(n1038) );
  INVX0 U9770 ( .INP(n9815), .ZN(n1037) );
  NAND2X0 U9771 ( .IN1(n9816), .IN2(n9817), .QN(g34980) );
  NAND2X0 U9772 ( .IN1(test_so14), .IN2(n9423), .QN(n9817) );
  NAND2X0 U9773 ( .IN1(n9818), .IN2(n9366), .QN(n9816) );
  NAND2X0 U9774 ( .IN1(n5842), .IN2(n9819), .QN(n9818) );
  NAND4X0 U9775 ( .IN1(n26), .IN2(n9820), .IN3(n9821), .IN4(n9822), .QN(n9819)
         );
  INVX0 U9776 ( .INP(g56), .ZN(n9822) );
  INVX0 U9777 ( .INP(n9823), .ZN(n26) );
  NAND2X0 U9778 ( .IN1(n9823), .IN2(g22), .QN(g34972) );
  NAND2X0 U9779 ( .IN1(n9824), .IN2(n9825), .QN(n9823) );
  NAND2X0 U9780 ( .IN1(n9826), .IN2(n9827), .QN(n9825) );
  INVX0 U9781 ( .INP(n9828), .ZN(n9824) );
  NOR2X0 U9782 ( .IN1(n9827), .IN2(n9826), .QN(n9828) );
  NAND2X0 U9783 ( .IN1(n9829), .IN2(n9830), .QN(n9826) );
  NAND2X0 U9784 ( .IN1(g34977), .IN2(n9831), .QN(n9830) );
  NAND2X0 U9785 ( .IN1(g34978), .IN2(n9832), .QN(n9829) );
  NOR2X0 U9786 ( .IN1(n9833), .IN2(n9834), .QN(n9827) );
  NOR2X0 U9787 ( .IN1(n9835), .IN2(g34975), .QN(n9834) );
  INVX0 U9788 ( .INP(n9836), .ZN(n9833) );
  NAND2X0 U9789 ( .IN1(n9835), .IN2(g34975), .QN(n9836) );
  NAND2X0 U9790 ( .IN1(n9837), .IN2(n9838), .QN(n9835) );
  NAND2X0 U9791 ( .IN1(n9839), .IN2(n9840), .QN(n9838) );
  INVX0 U9792 ( .INP(n9841), .ZN(n9837) );
  NOR2X0 U9793 ( .IN1(n9840), .IN2(n9839), .QN(n9841) );
  NAND2X0 U9794 ( .IN1(n9842), .IN2(n9843), .QN(n9839) );
  NAND2X0 U9795 ( .IN1(n9844), .IN2(n9845), .QN(n9843) );
  INVX0 U9796 ( .INP(n9846), .ZN(n9844) );
  NAND2X0 U9797 ( .IN1(n9846), .IN2(g34971), .QN(n9842) );
  NAND2X0 U9798 ( .IN1(n9847), .IN2(n9848), .QN(n9846) );
  INVX0 U9799 ( .INP(n9849), .ZN(n9848) );
  NOR2X0 U9800 ( .IN1(n9850), .IN2(n9851), .QN(n9849) );
  NAND2X0 U9801 ( .IN1(n9850), .IN2(n9851), .QN(n9847) );
  NAND2X0 U9802 ( .IN1(n9852), .IN2(g55), .QN(n9850) );
  INVX0 U9803 ( .INP(n9853), .ZN(n9852) );
  NOR2X0 U9804 ( .IN1(n9854), .IN2(n9855), .QN(n9840) );
  NOR2X0 U9805 ( .IN1(n9856), .IN2(g34970), .QN(n9855) );
  NOR2X0 U9806 ( .IN1(n9857), .IN2(n9858), .QN(n9854) );
  INVX0 U9807 ( .INP(n9856), .ZN(n9857) );
  NAND2X0 U9808 ( .IN1(n9859), .IN2(n9860), .QN(n9856) );
  NAND2X0 U9809 ( .IN1(g34974), .IN2(n9861), .QN(n9860) );
  NAND2X0 U9810 ( .IN1(g34976), .IN2(n9862), .QN(n9859) );
  NAND2X0 U9811 ( .IN1(n9851), .IN2(g22), .QN(g34927) );
  INVX0 U9812 ( .INP(g34979), .ZN(n9851) );
  NAND4X0 U9813 ( .IN1(n9863), .IN2(n9864), .IN3(n9865), .IN4(n9866), .QN(
        g34979) );
  NOR4X0 U9814 ( .IN1(n9867), .IN2(n9868), .IN3(n9869), .IN4(n9870), .QN(n9866) );
  NOR2X0 U9815 ( .IN1(n5415), .IN2(n9871), .QN(n9870) );
  NOR2X0 U9816 ( .IN1(n5635), .IN2(n9872), .QN(n9869) );
  NOR2X0 U9817 ( .IN1(n5308), .IN2(n9873), .QN(n9868) );
  NOR2X0 U9818 ( .IN1(n9874), .IN2(DFF_420_n1), .QN(n9867) );
  NOR2X0 U9819 ( .IN1(n9875), .IN2(n9876), .QN(n9865) );
  NOR2X0 U9820 ( .IN1(n9877), .IN2(n8902), .QN(n9876) );
  NAND2X0 U9821 ( .IN1(n1465), .IN2(n9878), .QN(n9864) );
  NAND2X0 U9822 ( .IN1(n9879), .IN2(n9880), .QN(n9878) );
  NOR4X0 U9823 ( .IN1(n9881), .IN2(n9882), .IN3(n9883), .IN4(n9884), .QN(n9880) );
  INVX0 U9824 ( .INP(n9885), .ZN(n9884) );
  NAND2X0 U9826 ( .IN1(n9886), .IN2(g29221), .QN(n9885) );
  NOR2X0 U9827 ( .IN1(n5293), .IN2(n9887), .QN(n9883) );
  NOR2X0 U9828 ( .IN1(n5470), .IN2(n9888), .QN(n9882) );
  NAND3X0 U9829 ( .IN1(n9889), .IN2(n9890), .IN3(n9891), .QN(n9881) );
  NAND2X0 U9830 ( .IN1(g127), .IN2(n9892), .QN(n9891) );
  NAND2X0 U9831 ( .IN1(test_so14), .IN2(n9893), .QN(n9890) );
  INVX0 U9832 ( .INP(n9894), .ZN(n9893) );
  NAND2X0 U9833 ( .IN1(g92), .IN2(n9895), .QN(n9889) );
  NOR4X0 U9834 ( .IN1(n9896), .IN2(n9897), .IN3(n9898), .IN4(n9899), .QN(n9879) );
  NOR2X0 U9835 ( .IN1(n8732), .IN2(n9900), .QN(n9899) );
  NOR2X0 U9836 ( .IN1(n5981), .IN2(n9901), .QN(n9898) );
  NOR2X0 U9837 ( .IN1(n8739), .IN2(n9902), .QN(n9897) );
  NAND3X0 U9838 ( .IN1(n9903), .IN2(n9904), .IN3(n9905), .QN(n9896) );
  NAND2X0 U9839 ( .IN1(n9906), .IN2(g2975), .QN(n9905) );
  NAND2X0 U9840 ( .IN1(n9907), .IN2(g568), .QN(n9904) );
  NAND2X0 U9841 ( .IN1(n9908), .IN2(g604), .QN(n9903) );
  NAND2X0 U9842 ( .IN1(n9909), .IN2(g2138), .QN(n9863) );
  NAND2X0 U9843 ( .IN1(n9831), .IN2(g22), .QN(g34925) );
  INVX0 U9844 ( .INP(g34978), .ZN(n9831) );
  NAND4X0 U9845 ( .IN1(n9910), .IN2(n9911), .IN3(n9912), .IN4(n9913), .QN(
        g34978) );
  NOR4X0 U9846 ( .IN1(n9914), .IN2(n9915), .IN3(n9916), .IN4(n9917), .QN(n9913) );
  NOR2X0 U9847 ( .IN1(n9871), .IN2(g952), .QN(n9917) );
  NOR2X0 U9848 ( .IN1(n9872), .IN2(g1296), .QN(n9916) );
  NOR2X0 U9849 ( .IN1(n5347), .IN2(n9873), .QN(n9915) );
  NOR2X0 U9850 ( .IN1(n9874), .IN2(DFF_1012_n1), .QN(n9914) );
  NOR2X0 U9851 ( .IN1(n9875), .IN2(n9918), .QN(n9912) );
  NOR2X0 U9852 ( .IN1(n5484), .IN2(n9877), .QN(n9918) );
  NAND2X0 U9853 ( .IN1(n1465), .IN2(n9919), .QN(n9911) );
  NAND4X0 U9854 ( .IN1(n9920), .IN2(n9921), .IN3(n9922), .IN4(n9923), .QN(
        n9919) );
  NOR4X0 U9855 ( .IN1(n9924), .IN2(n9925), .IN3(n9926), .IN4(n9927), .QN(n9923) );
  NOR2X0 U9856 ( .IN1(n5488), .IN2(n9928), .QN(n9927) );
  NOR2X0 U9857 ( .IN1(n5342), .IN2(n9929), .QN(n9926) );
  NOR2X0 U9858 ( .IN1(n5292), .IN2(n9887), .QN(n9925) );
  NAND3X0 U9859 ( .IN1(n9930), .IN2(n9931), .IN3(n9932), .QN(n9924) );
  NAND2X0 U9860 ( .IN1(n9907), .IN2(g572), .QN(n9932) );
  NAND2X0 U9861 ( .IN1(n8745), .IN2(n9886), .QN(n9931) );
  NAND2X0 U9862 ( .IN1(test_so2), .IN2(n9933), .QN(n9930) );
  NOR3X0 U9863 ( .IN1(n9934), .IN2(n9935), .IN3(n9936), .QN(n9922) );
  NOR2X0 U9864 ( .IN1(n8813), .IN2(n9937), .QN(n9936) );
  NOR2X0 U9865 ( .IN1(n5475), .IN2(n9938), .QN(n9935) );
  NOR2X0 U9866 ( .IN1(n5494), .IN2(n9901), .QN(n9934) );
  NAND2X0 U9867 ( .IN1(test_so22), .IN2(n9939), .QN(n9921) );
  NAND2X0 U9868 ( .IN1(n9940), .IN2(g2878), .QN(n9920) );
  NAND2X0 U9869 ( .IN1(n9909), .IN2(g2130), .QN(n9910) );
  INVX0 U9870 ( .INP(n9941), .ZN(n9909) );
  NAND2X0 U9871 ( .IN1(n9832), .IN2(g22), .QN(g34923) );
  INVX0 U9872 ( .INP(g34977), .ZN(n9832) );
  NAND4X0 U9873 ( .IN1(n9942), .IN2(n9943), .IN3(n9944), .IN4(n9945), .QN(
        g34977) );
  NOR4X0 U9874 ( .IN1(n9946), .IN2(n9947), .IN3(n9948), .IN4(n9949), .QN(n9945) );
  NOR2X0 U9875 ( .IN1(n5286), .IN2(n9871), .QN(n9949) );
  NOR2X0 U9876 ( .IN1(n2549), .IN2(n9872), .QN(n9948) );
  NOR2X0 U9877 ( .IN1(g4927), .IN2(n9950), .QN(n9947) );
  NOR2X0 U9878 ( .IN1(g4737), .IN2(n9951), .QN(n9946) );
  NOR2X0 U9879 ( .IN1(n9875), .IN2(n9952), .QN(n9944) );
  NOR2X0 U9880 ( .IN1(n5639), .IN2(n9877), .QN(n9952) );
  NAND2X0 U9881 ( .IN1(n1465), .IN2(n9953), .QN(n9943) );
  NAND2X0 U9882 ( .IN1(n9954), .IN2(n9955), .QN(n9953) );
  NOR4X0 U9883 ( .IN1(n9956), .IN2(n9957), .IN3(n9958), .IN4(n9959), .QN(n9955) );
  INVX0 U9884 ( .INP(n9960), .ZN(n9959) );
  NAND2X0 U9885 ( .IN1(g37), .IN2(n9895), .QN(n9960) );
  NOR2X0 U9887 ( .IN1(n8728), .IN2(n9928), .QN(n9957) );
  NAND3X0 U9888 ( .IN1(n9961), .IN2(n9962), .IN3(n9963), .QN(n9956) );
  NAND2X0 U9889 ( .IN1(n9933), .IN2(g758), .QN(n9963) );
  NAND2X0 U9890 ( .IN1(n9964), .IN2(g794), .QN(n9962) );
  NAND2X0 U9891 ( .IN1(n9886), .IN2(g534), .QN(n9961) );
  NOR4X0 U9892 ( .IN1(n9965), .IN2(n9966), .IN3(n9967), .IN4(n9968), .QN(n9954) );
  NOR2X0 U9893 ( .IN1(n8735), .IN2(n9900), .QN(n9968) );
  NOR2X0 U9894 ( .IN1(n5493), .IN2(n9901), .QN(n9967) );
  NOR2X0 U9895 ( .IN1(n8824), .IN2(n9902), .QN(n9966) );
  NAND3X0 U9896 ( .IN1(n9969), .IN2(n9970), .IN3(n9971), .QN(n9965) );
  NAND2X0 U9897 ( .IN1(n9906), .IN2(g2955), .QN(n9971) );
  NAND2X0 U9898 ( .IN1(n9907), .IN2(g586), .QN(n9970) );
  NAND2X0 U9899 ( .IN1(n9908), .IN2(g613), .QN(n9969) );
  INVX0 U9900 ( .INP(n9938), .ZN(n9908) );
  NAND2X0 U9901 ( .IN1(n9245), .IN2(n9972), .QN(n9942) );
  NAND2X0 U9902 ( .IN1(n9861), .IN2(g22), .QN(g34921) );
  INVX0 U9903 ( .INP(g34976), .ZN(n9861) );
  NAND4X0 U9904 ( .IN1(n9973), .IN2(n9974), .IN3(n9975), .IN4(n9976), .QN(
        g34976) );
  NOR4X0 U9905 ( .IN1(n9977), .IN2(n9978), .IN3(n9979), .IN4(n9980), .QN(n9976) );
  NOR2X0 U9906 ( .IN1(n5297), .IN2(n9950), .QN(n9980) );
  NOR2X0 U9907 ( .IN1(n5345), .IN2(n9951), .QN(n9979) );
  NOR2X0 U9908 ( .IN1(n5497), .IN2(n9873), .QN(n9978) );
  NOR2X0 U9909 ( .IN1(n9874), .IN2(DFF_150_n1), .QN(n9977) );
  NOR3X0 U9910 ( .IN1(n9981), .IN2(n9875), .IN3(n9982), .QN(n9975) );
  NOR2X0 U9911 ( .IN1(n9872), .IN2(n9983), .QN(n9982) );
  NOR2X0 U9912 ( .IN1(n9871), .IN2(n9984), .QN(n9981) );
  NAND2X0 U9913 ( .IN1(n1465), .IN2(n9985), .QN(n9974) );
  NAND4X0 U9914 ( .IN1(n9986), .IN2(n9987), .IN3(n9988), .IN4(n9989), .QN(
        n9985) );
  NOR4X0 U9915 ( .IN1(n9990), .IN2(n9991), .IN3(n9958), .IN4(n9992), .QN(n9989) );
  NOR2X0 U9916 ( .IN1(n8762), .IN2(n9928), .QN(n9992) );
  NOR2X0 U9917 ( .IN1(n5479), .IN2(n9887), .QN(n9991) );
  NAND3X0 U9918 ( .IN1(n9993), .IN2(n9994), .IN3(n9995), .QN(n9990) );
  NAND2X0 U9919 ( .IN1(n9907), .IN2(g577), .QN(n9995) );
  NAND2X0 U9920 ( .IN1(test_so41), .IN2(n9886), .QN(n9994) );
  NAND2X0 U9921 ( .IN1(n9933), .IN2(g763), .QN(n9993) );
  NOR3X0 U9922 ( .IN1(n9996), .IN2(n9997), .IN3(n9998), .QN(n9988) );
  NOR2X0 U9923 ( .IN1(n8737), .IN2(n9937), .QN(n9998) );
  NOR2X0 U9924 ( .IN1(n5339), .IN2(n9938), .QN(n9997) );
  INVX0 U9925 ( .INP(n9999), .ZN(n9996) );
  NAND2X0 U9926 ( .IN1(n10000), .IN2(test_so95), .QN(n9999) );
  NAND2X0 U9928 ( .IN1(n9939), .IN2(g2936), .QN(n9987) );
  NAND2X0 U9929 ( .IN1(n9940), .IN2(g2898), .QN(n9986) );
  INVX0 U9930 ( .INP(n10001), .ZN(n9973) );
  NOR2X0 U9931 ( .IN1(n9941), .IN2(n5498), .QN(n10001) );
  NAND2X0 U9932 ( .IN1(n10002), .IN2(g22), .QN(g34919) );
  INVX0 U9933 ( .INP(g34975), .ZN(n10002) );
  NAND4X0 U9934 ( .IN1(n10003), .IN2(n10004), .IN3(n10005), .IN4(n10006), .QN(
        g34975) );
  NOR4X0 U9935 ( .IN1(n10007), .IN2(n10008), .IN3(n10009), .IN4(n10010), .QN(
        n10006) );
  NOR2X0 U9936 ( .IN1(n5295), .IN2(n9950), .QN(n10010) );
  NOR2X0 U9937 ( .IN1(n5344), .IN2(n9951), .QN(n10009) );
  NOR2X0 U9938 ( .IN1(n5495), .IN2(n9873), .QN(n10008) );
  NOR2X0 U9939 ( .IN1(n9874), .IN2(DFF_829_n1), .QN(n10007) );
  NOR3X0 U9940 ( .IN1(n10011), .IN2(n9875), .IN3(n10012), .QN(n10005) );
  NOR2X0 U9941 ( .IN1(n9872), .IN2(n10013), .QN(n10012) );
  NOR2X0 U9942 ( .IN1(n9871), .IN2(n10014), .QN(n10011) );
  NAND2X0 U9943 ( .IN1(n1465), .IN2(n10015), .QN(n10004) );
  NAND4X0 U9944 ( .IN1(n10016), .IN2(n10017), .IN3(n10018), .IN4(n10019), .QN(
        n10015) );
  NOR4X0 U9945 ( .IN1(n10020), .IN2(n10021), .IN3(n10022), .IN4(n10023), .QN(
        n10019) );
  NOR2X0 U9946 ( .IN1(n8427), .IN2(n9887), .QN(n10023) );
  NOR2X0 U9947 ( .IN1(n9928), .IN2(g2994), .QN(n10022) );
  NOR2X0 U9948 ( .IN1(n5492), .IN2(n10024), .QN(n10021) );
  NAND2X0 U9949 ( .IN1(n10025), .IN2(n10026), .QN(n10020) );
  NAND2X0 U9950 ( .IN1(n9933), .IN2(g767), .QN(n10026) );
  NAND2X0 U9951 ( .IN1(n9907), .IN2(g582), .QN(n10025) );
  NOR3X0 U9952 ( .IN1(n10027), .IN2(n10028), .IN3(n10029), .QN(n10018) );
  NOR2X0 U9954 ( .IN1(n8815), .IN2(n9937), .QN(n10029) );
  NOR2X0 U9955 ( .IN1(n5672), .IN2(n9938), .QN(n10028) );
  NOR2X0 U9956 ( .IN1(n8729), .IN2(n9901), .QN(n10027) );
  NAND2X0 U9959 ( .IN1(n9939), .IN2(g2922), .QN(n10017) );
  NAND2X0 U9960 ( .IN1(n9940), .IN2(g2864), .QN(n10016) );
  INVX0 U9961 ( .INP(n10030), .ZN(n10003) );
  NOR2X0 U9962 ( .IN1(n9941), .IN2(n5643), .QN(n10030) );
  NAND2X0 U9963 ( .IN1(n9862), .IN2(g22), .QN(g34917) );
  INVX0 U9964 ( .INP(g34974), .ZN(n9862) );
  NAND4X0 U9965 ( .IN1(n10031), .IN2(n10032), .IN3(n10033), .IN4(n10034), .QN(
        g34974) );
  NOR4X0 U9966 ( .IN1(n10035), .IN2(n10036), .IN3(n10037), .IN4(n10038), .QN(
        n10034) );
  NOR2X0 U9967 ( .IN1(n5346), .IN2(n9950), .QN(n10038) );
  NOR2X0 U9969 ( .IN1(n5296), .IN2(n9951), .QN(n10037) );
  NOR2X0 U9970 ( .IN1(n9873), .IN2(n8884), .QN(n10036) );
  NOR2X0 U9971 ( .IN1(n9874), .IN2(DFF_477_n1), .QN(n10035) );
  NOR2X0 U9973 ( .IN1(n10039), .IN2(n10040), .QN(n10033) );
  NOR2X0 U9974 ( .IN1(n10041), .IN2(n10042), .QN(n10040) );
  NOR4X0 U9975 ( .IN1(n10043), .IN2(n10044), .IN3(n10045), .IN4(n10046), .QN(
        n10041) );
  NOR2X0 U9976 ( .IN1(n5288), .IN2(n9938), .QN(n10046) );
  NOR2X0 U9977 ( .IN1(n5472), .IN2(n10047), .QN(n10045) );
  NAND3X0 U9978 ( .IN1(n10048), .IN2(n10049), .IN3(n10050), .QN(n10044) );
  NAND2X0 U9979 ( .IN1(n9933), .IN2(g772), .QN(n10050) );
  NAND2X0 U9980 ( .IN1(n9892), .IN2(g2999), .QN(n10048) );
  NAND4X0 U9981 ( .IN1(n10051), .IN2(n10052), .IN3(n10053), .IN4(n10054), .QN(
        n10043) );
  NAND2X0 U9982 ( .IN1(n9906), .IN2(g2917), .QN(n10054) );
  NAND2X0 U9983 ( .IN1(n10000), .IN2(g2852), .QN(n10053) );
  NAND2X0 U9984 ( .IN1(n9939), .IN2(g2912), .QN(n10052) );
  NAND2X0 U9985 ( .IN1(n9940), .IN2(g2856), .QN(n10051) );
  NOR2X0 U9986 ( .IN1(n9871), .IN2(n10055), .QN(n10039) );
  NAND2X0 U9987 ( .IN1(n10056), .IN2(n10057), .QN(n10032) );
  INVX0 U9988 ( .INP(n10058), .ZN(n10056) );
  INVX0 U9989 ( .INP(n10059), .ZN(n10031) );
  NOR2X0 U9990 ( .IN1(n9941), .IN2(n5499), .QN(n10059) );
  NAND2X0 U9991 ( .IN1(n9845), .IN2(g22), .QN(g34915) );
  INVX0 U9993 ( .INP(g34971), .ZN(n9845) );
  NAND4X0 U9994 ( .IN1(n10060), .IN2(n10061), .IN3(n10062), .IN4(n10063), .QN(
        g34971) );
  NOR4X0 U9995 ( .IN1(n9875), .IN2(n10064), .IN3(n10065), .IN4(n10066), .QN(
        n10063) );
  NOR2X0 U9996 ( .IN1(n5307), .IN2(n9941), .QN(n10066) );
  NOR2X0 U9997 ( .IN1(n10067), .IN2(n10042), .QN(n10065) );
  NOR4X0 U9998 ( .IN1(n10068), .IN2(n10069), .IN3(n10070), .IN4(n10071), .QN(
        n10067) );
  NOR2X0 U9999 ( .IN1(n5983), .IN2(n9901), .QN(n10071) );
  NOR2X0 U10000 ( .IN1(n5550), .IN2(n9938), .QN(n10070) );
  NAND3X0 U10001 ( .IN1(n10072), .IN2(n10073), .IN3(n10074), .QN(n10069) );
  NAND2X0 U10002 ( .IN1(n9907), .IN2(g562), .QN(n10074) );
  INVX0 U10003 ( .INP(n10047), .ZN(n9907) );
  INVX0 U10004 ( .INP(n10075), .ZN(n10073) );
  NOR2X0 U10005 ( .IN1(n10024), .IN2(n8746), .QN(n10075) );
  NAND2X0 U10006 ( .IN1(n9933), .IN2(test_so60), .QN(n10072) );
  NAND4X0 U10007 ( .IN1(n10076), .IN2(n10077), .IN3(n10078), .IN4(n10079), 
        .QN(n10068) );
  NAND2X0 U10008 ( .IN1(g100), .IN2(n9895), .QN(n10079) );
  INVX0 U10009 ( .INP(n9929), .ZN(n9895) );
  NAND3X0 U10010 ( .IN1(n10080), .IN2(g28), .IN3(n10081), .QN(n9929) );
  NOR2X0 U10011 ( .IN1(n9958), .IN2(n10082), .QN(n10078) );
  NOR2X0 U10012 ( .IN1(n5842), .IN2(n9894), .QN(n10082) );
  NAND4X0 U10013 ( .IN1(n10083), .IN2(test_so25), .IN3(n5324), .IN4(n8809), 
        .QN(n9894) );
  NOR4X0 U10014 ( .IN1(n10084), .IN2(n5324), .IN3(n8809), .IN4(test_so25), 
        .QN(n9958) );
  NAND2X0 U10015 ( .IN1(n9892), .IN2(g2890), .QN(n10077) );
  INVX0 U10016 ( .INP(n9928), .ZN(n9892) );
  NAND2X0 U10017 ( .IN1(n10081), .IN2(n10085), .QN(n9928) );
  NAND2X0 U10018 ( .IN1(n9964), .IN2(g781), .QN(n10076) );
  NOR2X0 U10019 ( .IN1(n5640), .IN2(n9877), .QN(n10064) );
  NAND2X0 U10020 ( .IN1(n10086), .IN2(n10085), .QN(n9877) );
  NOR2X0 U10021 ( .IN1(n10042), .IN2(n10087), .QN(n9875) );
  INVX0 U10022 ( .INP(n10088), .ZN(n10087) );
  NAND2X0 U10023 ( .IN1(n10049), .IN2(n10089), .QN(n10088) );
  NAND2X0 U10024 ( .IN1(n9964), .IN2(n9409), .QN(n10089) );
  INVX0 U10025 ( .INP(n9887), .ZN(n9964) );
  NAND2X0 U10026 ( .IN1(n10085), .IN2(n10090), .QN(n9887) );
  NOR2X0 U10027 ( .IN1(n10091), .IN2(n10092), .QN(n10062) );
  NOR2X0 U10028 ( .IN1(n5377), .IN2(n9873), .QN(n10092) );
  NOR2X0 U10029 ( .IN1(n9874), .IN2(DFF_206_n1), .QN(n10091) );
  NAND2X0 U10030 ( .IN1(test_so64), .IN2(n10057), .QN(n10061) );
  INVX0 U10031 ( .INP(n10093), .ZN(n10060) );
  NOR2X0 U10032 ( .IN1(n9871), .IN2(n15962), .QN(n10093) );
  NAND2X0 U10033 ( .IN1(n9858), .IN2(g22), .QN(g34913) );
  INVX0 U10034 ( .INP(g34970), .ZN(n9858) );
  NAND4X0 U10035 ( .IN1(n10094), .IN2(n10095), .IN3(n10096), .IN4(n10097), 
        .QN(g34970) );
  NOR4X0 U10036 ( .IN1(n10098), .IN2(n10099), .IN3(n10100), .IN4(n10101), .QN(
        n10097) );
  NOR2X0 U10037 ( .IN1(n5408), .IN2(n9950), .QN(n10101) );
  NAND3X0 U10038 ( .IN1(n1465), .IN2(n10085), .IN3(n2527), .QN(n9950) );
  NOR2X0 U10039 ( .IN1(n5312), .IN2(n9951), .QN(n10100) );
  NAND3X0 U10040 ( .IN1(n1465), .IN2(n10102), .IN3(n2527), .QN(n9951) );
  NOR2X0 U10041 ( .IN1(n5641), .IN2(n9873), .QN(n10099) );
  NAND3X0 U10042 ( .IN1(n10080), .IN2(n5324), .IN3(n10086), .QN(n9873) );
  NOR2X0 U10043 ( .IN1(n9874), .IN2(DFF_514_n1), .QN(n10098) );
  INVX0 U10044 ( .INP(n9972), .ZN(n9874) );
  NOR2X0 U10045 ( .IN1(g53), .IN2(n1465), .QN(n9972) );
  NOR2X0 U10046 ( .IN1(n10103), .IN2(n10104), .QN(n10096) );
  NOR2X0 U10047 ( .IN1(n10105), .IN2(n10042), .QN(n10104) );
  NOR4X0 U10048 ( .IN1(n10106), .IN2(n10107), .IN3(n10108), .IN4(n10109), .QN(
        n10105) );
  NOR2X0 U10049 ( .IN1(n15963), .IN2(n9938), .QN(n10109) );
  NOR2X0 U10050 ( .IN1(n5476), .IN2(n10047), .QN(n10108) );
  NAND3X0 U10051 ( .IN1(n10110), .IN2(n10049), .IN3(n10111), .QN(n10107) );
  NAND2X0 U10052 ( .IN1(n9933), .IN2(g776), .QN(n10111) );
  INVX0 U10053 ( .INP(n9888), .ZN(n9933) );
  NAND2X0 U10054 ( .IN1(n9487), .IN2(n10112), .QN(n10049) );
  NAND3X0 U10055 ( .IN1(n10047), .IN2(n9938), .IN3(n9888), .QN(n10112) );
  NAND3X0 U10056 ( .IN1(n10090), .IN2(g28), .IN3(n10080), .QN(n9888) );
  NAND2X0 U10057 ( .IN1(n2552), .IN2(n10102), .QN(n9938) );
  NAND3X0 U10058 ( .IN1(n2552), .IN2(n5324), .IN3(n10080), .QN(n10047) );
  NOR4X0 U10059 ( .IN1(g8), .IN2(g6), .IN3(n5469), .IN4(test_so85), .QN(n10080) );
  NAND2X0 U10060 ( .IN1(n9886), .IN2(g538), .QN(n10110) );
  INVX0 U10061 ( .INP(n10024), .ZN(n9886) );
  NAND2X0 U10062 ( .IN1(n10102), .IN2(n10090), .QN(n10024) );
  INVX0 U10063 ( .INP(n10113), .ZN(n10090) );
  NAND2X0 U10064 ( .IN1(n5468), .IN2(n10114), .QN(n10113) );
  NAND4X0 U10065 ( .IN1(n10115), .IN2(n10116), .IN3(n10117), .IN4(n10118), 
        .QN(n10106) );
  NAND2X0 U10066 ( .IN1(n9906), .IN2(g2902), .QN(n10118) );
  INVX0 U10067 ( .INP(n9937), .ZN(n9906) );
  NAND3X0 U10068 ( .IN1(n5324), .IN2(n10114), .IN3(n10083), .QN(n9937) );
  NAND2X0 U10069 ( .IN1(n10000), .IN2(g2844), .QN(n10117) );
  INVX0 U10070 ( .INP(n9901), .ZN(n10000) );
  NAND3X0 U10071 ( .IN1(n10114), .IN2(g9), .IN3(n10102), .QN(n9901) );
  NAND2X0 U10072 ( .IN1(test_so1), .IN2(n9939), .QN(n10116) );
  INVX0 U10073 ( .INP(n9900), .ZN(n9939) );
  NAND3X0 U10074 ( .IN1(n10114), .IN2(g28), .IN3(n10083), .QN(n9900) );
  INVX0 U10075 ( .INP(n10084), .ZN(n10083) );
  NAND4X0 U10076 ( .IN1(test_so85), .IN2(n3395), .IN3(g9), .IN4(g8), .QN(
        n10084) );
  NAND2X0 U10077 ( .IN1(n9940), .IN2(g2848), .QN(n10115) );
  INVX0 U10078 ( .INP(n9902), .ZN(n9940) );
  NAND3X0 U10079 ( .IN1(n10114), .IN2(g9), .IN3(n10085), .QN(n9902) );
  NOR2X0 U10080 ( .IN1(g19), .IN2(test_so25), .QN(n10114) );
  NOR2X0 U10081 ( .IN1(n9871), .IN2(n10119), .QN(n10103) );
  NAND3X0 U10082 ( .IN1(n2552), .IN2(n10085), .IN3(n1465), .QN(n9871) );
  NOR2X0 U10083 ( .IN1(n10120), .IN2(n5324), .QN(n10085) );
  NAND2X0 U10084 ( .IN1(n10121), .IN2(n10057), .QN(n10095) );
  INVX0 U10085 ( .INP(n9872), .ZN(n10057) );
  NAND3X0 U10086 ( .IN1(n1465), .IN2(n10102), .IN3(n10081), .QN(n9872) );
  INVX0 U10087 ( .INP(n10122), .ZN(n10081) );
  NAND3X0 U10088 ( .IN1(n5468), .IN2(n8809), .IN3(test_so25), .QN(n10122) );
  INVX0 U10089 ( .INP(n10042), .ZN(n1465) );
  INVX0 U10090 ( .INP(n10123), .ZN(n10121) );
  INVX0 U10091 ( .INP(n10124), .ZN(n10094) );
  NOR2X0 U10092 ( .IN1(n9941), .IN2(n5644), .QN(n10124) );
  NAND2X0 U10093 ( .IN1(n10086), .IN2(n10102), .QN(n9941) );
  NOR2X0 U10094 ( .IN1(g28), .IN2(n10120), .QN(n10102) );
  NAND4X0 U10095 ( .IN1(n8810), .IN2(n8401), .IN3(n5469), .IN4(n8893), .QN(
        n10120) );
  NOR4X0 U10096 ( .IN1(n10042), .IN2(n5468), .IN3(n8809), .IN4(test_so25), 
        .QN(n10086) );
  NAND3X0 U10097 ( .IN1(n9853), .IN2(n9820), .IN3(n10125), .QN(n10042) );
  NOR2X0 U10098 ( .IN1(test_so74), .IN2(g57), .QN(n10125) );
  INVX0 U10099 ( .INP(g53), .ZN(n9820) );
  NOR2X0 U10100 ( .IN1(n9821), .IN2(g56), .QN(n9853) );
  INVX0 U10101 ( .INP(g54), .ZN(n9821) );
  NAND2X0 U10102 ( .IN1(n10126), .IN2(n10127), .QN(g34911) );
  NAND2X0 U10103 ( .IN1(n10128), .IN2(g807), .QN(n10127) );
  NAND2X0 U10104 ( .IN1(n9365), .IN2(n10129), .QN(n10128) );
  NAND2X0 U10105 ( .IN1(n2404), .IN2(g554), .QN(n10126) );
  NAND2X0 U10106 ( .IN1(n10130), .IN2(n10131), .QN(g34882) );
  NAND2X0 U10107 ( .IN1(n9487), .IN2(g4366), .QN(n10131) );
  NAND2X0 U10108 ( .IN1(n10132), .IN2(n9368), .QN(n10130) );
  NAND3X0 U10109 ( .IN1(n10133), .IN2(n10134), .IN3(n10135), .QN(n10132) );
  NAND3X0 U10110 ( .IN1(n5653), .IN2(n10136), .IN3(n10137), .QN(n10135) );
  INVX0 U10111 ( .INP(n10138), .ZN(n10136) );
  NOR2X0 U10112 ( .IN1(n10139), .IN2(g4358), .QN(n10138) );
  NAND3X0 U10113 ( .IN1(test_so81), .IN2(g4340), .IN3(g4358), .QN(n10134) );
  NAND3X0 U10114 ( .IN1(n10139), .IN2(n8867), .IN3(n5348), .QN(n10133) );
  NAND4X0 U10115 ( .IN1(n5653), .IN2(n8867), .IN3(n10140), .IN4(n10141), .QN(
        n10139) );
  NAND2X0 U10116 ( .IN1(n5540), .IN2(n10142), .QN(n10141) );
  NAND3X0 U10117 ( .IN1(n10143), .IN2(n10144), .IN3(n10145), .QN(n10142) );
  NAND2X0 U10118 ( .IN1(n8714), .IN2(g4322), .QN(n10144) );
  NAND3X0 U10119 ( .IN1(g90), .IN2(n5634), .IN3(n5506), .QN(n10143) );
  NAND3X0 U10120 ( .IN1(n5506), .IN2(g4311), .IN3(g4332), .QN(n10140) );
  NAND3X0 U10121 ( .IN1(n10146), .IN2(n10147), .IN3(n10148), .QN(g34881) );
  NAND2X0 U10122 ( .IN1(n9487), .IN2(g794), .QN(n10148) );
  NAND3X0 U10123 ( .IN1(n2404), .IN2(n10129), .IN3(g807), .QN(n10147) );
  INVX0 U10124 ( .INP(n2405), .ZN(n10129) );
  NAND2X0 U10125 ( .IN1(n2405), .IN2(n5479), .QN(n10146) );
  NAND3X0 U10126 ( .IN1(n10149), .IN2(n10150), .IN3(n10151), .QN(g34880) );
  NAND2X0 U10127 ( .IN1(n9487), .IN2(g626), .QN(n10151) );
  NAND3X0 U10128 ( .IN1(n2421), .IN2(n10152), .IN3(n9340), .QN(n10150) );
  INVX0 U10129 ( .INP(n2422), .ZN(n10152) );
  NAND2X0 U10130 ( .IN1(n2422), .IN2(n15963), .QN(n10149) );
  NAND3X0 U10131 ( .IN1(n10153), .IN2(n10154), .IN3(n10155), .QN(g34850) );
  NAND2X0 U10132 ( .IN1(n9487), .IN2(g790), .QN(n10155) );
  NAND3X0 U10133 ( .IN1(n2404), .IN2(n10156), .IN3(g794), .QN(n10154) );
  INVX0 U10134 ( .INP(n2419), .ZN(n10156) );
  NAND2X0 U10135 ( .IN1(n2419), .IN2(n5291), .QN(n10153) );
  NAND3X0 U10136 ( .IN1(n10157), .IN2(n10158), .IN3(n10159), .QN(g34849) );
  NAND2X0 U10137 ( .IN1(n9487), .IN2(g622), .QN(n10159) );
  NAND3X0 U10138 ( .IN1(n2421), .IN2(n10160), .IN3(g626), .QN(n10158) );
  INVX0 U10139 ( .INP(n2423), .ZN(n10160) );
  NAND2X0 U10140 ( .IN1(n2423), .IN2(n5288), .QN(n10157) );
  NOR2X0 U10141 ( .IN1(n8591), .IN2(n10161), .QN(g34839) );
  NOR3X0 U10142 ( .IN1(g4366), .IN2(n10162), .IN3(n10163), .QN(n10161) );
  NOR2X0 U10143 ( .IN1(n10164), .IN2(g4332), .QN(n10163) );
  NOR3X0 U10144 ( .IN1(g4311), .IN2(g73), .IN3(n10165), .QN(n10164) );
  NOR2X0 U10145 ( .IN1(n5540), .IN2(n10166), .QN(n10162) );
  NOR3X0 U10146 ( .IN1(n10167), .IN2(n10165), .IN3(g4311), .QN(n10166) );
  INVX0 U10147 ( .INP(n10168), .ZN(n10165) );
  NAND2X0 U10148 ( .IN1(n10169), .IN2(n10170), .QN(g34808) );
  NAND2X0 U10149 ( .IN1(n9487), .IN2(g2955), .QN(n10170) );
  NAND2X0 U10150 ( .IN1(n10171), .IN2(n9369), .QN(n10169) );
  NAND3X0 U10151 ( .IN1(g91), .IN2(n10172), .IN3(n8813), .QN(n10171) );
  NAND2X0 U10152 ( .IN1(n10173), .IN2(n10174), .QN(g34807) );
  INVX0 U10153 ( .INP(n10175), .ZN(n10174) );
  NOR2X0 U10154 ( .IN1(n9360), .IN2(n8737), .QN(n10175) );
  NAND2X0 U10155 ( .IN1(n10176), .IN2(n9369), .QN(n10173) );
  NAND4X0 U10156 ( .IN1(n10177), .IN2(n10178), .IN3(n10179), .IN4(n10180), 
        .QN(n10176) );
  NOR4X0 U10157 ( .IN1(n10181), .IN2(n10182), .IN3(g2955), .IN4(g2946), .QN(
        n10180) );
  NOR2X0 U10158 ( .IN1(n10183), .IN2(n10184), .QN(n10179) );
  NAND2X0 U10159 ( .IN1(n10185), .IN2(n10186), .QN(g34806) );
  NAND2X0 U10160 ( .IN1(n9486), .IN2(g2927), .QN(n10186) );
  NAND2X0 U10161 ( .IN1(n10187), .IN2(n9369), .QN(n10185) );
  NAND3X0 U10162 ( .IN1(n8819), .IN2(n8737), .IN3(n8820), .QN(n10187) );
  NOR2X0 U10163 ( .IN1(n9420), .IN2(n10188), .QN(g34805) );
  NOR2X0 U10164 ( .IN1(g2999), .IN2(g2932), .QN(n10188) );
  NAND2X0 U10165 ( .IN1(n10189), .IN2(n10190), .QN(g34804) );
  NAND2X0 U10166 ( .IN1(n9486), .IN2(g2965), .QN(n10190) );
  NAND2X0 U10167 ( .IN1(n10191), .IN2(n9369), .QN(n10189) );
  NAND3X0 U10168 ( .IN1(g962), .IN2(g1306), .IN3(n5750), .QN(n10191) );
  NAND2X0 U10169 ( .IN1(n10192), .IN2(n10193), .QN(g34803) );
  NAND2X0 U10170 ( .IN1(n9486), .IN2(g2917), .QN(n10193) );
  NAND2X0 U10171 ( .IN1(n10194), .IN2(n9369), .QN(n10192) );
  NAND3X0 U10172 ( .IN1(g44), .IN2(n8814), .IN3(n8815), .QN(n10194) );
  NAND2X0 U10173 ( .IN1(n10195), .IN2(n10196), .QN(g34802) );
  NAND2X0 U10174 ( .IN1(n9486), .IN2(g2902), .QN(n10196) );
  NAND2X0 U10175 ( .IN1(n10197), .IN2(n9369), .QN(n10195) );
  NAND3X0 U10176 ( .IN1(n10198), .IN2(n10199), .IN3(n8825), .QN(n10197) );
  NAND2X0 U10177 ( .IN1(n10200), .IN2(n10201), .QN(g34801) );
  NAND2X0 U10178 ( .IN1(n9486), .IN2(g2970), .QN(n10201) );
  NAND2X0 U10179 ( .IN1(n10202), .IN2(n9370), .QN(n10200) );
  NAND4X0 U10180 ( .IN1(n8823), .IN2(n8822), .IN3(n5595), .IN4(g691), .QN(
        n10202) );
  NAND2X0 U10181 ( .IN1(n10203), .IN2(n10204), .QN(g34799) );
  NAND2X0 U10182 ( .IN1(n9486), .IN2(g2873), .QN(n10204) );
  NAND2X0 U10183 ( .IN1(n10205), .IN2(n9370), .QN(n10203) );
  NAND2X0 U10184 ( .IN1(n8742), .IN2(g44), .QN(n10205) );
  NAND2X0 U10185 ( .IN1(n10206), .IN2(n10207), .QN(g34798) );
  NAND2X0 U10186 ( .IN1(n9486), .IN2(g2878), .QN(n10207) );
  NAND2X0 U10187 ( .IN1(n10208), .IN2(n9370), .QN(n10206) );
  NAND2X0 U10188 ( .IN1(n8739), .IN2(n8818), .QN(n10208) );
  NAND2X0 U10189 ( .IN1(n10209), .IN2(n10210), .QN(g34797) );
  INVX0 U10190 ( .INP(n10211), .ZN(n10210) );
  NOR2X0 U10191 ( .IN1(n9360), .IN2(n8824), .QN(n10211) );
  NAND2X0 U10192 ( .IN1(n10212), .IN2(n9370), .QN(n10209) );
  NAND2X0 U10193 ( .IN1(n8738), .IN2(g91), .QN(n10212) );
  NAND2X0 U10194 ( .IN1(n10213), .IN2(n10214), .QN(g34796) );
  NAND2X0 U10195 ( .IN1(n9485), .IN2(g2898), .QN(n10214) );
  NAND2X0 U10196 ( .IN1(n10215), .IN2(n9370), .QN(n10213) );
  NAND2X0 U10197 ( .IN1(n8824), .IN2(n10172), .QN(n10215) );
  NOR2X0 U10198 ( .IN1(n10216), .IN2(n10217), .QN(n10172) );
  NAND2X0 U10199 ( .IN1(n10218), .IN2(n10219), .QN(g34795) );
  NAND2X0 U10200 ( .IN1(n9485), .IN2(g2864), .QN(n10219) );
  NAND2X0 U10201 ( .IN1(n10220), .IN2(n9370), .QN(n10218) );
  NAND2X0 U10202 ( .IN1(n8740), .IN2(n10221), .QN(n10220) );
  INVX0 U10203 ( .INP(n10183), .ZN(n10221) );
  NAND4X0 U10204 ( .IN1(n5882), .IN2(n5861), .IN3(n10222), .IN4(n10223), .QN(
        n10183) );
  NAND2X0 U10205 ( .IN1(n10224), .IN2(n10225), .QN(g34794) );
  NAND2X0 U10206 ( .IN1(n9485), .IN2(g2856), .QN(n10225) );
  NAND2X0 U10207 ( .IN1(n10226), .IN2(n9370), .QN(n10224) );
  NAND2X0 U10208 ( .IN1(n5489), .IN2(n10227), .QN(n10226) );
  INVX0 U10209 ( .INP(n10184), .ZN(n10227) );
  NAND3X0 U10210 ( .IN1(n10228), .IN2(n10229), .IN3(n10230), .QN(n10184) );
  NAND2X0 U10211 ( .IN1(n10231), .IN2(n10232), .QN(g34793) );
  NAND2X0 U10212 ( .IN1(n9485), .IN2(g2848), .QN(n10232) );
  NAND2X0 U10213 ( .IN1(n10233), .IN2(n9370), .QN(n10231) );
  NAND3X0 U10214 ( .IN1(n10234), .IN2(n10177), .IN3(n8826), .QN(n10233) );
  NAND2X0 U10215 ( .IN1(n10235), .IN2(n10236), .QN(g34792) );
  NAND2X0 U10216 ( .IN1(n9485), .IN2(g29214), .QN(n10236) );
  NAND2X0 U10217 ( .IN1(n10237), .IN2(n9370), .QN(n10235) );
  NAND3X0 U10218 ( .IN1(n10238), .IN2(n10178), .IN3(n8821), .QN(n10237) );
  NAND3X0 U10219 ( .IN1(n10239), .IN2(n10240), .IN3(n10241), .QN(g34791) );
  NAND2X0 U10220 ( .IN1(n9485), .IN2(g785), .QN(n10241) );
  NAND3X0 U10221 ( .IN1(n2404), .IN2(n10242), .IN3(g790), .QN(n10240) );
  INVX0 U10222 ( .INP(n2425), .ZN(n10242) );
  NAND2X0 U10223 ( .IN1(n2425), .IN2(n5292), .QN(n10239) );
  NAND3X0 U10224 ( .IN1(n10243), .IN2(n10244), .IN3(n10245), .QN(g34790) );
  NAND2X0 U10225 ( .IN1(n9485), .IN2(g617), .QN(n10245) );
  NAND3X0 U10226 ( .IN1(n2421), .IN2(n10246), .IN3(g622), .QN(n10244) );
  INVX0 U10227 ( .INP(n2427), .ZN(n10246) );
  NAND2X0 U10228 ( .IN1(n2427), .IN2(n5672), .QN(n10243) );
  INVX0 U10229 ( .INP(n10247), .ZN(g34788) );
  NAND2X0 U10230 ( .IN1(g890), .IN2(n10248), .QN(n10247) );
  NAND2X0 U10231 ( .IN1(g479), .IN2(n3195), .QN(n10248) );
  NAND2X0 U10232 ( .IN1(n10249), .IN2(n10250), .QN(g34783) );
  NAND3X0 U10233 ( .IN1(n10251), .IN2(n10252), .IN3(n10253), .QN(n10250) );
  NAND3X0 U10234 ( .IN1(n10254), .IN2(n10255), .IN3(n10256), .QN(n10249) );
  NAND2X0 U10235 ( .IN1(n10257), .IN2(n10258), .QN(g34735) );
  INVX0 U10236 ( .INP(n10259), .ZN(n10258) );
  NOR2X0 U10237 ( .IN1(n9359), .IN2(n8372), .QN(n10259) );
  NAND2X0 U10238 ( .IN1(n10260), .IN2(n9370), .QN(n10257) );
  NAND2X0 U10239 ( .IN1(n5639), .IN2(n8741), .QN(n10260) );
  NAND2X0 U10240 ( .IN1(n10261), .IN2(n10262), .QN(g34734) );
  NAND2X0 U10241 ( .IN1(n9484), .IN2(g4172), .QN(n10262) );
  NAND2X0 U10242 ( .IN1(n10263), .IN2(n9371), .QN(n10261) );
  NAND2X0 U10243 ( .IN1(n5494), .IN2(n8820), .QN(n10263) );
  NOR2X0 U10244 ( .IN1(n9419), .IN2(n10264), .QN(g34733) );
  NOR2X0 U10245 ( .IN1(g4153), .IN2(g4172), .QN(n10264) );
  NAND2X0 U10246 ( .IN1(n10265), .IN2(n10266), .QN(g34732) );
  NAND2X0 U10247 ( .IN1(n9366), .IN2(g2994), .QN(n10266) );
  NAND2X0 U10248 ( .IN1(n9484), .IN2(g2999), .QN(n10265) );
  INVX0 U10249 ( .INP(n10267), .ZN(g34731) );
  NOR2X0 U10250 ( .IN1(n10268), .IN2(n10269), .QN(n10267) );
  NOR2X0 U10251 ( .IN1(n9358), .IN2(n5635), .QN(n10269) );
  NOR2X0 U10252 ( .IN1(n10270), .IN2(n9397), .QN(n10268) );
  NOR2X0 U10253 ( .IN1(n10271), .IN2(test_so64), .QN(n10270) );
  NAND2X0 U10254 ( .IN1(n10272), .IN2(n10273), .QN(g34730) );
  NAND2X0 U10255 ( .IN1(n9484), .IN2(g1296), .QN(n10273) );
  NAND2X0 U10256 ( .IN1(n10274), .IN2(n9371), .QN(n10272) );
  NAND2X0 U10257 ( .IN1(n8744), .IN2(n5635), .QN(n10274) );
  NAND3X0 U10258 ( .IN1(n10275), .IN2(n10276), .IN3(n10277), .QN(g34729) );
  INVX0 U10259 ( .INP(n2499), .ZN(n10277) );
  NAND2X0 U10260 ( .IN1(n5796), .IN2(n9371), .QN(n10276) );
  NAND2X0 U10261 ( .IN1(n9484), .IN2(g1291), .QN(n10275) );
  NAND2X0 U10262 ( .IN1(n10278), .IN2(n10279), .QN(g34728) );
  INVX0 U10263 ( .INP(n10280), .ZN(n10279) );
  NOR2X0 U10264 ( .IN1(n9358), .IN2(n5415), .QN(n10280) );
  NAND2X0 U10265 ( .IN1(n10281), .IN2(n9371), .QN(n10278) );
  NAND2X0 U10266 ( .IN1(n15962), .IN2(n10198), .QN(n10281) );
  NAND2X0 U10267 ( .IN1(n10282), .IN2(n10283), .QN(g34727) );
  NAND2X0 U10268 ( .IN1(n9484), .IN2(g952), .QN(n10283) );
  NAND2X0 U10269 ( .IN1(n10284), .IN2(n9371), .QN(n10282) );
  NAND2X0 U10270 ( .IN1(n5415), .IN2(n8748), .QN(n10284) );
  NAND3X0 U10271 ( .IN1(n10285), .IN2(n10286), .IN3(n10287), .QN(g34726) );
  INVX0 U10272 ( .INP(n2505), .ZN(n10287) );
  NAND2X0 U10273 ( .IN1(n5630), .IN2(n9371), .QN(n10286) );
  INVX0 U10274 ( .INP(n10288), .ZN(n10285) );
  NOR2X0 U10275 ( .IN1(n9356), .IN2(n5286), .QN(n10288) );
  NAND3X0 U10276 ( .IN1(n10289), .IN2(n10290), .IN3(n10291), .QN(g34725) );
  NAND2X0 U10277 ( .IN1(n9484), .IN2(g781), .QN(n10291) );
  NAND3X0 U10278 ( .IN1(n2404), .IN2(n10292), .IN3(g785), .QN(n10290) );
  INVX0 U10279 ( .INP(n2485), .ZN(n10292) );
  NAND2X0 U10280 ( .IN1(n2485), .IN2(n5293), .QN(n10289) );
  NAND3X0 U10281 ( .IN1(n10293), .IN2(n10294), .IN3(n10295), .QN(g34724) );
  NAND2X0 U10282 ( .IN1(n9484), .IN2(g613), .QN(n10295) );
  NAND3X0 U10283 ( .IN1(n2421), .IN2(n10296), .IN3(g617), .QN(n10294) );
  INVX0 U10284 ( .INP(n2487), .ZN(n10296) );
  NAND2X0 U10285 ( .IN1(n2487), .IN2(n5339), .QN(n10293) );
  NAND2X0 U10286 ( .IN1(n10297), .IN2(n10298), .QN(g34723) );
  NAND2X0 U10287 ( .IN1(test_so41), .IN2(n9513), .QN(n10298) );
  NAND2X0 U10288 ( .IN1(n10299), .IN2(n9371), .QN(n10297) );
  NAND2X0 U10289 ( .IN1(n5490), .IN2(n8822), .QN(n10299) );
  NAND2X0 U10290 ( .IN1(n10300), .IN2(n10301), .QN(g34722) );
  NAND2X0 U10291 ( .IN1(n9483), .IN2(g538), .QN(n10301) );
  NAND2X0 U10292 ( .IN1(n10302), .IN2(n9371), .QN(n10300) );
  NAND2X0 U10293 ( .IN1(n5492), .IN2(g691), .QN(n10302) );
  NAND2X0 U10294 ( .IN1(n10303), .IN2(n10304), .QN(g34721) );
  NAND2X0 U10295 ( .IN1(g29221), .IN2(n9513), .QN(n10304) );
  NAND2X0 U10296 ( .IN1(n10305), .IN2(n9371), .QN(n10303) );
  NAND2X0 U10297 ( .IN1(n8747), .IN2(n8746), .QN(n10305) );
  NAND2X0 U10298 ( .IN1(n10306), .IN2(n10307), .QN(g34720) );
  NAND2X0 U10299 ( .IN1(n9483), .IN2(g534), .QN(n10307) );
  NAND2X0 U10300 ( .IN1(n10308), .IN2(n9372), .QN(n10306) );
  NAND2X0 U10301 ( .IN1(n8745), .IN2(g29212), .QN(n10308) );
  NOR2X0 U10302 ( .IN1(n9414), .IN2(n10309), .QN(g34719) );
  NOR2X0 U10303 ( .IN1(g209), .IN2(g538), .QN(n10309) );
  NOR2X0 U10304 ( .IN1(n5497), .IN2(n9395), .QN(g34647) );
  NOR2X0 U10305 ( .IN1(n5644), .IN2(n9398), .QN(g34646) );
  NOR2X0 U10306 ( .IN1(n5499), .IN2(n9395), .QN(g34645) );
  NOR2X0 U10307 ( .IN1(n5643), .IN2(n9397), .QN(g34644) );
  NOR2X0 U10308 ( .IN1(n5498), .IN2(n9399), .QN(g34643) );
  NAND2X0 U10309 ( .IN1(n10310), .IN2(n10311), .QN(g34642) );
  NAND2X0 U10310 ( .IN1(n9364), .IN2(g4927), .QN(n10311) );
  NAND2X0 U10311 ( .IN1(n9483), .IN2(g4912), .QN(n10310) );
  NAND2X0 U10312 ( .IN1(n10312), .IN2(n10313), .QN(g34641) );
  NAND2X0 U10313 ( .IN1(n9364), .IN2(g4912), .QN(n10313) );
  NAND2X0 U10315 ( .IN1(n9483), .IN2(g4907), .QN(n10312) );
  NAND2X0 U10316 ( .IN1(n10314), .IN2(n10315), .QN(g34640) );
  NAND2X0 U10317 ( .IN1(n9364), .IN2(g4907), .QN(n10315) );
  NAND2X0 U10319 ( .IN1(n9483), .IN2(g4922), .QN(n10314) );
  NAND2X0 U10320 ( .IN1(n10316), .IN2(n10317), .QN(g34639) );
  NAND2X0 U10321 ( .IN1(n9364), .IN2(g4922), .QN(n10317) );
  NAND2X0 U10322 ( .IN1(n9483), .IN2(g4917), .QN(n10316) );
  NOR2X0 U10323 ( .IN1(n5408), .IN2(n9387), .QN(g34638) );
  NAND2X0 U10324 ( .IN1(n10318), .IN2(n10319), .QN(g34637) );
  NAND2X0 U10325 ( .IN1(n9364), .IN2(g4737), .QN(n10319) );
  NAND2X0 U10326 ( .IN1(n9483), .IN2(g4722), .QN(n10318) );
  NAND2X0 U10327 ( .IN1(n10320), .IN2(n10321), .QN(g34636) );
  NAND2X0 U10328 ( .IN1(n9364), .IN2(g4722), .QN(n10321) );
  NAND2X0 U10329 ( .IN1(n9482), .IN2(g4717), .QN(n10320) );
  NAND2X0 U10330 ( .IN1(n10322), .IN2(n10323), .QN(g34635) );
  NAND2X0 U10331 ( .IN1(n9364), .IN2(g4717), .QN(n10323) );
  NAND2X0 U10332 ( .IN1(n9482), .IN2(g4732), .QN(n10322) );
  NAND2X0 U10333 ( .IN1(n10324), .IN2(n10325), .QN(g34634) );
  NAND2X0 U10334 ( .IN1(n9363), .IN2(g4732), .QN(n10325) );
  NAND2X0 U10335 ( .IN1(n9482), .IN2(g4727), .QN(n10324) );
  NOR2X0 U10336 ( .IN1(n5312), .IN2(n9394), .QN(g34633) );
  NAND2X0 U10337 ( .IN1(n10326), .IN2(n10327), .QN(g34632) );
  NAND2X0 U10338 ( .IN1(n9363), .IN2(g4245), .QN(n10327) );
  NAND2X0 U10339 ( .IN1(test_so67), .IN2(n9512), .QN(n10326) );
  NAND2X0 U10340 ( .IN1(n10328), .IN2(n10329), .QN(g34631) );
  NAND2X0 U10341 ( .IN1(test_so67), .IN2(n9371), .QN(n10329) );
  NAND2X0 U10342 ( .IN1(n9482), .IN2(g4253), .QN(n10328) );
  NAND2X0 U10343 ( .IN1(n10330), .IN2(n10331), .QN(g34630) );
  NAND2X0 U10344 ( .IN1(n9363), .IN2(g4253), .QN(n10331) );
  INVX0 U10345 ( .INP(n10332), .ZN(n10330) );
  NOR2X0 U10346 ( .IN1(n9359), .IN2(n5639), .QN(n10332) );
  NAND2X0 U10347 ( .IN1(n10333), .IN2(n10334), .QN(g34629) );
  NAND2X0 U10348 ( .IN1(n9362), .IN2(g4157), .QN(n10334) );
  NAND2X0 U10349 ( .IN1(n9482), .IN2(g4146), .QN(n10333) );
  NAND2X0 U10350 ( .IN1(n10335), .IN2(n10336), .QN(g34628) );
  NAND2X0 U10351 ( .IN1(n9362), .IN2(g4146), .QN(n10336) );
  INVX0 U10352 ( .INP(n10337), .ZN(n10335) );
  NOR2X0 U10353 ( .IN1(n9360), .IN2(n5494), .QN(n10337) );
  NOR2X0 U10354 ( .IN1(n5641), .IN2(n9394), .QN(g34627) );
  NOR2X0 U10355 ( .IN1(n9413), .IN2(n8884), .QN(g34626) );
  NOR2X0 U10356 ( .IN1(n5495), .IN2(n9393), .QN(g34625) );
  NAND2X0 U10357 ( .IN1(n10338), .IN2(n10339), .QN(g34624) );
  NAND2X0 U10358 ( .IN1(n9362), .IN2(g2988), .QN(n10339) );
  NAND2X0 U10359 ( .IN1(n9482), .IN2(g2994), .QN(n10338) );
  NAND2X0 U10360 ( .IN1(n10340), .IN2(n10341), .QN(g34623) );
  NAND2X0 U10361 ( .IN1(n9362), .IN2(g2970), .QN(n10341) );
  NAND2X0 U10362 ( .IN1(test_so22), .IN2(n9511), .QN(n10340) );
  NAND2X0 U10363 ( .IN1(n10342), .IN2(n10343), .QN(g34622) );
  NAND2X0 U10364 ( .IN1(test_so22), .IN2(n9369), .QN(n10343) );
  NAND2X0 U10365 ( .IN1(n9482), .IN2(g2950), .QN(n10342) );
  NAND2X0 U10366 ( .IN1(n10344), .IN2(n10345), .QN(g34621) );
  NAND2X0 U10367 ( .IN1(n9363), .IN2(g2950), .QN(n10345) );
  NAND2X0 U10368 ( .IN1(n9481), .IN2(g2936), .QN(n10344) );
  NAND2X0 U10369 ( .IN1(n10346), .IN2(n10347), .QN(g34620) );
  NAND2X0 U10370 ( .IN1(n9362), .IN2(g2936), .QN(n10347) );
  NAND2X0 U10371 ( .IN1(n9481), .IN2(g2922), .QN(n10346) );
  NAND2X0 U10372 ( .IN1(n10348), .IN2(n10349), .QN(g34619) );
  NAND2X0 U10373 ( .IN1(n9362), .IN2(g2922), .QN(n10349) );
  NAND2X0 U10374 ( .IN1(n9481), .IN2(g2912), .QN(n10348) );
  NAND2X0 U10375 ( .IN1(n10350), .IN2(n10351), .QN(g34618) );
  NAND2X0 U10376 ( .IN1(n9363), .IN2(g2912), .QN(n10351) );
  NAND2X0 U10377 ( .IN1(test_so1), .IN2(n9513), .QN(n10350) );
  NAND2X0 U10378 ( .IN1(n10352), .IN2(n10353), .QN(g34617) );
  NAND2X0 U10379 ( .IN1(test_so1), .IN2(n9369), .QN(n10353) );
  INVX0 U10380 ( .INP(n10354), .ZN(n10352) );
  NOR2X0 U10381 ( .IN1(n9358), .IN2(n5842), .QN(n10354) );
  NAND2X0 U10382 ( .IN1(n10355), .IN2(n10356), .QN(g34616) );
  NAND2X0 U10383 ( .IN1(n9363), .IN2(g2868), .QN(n10356) );
  NAND2X0 U10384 ( .IN1(n9481), .IN2(g2988), .QN(n10355) );
  NAND2X0 U10385 ( .IN1(n10357), .IN2(n10358), .QN(g34615) );
  NAND2X0 U10386 ( .IN1(n9363), .IN2(g2873), .QN(n10358) );
  NAND2X0 U10387 ( .IN1(n9481), .IN2(g2868), .QN(n10357) );
  NAND2X0 U10388 ( .IN1(n10359), .IN2(n10360), .QN(g34614) );
  NAND2X0 U10389 ( .IN1(n9363), .IN2(g29214), .QN(n10360) );
  NAND2X0 U10390 ( .IN1(g37), .IN2(n9427), .QN(n10359) );
  NAND2X0 U10391 ( .IN1(n10361), .IN2(n10362), .QN(g34613) );
  NAND2X0 U10392 ( .IN1(test_so95), .IN2(n9426), .QN(n10362) );
  NAND2X0 U10393 ( .IN1(g37), .IN2(n9368), .QN(n10361) );
  NAND2X0 U10394 ( .IN1(n10363), .IN2(n10364), .QN(g34612) );
  NAND2X0 U10395 ( .IN1(test_so95), .IN2(n9366), .QN(n10364) );
  NAND2X0 U10396 ( .IN1(n9481), .IN2(g2860), .QN(n10363) );
  NAND2X0 U10397 ( .IN1(n10365), .IN2(n10366), .QN(g34611) );
  NAND2X0 U10398 ( .IN1(n9364), .IN2(g2860), .QN(n10366) );
  NAND2X0 U10399 ( .IN1(n9481), .IN2(g2852), .QN(n10365) );
  NAND2X0 U10400 ( .IN1(n10367), .IN2(n10368), .QN(g34610) );
  NAND2X0 U10401 ( .IN1(n9364), .IN2(g2852), .QN(n10368) );
  NAND2X0 U10402 ( .IN1(n9480), .IN2(g2844), .QN(n10367) );
  NAND2X0 U10403 ( .IN1(n10369), .IN2(n10370), .QN(g34609) );
  NAND2X0 U10404 ( .IN1(n9364), .IN2(g2844), .QN(n10370) );
  NAND2X0 U10405 ( .IN1(n9480), .IN2(g2890), .QN(n10369) );
  NAND2X0 U10406 ( .IN1(n10371), .IN2(n10372), .QN(g34608) );
  NAND2X0 U10407 ( .IN1(n9364), .IN2(g2704), .QN(n10372) );
  NAND2X0 U10408 ( .IN1(n9480), .IN2(g2697), .QN(n10371) );
  NAND2X0 U10409 ( .IN1(n10373), .IN2(n10374), .QN(g34607) );
  NAND2X0 U10410 ( .IN1(n9364), .IN2(g2697), .QN(n10374) );
  NAND2X0 U10411 ( .IN1(n9480), .IN2(g2689), .QN(n10373) );
  NOR2X0 U10412 ( .IN1(n5347), .IN2(n9393), .QN(g34606) );
  NAND2X0 U10413 ( .IN1(n10375), .IN2(n10376), .QN(g34605) );
  NAND2X0 U10414 ( .IN1(n9364), .IN2(g2145), .QN(n10376) );
  NAND2X0 U10415 ( .IN1(n9480), .IN2(g2138), .QN(n10375) );
  NAND2X0 U10416 ( .IN1(n10377), .IN2(n10378), .QN(g34604) );
  NAND2X0 U10417 ( .IN1(n9364), .IN2(g2138), .QN(n10378) );
  NAND2X0 U10418 ( .IN1(n9480), .IN2(g2130), .QN(n10377) );
  NOR2X0 U10419 ( .IN1(n5487), .IN2(n9392), .QN(g34603) );
  NOR2X0 U10420 ( .IN1(n2549), .IN2(n9391), .QN(g34602) );
  NOR2X0 U10421 ( .IN1(n5286), .IN2(n9391), .QN(g34601) );
  NAND3X0 U10422 ( .IN1(n10379), .IN2(n10380), .IN3(n10381), .QN(g34600) );
  NAND2X0 U10423 ( .IN1(n9480), .IN2(g776), .QN(n10381) );
  NAND3X0 U10424 ( .IN1(n2404), .IN2(n10382), .IN3(g781), .QN(n10380) );
  INVX0 U10425 ( .INP(n2507), .ZN(n10382) );
  NAND2X0 U10426 ( .IN1(n2507), .IN2(n5551), .QN(n10379) );
  NAND3X0 U10427 ( .IN1(n10383), .IN2(n10384), .IN3(n10385), .QN(g34599) );
  NAND2X0 U10428 ( .IN1(n9479), .IN2(g608), .QN(n10385) );
  NAND3X0 U10429 ( .IN1(n2421), .IN2(n10386), .IN3(g613), .QN(n10384) );
  INVX0 U10430 ( .INP(n2509), .ZN(n10386) );
  NAND2X0 U10431 ( .IN1(n2509), .IN2(n5474), .QN(n10383) );
  NAND2X0 U10432 ( .IN1(n10387), .IN2(n10388), .QN(g34598) );
  INVX0 U10433 ( .INP(n10389), .ZN(n10388) );
  NOR2X0 U10434 ( .IN1(n9358), .IN2(n8745), .QN(n10389) );
  NAND2X0 U10435 ( .IN1(g29221), .IN2(n9382), .QN(n10387) );
  NAND2X0 U10436 ( .IN1(n10390), .IN2(n10391), .QN(g34468) );
  NAND2X0 U10437 ( .IN1(n10392), .IN2(g4854), .QN(n10391) );
  NAND2X0 U10438 ( .IN1(n10393), .IN2(n9382), .QN(n10392) );
  NAND2X0 U10439 ( .IN1(n10394), .IN2(n10395), .QN(n10393) );
  INVX0 U10440 ( .INP(n10396), .ZN(n10390) );
  NOR2X0 U10441 ( .IN1(n10397), .IN2(n8832), .QN(n10396) );
  NAND2X0 U10442 ( .IN1(n10398), .IN2(n10399), .QN(g34467) );
  NAND3X0 U10443 ( .IN1(n10400), .IN2(n10401), .IN3(n10402), .QN(n10399) );
  NAND2X0 U10444 ( .IN1(n8363), .IN2(n10403), .QN(n10401) );
  NAND2X0 U10445 ( .IN1(n10395), .IN2(g4854), .QN(n10400) );
  INVX0 U10446 ( .INP(n10403), .ZN(n10395) );
  NAND2X0 U10447 ( .IN1(n2563), .IN2(g4849), .QN(n10403) );
  NAND2X0 U10448 ( .IN1(n9479), .IN2(g4849), .QN(n10398) );
  NAND2X0 U10449 ( .IN1(n10404), .IN2(n10405), .QN(g34466) );
  NAND2X0 U10450 ( .IN1(n10406), .IN2(g4878), .QN(n10405) );
  NAND2X0 U10451 ( .IN1(n10407), .IN2(n9382), .QN(n10406) );
  NAND2X0 U10452 ( .IN1(n8833), .IN2(n10394), .QN(n10407) );
  NAND3X0 U10453 ( .IN1(n10402), .IN2(g4843), .IN3(n5283), .QN(n10404) );
  NAND3X0 U10454 ( .IN1(n10408), .IN2(n10409), .IN3(n10410), .QN(g34465) );
  NAND2X0 U10455 ( .IN1(n9479), .IN2(g4843), .QN(n10410) );
  NAND3X0 U10456 ( .IN1(n10394), .IN2(n2563), .IN3(n8834), .QN(n10409) );
  NAND2X0 U10457 ( .IN1(n2567), .IN2(n10402), .QN(n10408) );
  INVX0 U10458 ( .INP(n10397), .ZN(n10402) );
  NAND2X0 U10459 ( .IN1(n10411), .IN2(n10412), .QN(g34464) );
  NAND2X0 U10460 ( .IN1(n10413), .IN2(g4664), .QN(n10412) );
  NAND2X0 U10461 ( .IN1(n10414), .IN2(n9381), .QN(n10413) );
  NAND2X0 U10462 ( .IN1(n10415), .IN2(n10416), .QN(n10414) );
  INVX0 U10463 ( .INP(n10417), .ZN(n10411) );
  NOR2X0 U10464 ( .IN1(n10418), .IN2(n8830), .QN(n10417) );
  NAND2X0 U10465 ( .IN1(n10419), .IN2(n10420), .QN(g34463) );
  NAND3X0 U10466 ( .IN1(n10421), .IN2(n10422), .IN3(n10423), .QN(n10420) );
  NAND2X0 U10467 ( .IN1(n8377), .IN2(n10424), .QN(n10422) );
  NAND2X0 U10468 ( .IN1(n10416), .IN2(g4664), .QN(n10421) );
  INVX0 U10469 ( .INP(n10424), .ZN(n10416) );
  NAND2X0 U10470 ( .IN1(n2573), .IN2(g4659), .QN(n10424) );
  NAND2X0 U10471 ( .IN1(n9479), .IN2(g4659), .QN(n10419) );
  NAND2X0 U10472 ( .IN1(n10425), .IN2(n10426), .QN(g34462) );
  NAND2X0 U10473 ( .IN1(n10427), .IN2(g4688), .QN(n10426) );
  NAND2X0 U10474 ( .IN1(n10428), .IN2(n9381), .QN(n10427) );
  NAND2X0 U10475 ( .IN1(n10415), .IN2(n8881), .QN(n10428) );
  NAND3X0 U10476 ( .IN1(n10423), .IN2(test_so19), .IN3(n5656), .QN(n10425) );
  NAND3X0 U10477 ( .IN1(n10429), .IN2(n10430), .IN3(n10431), .QN(g34461) );
  NAND2X0 U10478 ( .IN1(test_so19), .IN2(n9415), .QN(n10431) );
  NAND3X0 U10479 ( .IN1(n10415), .IN2(n2573), .IN3(n8831), .QN(n10430) );
  NAND2X0 U10480 ( .IN1(n2577), .IN2(n10423), .QN(n10429) );
  INVX0 U10481 ( .INP(n10418), .ZN(n10423) );
  NAND2X0 U10482 ( .IN1(n10432), .IN2(n10433), .QN(g34460) );
  NAND2X0 U10483 ( .IN1(n10434), .IN2(g4639), .QN(n10433) );
  NAND2X0 U10484 ( .IN1(n10435), .IN2(n9381), .QN(n10434) );
  NAND2X0 U10485 ( .IN1(n10436), .IN2(n8873), .QN(n10435) );
  NAND2X0 U10486 ( .IN1(n408), .IN2(test_so3), .QN(n10432) );
  INVX0 U10487 ( .INP(n10437), .ZN(n408) );
  NAND2X0 U10488 ( .IN1(n10438), .IN2(n10439), .QN(g34459) );
  NAND2X0 U10489 ( .IN1(n9479), .IN2(g4643), .QN(n10439) );
  NAND2X0 U10490 ( .IN1(n10440), .IN2(n9381), .QN(n10438) );
  NAND2X0 U10491 ( .IN1(n10441), .IN2(n10442), .QN(n10440) );
  NAND2X0 U10492 ( .IN1(n10443), .IN2(n10444), .QN(n10442) );
  NAND2X0 U10493 ( .IN1(n5653), .IN2(n10445), .QN(n10443) );
  NAND2X0 U10494 ( .IN1(test_so99), .IN2(n10446), .QN(n10445) );
  NAND2X0 U10495 ( .IN1(n10447), .IN2(n10448), .QN(g34458) );
  NAND2X0 U10496 ( .IN1(n10449), .IN2(g4633), .QN(n10448) );
  NAND2X0 U10497 ( .IN1(n10450), .IN2(n10451), .QN(n10449) );
  NAND3X0 U10498 ( .IN1(n9350), .IN2(n8876), .IN3(n10436), .QN(n10451) );
  INVX0 U10499 ( .INP(n10452), .ZN(n10450) );
  NAND2X0 U10500 ( .IN1(test_so99), .IN2(n10453), .QN(n10447) );
  NAND2X0 U10501 ( .IN1(n10454), .IN2(n9381), .QN(n10453) );
  NAND4X0 U10502 ( .IN1(n5844), .IN2(n10436), .IN3(test_so3), .IN4(g4639), 
        .QN(n10454) );
  NAND2X0 U10503 ( .IN1(n10455), .IN2(n10456), .QN(g34457) );
  NAND2X0 U10504 ( .IN1(test_so3), .IN2(n10457), .QN(n10456) );
  NAND2X0 U10505 ( .IN1(n10458), .IN2(n9380), .QN(n10457) );
  NAND3X0 U10506 ( .IN1(g4639), .IN2(n8876), .IN3(n10436), .QN(n10458) );
  NAND2X0 U10507 ( .IN1(test_so99), .IN2(n10452), .QN(n10455) );
  NAND2X0 U10508 ( .IN1(n10437), .IN2(n10459), .QN(n10452) );
  NAND3X0 U10509 ( .IN1(n9350), .IN2(n8873), .IN3(n10436), .QN(n10459) );
  NAND3X0 U10510 ( .IN1(n5382), .IN2(n10460), .IN3(n5727), .QN(n10437) );
  NAND2X0 U10511 ( .IN1(n10461), .IN2(n10462), .QN(g34456) );
  NAND2X0 U10512 ( .IN1(n10463), .IN2(g4608), .QN(n10462) );
  NAND2X0 U10513 ( .IN1(n10464), .IN2(n9380), .QN(n10463) );
  NAND2X0 U10514 ( .IN1(n2590), .IN2(n10465), .QN(n10464) );
  NAND2X0 U10515 ( .IN1(n10466), .IN2(g4616), .QN(n10461) );
  NAND2X0 U10516 ( .IN1(n10467), .IN2(n10468), .QN(g34455) );
  NAND2X0 U10517 ( .IN1(n10469), .IN2(g4322), .QN(n10468) );
  NAND2X0 U10518 ( .IN1(n10470), .IN2(n9380), .QN(n10469) );
  NAND3X0 U10519 ( .IN1(n10471), .IN2(n10441), .IN3(n2594), .QN(n10470) );
  NAND2X0 U10520 ( .IN1(n2595), .IN2(g4332), .QN(n10467) );
  NAND2X0 U10521 ( .IN1(n10472), .IN2(n10473), .QN(g34454) );
  NAND3X0 U10522 ( .IN1(n10474), .IN2(n10475), .IN3(n10466), .QN(n10473) );
  INVX0 U10523 ( .INP(n10476), .ZN(n10475) );
  NOR2X0 U10524 ( .IN1(g4608), .IN2(n2590), .QN(n10476) );
  NAND2X0 U10525 ( .IN1(n2590), .IN2(g4608), .QN(n10474) );
  NAND2X0 U10526 ( .IN1(n9479), .IN2(g4601), .QN(n10472) );
  NAND3X0 U10527 ( .IN1(n10477), .IN2(n10478), .IN3(n10479), .QN(g34453) );
  NAND2X0 U10528 ( .IN1(n9479), .IN2(g4593), .QN(n10479) );
  NAND3X0 U10529 ( .IN1(n10466), .IN2(n10480), .IN3(g4601), .QN(n10478) );
  INVX0 U10530 ( .INP(n2598), .ZN(n10480) );
  NAND3X0 U10531 ( .IN1(n2598), .IN2(n10465), .IN3(n5365), .QN(n10477) );
  NAND2X0 U10532 ( .IN1(n10481), .IN2(n10482), .QN(g34452) );
  NAND3X0 U10533 ( .IN1(n10483), .IN2(n10484), .IN3(n10466), .QN(n10482) );
  NAND2X0 U10534 ( .IN1(n5303), .IN2(n10485), .QN(n10484) );
  NAND2X0 U10535 ( .IN1(n101), .IN2(g4593), .QN(n10483) );
  NAND2X0 U10536 ( .IN1(n9478), .IN2(g4584), .QN(n10481) );
  NAND2X0 U10537 ( .IN1(n10486), .IN2(n10487), .QN(g34451) );
  NAND3X0 U10538 ( .IN1(n10488), .IN2(n10485), .IN3(n10466), .QN(n10487) );
  NOR2X0 U10539 ( .IN1(n10489), .IN2(n9390), .QN(n10466) );
  INVX0 U10540 ( .INP(n10465), .ZN(n10489) );
  NOR2X0 U10541 ( .IN1(n10490), .IN2(n10491), .QN(n10465) );
  NOR2X0 U10542 ( .IN1(n10485), .IN2(n5608), .QN(n10491) );
  INVX0 U10543 ( .INP(n101), .ZN(n10485) );
  NOR2X0 U10544 ( .IN1(n10471), .IN2(n5539), .QN(n101) );
  NAND2X0 U10545 ( .IN1(n5539), .IN2(n10471), .QN(n10488) );
  NAND2X0 U10546 ( .IN1(n9478), .IN2(g4332), .QN(n10486) );
  NAND3X0 U10547 ( .IN1(n10492), .IN2(n10493), .IN3(n10494), .QN(g34450) );
  NAND2X0 U10548 ( .IN1(n9478), .IN2(g4311), .QN(n10494) );
  NAND3X0 U10549 ( .IN1(n2595), .IN2(n10495), .IN3(g4322), .QN(n10493) );
  INVX0 U10550 ( .INP(n2594), .ZN(n10495) );
  INVX0 U10551 ( .INP(n10496), .ZN(n2595) );
  NAND2X0 U10552 ( .IN1(n10460), .IN2(n10471), .QN(n10496) );
  NAND3X0 U10553 ( .IN1(g4322), .IN2(g4332), .IN3(n103), .QN(n10471) );
  INVX0 U10554 ( .INP(n9799), .ZN(n103) );
  NAND2X0 U10555 ( .IN1(n10497), .IN2(g4358), .QN(n9799) );
  NAND3X0 U10556 ( .IN1(n2594), .IN2(n10441), .IN3(n5506), .QN(n10492) );
  NAND3X0 U10557 ( .IN1(n10498), .IN2(n10499), .IN3(n10500), .QN(g34448) );
  NAND2X0 U10558 ( .IN1(n9478), .IN2(g2827), .QN(n10500) );
  NAND3X0 U10559 ( .IN1(n9350), .IN2(g2819), .IN3(n10501), .QN(n10499) );
  NAND3X0 U10560 ( .IN1(n10502), .IN2(n10503), .IN3(n10504), .QN(n10498) );
  NAND2X0 U10561 ( .IN1(n10505), .IN2(g2827), .QN(n10503) );
  NAND3X0 U10562 ( .IN1(n10506), .IN2(n10507), .IN3(n10508), .QN(g34447) );
  NAND2X0 U10563 ( .IN1(n9478), .IN2(g2815), .QN(n10508) );
  NAND3X0 U10564 ( .IN1(n9350), .IN2(g2807), .IN3(n10509), .QN(n10507) );
  NAND3X0 U10565 ( .IN1(n10502), .IN2(n10510), .IN3(n10511), .QN(n10506) );
  NAND2X0 U10566 ( .IN1(n10505), .IN2(g2811), .QN(n10510) );
  NAND3X0 U10567 ( .IN1(n10512), .IN2(n10513), .IN3(n10514), .QN(g34446) );
  NAND2X0 U10568 ( .IN1(n9478), .IN2(g2819), .QN(n10514) );
  NAND3X0 U10569 ( .IN1(n9350), .IN2(g2815), .IN3(n10515), .QN(n10513) );
  NAND3X0 U10570 ( .IN1(n10502), .IN2(n10516), .IN3(n10517), .QN(n10512) );
  NAND2X0 U10571 ( .IN1(test_so37), .IN2(n10505), .QN(n10516) );
  NAND3X0 U10572 ( .IN1(n10518), .IN2(n10519), .IN3(n10520), .QN(g34445) );
  NAND2X0 U10573 ( .IN1(n9478), .IN2(g2807), .QN(n10520) );
  NAND3X0 U10574 ( .IN1(n9353), .IN2(g2803), .IN3(n10521), .QN(n10519) );
  NAND3X0 U10575 ( .IN1(n10502), .IN2(n10522), .IN3(n10523), .QN(n10518) );
  NAND2X0 U10576 ( .IN1(n10505), .IN2(g2799), .QN(n10522) );
  INVX0 U10577 ( .INP(n10524), .ZN(n10502) );
  NAND2X0 U10578 ( .IN1(n10525), .IN2(n9380), .QN(n10524) );
  NAND2X0 U10579 ( .IN1(n2760), .IN2(n9255), .QN(n10525) );
  NAND3X0 U10580 ( .IN1(n10526), .IN2(n10527), .IN3(n10528), .QN(g34444) );
  NAND2X0 U10581 ( .IN1(n9477), .IN2(g2795), .QN(n10528) );
  NAND3X0 U10582 ( .IN1(n9353), .IN2(g2787), .IN3(n10501), .QN(n10527) );
  INVX0 U10583 ( .INP(n10504), .ZN(n10501) );
  NAND3X0 U10584 ( .IN1(n10529), .IN2(n10530), .IN3(n10504), .QN(n10526) );
  NOR2X0 U10585 ( .IN1(n10531), .IN2(n10532), .QN(n10504) );
  NAND2X0 U10586 ( .IN1(n10505), .IN2(g2795), .QN(n10530) );
  NAND3X0 U10587 ( .IN1(n10533), .IN2(n10534), .IN3(n10535), .QN(g34443) );
  NAND2X0 U10588 ( .IN1(n9477), .IN2(g2783), .QN(n10535) );
  NAND3X0 U10589 ( .IN1(n9353), .IN2(g2775), .IN3(n10509), .QN(n10534) );
  INVX0 U10590 ( .INP(n10511), .ZN(n10509) );
  NAND3X0 U10591 ( .IN1(n10529), .IN2(n10536), .IN3(n10511), .QN(n10533) );
  NOR2X0 U10592 ( .IN1(n10537), .IN2(n10531), .QN(n10511) );
  NAND2X0 U10593 ( .IN1(n10505), .IN2(g2779), .QN(n10536) );
  NAND3X0 U10594 ( .IN1(n10538), .IN2(n10539), .IN3(n10540), .QN(g34442) );
  NAND2X0 U10595 ( .IN1(n9477), .IN2(g2787), .QN(n10540) );
  NAND3X0 U10596 ( .IN1(n9353), .IN2(g2783), .IN3(n10515), .QN(n10539) );
  INVX0 U10597 ( .INP(n10517), .ZN(n10515) );
  NAND3X0 U10598 ( .IN1(n10529), .IN2(n10541), .IN3(n10517), .QN(n10538) );
  NOR2X0 U10599 ( .IN1(n10542), .IN2(n10531), .QN(n10517) );
  NAND2X0 U10600 ( .IN1(n10505), .IN2(g2791), .QN(n10541) );
  NAND3X0 U10601 ( .IN1(n10543), .IN2(n10544), .IN3(n10545), .QN(g34441) );
  NAND2X0 U10602 ( .IN1(n9477), .IN2(g2775), .QN(n10545) );
  NAND3X0 U10603 ( .IN1(n9353), .IN2(g2771), .IN3(n10521), .QN(n10544) );
  INVX0 U10604 ( .INP(n10523), .ZN(n10521) );
  NAND3X0 U10605 ( .IN1(n10529), .IN2(n10546), .IN3(n10523), .QN(n10543) );
  NOR2X0 U10606 ( .IN1(n10531), .IN2(n10547), .QN(n10523) );
  NAND2X0 U10607 ( .IN1(n10505), .IN2(g2767), .QN(n10546) );
  INVX0 U10608 ( .INP(n10548), .ZN(n10529) );
  NAND2X0 U10609 ( .IN1(n10549), .IN2(n9380), .QN(n10548) );
  NAND2X0 U10610 ( .IN1(n2760), .IN2(n9265), .QN(n10549) );
  NAND2X0 U10611 ( .IN1(n10550), .IN2(n10551), .QN(g34440) );
  NAND2X0 U10612 ( .IN1(n9477), .IN2(g446), .QN(n10551) );
  NAND2X0 U10613 ( .IN1(n10552), .IN2(n9380), .QN(n10550) );
  NAND2X0 U10614 ( .IN1(n10553), .IN2(n10554), .QN(n10552) );
  NAND2X0 U10615 ( .IN1(n10555), .IN2(g862), .QN(n10554) );
  NAND2X0 U10616 ( .IN1(g896), .IN2(n10556), .QN(n10555) );
  NAND2X0 U10617 ( .IN1(n10557), .IN2(n10558), .QN(n10556) );
  NAND3X0 U10618 ( .IN1(n10559), .IN2(n10560), .IN3(n5821), .QN(n10557) );
  NAND2X0 U10619 ( .IN1(g890), .IN2(g896), .QN(n10553) );
  NAND3X0 U10620 ( .IN1(n10561), .IN2(n10562), .IN3(n10563), .QN(g34439) );
  NAND2X0 U10621 ( .IN1(n9477), .IN2(g772), .QN(n10563) );
  NAND3X0 U10622 ( .IN1(n2404), .IN2(n10564), .IN3(g776), .QN(n10562) );
  INVX0 U10623 ( .INP(n2554), .ZN(n10564) );
  NAND2X0 U10624 ( .IN1(n2554), .IN2(n5330), .QN(n10561) );
  NAND3X0 U10625 ( .IN1(n10565), .IN2(n10566), .IN3(n10567), .QN(g34438) );
  NAND2X0 U10626 ( .IN1(n9477), .IN2(g604), .QN(n10567) );
  NAND3X0 U10627 ( .IN1(n2421), .IN2(n10568), .IN3(g608), .QN(n10566) );
  INVX0 U10628 ( .INP(n2556), .ZN(n10568) );
  NAND2X0 U10629 ( .IN1(n2556), .IN2(n5475), .QN(n10565) );
  NOR4X0 U10630 ( .IN1(n10569), .IN2(g4064), .IN3(g4057), .IN4(g4125), .QN(
        g34435) );
  NOR3X0 U10631 ( .IN1(g4082), .IN2(n10570), .IN3(g4141), .QN(n10569) );
  NOR4X0 U10632 ( .IN1(n8708), .IN2(n10571), .IN3(g4098), .IN4(n8878), .QN(
        n10570) );
  NAND2X0 U10633 ( .IN1(n2730), .IN2(n10572), .QN(g34425) );
  INVX0 U10634 ( .INP(n8847), .ZN(n10572) );
  NAND2X0 U10635 ( .IN1(n10573), .IN2(n10574), .QN(n8847) );
  NAND2X0 U10636 ( .IN1(n10575), .IN2(g4358), .QN(n10574) );
  NAND2X0 U10637 ( .IN1(n10576), .IN2(n10577), .QN(n10575) );
  NAND2X0 U10638 ( .IN1(test_so81), .IN2(n10578), .QN(n10577) );
  NAND2X0 U10639 ( .IN1(n10579), .IN2(n10580), .QN(n10578) );
  NAND2X0 U10640 ( .IN1(n10581), .IN2(n10255), .QN(n10580) );
  NAND2X0 U10641 ( .IN1(n10582), .IN2(n10252), .QN(n10579) );
  NAND2X0 U10642 ( .IN1(n10583), .IN2(n8867), .QN(n10576) );
  NAND2X0 U10643 ( .IN1(n10584), .IN2(n10585), .QN(n10583) );
  NAND2X0 U10644 ( .IN1(n10586), .IN2(n10255), .QN(n10585) );
  NAND2X0 U10645 ( .IN1(n10587), .IN2(n10252), .QN(n10584) );
  NAND2X0 U10646 ( .IN1(n10588), .IN2(n5348), .QN(n10573) );
  NAND2X0 U10647 ( .IN1(n10589), .IN2(n10590), .QN(n10588) );
  NAND2X0 U10648 ( .IN1(test_so81), .IN2(n10591), .QN(n10590) );
  NAND2X0 U10649 ( .IN1(n10592), .IN2(n10593), .QN(n10591) );
  NAND2X0 U10650 ( .IN1(n10594), .IN2(n10255), .QN(n10593) );
  NAND2X0 U10651 ( .IN1(n10595), .IN2(n10252), .QN(n10592) );
  NAND2X0 U10652 ( .IN1(n10596), .IN2(n8867), .QN(n10589) );
  NAND2X0 U10653 ( .IN1(n10597), .IN2(n10598), .QN(n10596) );
  NAND2X0 U10654 ( .IN1(g31860), .IN2(n10255), .QN(n10598) );
  NAND2X0 U10655 ( .IN1(n9684), .IN2(n10252), .QN(n10597) );
  NOR2X0 U10656 ( .IN1(n10599), .IN2(n10600), .QN(n2730) );
  NOR2X0 U10657 ( .IN1(n10252), .IN2(n10255), .QN(n10600) );
  NAND3X0 U10658 ( .IN1(n10601), .IN2(n10602), .IN3(n10603), .QN(g34383) );
  INVX0 U10659 ( .INP(g34843), .ZN(n10602) );
  NAND4X0 U10660 ( .IN1(n10604), .IN2(n10605), .IN3(n10606), .IN4(n10607), 
        .QN(g34843) );
  NOR4X0 U10661 ( .IN1(n10608), .IN2(n10609), .IN3(n10610), .IN4(n10611), .QN(
        n10607) );
  NOR2X0 U10662 ( .IN1(n10612), .IN2(n10613), .QN(n10611) );
  NOR2X0 U10663 ( .IN1(n1013), .IN2(n10614), .QN(n10610) );
  INVX0 U10664 ( .INP(n10615), .ZN(n1013) );
  NOR2X0 U10665 ( .IN1(n999), .IN2(n10616), .QN(n10609) );
  INVX0 U10666 ( .INP(n10617), .ZN(n999) );
  NOR2X0 U10667 ( .IN1(n10618), .IN2(n10619), .QN(n10608) );
  NOR2X0 U10668 ( .IN1(n10620), .IN2(n10621), .QN(n10606) );
  NOR2X0 U10669 ( .IN1(n10622), .IN2(n10623), .QN(n10621) );
  NOR2X0 U10670 ( .IN1(n3146), .IN2(n10624), .QN(n10620) );
  NAND3X0 U10671 ( .IN1(n10625), .IN2(g1802), .IN3(n5504), .QN(n10605) );
  NAND2X0 U10672 ( .IN1(n10626), .IN2(n10627), .QN(n10604) );
  NAND4X0 U10673 ( .IN1(n10623), .IN2(n10628), .IN3(n10619), .IN4(n10629), 
        .QN(n10601) );
  INVX0 U10674 ( .INP(n10630), .ZN(n10629) );
  NAND4X0 U10675 ( .IN1(n10631), .IN2(n3165), .IN3(n3146), .IN4(n10612), .QN(
        n10630) );
  NAND2X0 U10676 ( .IN1(n10632), .IN2(n10633), .QN(g34269) );
  NAND2X0 U10677 ( .IN1(n9476), .IN2(g4961), .QN(n10633) );
  NAND3X0 U10678 ( .IN1(n10634), .IN2(n10635), .IN3(n10636), .QN(n10632) );
  NAND3X0 U10679 ( .IN1(n5614), .IN2(n10637), .IN3(n10638), .QN(n10635) );
  INVX0 U10680 ( .INP(n10639), .ZN(n10638) );
  NAND3X0 U10681 ( .IN1(n5770), .IN2(n10640), .IN3(n10639), .QN(n10634) );
  NAND2X0 U10682 ( .IN1(n10641), .IN2(n10642), .QN(g34268) );
  NAND2X0 U10683 ( .IN1(n9476), .IN2(g4950), .QN(n10642) );
  NAND3X0 U10684 ( .IN1(n10643), .IN2(n10644), .IN3(n10636), .QN(n10641) );
  NAND3X0 U10685 ( .IN1(n5875), .IN2(n10637), .IN3(n10645), .QN(n10644) );
  INVX0 U10686 ( .INP(n10646), .ZN(n10645) );
  NAND3X0 U10687 ( .IN1(n5772), .IN2(n10640), .IN3(n10646), .QN(n10643) );
  NAND2X0 U10688 ( .IN1(n10647), .IN2(n10648), .QN(g34267) );
  NAND2X0 U10689 ( .IN1(n10649), .IN2(n9380), .QN(n10648) );
  NAND2X0 U10690 ( .IN1(n10640), .IN2(n10650), .QN(n10649) );
  NAND3X0 U10691 ( .IN1(n10637), .IN2(g4933), .IN3(n10651), .QN(n10650) );
  NAND2X0 U10692 ( .IN1(n10652), .IN2(g4939), .QN(n10647) );
  NAND2X0 U10693 ( .IN1(n10653), .IN2(n9380), .QN(n10652) );
  NAND2X0 U10694 ( .IN1(n10654), .IN2(n10637), .QN(n10653) );
  NAND2X0 U10695 ( .IN1(n10655), .IN2(n10656), .QN(g34266) );
  NAND2X0 U10696 ( .IN1(n9476), .IN2(g4894), .QN(n10656) );
  NAND3X0 U10697 ( .IN1(n10657), .IN2(n10658), .IN3(n10636), .QN(n10655) );
  NOR2X0 U10698 ( .IN1(n10659), .IN2(n9389), .QN(n10636) );
  INVX0 U10699 ( .INP(n10660), .ZN(n10659) );
  NAND2X0 U10700 ( .IN1(n10661), .IN2(n10640), .QN(n10660) );
  NAND3X0 U10701 ( .IN1(n5863), .IN2(n10637), .IN3(n10662), .QN(n10658) );
  NAND3X0 U10702 ( .IN1(n5774), .IN2(n10640), .IN3(n10251), .QN(n10657) );
  NAND2X0 U10703 ( .IN1(n10661), .IN2(g71), .QN(n10640) );
  INVX0 U10704 ( .INP(n10637), .ZN(n10661) );
  NAND3X0 U10705 ( .IN1(n2668), .IN2(DFF_672_n1), .IN3(n5637), .QN(n10637) );
  NOR4X0 U10706 ( .IN1(g4864), .IN2(g4871), .IN3(g4836), .IN4(n10397), .QN(
        g34265) );
  NAND2X0 U10707 ( .IN1(n10394), .IN2(n9380), .QN(n10397) );
  NOR2X0 U10708 ( .IN1(n10663), .IN2(n10253), .QN(n10394) );
  NAND2X0 U10709 ( .IN1(n10664), .IN2(n10665), .QN(g34264) );
  NAND2X0 U10710 ( .IN1(n9476), .IN2(g4771), .QN(n10665) );
  NAND3X0 U10711 ( .IN1(n10666), .IN2(n10667), .IN3(n10668), .QN(n10664) );
  NAND3X0 U10712 ( .IN1(n5613), .IN2(n10669), .IN3(n10670), .QN(n10667) );
  INVX0 U10713 ( .INP(n10671), .ZN(n10670) );
  NAND3X0 U10714 ( .IN1(n5769), .IN2(n10672), .IN3(n10671), .QN(n10666) );
  NAND2X0 U10715 ( .IN1(n10673), .IN2(n10674), .QN(g34263) );
  NAND2X0 U10716 ( .IN1(n9476), .IN2(g4760), .QN(n10674) );
  NAND3X0 U10717 ( .IN1(n10675), .IN2(n10676), .IN3(n10668), .QN(n10673) );
  NAND3X0 U10718 ( .IN1(n5877), .IN2(n10669), .IN3(n10677), .QN(n10676) );
  INVX0 U10719 ( .INP(n10678), .ZN(n10677) );
  NAND3X0 U10720 ( .IN1(n5775), .IN2(n10672), .IN3(n10678), .QN(n10675) );
  NAND2X0 U10721 ( .IN1(n10679), .IN2(n10680), .QN(g34262) );
  NAND2X0 U10722 ( .IN1(n10681), .IN2(n9380), .QN(n10680) );
  NAND2X0 U10723 ( .IN1(n10672), .IN2(n10682), .QN(n10681) );
  NAND3X0 U10724 ( .IN1(n10669), .IN2(g4743), .IN3(n10683), .QN(n10682) );
  NAND2X0 U10725 ( .IN1(test_so18), .IN2(n10684), .QN(n10679) );
  NAND2X0 U10726 ( .IN1(n10685), .IN2(n9380), .QN(n10684) );
  NAND2X0 U10727 ( .IN1(n10686), .IN2(n10669), .QN(n10685) );
  NAND2X0 U10728 ( .IN1(n10687), .IN2(n10688), .QN(g34261) );
  NAND2X0 U10729 ( .IN1(n9476), .IN2(g4704), .QN(n10688) );
  NAND3X0 U10730 ( .IN1(n10689), .IN2(n10690), .IN3(n10668), .QN(n10687) );
  NOR2X0 U10731 ( .IN1(n10691), .IN2(n9387), .QN(n10668) );
  INVX0 U10732 ( .INP(n10692), .ZN(n10691) );
  NAND2X0 U10733 ( .IN1(n10693), .IN2(n10672), .QN(n10692) );
  NAND3X0 U10734 ( .IN1(n5862), .IN2(n10669), .IN3(n10694), .QN(n10690) );
  NAND3X0 U10735 ( .IN1(n5771), .IN2(n10672), .IN3(n10254), .QN(n10689) );
  NAND2X0 U10736 ( .IN1(n10693), .IN2(g101), .QN(n10672) );
  INVX0 U10737 ( .INP(n10669), .ZN(n10693) );
  NAND3X0 U10738 ( .IN1(n2668), .IN2(DFF_178_n1), .IN3(n5636), .QN(n10669) );
  NOR4X0 U10739 ( .IN1(g4674), .IN2(g4646), .IN3(g4681), .IN4(n10418), .QN(
        g34260) );
  NAND2X0 U10740 ( .IN1(n10415), .IN2(n9380), .QN(n10418) );
  NOR2X0 U10741 ( .IN1(n10256), .IN2(n10695), .QN(n10415) );
  NOR2X0 U10742 ( .IN1(n5844), .IN2(n10696), .QN(g34259) );
  NOR2X0 U10743 ( .IN1(n9418), .IN2(n10697), .QN(n10696) );
  NOR2X0 U10744 ( .IN1(n10698), .IN2(n10699), .QN(n10697) );
  INVX0 U10745 ( .INP(n10436), .ZN(n10699) );
  NOR2X0 U10746 ( .IN1(g4643), .IN2(n10490), .QN(n10436) );
  NAND3X0 U10747 ( .IN1(n10700), .IN2(n10701), .IN3(n10702), .QN(g34258) );
  NAND2X0 U10748 ( .IN1(test_so81), .IN2(n9412), .QN(n10702) );
  NAND3X0 U10749 ( .IN1(n10460), .IN2(n10703), .IN3(g4358), .QN(n10701) );
  INVX0 U10750 ( .INP(n10497), .ZN(n10703) );
  NAND3X0 U10751 ( .IN1(n10497), .IN2(n10441), .IN3(n5348), .QN(n10700) );
  NOR2X0 U10752 ( .IN1(n10444), .IN2(n8867), .QN(n10497) );
  NAND3X0 U10753 ( .IN1(n10704), .IN2(n10705), .IN3(n10706), .QN(g34257) );
  NAND2X0 U10754 ( .IN1(n9476), .IN2(g4340), .QN(n10706) );
  NAND3X0 U10755 ( .IN1(n10460), .IN2(test_so81), .IN3(n10444), .QN(n10705) );
  NOR2X0 U10756 ( .IN1(n10490), .IN2(n9387), .QN(n10460) );
  INVX0 U10757 ( .INP(n10441), .ZN(n10490) );
  NAND3X0 U10758 ( .IN1(n10441), .IN2(n8867), .IN3(n10707), .QN(n10704) );
  INVX0 U10759 ( .INP(n10444), .ZN(n10707) );
  NAND3X0 U10760 ( .IN1(n10446), .IN2(g4340), .IN3(test_so99), .QN(n10444) );
  NAND2X0 U10761 ( .IN1(n9281), .IN2(n10708), .QN(n10441) );
  NAND2X0 U10762 ( .IN1(n10145), .IN2(n1835), .QN(n10708) );
  NAND2X0 U10763 ( .IN1(n10709), .IN2(n10710), .QN(g34256) );
  INVX0 U10764 ( .INP(n10711), .ZN(n10710) );
  NOR2X0 U10765 ( .IN1(n9360), .IN2(n8591), .QN(n10711) );
  NAND2X0 U10766 ( .IN1(n10712), .IN2(n9380), .QN(n10709) );
  NAND3X0 U10767 ( .IN1(n10713), .IN2(n10714), .IN3(n5765), .QN(n10712) );
  NAND2X0 U10768 ( .IN1(n5671), .IN2(g4473), .QN(n10713) );
  NAND4X0 U10769 ( .IN1(n5671), .IN2(n10715), .IN3(n10714), .IN4(n9362), .QN(
        g34255) );
  NAND2X0 U10770 ( .IN1(test_so38), .IN2(g4473), .QN(n10715) );
  NAND2X0 U10771 ( .IN1(n10716), .IN2(n10717), .QN(g34254) );
  NAND2X0 U10772 ( .IN1(n10718), .IN2(g4473), .QN(n10717) );
  NAND4X0 U10773 ( .IN1(n9362), .IN2(g4643), .IN3(g4462), .IN4(n8864), .QN(
        n10718) );
  NAND2X0 U10774 ( .IN1(n10719), .IN2(n9380), .QN(n10716) );
  NOR2X0 U10775 ( .IN1(n9418), .IN2(n10720), .QN(g34253) );
  NOR3X0 U10776 ( .IN1(n8864), .IN2(n5671), .IN3(n10719), .QN(n10720) );
  INVX0 U10777 ( .INP(n10714), .ZN(n10719) );
  NAND3X0 U10778 ( .IN1(n10721), .IN2(g26960), .IN3(n5849), .QN(n10714) );
  NAND2X0 U10779 ( .IN1(n10145), .IN2(n10722), .QN(n10721) );
  NAND2X0 U10780 ( .IN1(n5846), .IN2(n2668), .QN(n10722) );
  NAND3X0 U10781 ( .IN1(n10723), .IN2(n10724), .IN3(n10725), .QN(g34252) );
  NAND2X0 U10782 ( .IN1(n9475), .IN2(g767), .QN(n10725) );
  NAND3X0 U10783 ( .IN1(n2404), .IN2(n10726), .IN3(g772), .QN(n10724) );
  INVX0 U10784 ( .INP(n2647), .ZN(n10726) );
  NAND2X0 U10785 ( .IN1(n2647), .IN2(n5334), .QN(n10723) );
  NAND3X0 U10786 ( .IN1(n10727), .IN2(n10728), .IN3(n10729), .QN(g34251) );
  NAND2X0 U10787 ( .IN1(n9475), .IN2(g599), .QN(n10729) );
  NAND3X0 U10788 ( .IN1(n2421), .IN2(n10730), .IN3(g604), .QN(n10728) );
  INVX0 U10789 ( .INP(n2649), .ZN(n10730) );
  NAND2X0 U10790 ( .IN1(n2649), .IN2(n5473), .QN(n10727) );
  NAND3X0 U10791 ( .IN1(n10731), .IN2(n10732), .IN3(n10733), .QN(g34250) );
  NAND2X0 U10792 ( .IN1(n9475), .IN2(g298), .QN(n10733) );
  NAND3X0 U10793 ( .IN1(n10734), .IN2(n10735), .IN3(g142), .QN(n10732) );
  INVX0 U10794 ( .INP(n2707), .ZN(n10735) );
  NAND2X0 U10795 ( .IN1(n5724), .IN2(n2707), .QN(n10731) );
  NAND3X0 U10796 ( .IN1(n10736), .IN2(n10737), .IN3(n10738), .QN(g34249) );
  NAND2X0 U10797 ( .IN1(n9475), .IN2(g157), .QN(n10738) );
  NAND3X0 U10798 ( .IN1(n10739), .IN2(n10740), .IN3(g160), .QN(n10737) );
  INVX0 U10799 ( .INP(n2710), .ZN(n10740) );
  NAND2X0 U10800 ( .IN1(n2710), .IN2(n5843), .QN(n10736) );
  NAND3X0 U10801 ( .IN1(n10741), .IN2(n10742), .IN3(n10603), .QN(g34201) );
  INVX0 U10802 ( .INP(g34781), .ZN(n10742) );
  NAND4X0 U10803 ( .IN1(n10743), .IN2(n10744), .IN3(n10745), .IN4(n10746), 
        .QN(g34781) );
  NOR4X0 U10804 ( .IN1(n10747), .IN2(n10748), .IN3(n10749), .IN4(n10750), .QN(
        n10746) );
  NOR3X0 U10805 ( .IN1(g2217), .IN2(n8756), .IN3(n3569), .QN(n10750) );
  NOR3X0 U10806 ( .IN1(g2351), .IN2(n3550), .IN3(n8869), .QN(n10749) );
  NOR3X0 U10807 ( .IN1(g2485), .IN2(n8758), .IN3(n3007), .QN(n10748) );
  NOR3X0 U10808 ( .IN1(g2619), .IN2(n8759), .IN3(n3006), .QN(n10747) );
  NOR2X0 U10809 ( .IN1(n10751), .IN2(n10752), .QN(n10745) );
  NOR2X0 U10810 ( .IN1(n3003), .IN2(n10753), .QN(n10752) );
  NOR3X0 U10811 ( .IN1(g1792), .IN2(n5596), .IN3(n1774), .QN(n10751) );
  NAND3X0 U10812 ( .IN1(n10754), .IN2(g2051), .IN3(n5507), .QN(n10744) );
  NAND3X0 U10813 ( .IN1(n10755), .IN2(g1917), .IN3(n5510), .QN(n10743) );
  NAND4X0 U10814 ( .IN1(n3588), .IN2(n3606), .IN3(n10756), .IN4(n10757), .QN(
        n10741) );
  NOR4X0 U10815 ( .IN1(n10758), .IN2(n10759), .IN3(n10760), .IN4(n10761), .QN(
        n10757) );
  NOR2X0 U10816 ( .IN1(n3005), .IN2(n10762), .QN(n10756) );
  NAND2X0 U10817 ( .IN1(n10763), .IN2(n10764), .QN(g34041) );
  NAND3X0 U10818 ( .IN1(n10765), .IN2(n10766), .IN3(n10767), .QN(n10764) );
  NAND2X0 U10819 ( .IN1(n5367), .IN2(n10768), .QN(n10766) );
  NAND2X0 U10820 ( .IN1(n10253), .IN2(g4983), .QN(n10765) );
  INVX0 U10821 ( .INP(n10768), .ZN(n10253) );
  INVX0 U10822 ( .INP(n10769), .ZN(n10763) );
  NOR2X0 U10823 ( .IN1(n9360), .IN2(n5637), .QN(n10769) );
  NAND3X0 U10824 ( .IN1(n10770), .IN2(n10771), .IN3(n10772), .QN(g34040) );
  NAND2X0 U10825 ( .IN1(n9475), .IN2(g4975), .QN(n10772) );
  NAND2X0 U10826 ( .IN1(n10773), .IN2(n10774), .QN(n10771) );
  NAND2X0 U10827 ( .IN1(n10775), .IN2(n10776), .QN(n10773) );
  NAND2X0 U10828 ( .IN1(n10777), .IN2(n9759), .QN(n10776) );
  NAND2X0 U10829 ( .IN1(n9758), .IN2(n9380), .QN(n10775) );
  NAND2X0 U10830 ( .IN1(n10767), .IN2(g4899), .QN(n10770) );
  NAND2X0 U10831 ( .IN1(n10778), .IN2(n10779), .QN(g34039) );
  NAND2X0 U10832 ( .IN1(test_so58), .IN2(n10780), .QN(n10779) );
  NAND2X0 U10833 ( .IN1(n10781), .IN2(n9380), .QN(n10780) );
  NAND2X0 U10834 ( .IN1(n10782), .IN2(n10783), .QN(n10781) );
  NAND2X0 U10835 ( .IN1(n10767), .IN2(g4966), .QN(n10778) );
  NAND3X0 U10836 ( .IN1(n10784), .IN2(n10785), .IN3(n10786), .QN(g34038) );
  NAND2X0 U10837 ( .IN1(n9488), .IN2(g4983), .QN(n10786) );
  NAND3X0 U10838 ( .IN1(n10782), .IN2(n10783), .IN3(n8863), .QN(n10785) );
  NAND3X0 U10839 ( .IN1(n10767), .IN2(n10787), .IN3(test_so58), .QN(n10784) );
  NAND3X0 U10840 ( .IN1(n10788), .IN2(n10789), .IN3(n10790), .QN(g34037) );
  NAND2X0 U10841 ( .IN1(n9475), .IN2(g4966), .QN(n10790) );
  NAND2X0 U10842 ( .IN1(n10767), .IN2(g4975), .QN(n10789) );
  NOR2X0 U10843 ( .IN1(n10791), .IN2(n9386), .QN(n10767) );
  INVX0 U10844 ( .INP(n10782), .ZN(n10791) );
  NOR2X0 U10845 ( .IN1(n10663), .IN2(n10777), .QN(n10782) );
  INVX0 U10846 ( .INP(n10774), .ZN(n10663) );
  NAND3X0 U10847 ( .IN1(n10777), .IN2(n10774), .IN3(n5360), .QN(n10788) );
  NOR2X0 U10848 ( .IN1(n10787), .IN2(n5706), .QN(n10777) );
  INVX0 U10849 ( .INP(n10783), .ZN(n10787) );
  NOR2X0 U10850 ( .IN1(n10768), .IN2(n5367), .QN(n10783) );
  NAND2X0 U10851 ( .IN1(n10792), .IN2(g4878), .QN(n10768) );
  NOR2X0 U10852 ( .IN1(n5443), .IN2(n10793), .QN(g34036) );
  NOR2X0 U10853 ( .IN1(n5318), .IN2(n10793), .QN(g34035) );
  NOR2X0 U10854 ( .IN1(n5713), .IN2(n10793), .QN(g34034) );
  NOR2X0 U10855 ( .IN1(n10774), .IN2(n9386), .QN(n10793) );
  NAND3X0 U10856 ( .IN1(n2760), .IN2(g63), .IN3(n10252), .QN(n10774) );
  NAND2X0 U10857 ( .IN1(n10794), .IN2(n10795), .QN(g34033) );
  NAND3X0 U10858 ( .IN1(n10796), .IN2(n10797), .IN3(n10798), .QN(n10795) );
  NAND2X0 U10859 ( .IN1(n5368), .IN2(n10799), .QN(n10797) );
  NAND2X0 U10860 ( .IN1(n10256), .IN2(g4793), .QN(n10796) );
  INVX0 U10861 ( .INP(n10799), .ZN(n10256) );
  INVX0 U10862 ( .INP(n10800), .ZN(n10794) );
  NOR2X0 U10863 ( .IN1(n9360), .IN2(n5636), .QN(n10800) );
  NAND3X0 U10864 ( .IN1(n10801), .IN2(n10802), .IN3(n10803), .QN(g34032) );
  NAND2X0 U10865 ( .IN1(n9475), .IN2(g4785), .QN(n10803) );
  NAND2X0 U10866 ( .IN1(n10804), .IN2(n10805), .QN(n10802) );
  NAND2X0 U10867 ( .IN1(n10806), .IN2(n10807), .QN(n10804) );
  NAND2X0 U10868 ( .IN1(n10808), .IN2(n9724), .QN(n10807) );
  NAND2X0 U10869 ( .IN1(n9723), .IN2(n9379), .QN(n10806) );
  NAND2X0 U10870 ( .IN1(n10798), .IN2(g4709), .QN(n10801) );
  NAND2X0 U10871 ( .IN1(n10809), .IN2(n10810), .QN(g34031) );
  NAND2X0 U10872 ( .IN1(test_so29), .IN2(n10811), .QN(n10810) );
  NAND2X0 U10873 ( .IN1(n10812), .IN2(n9379), .QN(n10811) );
  NAND2X0 U10874 ( .IN1(n10813), .IN2(n10814), .QN(n10812) );
  NAND2X0 U10875 ( .IN1(n10798), .IN2(g4776), .QN(n10809) );
  NAND3X0 U10876 ( .IN1(n10815), .IN2(n10816), .IN3(n10817), .QN(g34030) );
  NAND2X0 U10877 ( .IN1(n9474), .IN2(g4793), .QN(n10817) );
  NAND3X0 U10878 ( .IN1(n10813), .IN2(n10814), .IN3(n8862), .QN(n10816) );
  NAND3X0 U10879 ( .IN1(n10798), .IN2(n10818), .IN3(test_so29), .QN(n10815) );
  NAND3X0 U10880 ( .IN1(n10819), .IN2(n10820), .IN3(n10821), .QN(g34029) );
  NAND2X0 U10881 ( .IN1(n9474), .IN2(g4776), .QN(n10821) );
  NAND2X0 U10882 ( .IN1(n10798), .IN2(g4785), .QN(n10820) );
  NOR2X0 U10883 ( .IN1(n10822), .IN2(n9386), .QN(n10798) );
  INVX0 U10884 ( .INP(n10813), .ZN(n10822) );
  NOR2X0 U10885 ( .IN1(n10695), .IN2(n10808), .QN(n10813) );
  INVX0 U10886 ( .INP(n10805), .ZN(n10695) );
  NAND3X0 U10887 ( .IN1(n10808), .IN2(n10805), .IN3(n5361), .QN(n10819) );
  NOR2X0 U10888 ( .IN1(n10818), .IN2(n5707), .QN(n10808) );
  INVX0 U10889 ( .INP(n10814), .ZN(n10818) );
  NOR2X0 U10890 ( .IN1(n10799), .IN2(n5368), .QN(n10814) );
  NAND2X0 U10891 ( .IN1(n10823), .IN2(g4688), .QN(n10799) );
  NOR2X0 U10892 ( .IN1(n5440), .IN2(n2774), .QN(g34027) );
  NOR2X0 U10893 ( .IN1(n5712), .IN2(n2774), .QN(g34026) );
  NOR2X0 U10894 ( .IN1(n10805), .IN2(n9395), .QN(n2774) );
  NAND3X0 U10895 ( .IN1(n2760), .IN2(g63), .IN3(n10255), .QN(n10805) );
  NAND4X0 U10896 ( .IN1(n10824), .IN2(n10825), .IN3(n10826), .IN4(n10827), 
        .QN(g34024) );
  NAND2X0 U10897 ( .IN1(n9474), .IN2(g4492), .QN(n10827) );
  NAND2X0 U10898 ( .IN1(n10828), .IN2(n9379), .QN(n10826) );
  NAND2X0 U10899 ( .IN1(n10829), .IN2(n10830), .QN(n10828) );
  NAND2X0 U10900 ( .IN1(n10831), .IN2(g4512), .QN(n10830) );
  NAND2X0 U10901 ( .IN1(n10832), .IN2(n10145), .QN(n10829) );
  NAND4X0 U10902 ( .IN1(n10833), .IN2(n10834), .IN3(n10824), .IN4(n10825), 
        .QN(g34023) );
  NAND3X0 U10903 ( .IN1(n9354), .IN2(g2988), .IN3(n10145), .QN(n10824) );
  NAND3X0 U10904 ( .IN1(n9354), .IN2(g4552), .IN3(n10831), .QN(n10834) );
  NAND2X0 U10905 ( .IN1(n10835), .IN2(n9325), .QN(n10833) );
  NAND2X0 U10906 ( .IN1(n10836), .IN2(n9379), .QN(n10835) );
  NAND4X0 U10907 ( .IN1(n10145), .IN2(g4555), .IN3(g4558), .IN4(g4561), .QN(
        n10836) );
  NAND4X0 U10908 ( .IN1(n10837), .IN2(n9664), .IN3(n10838), .IN4(n10839), .QN(
        g34022) );
  NAND3X0 U10909 ( .IN1(n10840), .IN2(g2763), .IN3(n9342), .QN(n10839) );
  NAND2X0 U10910 ( .IN1(n9474), .IN2(g2759), .QN(n10838) );
  NAND2X0 U10911 ( .IN1(n10841), .IN2(n8337), .QN(n10837) );
  INVX0 U10912 ( .INP(n10840), .ZN(n10841) );
  NAND2X0 U10913 ( .IN1(n10842), .IN2(g2759), .QN(n10840) );
  NAND3X0 U10914 ( .IN1(n10843), .IN2(n10844), .IN3(n10845), .QN(g34021) );
  NAND2X0 U10915 ( .IN1(n9474), .IN2(g2648), .QN(n10845) );
  NAND2X0 U10916 ( .IN1(n10846), .IN2(n10847), .QN(n10844) );
  NAND2X0 U10917 ( .IN1(n10848), .IN2(g2567), .QN(n10843) );
  NAND2X0 U10918 ( .IN1(n10849), .IN2(n10850), .QN(g34020) );
  NAND2X0 U10919 ( .IN1(n10851), .IN2(g2629), .QN(n10850) );
  NAND2X0 U10920 ( .IN1(n10852), .IN2(n9379), .QN(n10851) );
  NAND2X0 U10921 ( .IN1(n10853), .IN2(g2643), .QN(n10852) );
  NAND2X0 U10922 ( .IN1(n10854), .IN2(n9379), .QN(n10849) );
  NAND2X0 U10923 ( .IN1(n10855), .IN2(n10856), .QN(n10854) );
  NAND2X0 U10924 ( .IN1(n10857), .IN2(n10858), .QN(n10856) );
  NAND2X0 U10925 ( .IN1(n10859), .IN2(n10860), .QN(n10858) );
  NAND2X0 U10926 ( .IN1(n8415), .IN2(n10861), .QN(n10860) );
  NAND2X0 U10927 ( .IN1(n10862), .IN2(g2643), .QN(n10855) );
  NAND2X0 U10928 ( .IN1(n10861), .IN2(n10863), .QN(n10862) );
  NAND2X0 U10929 ( .IN1(n10853), .IN2(g2555), .QN(n10863) );
  INVX0 U10930 ( .INP(n10857), .ZN(n10853) );
  NAND2X0 U10931 ( .IN1(n10864), .IN2(n10865), .QN(n10857) );
  NAND2X0 U10932 ( .IN1(n5755), .IN2(n10866), .QN(n10865) );
  NAND2X0 U10933 ( .IN1(n10867), .IN2(n10868), .QN(n10864) );
  NAND2X0 U10934 ( .IN1(n10869), .IN2(n10123), .QN(n10867) );
  NAND3X0 U10935 ( .IN1(n10870), .IN2(n10871), .IN3(n10872), .QN(g34019) );
  NAND2X0 U10936 ( .IN1(n9474), .IN2(g2571), .QN(n10872) );
  NAND3X0 U10937 ( .IN1(n10873), .IN2(n10861), .IN3(n10847), .QN(n10871) );
  INVX0 U10938 ( .INP(n10874), .ZN(n10847) );
  NAND2X0 U10939 ( .IN1(n10875), .IN2(g2583), .QN(n10870) );
  NAND2X0 U10940 ( .IN1(n10876), .IN2(n10877), .QN(n10875) );
  NAND2X0 U10941 ( .IN1(n10614), .IN2(n9378), .QN(n10877) );
  INVX0 U10942 ( .INP(n10873), .ZN(n10614) );
  INVX0 U10943 ( .INP(n10878), .ZN(n10876) );
  NAND3X0 U10944 ( .IN1(n10879), .IN2(n10880), .IN3(n10881), .QN(g34018) );
  INVX0 U10945 ( .INP(n10882), .ZN(n10881) );
  NOR2X0 U10946 ( .IN1(n10883), .IN2(n10874), .QN(n10882) );
  NAND3X0 U10947 ( .IN1(test_so61), .IN2(n10883), .IN3(n9342), .QN(n10880) );
  NAND2X0 U10948 ( .IN1(n10884), .IN2(n5351), .QN(n10883) );
  NAND2X0 U10949 ( .IN1(n9473), .IN2(g2583), .QN(n10879) );
  NAND3X0 U10950 ( .IN1(n10885), .IN2(n10886), .IN3(n10887), .QN(g34017) );
  INVX0 U10951 ( .INP(n10888), .ZN(n10887) );
  NOR2X0 U10952 ( .IN1(n10889), .IN2(n10874), .QN(n10888) );
  NAND3X0 U10953 ( .IN1(test_so66), .IN2(n10889), .IN3(n9342), .QN(n10886) );
  NAND2X0 U10954 ( .IN1(n10890), .IN2(g2629), .QN(n10889) );
  NAND2X0 U10955 ( .IN1(test_so61), .IN2(n9513), .QN(n10885) );
  NAND3X0 U10956 ( .IN1(n10891), .IN2(n10892), .IN3(n10893), .QN(g34016) );
  INVX0 U10957 ( .INP(n10894), .ZN(n10893) );
  NOR2X0 U10958 ( .IN1(n10895), .IN2(n10874), .QN(n10894) );
  NAND3X0 U10959 ( .IN1(n10895), .IN2(g2571), .IN3(n9342), .QN(n10892) );
  NAND2X0 U10960 ( .IN1(n10884), .IN2(n5521), .QN(n10895) );
  NAND2X0 U10961 ( .IN1(n9473), .IN2(g2563), .QN(n10891) );
  NAND3X0 U10962 ( .IN1(n10896), .IN2(n10897), .IN3(n10898), .QN(g34015) );
  INVX0 U10963 ( .INP(n10899), .ZN(n10898) );
  NOR2X0 U10964 ( .IN1(n10900), .IN2(n10874), .QN(n10899) );
  NAND3X0 U10965 ( .IN1(n10901), .IN2(n10902), .IN3(n9342), .QN(n10874) );
  NAND2X0 U10966 ( .IN1(n10866), .IN2(g1585), .QN(n10902) );
  INVX0 U10967 ( .INP(n10868), .ZN(n10866) );
  NAND3X0 U10968 ( .IN1(n10869), .IN2(n10123), .IN3(n10868), .QN(n10901) );
  NAND3X0 U10969 ( .IN1(n10900), .IN2(g2563), .IN3(n9342), .QN(n10897) );
  NAND2X0 U10970 ( .IN1(n10890), .IN2(n5524), .QN(n10900) );
  NAND2X0 U10971 ( .IN1(n9473), .IN2(g2567), .QN(n10896) );
  NAND3X0 U10972 ( .IN1(n10903), .IN2(n10904), .IN3(n10905), .QN(g34014) );
  NAND2X0 U10973 ( .IN1(n9473), .IN2(g2514), .QN(n10905) );
  NAND2X0 U10974 ( .IN1(n10906), .IN2(n10907), .QN(n10904) );
  NAND2X0 U10975 ( .IN1(n10908), .IN2(g2433), .QN(n10903) );
  NAND2X0 U10976 ( .IN1(n10909), .IN2(n10910), .QN(g34013) );
  NAND2X0 U10977 ( .IN1(n10911), .IN2(g2495), .QN(n10910) );
  NAND2X0 U10978 ( .IN1(n10912), .IN2(n9378), .QN(n10911) );
  NAND2X0 U10979 ( .IN1(n10913), .IN2(g2509), .QN(n10912) );
  NAND2X0 U10980 ( .IN1(n10914), .IN2(n9378), .QN(n10909) );
  NAND2X0 U10981 ( .IN1(n10915), .IN2(n10916), .QN(n10914) );
  NAND2X0 U10982 ( .IN1(n10917), .IN2(n10918), .QN(n10916) );
  NAND2X0 U10983 ( .IN1(n10919), .IN2(n10920), .QN(n10918) );
  NAND2X0 U10984 ( .IN1(n8414), .IN2(n10921), .QN(n10920) );
  NAND2X0 U10985 ( .IN1(n10922), .IN2(g2509), .QN(n10915) );
  NAND2X0 U10986 ( .IN1(n10921), .IN2(n10923), .QN(n10922) );
  NAND2X0 U10987 ( .IN1(test_so79), .IN2(n10913), .QN(n10923) );
  INVX0 U10988 ( .INP(n10917), .ZN(n10913) );
  NAND2X0 U10989 ( .IN1(n10924), .IN2(n10925), .QN(n10917) );
  NAND2X0 U10990 ( .IN1(n10926), .IN2(g1589), .QN(n10925) );
  NAND2X0 U10991 ( .IN1(n10927), .IN2(n10928), .QN(n10924) );
  NAND2X0 U10992 ( .IN1(n10869), .IN2(n10058), .QN(n10927) );
  NAND3X0 U10993 ( .IN1(n10929), .IN2(n10930), .IN3(n10931), .QN(g34012) );
  NAND2X0 U10994 ( .IN1(n9473), .IN2(g2437), .QN(n10931) );
  NAND3X0 U10995 ( .IN1(n10932), .IN2(n10921), .IN3(n10907), .QN(n10930) );
  INVX0 U10996 ( .INP(n10933), .ZN(n10907) );
  NAND2X0 U10997 ( .IN1(n10934), .IN2(g2449), .QN(n10929) );
  NAND2X0 U10998 ( .IN1(n10935), .IN2(n10936), .QN(n10934) );
  NAND2X0 U10999 ( .IN1(n10616), .IN2(n9378), .QN(n10936) );
  INVX0 U11000 ( .INP(n10932), .ZN(n10616) );
  INVX0 U11001 ( .INP(n10937), .ZN(n10935) );
  NAND3X0 U11002 ( .IN1(n10938), .IN2(n10939), .IN3(n10940), .QN(g34011) );
  INVX0 U11003 ( .INP(n10941), .ZN(n10940) );
  NOR2X0 U11004 ( .IN1(n10942), .IN2(n10933), .QN(n10941) );
  NAND3X0 U11005 ( .IN1(n10942), .IN2(n9274), .IN3(n9343), .QN(n10939) );
  NAND2X0 U11006 ( .IN1(n10943), .IN2(n8860), .QN(n10942) );
  NAND2X0 U11007 ( .IN1(n9473), .IN2(g2449), .QN(n10938) );
  NAND3X0 U11008 ( .IN1(n10944), .IN2(n10945), .IN3(n10946), .QN(g34010) );
  INVX0 U11009 ( .INP(n10947), .ZN(n10946) );
  NOR2X0 U11010 ( .IN1(n10948), .IN2(n10933), .QN(n10947) );
  NAND3X0 U11011 ( .IN1(n10948), .IN2(g2441), .IN3(n9343), .QN(n10945) );
  NAND2X0 U11012 ( .IN1(n10949), .IN2(g2495), .QN(n10948) );
  NAND2X0 U11013 ( .IN1(n9473), .IN2(n9274), .QN(n10944) );
  NAND3X0 U11014 ( .IN1(n10950), .IN2(n10951), .IN3(n10952), .QN(g34009) );
  INVX0 U11015 ( .INP(n10953), .ZN(n10952) );
  NOR2X0 U11016 ( .IN1(n10954), .IN2(n10933), .QN(n10953) );
  NAND3X0 U11017 ( .IN1(n10954), .IN2(g2437), .IN3(n9343), .QN(n10951) );
  NAND2X0 U11018 ( .IN1(n10943), .IN2(n5522), .QN(n10954) );
  NAND2X0 U11019 ( .IN1(n9472), .IN2(g2429), .QN(n10950) );
  NAND3X0 U11020 ( .IN1(n10955), .IN2(n10956), .IN3(n10957), .QN(g34008) );
  INVX0 U11021 ( .INP(n10958), .ZN(n10957) );
  NOR2X0 U11022 ( .IN1(n10959), .IN2(n10933), .QN(n10958) );
  NAND3X0 U11023 ( .IN1(n10960), .IN2(n10961), .IN3(n9343), .QN(n10933) );
  NAND3X0 U11024 ( .IN1(n10869), .IN2(n10058), .IN3(n10928), .QN(n10961) );
  NAND2X0 U11025 ( .IN1(n5757), .IN2(n10926), .QN(n10960) );
  INVX0 U11026 ( .INP(n10928), .ZN(n10926) );
  NAND3X0 U11027 ( .IN1(n10959), .IN2(g2429), .IN3(n9343), .QN(n10956) );
  NAND2X0 U11028 ( .IN1(n10949), .IN2(n5523), .QN(n10959) );
  NAND2X0 U11029 ( .IN1(n9472), .IN2(g2433), .QN(n10955) );
  NAND3X0 U11030 ( .IN1(n10962), .IN2(n10963), .IN3(n10964), .QN(g34007) );
  NAND2X0 U11031 ( .IN1(n9472), .IN2(g2380), .QN(n10964) );
  NAND2X0 U11032 ( .IN1(n10965), .IN2(n10966), .QN(n10963) );
  NAND2X0 U11033 ( .IN1(g2299), .IN2(n10967), .QN(n10962) );
  NAND2X0 U11034 ( .IN1(n10968), .IN2(n10969), .QN(g34006) );
  NAND2X0 U11035 ( .IN1(n10970), .IN2(g2361), .QN(n10969) );
  NAND2X0 U11036 ( .IN1(n10971), .IN2(n9378), .QN(n10970) );
  NAND2X0 U11037 ( .IN1(n10972), .IN2(g2375), .QN(n10971) );
  NAND2X0 U11038 ( .IN1(n10973), .IN2(n9377), .QN(n10968) );
  NAND2X0 U11039 ( .IN1(n10974), .IN2(n10975), .QN(n10973) );
  NAND2X0 U11040 ( .IN1(n10976), .IN2(n10977), .QN(n10975) );
  NAND2X0 U11041 ( .IN1(n10978), .IN2(n10979), .QN(n10977) );
  NAND2X0 U11042 ( .IN1(n8416), .IN2(n10980), .QN(n10979) );
  NAND2X0 U11043 ( .IN1(n10981), .IN2(g2375), .QN(n10974) );
  NAND2X0 U11044 ( .IN1(n10980), .IN2(n10982), .QN(n10981) );
  NAND2X0 U11045 ( .IN1(n10972), .IN2(g2287), .QN(n10982) );
  INVX0 U11046 ( .INP(n10976), .ZN(n10972) );
  NAND2X0 U11047 ( .IN1(n10983), .IN2(n10984), .QN(n10976) );
  NAND2X0 U11048 ( .IN1(n10985), .IN2(n5755), .QN(n10984) );
  NAND2X0 U11049 ( .IN1(n10986), .IN2(n10987), .QN(n10983) );
  NAND3X0 U11050 ( .IN1(n10988), .IN2(n10989), .IN3(n10990), .QN(g34005) );
  NAND2X0 U11051 ( .IN1(n10991), .IN2(n10965), .QN(n10990) );
  NAND3X0 U11052 ( .IN1(n10992), .IN2(g2315), .IN3(n9343), .QN(n10989) );
  INVX0 U11053 ( .INP(n10991), .ZN(n10992) );
  NOR2X0 U11054 ( .IN1(n10993), .IN2(n5537), .QN(n10991) );
  NAND2X0 U11055 ( .IN1(n9472), .IN2(g2303), .QN(n10988) );
  NAND3X0 U11056 ( .IN1(n10994), .IN2(n10995), .IN3(n10996), .QN(g34004) );
  NAND2X0 U11057 ( .IN1(n9472), .IN2(g2315), .QN(n10996) );
  NAND3X0 U11058 ( .IN1(n10965), .IN2(n5353), .IN3(n10997), .QN(n10995) );
  INVX0 U11059 ( .INP(n10998), .ZN(n10994) );
  NOR2X0 U11060 ( .IN1(n10999), .IN2(n15964), .QN(n10998) );
  NOR2X0 U11061 ( .IN1(n11000), .IN2(n11001), .QN(n10999) );
  NOR2X0 U11062 ( .IN1(n10997), .IN2(n9389), .QN(n11001) );
  NAND3X0 U11063 ( .IN1(n11002), .IN2(n11003), .IN3(n11004), .QN(g34003) );
  NAND2X0 U11064 ( .IN1(n11005), .IN2(n10965), .QN(n11004) );
  INVX0 U11065 ( .INP(n11006), .ZN(n11005) );
  NAND3X0 U11066 ( .IN1(n11006), .IN2(g2307), .IN3(n9344), .QN(n11003) );
  NAND3X0 U11067 ( .IN1(g2287), .IN2(g2361), .IN3(n10980), .QN(n11006) );
  NAND2X0 U11068 ( .IN1(n9472), .IN2(n9314), .QN(n11002) );
  NAND3X0 U11069 ( .IN1(n11007), .IN2(n11008), .IN3(n11009), .QN(g34002) );
  NAND2X0 U11070 ( .IN1(n11010), .IN2(n10965), .QN(n11009) );
  INVX0 U11071 ( .INP(n11011), .ZN(n11010) );
  NAND3X0 U11072 ( .IN1(n11011), .IN2(g2303), .IN3(n9344), .QN(n11008) );
  NAND2X0 U11073 ( .IN1(n10997), .IN2(n5537), .QN(n11011) );
  NAND2X0 U11074 ( .IN1(n9472), .IN2(g2295), .QN(n11007) );
  NAND3X0 U11075 ( .IN1(n11012), .IN2(n11013), .IN3(n11014), .QN(g34001) );
  NAND2X0 U11076 ( .IN1(n11015), .IN2(n10965), .QN(n11014) );
  NOR3X0 U11077 ( .IN1(n11016), .IN2(n11017), .IN3(n9383), .QN(n10965) );
  NOR2X0 U11078 ( .IN1(n10987), .IN2(n5757), .QN(n11017) );
  NOR2X0 U11079 ( .IN1(n10986), .IN2(n10985), .QN(n11016) );
  INVX0 U11080 ( .INP(n10987), .ZN(n10985) );
  NAND2X0 U11081 ( .IN1(n10869), .IN2(n10013), .QN(n10986) );
  NAND3X0 U11082 ( .IN1(n11018), .IN2(g2295), .IN3(n9344), .QN(n11013) );
  INVX0 U11083 ( .INP(n11015), .ZN(n11018) );
  NOR2X0 U11084 ( .IN1(n10993), .IN2(n5353), .QN(n11015) );
  NAND2X0 U11085 ( .IN1(g2299), .IN2(n9516), .QN(n11012) );
  NAND3X0 U11086 ( .IN1(n11019), .IN2(n11020), .IN3(n11021), .QN(g34000) );
  NAND2X0 U11087 ( .IN1(n9471), .IN2(g2246), .QN(n11021) );
  NAND2X0 U11088 ( .IN1(n11022), .IN2(n11023), .QN(n11020) );
  NAND2X0 U11089 ( .IN1(n11024), .IN2(g2165), .QN(n11019) );
  NAND2X0 U11090 ( .IN1(n11025), .IN2(n11026), .QN(g33999) );
  NAND2X0 U11091 ( .IN1(n11027), .IN2(g2227), .QN(n11026) );
  NAND2X0 U11092 ( .IN1(n11028), .IN2(n9377), .QN(n11027) );
  NAND2X0 U11093 ( .IN1(n11029), .IN2(g2241), .QN(n11028) );
  NAND2X0 U11094 ( .IN1(n11030), .IN2(n9377), .QN(n11025) );
  NAND2X0 U11095 ( .IN1(n11031), .IN2(n11032), .QN(n11030) );
  NAND2X0 U11096 ( .IN1(n11033), .IN2(n11034), .QN(n11032) );
  NAND2X0 U11097 ( .IN1(n11035), .IN2(n11036), .QN(n11034) );
  NAND2X0 U11098 ( .IN1(n8418), .IN2(n11037), .QN(n11036) );
  NAND2X0 U11099 ( .IN1(n11038), .IN2(g2241), .QN(n11031) );
  NAND2X0 U11100 ( .IN1(n11037), .IN2(n11039), .QN(n11038) );
  NAND2X0 U11101 ( .IN1(n11029), .IN2(g2153), .QN(n11039) );
  INVX0 U11102 ( .INP(n11033), .ZN(n11029) );
  NAND2X0 U11103 ( .IN1(n11040), .IN2(n11041), .QN(n11033) );
  NAND2X0 U11104 ( .IN1(n11042), .IN2(g1589), .QN(n11041) );
  NAND2X0 U11105 ( .IN1(n11043), .IN2(n11044), .QN(n11040) );
  NAND3X0 U11106 ( .IN1(n11045), .IN2(n11046), .IN3(n11047), .QN(g33998) );
  NAND2X0 U11107 ( .IN1(n11048), .IN2(n11022), .QN(n11047) );
  NAND3X0 U11108 ( .IN1(n11049), .IN2(g2181), .IN3(n9344), .QN(n11046) );
  INVX0 U11109 ( .INP(n11048), .ZN(n11049) );
  NOR2X0 U11110 ( .IN1(n11050), .IN2(n5538), .QN(n11048) );
  NAND2X0 U11111 ( .IN1(n9471), .IN2(g2169), .QN(n11045) );
  NAND3X0 U11112 ( .IN1(n11051), .IN2(n11052), .IN3(n11053), .QN(g33997) );
  NAND2X0 U11113 ( .IN1(n9471), .IN2(g2181), .QN(n11053) );
  NAND3X0 U11114 ( .IN1(n11022), .IN2(n5356), .IN3(n11054), .QN(n11052) );
  INVX0 U11115 ( .INP(n11055), .ZN(n11051) );
  NOR2X0 U11116 ( .IN1(n11056), .IN2(n15965), .QN(n11055) );
  NOR2X0 U11117 ( .IN1(n11057), .IN2(n11058), .QN(n11056) );
  NOR2X0 U11118 ( .IN1(n11054), .IN2(n9391), .QN(n11058) );
  NAND3X0 U11119 ( .IN1(n11059), .IN2(n11060), .IN3(n11061), .QN(g33996) );
  NAND2X0 U11120 ( .IN1(n11062), .IN2(n11022), .QN(n11061) );
  INVX0 U11121 ( .INP(n11063), .ZN(n11062) );
  NAND3X0 U11122 ( .IN1(n11063), .IN2(g2173), .IN3(n9344), .QN(n11060) );
  NAND3X0 U11123 ( .IN1(g2153), .IN2(g2227), .IN3(n11037), .QN(n11063) );
  NAND2X0 U11124 ( .IN1(n9471), .IN2(n9352), .QN(n11059) );
  NAND3X0 U11125 ( .IN1(n11064), .IN2(n11065), .IN3(n11066), .QN(g33995) );
  NAND2X0 U11126 ( .IN1(n11067), .IN2(n11022), .QN(n11066) );
  INVX0 U11127 ( .INP(n11068), .ZN(n11067) );
  NAND3X0 U11128 ( .IN1(n11068), .IN2(g2169), .IN3(n9344), .QN(n11065) );
  NAND2X0 U11129 ( .IN1(n11054), .IN2(n5538), .QN(n11068) );
  NAND2X0 U11130 ( .IN1(n9471), .IN2(g2161), .QN(n11064) );
  NAND3X0 U11131 ( .IN1(n11069), .IN2(n11070), .IN3(n11071), .QN(g33994) );
  NAND2X0 U11132 ( .IN1(n11072), .IN2(n11022), .QN(n11071) );
  NOR3X0 U11133 ( .IN1(n11073), .IN2(n11074), .IN3(n9383), .QN(n11022) );
  NOR2X0 U11134 ( .IN1(n11043), .IN2(n11042), .QN(n11074) );
  INVX0 U11135 ( .INP(n11044), .ZN(n11042) );
  NAND2X0 U11136 ( .IN1(n10869), .IN2(n9983), .QN(n11043) );
  NOR2X0 U11137 ( .IN1(n11075), .IN2(n5380), .QN(n10869) );
  INVX0 U11138 ( .INP(n11076), .ZN(n11075) );
  NOR2X0 U11139 ( .IN1(n11044), .IN2(g1585), .QN(n11073) );
  NAND3X0 U11140 ( .IN1(n11077), .IN2(g2161), .IN3(n9344), .QN(n11070) );
  INVX0 U11141 ( .INP(n11072), .ZN(n11077) );
  NOR2X0 U11142 ( .IN1(n11050), .IN2(n5356), .QN(n11072) );
  NAND2X0 U11143 ( .IN1(n9471), .IN2(g2165), .QN(n11069) );
  NAND3X0 U11144 ( .IN1(n11078), .IN2(n11079), .IN3(n11080), .QN(g33993) );
  NAND2X0 U11145 ( .IN1(n9471), .IN2(g2089), .QN(n11080) );
  NAND2X0 U11146 ( .IN1(n11081), .IN2(n11082), .QN(n11079) );
  NAND2X0 U11147 ( .IN1(n11083), .IN2(g2008), .QN(n11078) );
  NAND2X0 U11148 ( .IN1(n11084), .IN2(n11085), .QN(g33992) );
  NAND2X0 U11149 ( .IN1(n11086), .IN2(g2070), .QN(n11085) );
  NAND2X0 U11150 ( .IN1(n11087), .IN2(n9377), .QN(n11086) );
  NAND2X0 U11151 ( .IN1(n11088), .IN2(g2084), .QN(n11087) );
  NAND2X0 U11152 ( .IN1(n11089), .IN2(n9377), .QN(n11084) );
  NAND2X0 U11153 ( .IN1(n11090), .IN2(n11091), .QN(n11089) );
  NAND2X0 U11154 ( .IN1(n11092), .IN2(n11093), .QN(n11091) );
  NAND2X0 U11155 ( .IN1(n11094), .IN2(n11095), .QN(n11093) );
  NAND2X0 U11156 ( .IN1(n8413), .IN2(n11096), .QN(n11095) );
  NAND2X0 U11157 ( .IN1(n11097), .IN2(g2084), .QN(n11090) );
  NAND2X0 U11158 ( .IN1(n11096), .IN2(n11098), .QN(n11097) );
  NAND2X0 U11159 ( .IN1(n11088), .IN2(g1996), .QN(n11098) );
  INVX0 U11160 ( .INP(n11092), .ZN(n11088) );
  NAND2X0 U11161 ( .IN1(n11099), .IN2(n11100), .QN(n11092) );
  NAND2X0 U11162 ( .IN1(n5756), .IN2(n11101), .QN(n11100) );
  NAND2X0 U11163 ( .IN1(n11102), .IN2(n11103), .QN(n11099) );
  NAND3X0 U11164 ( .IN1(n11104), .IN2(n11105), .IN3(n11106), .QN(g33991) );
  NAND2X0 U11165 ( .IN1(n11107), .IN2(n11081), .QN(n11106) );
  NAND3X0 U11166 ( .IN1(n11108), .IN2(g2024), .IN3(n9345), .QN(n11105) );
  INVX0 U11167 ( .INP(n11107), .ZN(n11108) );
  NOR2X0 U11168 ( .IN1(n10618), .IN2(n11109), .QN(n11107) );
  NAND2X0 U11169 ( .IN1(n9470), .IN2(g2012), .QN(n11104) );
  NAND3X0 U11170 ( .IN1(n11110), .IN2(n11111), .IN3(n11112), .QN(g33990) );
  NAND2X0 U11171 ( .IN1(n11113), .IN2(n11081), .QN(n11112) );
  INVX0 U11172 ( .INP(n11114), .ZN(n11113) );
  NAND3X0 U11173 ( .IN1(n11114), .IN2(n9312), .IN3(n9344), .QN(n11111) );
  NAND2X0 U11174 ( .IN1(n11115), .IN2(n5355), .QN(n11114) );
  NAND2X0 U11175 ( .IN1(n9470), .IN2(g2024), .QN(n11110) );
  NAND3X0 U11176 ( .IN1(n11116), .IN2(n11117), .IN3(n11118), .QN(g33989) );
  NAND2X0 U11177 ( .IN1(n11119), .IN2(n11081), .QN(n11118) );
  INVX0 U11178 ( .INP(n11120), .ZN(n11119) );
  NAND3X0 U11179 ( .IN1(n11120), .IN2(g2016), .IN3(n9345), .QN(n11117) );
  NAND2X0 U11180 ( .IN1(n11121), .IN2(g2070), .QN(n11120) );
  NAND2X0 U11181 ( .IN1(n9470), .IN2(n9312), .QN(n11116) );
  NAND3X0 U11182 ( .IN1(n11122), .IN2(n11123), .IN3(n11124), .QN(g33988) );
  NAND2X0 U11183 ( .IN1(n11125), .IN2(n11081), .QN(n11124) );
  INVX0 U11184 ( .INP(n11126), .ZN(n11125) );
  NAND3X0 U11185 ( .IN1(n11126), .IN2(g2012), .IN3(n9345), .QN(n11123) );
  NAND2X0 U11186 ( .IN1(n11115), .IN2(n5535), .QN(n11126) );
  NAND2X0 U11187 ( .IN1(n9470), .IN2(g2004), .QN(n11122) );
  NAND3X0 U11188 ( .IN1(n11127), .IN2(n11128), .IN3(n11129), .QN(g33987) );
  NAND2X0 U11189 ( .IN1(n11130), .IN2(n11081), .QN(n11129) );
  NOR3X0 U11190 ( .IN1(n11131), .IN2(n11132), .IN3(n9383), .QN(n11081) );
  NOR2X0 U11191 ( .IN1(n11103), .IN2(n5526), .QN(n11132) );
  NOR2X0 U11192 ( .IN1(n11102), .IN2(n11101), .QN(n11131) );
  INVX0 U11193 ( .INP(n11103), .ZN(n11101) );
  NAND2X0 U11194 ( .IN1(n11133), .IN2(n10119), .QN(n11102) );
  INVX0 U11195 ( .INP(n11134), .ZN(n11130) );
  NAND3X0 U11196 ( .IN1(n11134), .IN2(g2004), .IN3(n9345), .QN(n11128) );
  NAND2X0 U11197 ( .IN1(n11121), .IN2(n5505), .QN(n11134) );
  NAND2X0 U11198 ( .IN1(n9470), .IN2(g2008), .QN(n11127) );
  NAND3X0 U11199 ( .IN1(n11135), .IN2(n11136), .IN3(n11137), .QN(g33986) );
  NAND2X0 U11200 ( .IN1(n9470), .IN2(g1955), .QN(n11137) );
  NAND2X0 U11201 ( .IN1(n11138), .IN2(n11139), .QN(n11136) );
  NAND2X0 U11202 ( .IN1(n11140), .IN2(g1874), .QN(n11135) );
  NAND2X0 U11203 ( .IN1(n11141), .IN2(n11142), .QN(g33985) );
  NAND2X0 U11204 ( .IN1(n11143), .IN2(g1936), .QN(n11142) );
  NAND2X0 U11205 ( .IN1(n11144), .IN2(n9377), .QN(n11143) );
  NAND2X0 U11206 ( .IN1(n11145), .IN2(g1950), .QN(n11144) );
  NAND2X0 U11207 ( .IN1(n11146), .IN2(n9376), .QN(n11141) );
  NAND2X0 U11208 ( .IN1(n11147), .IN2(n11148), .QN(n11146) );
  NAND2X0 U11209 ( .IN1(n11149), .IN2(n11150), .QN(n11148) );
  NAND2X0 U11210 ( .IN1(n11151), .IN2(n11152), .QN(n11150) );
  NAND2X0 U11211 ( .IN1(n8417), .IN2(n11153), .QN(n11152) );
  NAND2X0 U11212 ( .IN1(n11154), .IN2(g1950), .QN(n11147) );
  NAND2X0 U11213 ( .IN1(n11153), .IN2(n11155), .QN(n11154) );
  NAND2X0 U11214 ( .IN1(test_so8), .IN2(n11145), .QN(n11155) );
  INVX0 U11215 ( .INP(n11149), .ZN(n11145) );
  NAND2X0 U11216 ( .IN1(n11156), .IN2(n11157), .QN(n11149) );
  NAND2X0 U11217 ( .IN1(n11158), .IN2(g1246), .QN(n11157) );
  NAND2X0 U11218 ( .IN1(n11159), .IN2(n11160), .QN(n11156) );
  NAND3X0 U11219 ( .IN1(n11161), .IN2(n11162), .IN3(n11163), .QN(g33984) );
  NAND2X0 U11220 ( .IN1(n11164), .IN2(n11138), .QN(n11163) );
  NAND3X0 U11221 ( .IN1(n11165), .IN2(g1890), .IN3(n9345), .QN(n11162) );
  INVX0 U11222 ( .INP(n11164), .ZN(n11165) );
  NOR2X0 U11223 ( .IN1(n10622), .IN2(n11166), .QN(n11164) );
  NAND2X0 U11224 ( .IN1(n9470), .IN2(g1878), .QN(n11161) );
  NAND3X0 U11225 ( .IN1(n11167), .IN2(n11168), .IN3(n11169), .QN(g33983) );
  NAND2X0 U11226 ( .IN1(n11170), .IN2(n11138), .QN(n11169) );
  INVX0 U11227 ( .INP(n11171), .ZN(n11170) );
  NAND3X0 U11228 ( .IN1(n11171), .IN2(n9280), .IN3(n9345), .QN(n11168) );
  NAND2X0 U11229 ( .IN1(n11172), .IN2(n8861), .QN(n11171) );
  NAND2X0 U11230 ( .IN1(n9469), .IN2(g1890), .QN(n11167) );
  NAND3X0 U11231 ( .IN1(n11173), .IN2(n11174), .IN3(n11175), .QN(g33982) );
  NAND2X0 U11232 ( .IN1(n11176), .IN2(n11138), .QN(n11175) );
  INVX0 U11233 ( .INP(n11177), .ZN(n11176) );
  NAND3X0 U11234 ( .IN1(n11177), .IN2(g1882), .IN3(n9345), .QN(n11174) );
  NAND2X0 U11235 ( .IN1(n11178), .IN2(g1936), .QN(n11177) );
  NAND2X0 U11236 ( .IN1(n9469), .IN2(n9280), .QN(n11173) );
  NAND3X0 U11237 ( .IN1(n11179), .IN2(n11180), .IN3(n11181), .QN(g33981) );
  NAND2X0 U11238 ( .IN1(n11182), .IN2(n11138), .QN(n11181) );
  INVX0 U11239 ( .INP(n11183), .ZN(n11182) );
  NAND3X0 U11240 ( .IN1(n11183), .IN2(g1878), .IN3(n9345), .QN(n11180) );
  NAND2X0 U11241 ( .IN1(n11172), .IN2(n5534), .QN(n11183) );
  NAND2X0 U11242 ( .IN1(n9469), .IN2(g1870), .QN(n11179) );
  NAND3X0 U11243 ( .IN1(n11184), .IN2(n11185), .IN3(n11186), .QN(g33980) );
  NAND2X0 U11244 ( .IN1(n11187), .IN2(n11138), .QN(n11186) );
  NOR3X0 U11245 ( .IN1(n11188), .IN2(n11189), .IN3(n9383), .QN(n11138) );
  NOR2X0 U11246 ( .IN1(n11159), .IN2(n11158), .QN(n11189) );
  INVX0 U11247 ( .INP(n11160), .ZN(n11158) );
  NAND2X0 U11248 ( .IN1(n11133), .IN2(n10055), .QN(n11159) );
  NOR2X0 U11249 ( .IN1(g30332), .IN2(n11160), .QN(n11188) );
  INVX0 U11250 ( .INP(n11190), .ZN(n11187) );
  NAND3X0 U11251 ( .IN1(n11190), .IN2(g1870), .IN3(n9345), .QN(n11185) );
  NAND2X0 U11252 ( .IN1(n11178), .IN2(n5503), .QN(n11190) );
  NAND2X0 U11253 ( .IN1(n9469), .IN2(g1874), .QN(n11184) );
  NAND3X0 U11254 ( .IN1(n11191), .IN2(n11192), .IN3(n11193), .QN(g33979) );
  NAND2X0 U11255 ( .IN1(n9469), .IN2(g1821), .QN(n11193) );
  NAND2X0 U11256 ( .IN1(n11194), .IN2(n11195), .QN(n11192) );
  NAND2X0 U11257 ( .IN1(n11196), .IN2(g1740), .QN(n11191) );
  NAND2X0 U11258 ( .IN1(n11197), .IN2(n11198), .QN(g33978) );
  NAND2X0 U11259 ( .IN1(n11199), .IN2(g1802), .QN(n11198) );
  NAND2X0 U11260 ( .IN1(n11200), .IN2(n9376), .QN(n11199) );
  NAND2X0 U11261 ( .IN1(n11201), .IN2(g1816), .QN(n11200) );
  NAND2X0 U11262 ( .IN1(n11202), .IN2(n9375), .QN(n11197) );
  NAND2X0 U11263 ( .IN1(n11203), .IN2(n11204), .QN(n11202) );
  NAND2X0 U11264 ( .IN1(n11205), .IN2(n11206), .QN(n11204) );
  NAND2X0 U11265 ( .IN1(n11207), .IN2(n11208), .QN(n11206) );
  NAND2X0 U11266 ( .IN1(n8355), .IN2(n11209), .QN(n11208) );
  NAND2X0 U11267 ( .IN1(n11210), .IN2(g1816), .QN(n11203) );
  NAND2X0 U11268 ( .IN1(n11209), .IN2(n11211), .QN(n11210) );
  NAND2X0 U11269 ( .IN1(n11201), .IN2(g1728), .QN(n11211) );
  INVX0 U11270 ( .INP(n11205), .ZN(n11201) );
  NAND2X0 U11271 ( .IN1(n11212), .IN2(n11213), .QN(n11205) );
  NAND2X0 U11272 ( .IN1(n11214), .IN2(n5756), .QN(n11213) );
  NAND2X0 U11273 ( .IN1(n11215), .IN2(n11216), .QN(n11212) );
  NAND3X0 U11274 ( .IN1(n11217), .IN2(n11218), .IN3(n11219), .QN(g33977) );
  NAND2X0 U11275 ( .IN1(n11220), .IN2(n11194), .QN(n11219) );
  NAND3X0 U11276 ( .IN1(n11221), .IN2(g1756), .IN3(n9345), .QN(n11218) );
  INVX0 U11277 ( .INP(n11220), .ZN(n11221) );
  NOR2X0 U11278 ( .IN1(n11222), .IN2(n5536), .QN(n11220) );
  NAND2X0 U11279 ( .IN1(n9469), .IN2(g1744), .QN(n11217) );
  NAND3X0 U11280 ( .IN1(n11223), .IN2(n11224), .IN3(n11225), .QN(g33976) );
  NAND2X0 U11281 ( .IN1(n9469), .IN2(g1756), .QN(n11225) );
  NAND3X0 U11282 ( .IN1(n11194), .IN2(n5352), .IN3(n11226), .QN(n11224) );
  INVX0 U11283 ( .INP(n11227), .ZN(n11223) );
  NOR2X0 U11284 ( .IN1(n11228), .IN2(n5797), .QN(n11227) );
  NOR2X0 U11285 ( .IN1(n11229), .IN2(n11230), .QN(n11228) );
  NOR2X0 U11286 ( .IN1(n11226), .IN2(n9393), .QN(n11230) );
  NAND3X0 U11287 ( .IN1(n11231), .IN2(n11232), .IN3(n11233), .QN(g33975) );
  NAND2X0 U11288 ( .IN1(n11234), .IN2(n11194), .QN(n11233) );
  INVX0 U11289 ( .INP(n11235), .ZN(n11234) );
  NAND3X0 U11290 ( .IN1(n11235), .IN2(g1748), .IN3(n9346), .QN(n11232) );
  NAND3X0 U11291 ( .IN1(g1728), .IN2(g1802), .IN3(n11209), .QN(n11235) );
  NAND2X0 U11292 ( .IN1(n9468), .IN2(g1752), .QN(n11231) );
  NAND3X0 U11293 ( .IN1(n11236), .IN2(n11237), .IN3(n11238), .QN(g33974) );
  NAND2X0 U11294 ( .IN1(n11239), .IN2(n11194), .QN(n11238) );
  INVX0 U11295 ( .INP(n11240), .ZN(n11239) );
  NAND3X0 U11296 ( .IN1(n11240), .IN2(g1744), .IN3(n9346), .QN(n11237) );
  NAND2X0 U11297 ( .IN1(n11226), .IN2(n5536), .QN(n11240) );
  NAND2X0 U11298 ( .IN1(n9468), .IN2(g1736), .QN(n11236) );
  NAND3X0 U11299 ( .IN1(n11241), .IN2(n11242), .IN3(n11243), .QN(g33973) );
  NAND2X0 U11300 ( .IN1(n11244), .IN2(n11194), .QN(n11243) );
  NOR3X0 U11301 ( .IN1(n11245), .IN2(n11246), .IN3(n9384), .QN(n11194) );
  NOR2X0 U11302 ( .IN1(n11216), .IN2(n5526), .QN(n11246) );
  NOR2X0 U11303 ( .IN1(n11215), .IN2(n11214), .QN(n11245) );
  INVX0 U11304 ( .INP(n11216), .ZN(n11214) );
  NAND2X0 U11305 ( .IN1(n11133), .IN2(n10014), .QN(n11215) );
  NAND3X0 U11306 ( .IN1(n11247), .IN2(g1736), .IN3(n9346), .QN(n11242) );
  INVX0 U11307 ( .INP(n11244), .ZN(n11247) );
  NOR2X0 U11308 ( .IN1(n11222), .IN2(n5352), .QN(n11244) );
  NAND2X0 U11309 ( .IN1(n9468), .IN2(g1740), .QN(n11241) );
  NAND3X0 U11310 ( .IN1(n11248), .IN2(n11249), .IN3(n11250), .QN(g33972) );
  NAND2X0 U11311 ( .IN1(n9468), .IN2(g1687), .QN(n11250) );
  NAND2X0 U11312 ( .IN1(n11251), .IN2(n11252), .QN(n11249) );
  NAND2X0 U11313 ( .IN1(n11253), .IN2(g1604), .QN(n11248) );
  NAND2X0 U11314 ( .IN1(n11254), .IN2(n11255), .QN(g33971) );
  NAND2X0 U11315 ( .IN1(n11256), .IN2(g1668), .QN(n11255) );
  NAND2X0 U11316 ( .IN1(n11257), .IN2(n9375), .QN(n11256) );
  NAND2X0 U11317 ( .IN1(n11258), .IN2(g1682), .QN(n11257) );
  NAND2X0 U11318 ( .IN1(n11259), .IN2(n9375), .QN(n11254) );
  NAND2X0 U11319 ( .IN1(n11260), .IN2(n11261), .QN(n11259) );
  NAND2X0 U11320 ( .IN1(n11262), .IN2(n11263), .QN(n11261) );
  NAND2X0 U11321 ( .IN1(n11264), .IN2(n11265), .QN(n11263) );
  NAND2X0 U11322 ( .IN1(n8419), .IN2(n11266), .QN(n11265) );
  NAND2X0 U11323 ( .IN1(n11267), .IN2(g1682), .QN(n11260) );
  NAND2X0 U11324 ( .IN1(n11266), .IN2(n11268), .QN(n11267) );
  NAND2X0 U11325 ( .IN1(n11258), .IN2(g1592), .QN(n11268) );
  INVX0 U11326 ( .INP(n11262), .ZN(n11258) );
  NAND2X0 U11327 ( .IN1(n11269), .IN2(n11270), .QN(n11262) );
  NAND2X0 U11328 ( .IN1(n11271), .IN2(g1246), .QN(n11270) );
  NAND2X0 U11329 ( .IN1(n11272), .IN2(n11273), .QN(n11269) );
  NAND2X0 U11330 ( .IN1(n11133), .IN2(n9984), .QN(n11272) );
  NAND3X0 U11331 ( .IN1(n11274), .IN2(n11275), .IN3(n11276), .QN(g33970) );
  NAND2X0 U11332 ( .IN1(n11277), .IN2(n11252), .QN(n11276) );
  INVX0 U11333 ( .INP(n11278), .ZN(n11277) );
  NAND3X0 U11334 ( .IN1(n11278), .IN2(g1620), .IN3(n9346), .QN(n11275) );
  NAND2X0 U11335 ( .IN1(g25259), .IN2(n11266), .QN(n11278) );
  NAND2X0 U11336 ( .IN1(n9468), .IN2(g1608), .QN(n11274) );
  NAND3X0 U11337 ( .IN1(n11279), .IN2(n11280), .IN3(n11281), .QN(g33969) );
  NAND2X0 U11338 ( .IN1(n11282), .IN2(n11252), .QN(n11281) );
  INVX0 U11339 ( .INP(n11283), .ZN(n11282) );
  NAND3X0 U11340 ( .IN1(n11283), .IN2(n9303), .IN3(n9346), .QN(n11280) );
  NAND2X0 U11341 ( .IN1(n11284), .IN2(n5362), .QN(n11283) );
  NAND2X0 U11342 ( .IN1(n9468), .IN2(g1620), .QN(n11279) );
  NAND3X0 U11343 ( .IN1(n11285), .IN2(n11286), .IN3(n11287), .QN(g33968) );
  NAND2X0 U11344 ( .IN1(n11288), .IN2(n11252), .QN(n11287) );
  INVX0 U11345 ( .INP(n11289), .ZN(n11288) );
  NAND3X0 U11346 ( .IN1(n11289), .IN2(g1612), .IN3(n9346), .QN(n11286) );
  NAND2X0 U11347 ( .IN1(n11290), .IN2(g1668), .QN(n11289) );
  NAND2X0 U11348 ( .IN1(n9468), .IN2(n9303), .QN(n11285) );
  NAND3X0 U11349 ( .IN1(n11291), .IN2(n11292), .IN3(n11293), .QN(g33967) );
  NAND2X0 U11350 ( .IN1(n11294), .IN2(n11252), .QN(n11293) );
  INVX0 U11351 ( .INP(n11295), .ZN(n11294) );
  NAND3X0 U11352 ( .IN1(n11295), .IN2(g1608), .IN3(n9346), .QN(n11292) );
  NAND2X0 U11353 ( .IN1(n11284), .IN2(n5598), .QN(n11295) );
  NAND2X0 U11354 ( .IN1(n9467), .IN2(g1600), .QN(n11291) );
  NAND3X0 U11355 ( .IN1(n11296), .IN2(n11297), .IN3(n11298), .QN(g33966) );
  NAND2X0 U11356 ( .IN1(n11299), .IN2(n11252), .QN(n11298) );
  INVX0 U11357 ( .INP(n11300), .ZN(n11252) );
  NAND3X0 U11358 ( .IN1(n11301), .IN2(n11302), .IN3(n9346), .QN(n11300) );
  NAND3X0 U11359 ( .IN1(n11133), .IN2(n9984), .IN3(n11273), .QN(n11302) );
  NOR2X0 U11360 ( .IN1(n11303), .IN2(n5380), .QN(n11133) );
  INVX0 U11361 ( .INP(n11304), .ZN(n11303) );
  NAND2X0 U11362 ( .IN1(n11271), .IN2(n5526), .QN(n11301) );
  INVX0 U11363 ( .INP(n11273), .ZN(n11271) );
  INVX0 U11364 ( .INP(n11305), .ZN(n11299) );
  NAND3X0 U11365 ( .IN1(n11305), .IN2(g1600), .IN3(n9346), .QN(n11297) );
  NAND2X0 U11366 ( .IN1(n11290), .IN2(n5549), .QN(n11305) );
  NAND2X0 U11367 ( .IN1(n9467), .IN2(g1604), .QN(n11296) );
  NAND3X0 U11368 ( .IN1(n11306), .IN2(n11307), .IN3(n11308), .QN(g33965) );
  NAND2X0 U11369 ( .IN1(n9467), .IN2(g763), .QN(n11308) );
  NAND3X0 U11370 ( .IN1(n2404), .IN2(n11309), .IN3(g767), .QN(n11307) );
  INVX0 U11371 ( .INP(n2704), .ZN(n11309) );
  NAND2X0 U11372 ( .IN1(n2704), .IN2(n5333), .QN(n11306) );
  NAND3X0 U11373 ( .IN1(n11310), .IN2(n11311), .IN3(n11312), .QN(g33964) );
  NAND2X0 U11374 ( .IN1(n9467), .IN2(g595), .QN(n11312) );
  NAND3X0 U11375 ( .IN1(n2421), .IN2(n11313), .IN3(g599), .QN(n11311) );
  INVX0 U11376 ( .INP(n2706), .ZN(n11313) );
  NAND2X0 U11377 ( .IN1(n2706), .IN2(n5550), .QN(n11310) );
  NAND2X0 U11378 ( .IN1(n11314), .IN2(n11315), .QN(g33963) );
  NAND2X0 U11379 ( .IN1(n9467), .IN2(g29215), .QN(n11315) );
  NAND3X0 U11380 ( .IN1(n11316), .IN2(n11317), .IN3(n9346), .QN(n11314) );
  NAND3X0 U11381 ( .IN1(n11318), .IN2(n9794), .IN3(n11319), .QN(n11317) );
  NAND2X0 U11382 ( .IN1(g72), .IN2(g262), .QN(n11319) );
  NAND2X0 U11383 ( .IN1(n11320), .IN2(g269), .QN(n11318) );
  NAND2X0 U11384 ( .IN1(g73), .IN2(n11321), .QN(n11316) );
  NAND2X0 U11385 ( .IN1(n11320), .IN2(g255), .QN(n11321) );
  NAND2X0 U11386 ( .IN1(n11322), .IN2(n11323), .QN(g33962) );
  NAND2X0 U11387 ( .IN1(n9467), .IN2(g479), .QN(n11323) );
  NAND3X0 U11388 ( .IN1(n11324), .IN2(n11325), .IN3(n9346), .QN(n11322) );
  NAND3X0 U11389 ( .IN1(n11326), .IN2(n9794), .IN3(n11327), .QN(n11325) );
  NAND2X0 U11390 ( .IN1(g72), .IN2(g239), .QN(n11327) );
  NAND2X0 U11391 ( .IN1(n11320), .IN2(g246), .QN(n11326) );
  NAND2X0 U11392 ( .IN1(g73), .IN2(n11328), .QN(n11324) );
  NAND2X0 U11393 ( .IN1(n11329), .IN2(n11330), .QN(n11328) );
  NAND2X0 U11394 ( .IN1(n5597), .IN2(g72), .QN(n11330) );
  NAND2X0 U11395 ( .IN1(n8589), .IN2(n9791), .QN(n11329) );
  NAND3X0 U11396 ( .IN1(n11331), .IN2(n11332), .IN3(n11333), .QN(g33961) );
  NAND2X0 U11397 ( .IN1(n9467), .IN2(g294), .QN(n11333) );
  NAND3X0 U11398 ( .IN1(n10734), .IN2(n11334), .IN3(g298), .QN(n11332) );
  INVX0 U11399 ( .INP(n2989), .ZN(n11334) );
  NAND2X0 U11400 ( .IN1(n2989), .IN2(n5675), .QN(n11331) );
  NAND3X0 U11401 ( .IN1(n11335), .IN2(n11336), .IN3(n11337), .QN(g33960) );
  NAND2X0 U11402 ( .IN1(n9466), .IN2(g153), .QN(n11337) );
  NAND3X0 U11403 ( .IN1(n10739), .IN2(n11338), .IN3(g157), .QN(n11336) );
  INVX0 U11404 ( .INP(n2991), .ZN(n11338) );
  NAND2X0 U11405 ( .IN1(n2991), .IN2(n5678), .QN(n11335) );
  NAND4X0 U11406 ( .IN1(n2668), .IN2(n9750), .IN3(g8403), .IN4(g8283), .QN(
        g33935) );
  INVX0 U11407 ( .INP(g34649), .ZN(n9750) );
  NAND4X0 U11408 ( .IN1(n11339), .IN2(n11340), .IN3(n11341), .IN4(n11342), 
        .QN(g34649) );
  NAND2X0 U11409 ( .IN1(n9756), .IN2(g4888), .QN(n11342) );
  NAND2X0 U11410 ( .IN1(n9757), .IN2(g4955), .QN(n11341) );
  NAND2X0 U11411 ( .IN1(n9758), .IN2(g4944), .QN(n11340) );
  NAND2X0 U11412 ( .IN1(n9759), .IN2(g4933), .QN(n11339) );
  NAND3X0 U11413 ( .IN1(n2668), .IN2(g4507), .IN3(n5541), .QN(g33874) );
  NAND4X0 U11414 ( .IN1(n9661), .IN2(n10603), .IN3(n9771), .IN4(n9772), .QN(
        g33659) );
  NAND2X0 U11415 ( .IN1(n11343), .IN2(n11344), .QN(n9772) );
  NAND2X0 U11416 ( .IN1(n8593), .IN2(n9794), .QN(n11344) );
  NAND2X0 U11417 ( .IN1(g73), .IN2(g4104), .QN(n11343) );
  NAND2X0 U11418 ( .IN1(n11345), .IN2(n11346), .QN(n9771) );
  NAND2X0 U11419 ( .IN1(g72), .IN2(g4108), .QN(n11346) );
  NAND2X0 U11420 ( .IN1(n5715), .IN2(n9791), .QN(n11345) );
  INVX0 U11421 ( .INP(n10599), .ZN(n10603) );
  NAND2X0 U11422 ( .IN1(g113), .IN2(n2668), .QN(n10599) );
  INVX0 U11423 ( .INP(n11347), .ZN(n9661) );
  NAND2X0 U11424 ( .IN1(n11348), .IN2(n11349), .QN(n11347) );
  NAND2X0 U11425 ( .IN1(n5350), .IN2(n11350), .QN(n11349) );
  NAND3X0 U11426 ( .IN1(n11351), .IN2(n11352), .IN3(n11353), .QN(n11350) );
  NAND2X0 U11427 ( .IN1(n11354), .IN2(n11355), .QN(n11353) );
  NAND3X0 U11428 ( .IN1(n11356), .IN2(n11357), .IN3(g4093), .QN(n11352) );
  NAND2X0 U11429 ( .IN1(n5480), .IN2(n11358), .QN(n11357) );
  NAND2X0 U11430 ( .IN1(n11359), .IN2(g4087), .QN(n11356) );
  NAND2X0 U11431 ( .IN1(g32975), .IN2(n11360), .QN(n11351) );
  NAND2X0 U11432 ( .IN1(n11361), .IN2(g4098), .QN(n11348) );
  NAND3X0 U11433 ( .IN1(n11362), .IN2(n11363), .IN3(n11364), .QN(n11361) );
  NAND2X0 U11434 ( .IN1(n11365), .IN2(n11355), .QN(n11364) );
  NAND3X0 U11435 ( .IN1(n11366), .IN2(n11367), .IN3(g4093), .QN(n11363) );
  NAND2X0 U11436 ( .IN1(n5480), .IN2(n11368), .QN(n11367) );
  NAND2X0 U11437 ( .IN1(n11369), .IN2(g4087), .QN(n11366) );
  NAND2X0 U11438 ( .IN1(n11370), .IN2(n11360), .QN(n11362) );
  NAND4X0 U11439 ( .IN1(n2668), .IN2(n9717), .IN3(g8353), .IN4(g8235), .QN(
        g33636) );
  INVX0 U11440 ( .INP(g34657), .ZN(n9717) );
  NAND4X0 U11441 ( .IN1(n11371), .IN2(n11372), .IN3(n11373), .IN4(n11374), 
        .QN(g34657) );
  NAND2X0 U11442 ( .IN1(n9723), .IN2(g4754), .QN(n11374) );
  NAND2X0 U11443 ( .IN1(n9724), .IN2(g4743), .QN(n11373) );
  NAND2X0 U11444 ( .IN1(n9725), .IN2(g4765), .QN(n11372) );
  NAND2X0 U11445 ( .IN1(n9726), .IN2(g4698), .QN(n11371) );
  NAND2X0 U11446 ( .IN1(n11375), .IN2(n11376), .QN(n2668) );
  NAND2X0 U11447 ( .IN1(g99), .IN2(g37), .QN(n11376) );
  NAND3X0 U11448 ( .IN1(n11377), .IN2(n11378), .IN3(n11379), .QN(g33627) );
  NAND3X0 U11449 ( .IN1(n11380), .IN2(n11381), .IN3(n9685), .QN(n11379) );
  NAND2X0 U11450 ( .IN1(n9466), .IN2(g6741), .QN(n11378) );
  NAND2X0 U11451 ( .IN1(n11382), .IN2(n9375), .QN(n11377) );
  NAND2X0 U11452 ( .IN1(n11383), .IN2(n11384), .QN(n11382) );
  NAND2X0 U11453 ( .IN1(n8850), .IN2(g6682), .QN(n11384) );
  NAND2X0 U11454 ( .IN1(n9682), .IN2(n11380), .QN(n11383) );
  NAND3X0 U11455 ( .IN1(n11385), .IN2(n11386), .IN3(n11387), .QN(g33626) );
  NAND2X0 U11456 ( .IN1(n11388), .IN2(g6741), .QN(n11387) );
  NAND4X0 U11457 ( .IN1(n11380), .IN2(n11381), .IN3(n5398), .IN4(n9360), .QN(
        n11386) );
  NAND2X0 U11458 ( .IN1(n11389), .IN2(n10252), .QN(n11380) );
  NAND2X0 U11459 ( .IN1(n9466), .IN2(g6736), .QN(n11385) );
  NAND3X0 U11460 ( .IN1(n11390), .IN2(n11391), .IN3(n11392), .QN(g33625) );
  NAND3X0 U11461 ( .IN1(n11393), .IN2(n11394), .IN3(n11395), .QN(n11392) );
  NAND2X0 U11462 ( .IN1(n9466), .IN2(g6395), .QN(n11391) );
  NAND2X0 U11463 ( .IN1(n11396), .IN2(n9375), .QN(n11390) );
  NAND2X0 U11464 ( .IN1(n11397), .IN2(n11398), .QN(n11396) );
  NAND2X0 U11465 ( .IN1(n11399), .IN2(g6336), .QN(n11398) );
  NAND2X0 U11466 ( .IN1(n11400), .IN2(n11394), .QN(n11397) );
  NAND3X0 U11467 ( .IN1(n11401), .IN2(n11402), .IN3(n11403), .QN(g33624) );
  NAND2X0 U11468 ( .IN1(n11404), .IN2(g6395), .QN(n11403) );
  NAND4X0 U11469 ( .IN1(n11393), .IN2(n11394), .IN3(n5396), .IN4(n9360), .QN(
        n11402) );
  NAND2X0 U11470 ( .IN1(n11405), .IN2(n10255), .QN(n11394) );
  NAND2X0 U11471 ( .IN1(n9466), .IN2(g6390), .QN(n11401) );
  NAND3X0 U11472 ( .IN1(n11406), .IN2(n11407), .IN3(n11408), .QN(g33623) );
  NAND3X0 U11473 ( .IN1(n11409), .IN2(n11410), .IN3(n11411), .QN(n11408) );
  NAND2X0 U11474 ( .IN1(test_so57), .IN2(n9425), .QN(n11407) );
  NAND2X0 U11475 ( .IN1(n11412), .IN2(n9375), .QN(n11406) );
  NAND2X0 U11476 ( .IN1(n11413), .IN2(n11414), .QN(n11412) );
  NAND2X0 U11477 ( .IN1(n11415), .IN2(g5990), .QN(n11414) );
  NAND2X0 U11478 ( .IN1(n11416), .IN2(n11410), .QN(n11413) );
  NAND3X0 U11479 ( .IN1(n11417), .IN2(n11418), .IN3(n11419), .QN(g33622) );
  NAND2X0 U11480 ( .IN1(n11420), .IN2(test_so57), .QN(n11419) );
  NAND4X0 U11481 ( .IN1(n11410), .IN2(n8866), .IN3(n11409), .IN4(n9361), .QN(
        n11418) );
  NAND2X0 U11482 ( .IN1(n11421), .IN2(n10255), .QN(n11410) );
  NAND2X0 U11483 ( .IN1(test_so50), .IN2(n9411), .QN(n11417) );
  NAND3X0 U11484 ( .IN1(n11422), .IN2(n11423), .IN3(n11424), .QN(g33621) );
  NAND3X0 U11485 ( .IN1(n11425), .IN2(n11426), .IN3(n11427), .QN(n11424) );
  NAND2X0 U11486 ( .IN1(n9466), .IN2(g5703), .QN(n11423) );
  NAND2X0 U11487 ( .IN1(n11428), .IN2(n9375), .QN(n11422) );
  NAND2X0 U11488 ( .IN1(n11429), .IN2(n11430), .QN(n11428) );
  NAND2X0 U11489 ( .IN1(n11431), .IN2(g5644), .QN(n11430) );
  NAND2X0 U11490 ( .IN1(n11432), .IN2(n11426), .QN(n11429) );
  NAND3X0 U11491 ( .IN1(n11433), .IN2(n11434), .IN3(n11435), .QN(g33620) );
  NAND2X0 U11492 ( .IN1(n11436), .IN2(g5703), .QN(n11435) );
  NAND4X0 U11493 ( .IN1(n11425), .IN2(n11426), .IN3(n5397), .IN4(n9361), .QN(
        n11434) );
  NAND2X0 U11494 ( .IN1(n11437), .IN2(n10255), .QN(n11426) );
  NAND2X0 U11495 ( .IN1(n9466), .IN2(g5698), .QN(n11433) );
  NAND3X0 U11496 ( .IN1(n11438), .IN2(n11439), .IN3(n11440), .QN(g33619) );
  NAND3X0 U11497 ( .IN1(n11441), .IN2(g33959), .IN3(n9677), .QN(n11440) );
  NAND2X0 U11498 ( .IN1(n9465), .IN2(g5357), .QN(n11439) );
  NAND2X0 U11499 ( .IN1(n11442), .IN2(n9375), .QN(n11438) );
  NAND2X0 U11500 ( .IN1(n11443), .IN2(n11444), .QN(n11442) );
  NAND2X0 U11501 ( .IN1(n8845), .IN2(g5297), .QN(n11444) );
  NAND2X0 U11502 ( .IN1(n9675), .IN2(n11441), .QN(n11443) );
  NAND3X0 U11503 ( .IN1(n11445), .IN2(n11446), .IN3(n11447), .QN(g33618) );
  NAND2X0 U11504 ( .IN1(n11448), .IN2(g5357), .QN(n11447) );
  NAND4X0 U11505 ( .IN1(n11441), .IN2(g33959), .IN3(n5393), .IN4(n9361), .QN(
        n11446) );
  NAND2X0 U11506 ( .IN1(n11389), .IN2(n10255), .QN(n11441) );
  NOR2X0 U11507 ( .IN1(g4311), .IN2(n11449), .QN(n10255) );
  NOR2X0 U11508 ( .IN1(n11450), .IN2(test_so81), .QN(n11389) );
  NAND2X0 U11509 ( .IN1(n9465), .IN2(g5352), .QN(n11445) );
  NAND3X0 U11510 ( .IN1(n11451), .IN2(n10825), .IN3(n11452), .QN(g33617) );
  NAND2X0 U11511 ( .IN1(n11453), .IN2(g4552), .QN(n11452) );
  NAND4X0 U11512 ( .IN1(n11454), .IN2(n11455), .IN3(n11456), .IN4(n10825), 
        .QN(g33616) );
  NAND2X0 U11513 ( .IN1(n11457), .IN2(g4512), .QN(n11455) );
  INVX0 U11514 ( .INP(n11458), .ZN(n11454) );
  NOR2X0 U11515 ( .IN1(n9360), .IN2(n8714), .QN(n11458) );
  NAND2X0 U11516 ( .IN1(n3064), .IN2(n11459), .QN(g33615) );
  NAND2X0 U11517 ( .IN1(n11460), .IN2(g4108), .QN(n11459) );
  NAND2X0 U11518 ( .IN1(n11461), .IN2(n9375), .QN(n11460) );
  NAND2X0 U11519 ( .IN1(n9796), .IN2(n8593), .QN(n11461) );
  NAND3X0 U11520 ( .IN1(n11462), .IN2(n11463), .IN3(n11464), .QN(g33614) );
  NAND3X0 U11521 ( .IN1(n11465), .IN2(n11466), .IN3(n11467), .QN(n11464) );
  NAND2X0 U11522 ( .IN1(n9465), .IN2(g4054), .QN(n11463) );
  NAND2X0 U11523 ( .IN1(n11468), .IN2(n9375), .QN(n11462) );
  NAND2X0 U11524 ( .IN1(n11469), .IN2(n11470), .QN(n11468) );
  NAND2X0 U11525 ( .IN1(n11471), .IN2(g3990), .QN(n11470) );
  NAND2X0 U11526 ( .IN1(n11472), .IN2(n11466), .QN(n11469) );
  NAND3X0 U11527 ( .IN1(n11473), .IN2(n11474), .IN3(n11475), .QN(g33613) );
  NAND2X0 U11528 ( .IN1(n11476), .IN2(g4054), .QN(n11475) );
  NAND4X0 U11529 ( .IN1(n11465), .IN2(n11466), .IN3(n5395), .IN4(n9361), .QN(
        n11474) );
  NAND2X0 U11530 ( .IN1(n11405), .IN2(n10252), .QN(n11466) );
  NOR2X0 U11531 ( .IN1(n11477), .IN2(n8867), .QN(n11405) );
  NAND2X0 U11532 ( .IN1(n9465), .IN2(g4049), .QN(n11473) );
  NAND3X0 U11533 ( .IN1(n11478), .IN2(n11479), .IN3(n11480), .QN(g33612) );
  NAND3X0 U11534 ( .IN1(n11481), .IN2(n11482), .IN3(n11483), .QN(n11480) );
  NAND2X0 U11535 ( .IN1(n9465), .IN2(g3703), .QN(n11479) );
  NAND2X0 U11536 ( .IN1(n11484), .IN2(n9375), .QN(n11478) );
  NAND2X0 U11537 ( .IN1(n11485), .IN2(n11486), .QN(n11484) );
  NAND2X0 U11538 ( .IN1(n11487), .IN2(g3639), .QN(n11486) );
  NAND2X0 U11539 ( .IN1(n11488), .IN2(n11482), .QN(n11485) );
  NAND3X0 U11540 ( .IN1(n11489), .IN2(n11490), .IN3(n11491), .QN(g33611) );
  NAND2X0 U11541 ( .IN1(n11492), .IN2(g3703), .QN(n11491) );
  NAND4X0 U11542 ( .IN1(n11481), .IN2(n11482), .IN3(n5399), .IN4(n9361), .QN(
        n11490) );
  NAND2X0 U11543 ( .IN1(n11421), .IN2(n10252), .QN(n11482) );
  NOR2X0 U11544 ( .IN1(n11477), .IN2(test_so81), .QN(n11421) );
  INVX0 U11545 ( .INP(n3033), .ZN(n11477) );
  NAND2X0 U11546 ( .IN1(n9465), .IN2(g3698), .QN(n11489) );
  NAND2X0 U11547 ( .IN1(n11493), .IN2(n11494), .QN(g33610) );
  NAND2X0 U11548 ( .IN1(n9465), .IN2(g3352), .QN(n11494) );
  NAND2X0 U11549 ( .IN1(n11495), .IN2(n9375), .QN(n11493) );
  NAND2X0 U11550 ( .IN1(n11496), .IN2(n11497), .QN(n11495) );
  NAND2X0 U11551 ( .IN1(n11498), .IN2(g3288), .QN(n11497) );
  NAND3X0 U11552 ( .IN1(n11499), .IN2(n11500), .IN3(n11501), .QN(n11496) );
  NAND2X0 U11553 ( .IN1(n11502), .IN2(n11503), .QN(n11499) );
  NAND3X0 U11554 ( .IN1(n11504), .IN2(n11505), .IN3(n11506), .QN(g33609) );
  NAND2X0 U11555 ( .IN1(n11507), .IN2(g3352), .QN(n11506) );
  NAND4X0 U11556 ( .IN1(n5604), .IN2(n11500), .IN3(n11501), .IN4(n9361), .QN(
        n11505) );
  NAND2X0 U11557 ( .IN1(n11437), .IN2(n10252), .QN(n11500) );
  NOR2X0 U11558 ( .IN1(n11449), .IN2(n5323), .QN(n10252) );
  NAND2X0 U11559 ( .IN1(n11508), .IN2(n10168), .QN(n11449) );
  NAND2X0 U11560 ( .IN1(n11509), .IN2(n11510), .QN(n10168) );
  NAND2X0 U11561 ( .IN1(n5506), .IN2(n11320), .QN(n11510) );
  NAND2X0 U11562 ( .IN1(g72), .IN2(g4322), .QN(n11509) );
  NAND2X0 U11563 ( .IN1(n11511), .IN2(n11512), .QN(n11508) );
  NAND2X0 U11564 ( .IN1(n5540), .IN2(n9794), .QN(n11512) );
  NAND2X0 U11565 ( .IN1(g73), .IN2(g4332), .QN(n11511) );
  NOR2X0 U11566 ( .IN1(n11450), .IN2(n8867), .QN(n11437) );
  INVX0 U11567 ( .INP(n3023), .ZN(n11450) );
  NAND2X0 U11568 ( .IN1(n9464), .IN2(g3347), .QN(n11504) );
  NAND4X0 U11569 ( .IN1(n11513), .IN2(n9664), .IN3(n11514), .IN4(n11515), .QN(
        g33608) );
  NAND3X0 U11570 ( .IN1(n11516), .IN2(g2759), .IN3(n9321), .QN(n11515) );
  NAND2X0 U11571 ( .IN1(test_so30), .IN2(n9419), .QN(n11514) );
  NAND2X0 U11572 ( .IN1(n10842), .IN2(n8336), .QN(n11513) );
  INVX0 U11573 ( .INP(n11516), .ZN(n10842) );
  NAND2X0 U11574 ( .IN1(n2790), .IN2(test_so30), .QN(n11516) );
  NAND3X0 U11575 ( .IN1(n11517), .IN2(n11518), .IN3(n11519), .QN(g33607) );
  NAND2X0 U11576 ( .IN1(n9464), .IN2(g2555), .QN(n11519) );
  NAND3X0 U11577 ( .IN1(n11520), .IN2(n11521), .IN3(n3102), .QN(n11518) );
  NAND2X0 U11578 ( .IN1(n11522), .IN2(n11523), .QN(n11521) );
  NAND2X0 U11579 ( .IN1(n3111), .IN2(n9375), .QN(n11523) );
  NAND3X0 U11580 ( .IN1(n10873), .IN2(n10615), .IN3(n11524), .QN(n11522) );
  NOR2X0 U11581 ( .IN1(g504), .IN2(n10631), .QN(n10615) );
  NAND2X0 U11582 ( .IN1(n10873), .IN2(g112), .QN(n11520) );
  NOR2X0 U11583 ( .IN1(g2599), .IN2(n5521), .QN(n10873) );
  NAND2X0 U11584 ( .IN1(n11525), .IN2(g2606), .QN(n11517) );
  NAND2X0 U11585 ( .IN1(n11526), .IN2(n11527), .QN(n11525) );
  INVX0 U11586 ( .INP(n11528), .ZN(n11527) );
  NOR2X0 U11587 ( .IN1(n9419), .IN2(n3105), .QN(n11528) );
  NAND3X0 U11588 ( .IN1(n11529), .IN2(n11530), .IN3(n11531), .QN(g33606) );
  NAND2X0 U11589 ( .IN1(n10848), .IN2(g2675), .QN(n11531) );
  NAND3X0 U11590 ( .IN1(n5457), .IN2(n10846), .IN3(n9321), .QN(n11530) );
  NAND2X0 U11591 ( .IN1(n9464), .IN2(g2671), .QN(n11529) );
  NAND3X0 U11592 ( .IN1(n11532), .IN2(n11533), .IN3(n11534), .QN(g33605) );
  NAND2X0 U11593 ( .IN1(n10848), .IN2(g2671), .QN(n11534) );
  NAND2X0 U11594 ( .IN1(test_so48), .IN2(n11535), .QN(n11533) );
  NAND2X0 U11595 ( .IN1(n11536), .IN2(n9375), .QN(n11535) );
  NAND2X0 U11596 ( .IN1(n10846), .IN2(g2661), .QN(n11536) );
  NAND4X0 U11597 ( .IN1(n10846), .IN2(n9356), .IN3(n5418), .IN4(n8897), .QN(
        n11532) );
  NAND2X0 U11598 ( .IN1(n11537), .IN2(n11538), .QN(g33604) );
  NAND2X0 U11599 ( .IN1(test_so48), .IN2(n10848), .QN(n11538) );
  NAND2X0 U11600 ( .IN1(n11539), .IN2(g2661), .QN(n11537) );
  NAND2X0 U11601 ( .IN1(n11540), .IN2(n11541), .QN(g33603) );
  NAND2X0 U11602 ( .IN1(n10848), .IN2(g2648), .QN(n11541) );
  NAND2X0 U11603 ( .IN1(n11539), .IN2(g2643), .QN(n11540) );
  INVX0 U11604 ( .INP(n10848), .ZN(n11539) );
  NOR2X0 U11605 ( .IN1(n10846), .IN2(n9397), .QN(n10848) );
  INVX0 U11606 ( .INP(n10859), .ZN(n10846) );
  NAND3X0 U11607 ( .IN1(n5351), .IN2(n10861), .IN3(n5521), .QN(n10859) );
  NAND3X0 U11608 ( .IN1(n11542), .IN2(n11543), .IN3(n11544), .QN(g33602) );
  NAND2X0 U11609 ( .IN1(n9464), .IN2(g2599), .QN(n11544) );
  NAND2X0 U11610 ( .IN1(n10878), .IN2(g2629), .QN(n11543) );
  NAND2X0 U11611 ( .IN1(n10884), .IN2(n11545), .QN(n11542) );
  NOR2X0 U11612 ( .IN1(n5524), .IN2(n11546), .QN(n10884) );
  NAND3X0 U11613 ( .IN1(n11547), .IN2(n11548), .IN3(n11549), .QN(g33601) );
  NAND2X0 U11614 ( .IN1(n10878), .IN2(g2599), .QN(n11549) );
  NAND2X0 U11615 ( .IN1(n9464), .IN2(g2606), .QN(n11548) );
  NAND3X0 U11616 ( .IN1(n10890), .IN2(n11545), .IN3(n9321), .QN(n11547) );
  NOR2X0 U11617 ( .IN1(n5351), .IN2(n11546), .QN(n10890) );
  NAND2X0 U11618 ( .IN1(n11550), .IN2(n11551), .QN(g33600) );
  NAND4X0 U11619 ( .IN1(n5521), .IN2(n11552), .IN3(n9355), .IN4(n11545), .QN(
        n11551) );
  INVX0 U11620 ( .INP(n3111), .ZN(n11545) );
  NAND2X0 U11621 ( .IN1(n5351), .IN2(n11553), .QN(n11552) );
  NAND2X0 U11622 ( .IN1(n5524), .IN2(n10861), .QN(n11553) );
  NAND2X0 U11623 ( .IN1(n10878), .IN2(g2555), .QN(n11550) );
  NOR2X0 U11624 ( .IN1(n10861), .IN2(n9398), .QN(n10878) );
  INVX0 U11625 ( .INP(n11546), .ZN(n10861) );
  NOR2X0 U11626 ( .IN1(n10868), .IN2(n3102), .QN(n11546) );
  NOR2X0 U11627 ( .IN1(n11554), .IN2(n8721), .QN(n3102) );
  NOR2X0 U11628 ( .IN1(n11555), .IN2(g1514), .QN(n11554) );
  NAND3X0 U11629 ( .IN1(n11076), .IN2(n10123), .IN3(n11556), .QN(n10868) );
  NAND3X0 U11630 ( .IN1(g2689), .IN2(g2704), .IN3(g2697), .QN(n11556) );
  NAND2X0 U11631 ( .IN1(n2549), .IN2(g1300), .QN(n10123) );
  NAND3X0 U11632 ( .IN1(n11557), .IN2(n11558), .IN3(n11559), .QN(g33599) );
  NAND2X0 U11633 ( .IN1(test_so79), .IN2(n9511), .QN(n11559) );
  NAND3X0 U11634 ( .IN1(n11560), .IN2(n11561), .IN3(n716), .QN(n11558) );
  NAND2X0 U11635 ( .IN1(n11562), .IN2(n11563), .QN(n11561) );
  NAND2X0 U11636 ( .IN1(n3131), .IN2(n9375), .QN(n11563) );
  NAND3X0 U11637 ( .IN1(n10932), .IN2(n10617), .IN3(n11524), .QN(n11562) );
  NOR2X0 U11638 ( .IN1(n10631), .IN2(n5519), .QN(n10617) );
  NAND2X0 U11639 ( .IN1(n3116), .IN2(g518), .QN(n10631) );
  NAND2X0 U11640 ( .IN1(n10932), .IN2(g112), .QN(n11560) );
  NOR2X0 U11641 ( .IN1(g2465), .IN2(n5522), .QN(n10932) );
  NAND2X0 U11642 ( .IN1(n11564), .IN2(g2472), .QN(n11557) );
  NAND2X0 U11643 ( .IN1(n11526), .IN2(n11565), .QN(n11564) );
  INVX0 U11644 ( .INP(n11566), .ZN(n11565) );
  NOR2X0 U11645 ( .IN1(n9420), .IN2(n3125), .QN(n11566) );
  NAND3X0 U11646 ( .IN1(n11567), .IN2(n11568), .IN3(n11569), .QN(g33598) );
  NAND2X0 U11647 ( .IN1(n10908), .IN2(g2541), .QN(n11569) );
  NAND3X0 U11648 ( .IN1(n5461), .IN2(n10906), .IN3(n9321), .QN(n11568) );
  NAND2X0 U11649 ( .IN1(n9464), .IN2(g2537), .QN(n11567) );
  NAND3X0 U11650 ( .IN1(n11570), .IN2(n11571), .IN3(n11572), .QN(g33597) );
  NAND2X0 U11651 ( .IN1(n10908), .IN2(g2537), .QN(n11572) );
  NAND2X0 U11652 ( .IN1(n11573), .IN2(g2533), .QN(n11571) );
  NAND2X0 U11653 ( .IN1(n11574), .IN2(n9375), .QN(n11573) );
  NAND2X0 U11654 ( .IN1(n10906), .IN2(g2527), .QN(n11574) );
  NAND4X0 U11655 ( .IN1(n10906), .IN2(n9355), .IN3(n5420), .IN4(n5761), .QN(
        n11570) );
  NAND2X0 U11656 ( .IN1(n11575), .IN2(n11576), .QN(g33596) );
  NAND2X0 U11657 ( .IN1(n10908), .IN2(g2533), .QN(n11576) );
  NAND2X0 U11658 ( .IN1(n11577), .IN2(g2527), .QN(n11575) );
  NAND2X0 U11659 ( .IN1(n11578), .IN2(n11579), .QN(g33595) );
  NAND2X0 U11660 ( .IN1(n10908), .IN2(g2514), .QN(n11579) );
  NAND2X0 U11661 ( .IN1(n11577), .IN2(g2509), .QN(n11578) );
  INVX0 U11662 ( .INP(n10908), .ZN(n11577) );
  NOR2X0 U11663 ( .IN1(n10906), .IN2(n9398), .QN(n10908) );
  INVX0 U11664 ( .INP(n10919), .ZN(n10906) );
  NAND3X0 U11665 ( .IN1(n10921), .IN2(n8860), .IN3(n5522), .QN(n10919) );
  NAND3X0 U11666 ( .IN1(n11580), .IN2(n11581), .IN3(n11582), .QN(g33594) );
  NAND2X0 U11667 ( .IN1(n9464), .IN2(g2465), .QN(n11582) );
  NAND2X0 U11668 ( .IN1(n10937), .IN2(g2495), .QN(n11581) );
  NAND2X0 U11669 ( .IN1(n10943), .IN2(n11583), .QN(n11580) );
  NOR2X0 U11670 ( .IN1(n5523), .IN2(n11584), .QN(n10943) );
  NAND3X0 U11671 ( .IN1(n11585), .IN2(n11586), .IN3(n11587), .QN(g33593) );
  NAND2X0 U11672 ( .IN1(n10937), .IN2(g2465), .QN(n11587) );
  NAND2X0 U11673 ( .IN1(n9463), .IN2(g2472), .QN(n11586) );
  NAND3X0 U11674 ( .IN1(n10949), .IN2(n11583), .IN3(n9320), .QN(n11585) );
  NOR2X0 U11675 ( .IN1(n8860), .IN2(n11584), .QN(n10949) );
  NAND2X0 U11676 ( .IN1(n11588), .IN2(n11589), .QN(g33592) );
  NAND4X0 U11677 ( .IN1(n5522), .IN2(n11590), .IN3(n9355), .IN4(n11583), .QN(
        n11589) );
  INVX0 U11678 ( .INP(n3131), .ZN(n11583) );
  NAND2X0 U11679 ( .IN1(n8860), .IN2(n11591), .QN(n11590) );
  NAND2X0 U11680 ( .IN1(n5523), .IN2(n10921), .QN(n11591) );
  NAND2X0 U11681 ( .IN1(n10937), .IN2(test_so79), .QN(n11588) );
  NOR2X0 U11682 ( .IN1(n10921), .IN2(n9398), .QN(n10937) );
  INVX0 U11683 ( .INP(n11584), .ZN(n10921) );
  NOR2X0 U11684 ( .IN1(n10928), .IN2(n716), .QN(n11584) );
  NOR2X0 U11685 ( .IN1(n8442), .IN2(n11592), .QN(n716) );
  NOR3X0 U11686 ( .IN1(n11593), .IN2(n5364), .IN3(n8859), .QN(n11592) );
  NAND3X0 U11687 ( .IN1(n11076), .IN2(n10058), .IN3(n11594), .QN(n10928) );
  NAND3X0 U11688 ( .IN1(g2697), .IN2(g2689), .IN3(n5377), .QN(n11594) );
  NAND2X0 U11689 ( .IN1(n2549), .IN2(g1472), .QN(n10058) );
  NAND3X0 U11690 ( .IN1(n11595), .IN2(n11596), .IN3(n11597), .QN(g33591) );
  NAND2X0 U11691 ( .IN1(n9463), .IN2(g2287), .QN(n11597) );
  NAND3X0 U11692 ( .IN1(n11598), .IN2(n11599), .IN3(n353), .QN(n11596) );
  NAND2X0 U11693 ( .IN1(n11600), .IN2(n11601), .QN(n11599) );
  INVX0 U11694 ( .INP(n11602), .ZN(n11601) );
  NOR2X0 U11695 ( .IN1(n11603), .IN2(n9389), .QN(n11602) );
  NAND3X0 U11696 ( .IN1(n11604), .IN2(n11605), .IN3(n11524), .QN(n11600) );
  NAND2X0 U11697 ( .IN1(n11604), .IN2(g112), .QN(n11598) );
  INVX0 U11698 ( .INP(n10624), .ZN(n11604) );
  NAND2X0 U11699 ( .IN1(n5513), .IN2(g2361), .QN(n10624) );
  NAND2X0 U11700 ( .IN1(n11606), .IN2(g2338), .QN(n11595) );
  NAND2X0 U11701 ( .IN1(n11526), .IN2(n11607), .QN(n11606) );
  INVX0 U11702 ( .INP(n11608), .ZN(n11607) );
  NOR2X0 U11703 ( .IN1(n9420), .IN2(n3145), .QN(n11608) );
  NAND3X0 U11704 ( .IN1(n11609), .IN2(n11610), .IN3(n11611), .QN(g33590) );
  NAND2X0 U11705 ( .IN1(n10967), .IN2(g2407), .QN(n11611) );
  NAND3X0 U11706 ( .IN1(n5459), .IN2(n10966), .IN3(n9320), .QN(n11610) );
  NAND2X0 U11707 ( .IN1(test_so31), .IN2(n9408), .QN(n11609) );
  NAND3X0 U11708 ( .IN1(n11612), .IN2(n11613), .IN3(n11614), .QN(g33589) );
  NAND2X0 U11709 ( .IN1(test_so31), .IN2(n10967), .QN(n11614) );
  NAND2X0 U11710 ( .IN1(n11615), .IN2(g2399), .QN(n11613) );
  NAND2X0 U11711 ( .IN1(n11616), .IN2(n9375), .QN(n11615) );
  NAND2X0 U11712 ( .IN1(n10966), .IN2(g2393), .QN(n11616) );
  NAND4X0 U11713 ( .IN1(n10966), .IN2(n9356), .IN3(n5421), .IN4(n5762), .QN(
        n11612) );
  NAND2X0 U11714 ( .IN1(n11617), .IN2(n11618), .QN(g33588) );
  NAND2X0 U11715 ( .IN1(n10967), .IN2(g2399), .QN(n11618) );
  NAND2X0 U11716 ( .IN1(n11619), .IN2(g2393), .QN(n11617) );
  NAND2X0 U11717 ( .IN1(n11620), .IN2(n11621), .QN(g33587) );
  NAND2X0 U11718 ( .IN1(n10967), .IN2(g2380), .QN(n11621) );
  NAND2X0 U11719 ( .IN1(n11619), .IN2(g2375), .QN(n11620) );
  INVX0 U11720 ( .INP(n10967), .ZN(n11619) );
  NOR2X0 U11721 ( .IN1(n10966), .IN2(n9383), .QN(n10967) );
  INVX0 U11722 ( .INP(n10978), .ZN(n10966) );
  NAND3X0 U11723 ( .IN1(n5353), .IN2(n10980), .IN3(n5537), .QN(n10978) );
  NAND3X0 U11724 ( .IN1(n11622), .IN2(n11623), .IN3(n11624), .QN(g33586) );
  NAND2X0 U11725 ( .IN1(n10997), .IN2(n11603), .QN(n11624) );
  NOR2X0 U11726 ( .IN1(n5513), .IN2(n11625), .QN(n10997) );
  NAND2X0 U11727 ( .IN1(n9463), .IN2(g2331), .QN(n11623) );
  NAND3X0 U11728 ( .IN1(n11625), .IN2(g2361), .IN3(n9320), .QN(n11622) );
  NAND3X0 U11729 ( .IN1(n11626), .IN2(n11627), .IN3(n11628), .QN(g33585) );
  NAND3X0 U11730 ( .IN1(n11603), .IN2(n10980), .IN3(n11000), .QN(n11628) );
  NAND3X0 U11731 ( .IN1(n11625), .IN2(g2331), .IN3(n9320), .QN(n11627) );
  NAND2X0 U11732 ( .IN1(n9463), .IN2(g2338), .QN(n11626) );
  NAND2X0 U11733 ( .IN1(n11629), .IN2(n11630), .QN(g33584) );
  NAND2X0 U11734 ( .IN1(n11000), .IN2(n11625), .QN(n11630) );
  NOR2X0 U11735 ( .IN1(n9416), .IN2(n5353), .QN(n11000) );
  NAND4X0 U11736 ( .IN1(n5537), .IN2(n11631), .IN3(n11603), .IN4(n9361), .QN(
        n11629) );
  NAND2X0 U11737 ( .IN1(n3115), .IN2(n11605), .QN(n11603) );
  INVX0 U11738 ( .INP(n3146), .ZN(n11605) );
  NAND3X0 U11739 ( .IN1(n3116), .IN2(g504), .IN3(n5287), .QN(n3146) );
  NAND2X0 U11740 ( .IN1(n5353), .IN2(n10993), .QN(n11631) );
  NAND2X0 U11741 ( .IN1(n5513), .IN2(n10980), .QN(n10993) );
  INVX0 U11742 ( .INP(n11625), .ZN(n10980) );
  NOR2X0 U11743 ( .IN1(n10987), .IN2(n353), .QN(n11625) );
  NOR2X0 U11744 ( .IN1(n8443), .IN2(n11632), .QN(n353) );
  NOR2X0 U11745 ( .IN1(n11633), .IN2(n11593), .QN(n11632) );
  NAND3X0 U11746 ( .IN1(n11076), .IN2(n10013), .IN3(n11634), .QN(n10987) );
  NAND3X0 U11747 ( .IN1(g2689), .IN2(g2704), .IN3(n5308), .QN(n11634) );
  NAND2X0 U11748 ( .IN1(n2549), .IN2(g1448), .QN(n10013) );
  NAND3X0 U11749 ( .IN1(n11635), .IN2(n11636), .IN3(n11637), .QN(g33583) );
  NAND2X0 U11750 ( .IN1(n9463), .IN2(g2153), .QN(n11637) );
  NAND3X0 U11751 ( .IN1(n11638), .IN2(n11639), .IN3(n3160), .QN(n11636) );
  NAND2X0 U11752 ( .IN1(n11640), .IN2(n11641), .QN(n11639) );
  INVX0 U11753 ( .INP(n11642), .ZN(n11641) );
  NOR2X0 U11754 ( .IN1(n11643), .IN2(n9405), .QN(n11642) );
  NAND3X0 U11755 ( .IN1(n10626), .IN2(n10627), .IN3(n11524), .QN(n11640) );
  NAND2X0 U11756 ( .IN1(n10626), .IN2(g112), .QN(n11638) );
  NOR2X0 U11757 ( .IN1(g2197), .IN2(n5538), .QN(n10626) );
  NAND2X0 U11758 ( .IN1(n11644), .IN2(g2204), .QN(n11635) );
  NAND2X0 U11759 ( .IN1(n11526), .IN2(n11645), .QN(n11644) );
  INVX0 U11760 ( .INP(n11646), .ZN(n11645) );
  NOR2X0 U11761 ( .IN1(n9411), .IN2(n3164), .QN(n11646) );
  NAND3X0 U11762 ( .IN1(n11647), .IN2(n11648), .IN3(n11649), .QN(g33582) );
  NAND2X0 U11763 ( .IN1(n11024), .IN2(g2273), .QN(n11649) );
  NAND3X0 U11764 ( .IN1(n5458), .IN2(n11023), .IN3(n9320), .QN(n11648) );
  NAND2X0 U11765 ( .IN1(n9463), .IN2(g2269), .QN(n11647) );
  NAND3X0 U11766 ( .IN1(n11650), .IN2(n11651), .IN3(n11652), .QN(g33581) );
  NAND2X0 U11767 ( .IN1(n11024), .IN2(g2269), .QN(n11652) );
  NAND2X0 U11768 ( .IN1(test_so62), .IN2(n11653), .QN(n11651) );
  NAND2X0 U11769 ( .IN1(n11654), .IN2(n9374), .QN(n11653) );
  NAND2X0 U11770 ( .IN1(n11023), .IN2(g2259), .QN(n11654) );
  NAND4X0 U11771 ( .IN1(n11023), .IN2(n9355), .IN3(n5419), .IN4(n8898), .QN(
        n11650) );
  NAND2X0 U11772 ( .IN1(n11655), .IN2(n11656), .QN(g33580) );
  NAND2X0 U11773 ( .IN1(test_so62), .IN2(n11024), .QN(n11656) );
  NAND2X0 U11774 ( .IN1(n11657), .IN2(g2259), .QN(n11655) );
  NAND2X0 U11775 ( .IN1(n11658), .IN2(n11659), .QN(g33579) );
  NAND2X0 U11776 ( .IN1(n11024), .IN2(g2246), .QN(n11659) );
  NAND2X0 U11777 ( .IN1(n11657), .IN2(g2241), .QN(n11658) );
  INVX0 U11778 ( .INP(n11024), .ZN(n11657) );
  NOR2X0 U11779 ( .IN1(n11023), .IN2(n9406), .QN(n11024) );
  INVX0 U11780 ( .INP(n11035), .ZN(n11023) );
  NAND3X0 U11781 ( .IN1(n5356), .IN2(n11037), .IN3(n5538), .QN(n11035) );
  NAND3X0 U11782 ( .IN1(n11660), .IN2(n11661), .IN3(n11662), .QN(g33578) );
  NAND2X0 U11783 ( .IN1(n11054), .IN2(n11643), .QN(n11662) );
  NOR2X0 U11784 ( .IN1(n5514), .IN2(n11663), .QN(n11054) );
  NAND2X0 U11785 ( .IN1(n9463), .IN2(g2197), .QN(n11661) );
  NAND3X0 U11786 ( .IN1(n11663), .IN2(g2227), .IN3(n9319), .QN(n11660) );
  NAND3X0 U11787 ( .IN1(n11664), .IN2(n11665), .IN3(n11666), .QN(g33577) );
  NAND3X0 U11788 ( .IN1(n11643), .IN2(n11037), .IN3(n11057), .QN(n11666) );
  NAND3X0 U11789 ( .IN1(n11663), .IN2(g2197), .IN3(n9319), .QN(n11665) );
  NAND2X0 U11790 ( .IN1(n9462), .IN2(g2204), .QN(n11664) );
  NAND2X0 U11791 ( .IN1(n11667), .IN2(n11668), .QN(g33576) );
  NAND2X0 U11792 ( .IN1(n11057), .IN2(n11663), .QN(n11668) );
  NOR2X0 U11793 ( .IN1(n9411), .IN2(n5356), .QN(n11057) );
  NAND4X0 U11794 ( .IN1(n5538), .IN2(n11669), .IN3(n11643), .IN4(n9361), .QN(
        n11667) );
  NAND2X0 U11795 ( .IN1(n3115), .IN2(n10627), .QN(n11643) );
  INVX0 U11796 ( .INP(n3165), .ZN(n10627) );
  NAND3X0 U11797 ( .IN1(n5519), .IN2(n3116), .IN3(n5287), .QN(n3165) );
  NAND2X0 U11798 ( .IN1(n5356), .IN2(n11050), .QN(n11669) );
  NAND2X0 U11799 ( .IN1(n5514), .IN2(n11037), .QN(n11050) );
  INVX0 U11800 ( .INP(n11663), .ZN(n11037) );
  NOR2X0 U11801 ( .IN1(n11044), .IN2(n3160), .QN(n11663) );
  NOR2X0 U11802 ( .IN1(n11670), .IN2(n8444), .QN(n3160) );
  NOR2X0 U11803 ( .IN1(n11555), .IN2(n5364), .QN(n11670) );
  INVX0 U11804 ( .INP(n11671), .ZN(n11555) );
  NOR2X0 U11805 ( .IN1(n11593), .IN2(test_so49), .QN(n11671) );
  NAND4X0 U11806 ( .IN1(n8720), .IN2(n5768), .IN3(test_so68), .IN4(n11672), 
        .QN(n11593) );
  NOR3X0 U11807 ( .IN1(g1548), .IN2(n8450), .IN3(g1559), .QN(n11672) );
  NAND3X0 U11808 ( .IN1(n11076), .IN2(n9983), .IN3(n11673), .QN(n11044) );
  NAND3X0 U11809 ( .IN1(n5377), .IN2(g2689), .IN3(n5308), .QN(n11673) );
  NAND2X0 U11810 ( .IN1(n2549), .IN2(g1478), .QN(n9983) );
  NAND2X0 U11811 ( .IN1(n11375), .IN2(n11674), .QN(n11076) );
  NAND3X0 U11812 ( .IN1(n10199), .IN2(g691), .IN3(n5595), .QN(n11674) );
  NAND3X0 U11813 ( .IN1(n11675), .IN2(n11676), .IN3(n11677), .QN(g33575) );
  NAND2X0 U11814 ( .IN1(n9462), .IN2(g1996), .QN(n11677) );
  NAND2X0 U11815 ( .IN1(n11678), .IN2(n11679), .QN(n11676) );
  NAND2X0 U11816 ( .IN1(n11680), .IN2(n11681), .QN(n11679) );
  NAND3X0 U11817 ( .IN1(n10618), .IN2(n9317), .IN3(n11682), .QN(n11681) );
  INVX0 U11818 ( .INP(n11683), .ZN(n10618) );
  NAND2X0 U11819 ( .IN1(n8468), .IN2(n11684), .QN(n11680) );
  NAND2X0 U11820 ( .IN1(n11685), .IN2(n11686), .QN(n11684) );
  NAND3X0 U11821 ( .IN1(n11687), .IN2(n11683), .IN3(n11524), .QN(n11686) );
  NOR2X0 U11822 ( .IN1(g2040), .IN2(n5535), .QN(n11683) );
  NAND2X0 U11823 ( .IN1(n11682), .IN2(n9374), .QN(n11685) );
  INVX0 U11824 ( .INP(n11688), .ZN(n11682) );
  NAND2X0 U11825 ( .IN1(n11689), .IN2(g2047), .QN(n11675) );
  NAND2X0 U11826 ( .IN1(n11526), .IN2(n11690), .QN(n11689) );
  NAND2X0 U11827 ( .IN1(n11691), .IN2(n9374), .QN(n11690) );
  NAND2X0 U11828 ( .IN1(n11678), .IN2(n11687), .QN(n11691) );
  NAND3X0 U11829 ( .IN1(n11692), .IN2(n11693), .IN3(n11694), .QN(g33574) );
  NAND2X0 U11830 ( .IN1(n11083), .IN2(g2116), .QN(n11694) );
  NAND3X0 U11831 ( .IN1(n5463), .IN2(n11082), .IN3(n9319), .QN(n11693) );
  NAND2X0 U11832 ( .IN1(n9462), .IN2(g2112), .QN(n11692) );
  NAND3X0 U11833 ( .IN1(n11695), .IN2(n11696), .IN3(n11697), .QN(g33573) );
  NAND2X0 U11834 ( .IN1(n11083), .IN2(g2112), .QN(n11697) );
  NAND2X0 U11835 ( .IN1(n11698), .IN2(g2108), .QN(n11696) );
  NAND2X0 U11836 ( .IN1(n11699), .IN2(n9374), .QN(n11698) );
  NAND2X0 U11837 ( .IN1(n11082), .IN2(g2102), .QN(n11699) );
  NAND4X0 U11838 ( .IN1(n11082), .IN2(n9356), .IN3(n5666), .IN4(n5452), .QN(
        n11695) );
  NAND2X0 U11839 ( .IN1(n11700), .IN2(n11701), .QN(g33572) );
  NAND2X0 U11840 ( .IN1(n11083), .IN2(g2108), .QN(n11701) );
  NAND2X0 U11841 ( .IN1(n11702), .IN2(g2102), .QN(n11700) );
  NAND2X0 U11842 ( .IN1(n11703), .IN2(n11704), .QN(g33571) );
  NAND2X0 U11843 ( .IN1(n11083), .IN2(g2089), .QN(n11704) );
  NAND2X0 U11844 ( .IN1(n11702), .IN2(g2084), .QN(n11703) );
  INVX0 U11845 ( .INP(n11083), .ZN(n11702) );
  NOR2X0 U11846 ( .IN1(n11082), .IN2(n9406), .QN(n11083) );
  INVX0 U11847 ( .INP(n11094), .ZN(n11082) );
  NAND3X0 U11848 ( .IN1(n5355), .IN2(n11096), .IN3(n5535), .QN(n11094) );
  NAND3X0 U11849 ( .IN1(n11705), .IN2(n11706), .IN3(n11707), .QN(g33570) );
  NAND2X0 U11850 ( .IN1(n9462), .IN2(g2040), .QN(n11707) );
  NAND2X0 U11851 ( .IN1(n11708), .IN2(g2070), .QN(n11706) );
  NAND2X0 U11852 ( .IN1(n11115), .IN2(n11688), .QN(n11705) );
  NOR2X0 U11853 ( .IN1(n5505), .IN2(n11109), .QN(n11115) );
  NAND3X0 U11854 ( .IN1(n11709), .IN2(n11710), .IN3(n11711), .QN(g33569) );
  NAND2X0 U11855 ( .IN1(n11708), .IN2(g2040), .QN(n11711) );
  NAND2X0 U11856 ( .IN1(n9462), .IN2(g2047), .QN(n11710) );
  NAND3X0 U11857 ( .IN1(n11121), .IN2(n11688), .IN3(n9319), .QN(n11709) );
  NOR2X0 U11858 ( .IN1(n5355), .IN2(n11109), .QN(n11121) );
  NAND2X0 U11859 ( .IN1(n11712), .IN2(n11713), .QN(g33568) );
  NAND4X0 U11860 ( .IN1(n5535), .IN2(n11714), .IN3(n11688), .IN4(n9361), .QN(
        n11713) );
  NAND2X0 U11861 ( .IN1(n3115), .IN2(n11687), .QN(n11688) );
  INVX0 U11862 ( .INP(n10619), .ZN(n11687) );
  NAND3X0 U11863 ( .IN1(n5519), .IN2(g518), .IN3(n3195), .QN(n10619) );
  NAND2X0 U11864 ( .IN1(n5355), .IN2(n11715), .QN(n11714) );
  NAND2X0 U11865 ( .IN1(n5505), .IN2(n11096), .QN(n11715) );
  NAND2X0 U11866 ( .IN1(n11708), .IN2(g1996), .QN(n11712) );
  NOR2X0 U11867 ( .IN1(n11096), .IN2(n9404), .QN(n11708) );
  INVX0 U11868 ( .INP(n11109), .ZN(n11096) );
  NOR2X0 U11869 ( .IN1(n11103), .IN2(n11678), .QN(n11109) );
  NOR2X0 U11870 ( .IN1(n11716), .IN2(n8723), .QN(n11678) );
  NOR3X0 U11871 ( .IN1(g1171), .IN2(n11717), .IN3(g1183), .QN(n11716) );
  NAND3X0 U11872 ( .IN1(n11304), .IN2(n10119), .IN3(n11718), .QN(n11103) );
  NAND3X0 U11873 ( .IN1(g2145), .IN2(g2130), .IN3(g2138), .QN(n11718) );
  NAND2X0 U11874 ( .IN1(n5286), .IN2(g956), .QN(n10119) );
  NAND3X0 U11875 ( .IN1(n11719), .IN2(n11720), .IN3(n11721), .QN(g33567) );
  NAND2X0 U11876 ( .IN1(test_so8), .IN2(n9515), .QN(n11721) );
  NAND2X0 U11877 ( .IN1(n11722), .IN2(n11723), .QN(n11720) );
  NAND2X0 U11878 ( .IN1(n11724), .IN2(n11725), .QN(n11723) );
  NAND3X0 U11879 ( .IN1(n10622), .IN2(n9315), .IN3(n11726), .QN(n11725) );
  INVX0 U11880 ( .INP(n11727), .ZN(n10622) );
  NAND2X0 U11881 ( .IN1(n8468), .IN2(n11728), .QN(n11724) );
  NAND2X0 U11882 ( .IN1(n11729), .IN2(n11730), .QN(n11728) );
  NAND3X0 U11883 ( .IN1(n11731), .IN2(n11727), .IN3(n11524), .QN(n11730) );
  NOR2X0 U11884 ( .IN1(g1906), .IN2(n5534), .QN(n11727) );
  NAND2X0 U11885 ( .IN1(n11726), .IN2(n9374), .QN(n11729) );
  INVX0 U11886 ( .INP(n11732), .ZN(n11726) );
  NAND2X0 U11887 ( .IN1(n11733), .IN2(g1913), .QN(n11719) );
  NAND2X0 U11888 ( .IN1(n11526), .IN2(n11734), .QN(n11733) );
  NAND2X0 U11889 ( .IN1(n11735), .IN2(n9374), .QN(n11734) );
  NAND2X0 U11890 ( .IN1(n11722), .IN2(n11731), .QN(n11735) );
  NAND3X0 U11891 ( .IN1(n11736), .IN2(n11737), .IN3(n11738), .QN(g33566) );
  NAND2X0 U11892 ( .IN1(n11140), .IN2(g1982), .QN(n11738) );
  NAND3X0 U11893 ( .IN1(n5462), .IN2(n11139), .IN3(n9319), .QN(n11737) );
  NAND2X0 U11894 ( .IN1(n9462), .IN2(g1978), .QN(n11736) );
  NAND3X0 U11895 ( .IN1(n11739), .IN2(n11740), .IN3(n11741), .QN(g33565) );
  NAND2X0 U11896 ( .IN1(n11140), .IN2(g1978), .QN(n11741) );
  NAND2X0 U11897 ( .IN1(n11742), .IN2(g1974), .QN(n11740) );
  NAND2X0 U11898 ( .IN1(n11743), .IN2(n9374), .QN(n11742) );
  NAND2X0 U11899 ( .IN1(n11139), .IN2(g1968), .QN(n11743) );
  NAND4X0 U11900 ( .IN1(n11139), .IN2(n9356), .IN3(n5664), .IN4(n5450), .QN(
        n11739) );
  NAND2X0 U11901 ( .IN1(n11744), .IN2(n11745), .QN(g33564) );
  NAND2X0 U11902 ( .IN1(n11140), .IN2(g1974), .QN(n11745) );
  NAND2X0 U11903 ( .IN1(n11746), .IN2(g1968), .QN(n11744) );
  NAND2X0 U11904 ( .IN1(n11747), .IN2(n11748), .QN(g33563) );
  NAND2X0 U11905 ( .IN1(n11140), .IN2(g1955), .QN(n11748) );
  NAND2X0 U11906 ( .IN1(n11746), .IN2(g1950), .QN(n11747) );
  INVX0 U11907 ( .INP(n11140), .ZN(n11746) );
  NOR2X0 U11908 ( .IN1(n11139), .IN2(n9404), .QN(n11140) );
  INVX0 U11909 ( .INP(n11151), .ZN(n11139) );
  NAND3X0 U11910 ( .IN1(n11153), .IN2(n8861), .IN3(n5534), .QN(n11151) );
  NAND3X0 U11911 ( .IN1(n11749), .IN2(n11750), .IN3(n11751), .QN(g33562) );
  NAND2X0 U11912 ( .IN1(n9462), .IN2(g1906), .QN(n11751) );
  NAND2X0 U11913 ( .IN1(n11752), .IN2(g1936), .QN(n11750) );
  NAND2X0 U11914 ( .IN1(n11172), .IN2(n11732), .QN(n11749) );
  NOR2X0 U11915 ( .IN1(n5503), .IN2(n11166), .QN(n11172) );
  NAND3X0 U11916 ( .IN1(n11753), .IN2(n11754), .IN3(n11755), .QN(g33561) );
  NAND2X0 U11917 ( .IN1(n11752), .IN2(g1906), .QN(n11755) );
  NAND2X0 U11918 ( .IN1(n9497), .IN2(g1913), .QN(n11754) );
  NAND3X0 U11919 ( .IN1(n11178), .IN2(n11732), .IN3(n9318), .QN(n11753) );
  NOR2X0 U11920 ( .IN1(n8861), .IN2(n11166), .QN(n11178) );
  NAND2X0 U11921 ( .IN1(n11756), .IN2(n11757), .QN(g33560) );
  NAND4X0 U11922 ( .IN1(n5534), .IN2(n11758), .IN3(n11732), .IN4(n9362), .QN(
        n11757) );
  NAND2X0 U11923 ( .IN1(n3115), .IN2(n11731), .QN(n11732) );
  INVX0 U11924 ( .INP(n10623), .ZN(n11731) );
  NAND3X0 U11925 ( .IN1(g518), .IN2(g504), .IN3(n3195), .QN(n10623) );
  NAND2X0 U11926 ( .IN1(n8861), .IN2(n11759), .QN(n11758) );
  NAND2X0 U11927 ( .IN1(n5503), .IN2(n11153), .QN(n11759) );
  NAND2X0 U11928 ( .IN1(n11752), .IN2(test_so8), .QN(n11756) );
  NOR2X0 U11929 ( .IN1(n11153), .IN2(n9403), .QN(n11752) );
  INVX0 U11930 ( .INP(n11166), .ZN(n11153) );
  NOR2X0 U11931 ( .IN1(n11160), .IN2(n11722), .QN(n11166) );
  NOR2X0 U11932 ( .IN1(n11760), .IN2(n8438), .QN(n11722) );
  NOR2X0 U11933 ( .IN1(n11761), .IN2(n11717), .QN(n11760) );
  INVX0 U11934 ( .INP(n11762), .ZN(n11761) );
  NAND3X0 U11935 ( .IN1(n11304), .IN2(n10055), .IN3(n11763), .QN(n11160) );
  NAND3X0 U11936 ( .IN1(g2138), .IN2(g2130), .IN3(n5307), .QN(n11763) );
  NAND2X0 U11937 ( .IN1(n5286), .IN2(g1129), .QN(n10055) );
  NAND3X0 U11938 ( .IN1(n11764), .IN2(n11765), .IN3(n11766), .QN(g33559) );
  NAND2X0 U11939 ( .IN1(n9499), .IN2(g1728), .QN(n11766) );
  NAND4X0 U11940 ( .IN1(n11767), .IN2(n10625), .IN3(n11768), .IN4(n11769), 
        .QN(n11765) );
  NAND3X0 U11941 ( .IN1(g1802), .IN2(g112), .IN3(n5504), .QN(n11769) );
  NAND2X0 U11942 ( .IN1(n11770), .IN2(n11771), .QN(n11768) );
  NAND3X0 U11943 ( .IN1(n5504), .IN2(g1802), .IN3(n11524), .QN(n11771) );
  NAND2X0 U11944 ( .IN1(n3115), .IN2(n9374), .QN(n11770) );
  NAND2X0 U11945 ( .IN1(n11772), .IN2(g1779), .QN(n11764) );
  NAND2X0 U11946 ( .IN1(n11526), .IN2(n11773), .QN(n11772) );
  NAND2X0 U11947 ( .IN1(n11774), .IN2(n9374), .QN(n11773) );
  NAND2X0 U11948 ( .IN1(n11767), .IN2(n10625), .QN(n11774) );
  NAND3X0 U11949 ( .IN1(n11775), .IN2(n11776), .IN3(n11777), .QN(g33558) );
  NAND2X0 U11950 ( .IN1(n11196), .IN2(g1848), .QN(n11777) );
  NAND3X0 U11951 ( .IN1(n5464), .IN2(n11195), .IN3(n9319), .QN(n11776) );
  NAND2X0 U11952 ( .IN1(n9500), .IN2(g1844), .QN(n11775) );
  NAND3X0 U11953 ( .IN1(n11778), .IN2(n11779), .IN3(n11780), .QN(g33557) );
  NAND2X0 U11954 ( .IN1(n11196), .IN2(g1844), .QN(n11780) );
  NAND2X0 U11955 ( .IN1(n11781), .IN2(g1840), .QN(n11779) );
  NAND2X0 U11956 ( .IN1(n11782), .IN2(n9374), .QN(n11781) );
  NAND2X0 U11957 ( .IN1(n11195), .IN2(g1834), .QN(n11782) );
  NAND4X0 U11958 ( .IN1(n11195), .IN2(n9356), .IN3(n5665), .IN4(n5451), .QN(
        n11778) );
  NAND2X0 U11959 ( .IN1(n11783), .IN2(n11784), .QN(g33556) );
  NAND2X0 U11960 ( .IN1(n11196), .IN2(g1840), .QN(n11784) );
  NAND2X0 U11961 ( .IN1(n11785), .IN2(g1834), .QN(n11783) );
  NAND2X0 U11962 ( .IN1(n11786), .IN2(n11787), .QN(g33555) );
  NAND2X0 U11963 ( .IN1(n11196), .IN2(g1821), .QN(n11787) );
  NAND2X0 U11964 ( .IN1(n11785), .IN2(g1816), .QN(n11786) );
  INVX0 U11965 ( .INP(n11196), .ZN(n11785) );
  NOR2X0 U11966 ( .IN1(n11195), .IN2(n9403), .QN(n11196) );
  INVX0 U11967 ( .INP(n11207), .ZN(n11195) );
  NAND3X0 U11968 ( .IN1(n5352), .IN2(n11209), .IN3(n5536), .QN(n11207) );
  NAND3X0 U11969 ( .IN1(n11788), .IN2(n11789), .IN3(n11790), .QN(g33554) );
  NAND2X0 U11970 ( .IN1(n11226), .IN2(n11791), .QN(n11790) );
  NOR2X0 U11971 ( .IN1(n5504), .IN2(n11792), .QN(n11226) );
  NAND2X0 U11972 ( .IN1(n9498), .IN2(g1772), .QN(n11789) );
  NAND3X0 U11973 ( .IN1(n11792), .IN2(g1802), .IN3(n9318), .QN(n11788) );
  NAND3X0 U11974 ( .IN1(n11793), .IN2(n11794), .IN3(n11795), .QN(g33553) );
  NAND3X0 U11975 ( .IN1(n11791), .IN2(n11209), .IN3(n11229), .QN(n11795) );
  NAND3X0 U11976 ( .IN1(n11792), .IN2(g1772), .IN3(n9319), .QN(n11794) );
  NAND2X0 U11977 ( .IN1(n9483), .IN2(g1779), .QN(n11793) );
  NAND2X0 U11978 ( .IN1(n11796), .IN2(n11797), .QN(g33552) );
  NAND2X0 U11979 ( .IN1(n11229), .IN2(n11792), .QN(n11797) );
  NOR2X0 U11980 ( .IN1(n9414), .IN2(n5352), .QN(n11229) );
  NAND4X0 U11981 ( .IN1(n5536), .IN2(n11798), .IN3(n11791), .IN4(n9362), .QN(
        n11796) );
  NAND2X0 U11982 ( .IN1(n3115), .IN2(n10625), .QN(n11791) );
  INVX0 U11983 ( .INP(n10628), .ZN(n10625) );
  NAND3X0 U11984 ( .IN1(n5287), .IN2(g504), .IN3(n3195), .QN(n10628) );
  NAND2X0 U11985 ( .IN1(n5352), .IN2(n11222), .QN(n11798) );
  NAND2X0 U11986 ( .IN1(n5504), .IN2(n11209), .QN(n11222) );
  INVX0 U11987 ( .INP(n11792), .ZN(n11209) );
  NOR2X0 U11988 ( .IN1(n11216), .IN2(n11767), .QN(n11792) );
  NOR2X0 U11989 ( .IN1(n8895), .IN2(n11799), .QN(n11767) );
  NOR2X0 U11990 ( .IN1(n11800), .IN2(n11717), .QN(n11799) );
  NAND3X0 U11991 ( .IN1(n11304), .IN2(n10014), .IN3(n11801), .QN(n11216) );
  NAND3X0 U11992 ( .IN1(g2145), .IN2(g2130), .IN3(n5275), .QN(n11801) );
  NAND2X0 U11993 ( .IN1(n5286), .IN2(g1105), .QN(n10014) );
  NAND3X0 U11994 ( .IN1(n11802), .IN2(n11803), .IN3(n11804), .QN(g33551) );
  NAND2X0 U11995 ( .IN1(n9484), .IN2(g1592), .QN(n11804) );
  NAND3X0 U11996 ( .IN1(n11805), .IN2(n11806), .IN3(g33533), .QN(n11803) );
  NAND2X0 U11997 ( .IN1(n11807), .IN2(n11808), .QN(n11806) );
  NAND3X0 U11998 ( .IN1(n11809), .IN2(n9316), .IN3(n3115), .QN(n11808) );
  NAND2X0 U11999 ( .IN1(g25259), .IN2(g112), .QN(n11809) );
  NAND3X0 U12000 ( .IN1(n11524), .IN2(g25259), .IN3(n8468), .QN(n11807) );
  NAND2X0 U12001 ( .IN1(test_so75), .IN2(n11810), .QN(n11802) );
  NAND2X0 U12002 ( .IN1(n11526), .IN2(n11811), .QN(n11810) );
  NAND2X0 U12003 ( .IN1(n11812), .IN2(n9374), .QN(n11811) );
  NAND2X0 U12004 ( .IN1(g33533), .IN2(n11805), .QN(n11812) );
  NAND3X0 U12005 ( .IN1(n11813), .IN2(n11814), .IN3(n11815), .QN(g33550) );
  NAND2X0 U12006 ( .IN1(n11253), .IN2(g1714), .QN(n11815) );
  NAND3X0 U12007 ( .IN1(n5460), .IN2(n11251), .IN3(n9318), .QN(n11814) );
  NAND2X0 U12008 ( .IN1(n9485), .IN2(g1710), .QN(n11813) );
  NAND3X0 U12009 ( .IN1(n11816), .IN2(n11817), .IN3(n11818), .QN(g33549) );
  NAND2X0 U12010 ( .IN1(n11253), .IN2(g1710), .QN(n11818) );
  NAND2X0 U12011 ( .IN1(test_so15), .IN2(n11819), .QN(n11817) );
  NAND2X0 U12012 ( .IN1(n11820), .IN2(n9374), .QN(n11819) );
  NAND2X0 U12013 ( .IN1(n11251), .IN2(g1700), .QN(n11820) );
  NAND4X0 U12014 ( .IN1(n11251), .IN2(n9356), .IN3(n5417), .IN4(n8899), .QN(
        n11816) );
  NAND2X0 U12015 ( .IN1(n11821), .IN2(n11822), .QN(g33548) );
  NAND2X0 U12016 ( .IN1(test_so15), .IN2(n11253), .QN(n11822) );
  NAND2X0 U12017 ( .IN1(n11823), .IN2(g1700), .QN(n11821) );
  NAND2X0 U12018 ( .IN1(n11824), .IN2(n11825), .QN(g33547) );
  NAND2X0 U12019 ( .IN1(n11253), .IN2(g1687), .QN(n11825) );
  NAND2X0 U12020 ( .IN1(n11823), .IN2(g1682), .QN(n11824) );
  INVX0 U12021 ( .INP(n11253), .ZN(n11823) );
  NOR2X0 U12022 ( .IN1(n11251), .IN2(n9402), .QN(n11253) );
  INVX0 U12023 ( .INP(n11264), .ZN(n11251) );
  NAND3X0 U12024 ( .IN1(n5362), .IN2(n11266), .IN3(n5598), .QN(n11264) );
  NAND3X0 U12025 ( .IN1(n11826), .IN2(n11827), .IN3(n11828), .QN(g33546) );
  NAND2X0 U12026 ( .IN1(n9501), .IN2(g1636), .QN(n11828) );
  NAND2X0 U12027 ( .IN1(n11829), .IN2(g1668), .QN(n11827) );
  NAND2X0 U12028 ( .IN1(n11284), .IN2(n11830), .QN(n11826) );
  NOR2X0 U12029 ( .IN1(n5549), .IN2(n11831), .QN(n11284) );
  NAND3X0 U12030 ( .IN1(n11832), .IN2(n11833), .IN3(n11834), .QN(g33545) );
  NAND2X0 U12031 ( .IN1(n11829), .IN2(g1636), .QN(n11834) );
  NAND2X0 U12032 ( .IN1(test_so75), .IN2(n9516), .QN(n11833) );
  NAND3X0 U12033 ( .IN1(n11290), .IN2(n11830), .IN3(n9317), .QN(n11832) );
  NOR2X0 U12034 ( .IN1(n5362), .IN2(n11831), .QN(n11290) );
  NAND2X0 U12035 ( .IN1(n11835), .IN2(n11836), .QN(g33544) );
  NAND2X0 U12036 ( .IN1(n11829), .IN2(g1592), .QN(n11836) );
  NOR2X0 U12037 ( .IN1(n11266), .IN2(n9401), .QN(n11829) );
  NAND4X0 U12038 ( .IN1(n11266), .IN2(n9356), .IN3(n11830), .IN4(n11837), .QN(
        n11835) );
  NOR2X0 U12039 ( .IN1(n11838), .IN2(g1668), .QN(n11837) );
  INVX0 U12040 ( .INP(n11839), .ZN(n11838) );
  NAND2X0 U12041 ( .IN1(n3115), .IN2(n11805), .QN(n11830) );
  INVX0 U12042 ( .INP(n10612), .ZN(n11805) );
  NAND3X0 U12043 ( .IN1(n5287), .IN2(n5519), .IN3(n3195), .QN(n10612) );
  INVX0 U12044 ( .INP(n11831), .ZN(n11266) );
  NOR2X0 U12045 ( .IN1(n11273), .IN2(g33533), .QN(n11831) );
  NAND3X0 U12046 ( .IN1(n11304), .IN2(n9984), .IN3(n11840), .QN(n11273) );
  NAND3X0 U12047 ( .IN1(n5307), .IN2(g2130), .IN3(n5275), .QN(n11840) );
  NAND2X0 U12048 ( .IN1(n5286), .IN2(g1135), .QN(n9984) );
  NAND2X0 U12049 ( .IN1(n11375), .IN2(n11841), .QN(n11304) );
  NAND3X0 U12050 ( .IN1(n10198), .IN2(g691), .IN3(n5595), .QN(n11841) );
  INVX0 U12051 ( .INP(g134), .ZN(n11375) );
  NAND2X0 U12052 ( .IN1(n11842), .IN2(n11843), .QN(g33543) );
  NAND3X0 U12053 ( .IN1(n9353), .IN2(g1379), .IN3(n11844), .QN(n11843) );
  NAND2X0 U12054 ( .IN1(n11845), .IN2(n11846), .QN(n11844) );
  NAND2X0 U12055 ( .IN1(n8455), .IN2(n11847), .QN(n11846) );
  NAND2X0 U12056 ( .IN1(n11848), .IN2(g1373), .QN(n11842) );
  NAND2X0 U12057 ( .IN1(n11849), .IN2(n9374), .QN(n11848) );
  NAND3X0 U12058 ( .IN1(n11845), .IN2(n11847), .IN3(n8793), .QN(n11849) );
  NAND3X0 U12059 ( .IN1(n11850), .IN2(n11851), .IN3(n11852), .QN(g33542) );
  NAND2X0 U12060 ( .IN1(n9502), .IN2(g1270), .QN(n11852) );
  NAND3X0 U12061 ( .IN1(n11853), .IN2(n11854), .IN3(g1274), .QN(n11851) );
  NAND2X0 U12062 ( .IN1(n5730), .IN2(n11855), .QN(n11850) );
  INVX0 U12063 ( .INP(n11854), .ZN(n11855) );
  NAND2X0 U12064 ( .IN1(n11856), .IN2(n11857), .QN(g33541) );
  NAND3X0 U12065 ( .IN1(n9353), .IN2(g1036), .IN3(n11858), .QN(n11857) );
  NAND2X0 U12066 ( .IN1(n11859), .IN2(n11860), .QN(n11858) );
  NAND2X0 U12067 ( .IN1(n8457), .IN2(n11861), .QN(n11860) );
  NAND2X0 U12068 ( .IN1(n11862), .IN2(g1030), .QN(n11856) );
  NAND2X0 U12069 ( .IN1(n11863), .IN2(n9374), .QN(n11862) );
  NAND3X0 U12070 ( .IN1(n11859), .IN2(n11861), .IN3(n8792), .QN(n11863) );
  NAND3X0 U12071 ( .IN1(n11864), .IN2(n11865), .IN3(n11866), .QN(g33540) );
  NAND2X0 U12072 ( .IN1(n9503), .IN2(g925), .QN(n11866) );
  NAND3X0 U12073 ( .IN1(n11867), .IN2(n11868), .IN3(g930), .QN(n11865) );
  NAND2X0 U12074 ( .IN1(n5731), .IN2(n11869), .QN(n11864) );
  INVX0 U12075 ( .INP(n11868), .ZN(n11869) );
  NAND3X0 U12076 ( .IN1(n11870), .IN2(n11871), .IN3(n11872), .QN(g33539) );
  NAND2X0 U12077 ( .IN1(n9506), .IN2(g758), .QN(n11872) );
  NAND3X0 U12078 ( .IN1(n2404), .IN2(n11873), .IN3(g763), .QN(n11871) );
  INVX0 U12079 ( .INP(n2980), .ZN(n11873) );
  NAND2X0 U12080 ( .IN1(n2980), .IN2(n5332), .QN(n11870) );
  NAND3X0 U12081 ( .IN1(n11874), .IN2(n11875), .IN3(n11876), .QN(g33538) );
  NAND2X0 U12082 ( .IN1(n9505), .IN2(g590), .QN(n11876) );
  NAND3X0 U12083 ( .IN1(n2421), .IN2(n11877), .IN3(g595), .QN(n11875) );
  INVX0 U12084 ( .INP(n2982), .ZN(n11877) );
  NAND2X0 U12085 ( .IN1(n2982), .IN2(n5476), .QN(n11874) );
  NAND2X0 U12086 ( .IN1(n11878), .IN2(n11879), .QN(g33537) );
  INVX0 U12087 ( .INP(n11880), .ZN(n11879) );
  NOR2X0 U12088 ( .IN1(n9359), .IN2(n8822), .QN(n11880) );
  NAND3X0 U12089 ( .IN1(n2707), .IN2(g142), .IN3(n9318), .QN(n11878) );
  NOR2X0 U12090 ( .IN1(n5843), .IN2(n11881), .QN(g33536) );
  NOR2X0 U12091 ( .IN1(n2710), .IN2(n9401), .QN(n11881) );
  NAND3X0 U12092 ( .IN1(n11882), .IN2(n11883), .IN3(n11884), .QN(g33535) );
  NAND2X0 U12093 ( .IN1(n9504), .IN2(g291), .QN(n11884) );
  NAND3X0 U12094 ( .IN1(n10734), .IN2(n11885), .IN3(g294), .QN(n11883) );
  INVX0 U12095 ( .INP(n3276), .ZN(n11885) );
  NAND2X0 U12096 ( .IN1(n3276), .IN2(n5680), .QN(n11882) );
  NAND3X0 U12097 ( .IN1(n11886), .IN2(n11887), .IN3(n11888), .QN(g33534) );
  NAND2X0 U12098 ( .IN1(n9474), .IN2(g150), .QN(n11888) );
  NAND3X0 U12099 ( .IN1(n10739), .IN2(n11889), .IN3(g153), .QN(n11887) );
  INVX0 U12100 ( .INP(n3277), .ZN(n11889) );
  NAND2X0 U12101 ( .IN1(n3277), .IN2(n5677), .QN(n11886) );
  NOR2X0 U12102 ( .IN1(n8433), .IN2(n11890), .QN(g33533) );
  NOR3X0 U12103 ( .IN1(n11717), .IN2(n5363), .IN3(g1183), .QN(n11890) );
  NAND4X0 U12104 ( .IN1(n5547), .IN2(n5442), .IN3(n8722), .IN4(n11891), .QN(
        n11717) );
  NOR3X0 U12105 ( .IN1(n5320), .IN2(test_so76), .IN3(n8451), .QN(n11891) );
  NOR4X0 U12106 ( .IN1(n11892), .IN2(n11893), .IN3(n11894), .IN4(n11895), .QN(
        g33435) );
  NOR2X0 U12107 ( .IN1(n5403), .IN2(n10542), .QN(n11895) );
  NOR2X0 U12108 ( .IN1(n5544), .IN2(n10547), .QN(n11894) );
  NOR2X0 U12109 ( .IN1(n5378), .IN2(n10537), .QN(n11893) );
  NOR2X0 U12110 ( .IN1(n5610), .IN2(n10532), .QN(n11892) );
  NOR4X0 U12111 ( .IN1(n11896), .IN2(n11897), .IN3(n11898), .IN4(n11899), .QN(
        g33079) );
  NOR2X0 U12112 ( .IN1(n5404), .IN2(n10542), .QN(n11899) );
  NAND2X0 U12113 ( .IN1(n5301), .IN2(g2729), .QN(n10542) );
  NOR2X0 U12114 ( .IN1(n5545), .IN2(n10547), .QN(n11898) );
  NOR2X0 U12115 ( .IN1(n5379), .IN2(n10537), .QN(n11897) );
  NAND2X0 U12116 ( .IN1(n8469), .IN2(g2724), .QN(n10537) );
  NOR2X0 U12117 ( .IN1(n5609), .IN2(n10532), .QN(n11896) );
  NAND2X0 U12118 ( .IN1(n11900), .IN2(n11901), .QN(g33070) );
  NAND2X0 U12119 ( .IN1(n11902), .IN2(n11903), .QN(n11901) );
  NAND3X0 U12120 ( .IN1(n11904), .IN2(n11905), .IN3(n11906), .QN(n11902) );
  NAND2X0 U12121 ( .IN1(g25756), .IN2(n5646), .QN(n11906) );
  NAND2X0 U12122 ( .IN1(n11907), .IN2(n9374), .QN(n11904) );
  NAND2X0 U12123 ( .IN1(n9509), .IN2(g6565), .QN(n11900) );
  NAND2X0 U12124 ( .IN1(n11908), .IN2(n11909), .QN(g33069) );
  NAND2X0 U12125 ( .IN1(n11910), .IN2(g6561), .QN(n11909) );
  NAND2X0 U12126 ( .IN1(n11911), .IN2(n9374), .QN(n11910) );
  NAND2X0 U12127 ( .IN1(n5386), .IN2(n11903), .QN(n11911) );
  INVX0 U12128 ( .INP(n11912), .ZN(n11908) );
  NOR2X0 U12129 ( .IN1(n11913), .IN2(n5386), .QN(n11912) );
  NAND2X0 U12130 ( .IN1(n11914), .IN2(n11915), .QN(g33068) );
  NAND3X0 U12131 ( .IN1(n11903), .IN2(n9666), .IN3(n5646), .QN(n11915) );
  NAND2X0 U12132 ( .IN1(n9501), .IN2(g6555), .QN(n11914) );
  NAND2X0 U12133 ( .IN1(n11916), .IN2(n11917), .QN(g33067) );
  NAND2X0 U12134 ( .IN1(n11918), .IN2(n11903), .QN(n11917) );
  NAND2X0 U12135 ( .IN1(n764), .IN2(n11919), .QN(n11918) );
  NAND2X0 U12136 ( .IN1(n9366), .IN2(n9665), .QN(n11919) );
  INVX0 U12137 ( .INP(n11920), .ZN(n764) );
  NAND2X0 U12138 ( .IN1(n9501), .IN2(g6549), .QN(n11916) );
  NAND2X0 U12139 ( .IN1(n11921), .IN2(n11922), .QN(g33065) );
  NAND2X0 U12140 ( .IN1(n11923), .IN2(n11924), .QN(n11922) );
  NAND3X0 U12141 ( .IN1(n11925), .IN2(n11926), .IN3(n11927), .QN(n11923) );
  NAND2X0 U12142 ( .IN1(g25742), .IN2(n5651), .QN(n11927) );
  NAND2X0 U12143 ( .IN1(n9366), .IN2(n11928), .QN(n11925) );
  NAND2X0 U12144 ( .IN1(n9501), .IN2(g6219), .QN(n11921) );
  NAND2X0 U12145 ( .IN1(n11929), .IN2(n11930), .QN(g33064) );
  NAND2X0 U12146 ( .IN1(n11931), .IN2(g6215), .QN(n11930) );
  NAND2X0 U12147 ( .IN1(n11932), .IN2(n9374), .QN(n11931) );
  NAND2X0 U12148 ( .IN1(n5385), .IN2(n11924), .QN(n11932) );
  INVX0 U12149 ( .INP(n11933), .ZN(n11929) );
  NOR2X0 U12150 ( .IN1(n11934), .IN2(n5385), .QN(n11933) );
  NAND2X0 U12151 ( .IN1(n11935), .IN2(n11936), .QN(g33063) );
  NAND3X0 U12152 ( .IN1(n11924), .IN2(n9815), .IN3(n5651), .QN(n11936) );
  NAND2X0 U12153 ( .IN1(n9502), .IN2(g6209), .QN(n11935) );
  NAND2X0 U12154 ( .IN1(n11937), .IN2(n11938), .QN(g33062) );
  NAND2X0 U12155 ( .IN1(n11939), .IN2(n11924), .QN(n11938) );
  NAND2X0 U12156 ( .IN1(n1039), .IN2(n11940), .QN(n11939) );
  NAND2X0 U12157 ( .IN1(n9814), .IN2(n9374), .QN(n11940) );
  INVX0 U12158 ( .INP(n11941), .ZN(n1039) );
  NAND2X0 U12159 ( .IN1(n9502), .IN2(g6203), .QN(n11937) );
  NAND2X0 U12160 ( .IN1(n11942), .IN2(n11943), .QN(g33060) );
  NAND2X0 U12161 ( .IN1(n11944), .IN2(n11945), .QN(n11943) );
  NAND3X0 U12162 ( .IN1(n11946), .IN2(n11947), .IN3(n11948), .QN(n11944) );
  NAND2X0 U12163 ( .IN1(g25728), .IN2(n5649), .QN(n11948) );
  NAND2X0 U12164 ( .IN1(n9365), .IN2(n11949), .QN(n11946) );
  NAND2X0 U12165 ( .IN1(n9502), .IN2(g5873), .QN(n11942) );
  NAND2X0 U12166 ( .IN1(n11950), .IN2(n11951), .QN(g33059) );
  NAND2X0 U12167 ( .IN1(n11952), .IN2(g5869), .QN(n11951) );
  NAND2X0 U12168 ( .IN1(n11953), .IN2(n9374), .QN(n11952) );
  NAND2X0 U12169 ( .IN1(n5388), .IN2(n11945), .QN(n11953) );
  INVX0 U12170 ( .INP(n11954), .ZN(n11950) );
  NOR2X0 U12171 ( .IN1(n11955), .IN2(n5388), .QN(n11954) );
  NAND2X0 U12172 ( .IN1(n11956), .IN2(n11957), .QN(g33058) );
  NAND3X0 U12173 ( .IN1(n11945), .IN2(n9813), .IN3(n5649), .QN(n11957) );
  NAND2X0 U12174 ( .IN1(n9502), .IN2(g5863), .QN(n11956) );
  NAND2X0 U12175 ( .IN1(n11958), .IN2(n11959), .QN(g33057) );
  NAND2X0 U12176 ( .IN1(n11960), .IN2(n11945), .QN(n11959) );
  NAND2X0 U12177 ( .IN1(n1109), .IN2(n11961), .QN(n11960) );
  NAND2X0 U12178 ( .IN1(n9812), .IN2(n9373), .QN(n11961) );
  INVX0 U12179 ( .INP(n11962), .ZN(n1109) );
  NAND2X0 U12180 ( .IN1(n9502), .IN2(g5857), .QN(n11958) );
  NAND2X0 U12181 ( .IN1(n11963), .IN2(n11964), .QN(g33055) );
  NAND2X0 U12182 ( .IN1(n11965), .IN2(n11966), .QN(n11964) );
  NAND3X0 U12183 ( .IN1(n11967), .IN2(n11968), .IN3(n11969), .QN(n11965) );
  NAND2X0 U12184 ( .IN1(g25714), .IN2(n5647), .QN(n11969) );
  NAND2X0 U12185 ( .IN1(n9366), .IN2(n11970), .QN(n11967) );
  NAND2X0 U12186 ( .IN1(n9502), .IN2(g5527), .QN(n11963) );
  NAND2X0 U12187 ( .IN1(n11971), .IN2(n11972), .QN(g33054) );
  NAND2X0 U12188 ( .IN1(n11973), .IN2(g5523), .QN(n11972) );
  NAND2X0 U12189 ( .IN1(n11974), .IN2(n9373), .QN(n11973) );
  NAND2X0 U12190 ( .IN1(n5389), .IN2(n11966), .QN(n11974) );
  INVX0 U12191 ( .INP(n11975), .ZN(n11971) );
  NOR2X0 U12192 ( .IN1(n11976), .IN2(n5389), .QN(n11975) );
  NAND2X0 U12193 ( .IN1(n11977), .IN2(n11978), .QN(g33053) );
  NAND3X0 U12194 ( .IN1(n11966), .IN2(n9688), .IN3(n5647), .QN(n11978) );
  NAND2X0 U12195 ( .IN1(n9502), .IN2(g5517), .QN(n11977) );
  NAND2X0 U12196 ( .IN1(n11979), .IN2(n11980), .QN(g33052) );
  NAND2X0 U12197 ( .IN1(n11981), .IN2(n11966), .QN(n11980) );
  NAND2X0 U12198 ( .IN1(n498), .IN2(n11982), .QN(n11981) );
  NAND2X0 U12199 ( .IN1(n9366), .IN2(n9687), .QN(n11982) );
  INVX0 U12200 ( .INP(n11983), .ZN(n498) );
  NAND2X0 U12201 ( .IN1(n9503), .IN2(g5511), .QN(n11979) );
  NAND2X0 U12202 ( .IN1(n11984), .IN2(n11985), .QN(g33050) );
  NAND2X0 U12203 ( .IN1(n11986), .IN2(n11987), .QN(n11985) );
  NAND3X0 U12204 ( .IN1(n11988), .IN2(n11989), .IN3(n11990), .QN(n11986) );
  NAND2X0 U12205 ( .IN1(g25700), .IN2(n5650), .QN(n11990) );
  NAND2X0 U12206 ( .IN1(n9365), .IN2(n11991), .QN(n11988) );
  NAND2X0 U12207 ( .IN1(n9503), .IN2(g5180), .QN(n11984) );
  NAND2X0 U12208 ( .IN1(n11992), .IN2(n11993), .QN(g33049) );
  NAND2X0 U12209 ( .IN1(n11994), .IN2(g5176), .QN(n11993) );
  NAND2X0 U12210 ( .IN1(n11995), .IN2(n9373), .QN(n11994) );
  NAND2X0 U12211 ( .IN1(n5384), .IN2(n11987), .QN(n11995) );
  INVX0 U12212 ( .INP(n11996), .ZN(n11992) );
  NOR2X0 U12213 ( .IN1(n11997), .IN2(n5384), .QN(n11996) );
  NAND2X0 U12214 ( .IN1(n11998), .IN2(n11999), .QN(g33048) );
  NAND3X0 U12215 ( .IN1(n11987), .IN2(n9668), .IN3(n5650), .QN(n11999) );
  NAND2X0 U12216 ( .IN1(n9503), .IN2(g5170), .QN(n11998) );
  NAND2X0 U12217 ( .IN1(n12000), .IN2(n12001), .QN(g33047) );
  NAND2X0 U12218 ( .IN1(n12002), .IN2(n11987), .QN(n12001) );
  NAND2X0 U12219 ( .IN1(n758), .IN2(n12003), .QN(n12002) );
  NAND2X0 U12220 ( .IN1(n9364), .IN2(n9667), .QN(n12003) );
  INVX0 U12221 ( .INP(n12004), .ZN(n758) );
  NAND2X0 U12222 ( .IN1(n9503), .IN2(g5164), .QN(n12000) );
  NAND3X0 U12223 ( .IN1(n12005), .IN2(n12006), .IN3(n12007), .QN(g33046) );
  NAND2X0 U12224 ( .IN1(n9503), .IN2(g5052), .QN(n12007) );
  NAND2X0 U12225 ( .IN1(n5615), .IN2(n12008), .QN(n12006) );
  NAND2X0 U12226 ( .IN1(n12009), .IN2(n12010), .QN(n12008) );
  NAND3X0 U12227 ( .IN1(n12011), .IN2(n12010), .IN3(g5057), .QN(n12005) );
  NAND2X0 U12228 ( .IN1(n12012), .IN2(g5052), .QN(n12010) );
  NAND3X0 U12229 ( .IN1(n12013), .IN2(n12014), .IN3(n12015), .QN(g33045) );
  NAND2X0 U12230 ( .IN1(n11453), .IN2(g4567), .QN(n12015) );
  NAND3X0 U12231 ( .IN1(n12014), .IN2(n10825), .IN3(n12016), .QN(g33044) );
  NAND2X0 U12232 ( .IN1(test_so93), .IN2(n11453), .QN(n12016) );
  NAND3X0 U12233 ( .IN1(n12017), .IN2(n11451), .IN3(n12018), .QN(g33043) );
  NAND2X0 U12234 ( .IN1(test_so16), .IN2(n11453), .QN(n12018) );
  NAND3X0 U12235 ( .IN1(n12017), .IN2(n12014), .IN3(n12019), .QN(g33042) );
  NAND2X0 U12236 ( .IN1(n11453), .IN2(g4540), .QN(n12019) );
  NAND2X0 U12237 ( .IN1(n12020), .IN2(g4578), .QN(n12014) );
  NAND3X0 U12238 ( .IN1(n12013), .IN2(n11451), .IN3(n12021), .QN(g33041) );
  NAND2X0 U12239 ( .IN1(test_so56), .IN2(n11453), .QN(n12021) );
  NAND3X0 U12240 ( .IN1(n12022), .IN2(n10825), .IN3(n12023), .QN(g33040) );
  NAND2X0 U12241 ( .IN1(n11453), .IN2(g4504), .QN(n12023) );
  NAND2X0 U12242 ( .IN1(n12020), .IN2(n10831), .QN(n10825) );
  INVX0 U12243 ( .INP(n10145), .ZN(n10831) );
  NOR2X0 U12244 ( .IN1(g73), .IN2(g72), .QN(n10145) );
  NAND3X0 U12245 ( .IN1(n12013), .IN2(n11456), .IN3(n12024), .QN(g33039) );
  NAND2X0 U12246 ( .IN1(n11453), .IN2(g4501), .QN(n12024) );
  NAND3X0 U12247 ( .IN1(n12013), .IN2(n12022), .IN3(n12025), .QN(g33038) );
  NAND2X0 U12248 ( .IN1(n11453), .IN2(g4498), .QN(n12025) );
  NAND2X0 U12249 ( .IN1(n12020), .IN2(n12026), .QN(n12013) );
  NAND2X0 U12250 ( .IN1(g72), .IN2(n10167), .QN(n12026) );
  INVX0 U12251 ( .INP(g73), .ZN(n10167) );
  NAND3X0 U12252 ( .IN1(n12017), .IN2(n11456), .IN3(n12027), .QN(g33037) );
  NAND2X0 U12253 ( .IN1(n11453), .IN2(g4495), .QN(n12027) );
  NAND3X0 U12254 ( .IN1(n12017), .IN2(n12022), .IN3(n12028), .QN(g33036) );
  NAND2X0 U12255 ( .IN1(n11453), .IN2(g4480), .QN(n12028) );
  INVX0 U12256 ( .INP(n12029), .ZN(n12022) );
  NOR2X0 U12257 ( .IN1(n11453), .IN2(n8404), .QN(n12029) );
  INVX0 U12258 ( .INP(n12020), .ZN(n11453) );
  NAND2X0 U12259 ( .IN1(n12020), .IN2(n12030), .QN(n12017) );
  NAND2X0 U12260 ( .IN1(g73), .IN2(n11320), .QN(n12030) );
  INVX0 U12261 ( .INP(g72), .ZN(n11320) );
  NAND4X0 U12262 ( .IN1(n12031), .IN2(n12032), .IN3(n12033), .IN4(n12034), 
        .QN(g33035) );
  NAND3X0 U12263 ( .IN1(n12035), .IN2(g4108), .IN3(n9326), .QN(n12034) );
  NAND2X0 U12264 ( .IN1(n9503), .IN2(g4098), .QN(n12033) );
  NAND2X0 U12265 ( .IN1(n9796), .IN2(n5715), .QN(n12031) );
  INVX0 U12266 ( .INP(n12035), .ZN(n9796) );
  NAND2X0 U12267 ( .IN1(n12036), .IN2(n12037), .QN(g33034) );
  NAND2X0 U12268 ( .IN1(n12038), .IN2(n12039), .QN(n12037) );
  NAND3X0 U12269 ( .IN1(n12040), .IN2(n12041), .IN3(n12042), .QN(n12038) );
  NAND2X0 U12270 ( .IN1(g25676), .IN2(n8868), .QN(n12042) );
  NAND2X0 U12271 ( .IN1(n9366), .IN2(n12043), .QN(n12040) );
  NAND2X0 U12272 ( .IN1(n9503), .IN2(g3873), .QN(n12036) );
  NAND2X0 U12273 ( .IN1(n12044), .IN2(n12045), .QN(g33033) );
  NAND2X0 U12274 ( .IN1(test_so33), .IN2(n12046), .QN(n12045) );
  NAND2X0 U12275 ( .IN1(n12047), .IN2(n9373), .QN(n12046) );
  NAND2X0 U12276 ( .IN1(n5387), .IN2(n12039), .QN(n12047) );
  INVX0 U12277 ( .INP(n12048), .ZN(n12044) );
  NOR2X0 U12278 ( .IN1(n12049), .IN2(n5387), .QN(n12048) );
  NAND2X0 U12279 ( .IN1(n12050), .IN2(n12051), .QN(g33032) );
  NAND3X0 U12280 ( .IN1(n9811), .IN2(n8868), .IN3(n12039), .QN(n12051) );
  NAND2X0 U12281 ( .IN1(n9504), .IN2(g3863), .QN(n12050) );
  NAND2X0 U12282 ( .IN1(n12052), .IN2(n12053), .QN(g33031) );
  NAND2X0 U12283 ( .IN1(n12054), .IN2(n12039), .QN(n12053) );
  NAND2X0 U12284 ( .IN1(n1180), .IN2(n12055), .QN(n12054) );
  NAND2X0 U12285 ( .IN1(n9810), .IN2(n9373), .QN(n12055) );
  INVX0 U12286 ( .INP(n12056), .ZN(n1180) );
  NAND2X0 U12287 ( .IN1(n9504), .IN2(g3857), .QN(n12052) );
  NAND2X0 U12288 ( .IN1(n12057), .IN2(n12058), .QN(g33029) );
  NAND2X0 U12289 ( .IN1(n12059), .IN2(n12060), .QN(n12058) );
  NAND3X0 U12290 ( .IN1(n12061), .IN2(n12062), .IN3(n12063), .QN(n12059) );
  NAND2X0 U12291 ( .IN1(g25662), .IN2(n5645), .QN(n12063) );
  NAND2X0 U12292 ( .IN1(n9365), .IN2(n12064), .QN(n12061) );
  NAND2X0 U12293 ( .IN1(n9504), .IN2(g3522), .QN(n12057) );
  NAND2X0 U12294 ( .IN1(n12065), .IN2(n12066), .QN(g33028) );
  NAND2X0 U12295 ( .IN1(n12067), .IN2(g3518), .QN(n12066) );
  NAND2X0 U12296 ( .IN1(n12068), .IN2(n9373), .QN(n12067) );
  NAND2X0 U12297 ( .IN1(n5383), .IN2(n12060), .QN(n12068) );
  INVX0 U12298 ( .INP(n12069), .ZN(n12065) );
  NOR2X0 U12299 ( .IN1(n12070), .IN2(n5383), .QN(n12069) );
  NAND2X0 U12300 ( .IN1(n12071), .IN2(n12072), .QN(g33027) );
  NAND3X0 U12301 ( .IN1(n12060), .IN2(n9670), .IN3(n5645), .QN(n12072) );
  NAND2X0 U12302 ( .IN1(n9504), .IN2(g3512), .QN(n12071) );
  NAND2X0 U12303 ( .IN1(n12073), .IN2(n12074), .QN(g33026) );
  NAND2X0 U12304 ( .IN1(n12075), .IN2(n12060), .QN(n12074) );
  NAND2X0 U12305 ( .IN1(n75), .IN2(n12076), .QN(n12075) );
  NAND2X0 U12306 ( .IN1(n9365), .IN2(n9669), .QN(n12076) );
  INVX0 U12307 ( .INP(n12077), .ZN(n75) );
  NAND2X0 U12308 ( .IN1(n9504), .IN2(g3506), .QN(n12073) );
  NAND3X0 U12309 ( .IN1(n12078), .IN2(n12079), .IN3(n12080), .QN(g33024) );
  NAND2X0 U12310 ( .IN1(g25648), .IN2(n12081), .QN(n12080) );
  NAND2X0 U12311 ( .IN1(n9504), .IN2(g3171), .QN(n12079) );
  NAND3X0 U12312 ( .IN1(n12082), .IN2(n12083), .IN3(n9326), .QN(n12078) );
  NAND2X0 U12313 ( .IN1(n12084), .IN2(n536), .QN(n12082) );
  NAND2X0 U12314 ( .IN1(n12085), .IN2(n12086), .QN(g33023) );
  NAND3X0 U12315 ( .IN1(n9350), .IN2(g3171), .IN3(n12081), .QN(n12086) );
  NAND2X0 U12316 ( .IN1(n12087), .IN2(g3167), .QN(n12085) );
  NAND2X0 U12317 ( .IN1(n12088), .IN2(n9373), .QN(n12087) );
  NAND2X0 U12318 ( .IN1(n5603), .IN2(n12083), .QN(n12088) );
  NAND2X0 U12319 ( .IN1(n12089), .IN2(n12090), .QN(g33022) );
  NAND2X0 U12320 ( .IN1(n12081), .IN2(n9659), .QN(n12090) );
  INVX0 U12321 ( .INP(n12091), .ZN(n12081) );
  NAND2X0 U12322 ( .IN1(n9504), .IN2(g3161), .QN(n12089) );
  NAND2X0 U12323 ( .IN1(n12092), .IN2(n12093), .QN(g33021) );
  NAND2X0 U12324 ( .IN1(n12094), .IN2(n12083), .QN(n12093) );
  NAND2X0 U12325 ( .IN1(n90), .IN2(n12095), .QN(n12094) );
  NAND2X0 U12326 ( .IN1(n9365), .IN2(n9658), .QN(n12095) );
  INVX0 U12327 ( .INP(n12096), .ZN(n90) );
  NAND2X0 U12328 ( .IN1(n9505), .IN2(g3155), .QN(n12092) );
  NAND3X0 U12329 ( .IN1(n12097), .IN2(n12098), .IN3(n9664), .QN(g33019) );
  NAND2X0 U12330 ( .IN1(n9505), .IN2(g2748), .QN(n12098) );
  NAND2X0 U12331 ( .IN1(n12099), .IN2(n9373), .QN(n12097) );
  NAND2X0 U12332 ( .IN1(n12100), .IN2(n12101), .QN(n12099) );
  NAND2X0 U12333 ( .IN1(test_so30), .IN2(n12102), .QN(n12101) );
  INVX0 U12334 ( .INP(n2790), .ZN(n12102) );
  NAND2X0 U12335 ( .IN1(n2790), .IN2(n5300), .QN(n12100) );
  NAND4X0 U12336 ( .IN1(n12103), .IN2(n12104), .IN3(n12105), .IN4(n12106), 
        .QN(g33018) );
  NAND2X0 U12337 ( .IN1(n9505), .IN2(g2610), .QN(n12106) );
  NAND4X0 U12338 ( .IN1(n3511), .IN2(n11524), .IN3(n12107), .IN4(n8759), .QN(
        n12105) );
  NOR2X0 U12339 ( .IN1(n5508), .IN2(n12108), .QN(n12107) );
  NAND3X0 U12340 ( .IN1(n3512), .IN2(n12109), .IN3(n3517), .QN(n12104) );
  INVX0 U12341 ( .INP(n3513), .ZN(n12109) );
  NAND2X0 U12342 ( .IN1(n3524), .IN2(n10761), .QN(n3513) );
  INVX0 U12343 ( .INP(n3006), .ZN(n10761) );
  NAND3X0 U12344 ( .IN1(g2619), .IN2(g110), .IN3(n8759), .QN(n3512) );
  NAND2X0 U12345 ( .IN1(test_so40), .IN2(n12110), .QN(n12103) );
  NAND3X0 U12346 ( .IN1(n12111), .IN2(n11526), .IN3(n12112), .QN(n12110) );
  NAND2X0 U12347 ( .IN1(n3006), .IN2(n9373), .QN(n12112) );
  NAND2X0 U12348 ( .IN1(n3525), .IN2(n3505), .QN(n3006) );
  NAND4X0 U12349 ( .IN1(n12113), .IN2(n12114), .IN3(n12115), .IN4(n12116), 
        .QN(g33017) );
  NAND2X0 U12350 ( .IN1(n12117), .IN2(g2619), .QN(n12115) );
  NAND2X0 U12351 ( .IN1(n3517), .IN2(g2610), .QN(n12114) );
  NAND2X0 U12352 ( .IN1(test_so40), .IN2(n9512), .QN(n12113) );
  NAND3X0 U12353 ( .IN1(n12118), .IN2(n12119), .IN3(n12116), .QN(g33016) );
  NAND2X0 U12354 ( .IN1(n12117), .IN2(g2610), .QN(n12119) );
  NAND2X0 U12355 ( .IN1(n12111), .IN2(g2587), .QN(n12118) );
  NAND4X0 U12356 ( .IN1(n12120), .IN2(n12121), .IN3(n12122), .IN4(n12116), 
        .QN(g33015) );
  INVX0 U12357 ( .INP(n3519), .ZN(n12116) );
  NAND3X0 U12358 ( .IN1(n5508), .IN2(n12123), .IN3(n3517), .QN(n12122) );
  NAND2X0 U12359 ( .IN1(n12117), .IN2(g2587), .QN(n12121) );
  NAND2X0 U12360 ( .IN1(test_so34), .IN2(n9424), .QN(n12120) );
  NAND4X0 U12361 ( .IN1(n12124), .IN2(n12125), .IN3(n12126), .IN4(n12127), 
        .QN(g33014) );
  NAND2X0 U12362 ( .IN1(n9505), .IN2(g2476), .QN(n12127) );
  NAND4X0 U12363 ( .IN1(n3530), .IN2(n11524), .IN3(n12128), .IN4(n8758), .QN(
        n12126) );
  NOR2X0 U12364 ( .IN1(n5509), .IN2(n12129), .QN(n12128) );
  NAND3X0 U12365 ( .IN1(n3531), .IN2(n12130), .IN3(n3536), .QN(n12125) );
  INVX0 U12366 ( .INP(n3532), .ZN(n12130) );
  NAND2X0 U12367 ( .IN1(n3524), .IN2(n10760), .QN(n3532) );
  INVX0 U12368 ( .INP(n3007), .ZN(n10760) );
  NAND3X0 U12369 ( .IN1(g2485), .IN2(g110), .IN3(n8758), .QN(n3531) );
  NAND2X0 U12370 ( .IN1(n12131), .IN2(g2491), .QN(n12124) );
  NAND3X0 U12371 ( .IN1(n12132), .IN2(n11526), .IN3(n12133), .QN(n12131) );
  NAND2X0 U12372 ( .IN1(n3007), .IN2(n9373), .QN(n12133) );
  NAND3X0 U12373 ( .IN1(n5349), .IN2(g2748), .IN3(n3525), .QN(n3007) );
  NAND4X0 U12374 ( .IN1(n12134), .IN2(n12135), .IN3(n12136), .IN4(n12137), 
        .QN(g33013) );
  NAND2X0 U12375 ( .IN1(n12138), .IN2(g2485), .QN(n12136) );
  NAND2X0 U12376 ( .IN1(n3536), .IN2(g2476), .QN(n12135) );
  NAND2X0 U12377 ( .IN1(n9505), .IN2(g2491), .QN(n12134) );
  NAND3X0 U12378 ( .IN1(n12139), .IN2(n12140), .IN3(n12137), .QN(g33012) );
  NAND2X0 U12379 ( .IN1(n12138), .IN2(g2476), .QN(n12140) );
  NAND2X0 U12380 ( .IN1(n12132), .IN2(g2453), .QN(n12139) );
  NAND4X0 U12381 ( .IN1(n12141), .IN2(n12142), .IN3(n12143), .IN4(n12137), 
        .QN(g33011) );
  INVX0 U12382 ( .INP(n3538), .ZN(n12137) );
  NAND3X0 U12383 ( .IN1(n5509), .IN2(n12144), .IN3(n3536), .QN(n12143) );
  NAND2X0 U12384 ( .IN1(n12138), .IN2(g2453), .QN(n12142) );
  NAND2X0 U12385 ( .IN1(n9505), .IN2(g2461), .QN(n12141) );
  NAND4X0 U12386 ( .IN1(n12145), .IN2(n12146), .IN3(n12147), .IN4(n12148), 
        .QN(g33010) );
  NAND2X0 U12387 ( .IN1(test_so21), .IN2(n9417), .QN(n12148) );
  NAND4X0 U12388 ( .IN1(n3548), .IN2(n11524), .IN3(n12149), .IN4(n8869), .QN(
        n12147) );
  NOR2X0 U12389 ( .IN1(n5511), .IN2(n12150), .QN(n12149) );
  NAND3X0 U12390 ( .IN1(n3549), .IN2(n12151), .IN3(n3555), .QN(n12146) );
  INVX0 U12391 ( .INP(n3551), .ZN(n12151) );
  NAND2X0 U12392 ( .IN1(n3524), .IN2(n10759), .QN(n3551) );
  INVX0 U12393 ( .INP(n3550), .ZN(n10759) );
  NAND3X0 U12394 ( .IN1(g110), .IN2(n8869), .IN3(g2351), .QN(n3549) );
  NAND2X0 U12395 ( .IN1(n12152), .IN2(g2357), .QN(n12145) );
  NAND3X0 U12396 ( .IN1(n12153), .IN2(n11526), .IN3(n12154), .QN(n12152) );
  NAND2X0 U12397 ( .IN1(n3550), .IN2(n9373), .QN(n12154) );
  NAND3X0 U12398 ( .IN1(n5516), .IN2(g2741), .IN3(n3525), .QN(n3550) );
  NAND4X0 U12399 ( .IN1(n12155), .IN2(n12156), .IN3(n12157), .IN4(n12158), 
        .QN(g33009) );
  NAND2X0 U12400 ( .IN1(n12159), .IN2(g2351), .QN(n12157) );
  NAND2X0 U12401 ( .IN1(n3555), .IN2(test_so21), .QN(n12156) );
  NAND2X0 U12402 ( .IN1(n9505), .IN2(g2357), .QN(n12155) );
  NAND3X0 U12403 ( .IN1(n12160), .IN2(n12161), .IN3(n12158), .QN(g33008) );
  NAND2X0 U12404 ( .IN1(n12159), .IN2(test_so21), .QN(n12161) );
  NAND2X0 U12405 ( .IN1(n12153), .IN2(g2319), .QN(n12160) );
  NAND4X0 U12406 ( .IN1(n12162), .IN2(n12163), .IN3(n12164), .IN4(n12158), 
        .QN(g33007) );
  INVX0 U12407 ( .INP(n3557), .ZN(n12158) );
  NAND3X0 U12408 ( .IN1(n5511), .IN2(n12165), .IN3(n3555), .QN(n12164) );
  NAND2X0 U12409 ( .IN1(n12159), .IN2(g2319), .QN(n12163) );
  NAND2X0 U12410 ( .IN1(n9506), .IN2(g2327), .QN(n12162) );
  NAND4X0 U12411 ( .IN1(n12166), .IN2(n12167), .IN3(n12168), .IN4(n12169), 
        .QN(g33006) );
  NAND2X0 U12412 ( .IN1(n9506), .IN2(g2208), .QN(n12169) );
  NAND4X0 U12413 ( .IN1(n3567), .IN2(n11524), .IN3(n12170), .IN4(n8756), .QN(
        n12168) );
  NOR2X0 U12414 ( .IN1(n5512), .IN2(n12171), .QN(n12170) );
  NAND3X0 U12415 ( .IN1(n3568), .IN2(n12172), .IN3(n3574), .QN(n12167) );
  INVX0 U12416 ( .INP(n3570), .ZN(n12172) );
  NAND2X0 U12417 ( .IN1(n3524), .IN2(n10758), .QN(n3570) );
  INVX0 U12418 ( .INP(n3569), .ZN(n10758) );
  NAND3X0 U12419 ( .IN1(g2217), .IN2(g110), .IN3(n8756), .QN(n3568) );
  NAND2X0 U12420 ( .IN1(n12173), .IN2(g2223), .QN(n12166) );
  NAND3X0 U12421 ( .IN1(n12174), .IN2(n11526), .IN3(n12175), .QN(n12173) );
  NAND2X0 U12422 ( .IN1(n3569), .IN2(n9373), .QN(n12175) );
  NAND3X0 U12423 ( .IN1(n5516), .IN2(n5349), .IN3(n3525), .QN(n3569) );
  NAND4X0 U12424 ( .IN1(n12176), .IN2(n12177), .IN3(n12178), .IN4(n12179), 
        .QN(g33005) );
  NAND2X0 U12425 ( .IN1(n12180), .IN2(g2217), .QN(n12178) );
  NAND2X0 U12426 ( .IN1(n3574), .IN2(g2208), .QN(n12177) );
  NAND2X0 U12427 ( .IN1(n9506), .IN2(g2223), .QN(n12176) );
  NAND3X0 U12428 ( .IN1(n12181), .IN2(n12182), .IN3(n12179), .QN(g33004) );
  NAND2X0 U12429 ( .IN1(n12180), .IN2(g2208), .QN(n12182) );
  NAND2X0 U12430 ( .IN1(n12174), .IN2(g2185), .QN(n12181) );
  NAND4X0 U12431 ( .IN1(n12183), .IN2(n12184), .IN3(n12185), .IN4(n12179), 
        .QN(g33003) );
  INVX0 U12432 ( .INP(n3576), .ZN(n12179) );
  NAND3X0 U12433 ( .IN1(n5512), .IN2(n12186), .IN3(n3574), .QN(n12185) );
  NAND2X0 U12434 ( .IN1(n12180), .IN2(g2185), .QN(n12184) );
  NAND2X0 U12435 ( .IN1(n9506), .IN2(g2193), .QN(n12183) );
  NAND4X0 U12436 ( .IN1(n12187), .IN2(n12188), .IN3(n12189), .IN4(n12190), 
        .QN(g33002) );
  NAND2X0 U12437 ( .IN1(n9506), .IN2(g2051), .QN(n12190) );
  NAND4X0 U12438 ( .IN1(n3586), .IN2(n11524), .IN3(n12191), .IN4(n8760), .QN(
        n12189) );
  NOR2X0 U12439 ( .IN1(n5507), .IN2(n12192), .QN(n12191) );
  NAND3X0 U12440 ( .IN1(n3587), .IN2(n12193), .IN3(n3593), .QN(n12188) );
  INVX0 U12441 ( .INP(n3589), .ZN(n12193) );
  NAND2X0 U12442 ( .IN1(n3524), .IN2(n10754), .QN(n3589) );
  INVX0 U12443 ( .INP(n3588), .ZN(n10754) );
  NAND3X0 U12444 ( .IN1(g2060), .IN2(g110), .IN3(n8760), .QN(n3587) );
  NAND2X0 U12445 ( .IN1(n12194), .IN2(g2066), .QN(n12187) );
  NAND3X0 U12446 ( .IN1(n12195), .IN2(n11526), .IN3(n12196), .QN(n12194) );
  NAND2X0 U12447 ( .IN1(n3588), .IN2(n9373), .QN(n12196) );
  NAND3X0 U12448 ( .IN1(n826), .IN2(n5300), .IN3(n3505), .QN(n3588) );
  NAND4X0 U12449 ( .IN1(n12197), .IN2(n12198), .IN3(n12199), .IN4(n12200), 
        .QN(g33001) );
  NAND2X0 U12450 ( .IN1(n12201), .IN2(g2060), .QN(n12199) );
  NAND2X0 U12451 ( .IN1(n3593), .IN2(g2051), .QN(n12198) );
  NAND2X0 U12452 ( .IN1(n9506), .IN2(g2066), .QN(n12197) );
  NAND3X0 U12453 ( .IN1(n12202), .IN2(n12203), .IN3(n12200), .QN(g33000) );
  NAND2X0 U12454 ( .IN1(n12201), .IN2(g2051), .QN(n12203) );
  NAND2X0 U12455 ( .IN1(n12195), .IN2(g2028), .QN(n12202) );
  NAND4X0 U12456 ( .IN1(n12204), .IN2(n12205), .IN3(n12206), .IN4(n12200), 
        .QN(g32999) );
  INVX0 U12457 ( .INP(n3595), .ZN(n12200) );
  NAND3X0 U12458 ( .IN1(n5507), .IN2(n12207), .IN3(n3593), .QN(n12206) );
  NAND2X0 U12459 ( .IN1(n12201), .IN2(g2028), .QN(n12205) );
  NAND2X0 U12460 ( .IN1(test_so59), .IN2(n9420), .QN(n12204) );
  NAND4X0 U12461 ( .IN1(n12208), .IN2(n12209), .IN3(n12210), .IN4(n12211), 
        .QN(g32998) );
  NAND2X0 U12462 ( .IN1(n9506), .IN2(g1917), .QN(n12211) );
  NAND4X0 U12463 ( .IN1(n3604), .IN2(n11524), .IN3(n12212), .IN4(n8757), .QN(
        n12210) );
  NOR2X0 U12464 ( .IN1(n5510), .IN2(n12213), .QN(n12212) );
  NAND3X0 U12465 ( .IN1(n3605), .IN2(n12214), .IN3(n3611), .QN(n12209) );
  INVX0 U12466 ( .INP(n3607), .ZN(n12214) );
  NAND2X0 U12467 ( .IN1(n3524), .IN2(n10755), .QN(n3607) );
  INVX0 U12468 ( .INP(n3606), .ZN(n10755) );
  NAND3X0 U12469 ( .IN1(g1926), .IN2(g110), .IN3(n8757), .QN(n3605) );
  NAND2X0 U12470 ( .IN1(n12215), .IN2(g1932), .QN(n12208) );
  NAND3X0 U12471 ( .IN1(n12216), .IN2(n11526), .IN3(n12217), .QN(n12215) );
  NAND2X0 U12472 ( .IN1(n3606), .IN2(n9373), .QN(n12217) );
  NAND4X0 U12473 ( .IN1(n826), .IN2(n5349), .IN3(g2748), .IN4(n5300), .QN(
        n3606) );
  NAND4X0 U12474 ( .IN1(n12218), .IN2(n12219), .IN3(n12220), .IN4(n12221), 
        .QN(g32997) );
  NAND2X0 U12475 ( .IN1(n12222), .IN2(g1926), .QN(n12220) );
  NAND2X0 U12476 ( .IN1(n3611), .IN2(g1917), .QN(n12219) );
  NAND2X0 U12477 ( .IN1(n9507), .IN2(g1932), .QN(n12218) );
  NAND3X0 U12478 ( .IN1(n12223), .IN2(n12224), .IN3(n12221), .QN(g32996) );
  NAND2X0 U12479 ( .IN1(n12222), .IN2(g1917), .QN(n12224) );
  NAND2X0 U12480 ( .IN1(n12216), .IN2(g1894), .QN(n12223) );
  NAND4X0 U12481 ( .IN1(n12225), .IN2(n12226), .IN3(n12227), .IN4(n12221), 
        .QN(g32995) );
  INVX0 U12482 ( .INP(n3613), .ZN(n12221) );
  NAND3X0 U12483 ( .IN1(n5510), .IN2(n12228), .IN3(n3611), .QN(n12227) );
  NAND2X0 U12484 ( .IN1(n12222), .IN2(g1894), .QN(n12226) );
  NAND2X0 U12485 ( .IN1(n9507), .IN2(g1902), .QN(n12225) );
  NAND4X0 U12486 ( .IN1(n12229), .IN2(n12230), .IN3(n12231), .IN4(n12232), 
        .QN(g32994) );
  NAND2X0 U12487 ( .IN1(n9507), .IN2(g1783), .QN(n12232) );
  NAND4X0 U12488 ( .IN1(n3622), .IN2(n11524), .IN3(n12233), .IN4(n5596), .QN(
        n12231) );
  NOR2X0 U12489 ( .IN1(n5359), .IN2(n12234), .QN(n12233) );
  NAND3X0 U12490 ( .IN1(n3623), .IN2(n12235), .IN3(n3628), .QN(n12230) );
  INVX0 U12491 ( .INP(n3624), .ZN(n12235) );
  NAND2X0 U12492 ( .IN1(n3524), .IN2(n3005), .QN(n3624) );
  NAND3X0 U12493 ( .IN1(g1792), .IN2(g110), .IN3(n5596), .QN(n3623) );
  NAND2X0 U12494 ( .IN1(n12236), .IN2(g1798), .QN(n12229) );
  NAND3X0 U12495 ( .IN1(n12237), .IN2(n11526), .IN3(n12238), .QN(n12236) );
  NAND2X0 U12496 ( .IN1(n9365), .IN2(n1774), .QN(n12238) );
  INVX0 U12497 ( .INP(n3005), .ZN(n1774) );
  NAND4X0 U12498 ( .IN1(n12239), .IN2(n12240), .IN3(n12241), .IN4(n12242), 
        .QN(g32993) );
  NAND2X0 U12499 ( .IN1(n12243), .IN2(g1792), .QN(n12241) );
  NAND2X0 U12500 ( .IN1(n3628), .IN2(g1783), .QN(n12240) );
  NAND2X0 U12501 ( .IN1(n9507), .IN2(g1798), .QN(n12239) );
  NAND3X0 U12502 ( .IN1(n12244), .IN2(n12245), .IN3(n12242), .QN(g32992) );
  NAND2X0 U12503 ( .IN1(n12243), .IN2(g1783), .QN(n12245) );
  NAND2X0 U12504 ( .IN1(n12237), .IN2(g1760), .QN(n12244) );
  NAND4X0 U12505 ( .IN1(n12246), .IN2(n12247), .IN3(n12248), .IN4(n12242), 
        .QN(g32991) );
  INVX0 U12506 ( .INP(n3630), .ZN(n12242) );
  NAND3X0 U12507 ( .IN1(n5359), .IN2(n12249), .IN3(n3628), .QN(n12248) );
  NAND2X0 U12508 ( .IN1(n12243), .IN2(g1760), .QN(n12247) );
  NAND2X0 U12509 ( .IN1(n9507), .IN2(g1768), .QN(n12246) );
  NAND4X0 U12510 ( .IN1(n12250), .IN2(n12251), .IN3(n12252), .IN4(n12253), 
        .QN(g32990) );
  NAND2X0 U12511 ( .IN1(test_so94), .IN2(n9422), .QN(n12253) );
  NAND4X0 U12512 ( .IN1(n3640), .IN2(n11524), .IN3(n12254), .IN4(n8870), .QN(
        n12252) );
  NOR2X0 U12513 ( .IN1(n5525), .IN2(n12255), .QN(n12254) );
  NAND3X0 U12514 ( .IN1(n3641), .IN2(n12256), .IN3(n3646), .QN(n12251) );
  INVX0 U12515 ( .INP(n3642), .ZN(n12256) );
  NAND2X0 U12516 ( .IN1(n3524), .IN2(n10762), .QN(n3642) );
  INVX0 U12517 ( .INP(n3003), .ZN(n10762) );
  NAND3X0 U12518 ( .IN1(g110), .IN2(n8870), .IN3(g1657), .QN(n3641) );
  NAND2X0 U12519 ( .IN1(n12257), .IN2(g1664), .QN(n12250) );
  NAND3X0 U12520 ( .IN1(n11526), .IN2(n12258), .IN3(n12259), .QN(n12257) );
  NAND2X0 U12521 ( .IN1(n3003), .IN2(n9373), .QN(n12259) );
  NAND2X0 U12522 ( .IN1(n3653), .IN2(n826), .QN(n3003) );
  INVX0 U12523 ( .INP(n12260), .ZN(n826) );
  NAND2X0 U12524 ( .IN1(n12261), .IN2(n12262), .QN(n12260) );
  NAND2X0 U12525 ( .IN1(n12263), .IN2(n12264), .QN(n12262) );
  NAND2X0 U12526 ( .IN1(n8337), .IN2(n9794), .QN(n12264) );
  INVX0 U12527 ( .INP(g73), .ZN(n9794) );
  NAND2X0 U12528 ( .IN1(g73), .IN2(g2763), .QN(n12263) );
  NAND2X0 U12529 ( .IN1(n12265), .IN2(n12266), .QN(n12261) );
  NAND2X0 U12530 ( .IN1(n8336), .IN2(n9791), .QN(n12266) );
  INVX0 U12531 ( .INP(g72), .ZN(n9791) );
  NAND2X0 U12532 ( .IN1(g72), .IN2(g2759), .QN(n12265) );
  NAND2X0 U12533 ( .IN1(n9365), .IN2(n1835), .QN(n11526) );
  NAND4X0 U12534 ( .IN1(n12267), .IN2(n12268), .IN3(n12269), .IN4(n12270), 
        .QN(g32989) );
  NAND2X0 U12535 ( .IN1(n12271), .IN2(g1657), .QN(n12269) );
  NAND2X0 U12536 ( .IN1(n3646), .IN2(test_so94), .QN(n12268) );
  NAND2X0 U12537 ( .IN1(n9508), .IN2(g1664), .QN(n12267) );
  NAND3X0 U12538 ( .IN1(n12272), .IN2(n12273), .IN3(n12270), .QN(g32988) );
  NAND2X0 U12539 ( .IN1(n12271), .IN2(test_so94), .QN(n12273) );
  NAND2X0 U12540 ( .IN1(n12258), .IN2(g1624), .QN(n12272) );
  NAND4X0 U12541 ( .IN1(n12274), .IN2(n12275), .IN3(n12276), .IN4(n12270), 
        .QN(g32987) );
  INVX0 U12542 ( .INP(n3648), .ZN(n12270) );
  NAND3X0 U12543 ( .IN1(n5525), .IN2(n12277), .IN3(n3646), .QN(n12276) );
  NAND2X0 U12544 ( .IN1(n12271), .IN2(g1624), .QN(n12275) );
  NAND2X0 U12545 ( .IN1(n9507), .IN2(g1632), .QN(n12274) );
  NAND3X0 U12546 ( .IN1(n12278), .IN2(n12279), .IN3(n12280), .QN(g32986) );
  NAND3X0 U12547 ( .IN1(n11845), .IN2(n8455), .IN3(n12281), .QN(n12280) );
  INVX0 U12548 ( .INP(n12282), .ZN(n11845) );
  NAND3X0 U12549 ( .IN1(n12282), .IN2(g1373), .IN3(n9328), .QN(n12279) );
  NAND2X0 U12550 ( .IN1(n183), .IN2(n12283), .QN(n12282) );
  NAND2X0 U12551 ( .IN1(n8439), .IN2(n11847), .QN(n12283) );
  INVX0 U12552 ( .INP(n12284), .ZN(n183) );
  NAND2X0 U12553 ( .IN1(n9508), .IN2(g1367), .QN(n12278) );
  NOR2X0 U12554 ( .IN1(n5730), .IN2(n12285), .QN(g32985) );
  NOR2X0 U12555 ( .IN1(n9414), .IN2(n12286), .QN(n12285) );
  NOR2X0 U12556 ( .IN1(n10199), .IN2(n11854), .QN(n12286) );
  NAND2X0 U12557 ( .IN1(n3662), .IN2(g1270), .QN(n11854) );
  NAND3X0 U12558 ( .IN1(n12287), .IN2(n12288), .IN3(n12289), .QN(g32984) );
  NAND2X0 U12559 ( .IN1(n9509), .IN2(g1263), .QN(n12289) );
  NAND3X0 U12560 ( .IN1(n11853), .IN2(n12290), .IN3(g1270), .QN(n12288) );
  INVX0 U12561 ( .INP(n3662), .ZN(n12290) );
  NAND2X0 U12562 ( .IN1(n5716), .IN2(n3662), .QN(n12287) );
  NAND3X0 U12563 ( .IN1(n12291), .IN2(n12292), .IN3(n12293), .QN(g32983) );
  NAND3X0 U12564 ( .IN1(n11859), .IN2(n8457), .IN3(n12294), .QN(n12293) );
  INVX0 U12565 ( .INP(n12295), .ZN(n11859) );
  NAND3X0 U12566 ( .IN1(n12295), .IN2(g1030), .IN3(n9328), .QN(n12292) );
  NAND2X0 U12567 ( .IN1(n552), .IN2(n12296), .QN(n12295) );
  NAND2X0 U12568 ( .IN1(n8440), .IN2(n11861), .QN(n12296) );
  INVX0 U12569 ( .INP(n12297), .ZN(n552) );
  NAND2X0 U12570 ( .IN1(n9509), .IN2(g1024), .QN(n12291) );
  NOR2X0 U12571 ( .IN1(n5731), .IN2(n12298), .QN(g32982) );
  NOR2X0 U12572 ( .IN1(n9412), .IN2(n12299), .QN(n12298) );
  NOR2X0 U12573 ( .IN1(n10198), .IN2(n11868), .QN(n12299) );
  NAND2X0 U12574 ( .IN1(n3671), .IN2(g925), .QN(n11868) );
  NAND3X0 U12575 ( .IN1(n12300), .IN2(n12301), .IN3(n12302), .QN(g32981) );
  NAND2X0 U12576 ( .IN1(n9509), .IN2(g918), .QN(n12302) );
  NAND3X0 U12577 ( .IN1(n11867), .IN2(n12303), .IN3(g925), .QN(n12301) );
  INVX0 U12578 ( .INP(n3671), .ZN(n12303) );
  NAND2X0 U12579 ( .IN1(n5725), .IN2(n3671), .QN(n12300) );
  NOR3X0 U12580 ( .IN1(n9385), .IN2(n12304), .IN3(n12305), .QN(g32980) );
  NOR2X0 U12581 ( .IN1(n12306), .IN2(n10560), .QN(n12305) );
  INVX0 U12582 ( .INP(n2644), .ZN(n10560) );
  NOR2X0 U12583 ( .IN1(n10559), .IN2(g854), .QN(n12304) );
  INVX0 U12584 ( .INP(n12306), .ZN(n10559) );
  NAND4X0 U12585 ( .IN1(n5632), .IN2(g376), .IN3(g8719), .IN4(g370), .QN(
        n12306) );
  NAND3X0 U12586 ( .IN1(n12307), .IN2(n12308), .IN3(n12309), .QN(g32979) );
  NAND2X0 U12587 ( .IN1(test_so2), .IN2(n9418), .QN(n12309) );
  NAND3X0 U12588 ( .IN1(n2404), .IN2(n12310), .IN3(g758), .QN(n12308) );
  INVX0 U12589 ( .INP(n3272), .ZN(n12310) );
  NAND2X0 U12590 ( .IN1(n3272), .IN2(n5331), .QN(n12307) );
  NAND3X0 U12591 ( .IN1(n12311), .IN2(n12312), .IN3(n12313), .QN(g32978) );
  NAND2X0 U12592 ( .IN1(n9510), .IN2(g582), .QN(n12313) );
  NAND3X0 U12593 ( .IN1(n2421), .IN2(n12314), .IN3(g590), .QN(n12312) );
  INVX0 U12594 ( .INP(n3274), .ZN(n12314) );
  NAND2X0 U12595 ( .IN1(n3274), .IN2(n5472), .QN(n12311) );
  NAND3X0 U12596 ( .IN1(n12315), .IN2(n12316), .IN3(n12317), .QN(g32977) );
  NAND2X0 U12597 ( .IN1(test_so51), .IN2(n9513), .QN(n12317) );
  NAND3X0 U12598 ( .IN1(n10734), .IN2(n12318), .IN3(g291), .QN(n12316) );
  NAND2X0 U12599 ( .IN1(n54), .IN2(n5679), .QN(n12315) );
  INVX0 U12600 ( .INP(n12318), .ZN(n54) );
  NAND3X0 U12601 ( .IN1(test_so51), .IN2(n12319), .IN3(test_so55), .QN(n12318)
         );
  INVX0 U12602 ( .INP(n12320), .ZN(n12319) );
  NAND3X0 U12603 ( .IN1(n12321), .IN2(n12322), .IN3(n12323), .QN(g32976) );
  NAND2X0 U12604 ( .IN1(n9508), .IN2(g164), .QN(n12323) );
  NAND3X0 U12605 ( .IN1(n10739), .IN2(n12324), .IN3(g150), .QN(n12322) );
  INVX0 U12606 ( .INP(n3281), .ZN(n12324) );
  NAND2X0 U12607 ( .IN1(n3281), .IN2(n5676), .QN(n12321) );
  NOR4X0 U12608 ( .IN1(n12325), .IN2(n12326), .IN3(n12327), .IN4(n12328), .QN(
        g32185) );
  INVX0 U12609 ( .INP(n12329), .ZN(n12328) );
  NAND2X0 U12610 ( .IN1(g2902), .IN2(test_so1), .QN(n12329) );
  NOR2X0 U12611 ( .IN1(n8737), .IN2(n8736), .QN(n12327) );
  NOR2X0 U12612 ( .IN1(n8813), .IN2(n8894), .QN(n12326) );
  NAND4X0 U12613 ( .IN1(n12330), .IN2(n12331), .IN3(n12332), .IN4(n12333), 
        .QN(n12325) );
  NAND2X0 U12614 ( .IN1(g2975), .IN2(g2970), .QN(n12333) );
  NAND2X0 U12615 ( .IN1(g2950), .IN2(g2955), .QN(n12332) );
  NAND2X0 U12616 ( .IN1(g2912), .IN2(g2917), .QN(n12331) );
  NAND2X0 U12617 ( .IN1(g2922), .IN2(g2927), .QN(n12330) );
  NAND4X0 U12618 ( .IN1(n12334), .IN2(n12335), .IN3(n12336), .IN4(n12337), 
        .QN(g31904) );
  NAND4X0 U12619 ( .IN1(n12338), .IN2(n12339), .IN3(n12011), .IN4(g5033), .QN(
        n12337) );
  NAND2X0 U12620 ( .IN1(n8795), .IN2(n12340), .QN(n12336) );
  NAND2X0 U12621 ( .IN1(n9510), .IN2(g5029), .QN(n12335) );
  NAND2X0 U12622 ( .IN1(n12341), .IN2(n9373), .QN(n12334) );
  NAND4X0 U12623 ( .IN1(n12342), .IN2(n12009), .IN3(n12343), .IN4(n12344), 
        .QN(g31903) );
  NAND4X0 U12624 ( .IN1(n12345), .IN2(n12346), .IN3(n12011), .IN4(g5052), .QN(
        n12344) );
  INVX0 U12625 ( .INP(n12347), .ZN(n12346) );
  NAND2X0 U12626 ( .IN1(n5607), .IN2(n12012), .QN(n12343) );
  INVX0 U12627 ( .INP(n12345), .ZN(n12012) );
  NAND2X0 U12628 ( .IN1(n12348), .IN2(g5046), .QN(n12345) );
  NAND3X0 U12629 ( .IN1(n12347), .IN2(n9316), .IN3(n5607), .QN(n12009) );
  NAND2X0 U12630 ( .IN1(n9510), .IN2(g5046), .QN(n12342) );
  NAND3X0 U12631 ( .IN1(n12349), .IN2(n12350), .IN3(n12351), .QN(g31902) );
  NAND2X0 U12632 ( .IN1(n12352), .IN2(n9373), .QN(n12351) );
  NAND4X0 U12633 ( .IN1(n12011), .IN2(g5029), .IN3(n12353), .IN4(n12354), .QN(
        n12350) );
  NAND2X0 U12634 ( .IN1(n5369), .IN2(g5022), .QN(n12354) );
  NAND2X0 U12635 ( .IN1(g5016), .IN2(g5062), .QN(n12353) );
  NAND2X0 U12636 ( .IN1(n12355), .IN2(g5016), .QN(n12349) );
  NAND2X0 U12637 ( .IN1(n12356), .IN2(n9373), .QN(n12355) );
  NAND2X0 U12638 ( .IN1(n5601), .IN2(g5062), .QN(n12356) );
  NAND4X0 U12639 ( .IN1(n12357), .IN2(n12358), .IN3(n12359), .IN4(n12360), 
        .QN(g31901) );
  NAND4X0 U12640 ( .IN1(n12361), .IN2(n12362), .IN3(n12011), .IN4(g5046), .QN(
        n12360) );
  NAND2X0 U12641 ( .IN1(n12348), .IN2(n5578), .QN(n12359) );
  INVX0 U12642 ( .INP(n12362), .ZN(n12348) );
  NAND3X0 U12643 ( .IN1(g5041), .IN2(g5037), .IN3(n12363), .QN(n12362) );
  NAND2X0 U12644 ( .IN1(n9510), .IN2(g5041), .QN(n12358) );
  NAND2X0 U12645 ( .IN1(n12347), .IN2(n9373), .QN(n12357) );
  NOR2X0 U12646 ( .IN1(n12361), .IN2(g5046), .QN(n12347) );
  NAND3X0 U12647 ( .IN1(n5605), .IN2(n12341), .IN3(n5611), .QN(n12361) );
  NAND3X0 U12648 ( .IN1(n12364), .IN2(n12365), .IN3(n12366), .QN(g31900) );
  INVX0 U12649 ( .INP(n12367), .ZN(n12366) );
  NOR2X0 U12650 ( .IN1(n12368), .IN2(g5041), .QN(n12367) );
  NAND4X0 U12651 ( .IN1(n12369), .IN2(g5041), .IN3(n12011), .IN4(n5611), .QN(
        n12365) );
  NAND2X0 U12652 ( .IN1(n12370), .IN2(g5037), .QN(n12364) );
  NAND3X0 U12653 ( .IN1(n12371), .IN2(n12372), .IN3(n9329), .QN(n12370) );
  NAND3X0 U12654 ( .IN1(n12373), .IN2(n12374), .IN3(g5041), .QN(n12372) );
  INVX0 U12655 ( .INP(n12375), .ZN(n12373) );
  NAND2X0 U12656 ( .IN1(n5605), .IN2(n12363), .QN(n12371) );
  NAND4X0 U12657 ( .IN1(n12376), .IN2(n12368), .IN3(n12377), .IN4(n12378), 
        .QN(g31899) );
  NAND4X0 U12658 ( .IN1(n12369), .IN2(n12374), .IN3(n12011), .IN4(g5037), .QN(
        n12378) );
  NAND2X0 U12659 ( .IN1(n5611), .IN2(n12363), .QN(n12377) );
  INVX0 U12660 ( .INP(n12374), .ZN(n12363) );
  NAND2X0 U12661 ( .IN1(n12340), .IN2(g5033), .QN(n12374) );
  INVX0 U12662 ( .INP(n12339), .ZN(n12340) );
  NAND3X0 U12663 ( .IN1(g5029), .IN2(g5062), .IN3(g5016), .QN(n12339) );
  NAND3X0 U12664 ( .IN1(n12341), .IN2(n9316), .IN3(n5611), .QN(n12368) );
  INVX0 U12665 ( .INP(n12369), .ZN(n12341) );
  NAND2X0 U12666 ( .IN1(n8795), .IN2(n12352), .QN(n12369) );
  INVX0 U12667 ( .INP(n12338), .ZN(n12352) );
  NAND3X0 U12668 ( .IN1(n5369), .IN2(g5022), .IN3(n5601), .QN(n12338) );
  NAND2X0 U12669 ( .IN1(n9508), .IN2(g5033), .QN(n12376) );
  NAND3X0 U12670 ( .IN1(n12379), .IN2(n12380), .IN3(n12381), .QN(g31898) );
  NAND3X0 U12671 ( .IN1(n12011), .IN2(n12382), .IN3(n5369), .QN(n12381) );
  INVX0 U12672 ( .INP(n12383), .ZN(n12382) );
  NOR2X0 U12673 ( .IN1(n12375), .IN2(n9397), .QN(n12011) );
  NAND2X0 U12674 ( .IN1(n12384), .IN2(n12385), .QN(n12375) );
  NAND3X0 U12675 ( .IN1(n12383), .IN2(g5016), .IN3(n9329), .QN(n12380) );
  NOR2X0 U12676 ( .IN1(g5062), .IN2(g5022), .QN(n12383) );
  NAND2X0 U12677 ( .IN1(n9509), .IN2(g5022), .QN(n12379) );
  NAND3X0 U12678 ( .IN1(n12386), .IN2(n11451), .IN3(n12387), .QN(g31897) );
  NAND2X0 U12679 ( .IN1(n12020), .IN2(g4575), .QN(n11451) );
  NAND2X0 U12680 ( .IN1(n9508), .IN2(g4423), .QN(n12386) );
  NAND3X0 U12681 ( .IN1(n12388), .IN2(n11456), .IN3(n12387), .QN(g31896) );
  INVX0 U12682 ( .INP(n12389), .ZN(n12387) );
  NAND2X0 U12683 ( .IN1(n12390), .IN2(n12391), .QN(n12389) );
  NAND2X0 U12684 ( .IN1(n12020), .IN2(n12392), .QN(n12391) );
  NAND2X0 U12685 ( .IN1(g72), .IN2(g73), .QN(n12392) );
  NAND2X0 U12686 ( .IN1(n11457), .IN2(g4372), .QN(n12390) );
  INVX0 U12687 ( .INP(n12393), .ZN(n11457) );
  NAND2X0 U12688 ( .IN1(n12020), .IN2(test_so100), .QN(n11456) );
  NOR2X0 U12689 ( .IN1(n9418), .IN2(n5670), .QN(n12020) );
  INVX0 U12690 ( .INP(n12394), .ZN(n12388) );
  NOR2X0 U12691 ( .IN1(n9358), .IN2(n5849), .QN(n12394) );
  NAND2X0 U12692 ( .IN1(n10505), .IN2(n12395), .QN(g31895) );
  NAND2X0 U12693 ( .IN1(n9510), .IN2(g4382), .QN(n12395) );
  INVX0 U12694 ( .INP(n11524), .ZN(n10505) );
  NOR2X0 U12695 ( .IN1(n1835), .IN2(n9396), .QN(n11524) );
  INVX0 U12696 ( .INP(n2760), .ZN(n1835) );
  NAND3X0 U12697 ( .IN1(n12396), .IN2(n12032), .IN3(n12397), .QN(g31894) );
  NAND2X0 U12698 ( .IN1(n12398), .IN2(g4093), .QN(n12397) );
  NAND2X0 U12699 ( .IN1(n12399), .IN2(n9377), .QN(n12398) );
  NAND2X0 U12700 ( .IN1(n12035), .IN2(n9773), .QN(n12399) );
  NAND3X0 U12701 ( .IN1(n9349), .IN2(g4098), .IN3(n12035), .QN(n12396) );
  NAND3X0 U12702 ( .IN1(g4093), .IN2(g4098), .IN3(n9773), .QN(n12035) );
  NOR2X0 U12703 ( .IN1(n12400), .IN2(n5480), .QN(n9773) );
  NAND2X0 U12704 ( .IN1(n12401), .IN2(n12402), .QN(g31872) );
  NAND3X0 U12705 ( .IN1(n12403), .IN2(n12404), .IN3(n3730), .QN(n12402) );
  NAND2X0 U12706 ( .IN1(n5516), .IN2(n12405), .QN(n12404) );
  INVX0 U12707 ( .INP(n12406), .ZN(n12403) );
  NOR2X0 U12708 ( .IN1(n12405), .IN2(n5516), .QN(n12406) );
  NAND2X0 U12709 ( .IN1(n9507), .IN2(g2741), .QN(n12401) );
  NAND3X0 U12710 ( .IN1(n12407), .IN2(n12408), .IN3(n12409), .QN(g31871) );
  NAND2X0 U12711 ( .IN1(n3733), .IN2(n12281), .QN(n12409) );
  NAND2X0 U12712 ( .IN1(n9510), .IN2(g1361), .QN(n12408) );
  NAND3X0 U12713 ( .IN1(n12284), .IN2(g1367), .IN3(n9329), .QN(n12407) );
  NAND2X0 U12714 ( .IN1(n184), .IN2(n12410), .QN(n12284) );
  NAND2X0 U12715 ( .IN1(n8454), .IN2(n11847), .QN(n12410) );
  INVX0 U12716 ( .INP(n12411), .ZN(n184) );
  NAND3X0 U12717 ( .IN1(n12412), .IN2(n12413), .IN3(n12414), .QN(g31870) );
  NAND2X0 U12718 ( .IN1(n9509), .IN2(g1259), .QN(n12414) );
  NAND3X0 U12719 ( .IN1(n11853), .IN2(n12415), .IN3(g1263), .QN(n12413) );
  INVX0 U12720 ( .INP(n3664), .ZN(n12415) );
  NAND2X0 U12721 ( .IN1(n3664), .IN2(n5674), .QN(n12412) );
  NAND3X0 U12722 ( .IN1(n12416), .IN2(n12417), .IN3(n12418), .QN(g31869) );
  NAND2X0 U12723 ( .IN1(n3738), .IN2(n12294), .QN(n12418) );
  NAND2X0 U12724 ( .IN1(n9511), .IN2(g1018), .QN(n12417) );
  NAND3X0 U12725 ( .IN1(n12297), .IN2(g1024), .IN3(n9329), .QN(n12416) );
  NAND2X0 U12726 ( .IN1(n553), .IN2(n12419), .QN(n12297) );
  NAND2X0 U12727 ( .IN1(n8456), .IN2(n11861), .QN(n12419) );
  INVX0 U12728 ( .INP(n12420), .ZN(n553) );
  NAND3X0 U12729 ( .IN1(n12421), .IN2(n12422), .IN3(n12423), .QN(g31868) );
  NAND2X0 U12730 ( .IN1(n9511), .IN2(g914), .QN(n12423) );
  NAND3X0 U12731 ( .IN1(n11867), .IN2(n12424), .IN3(g918), .QN(n12422) );
  INVX0 U12732 ( .INP(n3673), .ZN(n12424) );
  NAND2X0 U12733 ( .IN1(n3673), .IN2(n5673), .QN(n12421) );
  NAND3X0 U12734 ( .IN1(n12425), .IN2(n12426), .IN3(n12427), .QN(g31867) );
  NAND2X0 U12735 ( .IN1(n9509), .IN2(g744), .QN(n12427) );
  NAND3X0 U12736 ( .IN1(n2404), .IN2(test_so2), .IN3(n12428), .QN(n12426) );
  INVX0 U12737 ( .INP(n12429), .ZN(n12425) );
  NOR2X0 U12738 ( .IN1(n12428), .IN2(test_so2), .QN(n12429) );
  INVX0 U12739 ( .INP(n3682), .ZN(n12428) );
  NAND3X0 U12740 ( .IN1(n12430), .IN2(n12431), .IN3(n12432), .QN(g31866) );
  NAND2X0 U12741 ( .IN1(n9508), .IN2(g577), .QN(n12432) );
  NAND3X0 U12742 ( .IN1(n2421), .IN2(n12433), .IN3(g582), .QN(n12431) );
  INVX0 U12743 ( .INP(n3684), .ZN(n12433) );
  NAND2X0 U12744 ( .IN1(n3684), .IN2(n5552), .QN(n12430) );
  NAND2X0 U12745 ( .IN1(n12434), .IN2(n12435), .QN(g31865) );
  INVX0 U12746 ( .INP(n12436), .ZN(n12435) );
  NOR2X0 U12747 ( .IN1(n8874), .IN2(n12437), .QN(n12436) );
  NOR2X0 U12748 ( .IN1(n12438), .IN2(n9510), .QN(n12437) );
  NOR2X0 U12749 ( .IN1(n12320), .IN2(test_so51), .QN(n12438) );
  NAND3X0 U12750 ( .IN1(n10734), .IN2(test_so51), .IN3(n8874), .QN(n12434) );
  NAND3X0 U12751 ( .IN1(n12439), .IN2(n12440), .IN3(n12441), .QN(g31864) );
  NAND2X0 U12752 ( .IN1(test_so73), .IN2(n9516), .QN(n12441) );
  NAND3X0 U12753 ( .IN1(n10739), .IN2(n12442), .IN3(g164), .QN(n12440) );
  INVX0 U12754 ( .INP(n3687), .ZN(n12442) );
  NAND2X0 U12755 ( .IN1(n3687), .IN2(n5561), .QN(n12439) );
  NOR3X0 U12756 ( .IN1(n12443), .IN2(n12444), .IN3(n8883), .QN(n3687) );
  NAND2X0 U12757 ( .IN1(n12445), .IN2(n12446), .QN(g31793) );
  NAND2X0 U12758 ( .IN1(n12447), .IN2(n10229), .QN(n12446) );
  NAND2X0 U12759 ( .IN1(n12448), .IN2(n9369), .QN(n12447) );
  NAND2X0 U12760 ( .IN1(n10228), .IN2(n12449), .QN(n12448) );
  NAND2X0 U12761 ( .IN1(n12450), .IN2(n12451), .QN(n12449) );
  NAND3X0 U12762 ( .IN1(n12452), .IN2(n12453), .IN3(n8356), .QN(n12451) );
  NAND2X0 U12763 ( .IN1(g6509), .IN2(n12454), .QN(n12453) );
  NAND4X0 U12764 ( .IN1(n8463), .IN2(n8462), .IN3(n8395), .IN4(n12455), .QN(
        n12450) );
  NAND2X0 U12765 ( .IN1(n12456), .IN2(n12457), .QN(n12455) );
  NAND3X0 U12766 ( .IN1(n12458), .IN2(n12459), .IN3(n8356), .QN(n12456) );
  NAND2X0 U12767 ( .IN1(n12460), .IN2(g6163), .QN(n12459) );
  NAND2X0 U12768 ( .IN1(g5817), .IN2(g5471), .QN(n12458) );
  INVX0 U12769 ( .INP(n12461), .ZN(n10228) );
  NAND3X0 U12770 ( .IN1(n12462), .IN2(n12463), .IN3(n10230), .QN(n12445) );
  NOR4X0 U12771 ( .IN1(g5124), .IN2(n12457), .IN3(g6509), .IN4(n12454), .QN(
        n10230) );
  NAND2X0 U12772 ( .IN1(n8463), .IN2(n8462), .QN(n12454) );
  INVX0 U12773 ( .INP(n12452), .ZN(n12457) );
  NOR2X0 U12774 ( .IN1(g6163), .IN2(n12460), .QN(n12452) );
  NAND2X0 U12775 ( .IN1(n8365), .IN2(n8358), .QN(n12460) );
  NAND2X0 U12776 ( .IN1(n12464), .IN2(n12461), .QN(n12463) );
  NAND2X0 U12777 ( .IN1(n8394), .IN2(n8374), .QN(n12461) );
  NAND2X0 U12778 ( .IN1(g3466), .IN2(g3115), .QN(n12462) );
  NAND2X0 U12779 ( .IN1(g113), .IN2(g2868), .QN(g31665) );
  NAND2X0 U12780 ( .IN1(g113), .IN2(g2873), .QN(g31656) );
  NAND3X0 U12781 ( .IN1(n12465), .IN2(n12466), .IN3(n12467), .QN(g30563) );
  NAND2X0 U12782 ( .IN1(n9510), .IN2(g6653), .QN(n12467) );
  NAND2X0 U12783 ( .IN1(n12468), .IN2(g6657), .QN(n12466) );
  NAND2X0 U12784 ( .IN1(n3765), .IN2(n11370), .QN(n12465) );
  NAND3X0 U12785 ( .IN1(n12469), .IN2(n12470), .IN3(n12471), .QN(g30562) );
  NAND2X0 U12786 ( .IN1(n12472), .IN2(n3765), .QN(n12471) );
  NAND3X0 U12787 ( .IN1(n12473), .IN2(g6605), .IN3(n9329), .QN(n12470) );
  INVX0 U12788 ( .INP(n12472), .ZN(n12473) );
  NOR2X0 U12789 ( .IN1(n1452), .IN2(n5646), .QN(n12472) );
  INVX0 U12790 ( .INP(n11907), .ZN(n1452) );
  NAND2X0 U12791 ( .IN1(n9508), .IN2(g6649), .QN(n12469) );
  NAND3X0 U12792 ( .IN1(n12474), .IN2(n12475), .IN3(n12476), .QN(g30561) );
  NAND2X0 U12793 ( .IN1(n12477), .IN2(n3765), .QN(n12476) );
  NAND3X0 U12794 ( .IN1(n11905), .IN2(g6597), .IN3(n9329), .QN(n12475) );
  INVX0 U12795 ( .INP(n12477), .ZN(n11905) );
  NOR2X0 U12796 ( .IN1(n1456), .IN2(n5646), .QN(n12477) );
  INVX0 U12797 ( .INP(n12478), .ZN(n1456) );
  NAND2X0 U12798 ( .IN1(n9501), .IN2(g6645), .QN(n12474) );
  NAND3X0 U12799 ( .IN1(n12479), .IN2(n12480), .IN3(n12481), .QN(g30560) );
  NAND2X0 U12800 ( .IN1(n12482), .IN2(n3765), .QN(n12481) );
  NAND3X0 U12801 ( .IN1(n12483), .IN2(g6589), .IN3(n9329), .QN(n12480) );
  INVX0 U12802 ( .INP(n12482), .ZN(n12483) );
  NOR2X0 U12803 ( .IN1(n1454), .IN2(n5646), .QN(n12482) );
  INVX0 U12804 ( .INP(n12484), .ZN(n1454) );
  NAND2X0 U12805 ( .IN1(n9501), .IN2(g6641), .QN(n12479) );
  NAND3X0 U12806 ( .IN1(n12485), .IN2(n12486), .IN3(n12487), .QN(g30559) );
  NAND2X0 U12807 ( .IN1(n3774), .IN2(n9806), .QN(n12487) );
  NAND2X0 U12808 ( .IN1(n9501), .IN2(g6637), .QN(n12486) );
  NAND3X0 U12809 ( .IN1(n12488), .IN2(g6653), .IN3(n9329), .QN(n12485) );
  NAND2X0 U12810 ( .IN1(n9806), .IN2(n9666), .QN(n12488) );
  NAND3X0 U12811 ( .IN1(n12489), .IN2(n12490), .IN3(n12491), .QN(g30558) );
  NAND2X0 U12812 ( .IN1(n3774), .IN2(n11907), .QN(n12491) );
  NAND2X0 U12813 ( .IN1(n9500), .IN2(g6633), .QN(n12490) );
  NAND3X0 U12814 ( .IN1(n12492), .IN2(g6649), .IN3(n9330), .QN(n12489) );
  NAND2X0 U12815 ( .IN1(n11907), .IN2(n9666), .QN(n12492) );
  NAND3X0 U12816 ( .IN1(n12493), .IN2(n12494), .IN3(n12495), .QN(g30557) );
  NAND2X0 U12817 ( .IN1(n3774), .IN2(n12478), .QN(n12495) );
  NAND2X0 U12818 ( .IN1(n9500), .IN2(g6629), .QN(n12494) );
  NAND3X0 U12819 ( .IN1(n12496), .IN2(g6645), .IN3(n9330), .QN(n12493) );
  NAND2X0 U12820 ( .IN1(n12478), .IN2(n9666), .QN(n12496) );
  NAND3X0 U12821 ( .IN1(n12497), .IN2(n12498), .IN3(n12499), .QN(g30556) );
  NAND2X0 U12822 ( .IN1(n3774), .IN2(n12484), .QN(n12499) );
  NAND2X0 U12823 ( .IN1(n9500), .IN2(g6625), .QN(n12498) );
  NAND3X0 U12824 ( .IN1(n12500), .IN2(g6641), .IN3(n9330), .QN(n12497) );
  NAND2X0 U12825 ( .IN1(n12484), .IN2(n9666), .QN(n12500) );
  NOR2X0 U12826 ( .IN1(n5571), .IN2(n8772), .QN(n9666) );
  NAND3X0 U12827 ( .IN1(n12501), .IN2(n12502), .IN3(n12503), .QN(g30555) );
  NAND2X0 U12828 ( .IN1(n3780), .IN2(n9806), .QN(n12503) );
  NAND2X0 U12829 ( .IN1(n9500), .IN2(g6621), .QN(n12502) );
  NAND3X0 U12830 ( .IN1(n12504), .IN2(g6637), .IN3(n9330), .QN(n12501) );
  NAND2X0 U12831 ( .IN1(n9806), .IN2(n9665), .QN(n12504) );
  NAND3X0 U12832 ( .IN1(n12505), .IN2(n12506), .IN3(n12507), .QN(g30554) );
  NAND2X0 U12833 ( .IN1(n3780), .IN2(n11907), .QN(n12507) );
  NAND2X0 U12834 ( .IN1(n9500), .IN2(g6617), .QN(n12506) );
  NAND3X0 U12835 ( .IN1(n12508), .IN2(g6633), .IN3(n9330), .QN(n12505) );
  NAND2X0 U12836 ( .IN1(n11907), .IN2(n9665), .QN(n12508) );
  NAND3X0 U12837 ( .IN1(n12509), .IN2(n12510), .IN3(n12511), .QN(g30553) );
  NAND2X0 U12838 ( .IN1(n3780), .IN2(n12478), .QN(n12511) );
  NAND2X0 U12839 ( .IN1(n9500), .IN2(g6613), .QN(n12510) );
  NAND3X0 U12840 ( .IN1(n12512), .IN2(g6629), .IN3(n9330), .QN(n12509) );
  NAND2X0 U12841 ( .IN1(n12478), .IN2(n9665), .QN(n12512) );
  NAND3X0 U12842 ( .IN1(n12513), .IN2(n12514), .IN3(n12515), .QN(g30552) );
  NAND2X0 U12843 ( .IN1(n3780), .IN2(n12484), .QN(n12515) );
  NAND2X0 U12844 ( .IN1(n9500), .IN2(g6609), .QN(n12514) );
  NAND3X0 U12845 ( .IN1(n12516), .IN2(g6625), .IN3(n9330), .QN(n12513) );
  NAND2X0 U12846 ( .IN1(n12484), .IN2(n9665), .QN(n12516) );
  NOR2X0 U12847 ( .IN1(g6549), .IN2(n8772), .QN(n9665) );
  NAND3X0 U12848 ( .IN1(n12517), .IN2(n12518), .IN3(n12519), .QN(g30551) );
  NAND2X0 U12849 ( .IN1(n3785), .IN2(n9806), .QN(n12519) );
  NAND2X0 U12850 ( .IN1(n9499), .IN2(g6601), .QN(n12518) );
  NAND3X0 U12851 ( .IN1(n12520), .IN2(g6621), .IN3(n9330), .QN(n12517) );
  NAND2X0 U12852 ( .IN1(n9806), .IN2(n11920), .QN(n12520) );
  NAND3X0 U12853 ( .IN1(n12521), .IN2(n12522), .IN3(n12523), .QN(g30550) );
  NAND2X0 U12854 ( .IN1(n3785), .IN2(n11907), .QN(n12523) );
  NAND2X0 U12855 ( .IN1(n9499), .IN2(g6593), .QN(n12522) );
  NAND3X0 U12856 ( .IN1(n12524), .IN2(g6617), .IN3(n9330), .QN(n12521) );
  NAND2X0 U12857 ( .IN1(n11907), .IN2(n11920), .QN(n12524) );
  NOR2X0 U12858 ( .IN1(g6565), .IN2(n5563), .QN(n11907) );
  NAND3X0 U12859 ( .IN1(n12525), .IN2(n12526), .IN3(n12527), .QN(g30549) );
  NAND2X0 U12860 ( .IN1(n3785), .IN2(n12478), .QN(n12527) );
  NAND2X0 U12861 ( .IN1(test_so71), .IN2(n9514), .QN(n12526) );
  NAND3X0 U12862 ( .IN1(n12528), .IN2(g6613), .IN3(n9330), .QN(n12525) );
  NAND2X0 U12863 ( .IN1(n12478), .IN2(n11920), .QN(n12528) );
  NOR2X0 U12864 ( .IN1(g6573), .IN2(n5386), .QN(n12478) );
  NAND3X0 U12865 ( .IN1(n12529), .IN2(n12530), .IN3(n12531), .QN(g30548) );
  NAND2X0 U12866 ( .IN1(n3785), .IN2(n12484), .QN(n12531) );
  NAND2X0 U12867 ( .IN1(n9499), .IN2(g6581), .QN(n12530) );
  NAND3X0 U12868 ( .IN1(n12532), .IN2(g6609), .IN3(n9330), .QN(n12529) );
  NAND2X0 U12869 ( .IN1(n12484), .IN2(n11920), .QN(n12532) );
  NOR2X0 U12870 ( .IN1(g6555), .IN2(n5571), .QN(n11920) );
  NOR2X0 U12871 ( .IN1(g6565), .IN2(g6573), .QN(n12484) );
  NAND3X0 U12872 ( .IN1(n12533), .IN2(n12534), .IN3(n12535), .QN(g30547) );
  NAND2X0 U12873 ( .IN1(n9499), .IN2(g6605), .QN(n12535) );
  NAND3X0 U12874 ( .IN1(n9349), .IN2(g6601), .IN3(n12536), .QN(n12534) );
  INVX0 U12875 ( .INP(n3790), .ZN(n12536) );
  NAND2X0 U12876 ( .IN1(n3790), .IN2(n3765), .QN(n12533) );
  NAND3X0 U12877 ( .IN1(n12537), .IN2(n12538), .IN3(n12539), .QN(g30546) );
  NAND2X0 U12878 ( .IN1(n9499), .IN2(g6597), .QN(n12539) );
  NAND3X0 U12879 ( .IN1(n9349), .IN2(g6593), .IN3(n12540), .QN(n12538) );
  INVX0 U12880 ( .INP(n3793), .ZN(n12540) );
  NAND2X0 U12881 ( .IN1(n3793), .IN2(n3765), .QN(n12537) );
  NAND3X0 U12882 ( .IN1(n12541), .IN2(n12542), .IN3(n12543), .QN(g30545) );
  NAND2X0 U12883 ( .IN1(n9499), .IN2(g6589), .QN(n12543) );
  NAND3X0 U12884 ( .IN1(test_so71), .IN2(n9315), .IN3(n12544), .QN(n12542) );
  INVX0 U12885 ( .INP(n3795), .ZN(n12544) );
  NAND2X0 U12886 ( .IN1(n3795), .IN2(n3765), .QN(n12541) );
  NAND3X0 U12887 ( .IN1(n12545), .IN2(n12546), .IN3(n12547), .QN(g30544) );
  NAND2X0 U12888 ( .IN1(n9499), .IN2(g6573), .QN(n12547) );
  NAND3X0 U12889 ( .IN1(n9347), .IN2(g6581), .IN3(n12548), .QN(n12546) );
  INVX0 U12890 ( .INP(n3797), .ZN(n12548) );
  NAND2X0 U12891 ( .IN1(n3797), .IN2(n3765), .QN(n12545) );
  NOR2X0 U12892 ( .IN1(g6549), .IN2(n11913), .QN(g30543) );
  NAND3X0 U12893 ( .IN1(n11903), .IN2(n9316), .IN3(n5646), .QN(n11913) );
  NAND2X0 U12894 ( .IN1(n3799), .IN2(n11360), .QN(n11903) );
  NAND3X0 U12895 ( .IN1(n12549), .IN2(n12550), .IN3(n12551), .QN(g30542) );
  NAND2X0 U12896 ( .IN1(n9498), .IN2(g6307), .QN(n12551) );
  NAND2X0 U12897 ( .IN1(n12552), .IN2(g6311), .QN(n12550) );
  NAND2X0 U12898 ( .IN1(n12553), .IN2(n3765), .QN(n12549) );
  NAND3X0 U12899 ( .IN1(n12554), .IN2(n12555), .IN3(n12556), .QN(g30541) );
  NAND2X0 U12900 ( .IN1(n12557), .IN2(n3765), .QN(n12556) );
  NAND3X0 U12901 ( .IN1(n12558), .IN2(g6259), .IN3(n9330), .QN(n12555) );
  INVX0 U12902 ( .INP(n12557), .ZN(n12558) );
  NOR2X0 U12903 ( .IN1(n47), .IN2(n5651), .QN(n12557) );
  INVX0 U12904 ( .INP(n11928), .ZN(n47) );
  NAND2X0 U12905 ( .IN1(n9498), .IN2(g6303), .QN(n12554) );
  NAND3X0 U12906 ( .IN1(n12559), .IN2(n12560), .IN3(n12561), .QN(g30540) );
  NAND2X0 U12907 ( .IN1(n12562), .IN2(n3765), .QN(n12561) );
  NAND3X0 U12908 ( .IN1(n11926), .IN2(g6251), .IN3(n9331), .QN(n12560) );
  INVX0 U12909 ( .INP(n12562), .ZN(n11926) );
  NOR2X0 U12910 ( .IN1(n43), .IN2(n5651), .QN(n12562) );
  INVX0 U12911 ( .INP(n12563), .ZN(n43) );
  NAND2X0 U12912 ( .IN1(n9498), .IN2(g6299), .QN(n12559) );
  NAND3X0 U12913 ( .IN1(n12564), .IN2(n12565), .IN3(n12566), .QN(g30539) );
  NAND2X0 U12914 ( .IN1(n12567), .IN2(n3765), .QN(n12566) );
  NAND3X0 U12915 ( .IN1(n12568), .IN2(g6243), .IN3(n9331), .QN(n12565) );
  INVX0 U12916 ( .INP(n12567), .ZN(n12568) );
  NOR2X0 U12917 ( .IN1(n45), .IN2(n5651), .QN(n12567) );
  INVX0 U12918 ( .INP(n12569), .ZN(n45) );
  NAND2X0 U12919 ( .IN1(n9498), .IN2(g6295), .QN(n12564) );
  NAND3X0 U12920 ( .IN1(n12570), .IN2(n12571), .IN3(n12572), .QN(g30538) );
  NAND2X0 U12921 ( .IN1(n3808), .IN2(n12573), .QN(n12572) );
  NAND2X0 U12922 ( .IN1(n9498), .IN2(g6291), .QN(n12571) );
  NAND3X0 U12923 ( .IN1(n12574), .IN2(g6307), .IN3(n9331), .QN(n12570) );
  NAND2X0 U12924 ( .IN1(n9815), .IN2(n12573), .QN(n12574) );
  NAND3X0 U12925 ( .IN1(n12575), .IN2(n12576), .IN3(n12577), .QN(g30537) );
  NAND2X0 U12926 ( .IN1(n3808), .IN2(n11928), .QN(n12577) );
  NAND2X0 U12927 ( .IN1(n9498), .IN2(g6287), .QN(n12576) );
  NAND3X0 U12928 ( .IN1(n12578), .IN2(g6303), .IN3(n9331), .QN(n12575) );
  NAND2X0 U12929 ( .IN1(n9815), .IN2(n11928), .QN(n12578) );
  NAND3X0 U12930 ( .IN1(n12579), .IN2(n12580), .IN3(n12581), .QN(g30536) );
  NAND2X0 U12931 ( .IN1(n3808), .IN2(n12563), .QN(n12581) );
  NAND2X0 U12932 ( .IN1(n9498), .IN2(g6283), .QN(n12580) );
  NAND3X0 U12933 ( .IN1(n12582), .IN2(g6299), .IN3(n9331), .QN(n12579) );
  NAND2X0 U12934 ( .IN1(n9815), .IN2(n12563), .QN(n12582) );
  NAND3X0 U12935 ( .IN1(n12583), .IN2(n12584), .IN3(n12585), .QN(g30535) );
  NAND2X0 U12936 ( .IN1(n3808), .IN2(n12569), .QN(n12585) );
  NAND2X0 U12937 ( .IN1(n9497), .IN2(g6279), .QN(n12584) );
  NAND3X0 U12938 ( .IN1(n12586), .IN2(g6295), .IN3(n9331), .QN(n12583) );
  NAND2X0 U12939 ( .IN1(n9815), .IN2(n12569), .QN(n12586) );
  NOR2X0 U12940 ( .IN1(n5574), .IN2(n8768), .QN(n9815) );
  NAND3X0 U12941 ( .IN1(n12587), .IN2(n12588), .IN3(n12589), .QN(g30534) );
  NAND2X0 U12942 ( .IN1(n3814), .IN2(n12573), .QN(n12589) );
  NAND2X0 U12943 ( .IN1(n9497), .IN2(g6275), .QN(n12588) );
  NAND3X0 U12944 ( .IN1(n12590), .IN2(g6291), .IN3(n9331), .QN(n12587) );
  NAND2X0 U12945 ( .IN1(n9814), .IN2(n12573), .QN(n12590) );
  NAND3X0 U12946 ( .IN1(n12591), .IN2(n12592), .IN3(n12593), .QN(g30533) );
  NAND2X0 U12947 ( .IN1(n3814), .IN2(n11928), .QN(n12593) );
  NAND2X0 U12948 ( .IN1(n9497), .IN2(g6271), .QN(n12592) );
  NAND3X0 U12949 ( .IN1(n12594), .IN2(g6287), .IN3(n9331), .QN(n12591) );
  NAND2X0 U12950 ( .IN1(n9814), .IN2(n11928), .QN(n12594) );
  NAND3X0 U12951 ( .IN1(n12595), .IN2(n12596), .IN3(n12597), .QN(g30532) );
  NAND2X0 U12952 ( .IN1(n3814), .IN2(n12563), .QN(n12597) );
  NAND2X0 U12953 ( .IN1(n9497), .IN2(g6267), .QN(n12596) );
  NAND3X0 U12954 ( .IN1(n12598), .IN2(g6283), .IN3(n9331), .QN(n12595) );
  NAND2X0 U12955 ( .IN1(n9814), .IN2(n12563), .QN(n12598) );
  NAND3X0 U12956 ( .IN1(n12599), .IN2(n12600), .IN3(n12601), .QN(g30531) );
  NAND2X0 U12957 ( .IN1(n3814), .IN2(n12569), .QN(n12601) );
  NAND2X0 U12958 ( .IN1(n9497), .IN2(g6263), .QN(n12600) );
  NAND3X0 U12959 ( .IN1(n12602), .IN2(g6279), .IN3(n9331), .QN(n12599) );
  NAND2X0 U12960 ( .IN1(n9814), .IN2(n12569), .QN(n12602) );
  NOR2X0 U12961 ( .IN1(g6203), .IN2(n8768), .QN(n9814) );
  NAND3X0 U12962 ( .IN1(n12603), .IN2(n12604), .IN3(n12605), .QN(g30530) );
  NAND2X0 U12963 ( .IN1(n3819), .IN2(n12573), .QN(n12605) );
  NAND2X0 U12964 ( .IN1(n9497), .IN2(g6255), .QN(n12604) );
  NAND3X0 U12965 ( .IN1(n12606), .IN2(g6275), .IN3(n9331), .QN(n12603) );
  NAND2X0 U12966 ( .IN1(n11941), .IN2(n12573), .QN(n12606) );
  NAND3X0 U12967 ( .IN1(n12607), .IN2(n12608), .IN3(n12609), .QN(g30529) );
  NAND2X0 U12968 ( .IN1(n3819), .IN2(n11928), .QN(n12609) );
  NAND2X0 U12969 ( .IN1(n9497), .IN2(g6247), .QN(n12608) );
  NAND3X0 U12970 ( .IN1(n12610), .IN2(g6271), .IN3(n9331), .QN(n12607) );
  NAND2X0 U12971 ( .IN1(n11941), .IN2(n11928), .QN(n12610) );
  NOR2X0 U12972 ( .IN1(g6219), .IN2(n5568), .QN(n11928) );
  NAND3X0 U12973 ( .IN1(n12611), .IN2(n12612), .IN3(n12613), .QN(g30528) );
  NAND2X0 U12974 ( .IN1(n3819), .IN2(n12563), .QN(n12613) );
  NAND2X0 U12975 ( .IN1(n9496), .IN2(g6239), .QN(n12612) );
  NAND3X0 U12976 ( .IN1(n12614), .IN2(g6267), .IN3(n9333), .QN(n12611) );
  NAND2X0 U12977 ( .IN1(n11941), .IN2(n12563), .QN(n12614) );
  NOR2X0 U12978 ( .IN1(g6227), .IN2(n5385), .QN(n12563) );
  NAND3X0 U12979 ( .IN1(n12615), .IN2(n12616), .IN3(n12617), .QN(g30527) );
  NAND2X0 U12980 ( .IN1(n3819), .IN2(n12569), .QN(n12617) );
  NAND2X0 U12981 ( .IN1(n9496), .IN2(g6235), .QN(n12616) );
  NAND3X0 U12982 ( .IN1(n12618), .IN2(g6263), .IN3(n9333), .QN(n12615) );
  NAND2X0 U12983 ( .IN1(n11941), .IN2(n12569), .QN(n12618) );
  NOR2X0 U12984 ( .IN1(g6227), .IN2(g6219), .QN(n12569) );
  NOR2X0 U12985 ( .IN1(g6209), .IN2(n5574), .QN(n11941) );
  NAND3X0 U12986 ( .IN1(n12619), .IN2(n12620), .IN3(n12621), .QN(g30526) );
  NAND2X0 U12987 ( .IN1(n9496), .IN2(g6259), .QN(n12621) );
  NAND3X0 U12988 ( .IN1(n9347), .IN2(g6255), .IN3(n12622), .QN(n12620) );
  INVX0 U12989 ( .INP(n3824), .ZN(n12622) );
  NAND2X0 U12990 ( .IN1(n3824), .IN2(n3765), .QN(n12619) );
  NAND3X0 U12991 ( .IN1(n12623), .IN2(n12624), .IN3(n12625), .QN(g30525) );
  NAND2X0 U12992 ( .IN1(n9496), .IN2(g6251), .QN(n12625) );
  NAND3X0 U12993 ( .IN1(n9347), .IN2(g6247), .IN3(n12626), .QN(n12624) );
  INVX0 U12994 ( .INP(n3827), .ZN(n12626) );
  NAND2X0 U12995 ( .IN1(n3827), .IN2(n3765), .QN(n12623) );
  NAND3X0 U12996 ( .IN1(n12627), .IN2(n12628), .IN3(n12629), .QN(g30524) );
  NAND2X0 U12997 ( .IN1(n9496), .IN2(g6243), .QN(n12629) );
  NAND3X0 U12998 ( .IN1(n9349), .IN2(g6239), .IN3(n12630), .QN(n12628) );
  INVX0 U12999 ( .INP(n3829), .ZN(n12630) );
  NAND2X0 U13000 ( .IN1(n3829), .IN2(n3765), .QN(n12627) );
  NAND3X0 U13001 ( .IN1(n12631), .IN2(n12632), .IN3(n12633), .QN(g30523) );
  NAND2X0 U13002 ( .IN1(n9496), .IN2(g6227), .QN(n12633) );
  NAND3X0 U13003 ( .IN1(n9347), .IN2(g6235), .IN3(n12634), .QN(n12632) );
  INVX0 U13004 ( .INP(n3831), .ZN(n12634) );
  NAND2X0 U13005 ( .IN1(n3831), .IN2(n3765), .QN(n12631) );
  NOR2X0 U13006 ( .IN1(g6203), .IN2(n11934), .QN(g30522) );
  NAND3X0 U13007 ( .IN1(n11924), .IN2(n9315), .IN3(n5651), .QN(n11934) );
  NAND3X0 U13008 ( .IN1(g4093), .IN2(g4087), .IN3(n3833), .QN(n11924) );
  NAND3X0 U13009 ( .IN1(n12635), .IN2(n12636), .IN3(n12637), .QN(g30521) );
  NAND2X0 U13010 ( .IN1(n9496), .IN2(g5961), .QN(n12637) );
  NAND2X0 U13011 ( .IN1(test_so13), .IN2(n12638), .QN(n12636) );
  NAND2X0 U13012 ( .IN1(n12639), .IN2(n3765), .QN(n12635) );
  NAND3X0 U13013 ( .IN1(n12640), .IN2(n12641), .IN3(n12642), .QN(g30520) );
  NAND2X0 U13014 ( .IN1(n12643), .IN2(n3765), .QN(n12642) );
  NAND3X0 U13015 ( .IN1(n12644), .IN2(g5913), .IN3(n9333), .QN(n12641) );
  INVX0 U13016 ( .INP(n12643), .ZN(n12644) );
  NOR2X0 U13017 ( .IN1(n729), .IN2(n5649), .QN(n12643) );
  INVX0 U13018 ( .INP(n11949), .ZN(n729) );
  NAND2X0 U13019 ( .IN1(n9495), .IN2(g5957), .QN(n12640) );
  NAND3X0 U13020 ( .IN1(n12645), .IN2(n12646), .IN3(n12647), .QN(g30519) );
  NAND2X0 U13021 ( .IN1(n12648), .IN2(n3765), .QN(n12647) );
  NAND3X0 U13022 ( .IN1(n11947), .IN2(g5905), .IN3(n9333), .QN(n12646) );
  INVX0 U13023 ( .INP(n12648), .ZN(n11947) );
  NOR2X0 U13024 ( .IN1(n725), .IN2(n5649), .QN(n12648) );
  INVX0 U13025 ( .INP(n12649), .ZN(n725) );
  NAND2X0 U13026 ( .IN1(n9495), .IN2(g5953), .QN(n12645) );
  NAND3X0 U13027 ( .IN1(n12650), .IN2(n12651), .IN3(n12652), .QN(g30518) );
  NAND2X0 U13028 ( .IN1(n12653), .IN2(n3765), .QN(n12652) );
  NAND3X0 U13029 ( .IN1(n12654), .IN2(g5897), .IN3(n9333), .QN(n12651) );
  INVX0 U13030 ( .INP(n12653), .ZN(n12654) );
  NOR2X0 U13031 ( .IN1(n727), .IN2(n5649), .QN(n12653) );
  INVX0 U13032 ( .INP(n12655), .ZN(n727) );
  NAND2X0 U13033 ( .IN1(n9495), .IN2(g5949), .QN(n12650) );
  NAND3X0 U13034 ( .IN1(n12656), .IN2(n12657), .IN3(n12658), .QN(g30517) );
  NAND2X0 U13035 ( .IN1(n3842), .IN2(n12659), .QN(n12658) );
  NAND2X0 U13036 ( .IN1(n9495), .IN2(g5945), .QN(n12657) );
  NAND3X0 U13037 ( .IN1(n12660), .IN2(g5961), .IN3(n9333), .QN(n12656) );
  NAND2X0 U13038 ( .IN1(n9813), .IN2(n12659), .QN(n12660) );
  NAND3X0 U13039 ( .IN1(n12661), .IN2(n12662), .IN3(n12663), .QN(g30516) );
  NAND2X0 U13040 ( .IN1(n3842), .IN2(n11949), .QN(n12663) );
  NAND2X0 U13041 ( .IN1(n9495), .IN2(g5941), .QN(n12662) );
  NAND3X0 U13042 ( .IN1(n12664), .IN2(g5957), .IN3(n9333), .QN(n12661) );
  NAND2X0 U13043 ( .IN1(n9813), .IN2(n11949), .QN(n12664) );
  NAND3X0 U13044 ( .IN1(n12665), .IN2(n12666), .IN3(n12667), .QN(g30515) );
  NAND2X0 U13045 ( .IN1(n3842), .IN2(n12649), .QN(n12667) );
  NAND2X0 U13046 ( .IN1(n9495), .IN2(g5937), .QN(n12666) );
  NAND3X0 U13047 ( .IN1(n12668), .IN2(g5953), .IN3(n9333), .QN(n12665) );
  NAND2X0 U13048 ( .IN1(n9813), .IN2(n12649), .QN(n12668) );
  NAND3X0 U13049 ( .IN1(n12669), .IN2(n12670), .IN3(n12671), .QN(g30514) );
  NAND2X0 U13050 ( .IN1(n3842), .IN2(n12655), .QN(n12671) );
  NAND2X0 U13051 ( .IN1(n9495), .IN2(g5933), .QN(n12670) );
  NAND3X0 U13052 ( .IN1(n12672), .IN2(g5949), .IN3(n9333), .QN(n12669) );
  NAND2X0 U13053 ( .IN1(n9813), .IN2(n12655), .QN(n12672) );
  NOR2X0 U13054 ( .IN1(n5573), .IN2(n8770), .QN(n9813) );
  NAND3X0 U13055 ( .IN1(n12673), .IN2(n12674), .IN3(n12675), .QN(g30513) );
  NAND2X0 U13056 ( .IN1(n3848), .IN2(n12659), .QN(n12675) );
  NAND2X0 U13057 ( .IN1(n9494), .IN2(g5929), .QN(n12674) );
  NAND3X0 U13058 ( .IN1(n12676), .IN2(g5945), .IN3(n9333), .QN(n12673) );
  NAND2X0 U13059 ( .IN1(n9812), .IN2(n12659), .QN(n12676) );
  NAND3X0 U13060 ( .IN1(n12677), .IN2(n12678), .IN3(n12679), .QN(g30512) );
  NAND2X0 U13061 ( .IN1(n3848), .IN2(n11949), .QN(n12679) );
  NAND2X0 U13062 ( .IN1(n9494), .IN2(g5925), .QN(n12678) );
  NAND3X0 U13063 ( .IN1(n12680), .IN2(g5941), .IN3(n9333), .QN(n12677) );
  NAND2X0 U13064 ( .IN1(n9812), .IN2(n11949), .QN(n12680) );
  NAND3X0 U13065 ( .IN1(n12681), .IN2(n12682), .IN3(n12683), .QN(g30511) );
  NAND2X0 U13066 ( .IN1(n3848), .IN2(n12649), .QN(n12683) );
  NAND2X0 U13067 ( .IN1(n9494), .IN2(g5921), .QN(n12682) );
  NAND3X0 U13068 ( .IN1(n12684), .IN2(g5937), .IN3(n9333), .QN(n12681) );
  NAND2X0 U13069 ( .IN1(n9812), .IN2(n12649), .QN(n12684) );
  NAND3X0 U13070 ( .IN1(n12685), .IN2(n12686), .IN3(n12687), .QN(g30510) );
  NAND2X0 U13071 ( .IN1(n3848), .IN2(n12655), .QN(n12687) );
  NAND2X0 U13072 ( .IN1(test_so28), .IN2(n9416), .QN(n12686) );
  NAND3X0 U13073 ( .IN1(n12688), .IN2(g5933), .IN3(n9334), .QN(n12685) );
  NAND2X0 U13074 ( .IN1(n9812), .IN2(n12655), .QN(n12688) );
  NOR2X0 U13075 ( .IN1(g5857), .IN2(n8770), .QN(n9812) );
  NAND3X0 U13076 ( .IN1(n12689), .IN2(n12690), .IN3(n12691), .QN(g30509) );
  NAND2X0 U13077 ( .IN1(n3853), .IN2(n12659), .QN(n12691) );
  NAND2X0 U13078 ( .IN1(g5909), .IN2(n9429), .QN(n12690) );
  NAND3X0 U13079 ( .IN1(n12692), .IN2(g5929), .IN3(n9334), .QN(n12689) );
  NAND2X0 U13080 ( .IN1(n11962), .IN2(n12659), .QN(n12692) );
  NAND3X0 U13081 ( .IN1(n12693), .IN2(n12694), .IN3(n12695), .QN(g30508) );
  NAND2X0 U13082 ( .IN1(n3853), .IN2(n11949), .QN(n12695) );
  NAND2X0 U13083 ( .IN1(n9494), .IN2(g5901), .QN(n12694) );
  NAND3X0 U13084 ( .IN1(n12696), .IN2(g5925), .IN3(n9334), .QN(n12693) );
  NAND2X0 U13085 ( .IN1(n11962), .IN2(n11949), .QN(n12696) );
  NOR2X0 U13086 ( .IN1(g5873), .IN2(n8872), .QN(n11949) );
  NAND3X0 U13087 ( .IN1(n12697), .IN2(n12698), .IN3(n12699), .QN(g30507) );
  NAND2X0 U13088 ( .IN1(n3853), .IN2(n12649), .QN(n12699) );
  NAND2X0 U13089 ( .IN1(n9494), .IN2(g5893), .QN(n12698) );
  NAND3X0 U13090 ( .IN1(n12700), .IN2(g5921), .IN3(n9334), .QN(n12697) );
  NAND2X0 U13091 ( .IN1(n11962), .IN2(n12649), .QN(n12700) );
  NOR2X0 U13092 ( .IN1(n5388), .IN2(test_so36), .QN(n12649) );
  NAND3X0 U13093 ( .IN1(n12701), .IN2(n12702), .IN3(n12703), .QN(g30506) );
  NAND2X0 U13094 ( .IN1(n3853), .IN2(n12655), .QN(n12703) );
  NAND2X0 U13095 ( .IN1(n9494), .IN2(g5889), .QN(n12702) );
  NAND3X0 U13096 ( .IN1(test_so28), .IN2(n12704), .IN3(n9334), .QN(n12701) );
  NAND2X0 U13097 ( .IN1(n11962), .IN2(n12655), .QN(n12704) );
  NOR2X0 U13098 ( .IN1(g5873), .IN2(test_so36), .QN(n12655) );
  NOR2X0 U13099 ( .IN1(g5863), .IN2(n5573), .QN(n11962) );
  NAND3X0 U13100 ( .IN1(n12705), .IN2(n12706), .IN3(n12707), .QN(g30505) );
  NAND2X0 U13101 ( .IN1(n9494), .IN2(g5913), .QN(n12707) );
  NAND3X0 U13102 ( .IN1(g5909), .IN2(n9313), .IN3(n12708), .QN(n12706) );
  INVX0 U13103 ( .INP(n3858), .ZN(n12708) );
  NAND2X0 U13104 ( .IN1(n3858), .IN2(n3765), .QN(n12705) );
  NAND3X0 U13105 ( .IN1(n12709), .IN2(n12710), .IN3(n12711), .QN(g30504) );
  NAND2X0 U13106 ( .IN1(n9493), .IN2(g5905), .QN(n12711) );
  NAND3X0 U13107 ( .IN1(n9347), .IN2(g5901), .IN3(n12712), .QN(n12710) );
  INVX0 U13108 ( .INP(n3861), .ZN(n12712) );
  NAND2X0 U13109 ( .IN1(n3861), .IN2(n3765), .QN(n12709) );
  NAND3X0 U13110 ( .IN1(n12713), .IN2(n12714), .IN3(n12715), .QN(g30503) );
  NAND2X0 U13111 ( .IN1(n9493), .IN2(g5897), .QN(n12715) );
  NAND3X0 U13112 ( .IN1(n9347), .IN2(g5893), .IN3(n12716), .QN(n12714) );
  INVX0 U13113 ( .INP(n3863), .ZN(n12716) );
  NAND2X0 U13114 ( .IN1(n3863), .IN2(n3765), .QN(n12713) );
  NAND3X0 U13115 ( .IN1(n12717), .IN2(n12718), .IN3(n12719), .QN(g30502) );
  NAND2X0 U13116 ( .IN1(test_so36), .IN2(n9512), .QN(n12719) );
  NAND3X0 U13117 ( .IN1(n9347), .IN2(g5889), .IN3(n12720), .QN(n12718) );
  INVX0 U13118 ( .INP(n3865), .ZN(n12720) );
  NAND2X0 U13119 ( .IN1(n3865), .IN2(n3765), .QN(n12717) );
  NOR2X0 U13120 ( .IN1(g5857), .IN2(n11955), .QN(g30501) );
  NAND3X0 U13121 ( .IN1(n11945), .IN2(n9313), .IN3(n5649), .QN(n11955) );
  NAND3X0 U13122 ( .IN1(n5480), .IN2(g4093), .IN3(n3833), .QN(n11945) );
  NAND3X0 U13123 ( .IN1(n12721), .IN2(n12722), .IN3(n12723), .QN(g30500) );
  NAND2X0 U13124 ( .IN1(n9493), .IN2(g5615), .QN(n12723) );
  NAND2X0 U13125 ( .IN1(n12724), .IN2(g5619), .QN(n12722) );
  NAND2X0 U13126 ( .IN1(n3765), .IN2(n11354), .QN(n12721) );
  NAND3X0 U13127 ( .IN1(n12725), .IN2(n12726), .IN3(n12727), .QN(g30499) );
  NAND2X0 U13128 ( .IN1(n12728), .IN2(n3765), .QN(n12727) );
  NAND3X0 U13129 ( .IN1(n12729), .IN2(g5567), .IN3(n9317), .QN(n12726) );
  INVX0 U13130 ( .INP(n12728), .ZN(n12729) );
  NOR2X0 U13131 ( .IN1(n955), .IN2(n5647), .QN(n12728) );
  INVX0 U13132 ( .INP(n11970), .ZN(n955) );
  NAND2X0 U13133 ( .IN1(n9493), .IN2(g5611), .QN(n12725) );
  NAND3X0 U13134 ( .IN1(n12730), .IN2(n12731), .IN3(n12732), .QN(g30498) );
  NAND2X0 U13135 ( .IN1(n12733), .IN2(n3765), .QN(n12732) );
  NAND3X0 U13136 ( .IN1(test_so6), .IN2(n11968), .IN3(n9343), .QN(n12731) );
  INVX0 U13137 ( .INP(n12733), .ZN(n11968) );
  NOR2X0 U13138 ( .IN1(n957), .IN2(n5647), .QN(n12733) );
  INVX0 U13139 ( .INP(n12734), .ZN(n957) );
  NAND2X0 U13140 ( .IN1(n9493), .IN2(g5607), .QN(n12730) );
  NAND3X0 U13141 ( .IN1(n12735), .IN2(n12736), .IN3(n12737), .QN(g30497) );
  NAND2X0 U13142 ( .IN1(n12738), .IN2(n3765), .QN(n12737) );
  NAND3X0 U13143 ( .IN1(n12739), .IN2(g5551), .IN3(n9329), .QN(n12736) );
  INVX0 U13144 ( .INP(n12738), .ZN(n12739) );
  NOR2X0 U13145 ( .IN1(n956), .IN2(n5647), .QN(n12738) );
  INVX0 U13146 ( .INP(n12740), .ZN(n956) );
  NAND2X0 U13147 ( .IN1(n9493), .IN2(g5603), .QN(n12735) );
  NAND3X0 U13148 ( .IN1(n12741), .IN2(n12742), .IN3(n12743), .QN(g30496) );
  NAND2X0 U13149 ( .IN1(n3875), .IN2(n9657), .QN(n12743) );
  NAND2X0 U13150 ( .IN1(n9493), .IN2(g5599), .QN(n12742) );
  NAND3X0 U13151 ( .IN1(n12744), .IN2(g5615), .IN3(n9329), .QN(n12741) );
  NAND2X0 U13152 ( .IN1(n9688), .IN2(n9657), .QN(n12744) );
  NAND3X0 U13153 ( .IN1(n12745), .IN2(n12746), .IN3(n12747), .QN(g30495) );
  NAND2X0 U13154 ( .IN1(n3875), .IN2(n11970), .QN(n12747) );
  NAND2X0 U13155 ( .IN1(n9492), .IN2(g5595), .QN(n12746) );
  NAND3X0 U13156 ( .IN1(n12748), .IN2(g5611), .IN3(n9329), .QN(n12745) );
  NAND2X0 U13157 ( .IN1(n9688), .IN2(n11970), .QN(n12748) );
  NAND3X0 U13158 ( .IN1(n12749), .IN2(n12750), .IN3(n12751), .QN(g30494) );
  NAND2X0 U13159 ( .IN1(n3875), .IN2(n12734), .QN(n12751) );
  NAND2X0 U13160 ( .IN1(test_so5), .IN2(n9511), .QN(n12750) );
  NAND3X0 U13161 ( .IN1(n12752), .IN2(g5607), .IN3(n9329), .QN(n12749) );
  NAND2X0 U13162 ( .IN1(n9688), .IN2(n12734), .QN(n12752) );
  NAND3X0 U13163 ( .IN1(n12753), .IN2(n12754), .IN3(n12755), .QN(g30493) );
  NAND2X0 U13164 ( .IN1(n3875), .IN2(n12740), .QN(n12755) );
  NAND2X0 U13165 ( .IN1(n9492), .IN2(g5587), .QN(n12754) );
  NAND3X0 U13166 ( .IN1(n12756), .IN2(g5603), .IN3(n9328), .QN(n12753) );
  NAND2X0 U13167 ( .IN1(n9688), .IN2(n12740), .QN(n12756) );
  NOR2X0 U13168 ( .IN1(n5575), .IN2(n8769), .QN(n9688) );
  NAND3X0 U13169 ( .IN1(n12757), .IN2(n12758), .IN3(n12759), .QN(g30492) );
  NAND2X0 U13170 ( .IN1(n3881), .IN2(n9657), .QN(n12759) );
  NAND2X0 U13171 ( .IN1(n9492), .IN2(g5583), .QN(n12758) );
  NAND3X0 U13172 ( .IN1(n12760), .IN2(g5599), .IN3(n9328), .QN(n12757) );
  NAND2X0 U13173 ( .IN1(n9687), .IN2(n9657), .QN(n12760) );
  NAND3X0 U13174 ( .IN1(n12761), .IN2(n12762), .IN3(n12763), .QN(g30491) );
  NAND2X0 U13175 ( .IN1(n3881), .IN2(n11970), .QN(n12763) );
  NAND2X0 U13176 ( .IN1(n9492), .IN2(g5579), .QN(n12762) );
  NAND3X0 U13177 ( .IN1(n12764), .IN2(g5595), .IN3(n9328), .QN(n12761) );
  NAND2X0 U13178 ( .IN1(n9687), .IN2(n11970), .QN(n12764) );
  NAND3X0 U13179 ( .IN1(n12765), .IN2(n12766), .IN3(n12767), .QN(g30490) );
  NAND2X0 U13180 ( .IN1(n3881), .IN2(n12734), .QN(n12767) );
  NAND2X0 U13181 ( .IN1(n9492), .IN2(g5575), .QN(n12766) );
  NAND3X0 U13182 ( .IN1(test_so5), .IN2(n12768), .IN3(n9328), .QN(n12765) );
  NAND2X0 U13183 ( .IN1(n9687), .IN2(n12734), .QN(n12768) );
  NAND3X0 U13184 ( .IN1(n12769), .IN2(n12770), .IN3(n12771), .QN(g30489) );
  NAND2X0 U13185 ( .IN1(n3881), .IN2(n12740), .QN(n12771) );
  NAND2X0 U13186 ( .IN1(n9492), .IN2(g5571), .QN(n12770) );
  NAND3X0 U13187 ( .IN1(n12772), .IN2(g5587), .IN3(n9328), .QN(n12769) );
  NAND2X0 U13188 ( .IN1(n9687), .IN2(n12740), .QN(n12772) );
  NOR2X0 U13189 ( .IN1(g5511), .IN2(n8769), .QN(n9687) );
  NAND3X0 U13190 ( .IN1(n12773), .IN2(n12774), .IN3(n12775), .QN(g30488) );
  NAND2X0 U13191 ( .IN1(n3886), .IN2(n9657), .QN(n12775) );
  NAND2X0 U13192 ( .IN1(n9492), .IN2(g5563), .QN(n12774) );
  NAND3X0 U13193 ( .IN1(n12776), .IN2(g5583), .IN3(n9328), .QN(n12773) );
  NAND2X0 U13194 ( .IN1(n11983), .IN2(n9657), .QN(n12776) );
  NAND3X0 U13195 ( .IN1(n12777), .IN2(n12778), .IN3(n12779), .QN(g30487) );
  NAND2X0 U13196 ( .IN1(n3886), .IN2(n11970), .QN(n12779) );
  NAND2X0 U13197 ( .IN1(n9491), .IN2(g5555), .QN(n12778) );
  NAND3X0 U13198 ( .IN1(n12780), .IN2(g5579), .IN3(n9328), .QN(n12777) );
  NAND2X0 U13199 ( .IN1(n11983), .IN2(n11970), .QN(n12780) );
  NOR2X0 U13200 ( .IN1(g5527), .IN2(n5566), .QN(n11970) );
  NAND3X0 U13201 ( .IN1(n12781), .IN2(n12782), .IN3(n12783), .QN(g30486) );
  NAND2X0 U13202 ( .IN1(n3886), .IN2(n12734), .QN(n12783) );
  NAND2X0 U13203 ( .IN1(n9491), .IN2(g5547), .QN(n12782) );
  NAND3X0 U13204 ( .IN1(n12784), .IN2(g5575), .IN3(n9328), .QN(n12781) );
  NAND2X0 U13205 ( .IN1(n11983), .IN2(n12734), .QN(n12784) );
  NOR2X0 U13206 ( .IN1(g5535), .IN2(n5389), .QN(n12734) );
  NAND3X0 U13207 ( .IN1(n12785), .IN2(n12786), .IN3(n12787), .QN(g30485) );
  NAND2X0 U13208 ( .IN1(n3886), .IN2(n12740), .QN(n12787) );
  NAND2X0 U13209 ( .IN1(n9491), .IN2(g5543), .QN(n12786) );
  NAND3X0 U13210 ( .IN1(n12788), .IN2(g5571), .IN3(n9328), .QN(n12785) );
  NAND2X0 U13211 ( .IN1(n11983), .IN2(n12740), .QN(n12788) );
  NOR2X0 U13212 ( .IN1(g5527), .IN2(g5535), .QN(n12740) );
  NOR2X0 U13213 ( .IN1(g5517), .IN2(n5575), .QN(n11983) );
  NAND3X0 U13214 ( .IN1(n12789), .IN2(n12790), .IN3(n12791), .QN(g30484) );
  NAND2X0 U13215 ( .IN1(n9491), .IN2(g5567), .QN(n12791) );
  NAND3X0 U13216 ( .IN1(n9350), .IN2(g5563), .IN3(n12792), .QN(n12790) );
  INVX0 U13217 ( .INP(n3891), .ZN(n12792) );
  NAND2X0 U13218 ( .IN1(n3891), .IN2(n3765), .QN(n12789) );
  NAND3X0 U13219 ( .IN1(n12793), .IN2(n12794), .IN3(n12795), .QN(g30483) );
  NAND2X0 U13220 ( .IN1(test_so6), .IN2(n9514), .QN(n12795) );
  NAND3X0 U13221 ( .IN1(n9350), .IN2(g5555), .IN3(n12796), .QN(n12794) );
  INVX0 U13222 ( .INP(n3894), .ZN(n12796) );
  NAND2X0 U13223 ( .IN1(n3894), .IN2(n3765), .QN(n12793) );
  NAND3X0 U13224 ( .IN1(n12797), .IN2(n12798), .IN3(n12799), .QN(g30482) );
  NAND2X0 U13225 ( .IN1(n9491), .IN2(g5551), .QN(n12799) );
  NAND3X0 U13226 ( .IN1(n9350), .IN2(g5547), .IN3(n12800), .QN(n12798) );
  INVX0 U13227 ( .INP(n3896), .ZN(n12800) );
  NAND2X0 U13228 ( .IN1(n3896), .IN2(n3765), .QN(n12797) );
  NAND3X0 U13229 ( .IN1(n12801), .IN2(n12802), .IN3(n12803), .QN(g30481) );
  NAND2X0 U13230 ( .IN1(n9491), .IN2(g5535), .QN(n12803) );
  NAND3X0 U13231 ( .IN1(n9350), .IN2(g5543), .IN3(n12804), .QN(n12802) );
  INVX0 U13232 ( .INP(n3898), .ZN(n12804) );
  NAND2X0 U13233 ( .IN1(n3898), .IN2(n3765), .QN(n12801) );
  NOR2X0 U13234 ( .IN1(g5511), .IN2(n11976), .QN(g30480) );
  NAND3X0 U13235 ( .IN1(n11966), .IN2(n9315), .IN3(n5647), .QN(n11976) );
  NAND2X0 U13236 ( .IN1(n3833), .IN2(n11355), .QN(n11966) );
  NAND3X0 U13237 ( .IN1(n12805), .IN2(n12806), .IN3(n12807), .QN(g30479) );
  NAND2X0 U13238 ( .IN1(n9491), .IN2(g5268), .QN(n12807) );
  NAND2X0 U13239 ( .IN1(n12808), .IN2(g5272), .QN(n12806) );
  NAND2X0 U13240 ( .IN1(n3765), .IN2(g32975), .QN(n12805) );
  NAND3X0 U13241 ( .IN1(n12809), .IN2(n12810), .IN3(n12811), .QN(g30478) );
  NAND2X0 U13242 ( .IN1(n12812), .IN2(n3765), .QN(n12811) );
  NAND3X0 U13243 ( .IN1(n12813), .IN2(g5220), .IN3(n9328), .QN(n12810) );
  INVX0 U13244 ( .INP(n12812), .ZN(n12813) );
  NOR2X0 U13245 ( .IN1(n194), .IN2(n5650), .QN(n12812) );
  INVX0 U13246 ( .INP(n11991), .ZN(n194) );
  NAND2X0 U13247 ( .IN1(n9490), .IN2(g5264), .QN(n12809) );
  NAND3X0 U13248 ( .IN1(n12814), .IN2(n12815), .IN3(n12816), .QN(g30477) );
  NAND2X0 U13249 ( .IN1(n12817), .IN2(n3765), .QN(n12816) );
  NAND3X0 U13250 ( .IN1(n11989), .IN2(g5212), .IN3(n9326), .QN(n12815) );
  INVX0 U13251 ( .INP(n12817), .ZN(n11989) );
  NOR2X0 U13252 ( .IN1(n190), .IN2(n5650), .QN(n12817) );
  INVX0 U13253 ( .INP(n12818), .ZN(n190) );
  NAND2X0 U13254 ( .IN1(n9490), .IN2(g5260), .QN(n12814) );
  NAND3X0 U13255 ( .IN1(n12819), .IN2(n12820), .IN3(n12821), .QN(g30476) );
  NAND2X0 U13256 ( .IN1(n12822), .IN2(n3765), .QN(n12821) );
  NAND3X0 U13257 ( .IN1(n12823), .IN2(g5204), .IN3(n9326), .QN(n12820) );
  INVX0 U13258 ( .INP(n12822), .ZN(n12823) );
  NOR2X0 U13259 ( .IN1(n192), .IN2(n5650), .QN(n12822) );
  INVX0 U13260 ( .INP(n12824), .ZN(n192) );
  NAND2X0 U13261 ( .IN1(n9490), .IN2(g5256), .QN(n12819) );
  NAND3X0 U13262 ( .IN1(n12825), .IN2(n12826), .IN3(n12827), .QN(g30475) );
  NAND2X0 U13263 ( .IN1(n3908), .IN2(n9800), .QN(n12827) );
  NAND2X0 U13264 ( .IN1(n9490), .IN2(g5252), .QN(n12826) );
  NAND3X0 U13265 ( .IN1(n12828), .IN2(g5268), .IN3(n9326), .QN(n12825) );
  NAND2X0 U13266 ( .IN1(n9800), .IN2(n9668), .QN(n12828) );
  NAND3X0 U13267 ( .IN1(n12829), .IN2(n12830), .IN3(n12831), .QN(g30474) );
  NAND2X0 U13268 ( .IN1(n3908), .IN2(n11991), .QN(n12831) );
  NAND2X0 U13269 ( .IN1(n9490), .IN2(g5248), .QN(n12830) );
  NAND3X0 U13270 ( .IN1(n12832), .IN2(g5264), .IN3(n9326), .QN(n12829) );
  NAND2X0 U13271 ( .IN1(n11991), .IN2(n9668), .QN(n12832) );
  NAND3X0 U13272 ( .IN1(n12833), .IN2(n12834), .IN3(n12835), .QN(g30473) );
  NAND2X0 U13273 ( .IN1(n3908), .IN2(n12818), .QN(n12835) );
  NAND2X0 U13274 ( .IN1(n9490), .IN2(g5244), .QN(n12834) );
  NAND3X0 U13275 ( .IN1(n12836), .IN2(g5260), .IN3(n9326), .QN(n12833) );
  NAND2X0 U13276 ( .IN1(n12818), .IN2(n9668), .QN(n12836) );
  NAND3X0 U13277 ( .IN1(n12837), .IN2(n12838), .IN3(n12839), .QN(g30472) );
  NAND2X0 U13278 ( .IN1(n3908), .IN2(n12824), .QN(n12839) );
  NAND2X0 U13279 ( .IN1(n9490), .IN2(g5240), .QN(n12838) );
  NAND3X0 U13280 ( .IN1(n12840), .IN2(g5256), .IN3(n9326), .QN(n12837) );
  NAND2X0 U13281 ( .IN1(n12824), .IN2(n9668), .QN(n12840) );
  NOR2X0 U13282 ( .IN1(n5570), .IN2(n8766), .QN(n9668) );
  NAND3X0 U13283 ( .IN1(n12841), .IN2(n12842), .IN3(n12843), .QN(g30471) );
  NAND2X0 U13284 ( .IN1(n3914), .IN2(n9800), .QN(n12843) );
  NAND2X0 U13285 ( .IN1(n9489), .IN2(g5236), .QN(n12842) );
  NAND3X0 U13286 ( .IN1(n12844), .IN2(g5252), .IN3(n9326), .QN(n12841) );
  NAND2X0 U13287 ( .IN1(n9800), .IN2(n9667), .QN(n12844) );
  NAND3X0 U13288 ( .IN1(n12845), .IN2(n12846), .IN3(n12847), .QN(g30470) );
  NAND2X0 U13289 ( .IN1(n3914), .IN2(n11991), .QN(n12847) );
  NAND2X0 U13290 ( .IN1(g5232), .IN2(n9515), .QN(n12846) );
  NAND3X0 U13291 ( .IN1(n12848), .IN2(g5248), .IN3(n9326), .QN(n12845) );
  NAND2X0 U13292 ( .IN1(n11991), .IN2(n9667), .QN(n12848) );
  NAND3X0 U13293 ( .IN1(n12849), .IN2(n12850), .IN3(n12851), .QN(g30469) );
  NAND2X0 U13294 ( .IN1(n3914), .IN2(n12818), .QN(n12851) );
  NAND2X0 U13295 ( .IN1(test_so82), .IN2(n9516), .QN(n12850) );
  NAND3X0 U13296 ( .IN1(n12852), .IN2(g5244), .IN3(n9326), .QN(n12849) );
  NAND2X0 U13297 ( .IN1(n12818), .IN2(n9667), .QN(n12852) );
  NAND3X0 U13298 ( .IN1(n12853), .IN2(n12854), .IN3(n12855), .QN(g30468) );
  NAND2X0 U13299 ( .IN1(n3914), .IN2(n12824), .QN(n12855) );
  NAND2X0 U13300 ( .IN1(n9489), .IN2(g5224), .QN(n12854) );
  NAND3X0 U13301 ( .IN1(n12856), .IN2(g5240), .IN3(n9326), .QN(n12853) );
  NAND2X0 U13302 ( .IN1(n12824), .IN2(n9667), .QN(n12856) );
  NOR2X0 U13303 ( .IN1(g5164), .IN2(n8766), .QN(n9667) );
  NAND3X0 U13304 ( .IN1(n12857), .IN2(n12858), .IN3(n12859), .QN(g30467) );
  NAND2X0 U13305 ( .IN1(n3919), .IN2(n9800), .QN(n12859) );
  NAND2X0 U13306 ( .IN1(n9489), .IN2(g5216), .QN(n12858) );
  NAND3X0 U13307 ( .IN1(n12860), .IN2(g5236), .IN3(n9323), .QN(n12857) );
  NAND2X0 U13308 ( .IN1(n9800), .IN2(n12004), .QN(n12860) );
  NAND3X0 U13309 ( .IN1(n12861), .IN2(n12862), .IN3(n12863), .QN(g30466) );
  NAND2X0 U13310 ( .IN1(n3919), .IN2(n11991), .QN(n12863) );
  NAND2X0 U13311 ( .IN1(n9489), .IN2(g5208), .QN(n12862) );
  NAND3X0 U13312 ( .IN1(g5232), .IN2(n12864), .IN3(n9323), .QN(n12861) );
  NAND2X0 U13313 ( .IN1(n11991), .IN2(n12004), .QN(n12864) );
  NOR2X0 U13314 ( .IN1(g5180), .IN2(n5567), .QN(n11991) );
  NAND3X0 U13315 ( .IN1(n12865), .IN2(n12866), .IN3(n12867), .QN(g30465) );
  NAND2X0 U13316 ( .IN1(n3919), .IN2(n12818), .QN(n12867) );
  NAND2X0 U13317 ( .IN1(n9489), .IN2(g5200), .QN(n12866) );
  NAND3X0 U13318 ( .IN1(test_so82), .IN2(n12868), .IN3(n9323), .QN(n12865) );
  NAND2X0 U13319 ( .IN1(n12818), .IN2(n12004), .QN(n12868) );
  NOR2X0 U13320 ( .IN1(g5188), .IN2(n5384), .QN(n12818) );
  NAND3X0 U13321 ( .IN1(n12869), .IN2(n12870), .IN3(n12871), .QN(g30464) );
  NAND2X0 U13322 ( .IN1(n3919), .IN2(n12824), .QN(n12871) );
  NAND2X0 U13323 ( .IN1(n9489), .IN2(g5196), .QN(n12870) );
  NAND3X0 U13324 ( .IN1(n12872), .IN2(g5224), .IN3(n9318), .QN(n12869) );
  NAND2X0 U13325 ( .IN1(n12824), .IN2(n12004), .QN(n12872) );
  NOR2X0 U13326 ( .IN1(g5170), .IN2(n5570), .QN(n12004) );
  NOR2X0 U13327 ( .IN1(g5188), .IN2(g5180), .QN(n12824) );
  NAND3X0 U13328 ( .IN1(n12873), .IN2(n12874), .IN3(n12875), .QN(g30463) );
  NAND2X0 U13329 ( .IN1(n9489), .IN2(g5220), .QN(n12875) );
  NAND3X0 U13330 ( .IN1(n9353), .IN2(g5216), .IN3(n12876), .QN(n12874) );
  INVX0 U13331 ( .INP(n3924), .ZN(n12876) );
  NAND2X0 U13332 ( .IN1(n3924), .IN2(n3765), .QN(n12873) );
  NAND3X0 U13333 ( .IN1(n12877), .IN2(n12878), .IN3(n12879), .QN(g30462) );
  NAND2X0 U13334 ( .IN1(n9488), .IN2(g5212), .QN(n12879) );
  NAND3X0 U13335 ( .IN1(n9353), .IN2(g5208), .IN3(n12880), .QN(n12878) );
  INVX0 U13336 ( .INP(n3927), .ZN(n12880) );
  NAND2X0 U13337 ( .IN1(n3927), .IN2(n3765), .QN(n12877) );
  NAND3X0 U13338 ( .IN1(n12881), .IN2(n12882), .IN3(n12883), .QN(g30461) );
  NAND2X0 U13339 ( .IN1(n9488), .IN2(g5204), .QN(n12883) );
  NAND3X0 U13340 ( .IN1(n9353), .IN2(g5200), .IN3(n12884), .QN(n12882) );
  INVX0 U13341 ( .INP(n3929), .ZN(n12884) );
  NAND2X0 U13342 ( .IN1(n3929), .IN2(n3765), .QN(n12881) );
  NAND3X0 U13343 ( .IN1(n12885), .IN2(n12886), .IN3(n12887), .QN(g30460) );
  NAND2X0 U13344 ( .IN1(n9488), .IN2(g5188), .QN(n12887) );
  NAND3X0 U13345 ( .IN1(n9353), .IN2(g5196), .IN3(n12888), .QN(n12886) );
  INVX0 U13346 ( .INP(n3931), .ZN(n12888) );
  NAND2X0 U13347 ( .IN1(n3931), .IN2(n3765), .QN(n12885) );
  NOR2X0 U13348 ( .IN1(g5164), .IN2(n11997), .QN(g30459) );
  NAND3X0 U13349 ( .IN1(n11987), .IN2(n9315), .IN3(n5650), .QN(n11997) );
  NAND2X0 U13350 ( .IN1(n3833), .IN2(n11360), .QN(n11987) );
  NAND3X0 U13351 ( .IN1(n12889), .IN2(n12890), .IN3(n9318), .QN(g30458) );
  NAND2X0 U13352 ( .IN1(n12891), .IN2(g113), .QN(n12890) );
  INVX0 U13353 ( .INP(n12892), .ZN(n12889) );
  NOR2X0 U13354 ( .IN1(n12891), .IN2(n5846), .QN(n12892) );
  NOR2X0 U13355 ( .IN1(g4459), .IN2(n8423), .QN(n12891) );
  NAND2X0 U13356 ( .IN1(n12893), .IN2(n12894), .QN(g30457) );
  NAND2X0 U13357 ( .IN1(n9488), .IN2(g4122), .QN(n12894) );
  NAND2X0 U13358 ( .IN1(n12895), .IN2(n9374), .QN(n12893) );
  NAND2X0 U13359 ( .IN1(n12896), .IN2(n12897), .QN(n12895) );
  NAND3X0 U13360 ( .IN1(n12898), .IN2(n12899), .IN3(n5981), .QN(n12897) );
  NAND2X0 U13361 ( .IN1(g126), .IN2(n12900), .QN(n12899) );
  INVX0 U13362 ( .INP(n12901), .ZN(n12900) );
  NAND2X0 U13363 ( .IN1(n12901), .IN2(n12902), .QN(n12898) );
  INVX0 U13364 ( .INP(g126), .ZN(n12902) );
  NAND3X0 U13365 ( .IN1(n12903), .IN2(n12904), .IN3(n5983), .QN(n12896) );
  NAND2X0 U13366 ( .IN1(g115), .IN2(n12905), .QN(n12904) );
  INVX0 U13367 ( .INP(n12906), .ZN(n12905) );
  NAND2X0 U13368 ( .IN1(n12906), .IN2(n12907), .QN(n12903) );
  INVX0 U13369 ( .INP(g115), .ZN(n12907) );
  NAND3X0 U13370 ( .IN1(n12908), .IN2(n12909), .IN3(n12910), .QN(g30456) );
  NAND2X0 U13371 ( .IN1(n9488), .IN2(g4087), .QN(n12910) );
  NAND3X0 U13372 ( .IN1(n11355), .IN2(g4169), .IN3(n12911), .QN(n12909) );
  NAND2X0 U13373 ( .IN1(n3941), .IN2(n12912), .QN(n12908) );
  NAND3X0 U13374 ( .IN1(n12913), .IN2(n12914), .IN3(n12915), .QN(g30455) );
  NAND2X0 U13375 ( .IN1(n9488), .IN2(g3961), .QN(n12915) );
  NAND2X0 U13376 ( .IN1(n12916), .IN2(g3965), .QN(n12914) );
  NAND2X0 U13377 ( .IN1(n12917), .IN2(n3765), .QN(n12913) );
  NAND3X0 U13378 ( .IN1(n12918), .IN2(n12919), .IN3(n12920), .QN(g30454) );
  NAND2X0 U13379 ( .IN1(n12921), .IN2(n3765), .QN(n12920) );
  NAND3X0 U13380 ( .IN1(n12922), .IN2(g3913), .IN3(n9317), .QN(n12919) );
  INVX0 U13381 ( .INP(n12921), .ZN(n12922) );
  NOR2X0 U13382 ( .IN1(n8868), .IN2(n845), .QN(n12921) );
  INVX0 U13383 ( .INP(n12043), .ZN(n845) );
  NAND2X0 U13384 ( .IN1(n9501), .IN2(g3957), .QN(n12918) );
  NAND3X0 U13385 ( .IN1(n12923), .IN2(n12924), .IN3(n12925), .QN(g30453) );
  NAND2X0 U13386 ( .IN1(n12926), .IN2(n3765), .QN(n12925) );
  NAND3X0 U13387 ( .IN1(n12041), .IN2(g3905), .IN3(n9317), .QN(n12924) );
  INVX0 U13388 ( .INP(n12926), .ZN(n12041) );
  NOR2X0 U13389 ( .IN1(n8868), .IN2(n841), .QN(n12926) );
  INVX0 U13390 ( .INP(n12927), .ZN(n841) );
  NAND2X0 U13391 ( .IN1(n9468), .IN2(g3953), .QN(n12923) );
  NAND3X0 U13392 ( .IN1(n12928), .IN2(n12929), .IN3(n12930), .QN(g30452) );
  NAND2X0 U13393 ( .IN1(n12931), .IN2(n3765), .QN(n12930) );
  NAND3X0 U13394 ( .IN1(n12932), .IN2(g3897), .IN3(n9317), .QN(n12929) );
  INVX0 U13395 ( .INP(n12931), .ZN(n12932) );
  NOR2X0 U13396 ( .IN1(n8868), .IN2(n843), .QN(n12931) );
  INVX0 U13397 ( .INP(n12933), .ZN(n843) );
  NAND2X0 U13398 ( .IN1(test_so65), .IN2(n9516), .QN(n12928) );
  NAND3X0 U13399 ( .IN1(n12934), .IN2(n12935), .IN3(n12936), .QN(g30451) );
  NAND2X0 U13400 ( .IN1(n3951), .IN2(n12937), .QN(n12936) );
  NAND2X0 U13401 ( .IN1(n9432), .IN2(g3945), .QN(n12935) );
  NAND3X0 U13402 ( .IN1(n12938), .IN2(g3961), .IN3(n9317), .QN(n12934) );
  NAND2X0 U13403 ( .IN1(n9811), .IN2(n12937), .QN(n12938) );
  NAND3X0 U13404 ( .IN1(n12939), .IN2(n12940), .IN3(n12941), .QN(g30450) );
  NAND2X0 U13405 ( .IN1(n3951), .IN2(n12043), .QN(n12941) );
  NAND2X0 U13406 ( .IN1(n9432), .IN2(g3941), .QN(n12940) );
  NAND3X0 U13407 ( .IN1(n12942), .IN2(g3957), .IN3(n9317), .QN(n12939) );
  NAND2X0 U13408 ( .IN1(n9811), .IN2(n12043), .QN(n12942) );
  NAND3X0 U13409 ( .IN1(n12943), .IN2(n12944), .IN3(n12945), .QN(g30449) );
  NAND2X0 U13410 ( .IN1(n3951), .IN2(n12927), .QN(n12945) );
  NAND2X0 U13411 ( .IN1(n9432), .IN2(g3937), .QN(n12944) );
  NAND3X0 U13412 ( .IN1(n12946), .IN2(g3953), .IN3(n9317), .QN(n12943) );
  NAND2X0 U13413 ( .IN1(n9811), .IN2(n12927), .QN(n12946) );
  NAND3X0 U13414 ( .IN1(n12947), .IN2(n12948), .IN3(n12949), .QN(g30448) );
  NAND2X0 U13415 ( .IN1(n3951), .IN2(n12933), .QN(n12949) );
  NAND2X0 U13416 ( .IN1(n9432), .IN2(g3933), .QN(n12948) );
  NAND3X0 U13417 ( .IN1(test_so65), .IN2(n12950), .IN3(n9318), .QN(n12947) );
  NAND2X0 U13418 ( .IN1(n9811), .IN2(n12933), .QN(n12950) );
  NOR2X0 U13419 ( .IN1(n5572), .IN2(n8771), .QN(n9811) );
  NAND3X0 U13420 ( .IN1(n12951), .IN2(n12952), .IN3(n12953), .QN(g30447) );
  NAND2X0 U13421 ( .IN1(n3957), .IN2(n12937), .QN(n12953) );
  NAND2X0 U13422 ( .IN1(n9432), .IN2(g3929), .QN(n12952) );
  NAND3X0 U13423 ( .IN1(n12954), .IN2(g3945), .IN3(n9317), .QN(n12951) );
  NAND2X0 U13424 ( .IN1(n9810), .IN2(n12937), .QN(n12954) );
  NAND3X0 U13425 ( .IN1(n12955), .IN2(n12956), .IN3(n12957), .QN(g30446) );
  NAND2X0 U13426 ( .IN1(n3957), .IN2(n12043), .QN(n12957) );
  NAND2X0 U13427 ( .IN1(n9432), .IN2(g3925), .QN(n12956) );
  NAND3X0 U13428 ( .IN1(n12958), .IN2(g3941), .IN3(n9317), .QN(n12955) );
  NAND2X0 U13429 ( .IN1(n9810), .IN2(n12043), .QN(n12958) );
  NAND3X0 U13430 ( .IN1(n12959), .IN2(n12960), .IN3(n12961), .QN(g30445) );
  NAND2X0 U13431 ( .IN1(n3957), .IN2(n12927), .QN(n12961) );
  NAND2X0 U13432 ( .IN1(n9433), .IN2(g3921), .QN(n12960) );
  NAND3X0 U13433 ( .IN1(n12962), .IN2(g3937), .IN3(n9318), .QN(n12959) );
  NAND2X0 U13434 ( .IN1(n9810), .IN2(n12927), .QN(n12962) );
  NAND3X0 U13435 ( .IN1(n12963), .IN2(n12964), .IN3(n12965), .QN(g30444) );
  NAND2X0 U13436 ( .IN1(n3957), .IN2(n12933), .QN(n12965) );
  NAND2X0 U13437 ( .IN1(n9433), .IN2(g3917), .QN(n12964) );
  NAND3X0 U13438 ( .IN1(n12966), .IN2(g3933), .IN3(n9318), .QN(n12963) );
  NAND2X0 U13439 ( .IN1(n9810), .IN2(n12933), .QN(n12966) );
  NOR2X0 U13440 ( .IN1(g3857), .IN2(n8771), .QN(n9810) );
  NAND3X0 U13441 ( .IN1(n12967), .IN2(n12968), .IN3(n12969), .QN(g30443) );
  NAND2X0 U13442 ( .IN1(n3962), .IN2(n12937), .QN(n12969) );
  NAND2X0 U13443 ( .IN1(n9433), .IN2(g3909), .QN(n12968) );
  NAND3X0 U13444 ( .IN1(n12970), .IN2(g3929), .IN3(n9318), .QN(n12967) );
  NAND2X0 U13445 ( .IN1(n12056), .IN2(n12937), .QN(n12970) );
  NAND3X0 U13446 ( .IN1(n12971), .IN2(n12972), .IN3(n12973), .QN(g30442) );
  NAND2X0 U13447 ( .IN1(n3962), .IN2(n12043), .QN(n12973) );
  NAND2X0 U13448 ( .IN1(n9433), .IN2(g3901), .QN(n12972) );
  NAND3X0 U13449 ( .IN1(n12974), .IN2(g3925), .IN3(n9318), .QN(n12971) );
  NAND2X0 U13450 ( .IN1(n12056), .IN2(n12043), .QN(n12974) );
  NOR2X0 U13451 ( .IN1(g3873), .IN2(n5564), .QN(n12043) );
  NAND3X0 U13452 ( .IN1(n12975), .IN2(n12976), .IN3(n12977), .QN(g30441) );
  NAND2X0 U13453 ( .IN1(n3962), .IN2(n12927), .QN(n12977) );
  NAND2X0 U13454 ( .IN1(n9434), .IN2(g3893), .QN(n12976) );
  NAND3X0 U13455 ( .IN1(n12978), .IN2(g3921), .IN3(n9318), .QN(n12975) );
  NAND2X0 U13456 ( .IN1(n12056), .IN2(n12927), .QN(n12978) );
  NOR2X0 U13457 ( .IN1(g3881), .IN2(n5387), .QN(n12927) );
  NAND3X0 U13458 ( .IN1(n12979), .IN2(n12980), .IN3(n12981), .QN(g30440) );
  NAND2X0 U13459 ( .IN1(n3962), .IN2(n12933), .QN(n12981) );
  NAND2X0 U13460 ( .IN1(test_so24), .IN2(n9515), .QN(n12980) );
  NAND3X0 U13461 ( .IN1(n12982), .IN2(g3917), .IN3(n9319), .QN(n12979) );
  NAND2X0 U13462 ( .IN1(n12056), .IN2(n12933), .QN(n12982) );
  NOR2X0 U13463 ( .IN1(g3881), .IN2(g3873), .QN(n12933) );
  NOR2X0 U13464 ( .IN1(g3863), .IN2(n5572), .QN(n12056) );
  NAND3X0 U13465 ( .IN1(n12983), .IN2(n12984), .IN3(n12985), .QN(g30439) );
  NAND2X0 U13466 ( .IN1(n9434), .IN2(g3913), .QN(n12985) );
  NAND3X0 U13467 ( .IN1(n9354), .IN2(g3909), .IN3(n12986), .QN(n12984) );
  INVX0 U13468 ( .INP(n3967), .ZN(n12986) );
  NAND2X0 U13469 ( .IN1(n3967), .IN2(n3765), .QN(n12983) );
  NAND3X0 U13470 ( .IN1(n12987), .IN2(n12988), .IN3(n12989), .QN(g30438) );
  NAND2X0 U13471 ( .IN1(n9434), .IN2(g3905), .QN(n12989) );
  NAND3X0 U13472 ( .IN1(n9353), .IN2(g3901), .IN3(n12990), .QN(n12988) );
  INVX0 U13473 ( .INP(n3970), .ZN(n12990) );
  NAND2X0 U13474 ( .IN1(n3970), .IN2(n3765), .QN(n12987) );
  NAND3X0 U13475 ( .IN1(n12991), .IN2(n12992), .IN3(n12993), .QN(g30437) );
  NAND2X0 U13476 ( .IN1(n9434), .IN2(g3897), .QN(n12993) );
  NAND3X0 U13477 ( .IN1(n9354), .IN2(g3893), .IN3(n12994), .QN(n12992) );
  INVX0 U13478 ( .INP(n3972), .ZN(n12994) );
  NAND2X0 U13479 ( .IN1(n3972), .IN2(n3765), .QN(n12991) );
  NAND3X0 U13480 ( .IN1(n12995), .IN2(n12996), .IN3(n12997), .QN(g30436) );
  NAND2X0 U13481 ( .IN1(n9435), .IN2(g3881), .QN(n12997) );
  NAND3X0 U13482 ( .IN1(test_so24), .IN2(n9317), .IN3(n12998), .QN(n12996) );
  INVX0 U13483 ( .INP(n3974), .ZN(n12998) );
  NAND2X0 U13484 ( .IN1(n3974), .IN2(n3765), .QN(n12995) );
  NOR2X0 U13485 ( .IN1(g3857), .IN2(n12049), .QN(g30435) );
  NAND3X0 U13486 ( .IN1(n9354), .IN2(n8868), .IN3(n12039), .QN(n12049) );
  NAND3X0 U13487 ( .IN1(g4093), .IN2(g4087), .IN3(n3799), .QN(n12039) );
  NAND3X0 U13488 ( .IN1(n12999), .IN2(n13000), .IN3(n13001), .QN(g30434) );
  NAND2X0 U13489 ( .IN1(n9435), .IN2(g3610), .QN(n13001) );
  NAND2X0 U13490 ( .IN1(n13002), .IN2(g3614), .QN(n13000) );
  NAND2X0 U13491 ( .IN1(n13003), .IN2(n3765), .QN(n12999) );
  NAND3X0 U13492 ( .IN1(n13004), .IN2(n13005), .IN3(n13006), .QN(g30433) );
  NAND2X0 U13493 ( .IN1(n13007), .IN2(n3765), .QN(n13006) );
  NAND3X0 U13494 ( .IN1(n13008), .IN2(g3562), .IN3(n9319), .QN(n13005) );
  INVX0 U13495 ( .INP(n13007), .ZN(n13008) );
  NOR2X0 U13496 ( .IN1(n430), .IN2(n5645), .QN(n13007) );
  INVX0 U13497 ( .INP(n12064), .ZN(n430) );
  NAND2X0 U13498 ( .IN1(n9435), .IN2(g3606), .QN(n13004) );
  NAND3X0 U13499 ( .IN1(n13009), .IN2(n13010), .IN3(n13011), .QN(g30432) );
  NAND2X0 U13500 ( .IN1(n13012), .IN2(n3765), .QN(n13011) );
  NAND3X0 U13501 ( .IN1(g3554), .IN2(n12062), .IN3(n9319), .QN(n13010) );
  INVX0 U13502 ( .INP(n13012), .ZN(n12062) );
  NOR2X0 U13503 ( .IN1(n434), .IN2(n5645), .QN(n13012) );
  INVX0 U13504 ( .INP(n13013), .ZN(n434) );
  NAND2X0 U13505 ( .IN1(test_so43), .IN2(n9515), .QN(n13009) );
  NAND3X0 U13506 ( .IN1(n13014), .IN2(n13015), .IN3(n13016), .QN(g30431) );
  NAND2X0 U13507 ( .IN1(n13017), .IN2(n3765), .QN(n13016) );
  NAND3X0 U13508 ( .IN1(n13018), .IN2(g3546), .IN3(n9319), .QN(n13015) );
  INVX0 U13509 ( .INP(n13017), .ZN(n13018) );
  NOR2X0 U13510 ( .IN1(n432), .IN2(n5645), .QN(n13017) );
  INVX0 U13511 ( .INP(n13019), .ZN(n432) );
  NAND2X0 U13512 ( .IN1(n9435), .IN2(g3598), .QN(n13014) );
  NAND3X0 U13513 ( .IN1(n13020), .IN2(n13021), .IN3(n13022), .QN(g30430) );
  NAND2X0 U13514 ( .IN1(n3984), .IN2(n13023), .QN(n13022) );
  NAND2X0 U13515 ( .IN1(n9435), .IN2(g3594), .QN(n13021) );
  NAND3X0 U13516 ( .IN1(n13024), .IN2(g3610), .IN3(n9319), .QN(n13020) );
  NAND2X0 U13517 ( .IN1(n13023), .IN2(n9670), .QN(n13024) );
  NAND3X0 U13518 ( .IN1(n13025), .IN2(n13026), .IN3(n13027), .QN(g30429) );
  NAND2X0 U13519 ( .IN1(n3984), .IN2(n12064), .QN(n13027) );
  NAND2X0 U13520 ( .IN1(n9435), .IN2(g3590), .QN(n13026) );
  NAND3X0 U13521 ( .IN1(n13028), .IN2(g3606), .IN3(n9320), .QN(n13025) );
  NAND2X0 U13522 ( .IN1(n12064), .IN2(n9670), .QN(n13028) );
  NAND3X0 U13523 ( .IN1(n13029), .IN2(n13030), .IN3(n13031), .QN(g30428) );
  NAND2X0 U13524 ( .IN1(n3984), .IN2(n13013), .QN(n13031) );
  NAND2X0 U13525 ( .IN1(n9436), .IN2(g3586), .QN(n13030) );
  NAND3X0 U13526 ( .IN1(test_so43), .IN2(n13032), .IN3(n9320), .QN(n13029) );
  NAND2X0 U13527 ( .IN1(n13013), .IN2(n9670), .QN(n13032) );
  NAND3X0 U13528 ( .IN1(n13033), .IN2(n13034), .IN3(n13035), .QN(g30427) );
  NAND2X0 U13529 ( .IN1(n3984), .IN2(n13019), .QN(n13035) );
  NAND2X0 U13530 ( .IN1(n9436), .IN2(g3582), .QN(n13034) );
  NAND3X0 U13531 ( .IN1(n13036), .IN2(g3598), .IN3(n9320), .QN(n13033) );
  NAND2X0 U13532 ( .IN1(n13019), .IN2(n9670), .QN(n13036) );
  NOR2X0 U13533 ( .IN1(n5576), .IN2(n8767), .QN(n9670) );
  NAND3X0 U13534 ( .IN1(n13037), .IN2(n13038), .IN3(n13039), .QN(g30426) );
  NAND2X0 U13535 ( .IN1(n3990), .IN2(n13023), .QN(n13039) );
  NAND2X0 U13536 ( .IN1(n9436), .IN2(g3578), .QN(n13038) );
  NAND3X0 U13537 ( .IN1(n13040), .IN2(g3594), .IN3(n9320), .QN(n13037) );
  NAND2X0 U13538 ( .IN1(n13023), .IN2(n9669), .QN(n13040) );
  NAND3X0 U13539 ( .IN1(n13041), .IN2(n13042), .IN3(n13043), .QN(g30425) );
  NAND2X0 U13540 ( .IN1(n3990), .IN2(n12064), .QN(n13043) );
  NAND2X0 U13541 ( .IN1(n9437), .IN2(g3574), .QN(n13042) );
  NAND3X0 U13542 ( .IN1(n13044), .IN2(g3590), .IN3(n9320), .QN(n13041) );
  NAND2X0 U13543 ( .IN1(n12064), .IN2(n9669), .QN(n13044) );
  NAND3X0 U13544 ( .IN1(n13045), .IN2(n13046), .IN3(n13047), .QN(g30424) );
  NAND2X0 U13545 ( .IN1(n3990), .IN2(n13013), .QN(n13047) );
  NAND2X0 U13546 ( .IN1(n9437), .IN2(g3570), .QN(n13046) );
  NAND3X0 U13547 ( .IN1(n13048), .IN2(g3586), .IN3(n9320), .QN(n13045) );
  NAND2X0 U13548 ( .IN1(n13013), .IN2(n9669), .QN(n13048) );
  NAND3X0 U13549 ( .IN1(n13049), .IN2(n13050), .IN3(n13051), .QN(g30423) );
  NAND2X0 U13550 ( .IN1(n3990), .IN2(n13019), .QN(n13051) );
  NAND2X0 U13551 ( .IN1(n9437), .IN2(g3566), .QN(n13050) );
  NAND3X0 U13552 ( .IN1(n13052), .IN2(g3582), .IN3(n9320), .QN(n13049) );
  NAND2X0 U13553 ( .IN1(n13019), .IN2(n9669), .QN(n13052) );
  NOR2X0 U13554 ( .IN1(g3506), .IN2(n8767), .QN(n9669) );
  NAND3X0 U13555 ( .IN1(n13053), .IN2(n13054), .IN3(n13055), .QN(g30422) );
  NAND2X0 U13556 ( .IN1(n3995), .IN2(n13023), .QN(n13055) );
  NAND2X0 U13557 ( .IN1(n9438), .IN2(g3558), .QN(n13054) );
  NAND3X0 U13558 ( .IN1(n13056), .IN2(g3578), .IN3(n9321), .QN(n13053) );
  NAND2X0 U13559 ( .IN1(n13023), .IN2(n12077), .QN(n13056) );
  NAND3X0 U13560 ( .IN1(n13057), .IN2(n13058), .IN3(n13059), .QN(g30421) );
  NAND2X0 U13561 ( .IN1(n3995), .IN2(n12064), .QN(n13059) );
  NAND2X0 U13562 ( .IN1(n9438), .IN2(g3550), .QN(n13058) );
  NAND3X0 U13563 ( .IN1(n13060), .IN2(g3574), .IN3(n9321), .QN(n13057) );
  NAND2X0 U13564 ( .IN1(n12064), .IN2(n12077), .QN(n13060) );
  NOR2X0 U13565 ( .IN1(g3522), .IN2(n5569), .QN(n12064) );
  NAND3X0 U13566 ( .IN1(n13061), .IN2(n13062), .IN3(n13063), .QN(g30420) );
  NAND2X0 U13567 ( .IN1(n3995), .IN2(n13013), .QN(n13063) );
  NAND2X0 U13568 ( .IN1(g3542), .IN2(n9513), .QN(n13062) );
  NAND3X0 U13569 ( .IN1(n13064), .IN2(g3570), .IN3(n9321), .QN(n13061) );
  NAND2X0 U13570 ( .IN1(n13013), .IN2(n12077), .QN(n13064) );
  NOR2X0 U13571 ( .IN1(g3530), .IN2(n5383), .QN(n13013) );
  NAND3X0 U13572 ( .IN1(n13065), .IN2(n13066), .IN3(n13067), .QN(g30419) );
  NAND2X0 U13573 ( .IN1(n3995), .IN2(n13019), .QN(n13067) );
  NAND2X0 U13574 ( .IN1(n9439), .IN2(g3538), .QN(n13066) );
  NAND3X0 U13575 ( .IN1(n13068), .IN2(g3566), .IN3(n9321), .QN(n13065) );
  NAND2X0 U13576 ( .IN1(n13019), .IN2(n12077), .QN(n13068) );
  NOR2X0 U13577 ( .IN1(g3512), .IN2(n5576), .QN(n12077) );
  NOR2X0 U13578 ( .IN1(g3522), .IN2(g3530), .QN(n13019) );
  NAND3X0 U13579 ( .IN1(n13069), .IN2(n13070), .IN3(n13071), .QN(g30418) );
  NAND2X0 U13580 ( .IN1(n9439), .IN2(g3562), .QN(n13071) );
  NAND3X0 U13581 ( .IN1(n9354), .IN2(g3558), .IN3(n13072), .QN(n13070) );
  INVX0 U13582 ( .INP(n4000), .ZN(n13072) );
  NAND2X0 U13583 ( .IN1(n4000), .IN2(n3765), .QN(n13069) );
  NAND3X0 U13584 ( .IN1(n13073), .IN2(n13074), .IN3(n13075), .QN(g30417) );
  NAND2X0 U13585 ( .IN1(g3554), .IN2(n9513), .QN(n13075) );
  NAND3X0 U13586 ( .IN1(n9354), .IN2(g3550), .IN3(n13076), .QN(n13074) );
  INVX0 U13587 ( .INP(n4003), .ZN(n13076) );
  NAND2X0 U13588 ( .IN1(n4003), .IN2(n3765), .QN(n13073) );
  NAND3X0 U13589 ( .IN1(n13077), .IN2(n13078), .IN3(n13079), .QN(g30416) );
  NAND2X0 U13590 ( .IN1(n9439), .IN2(g3546), .QN(n13079) );
  NAND3X0 U13591 ( .IN1(g3542), .IN2(n9315), .IN3(n13080), .QN(n13078) );
  INVX0 U13592 ( .INP(n4005), .ZN(n13080) );
  NAND2X0 U13593 ( .IN1(n4005), .IN2(n3765), .QN(n13077) );
  NAND3X0 U13594 ( .IN1(n13081), .IN2(n13082), .IN3(n13083), .QN(g30415) );
  NAND2X0 U13595 ( .IN1(n9440), .IN2(g3530), .QN(n13083) );
  NAND3X0 U13596 ( .IN1(n9354), .IN2(g3538), .IN3(n13084), .QN(n13082) );
  INVX0 U13597 ( .INP(n4007), .ZN(n13084) );
  NAND2X0 U13598 ( .IN1(n4007), .IN2(n3765), .QN(n13081) );
  NOR2X0 U13599 ( .IN1(g3506), .IN2(n12070), .QN(g30414) );
  NAND3X0 U13600 ( .IN1(n12060), .IN2(n9315), .IN3(n5645), .QN(n12070) );
  NAND3X0 U13601 ( .IN1(n5480), .IN2(g4093), .IN3(n3799), .QN(n12060) );
  NAND3X0 U13602 ( .IN1(n13085), .IN2(n13086), .IN3(n13087), .QN(g30413) );
  NAND2X0 U13603 ( .IN1(test_so84), .IN2(n9512), .QN(n13087) );
  NAND2X0 U13604 ( .IN1(n13088), .IN2(g3263), .QN(n13086) );
  NAND2X0 U13605 ( .IN1(n3765), .IN2(n11365), .QN(n13085) );
  NAND3X0 U13606 ( .IN1(n13089), .IN2(n13090), .IN3(n13091), .QN(g30412) );
  NAND2X0 U13607 ( .IN1(n13092), .IN2(n3765), .QN(n13091) );
  NAND3X0 U13608 ( .IN1(n13093), .IN2(g3211), .IN3(n9321), .QN(n13090) );
  INVX0 U13609 ( .INP(n13092), .ZN(n13093) );
  NOR2X0 U13610 ( .IN1(n536), .IN2(n5652), .QN(n13092) );
  INVX0 U13611 ( .INP(n13094), .ZN(n536) );
  NAND2X0 U13612 ( .IN1(n9440), .IN2(g3255), .QN(n13089) );
  NAND3X0 U13613 ( .IN1(n13095), .IN2(n13096), .IN3(n13097), .QN(g30411) );
  NAND2X0 U13614 ( .IN1(n13098), .IN2(n3765), .QN(n13097) );
  NAND3X0 U13615 ( .IN1(n12084), .IN2(g3203), .IN3(n9321), .QN(n13096) );
  INVX0 U13616 ( .INP(n13098), .ZN(n12084) );
  NOR2X0 U13617 ( .IN1(n538), .IN2(n5652), .QN(n13098) );
  INVX0 U13618 ( .INP(n13099), .ZN(n538) );
  NAND2X0 U13619 ( .IN1(n9441), .IN2(g3251), .QN(n13095) );
  NAND3X0 U13620 ( .IN1(n13100), .IN2(n13101), .IN3(n13102), .QN(g30410) );
  NAND2X0 U13621 ( .IN1(n13103), .IN2(n3765), .QN(n13102) );
  NAND3X0 U13622 ( .IN1(test_so88), .IN2(n13104), .IN3(n9321), .QN(n13101) );
  INVX0 U13623 ( .INP(n13103), .ZN(n13104) );
  NOR2X0 U13624 ( .IN1(n537), .IN2(n5652), .QN(n13103) );
  INVX0 U13625 ( .INP(n13105), .ZN(n537) );
  NAND2X0 U13626 ( .IN1(n9441), .IN2(g3247), .QN(n13100) );
  NAND3X0 U13627 ( .IN1(n13106), .IN2(n13107), .IN3(n13108), .QN(g30409) );
  NAND2X0 U13628 ( .IN1(n4015), .IN2(n9686), .QN(n13108) );
  NAND2X0 U13629 ( .IN1(g3243), .IN2(n9511), .QN(n13107) );
  NAND3X0 U13630 ( .IN1(test_so84), .IN2(n13109), .IN3(n9321), .QN(n13106) );
  NAND2X0 U13631 ( .IN1(n9686), .IN2(n9659), .QN(n13109) );
  NAND3X0 U13632 ( .IN1(n13110), .IN2(n13111), .IN3(n13112), .QN(g30408) );
  NAND2X0 U13633 ( .IN1(n4015), .IN2(n13094), .QN(n13112) );
  NAND2X0 U13634 ( .IN1(n9441), .IN2(g3239), .QN(n13111) );
  NAND3X0 U13635 ( .IN1(n13113), .IN2(g3255), .IN3(n9323), .QN(n13110) );
  NAND2X0 U13636 ( .IN1(n13094), .IN2(n9659), .QN(n13113) );
  NAND3X0 U13637 ( .IN1(n13114), .IN2(n13115), .IN3(n13116), .QN(g30407) );
  NAND2X0 U13638 ( .IN1(n4015), .IN2(n13099), .QN(n13116) );
  NAND2X0 U13639 ( .IN1(n9441), .IN2(g3235), .QN(n13115) );
  NAND3X0 U13640 ( .IN1(n13117), .IN2(g3251), .IN3(n9323), .QN(n13114) );
  NAND2X0 U13641 ( .IN1(n13099), .IN2(n9659), .QN(n13117) );
  NAND3X0 U13642 ( .IN1(n13118), .IN2(n13119), .IN3(n13120), .QN(g30406) );
  NAND2X0 U13643 ( .IN1(n4015), .IN2(n13105), .QN(n13120) );
  NAND2X0 U13644 ( .IN1(n9442), .IN2(g3231), .QN(n13119) );
  NAND3X0 U13645 ( .IN1(n13121), .IN2(g3247), .IN3(n9323), .QN(n13118) );
  NAND2X0 U13646 ( .IN1(n13105), .IN2(n9659), .QN(n13121) );
  NOR2X0 U13647 ( .IN1(n5366), .IN2(n8752), .QN(n9659) );
  NAND3X0 U13648 ( .IN1(n13122), .IN2(n13123), .IN3(n13124), .QN(g30405) );
  NAND2X0 U13649 ( .IN1(n4022), .IN2(n9686), .QN(n13124) );
  NAND2X0 U13650 ( .IN1(n9442), .IN2(g3227), .QN(n13123) );
  NAND3X0 U13651 ( .IN1(g3243), .IN2(n13125), .IN3(n9323), .QN(n13122) );
  NAND2X0 U13652 ( .IN1(n9686), .IN2(n9658), .QN(n13125) );
  NAND3X0 U13653 ( .IN1(n13126), .IN2(n13127), .IN3(n13128), .QN(g30404) );
  NAND2X0 U13654 ( .IN1(n4022), .IN2(n13094), .QN(n13128) );
  NAND2X0 U13655 ( .IN1(n9442), .IN2(g3223), .QN(n13127) );
  NAND3X0 U13656 ( .IN1(n13129), .IN2(g3239), .IN3(n9323), .QN(n13126) );
  NAND2X0 U13657 ( .IN1(n13094), .IN2(n9658), .QN(n13129) );
  NAND3X0 U13658 ( .IN1(n13130), .IN2(n13131), .IN3(n13132), .QN(g30403) );
  NAND2X0 U13659 ( .IN1(n4022), .IN2(n13099), .QN(n13132) );
  NAND2X0 U13660 ( .IN1(n9442), .IN2(g3219), .QN(n13131) );
  NAND3X0 U13661 ( .IN1(n13133), .IN2(g3235), .IN3(n9323), .QN(n13130) );
  NAND2X0 U13662 ( .IN1(n13099), .IN2(n9658), .QN(n13133) );
  NAND3X0 U13663 ( .IN1(n13134), .IN2(n13135), .IN3(n13136), .QN(g30402) );
  NAND2X0 U13664 ( .IN1(n4022), .IN2(n13105), .QN(n13136) );
  NAND2X0 U13665 ( .IN1(n9443), .IN2(g3215), .QN(n13135) );
  NAND3X0 U13666 ( .IN1(n13137), .IN2(g3231), .IN3(n9323), .QN(n13134) );
  NAND2X0 U13667 ( .IN1(n13105), .IN2(n9658), .QN(n13137) );
  NOR2X0 U13668 ( .IN1(g3155), .IN2(n8752), .QN(n9658) );
  NAND3X0 U13669 ( .IN1(n13138), .IN2(n13139), .IN3(n13140), .QN(g30401) );
  NAND2X0 U13670 ( .IN1(n4027), .IN2(n9686), .QN(n13140) );
  NAND2X0 U13671 ( .IN1(n9443), .IN2(g3207), .QN(n13139) );
  NAND3X0 U13672 ( .IN1(n13141), .IN2(g3227), .IN3(n9323), .QN(n13138) );
  NAND2X0 U13673 ( .IN1(n9686), .IN2(n12096), .QN(n13141) );
  NAND3X0 U13674 ( .IN1(n13142), .IN2(n13143), .IN3(n13144), .QN(g30400) );
  NAND2X0 U13675 ( .IN1(n4027), .IN2(n13094), .QN(n13144) );
  NAND2X0 U13676 ( .IN1(n9443), .IN2(g3199), .QN(n13143) );
  NAND3X0 U13677 ( .IN1(n13145), .IN2(g3223), .IN3(n9323), .QN(n13142) );
  NAND2X0 U13678 ( .IN1(n13094), .IN2(n12096), .QN(n13145) );
  NOR2X0 U13679 ( .IN1(g3171), .IN2(n5390), .QN(n13094) );
  NAND3X0 U13680 ( .IN1(n13146), .IN2(n13147), .IN3(n13148), .QN(g30399) );
  NAND2X0 U13681 ( .IN1(n4027), .IN2(n13099), .QN(n13148) );
  NAND2X0 U13682 ( .IN1(n9443), .IN2(g3191), .QN(n13147) );
  NAND3X0 U13683 ( .IN1(n13149), .IN2(g3219), .IN3(n9346), .QN(n13146) );
  NAND2X0 U13684 ( .IN1(n13099), .IN2(n12096), .QN(n13149) );
  NOR2X0 U13685 ( .IN1(g3179), .IN2(n5603), .QN(n13099) );
  NAND3X0 U13686 ( .IN1(n13150), .IN2(n13151), .IN3(n13152), .QN(g30398) );
  NAND2X0 U13687 ( .IN1(n4027), .IN2(n13105), .QN(n13152) );
  NAND2X0 U13688 ( .IN1(n9464), .IN2(g3187), .QN(n13151) );
  NAND3X0 U13689 ( .IN1(n13153), .IN2(g3215), .IN3(n9347), .QN(n13150) );
  NAND2X0 U13690 ( .IN1(n13105), .IN2(n12096), .QN(n13153) );
  NOR2X0 U13691 ( .IN1(g3161), .IN2(n5366), .QN(n12096) );
  NOR2X0 U13692 ( .IN1(g3171), .IN2(g3179), .QN(n13105) );
  NAND3X0 U13693 ( .IN1(n13154), .IN2(n13155), .IN3(n13156), .QN(g30397) );
  NAND2X0 U13694 ( .IN1(n9462), .IN2(g3211), .QN(n13156) );
  NAND3X0 U13695 ( .IN1(n9349), .IN2(g3207), .IN3(n13157), .QN(n13155) );
  INVX0 U13696 ( .INP(n4032), .ZN(n13157) );
  NAND2X0 U13697 ( .IN1(n4032), .IN2(n3765), .QN(n13154) );
  NAND3X0 U13698 ( .IN1(n13158), .IN2(n13159), .IN3(n13160), .QN(g30396) );
  NAND2X0 U13699 ( .IN1(n9461), .IN2(g3203), .QN(n13160) );
  NAND3X0 U13700 ( .IN1(n9354), .IN2(g3199), .IN3(n13161), .QN(n13159) );
  INVX0 U13701 ( .INP(n4035), .ZN(n13161) );
  NAND2X0 U13702 ( .IN1(n4035), .IN2(n3765), .QN(n13158) );
  NAND3X0 U13703 ( .IN1(n13162), .IN2(n13163), .IN3(n13164), .QN(g30395) );
  NAND2X0 U13704 ( .IN1(test_so88), .IN2(n9512), .QN(n13164) );
  NAND3X0 U13705 ( .IN1(n9354), .IN2(g3191), .IN3(n13165), .QN(n13163) );
  INVX0 U13706 ( .INP(n4037), .ZN(n13165) );
  NAND2X0 U13707 ( .IN1(n4037), .IN2(n3765), .QN(n13162) );
  NAND3X0 U13708 ( .IN1(n13166), .IN2(n13167), .IN3(n13168), .QN(g30394) );
  NAND2X0 U13709 ( .IN1(n9459), .IN2(g3179), .QN(n13168) );
  NAND3X0 U13710 ( .IN1(n9354), .IN2(g3187), .IN3(n13169), .QN(n13167) );
  INVX0 U13711 ( .INP(n4039), .ZN(n13169) );
  NAND2X0 U13712 ( .IN1(n4039), .IN2(n3765), .QN(n13166) );
  NOR3X0 U13713 ( .IN1(n12091), .IN2(n9384), .IN3(g3155), .QN(g30393) );
  NAND2X0 U13714 ( .IN1(n5652), .IN2(n12083), .QN(n12091) );
  NAND2X0 U13715 ( .IN1(n3799), .IN2(n11355), .QN(n12083) );
  NAND2X0 U13716 ( .IN1(n13170), .IN2(n13171), .QN(g30392) );
  NAND2X0 U13717 ( .IN1(n9473), .IN2(g2803), .QN(n13171) );
  NAND2X0 U13718 ( .IN1(n13172), .IN2(n13173), .QN(g30391) );
  NAND2X0 U13719 ( .IN1(n9457), .IN2(g2771), .QN(n13173) );
  NAND2X0 U13720 ( .IN1(n13170), .IN2(n13174), .QN(g30390) );
  NAND2X0 U13721 ( .IN1(g2834), .IN2(n9511), .QN(n13174) );
  NAND2X0 U13722 ( .IN1(n13175), .IN2(n9375), .QN(n13170) );
  NAND2X0 U13723 ( .IN1(n13176), .IN2(n13177), .QN(n13175) );
  NAND4X0 U13724 ( .IN1(n13178), .IN2(n13179), .IN3(n13180), .IN4(n13181), 
        .QN(n13177) );
  NOR2X0 U13725 ( .IN1(n13182), .IN2(n13183), .QN(n13180) );
  NOR2X0 U13726 ( .IN1(n13184), .IN2(g2236), .QN(n13183) );
  NOR2X0 U13727 ( .IN1(n1296), .IN2(g2370), .QN(n13182) );
  NAND2X0 U13728 ( .IN1(n8789), .IN2(n13185), .QN(n13179) );
  NAND2X0 U13729 ( .IN1(n8761), .IN2(n13186), .QN(n13178) );
  NAND4X0 U13730 ( .IN1(n13187), .IN2(n13188), .IN3(n13189), .IN4(n13190), 
        .QN(n13176) );
  NOR2X0 U13731 ( .IN1(n13191), .IN2(n13192), .QN(n13189) );
  NOR2X0 U13732 ( .IN1(n5545), .IN2(n13184), .QN(n13192) );
  NOR2X0 U13733 ( .IN1(n5379), .IN2(n1296), .QN(n13191) );
  NAND2X0 U13734 ( .IN1(n13185), .IN2(g2819), .QN(n13188) );
  NAND2X0 U13735 ( .IN1(n13186), .IN2(g2815), .QN(n13187) );
  NAND2X0 U13736 ( .IN1(n13172), .IN2(n13193), .QN(g30389) );
  NAND2X0 U13737 ( .IN1(g2831), .IN2(n9513), .QN(n13193) );
  NAND2X0 U13738 ( .IN1(n13194), .IN2(n9375), .QN(n13172) );
  NAND2X0 U13739 ( .IN1(n13195), .IN2(n13196), .QN(n13194) );
  NAND4X0 U13740 ( .IN1(n13197), .IN2(n13198), .IN3(n13199), .IN4(n13181), 
        .QN(n13196) );
  NOR2X0 U13741 ( .IN1(n13200), .IN2(n13201), .QN(n13199) );
  NOR2X0 U13742 ( .IN1(n13184), .IN2(g1677), .QN(n13201) );
  NOR2X0 U13743 ( .IN1(n1296), .IN2(g1811), .QN(n13200) );
  NAND2X0 U13744 ( .IN1(n8790), .IN2(n13185), .QN(n13198) );
  NAND2X0 U13745 ( .IN1(n13186), .IN2(n8905), .QN(n13197) );
  NAND4X0 U13746 ( .IN1(n13202), .IN2(n13203), .IN3(n13204), .IN4(n13190), 
        .QN(n13195) );
  INVX0 U13747 ( .INP(n13181), .ZN(n13190) );
  NAND3X0 U13748 ( .IN1(n3653), .IN2(n13205), .IN3(n5600), .QN(n13181) );
  NOR3X0 U13749 ( .IN1(g2741), .IN2(test_so30), .IN3(g2748), .QN(n3653) );
  NOR2X0 U13750 ( .IN1(n13206), .IN2(n13207), .QN(n13204) );
  NOR2X0 U13751 ( .IN1(n5544), .IN2(n13184), .QN(n13207) );
  INVX0 U13752 ( .INP(n13208), .ZN(n13184) );
  NOR2X0 U13753 ( .IN1(n5378), .IN2(n1296), .QN(n13206) );
  INVX0 U13754 ( .INP(n13209), .ZN(n1296) );
  NAND2X0 U13755 ( .IN1(n13185), .IN2(g2787), .QN(n13203) );
  NAND2X0 U13756 ( .IN1(n13186), .IN2(g2783), .QN(n13202) );
  NAND2X0 U13757 ( .IN1(n13210), .IN2(n13211), .QN(g30388) );
  NAND3X0 U13758 ( .IN1(n12405), .IN2(n13212), .IN3(n3730), .QN(n13211) );
  NAND2X0 U13759 ( .IN1(n5349), .IN2(n3506), .QN(n13212) );
  INVX0 U13760 ( .INP(n13213), .ZN(n3506) );
  NAND2X0 U13761 ( .IN1(n13213), .IN2(g2741), .QN(n12405) );
  NOR2X0 U13762 ( .IN1(n13214), .IN2(n5600), .QN(n13213) );
  NAND2X0 U13763 ( .IN1(n9456), .IN2(g2735), .QN(n13210) );
  NAND3X0 U13764 ( .IN1(n13215), .IN2(n13216), .IN3(n13217), .QN(g30387) );
  INVX0 U13765 ( .INP(n13218), .ZN(n13217) );
  NOR2X0 U13766 ( .IN1(n13219), .IN2(n15960), .QN(n13218) );
  INVX0 U13767 ( .INP(n13220), .ZN(n13216) );
  NOR2X0 U13768 ( .IN1(n13221), .IN2(n5777), .QN(n13220) );
  NOR2X0 U13769 ( .IN1(n13222), .IN2(n9388), .QN(n13221) );
  NOR2X0 U13770 ( .IN1(n13223), .IN2(n5457), .QN(n13222) );
  NAND3X0 U13771 ( .IN1(n13224), .IN2(n5457), .IN3(n5777), .QN(n13215) );
  NAND2X0 U13772 ( .IN1(n13225), .IN2(n13226), .QN(g30386) );
  INVX0 U13773 ( .INP(n13227), .ZN(n13226) );
  NOR2X0 U13774 ( .IN1(n13219), .IN2(n5777), .QN(n13227) );
  NAND2X0 U13775 ( .IN1(n13219), .IN2(g2675), .QN(n13225) );
  NAND3X0 U13776 ( .IN1(n13228), .IN2(n13229), .IN3(n13230), .QN(g30385) );
  NAND2X0 U13777 ( .IN1(n9455), .IN2(g2657), .QN(n13230) );
  NAND2X0 U13778 ( .IN1(n13231), .IN2(g2661), .QN(n13229) );
  INVX0 U13779 ( .INP(n13219), .ZN(n13231) );
  NAND2X0 U13780 ( .IN1(n13223), .IN2(n9375), .QN(n13219) );
  NAND2X0 U13781 ( .IN1(n13224), .IN2(n5418), .QN(n13228) );
  NAND3X0 U13782 ( .IN1(n13232), .IN2(n13233), .IN3(n13234), .QN(g30384) );
  NAND2X0 U13783 ( .IN1(n9463), .IN2(g2652), .QN(n13234) );
  NAND3X0 U13784 ( .IN1(n3517), .IN2(n13235), .IN3(n8849), .QN(n13233) );
  NAND2X0 U13785 ( .IN1(n13236), .IN2(n13237), .QN(n13235) );
  NAND2X0 U13786 ( .IN1(n8513), .IN2(g2648), .QN(n13237) );
  NAND2X0 U13787 ( .IN1(n8390), .IN2(g2652), .QN(n13236) );
  NAND2X0 U13788 ( .IN1(n13238), .IN2(g2657), .QN(n13232) );
  NAND2X0 U13789 ( .IN1(n12111), .IN2(n13239), .QN(n13238) );
  NAND2X0 U13790 ( .IN1(n9366), .IN2(n12123), .QN(n13239) );
  INVX0 U13791 ( .INP(n8849), .ZN(n12123) );
  NAND2X0 U13792 ( .IN1(n13240), .IN2(n13241), .QN(g30383) );
  NAND2X0 U13793 ( .IN1(test_so66), .IN2(n9428), .QN(n13241) );
  NAND2X0 U13794 ( .IN1(n13242), .IN2(n9376), .QN(n13240) );
  NAND2X0 U13795 ( .IN1(n13243), .IN2(n13244), .QN(n13242) );
  NAND2X0 U13796 ( .IN1(test_so34), .IN2(n13245), .QN(n13244) );
  NAND2X0 U13797 ( .IN1(n13246), .IN2(n13247), .QN(n13243) );
  NAND2X0 U13798 ( .IN1(n5351), .IN2(g2599), .QN(n13247) );
  INVX0 U13799 ( .INP(n13245), .ZN(n13246) );
  NAND3X0 U13800 ( .IN1(n13248), .IN2(g2610), .IN3(n5508), .QN(n13245) );
  NAND3X0 U13801 ( .IN1(n13249), .IN2(n13250), .IN3(n13251), .QN(g30382) );
  NAND2X0 U13802 ( .IN1(n13252), .IN2(n9295), .QN(n13251) );
  INVX0 U13803 ( .INP(n13253), .ZN(n13250) );
  NOR2X0 U13804 ( .IN1(n13254), .IN2(n5782), .QN(n13253) );
  NOR2X0 U13805 ( .IN1(n13255), .IN2(n9387), .QN(n13254) );
  NOR2X0 U13806 ( .IN1(n13256), .IN2(n5461), .QN(n13255) );
  NAND3X0 U13807 ( .IN1(n13257), .IN2(n5461), .IN3(n5782), .QN(n13249) );
  NAND2X0 U13808 ( .IN1(n13258), .IN2(n13259), .QN(g30381) );
  NAND2X0 U13809 ( .IN1(n13252), .IN2(g2547), .QN(n13259) );
  NAND2X0 U13810 ( .IN1(n13260), .IN2(g2541), .QN(n13258) );
  NAND3X0 U13811 ( .IN1(n13261), .IN2(n13262), .IN3(n13263), .QN(g30380) );
  NAND2X0 U13812 ( .IN1(n9469), .IN2(g2523), .QN(n13263) );
  NAND2X0 U13813 ( .IN1(n13252), .IN2(g2527), .QN(n13262) );
  INVX0 U13814 ( .INP(n13260), .ZN(n13252) );
  NAND2X0 U13815 ( .IN1(n13256), .IN2(n9376), .QN(n13260) );
  NAND2X0 U13816 ( .IN1(n13257), .IN2(n5420), .QN(n13261) );
  NAND3X0 U13817 ( .IN1(n13264), .IN2(n13265), .IN3(n13266), .QN(g30379) );
  NAND2X0 U13818 ( .IN1(n9430), .IN2(g2518), .QN(n13266) );
  NAND3X0 U13819 ( .IN1(n3536), .IN2(n13267), .IN3(n8855), .QN(n13265) );
  NAND2X0 U13820 ( .IN1(n13268), .IN2(n13269), .QN(n13267) );
  NAND2X0 U13821 ( .IN1(n8512), .IN2(g2514), .QN(n13269) );
  NAND2X0 U13822 ( .IN1(n8387), .IN2(g2518), .QN(n13268) );
  NAND2X0 U13823 ( .IN1(n13270), .IN2(g2523), .QN(n13264) );
  NAND2X0 U13824 ( .IN1(n12132), .IN2(n13271), .QN(n13270) );
  NAND2X0 U13825 ( .IN1(n9366), .IN2(n12144), .QN(n13271) );
  INVX0 U13826 ( .INP(n8855), .ZN(n12144) );
  NAND2X0 U13827 ( .IN1(n13272), .IN2(n13273), .QN(g30378) );
  NAND2X0 U13828 ( .IN1(n9471), .IN2(g2441), .QN(n13273) );
  NAND2X0 U13829 ( .IN1(n13274), .IN2(n9376), .QN(n13272) );
  NAND2X0 U13830 ( .IN1(n13275), .IN2(n13276), .QN(n13274) );
  NAND2X0 U13831 ( .IN1(n13277), .IN2(g2461), .QN(n13276) );
  NAND2X0 U13832 ( .IN1(n13278), .IN2(n13279), .QN(n13275) );
  NAND2X0 U13833 ( .IN1(g2465), .IN2(n8860), .QN(n13279) );
  INVX0 U13834 ( .INP(n13277), .ZN(n13278) );
  NAND3X0 U13835 ( .IN1(n13280), .IN2(g2476), .IN3(n5509), .QN(n13277) );
  NAND3X0 U13836 ( .IN1(n13281), .IN2(n13282), .IN3(n13283), .QN(g30377) );
  NAND2X0 U13837 ( .IN1(n13284), .IN2(n9324), .QN(n13283) );
  NAND2X0 U13838 ( .IN1(test_so89), .IN2(n13285), .QN(n13282) );
  NAND2X0 U13839 ( .IN1(n13286), .IN2(n9376), .QN(n13285) );
  INVX0 U13840 ( .INP(n13287), .ZN(n13286) );
  NOR2X0 U13841 ( .IN1(n13288), .IN2(n5459), .QN(n13287) );
  NAND3X0 U13842 ( .IN1(n13289), .IN2(n5459), .IN3(n8892), .QN(n13281) );
  NAND2X0 U13843 ( .IN1(n13290), .IN2(n13291), .QN(g30376) );
  NAND2X0 U13844 ( .IN1(test_so89), .IN2(n13284), .QN(n13291) );
  NAND2X0 U13845 ( .IN1(n13292), .IN2(g2407), .QN(n13290) );
  NAND3X0 U13846 ( .IN1(n13293), .IN2(n13294), .IN3(n13295), .QN(g30375) );
  NAND2X0 U13847 ( .IN1(n9453), .IN2(g2389), .QN(n13295) );
  NAND2X0 U13848 ( .IN1(n13284), .IN2(g2393), .QN(n13294) );
  INVX0 U13849 ( .INP(n13292), .ZN(n13284) );
  NAND2X0 U13850 ( .IN1(n13288), .IN2(n9376), .QN(n13292) );
  NAND2X0 U13851 ( .IN1(n13289), .IN2(n5421), .QN(n13293) );
  NAND3X0 U13852 ( .IN1(n13296), .IN2(n13297), .IN3(n13298), .QN(g30374) );
  NAND2X0 U13853 ( .IN1(n9454), .IN2(g2384), .QN(n13298) );
  NAND3X0 U13854 ( .IN1(n3555), .IN2(n13299), .IN3(n8851), .QN(n13297) );
  NAND2X0 U13855 ( .IN1(n13300), .IN2(n13301), .QN(n13299) );
  NAND2X0 U13856 ( .IN1(n8507), .IN2(g2380), .QN(n13301) );
  NAND2X0 U13857 ( .IN1(n8386), .IN2(g2384), .QN(n13300) );
  NAND2X0 U13858 ( .IN1(n13302), .IN2(g2389), .QN(n13296) );
  NAND2X0 U13859 ( .IN1(n12153), .IN2(n13303), .QN(n13302) );
  NAND2X0 U13860 ( .IN1(n9365), .IN2(n12165), .QN(n13303) );
  INVX0 U13861 ( .INP(n8851), .ZN(n12165) );
  NAND2X0 U13862 ( .IN1(n13304), .IN2(n13305), .QN(g30373) );
  NAND2X0 U13863 ( .IN1(n9458), .IN2(g2307), .QN(n13305) );
  NAND2X0 U13864 ( .IN1(n13306), .IN2(n9376), .QN(n13304) );
  NAND2X0 U13865 ( .IN1(n13307), .IN2(n13308), .QN(n13306) );
  NAND2X0 U13866 ( .IN1(n13309), .IN2(g2327), .QN(n13308) );
  NAND2X0 U13867 ( .IN1(n13310), .IN2(n13311), .QN(n13307) );
  NAND2X0 U13868 ( .IN1(n5353), .IN2(g2331), .QN(n13311) );
  INVX0 U13869 ( .INP(n13309), .ZN(n13310) );
  NAND3X0 U13870 ( .IN1(n13312), .IN2(test_so21), .IN3(n5511), .QN(n13309) );
  NAND3X0 U13871 ( .IN1(n13313), .IN2(n13314), .IN3(n13315), .QN(g30372) );
  INVX0 U13872 ( .INP(n13316), .ZN(n13315) );
  NOR2X0 U13873 ( .IN1(n13317), .IN2(n15967), .QN(n13316) );
  INVX0 U13874 ( .INP(n13318), .ZN(n13314) );
  NOR2X0 U13875 ( .IN1(n13319), .IN2(n5778), .QN(n13318) );
  NOR2X0 U13876 ( .IN1(n13320), .IN2(n9388), .QN(n13319) );
  NOR2X0 U13877 ( .IN1(n13321), .IN2(n5458), .QN(n13320) );
  NAND3X0 U13878 ( .IN1(n13322), .IN2(n5458), .IN3(n5778), .QN(n13313) );
  NAND2X0 U13879 ( .IN1(n13323), .IN2(n13324), .QN(g30371) );
  INVX0 U13880 ( .INP(n13325), .ZN(n13324) );
  NOR2X0 U13881 ( .IN1(n13317), .IN2(n5778), .QN(n13325) );
  NAND2X0 U13882 ( .IN1(n13317), .IN2(g2273), .QN(n13323) );
  NAND3X0 U13883 ( .IN1(n13326), .IN2(n13327), .IN3(n13328), .QN(g30370) );
  NAND2X0 U13884 ( .IN1(n9472), .IN2(g2255), .QN(n13328) );
  NAND2X0 U13885 ( .IN1(n13329), .IN2(g2259), .QN(n13327) );
  INVX0 U13886 ( .INP(n13317), .ZN(n13329) );
  NAND2X0 U13887 ( .IN1(n13321), .IN2(n9376), .QN(n13317) );
  NAND2X0 U13888 ( .IN1(n13322), .IN2(n5419), .QN(n13326) );
  NAND3X0 U13889 ( .IN1(n13330), .IN2(n13331), .IN3(n13332), .QN(g30369) );
  NAND2X0 U13890 ( .IN1(n9460), .IN2(g2250), .QN(n13332) );
  NAND3X0 U13891 ( .IN1(n3574), .IN2(n13333), .IN3(n8856), .QN(n13331) );
  NAND2X0 U13892 ( .IN1(n13334), .IN2(n13335), .QN(n13333) );
  NAND2X0 U13893 ( .IN1(n8503), .IN2(g2246), .QN(n13335) );
  NAND2X0 U13894 ( .IN1(n8389), .IN2(g2250), .QN(n13334) );
  NAND2X0 U13895 ( .IN1(n13336), .IN2(g2255), .QN(n13330) );
  NAND2X0 U13896 ( .IN1(n12174), .IN2(n13337), .QN(n13336) );
  NAND2X0 U13897 ( .IN1(n9366), .IN2(n12186), .QN(n13337) );
  INVX0 U13898 ( .INP(n8856), .ZN(n12186) );
  NAND2X0 U13899 ( .IN1(n13338), .IN2(n13339), .QN(g30368) );
  NAND2X0 U13900 ( .IN1(n9443), .IN2(g2173), .QN(n13339) );
  NAND2X0 U13901 ( .IN1(n13340), .IN2(n9376), .QN(n13338) );
  NAND2X0 U13902 ( .IN1(n13341), .IN2(n13342), .QN(n13340) );
  NAND2X0 U13903 ( .IN1(n13343), .IN2(g2193), .QN(n13342) );
  NAND2X0 U13904 ( .IN1(n13344), .IN2(n13345), .QN(n13341) );
  NAND2X0 U13905 ( .IN1(n5356), .IN2(g2197), .QN(n13345) );
  INVX0 U13906 ( .INP(n13343), .ZN(n13344) );
  NAND3X0 U13907 ( .IN1(n13346), .IN2(g2208), .IN3(n5512), .QN(n13343) );
  NAND3X0 U13908 ( .IN1(n13347), .IN2(n13348), .IN3(n13349), .QN(g30367) );
  NAND2X0 U13909 ( .IN1(n13350), .IN2(g2126), .QN(n13349) );
  INVX0 U13910 ( .INP(n13351), .ZN(n13348) );
  NOR2X0 U13911 ( .IN1(n13352), .IN2(n5784), .QN(n13351) );
  NOR2X0 U13912 ( .IN1(n13353), .IN2(n9390), .QN(n13352) );
  NOR2X0 U13913 ( .IN1(n13354), .IN2(n5463), .QN(n13353) );
  NAND3X0 U13914 ( .IN1(n13355), .IN2(n5463), .IN3(n5784), .QN(n13347) );
  NAND2X0 U13915 ( .IN1(n13356), .IN2(n13357), .QN(g30366) );
  NAND2X0 U13916 ( .IN1(n13350), .IN2(g2122), .QN(n13357) );
  NAND2X0 U13917 ( .IN1(n13358), .IN2(g2116), .QN(n13356) );
  NAND3X0 U13918 ( .IN1(n13359), .IN2(n13360), .IN3(n13361), .QN(g30365) );
  NAND2X0 U13919 ( .IN1(n9443), .IN2(g2098), .QN(n13361) );
  NAND2X0 U13920 ( .IN1(n13350), .IN2(g2102), .QN(n13360) );
  INVX0 U13921 ( .INP(n13358), .ZN(n13350) );
  NAND2X0 U13922 ( .IN1(n13354), .IN2(n9376), .QN(n13358) );
  NAND2X0 U13923 ( .IN1(n13355), .IN2(n5666), .QN(n13359) );
  NAND3X0 U13924 ( .IN1(n13362), .IN2(n13363), .IN3(n13364), .QN(g30364) );
  NAND2X0 U13925 ( .IN1(test_so78), .IN2(n9385), .QN(n13364) );
  NAND4X0 U13926 ( .IN1(n8858), .IN2(n3593), .IN3(n13365), .IN4(n13366), .QN(
        n13363) );
  NAND2X0 U13927 ( .IN1(test_so78), .IN2(g2089), .QN(n13366) );
  NAND2X0 U13928 ( .IN1(n8385), .IN2(n8885), .QN(n13365) );
  NAND2X0 U13929 ( .IN1(n13367), .IN2(g2098), .QN(n13362) );
  NAND2X0 U13930 ( .IN1(n12195), .IN2(n13368), .QN(n13367) );
  NAND2X0 U13931 ( .IN1(n9365), .IN2(n12207), .QN(n13368) );
  INVX0 U13932 ( .INP(n8858), .ZN(n12207) );
  NAND2X0 U13933 ( .IN1(n13369), .IN2(n13370), .QN(g30363) );
  NAND2X0 U13934 ( .IN1(n9443), .IN2(g2016), .QN(n13370) );
  NAND2X0 U13935 ( .IN1(n13371), .IN2(n9373), .QN(n13369) );
  NAND2X0 U13936 ( .IN1(n13372), .IN2(n13373), .QN(n13371) );
  NAND2X0 U13937 ( .IN1(test_so59), .IN2(n13374), .QN(n13373) );
  NAND2X0 U13938 ( .IN1(n13375), .IN2(n13376), .QN(n13372) );
  NAND2X0 U13939 ( .IN1(n5355), .IN2(g2040), .QN(n13376) );
  INVX0 U13940 ( .INP(n13374), .ZN(n13375) );
  NAND3X0 U13941 ( .IN1(n13377), .IN2(g2051), .IN3(n5507), .QN(n13374) );
  NAND3X0 U13942 ( .IN1(n13378), .IN2(n13379), .IN3(n13380), .QN(g30362) );
  NAND2X0 U13943 ( .IN1(n13381), .IN2(g1992), .QN(n13380) );
  INVX0 U13944 ( .INP(n13382), .ZN(n13379) );
  NOR2X0 U13945 ( .IN1(n13383), .IN2(n5783), .QN(n13382) );
  NOR2X0 U13946 ( .IN1(n13384), .IN2(n9391), .QN(n13383) );
  NOR2X0 U13947 ( .IN1(n13385), .IN2(n5462), .QN(n13384) );
  NAND3X0 U13948 ( .IN1(n13386), .IN2(n5462), .IN3(n5783), .QN(n13378) );
  NAND2X0 U13949 ( .IN1(n13387), .IN2(n13388), .QN(g30361) );
  NAND2X0 U13950 ( .IN1(n13381), .IN2(g1988), .QN(n13388) );
  NAND2X0 U13951 ( .IN1(n13389), .IN2(g1982), .QN(n13387) );
  NAND3X0 U13952 ( .IN1(n13390), .IN2(n13391), .IN3(n13392), .QN(g30360) );
  NAND2X0 U13953 ( .IN1(n9442), .IN2(g1964), .QN(n13392) );
  NAND2X0 U13954 ( .IN1(n13381), .IN2(g1968), .QN(n13391) );
  INVX0 U13955 ( .INP(n13389), .ZN(n13381) );
  NAND2X0 U13956 ( .IN1(n13385), .IN2(n9376), .QN(n13389) );
  NAND2X0 U13957 ( .IN1(n13386), .IN2(n5664), .QN(n13390) );
  NAND3X0 U13958 ( .IN1(n13393), .IN2(n13394), .IN3(n13395), .QN(g30359) );
  NAND2X0 U13959 ( .IN1(n9442), .IN2(g1959), .QN(n13395) );
  NAND3X0 U13960 ( .IN1(n3611), .IN2(n13396), .IN3(n8848), .QN(n13394) );
  NAND2X0 U13961 ( .IN1(n13397), .IN2(n13398), .QN(n13396) );
  NAND2X0 U13962 ( .IN1(n8511), .IN2(g1955), .QN(n13398) );
  NAND2X0 U13963 ( .IN1(n8383), .IN2(g1959), .QN(n13397) );
  NAND2X0 U13964 ( .IN1(n13399), .IN2(g1964), .QN(n13393) );
  NAND2X0 U13965 ( .IN1(n12216), .IN2(n13400), .QN(n13399) );
  NAND2X0 U13966 ( .IN1(n9366), .IN2(n12228), .QN(n13400) );
  INVX0 U13967 ( .INP(n8848), .ZN(n12228) );
  NAND2X0 U13968 ( .IN1(n13401), .IN2(n13402), .QN(g30358) );
  NAND2X0 U13969 ( .IN1(n9442), .IN2(g1882), .QN(n13402) );
  NAND2X0 U13970 ( .IN1(n13403), .IN2(n9376), .QN(n13401) );
  NAND2X0 U13971 ( .IN1(n13404), .IN2(n13405), .QN(n13403) );
  NAND2X0 U13972 ( .IN1(n13406), .IN2(g1902), .QN(n13405) );
  NAND2X0 U13973 ( .IN1(n13407), .IN2(n13408), .QN(n13404) );
  NAND2X0 U13974 ( .IN1(g1906), .IN2(n8861), .QN(n13408) );
  INVX0 U13975 ( .INP(n13406), .ZN(n13407) );
  NAND3X0 U13976 ( .IN1(n13409), .IN2(g1917), .IN3(n5510), .QN(n13406) );
  NAND3X0 U13977 ( .IN1(n13410), .IN2(n13411), .IN3(n13412), .QN(g30357) );
  INVX0 U13978 ( .INP(n13413), .ZN(n13412) );
  NOR2X0 U13979 ( .IN1(n13414), .IN2(n5892), .QN(n13413) );
  INVX0 U13980 ( .INP(n13415), .ZN(n13411) );
  NOR2X0 U13981 ( .IN1(n13416), .IN2(n5785), .QN(n13415) );
  NOR2X0 U13982 ( .IN1(n13417), .IN2(n9392), .QN(n13416) );
  NOR2X0 U13983 ( .IN1(n13418), .IN2(n5464), .QN(n13417) );
  NAND3X0 U13984 ( .IN1(n13419), .IN2(n5464), .IN3(n5785), .QN(n13410) );
  NAND2X0 U13985 ( .IN1(n13420), .IN2(n13421), .QN(g30356) );
  INVX0 U13986 ( .INP(n13422), .ZN(n13421) );
  NOR2X0 U13987 ( .IN1(n13414), .IN2(n5785), .QN(n13422) );
  NAND2X0 U13988 ( .IN1(n13414), .IN2(g1848), .QN(n13420) );
  NAND3X0 U13989 ( .IN1(n13423), .IN2(n13424), .IN3(n13425), .QN(g30355) );
  NAND2X0 U13990 ( .IN1(n9441), .IN2(g1830), .QN(n13425) );
  NAND2X0 U13991 ( .IN1(n13426), .IN2(g1834), .QN(n13424) );
  INVX0 U13992 ( .INP(n13414), .ZN(n13426) );
  NAND2X0 U13993 ( .IN1(n13418), .IN2(n9376), .QN(n13414) );
  NAND2X0 U13994 ( .IN1(n13419), .IN2(n5665), .QN(n13423) );
  NAND3X0 U13995 ( .IN1(n13427), .IN2(n13428), .IN3(n13429), .QN(g30354) );
  NAND2X0 U13996 ( .IN1(n9441), .IN2(g1825), .QN(n13429) );
  NAND3X0 U13997 ( .IN1(n3628), .IN2(n13430), .IN3(n8854), .QN(n13428) );
  NAND2X0 U13998 ( .IN1(n13431), .IN2(n13432), .QN(n13430) );
  NAND2X0 U13999 ( .IN1(n8505), .IN2(g1821), .QN(n13432) );
  NAND2X0 U14000 ( .IN1(n8384), .IN2(g1825), .QN(n13431) );
  NAND2X0 U14001 ( .IN1(n13433), .IN2(g1830), .QN(n13427) );
  NAND2X0 U14002 ( .IN1(n12237), .IN2(n13434), .QN(n13433) );
  NAND2X0 U14003 ( .IN1(n9365), .IN2(n12249), .QN(n13434) );
  INVX0 U14004 ( .INP(n8854), .ZN(n12249) );
  NAND2X0 U14005 ( .IN1(n13435), .IN2(n13436), .QN(g30353) );
  NAND2X0 U14006 ( .IN1(n9441), .IN2(g1748), .QN(n13436) );
  NAND2X0 U14007 ( .IN1(n13437), .IN2(n9376), .QN(n13435) );
  NAND2X0 U14008 ( .IN1(n13438), .IN2(n13439), .QN(n13437) );
  NAND2X0 U14009 ( .IN1(n13440), .IN2(g1768), .QN(n13439) );
  NAND2X0 U14010 ( .IN1(n13441), .IN2(n13442), .QN(n13438) );
  NAND2X0 U14011 ( .IN1(n5352), .IN2(g1772), .QN(n13442) );
  INVX0 U14012 ( .INP(n13440), .ZN(n13441) );
  NAND3X0 U14013 ( .IN1(n13443), .IN2(g1783), .IN3(n5359), .QN(n13440) );
  NAND3X0 U14014 ( .IN1(n13444), .IN2(n13445), .IN3(n13446), .QN(g30352) );
  NAND2X0 U14015 ( .IN1(n13447), .IN2(n9236), .QN(n13446) );
  NAND2X0 U14016 ( .IN1(n13448), .IN2(g1720), .QN(n13445) );
  NAND2X0 U14017 ( .IN1(n13449), .IN2(n9376), .QN(n13448) );
  NAND2X0 U14018 ( .IN1(n13450), .IN2(g1714), .QN(n13449) );
  NAND4X0 U14019 ( .IN1(n5460), .IN2(n9355), .IN3(n13450), .IN4(n5780), .QN(
        n13444) );
  NAND2X0 U14020 ( .IN1(n13451), .IN2(n13452), .QN(g30351) );
  NAND2X0 U14021 ( .IN1(n13447), .IN2(g1720), .QN(n13452) );
  NAND2X0 U14022 ( .IN1(n13453), .IN2(g1714), .QN(n13451) );
  INVX0 U14023 ( .INP(n13447), .ZN(n13453) );
  NAND3X0 U14024 ( .IN1(n13454), .IN2(n13455), .IN3(n13456), .QN(g30350) );
  NAND2X0 U14025 ( .IN1(n13447), .IN2(g1700), .QN(n13456) );
  NOR2X0 U14026 ( .IN1(n13450), .IN2(n9393), .QN(n13447) );
  NAND3X0 U14027 ( .IN1(n13450), .IN2(n5417), .IN3(n9345), .QN(n13455) );
  NAND2X0 U14028 ( .IN1(n9440), .IN2(g1696), .QN(n13454) );
  NAND3X0 U14029 ( .IN1(n13457), .IN2(n13458), .IN3(n13459), .QN(g30349) );
  NAND2X0 U14030 ( .IN1(n9440), .IN2(g1691), .QN(n13459) );
  NAND3X0 U14031 ( .IN1(n3646), .IN2(n13460), .IN3(n8857), .QN(n13458) );
  NAND2X0 U14032 ( .IN1(n13461), .IN2(n13462), .QN(n13460) );
  NAND2X0 U14033 ( .IN1(n8509), .IN2(g1687), .QN(n13462) );
  NAND2X0 U14034 ( .IN1(n8388), .IN2(g1691), .QN(n13461) );
  NAND2X0 U14035 ( .IN1(n13463), .IN2(g1696), .QN(n13457) );
  NAND2X0 U14036 ( .IN1(n12258), .IN2(n13464), .QN(n13463) );
  NAND2X0 U14037 ( .IN1(n9366), .IN2(n12277), .QN(n13464) );
  INVX0 U14038 ( .INP(n8857), .ZN(n12277) );
  NAND3X0 U14039 ( .IN1(n13465), .IN2(n13466), .IN3(n13467), .QN(g30348) );
  NAND2X0 U14040 ( .IN1(n9440), .IN2(g1612), .QN(n13467) );
  NAND3X0 U14041 ( .IN1(g25167), .IN2(n11839), .IN3(n3646), .QN(n13466) );
  NAND2X0 U14042 ( .IN1(n5362), .IN2(g1636), .QN(n11839) );
  NAND2X0 U14043 ( .IN1(n13468), .IN2(g1632), .QN(n13465) );
  NAND2X0 U14044 ( .IN1(n12258), .IN2(n13469), .QN(n13468) );
  NAND2X0 U14045 ( .IN1(n10753), .IN2(n9376), .QN(n13469) );
  INVX0 U14046 ( .INP(g25167), .ZN(n10753) );
  NAND2X0 U14047 ( .IN1(n13470), .IN2(n13471), .QN(g30347) );
  NAND3X0 U14048 ( .IN1(n13472), .IN2(n13473), .IN3(n13474), .QN(n13471) );
  NAND2X0 U14049 ( .IN1(n13475), .IN2(n13476), .QN(n13472) );
  NAND2X0 U14050 ( .IN1(n9365), .IN2(g1413), .QN(n13475) );
  NAND2X0 U14051 ( .IN1(n9440), .IN2(g1542), .QN(n13470) );
  NAND2X0 U14052 ( .IN1(n13477), .IN2(n13478), .QN(g30346) );
  NAND2X0 U14053 ( .IN1(n9440), .IN2(g1536), .QN(n13478) );
  NAND4X0 U14054 ( .IN1(n13476), .IN2(n13479), .IN3(n13474), .IN4(n9361), .QN(
        n13477) );
  NAND2X0 U14055 ( .IN1(n8764), .IN2(n13480), .QN(n13479) );
  INVX0 U14056 ( .INP(n13481), .ZN(n13476) );
  NAND2X0 U14057 ( .IN1(n13482), .IN2(n13483), .QN(g30345) );
  NAND2X0 U14058 ( .IN1(n13484), .IN2(n9376), .QN(n13483) );
  NAND2X0 U14059 ( .IN1(n13474), .IN2(n11633), .QN(n13484) );
  INVX0 U14060 ( .INP(n13485), .ZN(n13474) );
  NAND2X0 U14061 ( .IN1(n13486), .IN2(g1514), .QN(n13482) );
  NAND2X0 U14062 ( .IN1(n13487), .IN2(n9376), .QN(n13486) );
  NAND2X0 U14063 ( .IN1(n13488), .IN2(n13489), .QN(n13487) );
  NAND2X0 U14064 ( .IN1(test_so49), .IN2(g7946), .QN(n13489) );
  NAND2X0 U14065 ( .IN1(n5302), .IN2(n8859), .QN(n13488) );
  NOR2X0 U14066 ( .IN1(n9413), .IN2(n13490), .QN(g30344) );
  NOR3X0 U14067 ( .IN1(n13485), .IN2(n13491), .IN3(n13492), .QN(n13490) );
  NOR2X0 U14068 ( .IN1(n5364), .IN2(g7946), .QN(n13492) );
  NOR2X0 U14069 ( .IN1(n5302), .IN2(g1514), .QN(n13491) );
  NAND2X0 U14070 ( .IN1(n13493), .IN2(n13494), .QN(n13485) );
  NAND2X0 U14071 ( .IN1(n4172), .IN2(n13495), .QN(n13494) );
  INVX0 U14072 ( .INP(n13496), .ZN(n4172) );
  NAND4X0 U14073 ( .IN1(n8588), .IN2(n4895), .IN3(n13497), .IN4(g7946), .QN(
        n13496) );
  NOR2X0 U14074 ( .IN1(n5577), .IN2(n5381), .QN(n13497) );
  NAND3X0 U14075 ( .IN1(n13498), .IN2(n13499), .IN3(n13500), .QN(g30343) );
  NAND2X0 U14076 ( .IN1(n4175), .IN2(n12281), .QN(n13500) );
  NAND2X0 U14077 ( .IN1(n9439), .IN2(g1345), .QN(n13499) );
  NAND3X0 U14078 ( .IN1(n12411), .IN2(g1361), .IN3(n9345), .QN(n13498) );
  NAND2X0 U14079 ( .IN1(n13501), .IN2(n13502), .QN(n12411) );
  NAND2X0 U14080 ( .IN1(n8448), .IN2(n11847), .QN(n13502) );
  INVX0 U14081 ( .INP(n13503), .ZN(n11847) );
  NAND3X0 U14082 ( .IN1(n13504), .IN2(n13505), .IN3(n13506), .QN(g30342) );
  NAND2X0 U14083 ( .IN1(n9439), .IN2(g1256), .QN(n13506) );
  NAND3X0 U14084 ( .IN1(n11853), .IN2(n13507), .IN3(g1259), .QN(n13505) );
  INVX0 U14085 ( .INP(n3736), .ZN(n13507) );
  NAND2X0 U14086 ( .IN1(n3736), .IN2(n5553), .QN(n13504) );
  NAND2X0 U14087 ( .IN1(n13508), .IN2(n13509), .QN(g30341) );
  NAND3X0 U14088 ( .IN1(n13510), .IN2(n13511), .IN3(n13512), .QN(n13509) );
  NAND2X0 U14089 ( .IN1(n13513), .IN2(n13514), .QN(n13510) );
  NAND2X0 U14090 ( .IN1(n9365), .IN2(g1070), .QN(n13513) );
  NAND2X0 U14091 ( .IN1(n9439), .IN2(g1199), .QN(n13508) );
  NAND2X0 U14092 ( .IN1(n13515), .IN2(n13516), .QN(g30340) );
  NAND2X0 U14093 ( .IN1(n9439), .IN2(g1193), .QN(n13516) );
  NAND4X0 U14094 ( .IN1(n13514), .IN2(n13517), .IN3(n13512), .IN4(n9361), .QN(
        n13515) );
  NAND2X0 U14095 ( .IN1(n8763), .IN2(n13518), .QN(n13517) );
  INVX0 U14096 ( .INP(n13519), .ZN(n13514) );
  NAND2X0 U14097 ( .IN1(n13520), .IN2(n13521), .QN(g30339) );
  NAND2X0 U14098 ( .IN1(n13522), .IN2(n9376), .QN(n13521) );
  NAND2X0 U14099 ( .IN1(n13512), .IN2(n11800), .QN(n13522) );
  INVX0 U14100 ( .INP(n13523), .ZN(n13512) );
  NAND2X0 U14101 ( .IN1(n13524), .IN2(g1171), .QN(n13520) );
  NAND3X0 U14102 ( .IN1(n13525), .IN2(n13526), .IN3(n9344), .QN(n13524) );
  NAND2X0 U14103 ( .IN1(n5599), .IN2(g7916), .QN(n13526) );
  NAND2X0 U14104 ( .IN1(n5304), .IN2(g1183), .QN(n13525) );
  NOR2X0 U14105 ( .IN1(n9415), .IN2(n13527), .QN(g30338) );
  NOR3X0 U14106 ( .IN1(n13523), .IN2(n13528), .IN3(n13529), .QN(n13527) );
  NOR2X0 U14107 ( .IN1(n5363), .IN2(g7916), .QN(n13529) );
  NOR2X0 U14108 ( .IN1(n5304), .IN2(g1171), .QN(n13528) );
  NAND2X0 U14109 ( .IN1(n13530), .IN2(n13531), .QN(n13523) );
  NAND2X0 U14110 ( .IN1(n4190), .IN2(n13532), .QN(n13531) );
  INVX0 U14111 ( .INP(n13533), .ZN(n4190) );
  NAND4X0 U14112 ( .IN1(n5642), .IN2(n4920), .IN3(n13534), .IN4(g1178), .QN(
        n13533) );
  NAND3X0 U14113 ( .IN1(n13535), .IN2(n13536), .IN3(n13537), .QN(g30337) );
  NAND2X0 U14114 ( .IN1(n4193), .IN2(n12294), .QN(n13537) );
  NAND2X0 U14115 ( .IN1(n9438), .IN2(g1002), .QN(n13536) );
  NAND3X0 U14116 ( .IN1(n12420), .IN2(g1018), .IN3(n9344), .QN(n13535) );
  NAND2X0 U14117 ( .IN1(n13538), .IN2(n13539), .QN(n12420) );
  NAND2X0 U14118 ( .IN1(n8449), .IN2(n11861), .QN(n13539) );
  NAND3X0 U14119 ( .IN1(n13540), .IN2(n13541), .IN3(n13542), .QN(g30336) );
  NAND2X0 U14120 ( .IN1(n9438), .IN2(g911), .QN(n13542) );
  NAND3X0 U14121 ( .IN1(n11867), .IN2(n13543), .IN3(g914), .QN(n13541) );
  INVX0 U14122 ( .INP(n3741), .ZN(n13543) );
  NAND2X0 U14123 ( .IN1(n3741), .IN2(n5560), .QN(n13540) );
  NAND3X0 U14124 ( .IN1(n13544), .IN2(n13545), .IN3(n13546), .QN(g30335) );
  NAND2X0 U14125 ( .IN1(test_so60), .IN2(n9516), .QN(n13546) );
  NAND3X0 U14126 ( .IN1(n2404), .IN2(n13547), .IN3(g744), .QN(n13545) );
  NAND2X0 U14127 ( .IN1(n57), .IN2(n5470), .QN(n13544) );
  INVX0 U14128 ( .INP(n13547), .ZN(n57) );
  NAND3X0 U14129 ( .IN1(n13548), .IN2(n513), .IN3(test_so60), .QN(n13547) );
  NAND2X0 U14130 ( .IN1(n8791), .IN2(g11678), .QN(n513) );
  NAND3X0 U14131 ( .IN1(n13549), .IN2(n13550), .IN3(n13551), .QN(g30334) );
  NAND2X0 U14132 ( .IN1(n9438), .IN2(g586), .QN(n13551) );
  NAND3X0 U14133 ( .IN1(n2421), .IN2(n13552), .IN3(g577), .QN(n13550) );
  INVX0 U14134 ( .INP(n3745), .ZN(n13552) );
  NAND2X0 U14135 ( .IN1(n3745), .IN2(n5294), .QN(n13549) );
  NAND2X0 U14136 ( .IN1(n13553), .IN2(n13554), .QN(g30333) );
  NAND2X0 U14137 ( .IN1(n10739), .IN2(n13555), .QN(n13554) );
  NAND2X0 U14138 ( .IN1(n13556), .IN2(n13557), .QN(n13555) );
  NAND2X0 U14139 ( .IN1(test_so73), .IN2(n12444), .QN(n13557) );
  NAND2X0 U14140 ( .IN1(n13558), .IN2(n8883), .QN(n13556) );
  NOR2X0 U14141 ( .IN1(n12443), .IN2(n9394), .QN(n10739) );
  NAND3X0 U14142 ( .IN1(n13559), .IN2(g691), .IN3(n13560), .QN(n12443) );
  NAND2X0 U14143 ( .IN1(n13558), .IN2(n13561), .QN(n13560) );
  NAND2X0 U14144 ( .IN1(n13562), .IN2(n8871), .QN(n13561) );
  INVX0 U14145 ( .INP(n12444), .ZN(n13558) );
  NAND2X0 U14146 ( .IN1(n9438), .IN2(g142), .QN(n13553) );
  NAND3X0 U14147 ( .IN1(n13563), .IN2(n13564), .IN3(n13565), .QN(g29309) );
  NAND2X0 U14148 ( .IN1(n3765), .IN2(n13566), .QN(n13565) );
  NAND2X0 U14149 ( .IN1(g6541), .IN2(n13567), .QN(n13566) );
  NAND3X0 U14150 ( .IN1(n13568), .IN2(g6541), .IN3(n12468), .QN(n13563) );
  NAND3X0 U14151 ( .IN1(n13569), .IN2(n13570), .IN3(n13571), .QN(g29308) );
  NAND2X0 U14152 ( .IN1(n9438), .IN2(g6523), .QN(n13571) );
  NAND2X0 U14153 ( .IN1(n13572), .IN2(g6527), .QN(n13570) );
  NAND2X0 U14154 ( .IN1(n5659), .IN2(n13573), .QN(n13569) );
  NAND3X0 U14155 ( .IN1(n13574), .IN2(n13575), .IN3(n13576), .QN(g29307) );
  NAND2X0 U14156 ( .IN1(n13572), .IN2(g6523), .QN(n13576) );
  NAND2X0 U14157 ( .IN1(n13577), .IN2(g6519), .QN(n13575) );
  NAND2X0 U14158 ( .IN1(n13578), .IN2(n9377), .QN(n13577) );
  NAND2X0 U14159 ( .IN1(n13579), .IN2(g6513), .QN(n13578) );
  NAND3X0 U14160 ( .IN1(n5426), .IN2(n13573), .IN3(n5806), .QN(n13574) );
  NAND2X0 U14161 ( .IN1(n13580), .IN2(n13581), .QN(g29306) );
  NAND2X0 U14162 ( .IN1(n13572), .IN2(g6519), .QN(n13581) );
  NAND2X0 U14163 ( .IN1(n13582), .IN2(g6513), .QN(n13580) );
  NAND3X0 U14164 ( .IN1(n13583), .IN2(n13584), .IN3(n13585), .QN(g29305) );
  NAND2X0 U14165 ( .IN1(n13572), .IN2(g6509), .QN(n13585) );
  INVX0 U14166 ( .INP(n13582), .ZN(n13572) );
  NAND2X0 U14167 ( .IN1(n13586), .IN2(n9377), .QN(n13582) );
  NAND2X0 U14168 ( .IN1(n13587), .IN2(g6500), .QN(n13584) );
  NAND2X0 U14169 ( .IN1(n13588), .IN2(n9377), .QN(n13587) );
  NAND2X0 U14170 ( .IN1(n8422), .IN2(n13579), .QN(n13588) );
  NAND3X0 U14171 ( .IN1(n13573), .IN2(g6505), .IN3(n5748), .QN(n13583) );
  NOR2X0 U14172 ( .IN1(n13586), .IN2(n9394), .QN(n13573) );
  INVX0 U14173 ( .INP(n13579), .ZN(n13586) );
  NOR2X0 U14174 ( .IN1(n13589), .IN2(n8850), .QN(n13579) );
  NAND3X0 U14175 ( .IN1(n13590), .IN2(n13591), .IN3(n13592), .QN(g29304) );
  NAND2X0 U14176 ( .IN1(n11388), .IN2(g6500), .QN(n13592) );
  NAND2X0 U14177 ( .IN1(n9437), .IN2(g6505), .QN(n13591) );
  NAND3X0 U14178 ( .IN1(n11381), .IN2(n13593), .IN3(n9344), .QN(n13590) );
  NAND2X0 U14179 ( .IN1(n13594), .IN2(n13595), .QN(n13593) );
  INVX0 U14180 ( .INP(n13596), .ZN(n13595) );
  NOR2X0 U14181 ( .IN1(n13597), .IN2(n13598), .QN(n13596) );
  NAND2X0 U14182 ( .IN1(n13598), .IN2(n13597), .QN(n13594) );
  NAND2X0 U14183 ( .IN1(g6500), .IN2(n13589), .QN(n13597) );
  NAND3X0 U14184 ( .IN1(g6727), .IN2(g17722), .IN3(n9684), .QN(n13589) );
  NAND3X0 U14185 ( .IN1(n13599), .IN2(n13564), .IN3(n13600), .QN(g29303) );
  NAND2X0 U14186 ( .IN1(n3765), .IN2(n13601), .QN(n13600) );
  NAND2X0 U14187 ( .IN1(g6195), .IN2(n11359), .QN(n13601) );
  INVX0 U14188 ( .INP(n12553), .ZN(n11359) );
  NAND3X0 U14189 ( .IN1(n13568), .IN2(g6195), .IN3(n12552), .QN(n13599) );
  NAND3X0 U14190 ( .IN1(n13602), .IN2(n13603), .IN3(n13604), .QN(g29302) );
  NAND2X0 U14191 ( .IN1(n9437), .IN2(g6177), .QN(n13604) );
  NAND2X0 U14192 ( .IN1(n13605), .IN2(g6181), .QN(n13603) );
  NAND2X0 U14193 ( .IN1(n5667), .IN2(n13606), .QN(n13602) );
  NAND3X0 U14194 ( .IN1(n13607), .IN2(n13608), .IN3(n13609), .QN(g29301) );
  NAND2X0 U14195 ( .IN1(n13605), .IN2(g6177), .QN(n13609) );
  NAND2X0 U14196 ( .IN1(n13610), .IN2(g6173), .QN(n13608) );
  NAND2X0 U14197 ( .IN1(n13611), .IN2(n9377), .QN(n13610) );
  NAND2X0 U14198 ( .IN1(n13612), .IN2(g6167), .QN(n13611) );
  NAND3X0 U14199 ( .IN1(n5430), .IN2(n13606), .IN3(n5810), .QN(n13607) );
  NAND2X0 U14200 ( .IN1(n13613), .IN2(n13614), .QN(g29300) );
  NAND2X0 U14201 ( .IN1(n13605), .IN2(g6173), .QN(n13614) );
  NAND2X0 U14202 ( .IN1(n13615), .IN2(g6167), .QN(n13613) );
  NAND3X0 U14203 ( .IN1(n13616), .IN2(n13617), .IN3(n13618), .QN(g29299) );
  NAND2X0 U14204 ( .IN1(n13605), .IN2(g6163), .QN(n13618) );
  INVX0 U14205 ( .INP(n13615), .ZN(n13605) );
  NAND2X0 U14206 ( .IN1(n13619), .IN2(n9377), .QN(n13615) );
  NAND2X0 U14207 ( .IN1(n13620), .IN2(g6154), .QN(n13617) );
  NAND2X0 U14208 ( .IN1(n13621), .IN2(n9377), .QN(n13620) );
  NAND2X0 U14209 ( .IN1(n8421), .IN2(n13612), .QN(n13621) );
  NAND3X0 U14210 ( .IN1(n13606), .IN2(g6159), .IN3(n5747), .QN(n13616) );
  NOR2X0 U14211 ( .IN1(n13619), .IN2(n9394), .QN(n13606) );
  INVX0 U14212 ( .INP(n13612), .ZN(n13619) );
  NOR2X0 U14213 ( .IN1(n13622), .IN2(n11399), .QN(n13612) );
  NAND3X0 U14214 ( .IN1(n13623), .IN2(n13624), .IN3(n13625), .QN(g29298) );
  NAND2X0 U14215 ( .IN1(n11404), .IN2(g6154), .QN(n13625) );
  NAND2X0 U14216 ( .IN1(n9437), .IN2(g6159), .QN(n13624) );
  NAND3X0 U14217 ( .IN1(n11393), .IN2(n13626), .IN3(n9344), .QN(n13623) );
  NAND2X0 U14218 ( .IN1(n13627), .IN2(n13628), .QN(n13626) );
  INVX0 U14219 ( .INP(n13629), .ZN(n13628) );
  NOR2X0 U14220 ( .IN1(n13630), .IN2(n13631), .QN(n13629) );
  NAND2X0 U14221 ( .IN1(n13631), .IN2(n13630), .QN(n13627) );
  NAND2X0 U14222 ( .IN1(g6154), .IN2(n13622), .QN(n13630) );
  NAND3X0 U14223 ( .IN1(n10581), .IN2(g17685), .IN3(test_so69), .QN(n13622) );
  NAND3X0 U14224 ( .IN1(n13632), .IN2(n13564), .IN3(n13633), .QN(g29297) );
  NAND2X0 U14225 ( .IN1(n3765), .IN2(n13634), .QN(n13633) );
  NAND2X0 U14226 ( .IN1(g5849), .IN2(n11358), .QN(n13634) );
  INVX0 U14227 ( .INP(n12639), .ZN(n11358) );
  NAND3X0 U14228 ( .IN1(n13568), .IN2(g5849), .IN3(n12638), .QN(n13632) );
  NAND3X0 U14229 ( .IN1(n13635), .IN2(n13636), .IN3(n13637), .QN(g29296) );
  NAND2X0 U14230 ( .IN1(n9437), .IN2(g5831), .QN(n13637) );
  NAND2X0 U14231 ( .IN1(n13638), .IN2(g5835), .QN(n13636) );
  NAND2X0 U14232 ( .IN1(n5663), .IN2(n13639), .QN(n13635) );
  NAND3X0 U14233 ( .IN1(n13640), .IN2(n13641), .IN3(n13642), .QN(g29295) );
  NAND2X0 U14234 ( .IN1(n13638), .IN2(g5831), .QN(n13642) );
  NAND2X0 U14235 ( .IN1(n13643), .IN2(g5827), .QN(n13641) );
  NAND2X0 U14236 ( .IN1(n13644), .IN2(n9377), .QN(n13643) );
  NAND2X0 U14237 ( .IN1(n13645), .IN2(g5821), .QN(n13644) );
  NAND3X0 U14238 ( .IN1(n5429), .IN2(n13639), .IN3(n5809), .QN(n13640) );
  NAND2X0 U14239 ( .IN1(n13646), .IN2(n13647), .QN(g29294) );
  NAND2X0 U14240 ( .IN1(n13638), .IN2(g5827), .QN(n13647) );
  NAND2X0 U14241 ( .IN1(n13648), .IN2(g5821), .QN(n13646) );
  NAND3X0 U14242 ( .IN1(n13649), .IN2(n13650), .IN3(n13651), .QN(g29293) );
  NAND2X0 U14243 ( .IN1(n13638), .IN2(g5817), .QN(n13651) );
  INVX0 U14244 ( .INP(n13648), .ZN(n13638) );
  NAND2X0 U14245 ( .IN1(n13652), .IN2(n9377), .QN(n13648) );
  NAND2X0 U14246 ( .IN1(n13653), .IN2(g5808), .QN(n13650) );
  NAND2X0 U14247 ( .IN1(n13654), .IN2(n9377), .QN(n13653) );
  NAND2X0 U14248 ( .IN1(n13645), .IN2(Tj_TriggerIN7), .QN(n13654) );
  NAND3X0 U14249 ( .IN1(g5813), .IN2(n13639), .IN3(n5749), .QN(n13649) );
  NOR2X0 U14250 ( .IN1(n13652), .IN2(n9388), .QN(n13639) );
  INVX0 U14251 ( .INP(n13645), .ZN(n13652) );
  NOR2X0 U14252 ( .IN1(n13655), .IN2(n11415), .QN(n13645) );
  NAND3X0 U14253 ( .IN1(n13656), .IN2(n13657), .IN3(n13658), .QN(g29292) );
  NAND2X0 U14254 ( .IN1(n11420), .IN2(g5808), .QN(n13658) );
  NAND2X0 U14255 ( .IN1(g5813), .IN2(n9516), .QN(n13657) );
  NAND3X0 U14256 ( .IN1(n11409), .IN2(n13659), .IN3(n9343), .QN(n13656) );
  NAND2X0 U14257 ( .IN1(n13660), .IN2(n13661), .QN(n13659) );
  INVX0 U14258 ( .INP(n13662), .ZN(n13661) );
  NOR2X0 U14259 ( .IN1(n13663), .IN2(n13664), .QN(n13662) );
  NAND2X0 U14260 ( .IN1(n13664), .IN2(n13663), .QN(n13660) );
  NAND2X0 U14261 ( .IN1(g5808), .IN2(n13655), .QN(n13663) );
  NAND3X0 U14262 ( .IN1(g6035), .IN2(g17646), .IN3(n10586), .QN(n13655) );
  NAND3X0 U14263 ( .IN1(n13665), .IN2(n13564), .IN3(n13666), .QN(g29291) );
  NAND2X0 U14264 ( .IN1(n3765), .IN2(n13667), .QN(n13666) );
  NAND2X0 U14265 ( .IN1(g5503), .IN2(n13668), .QN(n13667) );
  NAND3X0 U14266 ( .IN1(n13568), .IN2(g5503), .IN3(n12724), .QN(n13665) );
  NAND3X0 U14267 ( .IN1(n13669), .IN2(n13670), .IN3(n13671), .QN(g29290) );
  NAND2X0 U14268 ( .IN1(n9436), .IN2(g5485), .QN(n13671) );
  NAND2X0 U14269 ( .IN1(n13672), .IN2(g5489), .QN(n13670) );
  NAND2X0 U14270 ( .IN1(n5660), .IN2(n13673), .QN(n13669) );
  NAND3X0 U14271 ( .IN1(n13674), .IN2(n13675), .IN3(n13676), .QN(g29289) );
  NAND2X0 U14272 ( .IN1(n13672), .IN2(g5485), .QN(n13676) );
  NAND2X0 U14273 ( .IN1(n13677), .IN2(g5481), .QN(n13675) );
  NAND2X0 U14274 ( .IN1(n13678), .IN2(n9377), .QN(n13677) );
  NAND2X0 U14275 ( .IN1(n13679), .IN2(g5475), .QN(n13678) );
  NAND3X0 U14276 ( .IN1(n5425), .IN2(n13673), .IN3(n5805), .QN(n13674) );
  NAND2X0 U14277 ( .IN1(n13680), .IN2(n13681), .QN(g29288) );
  NAND2X0 U14278 ( .IN1(n13672), .IN2(g5481), .QN(n13681) );
  NAND2X0 U14279 ( .IN1(n13682), .IN2(g5475), .QN(n13680) );
  NAND3X0 U14280 ( .IN1(n13683), .IN2(n13684), .IN3(n13685), .QN(g29287) );
  NAND2X0 U14281 ( .IN1(n13672), .IN2(g5471), .QN(n13685) );
  INVX0 U14282 ( .INP(n13682), .ZN(n13672) );
  NAND2X0 U14283 ( .IN1(n13686), .IN2(n9377), .QN(n13682) );
  NAND2X0 U14284 ( .IN1(n13687), .IN2(g5462), .QN(n13684) );
  NAND2X0 U14285 ( .IN1(n13688), .IN2(n9377), .QN(n13687) );
  NAND2X0 U14286 ( .IN1(n8408), .IN2(n13679), .QN(n13688) );
  NAND3X0 U14287 ( .IN1(n13673), .IN2(g5467), .IN3(n5744), .QN(n13683) );
  NOR2X0 U14288 ( .IN1(n13686), .IN2(n9421), .QN(n13673) );
  INVX0 U14289 ( .INP(n13679), .ZN(n13686) );
  NOR2X0 U14290 ( .IN1(n13689), .IN2(n11431), .QN(n13679) );
  NAND3X0 U14291 ( .IN1(n13690), .IN2(n13691), .IN3(n13692), .QN(g29286) );
  NAND2X0 U14292 ( .IN1(n11436), .IN2(g5462), .QN(n13692) );
  NAND2X0 U14293 ( .IN1(n9436), .IN2(g5467), .QN(n13691) );
  NAND3X0 U14294 ( .IN1(n11425), .IN2(n13693), .IN3(n9334), .QN(n13690) );
  NAND2X0 U14295 ( .IN1(n13694), .IN2(n13695), .QN(n13693) );
  INVX0 U14296 ( .INP(n13696), .ZN(n13695) );
  NOR2X0 U14297 ( .IN1(n13697), .IN2(n13698), .QN(n13696) );
  NAND2X0 U14298 ( .IN1(n13698), .IN2(n13697), .QN(n13694) );
  NAND2X0 U14299 ( .IN1(g5462), .IN2(n13689), .QN(n13697) );
  NAND3X0 U14300 ( .IN1(g5689), .IN2(g17604), .IN3(n10594), .QN(n13689) );
  NAND3X0 U14301 ( .IN1(n13699), .IN2(n13564), .IN3(n13700), .QN(g29285) );
  NAND2X0 U14302 ( .IN1(n3765), .IN2(n13701), .QN(n13700) );
  NAND2X0 U14303 ( .IN1(g5156), .IN2(n13702), .QN(n13701) );
  NAND3X0 U14304 ( .IN1(n13568), .IN2(g5156), .IN3(n12808), .QN(n13699) );
  NAND3X0 U14305 ( .IN1(n13703), .IN2(n13704), .IN3(n13705), .QN(g29284) );
  NAND2X0 U14306 ( .IN1(n9436), .IN2(g5138), .QN(n13705) );
  NAND2X0 U14307 ( .IN1(n13706), .IN2(g5142), .QN(n13704) );
  NAND2X0 U14308 ( .IN1(n5658), .IN2(n13707), .QN(n13703) );
  NAND3X0 U14309 ( .IN1(n13708), .IN2(n13709), .IN3(n13710), .QN(g29283) );
  NAND2X0 U14310 ( .IN1(n13706), .IN2(g5138), .QN(n13710) );
  NAND2X0 U14311 ( .IN1(n13711), .IN2(g5134), .QN(n13709) );
  NAND2X0 U14312 ( .IN1(n13712), .IN2(n9377), .QN(n13711) );
  NAND2X0 U14313 ( .IN1(test_so96), .IN2(n13713), .QN(n13712) );
  NAND3X0 U14314 ( .IN1(n13707), .IN2(n8877), .IN3(n5807), .QN(n13708) );
  NAND2X0 U14315 ( .IN1(n13714), .IN2(n13715), .QN(g29282) );
  NAND2X0 U14316 ( .IN1(n13706), .IN2(g5134), .QN(n13715) );
  NAND2X0 U14317 ( .IN1(test_so96), .IN2(n13716), .QN(n13714) );
  NAND3X0 U14318 ( .IN1(n13717), .IN2(n13718), .IN3(n13719), .QN(g29281) );
  NAND2X0 U14319 ( .IN1(n13706), .IN2(g5124), .QN(n13719) );
  INVX0 U14320 ( .INP(n13716), .ZN(n13706) );
  NAND2X0 U14321 ( .IN1(n13720), .IN2(n9378), .QN(n13716) );
  NAND2X0 U14322 ( .IN1(n13721), .IN2(g5115), .QN(n13718) );
  NAND2X0 U14323 ( .IN1(n13722), .IN2(n9378), .QN(n13721) );
  NAND2X0 U14324 ( .IN1(n8407), .IN2(n13713), .QN(n13722) );
  NAND3X0 U14325 ( .IN1(n13707), .IN2(g5120), .IN3(n5743), .QN(n13717) );
  NOR2X0 U14326 ( .IN1(n13720), .IN2(n9400), .QN(n13707) );
  INVX0 U14327 ( .INP(n13713), .ZN(n13720) );
  NOR2X0 U14328 ( .IN1(n13723), .IN2(n8845), .QN(n13713) );
  NAND3X0 U14329 ( .IN1(n13724), .IN2(n13725), .IN3(n13726), .QN(g29280) );
  NAND2X0 U14330 ( .IN1(n11448), .IN2(g5115), .QN(n13726) );
  NAND2X0 U14331 ( .IN1(n9436), .IN2(g5120), .QN(n13725) );
  NAND3X0 U14332 ( .IN1(g33959), .IN2(n13727), .IN3(n9343), .QN(n13724) );
  NAND2X0 U14333 ( .IN1(n13728), .IN2(n13729), .QN(n13727) );
  INVX0 U14334 ( .INP(n13730), .ZN(n13729) );
  NOR2X0 U14335 ( .IN1(n13731), .IN2(n13732), .QN(n13730) );
  NAND2X0 U14336 ( .IN1(n13732), .IN2(n13731), .QN(n13728) );
  NAND2X0 U14337 ( .IN1(g5115), .IN2(n13723), .QN(n13731) );
  NAND3X0 U14338 ( .IN1(g31860), .IN2(g17577), .IN3(test_so10), .QN(n13723) );
  NAND3X0 U14339 ( .IN1(n13733), .IN2(n13734), .IN3(n13735), .QN(g29275) );
  NAND2X0 U14340 ( .IN1(test_so11), .IN2(n9515), .QN(n13735) );
  NAND3X0 U14341 ( .IN1(n12912), .IN2(n12400), .IN3(g4087), .QN(n13734) );
  NAND3X0 U14342 ( .IN1(n12911), .IN2(g4169), .IN3(n5480), .QN(n13733) );
  INVX0 U14343 ( .INP(n12400), .ZN(n12911) );
  NAND2X0 U14344 ( .IN1(test_so11), .IN2(n13736), .QN(n12400) );
  NAND3X0 U14345 ( .IN1(n13737), .IN2(n13564), .IN3(n13738), .QN(g29274) );
  NAND2X0 U14346 ( .IN1(n3765), .IN2(n13739), .QN(n13738) );
  NAND2X0 U14347 ( .IN1(g3849), .IN2(n11369), .QN(n13739) );
  INVX0 U14348 ( .INP(n12917), .ZN(n11369) );
  NAND3X0 U14349 ( .IN1(n13568), .IN2(g3849), .IN3(n12916), .QN(n13737) );
  NAND3X0 U14350 ( .IN1(n13740), .IN2(n13741), .IN3(n13742), .QN(g29273) );
  NAND2X0 U14351 ( .IN1(n9435), .IN2(g3831), .QN(n13742) );
  NAND2X0 U14352 ( .IN1(n13743), .IN2(g3835), .QN(n13741) );
  NAND2X0 U14353 ( .IN1(n5662), .IN2(n13744), .QN(n13740) );
  NAND3X0 U14354 ( .IN1(n13745), .IN2(n13746), .IN3(n13747), .QN(g29272) );
  NAND2X0 U14355 ( .IN1(n13743), .IN2(g3831), .QN(n13747) );
  NAND2X0 U14356 ( .IN1(n13748), .IN2(g3827), .QN(n13746) );
  NAND2X0 U14357 ( .IN1(n13749), .IN2(n9378), .QN(n13748) );
  NAND2X0 U14358 ( .IN1(n13750), .IN2(g3821), .QN(n13749) );
  NAND3X0 U14359 ( .IN1(n5428), .IN2(n13744), .IN3(n5808), .QN(n13745) );
  NAND2X0 U14360 ( .IN1(n13751), .IN2(n13752), .QN(g29271) );
  NAND2X0 U14361 ( .IN1(n13743), .IN2(g3827), .QN(n13752) );
  INVX0 U14362 ( .INP(n13753), .ZN(n13743) );
  NAND2X0 U14363 ( .IN1(n13753), .IN2(g3821), .QN(n13751) );
  NAND2X0 U14364 ( .IN1(n13754), .IN2(n9378), .QN(n13753) );
  NAND3X0 U14365 ( .IN1(n13755), .IN2(n13756), .IN3(n13757), .QN(g29270) );
  NAND2X0 U14366 ( .IN1(n12464), .IN2(n13754), .QN(n13757) );
  INVX0 U14367 ( .INP(n10229), .ZN(n12464) );
  NAND2X0 U14368 ( .IN1(n9364), .IN2(g3817), .QN(n10229) );
  NAND2X0 U14369 ( .IN1(n13758), .IN2(g3808), .QN(n13756) );
  NAND2X0 U14370 ( .IN1(n13759), .IN2(n9378), .QN(n13758) );
  NAND2X0 U14371 ( .IN1(n8409), .IN2(n13750), .QN(n13759) );
  NAND3X0 U14372 ( .IN1(n13744), .IN2(g3813), .IN3(n5745), .QN(n13755) );
  NOR2X0 U14373 ( .IN1(n13754), .IN2(n9396), .QN(n13744) );
  INVX0 U14374 ( .INP(n13750), .ZN(n13754) );
  NOR2X0 U14375 ( .IN1(n13760), .IN2(n11471), .QN(n13750) );
  NAND3X0 U14376 ( .IN1(n13761), .IN2(n13762), .IN3(n13763), .QN(g29269) );
  NAND2X0 U14377 ( .IN1(n11476), .IN2(g3808), .QN(n13763) );
  NAND2X0 U14378 ( .IN1(n9434), .IN2(g3813), .QN(n13762) );
  NAND3X0 U14379 ( .IN1(n11465), .IN2(n13764), .IN3(n9342), .QN(n13761) );
  NAND2X0 U14380 ( .IN1(n13765), .IN2(n13766), .QN(n13764) );
  INVX0 U14381 ( .INP(n13767), .ZN(n13766) );
  NOR2X0 U14382 ( .IN1(n13768), .IN2(n13769), .QN(n13767) );
  NAND2X0 U14383 ( .IN1(n13769), .IN2(n13768), .QN(n13765) );
  NAND2X0 U14384 ( .IN1(g3808), .IN2(n13760), .QN(n13768) );
  NAND3X0 U14385 ( .IN1(g4040), .IN2(g16693), .IN3(n10582), .QN(n13760) );
  NAND3X0 U14386 ( .IN1(n13770), .IN2(n13564), .IN3(n13771), .QN(g29268) );
  NAND2X0 U14387 ( .IN1(n3765), .IN2(n13772), .QN(n13771) );
  NAND2X0 U14388 ( .IN1(g3498), .IN2(n11368), .QN(n13772) );
  INVX0 U14389 ( .INP(n13003), .ZN(n11368) );
  NAND3X0 U14390 ( .IN1(n13568), .IN2(g3498), .IN3(n13002), .QN(n13770) );
  NAND3X0 U14391 ( .IN1(n13773), .IN2(n13774), .IN3(n13775), .QN(g29267) );
  NAND2X0 U14392 ( .IN1(n9434), .IN2(g3480), .QN(n13775) );
  NAND2X0 U14393 ( .IN1(n13776), .IN2(g3484), .QN(n13774) );
  NAND2X0 U14394 ( .IN1(n5668), .IN2(n13777), .QN(n13773) );
  NAND3X0 U14395 ( .IN1(n13778), .IN2(n13779), .IN3(n13780), .QN(g29266) );
  NAND2X0 U14396 ( .IN1(n13776), .IN2(g3480), .QN(n13780) );
  NAND2X0 U14397 ( .IN1(n13781), .IN2(g3476), .QN(n13779) );
  NAND2X0 U14398 ( .IN1(n13782), .IN2(n9378), .QN(n13781) );
  NAND2X0 U14399 ( .IN1(n13783), .IN2(g3470), .QN(n13782) );
  NAND3X0 U14400 ( .IN1(n5424), .IN2(n13777), .IN3(n5786), .QN(n13778) );
  NAND2X0 U14401 ( .IN1(n13784), .IN2(n13785), .QN(g29265) );
  NAND2X0 U14402 ( .IN1(n13776), .IN2(g3476), .QN(n13785) );
  NAND2X0 U14403 ( .IN1(n13786), .IN2(g3470), .QN(n13784) );
  NAND3X0 U14404 ( .IN1(n13787), .IN2(n13788), .IN3(n13789), .QN(g29264) );
  NAND2X0 U14405 ( .IN1(n13776), .IN2(g3466), .QN(n13789) );
  INVX0 U14406 ( .INP(n13786), .ZN(n13776) );
  NAND2X0 U14407 ( .IN1(n13790), .IN2(n9378), .QN(n13786) );
  NAND2X0 U14408 ( .IN1(test_so4), .IN2(n13791), .QN(n13788) );
  NAND2X0 U14409 ( .IN1(n13792), .IN2(n9378), .QN(n13791) );
  NAND2X0 U14410 ( .IN1(n8410), .IN2(n13783), .QN(n13792) );
  NAND3X0 U14411 ( .IN1(n13777), .IN2(g3462), .IN3(n8891), .QN(n13787) );
  NOR2X0 U14412 ( .IN1(n13790), .IN2(n9397), .QN(n13777) );
  INVX0 U14413 ( .INP(n13783), .ZN(n13790) );
  NOR2X0 U14414 ( .IN1(n13793), .IN2(n11487), .QN(n13783) );
  NAND3X0 U14415 ( .IN1(n13794), .IN2(n13795), .IN3(n13796), .QN(g29263) );
  NAND2X0 U14416 ( .IN1(test_so4), .IN2(n11492), .QN(n13796) );
  NAND2X0 U14417 ( .IN1(n9433), .IN2(g3462), .QN(n13795) );
  NAND3X0 U14418 ( .IN1(n11481), .IN2(n13797), .IN3(n9342), .QN(n13794) );
  NAND2X0 U14419 ( .IN1(n13798), .IN2(n13799), .QN(n13797) );
  INVX0 U14420 ( .INP(n13800), .ZN(n13799) );
  NOR2X0 U14421 ( .IN1(n13801), .IN2(n13802), .QN(n13800) );
  NAND2X0 U14422 ( .IN1(n13802), .IN2(n13801), .QN(n13798) );
  NAND2X0 U14423 ( .IN1(test_so4), .IN2(n13793), .QN(n13801) );
  NAND3X0 U14424 ( .IN1(g3689), .IN2(g16656), .IN3(n10587), .QN(n13793) );
  NAND3X0 U14425 ( .IN1(n13803), .IN2(n13564), .IN3(n13804), .QN(g29262) );
  NAND2X0 U14426 ( .IN1(n3765), .IN2(n13805), .QN(n13804) );
  NAND2X0 U14427 ( .IN1(g3147), .IN2(n13806), .QN(n13805) );
  NAND2X0 U14428 ( .IN1(n3765), .IN2(n13568), .QN(n13564) );
  NAND3X0 U14429 ( .IN1(n13568), .IN2(g3147), .IN3(n13088), .QN(n13803) );
  INVX0 U14430 ( .INP(n4210), .ZN(n13568) );
  NAND2X0 U14431 ( .IN1(n8788), .IN2(g4180), .QN(n4210) );
  NAND3X0 U14432 ( .IN1(n13807), .IN2(n13808), .IN3(n13809), .QN(g29261) );
  NAND2X0 U14433 ( .IN1(n9433), .IN2(g3129), .QN(n13809) );
  NAND2X0 U14434 ( .IN1(n13810), .IN2(g3133), .QN(n13808) );
  NAND2X0 U14435 ( .IN1(n5661), .IN2(n13811), .QN(n13807) );
  NAND3X0 U14436 ( .IN1(n13812), .IN2(n13813), .IN3(n13814), .QN(g29260) );
  NAND2X0 U14437 ( .IN1(n13810), .IN2(g3129), .QN(n13814) );
  NAND2X0 U14438 ( .IN1(n13815), .IN2(g3125), .QN(n13813) );
  NAND2X0 U14439 ( .IN1(n13816), .IN2(n9378), .QN(n13815) );
  NAND2X0 U14440 ( .IN1(n13817), .IN2(g3119), .QN(n13816) );
  NAND3X0 U14441 ( .IN1(n5423), .IN2(n13811), .IN3(n5781), .QN(n13812) );
  NAND2X0 U14442 ( .IN1(n13818), .IN2(n13819), .QN(g29259) );
  NAND2X0 U14443 ( .IN1(n13810), .IN2(g3125), .QN(n13819) );
  NAND2X0 U14444 ( .IN1(n13820), .IN2(g3119), .QN(n13818) );
  NAND3X0 U14445 ( .IN1(n13821), .IN2(n13822), .IN3(n13823), .QN(g29258) );
  NAND2X0 U14446 ( .IN1(n13810), .IN2(g3115), .QN(n13823) );
  INVX0 U14447 ( .INP(n13820), .ZN(n13810) );
  NAND2X0 U14448 ( .IN1(n13824), .IN2(n9378), .QN(n13820) );
  NAND2X0 U14449 ( .IN1(n13825), .IN2(g3106), .QN(n13822) );
  NAND2X0 U14450 ( .IN1(n13826), .IN2(n9378), .QN(n13825) );
  NAND2X0 U14451 ( .IN1(n8406), .IN2(n13817), .QN(n13826) );
  NAND3X0 U14452 ( .IN1(n13811), .IN2(g3111), .IN3(n5742), .QN(n13821) );
  NOR2X0 U14453 ( .IN1(n13824), .IN2(n9398), .QN(n13811) );
  INVX0 U14454 ( .INP(n13817), .ZN(n13824) );
  NOR2X0 U14455 ( .IN1(n13827), .IN2(n11498), .QN(n13817) );
  NAND3X0 U14456 ( .IN1(n13828), .IN2(n13829), .IN3(n13830), .QN(g29257) );
  NAND2X0 U14457 ( .IN1(n11507), .IN2(g3106), .QN(n13830) );
  NAND2X0 U14458 ( .IN1(n9433), .IN2(g3111), .QN(n13829) );
  NAND3X0 U14459 ( .IN1(n11501), .IN2(n13831), .IN3(n9342), .QN(n13828) );
  NAND2X0 U14460 ( .IN1(n13832), .IN2(n13833), .QN(n13831) );
  INVX0 U14461 ( .INP(n13834), .ZN(n13833) );
  NOR2X0 U14462 ( .IN1(n13835), .IN2(n13836), .QN(n13834) );
  NAND2X0 U14463 ( .IN1(n13836), .IN2(n13835), .QN(n13832) );
  NAND2X0 U14464 ( .IN1(g3106), .IN2(n13827), .QN(n13835) );
  NAND3X0 U14465 ( .IN1(g3338), .IN2(g16624), .IN3(n10595), .QN(n13827) );
  NAND4X0 U14466 ( .IN1(n13837), .IN2(n9664), .IN3(n13838), .IN4(n13839), .QN(
        g29256) );
  NAND3X0 U14467 ( .IN1(n13214), .IN2(g2735), .IN3(n9342), .QN(n13839) );
  NAND2X0 U14468 ( .IN1(n9432), .IN2(g2729), .QN(n13838) );
  NAND2X0 U14469 ( .IN1(n5600), .IN2(n13840), .QN(n13837) );
  NAND2X0 U14470 ( .IN1(n13841), .IN2(n13842), .QN(g29255) );
  NAND2X0 U14471 ( .IN1(n13843), .IN2(g2652), .QN(n13842) );
  NAND2X0 U14472 ( .IN1(n12111), .IN2(n13844), .QN(n13843) );
  NAND2X0 U14473 ( .IN1(n4379), .IN2(n9378), .QN(n13844) );
  INVX0 U14474 ( .INP(n12117), .ZN(n12111) );
  NAND2X0 U14475 ( .IN1(n13845), .IN2(g2638), .QN(n13841) );
  NAND2X0 U14476 ( .IN1(n13846), .IN2(n9378), .QN(n13845) );
  INVX0 U14477 ( .INP(n13847), .ZN(n13846) );
  NOR2X0 U14478 ( .IN1(n12108), .IN2(n9698), .QN(n13847) );
  NOR2X0 U14479 ( .IN1(n8513), .IN2(n8849), .QN(n9698) );
  NAND4X0 U14480 ( .IN1(n13848), .IN2(n13849), .IN3(n13850), .IN4(n13851), 
        .QN(g29254) );
  NAND2X0 U14481 ( .IN1(n13224), .IN2(g2567), .QN(n13851) );
  NOR2X0 U14482 ( .IN1(n13223), .IN2(n9405), .QN(n13224) );
  NAND3X0 U14483 ( .IN1(g2587), .IN2(g2619), .IN3(n13248), .QN(n13223) );
  NAND2X0 U14484 ( .IN1(n3517), .IN2(n13852), .QN(n13850) );
  NAND3X0 U14485 ( .IN1(n13853), .IN2(n13854), .IN3(n13855), .QN(n13852) );
  NAND2X0 U14486 ( .IN1(n8849), .IN2(g2563), .QN(n13855) );
  NOR2X0 U14487 ( .IN1(g2587), .IN2(n8759), .QN(n8849) );
  NAND2X0 U14488 ( .IN1(n5508), .IN2(n13856), .QN(n13854) );
  NAND2X0 U14489 ( .IN1(n13857), .IN2(n13858), .QN(n13856) );
  NAND2X0 U14490 ( .IN1(test_so66), .IN2(n5372), .QN(n13858) );
  NAND2X0 U14491 ( .IN1(g2583), .IN2(g2610), .QN(n13857) );
  NAND2X0 U14492 ( .IN1(n8759), .IN2(n13859), .QN(n13853) );
  NAND2X0 U14493 ( .IN1(n13860), .IN2(n13861), .QN(n13859) );
  NAND2X0 U14494 ( .IN1(test_so61), .IN2(g2587), .QN(n13861) );
  NAND2X0 U14495 ( .IN1(g2619), .IN2(g2571), .QN(n13860) );
  NOR2X0 U14496 ( .IN1(n12108), .IN2(n9405), .QN(n3517) );
  NAND2X0 U14497 ( .IN1(n12117), .IN2(g2638), .QN(n13849) );
  NOR2X0 U14498 ( .IN1(n13248), .IN2(n9406), .QN(n12117) );
  INVX0 U14499 ( .INP(n12108), .ZN(n13248) );
  NAND3X0 U14500 ( .IN1(n13862), .IN2(n13863), .IN3(n13185), .QN(n12108) );
  NAND2X0 U14501 ( .IN1(n13205), .IN2(g2819), .QN(n13862) );
  NAND2X0 U14502 ( .IN1(n9431), .IN2(g2619), .QN(n13848) );
  NAND2X0 U14503 ( .IN1(n13864), .IN2(n13865), .QN(g29253) );
  NAND2X0 U14504 ( .IN1(n13866), .IN2(g2518), .QN(n13865) );
  NAND2X0 U14505 ( .IN1(n12132), .IN2(n13867), .QN(n13866) );
  NAND2X0 U14506 ( .IN1(n4391), .IN2(n9378), .QN(n13867) );
  INVX0 U14507 ( .INP(n12138), .ZN(n12132) );
  NAND2X0 U14508 ( .IN1(n13868), .IN2(g2504), .QN(n13864) );
  NAND2X0 U14509 ( .IN1(n13869), .IN2(n9378), .QN(n13868) );
  INVX0 U14510 ( .INP(n13870), .ZN(n13869) );
  NOR2X0 U14511 ( .IN1(n12129), .IN2(n9697), .QN(n13870) );
  NOR2X0 U14512 ( .IN1(n8512), .IN2(n8855), .QN(n9697) );
  NAND4X0 U14513 ( .IN1(n13871), .IN2(n13872), .IN3(n13873), .IN4(n13874), 
        .QN(g29252) );
  NAND2X0 U14514 ( .IN1(n13257), .IN2(g2433), .QN(n13874) );
  NOR2X0 U14515 ( .IN1(n13256), .IN2(n9405), .QN(n13257) );
  NAND3X0 U14516 ( .IN1(g2453), .IN2(g2485), .IN3(n13280), .QN(n13256) );
  NAND2X0 U14517 ( .IN1(n3536), .IN2(n13875), .QN(n13873) );
  NAND3X0 U14518 ( .IN1(n13876), .IN2(n13877), .IN3(n13878), .QN(n13875) );
  NAND2X0 U14519 ( .IN1(n8855), .IN2(g2429), .QN(n13878) );
  NOR2X0 U14520 ( .IN1(g2453), .IN2(n8758), .QN(n8855) );
  NAND2X0 U14521 ( .IN1(n5509), .IN2(n13879), .QN(n13877) );
  NAND2X0 U14522 ( .IN1(n13880), .IN2(n13881), .QN(n13879) );
  NAND2X0 U14523 ( .IN1(n5373), .IN2(g2441), .QN(n13881) );
  NAND2X0 U14524 ( .IN1(g2449), .IN2(g2476), .QN(n13880) );
  NAND2X0 U14525 ( .IN1(n8758), .IN2(n13882), .QN(n13876) );
  NAND2X0 U14526 ( .IN1(n13883), .IN2(n13884), .QN(n13882) );
  NAND2X0 U14527 ( .IN1(g2453), .IN2(n9274), .QN(n13884) );
  NAND2X0 U14528 ( .IN1(g2485), .IN2(g2437), .QN(n13883) );
  NOR2X0 U14529 ( .IN1(n12129), .IN2(n9404), .QN(n3536) );
  NAND2X0 U14530 ( .IN1(n12138), .IN2(g2504), .QN(n13872) );
  NOR2X0 U14531 ( .IN1(n13280), .IN2(n9403), .QN(n12138) );
  INVX0 U14532 ( .INP(n12129), .ZN(n13280) );
  NAND3X0 U14533 ( .IN1(n13885), .IN2(n13863), .IN3(n13186), .QN(n12129) );
  NAND2X0 U14534 ( .IN1(n13205), .IN2(g2815), .QN(n13885) );
  NAND2X0 U14535 ( .IN1(n9431), .IN2(g2485), .QN(n13871) );
  NAND2X0 U14536 ( .IN1(n13886), .IN2(n13887), .QN(g29251) );
  NAND2X0 U14537 ( .IN1(n13888), .IN2(g2384), .QN(n13887) );
  NAND2X0 U14538 ( .IN1(n12153), .IN2(n13889), .QN(n13888) );
  NAND2X0 U14539 ( .IN1(n4402), .IN2(n9379), .QN(n13889) );
  INVX0 U14540 ( .INP(n12159), .ZN(n12153) );
  NAND2X0 U14541 ( .IN1(n13890), .IN2(g2370), .QN(n13886) );
  NAND2X0 U14542 ( .IN1(n13891), .IN2(n9379), .QN(n13890) );
  INVX0 U14543 ( .INP(n13892), .ZN(n13891) );
  NOR2X0 U14544 ( .IN1(n12150), .IN2(n9696), .QN(n13892) );
  NOR2X0 U14545 ( .IN1(n8507), .IN2(n8851), .QN(n9696) );
  NAND4X0 U14546 ( .IN1(n13893), .IN2(n13894), .IN3(n13895), .IN4(n13896), 
        .QN(g29250) );
  NAND2X0 U14547 ( .IN1(n13289), .IN2(g2299), .QN(n13896) );
  NOR2X0 U14548 ( .IN1(n13288), .IN2(n9402), .QN(n13289) );
  NAND3X0 U14549 ( .IN1(g2319), .IN2(g2351), .IN3(n13312), .QN(n13288) );
  NAND2X0 U14550 ( .IN1(n3555), .IN2(n13897), .QN(n13895) );
  NAND3X0 U14551 ( .IN1(n13898), .IN2(n13899), .IN3(n13900), .QN(n13897) );
  NAND2X0 U14552 ( .IN1(n8851), .IN2(g2295), .QN(n13900) );
  NOR2X0 U14553 ( .IN1(n8869), .IN2(g2319), .QN(n8851) );
  NAND2X0 U14554 ( .IN1(n5511), .IN2(n13901), .QN(n13899) );
  NAND2X0 U14555 ( .IN1(n13902), .IN2(n13903), .QN(n13901) );
  NAND2X0 U14556 ( .IN1(n5375), .IN2(g2307), .QN(n13903) );
  NAND2X0 U14557 ( .IN1(test_so21), .IN2(g2315), .QN(n13902) );
  NAND2X0 U14558 ( .IN1(n13904), .IN2(n8869), .QN(n13898) );
  NAND2X0 U14559 ( .IN1(n13905), .IN2(n13906), .QN(n13904) );
  NAND2X0 U14560 ( .IN1(g2319), .IN2(n9314), .QN(n13906) );
  NAND2X0 U14561 ( .IN1(g2351), .IN2(g2303), .QN(n13905) );
  NOR2X0 U14562 ( .IN1(n12150), .IN2(n9402), .QN(n3555) );
  NAND2X0 U14563 ( .IN1(n12159), .IN2(g2370), .QN(n13894) );
  NOR2X0 U14564 ( .IN1(n13312), .IN2(n9402), .QN(n12159) );
  INVX0 U14565 ( .INP(n12150), .ZN(n13312) );
  NAND3X0 U14566 ( .IN1(n13863), .IN2(n13209), .IN3(n13907), .QN(n12150) );
  NAND2X0 U14567 ( .IN1(n13205), .IN2(g2807), .QN(n13907) );
  NAND2X0 U14568 ( .IN1(n9431), .IN2(g2351), .QN(n13893) );
  NAND2X0 U14569 ( .IN1(n13908), .IN2(n13909), .QN(g29249) );
  NAND2X0 U14570 ( .IN1(n13910), .IN2(g2250), .QN(n13909) );
  NAND2X0 U14571 ( .IN1(n12174), .IN2(n13911), .QN(n13910) );
  NAND2X0 U14572 ( .IN1(n4414), .IN2(n9379), .QN(n13911) );
  INVX0 U14573 ( .INP(n12180), .ZN(n12174) );
  NAND2X0 U14574 ( .IN1(n13912), .IN2(g2236), .QN(n13908) );
  NAND2X0 U14575 ( .IN1(n13913), .IN2(n9379), .QN(n13912) );
  INVX0 U14576 ( .INP(n13914), .ZN(n13913) );
  NOR2X0 U14577 ( .IN1(n12171), .IN2(n9695), .QN(n13914) );
  NOR2X0 U14578 ( .IN1(n8503), .IN2(n8856), .QN(n9695) );
  NAND4X0 U14579 ( .IN1(n13915), .IN2(n13916), .IN3(n13917), .IN4(n13918), 
        .QN(g29248) );
  NAND2X0 U14580 ( .IN1(n13322), .IN2(g2165), .QN(n13918) );
  NOR2X0 U14581 ( .IN1(n13321), .IN2(n9400), .QN(n13322) );
  NAND3X0 U14582 ( .IN1(g2185), .IN2(g2217), .IN3(n13346), .QN(n13321) );
  NAND2X0 U14583 ( .IN1(n3574), .IN2(n13919), .QN(n13917) );
  NAND3X0 U14584 ( .IN1(n13920), .IN2(n13921), .IN3(n13922), .QN(n13919) );
  NAND2X0 U14585 ( .IN1(n8856), .IN2(g2161), .QN(n13922) );
  NOR2X0 U14586 ( .IN1(g2185), .IN2(n8756), .QN(n8856) );
  NAND2X0 U14587 ( .IN1(n5512), .IN2(n13923), .QN(n13921) );
  NAND2X0 U14588 ( .IN1(n13924), .IN2(n13925), .QN(n13923) );
  NAND2X0 U14589 ( .IN1(n5376), .IN2(g2173), .QN(n13925) );
  NAND2X0 U14590 ( .IN1(g2181), .IN2(g2208), .QN(n13924) );
  NAND2X0 U14591 ( .IN1(n8756), .IN2(n13926), .QN(n13920) );
  NAND2X0 U14592 ( .IN1(n13927), .IN2(n13928), .QN(n13926) );
  NAND2X0 U14593 ( .IN1(g2185), .IN2(n9352), .QN(n13928) );
  NAND2X0 U14594 ( .IN1(g2217), .IN2(g2169), .QN(n13927) );
  NOR2X0 U14595 ( .IN1(n12171), .IN2(n9400), .QN(n3574) );
  NAND2X0 U14596 ( .IN1(n12180), .IN2(g2236), .QN(n13916) );
  NOR2X0 U14597 ( .IN1(n13346), .IN2(n9400), .QN(n12180) );
  INVX0 U14598 ( .INP(n12171), .ZN(n13346) );
  NAND3X0 U14599 ( .IN1(n13929), .IN2(n13863), .IN3(n13208), .QN(n12171) );
  NAND2X0 U14600 ( .IN1(n13205), .IN2(g2803), .QN(n13929) );
  NAND2X0 U14601 ( .IN1(n9431), .IN2(g2217), .QN(n13915) );
  NAND2X0 U14602 ( .IN1(n13930), .IN2(n13931), .QN(g29247) );
  NAND2X0 U14603 ( .IN1(n13932), .IN2(g2079), .QN(n13931) );
  NAND2X0 U14604 ( .IN1(n13933), .IN2(n9379), .QN(n13932) );
  INVX0 U14605 ( .INP(n13934), .ZN(n13933) );
  NOR2X0 U14606 ( .IN1(n12192), .IN2(n9694), .QN(n13934) );
  NOR2X0 U14607 ( .IN1(n8885), .IN2(n8858), .QN(n9694) );
  NAND2X0 U14608 ( .IN1(test_so78), .IN2(n13935), .QN(n13930) );
  NAND2X0 U14609 ( .IN1(n12195), .IN2(n13936), .QN(n13935) );
  NAND2X0 U14610 ( .IN1(n4425), .IN2(n9379), .QN(n13936) );
  INVX0 U14611 ( .INP(n12201), .ZN(n12195) );
  NAND4X0 U14612 ( .IN1(n13937), .IN2(n13938), .IN3(n13939), .IN4(n13940), 
        .QN(g29246) );
  NAND2X0 U14613 ( .IN1(n13355), .IN2(g2008), .QN(n13940) );
  NOR2X0 U14614 ( .IN1(n13354), .IN2(n9399), .QN(n13355) );
  NAND3X0 U14615 ( .IN1(g2028), .IN2(g2060), .IN3(n13377), .QN(n13354) );
  NAND2X0 U14616 ( .IN1(n3593), .IN2(n13941), .QN(n13939) );
  NAND3X0 U14617 ( .IN1(n13942), .IN2(n13943), .IN3(n13944), .QN(n13941) );
  NAND2X0 U14618 ( .IN1(n8858), .IN2(g2004), .QN(n13944) );
  NOR2X0 U14619 ( .IN1(g2028), .IN2(n8760), .QN(n8858) );
  NAND2X0 U14620 ( .IN1(n5507), .IN2(n13945), .QN(n13943) );
  NAND2X0 U14621 ( .IN1(n13946), .IN2(n13947), .QN(n13945) );
  NAND2X0 U14622 ( .IN1(n5371), .IN2(g2016), .QN(n13947) );
  NAND2X0 U14623 ( .IN1(g2024), .IN2(g2051), .QN(n13946) );
  NAND2X0 U14624 ( .IN1(n8760), .IN2(n13948), .QN(n13942) );
  NAND2X0 U14625 ( .IN1(n13949), .IN2(n13950), .QN(n13948) );
  NAND2X0 U14626 ( .IN1(g2028), .IN2(n9312), .QN(n13950) );
  NAND2X0 U14627 ( .IN1(g2060), .IN2(g2012), .QN(n13949) );
  NOR2X0 U14628 ( .IN1(n12192), .IN2(n9399), .QN(n3593) );
  NAND2X0 U14629 ( .IN1(n12201), .IN2(g2079), .QN(n13938) );
  NOR2X0 U14630 ( .IN1(n13377), .IN2(n9399), .QN(n12201) );
  INVX0 U14631 ( .INP(n12192), .ZN(n13377) );
  NAND3X0 U14632 ( .IN1(n13951), .IN2(n13863), .IN3(n13185), .QN(n12192) );
  NAND2X0 U14633 ( .IN1(n13205), .IN2(g2787), .QN(n13951) );
  NAND2X0 U14634 ( .IN1(n9430), .IN2(g2060), .QN(n13937) );
  NAND2X0 U14635 ( .IN1(n13952), .IN2(n13953), .QN(g29245) );
  NAND2X0 U14636 ( .IN1(n13954), .IN2(g1959), .QN(n13953) );
  NAND2X0 U14637 ( .IN1(n12216), .IN2(n13955), .QN(n13954) );
  NAND2X0 U14638 ( .IN1(n4436), .IN2(n9379), .QN(n13955) );
  INVX0 U14639 ( .INP(n12222), .ZN(n12216) );
  NAND2X0 U14640 ( .IN1(test_so53), .IN2(n13956), .QN(n13952) );
  NAND2X0 U14641 ( .IN1(n13957), .IN2(n9379), .QN(n13956) );
  INVX0 U14642 ( .INP(n13958), .ZN(n13957) );
  NOR2X0 U14643 ( .IN1(n12213), .IN2(n9693), .QN(n13958) );
  NOR2X0 U14644 ( .IN1(n8511), .IN2(n8848), .QN(n9693) );
  NAND4X0 U14645 ( .IN1(n13959), .IN2(n13960), .IN3(n13961), .IN4(n13962), 
        .QN(g29244) );
  NAND2X0 U14646 ( .IN1(n13386), .IN2(g1874), .QN(n13962) );
  NOR2X0 U14647 ( .IN1(n13385), .IN2(n9406), .QN(n13386) );
  NAND3X0 U14648 ( .IN1(g1894), .IN2(g1926), .IN3(n13409), .QN(n13385) );
  NAND2X0 U14649 ( .IN1(n3611), .IN2(n13963), .QN(n13961) );
  NAND3X0 U14650 ( .IN1(n13964), .IN2(n13965), .IN3(n13966), .QN(n13963) );
  NAND2X0 U14651 ( .IN1(n8848), .IN2(g1870), .QN(n13966) );
  NOR2X0 U14652 ( .IN1(g1894), .IN2(n8757), .QN(n8848) );
  NAND2X0 U14653 ( .IN1(n5510), .IN2(n13967), .QN(n13965) );
  NAND2X0 U14654 ( .IN1(n13968), .IN2(n13969), .QN(n13967) );
  NAND2X0 U14655 ( .IN1(n5374), .IN2(g1882), .QN(n13969) );
  NAND2X0 U14656 ( .IN1(g1890), .IN2(g1917), .QN(n13968) );
  NAND2X0 U14657 ( .IN1(n8757), .IN2(n13970), .QN(n13964) );
  NAND2X0 U14658 ( .IN1(n13971), .IN2(n13972), .QN(n13970) );
  NAND2X0 U14659 ( .IN1(g1894), .IN2(n9280), .QN(n13972) );
  NAND2X0 U14660 ( .IN1(g1926), .IN2(g1878), .QN(n13971) );
  NOR2X0 U14661 ( .IN1(n12213), .IN2(n9405), .QN(n3611) );
  NAND2X0 U14662 ( .IN1(n12222), .IN2(test_so53), .QN(n13960) );
  NOR2X0 U14663 ( .IN1(n13409), .IN2(n9390), .QN(n12222) );
  INVX0 U14664 ( .INP(n12213), .ZN(n13409) );
  NAND3X0 U14665 ( .IN1(n13973), .IN2(n13863), .IN3(n13186), .QN(n12213) );
  NAND2X0 U14666 ( .IN1(n13205), .IN2(g2783), .QN(n13973) );
  NAND2X0 U14667 ( .IN1(n9430), .IN2(g1926), .QN(n13959) );
  NAND2X0 U14668 ( .IN1(n13974), .IN2(n13975), .QN(g29243) );
  NAND2X0 U14669 ( .IN1(n13976), .IN2(g1825), .QN(n13975) );
  NAND2X0 U14670 ( .IN1(n12237), .IN2(n13977), .QN(n13976) );
  NAND2X0 U14671 ( .IN1(n4447), .IN2(n9379), .QN(n13977) );
  INVX0 U14672 ( .INP(n12243), .ZN(n12237) );
  NAND2X0 U14673 ( .IN1(n13978), .IN2(g1811), .QN(n13974) );
  NAND2X0 U14674 ( .IN1(n13979), .IN2(n9379), .QN(n13978) );
  INVX0 U14675 ( .INP(n13980), .ZN(n13979) );
  NOR2X0 U14676 ( .IN1(n12234), .IN2(n9692), .QN(n13980) );
  NOR2X0 U14677 ( .IN1(n8505), .IN2(n8854), .QN(n9692) );
  NAND4X0 U14678 ( .IN1(n13981), .IN2(n13982), .IN3(n13983), .IN4(n13984), 
        .QN(g29242) );
  NAND2X0 U14679 ( .IN1(n13419), .IN2(g1740), .QN(n13984) );
  NOR2X0 U14680 ( .IN1(n13418), .IN2(n9392), .QN(n13419) );
  NAND3X0 U14681 ( .IN1(g1792), .IN2(g1760), .IN3(n13443), .QN(n13418) );
  NAND2X0 U14682 ( .IN1(n3628), .IN2(n13985), .QN(n13983) );
  NAND3X0 U14683 ( .IN1(n13986), .IN2(n13987), .IN3(n13988), .QN(n13985) );
  NAND2X0 U14684 ( .IN1(n8854), .IN2(g1736), .QN(n13988) );
  NOR2X0 U14685 ( .IN1(g1760), .IN2(n5596), .QN(n8854) );
  NAND2X0 U14686 ( .IN1(n5359), .IN2(n13989), .QN(n13987) );
  NAND2X0 U14687 ( .IN1(n13990), .IN2(n13991), .QN(n13989) );
  NAND2X0 U14688 ( .IN1(g1783), .IN2(g1756), .QN(n13991) );
  NAND2X0 U14689 ( .IN1(n5602), .IN2(g1748), .QN(n13990) );
  NAND2X0 U14690 ( .IN1(n5596), .IN2(n13992), .QN(n13986) );
  NAND2X0 U14691 ( .IN1(n13993), .IN2(n13994), .QN(n13992) );
  NAND2X0 U14692 ( .IN1(g1792), .IN2(g1744), .QN(n13994) );
  NAND2X0 U14693 ( .IN1(g1760), .IN2(g1752), .QN(n13993) );
  NOR2X0 U14694 ( .IN1(n12234), .IN2(n9394), .QN(n3628) );
  NAND2X0 U14695 ( .IN1(n12243), .IN2(g1811), .QN(n13982) );
  NOR2X0 U14696 ( .IN1(n13443), .IN2(n9399), .QN(n12243) );
  INVX0 U14697 ( .INP(n12234), .ZN(n13443) );
  NAND3X0 U14698 ( .IN1(n13863), .IN2(n13209), .IN3(n13995), .QN(n12234) );
  NAND2X0 U14699 ( .IN1(n13205), .IN2(g2775), .QN(n13995) );
  NOR2X0 U14700 ( .IN1(g2719), .IN2(n5299), .QN(n13209) );
  NAND2X0 U14701 ( .IN1(n9431), .IN2(g1792), .QN(n13981) );
  NAND2X0 U14702 ( .IN1(n13996), .IN2(n13997), .QN(g29241) );
  NAND2X0 U14703 ( .IN1(n13998), .IN2(g1691), .QN(n13997) );
  NAND2X0 U14704 ( .IN1(n12258), .IN2(n13999), .QN(n13998) );
  NAND2X0 U14705 ( .IN1(n4458), .IN2(n9379), .QN(n13999) );
  NAND2X0 U14706 ( .IN1(n14000), .IN2(g1677), .QN(n13996) );
  NAND2X0 U14707 ( .IN1(n14001), .IN2(n9379), .QN(n14000) );
  INVX0 U14708 ( .INP(n14002), .ZN(n14001) );
  NOR2X0 U14709 ( .IN1(n12255), .IN2(n9691), .QN(n14002) );
  NOR2X0 U14710 ( .IN1(n8509), .IN2(n8857), .QN(n9691) );
  NAND4X0 U14711 ( .IN1(n14003), .IN2(n14004), .IN3(n14005), .IN4(n14006), 
        .QN(g29240) );
  NAND2X0 U14712 ( .IN1(n3646), .IN2(n14007), .QN(n14006) );
  NAND4X0 U14713 ( .IN1(n14008), .IN2(n14009), .IN3(n14010), .IN4(n14011), 
        .QN(n14007) );
  NAND3X0 U14714 ( .IN1(n5370), .IN2(g1612), .IN3(n5525), .QN(n14011) );
  NAND2X0 U14715 ( .IN1(n14012), .IN2(n8870), .QN(n14010) );
  NAND2X0 U14716 ( .IN1(n14013), .IN2(n14014), .QN(n14012) );
  NAND2X0 U14717 ( .IN1(g1624), .IN2(n9303), .QN(n14014) );
  NAND2X0 U14718 ( .IN1(g1657), .IN2(g1608), .QN(n14013) );
  NAND2X0 U14719 ( .IN1(g25167), .IN2(g1620), .QN(n14009) );
  NAND2X0 U14720 ( .IN1(n8857), .IN2(g1600), .QN(n14008) );
  NOR2X0 U14721 ( .IN1(n8870), .IN2(g1624), .QN(n8857) );
  NOR2X0 U14722 ( .IN1(n12255), .IN2(n9388), .QN(n3646) );
  NAND2X0 U14723 ( .IN1(n13450), .IN2(g1604), .QN(n14005) );
  NOR3X0 U14724 ( .IN1(n5370), .IN2(n5525), .IN3(n12255), .QN(n13450) );
  NAND2X0 U14725 ( .IN1(n12271), .IN2(g1677), .QN(n14004) );
  INVX0 U14726 ( .INP(n12258), .ZN(n12271) );
  NAND2X0 U14727 ( .IN1(n12255), .IN2(n9379), .QN(n12258) );
  NAND3X0 U14728 ( .IN1(n14015), .IN2(n13863), .IN3(n13208), .QN(n12255) );
  NOR2X0 U14729 ( .IN1(g2719), .IN2(g2715), .QN(n13208) );
  INVX0 U14730 ( .INP(n14016), .ZN(n13863) );
  NOR2X0 U14731 ( .IN1(n10547), .IN2(n4388), .QN(n14016) );
  INVX0 U14732 ( .INP(n13205), .ZN(n10547) );
  NAND2X0 U14733 ( .IN1(n13205), .IN2(g2771), .QN(n14015) );
  NOR2X0 U14734 ( .IN1(g2729), .IN2(g2724), .QN(n13205) );
  NAND2X0 U14735 ( .IN1(n9431), .IN2(g1657), .QN(n14003) );
  NAND3X0 U14736 ( .IN1(n14017), .IN2(n14018), .IN3(n14019), .QN(g29239) );
  NAND3X0 U14737 ( .IN1(n14020), .IN2(n13495), .IN3(n14021), .QN(n14019) );
  INVX0 U14738 ( .INP(n14022), .ZN(n14020) );
  NAND2X0 U14739 ( .IN1(n9434), .IN2(g1478), .QN(n14018) );
  NAND3X0 U14740 ( .IN1(n14023), .IN2(g1454), .IN3(n9342), .QN(n14017) );
  NAND2X0 U14741 ( .IN1(n14024), .IN2(n14022), .QN(n14023) );
  NAND2X0 U14742 ( .IN1(n14025), .IN2(n14026), .QN(n14022) );
  NAND2X0 U14743 ( .IN1(n5343), .IN2(n14027), .QN(n14026) );
  NAND2X0 U14744 ( .IN1(n14028), .IN2(g1448), .QN(n14025) );
  NAND3X0 U14745 ( .IN1(n14029), .IN2(n14030), .IN3(n14031), .QN(g29238) );
  NAND2X0 U14746 ( .IN1(n14032), .IN2(g1484), .QN(n14031) );
  NAND2X0 U14747 ( .IN1(n9507), .IN2(g1472), .QN(n14030) );
  NAND4X0 U14748 ( .IN1(n14033), .IN2(n14034), .IN3(n14035), .IN4(n9361), .QN(
        n14029) );
  NAND2X0 U14749 ( .IN1(n5865), .IN2(n14036), .QN(n14035) );
  NAND3X0 U14750 ( .IN1(n8717), .IN2(n5850), .IN3(n14037), .QN(n14036) );
  NAND2X0 U14751 ( .IN1(n5483), .IN2(n14027), .QN(n14034) );
  NAND2X0 U14752 ( .IN1(n14028), .IN2(g1300), .QN(n14033) );
  NAND3X0 U14753 ( .IN1(n14038), .IN2(n14039), .IN3(n14040), .QN(g29237) );
  NAND4X0 U14754 ( .IN1(n14041), .IN2(n14021), .IN3(test_so49), .IN4(g1514), 
        .QN(n14040) );
  INVX0 U14755 ( .INP(n14042), .ZN(n14041) );
  NAND2X0 U14756 ( .IN1(n9509), .IN2(g1448), .QN(n14039) );
  NAND3X0 U14757 ( .IN1(n14043), .IN2(g1467), .IN3(n9341), .QN(n14038) );
  NAND3X0 U14758 ( .IN1(test_so49), .IN2(n14042), .IN3(n14044), .QN(n14043) );
  NAND2X0 U14759 ( .IN1(n14045), .IN2(n14046), .QN(n14042) );
  NAND2X0 U14760 ( .IN1(n5290), .IN2(n14027), .QN(n14046) );
  NAND2X0 U14761 ( .IN1(n14028), .IN2(g1472), .QN(n14045) );
  NAND3X0 U14762 ( .IN1(n14047), .IN2(n14048), .IN3(n14049), .QN(g29236) );
  NAND4X0 U14763 ( .IN1(n14050), .IN2(n14021), .IN3(g1514), .IN4(n8859), .QN(
        n14049) );
  NOR4X0 U14764 ( .IN1(g1442), .IN2(g1489), .IN3(n9386), .IN4(n8798), .QN(
        n14021) );
  INVX0 U14765 ( .INP(n14051), .ZN(n14050) );
  NAND2X0 U14766 ( .IN1(n9493), .IN2(g1442), .QN(n14048) );
  NAND3X0 U14767 ( .IN1(n14052), .IN2(g1437), .IN3(n9341), .QN(n14047) );
  NAND3X0 U14768 ( .IN1(n14051), .IN2(n8859), .IN3(n14044), .QN(n14052) );
  NAND2X0 U14769 ( .IN1(n14053), .IN2(n14054), .QN(n14051) );
  NAND2X0 U14770 ( .IN1(n5289), .IN2(n14027), .QN(n14054) );
  NAND2X0 U14771 ( .IN1(n14028), .IN2(g1478), .QN(n14053) );
  INVX0 U14772 ( .INP(n14027), .ZN(n14028) );
  NAND2X0 U14773 ( .IN1(n10199), .IN2(DFF_1092_n1), .QN(n14027) );
  NAND3X0 U14774 ( .IN1(n14055), .IN2(n14056), .IN3(n14057), .QN(g29235) );
  NAND2X0 U14775 ( .IN1(n9492), .IN2(g1252), .QN(n14057) );
  NAND3X0 U14776 ( .IN1(n11853), .IN2(n14058), .IN3(g1256), .QN(n14056) );
  INVX0 U14777 ( .INP(n4178), .ZN(n14058) );
  NAND2X0 U14778 ( .IN1(n4178), .IN2(n5558), .QN(n14055) );
  NAND3X0 U14779 ( .IN1(n14059), .IN2(n14060), .IN3(n14061), .QN(g29234) );
  NAND3X0 U14780 ( .IN1(n14062), .IN2(n13532), .IN3(n14063), .QN(n14061) );
  INVX0 U14781 ( .INP(n14064), .ZN(n14062) );
  NAND2X0 U14782 ( .IN1(n9494), .IN2(g1135), .QN(n14060) );
  NAND3X0 U14783 ( .IN1(test_so90), .IN2(n14065), .IN3(n9341), .QN(n14059) );
  NAND2X0 U14784 ( .IN1(n14066), .IN2(n14064), .QN(n14065) );
  NAND2X0 U14785 ( .IN1(n14067), .IN2(n14068), .QN(n14064) );
  NAND2X0 U14786 ( .IN1(n5478), .IN2(n14069), .QN(n14068) );
  NAND2X0 U14787 ( .IN1(n14070), .IN2(g1105), .QN(n14067) );
  NAND3X0 U14788 ( .IN1(n14071), .IN2(n14072), .IN3(n14073), .QN(g29233) );
  NAND2X0 U14789 ( .IN1(n14074), .IN2(g1141), .QN(n14073) );
  NAND2X0 U14790 ( .IN1(n9496), .IN2(g1129), .QN(n14072) );
  NAND4X0 U14791 ( .IN1(n14075), .IN2(n14076), .IN3(n14077), .IN4(n9361), .QN(
        n14071) );
  NAND2X0 U14792 ( .IN1(n5691), .IN2(n14078), .QN(n14077) );
  NAND3X0 U14793 ( .IN1(n5851), .IN2(n8865), .IN3(n14079), .QN(n14078) );
  NAND2X0 U14794 ( .IN1(n5341), .IN2(n14069), .QN(n14076) );
  NAND2X0 U14795 ( .IN1(n14070), .IN2(g956), .QN(n14075) );
  NAND3X0 U14796 ( .IN1(n14080), .IN2(n14081), .IN3(n14082), .QN(g29232) );
  NAND3X0 U14797 ( .IN1(n14063), .IN2(n11762), .IN3(n14083), .QN(n14082) );
  INVX0 U14798 ( .INP(n14084), .ZN(n14083) );
  NAND2X0 U14799 ( .IN1(n9495), .IN2(g1105), .QN(n14081) );
  NAND3X0 U14800 ( .IN1(n14085), .IN2(g1124), .IN3(n9341), .QN(n14080) );
  NAND3X0 U14801 ( .IN1(n14084), .IN2(g13259), .IN3(n11762), .QN(n14085) );
  NAND2X0 U14802 ( .IN1(n14086), .IN2(n14087), .QN(n14084) );
  NAND2X0 U14803 ( .IN1(n5329), .IN2(n14069), .QN(n14087) );
  NAND2X0 U14804 ( .IN1(n14070), .IN2(g1129), .QN(n14086) );
  NAND3X0 U14805 ( .IN1(n14088), .IN2(n14089), .IN3(n14090), .QN(g29231) );
  NAND4X0 U14806 ( .IN1(n14091), .IN2(n14063), .IN3(n5599), .IN4(g1171), .QN(
        n14090) );
  NOR4X0 U14807 ( .IN1(g1146), .IN2(n9385), .IN3(n8804), .IN4(test_so7), .QN(
        n14063) );
  INVX0 U14808 ( .INP(n14092), .ZN(n14091) );
  NAND2X0 U14809 ( .IN1(test_so7), .IN2(n9515), .QN(n14089) );
  NAND3X0 U14810 ( .IN1(n14093), .IN2(g1094), .IN3(n9341), .QN(n14088) );
  NAND2X0 U14811 ( .IN1(n14094), .IN2(n14092), .QN(n14093) );
  NAND2X0 U14812 ( .IN1(n14095), .IN2(n14096), .QN(n14092) );
  NAND2X0 U14813 ( .IN1(n5328), .IN2(n14069), .QN(n14096) );
  NAND2X0 U14814 ( .IN1(n14070), .IN2(g1135), .QN(n14095) );
  INVX0 U14815 ( .INP(n14069), .ZN(n14070) );
  NAND2X0 U14816 ( .IN1(n10198), .IN2(DFF_24_n1), .QN(n14069) );
  NAND3X0 U14817 ( .IN1(n14097), .IN2(n14098), .IN3(n14099), .QN(g29230) );
  NAND2X0 U14818 ( .IN1(n9461), .IN2(g907), .QN(n14099) );
  NAND3X0 U14819 ( .IN1(n11867), .IN2(n14100), .IN3(g911), .QN(n14098) );
  INVX0 U14820 ( .INP(n4196), .ZN(n14100) );
  NAND2X0 U14821 ( .IN1(n4196), .IN2(n5559), .QN(n14097) );
  NAND3X0 U14822 ( .IN1(n14101), .IN2(n14102), .IN3(n14103), .QN(g29229) );
  NAND2X0 U14823 ( .IN1(n9461), .IN2(g827), .QN(n14103) );
  NAND2X0 U14824 ( .IN1(n4517), .IN2(g723), .QN(n14102) );
  NAND3X0 U14825 ( .IN1(n4516), .IN2(n14104), .IN3(n5826), .QN(n14101) );
  NAND2X0 U14826 ( .IN1(n14105), .IN2(n14106), .QN(g29228) );
  NAND2X0 U14827 ( .IN1(n2404), .IN2(n14107), .QN(n14106) );
  NAND2X0 U14828 ( .IN1(n14108), .IN2(n14109), .QN(n14107) );
  NAND2X0 U14829 ( .IN1(test_so60), .IN2(n14110), .QN(n14109) );
  NAND2X0 U14830 ( .IN1(n13548), .IN2(n8904), .QN(n14108) );
  INVX0 U14831 ( .INP(n14110), .ZN(n13548) );
  NAND2X0 U14832 ( .IN1(n14111), .IN2(n14112), .QN(n14110) );
  NAND2X0 U14833 ( .IN1(n5482), .IN2(g12184), .QN(n14112) );
  INVX0 U14834 ( .INP(n13559), .ZN(n14111) );
  INVX0 U14835 ( .INP(n14113), .ZN(n14105) );
  NOR2X0 U14836 ( .IN1(n9360), .IN2(n8791), .QN(n14113) );
  NAND3X0 U14837 ( .IN1(n14114), .IN2(n14115), .IN3(n14116), .QN(g29227) );
  NAND2X0 U14838 ( .IN1(n9461), .IN2(g676), .QN(n14116) );
  NAND3X0 U14839 ( .IN1(n4523), .IN2(n14117), .IN3(n8879), .QN(n14115) );
  NAND2X0 U14840 ( .IN1(n4524), .IN2(test_so70), .QN(n14114) );
  NAND3X0 U14841 ( .IN1(n14118), .IN2(n14119), .IN3(n14120), .QN(g29226) );
  NAND2X0 U14842 ( .IN1(n9461), .IN2(g671), .QN(n14120) );
  NAND3X0 U14843 ( .IN1(n4525), .IN2(n14121), .IN3(g676), .QN(n14119) );
  INVX0 U14844 ( .INP(n4526), .ZN(n14121) );
  NAND3X0 U14845 ( .IN1(n4526), .IN2(n14117), .IN3(n5751), .QN(n14118) );
  NAND2X0 U14846 ( .IN1(n14122), .IN2(n14123), .QN(g29225) );
  NAND3X0 U14847 ( .IN1(n14124), .IN2(n14125), .IN3(n4525), .QN(n14123) );
  NOR2X0 U14848 ( .IN1(n14126), .IN2(n9402), .QN(n4525) );
  INVX0 U14849 ( .INP(n14117), .ZN(n14126) );
  NOR2X0 U14850 ( .IN1(n5821), .IN2(n14127), .QN(n14117) );
  NOR4X0 U14851 ( .IN1(n4535), .IN2(n14128), .IN3(n8844), .IN4(n8441), .QN(
        n14127) );
  NAND2X0 U14852 ( .IN1(n14129), .IN2(n14130), .QN(n4535) );
  NAND2X0 U14853 ( .IN1(n8829), .IN2(g655), .QN(n14130) );
  NAND2X0 U14854 ( .IN1(n8827), .IN2(g718), .QN(n14129) );
  NAND2X0 U14855 ( .IN1(n8364), .IN2(n8844), .QN(n14125) );
  INVX0 U14856 ( .INP(n14131), .ZN(n8844) );
  NAND2X0 U14857 ( .IN1(n14131), .IN2(g671), .QN(n14124) );
  NAND2X0 U14858 ( .IN1(n9461), .IN2(g667), .QN(n14122) );
  NAND3X0 U14859 ( .IN1(n14132), .IN2(n14133), .IN3(n14134), .QN(g29224) );
  NAND2X0 U14860 ( .IN1(n9461), .IN2(g572), .QN(n14134) );
  NAND3X0 U14861 ( .IN1(n2421), .IN2(n14135), .IN3(g586), .QN(n14133) );
  INVX0 U14862 ( .INP(n4201), .ZN(n14135) );
  NAND2X0 U14863 ( .IN1(n4201), .IN2(n5336), .QN(n14132) );
  NAND3X0 U14864 ( .IN1(n14136), .IN2(n14137), .IN3(n14138), .QN(g29223) );
  NAND2X0 U14865 ( .IN1(n14139), .IN2(n5708), .QN(n14138) );
  NAND2X0 U14866 ( .IN1(n9461), .IN2(g482), .QN(n14137) );
  NAND2X0 U14867 ( .IN1(n14140), .IN2(n9379), .QN(n14136) );
  NAND2X0 U14868 ( .IN1(n14141), .IN2(n14142), .QN(n14140) );
  INVX0 U14869 ( .INP(n14143), .ZN(n14142) );
  NOR2X0 U14870 ( .IN1(n14139), .IN2(n5708), .QN(n14143) );
  NAND3X0 U14871 ( .IN1(n14144), .IN2(n14145), .IN3(n14146), .QN(g29222) );
  NAND2X0 U14872 ( .IN1(n14147), .IN2(g411), .QN(n14146) );
  INVX0 U14873 ( .INP(n14148), .ZN(n14145) );
  NOR2X0 U14874 ( .IN1(n14149), .IN2(n5358), .QN(n14148) );
  NOR2X0 U14875 ( .IN1(n14150), .IN2(n9399), .QN(n14149) );
  NOR2X0 U14876 ( .IN1(n14151), .IN2(n488), .QN(n14150) );
  NAND3X0 U14877 ( .IN1(n14152), .IN2(n488), .IN3(n5358), .QN(n14144) );
  NAND2X0 U14878 ( .IN1(n14153), .IN2(n14154), .QN(n488) );
  INVX0 U14879 ( .INP(n14155), .ZN(n14154) );
  NOR2X0 U14880 ( .IN1(n14156), .IN2(g417), .QN(n14155) );
  NAND2X0 U14881 ( .IN1(n14156), .IN2(g417), .QN(n14153) );
  NAND2X0 U14882 ( .IN1(n14157), .IN2(n14158), .QN(n14156) );
  NAND2X0 U14883 ( .IN1(n14159), .IN2(g392), .QN(n14158) );
  NAND2X0 U14884 ( .IN1(n14160), .IN2(n14161), .QN(n14159) );
  NAND2X0 U14885 ( .IN1(g401), .IN2(g405), .QN(n14161) );
  NAND2X0 U14886 ( .IN1(n8786), .IN2(g437), .QN(n14160) );
  NAND2X0 U14887 ( .IN1(n14162), .IN2(n8787), .QN(n14157) );
  NAND2X0 U14888 ( .IN1(n14163), .IN2(n14164), .QN(n14162) );
  NAND2X0 U14889 ( .IN1(n8786), .IN2(g424), .QN(n14164) );
  NAND2X0 U14890 ( .IN1(g437), .IN2(g405), .QN(n14163) );
  NAND3X0 U14891 ( .IN1(n14165), .IN2(n14166), .IN3(n14167), .QN(g28105) );
  NAND2X0 U14892 ( .IN1(n11388), .IN2(g5011), .QN(n14167) );
  NAND2X0 U14893 ( .IN1(n9460), .IN2(g6657), .QN(n14166) );
  NAND3X0 U14894 ( .IN1(n13598), .IN2(n11381), .IN3(n9341), .QN(n14165) );
  NAND2X0 U14895 ( .IN1(n14168), .IN2(n14169), .QN(n13598) );
  NAND2X0 U14896 ( .IN1(n5531), .IN2(n14170), .QN(n14169) );
  NAND4X0 U14897 ( .IN1(n14171), .IN2(n14172), .IN3(n14173), .IN4(n14174), 
        .QN(n14170) );
  NOR3X0 U14898 ( .IN1(n14175), .IN2(n14176), .IN3(n14177), .QN(n14174) );
  NOR2X0 U14899 ( .IN1(n14178), .IN2(n8882), .QN(n14177) );
  NOR2X0 U14900 ( .IN1(n14179), .IN2(n14180), .QN(n14178) );
  NOR2X0 U14901 ( .IN1(n8611), .IN2(n14181), .QN(n14179) );
  NOR2X0 U14902 ( .IN1(test_so80), .IN2(n14182), .QN(n14176) );
  NOR2X0 U14903 ( .IN1(n14183), .IN2(n14184), .QN(n14175) );
  INVX0 U14904 ( .INP(n9685), .ZN(n14184) );
  NOR2X0 U14905 ( .IN1(n14185), .IN2(n14186), .QN(n14183) );
  NOR2X0 U14906 ( .IN1(n8670), .IN2(n8669), .QN(n14186) );
  NOR2X0 U14907 ( .IN1(n8668), .IN2(n8667), .QN(n14185) );
  NAND2X0 U14908 ( .IN1(n9682), .IN2(n14187), .QN(n14173) );
  NAND2X0 U14909 ( .IN1(n14188), .IN2(n14189), .QN(n14187) );
  NAND2X0 U14910 ( .IN1(g6723), .IN2(g6605), .QN(n14189) );
  NAND2X0 U14911 ( .IN1(g13099), .IN2(g6593), .QN(n14188) );
  NAND3X0 U14912 ( .IN1(g14749), .IN2(g6633), .IN3(n9683), .QN(n14172) );
  NAND3X0 U14913 ( .IN1(g17871), .IN2(g6617), .IN3(n9684), .QN(n14171) );
  NAND2X0 U14914 ( .IN1(n14190), .IN2(g6727), .QN(n14168) );
  NAND4X0 U14915 ( .IN1(n14191), .IN2(n14192), .IN3(n14193), .IN4(n14194), 
        .QN(n14190) );
  INVX0 U14916 ( .INP(n14195), .ZN(n14194) );
  NAND3X0 U14917 ( .IN1(n14196), .IN2(n14197), .IN3(n14198), .QN(n14195) );
  NAND2X0 U14918 ( .IN1(n14199), .IN2(test_so80), .QN(n14198) );
  NAND2X0 U14919 ( .IN1(n14200), .IN2(n14182), .QN(n14199) );
  INVX0 U14920 ( .INP(n14201), .ZN(n14182) );
  NAND3X0 U14921 ( .IN1(n14202), .IN2(n14203), .IN3(n14204), .QN(n14201) );
  NAND3X0 U14922 ( .IN1(g14828), .IN2(g6613), .IN3(n9682), .QN(n14204) );
  NAND3X0 U14923 ( .IN1(g17688), .IN2(g6645), .IN3(n9683), .QN(n14203) );
  NAND3X0 U14924 ( .IN1(g17778), .IN2(g6629), .IN3(n9684), .QN(n14202) );
  NAND2X0 U14925 ( .IN1(n9685), .IN2(test_so71), .QN(n14200) );
  NAND2X0 U14926 ( .IN1(n8882), .IN2(n14180), .QN(n14197) );
  NAND3X0 U14927 ( .IN1(n14205), .IN2(n14206), .IN3(n14207), .QN(n14180) );
  NAND3X0 U14928 ( .IN1(g6637), .IN2(g17778), .IN3(n9685), .QN(n14207) );
  NAND3X0 U14929 ( .IN1(g14828), .IN2(g6621), .IN3(n9683), .QN(n14206) );
  NAND3X0 U14930 ( .IN1(g6653), .IN2(g17688), .IN3(n9682), .QN(n14205) );
  INVX0 U14931 ( .INP(n14208), .ZN(n14196) );
  NOR2X0 U14932 ( .IN1(n14209), .IN2(n14181), .QN(n14208) );
  INVX0 U14933 ( .INP(n9684), .ZN(n14181) );
  NOR2X0 U14934 ( .IN1(n5398), .IN2(n5590), .QN(n9684) );
  NOR2X0 U14935 ( .IN1(n14210), .IN2(n14211), .QN(n14209) );
  NOR2X0 U14936 ( .IN1(n8667), .IN2(n8485), .QN(n14211) );
  NOR2X0 U14937 ( .IN1(n8669), .IN2(n8484), .QN(n14210) );
  NAND2X0 U14938 ( .IN1(n9683), .IN2(n14212), .QN(n14193) );
  NAND2X0 U14939 ( .IN1(n14213), .IN2(n14214), .QN(n14212) );
  NAND2X0 U14940 ( .IN1(g6589), .IN2(g6723), .QN(n14214) );
  NAND2X0 U14941 ( .IN1(g6581), .IN2(g13099), .QN(n14213) );
  NOR2X0 U14942 ( .IN1(g6682), .IN2(g6741), .QN(n9683) );
  NAND3X0 U14943 ( .IN1(g14749), .IN2(g6625), .IN3(n9682), .QN(n14192) );
  NOR2X0 U14944 ( .IN1(g6741), .IN2(n5590), .QN(n9682) );
  NAND3X0 U14945 ( .IN1(g6609), .IN2(g17871), .IN3(n9685), .QN(n14191) );
  NOR2X0 U14946 ( .IN1(g6682), .IN2(n5398), .QN(n9685) );
  NAND3X0 U14947 ( .IN1(n14215), .IN2(n14216), .IN3(n14217), .QN(g28102) );
  NAND2X0 U14948 ( .IN1(n11404), .IN2(g4826), .QN(n14217) );
  NAND2X0 U14949 ( .IN1(n9460), .IN2(g6311), .QN(n14216) );
  NAND3X0 U14950 ( .IN1(n11393), .IN2(n13631), .IN3(n9341), .QN(n14215) );
  NAND2X0 U14951 ( .IN1(n14218), .IN2(n14219), .QN(n13631) );
  NAND2X0 U14952 ( .IN1(test_so69), .IN2(n14220), .QN(n14219) );
  NAND4X0 U14953 ( .IN1(n14221), .IN2(n14222), .IN3(n14223), .IN4(n14224), 
        .QN(n14220) );
  NOR3X0 U14954 ( .IN1(n14225), .IN2(n14226), .IN3(n14227), .QN(n14224) );
  NOR2X0 U14955 ( .IN1(n5437), .IN2(n14228), .QN(n14227) );
  NOR2X0 U14956 ( .IN1(n14229), .IN2(n14230), .QN(n14228) );
  NOR2X0 U14957 ( .IN1(n8493), .IN2(n14231), .QN(n14229) );
  INVX0 U14958 ( .INP(n14232), .ZN(n14226) );
  NAND2X0 U14959 ( .IN1(n14233), .IN2(n5437), .QN(n14232) );
  NOR2X0 U14960 ( .IN1(n14234), .IN2(n14235), .QN(n14225) );
  NOR2X0 U14961 ( .IN1(n14236), .IN2(n14237), .QN(n14234) );
  NOR2X0 U14962 ( .IN1(n8676), .IN2(n8491), .QN(n14237) );
  NOR2X0 U14963 ( .IN1(n8678), .IN2(n8490), .QN(n14236) );
  NAND2X0 U14964 ( .IN1(n14238), .IN2(n14239), .QN(n14223) );
  NAND2X0 U14965 ( .IN1(n14240), .IN2(n14241), .QN(n14239) );
  NAND2X0 U14966 ( .IN1(g6243), .IN2(g6377), .QN(n14241) );
  NAND2X0 U14967 ( .IN1(g6235), .IN2(g13085), .QN(n14240) );
  NAND3X0 U14968 ( .IN1(g6263), .IN2(g17845), .IN3(n11395), .QN(n14222) );
  NAND3X0 U14969 ( .IN1(g14705), .IN2(g6279), .IN3(n11400), .QN(n14221) );
  NAND2X0 U14970 ( .IN1(n14242), .IN2(n8889), .QN(n14218) );
  NAND4X0 U14971 ( .IN1(n14243), .IN2(n14244), .IN3(n14245), .IN4(n14246), 
        .QN(n14242) );
  NOR3X0 U14972 ( .IN1(n14247), .IN2(n14248), .IN3(n14249), .QN(n14246) );
  NOR2X0 U14973 ( .IN1(n5437), .IN2(n14250), .QN(n14249) );
  NOR2X0 U14974 ( .IN1(n14251), .IN2(n14233), .QN(n14250) );
  NAND3X0 U14975 ( .IN1(n14252), .IN2(n14253), .IN3(n14254), .QN(n14233) );
  NAND3X0 U14976 ( .IN1(g6307), .IN2(g17649), .IN3(n11400), .QN(n14254) );
  NAND3X0 U14977 ( .IN1(g6291), .IN2(g17760), .IN3(n11395), .QN(n14253) );
  NAND3X0 U14978 ( .IN1(g14779), .IN2(g6275), .IN3(n14238), .QN(n14252) );
  NOR2X0 U14979 ( .IN1(n8617), .IN2(n14235), .QN(n14251) );
  INVX0 U14980 ( .INP(n10581), .ZN(n14235) );
  INVX0 U14981 ( .INP(n14255), .ZN(n14248) );
  NAND2X0 U14982 ( .IN1(n14230), .IN2(n5437), .QN(n14255) );
  NAND3X0 U14983 ( .IN1(n14256), .IN2(n14257), .IN3(n14258), .QN(n14230) );
  NAND3X0 U14984 ( .IN1(g17760), .IN2(g6283), .IN3(n10581), .QN(n14258) );
  NAND3X0 U14985 ( .IN1(g17649), .IN2(g6299), .IN3(n14238), .QN(n14257) );
  NAND3X0 U14986 ( .IN1(g14779), .IN2(g6267), .IN3(n11400), .QN(n14256) );
  NOR2X0 U14987 ( .IN1(n14259), .IN2(n14260), .QN(n14247) );
  NOR2X0 U14988 ( .IN1(n14261), .IN2(n14262), .QN(n14259) );
  NOR2X0 U14989 ( .IN1(n8706), .IN2(n8705), .QN(n14262) );
  NOR2X0 U14990 ( .IN1(n8704), .IN2(n8703), .QN(n14261) );
  NAND2X0 U14991 ( .IN1(n11395), .IN2(n14263), .QN(n14245) );
  NAND2X0 U14992 ( .IN1(n14264), .IN2(n14265), .QN(n14263) );
  INVX0 U14993 ( .INP(n14266), .ZN(n14265) );
  NOR2X0 U14994 ( .IN1(n8676), .IN2(n8677), .QN(n14266) );
  NAND2X0 U14995 ( .IN1(g17685), .IN2(g6251), .QN(n14264) );
  NAND3X0 U14996 ( .IN1(g14705), .IN2(g6287), .IN3(n14238), .QN(n14244) );
  NAND3X0 U14997 ( .IN1(g17845), .IN2(g6271), .IN3(n10581), .QN(n14243) );
  NAND3X0 U14998 ( .IN1(n14267), .IN2(n14268), .IN3(n14269), .QN(g28099) );
  NAND2X0 U14999 ( .IN1(n11420), .IN2(g4831), .QN(n14269) );
  NAND2X0 U15000 ( .IN1(test_so13), .IN2(n9515), .QN(n14268) );
  NAND3X0 U15001 ( .IN1(n11409), .IN2(n13664), .IN3(n9341), .QN(n14267) );
  NAND2X0 U15002 ( .IN1(n14270), .IN2(n14271), .QN(n13664) );
  NAND2X0 U15003 ( .IN1(n5528), .IN2(n14272), .QN(n14271) );
  NAND4X0 U15004 ( .IN1(n14273), .IN2(n14274), .IN3(n14275), .IN4(n14276), 
        .QN(n14272) );
  NOR3X0 U15005 ( .IN1(n14277), .IN2(n14278), .IN3(n14279), .QN(n14276) );
  NOR2X0 U15006 ( .IN1(n5432), .IN2(n14280), .QN(n14279) );
  NOR2X0 U15007 ( .IN1(n14281), .IN2(n14282), .QN(n14280) );
  INVX0 U15008 ( .INP(n14283), .ZN(n14281) );
  NAND2X0 U15009 ( .IN1(n10586), .IN2(g5909), .QN(n14283) );
  NOR2X0 U15010 ( .IN1(n14284), .IN2(g12350), .QN(n14278) );
  NOR2X0 U15011 ( .IN1(n14285), .IN2(n14286), .QN(n14277) );
  NOR2X0 U15012 ( .IN1(n14287), .IN2(n14288), .QN(n14285) );
  NOR2X0 U15013 ( .IN1(n8686), .IN2(n8685), .QN(n14288) );
  NOR2X0 U15014 ( .IN1(n8684), .IN2(n8683), .QN(n14287) );
  NAND2X0 U15015 ( .IN1(n11411), .IN2(n14289), .QN(n14275) );
  NAND2X0 U15016 ( .IN1(n14290), .IN2(n14291), .QN(n14289) );
  NAND2X0 U15017 ( .IN1(g17715), .IN2(g5957), .QN(n14291) );
  NAND2X0 U15018 ( .IN1(g17646), .IN2(g5905), .QN(n14290) );
  NAND3X0 U15019 ( .IN1(g14673), .IN2(g5941), .IN3(n14292), .QN(n14274) );
  NAND3X0 U15020 ( .IN1(g17819), .IN2(g5925), .IN3(n10586), .QN(n14273) );
  NAND2X0 U15021 ( .IN1(n14293), .IN2(g6035), .QN(n14270) );
  NAND4X0 U15022 ( .IN1(n14294), .IN2(n14295), .IN3(n14296), .IN4(n14297), 
        .QN(n14293) );
  INVX0 U15023 ( .INP(n14298), .ZN(n14297) );
  NAND3X0 U15024 ( .IN1(n14299), .IN2(n14300), .IN3(n14301), .QN(n14298) );
  NAND2X0 U15025 ( .IN1(g12350), .IN2(n14302), .QN(n14301) );
  NAND2X0 U15026 ( .IN1(n14303), .IN2(n14284), .QN(n14302) );
  INVX0 U15027 ( .INP(n14304), .ZN(n14284) );
  NAND3X0 U15028 ( .IN1(n14305), .IN2(n14306), .IN3(n14307), .QN(n14304) );
  NAND3X0 U15029 ( .IN1(g17739), .IN2(g5937), .IN3(n10586), .QN(n14307) );
  NAND3X0 U15030 ( .IN1(g17607), .IN2(g5953), .IN3(n14292), .QN(n14306) );
  NAND3X0 U15031 ( .IN1(g14738), .IN2(g5921), .IN3(n11416), .QN(n14305) );
  NAND2X0 U15032 ( .IN1(g5893), .IN2(n11411), .QN(n14303) );
  NAND2X0 U15033 ( .IN1(n14282), .IN2(n5432), .QN(n14300) );
  NAND3X0 U15034 ( .IN1(n14308), .IN2(n14309), .IN3(n14310), .QN(n14282) );
  NAND3X0 U15035 ( .IN1(g5961), .IN2(g17607), .IN3(n11416), .QN(n14310) );
  NAND3X0 U15036 ( .IN1(g5945), .IN2(g17739), .IN3(n11411), .QN(n14309) );
  NAND3X0 U15037 ( .IN1(g14738), .IN2(g5929), .IN3(n14292), .QN(n14308) );
  NAND2X0 U15038 ( .IN1(n14311), .IN2(n10586), .QN(n14299) );
  NAND2X0 U15039 ( .IN1(n14312), .IN2(n14313), .QN(n14311) );
  NAND2X0 U15040 ( .IN1(g17646), .IN2(test_so13), .QN(n14313) );
  NAND2X0 U15041 ( .IN1(g17715), .IN2(g5949), .QN(n14312) );
  NAND2X0 U15042 ( .IN1(n14292), .IN2(n14314), .QN(n14296) );
  NAND2X0 U15043 ( .IN1(n14315), .IN2(n14316), .QN(n14314) );
  NAND2X0 U15044 ( .IN1(g5897), .IN2(g6031), .QN(n14316) );
  NAND2X0 U15045 ( .IN1(g5889), .IN2(g13068), .QN(n14315) );
  NAND3X0 U15046 ( .IN1(n11411), .IN2(g17819), .IN3(test_so28), .QN(n14295) );
  NAND3X0 U15047 ( .IN1(g14673), .IN2(g5933), .IN3(n11416), .QN(n14294) );
  NAND3X0 U15048 ( .IN1(n14317), .IN2(n14318), .IN3(n14319), .QN(g28096) );
  NAND2X0 U15049 ( .IN1(n11436), .IN2(g4821), .QN(n14319) );
  NAND2X0 U15050 ( .IN1(n9460), .IN2(g5619), .QN(n14318) );
  NAND3X0 U15051 ( .IN1(n11425), .IN2(n13698), .IN3(n9339), .QN(n14317) );
  NAND2X0 U15052 ( .IN1(n14320), .IN2(n14321), .QN(n13698) );
  NAND2X0 U15053 ( .IN1(n5529), .IN2(n14322), .QN(n14321) );
  NAND4X0 U15054 ( .IN1(n14323), .IN2(n14324), .IN3(n14325), .IN4(n14326), 
        .QN(n14322) );
  NOR3X0 U15055 ( .IN1(n14327), .IN2(n14328), .IN3(n14329), .QN(n14326) );
  NOR2X0 U15056 ( .IN1(n5439), .IN2(n14330), .QN(n14329) );
  NOR2X0 U15057 ( .IN1(n14331), .IN2(n14332), .QN(n14330) );
  NOR2X0 U15058 ( .IN1(n8605), .IN2(n14333), .QN(n14331) );
  NOR2X0 U15059 ( .IN1(n14334), .IN2(g12300), .QN(n14328) );
  NOR2X0 U15060 ( .IN1(n14335), .IN2(n14336), .QN(n14327) );
  NOR2X0 U15061 ( .IN1(n14337), .IN2(n14338), .QN(n14335) );
  NOR2X0 U15062 ( .IN1(n8690), .IN2(n8689), .QN(n14338) );
  NOR2X0 U15063 ( .IN1(n8688), .IN2(n8687), .QN(n14337) );
  NAND2X0 U15064 ( .IN1(n11427), .IN2(n14339), .QN(n14325) );
  NAND2X0 U15065 ( .IN1(n14340), .IN2(n14341), .QN(n14339) );
  INVX0 U15066 ( .INP(n14342), .ZN(n14341) );
  NOR2X0 U15067 ( .IN1(n8658), .IN2(n8659), .QN(n14342) );
  NAND2X0 U15068 ( .IN1(test_so6), .IN2(g17604), .QN(n14340) );
  NAND3X0 U15069 ( .IN1(g14635), .IN2(g5595), .IN3(n14343), .QN(n14324) );
  NAND3X0 U15070 ( .IN1(g17813), .IN2(g5579), .IN3(n10594), .QN(n14323) );
  NAND2X0 U15071 ( .IN1(n14344), .IN2(g5689), .QN(n14320) );
  NAND4X0 U15072 ( .IN1(n14345), .IN2(n14346), .IN3(n14347), .IN4(n14348), 
        .QN(n14344) );
  INVX0 U15073 ( .INP(n14349), .ZN(n14348) );
  NAND3X0 U15074 ( .IN1(n14350), .IN2(n14351), .IN3(n14352), .QN(n14349) );
  NAND2X0 U15075 ( .IN1(g12300), .IN2(n14353), .QN(n14352) );
  NAND2X0 U15076 ( .IN1(n14354), .IN2(n14334), .QN(n14353) );
  INVX0 U15077 ( .INP(n14355), .ZN(n14334) );
  NAND3X0 U15078 ( .IN1(n14356), .IN2(n14357), .IN3(n14358), .QN(n14355) );
  NAND3X0 U15079 ( .IN1(n10594), .IN2(g17711), .IN3(test_so5), .QN(n14358) );
  NAND3X0 U15080 ( .IN1(g17580), .IN2(g5607), .IN3(n14343), .QN(n14357) );
  NAND3X0 U15081 ( .IN1(g14694), .IN2(g5575), .IN3(n11432), .QN(n14356) );
  NAND2X0 U15082 ( .IN1(g5547), .IN2(n11427), .QN(n14354) );
  NAND2X0 U15083 ( .IN1(n14332), .IN2(n5439), .QN(n14351) );
  NAND3X0 U15084 ( .IN1(n14359), .IN2(n14360), .IN3(n14361), .QN(n14332) );
  NAND3X0 U15085 ( .IN1(g5615), .IN2(g17580), .IN3(n11432), .QN(n14361) );
  NAND3X0 U15086 ( .IN1(g5599), .IN2(g17711), .IN3(n11427), .QN(n14360) );
  NAND3X0 U15087 ( .IN1(g14694), .IN2(g5583), .IN3(n14343), .QN(n14359) );
  INVX0 U15088 ( .INP(n14362), .ZN(n14350) );
  NOR2X0 U15089 ( .IN1(n14363), .IN2(n14333), .QN(n14362) );
  INVX0 U15090 ( .INP(n10594), .ZN(n14333) );
  NOR2X0 U15091 ( .IN1(n14364), .IN2(n14365), .QN(n14363) );
  NOR2X0 U15092 ( .IN1(n8658), .IN2(n8481), .QN(n14365) );
  NOR2X0 U15093 ( .IN1(n8660), .IN2(n8480), .QN(n14364) );
  NAND2X0 U15094 ( .IN1(n14343), .IN2(n14366), .QN(n14347) );
  NAND2X0 U15095 ( .IN1(n14367), .IN2(n14368), .QN(n14366) );
  NAND2X0 U15096 ( .IN1(g5551), .IN2(g5685), .QN(n14368) );
  NAND2X0 U15097 ( .IN1(g5543), .IN2(g13049), .QN(n14367) );
  NAND3X0 U15098 ( .IN1(g5571), .IN2(g17813), .IN3(n11427), .QN(n14346) );
  NAND3X0 U15099 ( .IN1(g14635), .IN2(g5587), .IN3(n11432), .QN(n14345) );
  NAND3X0 U15100 ( .IN1(n14369), .IN2(n14370), .IN3(n14371), .QN(g28093) );
  NAND2X0 U15101 ( .IN1(n11448), .IN2(g29220), .QN(n14371) );
  NAND2X0 U15102 ( .IN1(n9460), .IN2(g5272), .QN(n14370) );
  NAND3X0 U15103 ( .IN1(n13732), .IN2(g33959), .IN3(n9339), .QN(n14369) );
  NAND2X0 U15104 ( .IN1(n14372), .IN2(n14373), .QN(n13732) );
  NAND2X0 U15105 ( .IN1(test_so10), .IN2(n14374), .QN(n14373) );
  NAND4X0 U15106 ( .IN1(n14375), .IN2(n14376), .IN3(n14377), .IN4(n14378), 
        .QN(n14374) );
  NOR3X0 U15107 ( .IN1(n14379), .IN2(n14380), .IN3(n14381), .QN(n14378) );
  NOR2X0 U15108 ( .IN1(n5438), .IN2(n14382), .QN(n14381) );
  NOR2X0 U15109 ( .IN1(n14383), .IN2(n14384), .QN(n14382) );
  NOR2X0 U15110 ( .IN1(n8497), .IN2(n14385), .QN(n14383) );
  INVX0 U15111 ( .INP(n14386), .ZN(n14380) );
  NAND2X0 U15112 ( .IN1(n14387), .IN2(n5438), .QN(n14386) );
  NOR2X0 U15113 ( .IN1(n14388), .IN2(n14389), .QN(n14379) );
  NOR2X0 U15114 ( .IN1(n14390), .IN2(n14391), .QN(n14388) );
  NOR2X0 U15115 ( .IN1(n8648), .IN2(n8495), .QN(n14391) );
  NOR2X0 U15116 ( .IN1(n8650), .IN2(n8494), .QN(n14390) );
  NAND2X0 U15117 ( .IN1(n9676), .IN2(n14392), .QN(n14377) );
  NAND2X0 U15118 ( .IN1(n14393), .IN2(n14394), .QN(n14392) );
  NAND2X0 U15119 ( .IN1(g5339), .IN2(g5204), .QN(n14394) );
  NAND2X0 U15120 ( .IN1(g13039), .IN2(g5196), .QN(n14393) );
  NAND3X0 U15121 ( .IN1(g14597), .IN2(g5240), .IN3(n9675), .QN(n14376) );
  NAND3X0 U15122 ( .IN1(g5224), .IN2(g17787), .IN3(n9677), .QN(n14375) );
  NAND2X0 U15123 ( .IN1(n14395), .IN2(n8888), .QN(n14372) );
  NAND4X0 U15124 ( .IN1(n14396), .IN2(n14397), .IN3(n14398), .IN4(n14399), 
        .QN(n14395) );
  NOR3X0 U15125 ( .IN1(n14400), .IN2(n14401), .IN3(n14402), .QN(n14399) );
  NOR2X0 U15126 ( .IN1(n5438), .IN2(n14403), .QN(n14402) );
  NOR2X0 U15127 ( .IN1(n14404), .IN2(n14387), .QN(n14403) );
  NAND3X0 U15128 ( .IN1(n14405), .IN2(n14406), .IN3(n14407), .QN(n14387) );
  NAND3X0 U15129 ( .IN1(g5252), .IN2(g17674), .IN3(n9677), .QN(n14407) );
  NAND3X0 U15130 ( .IN1(g5268), .IN2(g17519), .IN3(n9675), .QN(n14406) );
  NAND3X0 U15131 ( .IN1(g14662), .IN2(g5236), .IN3(n9676), .QN(n14405) );
  NOR2X0 U15132 ( .IN1(n8600), .IN2(n14389), .QN(n14404) );
  INVX0 U15133 ( .INP(g31860), .ZN(n14389) );
  INVX0 U15134 ( .INP(n14408), .ZN(n14401) );
  NAND2X0 U15135 ( .IN1(n14384), .IN2(n5438), .QN(n14408) );
  NAND3X0 U15136 ( .IN1(n14409), .IN2(n14410), .IN3(n14411), .QN(n14384) );
  NAND3X0 U15137 ( .IN1(g17674), .IN2(g5244), .IN3(g31860), .QN(n14411) );
  NAND3X0 U15138 ( .IN1(n9675), .IN2(g14662), .IN3(test_so82), .QN(n14410) );
  NAND3X0 U15139 ( .IN1(g17519), .IN2(g5260), .IN3(n9676), .QN(n14409) );
  NOR2X0 U15140 ( .IN1(n14412), .IN2(n14385), .QN(n14400) );
  INVX0 U15141 ( .INP(n9677), .ZN(n14385) );
  NOR2X0 U15142 ( .IN1(g5297), .IN2(n5393), .QN(n9677) );
  NOR2X0 U15143 ( .IN1(n14413), .IN2(n14414), .QN(n14412) );
  NOR2X0 U15144 ( .IN1(n8651), .IN2(n8650), .QN(n14414) );
  NOR2X0 U15145 ( .IN1(n8649), .IN2(n8648), .QN(n14413) );
  NAND2X0 U15146 ( .IN1(n9675), .IN2(n14415), .QN(n14398) );
  NAND2X0 U15147 ( .IN1(n14416), .IN2(n14417), .QN(n14415) );
  NAND2X0 U15148 ( .IN1(g5220), .IN2(g5339), .QN(n14417) );
  NAND2X0 U15149 ( .IN1(g5208), .IN2(g13039), .QN(n14416) );
  NOR2X0 U15150 ( .IN1(g5357), .IN2(n5588), .QN(n9675) );
  NAND3X0 U15151 ( .IN1(g14597), .IN2(g5248), .IN3(n9676), .QN(n14397) );
  NOR2X0 U15152 ( .IN1(g5297), .IN2(g5357), .QN(n9676) );
  NAND3X0 U15153 ( .IN1(g31860), .IN2(g17787), .IN3(g5232), .QN(n14396) );
  NOR2X0 U15154 ( .IN1(n5393), .IN2(n5588), .QN(g31860) );
  NAND2X0 U15155 ( .IN1(n14418), .IN2(n14419), .QN(g28092) );
  NAND2X0 U15156 ( .IN1(n9460), .IN2(g5057), .QN(n14419) );
  NAND2X0 U15157 ( .IN1(n12385), .IN2(n9380), .QN(n14418) );
  NAND2X0 U15158 ( .IN1(n14420), .IN2(n14421), .QN(n12385) );
  NOR3X0 U15159 ( .IN1(n5615), .IN2(n8773), .IN3(g5046), .QN(n14420) );
  NAND2X0 U15160 ( .IN1(n14422), .IN2(n14423), .QN(g28091) );
  NAND2X0 U15161 ( .IN1(n9460), .IN2(g5069), .QN(n14423) );
  NAND2X0 U15162 ( .IN1(n12384), .IN2(n9380), .QN(n14422) );
  NAND2X0 U15163 ( .IN1(n14424), .IN2(n14425), .QN(n12384) );
  INVX0 U15164 ( .INP(n14421), .ZN(n14425) );
  NOR2X0 U15165 ( .IN1(n14426), .IN2(n14427), .QN(n14421) );
  INVX0 U15166 ( .INP(n14428), .ZN(n14427) );
  NAND2X0 U15167 ( .IN1(g84), .IN2(g5041), .QN(n14428) );
  NOR2X0 U15168 ( .IN1(g84), .IN2(n5607), .QN(n14426) );
  NOR3X0 U15169 ( .IN1(n5578), .IN2(n8775), .IN3(g5057), .QN(n14424) );
  NAND2X0 U15170 ( .IN1(n14429), .IN2(n14430), .QN(g28090) );
  NAND3X0 U15171 ( .IN1(n14431), .IN2(n9313), .IN3(n10639), .QN(n14430) );
  NOR2X0 U15172 ( .IN1(n9741), .IN2(n9763), .QN(n10639) );
  INVX0 U15173 ( .INP(n9758), .ZN(n9763) );
  NAND2X0 U15174 ( .IN1(n5770), .IN2(n14432), .QN(n14431) );
  NAND2X0 U15175 ( .IN1(n11465), .IN2(n14433), .QN(n14432) );
  NAND4X0 U15176 ( .IN1(n14434), .IN2(n14435), .IN3(n14436), .IN4(n14437), 
        .QN(n14433) );
  NAND2X0 U15177 ( .IN1(n11472), .IN2(g4045), .QN(n14437) );
  NAND2X0 U15178 ( .IN1(n8587), .IN2(n14438), .QN(n14436) );
  NAND2X0 U15179 ( .IN1(n10582), .IN2(g4049), .QN(n14435) );
  NAND2X0 U15180 ( .IN1(n8586), .IN2(n11467), .QN(n14434) );
  NAND2X0 U15181 ( .IN1(n11476), .IN2(g4961), .QN(n14429) );
  NAND2X0 U15182 ( .IN1(n14439), .IN2(n14440), .QN(g28089) );
  NAND3X0 U15183 ( .IN1(n14441), .IN2(n9313), .IN3(n10646), .QN(n14440) );
  NOR2X0 U15184 ( .IN1(n9741), .IN2(n9764), .QN(n10646) );
  INVX0 U15185 ( .INP(n9759), .ZN(n9764) );
  NAND2X0 U15186 ( .IN1(n5772), .IN2(n14442), .QN(n14441) );
  NAND2X0 U15187 ( .IN1(n11481), .IN2(n14443), .QN(n14442) );
  NAND4X0 U15188 ( .IN1(n14444), .IN2(n14445), .IN3(n14446), .IN4(n14447), 
        .QN(n14443) );
  NAND2X0 U15189 ( .IN1(n11488), .IN2(g3694), .QN(n14447) );
  NAND2X0 U15190 ( .IN1(n8583), .IN2(n14448), .QN(n14446) );
  NAND2X0 U15191 ( .IN1(n10587), .IN2(g3698), .QN(n14445) );
  NAND2X0 U15192 ( .IN1(n8582), .IN2(n11483), .QN(n14444) );
  NAND2X0 U15193 ( .IN1(n11492), .IN2(g4950), .QN(n14439) );
  NAND2X0 U15194 ( .IN1(n14449), .IN2(n14450), .QN(g28088) );
  NAND3X0 U15195 ( .IN1(n14451), .IN2(n9313), .IN3(n10654), .QN(n14450) );
  INVX0 U15196 ( .INP(n10651), .ZN(n10654) );
  NAND2X0 U15197 ( .IN1(n14452), .IN2(n9756), .QN(n10651) );
  NAND2X0 U15198 ( .IN1(n5776), .IN2(n14453), .QN(n14451) );
  NAND2X0 U15199 ( .IN1(n11501), .IN2(n14454), .QN(n14453) );
  NAND4X0 U15200 ( .IN1(n14455), .IN2(n14456), .IN3(n14457), .IN4(n14458), 
        .QN(n14454) );
  NAND2X0 U15201 ( .IN1(n14459), .IN2(g3343), .QN(n14458) );
  NAND2X0 U15202 ( .IN1(n8578), .IN2(n14460), .QN(n14457) );
  NAND2X0 U15203 ( .IN1(n10595), .IN2(g3347), .QN(n14456) );
  NAND2X0 U15204 ( .IN1(n8577), .IN2(n14461), .QN(n14455) );
  NAND2X0 U15205 ( .IN1(n11507), .IN2(g4939), .QN(n14449) );
  NAND2X0 U15206 ( .IN1(n14462), .IN2(n14463), .QN(g28087) );
  NAND2X0 U15207 ( .IN1(n14464), .IN2(n10251), .QN(n14463) );
  INVX0 U15208 ( .INP(n10662), .ZN(n10251) );
  NAND2X0 U15209 ( .IN1(n14452), .IN2(n9757), .QN(n10662) );
  INVX0 U15210 ( .INP(n9741), .ZN(n14452) );
  NAND3X0 U15211 ( .IN1(g4966), .IN2(n8863), .IN3(g4983), .QN(n9741) );
  NOR2X0 U15212 ( .IN1(n9417), .IN2(n14465), .QN(n14464) );
  NOR2X0 U15213 ( .IN1(n4689), .IN2(g4894), .QN(n14465) );
  NAND2X0 U15214 ( .IN1(n11388), .IN2(g4894), .QN(n14462) );
  NOR2X0 U15215 ( .IN1(n11381), .IN2(n9400), .QN(n11388) );
  INVX0 U15216 ( .INP(n8850), .ZN(n11381) );
  NAND2X0 U15217 ( .IN1(g4836), .IN2(n14466), .QN(n8850) );
  NAND3X0 U15218 ( .IN1(n14467), .IN2(g4888), .IN3(n9756), .QN(n14466) );
  NOR2X0 U15219 ( .IN1(g4899), .IN2(g4975), .QN(n9756) );
  NAND2X0 U15220 ( .IN1(n14468), .IN2(n14469), .QN(g28086) );
  NAND3X0 U15221 ( .IN1(n14470), .IN2(n9313), .IN3(n10671), .QN(n14469) );
  NOR2X0 U15222 ( .IN1(n9708), .IN2(n9730), .QN(n10671) );
  INVX0 U15223 ( .INP(n9723), .ZN(n9730) );
  NAND2X0 U15224 ( .IN1(n5769), .IN2(n14471), .QN(n14470) );
  NAND2X0 U15225 ( .IN1(n11393), .IN2(n14472), .QN(n14471) );
  NAND4X0 U15226 ( .IN1(n14473), .IN2(n14474), .IN3(n14475), .IN4(n14476), 
        .QN(n14472) );
  NAND2X0 U15227 ( .IN1(n10581), .IN2(g6390), .QN(n14476) );
  NOR2X0 U15228 ( .IN1(n5396), .IN2(n5592), .QN(n10581) );
  NAND2X0 U15229 ( .IN1(n8579), .IN2(n11395), .QN(n14475) );
  INVX0 U15230 ( .INP(n14231), .ZN(n11395) );
  NAND2X0 U15231 ( .IN1(n5592), .IN2(g6395), .QN(n14231) );
  INVX0 U15232 ( .INP(n14477), .ZN(n14474) );
  NOR2X0 U15233 ( .IN1(n14260), .IN2(n8580), .QN(n14477) );
  INVX0 U15234 ( .INP(n11400), .ZN(n14260) );
  NOR2X0 U15235 ( .IN1(g6395), .IN2(n5592), .QN(n11400) );
  NAND2X0 U15236 ( .IN1(n8580), .IN2(n14238), .QN(n14473) );
  NOR2X0 U15237 ( .IN1(g6395), .IN2(g6336), .QN(n14238) );
  NAND2X0 U15238 ( .IN1(n11404), .IN2(g4771), .QN(n14468) );
  NOR2X0 U15239 ( .IN1(n11393), .IN2(n9400), .QN(n11404) );
  INVX0 U15240 ( .INP(n11399), .ZN(n11393) );
  NAND2X0 U15241 ( .IN1(g4688), .IN2(n14478), .QN(n11399) );
  NAND3X0 U15242 ( .IN1(n14479), .IN2(g4765), .IN3(n9725), .QN(n14478) );
  NAND2X0 U15243 ( .IN1(n14480), .IN2(n14481), .QN(g28085) );
  NAND3X0 U15244 ( .IN1(n14482), .IN2(n9313), .IN3(n10678), .QN(n14481) );
  NOR2X0 U15245 ( .IN1(n9708), .IN2(n9731), .QN(n10678) );
  INVX0 U15246 ( .INP(n9724), .ZN(n9731) );
  NAND2X0 U15247 ( .IN1(n5775), .IN2(n14483), .QN(n14482) );
  NAND2X0 U15248 ( .IN1(n11409), .IN2(n14484), .QN(n14483) );
  NAND4X0 U15249 ( .IN1(n14485), .IN2(n14486), .IN3(n14487), .IN4(n14488), 
        .QN(n14484) );
  NAND2X0 U15250 ( .IN1(n11411), .IN2(n8887), .QN(n14488) );
  NOR2X0 U15251 ( .IN1(g5990), .IN2(n8866), .QN(n11411) );
  NAND2X0 U15252 ( .IN1(test_so50), .IN2(n10586), .QN(n14487) );
  NOR2X0 U15253 ( .IN1(n8866), .IN2(n5589), .QN(n10586) );
  INVX0 U15254 ( .INP(n14489), .ZN(n14486) );
  NOR2X0 U15255 ( .IN1(n14286), .IN2(n8581), .QN(n14489) );
  INVX0 U15256 ( .INP(n11416), .ZN(n14286) );
  NOR2X0 U15257 ( .IN1(n5589), .IN2(test_so57), .QN(n11416) );
  NAND2X0 U15258 ( .IN1(n8581), .IN2(n14292), .QN(n14485) );
  NOR2X0 U15259 ( .IN1(g5990), .IN2(test_so57), .QN(n14292) );
  NAND2X0 U15260 ( .IN1(n11420), .IN2(g4760), .QN(n14480) );
  NOR2X0 U15261 ( .IN1(n11409), .IN2(n9401), .QN(n11420) );
  INVX0 U15262 ( .INP(n11415), .ZN(n11409) );
  NAND2X0 U15263 ( .IN1(g4681), .IN2(n14490), .QN(n11415) );
  NAND3X0 U15264 ( .IN1(n14479), .IN2(g4754), .IN3(n9723), .QN(n14490) );
  NOR2X0 U15265 ( .IN1(g4785), .IN2(n5518), .QN(n9723) );
  NAND2X0 U15266 ( .IN1(n14491), .IN2(n14492), .QN(g28084) );
  NAND3X0 U15267 ( .IN1(n14493), .IN2(n9313), .IN3(n10686), .QN(n14492) );
  INVX0 U15268 ( .INP(n10683), .ZN(n10686) );
  NAND2X0 U15269 ( .IN1(n14494), .IN2(n9726), .QN(n10683) );
  NAND2X0 U15270 ( .IN1(n8906), .IN2(n14495), .QN(n14493) );
  NAND2X0 U15271 ( .IN1(n11425), .IN2(n14496), .QN(n14495) );
  NAND4X0 U15272 ( .IN1(n14497), .IN2(n14498), .IN3(n14499), .IN4(n14500), 
        .QN(n14496) );
  NAND2X0 U15273 ( .IN1(n10594), .IN2(g5698), .QN(n14500) );
  NOR2X0 U15274 ( .IN1(n5397), .IN2(n5593), .QN(n10594) );
  NAND2X0 U15275 ( .IN1(n8584), .IN2(n11427), .QN(n14499) );
  NOR2X0 U15276 ( .IN1(g5644), .IN2(n5397), .QN(n11427) );
  INVX0 U15277 ( .INP(n14501), .ZN(n14498) );
  NOR2X0 U15278 ( .IN1(n14336), .IN2(n8585), .QN(n14501) );
  INVX0 U15279 ( .INP(n11432), .ZN(n14336) );
  NOR2X0 U15280 ( .IN1(g5703), .IN2(n5593), .QN(n11432) );
  NAND2X0 U15281 ( .IN1(n8585), .IN2(n14343), .QN(n14497) );
  NOR2X0 U15282 ( .IN1(g5703), .IN2(g5644), .QN(n14343) );
  NAND2X0 U15283 ( .IN1(n11436), .IN2(test_so18), .QN(n14491) );
  NOR2X0 U15284 ( .IN1(n11425), .IN2(n9401), .QN(n11436) );
  INVX0 U15285 ( .INP(n11431), .ZN(n11425) );
  NAND2X0 U15286 ( .IN1(g4674), .IN2(n14502), .QN(n11431) );
  NAND3X0 U15287 ( .IN1(n14479), .IN2(g4743), .IN3(n9724), .QN(n14502) );
  NOR2X0 U15288 ( .IN1(g4709), .IN2(n5361), .QN(n9724) );
  NAND2X0 U15289 ( .IN1(n14503), .IN2(n14504), .QN(g28083) );
  NAND2X0 U15290 ( .IN1(n14505), .IN2(n10254), .QN(n14504) );
  INVX0 U15291 ( .INP(n10694), .ZN(n10254) );
  NAND2X0 U15292 ( .IN1(n14494), .IN2(n9725), .QN(n10694) );
  NOR2X0 U15293 ( .IN1(n5361), .IN2(n5518), .QN(n9725) );
  INVX0 U15294 ( .INP(n9708), .ZN(n14494) );
  NAND3X0 U15295 ( .IN1(g4776), .IN2(n8862), .IN3(g4793), .QN(n9708) );
  NOR2X0 U15296 ( .IN1(n9416), .IN2(n14506), .QN(n14505) );
  NOR2X0 U15297 ( .IN1(n4708), .IN2(g4704), .QN(n14506) );
  NAND2X0 U15298 ( .IN1(n11448), .IN2(g4704), .QN(n14503) );
  NOR2X0 U15299 ( .IN1(g33959), .IN2(n9401), .QN(n11448) );
  INVX0 U15300 ( .INP(n8845), .ZN(g33959) );
  NAND2X0 U15301 ( .IN1(g4646), .IN2(n14507), .QN(n8845) );
  NAND3X0 U15302 ( .IN1(n14479), .IN2(g4698), .IN3(n9726), .QN(n14507) );
  NOR2X0 U15303 ( .IN1(g4709), .IN2(g4785), .QN(n9726) );
  INVX0 U15304 ( .INP(n14508), .ZN(n14479) );
  NAND4X0 U15305 ( .IN1(n5368), .IN2(n10823), .IN3(g4776), .IN4(n8862), .QN(
        n14508) );
  NOR3X0 U15306 ( .IN1(n8830), .IN2(n8831), .IN3(n8881), .QN(n10823) );
  NAND2X0 U15307 ( .IN1(n14509), .IN2(n14510), .QN(g28082) );
  NAND2X0 U15308 ( .IN1(n14511), .IN2(g4521), .QN(n14510) );
  NAND2X0 U15309 ( .IN1(n14512), .IN2(n9380), .QN(n14511) );
  NAND2X0 U15310 ( .IN1(n14513), .IN2(n14514), .QN(n14512) );
  NAND2X0 U15311 ( .IN1(n8725), .IN2(n14515), .QN(n14514) );
  NAND2X0 U15312 ( .IN1(n10832), .IN2(g4527), .QN(n14513) );
  NAND3X0 U15313 ( .IN1(n10137), .IN2(n9316), .IN3(n5752), .QN(n14509) );
  NAND3X0 U15314 ( .IN1(n14516), .IN2(n14517), .IN3(n14518), .QN(g28074) );
  NAND2X0 U15315 ( .IN1(n9460), .IN2(g4119), .QN(n14518) );
  NAND3X0 U15316 ( .IN1(n9353), .IN2(g4122), .IN3(n14519), .QN(n14517) );
  INVX0 U15317 ( .INP(n4714), .ZN(n14519) );
  NAND2X0 U15318 ( .IN1(n4714), .IN2(n4721), .QN(n14516) );
  NAND3X0 U15319 ( .IN1(n14520), .IN2(n14521), .IN3(n14522), .QN(g28073) );
  NAND2X0 U15320 ( .IN1(n14523), .IN2(n4721), .QN(n14522) );
  INVX0 U15321 ( .INP(n14524), .ZN(n14523) );
  NAND3X0 U15322 ( .IN1(n14524), .IN2(g4119), .IN3(n9339), .QN(n14521) );
  NAND3X0 U15323 ( .IN1(n5416), .IN2(g4057), .IN3(n4722), .QN(n14524) );
  NAND2X0 U15324 ( .IN1(n9459), .IN2(g4116), .QN(n14520) );
  NAND3X0 U15325 ( .IN1(n14525), .IN2(n14526), .IN3(n14527), .QN(g28072) );
  NAND2X0 U15326 ( .IN1(n14528), .IN2(n4721), .QN(n14527) );
  INVX0 U15327 ( .INP(n14529), .ZN(n14528) );
  NAND3X0 U15328 ( .IN1(n14529), .IN2(g4116), .IN3(n9339), .QN(n14526) );
  NAND3X0 U15329 ( .IN1(n5711), .IN2(g4064), .IN3(n4722), .QN(n14529) );
  INVX0 U15330 ( .INP(n14530), .ZN(n4722) );
  NAND2X0 U15331 ( .IN1(n9459), .IN2(g4112), .QN(n14525) );
  NAND2X0 U15332 ( .IN1(n14531), .IN2(n14532), .QN(g28071) );
  NAND2X0 U15333 ( .IN1(n14533), .IN2(g4112), .QN(n14532) );
  INVX0 U15334 ( .INP(n14534), .ZN(n14531) );
  NOR2X0 U15335 ( .IN1(n14533), .IN2(n8726), .QN(n14534) );
  NOR2X0 U15336 ( .IN1(n14535), .IN2(n9402), .QN(n14533) );
  NOR3X0 U15337 ( .IN1(g4057), .IN2(g4064), .IN3(n14530), .QN(n14535) );
  NAND4X0 U15338 ( .IN1(n8446), .IN2(n5612), .IN3(n14536), .IN4(n5350), .QN(
        n14530) );
  NOR2X0 U15339 ( .IN1(test_so11), .IN2(n10571), .QN(n14536) );
  INVX0 U15340 ( .INP(n11360), .ZN(n10571) );
  NOR2X0 U15341 ( .IN1(g4093), .IN2(g4087), .QN(n11360) );
  NAND4X0 U15342 ( .IN1(n14537), .IN2(n12032), .IN3(n14538), .IN4(n14539), 
        .QN(g28070) );
  NAND3X0 U15343 ( .IN1(test_so11), .IN2(n14540), .IN3(n9339), .QN(n14539) );
  NAND2X0 U15344 ( .IN1(n9459), .IN2(g4082), .QN(n14538) );
  NAND2X0 U15345 ( .IN1(n13736), .IN2(n8878), .QN(n14537) );
  INVX0 U15346 ( .INP(n14540), .ZN(n13736) );
  NAND3X0 U15347 ( .IN1(n14541), .IN2(n14542), .IN3(n14543), .QN(g28069) );
  NAND2X0 U15348 ( .IN1(n11476), .IN2(g4035), .QN(n14543) );
  NOR2X0 U15349 ( .IN1(n11465), .IN2(n9403), .QN(n11476) );
  NAND2X0 U15350 ( .IN1(n9459), .IN2(g3965), .QN(n14542) );
  NAND3X0 U15351 ( .IN1(n11465), .IN2(n13769), .IN3(n9338), .QN(n14541) );
  NAND2X0 U15352 ( .IN1(n14544), .IN2(n14545), .QN(n13769) );
  NAND2X0 U15353 ( .IN1(n5530), .IN2(n14546), .QN(n14545) );
  NAND4X0 U15354 ( .IN1(n14547), .IN2(n14548), .IN3(n14549), .IN4(n14550), 
        .QN(n14546) );
  NOR3X0 U15355 ( .IN1(n14551), .IN2(n14552), .IN3(n14553), .QN(n14550) );
  NOR2X0 U15356 ( .IN1(n5435), .IN2(n14554), .QN(n14553) );
  NOR2X0 U15357 ( .IN1(n14555), .IN2(n14556), .QN(n14554) );
  NOR2X0 U15358 ( .IN1(n8608), .IN2(n14557), .QN(n14555) );
  INVX0 U15359 ( .INP(n14558), .ZN(n14552) );
  NAND2X0 U15360 ( .IN1(n14559), .IN2(n5435), .QN(n14558) );
  NOR2X0 U15361 ( .IN1(n14560), .IN2(n14561), .QN(n14551) );
  NOR2X0 U15362 ( .IN1(n14562), .IN2(n14563), .QN(n14560) );
  NOR2X0 U15363 ( .IN1(n8665), .IN2(n8664), .QN(n14563) );
  NOR2X0 U15364 ( .IN1(n8663), .IN2(n8662), .QN(n14562) );
  NAND2X0 U15365 ( .IN1(n11472), .IN2(n14564), .QN(n14549) );
  NAND2X0 U15366 ( .IN1(n14565), .IN2(n14566), .QN(n14564) );
  NAND2X0 U15367 ( .IN1(g4031), .IN2(g3913), .QN(n14566) );
  NAND2X0 U15368 ( .IN1(g14518), .IN2(g3901), .QN(n14565) );
  NAND3X0 U15369 ( .IN1(g13906), .IN2(g3941), .IN3(n14438), .QN(n14548) );
  NAND3X0 U15370 ( .IN1(g16955), .IN2(g3925), .IN3(n10582), .QN(n14547) );
  NAND2X0 U15371 ( .IN1(n14567), .IN2(g4040), .QN(n14544) );
  NAND4X0 U15372 ( .IN1(n14568), .IN2(n14569), .IN3(n14570), .IN4(n14571), 
        .QN(n14567) );
  NOR3X0 U15373 ( .IN1(n14572), .IN2(n14573), .IN3(n14574), .QN(n14571) );
  NOR2X0 U15374 ( .IN1(n5435), .IN2(n14575), .QN(n14574) );
  NOR2X0 U15375 ( .IN1(n14576), .IN2(n14559), .QN(n14575) );
  NAND3X0 U15376 ( .IN1(n14577), .IN2(n14578), .IN3(n14579), .QN(n14559) );
  NAND3X0 U15377 ( .IN1(g13966), .IN2(g3921), .IN3(n11472), .QN(n14579) );
  NAND3X0 U15378 ( .IN1(g16659), .IN2(g3953), .IN3(n14438), .QN(n14578) );
  NAND3X0 U15379 ( .IN1(g16775), .IN2(g3937), .IN3(n10582), .QN(n14577) );
  NOR2X0 U15380 ( .IN1(n8502), .IN2(n14561), .QN(n14576) );
  INVX0 U15381 ( .INP(n14580), .ZN(n14573) );
  NAND2X0 U15382 ( .IN1(n14556), .IN2(n5435), .QN(n14580) );
  NAND3X0 U15383 ( .IN1(n14581), .IN2(n14582), .IN3(n14583), .QN(n14556) );
  NAND3X0 U15384 ( .IN1(g3945), .IN2(g16775), .IN3(n11467), .QN(n14583) );
  NAND3X0 U15385 ( .IN1(g13966), .IN2(g3929), .IN3(n14438), .QN(n14582) );
  NAND3X0 U15386 ( .IN1(g3961), .IN2(g16659), .IN3(n11472), .QN(n14581) );
  NOR2X0 U15387 ( .IN1(n14584), .IN2(n14557), .QN(n14572) );
  INVX0 U15388 ( .INP(n10582), .ZN(n14557) );
  NOR2X0 U15389 ( .IN1(n5395), .IN2(n5594), .QN(n10582) );
  NOR2X0 U15390 ( .IN1(n14585), .IN2(n14586), .QN(n14584) );
  NOR2X0 U15391 ( .IN1(n8662), .IN2(n8896), .QN(n14586) );
  NOR2X0 U15392 ( .IN1(n8664), .IN2(n8500), .QN(n14585) );
  NAND2X0 U15393 ( .IN1(n14438), .IN2(n14587), .QN(n14570) );
  NAND2X0 U15394 ( .IN1(n14588), .IN2(n14589), .QN(n14587) );
  NAND2X0 U15395 ( .IN1(g3897), .IN2(g4031), .QN(n14589) );
  NAND2X0 U15396 ( .IN1(test_so24), .IN2(g14518), .QN(n14588) );
  NOR2X0 U15397 ( .IN1(g4054), .IN2(g3990), .QN(n14438) );
  NAND3X0 U15398 ( .IN1(g13906), .IN2(g3933), .IN3(n11472), .QN(n14569) );
  NOR2X0 U15399 ( .IN1(g4054), .IN2(n5594), .QN(n11472) );
  NAND3X0 U15400 ( .IN1(g3917), .IN2(g16955), .IN3(n11467), .QN(n14568) );
  INVX0 U15401 ( .INP(n14561), .ZN(n11467) );
  NAND2X0 U15402 ( .IN1(n5594), .IN2(g4054), .QN(n14561) );
  INVX0 U15403 ( .INP(n11471), .ZN(n11465) );
  NAND2X0 U15404 ( .IN1(g4878), .IN2(n14590), .QN(n11471) );
  NAND3X0 U15405 ( .IN1(n14467), .IN2(g4955), .IN3(n9757), .QN(n14590) );
  NOR2X0 U15406 ( .IN1(n5360), .IN2(n5517), .QN(n9757) );
  NAND3X0 U15407 ( .IN1(n14591), .IN2(n14592), .IN3(n14593), .QN(g28066) );
  NAND2X0 U15408 ( .IN1(n11492), .IN2(g3684), .QN(n14593) );
  NOR2X0 U15409 ( .IN1(n11481), .IN2(n9403), .QN(n11492) );
  NAND2X0 U15410 ( .IN1(n9459), .IN2(g3614), .QN(n14592) );
  NAND3X0 U15411 ( .IN1(n11481), .IN2(n13802), .IN3(n9338), .QN(n14591) );
  NAND2X0 U15412 ( .IN1(n14594), .IN2(n14595), .QN(n13802) );
  NAND2X0 U15413 ( .IN1(n5532), .IN2(n14596), .QN(n14595) );
  NAND4X0 U15414 ( .IN1(n14597), .IN2(n14598), .IN3(n14599), .IN4(n14600), 
        .QN(n14596) );
  NOR3X0 U15415 ( .IN1(n14601), .IN2(n14602), .IN3(n14603), .QN(n14600) );
  NOR2X0 U15416 ( .IN1(n5433), .IN2(n14604), .QN(n14603) );
  NOR2X0 U15417 ( .IN1(n14605), .IN2(n14606), .QN(n14604) );
  NOR2X0 U15418 ( .IN1(n8614), .IN2(n14607), .QN(n14605) );
  NOR2X0 U15419 ( .IN1(n14608), .IN2(g11388), .QN(n14602) );
  NOR2X0 U15420 ( .IN1(n14609), .IN2(n14610), .QN(n14601) );
  NOR2X0 U15421 ( .IN1(n14611), .IN2(n14612), .QN(n14609) );
  NOR2X0 U15422 ( .IN1(n8673), .IN2(n8672), .QN(n14612) );
  INVX0 U15423 ( .INP(n14613), .ZN(n14611) );
  NAND2X0 U15424 ( .IN1(g16656), .IN2(g3554), .QN(n14613) );
  NAND2X0 U15425 ( .IN1(n11488), .IN2(n14614), .QN(n14599) );
  NAND2X0 U15426 ( .IN1(n14615), .IN2(n14616), .QN(n14614) );
  NAND2X0 U15427 ( .IN1(g3680), .IN2(g3562), .QN(n14616) );
  NAND2X0 U15428 ( .IN1(g14451), .IN2(g3550), .QN(n14615) );
  NAND3X0 U15429 ( .IN1(test_so26), .IN2(g3590), .IN3(n14448), .QN(n14598) );
  NAND3X0 U15430 ( .IN1(g16924), .IN2(g3574), .IN3(n10587), .QN(n14597) );
  NAND2X0 U15431 ( .IN1(n14617), .IN2(g3689), .QN(n14594) );
  NAND4X0 U15432 ( .IN1(n14618), .IN2(n14619), .IN3(n14620), .IN4(n14621), 
        .QN(n14617) );
  INVX0 U15433 ( .INP(n14622), .ZN(n14621) );
  NAND3X0 U15434 ( .IN1(n14623), .IN2(n14624), .IN3(n14625), .QN(n14622) );
  NAND2X0 U15435 ( .IN1(g11388), .IN2(n14626), .QN(n14625) );
  NAND2X0 U15436 ( .IN1(n14627), .IN2(n14608), .QN(n14626) );
  INVX0 U15437 ( .INP(n14628), .ZN(n14608) );
  NAND3X0 U15438 ( .IN1(n14629), .IN2(n14630), .IN3(n14631), .QN(n14628) );
  NAND3X0 U15439 ( .IN1(g13926), .IN2(g3570), .IN3(n11488), .QN(n14631) );
  NAND3X0 U15440 ( .IN1(test_so43), .IN2(g16627), .IN3(n14448), .QN(n14630) );
  NAND3X0 U15441 ( .IN1(g16744), .IN2(g3586), .IN3(n10587), .QN(n14629) );
  NAND2X0 U15442 ( .IN1(n11483), .IN2(g3542), .QN(n14627) );
  NAND2X0 U15443 ( .IN1(n14606), .IN2(n5433), .QN(n14624) );
  NAND3X0 U15444 ( .IN1(n14632), .IN2(n14633), .IN3(n14634), .QN(n14606) );
  NAND3X0 U15445 ( .IN1(g3594), .IN2(g16744), .IN3(n11483), .QN(n14634) );
  NAND3X0 U15446 ( .IN1(g13926), .IN2(g3578), .IN3(n14448), .QN(n14633) );
  NAND3X0 U15447 ( .IN1(g3610), .IN2(g16627), .IN3(n11488), .QN(n14632) );
  INVX0 U15448 ( .INP(n14635), .ZN(n14623) );
  NOR2X0 U15449 ( .IN1(n14636), .IN2(n14607), .QN(n14635) );
  INVX0 U15450 ( .INP(n10587), .ZN(n14607) );
  NOR2X0 U15451 ( .IN1(n5399), .IN2(n5591), .QN(n10587) );
  NOR2X0 U15452 ( .IN1(n14637), .IN2(n14638), .QN(n14636) );
  NOR2X0 U15453 ( .IN1(n8672), .IN2(n8488), .QN(n14638) );
  NOR2X0 U15454 ( .IN1(n8674), .IN2(n8487), .QN(n14637) );
  NAND2X0 U15455 ( .IN1(n14448), .IN2(n14639), .QN(n14620) );
  NAND2X0 U15456 ( .IN1(n14640), .IN2(n14641), .QN(n14639) );
  NAND2X0 U15457 ( .IN1(g3546), .IN2(g3680), .QN(n14641) );
  NAND2X0 U15458 ( .IN1(g3538), .IN2(g14451), .QN(n14640) );
  NOR2X0 U15459 ( .IN1(g3703), .IN2(g3639), .QN(n14448) );
  NAND3X0 U15460 ( .IN1(n11488), .IN2(g3582), .IN3(test_so26), .QN(n14619) );
  NOR2X0 U15461 ( .IN1(g3703), .IN2(n5591), .QN(n11488) );
  NAND3X0 U15462 ( .IN1(g3566), .IN2(g16924), .IN3(n11483), .QN(n14618) );
  INVX0 U15463 ( .INP(n14610), .ZN(n11483) );
  NAND2X0 U15464 ( .IN1(n5591), .IN2(g3703), .QN(n14610) );
  INVX0 U15465 ( .INP(n11487), .ZN(n11481) );
  NAND2X0 U15466 ( .IN1(g4871), .IN2(n14642), .QN(n11487) );
  NAND3X0 U15467 ( .IN1(n14467), .IN2(g4944), .IN3(n9758), .QN(n14642) );
  NOR2X0 U15468 ( .IN1(g4975), .IN2(n5517), .QN(n9758) );
  NAND3X0 U15469 ( .IN1(n14643), .IN2(n14644), .IN3(n14645), .QN(g28063) );
  NAND2X0 U15470 ( .IN1(n11507), .IN2(g3333), .QN(n14645) );
  NOR2X0 U15471 ( .IN1(n11501), .IN2(n9404), .QN(n11507) );
  NAND2X0 U15472 ( .IN1(n9459), .IN2(g3263), .QN(n14644) );
  NAND3X0 U15473 ( .IN1(n11501), .IN2(n13836), .IN3(n9338), .QN(n14643) );
  NAND2X0 U15474 ( .IN1(n14646), .IN2(n14647), .QN(n13836) );
  NAND2X0 U15475 ( .IN1(n5527), .IN2(n14648), .QN(n14647) );
  NAND4X0 U15476 ( .IN1(n14649), .IN2(n14650), .IN3(n14651), .IN4(n14652), 
        .QN(n14648) );
  NOR3X0 U15477 ( .IN1(n14653), .IN2(n14654), .IN3(n14655), .QN(n14652) );
  NOR2X0 U15478 ( .IN1(n5436), .IN2(n14656), .QN(n14655) );
  NOR2X0 U15479 ( .IN1(n14657), .IN2(n14658), .QN(n14656) );
  NOR2X0 U15480 ( .IN1(n8598), .IN2(n14659), .QN(n14657) );
  INVX0 U15481 ( .INP(n14660), .ZN(n14654) );
  NAND2X0 U15482 ( .IN1(n14661), .IN2(n5436), .QN(n14660) );
  NOR2X0 U15483 ( .IN1(n14662), .IN2(n11503), .QN(n14653) );
  NOR2X0 U15484 ( .IN1(n14663), .IN2(n14664), .QN(n14662) );
  NOR2X0 U15485 ( .IN1(n8646), .IN2(n8645), .QN(n14664) );
  NOR2X0 U15486 ( .IN1(n8644), .IN2(n8643), .QN(n14663) );
  NAND2X0 U15487 ( .IN1(n14459), .IN2(n14665), .QN(n14651) );
  NAND2X0 U15488 ( .IN1(n14666), .IN2(n14667), .QN(n14665) );
  NAND2X0 U15489 ( .IN1(test_so91), .IN2(g3211), .QN(n14667) );
  NAND2X0 U15490 ( .IN1(g14421), .IN2(g3199), .QN(n14666) );
  NAND3X0 U15491 ( .IN1(g13865), .IN2(g3239), .IN3(n14460), .QN(n14650) );
  NAND3X0 U15492 ( .IN1(g16874), .IN2(g3223), .IN3(n10595), .QN(n14649) );
  NAND2X0 U15493 ( .IN1(n14668), .IN2(g3338), .QN(n14646) );
  NAND4X0 U15494 ( .IN1(n14669), .IN2(n14670), .IN3(n14671), .IN4(n14672), 
        .QN(n14668) );
  NOR3X0 U15495 ( .IN1(n14673), .IN2(n14674), .IN3(n14675), .QN(n14672) );
  NOR2X0 U15496 ( .IN1(n5436), .IN2(n14676), .QN(n14675) );
  NOR2X0 U15497 ( .IN1(n14677), .IN2(n14661), .QN(n14676) );
  NAND3X0 U15498 ( .IN1(n14678), .IN2(n14679), .IN3(n14680), .QN(n14661) );
  NAND3X0 U15499 ( .IN1(g13895), .IN2(g3219), .IN3(n14459), .QN(n14680) );
  NAND3X0 U15500 ( .IN1(g16603), .IN2(g3251), .IN3(n14460), .QN(n14679) );
  NAND3X0 U15501 ( .IN1(g16718), .IN2(g3235), .IN3(n10595), .QN(n14678) );
  NOR2X0 U15502 ( .IN1(n8479), .IN2(n11503), .QN(n14677) );
  INVX0 U15503 ( .INP(n14461), .ZN(n11503) );
  INVX0 U15504 ( .INP(n14681), .ZN(n14674) );
  NAND2X0 U15505 ( .IN1(n14658), .IN2(n5436), .QN(n14681) );
  NAND3X0 U15506 ( .IN1(n14682), .IN2(n14683), .IN3(n14684), .QN(n14658) );
  NAND3X0 U15507 ( .IN1(g3243), .IN2(g16718), .IN3(n14461), .QN(n14684) );
  NAND3X0 U15508 ( .IN1(g13895), .IN2(g3227), .IN3(n14460), .QN(n14683) );
  NAND3X0 U15509 ( .IN1(test_so84), .IN2(g16603), .IN3(n14459), .QN(n14682) );
  NOR2X0 U15510 ( .IN1(n14685), .IN2(n14659), .QN(n14673) );
  INVX0 U15511 ( .INP(n10595), .ZN(n14659) );
  NOR2X0 U15512 ( .IN1(n5400), .IN2(n5604), .QN(n10595) );
  NOR2X0 U15513 ( .IN1(n14686), .IN2(n14687), .QN(n14685) );
  NOR2X0 U15514 ( .IN1(n8643), .IN2(n8477), .QN(n14687) );
  NOR2X0 U15515 ( .IN1(n8645), .IN2(n8476), .QN(n14686) );
  NAND2X0 U15516 ( .IN1(n14460), .IN2(n14688), .QN(n14671) );
  NAND2X0 U15517 ( .IN1(n14689), .IN2(n14690), .QN(n14688) );
  NAND2X0 U15518 ( .IN1(g3187), .IN2(g14421), .QN(n14690) );
  NAND2X0 U15519 ( .IN1(test_so91), .IN2(test_so88), .QN(n14689) );
  NOR2X0 U15520 ( .IN1(g3352), .IN2(g3288), .QN(n14460) );
  NAND3X0 U15521 ( .IN1(g13865), .IN2(g3231), .IN3(n14459), .QN(n14670) );
  INVX0 U15522 ( .INP(n11502), .ZN(n14459) );
  NAND2X0 U15523 ( .IN1(n5604), .IN2(g3288), .QN(n11502) );
  NAND3X0 U15524 ( .IN1(g3215), .IN2(g16874), .IN3(n14461), .QN(n14669) );
  NOR2X0 U15525 ( .IN1(g3288), .IN2(n5604), .QN(n14461) );
  INVX0 U15526 ( .INP(n11498), .ZN(n11501) );
  NAND2X0 U15527 ( .IN1(g4864), .IN2(n14691), .QN(n11498) );
  NAND3X0 U15528 ( .IN1(n14467), .IN2(g4933), .IN3(n9759), .QN(n14691) );
  NOR2X0 U15529 ( .IN1(g4899), .IN2(n5360), .QN(n9759) );
  INVX0 U15530 ( .INP(n14692), .ZN(n14467) );
  NAND4X0 U15531 ( .IN1(n5367), .IN2(n10792), .IN3(g4966), .IN4(n8863), .QN(
        n14692) );
  NOR3X0 U15532 ( .IN1(n8833), .IN2(n8834), .IN3(n8832), .QN(n10792) );
  NAND3X0 U15533 ( .IN1(n14693), .IN2(n9664), .IN3(n14694), .QN(g28060) );
  NAND2X0 U15534 ( .IN1(n14695), .IN2(g2724), .QN(n14694) );
  NAND2X0 U15535 ( .IN1(n14696), .IN2(n9380), .QN(n14695) );
  NAND2X0 U15536 ( .IN1(n13185), .IN2(n13214), .QN(n14696) );
  NAND3X0 U15537 ( .IN1(n9350), .IN2(g2729), .IN3(n13214), .QN(n14693) );
  INVX0 U15538 ( .INP(n13840), .ZN(n13214) );
  NOR2X0 U15539 ( .IN1(n10532), .IN2(n14697), .QN(n13840) );
  NAND2X0 U15540 ( .IN1(g2724), .IN2(g2729), .QN(n10532) );
  NAND3X0 U15541 ( .IN1(n14698), .IN2(n14699), .IN3(n14700), .QN(g28059) );
  NAND2X0 U15542 ( .IN1(n9459), .IN2(g1351), .QN(n14700) );
  NAND3X0 U15543 ( .IN1(n12281), .IN2(n8448), .IN3(n13501), .QN(n14699) );
  NOR2X0 U15544 ( .IN1(n13503), .IN2(n9404), .QN(n12281) );
  NAND4X0 U15545 ( .IN1(n5466), .IN2(n14701), .IN3(n14702), .IN4(n14703), .QN(
        n13503) );
  NAND2X0 U15546 ( .IN1(n14704), .IN2(n5322), .QN(n14703) );
  NAND3X0 U15547 ( .IN1(n14705), .IN2(g1351), .IN3(n14706), .QN(n14702) );
  NAND2X0 U15548 ( .IN1(n4798), .IN2(n14707), .QN(n14698) );
  NAND3X0 U15549 ( .IN1(n14708), .IN2(n14709), .IN3(n14710), .QN(g28058) );
  NAND2X0 U15550 ( .IN1(test_so77), .IN2(n9514), .QN(n14710) );
  NAND3X0 U15551 ( .IN1(n11853), .IN2(n14711), .IN3(g1252), .QN(n14709) );
  INVX0 U15552 ( .INP(n4490), .ZN(n14711) );
  NAND2X0 U15553 ( .IN1(n4490), .IN2(n5554), .QN(n14708) );
  NAND3X0 U15554 ( .IN1(n14712), .IN2(n14713), .IN3(n14714), .QN(g28057) );
  NAND2X0 U15555 ( .IN1(n9458), .IN2(g1008), .QN(n14714) );
  NAND3X0 U15556 ( .IN1(n12294), .IN2(n8449), .IN3(n13538), .QN(n14713) );
  NOR2X0 U15557 ( .IN1(n14715), .IN2(n9405), .QN(n12294) );
  INVX0 U15558 ( .INP(n11861), .ZN(n14715) );
  NOR4X0 U15559 ( .IN1(n14716), .IN2(test_so20), .IN3(n14717), .IN4(n14718), 
        .QN(n11861) );
  NOR2X0 U15560 ( .IN1(n14719), .IN2(n14720), .QN(n14718) );
  NOR2X0 U15561 ( .IN1(n14721), .IN2(g1008), .QN(n14717) );
  NAND2X0 U15562 ( .IN1(n4805), .IN2(n14722), .QN(n14712) );
  NAND3X0 U15563 ( .IN1(n14723), .IN2(n14724), .IN3(n14725), .QN(g28056) );
  NAND2X0 U15564 ( .IN1(n9458), .IN2(g936), .QN(n14725) );
  NAND3X0 U15565 ( .IN1(n11867), .IN2(n14726), .IN3(g907), .QN(n14724) );
  INVX0 U15566 ( .INP(n4514), .ZN(n14726) );
  NAND2X0 U15567 ( .IN1(n4514), .IN2(n5555), .QN(n14723) );
  NAND3X0 U15568 ( .IN1(n14727), .IN2(n14728), .IN3(n14729), .QN(g28055) );
  NAND2X0 U15569 ( .IN1(n9458), .IN2(g822), .QN(n14729) );
  NAND3X0 U15570 ( .IN1(n4518), .IN2(n14730), .IN3(g827), .QN(n14728) );
  INVX0 U15571 ( .INP(n4519), .ZN(n14730) );
  NAND3X0 U15572 ( .IN1(n4519), .IN2(n14104), .IN3(n5728), .QN(n14727) );
  NAND2X0 U15573 ( .IN1(n14731), .IN2(n14732), .QN(g28054) );
  NAND2X0 U15574 ( .IN1(n14733), .IN2(g728), .QN(n14732) );
  NAND2X0 U15575 ( .IN1(n14734), .IN2(g661), .QN(n14731) );
  NAND3X0 U15576 ( .IN1(n14735), .IN2(n14736), .IN3(n14737), .QN(g28053) );
  NAND2X0 U15577 ( .IN1(n9458), .IN2(g681), .QN(n14737) );
  INVX0 U15578 ( .INP(n14738), .ZN(n14736) );
  NAND2X0 U15579 ( .IN1(n14147), .IN2(test_so87), .QN(n14735) );
  NAND2X0 U15580 ( .IN1(n14739), .IN2(n14740), .QN(g28052) );
  NAND2X0 U15581 ( .IN1(n14733), .IN2(g661), .QN(n14740) );
  NAND2X0 U15582 ( .IN1(n14734), .IN2(g718), .QN(n14739) );
  NAND2X0 U15583 ( .IN1(n14741), .IN2(n14742), .QN(g28051) );
  NAND2X0 U15584 ( .IN1(n14733), .IN2(g718), .QN(n14742) );
  NAND2X0 U15585 ( .IN1(n14734), .IN2(g655), .QN(n14741) );
  NAND2X0 U15586 ( .IN1(n14743), .IN2(n14744), .QN(g28050) );
  NAND2X0 U15587 ( .IN1(n14733), .IN2(g655), .QN(n14744) );
  NAND2X0 U15588 ( .IN1(n14734), .IN2(g650), .QN(n14743) );
  NAND3X0 U15589 ( .IN1(n14745), .IN2(n14746), .IN3(n14747), .QN(g28049) );
  NAND2X0 U15590 ( .IN1(test_so87), .IN2(n9514), .QN(n14747) );
  NAND2X0 U15591 ( .IN1(n14738), .IN2(g681), .QN(n14746) );
  NAND2X0 U15592 ( .IN1(n14733), .IN2(g650), .QN(n14745) );
  NAND3X0 U15593 ( .IN1(n14748), .IN2(n14749), .IN3(n14750), .QN(g28048) );
  NAND2X0 U15594 ( .IN1(n9458), .IN2(g29212), .QN(n14750) );
  NAND2X0 U15595 ( .IN1(n14751), .IN2(g691), .QN(n14749) );
  NAND2X0 U15596 ( .IN1(n14752), .IN2(n14753), .QN(n14751) );
  NAND3X0 U15597 ( .IN1(g703), .IN2(n8879), .IN3(n9337), .QN(n14753) );
  NAND2X0 U15598 ( .IN1(n14754), .IN2(n14755), .QN(n14748) );
  INVX0 U15599 ( .INP(n4819), .ZN(n14755) );
  NAND4X0 U15600 ( .IN1(n5520), .IN2(n5112), .IN3(n14756), .IN4(g703), .QN(
        n4819) );
  INVX0 U15601 ( .INP(n14128), .ZN(n14756) );
  NAND4X0 U15602 ( .IN1(n14757), .IN2(n14758), .IN3(test_so87), .IN4(n14759), 
        .QN(n14128) );
  NOR2X0 U15603 ( .IN1(g645), .IN2(g650), .QN(n14759) );
  NAND2X0 U15604 ( .IN1(n8475), .IN2(g661), .QN(n14758) );
  NAND2X0 U15605 ( .IN1(n8474), .IN2(g728), .QN(n14757) );
  NAND2X0 U15606 ( .IN1(n14760), .IN2(n14761), .QN(g28047) );
  NAND2X0 U15607 ( .IN1(n14733), .IN2(g681), .QN(n14761) );
  NAND2X0 U15608 ( .IN1(n14734), .IN2(g645), .QN(n14760) );
  NAND2X0 U15609 ( .IN1(n14762), .IN2(n14763), .QN(g28046) );
  NAND2X0 U15610 ( .IN1(n14738), .IN2(g446), .QN(n14763) );
  NOR2X0 U15611 ( .IN1(n14764), .IN2(n9406), .QN(n14738) );
  NAND2X0 U15612 ( .IN1(n14733), .IN2(g645), .QN(n14762) );
  INVX0 U15613 ( .INP(n14734), .ZN(n14733) );
  NAND2X0 U15614 ( .IN1(n14764), .IN2(n9381), .QN(n14734) );
  NAND4X0 U15615 ( .IN1(n8816), .IN2(n14765), .IN3(n14766), .IN4(n14767), .QN(
        n14764) );
  INVX0 U15616 ( .INP(n14768), .ZN(n14767) );
  NOR2X0 U15617 ( .IN1(n14769), .IN2(n5520), .QN(n14768) );
  NAND2X0 U15618 ( .IN1(n5520), .IN2(n14770), .QN(n14766) );
  NAND3X0 U15619 ( .IN1(n5629), .IN2(g417), .IN3(n8784), .QN(n14770) );
  NAND3X0 U15620 ( .IN1(n14771), .IN2(n14772), .IN3(n14773), .QN(g28045) );
  NAND2X0 U15621 ( .IN1(n9458), .IN2(g568), .QN(n14773) );
  NAND3X0 U15622 ( .IN1(n2421), .IN2(n14774), .IN3(g572), .QN(n14772) );
  INVX0 U15623 ( .INP(n4537), .ZN(n14774) );
  NAND2X0 U15624 ( .IN1(n4537), .IN2(n5337), .QN(n14771) );
  NAND2X0 U15625 ( .IN1(n14775), .IN2(n14776), .QN(g28044) );
  NAND2X0 U15626 ( .IN1(n9458), .IN2(g528), .QN(n14776) );
  NAND2X0 U15627 ( .IN1(n14777), .IN2(n9381), .QN(n14775) );
  NAND2X0 U15628 ( .IN1(n14778), .IN2(n14141), .QN(n14777) );
  NAND2X0 U15629 ( .IN1(n14779), .IN2(n14780), .QN(n14778) );
  NAND2X0 U15630 ( .IN1(n5820), .IN2(n14781), .QN(n14780) );
  INVX0 U15631 ( .INP(n14139), .ZN(n14779) );
  NOR2X0 U15632 ( .IN1(n14781), .IN2(n5820), .QN(n14139) );
  NAND2X0 U15633 ( .IN1(n14782), .IN2(n14783), .QN(n14781) );
  NAND2X0 U15634 ( .IN1(n5327), .IN2(n14784), .QN(n14783) );
  NAND2X0 U15635 ( .IN1(n14785), .IN2(n14786), .QN(g28043) );
  NAND2X0 U15636 ( .IN1(n10734), .IN2(n8874), .QN(n14786) );
  NOR2X0 U15637 ( .IN1(n12320), .IN2(n9384), .QN(n10734) );
  NAND4X0 U15638 ( .IN1(n14787), .IN2(n9785), .IN3(n13559), .IN4(g691), .QN(
        n12320) );
  NAND4X0 U15639 ( .IN1(n14788), .IN2(n14789), .IN3(n14790), .IN4(n14791), 
        .QN(n13559) );
  NAND3X0 U15640 ( .IN1(g655), .IN2(g753), .IN3(g718), .QN(n14791) );
  NAND3X0 U15641 ( .IN1(n8828), .IN2(n8827), .IN3(n8829), .QN(n14790) );
  NAND2X0 U15642 ( .IN1(g807), .IN2(g554), .QN(n14789) );
  NAND2X0 U15643 ( .IN1(n5627), .IN2(n14792), .QN(n9785) );
  NAND4X0 U15644 ( .IN1(g262), .IN2(g269), .IN3(g255), .IN4(n14793), .QN(
        n14792) );
  NOR2X0 U15645 ( .IN1(n14794), .IN2(g232), .QN(n14793) );
  NAND2X0 U15646 ( .IN1(n9786), .IN2(g278), .QN(n14787) );
  NAND4X0 U15647 ( .IN1(n8471), .IN2(n8470), .IN3(n8472), .IN4(n14795), .QN(
        n9786) );
  NOR4X0 U15648 ( .IN1(n8590), .IN2(n8589), .IN3(n6008), .IN4(n5597), .QN(
        n14795) );
  NAND2X0 U15649 ( .IN1(n9457), .IN2(g278), .QN(n14785) );
  NAND3X0 U15650 ( .IN1(n5796), .IN2(n9315), .IN3(n5630), .QN(g28042) );
  NAND3X0 U15651 ( .IN1(n14796), .IN2(n9316), .IN3(n10271), .QN(g28041) );
  INVX0 U15652 ( .INP(n10199), .ZN(n10271) );
  NOR2X0 U15653 ( .IN1(n9807), .IN2(n8812), .QN(n10199) );
  INVX0 U15654 ( .INP(n10198), .ZN(n14796) );
  NOR2X0 U15655 ( .IN1(n14797), .IN2(n8811), .QN(n10198) );
  NAND2X0 U15656 ( .IN1(n14798), .IN2(n14799), .QN(g28030) );
  NAND3X0 U15657 ( .IN1(n5861), .IN2(n14800), .IN3(n5882), .QN(n14799) );
  NAND2X0 U15658 ( .IN1(n14801), .IN2(n14802), .QN(n14800) );
  NAND2X0 U15659 ( .IN1(n14803), .IN2(n10223), .QN(n14802) );
  NAND2X0 U15660 ( .IN1(n14804), .IN2(n14805), .QN(n14803) );
  NAND3X0 U15661 ( .IN1(n5872), .IN2(n14806), .IN3(n5886), .QN(n14805) );
  NAND2X0 U15662 ( .IN1(n14807), .IN2(n14808), .QN(n14806) );
  NAND2X0 U15663 ( .IN1(n14809), .IN2(n14810), .QN(n14808) );
  NAND2X0 U15664 ( .IN1(n14811), .IN2(n14812), .QN(n14809) );
  NAND4X0 U15665 ( .IN1(n5885), .IN2(n5869), .IN3(n14813), .IN4(n14814), .QN(
        n14812) );
  NAND3X0 U15666 ( .IN1(n5874), .IN2(n14815), .IN3(n5888), .QN(n14811) );
  NAND2X0 U15667 ( .IN1(n14816), .IN2(n14817), .QN(n14815) );
  NAND3X0 U15668 ( .IN1(n5869), .IN2(n14818), .IN3(n5885), .QN(n14817) );
  INVX0 U15669 ( .INP(n14819), .ZN(n14818) );
  NOR2X0 U15670 ( .IN1(n14814), .IN2(n14813), .QN(n14819) );
  NAND2X0 U15671 ( .IN1(n14813), .IN2(n14814), .QN(n14816) );
  NAND2X0 U15672 ( .IN1(n14820), .IN2(n14810), .QN(n14804) );
  NAND2X0 U15673 ( .IN1(n10222), .IN2(n10223), .QN(n14798) );
  NAND2X0 U15674 ( .IN1(n14821), .IN2(n9381), .QN(n10223) );
  NAND2X0 U15675 ( .IN1(n5889), .IN2(n5868), .QN(n14821) );
  INVX0 U15676 ( .INP(n14801), .ZN(n10222) );
  NAND3X0 U15677 ( .IN1(n14822), .IN2(n14810), .IN3(n14820), .QN(n14801) );
  INVX0 U15678 ( .INP(n14807), .ZN(n14820) );
  NAND3X0 U15679 ( .IN1(n14813), .IN2(n14814), .IN3(n14823), .QN(n14807) );
  NAND2X0 U15680 ( .IN1(n14824), .IN2(n9381), .QN(n14823) );
  NAND4X0 U15681 ( .IN1(n5888), .IN2(n5885), .IN3(n5874), .IN4(n5869), .QN(
        n14824) );
  INVX0 U15682 ( .INP(n14825), .ZN(n14814) );
  NOR2X0 U15683 ( .IN1(n14826), .IN2(n9391), .QN(n14825) );
  NOR2X0 U15684 ( .IN1(g5831), .IN2(test_so83), .QN(n14826) );
  NAND2X0 U15685 ( .IN1(n14827), .IN2(n9381), .QN(n14813) );
  NAND2X0 U15686 ( .IN1(n5884), .IN2(n5870), .QN(n14827) );
  NAND2X0 U15687 ( .IN1(n14828), .IN2(n9381), .QN(n14810) );
  NAND2X0 U15688 ( .IN1(n5883), .IN2(n5871), .QN(n14828) );
  NAND2X0 U15689 ( .IN1(n14829), .IN2(n9381), .QN(n14822) );
  NAND2X0 U15690 ( .IN1(n5886), .IN2(n5872), .QN(n14829) );
  NAND3X0 U15691 ( .IN1(n14830), .IN2(n14831), .IN3(n12393), .QN(g26971) );
  NAND2X0 U15692 ( .IN1(n5670), .IN2(n9381), .QN(n12393) );
  NAND2X0 U15693 ( .IN1(n15958), .IN2(n9381), .QN(n14831) );
  NAND2X0 U15694 ( .IN1(n9457), .IN2(g4512), .QN(n14830) );
  NAND2X0 U15695 ( .IN1(n14832), .IN2(n14833), .QN(g26970) );
  NAND2X0 U15696 ( .IN1(n9363), .IN2(g4473), .QN(n14833) );
  NAND2X0 U15697 ( .IN1(n9457), .IN2(g4459), .QN(n14832) );
  NAND2X0 U15698 ( .IN1(n14834), .IN2(n14835), .QN(g26969) );
  NAND2X0 U15699 ( .IN1(n9457), .IN2(g4462), .QN(n14835) );
  NAND3X0 U15700 ( .IN1(n8423), .IN2(n8864), .IN3(n9337), .QN(n14834) );
  NAND2X0 U15701 ( .IN1(n14836), .IN2(n14837), .QN(g26968) );
  NAND2X0 U15702 ( .IN1(n9457), .IN2(g4558), .QN(n14836) );
  NAND2X0 U15703 ( .IN1(n14838), .IN2(n14839), .QN(g26967) );
  NAND2X0 U15704 ( .IN1(n9457), .IN2(g4561), .QN(n14838) );
  NAND2X0 U15705 ( .IN1(n14840), .IN2(n14841), .QN(g26966) );
  NAND2X0 U15706 ( .IN1(n9457), .IN2(g4555), .QN(n14840) );
  NOR2X0 U15707 ( .IN1(n14842), .IN2(n14843), .QN(g26965) );
  NOR2X0 U15708 ( .IN1(n15959), .IN2(n14844), .QN(n14843) );
  INVX0 U15709 ( .INP(n14845), .ZN(n14842) );
  NAND2X0 U15710 ( .IN1(n14844), .IN2(n15959), .QN(n14845) );
  NAND2X0 U15711 ( .IN1(n9363), .IN2(g10306), .QN(n14844) );
  NAND2X0 U15712 ( .IN1(n14846), .IN2(n14847), .QN(g26964) );
  NAND3X0 U15713 ( .IN1(n14848), .IN2(n14849), .IN3(n9337), .QN(n14847) );
  NAND2X0 U15714 ( .IN1(n8714), .IN2(g4521), .QN(n14849) );
  NAND2X0 U15715 ( .IN1(n5752), .IN2(n14850), .QN(n14848) );
  NAND2X0 U15716 ( .IN1(n8725), .IN2(n10832), .QN(n14850) );
  INVX0 U15717 ( .INP(n14515), .ZN(n10832) );
  NAND2X0 U15718 ( .IN1(n14851), .IN2(g4527), .QN(n14846) );
  NAND2X0 U15719 ( .IN1(n14852), .IN2(n9381), .QN(n14851) );
  NAND2X0 U15720 ( .IN1(n5752), .IN2(n14515), .QN(n14852) );
  NAND4X0 U15721 ( .IN1(test_so27), .IN2(g4483), .IN3(g4489), .IN4(g4492), 
        .QN(n14515) );
  NAND2X0 U15722 ( .IN1(n14853), .IN2(n14839), .QN(g26963) );
  NAND2X0 U15723 ( .IN1(g6750), .IN2(n9381), .QN(n14839) );
  NAND2X0 U15724 ( .IN1(n9456), .IN2(g4489), .QN(n14853) );
  NAND2X0 U15725 ( .IN1(n14837), .IN2(n14854), .QN(g26962) );
  NAND2X0 U15726 ( .IN1(test_so27), .IN2(n9512), .QN(n14854) );
  NAND2X0 U15727 ( .IN1(g6749), .IN2(n9381), .QN(n14837) );
  NAND2X0 U15728 ( .IN1(n14855), .IN2(n14841), .QN(g26961) );
  NAND2X0 U15729 ( .IN1(g6748), .IN2(n9381), .QN(n14841) );
  NAND2X0 U15730 ( .IN1(n9456), .IN2(g4483), .QN(n14855) );
  NAND2X0 U15731 ( .IN1(n14856), .IN2(n14857), .QN(g26958) );
  NAND2X0 U15732 ( .IN1(n9456), .IN2(g4455), .QN(n14857) );
  NAND2X0 U15733 ( .IN1(n14858), .IN2(n14859), .QN(g26957) );
  NAND2X0 U15734 ( .IN1(n14860), .IN2(g4434), .QN(n14859) );
  NAND2X0 U15735 ( .IN1(n14861), .IN2(n9381), .QN(n14860) );
  NAND2X0 U15736 ( .IN1(n14862), .IN2(g4392), .QN(n14861) );
  NAND2X0 U15737 ( .IN1(test_so47), .IN2(n9381), .QN(n14858) );
  NAND2X0 U15738 ( .IN1(n15961), .IN2(n14863), .QN(g26956) );
  NAND3X0 U15739 ( .IN1(n14862), .IN2(g4430), .IN3(n14864), .QN(n14863) );
  NAND2X0 U15740 ( .IN1(n14865), .IN2(n14866), .QN(g26955) );
  NAND3X0 U15741 ( .IN1(n9350), .IN2(g4392), .IN3(n14862), .QN(n14866) );
  NAND2X0 U15742 ( .IN1(n14867), .IN2(g4438), .QN(n14865) );
  NAND3X0 U15743 ( .IN1(n14868), .IN2(n14869), .IN3(n14870), .QN(g26954) );
  NAND2X0 U15744 ( .IN1(test_so47), .IN2(n9514), .QN(n14870) );
  NAND2X0 U15745 ( .IN1(n14864), .IN2(n14862), .QN(n14869) );
  INVX0 U15746 ( .INP(n14871), .ZN(n14862) );
  NAND4X0 U15747 ( .IN1(n15961), .IN2(n8719), .IN3(n14872), .IN4(DFF_1225_n1), 
        .QN(n14871) );
  NOR2X0 U15748 ( .IN1(test_so47), .IN2(g7260), .QN(n14872) );
  NAND2X0 U15749 ( .IN1(n14873), .IN2(g4438), .QN(n14868) );
  NAND2X0 U15750 ( .IN1(n14874), .IN2(n14875), .QN(g26952) );
  NAND2X0 U15751 ( .IN1(n14876), .IN2(g4430), .QN(n14875) );
  NAND2X0 U15752 ( .IN1(n9363), .IN2(g4388), .QN(n14876) );
  NAND2X0 U15753 ( .IN1(n14877), .IN2(n9382), .QN(n14874) );
  NAND3X0 U15754 ( .IN1(n14878), .IN2(n14879), .IN3(n14880), .QN(n14877) );
  NAND2X0 U15755 ( .IN1(n8405), .IN2(g4388), .QN(n14880) );
  NAND2X0 U15756 ( .IN1(n8403), .IN2(g4401), .QN(n14879) );
  NAND2X0 U15757 ( .IN1(n8402), .IN2(g4434), .QN(n14878) );
  NAND2X0 U15758 ( .IN1(n14856), .IN2(n14881), .QN(g26950) );
  INVX0 U15759 ( .INP(n14882), .ZN(n14881) );
  NOR2X0 U15760 ( .IN1(n9358), .IN2(n8333), .QN(n14882) );
  NAND2X0 U15761 ( .IN1(n14883), .IN2(n9382), .QN(n14856) );
  NAND2X0 U15762 ( .IN1(n14884), .IN2(n14885), .QN(n14883) );
  NAND2X0 U15763 ( .IN1(n14886), .IN2(g4392), .QN(n14885) );
  NAND2X0 U15764 ( .IN1(n14887), .IN2(n14888), .QN(g26949) );
  NAND2X0 U15765 ( .IN1(n14889), .IN2(g4401), .QN(n14888) );
  NAND2X0 U15766 ( .IN1(n14890), .IN2(n9382), .QN(n14889) );
  NAND2X0 U15767 ( .IN1(n14891), .IN2(g4392), .QN(n14890) );
  NAND2X0 U15768 ( .IN1(n9363), .IN2(g4411), .QN(n14887) );
  NAND2X0 U15769 ( .IN1(n8838), .IN2(n14892), .QN(g26948) );
  NAND3X0 U15770 ( .IN1(n14891), .IN2(g4388), .IN3(n14864), .QN(n14892) );
  NAND2X0 U15771 ( .IN1(n14893), .IN2(n14894), .QN(g26947) );
  NAND2X0 U15772 ( .IN1(n9456), .IN2(g4388), .QN(n14894) );
  NAND2X0 U15773 ( .IN1(n14895), .IN2(n9382), .QN(n14893) );
  NAND2X0 U15774 ( .IN1(n14884), .IN2(n14896), .QN(n14895) );
  NAND2X0 U15775 ( .IN1(n14897), .IN2(n14886), .QN(n14896) );
  NAND2X0 U15776 ( .IN1(n14898), .IN2(n14899), .QN(n14897) );
  NAND2X0 U15777 ( .IN1(n8837), .IN2(g4382), .QN(n14899) );
  NAND2X0 U15778 ( .IN1(n5714), .IN2(g4375), .QN(n14898) );
  NAND3X0 U15779 ( .IN1(n5710), .IN2(n14891), .IN3(n8333), .QN(n14884) );
  NAND2X0 U15780 ( .IN1(n14900), .IN2(n14901), .QN(g26946) );
  NAND3X0 U15781 ( .IN1(n9350), .IN2(g4392), .IN3(n14891), .QN(n14901) );
  NAND2X0 U15782 ( .IN1(n14867), .IN2(g4375), .QN(n14900) );
  INVX0 U15783 ( .INP(n14873), .ZN(n14867) );
  NAND3X0 U15784 ( .IN1(n14902), .IN2(n14903), .IN3(n14904), .QN(g26945) );
  NAND2X0 U15785 ( .IN1(n9456), .IN2(g4411), .QN(n14904) );
  NAND2X0 U15786 ( .IN1(n14864), .IN2(n14891), .QN(n14903) );
  INVX0 U15787 ( .INP(n14886), .ZN(n14891) );
  NAND4X0 U15788 ( .IN1(n8838), .IN2(n8837), .IN3(n8839), .IN4(n14905), .QN(
        n14886) );
  NOR2X0 U15789 ( .IN1(g4411), .IN2(g7257), .QN(n14905) );
  NOR2X0 U15790 ( .IN1(g4392), .IN2(n9395), .QN(n14864) );
  NAND2X0 U15791 ( .IN1(n14873), .IN2(g4375), .QN(n14902) );
  NOR2X0 U15792 ( .IN1(g4382), .IN2(n9395), .QN(n14873) );
  NOR2X0 U15793 ( .IN1(n9414), .IN2(n14906), .QN(g26944) );
  NOR4X0 U15794 ( .IN1(n14907), .IN2(n14908), .IN3(n8867), .IN4(n10698), .QN(
        n14906) );
  INVX0 U15795 ( .INP(n10137), .ZN(n14908) );
  NOR2X0 U15796 ( .IN1(n14909), .IN2(g135), .QN(n10137) );
  INVX0 U15797 ( .INP(n14910), .ZN(n14909) );
  NAND3X0 U15798 ( .IN1(n14911), .IN2(n14912), .IN3(n14913), .QN(n14910) );
  NAND4X0 U15799 ( .IN1(n14914), .IN2(n5608), .IN3(n14915), .IN4(n14916), .QN(
        n14913) );
  NAND2X0 U15800 ( .IN1(n5539), .IN2(g4608), .QN(n14916) );
  NAND2X0 U15801 ( .IN1(n5274), .IN2(g4584), .QN(n14915) );
  NOR2X0 U15802 ( .IN1(n14917), .IN2(n14918), .QN(n14914) );
  NOR2X0 U15803 ( .IN1(n5365), .IN2(g4593), .QN(n14918) );
  NOR2X0 U15804 ( .IN1(n5303), .IN2(g4601), .QN(n14917) );
  NAND4X0 U15805 ( .IN1(n5365), .IN2(g4593), .IN3(n5274), .IN4(g4584), .QN(
        n14912) );
  NAND3X0 U15806 ( .IN1(n5303), .IN2(g4608), .IN3(n5539), .QN(n14911) );
  NAND3X0 U15807 ( .IN1(g4340), .IN2(g4633), .IN3(g4358), .QN(n14907) );
  NAND2X0 U15808 ( .IN1(n14919), .IN2(n14920), .QN(g26940) );
  NAND2X0 U15809 ( .IN1(n9456), .IN2(g4153), .QN(n14920) );
  NAND2X0 U15810 ( .IN1(n12906), .IN2(n9382), .QN(n14919) );
  NAND2X0 U15811 ( .IN1(n14921), .IN2(n14922), .QN(n12906) );
  NAND2X0 U15812 ( .IN1(g116), .IN2(g4157), .QN(n14922) );
  NAND2X0 U15813 ( .IN1(g114), .IN2(n5983), .QN(n14921) );
  NAND2X0 U15814 ( .IN1(n14923), .IN2(n14924), .QN(g26939) );
  NAND2X0 U15815 ( .IN1(n9456), .IN2(g4104), .QN(n14924) );
  NAND2X0 U15816 ( .IN1(n12901), .IN2(n9382), .QN(n14923) );
  NAND2X0 U15817 ( .IN1(n14925), .IN2(n14926), .QN(n12901) );
  NAND2X0 U15818 ( .IN1(g124), .IN2(g4146), .QN(n14926) );
  NAND2X0 U15819 ( .IN1(g120), .IN2(n5981), .QN(n14925) );
  NAND3X0 U15820 ( .IN1(n14927), .IN2(n12032), .IN3(n14928), .QN(g26938) );
  NAND2X0 U15821 ( .IN1(n14929), .IN2(g4141), .QN(n14928) );
  NAND2X0 U15822 ( .IN1(n14930), .IN2(n9382), .QN(n14929) );
  NAND2X0 U15823 ( .IN1(n14540), .IN2(n9808), .QN(n14930) );
  NAND3X0 U15824 ( .IN1(n9349), .IN2(g4082), .IN3(n14540), .QN(n14927) );
  NAND3X0 U15825 ( .IN1(g4141), .IN2(g4082), .IN3(n9808), .QN(n14540) );
  NAND3X0 U15826 ( .IN1(n14931), .IN2(n14932), .IN3(n14933), .QN(g26934) );
  NAND2X0 U15827 ( .IN1(n4888), .IN2(g2827), .QN(n14933) );
  INVX0 U15828 ( .INP(n14934), .ZN(n14932) );
  NOR2X0 U15829 ( .IN1(n14935), .IN2(test_so34), .QN(n14934) );
  NAND2X0 U15830 ( .IN1(test_so37), .IN2(n9414), .QN(n14931) );
  NAND3X0 U15831 ( .IN1(n14936), .IN2(n14937), .IN3(n14938), .QN(g26933) );
  NAND2X0 U15832 ( .IN1(n4888), .IN2(test_so37), .QN(n14938) );
  NAND2X0 U15833 ( .IN1(n5840), .IN2(n14939), .QN(n14937) );
  NAND2X0 U15834 ( .IN1(n9455), .IN2(g2811), .QN(n14936) );
  NAND3X0 U15835 ( .IN1(n14940), .IN2(n14941), .IN3(n14942), .QN(g26932) );
  NAND2X0 U15836 ( .IN1(n4888), .IN2(g2811), .QN(n14942) );
  NAND2X0 U15837 ( .IN1(n5841), .IN2(n14939), .QN(n14941) );
  NAND2X0 U15838 ( .IN1(n9455), .IN2(g2799), .QN(n14940) );
  NAND3X0 U15839 ( .IN1(n14943), .IN2(n14944), .IN3(n14945), .QN(g26931) );
  NAND2X0 U15840 ( .IN1(n4888), .IN2(g2799), .QN(n14945) );
  NAND2X0 U15841 ( .IN1(n5839), .IN2(n14939), .QN(n14944) );
  NAND2X0 U15842 ( .IN1(n9455), .IN2(g29219), .QN(n14943) );
  NAND3X0 U15843 ( .IN1(n14946), .IN2(n14947), .IN3(n14948), .QN(g26930) );
  NAND2X0 U15844 ( .IN1(n4888), .IN2(g2795), .QN(n14948) );
  INVX0 U15845 ( .INP(n14949), .ZN(n14947) );
  NOR2X0 U15846 ( .IN1(n14935), .IN2(test_so59), .QN(n14949) );
  NAND2X0 U15847 ( .IN1(n9455), .IN2(g2791), .QN(n14946) );
  NAND3X0 U15848 ( .IN1(n14950), .IN2(n14951), .IN3(n14952), .QN(g26929) );
  NAND2X0 U15849 ( .IN1(n4888), .IN2(g2791), .QN(n14952) );
  NAND2X0 U15850 ( .IN1(n5837), .IN2(n14939), .QN(n14951) );
  NAND2X0 U15851 ( .IN1(n9455), .IN2(g2779), .QN(n14950) );
  NAND3X0 U15852 ( .IN1(n14953), .IN2(n14954), .IN3(n14955), .QN(g26928) );
  NAND2X0 U15853 ( .IN1(n4888), .IN2(g2779), .QN(n14955) );
  NAND2X0 U15854 ( .IN1(n5834), .IN2(n14939), .QN(n14954) );
  NAND2X0 U15855 ( .IN1(n9455), .IN2(g2767), .QN(n14953) );
  NAND3X0 U15856 ( .IN1(n14956), .IN2(n14957), .IN3(n14958), .QN(g26927) );
  NAND2X0 U15857 ( .IN1(n4888), .IN2(g2767), .QN(n14958) );
  NAND2X0 U15858 ( .IN1(n5836), .IN2(n14939), .QN(n14957) );
  INVX0 U15859 ( .INP(n14935), .ZN(n14939) );
  NAND3X0 U15860 ( .IN1(n14959), .IN2(n10531), .IN3(n4888), .QN(n14935) );
  NAND3X0 U15861 ( .IN1(n3505), .IN2(g2735), .IN3(test_so30), .QN(n10531) );
  NOR2X0 U15862 ( .IN1(n5349), .IN2(n5516), .QN(n3505) );
  NAND2X0 U15863 ( .IN1(n5516), .IN2(n5300), .QN(n14959) );
  NAND2X0 U15864 ( .IN1(n9455), .IN2(g2763), .QN(n14956) );
  NAND2X0 U15865 ( .IN1(n14960), .IN2(n14961), .QN(g26926) );
  NAND3X0 U15866 ( .IN1(n14962), .IN2(n14963), .IN3(n3730), .QN(n14961) );
  NAND2X0 U15867 ( .IN1(n5301), .IN2(n14697), .QN(n14963) );
  INVX0 U15868 ( .INP(n13185), .ZN(n14697) );
  NAND2X0 U15869 ( .IN1(n13185), .IN2(g2724), .QN(n14962) );
  NOR2X0 U15870 ( .IN1(n5299), .IN2(n5465), .QN(n13185) );
  NAND2X0 U15871 ( .IN1(n9454), .IN2(g2719), .QN(n14960) );
  NAND2X0 U15872 ( .IN1(n14964), .IN2(n14965), .QN(g26925) );
  NAND2X0 U15873 ( .IN1(n9454), .IN2(g1532), .QN(n14965) );
  NAND2X0 U15874 ( .IN1(n14966), .IN2(n9382), .QN(n14964) );
  NAND2X0 U15875 ( .IN1(n13493), .IN2(n14967), .QN(n14966) );
  NAND2X0 U15876 ( .IN1(n13473), .IN2(g1536), .QN(n14967) );
  NAND2X0 U15877 ( .IN1(n13481), .IN2(g1413), .QN(n13473) );
  NOR2X0 U15878 ( .IN1(n13480), .IN2(n8764), .QN(n13481) );
  NAND3X0 U15879 ( .IN1(n14968), .IN2(g7946), .IN3(n13495), .QN(n13480) );
  NAND3X0 U15880 ( .IN1(g1339), .IN2(g1521), .IN3(n8588), .QN(n14968) );
  INVX0 U15881 ( .INP(n4173), .ZN(n13493) );
  NAND3X0 U15882 ( .IN1(n14969), .IN2(n14970), .IN3(n14971), .QN(g26924) );
  INVX0 U15883 ( .INP(n14972), .ZN(n14971) );
  NOR2X0 U15884 ( .IN1(n14973), .IN2(g1478), .QN(n14972) );
  NAND3X0 U15885 ( .IN1(n14973), .IN2(g1478), .IN3(n9337), .QN(n14970) );
  NAND4X0 U15886 ( .IN1(n14974), .IN2(n14044), .IN3(g1437), .IN4(n8859), .QN(
        n14973) );
  NAND2X0 U15887 ( .IN1(n9454), .IN2(g1437), .QN(n14969) );
  NAND3X0 U15888 ( .IN1(n14975), .IN2(n14976), .IN3(n14977), .QN(g26923) );
  INVX0 U15889 ( .INP(n14978), .ZN(n14977) );
  NOR2X0 U15890 ( .IN1(n14979), .IN2(g1472), .QN(n14978) );
  NAND3X0 U15891 ( .IN1(n14979), .IN2(g1472), .IN3(n9337), .QN(n14976) );
  NAND4X0 U15892 ( .IN1(n14974), .IN2(n14044), .IN3(test_so49), .IN4(g1467), 
        .QN(n14979) );
  NOR2X0 U15893 ( .IN1(n8798), .IN2(n5364), .QN(n14044) );
  NAND2X0 U15894 ( .IN1(n9454), .IN2(g1467), .QN(n14975) );
  NAND3X0 U15895 ( .IN1(n14980), .IN2(n14981), .IN3(n14982), .QN(g26922) );
  INVX0 U15896 ( .INP(n14983), .ZN(n14982) );
  NOR2X0 U15897 ( .IN1(n14984), .IN2(g1448), .QN(n14983) );
  NAND3X0 U15898 ( .IN1(n14984), .IN2(g1448), .IN3(n9337), .QN(n14981) );
  NAND3X0 U15899 ( .IN1(n14024), .IN2(g1454), .IN3(n14974), .QN(n14984) );
  NOR2X0 U15900 ( .IN1(n11633), .IN2(n8798), .QN(n14024) );
  INVX0 U15901 ( .INP(n13495), .ZN(n11633) );
  NOR2X0 U15902 ( .IN1(g1514), .IN2(n8859), .QN(n13495) );
  NAND2X0 U15903 ( .IN1(n9454), .IN2(g1454), .QN(n14980) );
  NAND2X0 U15904 ( .IN1(n14985), .IN2(n14986), .QN(g26921) );
  NAND2X0 U15905 ( .IN1(n9454), .IN2(g1395), .QN(n14986) );
  NAND4X0 U15906 ( .IN1(n14987), .IN2(n14988), .IN3(n8875), .IN4(n9362), .QN(
        n14985) );
  NAND2X0 U15907 ( .IN1(n8450), .IN2(n14989), .QN(n14988) );
  INVX0 U15908 ( .INP(n14990), .ZN(n14987) );
  NOR2X0 U15909 ( .IN1(n14989), .IN2(n8450), .QN(n14990) );
  NAND2X0 U15910 ( .IN1(n14991), .IN2(n14992), .QN(g26920) );
  NAND2X0 U15911 ( .IN1(n9454), .IN2(g1384), .QN(n14992) );
  NAND2X0 U15912 ( .IN1(n14993), .IN2(n9382), .QN(n14991) );
  NAND2X0 U15913 ( .IN1(n14994), .IN2(n14995), .QN(n14993) );
  NAND2X0 U15914 ( .IN1(n9801), .IN2(g1389), .QN(n14995) );
  NAND2X0 U15915 ( .IN1(n14996), .IN2(n14997), .QN(n9801) );
  NAND2X0 U15916 ( .IN1(n8340), .IN2(g1351), .QN(n14997) );
  NAND2X0 U15917 ( .IN1(n4913), .IN2(g1351), .QN(n14994) );
  NAND3X0 U15918 ( .IN1(n14998), .IN2(n14999), .IN3(n15000), .QN(g26919) );
  NAND2X0 U15919 ( .IN1(n9453), .IN2(g1266), .QN(n15000) );
  NAND3X0 U15920 ( .IN1(test_so77), .IN2(n11853), .IN3(n9809), .QN(n14999) );
  INVX0 U15921 ( .INP(n15001), .ZN(n14998) );
  NOR2X0 U15922 ( .IN1(n9809), .IN2(test_so77), .QN(n15001) );
  NAND3X0 U15923 ( .IN1(g1249), .IN2(g1266), .IN3(g12923), .QN(n9809) );
  NAND2X0 U15924 ( .IN1(n15002), .IN2(n15003), .QN(g26918) );
  NAND2X0 U15925 ( .IN1(n9453), .IN2(g1189), .QN(n15003) );
  NAND2X0 U15926 ( .IN1(n15004), .IN2(n9382), .QN(n15002) );
  NAND2X0 U15927 ( .IN1(n13530), .IN2(n15005), .QN(n15004) );
  NAND2X0 U15928 ( .IN1(n13511), .IN2(g1193), .QN(n15005) );
  NAND2X0 U15929 ( .IN1(n13519), .IN2(g1070), .QN(n13511) );
  NOR2X0 U15930 ( .IN1(n13518), .IN2(n8763), .QN(n13519) );
  NAND3X0 U15931 ( .IN1(n15006), .IN2(g7916), .IN3(n13532), .QN(n13518) );
  NAND3X0 U15932 ( .IN1(g1178), .IN2(g996), .IN3(n5642), .QN(n15006) );
  INVX0 U15933 ( .INP(n4191), .ZN(n13530) );
  NAND2X0 U15934 ( .IN1(n15007), .IN2(n15008), .QN(g26917) );
  NAND2X0 U15935 ( .IN1(n15009), .IN2(g1094), .QN(n15008) );
  NAND2X0 U15936 ( .IN1(n15010), .IN2(n9382), .QN(n15009) );
  NAND3X0 U15937 ( .IN1(n14094), .IN2(n5328), .IN3(n15011), .QN(n15010) );
  NAND3X0 U15938 ( .IN1(n9349), .IN2(g1135), .IN3(n15012), .QN(n15007) );
  NAND3X0 U15939 ( .IN1(n14094), .IN2(g1094), .IN3(n15011), .QN(n15012) );
  NOR3X0 U15940 ( .IN1(n5363), .IN2(n8804), .IN3(g1183), .QN(n14094) );
  NAND3X0 U15941 ( .IN1(n15013), .IN2(n15014), .IN3(n15015), .QN(g26916) );
  INVX0 U15942 ( .INP(n15016), .ZN(n15015) );
  NOR2X0 U15943 ( .IN1(n15017), .IN2(g1129), .QN(n15016) );
  NAND3X0 U15944 ( .IN1(n15017), .IN2(g1129), .IN3(n9337), .QN(n15014) );
  NAND4X0 U15945 ( .IN1(n15011), .IN2(n11762), .IN3(g1124), .IN4(g13259), .QN(
        n15017) );
  NAND2X0 U15946 ( .IN1(n9453), .IN2(g1124), .QN(n15013) );
  NAND3X0 U15947 ( .IN1(n15018), .IN2(n15019), .IN3(n15020), .QN(g26915) );
  INVX0 U15948 ( .INP(n15021), .ZN(n15020) );
  NOR2X0 U15949 ( .IN1(n15022), .IN2(g1105), .QN(n15021) );
  NAND3X0 U15950 ( .IN1(n15022), .IN2(g1105), .IN3(n9337), .QN(n15019) );
  NAND3X0 U15951 ( .IN1(test_so90), .IN2(n14066), .IN3(n15011), .QN(n15022) );
  NOR2X0 U15952 ( .IN1(n11800), .IN2(n8804), .QN(n14066) );
  INVX0 U15953 ( .INP(n13532), .ZN(n11800) );
  NOR2X0 U15954 ( .IN1(g1171), .IN2(n5599), .QN(n13532) );
  NAND2X0 U15955 ( .IN1(test_so90), .IN2(n9511), .QN(n15018) );
  NAND2X0 U15956 ( .IN1(n15023), .IN2(n15024), .QN(g26914) );
  NAND2X0 U15957 ( .IN1(n9453), .IN2(g1052), .QN(n15024) );
  NAND4X0 U15958 ( .IN1(n15025), .IN2(n15026), .IN3(n5320), .IN4(n9362), .QN(
        n15023) );
  NAND2X0 U15959 ( .IN1(n8451), .IN2(n15027), .QN(n15026) );
  INVX0 U15960 ( .INP(n15028), .ZN(n15025) );
  NOR2X0 U15961 ( .IN1(n15027), .IN2(n8451), .QN(n15028) );
  NAND3X0 U15962 ( .IN1(n15029), .IN2(n15030), .IN3(n15031), .QN(g26913) );
  NAND2X0 U15963 ( .IN1(n4938), .IN2(n15032), .QN(n15031) );
  NAND2X0 U15964 ( .IN1(n9453), .IN2(g1041), .QN(n15030) );
  NAND3X0 U15965 ( .IN1(n9663), .IN2(g1046), .IN3(n9335), .QN(n15029) );
  NAND2X0 U15966 ( .IN1(n15033), .IN2(n15034), .QN(n9663) );
  NAND2X0 U15967 ( .IN1(n8339), .IN2(g1008), .QN(n15034) );
  NAND3X0 U15968 ( .IN1(n15035), .IN2(n15036), .IN3(n15037), .QN(g26912) );
  NAND2X0 U15969 ( .IN1(n9453), .IN2(g921), .QN(n15037) );
  NAND3X0 U15970 ( .IN1(n11867), .IN2(n15038), .IN3(g936), .QN(n15036) );
  NAND2X0 U15971 ( .IN1(n266), .IN2(n5557), .QN(n15035) );
  INVX0 U15972 ( .INP(n15038), .ZN(n266) );
  NAND3X0 U15973 ( .IN1(g921), .IN2(g904), .IN3(g12919), .QN(n15038) );
  NAND2X0 U15974 ( .IN1(n15039), .IN2(n15040), .QN(g26910) );
  NAND2X0 U15975 ( .IN1(n15041), .IN2(g862), .QN(n15040) );
  NAND2X0 U15976 ( .IN1(n5305), .IN2(n9382), .QN(n15041) );
  NAND3X0 U15977 ( .IN1(n5305), .IN2(n9316), .IN3(n5682), .QN(n15039) );
  NAND2X0 U15978 ( .IN1(n15042), .IN2(n15043), .QN(g26909) );
  NAND2X0 U15979 ( .IN1(n9453), .IN2(g890), .QN(n15043) );
  NAND2X0 U15980 ( .IN1(n15044), .IN2(n9368), .QN(n15042) );
  NAND2X0 U15981 ( .IN1(n15045), .IN2(n15046), .QN(n15044) );
  NAND2X0 U15982 ( .IN1(n5431), .IN2(g862), .QN(n15046) );
  NAND2X0 U15983 ( .IN1(n5305), .IN2(g896), .QN(n15045) );
  NAND3X0 U15984 ( .IN1(n15047), .IN2(n15048), .IN3(n15049), .QN(g26908) );
  NAND2X0 U15985 ( .IN1(n4945), .IN2(g446), .QN(n15049) );
  NAND2X0 U15986 ( .IN1(n15050), .IN2(g872), .QN(n15048) );
  NAND2X0 U15987 ( .IN1(n9480), .IN2(g246), .QN(n15047) );
  NAND3X0 U15988 ( .IN1(n15051), .IN2(n15052), .IN3(n15053), .QN(g26907) );
  NAND2X0 U15989 ( .IN1(n4945), .IN2(g246), .QN(n15053) );
  NAND2X0 U15990 ( .IN1(n15050), .IN2(g14167), .QN(n15052) );
  NAND2X0 U15991 ( .IN1(n9444), .IN2(g269), .QN(n15051) );
  NAND3X0 U15992 ( .IN1(n15054), .IN2(n15055), .IN3(n15056), .QN(g26906) );
  NAND2X0 U15993 ( .IN1(n4945), .IN2(g269), .QN(n15056) );
  NAND2X0 U15994 ( .IN1(n15050), .IN2(g14147), .QN(n15055) );
  NAND2X0 U15995 ( .IN1(n9446), .IN2(g239), .QN(n15054) );
  NAND3X0 U15996 ( .IN1(n15057), .IN2(n15058), .IN3(n15059), .QN(g26905) );
  NAND2X0 U15997 ( .IN1(n4945), .IN2(g239), .QN(n15059) );
  NAND2X0 U15998 ( .IN1(n15050), .IN2(g14125), .QN(n15058) );
  NAND2X0 U15999 ( .IN1(n9445), .IN2(g262), .QN(n15057) );
  NAND3X0 U16000 ( .IN1(n15060), .IN2(n15061), .IN3(n15062), .QN(g26904) );
  NAND2X0 U16001 ( .IN1(n4945), .IN2(g262), .QN(n15062) );
  NAND2X0 U16002 ( .IN1(n15050), .IN2(g14096), .QN(n15061) );
  NAND2X0 U16003 ( .IN1(n9448), .IN2(g232), .QN(n15060) );
  NAND3X0 U16004 ( .IN1(n15063), .IN2(n15064), .IN3(n15065), .QN(g26903) );
  NAND2X0 U16005 ( .IN1(n4945), .IN2(g232), .QN(n15065) );
  NAND2X0 U16006 ( .IN1(n15050), .IN2(g14217), .QN(n15064) );
  NAND2X0 U16007 ( .IN1(n9449), .IN2(g255), .QN(n15063) );
  NAND3X0 U16008 ( .IN1(n15066), .IN2(n15067), .IN3(n15068), .QN(g26902) );
  NAND2X0 U16009 ( .IN1(n4945), .IN2(g255), .QN(n15068) );
  NAND2X0 U16010 ( .IN1(n15050), .IN2(g14201), .QN(n15067) );
  NAND2X0 U16011 ( .IN1(n9447), .IN2(g225), .QN(n15066) );
  NAND3X0 U16012 ( .IN1(n15069), .IN2(n15070), .IN3(n15071), .QN(g26901) );
  NAND2X0 U16013 ( .IN1(n4945), .IN2(g225), .QN(n15071) );
  NAND2X0 U16014 ( .IN1(n15050), .IN2(g14189), .QN(n15070) );
  NOR2X0 U16015 ( .IN1(n9411), .IN2(n4946), .QN(n15050) );
  NAND3X0 U16016 ( .IN1(n5431), .IN2(g890), .IN3(n5682), .QN(n4946) );
  NAND2X0 U16017 ( .IN1(n9486), .IN2(g872), .QN(n15069) );
  NAND3X0 U16018 ( .IN1(n15072), .IN2(n15073), .IN3(n15074), .QN(g26899) );
  NAND2X0 U16019 ( .IN1(n9488), .IN2(g832), .QN(n15074) );
  NAND3X0 U16020 ( .IN1(n4518), .IN2(n15075), .IN3(g822), .QN(n15073) );
  NAND3X0 U16021 ( .IN1(n905), .IN2(n14104), .IN3(n5422), .QN(n15072) );
  INVX0 U16022 ( .INP(n15075), .ZN(n905) );
  NAND3X0 U16023 ( .IN1(g817), .IN2(g832), .IN3(n4948), .QN(n15075) );
  NAND3X0 U16024 ( .IN1(n15076), .IN2(n15077), .IN3(n15078), .QN(g26898) );
  NAND2X0 U16025 ( .IN1(n9491), .IN2(g843), .QN(n15078) );
  NAND3X0 U16026 ( .IN1(n5733), .IN2(g837), .IN3(n15079), .QN(n15077) );
  NAND2X0 U16027 ( .IN1(n15080), .IN2(n15081), .QN(n15076) );
  NAND2X0 U16028 ( .IN1(n15082), .IN2(n15083), .QN(n15081) );
  NAND2X0 U16029 ( .IN1(n8431), .IN2(n9368), .QN(n15083) );
  INVX0 U16030 ( .INP(n15084), .ZN(n15080) );
  NAND2X0 U16031 ( .IN1(n15085), .IN2(n15086), .QN(g26897) );
  NAND2X0 U16032 ( .IN1(n15087), .IN2(g753), .QN(n15086) );
  INVX0 U16033 ( .INP(n15088), .ZN(n15085) );
  NOR2X0 U16034 ( .IN1(n15087), .IN2(n5732), .QN(n15088) );
  NOR2X0 U16035 ( .IN1(n14788), .IN2(n9392), .QN(n15087) );
  INVX0 U16036 ( .INP(n15089), .ZN(n14788) );
  NAND3X0 U16037 ( .IN1(n15090), .IN2(n15091), .IN3(n15092), .QN(g26896) );
  NAND2X0 U16038 ( .IN1(n4956), .IN2(n14131), .QN(n15092) );
  NAND2X0 U16039 ( .IN1(n15093), .IN2(g29212), .QN(n15091) );
  INVX0 U16040 ( .INP(n15094), .ZN(n15090) );
  NOR2X0 U16041 ( .IN1(n15093), .IN2(n8475), .QN(n15094) );
  NOR2X0 U16042 ( .IN1(n14131), .IN2(n9392), .QN(n15093) );
  NOR4X0 U16043 ( .IN1(n14784), .IN2(n14151), .IN3(g528), .IN4(n15095), .QN(
        n14131) );
  NAND2X0 U16044 ( .IN1(n5519), .IN2(test_so54), .QN(n15095) );
  NAND3X0 U16045 ( .IN1(n15096), .IN2(n15097), .IN3(n15098), .QN(g26895) );
  NAND2X0 U16046 ( .IN1(n9490), .IN2(g562), .QN(n15098) );
  NAND3X0 U16047 ( .IN1(n2421), .IN2(n15099), .IN3(g568), .QN(n15097) );
  NAND2X0 U16048 ( .IN1(n5), .IN2(n5335), .QN(n15096) );
  INVX0 U16049 ( .INP(n15099), .ZN(n5) );
  NAND3X0 U16050 ( .IN1(n15100), .IN2(g562), .IN3(n4959), .QN(n15099) );
  NAND2X0 U16051 ( .IN1(n15101), .IN2(n15102), .QN(g26894) );
  NAND2X0 U16052 ( .IN1(n9489), .IN2(g518), .QN(n15102) );
  NAND4X0 U16053 ( .IN1(n15103), .IN2(n15104), .IN3(n14141), .IN4(n9361), .QN(
        n15101) );
  NAND2X0 U16054 ( .IN1(n14782), .IN2(g528), .QN(n15104) );
  NAND2X0 U16055 ( .IN1(n5327), .IN2(n15105), .QN(n15103) );
  NAND2X0 U16056 ( .IN1(n14782), .IN2(n14784), .QN(n15105) );
  NAND2X0 U16057 ( .IN1(g482), .IN2(g490), .QN(n14784) );
  NOR3X0 U16058 ( .IN1(g513), .IN2(n5287), .IN3(n15106), .QN(n14782) );
  NAND2X0 U16059 ( .IN1(n15107), .IN2(n15108), .QN(g26893) );
  INVX0 U16060 ( .INP(n15109), .ZN(n15108) );
  NOR2X0 U16061 ( .IN1(n9358), .IN2(n8716), .QN(n15109) );
  NAND2X0 U16062 ( .IN1(n15110), .IN2(n9368), .QN(n15107) );
  NAND2X0 U16063 ( .IN1(n15111), .IN2(n15112), .QN(n15110) );
  NAND2X0 U16064 ( .IN1(g29211), .IN2(n8886), .QN(n15112) );
  NAND2X0 U16065 ( .IN1(test_so17), .IN2(n15113), .QN(n15111) );
  NAND2X0 U16066 ( .IN1(n15114), .IN2(n15115), .QN(g26892) );
  NAND3X0 U16067 ( .IN1(n9349), .IN2(n15113), .IN3(n8886), .QN(n15115) );
  NAND2X0 U16068 ( .IN1(n8716), .IN2(n8715), .QN(n15113) );
  NAND2X0 U16069 ( .IN1(test_so17), .IN2(n9516), .QN(n15114) );
  NAND2X0 U16070 ( .IN1(n15116), .IN2(n15117), .QN(g26891) );
  INVX0 U16071 ( .INP(n15118), .ZN(n15117) );
  NOR2X0 U16072 ( .IN1(n9356), .IN2(n5860), .QN(n15118) );
  NAND3X0 U16073 ( .IN1(n9349), .IN2(g7540), .IN3(n5860), .QN(n15116) );
  NAND2X0 U16074 ( .IN1(n15119), .IN2(n15120), .QN(g26890) );
  NAND2X0 U16075 ( .IN1(n5860), .IN2(n9368), .QN(n15120) );
  INVX0 U16076 ( .INP(n15121), .ZN(n15119) );
  NOR2X0 U16077 ( .IN1(n9358), .IN2(n8715), .QN(n15121) );
  NAND2X0 U16078 ( .IN1(n15122), .IN2(n15123), .QN(g26889) );
  NAND2X0 U16079 ( .IN1(n9474), .IN2(g29211), .QN(n15123) );
  NAND4X0 U16080 ( .IN1(g329), .IN2(DFF_709_n1), .IN3(n15124), .IN4(n9362), 
        .QN(n15122) );
  NAND2X0 U16081 ( .IN1(n15125), .IN2(n15126), .QN(g26888) );
  NAND2X0 U16082 ( .IN1(n9364), .IN2(g316), .QN(n15126) );
  NAND2X0 U16083 ( .IN1(n9476), .IN2(g29216), .QN(n15125) );
  NAND3X0 U16084 ( .IN1(n15127), .IN2(n15128), .IN3(n15129), .QN(g26887) );
  NAND2X0 U16085 ( .IN1(n9475), .IN2(g336), .QN(n15128) );
  NAND3X0 U16086 ( .IN1(n5317), .IN2(g324), .IN3(n9335), .QN(n15127) );
  NAND3X0 U16087 ( .IN1(n15130), .IN2(n15131), .IN3(n15132), .QN(g26886) );
  NAND2X0 U16088 ( .IN1(n15133), .IN2(n15134), .QN(n15132) );
  INVX0 U16089 ( .INP(n15129), .ZN(n15133) );
  NAND3X0 U16090 ( .IN1(n15124), .IN2(g336), .IN3(n9335), .QN(n15131) );
  NAND2X0 U16091 ( .IN1(n9479), .IN2(g311), .QN(n15130) );
  NAND2X0 U16092 ( .IN1(n15135), .IN2(n15136), .QN(g26884) );
  NAND2X0 U16093 ( .IN1(n9478), .IN2(g329), .QN(n15136) );
  NAND2X0 U16094 ( .IN1(n15137), .IN2(n9368), .QN(n15135) );
  NAND2X0 U16095 ( .IN1(n15138), .IN2(n15139), .QN(n15137) );
  NAND4X0 U16096 ( .IN1(n5766), .IN2(n5456), .IN3(n5282), .IN4(n5317), .QN(
        n15139) );
  NAND2X0 U16097 ( .IN1(n15134), .IN2(n15140), .QN(n15138) );
  NAND3X0 U16098 ( .IN1(n15141), .IN2(n15142), .IN3(n5456), .QN(n15140) );
  NAND2X0 U16099 ( .IN1(n5824), .IN2(g311), .QN(n15142) );
  NAND2X0 U16100 ( .IN1(g305), .IN2(g336), .QN(n15141) );
  NAND2X0 U16101 ( .IN1(n15143), .IN2(n15144), .QN(g26883) );
  NAND2X0 U16102 ( .IN1(n9477), .IN2(g324), .QN(n15144) );
  NAND2X0 U16103 ( .IN1(n15134), .IN2(n9368), .QN(n15143) );
  INVX0 U16104 ( .INP(n15124), .ZN(n15134) );
  NAND2X0 U16105 ( .IN1(n15145), .IN2(n15146), .QN(n15124) );
  NAND2X0 U16106 ( .IN1(n5282), .IN2(g324), .QN(n15146) );
  NAND2X0 U16107 ( .IN1(n5827), .IN2(n5317), .QN(n15145) );
  NAND3X0 U16108 ( .IN1(n15147), .IN2(n15148), .IN3(n15129), .QN(g26882) );
  NAND2X0 U16109 ( .IN1(n9363), .IN2(g305), .QN(n15129) );
  NAND2X0 U16110 ( .IN1(n9363), .IN2(g311), .QN(n15148) );
  NAND2X0 U16111 ( .IN1(n9481), .IN2(g316), .QN(n15147) );
  NAND2X0 U16112 ( .IN1(n15149), .IN2(n15150), .QN(g26881) );
  NAND2X0 U16113 ( .IN1(g6744), .IN2(n9368), .QN(n15150) );
  NAND2X0 U16114 ( .IN1(n9482), .IN2(g305), .QN(n15149) );
  NAND3X0 U16115 ( .IN1(n10216), .IN2(n9316), .IN3(n10217), .QN(g26877) );
  NAND4X0 U16116 ( .IN1(n5620), .IN2(n5619), .IN3(n15151), .IN4(n15152), .QN(
        n10217) );
  NOR4X0 U16117 ( .IN1(test_so40), .IN2(g2357), .IN3(g2338), .IN4(g2606), .QN(
        n15152) );
  NOR2X0 U16118 ( .IN1(g2491), .IN2(g2223), .QN(n15151) );
  NAND4X0 U16119 ( .IN1(n5833), .IN2(n5832), .IN3(n15153), .IN4(n15154), .QN(
        n10216) );
  NOR4X0 U16120 ( .IN1(test_so75), .IN2(g1664), .IN3(g1913), .IN4(g1932), .QN(
        n15154) );
  NOR2X0 U16121 ( .IN1(g1779), .IN2(g2047), .QN(n15153) );
  INVX0 U16122 ( .INP(n15155), .ZN(g26876) );
  NOR2X0 U16123 ( .IN1(n10177), .IN2(n10234), .QN(n15155) );
  INVX0 U16124 ( .INP(n10181), .ZN(n10234) );
  NAND4X0 U16125 ( .IN1(n15966), .IN2(n5892), .IN3(n15156), .IN4(n15157), .QN(
        n10181) );
  NOR4X0 U16126 ( .IN1(g1710), .IN2(g1978), .IN3(g1844), .IN4(g2112), .QN(
        n15157) );
  NOR2X0 U16127 ( .IN1(g1992), .IN2(g2126), .QN(n15156) );
  NAND2X0 U16128 ( .IN1(n15158), .IN2(n9368), .QN(n10177) );
  NAND4X0 U16129 ( .IN1(n15960), .IN2(n15967), .IN3(n15159), .IN4(n15160), 
        .QN(n15158) );
  NOR4X0 U16130 ( .IN1(test_so31), .IN2(g2671), .IN3(g2269), .IN4(g2537), .QN(
        n15160) );
  NOR2X0 U16131 ( .IN1(n9324), .IN2(n9295), .QN(n15159) );
  INVX0 U16132 ( .INP(n15161), .ZN(g26875) );
  NOR2X0 U16133 ( .IN1(n10178), .IN2(n10238), .QN(n15161) );
  INVX0 U16134 ( .INP(n10182), .ZN(n10238) );
  NAND4X0 U16135 ( .IN1(n5628), .IN2(n5413), .IN3(n5315), .IN4(n5280), .QN(
        n10182) );
  NAND2X0 U16136 ( .IN1(n15162), .IN2(n9369), .QN(n10178) );
  NAND4X0 U16137 ( .IN1(n5631), .IN2(n5414), .IN3(n5316), .IN4(n5281), .QN(
        n15162) );
  NAND2X0 U16138 ( .IN1(n15163), .IN2(n15164), .QN(g25764) );
  NAND2X0 U16139 ( .IN1(n12468), .IN2(g6505), .QN(n15164) );
  NAND2X0 U16140 ( .IN1(n15165), .IN2(g6541), .QN(n15163) );
  NAND3X0 U16141 ( .IN1(n15166), .IN2(n15167), .IN3(n15168), .QN(g25763) );
  INVX0 U16142 ( .INP(n15169), .ZN(n15168) );
  NOR2X0 U16143 ( .IN1(n15165), .IN2(n5884), .QN(n15169) );
  NAND2X0 U16144 ( .IN1(n15170), .IN2(g6533), .QN(n15167) );
  NAND2X0 U16145 ( .IN1(n15171), .IN2(n9368), .QN(n15170) );
  NAND2X0 U16146 ( .IN1(n11370), .IN2(g6527), .QN(n15171) );
  NAND4X0 U16147 ( .IN1(n11370), .IN2(n9356), .IN3(n5659), .IN4(n5445), .QN(
        n15166) );
  NAND2X0 U16148 ( .IN1(n15172), .IN2(n15173), .QN(g25762) );
  NAND2X0 U16149 ( .IN1(n12468), .IN2(g6533), .QN(n15173) );
  NAND2X0 U16150 ( .IN1(n15165), .IN2(g6527), .QN(n15172) );
  NAND3X0 U16151 ( .IN1(n15174), .IN2(n15175), .IN3(n15176), .QN(g25761) );
  NAND2X0 U16152 ( .IN1(n12468), .IN2(g6513), .QN(n15176) );
  INVX0 U16153 ( .INP(n15165), .ZN(n12468) );
  NAND2X0 U16154 ( .IN1(n13567), .IN2(n9368), .QN(n15165) );
  NAND3X0 U16155 ( .IN1(n5426), .IN2(n11370), .IN3(n9335), .QN(n15175) );
  INVX0 U16156 ( .INP(n13567), .ZN(n11370) );
  NAND2X0 U16157 ( .IN1(n9806), .IN2(g6561), .QN(n13567) );
  NOR2X0 U16158 ( .IN1(n5386), .IN2(n5563), .QN(n9806) );
  NAND2X0 U16159 ( .IN1(n9452), .IN2(g6509), .QN(n15174) );
  NAND2X0 U16160 ( .IN1(n15177), .IN2(n15178), .QN(g25758) );
  INVX0 U16161 ( .INP(n15179), .ZN(n15178) );
  NOR2X0 U16162 ( .IN1(n9359), .IN2(n8805), .QN(n15179) );
  NAND3X0 U16163 ( .IN1(n8373), .IN2(n15180), .IN3(n9335), .QN(n15177) );
  NAND2X0 U16164 ( .IN1(n5990), .IN2(n15181), .QN(n15180) );
  NAND2X0 U16165 ( .IN1(n8805), .IN2(g9743), .QN(n15181) );
  NAND2X0 U16166 ( .IN1(n15182), .IN2(n15183), .QN(g25757) );
  NAND2X0 U16167 ( .IN1(n9363), .IN2(g6727), .QN(n15183) );
  INVX0 U16168 ( .INP(n15184), .ZN(n15182) );
  NOR2X0 U16169 ( .IN1(n9359), .IN2(n5990), .QN(n15184) );
  NOR2X0 U16170 ( .IN1(n9413), .IN2(n5563), .QN(g25756) );
  NAND2X0 U16171 ( .IN1(n15185), .IN2(n15186), .QN(g25750) );
  NAND2X0 U16172 ( .IN1(n12552), .IN2(g6159), .QN(n15186) );
  NAND2X0 U16173 ( .IN1(n15187), .IN2(g6195), .QN(n15185) );
  NAND3X0 U16174 ( .IN1(n15188), .IN2(n15189), .IN3(n15190), .QN(g25749) );
  INVX0 U16175 ( .INP(n15191), .ZN(n15190) );
  NOR2X0 U16176 ( .IN1(n15187), .IN2(n5888), .QN(n15191) );
  NAND2X0 U16177 ( .IN1(n15192), .IN2(g6187), .QN(n15189) );
  NAND2X0 U16178 ( .IN1(n15193), .IN2(n9369), .QN(n15192) );
  NAND2X0 U16179 ( .IN1(n12553), .IN2(g6181), .QN(n15193) );
  NAND4X0 U16180 ( .IN1(n12553), .IN2(n9355), .IN3(n5667), .IN4(n5453), .QN(
        n15188) );
  NAND2X0 U16181 ( .IN1(n15194), .IN2(n15195), .QN(g25748) );
  NAND2X0 U16182 ( .IN1(n12552), .IN2(g6187), .QN(n15195) );
  NAND2X0 U16183 ( .IN1(n15187), .IN2(g6181), .QN(n15194) );
  INVX0 U16184 ( .INP(n12552), .ZN(n15187) );
  NAND3X0 U16185 ( .IN1(n15196), .IN2(n15197), .IN3(n15198), .QN(g25747) );
  NAND2X0 U16186 ( .IN1(n12552), .IN2(g6167), .QN(n15198) );
  NOR2X0 U16187 ( .IN1(n12553), .IN2(n9390), .QN(n12552) );
  NAND3X0 U16188 ( .IN1(n5430), .IN2(n12553), .IN3(n9335), .QN(n15197) );
  NOR2X0 U16189 ( .IN1(n52), .IN2(n5651), .QN(n12553) );
  INVX0 U16190 ( .INP(n12573), .ZN(n52) );
  NOR2X0 U16191 ( .IN1(n5385), .IN2(n5568), .QN(n12573) );
  NAND2X0 U16192 ( .IN1(n9452), .IN2(g6163), .QN(n15196) );
  NAND2X0 U16193 ( .IN1(n15199), .IN2(n15200), .QN(g25744) );
  INVX0 U16194 ( .INP(n15201), .ZN(n15200) );
  NOR2X0 U16195 ( .IN1(n9359), .IN2(n8806), .QN(n15201) );
  NAND3X0 U16196 ( .IN1(n8369), .IN2(n15202), .IN3(n9335), .QN(n15199) );
  NAND2X0 U16197 ( .IN1(n5988), .IN2(n15203), .QN(n15202) );
  NAND2X0 U16198 ( .IN1(test_so92), .IN2(n8806), .QN(n15203) );
  NAND2X0 U16199 ( .IN1(n15204), .IN2(n15205), .QN(g25743) );
  NAND2X0 U16200 ( .IN1(test_so69), .IN2(n9369), .QN(n15205) );
  INVX0 U16201 ( .INP(n15206), .ZN(n15204) );
  NOR2X0 U16202 ( .IN1(n9359), .IN2(n5988), .QN(n15206) );
  NOR2X0 U16203 ( .IN1(n9414), .IN2(n5568), .QN(g25742) );
  NAND2X0 U16204 ( .IN1(n15207), .IN2(n15208), .QN(g25736) );
  NAND2X0 U16205 ( .IN1(g5813), .IN2(n12638), .QN(n15208) );
  NAND2X0 U16206 ( .IN1(n15209), .IN2(g5849), .QN(n15207) );
  NAND3X0 U16207 ( .IN1(n15210), .IN2(n15211), .IN3(n15212), .QN(g25735) );
  NAND2X0 U16208 ( .IN1(test_so83), .IN2(n12638), .QN(n15212) );
  NAND2X0 U16209 ( .IN1(n15213), .IN2(g5841), .QN(n15211) );
  NAND2X0 U16210 ( .IN1(n15214), .IN2(n9369), .QN(n15213) );
  NAND2X0 U16211 ( .IN1(n12639), .IN2(g5835), .QN(n15214) );
  NAND4X0 U16212 ( .IN1(n12639), .IN2(n9355), .IN3(n5663), .IN4(n5449), .QN(
        n15210) );
  NAND2X0 U16213 ( .IN1(n15215), .IN2(n15216), .QN(g25734) );
  NAND2X0 U16214 ( .IN1(n12638), .IN2(g5841), .QN(n15216) );
  NAND2X0 U16215 ( .IN1(n15209), .IN2(g5835), .QN(n15215) );
  INVX0 U16216 ( .INP(n12638), .ZN(n15209) );
  NAND3X0 U16217 ( .IN1(n15217), .IN2(n15218), .IN3(n15219), .QN(g25733) );
  NAND2X0 U16218 ( .IN1(n12638), .IN2(g5821), .QN(n15219) );
  NOR2X0 U16219 ( .IN1(n12639), .IN2(n9389), .QN(n12638) );
  NAND3X0 U16220 ( .IN1(n5429), .IN2(n12639), .IN3(n9335), .QN(n15218) );
  NOR2X0 U16221 ( .IN1(n733), .IN2(n5649), .QN(n12639) );
  INVX0 U16222 ( .INP(n12659), .ZN(n733) );
  NOR2X0 U16223 ( .IN1(n8872), .IN2(n5388), .QN(n12659) );
  NAND2X0 U16224 ( .IN1(n9452), .IN2(g5817), .QN(n15217) );
  NAND2X0 U16225 ( .IN1(n15220), .IN2(n15221), .QN(g25730) );
  INVX0 U16226 ( .INP(n15222), .ZN(n15221) );
  NOR2X0 U16227 ( .IN1(n9360), .IN2(n8800), .QN(n15222) );
  NAND3X0 U16228 ( .IN1(n8379), .IN2(n15223), .IN3(n9335), .QN(n15220) );
  NAND2X0 U16229 ( .IN1(n5996), .IN2(n15224), .QN(n15223) );
  NAND2X0 U16230 ( .IN1(n8800), .IN2(g9617), .QN(n15224) );
  NAND2X0 U16231 ( .IN1(n15225), .IN2(n15226), .QN(g25729) );
  NAND2X0 U16232 ( .IN1(n9362), .IN2(g6035), .QN(n15226) );
  INVX0 U16233 ( .INP(n15227), .ZN(n15225) );
  NOR2X0 U16234 ( .IN1(n9359), .IN2(n5996), .QN(n15227) );
  NOR2X0 U16235 ( .IN1(n8872), .IN2(n9389), .QN(g25728) );
  NAND2X0 U16236 ( .IN1(n15228), .IN2(n15229), .QN(g25722) );
  NAND2X0 U16237 ( .IN1(n12724), .IN2(g5467), .QN(n15229) );
  NAND2X0 U16238 ( .IN1(n15230), .IN2(g5503), .QN(n15228) );
  NAND3X0 U16239 ( .IN1(n15231), .IN2(n15232), .IN3(n15233), .QN(g25721) );
  INVX0 U16240 ( .INP(n15234), .ZN(n15233) );
  NOR2X0 U16241 ( .IN1(n15230), .IN2(n5885), .QN(n15234) );
  NAND2X0 U16242 ( .IN1(n15235), .IN2(g5495), .QN(n15232) );
  NAND2X0 U16243 ( .IN1(n15236), .IN2(n9369), .QN(n15235) );
  NAND2X0 U16244 ( .IN1(n11354), .IN2(g5489), .QN(n15236) );
  NAND4X0 U16245 ( .IN1(n11354), .IN2(n9355), .IN3(n5660), .IN4(n5446), .QN(
        n15231) );
  NAND2X0 U16246 ( .IN1(n15237), .IN2(n15238), .QN(g25720) );
  NAND2X0 U16247 ( .IN1(n12724), .IN2(g5495), .QN(n15238) );
  NAND2X0 U16248 ( .IN1(n15230), .IN2(g5489), .QN(n15237) );
  NAND3X0 U16249 ( .IN1(n15239), .IN2(n15240), .IN3(n15241), .QN(g25719) );
  NAND2X0 U16250 ( .IN1(n12724), .IN2(g5475), .QN(n15241) );
  INVX0 U16251 ( .INP(n15230), .ZN(n12724) );
  NAND2X0 U16252 ( .IN1(n13668), .IN2(n9369), .QN(n15230) );
  NAND3X0 U16253 ( .IN1(n5425), .IN2(n11354), .IN3(n9335), .QN(n15240) );
  INVX0 U16254 ( .INP(n13668), .ZN(n11354) );
  NAND2X0 U16255 ( .IN1(n9657), .IN2(g5523), .QN(n13668) );
  NOR2X0 U16256 ( .IN1(n5389), .IN2(n5566), .QN(n9657) );
  NAND2X0 U16257 ( .IN1(n9452), .IN2(g5471), .QN(n15239) );
  NAND2X0 U16258 ( .IN1(n15242), .IN2(n15243), .QN(g25716) );
  INVX0 U16259 ( .INP(n15244), .ZN(n15243) );
  NOR2X0 U16260 ( .IN1(n9360), .IN2(n8802), .QN(n15244) );
  NAND3X0 U16261 ( .IN1(n15245), .IN2(n8375), .IN3(n9334), .QN(n15242) );
  NAND2X0 U16262 ( .IN1(n5992), .IN2(n15246), .QN(n15245) );
  NAND2X0 U16263 ( .IN1(n8802), .IN2(g9555), .QN(n15246) );
  NAND2X0 U16264 ( .IN1(n15247), .IN2(n15248), .QN(g25715) );
  NAND2X0 U16265 ( .IN1(n9362), .IN2(g5689), .QN(n15248) );
  INVX0 U16266 ( .INP(n15249), .ZN(n15247) );
  NOR2X0 U16267 ( .IN1(n9360), .IN2(n5992), .QN(n15249) );
  NOR2X0 U16268 ( .IN1(n9416), .IN2(n5566), .QN(g25714) );
  NAND2X0 U16269 ( .IN1(n15250), .IN2(n15251), .QN(g25708) );
  NAND2X0 U16270 ( .IN1(n12808), .IN2(g5120), .QN(n15251) );
  NAND2X0 U16271 ( .IN1(n15252), .IN2(g5156), .QN(n15250) );
  NAND3X0 U16272 ( .IN1(n15253), .IN2(n15254), .IN3(n15255), .QN(g25707) );
  INVX0 U16273 ( .INP(n15256), .ZN(n15255) );
  NOR2X0 U16274 ( .IN1(n15252), .IN2(n5883), .QN(n15256) );
  NAND2X0 U16275 ( .IN1(test_so98), .IN2(n15257), .QN(n15254) );
  NAND2X0 U16276 ( .IN1(n15258), .IN2(n9370), .QN(n15257) );
  NAND2X0 U16277 ( .IN1(g32975), .IN2(g5142), .QN(n15258) );
  NAND4X0 U16278 ( .IN1(g32975), .IN2(n9356), .IN3(n5658), .IN4(n8900), .QN(
        n15253) );
  NAND2X0 U16279 ( .IN1(n15259), .IN2(n15260), .QN(g25706) );
  NAND2X0 U16280 ( .IN1(test_so98), .IN2(n12808), .QN(n15260) );
  NAND2X0 U16281 ( .IN1(n15252), .IN2(g5142), .QN(n15259) );
  NAND3X0 U16282 ( .IN1(n15261), .IN2(n15262), .IN3(n15263), .QN(g25705) );
  NAND2X0 U16283 ( .IN1(test_so96), .IN2(n12808), .QN(n15263) );
  INVX0 U16284 ( .INP(n15252), .ZN(n12808) );
  NAND2X0 U16285 ( .IN1(n13702), .IN2(n9370), .QN(n15252) );
  NAND3X0 U16286 ( .IN1(g32975), .IN2(n8877), .IN3(n9334), .QN(n15262) );
  INVX0 U16287 ( .INP(n13702), .ZN(g32975) );
  NAND2X0 U16288 ( .IN1(n9800), .IN2(g5176), .QN(n13702) );
  NOR2X0 U16289 ( .IN1(n5384), .IN2(n5567), .QN(n9800) );
  NAND2X0 U16290 ( .IN1(n9452), .IN2(g5124), .QN(n15261) );
  NOR2X0 U16291 ( .IN1(n8412), .IN2(n15264), .QN(g25704) );
  NOR2X0 U16292 ( .IN1(n9417), .IN2(g5069), .QN(n15264) );
  NAND2X0 U16293 ( .IN1(n15265), .IN2(n15266), .QN(g25703) );
  NAND2X0 U16294 ( .IN1(n9452), .IN2(g5112), .QN(n15266) );
  NAND3X0 U16295 ( .IN1(n5689), .IN2(n15267), .IN3(n9334), .QN(n15265) );
  INVX0 U16296 ( .INP(n15268), .ZN(n15267) );
  NOR2X0 U16297 ( .IN1(g5022), .IN2(n15269), .QN(n15268) );
  NOR2X0 U16298 ( .IN1(g5112), .IN2(n5690), .QN(n15269) );
  NAND2X0 U16299 ( .IN1(n15270), .IN2(n15271), .QN(g25702) );
  NAND2X0 U16300 ( .IN1(test_so32), .IN2(n9514), .QN(n15271) );
  NAND3X0 U16301 ( .IN1(n5690), .IN2(n15272), .IN3(n9334), .QN(n15270) );
  INVX0 U16302 ( .INP(n15273), .ZN(n15272) );
  NOR2X0 U16303 ( .IN1(g5062), .IN2(n15274), .QN(n15273) );
  NOR2X0 U16304 ( .IN1(n5689), .IN2(test_so32), .QN(n15274) );
  NAND2X0 U16305 ( .IN1(n15275), .IN2(n15276), .QN(g25701) );
  NAND2X0 U16306 ( .IN1(test_so10), .IN2(n9370), .QN(n15276) );
  NAND2X0 U16307 ( .IN1(n9452), .IN2(g5062), .QN(n15275) );
  NOR2X0 U16308 ( .IN1(n9417), .IN2(n5567), .QN(g25700) );
  NAND3X0 U16309 ( .IN1(n15277), .IN2(n15278), .IN3(n15279), .QN(g25699) );
  NAND2X0 U16310 ( .IN1(n9451), .IN2(g5097), .QN(n15279) );
  INVX0 U16311 ( .INP(n15280), .ZN(n15278) );
  NOR3X0 U16312 ( .IN1(n9385), .IN2(n5014), .IN3(n5669), .QN(n15280) );
  NAND2X0 U16313 ( .IN1(n5014), .IN2(n5669), .QN(n15277) );
  NAND3X0 U16314 ( .IN1(n15281), .IN2(n15282), .IN3(n15283), .QN(g25698) );
  NAND2X0 U16315 ( .IN1(n9451), .IN2(g5092), .QN(n15283) );
  NAND3X0 U16316 ( .IN1(n9349), .IN2(n15284), .IN3(g5097), .QN(n15282) );
  INVX0 U16317 ( .INP(n5016), .ZN(n15284) );
  NAND2X0 U16318 ( .IN1(n5016), .IN2(n5753), .QN(n15281) );
  NAND2X0 U16319 ( .IN1(n15285), .IN2(n15286), .QN(g25697) );
  NAND2X0 U16320 ( .IN1(n15287), .IN2(g5084), .QN(n15286) );
  NAND2X0 U16321 ( .IN1(n9363), .IN2(g5092), .QN(n15287) );
  NAND3X0 U16322 ( .IN1(n9349), .IN2(g5092), .IN3(n5681), .QN(n15285) );
  NAND3X0 U16323 ( .IN1(n15288), .IN2(n15289), .IN3(n15290), .QN(g25696) );
  NAND3X0 U16324 ( .IN1(n9349), .IN2(g5077), .IN3(n8412), .QN(n15290) );
  INVX0 U16325 ( .INP(n15291), .ZN(n15289) );
  NOR2X0 U16326 ( .IN1(n15292), .IN2(n5893), .QN(n15291) );
  NAND3X0 U16327 ( .IN1(n15292), .IN2(n15293), .IN3(n5893), .QN(n15288) );
  NAND2X0 U16328 ( .IN1(n8411), .IN2(g5077), .QN(n15293) );
  NOR2X0 U16329 ( .IN1(g5084), .IN2(n9387), .QN(n15292) );
  NOR2X0 U16330 ( .IN1(n5455), .IN2(n15294), .QN(g25695) );
  NOR3X0 U16331 ( .IN1(n9385), .IN2(n15295), .IN3(n15296), .QN(n15294) );
  INVX0 U16332 ( .INP(n15297), .ZN(n15296) );
  NAND2X0 U16333 ( .IN1(n5681), .IN2(n8412), .QN(n15297) );
  NOR2X0 U16334 ( .IN1(n5681), .IN2(g5069), .QN(n15295) );
  NAND2X0 U16335 ( .IN1(n15298), .IN2(n15299), .QN(g25691) );
  NAND2X0 U16336 ( .IN1(n8852), .IN2(n15300), .QN(n15299) );
  NAND4X0 U16337 ( .IN1(n5416), .IN2(test_so11), .IN3(n5711), .IN4(n15301), 
        .QN(n15300) );
  INVX0 U16338 ( .INP(n15302), .ZN(n15301) );
  NAND4X0 U16339 ( .IN1(g4098), .IN2(n11355), .IN3(n5612), .IN4(n8446), .QN(
        n15302) );
  NOR2X0 U16340 ( .IN1(g4093), .IN2(n5480), .QN(n11355) );
  NAND2X0 U16341 ( .IN1(n9451), .IN2(g4125), .QN(n15298) );
  NAND2X0 U16342 ( .IN1(n15303), .IN2(n15304), .QN(g25690) );
  NAND2X0 U16343 ( .IN1(n9451), .IN2(g4169), .QN(n15304) );
  NAND3X0 U16344 ( .IN1(n8707), .IN2(g25689), .IN3(n9334), .QN(n15303) );
  NAND3X0 U16345 ( .IN1(n15305), .IN2(n15306), .IN3(n15307), .QN(g25687) );
  NAND2X0 U16346 ( .IN1(n9451), .IN2(g4057), .QN(n15307) );
  NAND3X0 U16347 ( .IN1(n9808), .IN2(g4169), .IN3(n5612), .QN(n15306) );
  NOR2X0 U16348 ( .IN1(n5711), .IN2(n5416), .QN(n9808) );
  NAND2X0 U16349 ( .IN1(n5026), .IN2(n12912), .QN(n15305) );
  NAND2X0 U16350 ( .IN1(n15308), .IN2(n15309), .QN(g25686) );
  NAND2X0 U16351 ( .IN1(n15310), .IN2(g4064), .QN(n15309) );
  NAND2X0 U16352 ( .IN1(n15311), .IN2(n9370), .QN(n15310) );
  NAND2X0 U16353 ( .IN1(n5711), .IN2(g4169), .QN(n15311) );
  NAND3X0 U16354 ( .IN1(n12912), .IN2(g4057), .IN3(n5416), .QN(n15308) );
  NOR2X0 U16355 ( .IN1(n9420), .IN2(n5729), .QN(n12912) );
  NAND3X0 U16356 ( .IN1(n15312), .IN2(n15313), .IN3(n12032), .QN(g25685) );
  INVX0 U16357 ( .INP(n8852), .ZN(n12032) );
  NOR2X0 U16358 ( .IN1(g4169), .IN2(n9387), .QN(n8852) );
  NAND2X0 U16359 ( .IN1(n5416), .IN2(n9371), .QN(n15313) );
  INVX0 U16360 ( .INP(n15314), .ZN(n15312) );
  NOR2X0 U16361 ( .IN1(n9359), .IN2(n8820), .QN(n15314) );
  NAND2X0 U16362 ( .IN1(n15315), .IN2(n15316), .QN(g25684) );
  NAND2X0 U16363 ( .IN1(n12916), .IN2(g3813), .QN(n15316) );
  NAND2X0 U16364 ( .IN1(n15317), .IN2(g3849), .QN(n15315) );
  NAND3X0 U16365 ( .IN1(n15318), .IN2(n15319), .IN3(n15320), .QN(g25683) );
  INVX0 U16366 ( .INP(n15321), .ZN(n15320) );
  NOR2X0 U16367 ( .IN1(n15317), .IN2(n5886), .QN(n15321) );
  NAND2X0 U16368 ( .IN1(test_so97), .IN2(n15322), .QN(n15319) );
  NAND2X0 U16369 ( .IN1(n15323), .IN2(n9371), .QN(n15322) );
  NAND2X0 U16370 ( .IN1(n12917), .IN2(g3835), .QN(n15323) );
  NAND4X0 U16371 ( .IN1(n12917), .IN2(n9356), .IN3(n5662), .IN4(n8901), .QN(
        n15318) );
  NAND2X0 U16372 ( .IN1(n15324), .IN2(n15325), .QN(g25682) );
  NAND2X0 U16373 ( .IN1(test_so97), .IN2(n12916), .QN(n15325) );
  NAND2X0 U16374 ( .IN1(n15317), .IN2(g3835), .QN(n15324) );
  INVX0 U16375 ( .INP(n12916), .ZN(n15317) );
  NAND3X0 U16376 ( .IN1(n15326), .IN2(n15327), .IN3(n15328), .QN(g25681) );
  NAND2X0 U16377 ( .IN1(n12916), .IN2(g3821), .QN(n15328) );
  NOR2X0 U16378 ( .IN1(n12917), .IN2(n9386), .QN(n12916) );
  NAND3X0 U16379 ( .IN1(n5428), .IN2(n12917), .IN3(n9342), .QN(n15327) );
  NOR2X0 U16380 ( .IN1(n8868), .IN2(n850), .QN(n12917) );
  INVX0 U16381 ( .INP(n12937), .ZN(n850) );
  NOR2X0 U16382 ( .IN1(n5387), .IN2(n5564), .QN(n12937) );
  NAND2X0 U16383 ( .IN1(n9451), .IN2(g3817), .QN(n15326) );
  NAND2X0 U16384 ( .IN1(n15329), .IN2(n15330), .QN(g25678) );
  INVX0 U16385 ( .INP(n15331), .ZN(n15330) );
  NOR2X0 U16386 ( .IN1(n9359), .IN2(n8801), .QN(n15331) );
  NAND3X0 U16387 ( .IN1(n8376), .IN2(n15332), .IN3(n9334), .QN(n15329) );
  NAND2X0 U16388 ( .IN1(n5994), .IN2(n15333), .QN(n15332) );
  NAND2X0 U16389 ( .IN1(n8801), .IN2(g8344), .QN(n15333) );
  NAND2X0 U16390 ( .IN1(n15334), .IN2(n15335), .QN(g25677) );
  NAND2X0 U16391 ( .IN1(n9363), .IN2(g4040), .QN(n15335) );
  INVX0 U16392 ( .INP(n15336), .ZN(n15334) );
  NOR2X0 U16393 ( .IN1(n9359), .IN2(n5994), .QN(n15336) );
  NOR2X0 U16394 ( .IN1(n9419), .IN2(n5564), .QN(g25676) );
  NAND2X0 U16395 ( .IN1(n15337), .IN2(n15338), .QN(g25670) );
  NAND2X0 U16396 ( .IN1(n13002), .IN2(g3462), .QN(n15338) );
  NAND2X0 U16397 ( .IN1(n15339), .IN2(g3498), .QN(n15337) );
  NAND3X0 U16398 ( .IN1(n15340), .IN2(n15341), .IN3(n15342), .QN(g25669) );
  INVX0 U16399 ( .INP(n15343), .ZN(n15342) );
  NOR2X0 U16400 ( .IN1(n15339), .IN2(n5889), .QN(n15343) );
  NAND2X0 U16401 ( .IN1(n15344), .IN2(g3490), .QN(n15341) );
  NAND2X0 U16402 ( .IN1(n15345), .IN2(n9371), .QN(n15344) );
  NAND2X0 U16403 ( .IN1(n13003), .IN2(g3484), .QN(n15345) );
  NAND4X0 U16404 ( .IN1(n13003), .IN2(n9355), .IN3(n5668), .IN4(n5454), .QN(
        n15340) );
  NAND2X0 U16405 ( .IN1(n15346), .IN2(n15347), .QN(g25668) );
  NAND2X0 U16406 ( .IN1(n13002), .IN2(g3490), .QN(n15347) );
  NAND2X0 U16407 ( .IN1(n15339), .IN2(g3484), .QN(n15346) );
  INVX0 U16408 ( .INP(n13002), .ZN(n15339) );
  NAND3X0 U16409 ( .IN1(n15348), .IN2(n15349), .IN3(n15350), .QN(g25667) );
  NAND2X0 U16410 ( .IN1(n13002), .IN2(g3470), .QN(n15350) );
  NOR2X0 U16411 ( .IN1(n13003), .IN2(n9388), .QN(n13002) );
  NAND3X0 U16412 ( .IN1(n5424), .IN2(n13003), .IN3(n9335), .QN(n15349) );
  NOR2X0 U16413 ( .IN1(n439), .IN2(n5645), .QN(n13003) );
  INVX0 U16414 ( .INP(n13023), .ZN(n439) );
  NOR2X0 U16415 ( .IN1(n5383), .IN2(n5569), .QN(n13023) );
  NAND2X0 U16416 ( .IN1(n9451), .IN2(g3466), .QN(n15348) );
  NAND2X0 U16417 ( .IN1(n15351), .IN2(n15352), .QN(g25664) );
  INVX0 U16418 ( .INP(n15353), .ZN(n15352) );
  NOR2X0 U16419 ( .IN1(n9358), .IN2(n8807), .QN(n15353) );
  NAND3X0 U16420 ( .IN1(n8359), .IN2(n15354), .IN3(n9335), .QN(n15351) );
  NAND2X0 U16421 ( .IN1(n5986), .IN2(n15355), .QN(n15354) );
  NAND2X0 U16422 ( .IN1(n8807), .IN2(g8279), .QN(n15355) );
  NAND2X0 U16423 ( .IN1(n15356), .IN2(n15357), .QN(g25663) );
  NAND2X0 U16424 ( .IN1(n9363), .IN2(g3689), .QN(n15357) );
  INVX0 U16425 ( .INP(n15358), .ZN(n15356) );
  NOR2X0 U16426 ( .IN1(n9358), .IN2(n5986), .QN(n15358) );
  NOR2X0 U16427 ( .IN1(n9418), .IN2(n5569), .QN(g25662) );
  NAND2X0 U16428 ( .IN1(n15359), .IN2(n15360), .QN(g25656) );
  NAND2X0 U16429 ( .IN1(n13088), .IN2(g3111), .QN(n15360) );
  NAND2X0 U16430 ( .IN1(n15361), .IN2(g3147), .QN(n15359) );
  NAND3X0 U16431 ( .IN1(n15362), .IN2(n15363), .IN3(n15364), .QN(g25655) );
  INVX0 U16432 ( .INP(n15365), .ZN(n15364) );
  NOR2X0 U16433 ( .IN1(n15361), .IN2(n5882), .QN(n15365) );
  NAND2X0 U16434 ( .IN1(n15366), .IN2(g3139), .QN(n15363) );
  NAND2X0 U16435 ( .IN1(n15367), .IN2(n9371), .QN(n15366) );
  NAND2X0 U16436 ( .IN1(n11365), .IN2(g3133), .QN(n15367) );
  NAND4X0 U16437 ( .IN1(n11365), .IN2(n9355), .IN3(n5661), .IN4(n5447), .QN(
        n15362) );
  NAND2X0 U16438 ( .IN1(n15368), .IN2(n15369), .QN(g25654) );
  NAND2X0 U16439 ( .IN1(n13088), .IN2(g3139), .QN(n15369) );
  NAND2X0 U16440 ( .IN1(n15361), .IN2(g3133), .QN(n15368) );
  NAND3X0 U16441 ( .IN1(n15370), .IN2(n15371), .IN3(n15372), .QN(g25653) );
  NAND2X0 U16442 ( .IN1(n13088), .IN2(g3119), .QN(n15372) );
  INVX0 U16443 ( .INP(n15361), .ZN(n13088) );
  NAND2X0 U16444 ( .IN1(n13806), .IN2(n9371), .QN(n15361) );
  NAND3X0 U16445 ( .IN1(n5423), .IN2(n11365), .IN3(n9337), .QN(n15371) );
  INVX0 U16446 ( .INP(n13806), .ZN(n11365) );
  NAND2X0 U16447 ( .IN1(n9686), .IN2(g3167), .QN(n13806) );
  NOR2X0 U16448 ( .IN1(n5390), .IN2(n5603), .QN(n9686) );
  NAND2X0 U16449 ( .IN1(n9450), .IN2(g3115), .QN(n15370) );
  NAND2X0 U16450 ( .IN1(n15373), .IN2(n15374), .QN(g25650) );
  INVX0 U16451 ( .INP(n15375), .ZN(n15374) );
  NOR2X0 U16452 ( .IN1(n9356), .IN2(n8799), .QN(n15375) );
  NAND3X0 U16453 ( .IN1(n8381), .IN2(n15376), .IN3(n9337), .QN(n15373) );
  NAND2X0 U16454 ( .IN1(n5998), .IN2(n15377), .QN(n15376) );
  NAND2X0 U16455 ( .IN1(n8799), .IN2(g8215), .QN(n15377) );
  NAND2X0 U16456 ( .IN1(n15378), .IN2(n15379), .QN(g25649) );
  NAND2X0 U16457 ( .IN1(n9364), .IN2(g3338), .QN(n15379) );
  INVX0 U16458 ( .INP(n15380), .ZN(n15378) );
  NOR2X0 U16459 ( .IN1(n9358), .IN2(n5998), .QN(n15380) );
  NOR2X0 U16460 ( .IN1(n9417), .IN2(n5390), .QN(g25648) );
  NAND3X0 U16461 ( .IN1(n15381), .IN2(n15382), .IN3(n15383), .QN(g25639) );
  INVX0 U16462 ( .INP(n5045), .ZN(n15383) );
  NAND2X0 U16463 ( .IN1(n9450), .IN2(g2715), .QN(n15382) );
  NAND2X0 U16464 ( .IN1(n13186), .IN2(n9371), .QN(n15381) );
  NOR2X0 U16465 ( .IN1(g2715), .IN2(n5465), .QN(n13186) );
  NAND2X0 U16466 ( .IN1(n15384), .IN2(n15385), .QN(g25638) );
  NAND2X0 U16467 ( .IN1(n9450), .IN2(g1564), .QN(n15385) );
  NAND2X0 U16468 ( .IN1(n15386), .IN2(n9371), .QN(n15384) );
  NAND2X0 U16469 ( .IN1(n15387), .IN2(n15388), .QN(n15386) );
  NAND2X0 U16470 ( .IN1(n15389), .IN2(g1559), .QN(n15388) );
  NAND3X0 U16471 ( .IN1(n15390), .IN2(n5768), .IN3(n5441), .QN(n15387) );
  NAND2X0 U16472 ( .IN1(n15391), .IN2(n15392), .QN(g25637) );
  NAND3X0 U16473 ( .IN1(n9347), .IN2(g1554), .IN3(n15389), .QN(n15392) );
  INVX0 U16474 ( .INP(n15390), .ZN(n15389) );
  NAND2X0 U16475 ( .IN1(n15393), .IN2(g1559), .QN(n15391) );
  NAND2X0 U16476 ( .IN1(n15394), .IN2(n9371), .QN(n15393) );
  NAND2X0 U16477 ( .IN1(n15390), .IN2(n5768), .QN(n15394) );
  NAND2X0 U16478 ( .IN1(n15395), .IN2(n15396), .QN(g25636) );
  NAND2X0 U16479 ( .IN1(n9450), .IN2(g1521), .QN(n15396) );
  NAND2X0 U16480 ( .IN1(n15397), .IN2(n9372), .QN(n15395) );
  NAND2X0 U16481 ( .IN1(n15398), .IN2(n15399), .QN(n15397) );
  INVX0 U16482 ( .INP(n15400), .ZN(n15399) );
  NOR2X0 U16483 ( .IN1(n15401), .IN2(n5381), .QN(n15400) );
  NAND2X0 U16484 ( .IN1(n15401), .IN2(g1306), .QN(n15398) );
  NAND3X0 U16485 ( .IN1(g7946), .IN2(g1514), .IN3(test_so49), .QN(n15401) );
  NAND2X0 U16486 ( .IN1(n15402), .IN2(n15403), .QN(g25635) );
  NAND2X0 U16487 ( .IN1(n15404), .IN2(g1484), .QN(n15403) );
  NAND2X0 U16488 ( .IN1(n15405), .IN2(n9372), .QN(n15404) );
  NAND3X0 U16489 ( .IN1(n5483), .IN2(n14037), .IN3(n14974), .QN(n15405) );
  NAND2X0 U16490 ( .IN1(n15406), .IN2(g1300), .QN(n15402) );
  NAND2X0 U16491 ( .IN1(n15407), .IN2(n15408), .QN(n15406) );
  NAND2X0 U16492 ( .IN1(n15409), .IN2(n9372), .QN(n15408) );
  NAND2X0 U16493 ( .IN1(n14974), .IN2(g1484), .QN(n15409) );
  NOR2X0 U16494 ( .IN1(n8717), .IN2(test_so12), .QN(n14974) );
  NOR3X0 U16495 ( .IN1(n15410), .IN2(test_so68), .IN3(n15411), .QN(g25634) );
  INVX0 U16496 ( .INP(n14989), .ZN(n15411) );
  NAND3X0 U16497 ( .IN1(g12923), .IN2(g1395), .IN3(n15412), .QN(n14989) );
  NOR2X0 U16498 ( .IN1(n15413), .IN2(n15414), .QN(n15410) );
  NOR2X0 U16499 ( .IN1(n8778), .IN2(n9392), .QN(n15414) );
  NOR2X0 U16500 ( .IN1(n15415), .IN2(n15416), .QN(n15413) );
  NAND2X0 U16501 ( .IN1(n15417), .IN2(n15418), .QN(g25633) );
  NAND2X0 U16502 ( .IN1(n9450), .IN2(g1379), .QN(n15418) );
  NAND2X0 U16503 ( .IN1(n15419), .IN2(n9372), .QN(n15417) );
  NAND2X0 U16504 ( .IN1(n15420), .IN2(n15421), .QN(n15419) );
  NAND2X0 U16505 ( .IN1(n15422), .IN2(g1384), .QN(n15421) );
  NAND3X0 U16506 ( .IN1(n14996), .IN2(g1351), .IN3(n8340), .QN(n15420) );
  NAND2X0 U16507 ( .IN1(n15423), .IN2(n15424), .QN(g25632) );
  NAND2X0 U16508 ( .IN1(n15425), .IN2(g1312), .QN(n15424) );
  NAND2X0 U16509 ( .IN1(n15422), .IN2(n9372), .QN(n15425) );
  INVX0 U16510 ( .INP(n14996), .ZN(n15422) );
  NAND4X0 U16511 ( .IN1(n15426), .IN2(n15427), .IN3(n9355), .IN4(g1351), .QN(
        n15423) );
  NAND2X0 U16512 ( .IN1(n14705), .IN2(n13501), .QN(n15427) );
  NAND2X0 U16513 ( .IN1(n14996), .IN2(g1389), .QN(n15426) );
  NOR2X0 U16514 ( .IN1(n9416), .IN2(n15428), .QN(g25631) );
  NOR2X0 U16515 ( .IN1(n15429), .IN2(n15430), .QN(n15428) );
  NOR2X0 U16516 ( .IN1(n5466), .IN2(n14996), .QN(n15430) );
  INVX0 U16517 ( .INP(n15431), .ZN(n15429) );
  NAND3X0 U16518 ( .IN1(n13501), .IN2(n15432), .IN3(n15433), .QN(n15431) );
  NAND2X0 U16519 ( .IN1(g1351), .IN2(n15434), .QN(n15433) );
  NAND2X0 U16520 ( .IN1(n14701), .IN2(n14705), .QN(n15434) );
  NOR2X0 U16521 ( .IN1(n8454), .IN2(n8455), .QN(n14705) );
  NAND2X0 U16522 ( .IN1(n14704), .IN2(g1389), .QN(n14701) );
  INVX0 U16523 ( .INP(n14706), .ZN(n14704) );
  NAND2X0 U16524 ( .IN1(n4896), .IN2(n5322), .QN(n15432) );
  NAND4X0 U16525 ( .IN1(n14706), .IN2(g1367), .IN3(g1345), .IN4(g1379), .QN(
        n4896) );
  INVX0 U16526 ( .INP(n14707), .ZN(n13501) );
  NAND2X0 U16527 ( .IN1(n15435), .IN2(n15436), .QN(g25630) );
  NAND2X0 U16528 ( .IN1(n15437), .IN2(g1249), .QN(n15436) );
  NAND2X0 U16529 ( .IN1(n15438), .IN2(n9372), .QN(n15437) );
  NAND2X0 U16530 ( .IN1(n8781), .IN2(g12923), .QN(n15438) );
  NAND2X0 U16531 ( .IN1(g24247), .IN2(g1266), .QN(n15435) );
  NAND2X0 U16532 ( .IN1(n15439), .IN2(n15440), .QN(g25629) );
  NAND2X0 U16533 ( .IN1(n9450), .IN2(g1221), .QN(n15440) );
  NAND2X0 U16534 ( .IN1(n15441), .IN2(n9372), .QN(n15439) );
  NAND2X0 U16535 ( .IN1(n15442), .IN2(n15443), .QN(n15441) );
  NAND2X0 U16536 ( .IN1(n15444), .IN2(g1216), .QN(n15443) );
  NAND3X0 U16537 ( .IN1(n15445), .IN2(n8880), .IN3(n5442), .QN(n15442) );
  NAND2X0 U16538 ( .IN1(n15446), .IN2(n15447), .QN(g25628) );
  NAND3X0 U16539 ( .IN1(n15444), .IN2(n9316), .IN3(test_so76), .QN(n15447) );
  NAND2X0 U16540 ( .IN1(n15448), .IN2(g1216), .QN(n15446) );
  NAND2X0 U16541 ( .IN1(n15449), .IN2(n9372), .QN(n15448) );
  NAND2X0 U16542 ( .IN1(n15445), .IN2(n8880), .QN(n15449) );
  NAND2X0 U16543 ( .IN1(n15450), .IN2(n15451), .QN(g25627) );
  NAND2X0 U16544 ( .IN1(n9450), .IN2(g1178), .QN(n15451) );
  NAND2X0 U16545 ( .IN1(n15452), .IN2(n9372), .QN(n15450) );
  NAND2X0 U16546 ( .IN1(n15453), .IN2(n15454), .QN(n15452) );
  NAND2X0 U16547 ( .IN1(n11762), .IN2(n13534), .QN(n15454) );
  NAND2X0 U16548 ( .IN1(n15455), .IN2(g962), .QN(n15453) );
  NAND2X0 U16549 ( .IN1(n11762), .IN2(g7916), .QN(n15455) );
  NOR2X0 U16550 ( .IN1(n5599), .IN2(n5363), .QN(n11762) );
  NAND2X0 U16551 ( .IN1(n15456), .IN2(n15457), .QN(g25626) );
  NAND2X0 U16552 ( .IN1(n15458), .IN2(g1141), .QN(n15457) );
  NAND2X0 U16553 ( .IN1(n15459), .IN2(n9372), .QN(n15458) );
  NAND3X0 U16554 ( .IN1(n5341), .IN2(n14079), .IN3(n15011), .QN(n15459) );
  NAND2X0 U16555 ( .IN1(n15460), .IN2(g956), .QN(n15456) );
  NAND2X0 U16556 ( .IN1(n15461), .IN2(n15462), .QN(n15460) );
  NAND2X0 U16557 ( .IN1(n15463), .IN2(n9372), .QN(n15462) );
  NAND2X0 U16558 ( .IN1(n15011), .IN2(g1141), .QN(n15463) );
  NOR2X0 U16559 ( .IN1(g1152), .IN2(n8865), .QN(n15011) );
  NOR3X0 U16560 ( .IN1(g979), .IN2(n15464), .IN3(n15465), .QN(g25625) );
  NOR2X0 U16561 ( .IN1(n15466), .IN2(n15467), .QN(n15465) );
  NOR2X0 U16562 ( .IN1(n8779), .IN2(n9388), .QN(n15467) );
  NOR2X0 U16563 ( .IN1(n15468), .IN2(n15469), .QN(n15466) );
  INVX0 U16564 ( .INP(n15027), .ZN(n15464) );
  NAND3X0 U16565 ( .IN1(g12919), .IN2(g1052), .IN3(n15470), .QN(n15027) );
  NAND3X0 U16566 ( .IN1(n15471), .IN2(n15472), .IN3(n15473), .QN(g25624) );
  NAND3X0 U16567 ( .IN1(n15033), .IN2(n8339), .IN3(n15032), .QN(n15473) );
  NAND3X0 U16568 ( .IN1(n15474), .IN2(g1041), .IN3(n9337), .QN(n15472) );
  NAND2X0 U16569 ( .IN1(n9449), .IN2(g1036), .QN(n15471) );
  NAND2X0 U16570 ( .IN1(n15475), .IN2(n15476), .QN(g25623) );
  NAND2X0 U16571 ( .IN1(test_so20), .IN2(n15477), .QN(n15476) );
  NAND2X0 U16572 ( .IN1(n15474), .IN2(n9372), .QN(n15477) );
  INVX0 U16573 ( .INP(n15033), .ZN(n15474) );
  NAND2X0 U16574 ( .IN1(n15032), .IN2(n15478), .QN(n15475) );
  NAND2X0 U16575 ( .IN1(n13538), .IN2(n15479), .QN(n15478) );
  NAND2X0 U16576 ( .IN1(n15480), .IN2(n15481), .QN(n15479) );
  INVX0 U16577 ( .INP(n14716), .ZN(n15481) );
  NAND2X0 U16578 ( .IN1(g1030), .IN2(g1018), .QN(n15480) );
  INVX0 U16579 ( .INP(n14722), .ZN(n13538) );
  NOR2X0 U16580 ( .IN1(n9415), .IN2(n5321), .QN(n15032) );
  NOR2X0 U16581 ( .IN1(n9415), .IN2(n15482), .QN(g25622) );
  NOR2X0 U16582 ( .IN1(n15483), .IN2(n15484), .QN(n15482) );
  NOR2X0 U16583 ( .IN1(n15033), .IN2(n8890), .QN(n15484) );
  NOR2X0 U16584 ( .IN1(n14722), .IN2(n15485), .QN(n15483) );
  NOR2X0 U16585 ( .IN1(n15486), .IN2(n15487), .QN(n15485) );
  NOR2X0 U16586 ( .IN1(n4921), .IN2(g1008), .QN(n15487) );
  NAND4X0 U16587 ( .IN1(n14721), .IN2(g1024), .IN3(g1002), .IN4(g1036), .QN(
        n4921) );
  NOR2X0 U16588 ( .IN1(n14716), .IN2(n14720), .QN(n15486) );
  NAND3X0 U16589 ( .IN1(g1018), .IN2(g1030), .IN3(g1008), .QN(n14720) );
  NOR2X0 U16590 ( .IN1(n14721), .IN2(n8835), .QN(n14716) );
  NAND2X0 U16591 ( .IN1(n15488), .IN2(n15489), .QN(g25621) );
  NAND2X0 U16592 ( .IN1(n15490), .IN2(g904), .QN(n15489) );
  NAND2X0 U16593 ( .IN1(n15491), .IN2(n9372), .QN(n15490) );
  NAND2X0 U16594 ( .IN1(n8782), .IN2(g12919), .QN(n15491) );
  NAND2X0 U16595 ( .IN1(g24231), .IN2(g921), .QN(n15488) );
  NOR2X0 U16596 ( .IN1(n5562), .IN2(n15492), .QN(g25619) );
  NOR2X0 U16597 ( .IN1(n9415), .IN2(n15493), .QN(n15492) );
  NOR2X0 U16598 ( .IN1(n15079), .IN2(n15494), .QN(n15493) );
  NOR2X0 U16599 ( .IN1(n15495), .IN2(g843), .QN(n15494) );
  INVX0 U16600 ( .INP(n15496), .ZN(n15079) );
  NAND2X0 U16601 ( .IN1(n15495), .IN2(g843), .QN(n15496) );
  NAND2X0 U16602 ( .IN1(n15497), .IN2(n15498), .QN(g25618) );
  NAND2X0 U16603 ( .IN1(n15499), .IN2(g817), .QN(n15498) );
  NAND2X0 U16604 ( .IN1(n15500), .IN2(n9372), .QN(n15499) );
  NAND3X0 U16605 ( .IN1(n4948), .IN2(n14104), .IN3(n8796), .QN(n15500) );
  NAND2X0 U16606 ( .IN1(n15501), .IN2(g832), .QN(n15497) );
  NAND2X0 U16607 ( .IN1(n15502), .IN2(n15503), .QN(n15501) );
  NAND2X0 U16608 ( .IN1(n14147), .IN2(n14104), .QN(n15503) );
  NAND2X0 U16609 ( .IN1(n5822), .IN2(n4518), .QN(n15502) );
  NOR2X0 U16610 ( .IN1(n15504), .IN2(n9390), .QN(n4518) );
  INVX0 U16611 ( .INP(n14104), .ZN(n15504) );
  NAND2X0 U16612 ( .IN1(n15505), .IN2(n15506), .QN(g25617) );
  NAND3X0 U16613 ( .IN1(n15507), .IN2(n15508), .IN3(n14104), .QN(n15506) );
  NAND2X0 U16614 ( .IN1(g847), .IN2(n15509), .QN(n14104) );
  NAND2X0 U16615 ( .IN1(n5733), .IN2(g837), .QN(n15509) );
  NAND2X0 U16616 ( .IN1(n15510), .IN2(g817), .QN(n15508) );
  NAND2X0 U16617 ( .IN1(n5822), .IN2(n15511), .QN(n15507) );
  NAND2X0 U16618 ( .IN1(n9449), .IN2(g812), .QN(n15505) );
  NOR2X0 U16619 ( .IN1(n9416), .IN2(n15512), .QN(g25616) );
  NOR3X0 U16620 ( .IN1(n15513), .IN2(n15514), .IN3(n15515), .QN(n15512) );
  NOR2X0 U16621 ( .IN1(g732), .IN2(n15516), .QN(n15515) );
  INVX0 U16622 ( .INP(n15517), .ZN(n15514) );
  NAND3X0 U16623 ( .IN1(g732), .IN2(n15089), .IN3(n15516), .QN(n15517) );
  NOR2X0 U16624 ( .IN1(n15516), .IN2(n15089), .QN(n15513) );
  NAND4X0 U16625 ( .IN1(n5327), .IN2(n14765), .IN3(n14769), .IN4(n15518), .QN(
        n15089) );
  NOR3X0 U16626 ( .IN1(g370), .IN2(g490), .IN3(g482), .QN(n15518) );
  NOR2X0 U16627 ( .IN1(g518), .IN2(test_so54), .QN(n14769) );
  NOR2X0 U16628 ( .IN1(n15519), .IN2(n15520), .QN(n15516) );
  INVX0 U16629 ( .INP(n15521), .ZN(n15520) );
  NAND2X0 U16630 ( .IN1(n15522), .IN2(n15523), .QN(n15521) );
  NOR2X0 U16631 ( .IN1(n15523), .IN2(n15522), .QN(n15519) );
  NAND2X0 U16632 ( .IN1(n15524), .IN2(n15525), .QN(n15522) );
  INVX0 U16633 ( .INP(n15526), .ZN(n15525) );
  NOR2X0 U16634 ( .IN1(n15527), .IN2(g262), .QN(n15526) );
  NAND2X0 U16635 ( .IN1(n15527), .IN2(g262), .QN(n15524) );
  NAND2X0 U16636 ( .IN1(n15528), .IN2(n15529), .QN(n15527) );
  NAND2X0 U16637 ( .IN1(n8589), .IN2(g269), .QN(n15529) );
  NAND2X0 U16638 ( .IN1(n8472), .IN2(g232), .QN(n15528) );
  NOR2X0 U16639 ( .IN1(n15530), .IN2(n15531), .QN(n15523) );
  INVX0 U16640 ( .INP(n15532), .ZN(n15531) );
  NAND2X0 U16641 ( .IN1(n8470), .IN2(n15533), .QN(n15532) );
  NOR2X0 U16642 ( .IN1(n15533), .IN2(n8470), .QN(n15530) );
  NAND3X0 U16643 ( .IN1(n15534), .IN2(n15535), .IN3(n14794), .QN(n15533) );
  NAND3X0 U16644 ( .IN1(n6008), .IN2(n5597), .IN3(n8590), .QN(n14794) );
  NAND2X0 U16645 ( .IN1(n15536), .IN2(g239), .QN(n15535) );
  NAND2X0 U16646 ( .IN1(n15537), .IN2(n15538), .QN(n15536) );
  NAND2X0 U16647 ( .IN1(n6008), .IN2(g225), .QN(n15538) );
  NAND2X0 U16648 ( .IN1(n5597), .IN2(g246), .QN(n15537) );
  NAND3X0 U16649 ( .IN1(g225), .IN2(g246), .IN3(n8590), .QN(n15534) );
  NAND2X0 U16650 ( .IN1(n15539), .IN2(n15540), .QN(g25615) );
  NAND2X0 U16651 ( .IN1(n15541), .IN2(g667), .QN(n15540) );
  NAND2X0 U16652 ( .IN1(n14752), .IN2(g686), .QN(n15539) );
  NAND3X0 U16653 ( .IN1(n15542), .IN2(n15543), .IN3(n15544), .QN(g25614) );
  NAND2X0 U16654 ( .IN1(n9449), .IN2(g691), .QN(n15544) );
  NAND2X0 U16655 ( .IN1(n15541), .IN2(g686), .QN(n15543) );
  NAND2X0 U16656 ( .IN1(n5111), .IN2(n15545), .QN(n15542) );
  NAND2X0 U16657 ( .IN1(n15546), .IN2(n15547), .QN(g25613) );
  NAND2X0 U16658 ( .IN1(g559), .IN2(n9413), .QN(n15547) );
  NAND4X0 U16659 ( .IN1(n2421), .IN2(n15548), .IN3(n15549), .IN4(n15550), .QN(
        n15546) );
  NAND2X0 U16660 ( .IN1(n8842), .IN2(n15551), .QN(n15550) );
  NAND2X0 U16661 ( .IN1(n15100), .IN2(g562), .QN(n15549) );
  INVX0 U16662 ( .INP(n15551), .ZN(n15100) );
  NAND2X0 U16663 ( .IN1(g29211), .IN2(n15552), .QN(n15551) );
  NAND2X0 U16664 ( .IN1(n8330), .IN2(g12368), .QN(n15552) );
  NAND2X0 U16665 ( .IN1(g626), .IN2(n9340), .QN(n15548) );
  NAND2X0 U16666 ( .IN1(n15553), .IN2(n15554), .QN(g25612) );
  NAND2X0 U16667 ( .IN1(n15555), .IN2(g513), .QN(n15554) );
  NAND2X0 U16668 ( .IN1(n15541), .IN2(g518), .QN(n15553) );
  NAND2X0 U16669 ( .IN1(n15556), .IN2(n15557), .QN(g25611) );
  NAND2X0 U16670 ( .IN1(n15555), .IN2(g504), .QN(n15557) );
  NAND2X0 U16671 ( .IN1(n15558), .IN2(n9372), .QN(n15555) );
  NAND2X0 U16672 ( .IN1(n15545), .IN2(n14141), .QN(n15558) );
  INVX0 U16673 ( .INP(n4962), .ZN(n14141) );
  NAND2X0 U16674 ( .IN1(n15541), .IN2(g513), .QN(n15556) );
  NAND3X0 U16675 ( .IN1(n15559), .IN2(n15560), .IN3(n15561), .QN(g25610) );
  NAND2X0 U16676 ( .IN1(n15541), .IN2(g504), .QN(n15560) );
  NAND2X0 U16677 ( .IN1(test_so54), .IN2(n14752), .QN(n15559) );
  NAND3X0 U16678 ( .IN1(n15562), .IN2(n15561), .IN3(n15563), .QN(g25609) );
  NAND2X0 U16679 ( .IN1(n14754), .IN2(n5287), .QN(n15563) );
  NAND2X0 U16680 ( .IN1(n4962), .IN2(n14754), .QN(n15561) );
  NOR2X0 U16681 ( .IN1(n15106), .IN2(n9389), .QN(n14754) );
  NAND2X0 U16682 ( .IN1(test_so54), .IN2(n15564), .QN(n15562) );
  NAND2X0 U16683 ( .IN1(n14752), .IN2(n15565), .QN(n15564) );
  NAND2X0 U16684 ( .IN1(n5548), .IN2(n9372), .QN(n15565) );
  INVX0 U16685 ( .INP(n15541), .ZN(n14752) );
  NOR2X0 U16686 ( .IN1(n15545), .IN2(n9391), .QN(n15541) );
  INVX0 U16687 ( .INP(n15106), .ZN(n15545) );
  NAND3X0 U16688 ( .IN1(g385), .IN2(g358), .IN3(n5633), .QN(n15106) );
  NAND3X0 U16689 ( .IN1(n15566), .IN2(n15567), .IN3(n15568), .QN(g25605) );
  NAND2X0 U16690 ( .IN1(n9449), .IN2(g168), .QN(n15568) );
  NAND3X0 U16691 ( .IN1(n14765), .IN2(g246), .IN3(n15569), .QN(n15567) );
  NAND2X0 U16692 ( .IN1(n15570), .IN2(g460), .QN(n15566) );
  NAND2X0 U16693 ( .IN1(n15571), .IN2(n15572), .QN(g25604) );
  NAND2X0 U16694 ( .IN1(g452), .IN2(n15570), .QN(n15572) );
  NAND2X0 U16695 ( .IN1(n15573), .IN2(g460), .QN(n15571) );
  NAND3X0 U16696 ( .IN1(n15574), .IN2(n15575), .IN3(n15576), .QN(g25602) );
  NAND2X0 U16697 ( .IN1(n9449), .IN2(g405), .QN(n15576) );
  NAND3X0 U16698 ( .IN1(n14765), .IN2(g446), .IN3(n15569), .QN(n15575) );
  NAND2X0 U16699 ( .IN1(n15570), .IN2(test_so72), .QN(n15574) );
  NAND2X0 U16700 ( .IN1(n15577), .IN2(n15578), .QN(g25601) );
  NAND2X0 U16701 ( .IN1(n15570), .IN2(g174), .QN(n15578) );
  NAND2X0 U16702 ( .IN1(test_so72), .IN2(n15573), .QN(n15577) );
  NAND2X0 U16703 ( .IN1(n15579), .IN2(n15580), .QN(g25600) );
  NAND2X0 U16704 ( .IN1(n15570), .IN2(g168), .QN(n15580) );
  INVX0 U16705 ( .INP(n15573), .ZN(n15570) );
  NAND2X0 U16706 ( .IN1(n15573), .IN2(g174), .QN(n15579) );
  NAND2X0 U16707 ( .IN1(n15581), .IN2(n9372), .QN(n15573) );
  NAND2X0 U16708 ( .IN1(n8816), .IN2(n14765), .QN(n15581) );
  INVX0 U16709 ( .INP(n1205), .ZN(n14765) );
  NAND2X0 U16710 ( .IN1(n10558), .IN2(n15582), .QN(g25599) );
  NAND2X0 U16711 ( .IN1(n9449), .IN2(g385), .QN(n15582) );
  NAND2X0 U16712 ( .IN1(n15583), .IN2(n15584), .QN(g25598) );
  NAND3X0 U16713 ( .IN1(n9347), .IN2(g385), .IN3(n1205), .QN(n15584) );
  NAND2X0 U16714 ( .IN1(n15585), .IN2(g376), .QN(n15583) );
  NAND2X0 U16715 ( .IN1(n15586), .IN2(n9366), .QN(n15585) );
  NAND2X0 U16716 ( .IN1(n1205), .IN2(g358), .QN(n15586) );
  NAND3X0 U16717 ( .IN1(g376), .IN2(g358), .IN3(g385), .QN(n1205) );
  NAND3X0 U16718 ( .IN1(n15587), .IN2(n15588), .IN3(n15589), .QN(g25597) );
  NAND2X0 U16719 ( .IN1(n15590), .IN2(n15569), .QN(n15589) );
  NOR2X0 U16720 ( .IN1(g370), .IN2(n9390), .QN(n15569) );
  INVX0 U16721 ( .INP(n10558), .ZN(n15590) );
  NAND3X0 U16722 ( .IN1(n10558), .IN2(g370), .IN3(n9337), .QN(n15588) );
  NAND3X0 U16723 ( .IN1(g376), .IN2(g8719), .IN3(g385), .QN(n10558) );
  NAND2X0 U16724 ( .IN1(n9449), .IN2(g358), .QN(n15587) );
  NAND2X0 U16725 ( .IN1(n15591), .IN2(n15592), .QN(g25596) );
  NAND2X0 U16726 ( .IN1(n9448), .IN2(g370), .QN(n15592) );
  NAND2X0 U16727 ( .IN1(n15593), .IN2(n9372), .QN(n15591) );
  NAND2X0 U16728 ( .IN1(n15594), .IN2(n15595), .QN(n15593) );
  NAND2X0 U16729 ( .IN1(n8473), .IN2(g376), .QN(n15595) );
  NAND2X0 U16730 ( .IN1(n5633), .IN2(g358), .QN(n15594) );
  NOR3X0 U16731 ( .IN1(g8719), .IN2(n9384), .IN3(g358), .QN(g25595) );
  NAND2X0 U16732 ( .IN1(n15596), .IN2(n15597), .QN(g25593) );
  NAND2X0 U16733 ( .IN1(n9448), .IN2(g191), .QN(n15597) );
  NAND2X0 U16734 ( .IN1(n15598), .IN2(n9372), .QN(n15596) );
  NAND2X0 U16735 ( .IN1(n15599), .IN2(n15600), .QN(n15598) );
  NAND2X0 U16736 ( .IN1(n15601), .IN2(g209), .QN(n15600) );
  NAND2X0 U16737 ( .IN1(n15602), .IN2(n15603), .QN(n15599) );
  NAND2X0 U16738 ( .IN1(n15604), .IN2(n15605), .QN(g25592) );
  INVX0 U16739 ( .INP(n15606), .ZN(n15605) );
  NOR2X0 U16740 ( .IN1(n9359), .IN2(n8747), .QN(n15606) );
  NAND3X0 U16741 ( .IN1(n15607), .IN2(n15608), .IN3(n9338), .QN(n15604) );
  INVX0 U16742 ( .INP(n15609), .ZN(n15608) );
  NOR2X0 U16743 ( .IN1(g8358), .IN2(n15610), .QN(n15609) );
  NAND2X0 U16744 ( .IN1(n15610), .IN2(g8358), .QN(n15607) );
  NOR2X0 U16745 ( .IN1(n15602), .IN2(n15601), .QN(n15610) );
  INVX0 U16746 ( .INP(n15603), .ZN(n15601) );
  NOR2X0 U16747 ( .IN1(n8903), .IN2(n8718), .QN(n15603) );
  NAND2X0 U16748 ( .IN1(n15611), .IN2(n15612), .QN(n15602) );
  NAND2X0 U16749 ( .IN1(n8453), .IN2(g8358), .QN(n15612) );
  NAND2X0 U16750 ( .IN1(n8452), .IN2(g191), .QN(n15611) );
  NAND2X0 U16751 ( .IN1(n15613), .IN2(n15614), .QN(g25591) );
  NAND2X0 U16752 ( .IN1(n8718), .IN2(n9371), .QN(n15614) );
  NAND2X0 U16753 ( .IN1(n9448), .IN2(g209), .QN(n15613) );
  INVX0 U16754 ( .INP(n10613), .ZN(g25259) );
  NAND2X0 U16755 ( .IN1(n5549), .IN2(g1668), .QN(n10613) );
  NOR2X0 U16756 ( .IN1(g1657), .IN2(n8870), .QN(g25167) );
  NOR2X0 U16757 ( .IN1(n8710), .IN2(n15615), .QN(g24355) );
  NOR2X0 U16758 ( .IN1(n9413), .IN2(n15616), .QN(n15615) );
  NAND2X0 U16759 ( .IN1(n15617), .IN2(n15618), .QN(g24354) );
  NAND2X0 U16760 ( .IN1(n9448), .IN2(g6727), .QN(n15618) );
  NAND3X0 U16761 ( .IN1(n8709), .IN2(n15616), .IN3(n9338), .QN(n15617) );
  NAND2X0 U16762 ( .IN1(n15619), .IN2(n15620), .QN(g24353) );
  NAND2X0 U16763 ( .IN1(n9448), .IN2(g6723), .QN(n15620) );
  NAND3X0 U16764 ( .IN1(n15621), .IN2(n15616), .IN3(n9338), .QN(n15619) );
  INVX0 U16765 ( .INP(n15622), .ZN(n15616) );
  NOR2X0 U16766 ( .IN1(n15623), .IN2(n5531), .QN(n15622) );
  NAND2X0 U16767 ( .IN1(n5531), .IN2(n15623), .QN(n15621) );
  NAND4X0 U16768 ( .IN1(test_so80), .IN2(g14828), .IN3(g17688), .IN4(g17778), 
        .QN(n15623) );
  NOR4X0 U16769 ( .IN1(n15624), .IN2(g13099), .IN3(n15625), .IN4(n15626), .QN(
        g24352) );
  NOR2X0 U16770 ( .IN1(test_so80), .IN2(n5700), .QN(n15626) );
  NOR2X0 U16771 ( .IN1(n8571), .IN2(g14828), .QN(n15625) );
  NAND3X0 U16772 ( .IN1(n8557), .IN2(n9316), .IN3(n8669), .QN(n15624) );
  NOR2X0 U16773 ( .IN1(n8580), .IN2(n15627), .QN(g24351) );
  NOR2X0 U16774 ( .IN1(n9412), .IN2(n15628), .QN(n15627) );
  NAND2X0 U16775 ( .IN1(n15629), .IN2(n15630), .QN(g24350) );
  NAND2X0 U16776 ( .IN1(test_so69), .IN2(n9512), .QN(n15630) );
  NAND3X0 U16777 ( .IN1(n8579), .IN2(n15628), .IN3(n9338), .QN(n15629) );
  NAND2X0 U16778 ( .IN1(n15631), .IN2(test_so69), .QN(n15628) );
  NAND2X0 U16779 ( .IN1(n15632), .IN2(n15633), .QN(g24349) );
  NAND2X0 U16780 ( .IN1(n9448), .IN2(g6377), .QN(n15633) );
  NAND2X0 U16781 ( .IN1(n15634), .IN2(n9371), .QN(n15632) );
  NAND2X0 U16782 ( .IN1(n15635), .IN2(n15636), .QN(n15634) );
  NAND2X0 U16783 ( .IN1(test_so69), .IN2(n15637), .QN(n15636) );
  NAND2X0 U16784 ( .IN1(n15631), .IN2(n8889), .QN(n15635) );
  INVX0 U16785 ( .INP(n15637), .ZN(n15631) );
  NAND4X0 U16786 ( .IN1(g12422), .IN2(g14779), .IN3(g17649), .IN4(g17760), 
        .QN(n15637) );
  NOR4X0 U16787 ( .IN1(n15638), .IN2(g13085), .IN3(n15639), .IN4(n15640), .QN(
        g24348) );
  NOR2X0 U16788 ( .IN1(n5703), .IN2(g12422), .QN(n15640) );
  NOR2X0 U16789 ( .IN1(n8575), .IN2(g14779), .QN(n15639) );
  NAND3X0 U16790 ( .IN1(n8560), .IN2(n9316), .IN3(n8678), .QN(n15638) );
  NOR2X0 U16791 ( .IN1(n8581), .IN2(n15641), .QN(g24347) );
  NOR2X0 U16792 ( .IN1(n9412), .IN2(n15642), .QN(n15641) );
  NAND2X0 U16793 ( .IN1(n15643), .IN2(n15644), .QN(g24346) );
  NAND2X0 U16794 ( .IN1(n9448), .IN2(g6035), .QN(n15644) );
  NAND3X0 U16795 ( .IN1(n15642), .IN2(n8887), .IN3(n9338), .QN(n15643) );
  NAND2X0 U16796 ( .IN1(n15645), .IN2(n15646), .QN(g24345) );
  NAND2X0 U16797 ( .IN1(n9447), .IN2(g6031), .QN(n15646) );
  NAND3X0 U16798 ( .IN1(n15647), .IN2(n15642), .IN3(n9338), .QN(n15645) );
  INVX0 U16799 ( .INP(n15648), .ZN(n15642) );
  NOR2X0 U16800 ( .IN1(n15649), .IN2(n5528), .QN(n15648) );
  NAND2X0 U16801 ( .IN1(n5528), .IN2(n15649), .QN(n15647) );
  NAND4X0 U16802 ( .IN1(g12350), .IN2(g14738), .IN3(g17607), .IN4(g17739), 
        .QN(n15649) );
  NOR4X0 U16803 ( .IN1(n15650), .IN2(g13068), .IN3(n15651), .IN4(n15652), .QN(
        g24344) );
  NOR2X0 U16804 ( .IN1(n5698), .IN2(g12350), .QN(n15652) );
  NOR2X0 U16805 ( .IN1(n8566), .IN2(g14738), .QN(n15651) );
  NAND3X0 U16806 ( .IN1(n8551), .IN2(n9316), .IN3(n8655), .QN(n15650) );
  NOR2X0 U16807 ( .IN1(n8585), .IN2(n15653), .QN(g24343) );
  NOR2X0 U16808 ( .IN1(n9412), .IN2(n15654), .QN(n15653) );
  NAND2X0 U16809 ( .IN1(n15655), .IN2(n15656), .QN(g24342) );
  NAND2X0 U16810 ( .IN1(n9447), .IN2(g5689), .QN(n15656) );
  NAND3X0 U16811 ( .IN1(n8584), .IN2(n15654), .IN3(n9338), .QN(n15655) );
  NAND2X0 U16812 ( .IN1(n15657), .IN2(n15658), .QN(g24341) );
  NAND2X0 U16813 ( .IN1(n9447), .IN2(g5685), .QN(n15658) );
  NAND3X0 U16814 ( .IN1(n15659), .IN2(n15654), .IN3(n9338), .QN(n15657) );
  INVX0 U16815 ( .INP(n15660), .ZN(n15654) );
  NOR2X0 U16816 ( .IN1(n15661), .IN2(n5529), .QN(n15660) );
  NAND2X0 U16817 ( .IN1(n5529), .IN2(n15661), .QN(n15659) );
  NAND4X0 U16818 ( .IN1(g12300), .IN2(g14694), .IN3(g17580), .IN4(g17711), 
        .QN(n15661) );
  NOR4X0 U16819 ( .IN1(n15662), .IN2(g13049), .IN3(n15663), .IN4(n15664), .QN(
        g24340) );
  NOR2X0 U16820 ( .IN1(n5705), .IN2(g12300), .QN(n15664) );
  NOR2X0 U16821 ( .IN1(n8568), .IN2(g14694), .QN(n15663) );
  NAND3X0 U16822 ( .IN1(n8553), .IN2(n9315), .IN3(n8660), .QN(n15662) );
  NOR2X0 U16823 ( .IN1(n8712), .IN2(n15665), .QN(g24339) );
  NOR2X0 U16824 ( .IN1(n9411), .IN2(n15666), .QN(n15665) );
  NAND2X0 U16825 ( .IN1(n15667), .IN2(n15668), .QN(g24338) );
  NAND2X0 U16826 ( .IN1(test_so10), .IN2(n9512), .QN(n15668) );
  NAND3X0 U16827 ( .IN1(n8711), .IN2(n15666), .IN3(n9338), .QN(n15667) );
  NAND2X0 U16828 ( .IN1(n15669), .IN2(test_so10), .QN(n15666) );
  NAND2X0 U16829 ( .IN1(n15670), .IN2(n15671), .QN(g24337) );
  NAND2X0 U16830 ( .IN1(n9447), .IN2(g5339), .QN(n15671) );
  NAND2X0 U16831 ( .IN1(n15672), .IN2(n9370), .QN(n15670) );
  NAND2X0 U16832 ( .IN1(n15673), .IN2(n15674), .QN(n15672) );
  NAND2X0 U16833 ( .IN1(test_so10), .IN2(n15675), .QN(n15674) );
  NAND2X0 U16834 ( .IN1(n15669), .IN2(n8888), .QN(n15673) );
  INVX0 U16835 ( .INP(n15675), .ZN(n15669) );
  NAND4X0 U16836 ( .IN1(g12238), .IN2(g14662), .IN3(g17519), .IN4(g17674), 
        .QN(n15675) );
  NOR4X0 U16837 ( .IN1(n15676), .IN2(g17577), .IN3(n15677), .IN4(n15678), .QN(
        g24336) );
  NOR2X0 U16838 ( .IN1(n5704), .IN2(g12238), .QN(n15678) );
  NOR2X0 U16839 ( .IN1(n8564), .IN2(g14662), .QN(n15677) );
  NAND3X0 U16840 ( .IN1(n8549), .IN2(n9315), .IN3(n8629), .QN(n15676) );
  NAND2X0 U16841 ( .IN1(n15679), .IN2(n15680), .QN(g24335) );
  NAND3X0 U16842 ( .IN1(n5653), .IN2(g4643), .IN3(n15681), .QN(n15680) );
  INVX0 U16843 ( .INP(n15682), .ZN(n15681) );
  INVX0 U16844 ( .INP(n15683), .ZN(n15679) );
  NOR2X0 U16845 ( .IN1(n9358), .IN2(n5541), .QN(n15683) );
  NAND2X0 U16846 ( .IN1(n15684), .IN2(n15685), .QN(g24334) );
  NAND4X0 U16847 ( .IN1(n5303), .IN2(n5365), .IN3(n15686), .IN4(n15687), .QN(
        n15685) );
  NOR4X0 U16848 ( .IN1(g4584), .IN2(g4608), .IN3(g4616), .IN4(n15682), .QN(
        n15687) );
  NAND4X0 U16849 ( .IN1(n9362), .IN2(n8867), .IN3(n5506), .IN4(n15688), .QN(
        n15682) );
  NOR3X0 U16850 ( .IN1(g4358), .IN2(g4332), .IN3(g4311), .QN(n15688) );
  NOR3X0 U16851 ( .IN1(n10698), .IN2(n5844), .IN3(n5653), .QN(n15686) );
  INVX0 U16852 ( .INP(n10446), .ZN(n10698) );
  NOR2X0 U16853 ( .IN1(n8873), .IN2(g4639), .QN(n10446) );
  NAND2X0 U16854 ( .IN1(n9447), .IN2(g4358), .QN(n15684) );
  NOR2X0 U16855 ( .IN1(n5710), .IN2(n9354), .QN(g24298) );
  NAND2X0 U16856 ( .IN1(n15689), .IN2(n15690), .QN(g24282) );
  NAND2X0 U16857 ( .IN1(n15691), .IN2(g4308), .QN(n15690) );
  NAND2X0 U16858 ( .IN1(n9366), .IN2(g9251), .QN(n15691) );
  NAND2X0 U16859 ( .IN1(g24281), .IN2(g9251), .QN(n15689) );
  NOR2X0 U16860 ( .IN1(g4308), .IN2(n9393), .QN(g24281) );
  NAND2X0 U16861 ( .IN1(n15692), .IN2(n15693), .QN(g24280) );
  NAND2X0 U16862 ( .IN1(n15694), .IN2(g4269), .QN(n15693) );
  NAND2X0 U16863 ( .IN1(n15695), .IN2(n9370), .QN(n15694) );
  NAND3X0 U16864 ( .IN1(g4264), .IN2(g4258), .IN3(n5764), .QN(n15695) );
  NAND2X0 U16865 ( .IN1(n15696), .IN2(g4273), .QN(n15692) );
  NAND2X0 U16866 ( .IN1(n15697), .IN2(n15698), .QN(n15696) );
  NAND2X0 U16867 ( .IN1(n5763), .IN2(n9370), .QN(n15698) );
  NAND3X0 U16868 ( .IN1(n15699), .IN2(n15700), .IN3(n15701), .QN(g24279) );
  NAND2X0 U16869 ( .IN1(n15702), .IN2(n15703), .QN(n15701) );
  INVX0 U16870 ( .INP(n15704), .ZN(n15700) );
  NOR2X0 U16871 ( .IN1(n9359), .IN2(n8514), .QN(n15704) );
  NAND2X0 U16872 ( .IN1(n15705), .IN2(n9370), .QN(n15699) );
  NAND2X0 U16873 ( .IN1(n15706), .IN2(n15707), .QN(n15705) );
  INVX0 U16874 ( .INP(n15708), .ZN(n15707) );
  NOR3X0 U16875 ( .IN1(n15703), .IN2(n15702), .IN3(n15709), .QN(n15708) );
  NOR2X0 U16876 ( .IN1(n8514), .IN2(n5726), .QN(n15702) );
  NAND2X0 U16877 ( .IN1(n15709), .IN2(n15703), .QN(n15706) );
  INVX0 U16878 ( .INP(n15710), .ZN(n15709) );
  NAND3X0 U16879 ( .IN1(n5726), .IN2(n15711), .IN3(n8514), .QN(n15710) );
  NAND4X0 U16880 ( .IN1(n15969), .IN2(n15970), .IN3(n15968), .IN4(n15712), 
        .QN(n15711) );
  NOR4X0 U16881 ( .IN1(g8915), .IN2(g8916), .IN3(g11770), .IN4(g8920), .QN(
        n15712) );
  NOR2X0 U16882 ( .IN1(n8587), .IN2(n15713), .QN(g24278) );
  NOR2X0 U16883 ( .IN1(n9411), .IN2(n15714), .QN(n15713) );
  NAND2X0 U16884 ( .IN1(n15715), .IN2(n15716), .QN(g24277) );
  NAND2X0 U16885 ( .IN1(n9447), .IN2(g4040), .QN(n15716) );
  NAND3X0 U16886 ( .IN1(n8586), .IN2(n15714), .IN3(n9339), .QN(n15715) );
  NAND2X0 U16887 ( .IN1(n15717), .IN2(n15718), .QN(g24276) );
  NAND2X0 U16888 ( .IN1(n9447), .IN2(g4031), .QN(n15718) );
  NAND3X0 U16889 ( .IN1(n15719), .IN2(n15714), .IN3(n9339), .QN(n15717) );
  INVX0 U16890 ( .INP(n15720), .ZN(n15714) );
  NOR2X0 U16891 ( .IN1(n15721), .IN2(n5530), .QN(n15720) );
  NAND2X0 U16892 ( .IN1(n5530), .IN2(n15721), .QN(n15719) );
  NAND4X0 U16893 ( .IN1(g11418), .IN2(g13966), .IN3(g16659), .IN4(g16775), 
        .QN(n15721) );
  NOR4X0 U16894 ( .IN1(n15722), .IN2(g14518), .IN3(n15723), .IN4(n15724), .QN(
        g24275) );
  NOR2X0 U16895 ( .IN1(n5701), .IN2(g11418), .QN(n15724) );
  NOR2X0 U16896 ( .IN1(n8569), .IN2(g13966), .QN(n15723) );
  NAND3X0 U16897 ( .IN1(n8555), .IN2(n9313), .IN3(n8664), .QN(n15722) );
  NOR2X0 U16898 ( .IN1(n8583), .IN2(n15725), .QN(g24274) );
  NOR2X0 U16899 ( .IN1(n9412), .IN2(n15726), .QN(n15725) );
  NAND2X0 U16900 ( .IN1(n15727), .IN2(n15728), .QN(g24273) );
  NAND2X0 U16901 ( .IN1(n9446), .IN2(g3689), .QN(n15728) );
  NAND3X0 U16902 ( .IN1(n8582), .IN2(n15726), .IN3(n9339), .QN(n15727) );
  NAND2X0 U16903 ( .IN1(n15729), .IN2(n15730), .QN(g24272) );
  NAND2X0 U16904 ( .IN1(n9446), .IN2(g3680), .QN(n15730) );
  NAND3X0 U16905 ( .IN1(n15731), .IN2(n15726), .IN3(n9339), .QN(n15729) );
  INVX0 U16906 ( .INP(n15732), .ZN(n15726) );
  NOR2X0 U16907 ( .IN1(n15733), .IN2(n5532), .QN(n15732) );
  NAND2X0 U16908 ( .IN1(n5532), .IN2(n15733), .QN(n15731) );
  NAND4X0 U16909 ( .IN1(g11388), .IN2(g13926), .IN3(g16627), .IN4(g16744), 
        .QN(n15733) );
  NOR4X0 U16910 ( .IN1(n15734), .IN2(g14451), .IN3(n15735), .IN4(n15736), .QN(
        g24271) );
  NOR2X0 U16911 ( .IN1(n5699), .IN2(g11388), .QN(n15736) );
  NOR2X0 U16912 ( .IN1(n8573), .IN2(g13926), .QN(n15735) );
  NAND3X0 U16913 ( .IN1(n8559), .IN2(n9315), .IN3(n8674), .QN(n15734) );
  NOR2X0 U16914 ( .IN1(n8578), .IN2(n15737), .QN(g24270) );
  NOR2X0 U16915 ( .IN1(n9413), .IN2(n15738), .QN(n15737) );
  NAND2X0 U16916 ( .IN1(n15739), .IN2(n15740), .QN(g24269) );
  NAND2X0 U16917 ( .IN1(n9446), .IN2(g3338), .QN(n15740) );
  NAND3X0 U16918 ( .IN1(n8577), .IN2(n15738), .IN3(n9339), .QN(n15739) );
  NAND2X0 U16919 ( .IN1(n15741), .IN2(n15742), .QN(g24268) );
  NAND2X0 U16920 ( .IN1(test_so91), .IN2(n9514), .QN(n15742) );
  NAND3X0 U16921 ( .IN1(n15743), .IN2(n15738), .IN3(n9339), .QN(n15741) );
  INVX0 U16922 ( .INP(n15744), .ZN(n15738) );
  NOR2X0 U16923 ( .IN1(n15745), .IN2(n5527), .QN(n15744) );
  NAND2X0 U16924 ( .IN1(n5527), .IN2(n15745), .QN(n15743) );
  NAND4X0 U16925 ( .IN1(g11349), .IN2(g13895), .IN3(g16603), .IN4(g16718), 
        .QN(n15745) );
  NOR4X0 U16926 ( .IN1(n15746), .IN2(g14421), .IN3(n15747), .IN4(n15748), .QN(
        g24267) );
  NOR2X0 U16927 ( .IN1(n5702), .IN2(g11349), .QN(n15748) );
  NOR2X0 U16928 ( .IN1(n8562), .IN2(g13895), .QN(n15747) );
  NAND3X0 U16929 ( .IN1(n8547), .IN2(n9315), .IN3(n8645), .QN(n15746) );
  NAND2X0 U16930 ( .IN1(n15749), .IN2(n15750), .QN(g24266) );
  NAND2X0 U16931 ( .IN1(n9446), .IN2(g2841), .QN(n15750) );
  NAND3X0 U16932 ( .IN1(test_so9), .IN2(n8368), .IN3(n9339), .QN(n15749) );
  NAND3X0 U16933 ( .IN1(n15751), .IN2(n15752), .IN3(n9664), .QN(g24263) );
  NAND2X0 U16934 ( .IN1(n5963), .IN2(n9370), .QN(n9664) );
  NAND2X0 U16935 ( .IN1(n5299), .IN2(n9370), .QN(n15752) );
  INVX0 U16936 ( .INP(n15753), .ZN(n15751) );
  NOR2X0 U16937 ( .IN1(n9360), .IN2(n8368), .QN(n15753) );
  NAND3X0 U16938 ( .IN1(n15754), .IN2(n15755), .IN3(n15756), .QN(g24262) );
  NAND2X0 U16939 ( .IN1(n15757), .IN2(n8720), .QN(n15756) );
  NAND3X0 U16940 ( .IN1(n15758), .IN2(g1564), .IN3(n9341), .QN(n15755) );
  NAND2X0 U16941 ( .IN1(n9446), .IN2(g1548), .QN(n15754) );
  NAND2X0 U16942 ( .IN1(n15416), .IN2(n15759), .QN(g24261) );
  NAND2X0 U16943 ( .IN1(n9446), .IN2(g1585), .QN(n15759) );
  NOR2X0 U16944 ( .IN1(n15760), .IN2(n15761), .QN(g24260) );
  NOR2X0 U16945 ( .IN1(n15762), .IN2(g1430), .QN(n15761) );
  NOR2X0 U16946 ( .IN1(n5546), .IN2(n9401), .QN(n15762) );
  NOR2X0 U16947 ( .IN1(n9415), .IN2(n15758), .QN(n15760) );
  NAND2X0 U16948 ( .IN1(n15416), .IN2(n15763), .QN(g24259) );
  NAND2X0 U16949 ( .IN1(n9446), .IN2(g1579), .QN(n15763) );
  NAND2X0 U16950 ( .IN1(n15764), .IN2(n15765), .QN(g24258) );
  NAND2X0 U16951 ( .IN1(n9365), .IN2(g496), .QN(n15765) );
  NAND2X0 U16952 ( .IN1(n9445), .IN2(g1554), .QN(n15764) );
  NOR2X0 U16953 ( .IN1(n15766), .IN2(n15767), .QN(g24257) );
  INVX0 U16954 ( .INP(n15768), .ZN(n15767) );
  NAND2X0 U16955 ( .IN1(g1333), .IN2(n15769), .QN(n15768) );
  NOR2X0 U16956 ( .IN1(n15769), .IN2(g1333), .QN(n15766) );
  NAND3X0 U16957 ( .IN1(n15770), .IN2(n15771), .IN3(n15772), .QN(g24256) );
  NAND2X0 U16958 ( .IN1(n15769), .IN2(n15773), .QN(n15772) );
  NOR2X0 U16959 ( .IN1(n15774), .IN2(n9396), .QN(n15769) );
  NAND3X0 U16960 ( .IN1(n15775), .IN2(n15774), .IN3(n9341), .QN(n15771) );
  NAND4X0 U16961 ( .IN1(n14996), .IN2(n9807), .IN3(n15776), .IN4(n15777), .QN(
        n15774) );
  NAND2X0 U16962 ( .IN1(test_so68), .IN2(g1579), .QN(n15777) );
  NAND2X0 U16963 ( .IN1(n8436), .IN2(n8875), .QN(n15776) );
  INVX0 U16964 ( .INP(n15773), .ZN(n15775) );
  NAND3X0 U16965 ( .IN1(n8797), .IN2(n15415), .IN3(n8798), .QN(n15773) );
  INVX0 U16966 ( .INP(n15412), .ZN(n15415) );
  NAND3X0 U16967 ( .IN1(n5302), .IN2(n5616), .IN3(n5401), .QN(n15412) );
  NAND2X0 U16968 ( .IN1(n9445), .IN2(g1339), .QN(n15770) );
  NAND3X0 U16969 ( .IN1(n15778), .IN2(n15779), .IN3(n15780), .QN(g24255) );
  INVX0 U16970 ( .INP(n15781), .ZN(n15780) );
  NOR2X0 U16971 ( .IN1(n15416), .IN2(n8442), .QN(n15781) );
  NAND3X0 U16972 ( .IN1(n8442), .IN2(g10527), .IN3(n9341), .QN(n15779) );
  NAND2X0 U16973 ( .IN1(n9445), .IN2(g1589), .QN(n15778) );
  INVX0 U16974 ( .INP(n15782), .ZN(g24254) );
  NAND4X0 U16975 ( .IN1(n8442), .IN2(n15783), .IN3(n8443), .IN4(n8444), .QN(
        n15782) );
  NOR2X0 U16976 ( .IN1(n15784), .IN2(n9395), .QN(n15783) );
  INVX0 U16977 ( .INP(n15785), .ZN(n15784) );
  NAND3X0 U16978 ( .IN1(n15786), .IN2(g1554), .IN3(n15390), .QN(n15785) );
  NOR2X0 U16979 ( .IN1(n15758), .IN2(n8720), .QN(n15390) );
  INVX0 U16980 ( .INP(n15757), .ZN(n15758) );
  NOR2X0 U16981 ( .IN1(n8721), .IN2(n5546), .QN(n15757) );
  NAND2X0 U16982 ( .IN1(n14996), .IN2(n9807), .QN(n15786) );
  NOR2X0 U16983 ( .IN1(g1312), .IN2(g1351), .QN(n9807) );
  NOR2X0 U16984 ( .IN1(n14706), .IN2(n14707), .QN(n14996) );
  NOR2X0 U16985 ( .IN1(g1333), .IN2(test_so68), .QN(n14707) );
  NAND2X0 U16986 ( .IN1(n15787), .IN2(n15788), .QN(n14706) );
  NAND2X0 U16987 ( .IN1(test_so68), .IN2(g1339), .QN(n15788) );
  NAND2X0 U16988 ( .IN1(n5381), .IN2(n8875), .QN(n15787) );
  NAND2X0 U16989 ( .IN1(n15789), .IN2(n15790), .QN(g24253) );
  NAND2X0 U16990 ( .IN1(n9445), .IN2(g1306), .QN(n15790) );
  NAND2X0 U16991 ( .IN1(n15791), .IN2(n9369), .QN(n15789) );
  NAND2X0 U16992 ( .IN1(n15792), .IN2(n15793), .QN(n15791) );
  NAND2X0 U16993 ( .IN1(n5302), .IN2(g1532), .QN(n15793) );
  NAND2X0 U16994 ( .IN1(g7946), .IN2(g1521), .QN(n15792) );
  NAND2X0 U16995 ( .IN1(n15794), .IN2(n15795), .QN(g24252) );
  NAND2X0 U16996 ( .IN1(test_so49), .IN2(n9515), .QN(n15795) );
  NAND2X0 U16997 ( .IN1(n15796), .IN2(n9369), .QN(n15794) );
  NAND2X0 U16998 ( .IN1(n15797), .IN2(n15798), .QN(n15796) );
  NAND2X0 U16999 ( .IN1(n5302), .IN2(g1521), .QN(n15798) );
  NAND2X0 U17000 ( .IN1(g7946), .IN2(g1339), .QN(n15797) );
  NAND2X0 U17001 ( .IN1(n15799), .IN2(n15800), .QN(g24251) );
  NAND2X0 U17002 ( .IN1(n14032), .IN2(g1442), .QN(n15800) );
  NAND2X0 U17003 ( .IN1(test_so12), .IN2(n15407), .QN(n15799) );
  NAND2X0 U17004 ( .IN1(n15801), .IN2(n15802), .QN(g24250) );
  NAND2X0 U17005 ( .IN1(test_so12), .IN2(n14032), .QN(n15802) );
  NAND2X0 U17006 ( .IN1(n15407), .IN2(g1489), .QN(n15801) );
  INVX0 U17007 ( .INP(n14032), .ZN(n15407) );
  NAND2X0 U17008 ( .IN1(n15803), .IN2(n15804), .QN(g24249) );
  NAND3X0 U17009 ( .IN1(n8717), .IN2(n9313), .IN3(n14037), .QN(n15804) );
  INVX0 U17010 ( .INP(n15805), .ZN(n15803) );
  NOR2X0 U17011 ( .IN1(n15806), .IN2(n5850), .QN(n15805) );
  NOR2X0 U17012 ( .IN1(n14032), .IN2(n15807), .QN(n15806) );
  NOR2X0 U17013 ( .IN1(n9418), .IN2(test_so12), .QN(n15807) );
  NOR2X0 U17014 ( .IN1(n14037), .IN2(n9396), .QN(n14032) );
  NOR3X0 U17015 ( .IN1(n8798), .IN2(test_so49), .IN3(g1514), .QN(n14037) );
  NAND3X0 U17016 ( .IN1(n15808), .IN2(n15809), .IN3(n15810), .QN(g24248) );
  NAND2X0 U17017 ( .IN1(n15811), .IN2(n15812), .QN(n15810) );
  NAND2X0 U17018 ( .IN1(n8450), .IN2(n15813), .QN(n15812) );
  INVX0 U17019 ( .INP(n15814), .ZN(n15811) );
  NOR2X0 U17020 ( .IN1(n15813), .IN2(n8450), .QN(n15814) );
  NAND2X0 U17021 ( .IN1(n5655), .IN2(n9369), .QN(n15813) );
  NAND2X0 U17022 ( .IN1(n11853), .IN2(g1395), .QN(n15809) );
  NAND2X0 U17023 ( .IN1(n5401), .IN2(n9369), .QN(n15808) );
  NOR2X0 U17024 ( .IN1(g1249), .IN2(n15416), .QN(g24247) );
  INVX0 U17025 ( .INP(n11853), .ZN(n15416) );
  NOR2X0 U17026 ( .IN1(n9417), .IN2(n5655), .QN(n11853) );
  NAND3X0 U17027 ( .IN1(n15815), .IN2(n15816), .IN3(n15817), .QN(g24246) );
  NAND2X0 U17028 ( .IN1(n15818), .IN2(n8722), .QN(n15817) );
  NAND3X0 U17029 ( .IN1(n15819), .IN2(g1221), .IN3(n9341), .QN(n15816) );
  NAND2X0 U17030 ( .IN1(n9445), .IN2(g1205), .QN(n15815) );
  NAND2X0 U17031 ( .IN1(n15469), .IN2(n15820), .QN(g24245) );
  NAND2X0 U17032 ( .IN1(n9445), .IN2(g30332), .QN(n15820) );
  NOR2X0 U17033 ( .IN1(n15821), .IN2(n15822), .QN(g24244) );
  NOR2X0 U17034 ( .IN1(n15823), .IN2(g1087), .QN(n15822) );
  NOR2X0 U17035 ( .IN1(n5547), .IN2(n9396), .QN(n15823) );
  NOR2X0 U17036 ( .IN1(n9419), .IN2(n15819), .QN(n15821) );
  INVX0 U17037 ( .INP(n15818), .ZN(n15819) );
  NAND2X0 U17038 ( .IN1(n15469), .IN2(n15824), .QN(g24243) );
  NAND2X0 U17039 ( .IN1(n9445), .IN2(g1236), .QN(n15824) );
  NAND2X0 U17040 ( .IN1(n15825), .IN2(n15826), .QN(g24242) );
  NAND2X0 U17041 ( .IN1(n9365), .IN2(g29215), .QN(n15826) );
  NAND2X0 U17042 ( .IN1(test_so76), .IN2(n9514), .QN(n15825) );
  NOR2X0 U17043 ( .IN1(n15827), .IN2(n15828), .QN(g24241) );
  INVX0 U17044 ( .INP(n15829), .ZN(n15828) );
  NAND2X0 U17045 ( .IN1(g990), .IN2(n15830), .QN(n15829) );
  NOR2X0 U17046 ( .IN1(n15830), .IN2(g990), .QN(n15827) );
  NAND3X0 U17047 ( .IN1(n15831), .IN2(n15832), .IN3(n15833), .QN(g24240) );
  NAND2X0 U17048 ( .IN1(n15830), .IN2(n15834), .QN(n15833) );
  NOR2X0 U17049 ( .IN1(n15835), .IN2(n9396), .QN(n15830) );
  NAND3X0 U17050 ( .IN1(n15836), .IN2(n15835), .IN3(n9343), .QN(n15832) );
  NAND3X0 U17051 ( .IN1(n15837), .IN2(n14797), .IN3(n15033), .QN(n15835) );
  NAND2X0 U17052 ( .IN1(n15838), .IN2(n15839), .QN(n15837) );
  NAND2X0 U17053 ( .IN1(n8435), .IN2(g979), .QN(n15839) );
  NAND2X0 U17054 ( .IN1(n5320), .IN2(g1236), .QN(n15838) );
  INVX0 U17055 ( .INP(n15834), .ZN(n15836) );
  NAND3X0 U17056 ( .IN1(n8803), .IN2(n15468), .IN3(n8804), .QN(n15834) );
  INVX0 U17057 ( .INP(n15470), .ZN(n15468) );
  NAND3X0 U17058 ( .IN1(n5304), .IN2(n5622), .IN3(n5392), .QN(n15470) );
  NAND2X0 U17059 ( .IN1(n9444), .IN2(g996), .QN(n15831) );
  NAND3X0 U17060 ( .IN1(n15840), .IN2(n15841), .IN3(n15842), .QN(g24239) );
  NAND2X0 U17061 ( .IN1(n11867), .IN2(g17400), .QN(n15842) );
  NAND3X0 U17062 ( .IN1(n8438), .IN2(g10500), .IN3(n9343), .QN(n15841) );
  NAND2X0 U17063 ( .IN1(n9444), .IN2(g1246), .QN(n15840) );
  INVX0 U17064 ( .INP(n15843), .ZN(g24238) );
  NAND4X0 U17065 ( .IN1(n15844), .IN2(n15845), .IN3(n8438), .IN4(n8433), .QN(
        n15843) );
  NOR2X0 U17066 ( .IN1(n9419), .IN2(test_so44), .QN(n15845) );
  NAND3X0 U17067 ( .IN1(test_so76), .IN2(n15846), .IN3(n15445), .QN(n15844) );
  INVX0 U17068 ( .INP(n15444), .ZN(n15445) );
  NAND2X0 U17069 ( .IN1(n15818), .IN2(g1221), .QN(n15444) );
  NOR2X0 U17070 ( .IN1(n8723), .IN2(n5547), .QN(n15818) );
  NAND2X0 U17071 ( .IN1(n14797), .IN2(n15033), .QN(n15846) );
  NOR2X0 U17072 ( .IN1(n14721), .IN2(n14722), .QN(n15033) );
  NOR2X0 U17073 ( .IN1(g990), .IN2(g979), .QN(n14722) );
  INVX0 U17074 ( .INP(n14719), .ZN(n14721) );
  NAND2X0 U17075 ( .IN1(n15847), .IN2(n15848), .QN(n14719) );
  NAND2X0 U17076 ( .IN1(n8808), .IN2(g979), .QN(n15848) );
  NAND2X0 U17077 ( .IN1(n5320), .IN2(g996), .QN(n15847) );
  INVX0 U17078 ( .INP(n4837), .ZN(n14797) );
  NAND2X0 U17079 ( .IN1(n5321), .IN2(n8890), .QN(n4837) );
  NAND2X0 U17080 ( .IN1(n15849), .IN2(n15850), .QN(g24237) );
  NAND2X0 U17081 ( .IN1(n9444), .IN2(g962), .QN(n15850) );
  NAND2X0 U17082 ( .IN1(n15851), .IN2(n9369), .QN(n15849) );
  NAND2X0 U17083 ( .IN1(n15852), .IN2(n15853), .QN(n15851) );
  NAND2X0 U17084 ( .IN1(n5304), .IN2(g1189), .QN(n15853) );
  NAND2X0 U17085 ( .IN1(g7916), .IN2(g1178), .QN(n15852) );
  NAND2X0 U17086 ( .IN1(n15854), .IN2(n15855), .QN(g24236) );
  NAND2X0 U17087 ( .IN1(n9444), .IN2(g1183), .QN(n15855) );
  NAND2X0 U17088 ( .IN1(n15856), .IN2(n9368), .QN(n15854) );
  NAND2X0 U17089 ( .IN1(n15857), .IN2(n15858), .QN(n15856) );
  NAND2X0 U17090 ( .IN1(n5304), .IN2(g1178), .QN(n15858) );
  INVX0 U17091 ( .INP(n13534), .ZN(n15857) );
  NOR2X0 U17092 ( .IN1(n5304), .IN2(n8808), .QN(n13534) );
  NAND2X0 U17093 ( .IN1(n15859), .IN2(n15860), .QN(g24235) );
  NAND2X0 U17094 ( .IN1(test_so7), .IN2(n14074), .QN(n15860) );
  NAND2X0 U17095 ( .IN1(n15461), .IN2(g1152), .QN(n15859) );
  NAND2X0 U17096 ( .IN1(n15861), .IN2(n15862), .QN(g24234) );
  NAND2X0 U17097 ( .IN1(n14074), .IN2(g1152), .QN(n15862) );
  NAND2X0 U17098 ( .IN1(n15461), .IN2(g1146), .QN(n15861) );
  NAND2X0 U17099 ( .IN1(n15863), .IN2(n15864), .QN(g24233) );
  NAND3X0 U17100 ( .IN1(n9347), .IN2(n8865), .IN3(n14079), .QN(n15864) );
  NAND2X0 U17101 ( .IN1(n15865), .IN2(g1146), .QN(n15863) );
  NAND2X0 U17102 ( .IN1(n15461), .IN2(n15866), .QN(n15865) );
  NAND2X0 U17103 ( .IN1(n5618), .IN2(n9368), .QN(n15866) );
  INVX0 U17104 ( .INP(n14074), .ZN(n15461) );
  NOR2X0 U17105 ( .IN1(n14079), .IN2(n9397), .QN(n14074) );
  NOR3X0 U17106 ( .IN1(g1171), .IN2(n8804), .IN3(g1183), .QN(n14079) );
  NAND3X0 U17107 ( .IN1(n15867), .IN2(n15868), .IN3(n15869), .QN(g24232) );
  NAND2X0 U17108 ( .IN1(n15870), .IN2(n15871), .QN(n15869) );
  NAND2X0 U17109 ( .IN1(n8451), .IN2(n15872), .QN(n15871) );
  INVX0 U17110 ( .INP(n15873), .ZN(n15870) );
  NOR2X0 U17111 ( .IN1(n15872), .IN2(n8451), .QN(n15873) );
  NAND2X0 U17112 ( .IN1(n5654), .IN2(n9368), .QN(n15872) );
  NAND2X0 U17113 ( .IN1(n11867), .IN2(g1052), .QN(n15868) );
  NAND2X0 U17114 ( .IN1(n5392), .IN2(n9368), .QN(n15867) );
  NOR2X0 U17115 ( .IN1(g904), .IN2(n15469), .QN(g24231) );
  INVX0 U17116 ( .INP(n11867), .ZN(n15469) );
  NOR2X0 U17117 ( .IN1(n9420), .IN2(n5654), .QN(n11867) );
  NAND2X0 U17118 ( .IN1(n15874), .IN2(n15875), .QN(g24216) );
  NAND2X0 U17119 ( .IN1(n14147), .IN2(g847), .QN(n15875) );
  NAND2X0 U17120 ( .IN1(n15510), .IN2(g854), .QN(n15874) );
  NAND2X0 U17121 ( .IN1(n15876), .IN2(n15877), .QN(g24215) );
  NAND2X0 U17122 ( .IN1(n15878), .IN2(g837), .QN(n15877) );
  NAND2X0 U17123 ( .IN1(n15510), .IN2(n15879), .QN(n15878) );
  NAND3X0 U17124 ( .IN1(n15880), .IN2(n9313), .IN3(n15881), .QN(n15879) );
  NAND2X0 U17125 ( .IN1(g827), .IN2(g832), .QN(n15881) );
  NAND2X0 U17126 ( .IN1(g847), .IN2(g812), .QN(n15880) );
  NAND2X0 U17127 ( .IN1(n15882), .IN2(g703), .QN(n15876) );
  NAND2X0 U17128 ( .IN1(n15883), .IN2(n9368), .QN(n15882) );
  NAND2X0 U17129 ( .IN1(n5562), .IN2(n15495), .QN(n15883) );
  NOR2X0 U17130 ( .IN1(n14151), .IN2(n5709), .QN(n15495) );
  NAND3X0 U17131 ( .IN1(n15884), .IN2(n15885), .IN3(n15886), .QN(g24214) );
  NAND2X0 U17132 ( .IN1(n15887), .IN2(g703), .QN(n15886) );
  NAND2X0 U17133 ( .IN1(n15082), .IN2(n15888), .QN(n15887) );
  NAND2X0 U17134 ( .IN1(n15084), .IN2(n9368), .QN(n15888) );
  NAND2X0 U17135 ( .IN1(g812), .IN2(g837), .QN(n15084) );
  NOR2X0 U17136 ( .IN1(n14147), .IN2(n15889), .QN(n15082) );
  NOR2X0 U17137 ( .IN1(g847), .IN2(n9398), .QN(n15889) );
  NAND2X0 U17138 ( .IN1(n9444), .IN2(g847), .QN(n15885) );
  NAND4X0 U17139 ( .IN1(g817), .IN2(g723), .IN3(n15890), .IN4(n5709), .QN(
        n15884) );
  NOR2X0 U17140 ( .IN1(n5422), .IN2(n15511), .QN(n15890) );
  INVX0 U17141 ( .INP(n14152), .ZN(n15511) );
  NAND2X0 U17142 ( .IN1(n15891), .IN2(n15892), .QN(g24211) );
  NAND2X0 U17143 ( .IN1(n2404), .IN2(n15893), .QN(n15892) );
  INVX0 U17144 ( .INP(n15894), .ZN(n15893) );
  NOR2X0 U17145 ( .IN1(test_so41), .IN2(n5520), .QN(n15894) );
  INVX0 U17146 ( .INP(n15895), .ZN(n15891) );
  NOR2X0 U17147 ( .IN1(n9358), .IN2(n5492), .QN(n15895) );
  NOR3X0 U17148 ( .IN1(n12444), .IN2(n9384), .IN3(n15896), .QN(g24210) );
  NOR2X0 U17149 ( .IN1(n15897), .IN2(n15898), .QN(n15896) );
  NOR2X0 U17150 ( .IN1(n5606), .IN2(n5402), .QN(n15898) );
  NOR2X0 U17151 ( .IN1(n13562), .IN2(n8871), .QN(n15897) );
  NOR2X0 U17152 ( .IN1(g168), .IN2(g174), .QN(n13562) );
  NAND3X0 U17153 ( .IN1(g518), .IN2(g203), .IN3(n5548), .QN(n12444) );
  NAND2X0 U17154 ( .IN1(n15899), .IN2(n15900), .QN(g24209) );
  NAND2X0 U17155 ( .IN1(n14152), .IN2(g446), .QN(n15900) );
  NAND2X0 U17156 ( .IN1(n14147), .IN2(g417), .QN(n15899) );
  NAND3X0 U17157 ( .IN1(n15901), .IN2(n15902), .IN3(n15903), .QN(g24208) );
  NAND2X0 U17158 ( .IN1(n9444), .IN2(g424), .QN(n15903) );
  NAND2X0 U17159 ( .IN1(n14152), .IN2(g246), .QN(n15902) );
  NAND2X0 U17160 ( .IN1(n14147), .IN2(g475), .QN(n15901) );
  NAND2X0 U17161 ( .IN1(n15904), .IN2(n15905), .QN(g24207) );
  NAND2X0 U17162 ( .IN1(n14147), .IN2(g441), .QN(n15905) );
  NAND2X0 U17163 ( .IN1(n15510), .IN2(g475), .QN(n15904) );
  NAND2X0 U17164 ( .IN1(n15906), .IN2(n15907), .QN(g24206) );
  NAND2X0 U17165 ( .IN1(n14147), .IN2(g437), .QN(n15907) );
  NAND2X0 U17166 ( .IN1(n15510), .IN2(g441), .QN(n15906) );
  NAND3X0 U17167 ( .IN1(n15908), .IN2(n15909), .IN3(n15910), .QN(g24205) );
  NAND2X0 U17168 ( .IN1(n9444), .IN2(g437), .QN(n15910) );
  NAND2X0 U17169 ( .IN1(n14152), .IN2(g269), .QN(n15909) );
  NAND2X0 U17170 ( .IN1(test_so23), .IN2(n14147), .QN(n15908) );
  NAND2X0 U17171 ( .IN1(n15911), .IN2(n15912), .QN(g24204) );
  NAND2X0 U17172 ( .IN1(n14147), .IN2(g429), .QN(n15912) );
  NAND2X0 U17173 ( .IN1(test_so23), .IN2(n15510), .QN(n15911) );
  NAND2X0 U17174 ( .IN1(n15913), .IN2(n15914), .QN(g24203) );
  NAND2X0 U17175 ( .IN1(n14147), .IN2(g401), .QN(n15914) );
  NAND2X0 U17176 ( .IN1(n15510), .IN2(g429), .QN(n15913) );
  NAND2X0 U17177 ( .IN1(n15915), .IN2(n15916), .QN(g24202) );
  NAND2X0 U17178 ( .IN1(n14147), .IN2(g424), .QN(n15916) );
  NAND2X0 U17179 ( .IN1(n15510), .IN2(g411), .QN(n15915) );
  NAND2X0 U17180 ( .IN1(n15917), .IN2(n15918), .QN(g24201) );
  NAND2X0 U17181 ( .IN1(n14147), .IN2(g405), .QN(n15918) );
  NAND2X0 U17182 ( .IN1(n15510), .IN2(g392), .QN(n15917) );
  INVX0 U17183 ( .INP(n14147), .ZN(n15510) );
  NAND3X0 U17184 ( .IN1(n15919), .IN2(n15920), .IN3(n15921), .QN(g24200) );
  NAND2X0 U17185 ( .IN1(n9465), .IN2(g401), .QN(n15921) );
  NAND3X0 U17186 ( .IN1(n5821), .IN2(g854), .IN3(n14152), .QN(n15920) );
  NOR2X0 U17187 ( .IN1(n14151), .IN2(n9393), .QN(n14152) );
  INVX0 U17188 ( .INP(n4948), .ZN(n14151) );
  NAND2X0 U17189 ( .IN1(n14147), .IN2(g392), .QN(n15919) );
  NOR2X0 U17190 ( .IN1(n9421), .IN2(n4948), .QN(n14147) );
  NOR2X0 U17191 ( .IN1(g22), .IN2(g25), .QN(g23190) );
  NAND2X0 U17192 ( .IN1(n15922), .IN2(n15923), .QN(g21901) );
  NAND2X0 U17193 ( .IN1(n9466), .IN2(g2946), .QN(n15923) );
  NAND2X0 U17194 ( .IN1(n15924), .IN2(n9366), .QN(n15922) );
  NAND2X0 U17195 ( .IN1(n15925), .IN2(n15926), .QN(n15924) );
  NAND2X0 U17196 ( .IN1(n5694), .IN2(g4180), .QN(n15926) );
  NAND2X0 U17197 ( .IN1(n5380), .IN2(n15927), .QN(n15925) );
  NAND2X0 U17198 ( .IN1(n5694), .IN2(n15928), .QN(n15927) );
  NAND4X0 U17199 ( .IN1(n15972), .IN2(n8460), .IN3(n15971), .IN4(n15929), .QN(
        n15928) );
  NOR4X0 U17200 ( .IN1(test_so86), .IN2(test_so39), .IN3(g8787), .IN4(g8788), 
        .QN(n15929) );
  NAND2X0 U17201 ( .IN1(n15930), .IN2(n15931), .QN(g21900) );
  INVX0 U17202 ( .INP(n15932), .ZN(n15931) );
  NOR2X0 U17203 ( .IN1(n9359), .IN2(n8425), .QN(n15932) );
  NAND3X0 U17204 ( .IN1(n8372), .IN2(n8371), .IN3(n9343), .QN(n15930) );
  NAND2X0 U17205 ( .IN1(n15933), .IN2(n15934), .QN(g21899) );
  NAND2X0 U17206 ( .IN1(n15935), .IN2(g4291), .QN(n15934) );
  NAND2X0 U17207 ( .IN1(n9365), .IN2(g9019), .QN(n15935) );
  NAND3X0 U17208 ( .IN1(n9349), .IN2(g9019), .IN3(n8749), .QN(n15933) );
  NAND2X0 U17209 ( .IN1(n15936), .IN2(n15937), .QN(g21898) );
  NAND2X0 U17210 ( .IN1(n8749), .IN2(n9368), .QN(n15937) );
  NAND2X0 U17211 ( .IN1(n9467), .IN2(g4284), .QN(n15936) );
  NAND2X0 U17212 ( .IN1(n15938), .IN2(n15939), .QN(g21897) );
  NAND2X0 U17213 ( .IN1(n15940), .IN2(g4281), .QN(n15939) );
  NAND2X0 U17214 ( .IN1(n9365), .IN2(g8839), .QN(n15940) );
  NAND3X0 U17215 ( .IN1(n9347), .IN2(g8839), .IN3(n8750), .QN(n15938) );
  NAND2X0 U17216 ( .IN1(n15941), .IN2(n15942), .QN(g21896) );
  NAND2X0 U17217 ( .IN1(n8750), .IN2(n9366), .QN(n15942) );
  NAND2X0 U17218 ( .IN1(n9470), .IN2(g4245), .QN(n15941) );
  NAND2X0 U17219 ( .IN1(n15943), .IN2(n15944), .QN(g21895) );
  NAND2X0 U17220 ( .IN1(n15945), .IN2(g4264), .QN(n15944) );
  NAND2X0 U17221 ( .IN1(n15946), .IN2(n9368), .QN(n15945) );
  NAND2X0 U17222 ( .IN1(n5763), .IN2(g4258), .QN(n15946) );
  INVX0 U17223 ( .INP(n15947), .ZN(n15943) );
  NOR2X0 U17224 ( .IN1(n15697), .IN2(n5763), .QN(n15947) );
  NOR2X0 U17225 ( .IN1(g21893), .IN2(n15948), .QN(n15697) );
  NOR2X0 U17226 ( .IN1(g4264), .IN2(n9403), .QN(n15948) );
  NAND2X0 U17227 ( .IN1(n15949), .IN2(n15950), .QN(g21894) );
  NAND2X0 U17228 ( .IN1(n15951), .IN2(g4258), .QN(n15950) );
  NAND2X0 U17229 ( .IN1(n9365), .IN2(g4264), .QN(n15951) );
  NAND2X0 U17230 ( .IN1(g21893), .IN2(g4264), .QN(n15949) );
  NOR2X0 U17231 ( .IN1(g4258), .IN2(n9404), .QN(g21893) );
  NAND2X0 U17232 ( .IN1(n15952), .IN2(n15953), .QN(g21892) );
  NAND2X0 U17233 ( .IN1(n8425), .IN2(n9366), .QN(n15953) );
  NAND2X0 U17234 ( .IN1(n9487), .IN2(g4273), .QN(n15952) );
  NAND2X0 U17235 ( .IN1(n15954), .IN2(n15955), .QN(g21891) );
  NAND2X0 U17236 ( .IN1(n9508), .IN2(g4180), .QN(n15955) );
  NAND2X0 U17237 ( .IN1(n15703), .IN2(n9366), .QN(n15954) );
  NAND2X0 U17238 ( .IN1(n15956), .IN2(n15957), .QN(n15703) );
  NAND2X0 U17239 ( .IN1(n8727), .IN2(g4253), .QN(n15957) );
  NAND2X0 U17240 ( .IN1(n8726), .IN2(n5484), .QN(n15956) );
  NOR2X0 U17241 ( .IN1(n9356), .IN2(DFF_1381_n1), .QN(g21727) );
  NOR2X0 U17242 ( .IN1(n5750), .IN2(n9355), .QN(g18597) );
  INVX0 U17243 ( .INP(g5), .ZN(g12833) );
  NOR2X0 U5116_U2 ( .IN1(g34783), .IN2(n2730), .QN(U5116_n1) );
  INVX0 U5116_U1 ( .INP(U5116_n1), .ZN(g34221) );
  NOR2X0 U5126_U2 ( .IN1(n1426), .IN2(n4896), .QN(U5126_n1) );
  INVX0 U5126_U1 ( .INP(U5126_n1), .ZN(n4895) );
  NOR2X0 U5127_U2 ( .IN1(n4837), .IN2(n4921), .QN(U5127_n1) );
  INVX0 U5127_U1 ( .INP(U5127_n1), .ZN(n4920) );
  NOR2X0 U5128_U2 ( .IN1(n822), .IN2(n1296), .QN(U5128_n1) );
  INVX0 U5128_U1 ( .INP(U5128_n1), .ZN(n5045) );
  NOR2X0 U5129_U2 ( .IN1(g559), .IN2(g9048), .QN(U5129_n1) );
  INVX0 U5129_U1 ( .INP(U5129_n1), .ZN(n4959) );
  INVX0 U5353_U2 ( .INP(n5960), .ZN(U5353_n1) );
  NOR2X0 U5353_U1 ( .IN1(n8850), .IN2(U5353_n1), .QN(n4689) );
  INVX0 U5355_U2 ( .INP(n5961), .ZN(U5355_n1) );
  NOR2X0 U5355_U1 ( .IN1(n8845), .IN2(U5355_n1), .QN(n4708) );
  INVX0 U5961_U2 ( .INP(n3593), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n3589), .IN2(U5961_n1), .QN(n3595) );
  INVX0 U5962_U2 ( .INP(n3574), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n3570), .IN2(U5962_n1), .QN(n3576) );
  INVX0 U5963_U2 ( .INP(n3517), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n3513), .IN2(U5963_n1), .QN(n3519) );
  INVX0 U5964_U2 ( .INP(n3628), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n3624), .IN2(U5964_n1), .QN(n3630) );
  INVX0 U5965_U2 ( .INP(n3555), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n3551), .IN2(U5965_n1), .QN(n3557) );
  INVX0 U5966_U2 ( .INP(n3646), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n3642), .IN2(U5966_n1), .QN(n3648) );
  INVX0 U5967_U2 ( .INP(n3536), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n3532), .IN2(U5967_n1), .QN(n3538) );
  INVX0 U5968_U2 ( .INP(n3611), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n3607), .IN2(U5968_n1), .QN(n3613) );
  INVX0 U6100_U2 ( .INP(n3635), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n9408), .IN2(U6100_n1), .QN(n4888) );
  INVX0 U6211_U2 ( .INP(n3623), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n1774), .IN2(U6211_n1), .QN(n3622) );
  INVX0 U6212_U2 ( .INP(n3587), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n3588), .IN2(U6212_n1), .QN(n3586) );
  INVX0 U6213_U2 ( .INP(n3605), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n3606), .IN2(U6213_n1), .QN(n3604) );
  INVX0 U6214_U2 ( .INP(n3568), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n3569), .IN2(U6214_n1), .QN(n3567) );
  INVX0 U6215_U2 ( .INP(n3549), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n3550), .IN2(U6215_n1), .QN(n3548) );
  INVX0 U6216_U2 ( .INP(n3512), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n3006), .IN2(U6216_n1), .QN(n3511) );
  INVX0 U6217_U2 ( .INP(n3531), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n3007), .IN2(U6217_n1), .QN(n3530) );
  INVX0 U6218_U2 ( .INP(n3641), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n3003), .IN2(U6218_n1), .QN(n3640) );
  INVX0 U6279_U2 ( .INP(n4537), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n5337), .IN2(U6279_n1), .QN(n4201) );
  INVX0 U6280_U2 ( .INP(n4201), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n5336), .IN2(U6280_n1), .QN(n3745) );
  INVX0 U6281_U2 ( .INP(n3745), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n5294), .IN2(U6281_n1), .QN(n3684) );
  INVX0 U6282_U2 ( .INP(n3684), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n5552), .IN2(U6282_n1), .QN(n3274) );
  INVX0 U6283_U2 ( .INP(n3274), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n5472), .IN2(U6283_n1), .QN(n2982) );
  INVX0 U6284_U2 ( .INP(n2982), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n5476), .IN2(U6284_n1), .QN(n2706) );
  INVX0 U6285_U2 ( .INP(n2706), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n5550), .IN2(U6285_n1), .QN(n2649) );
  INVX0 U6286_U2 ( .INP(n2649), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n5473), .IN2(U6286_n1), .QN(n2556) );
  INVX0 U6287_U2 ( .INP(n2556), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n5475), .IN2(U6287_n1), .QN(n2509) );
  INVX0 U6288_U2 ( .INP(n2509), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n5474), .IN2(U6288_n1), .QN(n2487) );
  INVX0 U6289_U2 ( .INP(n2487), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n5339), .IN2(U6289_n1), .QN(n2427) );
  INVX0 U6290_U2 ( .INP(n2427), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n5672), .IN2(U6290_n1), .QN(n2423) );
  INVX0 U6291_U2 ( .INP(n5), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n5335), .IN2(U6291_n1), .QN(n4537) );
  INVX0 U6292_U2 ( .INP(n4959), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n9408), .IN2(U6292_n1), .QN(n2421) );
  INVX0 U6338_U2 ( .INP(n4210), .ZN(U6338_n1) );
  NOR2X1 U6338_U1 ( .IN1(n9407), .IN2(U6338_n1), .QN(n3765) );
  INVX0 U6341_U2 ( .INP(n3765), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n1178), .IN2(U6341_n1), .QN(n3951) );
  INVX0 U6342_U2 ( .INP(n3765), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n763), .IN2(U6342_n1), .QN(n3774) );
  INVX0 U6343_U2 ( .INP(n3765), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n1107), .IN2(U6343_n1), .QN(n3842) );
  INVX0 U6344_U2 ( .INP(n3765), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n1037), .IN2(U6344_n1), .QN(n3808) );
  INVX0 U6345_U2 ( .INP(n3765), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n757), .IN2(U6345_n1), .QN(n3908) );
  INVX0 U6346_U2 ( .INP(n3765), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n73), .IN2(U6346_n1), .QN(n3984) );
  INVX0 U6347_U2 ( .INP(n3765), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n497), .IN2(U6347_n1), .QN(n3875) );
  INVX0 U6348_U2 ( .INP(n3765), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n89), .IN2(U6348_n1), .QN(n4015) );
  INVX0 U6349_U2 ( .INP(n3765), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n759), .IN2(U6349_n1), .QN(n3914) );
  INVX0 U6350_U2 ( .INP(n3765), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n765), .IN2(U6350_n1), .QN(n3780) );
  INVX0 U6351_U2 ( .INP(n3765), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n1179), .IN2(U6351_n1), .QN(n3957) );
  INVX0 U6352_U2 ( .INP(n3765), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n1108), .IN2(U6352_n1), .QN(n3848) );
  INVX0 U6353_U2 ( .INP(n3765), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n74), .IN2(U6353_n1), .QN(n3990) );
  INVX0 U6354_U2 ( .INP(n3765), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n1038), .IN2(U6354_n1), .QN(n3814) );
  INVX0 U6355_U2 ( .INP(n3765), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n499), .IN2(U6355_n1), .QN(n3881) );
  INVX0 U6356_U2 ( .INP(n3765), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n91), .IN2(U6356_n1), .QN(n4022) );
  INVX0 U6357_U2 ( .INP(n3765), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n90), .IN2(U6357_n1), .QN(n4027) );
  INVX0 U6358_U2 ( .INP(n3765), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n764), .IN2(U6358_n1), .QN(n3785) );
  INVX0 U6359_U2 ( .INP(n3765), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n1180), .IN2(U6359_n1), .QN(n3962) );
  INVX0 U6360_U2 ( .INP(n3765), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n1109), .IN2(U6360_n1), .QN(n3853) );
  INVX0 U6361_U2 ( .INP(n3765), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n498), .IN2(U6361_n1), .QN(n3886) );
  INVX0 U6362_U2 ( .INP(n3765), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n1039), .IN2(U6362_n1), .QN(n3819) );
  INVX0 U6363_U2 ( .INP(n3765), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n75), .IN2(U6363_n1), .QN(n3995) );
  INVX0 U6364_U2 ( .INP(n3765), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n758), .IN2(U6364_n1), .QN(n3919) );
  INVX0 U6365_U2 ( .INP(n3682), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n5471), .IN2(U6365_n1), .QN(n3272) );
  INVX0 U6366_U2 ( .INP(n3272), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n5331), .IN2(U6366_n1), .QN(n2980) );
  INVX0 U6367_U2 ( .INP(n2980), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n5332), .IN2(U6367_n1), .QN(n2704) );
  INVX0 U6368_U2 ( .INP(n2704), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n5333), .IN2(U6368_n1), .QN(n2647) );
  INVX0 U6369_U2 ( .INP(n2647), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n5334), .IN2(U6369_n1), .QN(n2554) );
  INVX0 U6370_U2 ( .INP(n2554), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n5330), .IN2(U6370_n1), .QN(n2507) );
  INVX0 U6371_U2 ( .INP(n2507), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n5551), .IN2(U6371_n1), .QN(n2485) );
  INVX0 U6372_U2 ( .INP(n2485), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n5293), .IN2(U6372_n1), .QN(n2425) );
  INVX0 U6373_U2 ( .INP(n2425), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n5292), .IN2(U6373_n1), .QN(n2419) );
  INVX0 U6374_U2 ( .INP(n57), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n5470), .IN2(U6374_n1), .QN(n3682) );
  INVX0 U6375_U2 ( .INP(n2419), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n5291), .IN2(U6375_n1), .QN(n2405) );
  INVX0 U6417_U2 ( .INP(n513), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n9409), .IN2(U6417_n1), .QN(n2404) );
  INVX0 U6446_U2 ( .INP(g110), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n1835), .IN2(U6446_n1), .QN(n3524) );
  INVX0 U6465_U2 ( .INP(n3653), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n5600), .IN2(U6465_n1), .QN(n4388) );
  INVX0 U6497_U2 ( .INP(n826), .ZN(U6497_n1) );
  NOR2X0 U6497_U1 ( .IN1(n3635), .IN2(U6497_n1), .QN(n3005) );
  INVX0 U6523_U2 ( .INP(n4946), .ZN(U6523_n1) );
  NOR2X0 U6523_U1 ( .IN1(n9409), .IN2(U6523_n1), .QN(n4945) );
  INVX0 U6542_U2 ( .INP(n826), .ZN(U6542_n1) );
  NOR2X0 U6542_U1 ( .IN1(n5300), .IN2(U6542_n1), .QN(n3525) );
  INVX0 U6552_U2 ( .INP(n3281), .ZN(U6552_n1) );
  NOR2X0 U6552_U1 ( .IN1(n5676), .IN2(U6552_n1), .QN(n3277) );
  INVX0 U6553_U2 ( .INP(n3276), .ZN(U6553_n1) );
  NOR2X0 U6553_U1 ( .IN1(n5680), .IN2(U6553_n1), .QN(n2989) );
  INVX0 U6554_U2 ( .INP(n3277), .ZN(U6554_n1) );
  NOR2X0 U6554_U1 ( .IN1(n5677), .IN2(U6554_n1), .QN(n2991) );
  INVX0 U6555_U2 ( .INP(n3687), .ZN(U6555_n1) );
  NOR2X0 U6555_U1 ( .IN1(n5561), .IN2(U6555_n1), .QN(n3281) );
  INVX0 U6556_U2 ( .INP(n54), .ZN(U6556_n1) );
  NOR2X0 U6556_U1 ( .IN1(n5679), .IN2(U6556_n1), .QN(n3276) );
  INVX0 U6559_U2 ( .INP(n2991), .ZN(U6559_n1) );
  NOR2X0 U6559_U1 ( .IN1(n5678), .IN2(U6559_n1), .QN(n2710) );
  INVX0 U6560_U2 ( .INP(n2989), .ZN(U6560_n1) );
  NOR2X0 U6560_U1 ( .IN1(n5675), .IN2(U6560_n1), .QN(n2707) );
  INVX0 U6561_U2 ( .INP(n3174), .ZN(U6561_n1) );
  NOR2X0 U6561_U1 ( .IN1(n5327), .IN2(U6561_n1), .QN(n3116) );
  INVX0 U6570_U2 ( .INP(n3362), .ZN(U6570_n1) );
  NOR2X0 U6570_U1 ( .IN1(n5477), .IN2(U6570_n1), .QN(n2527) );
  INVX0 U6911_U2 ( .INP(n3115), .ZN(U6911_n1) );
  NOR2X0 U6911_U1 ( .IN1(n1013), .IN2(U6911_n1), .QN(n3111) );
  INVX0 U6912_U2 ( .INP(n3115), .ZN(U6912_n1) );
  NOR2X0 U6912_U1 ( .IN1(n999), .IN2(U6912_n1), .QN(n3131) );
  INVX0 U6917_U2 ( .INP(n3933), .ZN(U6917_n1) );
  NOR2X0 U6917_U1 ( .IN1(n5350), .IN2(U6917_n1), .QN(n3799) );
  INVX0 U6926_U2 ( .INP(n3664), .ZN(U6926_n1) );
  NOR2X0 U6926_U1 ( .IN1(n5674), .IN2(U6926_n1), .QN(n3662) );
  INVX0 U6927_U2 ( .INP(n3673), .ZN(U6927_n1) );
  NOR2X0 U6927_U1 ( .IN1(n5673), .IN2(U6927_n1), .QN(n3671) );
  INVX0 U6929_U2 ( .INP(n3505), .ZN(U6929_n1) );
  NOR2X0 U6929_U1 ( .IN1(n3506), .IN2(U6929_n1), .QN(n2790) );
  INVX0 U6931_U2 ( .INP(n4490), .ZN(U6931_n1) );
  NOR2X0 U6931_U1 ( .IN1(n5554), .IN2(U6931_n1), .QN(n4178) );
  INVX0 U6932_U2 ( .INP(n4514), .ZN(U6932_n1) );
  NOR2X0 U6932_U1 ( .IN1(n5555), .IN2(U6932_n1), .QN(n4196) );
  INVX0 U6933_U2 ( .INP(n4178), .ZN(U6933_n1) );
  NOR2X0 U6933_U1 ( .IN1(n5558), .IN2(U6933_n1), .QN(n3736) );
  INVX0 U6934_U2 ( .INP(n4196), .ZN(U6934_n1) );
  NOR2X0 U6934_U1 ( .IN1(n5559), .IN2(U6934_n1), .QN(n3741) );
  INVX0 U6935_U2 ( .INP(n3736), .ZN(U6935_n1) );
  NOR2X0 U6935_U1 ( .IN1(n5553), .IN2(U6935_n1), .QN(n3664) );
  INVX0 U6936_U2 ( .INP(n3741), .ZN(U6936_n1) );
  NOR2X0 U6936_U1 ( .IN1(n5560), .IN2(U6936_n1), .QN(n3673) );
  INVX0 U6937_U2 ( .INP(n101), .ZN(U6937_n1) );
  NOR2X0 U6937_U1 ( .IN1(n5303), .IN2(U6937_n1), .QN(n2598) );
  INVX0 U6938_U2 ( .INP(n1266), .ZN(U6938_n1) );
  NOR2X0 U6938_U1 ( .IN1(n5556), .IN2(U6938_n1), .QN(n4490) );
  INVX0 U6939_U2 ( .INP(n266), .ZN(U6939_n1) );
  NOR2X0 U6939_U1 ( .IN1(n5557), .IN2(U6939_n1), .QN(n4514) );
  INVX0 U6940_U2 ( .INP(n905), .ZN(U6940_n1) );
  NOR2X0 U6940_U1 ( .IN1(n5422), .IN2(U6940_n1), .QN(n4519) );
  INVX0 U6941_U2 ( .INP(n103), .ZN(U6941_n1) );
  NOR2X0 U6941_U1 ( .IN1(n5323), .IN2(U6941_n1), .QN(n2594) );
  INVX0 U6944_U2 ( .INP(n3084), .ZN(U6944_n1) );
  NOR2X0 U6944_U1 ( .IN1(n5348), .IN2(U6944_n1), .QN(n3033) );
  INVX0 U6950_U2 ( .INP(n2598), .ZN(U6950_n1) );
  NOR2X0 U6950_U1 ( .IN1(n5365), .IN2(U6950_n1), .QN(n2590) );
  INVX0 U6954_U2 ( .INP(n716), .ZN(U6954_n1) );
  NOR2X0 U6954_U1 ( .IN1(n999), .IN2(U6954_n1), .QN(n3125) );
  INVX0 U6955_U2 ( .INP(n3102), .ZN(U6955_n1) );
  NOR2X0 U6955_U1 ( .IN1(n1013), .IN2(U6955_n1), .QN(n3105) );
  INVX0 U6956_U2 ( .INP(n353), .ZN(U6956_n1) );
  NOR2X0 U6956_U1 ( .IN1(n3146), .IN2(U6956_n1), .QN(n3145) );
  INVX0 U6957_U2 ( .INP(n3160), .ZN(U6957_n1) );
  NOR2X0 U6957_U1 ( .IN1(n3165), .IN2(U6957_n1), .QN(n3164) );
  INVX0 U7174_U2 ( .INP(n2423), .ZN(U7174_n1) );
  NOR2X0 U7174_U1 ( .IN1(n5288), .IN2(U7174_n1), .QN(n2422) );
  INVX0 U7248_U2 ( .INP(n4172), .ZN(U7248_n1) );
  NOR2X0 U7248_U1 ( .IN1(g1536), .IN2(U7248_n1), .QN(n4173) );
  INVX0 U7249_U2 ( .INP(n4190), .ZN(U7249_n1) );
  NOR2X0 U7249_U1 ( .IN1(g1193), .IN2(U7249_n1), .QN(n4191) );
  INVX0 U7402_U2 ( .INP(n4034), .ZN(U7402_n1) );
  NOR2X0 U7402_U1 ( .IN1(n538), .IN2(U7402_n1), .QN(n4037) );
  INVX0 U7405_U2 ( .INP(n4034), .ZN(U7405_n1) );
  NOR2X0 U7405_U1 ( .IN1(n537), .IN2(U7405_n1), .QN(n4039) );
  INVX0 U7413_U2 ( .INP(n3969), .ZN(U7413_n1) );
  NOR2X0 U7413_U1 ( .IN1(n841), .IN2(U7413_n1), .QN(n3972) );
  INVX0 U7416_U2 ( .INP(n3926), .ZN(U7416_n1) );
  NOR2X0 U7416_U1 ( .IN1(n190), .IN2(U7416_n1), .QN(n3929) );
  INVX0 U7427_U2 ( .INP(n3860), .ZN(U7427_n1) );
  NOR2X0 U7427_U1 ( .IN1(n725), .IN2(U7427_n1), .QN(n3863) );
  INVX0 U7438_U2 ( .INP(n4002), .ZN(U7438_n1) );
  NOR2X0 U7438_U1 ( .IN1(n430), .IN2(U7438_n1), .QN(n4003) );
  INVX0 U7449_U2 ( .INP(n4034), .ZN(U7449_n1) );
  NOR2X0 U7449_U1 ( .IN1(n540), .IN2(U7449_n1), .QN(n4032) );
  INVX0 U7455_U2 ( .INP(n4034), .ZN(U7455_n1) );
  NOR2X0 U7455_U1 ( .IN1(n536), .IN2(U7455_n1), .QN(n4035) );
  INVX0 U7464_U2 ( .INP(n3792), .ZN(U7464_n1) );
  NOR2X0 U7464_U1 ( .IN1(n1454), .IN2(U7464_n1), .QN(n3797) );
  INVX0 U7467_U2 ( .INP(n3792), .ZN(U7467_n1) );
  NOR2X0 U7467_U1 ( .IN1(n1460), .IN2(U7467_n1), .QN(n3790) );
  INVX0 U7482_U2 ( .INP(n3792), .ZN(U7482_n1) );
  NOR2X0 U7482_U1 ( .IN1(n1456), .IN2(U7482_n1), .QN(n3795) );
  INVX0 U7492_U2 ( .INP(n3893), .ZN(U7492_n1) );
  NOR2X0 U7492_U1 ( .IN1(n959), .IN2(U7492_n1), .QN(n3891) );
  INVX0 U7513_U2 ( .INP(n3826), .ZN(U7513_n1) );
  NOR2X0 U7513_U1 ( .IN1(n47), .IN2(U7513_n1), .QN(n3827) );
  INVX0 U7516_U2 ( .INP(n3893), .ZN(U7516_n1) );
  NOR2X0 U7516_U1 ( .IN1(n957), .IN2(U7516_n1), .QN(n3896) );
  INVX0 U7549_U2 ( .INP(n4002), .ZN(U7549_n1) );
  NOR2X0 U7549_U1 ( .IN1(n432), .IN2(U7549_n1), .QN(n4007) );
  INVX0 U7561_U2 ( .INP(n3926), .ZN(U7561_n1) );
  NOR2X0 U7561_U1 ( .IN1(n192), .IN2(U7561_n1), .QN(n3931) );
  INVX0 U7574_U2 ( .INP(n3792), .ZN(U7574_n1) );
  NOR2X0 U7574_U1 ( .IN1(n1452), .IN2(U7574_n1), .QN(n3793) );
  INVX0 U7577_U2 ( .INP(n3926), .ZN(U7577_n1) );
  NOR2X0 U7577_U1 ( .IN1(n199), .IN2(U7577_n1), .QN(n3924) );
  INVX0 U7585_U2 ( .INP(n3826), .ZN(U7585_n1) );
  NOR2X0 U7585_U1 ( .IN1(n45), .IN2(U7585_n1), .QN(n3831) );
  INVX0 U7595_U2 ( .INP(n3826), .ZN(U7595_n1) );
  NOR2X0 U7595_U1 ( .IN1(n43), .IN2(U7595_n1), .QN(n3829) );
  INVX0 U7614_U2 ( .INP(n3926), .ZN(U7614_n1) );
  NOR2X0 U7614_U1 ( .IN1(n194), .IN2(U7614_n1), .QN(n3927) );
  INVX0 U7621_U2 ( .INP(n3969), .ZN(U7621_n1) );
  NOR2X0 U7621_U1 ( .IN1(n843), .IN2(U7621_n1), .QN(n3974) );
  INVX0 U7629_U2 ( .INP(n3893), .ZN(U7629_n1) );
  NOR2X0 U7629_U1 ( .IN1(n956), .IN2(U7629_n1), .QN(n3898) );
  INVX0 U7636_U2 ( .INP(n3969), .ZN(U7636_n1) );
  NOR2X0 U7636_U1 ( .IN1(n845), .IN2(U7636_n1), .QN(n3970) );
  INVX0 U7639_U2 ( .INP(n4002), .ZN(U7639_n1) );
  NOR2X0 U7639_U1 ( .IN1(n439), .IN2(U7639_n1), .QN(n4000) );
  INVX0 U7649_U2 ( .INP(n3860), .ZN(U7649_n1) );
  NOR2X0 U7649_U1 ( .IN1(n727), .IN2(U7649_n1), .QN(n3865) );
  INVX0 U7652_U2 ( .INP(n3860), .ZN(U7652_n1) );
  NOR2X0 U7652_U1 ( .IN1(n729), .IN2(U7652_n1), .QN(n3861) );
  INVX0 U7668_U2 ( .INP(n3826), .ZN(U7668_n1) );
  NOR2X0 U7668_U1 ( .IN1(n52), .IN2(U7668_n1), .QN(n3824) );
  INVX0 U7673_U2 ( .INP(n3893), .ZN(U7673_n1) );
  NOR2X0 U7673_U1 ( .IN1(n955), .IN2(U7673_n1), .QN(n3894) );
  INVX0 U7690_U2 ( .INP(n3969), .ZN(U7690_n1) );
  NOR2X0 U7690_U1 ( .IN1(n850), .IN2(U7690_n1), .QN(n3967) );
  INVX0 U7707_U2 ( .INP(n3860), .ZN(U7707_n1) );
  NOR2X0 U7707_U1 ( .IN1(n733), .IN2(U7707_n1), .QN(n3858) );
  INVX0 U7712_U2 ( .INP(n4002), .ZN(U7712_n1) );
  NOR2X0 U7712_U1 ( .IN1(n434), .IN2(U7712_n1), .QN(n4005) );
  INVX0 U7792_U2 ( .INP(g952), .ZN(U7792_n1) );
  NOR2X0 U7792_U1 ( .IN1(n9409), .IN2(U7792_n1), .QN(n2505) );
  INVX0 U7794_U2 ( .INP(g1296), .ZN(U7794_n1) );
  NOR2X0 U7794_U1 ( .IN1(n9409), .IN2(U7794_n1), .QN(n2499) );
  INVX0 U7895_U2 ( .INP(n2668), .ZN(U7895_n1) );
  NOR2X0 U7895_U1 ( .IN1(g113), .IN2(U7895_n1), .QN(n2760) );
  INVX0 U7897_U2 ( .INP(g6), .ZN(U7897_n1) );
  NOR2X0 U7897_U1 ( .IN1(g31), .IN2(U7897_n1), .QN(n3395) );
  INVX0 U7977_U2 ( .INP(g661), .ZN(U7977_n1) );
  NOR2X0 U7977_U1 ( .IN1(n9407), .IN2(U7977_n1), .QN(n4956) );
  INVX0 U8034_U2 ( .INP(n1289), .ZN(U8034_n1) );
  NOR2X0 U8034_U1 ( .IN1(n5612), .IN2(U8034_n1), .QN(n5026) );
  INVX0 U8036_U2 ( .INP(n3729), .ZN(U8036_n1) );
  NOR2X0 U8036_U1 ( .IN1(n5340), .IN2(U8036_n1), .QN(n3941) );
  INVX0 U8050_U2 ( .INP(n183), .ZN(U8050_n1) );
  NOR2X0 U8050_U1 ( .IN1(g1367), .IN2(U8050_n1), .QN(n3733) );
  INVX0 U8055_U2 ( .INP(g1345), .ZN(U8055_n1) );
  NOR2X0 U8055_U1 ( .IN1(n9409), .IN2(U8055_n1), .QN(n4798) );
  INVX0 U8060_U2 ( .INP(g1002), .ZN(U8060_n1) );
  NOR2X0 U8060_U1 ( .IN1(n9407), .IN2(U8060_n1), .QN(n4805) );
  INVX0 U8070_U2 ( .INP(n184), .ZN(U8070_n1) );
  NOR2X0 U8070_U1 ( .IN1(g1361), .IN2(U8070_n1), .QN(n4175) );
  INVX0 U8074_U2 ( .INP(n553), .ZN(U8074_n1) );
  NOR2X0 U8074_U1 ( .IN1(g1018), .IN2(U8074_n1), .QN(n4193) );
  INVX0 U8088_U2 ( .INP(n552), .ZN(U8088_n1) );
  NOR2X0 U8088_U1 ( .IN1(g1024), .IN2(U8088_n1), .QN(n3738) );
  INVX0 U8112_U2 ( .INP(n4525), .ZN(U8112_n1) );
  NOR2X0 U8112_U1 ( .IN1(n4523), .IN2(U8112_n1), .QN(n4524) );
  INVX0 U8113_U2 ( .INP(n4526), .ZN(U8113_n1) );
  NOR2X0 U8113_U1 ( .IN1(n5751), .IN2(U8113_n1), .QN(n4523) );
  INVX0 U8147_U2 ( .INP(g4659), .ZN(U8147_n1) );
  NOR2X0 U8147_U1 ( .IN1(n2573), .IN2(U8147_n1), .QN(n2577) );
  INVX0 U8165_U2 ( .INP(g4849), .ZN(U8165_n1) );
  NOR2X0 U8165_U1 ( .IN1(n2563), .IN2(U8165_n1), .QN(n2567) );
  INVX0 U8185_U2 ( .INP(n869), .ZN(U8185_n1) );
  NOR2X0 U8185_U1 ( .IN1(g1046), .IN2(U8185_n1), .QN(n4938) );
  INVX0 U8192_U2 ( .INP(n176), .ZN(U8192_n1) );
  NOR2X0 U8192_U1 ( .IN1(g1389), .IN2(U8192_n1), .QN(n4913) );
  INVX0 U8210_U2 ( .INP(n4722), .ZN(U8210_n1) );
  NOR2X0 U8210_U1 ( .IN1(n1289), .IN2(U8210_n1), .QN(n4714) );
  INVX0 U8223_U2 ( .INP(n4518), .ZN(U8223_n1) );
  NOR2X0 U8223_U1 ( .IN1(n4516), .IN2(U8223_n1), .QN(n4517) );
  INVX0 U8224_U2 ( .INP(n4519), .ZN(U8224_n1) );
  NOR2X0 U8224_U1 ( .IN1(n5728), .IN2(U8224_n1), .QN(n4516) );
  INVX0 U8281_U2 ( .INP(n4819), .ZN(U8281_n1) );
  NOR2X0 U8281_U1 ( .IN1(n9410), .IN2(U8281_n1), .QN(n5111) );
  INVX0 U8307_U2 ( .INP(g29216), .ZN(U8307_n1) );
  NOR2X0 U8307_U1 ( .IN1(n9408), .IN2(U8307_n1), .QN(g26900) );
  INVX0 U8974_U2 ( .INP(n3362), .ZN(U8974_n1) );
  NOR2X0 U8974_U1 ( .IN1(test_so25), .IN2(U8974_n1), .QN(n2552) );
  INVX0 U8975_U2 ( .INP(n3174), .ZN(U8975_n1) );
  NOR2X0 U8975_U1 ( .IN1(g528), .IN2(U8975_n1), .QN(n3195) );
  INVX0 U9065_U2 ( .INP(g4145), .ZN(U9065_n1) );
  NOR2X0 U9065_U1 ( .IN1(n9408), .IN2(U9065_n1), .QN(n4721) );
  INVX0 U9070_U2 ( .INP(g2841), .ZN(U9070_n1) );
  NOR2X0 U9070_U1 ( .IN1(n9410), .IN2(U9070_n1), .QN(n3730) );
  INVX0 U9075_U2 ( .INP(g19), .ZN(U9075_n1) );
  NOR2X0 U9075_U1 ( .IN1(g9), .IN2(U9075_n1), .QN(n3362) );
  INVX0 U9076_U2 ( .INP(g113), .ZN(U9076_n1) );
  NOR2X0 U9076_U1 ( .IN1(n9407), .IN2(U9076_n1), .QN(g25694) );
  INVX0 U9080_U2 ( .INP(n4305), .ZN(U9080_n1) );
  NOR2X0 U9080_U1 ( .IN1(n9410), .IN2(U9080_n1), .QN(g29277) );
  INVX0 U9084_U2 ( .INP(g4423), .ZN(U9084_n1) );
  NOR2X0 U9084_U1 ( .IN1(n9410), .IN2(U9084_n1), .QN(g26953) );
  INVX0 U9085_U2 ( .INP(g64), .ZN(U9085_n1) );
  NOR2X0 U9085_U1 ( .IN1(n9408), .IN2(U9085_n1), .QN(g24212) );
  INVX0 U9086_U2 ( .INP(n4283), .ZN(U9086_n1) );
  NOR2X0 U9086_U1 ( .IN1(n9407), .IN2(U9086_n1), .QN(g29279) );
  INVX0 U9090_U2 ( .INP(g125), .ZN(U9090_n1) );
  NOR2X0 U9090_U1 ( .IN1(n9410), .IN2(U9090_n1), .QN(g25688) );
  INVX0 U9098_U2 ( .INP(g4681), .ZN(U9098_n1) );
  NOR2X0 U9098_U1 ( .IN1(n2774), .IN2(U9098_n1), .QN(g34028) );
  INVX0 U9099_U2 ( .INP(n2595), .ZN(U9099_n1) );
  NOR2X0 U9099_U1 ( .IN1(n2608), .IN2(U9099_n1), .QN(g34449) );
  INVX0 U9101_U2 ( .INP(g6745), .ZN(U9101_n1) );
  NOR2X0 U9101_U1 ( .IN1(n9406), .IN2(U9101_n1), .QN(g26880) );
  INVX0 U9107_U2 ( .INP(n4448), .ZN(U9107_n1) );
  NOR2X0 U9107_U1 ( .IN1(n8854), .IN2(U9107_n1), .QN(n4447) );
  INVX0 U9111_U2 ( .INP(n4403), .ZN(U9111_n1) );
  NOR2X0 U9111_U1 ( .IN1(n8851), .IN2(U9111_n1), .QN(n4402) );
  INVX0 U9116_U2 ( .INP(n4426), .ZN(U9116_n1) );
  NOR2X0 U9116_U1 ( .IN1(n8858), .IN2(U9116_n1), .QN(n4425) );
  INVX0 U9120_U2 ( .INP(n4437), .ZN(U9120_n1) );
  NOR2X0 U9120_U1 ( .IN1(n8848), .IN2(U9120_n1), .QN(n4436) );
  INVX0 U9124_U2 ( .INP(n4392), .ZN(U9124_n1) );
  NOR2X0 U9124_U1 ( .IN1(n8855), .IN2(U9124_n1), .QN(n4391) );
  INVX0 U9128_U2 ( .INP(n4380), .ZN(U9128_n1) );
  NOR2X0 U9128_U1 ( .IN1(n8849), .IN2(U9128_n1), .QN(n4379) );
  INVX0 U9132_U2 ( .INP(n4415), .ZN(U9132_n1) );
  NOR2X0 U9132_U1 ( .IN1(n8856), .IN2(U9132_n1), .QN(n4414) );
  INVX0 U9136_U2 ( .INP(n4459), .ZN(U9136_n1) );
  NOR2X0 U9136_U1 ( .IN1(n8857), .IN2(U9136_n1), .QN(n4458) );
  INVX0 U9315_U2 ( .INP(n5016), .ZN(U9315_n1) );
  NOR2X0 U9315_U1 ( .IN1(n5753), .IN2(U9315_n1), .QN(n5014) );
  INVX0 U9453_U2 ( .INP(n3065), .ZN(U9453_n1) );
  NOR2X0 U9453_U1 ( .IN1(n8852), .IN2(U9453_n1), .QN(n3064) );
  INVX0 U9825_U2 ( .INP(g112), .ZN(U9825_n1) );
  NOR2X0 U9825_U1 ( .IN1(n1835), .IN2(U9825_n1), .QN(n3115) );
  INVX0 U9886_U2 ( .INP(g370), .ZN(U9886_n1) );
  NOR2X0 U9886_U1 ( .IN1(n1205), .IN2(U9886_n1), .QN(n4948) );
  INVX0 U9927_U2 ( .INP(n3933), .ZN(U9927_n1) );
  NOR2X0 U9927_U1 ( .IN1(g4098), .IN2(U9927_n1), .QN(n3833) );
  INVX0 U9953_U2 ( .INP(g671), .ZN(U9953_n1) );
  NOR2X0 U9953_U1 ( .IN1(n8844), .IN2(U9953_n1), .QN(n4526) );
  INVX0 U9957_U2 ( .INP(g4843), .ZN(U9957_n1) );
  NOR2X0 U9957_U1 ( .IN1(n5283), .IN2(U9957_n1), .QN(n2563) );
  INVX0 U9958_U2 ( .INP(test_so19), .ZN(U9958_n1) );
  NOR2X0 U9958_U1 ( .IN1(n5656), .IN2(U9958_n1), .QN(n2573) );
  INVX0 U9968_U2 ( .INP(n3084), .ZN(U9968_n1) );
  NOR2X0 U9968_U1 ( .IN1(g4358), .IN2(U9968_n1), .QN(n3023) );
  INVX0 U9972_U2 ( .INP(g681), .ZN(U9972_n1) );
  NOR2X0 U9972_U1 ( .IN1(n4535), .IN2(U9972_n1), .QN(n5112) );
  INVX0 U9992_U2 ( .INP(n3675), .ZN(U9992_n1) );
  NOR2X0 U9992_U1 ( .IN1(n488), .IN2(U9992_n1), .QN(n2644) );
  INVX0 U10314_U2 ( .INP(g667), .ZN(U10314_n1) );
  NOR2X0 U10314_U1 ( .IN1(g686), .IN2(U10314_n1), .QN(n4962) );
  INVX0 U10318_U2 ( .INP(g5092), .ZN(U10318_n1) );
  NOR2X0 U10318_U1 ( .IN1(n5681), .IN2(U10318_n1), .QN(n5016) );
endmodule

