module add_mul_mix_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_, 
        c_9_, c_10_, c_11_, c_12_, c_13_, c_14_, c_15_, d_0_, d_1_, d_2_, d_3_, 
        d_4_, d_5_, d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, 
        d_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_, c_9_, c_10_,
         c_11_, c_12_, c_13_, c_14_, c_15_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_,
         d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, d_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958;

  XNOR2_X2 U2019 ( .A(n3826), .B(n3827), .ZN(n2148) );
  XNOR2_X2 U2020 ( .A(n3823), .B(n3824), .ZN(n2423) );
  XNOR2_X2 U2021 ( .A(n2491), .B(n2554), .ZN(n2040) );
  XNOR2_X2 U2022 ( .A(n3815), .B(n3816), .ZN(n3682) );
  XOR2_X2 U2023 ( .A(n2649), .B(n2650), .Z(n2432) );
  XNOR2_X1 U2024 ( .A(n1988), .B(n1989), .ZN(Result_9_) );
  OR2_X1 U2025 ( .A1(n1990), .A2(n1991), .ZN(n1988) );
  AND2_X1 U2026 ( .A1(n1992), .A2(n1993), .ZN(n1990) );
  OR2_X1 U2027 ( .A1(n1994), .A2(n1995), .ZN(n1992) );
  XOR2_X1 U2028 ( .A(n1996), .B(n1997), .Z(Result_8_) );
  XNOR2_X1 U2029 ( .A(n1998), .B(n1999), .ZN(Result_7_) );
  OR2_X1 U2030 ( .A1(n2000), .A2(n2001), .ZN(n1999) );
  AND2_X1 U2031 ( .A1(n2002), .A2(n2003), .ZN(n2000) );
  OR2_X1 U2032 ( .A1(n2004), .A2(n2005), .ZN(n2002) );
  XOR2_X1 U2033 ( .A(n2006), .B(n2007), .Z(Result_6_) );
  XOR2_X1 U2034 ( .A(n2008), .B(n2009), .Z(Result_5_) );
  AND2_X1 U2035 ( .A1(n2010), .A2(n2011), .ZN(n2009) );
  OR2_X1 U2036 ( .A1(n2012), .A2(n2013), .ZN(n2011) );
  AND2_X1 U2037 ( .A1(n2014), .A2(n2015), .ZN(n2013) );
  INV_X1 U2038 ( .A(n2016), .ZN(n2010) );
  XOR2_X1 U2039 ( .A(n2017), .B(n2018), .Z(Result_4_) );
  XOR2_X1 U2040 ( .A(n2019), .B(n2020), .Z(Result_3_) );
  AND2_X1 U2041 ( .A1(n2021), .A2(n2022), .ZN(n2020) );
  OR2_X1 U2042 ( .A1(n2023), .A2(n2024), .ZN(n2022) );
  AND2_X1 U2043 ( .A1(n2025), .A2(n2026), .ZN(n2024) );
  INV_X1 U2044 ( .A(n2027), .ZN(n2021) );
  AND2_X1 U2045 ( .A1(n2028), .A2(n2029), .ZN(Result_31_) );
  OR2_X1 U2046 ( .A1(n2030), .A2(n2031), .ZN(Result_30_) );
  AND2_X1 U2047 ( .A1(n2032), .A2(n2033), .ZN(n2031) );
  OR2_X1 U2048 ( .A1(n2034), .A2(n2035), .ZN(n2033) );
  AND2_X1 U2049 ( .A1(n2029), .A2(n2036), .ZN(n2034) );
  AND2_X1 U2050 ( .A1(n2028), .A2(n2037), .ZN(n2030) );
  OR2_X1 U2051 ( .A1(n2038), .A2(n2039), .ZN(n2037) );
  AND2_X1 U2052 ( .A1(n2040), .A2(n2041), .ZN(n2038) );
  XOR2_X1 U2053 ( .A(n2042), .B(n2043), .Z(Result_2_) );
  XNOR2_X1 U2054 ( .A(n2044), .B(n2045), .ZN(Result_29_) );
  XNOR2_X1 U2055 ( .A(n2046), .B(n2047), .ZN(n2044) );
  XNOR2_X1 U2056 ( .A(n2048), .B(n2049), .ZN(Result_28_) );
  XOR2_X1 U2057 ( .A(n2050), .B(n2051), .Z(n2049) );
  XNOR2_X1 U2058 ( .A(n2052), .B(n2053), .ZN(Result_27_) );
  XOR2_X1 U2059 ( .A(n2054), .B(n2055), .Z(n2053) );
  XNOR2_X1 U2060 ( .A(n2056), .B(n2057), .ZN(Result_26_) );
  XOR2_X1 U2061 ( .A(n2058), .B(n2059), .Z(n2057) );
  XNOR2_X1 U2062 ( .A(n2060), .B(n2061), .ZN(Result_25_) );
  XOR2_X1 U2063 ( .A(n2062), .B(n2063), .Z(n2061) );
  XNOR2_X1 U2064 ( .A(n2064), .B(n2065), .ZN(Result_24_) );
  XOR2_X1 U2065 ( .A(n2066), .B(n2067), .Z(n2065) );
  XNOR2_X1 U2066 ( .A(n2068), .B(n2069), .ZN(Result_23_) );
  XOR2_X1 U2067 ( .A(n2070), .B(n2071), .Z(n2069) );
  XNOR2_X1 U2068 ( .A(n2072), .B(n2073), .ZN(Result_22_) );
  XOR2_X1 U2069 ( .A(n2074), .B(n2075), .Z(n2073) );
  XNOR2_X1 U2070 ( .A(n2076), .B(n2077), .ZN(Result_21_) );
  XOR2_X1 U2071 ( .A(n2078), .B(n2079), .Z(n2077) );
  XNOR2_X1 U2072 ( .A(n2080), .B(n2081), .ZN(Result_20_) );
  XOR2_X1 U2073 ( .A(n2082), .B(n2083), .Z(n2081) );
  XOR2_X1 U2074 ( .A(n2084), .B(n2085), .Z(Result_1_) );
  AND2_X1 U2075 ( .A1(n2086), .A2(n2087), .ZN(n2085) );
  OR2_X1 U2076 ( .A1(n2088), .A2(n2089), .ZN(n2087) );
  AND2_X1 U2077 ( .A1(n2090), .A2(n2091), .ZN(n2088) );
  INV_X1 U2078 ( .A(n2092), .ZN(n2086) );
  XNOR2_X1 U2079 ( .A(n2093), .B(n2094), .ZN(Result_19_) );
  XOR2_X1 U2080 ( .A(n2095), .B(n2096), .Z(n2094) );
  XNOR2_X1 U2081 ( .A(n2097), .B(n2098), .ZN(Result_18_) );
  XOR2_X1 U2082 ( .A(n2099), .B(n2100), .Z(n2098) );
  XNOR2_X1 U2083 ( .A(n2101), .B(n2102), .ZN(Result_17_) );
  XOR2_X1 U2084 ( .A(n2103), .B(n2104), .Z(n2102) );
  XNOR2_X1 U2085 ( .A(n2105), .B(n2106), .ZN(Result_16_) );
  XOR2_X1 U2086 ( .A(n2107), .B(n2108), .Z(n2106) );
  XNOR2_X1 U2087 ( .A(n2109), .B(n2110), .ZN(Result_15_) );
  AND2_X1 U2088 ( .A1(n2111), .A2(n2112), .ZN(Result_14_) );
  INV_X1 U2089 ( .A(n2113), .ZN(n2112) );
  OR2_X1 U2090 ( .A1(n2114), .A2(n2115), .ZN(n2111) );
  AND2_X1 U2091 ( .A1(n2116), .A2(n2110), .ZN(n2114) );
  XOR2_X1 U2092 ( .A(n2117), .B(n2118), .Z(Result_13_) );
  OR2_X1 U2093 ( .A1(n2113), .A2(n2119), .ZN(n2117) );
  XNOR2_X1 U2094 ( .A(n2120), .B(n2121), .ZN(Result_12_) );
  OR2_X1 U2095 ( .A1(n2122), .A2(n2123), .ZN(n2120) );
  AND2_X1 U2096 ( .A1(n2124), .A2(n2125), .ZN(n2122) );
  OR2_X1 U2097 ( .A1(n2126), .A2(n2127), .ZN(n2125) );
  XNOR2_X1 U2098 ( .A(n2128), .B(n2129), .ZN(Result_11_) );
  OR2_X1 U2099 ( .A1(n2130), .A2(n2131), .ZN(n2128) );
  AND2_X1 U2100 ( .A1(n2132), .A2(n2133), .ZN(n2130) );
  OR2_X1 U2101 ( .A1(n2134), .A2(n2135), .ZN(n2133) );
  XNOR2_X1 U2102 ( .A(n2136), .B(n2137), .ZN(Result_10_) );
  OR2_X1 U2103 ( .A1(n2138), .A2(n2139), .ZN(n2136) );
  AND2_X1 U2104 ( .A1(n2140), .A2(n2141), .ZN(n2138) );
  OR2_X1 U2105 ( .A1(n2142), .A2(n2143), .ZN(n2141) );
  OR3_X1 U2106 ( .A1(n2092), .A2(n2144), .A3(n2145), .ZN(Result_0_) );
  INV_X1 U2107 ( .A(n2146), .ZN(n2145) );
  OR2_X1 U2108 ( .A1(n2147), .A2(n2148), .ZN(n2146) );
  AND2_X1 U2109 ( .A1(n2084), .A2(n2089), .ZN(n2144) );
  AND2_X1 U2110 ( .A1(n2042), .A2(n2043), .ZN(n2084) );
  XNOR2_X1 U2111 ( .A(n2091), .B(n2149), .ZN(n2043) );
  OR2_X1 U2112 ( .A1(n2150), .A2(n2151), .ZN(n2042) );
  OR2_X1 U2113 ( .A1(n2152), .A2(n2027), .ZN(n2150) );
  AND3_X1 U2114 ( .A1(n2026), .A2(n2025), .A3(n2023), .ZN(n2027) );
  INV_X1 U2115 ( .A(n2153), .ZN(n2025) );
  AND2_X1 U2116 ( .A1(n2019), .A2(n2023), .ZN(n2152) );
  INV_X1 U2117 ( .A(n2154), .ZN(n2023) );
  OR2_X1 U2118 ( .A1(n2155), .A2(n2151), .ZN(n2154) );
  INV_X1 U2119 ( .A(n2156), .ZN(n2151) );
  OR2_X1 U2120 ( .A1(n2157), .A2(n2158), .ZN(n2156) );
  AND2_X1 U2121 ( .A1(n2157), .A2(n2158), .ZN(n2155) );
  OR2_X1 U2122 ( .A1(n2159), .A2(n2160), .ZN(n2158) );
  AND2_X1 U2123 ( .A1(n2161), .A2(n2162), .ZN(n2160) );
  AND2_X1 U2124 ( .A1(n2163), .A2(n2164), .ZN(n2159) );
  OR2_X1 U2125 ( .A1(n2162), .A2(n2161), .ZN(n2164) );
  XOR2_X1 U2126 ( .A(n2165), .B(n2166), .Z(n2157) );
  XOR2_X1 U2127 ( .A(n2167), .B(n2168), .Z(n2166) );
  AND2_X1 U2128 ( .A1(n2017), .A2(n2018), .ZN(n2019) );
  XNOR2_X1 U2129 ( .A(n2026), .B(n2153), .ZN(n2018) );
  OR2_X1 U2130 ( .A1(n2169), .A2(n2170), .ZN(n2153) );
  AND2_X1 U2131 ( .A1(n2171), .A2(n2172), .ZN(n2170) );
  AND2_X1 U2132 ( .A1(n2173), .A2(n2174), .ZN(n2169) );
  OR2_X1 U2133 ( .A1(n2172), .A2(n2171), .ZN(n2174) );
  XNOR2_X1 U2134 ( .A(n2163), .B(n2175), .ZN(n2026) );
  XOR2_X1 U2135 ( .A(n2162), .B(n2161), .Z(n2175) );
  OR2_X1 U2136 ( .A1(n2176), .A2(n2148), .ZN(n2161) );
  OR2_X1 U2137 ( .A1(n2177), .A2(n2178), .ZN(n2162) );
  AND2_X1 U2138 ( .A1(n2179), .A2(n2180), .ZN(n2178) );
  AND2_X1 U2139 ( .A1(n2181), .A2(n2182), .ZN(n2177) );
  OR2_X1 U2140 ( .A1(n2180), .A2(n2179), .ZN(n2182) );
  XOR2_X1 U2141 ( .A(n2183), .B(n2184), .Z(n2163) );
  XOR2_X1 U2142 ( .A(n2185), .B(n2186), .Z(n2184) );
  OR2_X1 U2143 ( .A1(n2187), .A2(n2188), .ZN(n2017) );
  OR2_X1 U2144 ( .A1(n2189), .A2(n2016), .ZN(n2187) );
  AND3_X1 U2145 ( .A1(n2015), .A2(n2014), .A3(n2012), .ZN(n2016) );
  INV_X1 U2146 ( .A(n2190), .ZN(n2014) );
  AND2_X1 U2147 ( .A1(n2008), .A2(n2012), .ZN(n2189) );
  INV_X1 U2148 ( .A(n2191), .ZN(n2012) );
  OR2_X1 U2149 ( .A1(n2192), .A2(n2188), .ZN(n2191) );
  INV_X1 U2150 ( .A(n2193), .ZN(n2188) );
  OR2_X1 U2151 ( .A1(n2194), .A2(n2195), .ZN(n2193) );
  AND2_X1 U2152 ( .A1(n2194), .A2(n2195), .ZN(n2192) );
  OR2_X1 U2153 ( .A1(n2196), .A2(n2197), .ZN(n2195) );
  AND2_X1 U2154 ( .A1(n2198), .A2(n2199), .ZN(n2197) );
  AND2_X1 U2155 ( .A1(n2200), .A2(n2201), .ZN(n2196) );
  OR2_X1 U2156 ( .A1(n2199), .A2(n2198), .ZN(n2201) );
  XOR2_X1 U2157 ( .A(n2173), .B(n2202), .Z(n2194) );
  XOR2_X1 U2158 ( .A(n2172), .B(n2171), .Z(n2202) );
  OR2_X1 U2159 ( .A1(n2203), .A2(n2148), .ZN(n2171) );
  OR2_X1 U2160 ( .A1(n2204), .A2(n2205), .ZN(n2172) );
  AND2_X1 U2161 ( .A1(n2206), .A2(n2207), .ZN(n2205) );
  AND2_X1 U2162 ( .A1(n2208), .A2(n2209), .ZN(n2204) );
  OR2_X1 U2163 ( .A1(n2207), .A2(n2206), .ZN(n2209) );
  XOR2_X1 U2164 ( .A(n2181), .B(n2210), .Z(n2173) );
  XOR2_X1 U2165 ( .A(n2180), .B(n2179), .Z(n2210) );
  OR2_X1 U2166 ( .A1(n2176), .A2(n2211), .ZN(n2179) );
  OR2_X1 U2167 ( .A1(n2212), .A2(n2213), .ZN(n2180) );
  AND2_X1 U2168 ( .A1(n2214), .A2(n2215), .ZN(n2213) );
  AND2_X1 U2169 ( .A1(n2216), .A2(n2217), .ZN(n2212) );
  OR2_X1 U2170 ( .A1(n2215), .A2(n2214), .ZN(n2217) );
  XOR2_X1 U2171 ( .A(n2218), .B(n2219), .Z(n2181) );
  XOR2_X1 U2172 ( .A(n2220), .B(n2221), .Z(n2219) );
  AND2_X1 U2173 ( .A1(n2006), .A2(n2007), .ZN(n2008) );
  XNOR2_X1 U2174 ( .A(n2015), .B(n2190), .ZN(n2007) );
  OR2_X1 U2175 ( .A1(n2222), .A2(n2223), .ZN(n2190) );
  AND2_X1 U2176 ( .A1(n2224), .A2(n2225), .ZN(n2223) );
  AND2_X1 U2177 ( .A1(n2226), .A2(n2227), .ZN(n2222) );
  OR2_X1 U2178 ( .A1(n2225), .A2(n2224), .ZN(n2227) );
  XNOR2_X1 U2179 ( .A(n2200), .B(n2228), .ZN(n2015) );
  XOR2_X1 U2180 ( .A(n2199), .B(n2198), .Z(n2228) );
  OR2_X1 U2181 ( .A1(n2229), .A2(n2148), .ZN(n2198) );
  OR2_X1 U2182 ( .A1(n2230), .A2(n2231), .ZN(n2199) );
  AND2_X1 U2183 ( .A1(n2232), .A2(n2233), .ZN(n2231) );
  AND2_X1 U2184 ( .A1(n2234), .A2(n2235), .ZN(n2230) );
  OR2_X1 U2185 ( .A1(n2233), .A2(n2232), .ZN(n2235) );
  XOR2_X1 U2186 ( .A(n2208), .B(n2236), .Z(n2200) );
  XOR2_X1 U2187 ( .A(n2207), .B(n2206), .Z(n2236) );
  OR2_X1 U2188 ( .A1(n2203), .A2(n2211), .ZN(n2206) );
  OR2_X1 U2189 ( .A1(n2237), .A2(n2238), .ZN(n2207) );
  AND2_X1 U2190 ( .A1(n2239), .A2(n2240), .ZN(n2238) );
  AND2_X1 U2191 ( .A1(n2241), .A2(n2242), .ZN(n2237) );
  OR2_X1 U2192 ( .A1(n2240), .A2(n2239), .ZN(n2242) );
  XOR2_X1 U2193 ( .A(n2216), .B(n2243), .Z(n2208) );
  XOR2_X1 U2194 ( .A(n2215), .B(n2214), .Z(n2243) );
  OR2_X1 U2195 ( .A1(n2176), .A2(n2244), .ZN(n2214) );
  OR2_X1 U2196 ( .A1(n2245), .A2(n2246), .ZN(n2215) );
  AND2_X1 U2197 ( .A1(n2247), .A2(n2248), .ZN(n2246) );
  AND2_X1 U2198 ( .A1(n2249), .A2(n2250), .ZN(n2245) );
  OR2_X1 U2199 ( .A1(n2248), .A2(n2247), .ZN(n2250) );
  XOR2_X1 U2200 ( .A(n2251), .B(n2252), .Z(n2216) );
  XOR2_X1 U2201 ( .A(n2253), .B(n2254), .Z(n2252) );
  OR2_X1 U2202 ( .A1(n2255), .A2(n2256), .ZN(n2006) );
  OR2_X1 U2203 ( .A1(n2257), .A2(n2001), .ZN(n2255) );
  INV_X1 U2204 ( .A(n2258), .ZN(n2001) );
  OR3_X1 U2205 ( .A1(n2004), .A2(n2005), .A3(n2003), .ZN(n2258) );
  AND2_X1 U2206 ( .A1(n1998), .A2(n2259), .ZN(n2257) );
  INV_X1 U2207 ( .A(n2003), .ZN(n2259) );
  OR2_X1 U2208 ( .A1(n2260), .A2(n2256), .ZN(n2003) );
  INV_X1 U2209 ( .A(n2261), .ZN(n2256) );
  OR2_X1 U2210 ( .A1(n2262), .A2(n2263), .ZN(n2261) );
  AND2_X1 U2211 ( .A1(n2262), .A2(n2263), .ZN(n2260) );
  OR2_X1 U2212 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
  AND2_X1 U2213 ( .A1(n2266), .A2(n2267), .ZN(n2265) );
  AND2_X1 U2214 ( .A1(n2268), .A2(n2269), .ZN(n2264) );
  OR2_X1 U2215 ( .A1(n2267), .A2(n2266), .ZN(n2269) );
  XOR2_X1 U2216 ( .A(n2226), .B(n2270), .Z(n2262) );
  XOR2_X1 U2217 ( .A(n2225), .B(n2224), .Z(n2270) );
  OR2_X1 U2218 ( .A1(n2271), .A2(n2148), .ZN(n2224) );
  OR2_X1 U2219 ( .A1(n2272), .A2(n2273), .ZN(n2225) );
  AND2_X1 U2220 ( .A1(n2274), .A2(n2275), .ZN(n2273) );
  AND2_X1 U2221 ( .A1(n2276), .A2(n2277), .ZN(n2272) );
  OR2_X1 U2222 ( .A1(n2275), .A2(n2274), .ZN(n2277) );
  XOR2_X1 U2223 ( .A(n2234), .B(n2278), .Z(n2226) );
  XOR2_X1 U2224 ( .A(n2233), .B(n2232), .Z(n2278) );
  OR2_X1 U2225 ( .A1(n2229), .A2(n2211), .ZN(n2232) );
  OR2_X1 U2226 ( .A1(n2279), .A2(n2280), .ZN(n2233) );
  AND2_X1 U2227 ( .A1(n2281), .A2(n2282), .ZN(n2280) );
  AND2_X1 U2228 ( .A1(n2283), .A2(n2284), .ZN(n2279) );
  OR2_X1 U2229 ( .A1(n2282), .A2(n2281), .ZN(n2284) );
  XOR2_X1 U2230 ( .A(n2241), .B(n2285), .Z(n2234) );
  XOR2_X1 U2231 ( .A(n2240), .B(n2239), .Z(n2285) );
  OR2_X1 U2232 ( .A1(n2203), .A2(n2244), .ZN(n2239) );
  OR2_X1 U2233 ( .A1(n2286), .A2(n2287), .ZN(n2240) );
  AND2_X1 U2234 ( .A1(n2288), .A2(n2289), .ZN(n2287) );
  AND2_X1 U2235 ( .A1(n2290), .A2(n2291), .ZN(n2286) );
  OR2_X1 U2236 ( .A1(n2289), .A2(n2288), .ZN(n2291) );
  XOR2_X1 U2237 ( .A(n2249), .B(n2292), .Z(n2241) );
  XOR2_X1 U2238 ( .A(n2248), .B(n2247), .Z(n2292) );
  OR2_X1 U2239 ( .A1(n2176), .A2(n2293), .ZN(n2247) );
  OR2_X1 U2240 ( .A1(n2294), .A2(n2295), .ZN(n2248) );
  AND2_X1 U2241 ( .A1(n2296), .A2(n2297), .ZN(n2295) );
  AND2_X1 U2242 ( .A1(n2298), .A2(n2299), .ZN(n2294) );
  OR2_X1 U2243 ( .A1(n2297), .A2(n2296), .ZN(n2299) );
  XOR2_X1 U2244 ( .A(n2300), .B(n2301), .Z(n2249) );
  XOR2_X1 U2245 ( .A(n2302), .B(n2303), .Z(n2301) );
  AND2_X1 U2246 ( .A1(n1996), .A2(n1997), .ZN(n1998) );
  XOR2_X1 U2247 ( .A(n2004), .B(n2005), .Z(n1997) );
  OR2_X1 U2248 ( .A1(n2304), .A2(n2305), .ZN(n2005) );
  AND2_X1 U2249 ( .A1(n2306), .A2(n2307), .ZN(n2305) );
  AND2_X1 U2250 ( .A1(n2308), .A2(n2309), .ZN(n2304) );
  OR2_X1 U2251 ( .A1(n2307), .A2(n2306), .ZN(n2309) );
  XOR2_X1 U2252 ( .A(n2268), .B(n2310), .Z(n2004) );
  XOR2_X1 U2253 ( .A(n2267), .B(n2266), .Z(n2310) );
  OR2_X1 U2254 ( .A1(n2311), .A2(n2148), .ZN(n2266) );
  OR2_X1 U2255 ( .A1(n2312), .A2(n2313), .ZN(n2267) );
  AND2_X1 U2256 ( .A1(n2314), .A2(n2315), .ZN(n2313) );
  AND2_X1 U2257 ( .A1(n2316), .A2(n2317), .ZN(n2312) );
  OR2_X1 U2258 ( .A1(n2315), .A2(n2314), .ZN(n2317) );
  XOR2_X1 U2259 ( .A(n2276), .B(n2318), .Z(n2268) );
  XOR2_X1 U2260 ( .A(n2275), .B(n2274), .Z(n2318) );
  OR2_X1 U2261 ( .A1(n2271), .A2(n2211), .ZN(n2274) );
  OR2_X1 U2262 ( .A1(n2319), .A2(n2320), .ZN(n2275) );
  AND2_X1 U2263 ( .A1(n2321), .A2(n2322), .ZN(n2320) );
  AND2_X1 U2264 ( .A1(n2323), .A2(n2324), .ZN(n2319) );
  OR2_X1 U2265 ( .A1(n2322), .A2(n2321), .ZN(n2324) );
  XOR2_X1 U2266 ( .A(n2283), .B(n2325), .Z(n2276) );
  XOR2_X1 U2267 ( .A(n2282), .B(n2281), .Z(n2325) );
  OR2_X1 U2268 ( .A1(n2229), .A2(n2244), .ZN(n2281) );
  OR2_X1 U2269 ( .A1(n2326), .A2(n2327), .ZN(n2282) );
  AND2_X1 U2270 ( .A1(n2328), .A2(n2329), .ZN(n2327) );
  AND2_X1 U2271 ( .A1(n2330), .A2(n2331), .ZN(n2326) );
  OR2_X1 U2272 ( .A1(n2329), .A2(n2328), .ZN(n2331) );
  XOR2_X1 U2273 ( .A(n2290), .B(n2332), .Z(n2283) );
  XOR2_X1 U2274 ( .A(n2289), .B(n2288), .Z(n2332) );
  OR2_X1 U2275 ( .A1(n2203), .A2(n2293), .ZN(n2288) );
  OR2_X1 U2276 ( .A1(n2333), .A2(n2334), .ZN(n2289) );
  AND2_X1 U2277 ( .A1(n2335), .A2(n2336), .ZN(n2334) );
  AND2_X1 U2278 ( .A1(n2337), .A2(n2338), .ZN(n2333) );
  OR2_X1 U2279 ( .A1(n2336), .A2(n2335), .ZN(n2338) );
  XOR2_X1 U2280 ( .A(n2298), .B(n2339), .Z(n2290) );
  XOR2_X1 U2281 ( .A(n2297), .B(n2296), .Z(n2339) );
  OR2_X1 U2282 ( .A1(n2176), .A2(n2340), .ZN(n2296) );
  OR2_X1 U2283 ( .A1(n2341), .A2(n2342), .ZN(n2297) );
  AND2_X1 U2284 ( .A1(n2343), .A2(n2344), .ZN(n2342) );
  AND2_X1 U2285 ( .A1(n2345), .A2(n2346), .ZN(n2341) );
  OR2_X1 U2286 ( .A1(n2344), .A2(n2343), .ZN(n2346) );
  XOR2_X1 U2287 ( .A(n2347), .B(n2348), .Z(n2298) );
  XOR2_X1 U2288 ( .A(n2349), .B(n2350), .Z(n2348) );
  OR2_X1 U2289 ( .A1(n2351), .A2(n2352), .ZN(n1996) );
  OR2_X1 U2290 ( .A1(n2353), .A2(n1991), .ZN(n2351) );
  INV_X1 U2291 ( .A(n2354), .ZN(n1991) );
  OR3_X1 U2292 ( .A1(n1994), .A2(n1995), .A3(n1993), .ZN(n2354) );
  AND2_X1 U2293 ( .A1(n2355), .A2(n1989), .ZN(n2353) );
  OR2_X1 U2294 ( .A1(n2356), .A2(n2139), .ZN(n1989) );
  INV_X1 U2295 ( .A(n2357), .ZN(n2139) );
  OR3_X1 U2296 ( .A1(n2142), .A2(n2140), .A3(n2143), .ZN(n2357) );
  AND2_X1 U2297 ( .A1(n2358), .A2(n2137), .ZN(n2356) );
  OR2_X1 U2298 ( .A1(n2359), .A2(n2131), .ZN(n2137) );
  INV_X1 U2299 ( .A(n2360), .ZN(n2131) );
  OR3_X1 U2300 ( .A1(n2134), .A2(n2132), .A3(n2135), .ZN(n2360) );
  INV_X1 U2301 ( .A(n2361), .ZN(n2132) );
  AND2_X1 U2302 ( .A1(n2361), .A2(n2129), .ZN(n2359) );
  OR2_X1 U2303 ( .A1(n2362), .A2(n2123), .ZN(n2129) );
  INV_X1 U2304 ( .A(n2363), .ZN(n2123) );
  OR3_X1 U2305 ( .A1(n2126), .A2(n2124), .A3(n2127), .ZN(n2363) );
  INV_X1 U2306 ( .A(n2364), .ZN(n2124) );
  AND2_X1 U2307 ( .A1(n2364), .A2(n2121), .ZN(n2362) );
  OR2_X1 U2308 ( .A1(n2365), .A2(n2366), .ZN(n2121) );
  AND2_X1 U2309 ( .A1(n2119), .A2(n2118), .ZN(n2366) );
  INV_X1 U2310 ( .A(n2367), .ZN(n2119) );
  OR2_X1 U2311 ( .A1(n2368), .A2(n2369), .ZN(n2367) );
  AND2_X1 U2312 ( .A1(n2113), .A2(n2118), .ZN(n2365) );
  XOR2_X1 U2313 ( .A(n2126), .B(n2127), .Z(n2118) );
  OR2_X1 U2314 ( .A1(n2370), .A2(n2371), .ZN(n2127) );
  AND2_X1 U2315 ( .A1(n2372), .A2(n2373), .ZN(n2371) );
  AND2_X1 U2316 ( .A1(n2374), .A2(n2375), .ZN(n2370) );
  OR2_X1 U2317 ( .A1(n2373), .A2(n2372), .ZN(n2375) );
  XOR2_X1 U2318 ( .A(n2376), .B(n2377), .Z(n2126) );
  XOR2_X1 U2319 ( .A(n2378), .B(n2379), .Z(n2377) );
  AND3_X1 U2320 ( .A1(n2110), .A2(n2115), .A3(n2116), .ZN(n2113) );
  INV_X1 U2321 ( .A(n2109), .ZN(n2116) );
  OR2_X1 U2322 ( .A1(n2380), .A2(n2381), .ZN(n2109) );
  AND2_X1 U2323 ( .A1(n2108), .A2(n2107), .ZN(n2381) );
  AND2_X1 U2324 ( .A1(n2105), .A2(n2382), .ZN(n2380) );
  OR2_X1 U2325 ( .A1(n2108), .A2(n2107), .ZN(n2382) );
  OR2_X1 U2326 ( .A1(n2383), .A2(n2384), .ZN(n2107) );
  AND2_X1 U2327 ( .A1(n2104), .A2(n2103), .ZN(n2384) );
  AND2_X1 U2328 ( .A1(n2101), .A2(n2385), .ZN(n2383) );
  OR2_X1 U2329 ( .A1(n2104), .A2(n2103), .ZN(n2385) );
  OR2_X1 U2330 ( .A1(n2386), .A2(n2387), .ZN(n2103) );
  AND2_X1 U2331 ( .A1(n2100), .A2(n2099), .ZN(n2387) );
  AND2_X1 U2332 ( .A1(n2097), .A2(n2388), .ZN(n2386) );
  OR2_X1 U2333 ( .A1(n2100), .A2(n2099), .ZN(n2388) );
  OR2_X1 U2334 ( .A1(n2389), .A2(n2390), .ZN(n2099) );
  AND2_X1 U2335 ( .A1(n2096), .A2(n2095), .ZN(n2390) );
  AND2_X1 U2336 ( .A1(n2093), .A2(n2391), .ZN(n2389) );
  OR2_X1 U2337 ( .A1(n2096), .A2(n2095), .ZN(n2391) );
  OR2_X1 U2338 ( .A1(n2392), .A2(n2393), .ZN(n2095) );
  AND2_X1 U2339 ( .A1(n2083), .A2(n2082), .ZN(n2393) );
  AND2_X1 U2340 ( .A1(n2080), .A2(n2394), .ZN(n2392) );
  OR2_X1 U2341 ( .A1(n2083), .A2(n2082), .ZN(n2394) );
  OR2_X1 U2342 ( .A1(n2395), .A2(n2396), .ZN(n2082) );
  AND2_X1 U2343 ( .A1(n2079), .A2(n2078), .ZN(n2396) );
  AND2_X1 U2344 ( .A1(n2076), .A2(n2397), .ZN(n2395) );
  OR2_X1 U2345 ( .A1(n2079), .A2(n2078), .ZN(n2397) );
  OR2_X1 U2346 ( .A1(n2398), .A2(n2399), .ZN(n2078) );
  AND2_X1 U2347 ( .A1(n2075), .A2(n2074), .ZN(n2399) );
  AND2_X1 U2348 ( .A1(n2072), .A2(n2400), .ZN(n2398) );
  OR2_X1 U2349 ( .A1(n2075), .A2(n2074), .ZN(n2400) );
  OR2_X1 U2350 ( .A1(n2401), .A2(n2402), .ZN(n2074) );
  AND2_X1 U2351 ( .A1(n2071), .A2(n2070), .ZN(n2402) );
  AND2_X1 U2352 ( .A1(n2068), .A2(n2403), .ZN(n2401) );
  OR2_X1 U2353 ( .A1(n2071), .A2(n2070), .ZN(n2403) );
  OR2_X1 U2354 ( .A1(n2404), .A2(n2405), .ZN(n2070) );
  AND2_X1 U2355 ( .A1(n2067), .A2(n2066), .ZN(n2405) );
  AND2_X1 U2356 ( .A1(n2064), .A2(n2406), .ZN(n2404) );
  OR2_X1 U2357 ( .A1(n2067), .A2(n2066), .ZN(n2406) );
  OR2_X1 U2358 ( .A1(n2407), .A2(n2408), .ZN(n2066) );
  AND2_X1 U2359 ( .A1(n2063), .A2(n2062), .ZN(n2408) );
  AND2_X1 U2360 ( .A1(n2060), .A2(n2409), .ZN(n2407) );
  OR2_X1 U2361 ( .A1(n2063), .A2(n2062), .ZN(n2409) );
  OR2_X1 U2362 ( .A1(n2410), .A2(n2411), .ZN(n2062) );
  AND2_X1 U2363 ( .A1(n2059), .A2(n2058), .ZN(n2411) );
  AND2_X1 U2364 ( .A1(n2056), .A2(n2412), .ZN(n2410) );
  OR2_X1 U2365 ( .A1(n2059), .A2(n2058), .ZN(n2412) );
  OR2_X1 U2366 ( .A1(n2413), .A2(n2414), .ZN(n2058) );
  AND2_X1 U2367 ( .A1(n2055), .A2(n2054), .ZN(n2414) );
  AND2_X1 U2368 ( .A1(n2052), .A2(n2415), .ZN(n2413) );
  OR2_X1 U2369 ( .A1(n2055), .A2(n2054), .ZN(n2415) );
  OR2_X1 U2370 ( .A1(n2416), .A2(n2417), .ZN(n2054) );
  AND2_X1 U2371 ( .A1(n2051), .A2(n2050), .ZN(n2417) );
  AND2_X1 U2372 ( .A1(n2048), .A2(n2418), .ZN(n2416) );
  OR2_X1 U2373 ( .A1(n2051), .A2(n2050), .ZN(n2418) );
  OR2_X1 U2374 ( .A1(n2419), .A2(n2420), .ZN(n2050) );
  AND2_X1 U2375 ( .A1(n2045), .A2(n2047), .ZN(n2420) );
  AND2_X1 U2376 ( .A1(n2421), .A2(n2422), .ZN(n2419) );
  OR2_X1 U2377 ( .A1(n2045), .A2(n2047), .ZN(n2422) );
  OR2_X1 U2378 ( .A1(n2423), .A2(n2036), .ZN(n2047) );
  OR3_X1 U2379 ( .A1(n2040), .A2(n2036), .A3(n2424), .ZN(n2045) );
  INV_X1 U2380 ( .A(n2046), .ZN(n2421) );
  OR2_X1 U2381 ( .A1(n2425), .A2(n2426), .ZN(n2046) );
  AND2_X1 U2382 ( .A1(n2427), .A2(n2428), .ZN(n2426) );
  OR2_X1 U2383 ( .A1(n2429), .A2(n2035), .ZN(n2428) );
  AND2_X1 U2384 ( .A1(n2029), .A2(n2040), .ZN(n2429) );
  AND2_X1 U2385 ( .A1(n2032), .A2(n2430), .ZN(n2425) );
  OR2_X1 U2386 ( .A1(n2431), .A2(n2039), .ZN(n2430) );
  AND2_X1 U2387 ( .A1(n2432), .A2(n2041), .ZN(n2431) );
  INV_X1 U2388 ( .A(n2040), .ZN(n2032) );
  OR2_X1 U2389 ( .A1(n2433), .A2(n2036), .ZN(n2051) );
  XOR2_X1 U2390 ( .A(n2434), .B(n2435), .Z(n2048) );
  XNOR2_X1 U2391 ( .A(n2436), .B(n2437), .ZN(n2434) );
  OR2_X1 U2392 ( .A1(n2438), .A2(n2036), .ZN(n2055) );
  XOR2_X1 U2393 ( .A(n2439), .B(n2440), .Z(n2052) );
  XOR2_X1 U2394 ( .A(n2441), .B(n2442), .Z(n2440) );
  OR2_X1 U2395 ( .A1(n2443), .A2(n2036), .ZN(n2059) );
  XOR2_X1 U2396 ( .A(n2444), .B(n2445), .Z(n2056) );
  XOR2_X1 U2397 ( .A(n2446), .B(n2447), .Z(n2445) );
  OR2_X1 U2398 ( .A1(n2448), .A2(n2036), .ZN(n2063) );
  XOR2_X1 U2399 ( .A(n2449), .B(n2450), .Z(n2060) );
  XOR2_X1 U2400 ( .A(n2451), .B(n2452), .Z(n2450) );
  OR2_X1 U2401 ( .A1(n2453), .A2(n2036), .ZN(n2067) );
  XOR2_X1 U2402 ( .A(n2454), .B(n2455), .Z(n2064) );
  XOR2_X1 U2403 ( .A(n2456), .B(n2457), .Z(n2455) );
  OR2_X1 U2404 ( .A1(n2458), .A2(n2036), .ZN(n2071) );
  XOR2_X1 U2405 ( .A(n2459), .B(n2460), .Z(n2068) );
  XOR2_X1 U2406 ( .A(n2461), .B(n2462), .Z(n2460) );
  OR2_X1 U2407 ( .A1(n2463), .A2(n2036), .ZN(n2075) );
  XOR2_X1 U2408 ( .A(n2464), .B(n2465), .Z(n2072) );
  XOR2_X1 U2409 ( .A(n2466), .B(n2467), .Z(n2465) );
  OR2_X1 U2410 ( .A1(n2468), .A2(n2036), .ZN(n2079) );
  XOR2_X1 U2411 ( .A(n2469), .B(n2470), .Z(n2076) );
  XOR2_X1 U2412 ( .A(n2471), .B(n2472), .Z(n2470) );
  OR2_X1 U2413 ( .A1(n2340), .A2(n2036), .ZN(n2083) );
  XOR2_X1 U2414 ( .A(n2473), .B(n2474), .Z(n2080) );
  XOR2_X1 U2415 ( .A(n2475), .B(n2476), .Z(n2474) );
  OR2_X1 U2416 ( .A1(n2293), .A2(n2036), .ZN(n2096) );
  XOR2_X1 U2417 ( .A(n2477), .B(n2478), .Z(n2093) );
  XOR2_X1 U2418 ( .A(n2479), .B(n2480), .Z(n2478) );
  OR2_X1 U2419 ( .A1(n2244), .A2(n2036), .ZN(n2100) );
  XOR2_X1 U2420 ( .A(n2481), .B(n2482), .Z(n2097) );
  XOR2_X1 U2421 ( .A(n2483), .B(n2484), .Z(n2482) );
  OR2_X1 U2422 ( .A1(n2211), .A2(n2036), .ZN(n2104) );
  XOR2_X1 U2423 ( .A(n2485), .B(n2486), .Z(n2101) );
  XOR2_X1 U2424 ( .A(n2487), .B(n2488), .Z(n2486) );
  OR2_X1 U2425 ( .A1(n2036), .A2(n2148), .ZN(n2108) );
  INV_X1 U2426 ( .A(n2028), .ZN(n2036) );
  AND2_X1 U2427 ( .A1(n2489), .A2(n2490), .ZN(n2028) );
  INV_X1 U2428 ( .A(n2491), .ZN(n2490) );
  OR2_X1 U2429 ( .A1(c_15_), .A2(d_15_), .ZN(n2489) );
  XOR2_X1 U2430 ( .A(n2492), .B(n2493), .Z(n2105) );
  XOR2_X1 U2431 ( .A(n2494), .B(n2495), .Z(n2493) );
  XOR2_X1 U2432 ( .A(n2368), .B(n2369), .Z(n2115) );
  OR2_X1 U2433 ( .A1(n2496), .A2(n2497), .ZN(n2369) );
  AND2_X1 U2434 ( .A1(n2498), .A2(n2499), .ZN(n2497) );
  AND2_X1 U2435 ( .A1(n2500), .A2(n2501), .ZN(n2496) );
  OR2_X1 U2436 ( .A1(n2498), .A2(n2499), .ZN(n2501) );
  XOR2_X1 U2437 ( .A(n2374), .B(n2502), .Z(n2368) );
  XOR2_X1 U2438 ( .A(n2373), .B(n2372), .Z(n2502) );
  OR2_X1 U2439 ( .A1(n2432), .A2(n2148), .ZN(n2372) );
  OR2_X1 U2440 ( .A1(n2503), .A2(n2504), .ZN(n2373) );
  AND2_X1 U2441 ( .A1(n2505), .A2(n2506), .ZN(n2504) );
  AND2_X1 U2442 ( .A1(n2507), .A2(n2508), .ZN(n2503) );
  OR2_X1 U2443 ( .A1(n2506), .A2(n2505), .ZN(n2508) );
  XOR2_X1 U2444 ( .A(n2509), .B(n2510), .Z(n2374) );
  XOR2_X1 U2445 ( .A(n2511), .B(n2512), .Z(n2510) );
  XNOR2_X1 U2446 ( .A(n2500), .B(n2513), .ZN(n2110) );
  XOR2_X1 U2447 ( .A(n2499), .B(n2498), .Z(n2513) );
  OR2_X1 U2448 ( .A1(n2040), .A2(n2148), .ZN(n2498) );
  OR2_X1 U2449 ( .A1(n2514), .A2(n2515), .ZN(n2499) );
  AND2_X1 U2450 ( .A1(n2495), .A2(n2494), .ZN(n2515) );
  AND2_X1 U2451 ( .A1(n2492), .A2(n2516), .ZN(n2514) );
  OR2_X1 U2452 ( .A1(n2494), .A2(n2495), .ZN(n2516) );
  OR2_X1 U2453 ( .A1(n2211), .A2(n2040), .ZN(n2495) );
  OR2_X1 U2454 ( .A1(n2517), .A2(n2518), .ZN(n2494) );
  AND2_X1 U2455 ( .A1(n2488), .A2(n2487), .ZN(n2518) );
  AND2_X1 U2456 ( .A1(n2485), .A2(n2519), .ZN(n2517) );
  OR2_X1 U2457 ( .A1(n2487), .A2(n2488), .ZN(n2519) );
  OR2_X1 U2458 ( .A1(n2244), .A2(n2040), .ZN(n2488) );
  OR2_X1 U2459 ( .A1(n2520), .A2(n2521), .ZN(n2487) );
  AND2_X1 U2460 ( .A1(n2484), .A2(n2483), .ZN(n2521) );
  AND2_X1 U2461 ( .A1(n2481), .A2(n2522), .ZN(n2520) );
  OR2_X1 U2462 ( .A1(n2483), .A2(n2484), .ZN(n2522) );
  OR2_X1 U2463 ( .A1(n2293), .A2(n2040), .ZN(n2484) );
  OR2_X1 U2464 ( .A1(n2523), .A2(n2524), .ZN(n2483) );
  AND2_X1 U2465 ( .A1(n2480), .A2(n2479), .ZN(n2524) );
  AND2_X1 U2466 ( .A1(n2477), .A2(n2525), .ZN(n2523) );
  OR2_X1 U2467 ( .A1(n2479), .A2(n2480), .ZN(n2525) );
  OR2_X1 U2468 ( .A1(n2340), .A2(n2040), .ZN(n2480) );
  OR2_X1 U2469 ( .A1(n2526), .A2(n2527), .ZN(n2479) );
  AND2_X1 U2470 ( .A1(n2476), .A2(n2475), .ZN(n2527) );
  AND2_X1 U2471 ( .A1(n2473), .A2(n2528), .ZN(n2526) );
  OR2_X1 U2472 ( .A1(n2475), .A2(n2476), .ZN(n2528) );
  OR2_X1 U2473 ( .A1(n2468), .A2(n2040), .ZN(n2476) );
  OR2_X1 U2474 ( .A1(n2529), .A2(n2530), .ZN(n2475) );
  AND2_X1 U2475 ( .A1(n2472), .A2(n2471), .ZN(n2530) );
  AND2_X1 U2476 ( .A1(n2469), .A2(n2531), .ZN(n2529) );
  OR2_X1 U2477 ( .A1(n2471), .A2(n2472), .ZN(n2531) );
  OR2_X1 U2478 ( .A1(n2463), .A2(n2040), .ZN(n2472) );
  OR2_X1 U2479 ( .A1(n2532), .A2(n2533), .ZN(n2471) );
  AND2_X1 U2480 ( .A1(n2467), .A2(n2466), .ZN(n2533) );
  AND2_X1 U2481 ( .A1(n2464), .A2(n2534), .ZN(n2532) );
  OR2_X1 U2482 ( .A1(n2466), .A2(n2467), .ZN(n2534) );
  OR2_X1 U2483 ( .A1(n2458), .A2(n2040), .ZN(n2467) );
  OR2_X1 U2484 ( .A1(n2535), .A2(n2536), .ZN(n2466) );
  AND2_X1 U2485 ( .A1(n2462), .A2(n2461), .ZN(n2536) );
  AND2_X1 U2486 ( .A1(n2459), .A2(n2537), .ZN(n2535) );
  OR2_X1 U2487 ( .A1(n2461), .A2(n2462), .ZN(n2537) );
  OR2_X1 U2488 ( .A1(n2453), .A2(n2040), .ZN(n2462) );
  OR2_X1 U2489 ( .A1(n2538), .A2(n2539), .ZN(n2461) );
  AND2_X1 U2490 ( .A1(n2457), .A2(n2456), .ZN(n2539) );
  AND2_X1 U2491 ( .A1(n2454), .A2(n2540), .ZN(n2538) );
  OR2_X1 U2492 ( .A1(n2456), .A2(n2457), .ZN(n2540) );
  OR2_X1 U2493 ( .A1(n2448), .A2(n2040), .ZN(n2457) );
  OR2_X1 U2494 ( .A1(n2541), .A2(n2542), .ZN(n2456) );
  AND2_X1 U2495 ( .A1(n2452), .A2(n2451), .ZN(n2542) );
  AND2_X1 U2496 ( .A1(n2449), .A2(n2543), .ZN(n2541) );
  OR2_X1 U2497 ( .A1(n2451), .A2(n2452), .ZN(n2543) );
  OR2_X1 U2498 ( .A1(n2443), .A2(n2040), .ZN(n2452) );
  OR2_X1 U2499 ( .A1(n2544), .A2(n2545), .ZN(n2451) );
  AND2_X1 U2500 ( .A1(n2447), .A2(n2446), .ZN(n2545) );
  AND2_X1 U2501 ( .A1(n2444), .A2(n2546), .ZN(n2544) );
  OR2_X1 U2502 ( .A1(n2446), .A2(n2447), .ZN(n2546) );
  OR2_X1 U2503 ( .A1(n2438), .A2(n2040), .ZN(n2447) );
  OR2_X1 U2504 ( .A1(n2547), .A2(n2548), .ZN(n2446) );
  AND2_X1 U2505 ( .A1(n2442), .A2(n2441), .ZN(n2548) );
  AND2_X1 U2506 ( .A1(n2439), .A2(n2549), .ZN(n2547) );
  OR2_X1 U2507 ( .A1(n2441), .A2(n2442), .ZN(n2549) );
  OR2_X1 U2508 ( .A1(n2433), .A2(n2040), .ZN(n2442) );
  OR2_X1 U2509 ( .A1(n2550), .A2(n2551), .ZN(n2441) );
  AND2_X1 U2510 ( .A1(n2435), .A2(n2437), .ZN(n2551) );
  AND2_X1 U2511 ( .A1(n2552), .A2(n2553), .ZN(n2550) );
  OR2_X1 U2512 ( .A1(n2437), .A2(n2435), .ZN(n2553) );
  OR2_X1 U2513 ( .A1(n2040), .A2(n2423), .ZN(n2435) );
  OR3_X1 U2514 ( .A1(n2040), .A2(n2432), .A3(n2424), .ZN(n2437) );
  XOR2_X1 U2515 ( .A(d_14_), .B(c_14_), .Z(n2554) );
  INV_X1 U2516 ( .A(n2436), .ZN(n2552) );
  OR2_X1 U2517 ( .A1(n2555), .A2(n2556), .ZN(n2436) );
  AND2_X1 U2518 ( .A1(n2557), .A2(n2558), .ZN(n2556) );
  OR2_X1 U2519 ( .A1(n2559), .A2(n2035), .ZN(n2558) );
  AND2_X1 U2520 ( .A1(n2029), .A2(n2432), .ZN(n2559) );
  AND2_X1 U2521 ( .A1(n2427), .A2(n2560), .ZN(n2555) );
  OR2_X1 U2522 ( .A1(n2561), .A2(n2039), .ZN(n2560) );
  AND2_X1 U2523 ( .A1(n2562), .A2(n2041), .ZN(n2561) );
  INV_X1 U2524 ( .A(n2432), .ZN(n2427) );
  XOR2_X1 U2525 ( .A(n2563), .B(n2564), .Z(n2439) );
  XNOR2_X1 U2526 ( .A(n2565), .B(n2566), .ZN(n2563) );
  XOR2_X1 U2527 ( .A(n2567), .B(n2568), .Z(n2444) );
  XOR2_X1 U2528 ( .A(n2569), .B(n2570), .Z(n2568) );
  XOR2_X1 U2529 ( .A(n2571), .B(n2572), .Z(n2449) );
  XOR2_X1 U2530 ( .A(n2573), .B(n2574), .Z(n2572) );
  XOR2_X1 U2531 ( .A(n2575), .B(n2576), .Z(n2454) );
  XOR2_X1 U2532 ( .A(n2577), .B(n2578), .Z(n2576) );
  XOR2_X1 U2533 ( .A(n2579), .B(n2580), .Z(n2459) );
  XOR2_X1 U2534 ( .A(n2581), .B(n2582), .Z(n2580) );
  XOR2_X1 U2535 ( .A(n2583), .B(n2584), .Z(n2464) );
  XOR2_X1 U2536 ( .A(n2585), .B(n2586), .Z(n2584) );
  XOR2_X1 U2537 ( .A(n2587), .B(n2588), .Z(n2469) );
  XOR2_X1 U2538 ( .A(n2589), .B(n2590), .Z(n2588) );
  XOR2_X1 U2539 ( .A(n2591), .B(n2592), .Z(n2473) );
  XOR2_X1 U2540 ( .A(n2593), .B(n2594), .Z(n2592) );
  XOR2_X1 U2541 ( .A(n2595), .B(n2596), .Z(n2477) );
  XOR2_X1 U2542 ( .A(n2597), .B(n2598), .Z(n2596) );
  XOR2_X1 U2543 ( .A(n2599), .B(n2600), .Z(n2481) );
  XOR2_X1 U2544 ( .A(n2601), .B(n2602), .Z(n2600) );
  XOR2_X1 U2545 ( .A(n2603), .B(n2604), .Z(n2485) );
  XOR2_X1 U2546 ( .A(n2605), .B(n2606), .Z(n2604) );
  XOR2_X1 U2547 ( .A(n2607), .B(n2608), .Z(n2492) );
  XOR2_X1 U2548 ( .A(n2609), .B(n2610), .Z(n2608) );
  XOR2_X1 U2549 ( .A(n2507), .B(n2611), .Z(n2500) );
  XOR2_X1 U2550 ( .A(n2506), .B(n2505), .Z(n2611) );
  OR2_X1 U2551 ( .A1(n2211), .A2(n2432), .ZN(n2505) );
  OR2_X1 U2552 ( .A1(n2612), .A2(n2613), .ZN(n2506) );
  AND2_X1 U2553 ( .A1(n2610), .A2(n2609), .ZN(n2613) );
  AND2_X1 U2554 ( .A1(n2607), .A2(n2614), .ZN(n2612) );
  OR2_X1 U2555 ( .A1(n2609), .A2(n2610), .ZN(n2614) );
  OR2_X1 U2556 ( .A1(n2244), .A2(n2432), .ZN(n2610) );
  OR2_X1 U2557 ( .A1(n2615), .A2(n2616), .ZN(n2609) );
  AND2_X1 U2558 ( .A1(n2606), .A2(n2605), .ZN(n2616) );
  AND2_X1 U2559 ( .A1(n2603), .A2(n2617), .ZN(n2615) );
  OR2_X1 U2560 ( .A1(n2605), .A2(n2606), .ZN(n2617) );
  OR2_X1 U2561 ( .A1(n2293), .A2(n2432), .ZN(n2606) );
  OR2_X1 U2562 ( .A1(n2618), .A2(n2619), .ZN(n2605) );
  AND2_X1 U2563 ( .A1(n2602), .A2(n2601), .ZN(n2619) );
  AND2_X1 U2564 ( .A1(n2599), .A2(n2620), .ZN(n2618) );
  OR2_X1 U2565 ( .A1(n2601), .A2(n2602), .ZN(n2620) );
  OR2_X1 U2566 ( .A1(n2340), .A2(n2432), .ZN(n2602) );
  OR2_X1 U2567 ( .A1(n2621), .A2(n2622), .ZN(n2601) );
  AND2_X1 U2568 ( .A1(n2598), .A2(n2597), .ZN(n2622) );
  AND2_X1 U2569 ( .A1(n2595), .A2(n2623), .ZN(n2621) );
  OR2_X1 U2570 ( .A1(n2597), .A2(n2598), .ZN(n2623) );
  OR2_X1 U2571 ( .A1(n2468), .A2(n2432), .ZN(n2598) );
  OR2_X1 U2572 ( .A1(n2624), .A2(n2625), .ZN(n2597) );
  AND2_X1 U2573 ( .A1(n2594), .A2(n2593), .ZN(n2625) );
  AND2_X1 U2574 ( .A1(n2591), .A2(n2626), .ZN(n2624) );
  OR2_X1 U2575 ( .A1(n2593), .A2(n2594), .ZN(n2626) );
  OR2_X1 U2576 ( .A1(n2463), .A2(n2432), .ZN(n2594) );
  OR2_X1 U2577 ( .A1(n2627), .A2(n2628), .ZN(n2593) );
  AND2_X1 U2578 ( .A1(n2590), .A2(n2589), .ZN(n2628) );
  AND2_X1 U2579 ( .A1(n2587), .A2(n2629), .ZN(n2627) );
  OR2_X1 U2580 ( .A1(n2589), .A2(n2590), .ZN(n2629) );
  OR2_X1 U2581 ( .A1(n2458), .A2(n2432), .ZN(n2590) );
  OR2_X1 U2582 ( .A1(n2630), .A2(n2631), .ZN(n2589) );
  AND2_X1 U2583 ( .A1(n2586), .A2(n2585), .ZN(n2631) );
  AND2_X1 U2584 ( .A1(n2583), .A2(n2632), .ZN(n2630) );
  OR2_X1 U2585 ( .A1(n2585), .A2(n2586), .ZN(n2632) );
  OR2_X1 U2586 ( .A1(n2453), .A2(n2432), .ZN(n2586) );
  OR2_X1 U2587 ( .A1(n2633), .A2(n2634), .ZN(n2585) );
  AND2_X1 U2588 ( .A1(n2582), .A2(n2581), .ZN(n2634) );
  AND2_X1 U2589 ( .A1(n2579), .A2(n2635), .ZN(n2633) );
  OR2_X1 U2590 ( .A1(n2581), .A2(n2582), .ZN(n2635) );
  OR2_X1 U2591 ( .A1(n2448), .A2(n2432), .ZN(n2582) );
  OR2_X1 U2592 ( .A1(n2636), .A2(n2637), .ZN(n2581) );
  AND2_X1 U2593 ( .A1(n2578), .A2(n2577), .ZN(n2637) );
  AND2_X1 U2594 ( .A1(n2575), .A2(n2638), .ZN(n2636) );
  OR2_X1 U2595 ( .A1(n2577), .A2(n2578), .ZN(n2638) );
  OR2_X1 U2596 ( .A1(n2443), .A2(n2432), .ZN(n2578) );
  OR2_X1 U2597 ( .A1(n2639), .A2(n2640), .ZN(n2577) );
  AND2_X1 U2598 ( .A1(n2574), .A2(n2573), .ZN(n2640) );
  AND2_X1 U2599 ( .A1(n2571), .A2(n2641), .ZN(n2639) );
  OR2_X1 U2600 ( .A1(n2573), .A2(n2574), .ZN(n2641) );
  OR2_X1 U2601 ( .A1(n2438), .A2(n2432), .ZN(n2574) );
  OR2_X1 U2602 ( .A1(n2642), .A2(n2643), .ZN(n2573) );
  AND2_X1 U2603 ( .A1(n2570), .A2(n2569), .ZN(n2643) );
  AND2_X1 U2604 ( .A1(n2567), .A2(n2644), .ZN(n2642) );
  OR2_X1 U2605 ( .A1(n2569), .A2(n2570), .ZN(n2644) );
  OR2_X1 U2606 ( .A1(n2433), .A2(n2432), .ZN(n2570) );
  OR2_X1 U2607 ( .A1(n2645), .A2(n2646), .ZN(n2569) );
  AND2_X1 U2608 ( .A1(n2564), .A2(n2566), .ZN(n2646) );
  AND2_X1 U2609 ( .A1(n2647), .A2(n2648), .ZN(n2645) );
  OR2_X1 U2610 ( .A1(n2566), .A2(n2564), .ZN(n2648) );
  OR2_X1 U2611 ( .A1(n2432), .A2(n2423), .ZN(n2564) );
  OR3_X1 U2612 ( .A1(n2562), .A2(n2432), .A3(n2424), .ZN(n2566) );
  XNOR2_X1 U2613 ( .A(n2651), .B(c_13_), .ZN(n2650) );
  INV_X1 U2614 ( .A(n2565), .ZN(n2647) );
  OR2_X1 U2615 ( .A1(n2652), .A2(n2653), .ZN(n2565) );
  AND2_X1 U2616 ( .A1(n2654), .A2(n2655), .ZN(n2653) );
  OR2_X1 U2617 ( .A1(n2656), .A2(n2035), .ZN(n2655) );
  AND2_X1 U2618 ( .A1(n2562), .A2(n2029), .ZN(n2656) );
  AND2_X1 U2619 ( .A1(n2557), .A2(n2657), .ZN(n2652) );
  OR2_X1 U2620 ( .A1(n2658), .A2(n2039), .ZN(n2657) );
  AND2_X1 U2621 ( .A1(n2659), .A2(n2041), .ZN(n2658) );
  XOR2_X1 U2622 ( .A(n2660), .B(n2661), .Z(n2567) );
  XNOR2_X1 U2623 ( .A(n2662), .B(n2663), .ZN(n2660) );
  XOR2_X1 U2624 ( .A(n2664), .B(n2665), .Z(n2571) );
  XOR2_X1 U2625 ( .A(n2666), .B(n2667), .Z(n2665) );
  XOR2_X1 U2626 ( .A(n2668), .B(n2669), .Z(n2575) );
  XOR2_X1 U2627 ( .A(n2670), .B(n2671), .Z(n2669) );
  XOR2_X1 U2628 ( .A(n2672), .B(n2673), .Z(n2579) );
  XOR2_X1 U2629 ( .A(n2674), .B(n2675), .Z(n2673) );
  XOR2_X1 U2630 ( .A(n2676), .B(n2677), .Z(n2583) );
  XOR2_X1 U2631 ( .A(n2678), .B(n2679), .Z(n2677) );
  XOR2_X1 U2632 ( .A(n2680), .B(n2681), .Z(n2587) );
  XOR2_X1 U2633 ( .A(n2682), .B(n2683), .Z(n2681) );
  XOR2_X1 U2634 ( .A(n2684), .B(n2685), .Z(n2591) );
  XOR2_X1 U2635 ( .A(n2686), .B(n2687), .Z(n2685) );
  XOR2_X1 U2636 ( .A(n2688), .B(n2689), .Z(n2595) );
  XOR2_X1 U2637 ( .A(n2690), .B(n2691), .Z(n2689) );
  XOR2_X1 U2638 ( .A(n2692), .B(n2693), .Z(n2599) );
  XOR2_X1 U2639 ( .A(n2694), .B(n2695), .Z(n2693) );
  XOR2_X1 U2640 ( .A(n2696), .B(n2697), .Z(n2603) );
  XOR2_X1 U2641 ( .A(n2698), .B(n2699), .Z(n2697) );
  XOR2_X1 U2642 ( .A(n2700), .B(n2701), .Z(n2607) );
  XOR2_X1 U2643 ( .A(n2702), .B(n2703), .Z(n2701) );
  XOR2_X1 U2644 ( .A(n2704), .B(n2705), .Z(n2507) );
  XOR2_X1 U2645 ( .A(n2706), .B(n2707), .Z(n2705) );
  XOR2_X1 U2646 ( .A(n2134), .B(n2135), .Z(n2364) );
  OR2_X1 U2647 ( .A1(n2708), .A2(n2709), .ZN(n2135) );
  AND2_X1 U2648 ( .A1(n2379), .A2(n2378), .ZN(n2709) );
  AND2_X1 U2649 ( .A1(n2376), .A2(n2710), .ZN(n2708) );
  OR2_X1 U2650 ( .A1(n2378), .A2(n2379), .ZN(n2710) );
  OR2_X1 U2651 ( .A1(n2562), .A2(n2148), .ZN(n2379) );
  OR2_X1 U2652 ( .A1(n2711), .A2(n2712), .ZN(n2378) );
  AND2_X1 U2653 ( .A1(n2512), .A2(n2511), .ZN(n2712) );
  AND2_X1 U2654 ( .A1(n2509), .A2(n2713), .ZN(n2711) );
  OR2_X1 U2655 ( .A1(n2511), .A2(n2512), .ZN(n2713) );
  OR2_X1 U2656 ( .A1(n2562), .A2(n2211), .ZN(n2512) );
  OR2_X1 U2657 ( .A1(n2714), .A2(n2715), .ZN(n2511) );
  AND2_X1 U2658 ( .A1(n2707), .A2(n2706), .ZN(n2715) );
  AND2_X1 U2659 ( .A1(n2704), .A2(n2716), .ZN(n2714) );
  OR2_X1 U2660 ( .A1(n2706), .A2(n2707), .ZN(n2716) );
  OR2_X1 U2661 ( .A1(n2562), .A2(n2244), .ZN(n2707) );
  OR2_X1 U2662 ( .A1(n2717), .A2(n2718), .ZN(n2706) );
  AND2_X1 U2663 ( .A1(n2703), .A2(n2702), .ZN(n2718) );
  AND2_X1 U2664 ( .A1(n2700), .A2(n2719), .ZN(n2717) );
  OR2_X1 U2665 ( .A1(n2702), .A2(n2703), .ZN(n2719) );
  OR2_X1 U2666 ( .A1(n2293), .A2(n2562), .ZN(n2703) );
  OR2_X1 U2667 ( .A1(n2720), .A2(n2721), .ZN(n2702) );
  AND2_X1 U2668 ( .A1(n2699), .A2(n2698), .ZN(n2721) );
  AND2_X1 U2669 ( .A1(n2696), .A2(n2722), .ZN(n2720) );
  OR2_X1 U2670 ( .A1(n2698), .A2(n2699), .ZN(n2722) );
  OR2_X1 U2671 ( .A1(n2340), .A2(n2562), .ZN(n2699) );
  OR2_X1 U2672 ( .A1(n2723), .A2(n2724), .ZN(n2698) );
  AND2_X1 U2673 ( .A1(n2695), .A2(n2694), .ZN(n2724) );
  AND2_X1 U2674 ( .A1(n2692), .A2(n2725), .ZN(n2723) );
  OR2_X1 U2675 ( .A1(n2694), .A2(n2695), .ZN(n2725) );
  OR2_X1 U2676 ( .A1(n2468), .A2(n2562), .ZN(n2695) );
  OR2_X1 U2677 ( .A1(n2726), .A2(n2727), .ZN(n2694) );
  AND2_X1 U2678 ( .A1(n2691), .A2(n2690), .ZN(n2727) );
  AND2_X1 U2679 ( .A1(n2688), .A2(n2728), .ZN(n2726) );
  OR2_X1 U2680 ( .A1(n2690), .A2(n2691), .ZN(n2728) );
  OR2_X1 U2681 ( .A1(n2463), .A2(n2562), .ZN(n2691) );
  OR2_X1 U2682 ( .A1(n2729), .A2(n2730), .ZN(n2690) );
  AND2_X1 U2683 ( .A1(n2687), .A2(n2686), .ZN(n2730) );
  AND2_X1 U2684 ( .A1(n2684), .A2(n2731), .ZN(n2729) );
  OR2_X1 U2685 ( .A1(n2686), .A2(n2687), .ZN(n2731) );
  OR2_X1 U2686 ( .A1(n2458), .A2(n2562), .ZN(n2687) );
  OR2_X1 U2687 ( .A1(n2732), .A2(n2733), .ZN(n2686) );
  AND2_X1 U2688 ( .A1(n2683), .A2(n2682), .ZN(n2733) );
  AND2_X1 U2689 ( .A1(n2680), .A2(n2734), .ZN(n2732) );
  OR2_X1 U2690 ( .A1(n2682), .A2(n2683), .ZN(n2734) );
  OR2_X1 U2691 ( .A1(n2453), .A2(n2562), .ZN(n2683) );
  OR2_X1 U2692 ( .A1(n2735), .A2(n2736), .ZN(n2682) );
  AND2_X1 U2693 ( .A1(n2679), .A2(n2678), .ZN(n2736) );
  AND2_X1 U2694 ( .A1(n2676), .A2(n2737), .ZN(n2735) );
  OR2_X1 U2695 ( .A1(n2678), .A2(n2679), .ZN(n2737) );
  OR2_X1 U2696 ( .A1(n2448), .A2(n2562), .ZN(n2679) );
  OR2_X1 U2697 ( .A1(n2738), .A2(n2739), .ZN(n2678) );
  AND2_X1 U2698 ( .A1(n2675), .A2(n2674), .ZN(n2739) );
  AND2_X1 U2699 ( .A1(n2672), .A2(n2740), .ZN(n2738) );
  OR2_X1 U2700 ( .A1(n2674), .A2(n2675), .ZN(n2740) );
  OR2_X1 U2701 ( .A1(n2443), .A2(n2562), .ZN(n2675) );
  OR2_X1 U2702 ( .A1(n2741), .A2(n2742), .ZN(n2674) );
  AND2_X1 U2703 ( .A1(n2671), .A2(n2670), .ZN(n2742) );
  AND2_X1 U2704 ( .A1(n2668), .A2(n2743), .ZN(n2741) );
  OR2_X1 U2705 ( .A1(n2670), .A2(n2671), .ZN(n2743) );
  OR2_X1 U2706 ( .A1(n2438), .A2(n2562), .ZN(n2671) );
  OR2_X1 U2707 ( .A1(n2744), .A2(n2745), .ZN(n2670) );
  AND2_X1 U2708 ( .A1(n2667), .A2(n2666), .ZN(n2745) );
  AND2_X1 U2709 ( .A1(n2664), .A2(n2746), .ZN(n2744) );
  OR2_X1 U2710 ( .A1(n2666), .A2(n2667), .ZN(n2746) );
  OR2_X1 U2711 ( .A1(n2433), .A2(n2562), .ZN(n2667) );
  OR2_X1 U2712 ( .A1(n2747), .A2(n2748), .ZN(n2666) );
  AND2_X1 U2713 ( .A1(n2661), .A2(n2663), .ZN(n2748) );
  AND2_X1 U2714 ( .A1(n2749), .A2(n2750), .ZN(n2747) );
  OR2_X1 U2715 ( .A1(n2663), .A2(n2661), .ZN(n2750) );
  OR2_X1 U2716 ( .A1(n2562), .A2(n2423), .ZN(n2661) );
  OR3_X1 U2717 ( .A1(n2659), .A2(n2562), .A3(n2424), .ZN(n2663) );
  INV_X1 U2718 ( .A(n2557), .ZN(n2562) );
  XOR2_X1 U2719 ( .A(n2751), .B(n2752), .Z(n2557) );
  XNOR2_X1 U2720 ( .A(c_12_), .B(d_12_), .ZN(n2751) );
  INV_X1 U2721 ( .A(n2662), .ZN(n2749) );
  OR2_X1 U2722 ( .A1(n2753), .A2(n2754), .ZN(n2662) );
  AND2_X1 U2723 ( .A1(n2755), .A2(n2756), .ZN(n2754) );
  OR2_X1 U2724 ( .A1(n2757), .A2(n2035), .ZN(n2756) );
  AND2_X1 U2725 ( .A1(n2659), .A2(n2029), .ZN(n2757) );
  AND2_X1 U2726 ( .A1(n2654), .A2(n2758), .ZN(n2753) );
  OR2_X1 U2727 ( .A1(n2759), .A2(n2039), .ZN(n2758) );
  AND2_X1 U2728 ( .A1(n2760), .A2(n2041), .ZN(n2759) );
  XOR2_X1 U2729 ( .A(n2761), .B(n2762), .Z(n2664) );
  XNOR2_X1 U2730 ( .A(n2763), .B(n2764), .ZN(n2761) );
  XOR2_X1 U2731 ( .A(n2765), .B(n2766), .Z(n2668) );
  XOR2_X1 U2732 ( .A(n2767), .B(n2768), .Z(n2766) );
  XOR2_X1 U2733 ( .A(n2769), .B(n2770), .Z(n2672) );
  XOR2_X1 U2734 ( .A(n2771), .B(n2772), .Z(n2770) );
  XOR2_X1 U2735 ( .A(n2773), .B(n2774), .Z(n2676) );
  XOR2_X1 U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  XOR2_X1 U2737 ( .A(n2777), .B(n2778), .Z(n2680) );
  XOR2_X1 U2738 ( .A(n2779), .B(n2780), .Z(n2778) );
  XOR2_X1 U2739 ( .A(n2781), .B(n2782), .Z(n2684) );
  XOR2_X1 U2740 ( .A(n2783), .B(n2784), .Z(n2782) );
  XOR2_X1 U2741 ( .A(n2785), .B(n2786), .Z(n2688) );
  XOR2_X1 U2742 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR2_X1 U2743 ( .A(n2789), .B(n2790), .Z(n2692) );
  XOR2_X1 U2744 ( .A(n2791), .B(n2792), .Z(n2790) );
  XOR2_X1 U2745 ( .A(n2793), .B(n2794), .Z(n2696) );
  XOR2_X1 U2746 ( .A(n2795), .B(n2796), .Z(n2794) );
  XOR2_X1 U2747 ( .A(n2797), .B(n2798), .Z(n2700) );
  XOR2_X1 U2748 ( .A(n2799), .B(n2800), .Z(n2798) );
  XOR2_X1 U2749 ( .A(n2801), .B(n2802), .Z(n2704) );
  XOR2_X1 U2750 ( .A(n2803), .B(n2804), .Z(n2802) );
  XOR2_X1 U2751 ( .A(n2805), .B(n2806), .Z(n2509) );
  XOR2_X1 U2752 ( .A(n2807), .B(n2808), .Z(n2806) );
  XOR2_X1 U2753 ( .A(n2809), .B(n2810), .Z(n2376) );
  XOR2_X1 U2754 ( .A(n2811), .B(n2812), .Z(n2810) );
  XOR2_X1 U2755 ( .A(n2813), .B(n2814), .Z(n2134) );
  XOR2_X1 U2756 ( .A(n2815), .B(n2816), .Z(n2814) );
  XOR2_X1 U2757 ( .A(n2142), .B(n2143), .Z(n2361) );
  OR2_X1 U2758 ( .A1(n2817), .A2(n2818), .ZN(n2143) );
  AND2_X1 U2759 ( .A1(n2816), .A2(n2815), .ZN(n2818) );
  AND2_X1 U2760 ( .A1(n2813), .A2(n2819), .ZN(n2817) );
  OR2_X1 U2761 ( .A1(n2815), .A2(n2816), .ZN(n2819) );
  OR2_X1 U2762 ( .A1(n2659), .A2(n2148), .ZN(n2816) );
  OR2_X1 U2763 ( .A1(n2820), .A2(n2821), .ZN(n2815) );
  AND2_X1 U2764 ( .A1(n2812), .A2(n2811), .ZN(n2821) );
  AND2_X1 U2765 ( .A1(n2809), .A2(n2822), .ZN(n2820) );
  OR2_X1 U2766 ( .A1(n2811), .A2(n2812), .ZN(n2822) );
  OR2_X1 U2767 ( .A1(n2659), .A2(n2211), .ZN(n2812) );
  OR2_X1 U2768 ( .A1(n2823), .A2(n2824), .ZN(n2811) );
  AND2_X1 U2769 ( .A1(n2808), .A2(n2807), .ZN(n2824) );
  AND2_X1 U2770 ( .A1(n2805), .A2(n2825), .ZN(n2823) );
  OR2_X1 U2771 ( .A1(n2807), .A2(n2808), .ZN(n2825) );
  OR2_X1 U2772 ( .A1(n2659), .A2(n2244), .ZN(n2808) );
  OR2_X1 U2773 ( .A1(n2826), .A2(n2827), .ZN(n2807) );
  AND2_X1 U2774 ( .A1(n2804), .A2(n2803), .ZN(n2827) );
  AND2_X1 U2775 ( .A1(n2801), .A2(n2828), .ZN(n2826) );
  OR2_X1 U2776 ( .A1(n2803), .A2(n2804), .ZN(n2828) );
  OR2_X1 U2777 ( .A1(n2659), .A2(n2293), .ZN(n2804) );
  OR2_X1 U2778 ( .A1(n2829), .A2(n2830), .ZN(n2803) );
  AND2_X1 U2779 ( .A1(n2800), .A2(n2799), .ZN(n2830) );
  AND2_X1 U2780 ( .A1(n2797), .A2(n2831), .ZN(n2829) );
  OR2_X1 U2781 ( .A1(n2799), .A2(n2800), .ZN(n2831) );
  OR2_X1 U2782 ( .A1(n2340), .A2(n2659), .ZN(n2800) );
  OR2_X1 U2783 ( .A1(n2832), .A2(n2833), .ZN(n2799) );
  AND2_X1 U2784 ( .A1(n2796), .A2(n2795), .ZN(n2833) );
  AND2_X1 U2785 ( .A1(n2793), .A2(n2834), .ZN(n2832) );
  OR2_X1 U2786 ( .A1(n2795), .A2(n2796), .ZN(n2834) );
  OR2_X1 U2787 ( .A1(n2468), .A2(n2659), .ZN(n2796) );
  OR2_X1 U2788 ( .A1(n2835), .A2(n2836), .ZN(n2795) );
  AND2_X1 U2789 ( .A1(n2792), .A2(n2791), .ZN(n2836) );
  AND2_X1 U2790 ( .A1(n2789), .A2(n2837), .ZN(n2835) );
  OR2_X1 U2791 ( .A1(n2791), .A2(n2792), .ZN(n2837) );
  OR2_X1 U2792 ( .A1(n2463), .A2(n2659), .ZN(n2792) );
  OR2_X1 U2793 ( .A1(n2838), .A2(n2839), .ZN(n2791) );
  AND2_X1 U2794 ( .A1(n2788), .A2(n2787), .ZN(n2839) );
  AND2_X1 U2795 ( .A1(n2785), .A2(n2840), .ZN(n2838) );
  OR2_X1 U2796 ( .A1(n2787), .A2(n2788), .ZN(n2840) );
  OR2_X1 U2797 ( .A1(n2458), .A2(n2659), .ZN(n2788) );
  OR2_X1 U2798 ( .A1(n2841), .A2(n2842), .ZN(n2787) );
  AND2_X1 U2799 ( .A1(n2784), .A2(n2783), .ZN(n2842) );
  AND2_X1 U2800 ( .A1(n2781), .A2(n2843), .ZN(n2841) );
  OR2_X1 U2801 ( .A1(n2783), .A2(n2784), .ZN(n2843) );
  OR2_X1 U2802 ( .A1(n2453), .A2(n2659), .ZN(n2784) );
  OR2_X1 U2803 ( .A1(n2844), .A2(n2845), .ZN(n2783) );
  AND2_X1 U2804 ( .A1(n2780), .A2(n2779), .ZN(n2845) );
  AND2_X1 U2805 ( .A1(n2777), .A2(n2846), .ZN(n2844) );
  OR2_X1 U2806 ( .A1(n2779), .A2(n2780), .ZN(n2846) );
  OR2_X1 U2807 ( .A1(n2448), .A2(n2659), .ZN(n2780) );
  OR2_X1 U2808 ( .A1(n2847), .A2(n2848), .ZN(n2779) );
  AND2_X1 U2809 ( .A1(n2776), .A2(n2775), .ZN(n2848) );
  AND2_X1 U2810 ( .A1(n2773), .A2(n2849), .ZN(n2847) );
  OR2_X1 U2811 ( .A1(n2775), .A2(n2776), .ZN(n2849) );
  OR2_X1 U2812 ( .A1(n2443), .A2(n2659), .ZN(n2776) );
  OR2_X1 U2813 ( .A1(n2850), .A2(n2851), .ZN(n2775) );
  AND2_X1 U2814 ( .A1(n2772), .A2(n2771), .ZN(n2851) );
  AND2_X1 U2815 ( .A1(n2769), .A2(n2852), .ZN(n2850) );
  OR2_X1 U2816 ( .A1(n2771), .A2(n2772), .ZN(n2852) );
  OR2_X1 U2817 ( .A1(n2438), .A2(n2659), .ZN(n2772) );
  OR2_X1 U2818 ( .A1(n2853), .A2(n2854), .ZN(n2771) );
  AND2_X1 U2819 ( .A1(n2768), .A2(n2767), .ZN(n2854) );
  AND2_X1 U2820 ( .A1(n2765), .A2(n2855), .ZN(n2853) );
  OR2_X1 U2821 ( .A1(n2767), .A2(n2768), .ZN(n2855) );
  OR2_X1 U2822 ( .A1(n2433), .A2(n2659), .ZN(n2768) );
  OR2_X1 U2823 ( .A1(n2856), .A2(n2857), .ZN(n2767) );
  AND2_X1 U2824 ( .A1(n2762), .A2(n2764), .ZN(n2857) );
  AND2_X1 U2825 ( .A1(n2858), .A2(n2859), .ZN(n2856) );
  OR2_X1 U2826 ( .A1(n2764), .A2(n2762), .ZN(n2859) );
  OR2_X1 U2827 ( .A1(n2659), .A2(n2423), .ZN(n2762) );
  OR3_X1 U2828 ( .A1(n2760), .A2(n2659), .A3(n2424), .ZN(n2764) );
  INV_X1 U2829 ( .A(n2654), .ZN(n2659) );
  XOR2_X1 U2830 ( .A(n2860), .B(n2861), .Z(n2654) );
  XNOR2_X1 U2831 ( .A(c_11_), .B(d_11_), .ZN(n2860) );
  INV_X1 U2832 ( .A(n2763), .ZN(n2858) );
  OR2_X1 U2833 ( .A1(n2862), .A2(n2863), .ZN(n2763) );
  AND2_X1 U2834 ( .A1(n2864), .A2(n2865), .ZN(n2863) );
  OR2_X1 U2835 ( .A1(n2866), .A2(n2035), .ZN(n2865) );
  AND2_X1 U2836 ( .A1(n2760), .A2(n2029), .ZN(n2866) );
  AND2_X1 U2837 ( .A1(n2755), .A2(n2867), .ZN(n2862) );
  OR2_X1 U2838 ( .A1(n2868), .A2(n2039), .ZN(n2867) );
  AND2_X1 U2839 ( .A1(n2869), .A2(n2041), .ZN(n2868) );
  XOR2_X1 U2840 ( .A(n2870), .B(n2871), .Z(n2765) );
  XNOR2_X1 U2841 ( .A(n2872), .B(n2873), .ZN(n2870) );
  XOR2_X1 U2842 ( .A(n2874), .B(n2875), .Z(n2769) );
  XOR2_X1 U2843 ( .A(n2876), .B(n2877), .Z(n2875) );
  XOR2_X1 U2844 ( .A(n2878), .B(n2879), .Z(n2773) );
  XOR2_X1 U2845 ( .A(n2880), .B(n2881), .Z(n2879) );
  XOR2_X1 U2846 ( .A(n2882), .B(n2883), .Z(n2777) );
  XOR2_X1 U2847 ( .A(n2884), .B(n2885), .Z(n2883) );
  XOR2_X1 U2848 ( .A(n2886), .B(n2887), .Z(n2781) );
  XOR2_X1 U2849 ( .A(n2888), .B(n2889), .Z(n2887) );
  XOR2_X1 U2850 ( .A(n2890), .B(n2891), .Z(n2785) );
  XOR2_X1 U2851 ( .A(n2892), .B(n2893), .Z(n2891) );
  XOR2_X1 U2852 ( .A(n2894), .B(n2895), .Z(n2789) );
  XOR2_X1 U2853 ( .A(n2896), .B(n2897), .Z(n2895) );
  XOR2_X1 U2854 ( .A(n2898), .B(n2899), .Z(n2793) );
  XOR2_X1 U2855 ( .A(n2900), .B(n2901), .Z(n2899) );
  XOR2_X1 U2856 ( .A(n2902), .B(n2903), .Z(n2797) );
  XOR2_X1 U2857 ( .A(n2904), .B(n2905), .Z(n2903) );
  XOR2_X1 U2858 ( .A(n2906), .B(n2907), .Z(n2801) );
  XOR2_X1 U2859 ( .A(n2908), .B(n2909), .Z(n2907) );
  XOR2_X1 U2860 ( .A(n2910), .B(n2911), .Z(n2805) );
  XOR2_X1 U2861 ( .A(n2912), .B(n2913), .Z(n2911) );
  XOR2_X1 U2862 ( .A(n2914), .B(n2915), .Z(n2809) );
  XOR2_X1 U2863 ( .A(n2916), .B(n2917), .Z(n2915) );
  XOR2_X1 U2864 ( .A(n2918), .B(n2919), .Z(n2813) );
  XOR2_X1 U2865 ( .A(n2920), .B(n2921), .Z(n2919) );
  XOR2_X1 U2866 ( .A(n2922), .B(n2923), .Z(n2142) );
  XOR2_X1 U2867 ( .A(n2924), .B(n2925), .Z(n2923) );
  INV_X1 U2868 ( .A(n2140), .ZN(n2358) );
  XNOR2_X1 U2869 ( .A(n1994), .B(n1995), .ZN(n2140) );
  OR2_X1 U2870 ( .A1(n2926), .A2(n2927), .ZN(n1995) );
  AND2_X1 U2871 ( .A1(n2925), .A2(n2924), .ZN(n2927) );
  AND2_X1 U2872 ( .A1(n2922), .A2(n2928), .ZN(n2926) );
  OR2_X1 U2873 ( .A1(n2924), .A2(n2925), .ZN(n2928) );
  OR2_X1 U2874 ( .A1(n2760), .A2(n2148), .ZN(n2925) );
  OR2_X1 U2875 ( .A1(n2929), .A2(n2930), .ZN(n2924) );
  AND2_X1 U2876 ( .A1(n2921), .A2(n2920), .ZN(n2930) );
  AND2_X1 U2877 ( .A1(n2918), .A2(n2931), .ZN(n2929) );
  OR2_X1 U2878 ( .A1(n2920), .A2(n2921), .ZN(n2931) );
  OR2_X1 U2879 ( .A1(n2760), .A2(n2211), .ZN(n2921) );
  OR2_X1 U2880 ( .A1(n2932), .A2(n2933), .ZN(n2920) );
  AND2_X1 U2881 ( .A1(n2917), .A2(n2916), .ZN(n2933) );
  AND2_X1 U2882 ( .A1(n2914), .A2(n2934), .ZN(n2932) );
  OR2_X1 U2883 ( .A1(n2916), .A2(n2917), .ZN(n2934) );
  OR2_X1 U2884 ( .A1(n2760), .A2(n2244), .ZN(n2917) );
  OR2_X1 U2885 ( .A1(n2935), .A2(n2936), .ZN(n2916) );
  AND2_X1 U2886 ( .A1(n2910), .A2(n2913), .ZN(n2936) );
  AND2_X1 U2887 ( .A1(n2937), .A2(n2912), .ZN(n2935) );
  OR2_X1 U2888 ( .A1(n2938), .A2(n2939), .ZN(n2912) );
  AND2_X1 U2889 ( .A1(n2909), .A2(n2908), .ZN(n2939) );
  AND2_X1 U2890 ( .A1(n2906), .A2(n2940), .ZN(n2938) );
  OR2_X1 U2891 ( .A1(n2908), .A2(n2909), .ZN(n2940) );
  OR2_X1 U2892 ( .A1(n2760), .A2(n2340), .ZN(n2909) );
  OR2_X1 U2893 ( .A1(n2941), .A2(n2942), .ZN(n2908) );
  AND2_X1 U2894 ( .A1(n2902), .A2(n2905), .ZN(n2942) );
  AND2_X1 U2895 ( .A1(n2943), .A2(n2904), .ZN(n2941) );
  OR2_X1 U2896 ( .A1(n2944), .A2(n2945), .ZN(n2904) );
  AND2_X1 U2897 ( .A1(n2898), .A2(n2901), .ZN(n2945) );
  AND2_X1 U2898 ( .A1(n2946), .A2(n2900), .ZN(n2944) );
  OR2_X1 U2899 ( .A1(n2947), .A2(n2948), .ZN(n2900) );
  AND2_X1 U2900 ( .A1(n2894), .A2(n2897), .ZN(n2948) );
  AND2_X1 U2901 ( .A1(n2949), .A2(n2896), .ZN(n2947) );
  OR2_X1 U2902 ( .A1(n2950), .A2(n2951), .ZN(n2896) );
  AND2_X1 U2903 ( .A1(n2890), .A2(n2893), .ZN(n2951) );
  AND2_X1 U2904 ( .A1(n2952), .A2(n2892), .ZN(n2950) );
  OR2_X1 U2905 ( .A1(n2953), .A2(n2954), .ZN(n2892) );
  AND2_X1 U2906 ( .A1(n2886), .A2(n2889), .ZN(n2954) );
  AND2_X1 U2907 ( .A1(n2955), .A2(n2888), .ZN(n2953) );
  OR2_X1 U2908 ( .A1(n2956), .A2(n2957), .ZN(n2888) );
  AND2_X1 U2909 ( .A1(n2882), .A2(n2885), .ZN(n2957) );
  AND2_X1 U2910 ( .A1(n2958), .A2(n2884), .ZN(n2956) );
  OR2_X1 U2911 ( .A1(n2959), .A2(n2960), .ZN(n2884) );
  AND2_X1 U2912 ( .A1(n2878), .A2(n2881), .ZN(n2960) );
  AND2_X1 U2913 ( .A1(n2961), .A2(n2880), .ZN(n2959) );
  OR2_X1 U2914 ( .A1(n2962), .A2(n2963), .ZN(n2880) );
  AND2_X1 U2915 ( .A1(n2874), .A2(n2877), .ZN(n2963) );
  AND2_X1 U2916 ( .A1(n2964), .A2(n2876), .ZN(n2962) );
  OR2_X1 U2917 ( .A1(n2965), .A2(n2966), .ZN(n2876) );
  AND2_X1 U2918 ( .A1(n2871), .A2(n2873), .ZN(n2966) );
  AND2_X1 U2919 ( .A1(n2967), .A2(n2968), .ZN(n2965) );
  OR2_X1 U2920 ( .A1(n2873), .A2(n2871), .ZN(n2968) );
  OR2_X1 U2921 ( .A1(n2760), .A2(n2423), .ZN(n2871) );
  OR3_X1 U2922 ( .A1(n2869), .A2(n2760), .A3(n2424), .ZN(n2873) );
  INV_X1 U2923 ( .A(n2872), .ZN(n2967) );
  OR2_X1 U2924 ( .A1(n2969), .A2(n2970), .ZN(n2872) );
  AND2_X1 U2925 ( .A1(n2971), .A2(n2972), .ZN(n2970) );
  OR2_X1 U2926 ( .A1(n2973), .A2(n2035), .ZN(n2972) );
  AND2_X1 U2927 ( .A1(n2869), .A2(n2029), .ZN(n2973) );
  AND2_X1 U2928 ( .A1(n2864), .A2(n2974), .ZN(n2969) );
  OR2_X1 U2929 ( .A1(n2975), .A2(n2039), .ZN(n2974) );
  AND2_X1 U2930 ( .A1(n2976), .A2(n2041), .ZN(n2975) );
  OR2_X1 U2931 ( .A1(n2877), .A2(n2874), .ZN(n2964) );
  XOR2_X1 U2932 ( .A(n2977), .B(n2978), .Z(n2874) );
  XNOR2_X1 U2933 ( .A(n2979), .B(n2980), .ZN(n2977) );
  OR2_X1 U2934 ( .A1(n2433), .A2(n2760), .ZN(n2877) );
  OR2_X1 U2935 ( .A1(n2881), .A2(n2878), .ZN(n2961) );
  XOR2_X1 U2936 ( .A(n2981), .B(n2982), .Z(n2878) );
  XOR2_X1 U2937 ( .A(n2983), .B(n2984), .Z(n2982) );
  OR2_X1 U2938 ( .A1(n2438), .A2(n2760), .ZN(n2881) );
  OR2_X1 U2939 ( .A1(n2885), .A2(n2882), .ZN(n2958) );
  XOR2_X1 U2940 ( .A(n2985), .B(n2986), .Z(n2882) );
  XOR2_X1 U2941 ( .A(n2987), .B(n2988), .Z(n2986) );
  OR2_X1 U2942 ( .A1(n2443), .A2(n2760), .ZN(n2885) );
  OR2_X1 U2943 ( .A1(n2889), .A2(n2886), .ZN(n2955) );
  XOR2_X1 U2944 ( .A(n2989), .B(n2990), .Z(n2886) );
  XOR2_X1 U2945 ( .A(n2991), .B(n2992), .Z(n2990) );
  OR2_X1 U2946 ( .A1(n2448), .A2(n2760), .ZN(n2889) );
  OR2_X1 U2947 ( .A1(n2893), .A2(n2890), .ZN(n2952) );
  XOR2_X1 U2948 ( .A(n2993), .B(n2994), .Z(n2890) );
  XOR2_X1 U2949 ( .A(n2995), .B(n2996), .Z(n2994) );
  OR2_X1 U2950 ( .A1(n2453), .A2(n2760), .ZN(n2893) );
  OR2_X1 U2951 ( .A1(n2897), .A2(n2894), .ZN(n2949) );
  XOR2_X1 U2952 ( .A(n2997), .B(n2998), .Z(n2894) );
  XOR2_X1 U2953 ( .A(n2999), .B(n3000), .Z(n2998) );
  OR2_X1 U2954 ( .A1(n2458), .A2(n2760), .ZN(n2897) );
  OR2_X1 U2955 ( .A1(n2901), .A2(n2898), .ZN(n2946) );
  XOR2_X1 U2956 ( .A(n3001), .B(n3002), .Z(n2898) );
  XOR2_X1 U2957 ( .A(n3003), .B(n3004), .Z(n3002) );
  OR2_X1 U2958 ( .A1(n2463), .A2(n2760), .ZN(n2901) );
  OR2_X1 U2959 ( .A1(n2905), .A2(n2902), .ZN(n2943) );
  XOR2_X1 U2960 ( .A(n3005), .B(n3006), .Z(n2902) );
  XOR2_X1 U2961 ( .A(n3007), .B(n3008), .Z(n3006) );
  OR2_X1 U2962 ( .A1(n2468), .A2(n2760), .ZN(n2905) );
  XOR2_X1 U2963 ( .A(n3009), .B(n3010), .Z(n2906) );
  XOR2_X1 U2964 ( .A(n3011), .B(n3012), .Z(n3010) );
  OR2_X1 U2965 ( .A1(n2913), .A2(n2910), .ZN(n2937) );
  XOR2_X1 U2966 ( .A(n3013), .B(n3014), .Z(n2910) );
  XOR2_X1 U2967 ( .A(n3015), .B(n3016), .Z(n3014) );
  OR2_X1 U2968 ( .A1(n2760), .A2(n2293), .ZN(n2913) );
  INV_X1 U2969 ( .A(n2755), .ZN(n2760) );
  XOR2_X1 U2970 ( .A(n3017), .B(n3018), .Z(n2755) );
  XNOR2_X1 U2971 ( .A(c_10_), .B(d_10_), .ZN(n3017) );
  XOR2_X1 U2972 ( .A(n3019), .B(n3020), .Z(n2914) );
  XOR2_X1 U2973 ( .A(n3021), .B(n3022), .Z(n3020) );
  XOR2_X1 U2974 ( .A(n3023), .B(n3024), .Z(n2918) );
  XOR2_X1 U2975 ( .A(n3025), .B(n3026), .Z(n3024) );
  XOR2_X1 U2976 ( .A(n3027), .B(n3028), .Z(n2922) );
  XOR2_X1 U2977 ( .A(n3029), .B(n3030), .Z(n3028) );
  XNOR2_X1 U2978 ( .A(n3031), .B(n3032), .ZN(n1994) );
  XNOR2_X1 U2979 ( .A(n3033), .B(n3034), .ZN(n3031) );
  INV_X1 U2980 ( .A(n1993), .ZN(n2355) );
  OR2_X1 U2981 ( .A1(n3035), .A2(n2352), .ZN(n1993) );
  INV_X1 U2982 ( .A(n3036), .ZN(n2352) );
  OR2_X1 U2983 ( .A1(n3037), .A2(n3038), .ZN(n3036) );
  AND2_X1 U2984 ( .A1(n3037), .A2(n3038), .ZN(n3035) );
  OR2_X1 U2985 ( .A1(n3039), .A2(n3040), .ZN(n3038) );
  AND2_X1 U2986 ( .A1(n3034), .A2(n3033), .ZN(n3040) );
  AND2_X1 U2987 ( .A1(n3032), .A2(n3041), .ZN(n3039) );
  OR2_X1 U2988 ( .A1(n3033), .A2(n3034), .ZN(n3041) );
  OR2_X1 U2989 ( .A1(n2869), .A2(n2148), .ZN(n3034) );
  OR2_X1 U2990 ( .A1(n3042), .A2(n3043), .ZN(n3033) );
  AND2_X1 U2991 ( .A1(n3030), .A2(n3029), .ZN(n3043) );
  AND2_X1 U2992 ( .A1(n3027), .A2(n3044), .ZN(n3042) );
  OR2_X1 U2993 ( .A1(n3029), .A2(n3030), .ZN(n3044) );
  OR2_X1 U2994 ( .A1(n2869), .A2(n2211), .ZN(n3030) );
  OR2_X1 U2995 ( .A1(n3045), .A2(n3046), .ZN(n3029) );
  AND2_X1 U2996 ( .A1(n3026), .A2(n3025), .ZN(n3046) );
  AND2_X1 U2997 ( .A1(n3023), .A2(n3047), .ZN(n3045) );
  OR2_X1 U2998 ( .A1(n3025), .A2(n3026), .ZN(n3047) );
  OR2_X1 U2999 ( .A1(n2869), .A2(n2244), .ZN(n3026) );
  OR2_X1 U3000 ( .A1(n3048), .A2(n3049), .ZN(n3025) );
  AND2_X1 U3001 ( .A1(n3022), .A2(n3021), .ZN(n3049) );
  AND2_X1 U3002 ( .A1(n3019), .A2(n3050), .ZN(n3048) );
  OR2_X1 U3003 ( .A1(n3021), .A2(n3022), .ZN(n3050) );
  OR2_X1 U3004 ( .A1(n2869), .A2(n2293), .ZN(n3022) );
  OR2_X1 U3005 ( .A1(n3051), .A2(n3052), .ZN(n3021) );
  AND2_X1 U3006 ( .A1(n3013), .A2(n3016), .ZN(n3052) );
  AND2_X1 U3007 ( .A1(n3053), .A2(n3015), .ZN(n3051) );
  OR2_X1 U3008 ( .A1(n3054), .A2(n3055), .ZN(n3015) );
  AND2_X1 U3009 ( .A1(n3012), .A2(n3011), .ZN(n3055) );
  AND2_X1 U3010 ( .A1(n3009), .A2(n3056), .ZN(n3054) );
  OR2_X1 U3011 ( .A1(n3011), .A2(n3012), .ZN(n3056) );
  OR2_X1 U3012 ( .A1(n2869), .A2(n2468), .ZN(n3012) );
  OR2_X1 U3013 ( .A1(n3057), .A2(n3058), .ZN(n3011) );
  AND2_X1 U3014 ( .A1(n3005), .A2(n3008), .ZN(n3058) );
  AND2_X1 U3015 ( .A1(n3059), .A2(n3007), .ZN(n3057) );
  OR2_X1 U3016 ( .A1(n3060), .A2(n3061), .ZN(n3007) );
  AND2_X1 U3017 ( .A1(n3001), .A2(n3004), .ZN(n3061) );
  AND2_X1 U3018 ( .A1(n3062), .A2(n3003), .ZN(n3060) );
  OR2_X1 U3019 ( .A1(n3063), .A2(n3064), .ZN(n3003) );
  AND2_X1 U3020 ( .A1(n2997), .A2(n3000), .ZN(n3064) );
  AND2_X1 U3021 ( .A1(n3065), .A2(n2999), .ZN(n3063) );
  OR2_X1 U3022 ( .A1(n3066), .A2(n3067), .ZN(n2999) );
  AND2_X1 U3023 ( .A1(n2993), .A2(n2996), .ZN(n3067) );
  AND2_X1 U3024 ( .A1(n3068), .A2(n2995), .ZN(n3066) );
  OR2_X1 U3025 ( .A1(n3069), .A2(n3070), .ZN(n2995) );
  AND2_X1 U3026 ( .A1(n2989), .A2(n2992), .ZN(n3070) );
  AND2_X1 U3027 ( .A1(n3071), .A2(n2991), .ZN(n3069) );
  OR2_X1 U3028 ( .A1(n3072), .A2(n3073), .ZN(n2991) );
  AND2_X1 U3029 ( .A1(n2985), .A2(n2988), .ZN(n3073) );
  AND2_X1 U3030 ( .A1(n3074), .A2(n2987), .ZN(n3072) );
  OR2_X1 U3031 ( .A1(n3075), .A2(n3076), .ZN(n2987) );
  AND2_X1 U3032 ( .A1(n2981), .A2(n2984), .ZN(n3076) );
  AND2_X1 U3033 ( .A1(n3077), .A2(n2983), .ZN(n3075) );
  OR2_X1 U3034 ( .A1(n3078), .A2(n3079), .ZN(n2983) );
  AND2_X1 U3035 ( .A1(n2978), .A2(n2980), .ZN(n3079) );
  AND2_X1 U3036 ( .A1(n3080), .A2(n3081), .ZN(n3078) );
  OR2_X1 U3037 ( .A1(n2980), .A2(n2978), .ZN(n3081) );
  OR2_X1 U3038 ( .A1(n2869), .A2(n2423), .ZN(n2978) );
  OR3_X1 U3039 ( .A1(n2976), .A2(n2869), .A3(n2424), .ZN(n2980) );
  INV_X1 U3040 ( .A(n2979), .ZN(n3080) );
  OR2_X1 U3041 ( .A1(n3082), .A2(n3083), .ZN(n2979) );
  AND2_X1 U3042 ( .A1(n3084), .A2(n3085), .ZN(n3083) );
  OR2_X1 U3043 ( .A1(n3086), .A2(n2035), .ZN(n3085) );
  AND2_X1 U3044 ( .A1(n2976), .A2(n2029), .ZN(n3086) );
  AND2_X1 U3045 ( .A1(n2971), .A2(n3087), .ZN(n3082) );
  OR2_X1 U3046 ( .A1(n3088), .A2(n2039), .ZN(n3087) );
  AND2_X1 U3047 ( .A1(n2311), .A2(n2041), .ZN(n3088) );
  OR2_X1 U3048 ( .A1(n2984), .A2(n2981), .ZN(n3077) );
  XOR2_X1 U3049 ( .A(n3089), .B(n3090), .Z(n2981) );
  XNOR2_X1 U3050 ( .A(n3091), .B(n3092), .ZN(n3089) );
  OR2_X1 U3051 ( .A1(n2433), .A2(n2869), .ZN(n2984) );
  OR2_X1 U3052 ( .A1(n2988), .A2(n2985), .ZN(n3074) );
  XOR2_X1 U3053 ( .A(n3093), .B(n3094), .Z(n2985) );
  XOR2_X1 U3054 ( .A(n3095), .B(n3096), .Z(n3094) );
  OR2_X1 U3055 ( .A1(n2438), .A2(n2869), .ZN(n2988) );
  OR2_X1 U3056 ( .A1(n2992), .A2(n2989), .ZN(n3071) );
  XOR2_X1 U3057 ( .A(n3097), .B(n3098), .Z(n2989) );
  XOR2_X1 U3058 ( .A(n3099), .B(n3100), .Z(n3098) );
  OR2_X1 U3059 ( .A1(n2443), .A2(n2869), .ZN(n2992) );
  OR2_X1 U3060 ( .A1(n2996), .A2(n2993), .ZN(n3068) );
  XOR2_X1 U3061 ( .A(n3101), .B(n3102), .Z(n2993) );
  XOR2_X1 U3062 ( .A(n3103), .B(n3104), .Z(n3102) );
  OR2_X1 U3063 ( .A1(n2448), .A2(n2869), .ZN(n2996) );
  OR2_X1 U3064 ( .A1(n3000), .A2(n2997), .ZN(n3065) );
  XOR2_X1 U3065 ( .A(n3105), .B(n3106), .Z(n2997) );
  XOR2_X1 U3066 ( .A(n3107), .B(n3108), .Z(n3106) );
  OR2_X1 U3067 ( .A1(n2453), .A2(n2869), .ZN(n3000) );
  OR2_X1 U3068 ( .A1(n3004), .A2(n3001), .ZN(n3062) );
  XOR2_X1 U3069 ( .A(n3109), .B(n3110), .Z(n3001) );
  XOR2_X1 U3070 ( .A(n3111), .B(n3112), .Z(n3110) );
  OR2_X1 U3071 ( .A1(n2458), .A2(n2869), .ZN(n3004) );
  OR2_X1 U3072 ( .A1(n3008), .A2(n3005), .ZN(n3059) );
  XOR2_X1 U3073 ( .A(n3113), .B(n3114), .Z(n3005) );
  XOR2_X1 U3074 ( .A(n3115), .B(n3116), .Z(n3114) );
  OR2_X1 U3075 ( .A1(n2463), .A2(n2869), .ZN(n3008) );
  XOR2_X1 U3076 ( .A(n3117), .B(n3118), .Z(n3009) );
  XOR2_X1 U3077 ( .A(n3119), .B(n3120), .Z(n3118) );
  OR2_X1 U3078 ( .A1(n3016), .A2(n3013), .ZN(n3053) );
  XOR2_X1 U3079 ( .A(n3121), .B(n3122), .Z(n3013) );
  XOR2_X1 U3080 ( .A(n3123), .B(n3124), .Z(n3122) );
  OR2_X1 U3081 ( .A1(n2869), .A2(n2340), .ZN(n3016) );
  INV_X1 U3082 ( .A(n2864), .ZN(n2869) );
  XOR2_X1 U3083 ( .A(n3125), .B(n3126), .Z(n2864) );
  XNOR2_X1 U3084 ( .A(c_9_), .B(d_9_), .ZN(n3125) );
  XOR2_X1 U3085 ( .A(n3127), .B(n3128), .Z(n3019) );
  XOR2_X1 U3086 ( .A(n3129), .B(n3130), .Z(n3128) );
  XOR2_X1 U3087 ( .A(n3131), .B(n3132), .Z(n3023) );
  XOR2_X1 U3088 ( .A(n3133), .B(n3134), .Z(n3132) );
  XOR2_X1 U3089 ( .A(n3135), .B(n3136), .Z(n3027) );
  XOR2_X1 U3090 ( .A(n3137), .B(n3138), .Z(n3136) );
  XNOR2_X1 U3091 ( .A(n3139), .B(n3140), .ZN(n3032) );
  XNOR2_X1 U3092 ( .A(n3141), .B(n3142), .ZN(n3139) );
  XNOR2_X1 U3093 ( .A(n3143), .B(n2308), .ZN(n3037) );
  XOR2_X1 U3094 ( .A(n2316), .B(n3144), .Z(n2308) );
  XOR2_X1 U3095 ( .A(n2315), .B(n2314), .Z(n3144) );
  OR2_X1 U3096 ( .A1(n2311), .A2(n2211), .ZN(n2314) );
  OR2_X1 U3097 ( .A1(n3145), .A2(n3146), .ZN(n2315) );
  AND2_X1 U3098 ( .A1(n3147), .A2(n3148), .ZN(n3146) );
  AND2_X1 U3099 ( .A1(n3149), .A2(n3150), .ZN(n3145) );
  OR2_X1 U3100 ( .A1(n3148), .A2(n3147), .ZN(n3150) );
  XOR2_X1 U3101 ( .A(n2323), .B(n3151), .Z(n2316) );
  XOR2_X1 U3102 ( .A(n2322), .B(n2321), .Z(n3151) );
  OR2_X1 U3103 ( .A1(n2271), .A2(n2244), .ZN(n2321) );
  OR2_X1 U3104 ( .A1(n3152), .A2(n3153), .ZN(n2322) );
  AND2_X1 U3105 ( .A1(n3154), .A2(n3155), .ZN(n3153) );
  AND2_X1 U3106 ( .A1(n3156), .A2(n3157), .ZN(n3152) );
  OR2_X1 U3107 ( .A1(n3155), .A2(n3154), .ZN(n3157) );
  XOR2_X1 U3108 ( .A(n2330), .B(n3158), .Z(n2323) );
  XOR2_X1 U3109 ( .A(n2329), .B(n2328), .Z(n3158) );
  OR2_X1 U3110 ( .A1(n2229), .A2(n2293), .ZN(n2328) );
  OR2_X1 U3111 ( .A1(n3159), .A2(n3160), .ZN(n2329) );
  AND2_X1 U3112 ( .A1(n3161), .A2(n3162), .ZN(n3160) );
  AND2_X1 U3113 ( .A1(n3163), .A2(n3164), .ZN(n3159) );
  OR2_X1 U3114 ( .A1(n3162), .A2(n3161), .ZN(n3164) );
  XOR2_X1 U3115 ( .A(n2337), .B(n3165), .Z(n2330) );
  XOR2_X1 U3116 ( .A(n2336), .B(n2335), .Z(n3165) );
  OR2_X1 U3117 ( .A1(n2203), .A2(n2340), .ZN(n2335) );
  OR2_X1 U3118 ( .A1(n3166), .A2(n3167), .ZN(n2336) );
  AND2_X1 U3119 ( .A1(n3168), .A2(n3169), .ZN(n3167) );
  AND2_X1 U3120 ( .A1(n3170), .A2(n3171), .ZN(n3166) );
  OR2_X1 U3121 ( .A1(n3169), .A2(n3168), .ZN(n3171) );
  XOR2_X1 U3122 ( .A(n2345), .B(n3172), .Z(n2337) );
  XOR2_X1 U3123 ( .A(n2344), .B(n2343), .Z(n3172) );
  OR2_X1 U3124 ( .A1(n2176), .A2(n2468), .ZN(n2343) );
  OR2_X1 U3125 ( .A1(n3173), .A2(n3174), .ZN(n2344) );
  AND2_X1 U3126 ( .A1(n3175), .A2(n3176), .ZN(n3174) );
  AND2_X1 U3127 ( .A1(n3177), .A2(n3178), .ZN(n3173) );
  OR2_X1 U3128 ( .A1(n3176), .A2(n3175), .ZN(n3178) );
  XOR2_X1 U3129 ( .A(n3179), .B(n3180), .Z(n2345) );
  XOR2_X1 U3130 ( .A(n3181), .B(n3182), .Z(n3180) );
  XNOR2_X1 U3131 ( .A(n2307), .B(n2306), .ZN(n3143) );
  OR2_X1 U3132 ( .A1(n2976), .A2(n2148), .ZN(n2306) );
  OR2_X1 U3133 ( .A1(n3183), .A2(n3184), .ZN(n2307) );
  AND2_X1 U3134 ( .A1(n3142), .A2(n3141), .ZN(n3184) );
  AND2_X1 U3135 ( .A1(n3140), .A2(n3185), .ZN(n3183) );
  OR2_X1 U3136 ( .A1(n3141), .A2(n3142), .ZN(n3185) );
  OR2_X1 U3137 ( .A1(n2976), .A2(n2211), .ZN(n3142) );
  OR2_X1 U3138 ( .A1(n3186), .A2(n3187), .ZN(n3141) );
  AND2_X1 U3139 ( .A1(n3138), .A2(n3137), .ZN(n3187) );
  AND2_X1 U3140 ( .A1(n3135), .A2(n3188), .ZN(n3186) );
  OR2_X1 U3141 ( .A1(n3137), .A2(n3138), .ZN(n3188) );
  OR2_X1 U3142 ( .A1(n2976), .A2(n2244), .ZN(n3138) );
  OR2_X1 U3143 ( .A1(n3189), .A2(n3190), .ZN(n3137) );
  AND2_X1 U3144 ( .A1(n3134), .A2(n3133), .ZN(n3190) );
  AND2_X1 U3145 ( .A1(n3131), .A2(n3191), .ZN(n3189) );
  OR2_X1 U3146 ( .A1(n3133), .A2(n3134), .ZN(n3191) );
  OR2_X1 U3147 ( .A1(n2976), .A2(n2293), .ZN(n3134) );
  OR2_X1 U3148 ( .A1(n3192), .A2(n3193), .ZN(n3133) );
  AND2_X1 U3149 ( .A1(n3130), .A2(n3129), .ZN(n3193) );
  AND2_X1 U3150 ( .A1(n3127), .A2(n3194), .ZN(n3192) );
  OR2_X1 U3151 ( .A1(n3129), .A2(n3130), .ZN(n3194) );
  OR2_X1 U3152 ( .A1(n2976), .A2(n2340), .ZN(n3130) );
  OR2_X1 U3153 ( .A1(n3195), .A2(n3196), .ZN(n3129) );
  AND2_X1 U3154 ( .A1(n3121), .A2(n3124), .ZN(n3196) );
  AND2_X1 U3155 ( .A1(n3197), .A2(n3123), .ZN(n3195) );
  OR2_X1 U3156 ( .A1(n3198), .A2(n3199), .ZN(n3123) );
  AND2_X1 U3157 ( .A1(n3120), .A2(n3119), .ZN(n3199) );
  AND2_X1 U3158 ( .A1(n3117), .A2(n3200), .ZN(n3198) );
  OR2_X1 U3159 ( .A1(n3119), .A2(n3120), .ZN(n3200) );
  OR2_X1 U3160 ( .A1(n2976), .A2(n2463), .ZN(n3120) );
  OR2_X1 U3161 ( .A1(n3201), .A2(n3202), .ZN(n3119) );
  AND2_X1 U3162 ( .A1(n3113), .A2(n3116), .ZN(n3202) );
  AND2_X1 U3163 ( .A1(n3203), .A2(n3115), .ZN(n3201) );
  OR2_X1 U3164 ( .A1(n3204), .A2(n3205), .ZN(n3115) );
  AND2_X1 U3165 ( .A1(n3109), .A2(n3112), .ZN(n3205) );
  AND2_X1 U3166 ( .A1(n3206), .A2(n3111), .ZN(n3204) );
  OR2_X1 U3167 ( .A1(n3207), .A2(n3208), .ZN(n3111) );
  AND2_X1 U3168 ( .A1(n3105), .A2(n3108), .ZN(n3208) );
  AND2_X1 U3169 ( .A1(n3209), .A2(n3107), .ZN(n3207) );
  OR2_X1 U3170 ( .A1(n3210), .A2(n3211), .ZN(n3107) );
  AND2_X1 U3171 ( .A1(n3101), .A2(n3104), .ZN(n3211) );
  AND2_X1 U3172 ( .A1(n3212), .A2(n3103), .ZN(n3210) );
  OR2_X1 U3173 ( .A1(n3213), .A2(n3214), .ZN(n3103) );
  AND2_X1 U3174 ( .A1(n3097), .A2(n3100), .ZN(n3214) );
  AND2_X1 U3175 ( .A1(n3215), .A2(n3099), .ZN(n3213) );
  OR2_X1 U3176 ( .A1(n3216), .A2(n3217), .ZN(n3099) );
  AND2_X1 U3177 ( .A1(n3093), .A2(n3096), .ZN(n3217) );
  AND2_X1 U3178 ( .A1(n3218), .A2(n3095), .ZN(n3216) );
  OR2_X1 U3179 ( .A1(n3219), .A2(n3220), .ZN(n3095) );
  AND2_X1 U3180 ( .A1(n3090), .A2(n3092), .ZN(n3220) );
  AND2_X1 U3181 ( .A1(n3221), .A2(n3222), .ZN(n3219) );
  OR2_X1 U3182 ( .A1(n3092), .A2(n3090), .ZN(n3222) );
  OR2_X1 U3183 ( .A1(n2976), .A2(n2423), .ZN(n3090) );
  OR3_X1 U3184 ( .A1(n2311), .A2(n2976), .A3(n2424), .ZN(n3092) );
  INV_X1 U3185 ( .A(n3091), .ZN(n3221) );
  OR2_X1 U3186 ( .A1(n3223), .A2(n3224), .ZN(n3091) );
  AND2_X1 U3187 ( .A1(n3225), .A2(n3226), .ZN(n3224) );
  OR2_X1 U3188 ( .A1(n3227), .A2(n2035), .ZN(n3226) );
  AND2_X1 U3189 ( .A1(n2311), .A2(n2029), .ZN(n3227) );
  AND2_X1 U3190 ( .A1(n3084), .A2(n3228), .ZN(n3223) );
  OR2_X1 U3191 ( .A1(n3229), .A2(n2039), .ZN(n3228) );
  AND2_X1 U3192 ( .A1(n2271), .A2(n2041), .ZN(n3229) );
  OR2_X1 U3193 ( .A1(n3096), .A2(n3093), .ZN(n3218) );
  XOR2_X1 U3194 ( .A(n3230), .B(n3231), .Z(n3093) );
  XNOR2_X1 U3195 ( .A(n3232), .B(n3233), .ZN(n3230) );
  OR2_X1 U3196 ( .A1(n2433), .A2(n2976), .ZN(n3096) );
  OR2_X1 U3197 ( .A1(n3100), .A2(n3097), .ZN(n3215) );
  XOR2_X1 U3198 ( .A(n3234), .B(n3235), .Z(n3097) );
  XOR2_X1 U3199 ( .A(n3236), .B(n3237), .Z(n3235) );
  OR2_X1 U3200 ( .A1(n2438), .A2(n2976), .ZN(n3100) );
  OR2_X1 U3201 ( .A1(n3104), .A2(n3101), .ZN(n3212) );
  XOR2_X1 U3202 ( .A(n3238), .B(n3239), .Z(n3101) );
  XOR2_X1 U3203 ( .A(n3240), .B(n3241), .Z(n3239) );
  OR2_X1 U3204 ( .A1(n2443), .A2(n2976), .ZN(n3104) );
  OR2_X1 U3205 ( .A1(n3108), .A2(n3105), .ZN(n3209) );
  XOR2_X1 U3206 ( .A(n3242), .B(n3243), .Z(n3105) );
  XOR2_X1 U3207 ( .A(n3244), .B(n3245), .Z(n3243) );
  OR2_X1 U3208 ( .A1(n2448), .A2(n2976), .ZN(n3108) );
  OR2_X1 U3209 ( .A1(n3112), .A2(n3109), .ZN(n3206) );
  XOR2_X1 U3210 ( .A(n3246), .B(n3247), .Z(n3109) );
  XOR2_X1 U3211 ( .A(n3248), .B(n3249), .Z(n3247) );
  OR2_X1 U3212 ( .A1(n2453), .A2(n2976), .ZN(n3112) );
  OR2_X1 U3213 ( .A1(n3116), .A2(n3113), .ZN(n3203) );
  XOR2_X1 U3214 ( .A(n3250), .B(n3251), .Z(n3113) );
  XOR2_X1 U3215 ( .A(n3252), .B(n3253), .Z(n3251) );
  OR2_X1 U3216 ( .A1(n2458), .A2(n2976), .ZN(n3116) );
  XOR2_X1 U3217 ( .A(n3254), .B(n3255), .Z(n3117) );
  XOR2_X1 U3218 ( .A(n3256), .B(n3257), .Z(n3255) );
  OR2_X1 U3219 ( .A1(n3124), .A2(n3121), .ZN(n3197) );
  XOR2_X1 U3220 ( .A(n3258), .B(n3259), .Z(n3121) );
  XOR2_X1 U3221 ( .A(n3260), .B(n3261), .Z(n3259) );
  OR2_X1 U3222 ( .A1(n2976), .A2(n2468), .ZN(n3124) );
  INV_X1 U3223 ( .A(n2971), .ZN(n2976) );
  XOR2_X1 U3224 ( .A(n3262), .B(n3263), .Z(n2971) );
  XNOR2_X1 U3225 ( .A(c_8_), .B(d_8_), .ZN(n3262) );
  XOR2_X1 U3226 ( .A(n3264), .B(n3265), .Z(n3127) );
  XOR2_X1 U3227 ( .A(n3266), .B(n3267), .Z(n3265) );
  XOR2_X1 U3228 ( .A(n3268), .B(n3269), .Z(n3131) );
  XOR2_X1 U3229 ( .A(n3270), .B(n3271), .Z(n3269) );
  XNOR2_X1 U3230 ( .A(n3272), .B(n3273), .ZN(n3135) );
  XNOR2_X1 U3231 ( .A(n3274), .B(n3275), .ZN(n3272) );
  XOR2_X1 U3232 ( .A(n3149), .B(n3276), .Z(n3140) );
  XOR2_X1 U3233 ( .A(n3148), .B(n3147), .Z(n3276) );
  OR2_X1 U3234 ( .A1(n2311), .A2(n2244), .ZN(n3147) );
  OR2_X1 U3235 ( .A1(n3277), .A2(n3278), .ZN(n3148) );
  AND2_X1 U3236 ( .A1(n3275), .A2(n3274), .ZN(n3278) );
  AND2_X1 U3237 ( .A1(n3273), .A2(n3279), .ZN(n3277) );
  OR2_X1 U3238 ( .A1(n3274), .A2(n3275), .ZN(n3279) );
  OR2_X1 U3239 ( .A1(n2311), .A2(n2293), .ZN(n3275) );
  OR2_X1 U3240 ( .A1(n3280), .A2(n3281), .ZN(n3274) );
  AND2_X1 U3241 ( .A1(n3271), .A2(n3270), .ZN(n3281) );
  AND2_X1 U3242 ( .A1(n3268), .A2(n3282), .ZN(n3280) );
  OR2_X1 U3243 ( .A1(n3270), .A2(n3271), .ZN(n3282) );
  OR2_X1 U3244 ( .A1(n2311), .A2(n2340), .ZN(n3271) );
  OR2_X1 U3245 ( .A1(n3283), .A2(n3284), .ZN(n3270) );
  AND2_X1 U3246 ( .A1(n3267), .A2(n3266), .ZN(n3284) );
  AND2_X1 U3247 ( .A1(n3264), .A2(n3285), .ZN(n3283) );
  OR2_X1 U3248 ( .A1(n3266), .A2(n3267), .ZN(n3285) );
  OR2_X1 U3249 ( .A1(n2311), .A2(n2468), .ZN(n3267) );
  OR2_X1 U3250 ( .A1(n3286), .A2(n3287), .ZN(n3266) );
  AND2_X1 U3251 ( .A1(n3258), .A2(n3261), .ZN(n3287) );
  AND2_X1 U3252 ( .A1(n3288), .A2(n3260), .ZN(n3286) );
  OR2_X1 U3253 ( .A1(n3289), .A2(n3290), .ZN(n3260) );
  AND2_X1 U3254 ( .A1(n3257), .A2(n3256), .ZN(n3290) );
  AND2_X1 U3255 ( .A1(n3254), .A2(n3291), .ZN(n3289) );
  OR2_X1 U3256 ( .A1(n3256), .A2(n3257), .ZN(n3291) );
  OR2_X1 U3257 ( .A1(n2311), .A2(n2458), .ZN(n3257) );
  OR2_X1 U3258 ( .A1(n3292), .A2(n3293), .ZN(n3256) );
  AND2_X1 U3259 ( .A1(n3250), .A2(n3253), .ZN(n3293) );
  AND2_X1 U3260 ( .A1(n3294), .A2(n3252), .ZN(n3292) );
  OR2_X1 U3261 ( .A1(n3295), .A2(n3296), .ZN(n3252) );
  AND2_X1 U3262 ( .A1(n3246), .A2(n3249), .ZN(n3296) );
  AND2_X1 U3263 ( .A1(n3297), .A2(n3248), .ZN(n3295) );
  OR2_X1 U3264 ( .A1(n3298), .A2(n3299), .ZN(n3248) );
  AND2_X1 U3265 ( .A1(n3242), .A2(n3245), .ZN(n3299) );
  AND2_X1 U3266 ( .A1(n3300), .A2(n3244), .ZN(n3298) );
  OR2_X1 U3267 ( .A1(n3301), .A2(n3302), .ZN(n3244) );
  AND2_X1 U3268 ( .A1(n3238), .A2(n3241), .ZN(n3302) );
  AND2_X1 U3269 ( .A1(n3303), .A2(n3240), .ZN(n3301) );
  OR2_X1 U3270 ( .A1(n3304), .A2(n3305), .ZN(n3240) );
  AND2_X1 U3271 ( .A1(n3234), .A2(n3237), .ZN(n3305) );
  AND2_X1 U3272 ( .A1(n3306), .A2(n3236), .ZN(n3304) );
  OR2_X1 U3273 ( .A1(n3307), .A2(n3308), .ZN(n3236) );
  AND2_X1 U3274 ( .A1(n3231), .A2(n3233), .ZN(n3308) );
  AND2_X1 U3275 ( .A1(n3309), .A2(n3310), .ZN(n3307) );
  OR2_X1 U3276 ( .A1(n3233), .A2(n3231), .ZN(n3310) );
  OR2_X1 U3277 ( .A1(n2311), .A2(n2423), .ZN(n3231) );
  OR3_X1 U3278 ( .A1(n2271), .A2(n2311), .A3(n2424), .ZN(n3233) );
  INV_X1 U3279 ( .A(n3232), .ZN(n3309) );
  OR2_X1 U3280 ( .A1(n3311), .A2(n3312), .ZN(n3232) );
  AND2_X1 U3281 ( .A1(n3313), .A2(n3314), .ZN(n3312) );
  OR2_X1 U3282 ( .A1(n3315), .A2(n2035), .ZN(n3314) );
  AND2_X1 U3283 ( .A1(n2271), .A2(n2029), .ZN(n3315) );
  AND2_X1 U3284 ( .A1(n3225), .A2(n3316), .ZN(n3311) );
  OR2_X1 U3285 ( .A1(n3317), .A2(n2039), .ZN(n3316) );
  AND2_X1 U3286 ( .A1(n2229), .A2(n2041), .ZN(n3317) );
  OR2_X1 U3287 ( .A1(n3237), .A2(n3234), .ZN(n3306) );
  XOR2_X1 U3288 ( .A(n3318), .B(n3319), .Z(n3234) );
  XNOR2_X1 U3289 ( .A(n3320), .B(n3321), .ZN(n3318) );
  OR2_X1 U3290 ( .A1(n2433), .A2(n2311), .ZN(n3237) );
  OR2_X1 U3291 ( .A1(n3241), .A2(n3238), .ZN(n3303) );
  XOR2_X1 U3292 ( .A(n3322), .B(n3323), .Z(n3238) );
  XOR2_X1 U3293 ( .A(n3324), .B(n3325), .Z(n3323) );
  OR2_X1 U3294 ( .A1(n2438), .A2(n2311), .ZN(n3241) );
  OR2_X1 U3295 ( .A1(n3245), .A2(n3242), .ZN(n3300) );
  XOR2_X1 U3296 ( .A(n3326), .B(n3327), .Z(n3242) );
  XOR2_X1 U3297 ( .A(n3328), .B(n3329), .Z(n3327) );
  OR2_X1 U3298 ( .A1(n2443), .A2(n2311), .ZN(n3245) );
  OR2_X1 U3299 ( .A1(n3249), .A2(n3246), .ZN(n3297) );
  XOR2_X1 U3300 ( .A(n3330), .B(n3331), .Z(n3246) );
  XOR2_X1 U3301 ( .A(n3332), .B(n3333), .Z(n3331) );
  OR2_X1 U3302 ( .A1(n2448), .A2(n2311), .ZN(n3249) );
  OR2_X1 U3303 ( .A1(n3253), .A2(n3250), .ZN(n3294) );
  XOR2_X1 U3304 ( .A(n3334), .B(n3335), .Z(n3250) );
  XOR2_X1 U3305 ( .A(n3336), .B(n3337), .Z(n3335) );
  OR2_X1 U3306 ( .A1(n2453), .A2(n2311), .ZN(n3253) );
  XOR2_X1 U3307 ( .A(n3338), .B(n3339), .Z(n3254) );
  XOR2_X1 U3308 ( .A(n3340), .B(n3341), .Z(n3339) );
  OR2_X1 U3309 ( .A1(n3261), .A2(n3258), .ZN(n3288) );
  XOR2_X1 U3310 ( .A(n3342), .B(n3343), .Z(n3258) );
  XOR2_X1 U3311 ( .A(n3344), .B(n3345), .Z(n3343) );
  OR2_X1 U3312 ( .A1(n2311), .A2(n2463), .ZN(n3261) );
  INV_X1 U3313 ( .A(n3084), .ZN(n2311) );
  XOR2_X1 U3314 ( .A(n3346), .B(n3347), .Z(n3084) );
  XNOR2_X1 U3315 ( .A(c_7_), .B(d_7_), .ZN(n3346) );
  XOR2_X1 U3316 ( .A(n3348), .B(n3349), .Z(n3264) );
  XOR2_X1 U3317 ( .A(n3350), .B(n3351), .Z(n3349) );
  XOR2_X1 U3318 ( .A(n3352), .B(n3353), .Z(n3268) );
  XOR2_X1 U3319 ( .A(n3354), .B(n3355), .Z(n3353) );
  XOR2_X1 U3320 ( .A(n3356), .B(n3357), .Z(n3273) );
  XOR2_X1 U3321 ( .A(n3358), .B(n3359), .Z(n3357) );
  XOR2_X1 U3322 ( .A(n3156), .B(n3360), .Z(n3149) );
  XOR2_X1 U3323 ( .A(n3155), .B(n3154), .Z(n3360) );
  OR2_X1 U3324 ( .A1(n2271), .A2(n2293), .ZN(n3154) );
  OR2_X1 U3325 ( .A1(n3361), .A2(n3362), .ZN(n3155) );
  AND2_X1 U3326 ( .A1(n3359), .A2(n3358), .ZN(n3362) );
  AND2_X1 U3327 ( .A1(n3356), .A2(n3363), .ZN(n3361) );
  OR2_X1 U3328 ( .A1(n3358), .A2(n3359), .ZN(n3363) );
  OR2_X1 U3329 ( .A1(n2271), .A2(n2340), .ZN(n3359) );
  OR2_X1 U3330 ( .A1(n3364), .A2(n3365), .ZN(n3358) );
  AND2_X1 U3331 ( .A1(n3355), .A2(n3354), .ZN(n3365) );
  AND2_X1 U3332 ( .A1(n3352), .A2(n3366), .ZN(n3364) );
  OR2_X1 U3333 ( .A1(n3354), .A2(n3355), .ZN(n3366) );
  OR2_X1 U3334 ( .A1(n2271), .A2(n2468), .ZN(n3355) );
  OR2_X1 U3335 ( .A1(n3367), .A2(n3368), .ZN(n3354) );
  AND2_X1 U3336 ( .A1(n3351), .A2(n3350), .ZN(n3368) );
  AND2_X1 U3337 ( .A1(n3348), .A2(n3369), .ZN(n3367) );
  OR2_X1 U3338 ( .A1(n3350), .A2(n3351), .ZN(n3369) );
  OR2_X1 U3339 ( .A1(n2271), .A2(n2463), .ZN(n3351) );
  OR2_X1 U3340 ( .A1(n3370), .A2(n3371), .ZN(n3350) );
  AND2_X1 U3341 ( .A1(n3342), .A2(n3345), .ZN(n3371) );
  AND2_X1 U3342 ( .A1(n3372), .A2(n3344), .ZN(n3370) );
  OR2_X1 U3343 ( .A1(n3373), .A2(n3374), .ZN(n3344) );
  AND2_X1 U3344 ( .A1(n3341), .A2(n3340), .ZN(n3374) );
  AND2_X1 U3345 ( .A1(n3338), .A2(n3375), .ZN(n3373) );
  OR2_X1 U3346 ( .A1(n3340), .A2(n3341), .ZN(n3375) );
  OR2_X1 U3347 ( .A1(n2271), .A2(n2453), .ZN(n3341) );
  OR2_X1 U3348 ( .A1(n3376), .A2(n3377), .ZN(n3340) );
  AND2_X1 U3349 ( .A1(n3334), .A2(n3337), .ZN(n3377) );
  AND2_X1 U3350 ( .A1(n3378), .A2(n3336), .ZN(n3376) );
  OR2_X1 U3351 ( .A1(n3379), .A2(n3380), .ZN(n3336) );
  AND2_X1 U3352 ( .A1(n3330), .A2(n3333), .ZN(n3380) );
  AND2_X1 U3353 ( .A1(n3381), .A2(n3332), .ZN(n3379) );
  OR2_X1 U3354 ( .A1(n3382), .A2(n3383), .ZN(n3332) );
  AND2_X1 U3355 ( .A1(n3326), .A2(n3329), .ZN(n3383) );
  AND2_X1 U3356 ( .A1(n3384), .A2(n3328), .ZN(n3382) );
  OR2_X1 U3357 ( .A1(n3385), .A2(n3386), .ZN(n3328) );
  AND2_X1 U3358 ( .A1(n3322), .A2(n3325), .ZN(n3386) );
  AND2_X1 U3359 ( .A1(n3387), .A2(n3324), .ZN(n3385) );
  OR2_X1 U3360 ( .A1(n3388), .A2(n3389), .ZN(n3324) );
  AND2_X1 U3361 ( .A1(n3319), .A2(n3321), .ZN(n3389) );
  AND2_X1 U3362 ( .A1(n3390), .A2(n3391), .ZN(n3388) );
  OR2_X1 U3363 ( .A1(n3321), .A2(n3319), .ZN(n3391) );
  OR2_X1 U3364 ( .A1(n2271), .A2(n2423), .ZN(n3319) );
  OR3_X1 U3365 ( .A1(n2229), .A2(n2271), .A3(n2424), .ZN(n3321) );
  INV_X1 U3366 ( .A(n3320), .ZN(n3390) );
  OR2_X1 U3367 ( .A1(n3392), .A2(n3393), .ZN(n3320) );
  AND2_X1 U3368 ( .A1(n3394), .A2(n3395), .ZN(n3393) );
  OR2_X1 U3369 ( .A1(n3396), .A2(n2035), .ZN(n3395) );
  AND2_X1 U3370 ( .A1(n2229), .A2(n2029), .ZN(n3396) );
  AND2_X1 U3371 ( .A1(n3313), .A2(n3397), .ZN(n3392) );
  OR2_X1 U3372 ( .A1(n3398), .A2(n2039), .ZN(n3397) );
  AND2_X1 U3373 ( .A1(n2203), .A2(n2041), .ZN(n3398) );
  OR2_X1 U3374 ( .A1(n3325), .A2(n3322), .ZN(n3387) );
  XOR2_X1 U3375 ( .A(n3399), .B(n3400), .Z(n3322) );
  XNOR2_X1 U3376 ( .A(n3401), .B(n3402), .ZN(n3399) );
  OR2_X1 U3377 ( .A1(n2433), .A2(n2271), .ZN(n3325) );
  OR2_X1 U3378 ( .A1(n3329), .A2(n3326), .ZN(n3384) );
  XOR2_X1 U3379 ( .A(n3403), .B(n3404), .Z(n3326) );
  XOR2_X1 U3380 ( .A(n3405), .B(n3406), .Z(n3404) );
  OR2_X1 U3381 ( .A1(n2438), .A2(n2271), .ZN(n3329) );
  OR2_X1 U3382 ( .A1(n3333), .A2(n3330), .ZN(n3381) );
  XOR2_X1 U3383 ( .A(n3407), .B(n3408), .Z(n3330) );
  XOR2_X1 U3384 ( .A(n3409), .B(n3410), .Z(n3408) );
  OR2_X1 U3385 ( .A1(n2443), .A2(n2271), .ZN(n3333) );
  OR2_X1 U3386 ( .A1(n3337), .A2(n3334), .ZN(n3378) );
  XOR2_X1 U3387 ( .A(n3411), .B(n3412), .Z(n3334) );
  XOR2_X1 U3388 ( .A(n3413), .B(n3414), .Z(n3412) );
  OR2_X1 U3389 ( .A1(n2448), .A2(n2271), .ZN(n3337) );
  XOR2_X1 U3390 ( .A(n3415), .B(n3416), .Z(n3338) );
  XOR2_X1 U3391 ( .A(n3417), .B(n3418), .Z(n3416) );
  OR2_X1 U3392 ( .A1(n3345), .A2(n3342), .ZN(n3372) );
  XOR2_X1 U3393 ( .A(n3419), .B(n3420), .Z(n3342) );
  XOR2_X1 U3394 ( .A(n3421), .B(n3422), .Z(n3420) );
  OR2_X1 U3395 ( .A1(n2271), .A2(n2458), .ZN(n3345) );
  INV_X1 U3396 ( .A(n3225), .ZN(n2271) );
  XOR2_X1 U3397 ( .A(n3423), .B(n3424), .Z(n3225) );
  XNOR2_X1 U3398 ( .A(c_6_), .B(d_6_), .ZN(n3423) );
  XOR2_X1 U3399 ( .A(n3425), .B(n3426), .Z(n3348) );
  XOR2_X1 U3400 ( .A(n3427), .B(n3428), .Z(n3426) );
  XOR2_X1 U3401 ( .A(n3429), .B(n3430), .Z(n3352) );
  XOR2_X1 U3402 ( .A(n3431), .B(n3432), .Z(n3430) );
  XOR2_X1 U3403 ( .A(n3433), .B(n3434), .Z(n3356) );
  XOR2_X1 U3404 ( .A(n3435), .B(n3436), .Z(n3434) );
  XOR2_X1 U3405 ( .A(n3163), .B(n3437), .Z(n3156) );
  XOR2_X1 U3406 ( .A(n3162), .B(n3161), .Z(n3437) );
  OR2_X1 U3407 ( .A1(n2229), .A2(n2340), .ZN(n3161) );
  OR2_X1 U3408 ( .A1(n3438), .A2(n3439), .ZN(n3162) );
  AND2_X1 U3409 ( .A1(n3436), .A2(n3435), .ZN(n3439) );
  AND2_X1 U3410 ( .A1(n3433), .A2(n3440), .ZN(n3438) );
  OR2_X1 U3411 ( .A1(n3435), .A2(n3436), .ZN(n3440) );
  OR2_X1 U3412 ( .A1(n2229), .A2(n2468), .ZN(n3436) );
  OR2_X1 U3413 ( .A1(n3441), .A2(n3442), .ZN(n3435) );
  AND2_X1 U3414 ( .A1(n3432), .A2(n3431), .ZN(n3442) );
  AND2_X1 U3415 ( .A1(n3429), .A2(n3443), .ZN(n3441) );
  OR2_X1 U3416 ( .A1(n3431), .A2(n3432), .ZN(n3443) );
  OR2_X1 U3417 ( .A1(n2229), .A2(n2463), .ZN(n3432) );
  OR2_X1 U3418 ( .A1(n3444), .A2(n3445), .ZN(n3431) );
  AND2_X1 U3419 ( .A1(n3428), .A2(n3427), .ZN(n3445) );
  AND2_X1 U3420 ( .A1(n3425), .A2(n3446), .ZN(n3444) );
  OR2_X1 U3421 ( .A1(n3427), .A2(n3428), .ZN(n3446) );
  OR2_X1 U3422 ( .A1(n2229), .A2(n2458), .ZN(n3428) );
  OR2_X1 U3423 ( .A1(n3447), .A2(n3448), .ZN(n3427) );
  AND2_X1 U3424 ( .A1(n3419), .A2(n3422), .ZN(n3448) );
  AND2_X1 U3425 ( .A1(n3449), .A2(n3421), .ZN(n3447) );
  OR2_X1 U3426 ( .A1(n3450), .A2(n3451), .ZN(n3421) );
  AND2_X1 U3427 ( .A1(n3418), .A2(n3417), .ZN(n3451) );
  AND2_X1 U3428 ( .A1(n3415), .A2(n3452), .ZN(n3450) );
  OR2_X1 U3429 ( .A1(n3417), .A2(n3418), .ZN(n3452) );
  OR2_X1 U3430 ( .A1(n2229), .A2(n2448), .ZN(n3418) );
  OR2_X1 U3431 ( .A1(n3453), .A2(n3454), .ZN(n3417) );
  AND2_X1 U3432 ( .A1(n3411), .A2(n3414), .ZN(n3454) );
  AND2_X1 U3433 ( .A1(n3455), .A2(n3413), .ZN(n3453) );
  OR2_X1 U3434 ( .A1(n3456), .A2(n3457), .ZN(n3413) );
  AND2_X1 U3435 ( .A1(n3407), .A2(n3410), .ZN(n3457) );
  AND2_X1 U3436 ( .A1(n3458), .A2(n3409), .ZN(n3456) );
  OR2_X1 U3437 ( .A1(n3459), .A2(n3460), .ZN(n3409) );
  AND2_X1 U3438 ( .A1(n3403), .A2(n3406), .ZN(n3460) );
  AND2_X1 U3439 ( .A1(n3461), .A2(n3405), .ZN(n3459) );
  OR2_X1 U3440 ( .A1(n3462), .A2(n3463), .ZN(n3405) );
  AND2_X1 U3441 ( .A1(n3400), .A2(n3402), .ZN(n3463) );
  AND2_X1 U3442 ( .A1(n3464), .A2(n3465), .ZN(n3462) );
  OR2_X1 U3443 ( .A1(n3402), .A2(n3400), .ZN(n3465) );
  OR2_X1 U3444 ( .A1(n2229), .A2(n2423), .ZN(n3400) );
  OR3_X1 U3445 ( .A1(n2203), .A2(n2229), .A3(n2424), .ZN(n3402) );
  INV_X1 U3446 ( .A(n3401), .ZN(n3464) );
  OR2_X1 U3447 ( .A1(n3466), .A2(n3467), .ZN(n3401) );
  AND2_X1 U3448 ( .A1(n3468), .A2(n3469), .ZN(n3467) );
  OR2_X1 U3449 ( .A1(n3470), .A2(n2035), .ZN(n3469) );
  AND2_X1 U3450 ( .A1(n2203), .A2(n2029), .ZN(n3470) );
  AND2_X1 U3451 ( .A1(n3394), .A2(n3471), .ZN(n3466) );
  OR2_X1 U3452 ( .A1(n3472), .A2(n2039), .ZN(n3471) );
  AND2_X1 U3453 ( .A1(n2176), .A2(n2041), .ZN(n3472) );
  OR2_X1 U3454 ( .A1(n3406), .A2(n3403), .ZN(n3461) );
  XOR2_X1 U3455 ( .A(n3473), .B(n3474), .Z(n3403) );
  XNOR2_X1 U3456 ( .A(n3475), .B(n3476), .ZN(n3473) );
  OR2_X1 U3457 ( .A1(n2433), .A2(n2229), .ZN(n3406) );
  OR2_X1 U3458 ( .A1(n3410), .A2(n3407), .ZN(n3458) );
  XOR2_X1 U3459 ( .A(n3477), .B(n3478), .Z(n3407) );
  XOR2_X1 U3460 ( .A(n3479), .B(n3480), .Z(n3478) );
  OR2_X1 U3461 ( .A1(n2438), .A2(n2229), .ZN(n3410) );
  OR2_X1 U3462 ( .A1(n3414), .A2(n3411), .ZN(n3455) );
  XOR2_X1 U3463 ( .A(n3481), .B(n3482), .Z(n3411) );
  XOR2_X1 U3464 ( .A(n3483), .B(n3484), .Z(n3482) );
  OR2_X1 U3465 ( .A1(n2443), .A2(n2229), .ZN(n3414) );
  XOR2_X1 U3466 ( .A(n3485), .B(n3486), .Z(n3415) );
  XOR2_X1 U3467 ( .A(n3487), .B(n3488), .Z(n3486) );
  OR2_X1 U3468 ( .A1(n3422), .A2(n3419), .ZN(n3449) );
  XOR2_X1 U3469 ( .A(n3489), .B(n3490), .Z(n3419) );
  XOR2_X1 U3470 ( .A(n3491), .B(n3492), .Z(n3490) );
  OR2_X1 U3471 ( .A1(n2229), .A2(n2453), .ZN(n3422) );
  INV_X1 U3472 ( .A(n3313), .ZN(n2229) );
  XOR2_X1 U3473 ( .A(n3493), .B(n3494), .Z(n3313) );
  XNOR2_X1 U3474 ( .A(c_5_), .B(d_5_), .ZN(n3493) );
  XOR2_X1 U3475 ( .A(n3495), .B(n3496), .Z(n3425) );
  XOR2_X1 U3476 ( .A(n3497), .B(n3498), .Z(n3496) );
  XOR2_X1 U3477 ( .A(n3499), .B(n3500), .Z(n3429) );
  XOR2_X1 U3478 ( .A(n3501), .B(n3502), .Z(n3500) );
  XOR2_X1 U3479 ( .A(n3503), .B(n3504), .Z(n3433) );
  XOR2_X1 U3480 ( .A(n3505), .B(n3506), .Z(n3504) );
  XOR2_X1 U3481 ( .A(n3170), .B(n3507), .Z(n3163) );
  XOR2_X1 U3482 ( .A(n3169), .B(n3168), .Z(n3507) );
  OR2_X1 U3483 ( .A1(n2203), .A2(n2468), .ZN(n3168) );
  OR2_X1 U3484 ( .A1(n3508), .A2(n3509), .ZN(n3169) );
  AND2_X1 U3485 ( .A1(n3506), .A2(n3505), .ZN(n3509) );
  AND2_X1 U3486 ( .A1(n3503), .A2(n3510), .ZN(n3508) );
  OR2_X1 U3487 ( .A1(n3505), .A2(n3506), .ZN(n3510) );
  OR2_X1 U3488 ( .A1(n2203), .A2(n2463), .ZN(n3506) );
  OR2_X1 U3489 ( .A1(n3511), .A2(n3512), .ZN(n3505) );
  AND2_X1 U3490 ( .A1(n3502), .A2(n3501), .ZN(n3512) );
  AND2_X1 U3491 ( .A1(n3499), .A2(n3513), .ZN(n3511) );
  OR2_X1 U3492 ( .A1(n3501), .A2(n3502), .ZN(n3513) );
  OR2_X1 U3493 ( .A1(n2203), .A2(n2458), .ZN(n3502) );
  OR2_X1 U3494 ( .A1(n3514), .A2(n3515), .ZN(n3501) );
  AND2_X1 U3495 ( .A1(n3498), .A2(n3497), .ZN(n3515) );
  AND2_X1 U3496 ( .A1(n3495), .A2(n3516), .ZN(n3514) );
  OR2_X1 U3497 ( .A1(n3497), .A2(n3498), .ZN(n3516) );
  OR2_X1 U3498 ( .A1(n2203), .A2(n2453), .ZN(n3498) );
  OR2_X1 U3499 ( .A1(n3517), .A2(n3518), .ZN(n3497) );
  AND2_X1 U3500 ( .A1(n3489), .A2(n3492), .ZN(n3518) );
  AND2_X1 U3501 ( .A1(n3519), .A2(n3491), .ZN(n3517) );
  OR2_X1 U3502 ( .A1(n3520), .A2(n3521), .ZN(n3491) );
  AND2_X1 U3503 ( .A1(n3488), .A2(n3487), .ZN(n3521) );
  AND2_X1 U3504 ( .A1(n3485), .A2(n3522), .ZN(n3520) );
  OR2_X1 U3505 ( .A1(n3487), .A2(n3488), .ZN(n3522) );
  OR2_X1 U3506 ( .A1(n2203), .A2(n2443), .ZN(n3488) );
  OR2_X1 U3507 ( .A1(n3523), .A2(n3524), .ZN(n3487) );
  AND2_X1 U3508 ( .A1(n3481), .A2(n3484), .ZN(n3524) );
  AND2_X1 U3509 ( .A1(n3525), .A2(n3483), .ZN(n3523) );
  OR2_X1 U3510 ( .A1(n3526), .A2(n3527), .ZN(n3483) );
  AND2_X1 U3511 ( .A1(n3477), .A2(n3480), .ZN(n3527) );
  AND2_X1 U3512 ( .A1(n3528), .A2(n3479), .ZN(n3526) );
  OR2_X1 U3513 ( .A1(n3529), .A2(n3530), .ZN(n3479) );
  AND2_X1 U3514 ( .A1(n3474), .A2(n3476), .ZN(n3530) );
  AND2_X1 U3515 ( .A1(n3531), .A2(n3532), .ZN(n3529) );
  OR2_X1 U3516 ( .A1(n3476), .A2(n3474), .ZN(n3532) );
  OR2_X1 U3517 ( .A1(n2203), .A2(n2423), .ZN(n3474) );
  OR3_X1 U3518 ( .A1(n2176), .A2(n2203), .A3(n2424), .ZN(n3476) );
  INV_X1 U3519 ( .A(n3475), .ZN(n3531) );
  OR2_X1 U3520 ( .A1(n3533), .A2(n3534), .ZN(n3475) );
  AND2_X1 U3521 ( .A1(n3535), .A2(n3536), .ZN(n3534) );
  OR2_X1 U3522 ( .A1(n3537), .A2(n2035), .ZN(n3536) );
  AND2_X1 U3523 ( .A1(n2176), .A2(n2029), .ZN(n3537) );
  AND2_X1 U3524 ( .A1(n3468), .A2(n3538), .ZN(n3533) );
  OR2_X1 U3525 ( .A1(n3539), .A2(n2039), .ZN(n3538) );
  AND2_X1 U3526 ( .A1(n3540), .A2(n2041), .ZN(n3539) );
  OR2_X1 U3527 ( .A1(n3480), .A2(n3477), .ZN(n3528) );
  XOR2_X1 U3528 ( .A(n3541), .B(n3542), .Z(n3477) );
  XNOR2_X1 U3529 ( .A(n3543), .B(n3544), .ZN(n3541) );
  OR2_X1 U3530 ( .A1(n2433), .A2(n2203), .ZN(n3480) );
  OR2_X1 U3531 ( .A1(n3484), .A2(n3481), .ZN(n3525) );
  XOR2_X1 U3532 ( .A(n3545), .B(n3546), .Z(n3481) );
  XOR2_X1 U3533 ( .A(n3547), .B(n3548), .Z(n3546) );
  OR2_X1 U3534 ( .A1(n2438), .A2(n2203), .ZN(n3484) );
  XOR2_X1 U3535 ( .A(n3549), .B(n3550), .Z(n3485) );
  XOR2_X1 U3536 ( .A(n3551), .B(n3552), .Z(n3550) );
  OR2_X1 U3537 ( .A1(n3492), .A2(n3489), .ZN(n3519) );
  XOR2_X1 U3538 ( .A(n3553), .B(n3554), .Z(n3489) );
  XOR2_X1 U3539 ( .A(n3555), .B(n3556), .Z(n3554) );
  OR2_X1 U3540 ( .A1(n2203), .A2(n2448), .ZN(n3492) );
  INV_X1 U3541 ( .A(n3394), .ZN(n2203) );
  XOR2_X1 U3542 ( .A(n3557), .B(n3558), .Z(n3394) );
  XNOR2_X1 U3543 ( .A(c_4_), .B(d_4_), .ZN(n3557) );
  XOR2_X1 U3544 ( .A(n3559), .B(n3560), .Z(n3495) );
  XOR2_X1 U3545 ( .A(n3561), .B(n3562), .Z(n3560) );
  XOR2_X1 U3546 ( .A(n3563), .B(n3564), .Z(n3499) );
  XOR2_X1 U3547 ( .A(n3565), .B(n3566), .Z(n3564) );
  XOR2_X1 U3548 ( .A(n3567), .B(n3568), .Z(n3503) );
  XOR2_X1 U3549 ( .A(n3569), .B(n3570), .Z(n3568) );
  XOR2_X1 U3550 ( .A(n3177), .B(n3571), .Z(n3170) );
  XOR2_X1 U3551 ( .A(n3176), .B(n3175), .Z(n3571) );
  OR2_X1 U3552 ( .A1(n2176), .A2(n2463), .ZN(n3175) );
  OR2_X1 U3553 ( .A1(n3572), .A2(n3573), .ZN(n3176) );
  AND2_X1 U3554 ( .A1(n3570), .A2(n3569), .ZN(n3573) );
  AND2_X1 U3555 ( .A1(n3567), .A2(n3574), .ZN(n3572) );
  OR2_X1 U3556 ( .A1(n3569), .A2(n3570), .ZN(n3574) );
  OR2_X1 U3557 ( .A1(n2176), .A2(n2458), .ZN(n3570) );
  OR2_X1 U3558 ( .A1(n3575), .A2(n3576), .ZN(n3569) );
  AND2_X1 U3559 ( .A1(n3566), .A2(n3565), .ZN(n3576) );
  AND2_X1 U3560 ( .A1(n3563), .A2(n3577), .ZN(n3575) );
  OR2_X1 U3561 ( .A1(n3565), .A2(n3566), .ZN(n3577) );
  OR2_X1 U3562 ( .A1(n2176), .A2(n2453), .ZN(n3566) );
  OR2_X1 U3563 ( .A1(n3578), .A2(n3579), .ZN(n3565) );
  AND2_X1 U3564 ( .A1(n3562), .A2(n3561), .ZN(n3579) );
  AND2_X1 U3565 ( .A1(n3559), .A2(n3580), .ZN(n3578) );
  OR2_X1 U3566 ( .A1(n3561), .A2(n3562), .ZN(n3580) );
  OR2_X1 U3567 ( .A1(n2176), .A2(n2448), .ZN(n3562) );
  OR2_X1 U3568 ( .A1(n3581), .A2(n3582), .ZN(n3561) );
  AND2_X1 U3569 ( .A1(n3553), .A2(n3556), .ZN(n3582) );
  AND2_X1 U3570 ( .A1(n3583), .A2(n3555), .ZN(n3581) );
  OR2_X1 U3571 ( .A1(n3584), .A2(n3585), .ZN(n3555) );
  AND2_X1 U3572 ( .A1(n3552), .A2(n3551), .ZN(n3585) );
  AND2_X1 U3573 ( .A1(n3549), .A2(n3586), .ZN(n3584) );
  OR2_X1 U3574 ( .A1(n3551), .A2(n3552), .ZN(n3586) );
  OR2_X1 U3575 ( .A1(n2176), .A2(n2438), .ZN(n3552) );
  OR2_X1 U3576 ( .A1(n3587), .A2(n3588), .ZN(n3551) );
  AND2_X1 U3577 ( .A1(n3545), .A2(n3548), .ZN(n3588) );
  AND2_X1 U3578 ( .A1(n3589), .A2(n3547), .ZN(n3587) );
  OR2_X1 U3579 ( .A1(n3590), .A2(n3591), .ZN(n3547) );
  AND2_X1 U3580 ( .A1(n3542), .A2(n3544), .ZN(n3591) );
  AND2_X1 U3581 ( .A1(n3592), .A2(n3593), .ZN(n3590) );
  OR2_X1 U3582 ( .A1(n3544), .A2(n3542), .ZN(n3593) );
  OR2_X1 U3583 ( .A1(n2176), .A2(n2423), .ZN(n3542) );
  OR3_X1 U3584 ( .A1(n3540), .A2(n2176), .A3(n2424), .ZN(n3544) );
  INV_X1 U3585 ( .A(n3543), .ZN(n3592) );
  OR2_X1 U3586 ( .A1(n3594), .A2(n3595), .ZN(n3543) );
  AND2_X1 U3587 ( .A1(n3596), .A2(n3597), .ZN(n3595) );
  OR2_X1 U3588 ( .A1(n3598), .A2(n2035), .ZN(n3597) );
  AND2_X1 U3589 ( .A1(n3540), .A2(n2029), .ZN(n3598) );
  AND2_X1 U3590 ( .A1(n3535), .A2(n3599), .ZN(n3594) );
  OR2_X1 U3591 ( .A1(n3600), .A2(n2039), .ZN(n3599) );
  AND2_X1 U3592 ( .A1(n3601), .A2(n2041), .ZN(n3600) );
  OR2_X1 U3593 ( .A1(n3548), .A2(n3545), .ZN(n3589) );
  XOR2_X1 U3594 ( .A(n3602), .B(n3603), .Z(n3545) );
  XNOR2_X1 U3595 ( .A(n3604), .B(n3605), .ZN(n3602) );
  OR2_X1 U3596 ( .A1(n2433), .A2(n2176), .ZN(n3548) );
  XNOR2_X1 U3597 ( .A(n3606), .B(n3607), .ZN(n3549) );
  XNOR2_X1 U3598 ( .A(n3608), .B(n3609), .ZN(n3606) );
  OR2_X1 U3599 ( .A1(n3556), .A2(n3553), .ZN(n3583) );
  XOR2_X1 U3600 ( .A(n3610), .B(n3611), .Z(n3553) );
  XOR2_X1 U3601 ( .A(n3612), .B(n3613), .Z(n3611) );
  OR2_X1 U3602 ( .A1(n2176), .A2(n2443), .ZN(n3556) );
  INV_X1 U3603 ( .A(n3468), .ZN(n2176) );
  XOR2_X1 U3604 ( .A(n3614), .B(n3615), .Z(n3468) );
  XNOR2_X1 U3605 ( .A(c_3_), .B(d_3_), .ZN(n3614) );
  XOR2_X1 U3606 ( .A(n3616), .B(n3617), .Z(n3559) );
  XOR2_X1 U3607 ( .A(n3618), .B(n3619), .Z(n3617) );
  XOR2_X1 U3608 ( .A(n3620), .B(n3621), .Z(n3563) );
  XOR2_X1 U3609 ( .A(n3622), .B(n3623), .Z(n3621) );
  XOR2_X1 U3610 ( .A(n3624), .B(n3625), .Z(n3567) );
  XOR2_X1 U3611 ( .A(n3626), .B(n3627), .Z(n3625) );
  XOR2_X1 U3612 ( .A(n3628), .B(n3629), .Z(n3177) );
  XOR2_X1 U3613 ( .A(n3630), .B(n3631), .Z(n3629) );
  AND3_X1 U3614 ( .A1(n2091), .A2(n2089), .A3(n2090), .ZN(n2092) );
  INV_X1 U3615 ( .A(n2149), .ZN(n2090) );
  OR2_X1 U3616 ( .A1(n3632), .A2(n3633), .ZN(n2149) );
  AND2_X1 U3617 ( .A1(n2168), .A2(n2167), .ZN(n3633) );
  AND2_X1 U3618 ( .A1(n2165), .A2(n3634), .ZN(n3632) );
  OR2_X1 U3619 ( .A1(n2167), .A2(n2168), .ZN(n3634) );
  OR2_X1 U3620 ( .A1(n3540), .A2(n2148), .ZN(n2168) );
  OR2_X1 U3621 ( .A1(n3635), .A2(n3636), .ZN(n2167) );
  AND2_X1 U3622 ( .A1(n2186), .A2(n2185), .ZN(n3636) );
  AND2_X1 U3623 ( .A1(n2183), .A2(n3637), .ZN(n3635) );
  OR2_X1 U3624 ( .A1(n2185), .A2(n2186), .ZN(n3637) );
  OR2_X1 U3625 ( .A1(n3540), .A2(n2211), .ZN(n2186) );
  OR2_X1 U3626 ( .A1(n3638), .A2(n3639), .ZN(n2185) );
  AND2_X1 U3627 ( .A1(n2221), .A2(n2220), .ZN(n3639) );
  AND2_X1 U3628 ( .A1(n2218), .A2(n3640), .ZN(n3638) );
  OR2_X1 U3629 ( .A1(n2220), .A2(n2221), .ZN(n3640) );
  OR2_X1 U3630 ( .A1(n3540), .A2(n2244), .ZN(n2221) );
  OR2_X1 U3631 ( .A1(n3641), .A2(n3642), .ZN(n2220) );
  AND2_X1 U3632 ( .A1(n2254), .A2(n2253), .ZN(n3642) );
  AND2_X1 U3633 ( .A1(n2251), .A2(n3643), .ZN(n3641) );
  OR2_X1 U3634 ( .A1(n2253), .A2(n2254), .ZN(n3643) );
  OR2_X1 U3635 ( .A1(n3540), .A2(n2293), .ZN(n2254) );
  OR2_X1 U3636 ( .A1(n3644), .A2(n3645), .ZN(n2253) );
  AND2_X1 U3637 ( .A1(n2303), .A2(n2302), .ZN(n3645) );
  AND2_X1 U3638 ( .A1(n2300), .A2(n3646), .ZN(n3644) );
  OR2_X1 U3639 ( .A1(n2302), .A2(n2303), .ZN(n3646) );
  OR2_X1 U3640 ( .A1(n3540), .A2(n2340), .ZN(n2303) );
  OR2_X1 U3641 ( .A1(n3647), .A2(n3648), .ZN(n2302) );
  AND2_X1 U3642 ( .A1(n2350), .A2(n2349), .ZN(n3648) );
  AND2_X1 U3643 ( .A1(n2347), .A2(n3649), .ZN(n3647) );
  OR2_X1 U3644 ( .A1(n2349), .A2(n2350), .ZN(n3649) );
  OR2_X1 U3645 ( .A1(n3540), .A2(n2468), .ZN(n2350) );
  OR2_X1 U3646 ( .A1(n3650), .A2(n3651), .ZN(n2349) );
  AND2_X1 U3647 ( .A1(n3182), .A2(n3181), .ZN(n3651) );
  AND2_X1 U3648 ( .A1(n3179), .A2(n3652), .ZN(n3650) );
  OR2_X1 U3649 ( .A1(n3181), .A2(n3182), .ZN(n3652) );
  OR2_X1 U3650 ( .A1(n3540), .A2(n2463), .ZN(n3182) );
  OR2_X1 U3651 ( .A1(n3653), .A2(n3654), .ZN(n3181) );
  AND2_X1 U3652 ( .A1(n3631), .A2(n3630), .ZN(n3654) );
  AND2_X1 U3653 ( .A1(n3628), .A2(n3655), .ZN(n3653) );
  OR2_X1 U3654 ( .A1(n3630), .A2(n3631), .ZN(n3655) );
  OR2_X1 U3655 ( .A1(n3540), .A2(n2458), .ZN(n3631) );
  OR2_X1 U3656 ( .A1(n3656), .A2(n3657), .ZN(n3630) );
  AND2_X1 U3657 ( .A1(n3627), .A2(n3626), .ZN(n3657) );
  AND2_X1 U3658 ( .A1(n3624), .A2(n3658), .ZN(n3656) );
  OR2_X1 U3659 ( .A1(n3626), .A2(n3627), .ZN(n3658) );
  OR2_X1 U3660 ( .A1(n3540), .A2(n2453), .ZN(n3627) );
  OR2_X1 U3661 ( .A1(n3659), .A2(n3660), .ZN(n3626) );
  AND2_X1 U3662 ( .A1(n3623), .A2(n3622), .ZN(n3660) );
  AND2_X1 U3663 ( .A1(n3620), .A2(n3661), .ZN(n3659) );
  OR2_X1 U3664 ( .A1(n3622), .A2(n3623), .ZN(n3661) );
  OR2_X1 U3665 ( .A1(n3540), .A2(n2448), .ZN(n3623) );
  OR2_X1 U3666 ( .A1(n3662), .A2(n3663), .ZN(n3622) );
  AND2_X1 U3667 ( .A1(n3619), .A2(n3618), .ZN(n3663) );
  AND2_X1 U3668 ( .A1(n3616), .A2(n3664), .ZN(n3662) );
  OR2_X1 U3669 ( .A1(n3618), .A2(n3619), .ZN(n3664) );
  OR2_X1 U3670 ( .A1(n3540), .A2(n2443), .ZN(n3619) );
  OR2_X1 U3671 ( .A1(n3665), .A2(n3666), .ZN(n3618) );
  AND2_X1 U3672 ( .A1(n3610), .A2(n3613), .ZN(n3666) );
  AND2_X1 U3673 ( .A1(n3667), .A2(n3612), .ZN(n3665) );
  OR2_X1 U3674 ( .A1(n3668), .A2(n3669), .ZN(n3612) );
  AND2_X1 U3675 ( .A1(n3609), .A2(n3608), .ZN(n3669) );
  AND2_X1 U3676 ( .A1(n3607), .A2(n3670), .ZN(n3668) );
  OR2_X1 U3677 ( .A1(n3608), .A2(n3609), .ZN(n3670) );
  OR2_X1 U3678 ( .A1(n3540), .A2(n2433), .ZN(n3609) );
  OR2_X1 U3679 ( .A1(n3671), .A2(n3672), .ZN(n3608) );
  AND2_X1 U3680 ( .A1(n3603), .A2(n3605), .ZN(n3672) );
  AND2_X1 U3681 ( .A1(n3673), .A2(n3674), .ZN(n3671) );
  OR2_X1 U3682 ( .A1(n3605), .A2(n3603), .ZN(n3674) );
  OR2_X1 U3683 ( .A1(n3540), .A2(n2423), .ZN(n3603) );
  OR3_X1 U3684 ( .A1(n3601), .A2(n3540), .A3(n2424), .ZN(n3605) );
  OR2_X1 U3685 ( .A1(n3675), .A2(n3676), .ZN(n2424) );
  INV_X1 U3686 ( .A(n3604), .ZN(n3673) );
  OR2_X1 U3687 ( .A1(n3677), .A2(n3678), .ZN(n3604) );
  AND2_X1 U3688 ( .A1(n3679), .A2(n3680), .ZN(n3678) );
  OR2_X1 U3689 ( .A1(n3681), .A2(n2035), .ZN(n3680) );
  AND2_X1 U3690 ( .A1(n2029), .A2(n3675), .ZN(n2035) );
  AND2_X1 U3691 ( .A1(n3601), .A2(n2029), .ZN(n3681) );
  INV_X1 U3692 ( .A(n3682), .ZN(n3679) );
  AND2_X1 U3693 ( .A1(n3596), .A2(n3683), .ZN(n3677) );
  OR2_X1 U3694 ( .A1(n3684), .A2(n2039), .ZN(n3683) );
  AND2_X1 U3695 ( .A1(n3676), .A2(n2041), .ZN(n2039) );
  INV_X1 U3696 ( .A(n2029), .ZN(n3676) );
  AND2_X1 U3697 ( .A1(n3682), .A2(n2041), .ZN(n3684) );
  INV_X1 U3698 ( .A(n3675), .ZN(n2041) );
  XOR2_X1 U3699 ( .A(n3685), .B(n3686), .Z(n3607) );
  OR2_X1 U3700 ( .A1(n3687), .A2(n3688), .ZN(n3685) );
  AND2_X1 U3701 ( .A1(n3689), .A2(n3690), .ZN(n3687) );
  OR2_X1 U3702 ( .A1(n3601), .A2(n2423), .ZN(n3689) );
  OR2_X1 U3703 ( .A1(n3613), .A2(n3610), .ZN(n3667) );
  XOR2_X1 U3704 ( .A(n3691), .B(n3692), .Z(n3610) );
  XNOR2_X1 U3705 ( .A(n3693), .B(n3694), .ZN(n3691) );
  OR2_X1 U3706 ( .A1(n3540), .A2(n2438), .ZN(n3613) );
  INV_X1 U3707 ( .A(n3535), .ZN(n3540) );
  XOR2_X1 U3708 ( .A(n3695), .B(n3696), .Z(n3535) );
  XNOR2_X1 U3709 ( .A(c_2_), .B(d_2_), .ZN(n3695) );
  XNOR2_X1 U3710 ( .A(n3697), .B(n3698), .ZN(n3616) );
  XNOR2_X1 U3711 ( .A(n3699), .B(n3700), .ZN(n3697) );
  XNOR2_X1 U3712 ( .A(n3701), .B(n3702), .ZN(n3620) );
  XNOR2_X1 U3713 ( .A(n3703), .B(n3704), .ZN(n3701) );
  XNOR2_X1 U3714 ( .A(n3705), .B(n3706), .ZN(n3624) );
  XNOR2_X1 U3715 ( .A(n3707), .B(n3708), .ZN(n3705) );
  XOR2_X1 U3716 ( .A(n3709), .B(n3710), .Z(n3628) );
  XOR2_X1 U3717 ( .A(n3711), .B(n3712), .Z(n3710) );
  XOR2_X1 U3718 ( .A(n3713), .B(n3714), .Z(n3179) );
  XOR2_X1 U3719 ( .A(n3715), .B(n3716), .Z(n3714) );
  XOR2_X1 U3720 ( .A(n3717), .B(n3718), .Z(n2347) );
  XOR2_X1 U3721 ( .A(n3719), .B(n3720), .Z(n3718) );
  XOR2_X1 U3722 ( .A(n3721), .B(n3722), .Z(n2300) );
  XOR2_X1 U3723 ( .A(n3723), .B(n3724), .Z(n3722) );
  XOR2_X1 U3724 ( .A(n3725), .B(n3726), .Z(n2251) );
  XOR2_X1 U3725 ( .A(n3727), .B(n3728), .Z(n3726) );
  XOR2_X1 U3726 ( .A(n3729), .B(n3730), .Z(n2218) );
  XOR2_X1 U3727 ( .A(n3731), .B(n3732), .Z(n3730) );
  XOR2_X1 U3728 ( .A(n3733), .B(n3734), .Z(n2183) );
  XOR2_X1 U3729 ( .A(n3735), .B(n3736), .Z(n3734) );
  XOR2_X1 U3730 ( .A(n3737), .B(n3738), .Z(n2165) );
  XOR2_X1 U3731 ( .A(n3739), .B(n3740), .Z(n3738) );
  XOR2_X1 U3732 ( .A(n3741), .B(n2147), .Z(n2089) );
  OR2_X1 U3733 ( .A1(n3742), .A2(n3743), .ZN(n2147) );
  AND2_X1 U3734 ( .A1(n3744), .A2(n3745), .ZN(n3743) );
  AND2_X1 U3735 ( .A1(n3746), .A2(n3747), .ZN(n3742) );
  OR2_X1 U3736 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  OR2_X1 U3737 ( .A1(n2148), .A2(n3682), .ZN(n3741) );
  XNOR2_X1 U3738 ( .A(n3744), .B(n3748), .ZN(n2091) );
  XOR2_X1 U3739 ( .A(n3745), .B(n3747), .Z(n3748) );
  OR2_X1 U3740 ( .A1(n2211), .A2(n3682), .ZN(n3747) );
  OR2_X1 U3741 ( .A1(n3749), .A2(n3750), .ZN(n3745) );
  AND2_X1 U3742 ( .A1(n3737), .A2(n3739), .ZN(n3750) );
  AND2_X1 U3743 ( .A1(n3751), .A2(n3740), .ZN(n3749) );
  OR2_X1 U3744 ( .A1(n3601), .A2(n2211), .ZN(n3740) );
  XNOR2_X1 U3745 ( .A(n3752), .B(n3753), .ZN(n2211) );
  XNOR2_X1 U3746 ( .A(a_1_), .B(b_1_), .ZN(n3752) );
  OR2_X1 U3747 ( .A1(n3739), .A2(n3737), .ZN(n3751) );
  OR2_X1 U3748 ( .A1(n2244), .A2(n3682), .ZN(n3737) );
  OR2_X1 U3749 ( .A1(n3754), .A2(n3755), .ZN(n3739) );
  AND2_X1 U3750 ( .A1(n3733), .A2(n3735), .ZN(n3755) );
  AND2_X1 U3751 ( .A1(n3756), .A2(n3736), .ZN(n3754) );
  OR2_X1 U3752 ( .A1(n2293), .A2(n3682), .ZN(n3736) );
  OR2_X1 U3753 ( .A1(n3735), .A2(n3733), .ZN(n3756) );
  OR2_X1 U3754 ( .A1(n3601), .A2(n2244), .ZN(n3733) );
  XNOR2_X1 U3755 ( .A(n3757), .B(n3758), .ZN(n2244) );
  XNOR2_X1 U3756 ( .A(a_2_), .B(b_2_), .ZN(n3757) );
  OR2_X1 U3757 ( .A1(n3759), .A2(n3760), .ZN(n3735) );
  AND2_X1 U3758 ( .A1(n3729), .A2(n3731), .ZN(n3760) );
  AND2_X1 U3759 ( .A1(n3761), .A2(n3732), .ZN(n3759) );
  OR2_X1 U3760 ( .A1(n2340), .A2(n3682), .ZN(n3732) );
  OR2_X1 U3761 ( .A1(n3731), .A2(n3729), .ZN(n3761) );
  OR2_X1 U3762 ( .A1(n3601), .A2(n2293), .ZN(n3729) );
  XNOR2_X1 U3763 ( .A(n3762), .B(n3763), .ZN(n2293) );
  XNOR2_X1 U3764 ( .A(a_3_), .B(b_3_), .ZN(n3762) );
  OR2_X1 U3765 ( .A1(n3764), .A2(n3765), .ZN(n3731) );
  AND2_X1 U3766 ( .A1(n3725), .A2(n3727), .ZN(n3765) );
  AND2_X1 U3767 ( .A1(n3766), .A2(n3728), .ZN(n3764) );
  OR2_X1 U3768 ( .A1(n2468), .A2(n3682), .ZN(n3728) );
  OR2_X1 U3769 ( .A1(n3727), .A2(n3725), .ZN(n3766) );
  OR2_X1 U3770 ( .A1(n3601), .A2(n2340), .ZN(n3725) );
  XNOR2_X1 U3771 ( .A(n3767), .B(n3768), .ZN(n2340) );
  XNOR2_X1 U3772 ( .A(a_4_), .B(b_4_), .ZN(n3767) );
  OR2_X1 U3773 ( .A1(n3769), .A2(n3770), .ZN(n3727) );
  AND2_X1 U3774 ( .A1(n3721), .A2(n3723), .ZN(n3770) );
  AND2_X1 U3775 ( .A1(n3771), .A2(n3724), .ZN(n3769) );
  OR2_X1 U3776 ( .A1(n2463), .A2(n3682), .ZN(n3724) );
  OR2_X1 U3777 ( .A1(n3723), .A2(n3721), .ZN(n3771) );
  OR2_X1 U3778 ( .A1(n3601), .A2(n2468), .ZN(n3721) );
  XNOR2_X1 U3779 ( .A(n3772), .B(n3773), .ZN(n2468) );
  XNOR2_X1 U3780 ( .A(a_5_), .B(b_5_), .ZN(n3772) );
  OR2_X1 U3781 ( .A1(n3774), .A2(n3775), .ZN(n3723) );
  AND2_X1 U3782 ( .A1(n3717), .A2(n3719), .ZN(n3775) );
  AND2_X1 U3783 ( .A1(n3776), .A2(n3720), .ZN(n3774) );
  OR2_X1 U3784 ( .A1(n2458), .A2(n3682), .ZN(n3720) );
  OR2_X1 U3785 ( .A1(n3719), .A2(n3717), .ZN(n3776) );
  OR2_X1 U3786 ( .A1(n3601), .A2(n2463), .ZN(n3717) );
  XNOR2_X1 U3787 ( .A(n3777), .B(n3778), .ZN(n2463) );
  XNOR2_X1 U3788 ( .A(a_6_), .B(b_6_), .ZN(n3777) );
  OR2_X1 U3789 ( .A1(n3779), .A2(n3780), .ZN(n3719) );
  AND2_X1 U3790 ( .A1(n3713), .A2(n3715), .ZN(n3780) );
  AND2_X1 U3791 ( .A1(n3781), .A2(n3716), .ZN(n3779) );
  OR2_X1 U3792 ( .A1(n2453), .A2(n3682), .ZN(n3716) );
  OR2_X1 U3793 ( .A1(n3715), .A2(n3713), .ZN(n3781) );
  OR2_X1 U3794 ( .A1(n3601), .A2(n2458), .ZN(n3713) );
  XNOR2_X1 U3795 ( .A(n3782), .B(n3783), .ZN(n2458) );
  XNOR2_X1 U3796 ( .A(a_7_), .B(b_7_), .ZN(n3782) );
  OR2_X1 U3797 ( .A1(n3784), .A2(n3785), .ZN(n3715) );
  AND2_X1 U3798 ( .A1(n3709), .A2(n3711), .ZN(n3785) );
  AND2_X1 U3799 ( .A1(n3786), .A2(n3712), .ZN(n3784) );
  OR2_X1 U3800 ( .A1(n2448), .A2(n3682), .ZN(n3712) );
  OR2_X1 U3801 ( .A1(n3711), .A2(n3709), .ZN(n3786) );
  OR2_X1 U3802 ( .A1(n3601), .A2(n2453), .ZN(n3709) );
  XNOR2_X1 U3803 ( .A(n3787), .B(n3788), .ZN(n2453) );
  XNOR2_X1 U3804 ( .A(a_8_), .B(b_8_), .ZN(n3787) );
  OR2_X1 U3805 ( .A1(n3789), .A2(n3790), .ZN(n3711) );
  AND2_X1 U3806 ( .A1(n3706), .A2(n3708), .ZN(n3790) );
  AND2_X1 U3807 ( .A1(n3791), .A2(n3707), .ZN(n3789) );
  OR2_X1 U3808 ( .A1(n2443), .A2(n3682), .ZN(n3707) );
  OR2_X1 U3809 ( .A1(n3708), .A2(n3706), .ZN(n3791) );
  OR2_X1 U3810 ( .A1(n3601), .A2(n2448), .ZN(n3706) );
  XNOR2_X1 U3811 ( .A(n3792), .B(n3793), .ZN(n2448) );
  XNOR2_X1 U3812 ( .A(a_9_), .B(b_9_), .ZN(n3792) );
  OR2_X1 U3813 ( .A1(n3794), .A2(n3795), .ZN(n3708) );
  AND2_X1 U3814 ( .A1(n3702), .A2(n3704), .ZN(n3795) );
  AND2_X1 U3815 ( .A1(n3796), .A2(n3703), .ZN(n3794) );
  OR2_X1 U3816 ( .A1(n2438), .A2(n3682), .ZN(n3703) );
  OR2_X1 U3817 ( .A1(n3704), .A2(n3702), .ZN(n3796) );
  OR2_X1 U3818 ( .A1(n3601), .A2(n2443), .ZN(n3702) );
  XNOR2_X1 U3819 ( .A(n3797), .B(n3798), .ZN(n2443) );
  XNOR2_X1 U3820 ( .A(a_10_), .B(b_10_), .ZN(n3797) );
  OR2_X1 U3821 ( .A1(n3799), .A2(n3800), .ZN(n3704) );
  AND2_X1 U3822 ( .A1(n3698), .A2(n3700), .ZN(n3800) );
  AND2_X1 U3823 ( .A1(n3801), .A2(n3699), .ZN(n3799) );
  OR2_X1 U3824 ( .A1(n2433), .A2(n3682), .ZN(n3699) );
  OR2_X1 U3825 ( .A1(n3700), .A2(n3698), .ZN(n3801) );
  OR2_X1 U3826 ( .A1(n3601), .A2(n2438), .ZN(n3698) );
  XNOR2_X1 U3827 ( .A(n3802), .B(n3803), .ZN(n2438) );
  XNOR2_X1 U3828 ( .A(a_11_), .B(b_11_), .ZN(n3802) );
  OR2_X1 U3829 ( .A1(n3804), .A2(n3805), .ZN(n3700) );
  AND2_X1 U3830 ( .A1(n3692), .A2(n3694), .ZN(n3805) );
  AND2_X1 U3831 ( .A1(n3806), .A2(n3807), .ZN(n3804) );
  OR2_X1 U3832 ( .A1(n3694), .A2(n3692), .ZN(n3807) );
  OR2_X1 U3833 ( .A1(n3601), .A2(n2433), .ZN(n3692) );
  XNOR2_X1 U3834 ( .A(n3808), .B(n3809), .ZN(n2433) );
  XNOR2_X1 U3835 ( .A(a_12_), .B(b_12_), .ZN(n3808) );
  OR2_X1 U3836 ( .A1(n2423), .A2(n3682), .ZN(n3694) );
  INV_X1 U3837 ( .A(n3693), .ZN(n3806) );
  OR2_X1 U3838 ( .A1(n3688), .A2(n3686), .ZN(n3693) );
  AND3_X1 U3839 ( .A1(n3596), .A2(n2029), .A3(n3810), .ZN(n3686) );
  AND2_X1 U3840 ( .A1(n3811), .A2(n3812), .ZN(n2029) );
  OR2_X1 U3841 ( .A1(b_15_), .A2(a_15_), .ZN(n3812) );
  INV_X1 U3842 ( .A(n3813), .ZN(n3811) );
  AND3_X1 U3843 ( .A1(n3596), .A2(n3814), .A3(n3810), .ZN(n3688) );
  INV_X1 U3844 ( .A(n3690), .ZN(n3810) );
  OR2_X1 U3845 ( .A1(n3675), .A2(n3682), .ZN(n3690) );
  XOR2_X1 U3846 ( .A(d_0_), .B(c_0_), .Z(n3816) );
  OR2_X1 U3847 ( .A1(n3817), .A2(n3818), .ZN(n3815) );
  AND2_X1 U3848 ( .A1(n3819), .A2(c_1_), .ZN(n3818) );
  AND2_X1 U3849 ( .A1(d_1_), .A2(n3820), .ZN(n3817) );
  OR2_X1 U3850 ( .A1(n3819), .A2(c_1_), .ZN(n3820) );
  INV_X1 U3851 ( .A(n3821), .ZN(n3819) );
  XNOR2_X1 U3852 ( .A(n3813), .B(n3822), .ZN(n3675) );
  XOR2_X1 U3853 ( .A(b_14_), .B(a_14_), .Z(n3822) );
  INV_X1 U3854 ( .A(n2423), .ZN(n3814) );
  XNOR2_X1 U3855 ( .A(n3825), .B(a_13_), .ZN(n3824) );
  OR2_X1 U3856 ( .A1(n3601), .A2(n2148), .ZN(n3744) );
  XOR2_X1 U3857 ( .A(b_0_), .B(a_0_), .Z(n3827) );
  OR2_X1 U3858 ( .A1(n3828), .A2(n3829), .ZN(n3826) );
  AND2_X1 U3859 ( .A1(n3830), .A2(a_1_), .ZN(n3829) );
  AND2_X1 U3860 ( .A1(b_1_), .A2(n3831), .ZN(n3828) );
  OR2_X1 U3861 ( .A1(n3830), .A2(a_1_), .ZN(n3831) );
  INV_X1 U3862 ( .A(n3753), .ZN(n3830) );
  OR2_X1 U3863 ( .A1(n3832), .A2(n3833), .ZN(n3753) );
  AND2_X1 U3864 ( .A1(n3758), .A2(n3834), .ZN(n3833) );
  AND2_X1 U3865 ( .A1(n3835), .A2(n3836), .ZN(n3832) );
  INV_X1 U3866 ( .A(b_2_), .ZN(n3836) );
  OR2_X1 U3867 ( .A1(n3834), .A2(n3758), .ZN(n3835) );
  OR2_X1 U3868 ( .A1(n3837), .A2(n3838), .ZN(n3758) );
  AND2_X1 U3869 ( .A1(n3763), .A2(n3839), .ZN(n3838) );
  AND2_X1 U3870 ( .A1(n3840), .A2(n3841), .ZN(n3837) );
  INV_X1 U3871 ( .A(b_3_), .ZN(n3841) );
  OR2_X1 U3872 ( .A1(n3839), .A2(n3763), .ZN(n3840) );
  OR2_X1 U3873 ( .A1(n3842), .A2(n3843), .ZN(n3763) );
  AND2_X1 U3874 ( .A1(n3768), .A2(n3844), .ZN(n3843) );
  AND2_X1 U3875 ( .A1(n3845), .A2(n3846), .ZN(n3842) );
  INV_X1 U3876 ( .A(b_4_), .ZN(n3846) );
  OR2_X1 U3877 ( .A1(n3844), .A2(n3768), .ZN(n3845) );
  OR2_X1 U3878 ( .A1(n3847), .A2(n3848), .ZN(n3768) );
  AND2_X1 U3879 ( .A1(n3773), .A2(n3849), .ZN(n3848) );
  AND2_X1 U3880 ( .A1(n3850), .A2(n3851), .ZN(n3847) );
  INV_X1 U3881 ( .A(b_5_), .ZN(n3851) );
  OR2_X1 U3882 ( .A1(n3849), .A2(n3773), .ZN(n3850) );
  OR2_X1 U3883 ( .A1(n3852), .A2(n3853), .ZN(n3773) );
  AND2_X1 U3884 ( .A1(n3778), .A2(n3854), .ZN(n3853) );
  AND2_X1 U3885 ( .A1(n3855), .A2(n3856), .ZN(n3852) );
  INV_X1 U3886 ( .A(b_6_), .ZN(n3856) );
  OR2_X1 U3887 ( .A1(n3854), .A2(n3778), .ZN(n3855) );
  OR2_X1 U3888 ( .A1(n3857), .A2(n3858), .ZN(n3778) );
  AND2_X1 U3889 ( .A1(n3783), .A2(n3859), .ZN(n3858) );
  AND2_X1 U3890 ( .A1(n3860), .A2(n3861), .ZN(n3857) );
  INV_X1 U3891 ( .A(b_7_), .ZN(n3861) );
  OR2_X1 U3892 ( .A1(n3859), .A2(n3783), .ZN(n3860) );
  OR2_X1 U3893 ( .A1(n3862), .A2(n3863), .ZN(n3783) );
  AND2_X1 U3894 ( .A1(n3788), .A2(n3864), .ZN(n3863) );
  AND2_X1 U3895 ( .A1(n3865), .A2(n3866), .ZN(n3862) );
  INV_X1 U3896 ( .A(b_8_), .ZN(n3866) );
  OR2_X1 U3897 ( .A1(n3864), .A2(n3788), .ZN(n3865) );
  OR2_X1 U3898 ( .A1(n3867), .A2(n3868), .ZN(n3788) );
  AND2_X1 U3899 ( .A1(n3793), .A2(n3869), .ZN(n3868) );
  AND2_X1 U3900 ( .A1(n3870), .A2(n3871), .ZN(n3867) );
  INV_X1 U3901 ( .A(b_9_), .ZN(n3871) );
  OR2_X1 U3902 ( .A1(n3869), .A2(n3793), .ZN(n3870) );
  OR2_X1 U3903 ( .A1(n3872), .A2(n3873), .ZN(n3793) );
  AND2_X1 U3904 ( .A1(n3798), .A2(n3874), .ZN(n3873) );
  AND2_X1 U3905 ( .A1(n3875), .A2(n3876), .ZN(n3872) );
  INV_X1 U3906 ( .A(b_10_), .ZN(n3876) );
  OR2_X1 U3907 ( .A1(n3874), .A2(n3798), .ZN(n3875) );
  OR2_X1 U3908 ( .A1(n3877), .A2(n3878), .ZN(n3798) );
  AND2_X1 U3909 ( .A1(n3803), .A2(n3879), .ZN(n3878) );
  AND2_X1 U3910 ( .A1(n3880), .A2(n3881), .ZN(n3877) );
  INV_X1 U3911 ( .A(b_11_), .ZN(n3881) );
  OR2_X1 U3912 ( .A1(n3879), .A2(n3803), .ZN(n3880) );
  OR2_X1 U3913 ( .A1(n3882), .A2(n3883), .ZN(n3803) );
  AND2_X1 U3914 ( .A1(n3809), .A2(n3884), .ZN(n3883) );
  AND2_X1 U3915 ( .A1(n3885), .A2(n3886), .ZN(n3882) );
  INV_X1 U3916 ( .A(b_12_), .ZN(n3886) );
  OR2_X1 U3917 ( .A1(n3884), .A2(n3809), .ZN(n3885) );
  OR2_X1 U3918 ( .A1(n3887), .A2(n3888), .ZN(n3809) );
  AND2_X1 U3919 ( .A1(n3889), .A2(n3890), .ZN(n3888) );
  AND2_X1 U3920 ( .A1(n3891), .A2(n3825), .ZN(n3887) );
  INV_X1 U3921 ( .A(b_13_), .ZN(n3825) );
  OR2_X1 U3922 ( .A1(n3889), .A2(n3890), .ZN(n3891) );
  INV_X1 U3923 ( .A(a_13_), .ZN(n3890) );
  INV_X1 U3924 ( .A(n3823), .ZN(n3889) );
  OR2_X1 U3925 ( .A1(n3892), .A2(n3893), .ZN(n3823) );
  AND2_X1 U3926 ( .A1(n3813), .A2(a_14_), .ZN(n3893) );
  AND2_X1 U3927 ( .A1(b_14_), .A2(n3894), .ZN(n3892) );
  OR2_X1 U3928 ( .A1(n3813), .A2(a_14_), .ZN(n3894) );
  AND2_X1 U3929 ( .A1(a_15_), .A2(b_15_), .ZN(n3813) );
  INV_X1 U3930 ( .A(a_12_), .ZN(n3884) );
  INV_X1 U3931 ( .A(a_11_), .ZN(n3879) );
  INV_X1 U3932 ( .A(a_10_), .ZN(n3874) );
  INV_X1 U3933 ( .A(a_9_), .ZN(n3869) );
  INV_X1 U3934 ( .A(a_8_), .ZN(n3864) );
  INV_X1 U3935 ( .A(a_7_), .ZN(n3859) );
  INV_X1 U3936 ( .A(a_6_), .ZN(n3854) );
  INV_X1 U3937 ( .A(a_5_), .ZN(n3849) );
  INV_X1 U3938 ( .A(a_4_), .ZN(n3844) );
  INV_X1 U3939 ( .A(a_3_), .ZN(n3839) );
  INV_X1 U3940 ( .A(a_2_), .ZN(n3834) );
  INV_X1 U3941 ( .A(n3596), .ZN(n3601) );
  XOR2_X1 U3942 ( .A(n3895), .B(n3821), .Z(n3596) );
  OR2_X1 U3943 ( .A1(n3896), .A2(n3897), .ZN(n3821) );
  AND2_X1 U3944 ( .A1(n3696), .A2(n3898), .ZN(n3897) );
  AND2_X1 U3945 ( .A1(n3899), .A2(n3900), .ZN(n3896) );
  INV_X1 U3946 ( .A(d_2_), .ZN(n3900) );
  OR2_X1 U3947 ( .A1(n3898), .A2(n3696), .ZN(n3899) );
  OR2_X1 U3948 ( .A1(n3901), .A2(n3902), .ZN(n3696) );
  AND2_X1 U3949 ( .A1(n3615), .A2(n3903), .ZN(n3902) );
  AND2_X1 U3950 ( .A1(n3904), .A2(n3905), .ZN(n3901) );
  INV_X1 U3951 ( .A(d_3_), .ZN(n3905) );
  OR2_X1 U3952 ( .A1(n3903), .A2(n3615), .ZN(n3904) );
  OR2_X1 U3953 ( .A1(n3906), .A2(n3907), .ZN(n3615) );
  AND2_X1 U3954 ( .A1(n3558), .A2(n3908), .ZN(n3907) );
  AND2_X1 U3955 ( .A1(n3909), .A2(n3910), .ZN(n3906) );
  INV_X1 U3956 ( .A(d_4_), .ZN(n3910) );
  OR2_X1 U3957 ( .A1(n3908), .A2(n3558), .ZN(n3909) );
  OR2_X1 U3958 ( .A1(n3911), .A2(n3912), .ZN(n3558) );
  AND2_X1 U3959 ( .A1(n3494), .A2(n3913), .ZN(n3912) );
  AND2_X1 U3960 ( .A1(n3914), .A2(n3915), .ZN(n3911) );
  INV_X1 U3961 ( .A(d_5_), .ZN(n3915) );
  OR2_X1 U3962 ( .A1(n3913), .A2(n3494), .ZN(n3914) );
  OR2_X1 U3963 ( .A1(n3916), .A2(n3917), .ZN(n3494) );
  AND2_X1 U3964 ( .A1(n3424), .A2(n3918), .ZN(n3917) );
  AND2_X1 U3965 ( .A1(n3919), .A2(n3920), .ZN(n3916) );
  INV_X1 U3966 ( .A(d_6_), .ZN(n3920) );
  OR2_X1 U3967 ( .A1(n3918), .A2(n3424), .ZN(n3919) );
  OR2_X1 U3968 ( .A1(n3921), .A2(n3922), .ZN(n3424) );
  AND2_X1 U3969 ( .A1(n3347), .A2(n3923), .ZN(n3922) );
  AND2_X1 U3970 ( .A1(n3924), .A2(n3925), .ZN(n3921) );
  INV_X1 U3971 ( .A(d_7_), .ZN(n3925) );
  OR2_X1 U3972 ( .A1(n3923), .A2(n3347), .ZN(n3924) );
  OR2_X1 U3973 ( .A1(n3926), .A2(n3927), .ZN(n3347) );
  AND2_X1 U3974 ( .A1(n3263), .A2(n3928), .ZN(n3927) );
  AND2_X1 U3975 ( .A1(n3929), .A2(n3930), .ZN(n3926) );
  INV_X1 U3976 ( .A(d_8_), .ZN(n3930) );
  OR2_X1 U3977 ( .A1(n3928), .A2(n3263), .ZN(n3929) );
  OR2_X1 U3978 ( .A1(n3931), .A2(n3932), .ZN(n3263) );
  AND2_X1 U3979 ( .A1(n3126), .A2(n3933), .ZN(n3932) );
  AND2_X1 U3980 ( .A1(n3934), .A2(n3935), .ZN(n3931) );
  INV_X1 U3981 ( .A(d_9_), .ZN(n3935) );
  OR2_X1 U3982 ( .A1(n3933), .A2(n3126), .ZN(n3934) );
  OR2_X1 U3983 ( .A1(n3936), .A2(n3937), .ZN(n3126) );
  AND2_X1 U3984 ( .A1(n3018), .A2(n3938), .ZN(n3937) );
  AND2_X1 U3985 ( .A1(n3939), .A2(n3940), .ZN(n3936) );
  INV_X1 U3986 ( .A(d_10_), .ZN(n3940) );
  OR2_X1 U3987 ( .A1(n3938), .A2(n3018), .ZN(n3939) );
  OR2_X1 U3988 ( .A1(n3941), .A2(n3942), .ZN(n3018) );
  AND2_X1 U3989 ( .A1(n2861), .A2(n3943), .ZN(n3942) );
  AND2_X1 U3990 ( .A1(n3944), .A2(n3945), .ZN(n3941) );
  INV_X1 U3991 ( .A(d_11_), .ZN(n3945) );
  OR2_X1 U3992 ( .A1(n3943), .A2(n2861), .ZN(n3944) );
  OR2_X1 U3993 ( .A1(n3946), .A2(n3947), .ZN(n2861) );
  AND2_X1 U3994 ( .A1(n2752), .A2(n3948), .ZN(n3947) );
  AND2_X1 U3995 ( .A1(n3949), .A2(n3950), .ZN(n3946) );
  INV_X1 U3996 ( .A(d_12_), .ZN(n3950) );
  OR2_X1 U3997 ( .A1(n3948), .A2(n2752), .ZN(n3949) );
  OR2_X1 U3998 ( .A1(n3951), .A2(n3952), .ZN(n2752) );
  AND2_X1 U3999 ( .A1(n2649), .A2(n3953), .ZN(n3952) );
  AND2_X1 U4000 ( .A1(n3954), .A2(n2651), .ZN(n3951) );
  INV_X1 U4001 ( .A(d_13_), .ZN(n2651) );
  OR2_X1 U4002 ( .A1(n2649), .A2(n3953), .ZN(n3954) );
  INV_X1 U4003 ( .A(c_13_), .ZN(n3953) );
  INV_X1 U4004 ( .A(n3955), .ZN(n2649) );
  OR2_X1 U4005 ( .A1(n3956), .A2(n3957), .ZN(n3955) );
  AND2_X1 U4006 ( .A1(c_14_), .A2(n2491), .ZN(n3957) );
  AND2_X1 U4007 ( .A1(d_14_), .A2(n3958), .ZN(n3956) );
  OR2_X1 U4008 ( .A1(n2491), .A2(c_14_), .ZN(n3958) );
  AND2_X1 U4009 ( .A1(c_15_), .A2(d_15_), .ZN(n2491) );
  INV_X1 U4010 ( .A(c_12_), .ZN(n3948) );
  INV_X1 U4011 ( .A(c_11_), .ZN(n3943) );
  INV_X1 U4012 ( .A(c_10_), .ZN(n3938) );
  INV_X1 U4013 ( .A(c_9_), .ZN(n3933) );
  INV_X1 U4014 ( .A(c_8_), .ZN(n3928) );
  INV_X1 U4015 ( .A(c_7_), .ZN(n3923) );
  INV_X1 U4016 ( .A(c_6_), .ZN(n3918) );
  INV_X1 U4017 ( .A(c_5_), .ZN(n3913) );
  INV_X1 U4018 ( .A(c_4_), .ZN(n3908) );
  INV_X1 U4019 ( .A(c_3_), .ZN(n3903) );
  INV_X1 U4020 ( .A(c_2_), .ZN(n3898) );
  XNOR2_X1 U4021 ( .A(c_1_), .B(d_1_), .ZN(n3895) );
endmodule

