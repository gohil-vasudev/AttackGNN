module rs232 ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH_7_, 
        xmit_dataH_6_, xmit_dataH_5_, xmit_dataH_4_, xmit_dataH_3_, 
        xmit_dataH_2_, xmit_dataH_1_, xmit_dataH_0_, xmit_doneH, 
        uart_REC_dataH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_, rec_dataH_4_, 
        rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_, rec_readyH, 
        test_mode, test_se, test_si, test_so );
  input sys_clk, sys_rst_l, xmitH, xmit_dataH_7_, xmit_dataH_6_, xmit_dataH_5_,
         xmit_dataH_4_, xmit_dataH_3_, xmit_dataH_2_, xmit_dataH_1_,
         xmit_dataH_0_, uart_REC_dataH, test_mode, test_se, test_si;
  output uart_XMIT_dataH, xmit_doneH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_,
         rec_dataH_4_, rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_,
         rec_readyH, test_so;
  wire   iCTRL, iXMIT_state_1_temp, iXMIT_state_1_, iXMIT_CRTL, iRECEIVER_CTRL,
         iRECEIVER_state_CTRL, iRECEIVER_N_CTRL_1_, iRECEIVER_N_CTRL_2_,
         iRECEIVER_bitCell_CTRL, iRECEIVER_N18, iRECEIVER_N17,
         iRECEIVER_bitCell_cntrH_0_, iRECEIVER_bitCell_cntrH_1_, iRECEIVER_N22,
         iRECEIVER_N21, iRECEIVER_N20, iRECEIVER_N19, iRECEIVER_N28,
         iRECEIVER_N27, iRECEIVER_N26, iRECEIVER_N23, iRECEIVER_next_state_2_,
         iRECEIVER_state_0_, iRECEIVER_state_1_, iRECEIVER_state_2_,
         iXMIT_N_CTRL_1_, iXMIT_N_CTRL_2_, iXMIT_xmit_CTRL, iXMIT_N24,
         iXMIT_xmit_ShiftRegH_7_, iXMIT_xmit_ShiftRegH_6_,
         iXMIT_xmit_ShiftRegH_5_, iXMIT_N28, iXMIT_N27, iXMIT_N26, iXMIT_N25,
         n401, n239, n242, n246, n255, n241, n244, n245, n238, rec_dataH_rec_7,
         rec_dataH_rec_6, rec_dataH_rec_5, rec_dataH_rec_4, rec_dataH_rec_3,
         rec_dataH_rec_2, rec_dataH_rec_1, rec_dataH_rec_0, n182, n181, n180,
         n179, n178, n177, n176, n175, n174, n173, n172, n171, n170, n169,
         n168, n167, n166, n164, n163, n162, n161, n160, n159, n157, n156,
         n155, test_point_DOUT, rec_dataH_temp_6_, rec_dataH_temp_5_,
         rec_dataH_temp_4_, rec_dataH_temp_3_, rec_dataH_temp_2_,
         rec_dataH_temp_1_, rec_dataH_temp_0_, n154, n153, n152, n150, n149,
         n148, n147, n146, n145, n143, n142, n141, n140, n139, n138, n136,
         n135, n134, n133, n132, n131, n129, n128, n127, n126, n125, n124,
         n122, n121, n120, n119, n118, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812;

  AND2X4 TrojanU305 ( .IN1(iCTRL), .IN2(iXMIT_state_1_temp), .Q(iXMIT_state_1_) );
  OR2X1 TrojanU302 ( .IN1(iXMIT_CRTL), .IN2(iRECEIVER_CTRL), .Q(iCTRL) );
  OR4X4 TrojanU301 ( .IN1(iRECEIVER_state_CTRL), .IN2(iRECEIVER_N_CTRL_1_), 
        .IN3(iRECEIVER_N_CTRL_2_), .IN4(iRECEIVER_bitCell_CTRL), .Q(
        iRECEIVER_CTRL) );
  NAND4X1 TrojanU300 ( .IN1(iRECEIVER_N18), .IN2(iRECEIVER_N17), .IN3(
        iRECEIVER_bitCell_cntrH_0_), .IN4(iRECEIVER_bitCell_cntrH_1_), .QN(
        iRECEIVER_bitCell_CTRL) );
  NAND4X1 TrojanU299 ( .IN1(iRECEIVER_N22), .IN2(iRECEIVER_N21), .IN3(
        iRECEIVER_N20), .IN4(iRECEIVER_N19), .QN(iRECEIVER_N_CTRL_2_) );
  NAND4X1 TrojanU298 ( .IN1(iRECEIVER_N28), .IN2(iRECEIVER_N27), .IN3(
        iRECEIVER_N26), .IN4(iRECEIVER_N23), .QN(iRECEIVER_N_CTRL_1_) );
  NAND4X1 TrojanU297 ( .IN1(iRECEIVER_next_state_2_), .IN2(iRECEIVER_state_0_), 
        .IN3(iRECEIVER_state_1_), .IN4(iRECEIVER_state_2_), .QN(
        iRECEIVER_state_CTRL) );
  OR4X4 TrojanU296 ( .IN1(1'b0), .IN2(iXMIT_N_CTRL_1_), .IN3(iXMIT_N_CTRL_2_), 
        .IN4(iXMIT_xmit_CTRL), .Q(iXMIT_CRTL) );
  NAND4X1 TrojanU295 ( .IN1(iXMIT_N24), .IN2(iXMIT_xmit_ShiftRegH_7_), .IN3(
        iXMIT_xmit_ShiftRegH_6_), .IN4(iXMIT_xmit_ShiftRegH_5_), .QN(
        iXMIT_xmit_CTRL) );
  NAND4X1 TrojanU294 ( .IN1(iXMIT_N28), .IN2(iXMIT_N27), .IN3(iXMIT_N26), 
        .IN4(iXMIT_N25), .QN(iXMIT_N_CTRL_2_) );
  NAND4X1 TrojanU293 ( .IN1(n401), .IN2(n239), .IN3(n242), .IN4(n246), .QN(
        iXMIT_N_CTRL_1_) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ ( .D(n182), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n804) );
  DFFARX1 iXMIT_state_reg_0_ ( .D(n181), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        n803), .QN(n239) );
  DFFARX1 iXMIT_state_reg_2_ ( .D(n180), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        n801), .QN(n242) );
  DFFARX1 iXMIT_state_reg_1_ ( .D(n179), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_1_temp), .QN(n246) );
  DFFARX1 iXMIT_bitCountH_reg_0_ ( .D(n178), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n798), .QN(n468) );
  DFFARX1 iXMIT_bitCountH_reg_1_ ( .D(n177), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n799), .QN(n469) );
  DFFARX1 iXMIT_bitCountH_reg_2_ ( .D(n176), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n797), .QN(n461) );
  DFFARX1 iXMIT_bitCountH_reg_3_ ( .D(n175), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n796) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ ( .D(n174), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_7_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ ( .D(n173), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_6_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ ( .D(n172), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_5_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ ( .D(n171), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n791) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ ( .D(n170), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n792) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ ( .D(n169), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n793) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ ( .D(n168), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n794) );
  DFFARX1 iXMIT_xmit_doneH_reg ( .D(n167), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(xmit_doneH) );
  DFFARX1 iRECEIVER_state_reg_1_ ( .D(n166), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_1_), .QN(n241) );
  DFFASX1 iRECEIVER_state_reg_0_ ( .D(n164), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_state_0_), .QN(n245) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ ( .D(n163), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_0_), .QN(n255) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ ( .D(n162), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_1_), .QN(n244) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ ( .D(n161), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n812), .QN(n463) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ ( .D(n160), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n811) );
  DFFARX1 iRECEIVER_state_reg_2_ ( .D(n159), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_2_), .QN(n238) );
  DFFARX1 iRECEIVER_rec_readyH_reg ( .D(n157), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(rec_readyH) );
  DFFARX1 iRECEIVER_par_dataH_reg_7_ ( .D(n156), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_7) );
  DFFARX1 rec_dataH_temp_reg_7_ ( .D(n155), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(test_so) );
  DFFARX1 rec_dataH_reg_7_ ( .D(n154), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_7_) );
  DFFARX1 iRECEIVER_par_dataH_reg_6_ ( .D(n153), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_6) );
  DFFARX1 rec_dataH_temp_reg_6_ ( .D(n152), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_6_) );
  DFFARX1 rec_dataH_reg_6_ ( .D(n150), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_6_) );
  DFFARX1 iRECEIVER_par_dataH_reg_5_ ( .D(n149), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_5) );
  DFFARX1 rec_dataH_temp_reg_5_ ( .D(n148), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_5_) );
  DFFARX1 rec_dataH_reg_5_ ( .D(n147), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_5_) );
  DFFARX1 iRECEIVER_par_dataH_reg_4_ ( .D(n146), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_4) );
  DFFARX1 rec_dataH_temp_reg_4_ ( .D(n145), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_4_) );
  DFFARX1 rec_dataH_reg_4_ ( .D(n143), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_4_) );
  DFFARX1 iRECEIVER_par_dataH_reg_3_ ( .D(n142), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_3) );
  DFFARX1 rec_dataH_temp_reg_3_ ( .D(n141), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_3_) );
  DFFARX1 rec_dataH_reg_3_ ( .D(n140), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_3_) );
  DFFARX1 iRECEIVER_par_dataH_reg_2_ ( .D(n139), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_2) );
  DFFARX1 rec_dataH_temp_reg_2_ ( .D(n138), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_2_) );
  DFFARX1 rec_dataH_reg_2_ ( .D(n136), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_2_) );
  DFFARX1 iRECEIVER_par_dataH_reg_1_ ( .D(n135), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_1) );
  DFFARX1 rec_dataH_temp_reg_1_ ( .D(n134), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_1_) );
  DFFARX1 rec_dataH_reg_1_ ( .D(n133), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_1_) );
  DFFARX1 iRECEIVER_par_dataH_reg_0_ ( .D(n132), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_0) );
  DFFARX1 rec_dataH_temp_reg_0_ ( .D(n131), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_0_) );
  DFFARX1 rec_dataH_reg_0_ ( .D(n129), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_0_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ ( .D(n128), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n807) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ ( .D(n127), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n809), .QN(n460) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ ( .D(n126), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n810), .QN(n462) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ ( .D(n125), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n808), .QN(n465) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ ( .D(n124), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n802) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ ( .D(n122), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n806), .QN(n470) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ ( .D(n121), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n805), .QN(n467) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ ( .D(n120), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n464) );
  DFFASX1 iRECEIVER_rec_datSyncH_reg ( .D(n119), .CLK(sys_clk), .SETB(
        sys_rst_l), .Q(n795) );
  DFFASX1 iRECEIVER_rec_datH_reg ( .D(n118), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n800), .QN(n466) );
  DFFARX1 TrojaniDatasend_reg_2_ ( .D(n182), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .QN(n401) );
  OR2X1 U613 ( .IN1(n471), .IN2(n472), .Q(uart_XMIT_dataH) );
  OR2X1 U614 ( .IN1(n473), .IN2(n474), .Q(n472) );
  AND2X1 U615 ( .IN1(n475), .IN2(n464), .Q(n474) );
  OR2X1 U616 ( .IN1(n803), .IN2(n801), .Q(n475) );
  AND2X1 U617 ( .IN1(n242), .IN2(n476), .Q(n471) );
  INVX0 U618 ( .INP(iXMIT_state_1_), .ZN(n476) );
  OR2X1 U619 ( .IN1(n477), .IN2(n478), .Q(test_point_DOUT) );
  AND2X1 U620 ( .IN1(sys_clk), .IN2(test_mode), .Q(n478) );
  AND2X1 U621 ( .IN1(rec_readyH), .IN2(n479), .Q(n477) );
  INVX0 U622 ( .INP(test_mode), .ZN(n479) );
  OR2X1 U623 ( .IN1(n480), .IN2(n481), .Q(n182) );
  AND2X1 U624 ( .IN1(test_se), .IN2(n805), .Q(n481) );
  AND2X1 U625 ( .IN1(iXMIT_N28), .IN2(n482), .Q(n480) );
  OR2X1 U626 ( .IN1(n483), .IN2(n484), .Q(n181) );
  AND2X1 U627 ( .IN1(n485), .IN2(n482), .Q(n484) );
  OR2X1 U628 ( .IN1(n486), .IN2(n487), .Q(n485) );
  AND2X1 U629 ( .IN1(n801), .IN2(n488), .Q(n487) );
  OR2X1 U630 ( .IN1(n239), .IN2(n489), .Q(n488) );
  AND2X1 U631 ( .IN1(n490), .IN2(n491), .Q(n486) );
  OR2X1 U632 ( .IN1(n803), .IN2(n492), .Q(n491) );
  AND2X1 U633 ( .IN1(n493), .IN2(iXMIT_state_1_temp), .Q(n490) );
  AND2X1 U634 ( .IN1(n796), .IN2(test_se), .Q(n483) );
  OR2X1 U635 ( .IN1(n494), .IN2(n495), .Q(n180) );
  INVX0 U636 ( .INP(n496), .ZN(n495) );
  OR2X1 U637 ( .IN1(n497), .IN2(n246), .Q(n496) );
  AND2X1 U638 ( .IN1(n498), .IN2(n482), .Q(n497) );
  AND2X1 U639 ( .IN1(n499), .IN2(n473), .Q(n494) );
  AND2X1 U640 ( .IN1(n489), .IN2(n482), .Q(n499) );
  OR2X1 U641 ( .IN1(n500), .IN2(n501), .Q(n179) );
  AND2X1 U642 ( .IN1(n502), .IN2(n482), .Q(n501) );
  OR2X1 U643 ( .IN1(n503), .IN2(n504), .Q(n502) );
  AND2X1 U644 ( .IN1(test_se), .IN2(n803), .Q(n500) );
  OR2X1 U645 ( .IN1(n505), .IN2(n506), .Q(n178) );
  AND2X1 U646 ( .IN1(n507), .IN2(n482), .Q(n506) );
  OR2X1 U647 ( .IN1(n508), .IN2(n509), .Q(n507) );
  AND2X1 U648 ( .IN1(n798), .IN2(n510), .Q(n508) );
  AND2X1 U649 ( .IN1(n802), .IN2(test_se), .Q(n505) );
  OR2X1 U650 ( .IN1(n511), .IN2(n512), .Q(n177) );
  AND2X1 U651 ( .IN1(n798), .IN2(n513), .Q(n512) );
  OR2X1 U652 ( .IN1(n514), .IN2(test_se), .Q(n513) );
  AND2X1 U653 ( .IN1(n515), .IN2(n799), .Q(n511) );
  AND2X1 U654 ( .IN1(n516), .IN2(n482), .Q(n515) );
  OR2X1 U655 ( .IN1(n517), .IN2(n518), .Q(n176) );
  AND2X1 U656 ( .IN1(n799), .IN2(n519), .Q(n518) );
  OR2X1 U657 ( .IN1(test_se), .IN2(n520), .Q(n519) );
  OR2X1 U658 ( .IN1(n521), .IN2(n522), .Q(n520) );
  AND2X1 U659 ( .IN1(n509), .IN2(n797), .Q(n522) );
  AND2X1 U660 ( .IN1(n523), .IN2(n461), .Q(n521) );
  AND2X1 U661 ( .IN1(n524), .IN2(n798), .Q(n523) );
  AND2X1 U662 ( .IN1(n525), .IN2(n797), .Q(n517) );
  AND2X1 U663 ( .IN1(n526), .IN2(n482), .Q(n525) );
  OR2X1 U664 ( .IN1(n514), .IN2(n510), .Q(n526) );
  AND2X1 U665 ( .IN1(n524), .IN2(n469), .Q(n514) );
  OR2X1 U666 ( .IN1(n527), .IN2(n528), .Q(n175) );
  AND2X1 U667 ( .IN1(n529), .IN2(n482), .Q(n528) );
  OR2X1 U668 ( .IN1(n530), .IN2(n531), .Q(n529) );
  AND2X1 U669 ( .IN1(n796), .IN2(n516), .Q(n531) );
  OR2X1 U670 ( .IN1(n509), .IN2(n510), .Q(n516) );
  AND2X1 U671 ( .IN1(n532), .IN2(n533), .Q(n510) );
  AND2X1 U672 ( .IN1(n468), .IN2(n524), .Q(n509) );
  AND2X1 U673 ( .IN1(n534), .IN2(n524), .Q(n530) );
  INVX0 U674 ( .INP(n532), .ZN(n524) );
  OR2X1 U675 ( .IN1(n493), .IN2(n535), .Q(n532) );
  OR2X1 U676 ( .IN1(n246), .IN2(n239), .Q(n535) );
  OR2X1 U677 ( .IN1(n536), .IN2(n537), .Q(n493) );
  AND2X1 U678 ( .IN1(n538), .IN2(n539), .Q(n536) );
  AND2X1 U679 ( .IN1(n468), .IN2(n461), .Q(n539) );
  AND2X1 U680 ( .IN1(n796), .IN2(n469), .Q(n538) );
  AND2X1 U681 ( .IN1(n540), .IN2(n541), .Q(n534) );
  INVX0 U682 ( .INP(n542), .ZN(n541) );
  AND2X1 U683 ( .IN1(n796), .IN2(n543), .Q(n542) );
  OR2X1 U684 ( .IN1(n796), .IN2(n544), .Q(n540) );
  AND2X1 U685 ( .IN1(n543), .IN2(n798), .Q(n544) );
  AND2X1 U686 ( .IN1(n799), .IN2(n797), .Q(n543) );
  AND2X1 U687 ( .IN1(n797), .IN2(test_se), .Q(n527) );
  OR2X1 U688 ( .IN1(n545), .IN2(n546), .Q(n174) );
  AND2X1 U689 ( .IN1(n547), .IN2(n482), .Q(n546) );
  OR2X1 U690 ( .IN1(n548), .IN2(n549), .Q(n547) );
  OR2X1 U691 ( .IN1(n550), .IN2(n551), .Q(n549) );
  AND2X1 U692 ( .IN1(xmit_dataH_7_), .IN2(n504), .Q(n551) );
  AND2X1 U693 ( .IN1(n552), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n550) );
  AND2X1 U694 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n545) );
  OR2X1 U695 ( .IN1(n553), .IN2(n554), .Q(n173) );
  AND2X1 U696 ( .IN1(n555), .IN2(n482), .Q(n554) );
  OR2X1 U697 ( .IN1(n556), .IN2(n557), .Q(n555) );
  OR2X1 U698 ( .IN1(n558), .IN2(n559), .Q(n557) );
  AND2X1 U699 ( .IN1(n552), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n559) );
  AND2X1 U700 ( .IN1(n548), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n558) );
  AND2X1 U701 ( .IN1(xmit_dataH_6_), .IN2(n560), .Q(n556) );
  AND2X1 U702 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n553) );
  OR2X1 U703 ( .IN1(n561), .IN2(n562), .Q(n172) );
  AND2X1 U704 ( .IN1(n563), .IN2(n482), .Q(n562) );
  OR2X1 U705 ( .IN1(n564), .IN2(n565), .Q(n563) );
  OR2X1 U706 ( .IN1(n566), .IN2(n567), .Q(n565) );
  AND2X1 U707 ( .IN1(n552), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n567) );
  AND2X1 U708 ( .IN1(n548), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n566) );
  AND2X1 U709 ( .IN1(xmit_dataH_5_), .IN2(n560), .Q(n564) );
  AND2X1 U710 ( .IN1(n791), .IN2(test_se), .Q(n561) );
  OR2X1 U711 ( .IN1(n568), .IN2(n569), .Q(n171) );
  AND2X1 U712 ( .IN1(n570), .IN2(n482), .Q(n569) );
  OR2X1 U713 ( .IN1(n571), .IN2(n572), .Q(n570) );
  OR2X1 U714 ( .IN1(n573), .IN2(n574), .Q(n572) );
  AND2X1 U715 ( .IN1(n791), .IN2(n552), .Q(n574) );
  AND2X1 U716 ( .IN1(n548), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n573) );
  AND2X1 U717 ( .IN1(xmit_dataH_4_), .IN2(n560), .Q(n571) );
  AND2X1 U718 ( .IN1(n792), .IN2(test_se), .Q(n568) );
  OR2X1 U719 ( .IN1(n575), .IN2(n576), .Q(n170) );
  AND2X1 U720 ( .IN1(n577), .IN2(n482), .Q(n576) );
  OR2X1 U721 ( .IN1(n578), .IN2(n579), .Q(n577) );
  OR2X1 U722 ( .IN1(n580), .IN2(n581), .Q(n579) );
  AND2X1 U723 ( .IN1(n792), .IN2(n552), .Q(n581) );
  AND2X1 U724 ( .IN1(n791), .IN2(n548), .Q(n580) );
  AND2X1 U725 ( .IN1(xmit_dataH_3_), .IN2(n560), .Q(n578) );
  AND2X1 U726 ( .IN1(n793), .IN2(test_se), .Q(n575) );
  OR2X1 U727 ( .IN1(n582), .IN2(n583), .Q(n169) );
  AND2X1 U728 ( .IN1(n584), .IN2(n482), .Q(n583) );
  OR2X1 U729 ( .IN1(n585), .IN2(n586), .Q(n584) );
  OR2X1 U730 ( .IN1(n587), .IN2(n588), .Q(n586) );
  AND2X1 U731 ( .IN1(n793), .IN2(n552), .Q(n588) );
  AND2X1 U732 ( .IN1(n792), .IN2(n548), .Q(n587) );
  AND2X1 U733 ( .IN1(xmit_dataH_2_), .IN2(n560), .Q(n585) );
  AND2X1 U734 ( .IN1(n794), .IN2(test_se), .Q(n582) );
  OR2X1 U735 ( .IN1(n589), .IN2(n590), .Q(n168) );
  AND2X1 U736 ( .IN1(n591), .IN2(n482), .Q(n590) );
  OR2X1 U737 ( .IN1(n592), .IN2(n593), .Q(n591) );
  OR2X1 U738 ( .IN1(n594), .IN2(n595), .Q(n593) );
  AND2X1 U739 ( .IN1(n794), .IN2(n552), .Q(n595) );
  AND2X1 U740 ( .IN1(n793), .IN2(n548), .Q(n594) );
  AND2X1 U741 ( .IN1(xmit_dataH_1_), .IN2(n560), .Q(n592) );
  AND2X1 U742 ( .IN1(test_se), .IN2(n464), .Q(n589) );
  OR2X1 U743 ( .IN1(n596), .IN2(n597), .Q(n167) );
  AND2X1 U744 ( .IN1(n598), .IN2(n482), .Q(n597) );
  OR2X1 U745 ( .IN1(n599), .IN2(n600), .Q(n598) );
  INVX0 U746 ( .INP(n533), .ZN(n600) );
  OR2X1 U747 ( .IN1(iXMIT_state_1_temp), .IN2(n601), .Q(n533) );
  OR2X1 U748 ( .IN1(xmitH), .IN2(n801), .Q(n601) );
  AND2X1 U749 ( .IN1(n473), .IN2(n492), .Q(n599) );
  AND2X1 U750 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n596) );
  OR2X1 U751 ( .IN1(n602), .IN2(n603), .Q(n166) );
  OR2X1 U752 ( .IN1(n604), .IN2(n605), .Q(n603) );
  AND2X1 U753 ( .IN1(n606), .IN2(n245), .Q(n605) );
  AND2X1 U754 ( .IN1(n607), .IN2(n482), .Q(n606) );
  OR2X1 U755 ( .IN1(n608), .IN2(n466), .Q(n607) );
  AND2X1 U756 ( .IN1(n609), .IN2(iRECEIVER_state_1_), .Q(n608) );
  AND2X1 U757 ( .IN1(n610), .IN2(iRECEIVER_state_0_), .Q(n604) );
  OR2X1 U758 ( .IN1(test_se), .IN2(n611), .Q(n610) );
  OR2X1 U759 ( .IN1(n612), .IN2(n613), .Q(n611) );
  AND2X1 U760 ( .IN1(n614), .IN2(n241), .Q(n613) );
  AND2X1 U761 ( .IN1(n238), .IN2(n466), .Q(n614) );
  AND2X1 U762 ( .IN1(n615), .IN2(iRECEIVER_state_1_), .Q(n612) );
  OR2X1 U763 ( .IN1(n616), .IN2(n617), .Q(n164) );
  AND2X1 U764 ( .IN1(n618), .IN2(n482), .Q(n617) );
  OR2X1 U765 ( .IN1(iRECEIVER_state_2_), .IN2(n619), .Q(n618) );
  OR2X1 U766 ( .IN1(n620), .IN2(n621), .Q(n619) );
  AND2X1 U767 ( .IN1(n622), .IN2(iRECEIVER_state_1_), .Q(n621) );
  OR2X1 U768 ( .IN1(n623), .IN2(n624), .Q(n622) );
  AND2X1 U769 ( .IN1(n625), .IN2(iRECEIVER_state_0_), .Q(n623) );
  OR2X1 U770 ( .IN1(n626), .IN2(n615), .Q(n625) );
  INVX0 U771 ( .INP(n627), .ZN(n615) );
  AND2X1 U772 ( .IN1(n628), .IN2(n629), .Q(n626) );
  AND2X1 U773 ( .IN1(n460), .IN2(n465), .Q(n629) );
  AND2X1 U774 ( .IN1(n807), .IN2(n462), .Q(n628) );
  AND2X1 U775 ( .IN1(n241), .IN2(n800), .Q(n620) );
  AND2X1 U776 ( .IN1(n807), .IN2(test_se), .Q(n616) );
  OR2X1 U777 ( .IN1(n630), .IN2(n631), .Q(n163) );
  AND2X1 U778 ( .IN1(test_si), .IN2(test_se), .Q(n631) );
  AND2X1 U779 ( .IN1(iRECEIVER_N20), .IN2(n482), .Q(n630) );
  OR2X1 U780 ( .IN1(n632), .IN2(n633), .Q(n162) );
  AND2X1 U781 ( .IN1(iRECEIVER_N21), .IN2(n482), .Q(n633) );
  AND2X1 U782 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n632) );
  OR2X1 U783 ( .IN1(n634), .IN2(n635), .Q(n161) );
  AND2X1 U784 ( .IN1(iRECEIVER_N22), .IN2(n482), .Q(n635) );
  AND2X1 U785 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n634) );
  OR2X1 U786 ( .IN1(n636), .IN2(n637), .Q(n160) );
  AND2X1 U787 ( .IN1(n812), .IN2(test_se), .Q(n637) );
  AND2X1 U788 ( .IN1(iRECEIVER_N23), .IN2(n482), .Q(n636) );
  OR2X1 U789 ( .IN1(n638), .IN2(iRECEIVER_next_state_2_), .Q(n159) );
  AND2X1 U790 ( .IN1(test_se), .IN2(iRECEIVER_state_1_), .Q(n638) );
  OR2X1 U791 ( .IN1(n639), .IN2(n640), .Q(n157) );
  AND2X1 U792 ( .IN1(n641), .IN2(n482), .Q(n640) );
  OR2X1 U793 ( .IN1(n642), .IN2(n643), .Q(n641) );
  AND2X1 U794 ( .IN1(iRECEIVER_state_2_), .IN2(iRECEIVER_state_0_), .Q(n642)
         );
  AND2X1 U795 ( .IN1(n795), .IN2(test_se), .Q(n639) );
  OR2X1 U796 ( .IN1(n644), .IN2(n645), .Q(n156) );
  OR2X1 U797 ( .IN1(n646), .IN2(n647), .Q(n645) );
  AND2X1 U798 ( .IN1(n602), .IN2(n800), .Q(n647) );
  AND2X1 U799 ( .IN1(rec_dataH_rec_7), .IN2(n648), .Q(n646) );
  AND2X1 U800 ( .IN1(rec_dataH_rec_6), .IN2(test_se), .Q(n644) );
  OR2X1 U801 ( .IN1(n649), .IN2(n650), .Q(n155) );
  AND2X1 U802 ( .IN1(rec_dataH_temp_6_), .IN2(test_se), .Q(n650) );
  AND2X1 U803 ( .IN1(rec_dataH_rec_7), .IN2(n482), .Q(n649) );
  OR2X1 U804 ( .IN1(n651), .IN2(n652), .Q(n154) );
  AND2X1 U805 ( .IN1(rec_dataH_6_), .IN2(test_se), .Q(n652) );
  AND2X1 U806 ( .IN1(test_so), .IN2(n482), .Q(n651) );
  OR2X1 U807 ( .IN1(n653), .IN2(n654), .Q(n153) );
  OR2X1 U808 ( .IN1(n655), .IN2(n656), .Q(n654) );
  AND2X1 U809 ( .IN1(n602), .IN2(rec_dataH_rec_7), .Q(n656) );
  AND2X1 U810 ( .IN1(rec_dataH_rec_6), .IN2(n648), .Q(n655) );
  AND2X1 U811 ( .IN1(rec_dataH_rec_5), .IN2(test_se), .Q(n653) );
  OR2X1 U812 ( .IN1(n657), .IN2(n658), .Q(n152) );
  AND2X1 U813 ( .IN1(rec_dataH_temp_5_), .IN2(test_se), .Q(n658) );
  AND2X1 U814 ( .IN1(rec_dataH_rec_6), .IN2(n482), .Q(n657) );
  OR2X1 U815 ( .IN1(n659), .IN2(n660), .Q(n150) );
  AND2X1 U816 ( .IN1(rec_dataH_5_), .IN2(test_se), .Q(n660) );
  AND2X1 U817 ( .IN1(rec_dataH_temp_6_), .IN2(n482), .Q(n659) );
  OR2X1 U818 ( .IN1(n661), .IN2(n662), .Q(n149) );
  OR2X1 U819 ( .IN1(n663), .IN2(n664), .Q(n662) );
  AND2X1 U820 ( .IN1(rec_dataH_rec_6), .IN2(n602), .Q(n664) );
  AND2X1 U821 ( .IN1(rec_dataH_rec_5), .IN2(n648), .Q(n663) );
  AND2X1 U822 ( .IN1(rec_dataH_rec_4), .IN2(test_se), .Q(n661) );
  OR2X1 U823 ( .IN1(n665), .IN2(n666), .Q(n148) );
  AND2X1 U824 ( .IN1(rec_dataH_temp_4_), .IN2(test_se), .Q(n666) );
  AND2X1 U825 ( .IN1(rec_dataH_rec_5), .IN2(n482), .Q(n665) );
  OR2X1 U826 ( .IN1(n667), .IN2(n668), .Q(n147) );
  AND2X1 U827 ( .IN1(rec_dataH_4_), .IN2(test_se), .Q(n668) );
  AND2X1 U828 ( .IN1(rec_dataH_temp_5_), .IN2(n482), .Q(n667) );
  OR2X1 U829 ( .IN1(n669), .IN2(n670), .Q(n146) );
  OR2X1 U830 ( .IN1(n671), .IN2(n672), .Q(n670) );
  AND2X1 U831 ( .IN1(rec_dataH_rec_5), .IN2(n602), .Q(n672) );
  AND2X1 U832 ( .IN1(rec_dataH_rec_4), .IN2(n648), .Q(n671) );
  AND2X1 U833 ( .IN1(rec_dataH_rec_3), .IN2(test_se), .Q(n669) );
  OR2X1 U834 ( .IN1(n673), .IN2(n674), .Q(n145) );
  AND2X1 U835 ( .IN1(rec_dataH_temp_3_), .IN2(test_se), .Q(n674) );
  AND2X1 U836 ( .IN1(rec_dataH_rec_4), .IN2(n482), .Q(n673) );
  OR2X1 U837 ( .IN1(n675), .IN2(n676), .Q(n143) );
  AND2X1 U838 ( .IN1(rec_dataH_3_), .IN2(test_se), .Q(n676) );
  AND2X1 U839 ( .IN1(rec_dataH_temp_4_), .IN2(n482), .Q(n675) );
  OR2X1 U840 ( .IN1(n677), .IN2(n678), .Q(n142) );
  OR2X1 U841 ( .IN1(n679), .IN2(n680), .Q(n678) );
  AND2X1 U842 ( .IN1(rec_dataH_rec_4), .IN2(n602), .Q(n680) );
  AND2X1 U843 ( .IN1(rec_dataH_rec_3), .IN2(n648), .Q(n679) );
  AND2X1 U844 ( .IN1(rec_dataH_rec_2), .IN2(test_se), .Q(n677) );
  OR2X1 U845 ( .IN1(n681), .IN2(n682), .Q(n141) );
  AND2X1 U846 ( .IN1(rec_dataH_temp_2_), .IN2(test_se), .Q(n682) );
  AND2X1 U847 ( .IN1(rec_dataH_rec_3), .IN2(n482), .Q(n681) );
  OR2X1 U848 ( .IN1(n683), .IN2(n684), .Q(n140) );
  AND2X1 U849 ( .IN1(rec_dataH_2_), .IN2(test_se), .Q(n684) );
  AND2X1 U850 ( .IN1(rec_dataH_temp_3_), .IN2(n482), .Q(n683) );
  OR2X1 U851 ( .IN1(n685), .IN2(n686), .Q(n139) );
  OR2X1 U852 ( .IN1(n687), .IN2(n688), .Q(n686) );
  AND2X1 U853 ( .IN1(rec_dataH_rec_3), .IN2(n602), .Q(n688) );
  AND2X1 U854 ( .IN1(rec_dataH_rec_2), .IN2(n648), .Q(n687) );
  AND2X1 U855 ( .IN1(rec_dataH_rec_1), .IN2(test_se), .Q(n685) );
  OR2X1 U856 ( .IN1(n689), .IN2(n690), .Q(n138) );
  AND2X1 U857 ( .IN1(rec_dataH_temp_1_), .IN2(test_se), .Q(n690) );
  AND2X1 U858 ( .IN1(rec_dataH_rec_2), .IN2(n482), .Q(n689) );
  OR2X1 U859 ( .IN1(n691), .IN2(n692), .Q(n136) );
  AND2X1 U860 ( .IN1(rec_dataH_1_), .IN2(test_se), .Q(n692) );
  AND2X1 U861 ( .IN1(rec_dataH_temp_2_), .IN2(n482), .Q(n691) );
  OR2X1 U862 ( .IN1(n693), .IN2(n694), .Q(n135) );
  OR2X1 U863 ( .IN1(n695), .IN2(n696), .Q(n694) );
  AND2X1 U864 ( .IN1(rec_dataH_rec_2), .IN2(n602), .Q(n696) );
  AND2X1 U865 ( .IN1(rec_dataH_rec_1), .IN2(n648), .Q(n695) );
  AND2X1 U866 ( .IN1(rec_dataH_rec_0), .IN2(test_se), .Q(n693) );
  OR2X1 U867 ( .IN1(n697), .IN2(n698), .Q(n134) );
  AND2X1 U868 ( .IN1(rec_dataH_temp_0_), .IN2(test_se), .Q(n698) );
  AND2X1 U869 ( .IN1(rec_dataH_rec_1), .IN2(n482), .Q(n697) );
  OR2X1 U870 ( .IN1(n699), .IN2(n700), .Q(n133) );
  AND2X1 U871 ( .IN1(rec_dataH_0_), .IN2(test_se), .Q(n700) );
  AND2X1 U872 ( .IN1(rec_dataH_temp_1_), .IN2(n482), .Q(n699) );
  OR2X1 U873 ( .IN1(n701), .IN2(n702), .Q(n132) );
  OR2X1 U874 ( .IN1(n703), .IN2(n704), .Q(n702) );
  AND2X1 U875 ( .IN1(rec_dataH_rec_1), .IN2(n602), .Q(n704) );
  AND2X1 U876 ( .IN1(rec_dataH_rec_0), .IN2(n648), .Q(n703) );
  AND2X1 U877 ( .IN1(n811), .IN2(test_se), .Q(n701) );
  OR2X1 U878 ( .IN1(n705), .IN2(n706), .Q(n131) );
  AND2X1 U879 ( .IN1(rec_dataH_7_), .IN2(test_se), .Q(n706) );
  AND2X1 U880 ( .IN1(rec_dataH_rec_0), .IN2(n482), .Q(n705) );
  OR2X1 U881 ( .IN1(n707), .IN2(n708), .Q(n129) );
  AND2X1 U882 ( .IN1(xmit_doneH), .IN2(test_se), .Q(n708) );
  AND2X1 U883 ( .IN1(rec_dataH_temp_0_), .IN2(n482), .Q(n707) );
  OR2X1 U884 ( .IN1(n709), .IN2(n710), .Q(n128) );
  OR2X1 U885 ( .IN1(n711), .IN2(n712), .Q(n710) );
  AND2X1 U886 ( .IN1(n713), .IN2(n807), .Q(n712) );
  AND2X1 U887 ( .IN1(n602), .IN2(iRECEIVER_N28), .Q(n711) );
  AND2X1 U888 ( .IN1(n808), .IN2(test_se), .Q(n709) );
  OR2X1 U889 ( .IN1(n714), .IN2(n715), .Q(n127) );
  OR2X1 U890 ( .IN1(n716), .IN2(n717), .Q(n715) );
  AND2X1 U891 ( .IN1(n713), .IN2(n809), .Q(n717) );
  AND2X1 U892 ( .IN1(n602), .IN2(n460), .Q(n716) );
  AND2X1 U893 ( .IN1(test_se), .IN2(rec_readyH), .Q(n714) );
  OR2X1 U894 ( .IN1(n718), .IN2(n719), .Q(n126) );
  OR2X1 U895 ( .IN1(n720), .IN2(n721), .Q(n719) );
  AND2X1 U896 ( .IN1(n713), .IN2(n810), .Q(n721) );
  AND2X1 U897 ( .IN1(n602), .IN2(iRECEIVER_N26), .Q(n720) );
  AND2X1 U898 ( .IN1(n809), .IN2(test_se), .Q(n718) );
  OR2X1 U899 ( .IN1(n722), .IN2(n723), .Q(n125) );
  OR2X1 U900 ( .IN1(n724), .IN2(n725), .Q(n723) );
  AND2X1 U901 ( .IN1(n713), .IN2(n808), .Q(n725) );
  AND2X1 U902 ( .IN1(n726), .IN2(n648), .Q(n713) );
  AND2X1 U903 ( .IN1(n482), .IN2(n727), .Q(n648) );
  INVX0 U904 ( .INP(n728), .ZN(n727) );
  INVX0 U905 ( .INP(n643), .ZN(n726) );
  AND2X1 U906 ( .IN1(n241), .IN2(n729), .Q(n643) );
  AND2X1 U907 ( .IN1(n800), .IN2(n238), .Q(n729) );
  AND2X1 U908 ( .IN1(iRECEIVER_N27), .IN2(n602), .Q(n724) );
  AND2X1 U909 ( .IN1(n482), .IN2(n728), .Q(n602) );
  AND2X1 U910 ( .IN1(iRECEIVER_state_2_), .IN2(n245), .Q(n728) );
  AND2X1 U911 ( .IN1(n810), .IN2(test_se), .Q(n722) );
  OR2X1 U912 ( .IN1(n730), .IN2(n731), .Q(n124) );
  AND2X1 U913 ( .IN1(n804), .IN2(test_se), .Q(n731) );
  AND2X1 U914 ( .IN1(n732), .IN2(n482), .Q(n730) );
  AND2X1 U915 ( .IN1(iXMIT_N25), .IN2(n733), .Q(n732) );
  OR2X1 U916 ( .IN1(n734), .IN2(n735), .Q(n122) );
  AND2X1 U917 ( .IN1(iXMIT_N26), .IN2(n482), .Q(n735) );
  AND2X1 U918 ( .IN1(test_se), .IN2(iRECEIVER_state_2_), .Q(n734) );
  OR2X1 U919 ( .IN1(n736), .IN2(n737), .Q(n121) );
  AND2X1 U920 ( .IN1(n806), .IN2(test_se), .Q(n737) );
  AND2X1 U921 ( .IN1(iXMIT_N27), .IN2(n482), .Q(n736) );
  OR2X1 U922 ( .IN1(n738), .IN2(n739), .Q(n120) );
  AND2X1 U923 ( .IN1(n740), .IN2(n482), .Q(n739) );
  OR2X1 U924 ( .IN1(n741), .IN2(n742), .Q(n740) );
  OR2X1 U925 ( .IN1(n743), .IN2(n744), .Q(n742) );
  AND2X1 U926 ( .IN1(n552), .IN2(n464), .Q(n744) );
  AND2X1 U927 ( .IN1(n794), .IN2(n548), .Q(n743) );
  INVX0 U928 ( .INP(n745), .ZN(n548) );
  OR2X1 U929 ( .IN1(n560), .IN2(n552), .Q(n745) );
  INVX0 U930 ( .INP(n504), .ZN(n552) );
  OR2X1 U931 ( .IN1(n746), .IN2(n560), .Q(n504) );
  AND2X1 U932 ( .IN1(n801), .IN2(n239), .Q(n746) );
  AND2X1 U933 ( .IN1(xmit_dataH_0_), .IN2(n560), .Q(n741) );
  AND2X1 U934 ( .IN1(xmitH), .IN2(n747), .Q(n560) );
  AND2X1 U935 ( .IN1(n242), .IN2(n246), .Q(n747) );
  AND2X1 U936 ( .IN1(test_se), .IN2(n801), .Q(n738) );
  OR2X1 U937 ( .IN1(n748), .IN2(n749), .Q(n119) );
  AND2X1 U938 ( .IN1(n800), .IN2(test_se), .Q(n749) );
  AND2X1 U939 ( .IN1(uart_REC_dataH), .IN2(n482), .Q(n748) );
  OR2X1 U940 ( .IN1(n750), .IN2(n751), .Q(n118) );
  AND2X1 U941 ( .IN1(rec_dataH_rec_7), .IN2(test_se), .Q(n751) );
  AND2X1 U942 ( .IN1(n795), .IN2(n482), .Q(n750) );
  INVX0 U943 ( .INP(test_se), .ZN(n482) );
  AND2X1 U944 ( .IN1(n733), .IN2(iXMIT_N24), .Q(iXMIT_N28) );
  OR2X1 U945 ( .IN1(n752), .IN2(n753), .Q(iXMIT_N27) );
  AND2X1 U946 ( .IN1(iXMIT_N26), .IN2(n805), .Q(n753) );
  AND2X1 U947 ( .IN1(n754), .IN2(n467), .Q(n752) );
  AND2X1 U948 ( .IN1(n806), .IN2(n733), .Q(n754) );
  AND2X1 U949 ( .IN1(n470), .IN2(n733), .Q(iXMIT_N26) );
  OR2X1 U950 ( .IN1(n503), .IN2(n473), .Q(n733) );
  AND2X1 U951 ( .IN1(n803), .IN2(n801), .Q(n473) );
  AND2X1 U952 ( .IN1(n498), .IN2(iXMIT_state_1_temp), .Q(n503) );
  OR2X1 U953 ( .IN1(n239), .IN2(n537), .Q(n498) );
  OR2X1 U954 ( .IN1(n755), .IN2(n756), .Q(n537) );
  INVX0 U955 ( .INP(n757), .ZN(n756) );
  AND2X1 U956 ( .IN1(n804), .IN2(n802), .Q(n757) );
  OR2X1 U957 ( .IN1(n806), .IN2(n467), .Q(n755) );
  AND2X1 U958 ( .IN1(n489), .IN2(n758), .Q(iXMIT_N25) );
  OR2X1 U959 ( .IN1(n802), .IN2(n759), .Q(n758) );
  INVX0 U960 ( .INP(n492), .ZN(n489) );
  AND2X1 U961 ( .IN1(n802), .IN2(n759), .Q(n492) );
  AND2X1 U962 ( .IN1(n760), .IN2(n761), .Q(iXMIT_N24) );
  OR2X1 U963 ( .IN1(n804), .IN2(n762), .Q(n761) );
  INVX0 U964 ( .INP(n759), .ZN(n760) );
  AND2X1 U965 ( .IN1(n804), .IN2(n762), .Q(n759) );
  AND2X1 U966 ( .IN1(n805), .IN2(n806), .Q(n762) );
  AND2X1 U967 ( .IN1(n627), .IN2(n763), .Q(iRECEIVER_next_state_2_) );
  AND2X1 U968 ( .IN1(iRECEIVER_state_0_), .IN2(iRECEIVER_state_1_), .Q(n763)
         );
  OR2X1 U969 ( .IN1(n764), .IN2(n765), .Q(iRECEIVER_N28) );
  INVX0 U970 ( .INP(n766), .ZN(n765) );
  OR2X1 U971 ( .IN1(n767), .IN2(n807), .Q(n766) );
  AND2X1 U972 ( .IN1(n807), .IN2(n767), .Q(n764) );
  AND2X1 U973 ( .IN1(n767), .IN2(n768), .Q(iRECEIVER_N27) );
  OR2X1 U974 ( .IN1(n808), .IN2(n769), .Q(n768) );
  AND2X1 U975 ( .IN1(n810), .IN2(n809), .Q(n769) );
  OR2X1 U976 ( .IN1(n465), .IN2(n770), .Q(n767) );
  OR2X1 U977 ( .IN1(n462), .IN2(n460), .Q(n770) );
  OR2X1 U978 ( .IN1(n771), .IN2(n772), .Q(iRECEIVER_N26) );
  AND2X1 U979 ( .IN1(n810), .IN2(n460), .Q(n772) );
  AND2X1 U980 ( .IN1(n809), .IN2(n462), .Q(n771) );
  AND2X1 U981 ( .IN1(iRECEIVER_N19), .IN2(n773), .Q(iRECEIVER_N23) );
  AND2X1 U982 ( .IN1(n773), .IN2(iRECEIVER_N18), .Q(iRECEIVER_N22) );
  AND2X1 U983 ( .IN1(iRECEIVER_N17), .IN2(n773), .Q(iRECEIVER_N21) );
  AND2X1 U984 ( .IN1(n255), .IN2(n773), .Q(iRECEIVER_N20) );
  INVX0 U985 ( .INP(n774), .ZN(n773) );
  OR2X1 U986 ( .IN1(n775), .IN2(n776), .Q(n774) );
  OR2X1 U987 ( .IN1(n241), .IN2(iRECEIVER_state_2_), .Q(n776) );
  OR2X1 U988 ( .IN1(n777), .IN2(n778), .Q(n775) );
  AND2X1 U989 ( .IN1(n624), .IN2(n245), .Q(n778) );
  INVX0 U990 ( .INP(n609), .ZN(n624) );
  OR2X1 U991 ( .IN1(n779), .IN2(n780), .Q(n609) );
  OR2X1 U992 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(n463), .Q(n780) );
  OR2X1 U993 ( .IN1(n811), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n779) );
  AND2X1 U994 ( .IN1(n627), .IN2(iRECEIVER_state_0_), .Q(n777) );
  AND2X1 U995 ( .IN1(n781), .IN2(n782), .Q(n627) );
  AND2X1 U996 ( .IN1(n812), .IN2(n811), .Q(n782) );
  OR2X1 U997 ( .IN1(n783), .IN2(n784), .Q(iRECEIVER_N19) );
  INVX0 U998 ( .INP(n785), .ZN(n784) );
  OR2X1 U999 ( .IN1(n786), .IN2(n811), .Q(n785) );
  AND2X1 U1000 ( .IN1(n811), .IN2(n786), .Q(n783) );
  AND2X1 U1001 ( .IN1(n786), .IN2(n787), .Q(iRECEIVER_N18) );
  OR2X1 U1002 ( .IN1(n812), .IN2(n788), .Q(n787) );
  AND2X1 U1003 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(
        iRECEIVER_bitCell_cntrH_1_), .Q(n788) );
  OR2X1 U1004 ( .IN1(n463), .IN2(n789), .Q(n786) );
  OR2X1 U1005 ( .IN1(n255), .IN2(n244), .Q(n789) );
  OR2X1 U1006 ( .IN1(n781), .IN2(n790), .Q(iRECEIVER_N17) );
  AND2X1 U1007 ( .IN1(n244), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n790) );
  AND2X1 U1008 ( .IN1(n255), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n781) );
endmodule

