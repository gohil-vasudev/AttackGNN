module s38417 ( CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, 
        g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, 
        g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, 
        g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, 
        g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, 
        g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, 
        g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
        g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
        g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
        g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
        g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
        g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
        g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
        g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, test_se, 
        test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, 
        test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, 
        test_si8, test_so8, test_si9, test_so9, test_si10, test_so10, 
        test_si11, test_so11, test_si12, test_so12, test_si13, test_so13, 
        test_si14, test_so14, test_si15, test_so15, test_si16, test_so16, 
        test_si17, test_so17, test_si18, test_so18, test_si19, test_so19, 
        test_si20, test_so20, test_si21, test_so21, test_si22, test_so22, 
        test_si23, test_so23, test_si24, test_so24, test_si25, test_so25, 
        test_si26, test_so26, test_si27, test_so27, test_si28, test_so28, 
        test_si29, test_so29, test_si30, test_so30, test_si31, test_so31, 
        test_si32, test_so32, test_si33, test_so33, test_si34, test_so34, 
        test_si35, test_so35, test_si36, test_so36, test_si37, test_so37, 
        test_si38, test_so38, test_si39, test_so39, test_si40, test_so40, 
        test_si41, test_so41, test_si42, test_so42, test_si43, test_so43, 
        test_si44, test_so44, test_si45, test_so45, test_si46, test_so46, 
        test_si47, test_so47, test_si48, test_so48, test_si49, test_so49, 
        test_si50, test_so50, test_si51, test_so51, test_si52, test_so52, 
        test_si53, test_so53, test_si54, test_so54, test_si55, test_so55, 
        test_si56, test_so56, test_si57, test_so57, test_si58, test_so58, 
        test_si59, test_so59, test_si60, test_so60, test_si61, test_so61, 
        test_si62, test_so62, test_si63, test_so63, test_si64, test_so64, 
        test_si65, test_so65, test_si66, test_so66, test_si67, test_so67, 
        test_si68, test_so68, test_si69, test_so69, test_si70, test_so70, 
        test_si71, test_so71, test_si72, test_so72, test_si73, test_so73, 
        test_si74, test_so74, test_si75, test_so75, test_si76, test_so76, 
        test_si77, test_so77, test_si78, test_so78, test_si79, test_so79, 
        test_si80, test_so80, test_si81, test_so81, test_si82, test_so82, 
        test_si83, test_so83, test_si84, test_so84, test_si85, test_so85, 
        test_si86, test_so86, test_si87, test_so87, test_si88, test_so88, 
        test_si89, test_so89, test_si90, test_so90, test_si91, test_so91, 
        test_si92, test_so92, test_si93, test_so93, test_si94, test_so94, 
        test_si95, test_so95, test_si96, test_so96, test_si97, test_so97, 
        test_si98, test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;
  wire   test_so3, test_so4, test_so5, test_so23, test_so57, test_so63,
         test_so73, test_so99, test_so100, n2230, n2217, n2231, n2374, n2361,
         n2375, DFF_2_n1, n4264, n2445, n2446, n2440, n2426, n2670, n2671,
         n2669, n2685, n2686, n2684, n2718, n2719, n2717, g2124, n2981, g1430,
         n2984, g744, n2987, g56, n2990, n3742, n3741, n8104, g16802, n8103,
         g16823, n8102, g2950, n4423, n4274, g2883, n4330, g22026, g2888,
         g23358, g2896, n4431, g24473, g2892, g25201, g2903, n4305, g26037,
         g2900, n4291, g26798, g2908, n4355, g2912, n4482, g23357, g2917,
         n4479, g24476, g2924, n4349, g25199, g2920, n4280, n4281, n8099,
         n8098, DFF_18_n1, n4279, g2879, n4351, g2934, g2935, g2938, g2941,
         g2944, g2947, g2953, g2956, g2959, g2962, g2963, g2969, g2972, g2975,
         g2978, g2981, g2874, g18754, g1506, n4288, g18781, g1501, n4565,
         g18803, g1496, n4557, g18821, g1491, n4326, g18835, g1486, n4390,
         g18852, g1481, n4320, g18866, g1476, n4374, g18883, g1471, n4378,
         g21880, g2877, g19154, g813, n4289, g19163, g809, n4567, g19173, g805,
         n4559, g19184, g801, n4327, g20310, g797, n4391, g20343, g793, n4321,
         g20376, g789, n4375, g20417, g785, n4379, g21878, g2873, g19153, g125,
         n4290, g19162, g121, n4569, g19172, g117, n4561, g19144, g113, n4328,
         g19149, g109, n4392, g19157, g105, n4322, g19167, g101, n4376, g19178,
         g97, n4380, g20874, g2857, g18885, g2200, n4287, g18975, g2195, n4563,
         g18968, g2190, n4555, g18942, g2185, n4325, g18906, g2180, n4389,
         g18867, g2175, n4319, g18836, g2170, n4373, g18957, g2165, n4377,
         g21882, g2878, n4598, n4382, n4383, g3109, n4494, g18669, g18719,
         g3211, g18782, g3084, g17222, g3085, g17225, g3086, g17234, g3087,
         g17224, g3091, g17228, g3092, g17246, g3093, g17226, g3094, g17235,
         g3095, g17269, g3096, g25450, g3097, g25451, g3098, g25452, g3099,
         g28420, g3100, g28421, g28425, g3102, g29936, g3103, g29939, g3104,
         g29941, g3105, g30796, g3106, g30798, g3107, g30801, g3108, g17229,
         g3155, g17247, g3158, g17302, g3161, g17236, g3164, g17270, g3167,
         g17340, g3170, g17248, g3173, g17303, g3176, g17383, g17271, g3182,
         g17341, g3185, g17429, g3088, n8090, n8089, g3197, n8088, g3201,
         n4406, g3204, g3207, n4329, g3188, n4405, g3133, n8087, g3128, n8086,
         n8084, DFF_144_n1, g3124, n8083, DFF_146_n1, n8082, n8081, n8080,
         g3112, g3110, g3111, n8079, n8078, n8077, n8076, g3151, n4424, g3142,
         n4301, g185, n4384, n4318, n4512, g165, n4369, g22100, g130, g22122,
         g131, g22141, g129, g22123, g133, g22142, g134, g22161, g132, g22025,
         g142, g22027, g143, g22030, g141, g22028, g145, g22031, g146, g22037,
         g22032, g148, g22038, g149, g22047, g147, g22039, g151, g22048, g152,
         g22063, g150, g22049, g154, g22064, g155, g22079, g153, g22065, g157,
         g22080, g158, g22101, g156, g22081, g160, g22102, g161, g22124, g159,
         g22103, g22125, g164, g22143, g162, g25204, g169, g25206, g170,
         g25211, g168, g25207, g172, g25212, g173, g25218, g171, g25213, g175,
         g25219, g176, g25228, g174, g25220, g178, g25229, g179, g25239, g177,
         g30261, g186, g30267, g30275, g192, g30637, g231, g30640, g234,
         g30645, g237, g30668, g195, g30674, g198, g30680, g201, g30641, g240,
         g30646, g243, g30653, g246, g30276, g204, g30284, g207, g30292, g210,
         g30254, g249, g30257, g252, g30262, g30245, g213, g30246, g216,
         g30248, g219, g30258, g258, g30263, g261, g30268, g264, g30635, g222,
         g30636, g225, g30639, g228, g30661, g267, g30669, g270, g30675, g273,
         g25027, g92, g25932, g88, g26529, g83, g27120, g27594, g74, g28145,
         g70, g28634, g65, g29109, g61, g29353, g29579, g52, g13110, g180,
         g181, n4506, g309, n4388, g27253, g354, g27255, g343, g27258, g27256,
         g369, g27259, g358, g27265, g361, g27260, g384, g27266, g373, g27277,
         g376, g27267, g398, g27278, g388, g27293, g391, g28732, g408, g28735,
         g411, g28744, g414, g29194, g417, g29197, g420, g29201, g423, g28736,
         g28745, g428, g28754, g426, g26803, g429, g26804, g432, g26807, g435,
         g26805, g438, g26808, g441, g26812, g444, g27759, g448, g27760, g449,
         g27762, g447, g29606, g312, g29608, g313, g29611, g314, g30699, g315,
         g30700, g30702, g317, g30455, g318, g30468, g319, g30482, g320,
         g29167, g322, g29169, g323, g29172, g321, g26655, g403, g26659, g404,
         g26664, g402, g450, n8066, DFF_299_n1, g452, n8065, DFF_301_n1, g454,
         DFF_303_n1, g280, n8062, DFF_305_n1, g282, n8061, DFF_307_n1, g284,
         n8060, DFF_309_n1, g286, n8059, DFF_311_n1, g288, n8058, DFF_313_n1,
         g290, n8057, n4485, n4282, n8056, g21346, g305, n4278, n8055,
         DFF_328_n1, g349, g350, g351, g352, g353, g357, g364, g365, g366,
         g367, g368, g372, g379, g380, g381, g383, g387, g394, g395, g396,
         g397, g324, g337, n4298, n4372, g550, n4313, g21842, g554, g18678,
         g557, n4360, g18726, g513, g523, g524, g455, g564, g569, g458, g570,
         g571, g461, g572, g573, g465, g574, g565, g566, g567, g471, g568,
         g489, n4461, g485, n4466, g23067, g486, g23093, g487, g23117, g488,
         g23385, g23399, g24174, g24178, g477, g24207, g478, g24216, g479,
         g23092, g480, g23000, g484, g23022, g464, g24206, g24215, g24228,
         g528, g535, g542, g13149, g543, g544, g21851, g548, g13111, g549,
         g499, n4541, g13160, g558, g559, g27261, g576, g27268, g577, g27279,
         g575, g27269, g579, g27280, g27294, g578, g27281, g582, g27295, g583,
         g27311, g581, g27296, g585, g27312, g586, g27327, g584, g24491, g587,
         g24498, g590, g24507, g593, g24499, g596, g24508, g599, g24519, g602,
         g28345, g614, g28349, g617, g28353, g28342, g605, g28344, g608,
         g28348, g611, g26541, g490, g26545, g493, g26553, g496, g506, n4570,
         g22578, n4571, g525, n8047, n8046, n8045, n8044, n8043, g536, g537,
         g24059, g538, n4492, n8040, n4359, g629, n4295, g16654, g630, g20314,
         g659, g20682, g640, n4404, g23136, g633, n4478, g23324, g653, n4422,
         g24426, g646, n4414, g25185, g660, n4403, g26660, g672, n4413, g26776,
         g27672, g679, n4477, g28199, g686, n4396, g28668, g692, n4418, g20875,
         g699, g20879, g700, g20891, g698, g20880, g702, g20892, g703, g20901,
         g701, g20893, g705, g20902, g706, g20921, g704, g20903, g708, g20922,
         g709, g20944, g707, g20923, g20945, g712, g20966, g710, g20946, g714,
         g20967, g715, g20989, g713, g20968, g717, g20990, g718, g21009, g716,
         g20991, g720, g21010, g721, g21031, g719, g21011, g723, g21032, g724,
         g21051, g722, g20876, g726, g20881, g20894, g725, g20924, g729,
         g20947, g730, g20969, g728, g20948, g732, g20970, g733, g20992, g731,
         g25260, g735, g25262, g736, g25266, g734, g22218, g738, g22231, g739,
         g22242, g737, n4323, n4312, g22126, g818, g22145, g819, g22162, g817,
         g22146, g821, g22163, g822, g22177, g820, g22029, g830, g22033, g831,
         g22040, g829, g22034, g833, g22041, g834, g22054, g832, g22042, g836,
         g22055, g837, g22066, g835, g22056, g22067, g840, g22087, g838,
         g22068, g842, g22088, g843, g22104, g841, g22089, g845, g22105, g846,
         g22127, g844, g22106, g848, g22128, g849, g22147, g847, g22129, g851,
         g22148, g852, g22164, g850, g25209, g857, g25214, g25221, g856,
         g25215, g860, g25222, g861, g25230, g859, g25223, g863, g25231, g864,
         g25240, g862, g25232, g866, g25241, g867, g25248, g865, g30269, g873,
         g30277, g876, g30285, g879, g30643, g918, g30648, g921, g30654,
         g30676, g882, g30681, g885, g30687, g888, g30649, g927, g30655, g930,
         g30662, g933, g30286, g891, g30293, g894, g30298, g897, g30259, g936,
         g30264, g939, g30270, g942, g30247, g900, g30249, g903, g30251, g906,
         g30265, g30271, g948, g30278, g951, g30638, g909, g30642, g912,
         g30647, g915, g30670, g954, g30677, g957, g30682, g960, g25042, g780,
         g25935, g776, g26530, g771, g27123, g767, g27603, g762, g28146, g758,
         g28635, g753, g29110, g29354, g29580, g740, g868, g869, n4363, n4364,
         g1088, n4381, g996, n4387, g27257, g1041, g27262, g1030, g27270,
         g1033, g27263, g1056, g27271, g1045, g27282, g1048, g27272, g27283,
         g1060, g27297, g1063, g27284, g1085, g27298, g1075, g27313, g1078,
         g28738, g1095, g28746, g1098, g28758, g1101, g29198, g1104, g29204,
         g1107, g29209, g1110, g28747, g1114, g28759, g1115, g28767, g1113,
         g26806, g1116, g26809, g26813, g1122, g26810, g1125, g26814, g1128,
         g26818, g1131, g27761, g1135, g27763, g1136, g27765, g1134, g29609,
         g999, g29612, g1000, g29616, g1001, g30701, g1002, g30703, g1003,
         g30705, g1004, g30470, g1005, g30485, g1006, g30500, g29170, g1009,
         g29173, g1010, g29179, g1008, g26661, g1090, g26665, g1091, g26669,
         g1089, g1137, n8027, DFF_649_n1, g1139, n8026, DFF_651_n1, g1141,
         n8025, DFF_653_n1, g967, n8024, DFF_655_n1, g969, DFF_657_n1, g971,
         n8021, DFF_659_n1, g973, n8020, DFF_661_n1, g975, n8019, DFF_663_n1,
         g977, n8018, n4486, n4283, g986, n4432, g992, n4277, n8017, g1029,
         g1036, g1037, g1038, g1040, g1044, g1051, g1052, g1053, g1054, g1055,
         g1059, g1066, g1067, g1068, g1069, g1070, g1074, g1081, g1083, g1084,
         g1011, g1024, n4371, n4316, g1236, n4300, g21843, g1240, g18707,
         g1243, n4353, g18763, g1196, n4304, g1199, g1209, g1210, g1142, g1255,
         g1145, g1256, g1257, g1148, g1258, g1259, g1152, g1260, g1251, g1155,
         g1252, g1253, g1158, g1254, g1176, n4460, n4459, g1172, n4465, g23081,
         g1173, g23111, g23126, g1175, g23392, g23406, g24179, g24181, g1164,
         g24213, g1165, g24223, g1166, g23110, g1167, g23014, g1171, g23039,
         g1151, g24212, g24222, g24235, g1214, g1221, g13155, g1229, n4549,
         n4361, g13124, g1235, g1186, n4548, g13171, g1244, g1245, g27273,
         g1262, g27285, g1263, g27299, g1261, g27286, g1265, g27300, g1266,
         g27314, g1264, g27301, g1268, g27315, g1269, g27328, g27316, g1271,
         g27329, g1272, g27339, g1270, g24501, g1273, g24510, g1276, g24521,
         g1279, g24511, g1282, g24522, g1285, g24532, g1288, g28351, g1300,
         g28355, g1303, g28360, g1306, g28346, g1291, g28350, g1294, g28354,
         g1297, g26547, g26557, g1180, g26569, g1183, g1192, n4454, g22615,
         n8009, DFF_783_n1, DFF_792_n1, g1211, n8008, n8007, n8006, n8005,
         n8004, n8003, g1222, g1223, g24072, g1224, n4489, n4358, g1315, n4294,
         g16671, g1316, g20333, g1345, g20717, g1326, n4402, g21969, g1319,
         n4476, g23329, g1339, n4421, g24430, g1332, n4412, g25189, g1346,
         n4401, g26666, g1358, n4411, g26781, g1352, n4469, g27678, g1365,
         n4475, g27718, g1372, n4395, g28321, g1378, n4417, g20882, g20896,
         g1386, g20910, g1384, g20897, g1388, g20911, g1389, g20925, g1387,
         g20912, g1391, g20926, g1392, g20949, g1390, g20927, g1394, g20950,
         g1395, g20972, g1393, g20951, g1397, g20973, g1398, g20993, g1396,
         g20974, g1400, g20994, g21015, g1399, g20995, g1403, g21016, g1404,
         g21033, g1402, g21017, g1406, g21034, g1407, g21052, g1405, g21035,
         g1409, g21053, g1410, g21070, g1408, g20883, g1412, g20898, g1413,
         g20913, g1411, g20952, g1415, g20975, g1416, g20996, g20976, g1418,
         g20997, g1419, g21018, g1417, g25263, g1421, g25267, g1422, g25270,
         g1420, g22234, g1424, g22247, g1425, g22263, g1423, n4317, n4515,
         g1547, n4368, g22149, g1512, g22166, g1513, g22178, g1511, g22167,
         g22179, g1516, g22191, g1514, g22035, g1524, g22043, g1525, g22057,
         g1523, g22044, g1527, g22058, g1528, g22073, g1526, g22059, g1530,
         g22074, g1531, g22090, g1529, g22075, g1533, g22091, g1534, g22112,
         g1532, g22092, g1536, g22113, g22130, g1535, g22114, g1539, g22131,
         g1540, g22150, g1538, g22132, g1542, g22151, g1543, g22168, g1541,
         g22152, g1545, g22169, g1546, g22180, g1544, g25217, g1551, g25224,
         g1552, g25233, g1550, g25225, g1554, g25234, g1555, g25242, g25235,
         g1557, g25243, g1558, g25249, g1556, g25244, g1560, g25250, g1561,
         g25255, g1559, g30279, g1567, g30287, g1570, g30294, g1573, g30651,
         g1612, g30657, g1615, g30663, g1618, g30683, g1576, g30688, g1579,
         g30692, g1582, g30658, g30664, g1624, g30671, g1627, g30295, g1585,
         g30299, g1588, g30302, g1591, g30266, g1630, g30272, g1633, g30280,
         g1636, g30250, g1594, g30252, g1597, g30255, g1600, g30273, g1639,
         g30281, g1642, g30288, g1645, g30644, g1603, g30650, g30656, g1609,
         g30678, g1648, g30684, g1651, g30689, g1654, g25056, g1466, g25938,
         g1462, g26531, g1457, g27129, g1453, g27612, g1448, g28147, g1444,
         g28636, g1439, g29111, g1435, g29355, g29581, g1426, g1562, g1563,
         n4518, g1690, n4386, g27264, g1735, g27274, g1724, g27287, g1727,
         g27275, g1750, g27288, g1739, g27302, g1742, g27289, g1765, g27303,
         g1754, g27317, g1757, g27304, g1779, g27318, g27330, g1772, g28749,
         g1789, g28760, g1792, g28771, g1795, g29205, g1798, g29212, g1801,
         g29218, g1804, g28761, g1808, g28772, g1809, g28778, g1807, g26811,
         g1810, g26815, g1813, g26820, g1816, g26816, g1819, g26821, g1822,
         g26824, g27764, g1829, g27766, g1830, g27768, g1828, g29613, g1693,
         g29617, g1694, g29620, g1695, g30704, g1696, g30706, g1697, g30708,
         g1698, g30487, g1699, g30503, g1700, g30338, g1701, g29178, g1703,
         g29181, g1704, g29184, g1702, g26667, g26670, g1785, g26675, g1783,
         g1831, n7988, DFF_999_n1, g1833, n7987, DFF_1001_n1, g1835, n7986,
         DFF_1003_n1, g1661, n7985, DFF_1005_n1, g1663, n7984, DFF_1007_n1,
         g1665, n7983, DFF_1009_n1, g1667, DFF_1011_n1, g1669, n7980,
         DFF_1013_n1, g1671, n7979, n4484, n4284, g1680, n4488, g1686, n4276,
         n7978, g1723, g1730, g1731, g1732, g1733, g1734, g1738, g1745, g1747,
         g1748, g1749, g1753, g1760, g1761, g1762, g1763, g1764, g1768, g1775,
         g1776, g1777, g1778, g1705, g1718, n4296, n4315, g1930, n4366, g21845,
         g1934, g18743, g1937, n4311, g18794, g1890, n4297, g1893, g1903,
         g1904, g1836, g1944, g1949, g1950, g1951, g1842, g1953, g1846, g1954,
         g1945, g1849, g1946, g1947, g1852, g1948, g1870, n4458, n4457, g1866,
         n4464, g23097, g1867, g23124, g1868, g23137, g1869, g23400, g23413,
         g24182, g24208, g1858, g24219, g1859, g24231, g1860, g23123, g1861,
         g23030, g1865, g23058, g1845, g24218, g24230, g24243, g1908, g1915,
         g1922, g13164, g1923, DFF_1099_n1, n7971, DFF_1100_n1, g13135, g1929,
         g1880, n4545, g13182, g1938, g1939, g27290, g1956, g27305, g1957,
         g27319, g1955, g27306, g1959, g27320, g1960, g27331, g1958, g27321,
         g1962, g27332, g1963, g27340, g1961, g27333, g27341, g1966, g27346,
         g1964, g24513, g1967, g24524, g1970, g24534, g1973, g24525, g1976,
         g24535, g1979, g24545, g1982, g28357, g1994, g28362, g1997, g28366,
         g2000, g28352, g1985, g28356, g1988, g28361, g1991, g26559, g26573,
         g1874, g26592, g1877, g1886, n4493, g22651, n7968, DFF_1133_n1,
         DFF_1142_n1, g1905, n7967, n7966, n7965, n7964, n7963, n7962, g1916,
         g1917, g24083, n7960, n4357, g2009, n4293, g16692, g2010, g20353,
         g2039, g20752, g2020, n4400, g21972, g2013, n4474, g23339, g2033,
         n4420, g24434, g2026, n4410, g25194, g2040, n4399, g26671, g2052,
         n4409, g26789, g2046, n4468, g27682, g2059, n4473, g27722, g28325,
         g2072, n4416, g20899, g2079, g20915, g2080, g20934, g2078, g20916,
         g2082, g20935, g2083, g20953, g2081, g20936, g2085, g20954, g2086,
         g20977, g2084, g20955, g2088, g20978, g2089, g20999, g2087, g20979,
         g2091, g21000, g21019, g2090, g21001, g2094, g21020, g2095, g21039,
         g2093, g21021, g2097, g21040, g2098, g21054, g2096, g21041, g2100,
         g21055, g2101, g21071, g2099, g21056, g2103, g21072, g2104, g21080,
         g2102, g20900, g2106, g20917, g20937, g2105, g20980, g2109, g21002,
         g2110, g21022, g2108, g21003, g2112, g21023, g2113, g21042, g2111,
         g25268, g2115, g25271, g2116, g25279, g2114, g22249, g2118, g22267,
         g2119, g22280, g2117, n4324, g2241, n4367, g22170, g2206, g22182,
         g2207, g22192, g2205, g22183, g2209, g22193, g2210, g22200, g2208,
         g22045, g2218, g22060, g2219, g22076, g2217, g22061, g2221, g22077,
         g2222, g22097, g2220, g22078, g2224, g22098, g22115, g2223, g22099,
         g2227, g22116, g2228, g22138, g2226, g22117, g2230, g22139, g2231,
         g22153, g2229, g22140, g2233, g22154, g2234, g22171, g2232, g22155,
         g2236, g22172, g2237, g22184, g2235, g22173, g2239, g22185, g22194,
         g2238, g25227, g2245, g25236, g2246, g25245, g2244, g25237, g2248,
         g25246, g2249, g25251, g2247, g25247, g2251, g25252, g2252, g25256,
         g2250, g25253, g2254, g25257, g2255, g25259, g2253, g30289, g2261,
         g30296, g30300, g2267, g30660, g2306, g30666, g2309, g30672, g2312,
         g30690, g2270, g30693, g2273, g30695, g2276, g30667, g2315, g30673,
         g2318, g30679, g2321, g30301, g2279, g30303, g2282, g30304, g2285,
         g30274, g2324, g30282, g30290, g2330, g30253, g2288, g30256, g2291,
         g30260, g2294, g30283, g2333, g30291, g2336, g30297, g2339, g30652,
         g2297, g30659, g2300, g30665, g2303, g30686, g2342, g30691, g2345,
         g30694, g2348, g25067, g2160, g25940, g26532, g2151, g27131, g2147,
         g27621, g2142, g28148, g2138, g28637, g2133, g29112, g2129, g29357,
         g29582, g2120, g2256, g2257, n4516, g27276, g2429, g27291, g2418,
         g27307, g2421, g27292, g2444, g27308, g2433, g27322, g2436, g27309,
         g2459, g27323, g2448, g27334, g2451, g27324, g2473, g27335, g2463,
         g27342, g2466, g28763, g2483, g28773, g2486, g28782, g29213, g2492,
         g29221, g2495, g29226, g2498, g28774, g2502, g28783, g2503, g28788,
         g2501, g26817, g2504, g26822, g2507, g26825, g2510, g26823, g2513,
         g26826, g2516, g26827, g2519, g27767, g2523, g27769, g2524, g27771,
         g29618, g2387, g29621, g2388, g29623, g2389, g30707, g2390, g30709,
         g2391, g30566, g2392, g30505, g2393, g30341, g2394, g30356, g2395,
         g29182, g2397, g29185, g2398, g29187, g2396, g26672, g2478, g26676,
         g2479, g26025, g2525, n7946, DFF_1349_n1, g2527, n7945, DFF_1351_n1,
         g2529, n7944, DFF_1353_n1, g2355, n7943, DFF_1355_n1, g2357, n7942,
         DFF_1357_n1, g2359, n7941, DFF_1359_n1, g2361, n7940, DFF_1361_n1,
         n7938, DFF_1363_n1, g2365, n7937, n4483, n4285, g2374, n4487, g30055,
         g2380, n4275, n7936, DFF_1378_n1, g2417, g2424, g2425, g2426, g2427,
         g2428, g2432, g2439, g2441, g2442, g2443, g2447, g2454, g2455, g2456,
         g2457, g2458, g2462, g2469, g2470, g2471, g2472, g2412, n4314, n4370,
         g2624, n4299, g21847, g2628, g18780, g2631, n4352, g18820, g2584,
         n4303, g2587, g2597, g2598, g2530, g2638, g2643, g2533, g2645, g2536,
         g2646, g2647, g2540, g2648, g2639, g2543, g2640, g2641, g2546, g2642,
         g2564, n4456, n4455, g2560, n4463, g23114, g2561, g23133, g2562,
         g21970, g23407, g23418, g24209, g24214, g2552, g24226, g2553, g24238,
         g2554, g23132, g2555, g23047, g2559, g23076, g2539, g24225, g24237,
         g24250, g2602, g2609, g13175, g2617, n7930, g30072, n7929, g13143,
         g2623, g2574, n4543, g13194, g2632, g2633, g27310, g2650, g27325,
         g2651, g27336, g2649, g27326, g2653, g27337, g2654, g27343, g2652,
         g27338, g2656, g27344, g27347, g2655, g27345, g2659, g27348, g2660,
         g27354, g2658, g24527, g2661, g24537, g2664, g24547, g2667, g24538,
         g2670, g24548, g2673, g24557, g2676, g28364, g2688, g28368, g2691,
         g28371, g2694, g28358, g2679, g28363, g28367, g2685, g26575, g2565,
         g26596, g2568, g26616, g2571, g2580, g22687, n7926, g30061, g2599,
         n7925, n7924, n7923, n7922, n7921, n7920, g2611, g24092, g2612, n4490,
         n7918, n4356, g2703, n4292, g16718, g2704, g20375, g2733, g20789,
         g2714, n4398, g21974, g2707, n4472, g23348, g2727, n4419, g24438,
         g2720, n4408, g25197, g2734, n4397, g26677, g2746, n4407, g26795,
         g27243, g2753, n4471, g27724, g2760, n4393, g28328, g2766, n4415,
         g20918, g2773, g20939, g2774, g20962, g2772, g20940, g2776, g20963,
         g2777, g20981, g2775, g20964, g2779, g20982, g2780, g21004, g2778,
         g20983, g2782, g21005, g2783, g21025, g21006, g2785, g21026, g2786,
         g21043, g2784, g21027, g2788, g21044, g2789, g21060, g2787, g21045,
         g2791, g21061, g2792, g21073, g2790, g21062, g2794, g21074, g2795,
         g21081, g2793, g21075, g2797, g21082, g2798, g21094, g20919, g2800,
         g20941, g2801, g20965, g2799, g21007, g2803, g21028, g2804, g21046,
         g2802, g21029, g2806, g21047, g2807, g21063, g2805, g25272, g2809,
         g25280, g2810, g25288, g2808, g22269, g2812, g22284, g2813, g22299,
         g20877, n7913, g20884, n7912, n4263, n4269, g3043, n4268, g3044,
         n4267, g3045, n4266, g3046, n4265, g3047, n4272, g3048, n4271, g3049,
         n4270, g3050, n4259, g3051, n4236, g3052, n4239, g3053, n4237, n4234,
         g3056, n4233, g3057, n4238, g3058, n4235, g3059, n4240, g3060, n4232,
         g3061, n4245, g3062, n4248, g3063, n4246, g3064, n4243, g3065, n4242,
         g3066, n4247, g3067, n4244, g3068, n4249, g3069, n4241, n4254, g3071,
         n4257, g3072, n4255, g3073, n4252, g3074, n4251, g3075, n4256, g3076,
         n4253, g3077, n4258, g3078, n4250, g2997, g25265, g2993, g26048,
         n7909, g23330, g3006, g24445, g3002, g25191, g3013, g26031, g26786,
         g3024, n4262, g3018, n4481, g23359, g3028, n4350, g24446, g3036,
         n4480, g25202, g3032, n7907, DFF_1612_n1, g2987, n4365, g16824,
         g16844, g16853, g16860, g16803, DFF_1618_n1, g16835, g16851, g16857,
         g16866, g3083, n4261, N995, n4577, g16845, g16854, g16861, g16880,
         DFF_1628_n1, g18755, g18804, g18837, g18868, g18907, g2990, N690,
         n4578, n4260, n4309, n4308, n4307, n4306, n4524, n4525, n4511, n4509,
         n4499, n4520, n3683, n3887, n3686, n3890, n3692, n3896, n4513, n3897,
         n3424, n3427, n3433, n4529, n4530, n4522, n4523, n4521, n3171, n3159,
         n3163, n3893, n3689, n3430, n4527, n4528, n4526, n3167, n3894, n3888,
         n3891, n2302, n2289, n2303, n2275, n4066, n4065, n4606, n4618, n4640,
         n2489, n2542, n2617, n2279, n2207, n2381, n2309, n2237, n2459, n3936,
         n3260, n3252, n3254, n3301, n3293, n3341, n3334, n3380, n4102, n3374,
         n3038, n3070, n3102, n3130, n2800, n2798, n2616, n2594, n3940, n3705,
         n3933, n3939, n3700, n4058, n4123, n4101, n4182, n4073, n4057,
         n4122_Tj_Payload, n4122, n4160_Tj_Payload, n4149_Tj_Payload, n4149,
         n4161_Tj_Payload, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4, Tj_OUT1234,
         Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678, Tj_Trigger, n8, n122,
         n282, n305, n306, n308, n312, n338, n405, n407, n465, n467, n484,
         n486, n488, n490, n492, n515, n516, n517, n519, n590, n640, n710,
         n712, n714, n716, n785, n811, n869, n932, n1003, n1005, n1073, n1096,
         n1221, n1289, n1291, n1348, n1359, n1386, n8268, n8269, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8545, n8546, n8602,
         n8627, n8630, n8631, n8632, n8633, n8634, n8652, n8655, n8656, n8657,
         n8658, n8659, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8824, n8825, n8826, n8827, n8828, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8983, n8984, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n9012, n9013, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9063, n9065, n9067, n9068, n9069,
         n9071, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, U4467_n1, U4904_n1, U4930_n1, U5128_n1, U5141_n1,
         U5749_n1, U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1, U5755_n1,
         U5756_n1, U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1, U5762_n1,
         U5763_n1, U5764_n1, U5882_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1,
         U6140_n1, U6460_n1, U6470_n1, U6562_n1, U6563_n1, U6718_n1, U7116_n1,
         U7118_n1, U7293_n1;
  assign g8251 = test_so3;
  assign g7519 = test_so4;
  assign g4450 = test_so5;
  assign g7909 = test_so23;
  assign g5612 = test_so57;
  assign g5695 = test_so63;
  assign g7084 = test_so73;
  assign g8270 = test_so99;
  assign g8258 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(g51), .SI(test_si1), .SE(n9132), .CLK(n9319), .Q(
        n8104), .QN(n16489) );
  SDFFX1 DFF_1_Q_reg ( .D(g16802), .SI(n8104), .SE(n9132), .CLK(n9319), .Q(
        n8103) );
  SDFFX1 DFF_2_Q_reg ( .D(g16823), .SI(n8103), .SE(n9132), .CLK(n9319), .Q(
        n8102), .QN(DFF_2_n1) );
  SDFFX1 DFF_3_Q_reg ( .D(n4264), .SI(n8102), .SE(n9132), .CLK(n9319), .Q(
        g2950), .QN(n4423) );
  SDFFX1 DFF_4_Q_reg ( .D(n4274), .SI(g2950), .SE(n9133), .CLK(n9320), .Q(
        g2883), .QN(n4330) );
  SDFFX1 DFF_5_Q_reg ( .D(g22026), .SI(g2883), .SE(n9133), .CLK(n9320), .Q(
        g2888), .QN(n9081) );
  SDFFX1 DFF_6_Q_reg ( .D(g23358), .SI(g2888), .SE(n9157), .CLK(n9344), .Q(
        g2896), .QN(n4431) );
  SDFFX1 DFF_7_Q_reg ( .D(g24473), .SI(g2896), .SE(n9157), .CLK(n9344), .Q(
        g2892), .QN(n9102) );
  SDFFX1 DFF_8_Q_reg ( .D(g25201), .SI(g2892), .SE(n9157), .CLK(n9344), .Q(
        g2903), .QN(n4305) );
  SDFFX1 DFF_9_Q_reg ( .D(g26037), .SI(g2903), .SE(n9157), .CLK(n9344), .Q(
        g2900), .QN(n4291) );
  SDFFX1 DFF_10_Q_reg ( .D(g26798), .SI(g2900), .SE(n9157), .CLK(n9344), .Q(
        g2908), .QN(n4355) );
  SDFFX1 DFF_11_Q_reg ( .D(n8), .SI(g2908), .SE(n9157), .CLK(n9344), .Q(g2912), 
        .QN(n4482) );
  SDFFX1 DFF_12_Q_reg ( .D(g23357), .SI(g2912), .SE(n9158), .CLK(n9345), .Q(
        g2917), .QN(n4479) );
  SDFFX1 DFF_13_Q_reg ( .D(g24476), .SI(g2917), .SE(n9158), .CLK(n9345), .Q(
        g2924), .QN(n4349) );
  SDFFX1 DFF_14_Q_reg ( .D(g25199), .SI(g2924), .SE(n9158), .CLK(n9345), .Q(
        g2920), .QN(n8822) );
  SDFFX1 DFF_15_Q_reg ( .D(n4280), .SI(g2920), .SE(n9158), .CLK(n9345), .Q(
        test_so1) );
  SDFFX1 DFF_16_Q_reg ( .D(n4281), .SI(test_si2), .SE(n9130), .CLK(n9317), .Q(
        n8099) );
  SDFFX1 DFF_17_Q_reg ( .D(g51), .SI(n8099), .SE(n9130), .CLK(n9317), .Q(g8021) );
  SDFFX1 DFF_18_Q_reg ( .D(g8021), .SI(g8021), .SE(n9130), .CLK(n9317), .Q(
        n8098), .QN(DFF_18_n1) );
  SDFFX1 DFF_19_Q_reg ( .D(n4279), .SI(n8098), .SE(n9130), .CLK(n9317), .Q(
        g2879), .QN(n4351) );
  SDFFX1 DFF_20_Q_reg ( .D(g3212), .SI(g2879), .SE(n9130), .CLK(n9317), .Q(
        g2934) );
  SDFFX1 DFF_21_Q_reg ( .D(g3228), .SI(g2934), .SE(n9130), .CLK(n9317), .Q(
        g2935), .QN(n9061) );
  SDFFX1 DFF_22_Q_reg ( .D(g3227), .SI(g2935), .SE(n9131), .CLK(n9318), .Q(
        g2938) );
  SDFFX1 DFF_23_Q_reg ( .D(g3226), .SI(g2938), .SE(n9131), .CLK(n9318), .Q(
        g2941), .QN(n9059) );
  SDFFX1 DFF_24_Q_reg ( .D(g3225), .SI(g2941), .SE(n9131), .CLK(n9318), .Q(
        g2944), .QN(n9065) );
  SDFFX1 DFF_25_Q_reg ( .D(g3224), .SI(g2944), .SE(n9131), .CLK(n9318), .Q(
        g2947), .QN(n9063) );
  SDFFX1 DFF_26_Q_reg ( .D(g3223), .SI(g2947), .SE(n9131), .CLK(n9318), .Q(
        g2953) );
  SDFFX1 DFF_27_Q_reg ( .D(g3222), .SI(g2953), .SE(n9131), .CLK(n9318), .Q(
        g2956) );
  SDFFX1 DFF_28_Q_reg ( .D(g3221), .SI(g2956), .SE(n9131), .CLK(n9318), .Q(
        g2959), .QN(n9060) );
  SDFFX1 DFF_29_Q_reg ( .D(g3232), .SI(g2959), .SE(n9131), .CLK(n9318), .Q(
        g2962), .QN(n9079) );
  SDFFX1 DFF_30_Q_reg ( .D(g3220), .SI(g2962), .SE(n9131), .CLK(n9318), .Q(
        g2963), .QN(n9069) );
  SDFFX1 DFF_31_Q_reg ( .D(g3219), .SI(g2963), .SE(n9131), .CLK(n9318), .Q(
        test_so2) );
  SDFFX1 DFF_32_Q_reg ( .D(g3218), .SI(test_si3), .SE(n9130), .CLK(n9317), .Q(
        g2969) );
  SDFFX1 DFF_33_Q_reg ( .D(g3217), .SI(g2969), .SE(n9130), .CLK(n9317), .Q(
        g2972) );
  SDFFX1 DFF_34_Q_reg ( .D(g3216), .SI(g2972), .SE(n9130), .CLK(n9317), .Q(
        g2975), .QN(n9071) );
  SDFFX1 DFF_35_Q_reg ( .D(g3215), .SI(g2975), .SE(n9130), .CLK(n9317), .Q(
        g2978), .QN(n9067) );
  SDFFX1 DFF_36_Q_reg ( .D(g3214), .SI(g2978), .SE(n9130), .CLK(n9317), .Q(
        g2981) );
  SDFFX1 DFF_37_Q_reg ( .D(g3213), .SI(g2981), .SE(n9130), .CLK(n9317), .Q(
        g2874), .QN(n9068) );
  SDFFX1 DFF_38_Q_reg ( .D(g18754), .SI(g2874), .SE(n9131), .CLK(n9318), .Q(
        g1506), .QN(n4288) );
  SDFFX1 DFF_39_Q_reg ( .D(g18781), .SI(g1506), .SE(n9131), .CLK(n9318), .Q(
        g1501), .QN(n4565) );
  SDFFX1 DFF_40_Q_reg ( .D(g18803), .SI(g1501), .SE(n9132), .CLK(n9319), .Q(
        g1496), .QN(n4557) );
  SDFFX1 DFF_41_Q_reg ( .D(g18821), .SI(g1496), .SE(n9132), .CLK(n9319), .Q(
        g1491), .QN(n4326) );
  SDFFX1 DFF_42_Q_reg ( .D(g18835), .SI(g1491), .SE(n9132), .CLK(n9319), .Q(
        g1486), .QN(n4390) );
  SDFFX1 DFF_43_Q_reg ( .D(g18852), .SI(g1486), .SE(n9132), .CLK(n9319), .Q(
        g1481), .QN(n4320) );
  SDFFX1 DFF_44_Q_reg ( .D(g18866), .SI(g1481), .SE(n9132), .CLK(n9319), .Q(
        g1476), .QN(n4374) );
  SDFFX1 DFF_45_Q_reg ( .D(g18883), .SI(g1476), .SE(n9132), .CLK(n9319), .Q(
        g1471), .QN(n4378) );
  SDFFX1 DFF_46_Q_reg ( .D(g21880), .SI(g1471), .SE(n9138), .CLK(n9325), .Q(
        g2877) );
  SDFFX1 DFF_47_Q_reg ( .D(g19154), .SI(g2877), .SE(n9139), .CLK(n9326), .Q(
        test_so3) );
  SDFFX1 DFF_48_Q_reg ( .D(test_so3), .SI(test_si4), .SE(n9139), .CLK(n9326), 
        .Q(g813), .QN(n4289) );
  SDFFX1 DFF_49_Q_reg ( .D(g19163), .SI(g813), .SE(n9139), .CLK(n9326), .Q(
        g4090) );
  SDFFX1 DFF_50_Q_reg ( .D(g4090), .SI(g4090), .SE(n9139), .CLK(n9326), .Q(
        g809), .QN(n4567) );
  SDFFX1 DFF_51_Q_reg ( .D(g19173), .SI(g809), .SE(n9139), .CLK(n9326), .Q(
        g4323) );
  SDFFX1 DFF_52_Q_reg ( .D(g4323), .SI(g4323), .SE(n9139), .CLK(n9326), .Q(
        g805), .QN(n4559) );
  SDFFX1 DFF_53_Q_reg ( .D(g19184), .SI(g805), .SE(n9139), .CLK(n9326), .Q(
        g4590) );
  SDFFX1 DFF_54_Q_reg ( .D(g4590), .SI(g4590), .SE(n9139), .CLK(n9326), .Q(
        g801), .QN(n4327) );
  SDFFX1 DFF_55_Q_reg ( .D(g20310), .SI(g801), .SE(n9139), .CLK(n9326), .Q(
        g6225) );
  SDFFX1 DFF_56_Q_reg ( .D(g6225), .SI(g6225), .SE(n9139), .CLK(n9326), .Q(
        g797), .QN(n4391) );
  SDFFX1 DFF_57_Q_reg ( .D(g20343), .SI(g797), .SE(n9139), .CLK(n9326), .Q(
        g6442) );
  SDFFX1 DFF_58_Q_reg ( .D(g6442), .SI(g6442), .SE(n9139), .CLK(n9326), .Q(
        g793), .QN(n4321) );
  SDFFX1 DFF_59_Q_reg ( .D(g20376), .SI(g793), .SE(n9140), .CLK(n9327), .Q(
        g6895) );
  SDFFX1 DFF_60_Q_reg ( .D(g6895), .SI(g6895), .SE(n9140), .CLK(n9327), .Q(
        g789), .QN(n4375) );
  SDFFX1 DFF_61_Q_reg ( .D(g20417), .SI(g789), .SE(n9140), .CLK(n9327), .Q(
        g7334) );
  SDFFX1 DFF_62_Q_reg ( .D(g7334), .SI(g7334), .SE(n9140), .CLK(n9327), .Q(
        g785), .QN(n4379) );
  SDFFX1 DFF_63_Q_reg ( .D(g21878), .SI(g785), .SE(n9140), .CLK(n9327), .Q(
        test_so4) );
  SDFFX1 DFF_64_Q_reg ( .D(test_so4), .SI(test_si5), .SE(n9140), .CLK(n9327), 
        .Q(g2873) );
  SDFFX1 DFF_65_Q_reg ( .D(g19153), .SI(g2873), .SE(n9141), .CLK(n9328), .Q(
        g8249) );
  SDFFX1 DFF_66_Q_reg ( .D(g8249), .SI(g8249), .SE(n9141), .CLK(n9328), .Q(
        g125), .QN(n4290) );
  SDFFX1 DFF_67_Q_reg ( .D(g19162), .SI(g125), .SE(n9141), .CLK(n9328), .Q(
        g4088) );
  SDFFX1 DFF_68_Q_reg ( .D(g4088), .SI(g4088), .SE(n9141), .CLK(n9328), .Q(
        g121), .QN(n4569) );
  SDFFX1 DFF_69_Q_reg ( .D(g19172), .SI(g121), .SE(n9141), .CLK(n9328), .Q(
        g4321) );
  SDFFX1 DFF_70_Q_reg ( .D(g4321), .SI(g4321), .SE(n9141), .CLK(n9328), .Q(
        g117), .QN(n4561) );
  SDFFX1 DFF_71_Q_reg ( .D(g19144), .SI(g117), .SE(n9141), .CLK(n9328), .Q(
        g8023) );
  SDFFX1 DFF_72_Q_reg ( .D(g8023), .SI(g8023), .SE(n9141), .CLK(n9328), .Q(
        g113), .QN(n4328) );
  SDFFX1 DFF_73_Q_reg ( .D(g19149), .SI(g113), .SE(n9141), .CLK(n9328), .Q(
        g8175) );
  SDFFX1 DFF_74_Q_reg ( .D(g8175), .SI(g8175), .SE(n9141), .CLK(n9328), .Q(
        g109), .QN(n4392) );
  SDFFX1 DFF_75_Q_reg ( .D(g19157), .SI(g109), .SE(n9142), .CLK(n9329), .Q(
        g3993) );
  SDFFX1 DFF_76_Q_reg ( .D(g3993), .SI(g3993), .SE(n9142), .CLK(n9329), .Q(
        g105), .QN(n4322) );
  SDFFX1 DFF_77_Q_reg ( .D(g19167), .SI(g105), .SE(n9142), .CLK(n9329), .Q(
        g4200) );
  SDFFX1 DFF_78_Q_reg ( .D(g4200), .SI(g4200), .SE(n9142), .CLK(n9329), .Q(
        g101), .QN(n4376) );
  SDFFX1 DFF_79_Q_reg ( .D(g19178), .SI(g101), .SE(n9142), .CLK(n9329), .Q(
        test_so5) );
  SDFFX1 DFF_80_Q_reg ( .D(test_so5), .SI(test_si6), .SE(n9142), .CLK(n9329), 
        .Q(g97), .QN(n4380) );
  SDFFX1 DFF_81_Q_reg ( .D(g20874), .SI(g97), .SE(n9142), .CLK(n9329), .Q(
        g8096) );
  SDFFX1 DFF_82_Q_reg ( .D(g8096), .SI(g8096), .SE(n9142), .CLK(n9329), .Q(
        g2857) );
  SDFFX1 DFF_83_Q_reg ( .D(g18885), .SI(g2857), .SE(n9142), .CLK(n9329), .Q(
        g2200), .QN(n4287) );
  SDFFX1 DFF_84_Q_reg ( .D(g18975), .SI(g2200), .SE(n9142), .CLK(n9329), .Q(
        g2195), .QN(n4563) );
  SDFFX1 DFF_85_Q_reg ( .D(g18968), .SI(g2195), .SE(n9142), .CLK(n9329), .Q(
        g2190), .QN(n4555) );
  SDFFX1 DFF_86_Q_reg ( .D(g18942), .SI(g2190), .SE(n9142), .CLK(n9329), .Q(
        g2185), .QN(n4325) );
  SDFFX1 DFF_87_Q_reg ( .D(g18906), .SI(g2185), .SE(n9143), .CLK(n9330), .Q(
        g2180), .QN(n4389) );
  SDFFX1 DFF_88_Q_reg ( .D(g18867), .SI(g2180), .SE(n9143), .CLK(n9330), .Q(
        g2175), .QN(n4319) );
  SDFFX1 DFF_89_Q_reg ( .D(g18836), .SI(g2175), .SE(n9143), .CLK(n9330), .Q(
        g2170), .QN(n4373) );
  SDFFX1 DFF_90_Q_reg ( .D(g18957), .SI(g2170), .SE(n9143), .CLK(n9330), .Q(
        g2165), .QN(n4377) );
  SDFFX1 DFF_91_Q_reg ( .D(g21882), .SI(g2165), .SE(n9149), .CLK(n9336), .Q(
        g2878) );
  SDFFX1 DFF_92_Q_reg ( .D(n4598), .SI(g2878), .SE(n9255), .CLK(n9442), .Q(
        g8106), .QN(n4382) );
  SDFFX1 DFF_93_Q_reg ( .D(g8106), .SI(g8106), .SE(n9256), .CLK(n9443), .Q(
        g8030), .QN(n4383) );
  SDFFX1 DFF_94_Q_reg ( .D(g8030), .SI(g8030), .SE(n9256), .CLK(n9443), .Q(
        g3109), .QN(n4494) );
  SDFFX1 DFF_95_Q_reg ( .D(g18669), .SI(g3109), .SE(n9257), .CLK(n9444), .Q(
        test_so6) );
  SDFFX1 DFF_96_Q_reg ( .D(g18719), .SI(test_si7), .SE(n9256), .CLK(n9443), 
        .Q(g3211) );
  SDFFX1 DFF_97_Q_reg ( .D(g18782), .SI(g3211), .SE(n9256), .CLK(n9443), .Q(
        g3084) );
  SDFFX1 DFF_98_Q_reg ( .D(g17222), .SI(g3084), .SE(n9256), .CLK(n9443), .Q(
        g3085) );
  SDFFX1 DFF_99_Q_reg ( .D(g17225), .SI(g3085), .SE(n9256), .CLK(n9443), .Q(
        g3086) );
  SDFFX1 DFF_100_Q_reg ( .D(g17234), .SI(g3086), .SE(n9256), .CLK(n9443), .Q(
        g3087) );
  SDFFX1 DFF_101_Q_reg ( .D(g17224), .SI(g3087), .SE(n9256), .CLK(n9443), .Q(
        g3091) );
  SDFFX1 DFF_102_Q_reg ( .D(g17228), .SI(g3091), .SE(n9256), .CLK(n9443), .Q(
        g3092) );
  SDFFX1 DFF_103_Q_reg ( .D(g17246), .SI(g3092), .SE(n9256), .CLK(n9443), .Q(
        g3093) );
  SDFFX1 DFF_104_Q_reg ( .D(g17226), .SI(g3093), .SE(n9256), .CLK(n9443), .Q(
        g3094) );
  SDFFX1 DFF_105_Q_reg ( .D(g17235), .SI(g3094), .SE(n9257), .CLK(n9444), .Q(
        g3095) );
  SDFFX1 DFF_106_Q_reg ( .D(g17269), .SI(g3095), .SE(n9257), .CLK(n9444), .Q(
        g3096) );
  SDFFX1 DFF_107_Q_reg ( .D(g25450), .SI(g3096), .SE(n9257), .CLK(n9444), .Q(
        g3097) );
  SDFFX1 DFF_108_Q_reg ( .D(g25451), .SI(g3097), .SE(n9257), .CLK(n9444), .Q(
        g3098) );
  SDFFX1 DFF_109_Q_reg ( .D(g25452), .SI(g3098), .SE(n9257), .CLK(n9444), .Q(
        g3099) );
  SDFFX1 DFF_110_Q_reg ( .D(g28420), .SI(g3099), .SE(n9257), .CLK(n9444), .Q(
        g3100) );
  SDFFX1 DFF_111_Q_reg ( .D(g28421), .SI(g3100), .SE(n9257), .CLK(n9444), .Q(
        test_so7) );
  SDFFX1 DFF_112_Q_reg ( .D(g28425), .SI(test_si8), .SE(n9256), .CLK(n9443), 
        .Q(g3102) );
  SDFFX1 DFF_113_Q_reg ( .D(g29936), .SI(g3102), .SE(n9258), .CLK(n9445), .Q(
        g3103) );
  SDFFX1 DFF_114_Q_reg ( .D(g29939), .SI(g3103), .SE(n9258), .CLK(n9445), .Q(
        g3104) );
  SDFFX1 DFF_115_Q_reg ( .D(g29941), .SI(g3104), .SE(n9258), .CLK(n9445), .Q(
        g3105) );
  SDFFX1 DFF_116_Q_reg ( .D(g30796), .SI(g3105), .SE(n9258), .CLK(n9445), .Q(
        g3106) );
  SDFFX1 DFF_117_Q_reg ( .D(g30798), .SI(g3106), .SE(n9258), .CLK(n9445), .Q(
        g3107) );
  SDFFX1 DFF_118_Q_reg ( .D(g30801), .SI(g3107), .SE(n9258), .CLK(n9445), .Q(
        g3108) );
  SDFFX1 DFF_119_Q_reg ( .D(g17229), .SI(g3108), .SE(n9258), .CLK(n9445), .Q(
        g3155) );
  SDFFX1 DFF_120_Q_reg ( .D(g17247), .SI(g3155), .SE(n9258), .CLK(n9445), .Q(
        g3158) );
  SDFFX1 DFF_121_Q_reg ( .D(g17302), .SI(g3158), .SE(n9258), .CLK(n9445), .Q(
        g3161) );
  SDFFX1 DFF_122_Q_reg ( .D(g17236), .SI(g3161), .SE(n9258), .CLK(n9445), .Q(
        g3164) );
  SDFFX1 DFF_123_Q_reg ( .D(g17270), .SI(g3164), .SE(n9258), .CLK(n9445), .Q(
        g3167) );
  SDFFX1 DFF_124_Q_reg ( .D(g17340), .SI(g3167), .SE(n9258), .CLK(n9445), .Q(
        g3170) );
  SDFFX1 DFF_125_Q_reg ( .D(g17248), .SI(g3170), .SE(n9259), .CLK(n9446), .Q(
        g3173) );
  SDFFX1 DFF_126_Q_reg ( .D(g17303), .SI(g3173), .SE(n9259), .CLK(n9446), .Q(
        g3176) );
  SDFFX1 DFF_127_Q_reg ( .D(g17383), .SI(g3176), .SE(n9259), .CLK(n9446), .Q(
        test_so8) );
  SDFFX1 DFF_128_Q_reg ( .D(g17271), .SI(test_si9), .SE(n9257), .CLK(n9444), 
        .Q(g3182) );
  SDFFX1 DFF_129_Q_reg ( .D(g17341), .SI(g3182), .SE(n9257), .CLK(n9444), .Q(
        g3185) );
  SDFFX1 DFF_130_Q_reg ( .D(g17429), .SI(g3185), .SE(n9257), .CLK(n9444), .Q(
        g3088) );
  SDFFX1 DFF_131_Q_reg ( .D(g24734), .SI(g3088), .SE(n9257), .CLK(n9444), .Q(
        n8090) );
  SDFFX1 DFF_132_Q_reg ( .D(g25442), .SI(n8090), .SE(n9136), .CLK(n9323), .Q(
        n8089) );
  SDFFX1 DFF_133_Q_reg ( .D(g25435), .SI(n8089), .SE(n9136), .CLK(n9323), .Q(
        g3197) );
  SDFFX1 DFF_134_Q_reg ( .D(g25420), .SI(g3197), .SE(n9136), .CLK(n9323), .Q(
        n8088) );
  SDFFX1 DFF_135_Q_reg ( .D(g26149), .SI(n8088), .SE(n9136), .CLK(n9323), .Q(
        g3201), .QN(n4406) );
  SDFFX1 DFF_136_Q_reg ( .D(g26135), .SI(g3201), .SE(n9136), .CLK(n9323), .Q(
        g3204) );
  SDFFX1 DFF_137_Q_reg ( .D(g26104), .SI(g3204), .SE(n9136), .CLK(n9323), .Q(
        g3207), .QN(n4329) );
  SDFFX1 DFF_138_Q_reg ( .D(g27380), .SI(g3207), .SE(n9136), .CLK(n9323), .Q(
        g3188), .QN(n4405) );
  SDFFX1 DFF_139_Q_reg ( .D(n122), .SI(g3188), .SE(n9136), .CLK(n9323), .Q(
        g3133), .QN(n8545) );
  SDFFX1 DFF_140_Q_reg ( .D(g26104), .SI(g3133), .SE(n9136), .CLK(n9323), .Q(
        n8087) );
  SDFFX1 DFF_141_Q_reg ( .D(n282), .SI(n8087), .SE(n9136), .CLK(n9323), .Q(
        g3128), .QN(n8731) );
  SDFFX1 DFF_142_Q_reg ( .D(g26149), .SI(g3128), .SE(n9136), .CLK(n9323), .Q(
        n8086) );
  SDFFX1 DFF_143_Q_reg ( .D(g25420), .SI(n8086), .SE(n9137), .CLK(n9324), .Q(
        test_so9) );
  SDFFX1 DFF_144_Q_reg ( .D(n308), .SI(test_si10), .SE(n9137), .CLK(n9324), 
        .Q(n8084), .QN(DFF_144_n1) );
  SDFFX1 DFF_145_Q_reg ( .D(g25442), .SI(n8084), .SE(n9137), .CLK(n9324), .Q(
        g3124) );
  SDFFX1 DFF_146_Q_reg ( .D(n312), .SI(g3124), .SE(n9137), .CLK(n9324), .Q(
        n8083), .QN(DFF_146_n1) );
  SDFFX1 DFF_147_Q_reg ( .D(g26104), .SI(n8083), .SE(n9137), .CLK(n9324), .Q(
        n8082) );
  SDFFX1 DFF_148_Q_reg ( .D(g26135), .SI(n8082), .SE(n9137), .CLK(n9324), .Q(
        n8081) );
  SDFFX1 DFF_149_Q_reg ( .D(g26149), .SI(n8081), .SE(n9137), .CLK(n9324), .Q(
        n8080) );
  SDFFX1 DFF_150_Q_reg ( .D(g25420), .SI(n8080), .SE(n9137), .CLK(n9324), .Q(
        g3112) );
  SDFFX1 DFF_151_Q_reg ( .D(g25435), .SI(g3112), .SE(n9137), .CLK(n9324), .Q(
        g3110) );
  SDFFX1 DFF_152_Q_reg ( .D(g25442), .SI(g3110), .SE(n9137), .CLK(n9324), .Q(
        g3111) );
  SDFFX1 DFF_153_Q_reg ( .D(g27380), .SI(g3111), .SE(n9137), .CLK(n9324), .Q(
        n8079), .QN(n16494) );
  SDFFX1 DFF_154_Q_reg ( .D(g26104), .SI(n8079), .SE(n9137), .CLK(n9324), .Q(
        n8078), .QN(n16492) );
  SDFFX1 DFF_155_Q_reg ( .D(g26135), .SI(n8078), .SE(n9138), .CLK(n9325), .Q(
        n8077) );
  SDFFX1 DFF_156_Q_reg ( .D(g26149), .SI(n8077), .SE(n9138), .CLK(n9325), .Q(
        n8076) );
  SDFFX1 DFF_157_Q_reg ( .D(g27380), .SI(n8076), .SE(n9138), .CLK(n9325), .Q(
        g3151), .QN(n4424) );
  SDFFX1 DFF_158_Q_reg ( .D(g26104), .SI(g3151), .SE(n9138), .CLK(n9325), .Q(
        g3142), .QN(n4301) );
  SDFFX1 DFF_159_Q_reg ( .D(g26135), .SI(g3142), .SE(n9138), .CLK(n9325), .Q(
        test_so10), .QN(n9128) );
  SDFFX1 DFF_160_Q_reg ( .D(n122), .SI(test_si11), .SE(n9135), .CLK(n9322), 
        .Q(g185), .QN(n4384) );
  SDFFX1 DFF_161_Q_reg ( .D(g2950), .SI(g185), .SE(n9135), .CLK(n9322), .Q(
        g6231), .QN(n4318) );
  SDFFX1 DFF_162_Q_reg ( .D(g6231), .SI(g6231), .SE(n9135), .CLK(n9322), .Q(
        g6313), .QN(n4512) );
  SDFFX1 DFF_163_Q_reg ( .D(g6313), .SI(g6313), .SE(n9136), .CLK(n9323), .Q(
        g165), .QN(n4369) );
  SDFFX1 DFF_164_Q_reg ( .D(g22100), .SI(g165), .SE(n9144), .CLK(n9331), .Q(
        g130) );
  SDFFX1 DFF_165_Q_reg ( .D(g22122), .SI(g130), .SE(n9144), .CLK(n9331), .Q(
        g131) );
  SDFFX1 DFF_166_Q_reg ( .D(g22141), .SI(g131), .SE(n9144), .CLK(n9331), .Q(
        g129) );
  SDFFX1 DFF_167_Q_reg ( .D(g22123), .SI(g129), .SE(n9133), .CLK(n9320), .Q(
        g133) );
  SDFFX1 DFF_168_Q_reg ( .D(g22142), .SI(g133), .SE(n9145), .CLK(n9332), .Q(
        g134) );
  SDFFX1 DFF_169_Q_reg ( .D(g22161), .SI(g134), .SE(n9145), .CLK(n9332), .Q(
        g132) );
  SDFFX1 DFF_170_Q_reg ( .D(g22025), .SI(g132), .SE(n9145), .CLK(n9332), .Q(
        g142) );
  SDFFX1 DFF_171_Q_reg ( .D(g22027), .SI(g142), .SE(n9145), .CLK(n9332), .Q(
        g143) );
  SDFFX1 DFF_172_Q_reg ( .D(g22030), .SI(g143), .SE(n9145), .CLK(n9332), .Q(
        g141) );
  SDFFX1 DFF_173_Q_reg ( .D(g22028), .SI(g141), .SE(n9145), .CLK(n9332), .Q(
        g145) );
  SDFFX1 DFF_174_Q_reg ( .D(g22031), .SI(g145), .SE(n9145), .CLK(n9332), .Q(
        g146) );
  SDFFX1 DFF_175_Q_reg ( .D(g22037), .SI(g146), .SE(n9145), .CLK(n9332), .Q(
        test_so11) );
  SDFFX1 DFF_176_Q_reg ( .D(g22032), .SI(test_si12), .SE(n9145), .CLK(n9332), 
        .Q(g148) );
  SDFFX1 DFF_177_Q_reg ( .D(g22038), .SI(g148), .SE(n9145), .CLK(n9332), .Q(
        g149) );
  SDFFX1 DFF_178_Q_reg ( .D(g22047), .SI(g149), .SE(n9145), .CLK(n9332), .Q(
        g147) );
  SDFFX1 DFF_179_Q_reg ( .D(g22039), .SI(g147), .SE(n9147), .CLK(n9334), .Q(
        g151) );
  SDFFX1 DFF_180_Q_reg ( .D(g22048), .SI(g151), .SE(n9147), .CLK(n9334), .Q(
        g152) );
  SDFFX1 DFF_181_Q_reg ( .D(g22063), .SI(g152), .SE(n9147), .CLK(n9334), .Q(
        g150) );
  SDFFX1 DFF_182_Q_reg ( .D(g22049), .SI(g150), .SE(n9147), .CLK(n9334), .Q(
        g154) );
  SDFFX1 DFF_183_Q_reg ( .D(g22064), .SI(g154), .SE(n9147), .CLK(n9334), .Q(
        g155) );
  SDFFX1 DFF_184_Q_reg ( .D(g22079), .SI(g155), .SE(n9147), .CLK(n9334), .Q(
        g153) );
  SDFFX1 DFF_185_Q_reg ( .D(g22065), .SI(g153), .SE(n9149), .CLK(n9336), .Q(
        g157) );
  SDFFX1 DFF_186_Q_reg ( .D(g22080), .SI(g157), .SE(n9149), .CLK(n9336), .Q(
        g158) );
  SDFFX1 DFF_187_Q_reg ( .D(g22101), .SI(g158), .SE(n9149), .CLK(n9336), .Q(
        g156) );
  SDFFX1 DFF_188_Q_reg ( .D(g22081), .SI(g156), .SE(n9149), .CLK(n9336), .Q(
        g160) );
  SDFFX1 DFF_189_Q_reg ( .D(g22102), .SI(g160), .SE(n9149), .CLK(n9336), .Q(
        g161) );
  SDFFX1 DFF_190_Q_reg ( .D(g22124), .SI(g161), .SE(n9149), .CLK(n9336), .Q(
        g159) );
  SDFFX1 DFF_191_Q_reg ( .D(g22103), .SI(g159), .SE(n9149), .CLK(n9336), .Q(
        test_so12) );
  SDFFX1 DFF_192_Q_reg ( .D(g22125), .SI(test_si13), .SE(n9148), .CLK(n9335), 
        .Q(g164) );
  SDFFX1 DFF_193_Q_reg ( .D(g22143), .SI(g164), .SE(n9148), .CLK(n9335), .Q(
        g162) );
  SDFFX1 DFF_194_Q_reg ( .D(g25204), .SI(g162), .SE(n9148), .CLK(n9335), .Q(
        g169), .QN(n8730) );
  SDFFX1 DFF_195_Q_reg ( .D(g25206), .SI(g169), .SE(n9149), .CLK(n9336), .Q(
        g170), .QN(n8729) );
  SDFFX1 DFF_196_Q_reg ( .D(g25211), .SI(g170), .SE(n9147), .CLK(n9334), .Q(
        g168), .QN(n8728) );
  SDFFX1 DFF_197_Q_reg ( .D(g25207), .SI(g168), .SE(n9148), .CLK(n9335), .Q(
        g172), .QN(n8727) );
  SDFFX1 DFF_198_Q_reg ( .D(g25212), .SI(g172), .SE(n9148), .CLK(n9335), .Q(
        g173), .QN(n8726) );
  SDFFX1 DFF_199_Q_reg ( .D(g25218), .SI(g173), .SE(n9148), .CLK(n9335), .Q(
        g171), .QN(n8725) );
  SDFFX1 DFF_200_Q_reg ( .D(g25213), .SI(g171), .SE(n9148), .CLK(n9335), .Q(
        g175), .QN(n8724) );
  SDFFX1 DFF_201_Q_reg ( .D(g25219), .SI(g175), .SE(n9148), .CLK(n9335), .Q(
        g176), .QN(n8723) );
  SDFFX1 DFF_202_Q_reg ( .D(g25228), .SI(g176), .SE(n9148), .CLK(n9335), .Q(
        g174), .QN(n8722) );
  SDFFX1 DFF_203_Q_reg ( .D(g25220), .SI(g174), .SE(n9148), .CLK(n9335), .Q(
        g178), .QN(n8721) );
  SDFFX1 DFF_204_Q_reg ( .D(g25229), .SI(g178), .SE(n9148), .CLK(n9335), .Q(
        g179), .QN(n8720) );
  SDFFX1 DFF_205_Q_reg ( .D(g25239), .SI(g179), .SE(n9148), .CLK(n9335), .Q(
        g177), .QN(n8719) );
  SDFFX1 DFF_206_Q_reg ( .D(g30261), .SI(g177), .SE(n9159), .CLK(n9346), .Q(
        g186) );
  SDFFX1 DFF_207_Q_reg ( .D(g30267), .SI(g186), .SE(n9159), .CLK(n9346), .Q(
        test_so13) );
  SDFFX1 DFF_208_Q_reg ( .D(g30275), .SI(test_si14), .SE(n9159), .CLK(n9346), 
        .Q(g192) );
  SDFFX1 DFF_209_Q_reg ( .D(g30637), .SI(g192), .SE(n9159), .CLK(n9346), .Q(
        g231) );
  SDFFX1 DFF_210_Q_reg ( .D(g30640), .SI(g231), .SE(n9159), .CLK(n9346), .Q(
        g234) );
  SDFFX1 DFF_211_Q_reg ( .D(g30645), .SI(g234), .SE(n9159), .CLK(n9346), .Q(
        g237) );
  SDFFX1 DFF_212_Q_reg ( .D(g30668), .SI(g237), .SE(n9159), .CLK(n9346), .Q(
        g195) );
  SDFFX1 DFF_213_Q_reg ( .D(g30674), .SI(g195), .SE(n9159), .CLK(n9346), .Q(
        g198) );
  SDFFX1 DFF_214_Q_reg ( .D(g30680), .SI(g198), .SE(n9134), .CLK(n9321), .Q(
        g201) );
  SDFFX1 DFF_215_Q_reg ( .D(g30641), .SI(g201), .SE(n9160), .CLK(n9347), .Q(
        g240) );
  SDFFX1 DFF_216_Q_reg ( .D(g30646), .SI(g240), .SE(n9160), .CLK(n9347), .Q(
        g243) );
  SDFFX1 DFF_217_Q_reg ( .D(g30653), .SI(g243), .SE(n9161), .CLK(n9348), .Q(
        g246) );
  SDFFX1 DFF_218_Q_reg ( .D(g30276), .SI(g246), .SE(n9161), .CLK(n9348), .Q(
        g204) );
  SDFFX1 DFF_219_Q_reg ( .D(g30284), .SI(g204), .SE(n9161), .CLK(n9348), .Q(
        g207) );
  SDFFX1 DFF_220_Q_reg ( .D(g30292), .SI(g207), .SE(n9161), .CLK(n9348), .Q(
        g210) );
  SDFFX1 DFF_221_Q_reg ( .D(g30254), .SI(g210), .SE(n9161), .CLK(n9348), .Q(
        g249) );
  SDFFX1 DFF_222_Q_reg ( .D(g30257), .SI(g249), .SE(n9161), .CLK(n9348), .Q(
        g252) );
  SDFFX1 DFF_223_Q_reg ( .D(g30262), .SI(g252), .SE(n9161), .CLK(n9348), .Q(
        test_so14) );
  SDFFX1 DFF_224_Q_reg ( .D(g30245), .SI(test_si15), .SE(n9161), .CLK(n9348), 
        .Q(g213) );
  SDFFX1 DFF_225_Q_reg ( .D(g30246), .SI(g213), .SE(n9161), .CLK(n9348), .Q(
        g216) );
  SDFFX1 DFF_226_Q_reg ( .D(g30248), .SI(g216), .SE(n9161), .CLK(n9348), .Q(
        g219) );
  SDFFX1 DFF_227_Q_reg ( .D(g30258), .SI(g219), .SE(n9161), .CLK(n9348), .Q(
        g258) );
  SDFFX1 DFF_228_Q_reg ( .D(g30263), .SI(g258), .SE(n9161), .CLK(n9348), .Q(
        g261) );
  SDFFX1 DFF_229_Q_reg ( .D(g30268), .SI(g261), .SE(n9162), .CLK(n9349), .Q(
        g264) );
  SDFFX1 DFF_230_Q_reg ( .D(g30635), .SI(g264), .SE(n9162), .CLK(n9349), .Q(
        g222) );
  SDFFX1 DFF_231_Q_reg ( .D(g30636), .SI(g222), .SE(n9162), .CLK(n9349), .Q(
        g225) );
  SDFFX1 DFF_232_Q_reg ( .D(g30639), .SI(g225), .SE(n9162), .CLK(n9349), .Q(
        g228) );
  SDFFX1 DFF_233_Q_reg ( .D(g30661), .SI(g228), .SE(n9162), .CLK(n9349), .Q(
        g267) );
  SDFFX1 DFF_234_Q_reg ( .D(g30669), .SI(g267), .SE(n9162), .CLK(n9349), .Q(
        g270) );
  SDFFX1 DFF_235_Q_reg ( .D(g30675), .SI(g270), .SE(n9159), .CLK(n9346), .Q(
        g273) );
  SDFFX1 DFF_236_Q_reg ( .D(g25027), .SI(g273), .SE(n9160), .CLK(n9347), .Q(
        g92), .QN(n8821) );
  SDFFX1 DFF_237_Q_reg ( .D(g25932), .SI(g92), .SE(n9160), .CLK(n9347), .Q(g88), .QN(n9113) );
  SDFFX1 DFF_238_Q_reg ( .D(g26529), .SI(g88), .SE(n9160), .CLK(n9347), .Q(g83), .QN(n8820) );
  SDFFX1 DFF_239_Q_reg ( .D(g27120), .SI(g83), .SE(n9160), .CLK(n9347), .Q(
        test_so15) );
  SDFFX1 DFF_240_Q_reg ( .D(g27594), .SI(test_si16), .SE(n9160), .CLK(n9347), 
        .Q(g74), .QN(n8819) );
  SDFFX1 DFF_241_Q_reg ( .D(g28145), .SI(g74), .SE(n9160), .CLK(n9347), .Q(g70), .QN(n9096) );
  SDFFX1 DFF_242_Q_reg ( .D(g28634), .SI(g70), .SE(n9160), .CLK(n9347), .Q(g65), .QN(n8818) );
  SDFFX1 DFF_243_Q_reg ( .D(g29109), .SI(g65), .SE(n9160), .CLK(n9347), .Q(g61), .QN(n9105) );
  SDFFX1 DFF_244_Q_reg ( .D(g29353), .SI(g61), .SE(n9160), .CLK(n9347), .Q(g56), .QN(n8440) );
  SDFFX1 DFF_245_Q_reg ( .D(g29579), .SI(g56), .SE(n9160), .CLK(n9347), .Q(g52), .QN(n8286) );
  SDFFX1 DFF_246_Q_reg ( .D(g13110), .SI(g52), .SE(n9133), .CLK(n9320), .Q(
        g180) );
  SDFFX1 DFF_247_Q_reg ( .D(g180), .SI(g180), .SE(n9133), .CLK(n9320), .Q(
        g5549) );
  SDFFX1 DFF_248_Q_reg ( .D(g5549), .SI(g5549), .SE(n9133), .CLK(n9320), .Q(
        g181), .QN(n9088) );
  SDFFX1 DFF_251_Q_reg ( .D(g6447), .SI(g6447), .SE(n9133), .CLK(n9320), .Q(
        n4640), .QN(n4506) );
  SDFFX1 DFF_252_Q_reg ( .D(g5549), .SI(n4640), .SE(n9133), .CLK(n9320), .Q(
        g309), .QN(n4388) );
  SDFFX1 DFF_253_Q_reg ( .D(g27253), .SI(g309), .SE(n9165), .CLK(n9352), .Q(
        g354), .QN(n8772) );
  SDFFX1 DFF_254_Q_reg ( .D(g27255), .SI(g354), .SE(n9165), .CLK(n9352), .Q(
        g343), .QN(n8771) );
  SDFFX1 DFF_255_Q_reg ( .D(g27258), .SI(g343), .SE(n9165), .CLK(n9352), .Q(
        test_so16) );
  SDFFX1 DFF_256_Q_reg ( .D(g27256), .SI(test_si17), .SE(n9164), .CLK(n9351), 
        .Q(g369), .QN(n8750) );
  SDFFX1 DFF_257_Q_reg ( .D(g27259), .SI(g369), .SE(n9164), .CLK(n9351), .Q(
        g358), .QN(n8749) );
  SDFFX1 DFF_258_Q_reg ( .D(g27265), .SI(g358), .SE(n9164), .CLK(n9351), .Q(
        g361), .QN(n8748) );
  SDFFX1 DFF_259_Q_reg ( .D(g27260), .SI(g361), .SE(n9165), .CLK(n9352), .Q(
        g384), .QN(n8494) );
  SDFFX1 DFF_260_Q_reg ( .D(g27266), .SI(g384), .SE(n9165), .CLK(n9352), .Q(
        g373), .QN(n8496) );
  SDFFX1 DFF_261_Q_reg ( .D(g27277), .SI(g373), .SE(n9164), .CLK(n9351), .Q(
        g376), .QN(n8495) );
  SDFFX1 DFF_262_Q_reg ( .D(g27267), .SI(g376), .SE(n9166), .CLK(n9353), .Q(
        g398), .QN(n8761) );
  SDFFX1 DFF_263_Q_reg ( .D(g27278), .SI(g398), .SE(n9167), .CLK(n9354), .Q(
        g388), .QN(n8760) );
  SDFFX1 DFF_264_Q_reg ( .D(g27293), .SI(g388), .SE(n9158), .CLK(n9345), .Q(
        g391), .QN(n8759) );
  SDFFX1 DFF_265_Q_reg ( .D(g28732), .SI(g391), .SE(n9158), .CLK(n9345), .Q(
        g408) );
  SDFFX1 DFF_266_Q_reg ( .D(g28735), .SI(g408), .SE(n9164), .CLK(n9351), .Q(
        g411) );
  SDFFX1 DFF_267_Q_reg ( .D(g28744), .SI(g411), .SE(n9164), .CLK(n9351), .Q(
        g414) );
  SDFFX1 DFF_268_Q_reg ( .D(g29194), .SI(g414), .SE(n9164), .CLK(n9351), .Q(
        g417) );
  SDFFX1 DFF_269_Q_reg ( .D(g29197), .SI(g417), .SE(n9164), .CLK(n9351), .Q(
        g420) );
  SDFFX1 DFF_270_Q_reg ( .D(g29201), .SI(g420), .SE(n9158), .CLK(n9345), .Q(
        g423) );
  SDFFX1 DFF_271_Q_reg ( .D(g28736), .SI(g423), .SE(n9158), .CLK(n9345), .Q(
        test_so17) );
  SDFFX1 DFF_272_Q_reg ( .D(g28745), .SI(test_si18), .SE(n9158), .CLK(n9345), 
        .Q(g428), .QN(n8804) );
  SDFFX1 DFF_273_Q_reg ( .D(g28754), .SI(g428), .SE(n9158), .CLK(n9345), .Q(
        g426), .QN(n8803) );
  SDFFX1 DFF_274_Q_reg ( .D(g26803), .SI(g426), .SE(n9158), .CLK(n9345), .Q(
        g429) );
  SDFFX1 DFF_275_Q_reg ( .D(g26804), .SI(g429), .SE(n9158), .CLK(n9345), .Q(
        g432) );
  SDFFX1 DFF_276_Q_reg ( .D(g26807), .SI(g432), .SE(n9159), .CLK(n9346), .Q(
        g435) );
  SDFFX1 DFF_277_Q_reg ( .D(g26805), .SI(g435), .SE(n9163), .CLK(n9350), .Q(
        g438) );
  SDFFX1 DFF_278_Q_reg ( .D(g26808), .SI(g438), .SE(n9163), .CLK(n9350), .Q(
        g441) );
  SDFFX1 DFF_279_Q_reg ( .D(g26812), .SI(g441), .SE(n9164), .CLK(n9351), .Q(
        g444) );
  SDFFX1 DFF_280_Q_reg ( .D(g27759), .SI(g444), .SE(n9164), .CLK(n9351), .Q(
        g448), .QN(n8802) );
  SDFFX1 DFF_281_Q_reg ( .D(g27760), .SI(g448), .SE(n9164), .CLK(n9351), .Q(
        g449), .QN(n8801) );
  SDFFX1 DFF_282_Q_reg ( .D(g27762), .SI(g449), .SE(n9159), .CLK(n9346), .Q(
        g447), .QN(n8800) );
  SDFFX1 DFF_283_Q_reg ( .D(g29606), .SI(g447), .SE(n9159), .CLK(n9346), .Q(
        g312), .QN(n8407) );
  SDFFX1 DFF_284_Q_reg ( .D(g29608), .SI(g312), .SE(n9163), .CLK(n9350), .Q(
        g313), .QN(n8406) );
  SDFFX1 DFF_285_Q_reg ( .D(g29611), .SI(g313), .SE(n9163), .CLK(n9350), .Q(
        g314), .QN(n8405) );
  SDFFX1 DFF_286_Q_reg ( .D(g30699), .SI(g314), .SE(n9163), .CLK(n9350), .Q(
        g315), .QN(n8404) );
  SDFFX1 DFF_287_Q_reg ( .D(g30700), .SI(g315), .SE(n9163), .CLK(n9350), .Q(
        test_so18) );
  SDFFX1 DFF_288_Q_reg ( .D(g30702), .SI(test_si19), .SE(n9133), .CLK(n9320), 
        .Q(g317), .QN(n8403) );
  SDFFX1 DFF_289_Q_reg ( .D(g30455), .SI(g317), .SE(n9133), .CLK(n9320), .Q(
        g318), .QN(n8402) );
  SDFFX1 DFF_290_Q_reg ( .D(g30468), .SI(g318), .SE(n9134), .CLK(n9321), .Q(
        g319), .QN(n8401) );
  SDFFX1 DFF_291_Q_reg ( .D(g30482), .SI(g319), .SE(n9134), .CLK(n9321), .Q(
        g320), .QN(n8400) );
  SDFFX1 DFF_292_Q_reg ( .D(g29167), .SI(g320), .SE(n9162), .CLK(n9349), .Q(
        g322) );
  SDFFX1 DFF_293_Q_reg ( .D(g29169), .SI(g322), .SE(n9162), .CLK(n9349), .Q(
        g323) );
  SDFFX1 DFF_294_Q_reg ( .D(g29172), .SI(g323), .SE(n9162), .CLK(n9349), .Q(
        g321) );
  SDFFX1 DFF_295_Q_reg ( .D(g26655), .SI(g321), .SE(n9162), .CLK(n9349), .Q(
        g403), .QN(n8799) );
  SDFFX1 DFF_296_Q_reg ( .D(g26659), .SI(g403), .SE(n9162), .CLK(n9349), .Q(
        g404), .QN(n8798) );
  SDFFX1 DFF_297_Q_reg ( .D(g26664), .SI(g404), .SE(n9162), .CLK(n9349), .Q(
        g402), .QN(n8797) );
  SDFFX1 DFF_298_Q_reg ( .D(n4290), .SI(g402), .SE(n9163), .CLK(n9350), .Q(
        g450) );
  SDFFX1 DFF_299_Q_reg ( .D(g450), .SI(g450), .SE(n9163), .CLK(n9350), .Q(
        n8066), .QN(DFF_299_n1) );
  SDFFX1 DFF_300_Q_reg ( .D(n4569), .SI(n8066), .SE(n9163), .CLK(n9350), .Q(
        g452) );
  SDFFX1 DFF_301_Q_reg ( .D(g452), .SI(g452), .SE(n9163), .CLK(n9350), .Q(
        n8065), .QN(DFF_301_n1) );
  SDFFX1 DFF_302_Q_reg ( .D(n4561), .SI(n8065), .SE(n9163), .CLK(n9350), .Q(
        g454) );
  SDFFX1 DFF_303_Q_reg ( .D(g454), .SI(g454), .SE(n9163), .CLK(n9350), .Q(
        test_so19), .QN(DFF_303_n1) );
  SDFFX1 DFF_304_Q_reg ( .D(n4328), .SI(test_si20), .SE(n9145), .CLK(n9332), 
        .Q(g280) );
  SDFFX1 DFF_305_Q_reg ( .D(g280), .SI(g280), .SE(n9146), .CLK(n9333), .Q(
        n8062), .QN(DFF_305_n1) );
  SDFFX1 DFF_306_Q_reg ( .D(n4392), .SI(n8062), .SE(n9146), .CLK(n9333), .Q(
        g282) );
  SDFFX1 DFF_307_Q_reg ( .D(g282), .SI(g282), .SE(n9146), .CLK(n9333), .Q(
        n8061), .QN(DFF_307_n1) );
  SDFFX1 DFF_308_Q_reg ( .D(n4322), .SI(n8061), .SE(n9146), .CLK(n9333), .Q(
        g284) );
  SDFFX1 DFF_309_Q_reg ( .D(g284), .SI(g284), .SE(n9146), .CLK(n9333), .Q(
        n8060), .QN(DFF_309_n1) );
  SDFFX1 DFF_310_Q_reg ( .D(n4376), .SI(n8060), .SE(n9146), .CLK(n9333), .Q(
        g286) );
  SDFFX1 DFF_311_Q_reg ( .D(g286), .SI(g286), .SE(n9146), .CLK(n9333), .Q(
        n8059), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(n4380), .SI(n8059), .SE(n9146), .CLK(n9333), .Q(
        g288) );
  SDFFX1 DFF_313_Q_reg ( .D(g288), .SI(g288), .SE(n9146), .CLK(n9333), .Q(
        n8058), .QN(DFF_313_n1) );
  SDFFX1 DFF_314_Q_reg ( .D(g2857), .SI(n8058), .SE(n9146), .CLK(n9333), .Q(
        g290) );
  SDFFX1 DFF_315_Q_reg ( .D(g290), .SI(g290), .SE(n9146), .CLK(n9333), .Q(
        n8057), .QN(n4485) );
  SDFFX1 DFF_316_Q_reg ( .D(n4282), .SI(n8057), .SE(n9164), .CLK(n9351), .Q(
        n8056), .QN(n16490) );
  SDFFX1 DFF_317_Q_reg ( .D(g21346), .SI(n8056), .SE(n9134), .CLK(n9321), .Q(
        g305), .QN(n8546) );
  SDFFX1 DFF_328_Q_reg ( .D(n4278), .SI(g305), .SE(n9134), .CLK(n9321), .Q(
        n8055), .QN(DFF_328_n1) );
  SDFFX1 DFF_329_Q_reg ( .D(g354), .SI(n8055), .SE(n9165), .CLK(n9352), .Q(
        test_so20) );
  SDFFX1 DFF_330_Q_reg ( .D(test_so20), .SI(test_si21), .SE(n9165), .CLK(n9352), .Q(g349) );
  SDFFX1 DFF_331_Q_reg ( .D(g343), .SI(g349), .SE(n9165), .CLK(n9352), .Q(g350) );
  SDFFX1 DFF_332_Q_reg ( .D(g350), .SI(g350), .SE(n9165), .CLK(n9352), .Q(g351) );
  SDFFX1 DFF_333_Q_reg ( .D(test_so16), .SI(g351), .SE(n9165), .CLK(n9352), 
        .Q(g352) );
  SDFFX1 DFF_334_Q_reg ( .D(g352), .SI(g352), .SE(n9165), .CLK(n9352), .Q(g353) );
  SDFFX1 DFF_335_Q_reg ( .D(g369), .SI(g353), .SE(n9165), .CLK(n9352), .Q(g357) );
  SDFFX1 DFF_336_Q_reg ( .D(g357), .SI(g357), .SE(n9166), .CLK(n9353), .Q(g364) );
  SDFFX1 DFF_337_Q_reg ( .D(g358), .SI(g364), .SE(n9166), .CLK(n9353), .Q(g365) );
  SDFFX1 DFF_338_Q_reg ( .D(g365), .SI(g365), .SE(n9166), .CLK(n9353), .Q(g366) );
  SDFFX1 DFF_339_Q_reg ( .D(g361), .SI(g366), .SE(n9166), .CLK(n9353), .Q(g367) );
  SDFFX1 DFF_340_Q_reg ( .D(g367), .SI(g367), .SE(n9166), .CLK(n9353), .Q(g368) );
  SDFFX1 DFF_341_Q_reg ( .D(g384), .SI(g368), .SE(n9166), .CLK(n9353), .Q(g372) );
  SDFFX1 DFF_342_Q_reg ( .D(g372), .SI(g372), .SE(n9166), .CLK(n9353), .Q(g379) );
  SDFFX1 DFF_343_Q_reg ( .D(g373), .SI(g379), .SE(n9166), .CLK(n9353), .Q(g380) );
  SDFFX1 DFF_344_Q_reg ( .D(g380), .SI(g380), .SE(n9166), .CLK(n9353), .Q(g381) );
  SDFFX1 DFF_345_Q_reg ( .D(g376), .SI(g381), .SE(n9166), .CLK(n9353), .Q(
        test_so21) );
  SDFFX1 DFF_346_Q_reg ( .D(test_so21), .SI(test_si22), .SE(n9166), .CLK(n9353), .Q(g383) );
  SDFFX1 DFF_347_Q_reg ( .D(g398), .SI(g383), .SE(n9167), .CLK(n9354), .Q(g387) );
  SDFFX1 DFF_348_Q_reg ( .D(g387), .SI(g387), .SE(n9167), .CLK(n9354), .Q(g394) );
  SDFFX1 DFF_349_Q_reg ( .D(g388), .SI(g394), .SE(n9167), .CLK(n9354), .Q(g395) );
  SDFFX1 DFF_350_Q_reg ( .D(g395), .SI(g395), .SE(n9167), .CLK(n9354), .Q(g396) );
  SDFFX1 DFF_351_Q_reg ( .D(g391), .SI(g396), .SE(n9167), .CLK(n9354), .Q(g397) );
  SDFFX1 DFF_352_Q_reg ( .D(g397), .SI(g397), .SE(n9167), .CLK(n9354), .Q(g324) );
  SDFFX1 DFF_353_Q_reg ( .D(n4598), .SI(g324), .SE(n9167), .CLK(n9354), .Q(
        g5629) );
  SDFFX1 DFF_354_Q_reg ( .D(g5629), .SI(g5629), .SE(n9167), .CLK(n9354), .Q(
        g5648) );
  SDFFX1 DFF_355_Q_reg ( .D(g5648), .SI(g5648), .SE(n9167), .CLK(n9354), .Q(
        g337) );
  SDFFX1 DFF_356_Q_reg ( .D(n4598), .SI(g337), .SE(n9167), .CLK(n9354), .Q(
        g6485), .QN(n4298) );
  SDFFX1 DFF_357_Q_reg ( .D(g6485), .SI(g6485), .SE(n9167), .CLK(n9354), .Q(
        g6642), .QN(n4372) );
  SDFFX1 DFF_358_Q_reg ( .D(g6642), .SI(g6642), .SE(n9168), .CLK(n9355), .Q(
        g550), .QN(n4313) );
  SDFFX1 DFF_359_Q_reg ( .D(g21842), .SI(g550), .SE(n9168), .CLK(n9355), .Q(
        g554), .QN(n9053) );
  SDFFX1 DFF_360_Q_reg ( .D(g18678), .SI(g554), .SE(n9168), .CLK(n9355), .Q(
        g557), .QN(n4360) );
  SDFFX1 DFF_361_Q_reg ( .D(g18726), .SI(g557), .SE(n9168), .CLK(n9355), .Q(
        test_so22), .QN(n9126) );
  SDFFX1 DFF_362_Q_reg ( .D(n519), .SI(test_si23), .SE(n9172), .CLK(n9359), 
        .Q(g513) );
  SDFFX1 DFF_363_Q_reg ( .D(g513), .SI(g513), .SE(n9172), .CLK(n9359), .Q(g523) );
  SDFFX1 DFF_364_Q_reg ( .D(g523), .SI(g523), .SE(n9172), .CLK(n9359), .Q(g524) );
  SDFFX1 DFF_365_Q_reg ( .D(g455), .SI(g524), .SE(n9172), .CLK(n9359), .Q(g564) );
  SDFFX1 DFF_366_Q_reg ( .D(g564), .SI(g564), .SE(n9172), .CLK(n9359), .Q(g569) );
  SDFFX1 DFF_367_Q_reg ( .D(g458), .SI(g569), .SE(n9172), .CLK(n9359), .Q(g570) );
  SDFFX1 DFF_368_Q_reg ( .D(g570), .SI(g570), .SE(n9172), .CLK(n9359), .Q(g571) );
  SDFFX1 DFF_369_Q_reg ( .D(g461), .SI(g571), .SE(n9172), .CLK(n9359), .Q(g572) );
  SDFFX1 DFF_370_Q_reg ( .D(g572), .SI(g572), .SE(n9172), .CLK(n9359), .Q(g573) );
  SDFFX1 DFF_371_Q_reg ( .D(g465), .SI(g573), .SE(n9172), .CLK(n9359), .Q(g574) );
  SDFFX1 DFF_372_Q_reg ( .D(g574), .SI(g574), .SE(n9172), .CLK(n9359), .Q(g565) );
  SDFFX1 DFF_373_Q_reg ( .D(test_so24), .SI(g565), .SE(n9172), .CLK(n9359), 
        .Q(g566) );
  SDFFX1 DFF_374_Q_reg ( .D(g566), .SI(g566), .SE(n9173), .CLK(n9360), .Q(g567) );
  SDFFX1 DFF_375_Q_reg ( .D(g471), .SI(g567), .SE(n9173), .CLK(n9360), .Q(g568) );
  SDFFX1 DFF_376_Q_reg ( .D(g568), .SI(g568), .SE(n9173), .CLK(n9360), .Q(g489) );
  SDFFX1 DFF_377_Q_reg ( .D(g2950), .SI(g489), .SE(n9173), .CLK(n9360), .Q(
        test_so23), .QN(n9120) );
  SDFFX1 DFF_378_Q_reg ( .D(test_so23), .SI(test_si24), .SE(n9173), .CLK(n9360), .Q(g7956), .QN(n4461) );
  SDFFX1 DFF_379_Q_reg ( .D(g7956), .SI(g7956), .SE(n9173), .CLK(n9360), .Q(
        g485), .QN(n4466) );
  SDFFX1 DFF_380_Q_reg ( .D(g23067), .SI(g485), .SE(n9173), .CLK(n9360), .Q(
        g486) );
  SDFFX1 DFF_381_Q_reg ( .D(g23093), .SI(g486), .SE(n9173), .CLK(n9360), .Q(
        g487) );
  SDFFX1 DFF_382_Q_reg ( .D(g23117), .SI(g487), .SE(n9173), .CLK(n9360), .Q(
        g488) );
  SDFFX1 DFF_383_Q_reg ( .D(g23385), .SI(g488), .SE(n9173), .CLK(n9360), .Q(
        g455) );
  SDFFX1 DFF_384_Q_reg ( .D(g23399), .SI(g455), .SE(n9173), .CLK(n9360), .Q(
        g458) );
  SDFFX1 DFF_385_Q_reg ( .D(g24174), .SI(g458), .SE(n9174), .CLK(n9361), .Q(
        g461) );
  SDFFX1 DFF_386_Q_reg ( .D(g24178), .SI(g461), .SE(n9174), .CLK(n9361), .Q(
        g477) );
  SDFFX1 DFF_387_Q_reg ( .D(g24207), .SI(g477), .SE(n9174), .CLK(n9361), .Q(
        g478) );
  SDFFX1 DFF_388_Q_reg ( .D(g24216), .SI(g478), .SE(n9174), .CLK(n9361), .Q(
        g479) );
  SDFFX1 DFF_389_Q_reg ( .D(g23092), .SI(g479), .SE(n9174), .CLK(n9361), .Q(
        g480) );
  SDFFX1 DFF_390_Q_reg ( .D(g23000), .SI(g480), .SE(n9174), .CLK(n9361), .Q(
        g484) );
  SDFFX1 DFF_391_Q_reg ( .D(g23022), .SI(g484), .SE(n9174), .CLK(n9361), .Q(
        g464) );
  SDFFX1 DFF_392_Q_reg ( .D(g24206), .SI(g464), .SE(n9174), .CLK(n9361), .Q(
        g465) );
  SDFFX1 DFF_393_Q_reg ( .D(g24215), .SI(g465), .SE(n9174), .CLK(n9361), .Q(
        test_so24) );
  SDFFX1 DFF_394_Q_reg ( .D(g24228), .SI(test_si25), .SE(n9173), .CLK(n9360), 
        .Q(g471) );
  SDFFX1 DFF_395_Q_reg ( .D(n492), .SI(g471), .SE(n9174), .CLK(n9361), .Q(g528) );
  SDFFX1 DFF_396_Q_reg ( .D(g528), .SI(g528), .SE(n9174), .CLK(n9361), .Q(g535) );
  SDFFX1 DFF_397_Q_reg ( .D(g535), .SI(g535), .SE(n9174), .CLK(n9361), .Q(g542) );
  SDFFX1 DFF_398_Q_reg ( .D(g13149), .SI(g542), .SE(n9175), .CLK(n9362), .Q(
        g543) );
  SDFFX1 DFF_399_Q_reg ( .D(g543), .SI(g543), .SE(n9175), .CLK(n9362), .Q(g544) );
  SDFFX1 DFF_400_Q_reg ( .D(g21851), .SI(g544), .SE(n9175), .CLK(n9362), .Q(
        g548) );
  SDFFX1 DFF_401_Q_reg ( .D(g13111), .SI(g548), .SE(n9175), .CLK(n9362), .Q(
        g549) );
  SDFFX1 DFF_402_Q_reg ( .D(g549), .SI(g549), .SE(n9175), .CLK(n9362), .Q(g499), .QN(n4541) );
  SDFFX1 DFF_403_Q_reg ( .D(g13160), .SI(g499), .SE(n9175), .CLK(n9362), .Q(
        g558) );
  SDFFX1 DFF_404_Q_reg ( .D(g558), .SI(g558), .SE(n9175), .CLK(n9362), .Q(g559) );
  SDFFX1 DFF_405_Q_reg ( .D(g27261), .SI(g559), .SE(n9176), .CLK(n9363), .Q(
        g576), .QN(n8450) );
  SDFFX1 DFF_406_Q_reg ( .D(g27268), .SI(g576), .SE(n9176), .CLK(n9363), .Q(
        g577), .QN(n8452) );
  SDFFX1 DFF_407_Q_reg ( .D(g27279), .SI(g577), .SE(n9176), .CLK(n9363), .Q(
        g575), .QN(n8451) );
  SDFFX1 DFF_408_Q_reg ( .D(g27269), .SI(g575), .SE(n9176), .CLK(n9363), .Q(
        g579), .QN(n8462) );
  SDFFX1 DFF_409_Q_reg ( .D(g27280), .SI(g579), .SE(n9176), .CLK(n9363), .Q(
        test_so25) );
  SDFFX1 DFF_410_Q_reg ( .D(g27294), .SI(test_si26), .SE(n9176), .CLK(n9363), 
        .Q(g578), .QN(n8463) );
  SDFFX1 DFF_411_Q_reg ( .D(g27281), .SI(g578), .SE(n9176), .CLK(n9363), .Q(
        g582), .QN(n8294) );
  SDFFX1 DFF_412_Q_reg ( .D(g27295), .SI(g582), .SE(n9176), .CLK(n9363), .Q(
        g583), .QN(n8296) );
  SDFFX1 DFF_413_Q_reg ( .D(g27311), .SI(g583), .SE(n9176), .CLK(n9363), .Q(
        g581), .QN(n8295) );
  SDFFX1 DFF_414_Q_reg ( .D(g27296), .SI(g581), .SE(n9175), .CLK(n9362), .Q(
        g585), .QN(n8472) );
  SDFFX1 DFF_415_Q_reg ( .D(g27312), .SI(g585), .SE(n9176), .CLK(n9363), .Q(
        g586), .QN(n8474) );
  SDFFX1 DFF_416_Q_reg ( .D(g27327), .SI(g586), .SE(n9176), .CLK(n9363), .Q(
        g584), .QN(n8473) );
  SDFFX1 DFF_417_Q_reg ( .D(g24491), .SI(g584), .SE(n9176), .CLK(n9363), .Q(
        g587) );
  SDFFX1 DFF_418_Q_reg ( .D(g24498), .SI(g587), .SE(n9177), .CLK(n9364), .Q(
        g590) );
  SDFFX1 DFF_419_Q_reg ( .D(g24507), .SI(g590), .SE(n9177), .CLK(n9364), .Q(
        g593) );
  SDFFX1 DFF_420_Q_reg ( .D(g24499), .SI(g593), .SE(n9177), .CLK(n9364), .Q(
        g596) );
  SDFFX1 DFF_421_Q_reg ( .D(g24508), .SI(g596), .SE(n9177), .CLK(n9364), .Q(
        g599) );
  SDFFX1 DFF_422_Q_reg ( .D(g24519), .SI(g599), .SE(n9177), .CLK(n9364), .Q(
        g602) );
  SDFFX1 DFF_423_Q_reg ( .D(g28345), .SI(g602), .SE(n9177), .CLK(n9364), .Q(
        g614) );
  SDFFX1 DFF_424_Q_reg ( .D(g28349), .SI(g614), .SE(n9177), .CLK(n9364), .Q(
        g617) );
  SDFFX1 DFF_425_Q_reg ( .D(g28353), .SI(g617), .SE(n9175), .CLK(n9362), .Q(
        test_so26) );
  SDFFX1 DFF_426_Q_reg ( .D(g28342), .SI(test_si27), .SE(n9177), .CLK(n9364), 
        .Q(g605) );
  SDFFX1 DFF_427_Q_reg ( .D(g28344), .SI(g605), .SE(n9177), .CLK(n9364), .Q(
        g608) );
  SDFFX1 DFF_428_Q_reg ( .D(g28348), .SI(g608), .SE(n9177), .CLK(n9364), .Q(
        g611) );
  SDFFX1 DFF_429_Q_reg ( .D(g26541), .SI(g611), .SE(n9177), .CLK(n9364), .Q(
        g490) );
  SDFFX1 DFF_430_Q_reg ( .D(g26545), .SI(g490), .SE(n9177), .CLK(n9364), .Q(
        g493) );
  SDFFX1 DFF_431_Q_reg ( .D(g26553), .SI(g493), .SE(n9178), .CLK(n9365), .Q(
        g496) );
  SDFFX1 DFF_432_Q_reg ( .D(g499), .SI(g496), .SE(n9178), .CLK(n9365), .Q(g506), .QN(n4570) );
  SDFFX1 DFF_433_Q_reg ( .D(g22578), .SI(g506), .SE(n9178), .CLK(n9365), .Q(
        n4571) );
  SDFFX1 DFF_442_Q_reg ( .D(n517), .SI(n4571), .SE(n9178), .CLK(n9365), .Q(
        g16297) );
  SDFFX1 DFF_443_Q_reg ( .D(g16297), .SI(g16297), .SE(n9178), .CLK(n9365), .Q(
        g525), .QN(n8828) );
  SDFFX1 DFF_444_Q_reg ( .D(DFF_299_n1), .SI(g525), .SE(n9178), .CLK(n9365), 
        .Q(n8047) );
  SDFFX1 DFF_445_Q_reg ( .D(DFF_301_n1), .SI(n8047), .SE(n9178), .CLK(n9365), 
        .Q(n8046) );
  SDFFX1 DFF_446_Q_reg ( .D(DFF_303_n1), .SI(n8046), .SE(n9179), .CLK(n9366), 
        .Q(n8045) );
  SDFFX1 DFF_447_Q_reg ( .D(DFF_305_n1), .SI(n8045), .SE(n9179), .CLK(n9366), 
        .Q(n8044) );
  SDFFX1 DFF_448_Q_reg ( .D(DFF_307_n1), .SI(n8044), .SE(n9179), .CLK(n9366), 
        .Q(n8043) );
  SDFFX1 DFF_449_Q_reg ( .D(DFF_309_n1), .SI(n8043), .SE(n9179), .CLK(n9366), 
        .Q(test_so27) );
  SDFFX1 DFF_450_Q_reg ( .D(DFF_311_n1), .SI(test_si28), .SE(n9147), .CLK(
        n9334), .Q(g536) );
  SDFFX1 DFF_451_Q_reg ( .D(DFF_313_n1), .SI(g536), .SE(n9147), .CLK(n9334), 
        .Q(g537) );
  SDFFX1 DFF_452_Q_reg ( .D(g24059), .SI(g537), .SE(n9134), .CLK(n9321), .Q(
        g538), .QN(n4492) );
  SDFFX1 DFF_453_Q_reg ( .D(n4485), .SI(g538), .SE(n9146), .CLK(n9333), .Q(
        n8040) );
  SDFFX1 DFF_455_Q_reg ( .D(g6677), .SI(g6677), .SE(n9147), .CLK(n9334), .Q(
        g6911), .QN(n4359) );
  SDFFX1 DFF_456_Q_reg ( .D(g6911), .SI(g6911), .SE(n9147), .CLK(n9334), .Q(
        g629), .QN(n4295) );
  SDFFX1 DFF_457_Q_reg ( .D(g16654), .SI(g629), .SE(n9168), .CLK(n9355), .Q(
        g630), .QN(n9082) );
  SDFFX1 DFF_458_Q_reg ( .D(g20314), .SI(g630), .SE(n9168), .CLK(n9355), .Q(
        g659) );
  SDFFX1 DFF_459_Q_reg ( .D(g20682), .SI(g659), .SE(n9168), .CLK(n9355), .Q(
        g640), .QN(n4404) );
  SDFFX1 DFF_460_Q_reg ( .D(g23136), .SI(g640), .SE(n9168), .CLK(n9355), .Q(
        g633), .QN(n4478) );
  SDFFX1 DFF_461_Q_reg ( .D(g23324), .SI(g633), .SE(n9168), .CLK(n9355), .Q(
        g653), .QN(n4422) );
  SDFFX1 DFF_462_Q_reg ( .D(g24426), .SI(g653), .SE(n9168), .CLK(n9355), .Q(
        g646), .QN(n4414) );
  SDFFX1 DFF_463_Q_reg ( .D(g25185), .SI(g646), .SE(n9169), .CLK(n9356), .Q(
        g660), .QN(n4403) );
  SDFFX1 DFF_464_Q_reg ( .D(g26660), .SI(g660), .SE(n9169), .CLK(n9356), .Q(
        g672), .QN(n4413) );
  SDFFX1 DFF_465_Q_reg ( .D(g26776), .SI(g672), .SE(n9169), .CLK(n9356), .Q(
        test_so28), .QN(n9123) );
  SDFFX1 DFF_466_Q_reg ( .D(g27672), .SI(test_si29), .SE(n9169), .CLK(n9356), 
        .Q(g679), .QN(n4477) );
  SDFFX1 DFF_467_Q_reg ( .D(g28199), .SI(g679), .SE(n9170), .CLK(n9357), .Q(
        g686), .QN(n4396) );
  SDFFX1 DFF_468_Q_reg ( .D(g28668), .SI(g686), .SE(n9170), .CLK(n9357), .Q(
        g692), .QN(n4418) );
  SDFFX1 DFF_469_Q_reg ( .D(g20875), .SI(g692), .SE(n9170), .CLK(n9357), .Q(
        g699), .QN(n8940) );
  SDFFX1 DFF_470_Q_reg ( .D(g20879), .SI(g699), .SE(n9170), .CLK(n9357), .Q(
        g700), .QN(n8939) );
  SDFFX1 DFF_471_Q_reg ( .D(g20891), .SI(g700), .SE(n9170), .CLK(n9357), .Q(
        g698), .QN(n8978) );
  SDFFX1 DFF_472_Q_reg ( .D(g20880), .SI(g698), .SE(n9170), .CLK(n9357), .Q(
        g702), .QN(n8938) );
  SDFFX1 DFF_473_Q_reg ( .D(g20892), .SI(g702), .SE(n9171), .CLK(n9358), .Q(
        g703), .QN(n8937) );
  SDFFX1 DFF_474_Q_reg ( .D(g20901), .SI(g703), .SE(n9171), .CLK(n9358), .Q(
        g701), .QN(n8977) );
  SDFFX1 DFF_475_Q_reg ( .D(g20893), .SI(g701), .SE(n9171), .CLK(n9358), .Q(
        g705), .QN(n8936) );
  SDFFX1 DFF_476_Q_reg ( .D(g20902), .SI(g705), .SE(n9171), .CLK(n9358), .Q(
        g706), .QN(n8935) );
  SDFFX1 DFF_477_Q_reg ( .D(g20921), .SI(g706), .SE(n9171), .CLK(n9358), .Q(
        g704), .QN(n8976) );
  SDFFX1 DFF_478_Q_reg ( .D(g20903), .SI(g704), .SE(n9171), .CLK(n9358), .Q(
        g708), .QN(n8934) );
  SDFFX1 DFF_479_Q_reg ( .D(g20922), .SI(g708), .SE(n9171), .CLK(n9358), .Q(
        g709), .QN(n8933) );
  SDFFX1 DFF_480_Q_reg ( .D(g20944), .SI(g709), .SE(n9171), .CLK(n9358), .Q(
        g707), .QN(n8975) );
  SDFFX1 DFF_481_Q_reg ( .D(g20923), .SI(g707), .SE(n9171), .CLK(n9358), .Q(
        test_so29) );
  SDFFX1 DFF_482_Q_reg ( .D(g20945), .SI(test_si30), .SE(n9169), .CLK(n9356), 
        .Q(g712), .QN(n8932) );
  SDFFX1 DFF_483_Q_reg ( .D(g20966), .SI(g712), .SE(n9169), .CLK(n9356), .Q(
        g710), .QN(n8974) );
  SDFFX1 DFF_484_Q_reg ( .D(g20946), .SI(g710), .SE(n9169), .CLK(n9356), .Q(
        g714), .QN(n8931) );
  SDFFX1 DFF_485_Q_reg ( .D(g20967), .SI(g714), .SE(n9169), .CLK(n9356), .Q(
        g715), .QN(n8930) );
  SDFFX1 DFF_486_Q_reg ( .D(g20989), .SI(g715), .SE(n9169), .CLK(n9356), .Q(
        g713), .QN(n8973) );
  SDFFX1 DFF_487_Q_reg ( .D(g20968), .SI(g713), .SE(n9169), .CLK(n9356), .Q(
        g717), .QN(n8929) );
  SDFFX1 DFF_488_Q_reg ( .D(g20990), .SI(g717), .SE(n9169), .CLK(n9356), .Q(
        g718), .QN(n8928) );
  SDFFX1 DFF_489_Q_reg ( .D(g21009), .SI(g718), .SE(n9169), .CLK(n9356), .Q(
        g716), .QN(n8972) );
  SDFFX1 DFF_490_Q_reg ( .D(g20991), .SI(g716), .SE(n9170), .CLK(n9357), .Q(
        g720), .QN(n8927) );
  SDFFX1 DFF_491_Q_reg ( .D(g21010), .SI(g720), .SE(n9170), .CLK(n9357), .Q(
        g721), .QN(n8926) );
  SDFFX1 DFF_492_Q_reg ( .D(g21031), .SI(g721), .SE(n9170), .CLK(n9357), .Q(
        g719), .QN(n8971) );
  SDFFX1 DFF_493_Q_reg ( .D(g21011), .SI(g719), .SE(n9170), .CLK(n9357), .Q(
        g723), .QN(n8925) );
  SDFFX1 DFF_494_Q_reg ( .D(g21032), .SI(g723), .SE(n9170), .CLK(n9357), .Q(
        g724), .QN(n8924) );
  SDFFX1 DFF_495_Q_reg ( .D(g21051), .SI(g724), .SE(n9170), .CLK(n9357), .Q(
        g722), .QN(n8970) );
  SDFFX1 DFF_496_Q_reg ( .D(g20876), .SI(g722), .SE(n9171), .CLK(n9358), .Q(
        g726), .QN(n8923) );
  SDFFX1 DFF_497_Q_reg ( .D(g20881), .SI(g726), .SE(n9171), .CLK(n9358), .Q(
        test_so30) );
  SDFFX1 DFF_498_Q_reg ( .D(g20894), .SI(test_si31), .SE(n9171), .CLK(n9358), 
        .Q(g725), .QN(n8969) );
  SDFFX1 DFF_499_Q_reg ( .D(g20924), .SI(g725), .SE(n9175), .CLK(n9362), .Q(
        g729), .QN(n8684) );
  SDFFX1 DFF_500_Q_reg ( .D(g20947), .SI(g729), .SE(n9175), .CLK(n9362), .Q(
        g730), .QN(n8676) );
  SDFFX1 DFF_501_Q_reg ( .D(g20969), .SI(g730), .SE(n9175), .CLK(n9362), .Q(
        g728), .QN(n8738) );
  SDFFX1 DFF_502_Q_reg ( .D(g20948), .SI(g728), .SE(n9178), .CLK(n9365), .Q(
        g732), .QN(n8683) );
  SDFFX1 DFF_503_Q_reg ( .D(g20970), .SI(g732), .SE(n9178), .CLK(n9365), .Q(
        g733), .QN(n8675) );
  SDFFX1 DFF_504_Q_reg ( .D(g20992), .SI(g733), .SE(n9178), .CLK(n9365), .Q(
        g731), .QN(n8737) );
  SDFFX1 DFF_505_Q_reg ( .D(g25260), .SI(g731), .SE(n9178), .CLK(n9365), .Q(
        g735) );
  SDFFX1 DFF_506_Q_reg ( .D(g25262), .SI(g735), .SE(n9178), .CLK(n9365), .Q(
        g736) );
  SDFFX1 DFF_507_Q_reg ( .D(g25266), .SI(g736), .SE(n9134), .CLK(n9321), .Q(
        g734) );
  SDFFX1 DFF_508_Q_reg ( .D(g22218), .SI(g734), .SE(n9168), .CLK(n9355), .Q(
        g738) );
  SDFFX1 DFF_509_Q_reg ( .D(g22231), .SI(g738), .SE(n9168), .CLK(n9355), .Q(
        g739) );
  SDFFX1 DFF_510_Q_reg ( .D(g22242), .SI(g739), .SE(n9179), .CLK(n9366), .Q(
        g737) );
  SDFFX1 DFF_511_Q_reg ( .D(g2950), .SI(g737), .SE(n9179), .CLK(n9366), .Q(
        g6368), .QN(n4323) );
  SDFFX1 DFF_512_Q_reg ( .D(g6368), .SI(g6368), .SE(n9179), .CLK(n9366), .Q(
        g6518), .QN(n4312) );
  SDFFX1 DFF_513_Q_reg ( .D(g6518), .SI(g6518), .SE(n9179), .CLK(n9366), .Q(
        test_so31), .QN(n9118) );
  SDFFX1 DFF_514_Q_reg ( .D(g22126), .SI(test_si32), .SE(n9180), .CLK(n9367), 
        .Q(g818), .QN(n9026) );
  SDFFX1 DFF_515_Q_reg ( .D(g22145), .SI(g818), .SE(n9184), .CLK(n9371), .Q(
        g819), .QN(n9025) );
  SDFFX1 DFF_516_Q_reg ( .D(g22162), .SI(g819), .SE(n9184), .CLK(n9371), .Q(
        g817), .QN(n8659) );
  SDFFX1 DFF_517_Q_reg ( .D(g22146), .SI(g817), .SE(n9184), .CLK(n9371), .Q(
        g821), .QN(n9024) );
  SDFFX1 DFF_518_Q_reg ( .D(g22163), .SI(g821), .SE(n9184), .CLK(n9371), .Q(
        g822), .QN(n9023) );
  SDFFX1 DFF_519_Q_reg ( .D(g22177), .SI(g822), .SE(n9184), .CLK(n9371), .Q(
        g820), .QN(n8658) );
  SDFFX1 DFF_520_Q_reg ( .D(g22029), .SI(g820), .SE(n9185), .CLK(n9372), .Q(
        g830), .QN(n9022) );
  SDFFX1 DFF_521_Q_reg ( .D(g22033), .SI(g830), .SE(n9185), .CLK(n9372), .Q(
        g831), .QN(n9021) );
  SDFFX1 DFF_522_Q_reg ( .D(g22040), .SI(g831), .SE(n9185), .CLK(n9372), .Q(
        g829), .QN(n8657) );
  SDFFX1 DFF_523_Q_reg ( .D(g22034), .SI(g829), .SE(n9185), .CLK(n9372), .Q(
        g833), .QN(n9020) );
  SDFFX1 DFF_524_Q_reg ( .D(g22041), .SI(g833), .SE(n9185), .CLK(n9372), .Q(
        g834), .QN(n9019) );
  SDFFX1 DFF_525_Q_reg ( .D(g22054), .SI(g834), .SE(n9185), .CLK(n9372), .Q(
        g832), .QN(n8656) );
  SDFFX1 DFF_526_Q_reg ( .D(g22042), .SI(g832), .SE(n9185), .CLK(n9372), .Q(
        g836), .QN(n9018) );
  SDFFX1 DFF_527_Q_reg ( .D(g22055), .SI(g836), .SE(n9185), .CLK(n9372), .Q(
        g837), .QN(n9017) );
  SDFFX1 DFF_528_Q_reg ( .D(g22066), .SI(g837), .SE(n9185), .CLK(n9372), .Q(
        g835), .QN(n8655) );
  SDFFX1 DFF_529_Q_reg ( .D(g22056), .SI(g835), .SE(n9185), .CLK(n9372), .Q(
        test_so32) );
  SDFFX1 DFF_530_Q_reg ( .D(g22067), .SI(test_si33), .SE(n9185), .CLK(n9372), 
        .Q(g840) );
  SDFFX1 DFF_531_Q_reg ( .D(g22087), .SI(g840), .SE(n9185), .CLK(n9372), .Q(
        g838) );
  SDFFX1 DFF_532_Q_reg ( .D(g22068), .SI(g838), .SE(n9186), .CLK(n9373), .Q(
        g842) );
  SDFFX1 DFF_533_Q_reg ( .D(g22088), .SI(g842), .SE(n9186), .CLK(n9373), .Q(
        g843) );
  SDFFX1 DFF_534_Q_reg ( .D(g22104), .SI(g843), .SE(n9186), .CLK(n9373), .Q(
        g841) );
  SDFFX1 DFF_535_Q_reg ( .D(g22089), .SI(g841), .SE(n9186), .CLK(n9373), .Q(
        g845), .QN(n9013) );
  SDFFX1 DFF_536_Q_reg ( .D(g22105), .SI(g845), .SE(n9186), .CLK(n9373), .Q(
        g846), .QN(n9012) );
  SDFFX1 DFF_537_Q_reg ( .D(g22127), .SI(g846), .SE(n9186), .CLK(n9373), .Q(
        g844), .QN(n8652) );
  SDFFX1 DFF_538_Q_reg ( .D(g22106), .SI(g844), .SE(n9186), .CLK(n9373), .Q(
        g848) );
  SDFFX1 DFF_539_Q_reg ( .D(g22128), .SI(g848), .SE(n9186), .CLK(n9373), .Q(
        g849) );
  SDFFX1 DFF_540_Q_reg ( .D(g22147), .SI(g849), .SE(n9186), .CLK(n9373), .Q(
        g847) );
  SDFFX1 DFF_541_Q_reg ( .D(g22129), .SI(g847), .SE(n9180), .CLK(n9367), .Q(
        g851) );
  SDFFX1 DFF_542_Q_reg ( .D(g22148), .SI(g851), .SE(n9186), .CLK(n9373), .Q(
        g852) );
  SDFFX1 DFF_543_Q_reg ( .D(g22164), .SI(g852), .SE(n9186), .CLK(n9373), .Q(
        g850) );
  SDFFX1 DFF_544_Q_reg ( .D(g25209), .SI(g850), .SE(n9186), .CLK(n9373), .Q(
        g857), .QN(n8718) );
  SDFFX1 DFF_545_Q_reg ( .D(g25214), .SI(g857), .SE(n9187), .CLK(n9374), .Q(
        test_so33) );
  SDFFX1 DFF_546_Q_reg ( .D(g25221), .SI(test_si34), .SE(n9179), .CLK(n9366), 
        .Q(g856), .QN(n8717) );
  SDFFX1 DFF_547_Q_reg ( .D(g25215), .SI(g856), .SE(n9179), .CLK(n9366), .Q(
        g860), .QN(n8716) );
  SDFFX1 DFF_548_Q_reg ( .D(g25222), .SI(g860), .SE(n9179), .CLK(n9366), .Q(
        g861), .QN(n8715) );
  SDFFX1 DFF_549_Q_reg ( .D(g25230), .SI(g861), .SE(n9179), .CLK(n9366), .Q(
        g859), .QN(n8714) );
  SDFFX1 DFF_550_Q_reg ( .D(g25223), .SI(g859), .SE(n9180), .CLK(n9367), .Q(
        g863), .QN(n8713) );
  SDFFX1 DFF_551_Q_reg ( .D(g25231), .SI(g863), .SE(n9180), .CLK(n9367), .Q(
        g864), .QN(n8712) );
  SDFFX1 DFF_552_Q_reg ( .D(g25240), .SI(g864), .SE(n9180), .CLK(n9367), .Q(
        g862), .QN(n8711) );
  SDFFX1 DFF_553_Q_reg ( .D(g25232), .SI(g862), .SE(n9180), .CLK(n9367), .Q(
        g866), .QN(n8710) );
  SDFFX1 DFF_554_Q_reg ( .D(g25241), .SI(g866), .SE(n9180), .CLK(n9367), .Q(
        g867) );
  SDFFX1 DFF_555_Q_reg ( .D(g25248), .SI(g867), .SE(n9180), .CLK(n9367), .Q(
        g865), .QN(n8708) );
  SDFFX1 DFF_556_Q_reg ( .D(g30269), .SI(g865), .SE(n9189), .CLK(n9376), .Q(
        g873) );
  SDFFX1 DFF_557_Q_reg ( .D(g30277), .SI(g873), .SE(n9190), .CLK(n9377), .Q(
        g876) );
  SDFFX1 DFF_558_Q_reg ( .D(g30285), .SI(g876), .SE(n9190), .CLK(n9377), .Q(
        g879) );
  SDFFX1 DFF_559_Q_reg ( .D(g30643), .SI(g879), .SE(n9190), .CLK(n9377), .Q(
        g918) );
  SDFFX1 DFF_560_Q_reg ( .D(g30648), .SI(g918), .SE(n9190), .CLK(n9377), .Q(
        g921) );
  SDFFX1 DFF_561_Q_reg ( .D(g30654), .SI(g921), .SE(n9190), .CLK(n9377), .Q(
        test_so34) );
  SDFFX1 DFF_562_Q_reg ( .D(g30676), .SI(test_si35), .SE(n9180), .CLK(n9367), 
        .Q(g882) );
  SDFFX1 DFF_563_Q_reg ( .D(g30681), .SI(g882), .SE(n9181), .CLK(n9368), .Q(
        g885) );
  SDFFX1 DFF_564_Q_reg ( .D(g30687), .SI(g885), .SE(n9181), .CLK(n9368), .Q(
        g888) );
  SDFFX1 DFF_565_Q_reg ( .D(g30649), .SI(g888), .SE(n9181), .CLK(n9368), .Q(
        g927) );
  SDFFX1 DFF_566_Q_reg ( .D(g30655), .SI(g927), .SE(n9181), .CLK(n9368), .Q(
        g930) );
  SDFFX1 DFF_567_Q_reg ( .D(g30662), .SI(g930), .SE(n9180), .CLK(n9367), .Q(
        g933) );
  SDFFX1 DFF_568_Q_reg ( .D(g30286), .SI(g933), .SE(n9181), .CLK(n9368), .Q(
        g891) );
  SDFFX1 DFF_569_Q_reg ( .D(g30293), .SI(g891), .SE(n9181), .CLK(n9368), .Q(
        g894) );
  SDFFX1 DFF_570_Q_reg ( .D(g30298), .SI(g894), .SE(n9181), .CLK(n9368), .Q(
        g897) );
  SDFFX1 DFF_571_Q_reg ( .D(g30259), .SI(g897), .SE(n9181), .CLK(n9368), .Q(
        g936) );
  SDFFX1 DFF_572_Q_reg ( .D(g30264), .SI(g936), .SE(n9181), .CLK(n9368), .Q(
        g939) );
  SDFFX1 DFF_573_Q_reg ( .D(g30270), .SI(g939), .SE(n9181), .CLK(n9368), .Q(
        g942) );
  SDFFX1 DFF_574_Q_reg ( .D(g30247), .SI(g942), .SE(n9181), .CLK(n9368), .Q(
        g900) );
  SDFFX1 DFF_575_Q_reg ( .D(g30249), .SI(g900), .SE(n9181), .CLK(n9368), .Q(
        g903) );
  SDFFX1 DFF_576_Q_reg ( .D(g30251), .SI(g903), .SE(n9182), .CLK(n9369), .Q(
        g906) );
  SDFFX1 DFF_577_Q_reg ( .D(g30265), .SI(g906), .SE(n9182), .CLK(n9369), .Q(
        test_so35) );
  SDFFX1 DFF_578_Q_reg ( .D(g30271), .SI(test_si36), .SE(n9182), .CLK(n9369), 
        .Q(g948) );
  SDFFX1 DFF_579_Q_reg ( .D(g30278), .SI(g948), .SE(n9182), .CLK(n9369), .Q(
        g951) );
  SDFFX1 DFF_580_Q_reg ( .D(g30638), .SI(g951), .SE(n9182), .CLK(n9369), .Q(
        g909) );
  SDFFX1 DFF_581_Q_reg ( .D(g30642), .SI(g909), .SE(n9182), .CLK(n9369), .Q(
        g912) );
  SDFFX1 DFF_582_Q_reg ( .D(g30647), .SI(g912), .SE(n9182), .CLK(n9369), .Q(
        g915) );
  SDFFX1 DFF_583_Q_reg ( .D(g30670), .SI(g915), .SE(n9182), .CLK(n9369), .Q(
        g954) );
  SDFFX1 DFF_584_Q_reg ( .D(g30677), .SI(g954), .SE(n9182), .CLK(n9369), .Q(
        g957) );
  SDFFX1 DFF_585_Q_reg ( .D(g30682), .SI(g957), .SE(n9182), .CLK(n9369), .Q(
        g960) );
  SDFFX1 DFF_586_Q_reg ( .D(g25042), .SI(g960), .SE(n9182), .CLK(n9369), .Q(
        g780), .QN(n8817) );
  SDFFX1 DFF_587_Q_reg ( .D(g25935), .SI(g780), .SE(n9182), .CLK(n9369), .Q(
        g776), .QN(n9101) );
  SDFFX1 DFF_588_Q_reg ( .D(g26530), .SI(g776), .SE(n9183), .CLK(n9370), .Q(
        g771), .QN(n8816) );
  SDFFX1 DFF_589_Q_reg ( .D(g27123), .SI(g771), .SE(n9183), .CLK(n9370), .Q(
        g767), .QN(n9100) );
  SDFFX1 DFF_590_Q_reg ( .D(g27603), .SI(g767), .SE(n9183), .CLK(n9370), .Q(
        g762), .QN(n8815) );
  SDFFX1 DFF_591_Q_reg ( .D(g28146), .SI(g762), .SE(n9183), .CLK(n9370), .Q(
        g758), .QN(n9099) );
  SDFFX1 DFF_592_Q_reg ( .D(g28635), .SI(g758), .SE(n9183), .CLK(n9370), .Q(
        g753), .QN(n8814) );
  SDFFX1 DFF_593_Q_reg ( .D(g29110), .SI(g753), .SE(n9183), .CLK(n9370), .Q(
        test_so36) );
  SDFFX1 DFF_594_Q_reg ( .D(g29354), .SI(test_si37), .SE(n9183), .CLK(n9370), 
        .Q(g744), .QN(n8439) );
  SDFFX1 DFF_595_Q_reg ( .D(g29580), .SI(g744), .SE(n9183), .CLK(n9370), .Q(
        g740), .QN(n8285) );
  SDFFX1 DFF_596_Q_reg ( .D(g13110), .SI(g740), .SE(n9183), .CLK(n9370), .Q(
        g868) );
  SDFFX1 DFF_597_Q_reg ( .D(g868), .SI(g868), .SE(n9183), .CLK(n9370), .Q(
        g5595) );
  SDFFX1 DFF_598_Q_reg ( .D(g5595), .SI(g5595), .SE(n9183), .CLK(n9370), .Q(
        g869), .QN(n9089) );
  SDFFX1 DFF_599_Q_reg ( .D(g2950), .SI(g869), .SE(n9183), .CLK(n9370), .Q(
        g5472), .QN(n4363) );
  SDFFX1 DFF_600_Q_reg ( .D(g5472), .SI(g5472), .SE(n9184), .CLK(n9371), .Q(
        g6712), .QN(n4364) );
  SDFFX1 DFF_601_Q_reg ( .D(g6712), .SI(g6712), .SE(n9184), .CLK(n9371), .Q(
        g1088), .QN(n4381) );
  SDFFX1 DFF_602_Q_reg ( .D(g5595), .SI(g1088), .SE(n9184), .CLK(n9371), .Q(
        g996), .QN(n4387) );
  SDFFX1 DFF_603_Q_reg ( .D(g27257), .SI(g996), .SE(n9189), .CLK(n9376), .Q(
        g1041), .QN(n8770) );
  SDFFX1 DFF_604_Q_reg ( .D(g27262), .SI(g1041), .SE(n9189), .CLK(n9376), .Q(
        g1030), .QN(n8769) );
  SDFFX1 DFF_605_Q_reg ( .D(g27270), .SI(g1030), .SE(n9189), .CLK(n9376), .Q(
        g1033), .QN(n8768) );
  SDFFX1 DFF_606_Q_reg ( .D(g27263), .SI(g1033), .SE(n9189), .CLK(n9376), .Q(
        g1056), .QN(n8747) );
  SDFFX1 DFF_607_Q_reg ( .D(g27271), .SI(g1056), .SE(n9189), .CLK(n9376), .Q(
        g1045), .QN(n8746) );
  SDFFX1 DFF_608_Q_reg ( .D(g27282), .SI(g1045), .SE(n9189), .CLK(n9376), .Q(
        g1048), .QN(n8745) );
  SDFFX1 DFF_609_Q_reg ( .D(g27272), .SI(g1048), .SE(n9189), .CLK(n9376), .Q(
        test_so37) );
  SDFFX1 DFF_610_Q_reg ( .D(g27283), .SI(test_si38), .SE(n9189), .CLK(n9376), 
        .Q(g1060), .QN(n8492) );
  SDFFX1 DFF_611_Q_reg ( .D(g27297), .SI(g1060), .SE(n9189), .CLK(n9376), .Q(
        g1063), .QN(n8493) );
  SDFFX1 DFF_612_Q_reg ( .D(g27284), .SI(g1063), .SE(n9189), .CLK(n9376), .Q(
        g1085), .QN(n8758) );
  SDFFX1 DFF_613_Q_reg ( .D(g27298), .SI(g1085), .SE(n9189), .CLK(n9376), .Q(
        g1075), .QN(n8757) );
  SDFFX1 DFF_614_Q_reg ( .D(g27313), .SI(g1075), .SE(n9187), .CLK(n9374), .Q(
        g1078), .QN(n8756) );
  SDFFX1 DFF_615_Q_reg ( .D(g28738), .SI(g1078), .SE(n9187), .CLK(n9374), .Q(
        g1095) );
  SDFFX1 DFF_616_Q_reg ( .D(g28746), .SI(g1095), .SE(n9188), .CLK(n9375), .Q(
        g1098) );
  SDFFX1 DFF_617_Q_reg ( .D(g28758), .SI(g1098), .SE(n9188), .CLK(n9375), .Q(
        g1101) );
  SDFFX1 DFF_618_Q_reg ( .D(g29198), .SI(g1101), .SE(n9188), .CLK(n9375), .Q(
        g1104) );
  SDFFX1 DFF_619_Q_reg ( .D(g29204), .SI(g1104), .SE(n9188), .CLK(n9375), .Q(
        g1107) );
  SDFFX1 DFF_620_Q_reg ( .D(g29209), .SI(g1107), .SE(n9187), .CLK(n9374), .Q(
        g1110) );
  SDFFX1 DFF_621_Q_reg ( .D(g28747), .SI(g1110), .SE(n9187), .CLK(n9374), .Q(
        g1114), .QN(n8796) );
  SDFFX1 DFF_622_Q_reg ( .D(g28759), .SI(g1114), .SE(n9187), .CLK(n9374), .Q(
        g1115), .QN(n8781) );
  SDFFX1 DFF_623_Q_reg ( .D(g28767), .SI(g1115), .SE(n9187), .CLK(n9374), .Q(
        g1113), .QN(n8795) );
  SDFFX1 DFF_624_Q_reg ( .D(g26806), .SI(g1113), .SE(n9187), .CLK(n9374), .Q(
        g1116) );
  SDFFX1 DFF_625_Q_reg ( .D(g26809), .SI(g1116), .SE(n9187), .CLK(n9374), .Q(
        test_so38) );
  SDFFX1 DFF_626_Q_reg ( .D(g26813), .SI(test_si39), .SE(n9187), .CLK(n9374), 
        .Q(g1122) );
  SDFFX1 DFF_627_Q_reg ( .D(g26810), .SI(g1122), .SE(n9188), .CLK(n9375), .Q(
        g1125) );
  SDFFX1 DFF_628_Q_reg ( .D(g26814), .SI(g1125), .SE(n9188), .CLK(n9375), .Q(
        g1128) );
  SDFFX1 DFF_629_Q_reg ( .D(g26818), .SI(g1128), .SE(n9188), .CLK(n9375), .Q(
        g1131) );
  SDFFX1 DFF_630_Q_reg ( .D(g27761), .SI(g1131), .SE(n9188), .CLK(n9375), .Q(
        g1135), .QN(n8794) );
  SDFFX1 DFF_631_Q_reg ( .D(g27763), .SI(g1135), .SE(n9188), .CLK(n9375), .Q(
        g1136), .QN(n8780) );
  SDFFX1 DFF_632_Q_reg ( .D(g27765), .SI(g1136), .SE(n9187), .CLK(n9374), .Q(
        g1134), .QN(n8793) );
  SDFFX1 DFF_633_Q_reg ( .D(g29609), .SI(g1134), .SE(n9188), .CLK(n9375), .Q(
        g999), .QN(n8399) );
  SDFFX1 DFF_634_Q_reg ( .D(g29612), .SI(g999), .SE(n9188), .CLK(n9375), .Q(
        g1000), .QN(n8382) );
  SDFFX1 DFF_635_Q_reg ( .D(g29616), .SI(g1000), .SE(n9187), .CLK(n9374), .Q(
        g1001), .QN(n8398) );
  SDFFX1 DFF_636_Q_reg ( .D(g30701), .SI(g1001), .SE(n9180), .CLK(n9367), .Q(
        g1002), .QN(n8397) );
  SDFFX1 DFF_637_Q_reg ( .D(g30703), .SI(g1002), .SE(n9184), .CLK(n9371), .Q(
        g1003), .QN(n8381) );
  SDFFX1 DFF_638_Q_reg ( .D(g30705), .SI(g1003), .SE(n9184), .CLK(n9371), .Q(
        g1004), .QN(n8396) );
  SDFFX1 DFF_639_Q_reg ( .D(g30470), .SI(g1004), .SE(n9180), .CLK(n9367), .Q(
        g1005), .QN(n8395) );
  SDFFX1 DFF_640_Q_reg ( .D(g30485), .SI(g1005), .SE(n9184), .CLK(n9371), .Q(
        g1006), .QN(n8380) );
  SDFFX1 DFF_641_Q_reg ( .D(g30500), .SI(g1006), .SE(n9184), .CLK(n9371), .Q(
        test_so39) );
  SDFFX1 DFF_642_Q_reg ( .D(g29170), .SI(test_si40), .SE(n9190), .CLK(n9377), 
        .Q(g1009) );
  SDFFX1 DFF_643_Q_reg ( .D(g29173), .SI(g1009), .SE(n9190), .CLK(n9377), .Q(
        g1010) );
  SDFFX1 DFF_644_Q_reg ( .D(g29179), .SI(g1010), .SE(n9190), .CLK(n9377), .Q(
        g1008) );
  SDFFX1 DFF_645_Q_reg ( .D(g26661), .SI(g1008), .SE(n9190), .CLK(n9377), .Q(
        g1090), .QN(n8792) );
  SDFFX1 DFF_646_Q_reg ( .D(g26665), .SI(g1090), .SE(n9190), .CLK(n9377), .Q(
        g1091), .QN(n8779) );
  SDFFX1 DFF_647_Q_reg ( .D(g26669), .SI(g1091), .SE(n9190), .CLK(n9377), .Q(
        g1089), .QN(n8791) );
  SDFFX1 DFF_648_Q_reg ( .D(n4289), .SI(g1089), .SE(n9190), .CLK(n9377), .Q(
        g1137) );
  SDFFX1 DFF_649_Q_reg ( .D(g1137), .SI(g1137), .SE(n9191), .CLK(n9378), .Q(
        n8027), .QN(DFF_649_n1) );
  SDFFX1 DFF_650_Q_reg ( .D(n4567), .SI(n8027), .SE(n9191), .CLK(n9378), .Q(
        g1139) );
  SDFFX1 DFF_651_Q_reg ( .D(g1139), .SI(g1139), .SE(n9191), .CLK(n9378), .Q(
        n8026), .QN(DFF_651_n1) );
  SDFFX1 DFF_652_Q_reg ( .D(n4559), .SI(n8026), .SE(n9191), .CLK(n9378), .Q(
        g1141) );
  SDFFX1 DFF_653_Q_reg ( .D(g1141), .SI(g1141), .SE(n9191), .CLK(n9378), .Q(
        n8025), .QN(DFF_653_n1) );
  SDFFX1 DFF_654_Q_reg ( .D(n4327), .SI(n8025), .SE(n9191), .CLK(n9378), .Q(
        g967) );
  SDFFX1 DFF_655_Q_reg ( .D(g967), .SI(g967), .SE(n9191), .CLK(n9378), .Q(
        n8024), .QN(DFF_655_n1) );
  SDFFX1 DFF_656_Q_reg ( .D(n4391), .SI(n8024), .SE(n9191), .CLK(n9378), .Q(
        g969) );
  SDFFX1 DFF_657_Q_reg ( .D(g969), .SI(g969), .SE(n9191), .CLK(n9378), .Q(
        test_so40), .QN(DFF_657_n1) );
  SDFFX1 DFF_658_Q_reg ( .D(n4321), .SI(test_si41), .SE(n9140), .CLK(n9327), 
        .Q(g971) );
  SDFFX1 DFF_659_Q_reg ( .D(g971), .SI(g971), .SE(n9140), .CLK(n9327), .Q(
        n8021), .QN(DFF_659_n1) );
  SDFFX1 DFF_660_Q_reg ( .D(n4375), .SI(n8021), .SE(n9140), .CLK(n9327), .Q(
        g973) );
  SDFFX1 DFF_661_Q_reg ( .D(g973), .SI(g973), .SE(n9140), .CLK(n9327), .Q(
        n8020), .QN(DFF_661_n1) );
  SDFFX1 DFF_662_Q_reg ( .D(n4379), .SI(n8020), .SE(n9140), .CLK(n9327), .Q(
        g975) );
  SDFFX1 DFF_663_Q_reg ( .D(g975), .SI(g975), .SE(n9140), .CLK(n9327), .Q(
        n8019), .QN(DFF_663_n1) );
  SDFFX1 DFF_664_Q_reg ( .D(g2873), .SI(n8019), .SE(n9141), .CLK(n9328), .Q(
        g977) );
  SDFFX1 DFF_665_Q_reg ( .D(g977), .SI(g977), .SE(n9141), .CLK(n9328), .Q(
        n8018), .QN(n4486) );
  SDFFX1 DFF_666_Q_reg ( .D(n4283), .SI(n8018), .SE(n9188), .CLK(n9375), .Q(
        g986), .QN(n4432) );
  SDFFX1 DFF_667_Q_reg ( .D(n467), .SI(g986), .SE(n9191), .CLK(n9378), .Q(g992), .QN(n8824) );
  SDFFX1 DFF_678_Q_reg ( .D(n4277), .SI(g992), .SE(n9191), .CLK(n9378), .Q(
        n8017) );
  SDFFX1 DFF_679_Q_reg ( .D(g1041), .SI(n8017), .SE(n9191), .CLK(n9378), .Q(
        g1029) );
  SDFFX1 DFF_680_Q_reg ( .D(g1029), .SI(g1029), .SE(n9192), .CLK(n9379), .Q(
        g1036) );
  SDFFX1 DFF_681_Q_reg ( .D(g1030), .SI(g1036), .SE(n9192), .CLK(n9379), .Q(
        g1037) );
  SDFFX1 DFF_682_Q_reg ( .D(g1037), .SI(g1037), .SE(n9192), .CLK(n9379), .Q(
        g1038) );
  SDFFX1 DFF_683_Q_reg ( .D(g1033), .SI(g1038), .SE(n9192), .CLK(n9379), .Q(
        test_so41) );
  SDFFX1 DFF_684_Q_reg ( .D(test_so41), .SI(test_si42), .SE(n9192), .CLK(n9379), .Q(g1040) );
  SDFFX1 DFF_685_Q_reg ( .D(g1056), .SI(g1040), .SE(n9192), .CLK(n9379), .Q(
        g1044) );
  SDFFX1 DFF_686_Q_reg ( .D(g1044), .SI(g1044), .SE(n9192), .CLK(n9379), .Q(
        g1051) );
  SDFFX1 DFF_687_Q_reg ( .D(g1045), .SI(g1051), .SE(n9192), .CLK(n9379), .Q(
        g1052) );
  SDFFX1 DFF_688_Q_reg ( .D(g1052), .SI(g1052), .SE(n9192), .CLK(n9379), .Q(
        g1053) );
  SDFFX1 DFF_689_Q_reg ( .D(g1048), .SI(g1053), .SE(n9192), .CLK(n9379), .Q(
        g1054) );
  SDFFX1 DFF_690_Q_reg ( .D(g1054), .SI(g1054), .SE(n9192), .CLK(n9379), .Q(
        g1055) );
  SDFFX1 DFF_691_Q_reg ( .D(test_so37), .SI(g1055), .SE(n9192), .CLK(n9379), 
        .Q(g1059) );
  SDFFX1 DFF_692_Q_reg ( .D(g1059), .SI(g1059), .SE(n9193), .CLK(n9380), .Q(
        g1066) );
  SDFFX1 DFF_693_Q_reg ( .D(g1060), .SI(g1066), .SE(n9193), .CLK(n9380), .Q(
        g1067) );
  SDFFX1 DFF_694_Q_reg ( .D(g1067), .SI(g1067), .SE(n9193), .CLK(n9380), .Q(
        g1068) );
  SDFFX1 DFF_695_Q_reg ( .D(g1063), .SI(g1068), .SE(n9193), .CLK(n9380), .Q(
        g1069) );
  SDFFX1 DFF_696_Q_reg ( .D(g1069), .SI(g1069), .SE(n9193), .CLK(n9380), .Q(
        g1070) );
  SDFFX1 DFF_697_Q_reg ( .D(g1085), .SI(g1070), .SE(n9193), .CLK(n9380), .Q(
        g1074) );
  SDFFX1 DFF_698_Q_reg ( .D(g1074), .SI(g1074), .SE(n9193), .CLK(n9380), .Q(
        g1081) );
  SDFFX1 DFF_699_Q_reg ( .D(g1075), .SI(g1081), .SE(n9193), .CLK(n9380), .Q(
        test_so42) );
  SDFFX1 DFF_700_Q_reg ( .D(test_so42), .SI(test_si43), .SE(n9193), .CLK(n9380), .Q(g1083) );
  SDFFX1 DFF_701_Q_reg ( .D(g1078), .SI(g1083), .SE(n9193), .CLK(n9380), .Q(
        g1084) );
  SDFFX1 DFF_702_Q_reg ( .D(g1084), .SI(g1084), .SE(n9193), .CLK(n9380), .Q(
        g1011) );
  SDFFX1 DFF_703_Q_reg ( .D(n4598), .SI(g1011), .SE(n9193), .CLK(n9380), .Q(
        g5657) );
  SDFFX1 DFF_704_Q_reg ( .D(g5657), .SI(g5657), .SE(n9194), .CLK(n9381), .Q(
        g5686) );
  SDFFX1 DFF_705_Q_reg ( .D(g5686), .SI(g5686), .SE(n9194), .CLK(n9381), .Q(
        g1024) );
  SDFFX1 DFF_706_Q_reg ( .D(n4598), .SI(g1024), .SE(n9194), .CLK(n9381), .Q(
        g6750), .QN(n4371) );
  SDFFX1 DFF_707_Q_reg ( .D(g6750), .SI(g6750), .SE(n9194), .CLK(n9381), .Q(
        g6944), .QN(n4316) );
  SDFFX1 DFF_708_Q_reg ( .D(g6944), .SI(g6944), .SE(n9194), .CLK(n9381), .Q(
        g1236), .QN(n4300) );
  SDFFX1 DFF_709_Q_reg ( .D(g21843), .SI(g1236), .SE(n9194), .CLK(n9381), .Q(
        g1240), .QN(n9052) );
  SDFFX1 DFF_710_Q_reg ( .D(g18707), .SI(g1240), .SE(n9194), .CLK(n9381), .Q(
        g1243), .QN(n4353) );
  SDFFX1 DFF_711_Q_reg ( .D(g18763), .SI(g1243), .SE(n9194), .CLK(n9381), .Q(
        g1196), .QN(n4304) );
  SDFFX1 DFF_712_Q_reg ( .D(n785), .SI(g1196), .SE(n9195), .CLK(n9382), .Q(
        g1199) );
  SDFFX1 DFF_713_Q_reg ( .D(g1199), .SI(g1199), .SE(n9195), .CLK(n9382), .Q(
        g1209) );
  SDFFX1 DFF_714_Q_reg ( .D(g1209), .SI(g1209), .SE(n9195), .CLK(n9382), .Q(
        g1210) );
  SDFFX1 DFF_715_Q_reg ( .D(g1142), .SI(g1210), .SE(n9195), .CLK(n9382), .Q(
        test_so43) );
  SDFFX1 DFF_716_Q_reg ( .D(test_so43), .SI(test_si44), .SE(n9196), .CLK(n9383), .Q(g1255) );
  SDFFX1 DFF_717_Q_reg ( .D(g1145), .SI(g1255), .SE(n9196), .CLK(n9383), .Q(
        g1256) );
  SDFFX1 DFF_718_Q_reg ( .D(g1256), .SI(g1256), .SE(n9196), .CLK(n9383), .Q(
        g1257) );
  SDFFX1 DFF_719_Q_reg ( .D(g1148), .SI(g1257), .SE(n9196), .CLK(n9383), .Q(
        g1258) );
  SDFFX1 DFF_720_Q_reg ( .D(g1258), .SI(g1258), .SE(n9196), .CLK(n9383), .Q(
        g1259) );
  SDFFX1 DFF_721_Q_reg ( .D(g1152), .SI(g1259), .SE(n9196), .CLK(n9383), .Q(
        g1260) );
  SDFFX1 DFF_722_Q_reg ( .D(g1260), .SI(g1260), .SE(n9196), .CLK(n9383), .Q(
        g1251) );
  SDFFX1 DFF_723_Q_reg ( .D(g1155), .SI(g1251), .SE(n9196), .CLK(n9383), .Q(
        g1252) );
  SDFFX1 DFF_724_Q_reg ( .D(g1252), .SI(g1252), .SE(n9196), .CLK(n9383), .Q(
        g1253) );
  SDFFX1 DFF_725_Q_reg ( .D(g1158), .SI(g1253), .SE(n9196), .CLK(n9383), .Q(
        g1254) );
  SDFFX1 DFF_726_Q_reg ( .D(g1254), .SI(g1254), .SE(n9196), .CLK(n9383), .Q(
        g1176) );
  SDFFX1 DFF_727_Q_reg ( .D(g2950), .SI(g1176), .SE(n9196), .CLK(n9383), .Q(
        g7961), .QN(n4460) );
  SDFFX1 DFF_728_Q_reg ( .D(g7961), .SI(g7961), .SE(n9197), .CLK(n9384), .Q(
        g8007), .QN(n4459) );
  SDFFX1 DFF_729_Q_reg ( .D(g8007), .SI(g8007), .SE(n9197), .CLK(n9384), .Q(
        g1172), .QN(n4465) );
  SDFFX1 DFF_730_Q_reg ( .D(g23081), .SI(g1172), .SE(n9198), .CLK(n9385), .Q(
        g1173) );
  SDFFX1 DFF_731_Q_reg ( .D(g23111), .SI(g1173), .SE(n9198), .CLK(n9385), .Q(
        test_so44) );
  SDFFX1 DFF_732_Q_reg ( .D(g23126), .SI(test_si45), .SE(n9197), .CLK(n9384), 
        .Q(g1175) );
  SDFFX1 DFF_733_Q_reg ( .D(g23392), .SI(g1175), .SE(n9197), .CLK(n9384), .Q(
        g1142) );
  SDFFX1 DFF_734_Q_reg ( .D(g23406), .SI(g1142), .SE(n9197), .CLK(n9384), .Q(
        g1145) );
  SDFFX1 DFF_735_Q_reg ( .D(g24179), .SI(g1145), .SE(n9197), .CLK(n9384), .Q(
        g1148) );
  SDFFX1 DFF_736_Q_reg ( .D(g24181), .SI(g1148), .SE(n9197), .CLK(n9384), .Q(
        g1164) );
  SDFFX1 DFF_737_Q_reg ( .D(g24213), .SI(g1164), .SE(n9197), .CLK(n9384), .Q(
        g1165) );
  SDFFX1 DFF_738_Q_reg ( .D(g24223), .SI(g1165), .SE(n9197), .CLK(n9384), .Q(
        g1166) );
  SDFFX1 DFF_739_Q_reg ( .D(g23110), .SI(g1166), .SE(n9197), .CLK(n9384), .Q(
        g1167) );
  SDFFX1 DFF_740_Q_reg ( .D(g23014), .SI(g1167), .SE(n9197), .CLK(n9384), .Q(
        g1171) );
  SDFFX1 DFF_741_Q_reg ( .D(g23039), .SI(g1171), .SE(n9197), .CLK(n9384), .Q(
        g1151) );
  SDFFX1 DFF_742_Q_reg ( .D(g24212), .SI(g1151), .SE(n9198), .CLK(n9385), .Q(
        g1152) );
  SDFFX1 DFF_743_Q_reg ( .D(g24222), .SI(g1152), .SE(n9198), .CLK(n9385), .Q(
        g1155) );
  SDFFX1 DFF_744_Q_reg ( .D(g24235), .SI(g1155), .SE(n9198), .CLK(n9385), .Q(
        g1158) );
  SDFFX1 DFF_745_Q_reg ( .D(n811), .SI(g1158), .SE(n9198), .CLK(n9385), .Q(
        g1214) );
  SDFFX1 DFF_746_Q_reg ( .D(g1214), .SI(g1214), .SE(n9198), .CLK(n9385), .Q(
        g1221) );
  SDFFX1 DFF_747_Q_reg ( .D(g1221), .SI(g1221), .SE(n9198), .CLK(n9385), .Q(
        test_so45) );
  SDFFX1 DFF_748_Q_reg ( .D(g13155), .SI(test_si46), .SE(n9198), .CLK(n9385), 
        .Q(g1229) );
  SDFFX1 DFF_749_Q_reg ( .D(g1229), .SI(g1229), .SE(n9198), .CLK(n9385), .Q(
        n4549), .QN(n8268) );
  SDFFX1 DFF_750_Q_reg ( .D(n486), .SI(n4549), .SE(n9199), .CLK(n9386), .Q(
        n4361), .QN(n8269) );
  SDFFX1 DFF_751_Q_reg ( .D(g13124), .SI(n4361), .SE(n9198), .CLK(n9385), .Q(
        g1235) );
  SDFFX1 DFF_752_Q_reg ( .D(g1235), .SI(g1235), .SE(n9198), .CLK(n9385), .Q(
        g1186), .QN(n4548) );
  SDFFX1 DFF_753_Q_reg ( .D(g13171), .SI(g1186), .SE(n9199), .CLK(n9386), .Q(
        g1244) );
  SDFFX1 DFF_754_Q_reg ( .D(g1244), .SI(g1244), .SE(n9199), .CLK(n9386), .Q(
        g1245) );
  SDFFX1 DFF_755_Q_reg ( .D(g27273), .SI(g1245), .SE(n9199), .CLK(n9386), .Q(
        g1262), .QN(n8447) );
  SDFFX1 DFF_756_Q_reg ( .D(g27285), .SI(g1262), .SE(n9199), .CLK(n9386), .Q(
        g1263), .QN(n8449) );
  SDFFX1 DFF_757_Q_reg ( .D(g27299), .SI(g1263), .SE(n9199), .CLK(n9386), .Q(
        g1261), .QN(n8448) );
  SDFFX1 DFF_758_Q_reg ( .D(g27286), .SI(g1261), .SE(n9200), .CLK(n9387), .Q(
        g1265), .QN(n8459) );
  SDFFX1 DFF_759_Q_reg ( .D(g27300), .SI(g1265), .SE(n9200), .CLK(n9387), .Q(
        g1266), .QN(n8461) );
  SDFFX1 DFF_760_Q_reg ( .D(g27314), .SI(g1266), .SE(n9199), .CLK(n9386), .Q(
        g1264), .QN(n8460) );
  SDFFX1 DFF_761_Q_reg ( .D(g27301), .SI(g1264), .SE(n9199), .CLK(n9386), .Q(
        g1268), .QN(n8292) );
  SDFFX1 DFF_762_Q_reg ( .D(g27315), .SI(g1268), .SE(n9199), .CLK(n9386), .Q(
        g1269), .QN(n8293) );
  SDFFX1 DFF_763_Q_reg ( .D(g27328), .SI(g1269), .SE(n9199), .CLK(n9386), .Q(
        test_so46) );
  SDFFX1 DFF_764_Q_reg ( .D(g27316), .SI(test_si47), .SE(n9199), .CLK(n9386), 
        .Q(g1271), .QN(n8469) );
  SDFFX1 DFF_765_Q_reg ( .D(g27329), .SI(g1271), .SE(n9200), .CLK(n9387), .Q(
        g1272), .QN(n8471) );
  SDFFX1 DFF_766_Q_reg ( .D(g27339), .SI(g1272), .SE(n9200), .CLK(n9387), .Q(
        g1270), .QN(n8470) );
  SDFFX1 DFF_767_Q_reg ( .D(g24501), .SI(g1270), .SE(n9200), .CLK(n9387), .Q(
        g1273) );
  SDFFX1 DFF_768_Q_reg ( .D(g24510), .SI(g1273), .SE(n9200), .CLK(n9387), .Q(
        g1276) );
  SDFFX1 DFF_769_Q_reg ( .D(g24521), .SI(g1276), .SE(n9200), .CLK(n9387), .Q(
        g1279) );
  SDFFX1 DFF_770_Q_reg ( .D(g24511), .SI(g1279), .SE(n9200), .CLK(n9387), .Q(
        g1282) );
  SDFFX1 DFF_771_Q_reg ( .D(g24522), .SI(g1282), .SE(n9200), .CLK(n9387), .Q(
        g1285) );
  SDFFX1 DFF_772_Q_reg ( .D(g24532), .SI(g1285), .SE(n9200), .CLK(n9387), .Q(
        g1288) );
  SDFFX1 DFF_773_Q_reg ( .D(g28351), .SI(g1288), .SE(n9200), .CLK(n9387), .Q(
        g1300) );
  SDFFX1 DFF_774_Q_reg ( .D(g28355), .SI(g1300), .SE(n9200), .CLK(n9387), .Q(
        g1303) );
  SDFFX1 DFF_775_Q_reg ( .D(g28360), .SI(g1303), .SE(n9199), .CLK(n9386), .Q(
        g1306) );
  SDFFX1 DFF_776_Q_reg ( .D(g28346), .SI(g1306), .SE(n9201), .CLK(n9388), .Q(
        g1291) );
  SDFFX1 DFF_777_Q_reg ( .D(g28350), .SI(g1291), .SE(n9201), .CLK(n9388), .Q(
        g1294) );
  SDFFX1 DFF_778_Q_reg ( .D(g28354), .SI(g1294), .SE(n9201), .CLK(n9388), .Q(
        g1297) );
  SDFFX1 DFF_779_Q_reg ( .D(g26547), .SI(g1297), .SE(n9201), .CLK(n9388), .Q(
        test_so47) );
  SDFFX1 DFF_780_Q_reg ( .D(g26557), .SI(test_si48), .SE(n9201), .CLK(n9388), 
        .Q(g1180) );
  SDFFX1 DFF_781_Q_reg ( .D(g26569), .SI(g1180), .SE(n9201), .CLK(n9388), .Q(
        g1183) );
  SDFFX1 DFF_782_Q_reg ( .D(g1186), .SI(g1183), .SE(n9201), .CLK(n9388), .Q(
        g1192), .QN(n4454) );
  SDFFX1 DFF_783_Q_reg ( .D(g22615), .SI(g1192), .SE(n9201), .CLK(n9388), .Q(
        n8009), .QN(DFF_783_n1) );
  SDFFX1 DFF_792_Q_reg ( .D(n516), .SI(n8009), .SE(n9201), .CLK(n9388), .Q(
        g16355), .QN(DFF_792_n1) );
  SDFFX1 DFF_793_Q_reg ( .D(g16355), .SI(g16355), .SE(n9202), .CLK(n9389), .Q(
        g1211), .QN(n8827) );
  SDFFX1 DFF_794_Q_reg ( .D(DFF_649_n1), .SI(g1211), .SE(n9202), .CLK(n9389), 
        .Q(n8008) );
  SDFFX1 DFF_795_Q_reg ( .D(DFF_651_n1), .SI(n8008), .SE(n9202), .CLK(n9389), 
        .Q(n8007) );
  SDFFX1 DFF_796_Q_reg ( .D(DFF_653_n1), .SI(n8007), .SE(n9202), .CLK(n9389), 
        .Q(n8006) );
  SDFFX1 DFF_797_Q_reg ( .D(DFF_655_n1), .SI(n8006), .SE(n9202), .CLK(n9389), 
        .Q(n8005) );
  SDFFX1 DFF_798_Q_reg ( .D(DFF_657_n1), .SI(n8005), .SE(n9202), .CLK(n9389), 
        .Q(n8004) );
  SDFFX1 DFF_799_Q_reg ( .D(DFF_659_n1), .SI(n8004), .SE(n9202), .CLK(n9389), 
        .Q(n8003) );
  SDFFX1 DFF_800_Q_reg ( .D(DFF_661_n1), .SI(n8003), .SE(n9202), .CLK(n9389), 
        .Q(g1222) );
  SDFFX1 DFF_801_Q_reg ( .D(DFF_663_n1), .SI(g1222), .SE(n9202), .CLK(n9389), 
        .Q(g1223) );
  SDFFX1 DFF_802_Q_reg ( .D(g24072), .SI(g1223), .SE(n9202), .CLK(n9389), .Q(
        g1224), .QN(n4489) );
  SDFFX1 DFF_803_Q_reg ( .D(n4486), .SI(g1224), .SE(n9202), .CLK(n9389), .Q(
        test_so48) );
  SDFFX1 DFF_805_Q_reg ( .D(g6979), .SI(g6979), .SE(n9129), .CLK(n9316), .Q(
        g7161), .QN(n4358) );
  SDFFX1 DFF_806_Q_reg ( .D(g7161), .SI(g7161), .SE(n9129), .CLK(n9316), .Q(
        g1315), .QN(n4294) );
  SDFFX1 DFF_807_Q_reg ( .D(g16671), .SI(g1315), .SE(n9194), .CLK(n9381), .Q(
        g1316), .QN(n9083) );
  SDFFX1 DFF_808_Q_reg ( .D(g20333), .SI(g1316), .SE(n9194), .CLK(n9381), .Q(
        g1345) );
  SDFFX1 DFF_809_Q_reg ( .D(g20717), .SI(g1345), .SE(n9194), .CLK(n9381), .Q(
        g1326), .QN(n4402) );
  SDFFX1 DFF_810_Q_reg ( .D(g21969), .SI(g1326), .SE(n9194), .CLK(n9381), .Q(
        g1319), .QN(n4476) );
  SDFFX1 DFF_811_Q_reg ( .D(g23329), .SI(g1319), .SE(n9195), .CLK(n9382), .Q(
        g1339), .QN(n4421) );
  SDFFX1 DFF_812_Q_reg ( .D(g24430), .SI(g1339), .SE(n9195), .CLK(n9382), .Q(
        g1332), .QN(n4412) );
  SDFFX1 DFF_813_Q_reg ( .D(g25189), .SI(g1332), .SE(n9195), .CLK(n9382), .Q(
        g1346), .QN(n4401) );
  SDFFX1 DFF_814_Q_reg ( .D(g26666), .SI(g1346), .SE(n9195), .CLK(n9382), .Q(
        g1358), .QN(n4411) );
  SDFFX1 DFF_815_Q_reg ( .D(g26781), .SI(g1358), .SE(n9195), .CLK(n9382), .Q(
        g1352), .QN(n4469) );
  SDFFX1 DFF_816_Q_reg ( .D(g27678), .SI(g1352), .SE(n9195), .CLK(n9382), .Q(
        g1365), .QN(n4475) );
  SDFFX1 DFF_817_Q_reg ( .D(g27718), .SI(g1365), .SE(n9195), .CLK(n9382), .Q(
        g1372), .QN(n4395) );
  SDFFX1 DFF_818_Q_reg ( .D(g28321), .SI(g1372), .SE(n9195), .CLK(n9382), .Q(
        g1378), .QN(n4417) );
  SDFFX1 DFF_819_Q_reg ( .D(g20882), .SI(g1378), .SE(n9202), .CLK(n9389), .Q(
        test_so49) );
  SDFFX1 DFF_820_Q_reg ( .D(g20896), .SI(test_si50), .SE(n9203), .CLK(n9390), 
        .Q(g1386), .QN(n8922) );
  SDFFX1 DFF_821_Q_reg ( .D(g20910), .SI(g1386), .SE(n9203), .CLK(n9390), .Q(
        g1384), .QN(n8968) );
  SDFFX1 DFF_822_Q_reg ( .D(g20897), .SI(g1384), .SE(n9203), .CLK(n9390), .Q(
        g1388), .QN(n8921) );
  SDFFX1 DFF_823_Q_reg ( .D(g20911), .SI(g1388), .SE(n9203), .CLK(n9390), .Q(
        g1389), .QN(n8920) );
  SDFFX1 DFF_824_Q_reg ( .D(g20925), .SI(g1389), .SE(n9203), .CLK(n9390), .Q(
        g1387), .QN(n8967) );
  SDFFX1 DFF_825_Q_reg ( .D(g20912), .SI(g1387), .SE(n9203), .CLK(n9390), .Q(
        g1391), .QN(n8919) );
  SDFFX1 DFF_826_Q_reg ( .D(g20926), .SI(g1391), .SE(n9203), .CLK(n9390), .Q(
        g1392), .QN(n8918) );
  SDFFX1 DFF_827_Q_reg ( .D(g20949), .SI(g1392), .SE(n9203), .CLK(n9390), .Q(
        g1390), .QN(n8966) );
  SDFFX1 DFF_828_Q_reg ( .D(g20927), .SI(g1390), .SE(n9203), .CLK(n9390), .Q(
        g1394), .QN(n8917) );
  SDFFX1 DFF_829_Q_reg ( .D(g20950), .SI(g1394), .SE(n9203), .CLK(n9390), .Q(
        g1395), .QN(n8916) );
  SDFFX1 DFF_830_Q_reg ( .D(g20972), .SI(g1395), .SE(n9203), .CLK(n9390), .Q(
        g1393), .QN(n8965) );
  SDFFX1 DFF_831_Q_reg ( .D(g20951), .SI(g1393), .SE(n9203), .CLK(n9390), .Q(
        g1397), .QN(n8915) );
  SDFFX1 DFF_832_Q_reg ( .D(g20973), .SI(g1397), .SE(n9204), .CLK(n9391), .Q(
        g1398), .QN(n8914) );
  SDFFX1 DFF_833_Q_reg ( .D(g20993), .SI(g1398), .SE(n9204), .CLK(n9391), .Q(
        g1396), .QN(n8964) );
  SDFFX1 DFF_834_Q_reg ( .D(g20974), .SI(g1396), .SE(n9204), .CLK(n9391), .Q(
        g1400), .QN(n8913) );
  SDFFX1 DFF_835_Q_reg ( .D(g20994), .SI(g1400), .SE(n9204), .CLK(n9391), .Q(
        test_so50) );
  SDFFX1 DFF_836_Q_reg ( .D(g21015), .SI(test_si51), .SE(n9204), .CLK(n9391), 
        .Q(g1399), .QN(n8963) );
  SDFFX1 DFF_837_Q_reg ( .D(g20995), .SI(g1399), .SE(n9204), .CLK(n9391), .Q(
        g1403), .QN(n8912) );
  SDFFX1 DFF_838_Q_reg ( .D(g21016), .SI(g1403), .SE(n9204), .CLK(n9391), .Q(
        g1404), .QN(n8911) );
  SDFFX1 DFF_839_Q_reg ( .D(g21033), .SI(g1404), .SE(n9204), .CLK(n9391), .Q(
        g1402), .QN(n8962) );
  SDFFX1 DFF_840_Q_reg ( .D(g21017), .SI(g1402), .SE(n9204), .CLK(n9391), .Q(
        g1406), .QN(n8910) );
  SDFFX1 DFF_841_Q_reg ( .D(g21034), .SI(g1406), .SE(n9204), .CLK(n9391), .Q(
        g1407), .QN(n8909) );
  SDFFX1 DFF_842_Q_reg ( .D(g21052), .SI(g1407), .SE(n9204), .CLK(n9391), .Q(
        g1405), .QN(n8961) );
  SDFFX1 DFF_843_Q_reg ( .D(g21035), .SI(g1405), .SE(n9204), .CLK(n9391), .Q(
        g1409), .QN(n8908) );
  SDFFX1 DFF_844_Q_reg ( .D(g21053), .SI(g1409), .SE(n9205), .CLK(n9392), .Q(
        g1410), .QN(n8907) );
  SDFFX1 DFF_845_Q_reg ( .D(g21070), .SI(g1410), .SE(n9205), .CLK(n9392), .Q(
        g1408), .QN(n8960) );
  SDFFX1 DFF_846_Q_reg ( .D(g20883), .SI(g1408), .SE(n9205), .CLK(n9392), .Q(
        g1412), .QN(n8906) );
  SDFFX1 DFF_847_Q_reg ( .D(g20898), .SI(g1412), .SE(n9205), .CLK(n9392), .Q(
        g1413), .QN(n8905) );
  SDFFX1 DFF_848_Q_reg ( .D(g20913), .SI(g1413), .SE(n9205), .CLK(n9392), .Q(
        g1411), .QN(n8959) );
  SDFFX1 DFF_849_Q_reg ( .D(g20952), .SI(g1411), .SE(n9205), .CLK(n9392), .Q(
        g1415), .QN(n8682) );
  SDFFX1 DFF_850_Q_reg ( .D(g20975), .SI(g1415), .SE(n9205), .CLK(n9392), .Q(
        g1416), .QN(n8674) );
  SDFFX1 DFF_851_Q_reg ( .D(g20996), .SI(g1416), .SE(n9205), .CLK(n9392), .Q(
        test_so51) );
  SDFFX1 DFF_852_Q_reg ( .D(g20976), .SI(test_si52), .SE(n9201), .CLK(n9388), 
        .Q(g1418), .QN(n8681) );
  SDFFX1 DFF_853_Q_reg ( .D(g20997), .SI(g1418), .SE(n9201), .CLK(n9388), .Q(
        g1419), .QN(n8673) );
  SDFFX1 DFF_854_Q_reg ( .D(g21018), .SI(g1419), .SE(n9201), .CLK(n9388), .Q(
        g1417), .QN(n8736) );
  SDFFX1 DFF_855_Q_reg ( .D(g25263), .SI(g1417), .SE(n9205), .CLK(n9392), .Q(
        g1421) );
  SDFFX1 DFF_856_Q_reg ( .D(g25267), .SI(g1421), .SE(n9205), .CLK(n9392), .Q(
        g1422) );
  SDFFX1 DFF_857_Q_reg ( .D(g25270), .SI(g1422), .SE(n9205), .CLK(n9392), .Q(
        g1420) );
  SDFFX1 DFF_858_Q_reg ( .D(g22234), .SI(g1420), .SE(n9205), .CLK(n9392), .Q(
        g1424) );
  SDFFX1 DFF_859_Q_reg ( .D(g22247), .SI(g1424), .SE(n9206), .CLK(n9393), .Q(
        g1425) );
  SDFFX1 DFF_860_Q_reg ( .D(g22263), .SI(g1425), .SE(n9206), .CLK(n9393), .Q(
        g1423) );
  SDFFX1 DFF_861_Q_reg ( .D(g2950), .SI(g1423), .SE(n9206), .CLK(n9393), .Q(
        g6573), .QN(n4317) );
  SDFFX1 DFF_862_Q_reg ( .D(g6573), .SI(g6573), .SE(n9206), .CLK(n9393), .Q(
        g6782), .QN(n4515) );
  SDFFX1 DFF_863_Q_reg ( .D(g6782), .SI(g6782), .SE(n9206), .CLK(n9393), .Q(
        g1547), .QN(n4368) );
  SDFFX1 DFF_864_Q_reg ( .D(g22149), .SI(g1547), .SE(n9206), .CLK(n9393), .Q(
        g1512) );
  SDFFX1 DFF_865_Q_reg ( .D(g22166), .SI(g1512), .SE(n9209), .CLK(n9396), .Q(
        g1513) );
  SDFFX1 DFF_866_Q_reg ( .D(g22178), .SI(g1513), .SE(n9209), .CLK(n9396), .Q(
        g1511) );
  SDFFX1 DFF_867_Q_reg ( .D(g22167), .SI(g1511), .SE(n9207), .CLK(n9394), .Q(
        test_so52) );
  SDFFX1 DFF_868_Q_reg ( .D(g22179), .SI(test_si53), .SE(n9210), .CLK(n9397), 
        .Q(g1516) );
  SDFFX1 DFF_869_Q_reg ( .D(g22191), .SI(g1516), .SE(n9210), .CLK(n9397), .Q(
        g1514) );
  SDFFX1 DFF_870_Q_reg ( .D(g22035), .SI(g1514), .SE(n9210), .CLK(n9397), .Q(
        g1524) );
  SDFFX1 DFF_871_Q_reg ( .D(g22043), .SI(g1524), .SE(n9210), .CLK(n9397), .Q(
        g1525) );
  SDFFX1 DFF_872_Q_reg ( .D(g22057), .SI(g1525), .SE(n9211), .CLK(n9398), .Q(
        g1523) );
  SDFFX1 DFF_873_Q_reg ( .D(g22044), .SI(g1523), .SE(n9211), .CLK(n9398), .Q(
        g1527) );
  SDFFX1 DFF_874_Q_reg ( .D(g22058), .SI(g1527), .SE(n9211), .CLK(n9398), .Q(
        g1528) );
  SDFFX1 DFF_875_Q_reg ( .D(g22073), .SI(g1528), .SE(n9211), .CLK(n9398), .Q(
        g1526) );
  SDFFX1 DFF_876_Q_reg ( .D(g22059), .SI(g1526), .SE(n9211), .CLK(n9398), .Q(
        g1530) );
  SDFFX1 DFF_877_Q_reg ( .D(g22074), .SI(g1530), .SE(n9211), .CLK(n9398), .Q(
        g1531) );
  SDFFX1 DFF_878_Q_reg ( .D(g22090), .SI(g1531), .SE(n9211), .CLK(n9398), .Q(
        g1529) );
  SDFFX1 DFF_879_Q_reg ( .D(g22075), .SI(g1529), .SE(n9211), .CLK(n9398), .Q(
        g1533) );
  SDFFX1 DFF_880_Q_reg ( .D(g22091), .SI(g1533), .SE(n9211), .CLK(n9398), .Q(
        g1534) );
  SDFFX1 DFF_881_Q_reg ( .D(g22112), .SI(g1534), .SE(n9211), .CLK(n9398), .Q(
        g1532) );
  SDFFX1 DFF_882_Q_reg ( .D(g22092), .SI(g1532), .SE(n9211), .CLK(n9398), .Q(
        g1536) );
  SDFFX1 DFF_883_Q_reg ( .D(g22113), .SI(g1536), .SE(n9211), .CLK(n9398), .Q(
        test_so53) );
  SDFFX1 DFF_884_Q_reg ( .D(g22130), .SI(test_si54), .SE(n9209), .CLK(n9396), 
        .Q(g1535) );
  SDFFX1 DFF_885_Q_reg ( .D(g22114), .SI(g1535), .SE(n9209), .CLK(n9396), .Q(
        g1539) );
  SDFFX1 DFF_886_Q_reg ( .D(g22131), .SI(g1539), .SE(n9209), .CLK(n9396), .Q(
        g1540) );
  SDFFX1 DFF_887_Q_reg ( .D(g22150), .SI(g1540), .SE(n9209), .CLK(n9396), .Q(
        g1538) );
  SDFFX1 DFF_888_Q_reg ( .D(g22132), .SI(g1538), .SE(n9209), .CLK(n9396), .Q(
        g1542) );
  SDFFX1 DFF_889_Q_reg ( .D(g22151), .SI(g1542), .SE(n9209), .CLK(n9396), .Q(
        g1543) );
  SDFFX1 DFF_890_Q_reg ( .D(g22168), .SI(g1543), .SE(n9209), .CLK(n9396), .Q(
        g1541) );
  SDFFX1 DFF_891_Q_reg ( .D(g22152), .SI(g1541), .SE(n9210), .CLK(n9397), .Q(
        g1545) );
  SDFFX1 DFF_892_Q_reg ( .D(g22169), .SI(g1545), .SE(n9209), .CLK(n9396), .Q(
        g1546) );
  SDFFX1 DFF_893_Q_reg ( .D(g22180), .SI(g1546), .SE(n9210), .CLK(n9397), .Q(
        g1544) );
  SDFFX1 DFF_894_Q_reg ( .D(g25217), .SI(g1544), .SE(n9210), .CLK(n9397), .Q(
        g1551), .QN(n8707) );
  SDFFX1 DFF_895_Q_reg ( .D(g25224), .SI(g1551), .SE(n9210), .CLK(n9397), .Q(
        g1552), .QN(n8706) );
  SDFFX1 DFF_896_Q_reg ( .D(g25233), .SI(g1552), .SE(n9210), .CLK(n9397), .Q(
        g1550), .QN(n8705) );
  SDFFX1 DFF_897_Q_reg ( .D(g25225), .SI(g1550), .SE(n9210), .CLK(n9397), .Q(
        g1554), .QN(n8704) );
  SDFFX1 DFF_898_Q_reg ( .D(g25234), .SI(g1554), .SE(n9210), .CLK(n9397), .Q(
        g1555), .QN(n8703) );
  SDFFX1 DFF_899_Q_reg ( .D(g25242), .SI(g1555), .SE(n9210), .CLK(n9397), .Q(
        test_so54) );
  SDFFX1 DFF_900_Q_reg ( .D(g25235), .SI(test_si55), .SE(n9206), .CLK(n9393), 
        .Q(g1557), .QN(n8702) );
  SDFFX1 DFF_901_Q_reg ( .D(g25243), .SI(g1557), .SE(n9206), .CLK(n9393), .Q(
        g1558), .QN(n8701) );
  SDFFX1 DFF_902_Q_reg ( .D(g25249), .SI(g1558), .SE(n9206), .CLK(n9393), .Q(
        g1556), .QN(n8700) );
  SDFFX1 DFF_903_Q_reg ( .D(g25244), .SI(g1556), .SE(n9206), .CLK(n9393), .Q(
        g1560), .QN(n8699) );
  SDFFX1 DFF_904_Q_reg ( .D(g25250), .SI(g1560), .SE(n9206), .CLK(n9393), .Q(
        g1561), .QN(n8698) );
  SDFFX1 DFF_905_Q_reg ( .D(g25255), .SI(g1561), .SE(n9206), .CLK(n9393), .Q(
        g1559) );
  SDFFX1 DFF_906_Q_reg ( .D(g30279), .SI(g1559), .SE(n9216), .CLK(n9403), .Q(
        g1567) );
  SDFFX1 DFF_907_Q_reg ( .D(g30287), .SI(g1567), .SE(n9216), .CLK(n9403), .Q(
        g1570) );
  SDFFX1 DFF_908_Q_reg ( .D(g30294), .SI(g1570), .SE(n9216), .CLK(n9403), .Q(
        g1573) );
  SDFFX1 DFF_909_Q_reg ( .D(g30651), .SI(g1573), .SE(n9216), .CLK(n9403), .Q(
        g1612) );
  SDFFX1 DFF_910_Q_reg ( .D(g30657), .SI(g1612), .SE(n9216), .CLK(n9403), .Q(
        g1615) );
  SDFFX1 DFF_911_Q_reg ( .D(g30663), .SI(g1615), .SE(n9216), .CLK(n9403), .Q(
        g1618) );
  SDFFX1 DFF_912_Q_reg ( .D(g30683), .SI(g1618), .SE(n9217), .CLK(n9404), .Q(
        g1576) );
  SDFFX1 DFF_913_Q_reg ( .D(g30688), .SI(g1576), .SE(n9217), .CLK(n9404), .Q(
        g1579) );
  SDFFX1 DFF_914_Q_reg ( .D(g30692), .SI(g1579), .SE(n9212), .CLK(n9399), .Q(
        g1582) );
  SDFFX1 DFF_915_Q_reg ( .D(g30658), .SI(g1582), .SE(n9212), .CLK(n9399), .Q(
        test_so55) );
  SDFFX1 DFF_916_Q_reg ( .D(g30664), .SI(test_si56), .SE(n9212), .CLK(n9399), 
        .Q(g1624) );
  SDFFX1 DFF_917_Q_reg ( .D(g30671), .SI(g1624), .SE(n9212), .CLK(n9399), .Q(
        g1627) );
  SDFFX1 DFF_918_Q_reg ( .D(g30295), .SI(g1627), .SE(n9212), .CLK(n9399), .Q(
        g1585) );
  SDFFX1 DFF_919_Q_reg ( .D(g30299), .SI(g1585), .SE(n9212), .CLK(n9399), .Q(
        g1588) );
  SDFFX1 DFF_920_Q_reg ( .D(g30302), .SI(g1588), .SE(n9212), .CLK(n9399), .Q(
        g1591) );
  SDFFX1 DFF_921_Q_reg ( .D(g30266), .SI(g1591), .SE(n9212), .CLK(n9399), .Q(
        g1630) );
  SDFFX1 DFF_922_Q_reg ( .D(g30272), .SI(g1630), .SE(n9212), .CLK(n9399), .Q(
        g1633) );
  SDFFX1 DFF_923_Q_reg ( .D(g30280), .SI(g1633), .SE(n9212), .CLK(n9399), .Q(
        g1636) );
  SDFFX1 DFF_924_Q_reg ( .D(g30250), .SI(g1636), .SE(n9212), .CLK(n9399), .Q(
        g1594) );
  SDFFX1 DFF_925_Q_reg ( .D(g30252), .SI(g1594), .SE(n9212), .CLK(n9399), .Q(
        g1597) );
  SDFFX1 DFF_926_Q_reg ( .D(g30255), .SI(g1597), .SE(n9213), .CLK(n9400), .Q(
        g1600) );
  SDFFX1 DFF_927_Q_reg ( .D(g30273), .SI(g1600), .SE(n9213), .CLK(n9400), .Q(
        g1639) );
  SDFFX1 DFF_928_Q_reg ( .D(g30281), .SI(g1639), .SE(n9213), .CLK(n9400), .Q(
        g1642) );
  SDFFX1 DFF_929_Q_reg ( .D(g30288), .SI(g1642), .SE(n9213), .CLK(n9400), .Q(
        g1645) );
  SDFFX1 DFF_930_Q_reg ( .D(g30644), .SI(g1645), .SE(n9213), .CLK(n9400), .Q(
        g1603) );
  SDFFX1 DFF_931_Q_reg ( .D(g30650), .SI(g1603), .SE(n9213), .CLK(n9400), .Q(
        test_so56) );
  SDFFX1 DFF_932_Q_reg ( .D(g30656), .SI(test_si57), .SE(n9207), .CLK(n9394), 
        .Q(g1609) );
  SDFFX1 DFF_933_Q_reg ( .D(g30678), .SI(g1609), .SE(n9207), .CLK(n9394), .Q(
        g1648) );
  SDFFX1 DFF_934_Q_reg ( .D(g30684), .SI(g1648), .SE(n9207), .CLK(n9394), .Q(
        g1651) );
  SDFFX1 DFF_935_Q_reg ( .D(g30689), .SI(g1651), .SE(n9207), .CLK(n9394), .Q(
        g1654) );
  SDFFX1 DFF_936_Q_reg ( .D(g25056), .SI(g1654), .SE(n9207), .CLK(n9394), .Q(
        g1466), .QN(n8813) );
  SDFFX1 DFF_937_Q_reg ( .D(g25938), .SI(g1466), .SE(n9207), .CLK(n9394), .Q(
        g1462), .QN(n9114) );
  SDFFX1 DFF_938_Q_reg ( .D(g26531), .SI(g1462), .SE(n9207), .CLK(n9394), .Q(
        g1457), .QN(n8812) );
  SDFFX1 DFF_939_Q_reg ( .D(g27129), .SI(g1457), .SE(n9207), .CLK(n9394), .Q(
        g1453), .QN(n9115) );
  SDFFX1 DFF_940_Q_reg ( .D(g27612), .SI(g1453), .SE(n9207), .CLK(n9394), .Q(
        g1448), .QN(n8811) );
  SDFFX1 DFF_941_Q_reg ( .D(g28147), .SI(g1448), .SE(n9208), .CLK(n9395), .Q(
        g1444), .QN(n9097) );
  SDFFX1 DFF_942_Q_reg ( .D(g28636), .SI(g1444), .SE(n9208), .CLK(n9395), .Q(
        g1439), .QN(n8810) );
  SDFFX1 DFF_943_Q_reg ( .D(g29111), .SI(g1439), .SE(n9208), .CLK(n9395), .Q(
        g1435), .QN(n9103) );
  SDFFX1 DFF_944_Q_reg ( .D(g29355), .SI(g1435), .SE(n9208), .CLK(n9395), .Q(
        g1430), .QN(n8438) );
  SDFFX1 DFF_945_Q_reg ( .D(g29581), .SI(g1430), .SE(n9208), .CLK(n9395), .Q(
        g1426), .QN(n8284) );
  SDFFX1 DFF_946_Q_reg ( .D(g13110), .SI(g1426), .SE(n9208), .CLK(n9395), .Q(
        g1562) );
  SDFFX1 DFF_947_Q_reg ( .D(g1562), .SI(g1562), .SE(n9208), .CLK(n9395), .Q(
        test_so57) );
  SDFFX1 DFF_948_Q_reg ( .D(test_so57), .SI(test_si58), .SE(n9208), .CLK(n9395), .Q(g1563), .QN(n9090) );
  SDFFX1 DFF_949_Q_reg ( .D(g2950), .SI(g1563), .SE(n9208), .CLK(n9395), .Q(
        g5511), .QN(n4518) );
  SDFFX1 DFF_952_Q_reg ( .D(test_so57), .SI(n4618), .SE(n9208), .CLK(n9395), 
        .Q(g1690), .QN(n4386) );
  SDFFX1 DFF_953_Q_reg ( .D(g27264), .SI(g1690), .SE(n9215), .CLK(n9402), .Q(
        g1735), .QN(n8767) );
  SDFFX1 DFF_954_Q_reg ( .D(g27274), .SI(g1735), .SE(n9216), .CLK(n9403), .Q(
        g1724), .QN(n8766) );
  SDFFX1 DFF_955_Q_reg ( .D(g27287), .SI(g1724), .SE(n9216), .CLK(n9403), .Q(
        g1727), .QN(n8765) );
  SDFFX1 DFF_956_Q_reg ( .D(g27275), .SI(g1727), .SE(n9216), .CLK(n9403), .Q(
        g1750), .QN(n8744) );
  SDFFX1 DFF_957_Q_reg ( .D(g27288), .SI(g1750), .SE(n9216), .CLK(n9403), .Q(
        g1739), .QN(n8743) );
  SDFFX1 DFF_958_Q_reg ( .D(g27302), .SI(g1739), .SE(n9215), .CLK(n9402), .Q(
        g1742), .QN(n8742) );
  SDFFX1 DFF_959_Q_reg ( .D(g27289), .SI(g1742), .SE(n9215), .CLK(n9402), .Q(
        g1765), .QN(n8489) );
  SDFFX1 DFF_960_Q_reg ( .D(g27303), .SI(g1765), .SE(n9215), .CLK(n9402), .Q(
        g1754), .QN(n8491) );
  SDFFX1 DFF_961_Q_reg ( .D(g27317), .SI(g1754), .SE(n9215), .CLK(n9402), .Q(
        g1757), .QN(n8490) );
  SDFFX1 DFF_962_Q_reg ( .D(g27304), .SI(g1757), .SE(n9216), .CLK(n9403), .Q(
        g1779), .QN(n8755) );
  SDFFX1 DFF_963_Q_reg ( .D(g27318), .SI(g1779), .SE(n9216), .CLK(n9403), .Q(
        test_so58) );
  SDFFX1 DFF_964_Q_reg ( .D(g27330), .SI(test_si59), .SE(n9213), .CLK(n9400), 
        .Q(g1772), .QN(n8754) );
  SDFFX1 DFF_965_Q_reg ( .D(g28749), .SI(g1772), .SE(n9213), .CLK(n9400), .Q(
        g1789) );
  SDFFX1 DFF_966_Q_reg ( .D(g28760), .SI(g1789), .SE(n9215), .CLK(n9402), .Q(
        g1792) );
  SDFFX1 DFF_967_Q_reg ( .D(g28771), .SI(g1792), .SE(n9215), .CLK(n9402), .Q(
        g1795) );
  SDFFX1 DFF_968_Q_reg ( .D(g29205), .SI(g1795), .SE(n9215), .CLK(n9402), .Q(
        g1798) );
  SDFFX1 DFF_969_Q_reg ( .D(g29212), .SI(g1798), .SE(n9215), .CLK(n9402), .Q(
        g1801) );
  SDFFX1 DFF_970_Q_reg ( .D(g29218), .SI(g1801), .SE(n9213), .CLK(n9400), .Q(
        g1804) );
  SDFFX1 DFF_971_Q_reg ( .D(g28761), .SI(g1804), .SE(n9214), .CLK(n9401), .Q(
        g1808), .QN(n8790) );
  SDFFX1 DFF_972_Q_reg ( .D(g28772), .SI(g1808), .SE(n9214), .CLK(n9401), .Q(
        g1809), .QN(n8778) );
  SDFFX1 DFF_973_Q_reg ( .D(g28778), .SI(g1809), .SE(n9214), .CLK(n9401), .Q(
        g1807), .QN(n8789) );
  SDFFX1 DFF_974_Q_reg ( .D(g26811), .SI(g1807), .SE(n9214), .CLK(n9401), .Q(
        g1810) );
  SDFFX1 DFF_975_Q_reg ( .D(g26815), .SI(g1810), .SE(n9214), .CLK(n9401), .Q(
        g1813) );
  SDFFX1 DFF_976_Q_reg ( .D(g26820), .SI(g1813), .SE(n9214), .CLK(n9401), .Q(
        g1816) );
  SDFFX1 DFF_977_Q_reg ( .D(g26816), .SI(g1816), .SE(n9214), .CLK(n9401), .Q(
        g1819) );
  SDFFX1 DFF_978_Q_reg ( .D(g26821), .SI(g1819), .SE(n9215), .CLK(n9402), .Q(
        g1822) );
  SDFFX1 DFF_979_Q_reg ( .D(g26824), .SI(g1822), .SE(n9215), .CLK(n9402), .Q(
        test_so59) );
  SDFFX1 DFF_980_Q_reg ( .D(g27764), .SI(test_si60), .SE(n9214), .CLK(n9401), 
        .Q(g1829), .QN(n8788) );
  SDFFX1 DFF_981_Q_reg ( .D(g27766), .SI(g1829), .SE(n9214), .CLK(n9401), .Q(
        g1830), .QN(n8777) );
  SDFFX1 DFF_982_Q_reg ( .D(g27768), .SI(g1830), .SE(n9214), .CLK(n9401), .Q(
        g1828), .QN(n8787) );
  SDFFX1 DFF_983_Q_reg ( .D(g29613), .SI(g1828), .SE(n9214), .CLK(n9401), .Q(
        g1693), .QN(n8394) );
  SDFFX1 DFF_984_Q_reg ( .D(g29617), .SI(g1693), .SE(n9214), .CLK(n9401), .Q(
        g1694), .QN(n8379) );
  SDFFX1 DFF_985_Q_reg ( .D(g29620), .SI(g1694), .SE(n9213), .CLK(n9400), .Q(
        g1695), .QN(n8393) );
  SDFFX1 DFF_986_Q_reg ( .D(g30704), .SI(g1695), .SE(n9213), .CLK(n9400), .Q(
        g1696), .QN(n8392) );
  SDFFX1 DFF_987_Q_reg ( .D(g30706), .SI(g1696), .SE(n9213), .CLK(n9400), .Q(
        g1697), .QN(n8378) );
  SDFFX1 DFF_988_Q_reg ( .D(g30708), .SI(g1697), .SE(n9207), .CLK(n9394), .Q(
        g1698), .QN(n8391) );
  SDFFX1 DFF_989_Q_reg ( .D(g30487), .SI(g1698), .SE(n9209), .CLK(n9396), .Q(
        g1699), .QN(n8390) );
  SDFFX1 DFF_990_Q_reg ( .D(g30503), .SI(g1699), .SE(n9207), .CLK(n9394), .Q(
        g1700), .QN(n8377) );
  SDFFX1 DFF_991_Q_reg ( .D(g30338), .SI(g1700), .SE(n9209), .CLK(n9396), .Q(
        g1701), .QN(n8389) );
  SDFFX1 DFF_992_Q_reg ( .D(g29178), .SI(g1701), .SE(n9217), .CLK(n9404), .Q(
        g1703) );
  SDFFX1 DFF_993_Q_reg ( .D(g29181), .SI(g1703), .SE(n9217), .CLK(n9404), .Q(
        g1704) );
  SDFFX1 DFF_994_Q_reg ( .D(g29184), .SI(g1704), .SE(n9217), .CLK(n9404), .Q(
        g1702) );
  SDFFX1 DFF_995_Q_reg ( .D(g26667), .SI(g1702), .SE(n9217), .CLK(n9404), .Q(
        test_so60) );
  SDFFX1 DFF_996_Q_reg ( .D(g26670), .SI(test_si61), .SE(n9217), .CLK(n9404), 
        .Q(g1785), .QN(n8776) );
  SDFFX1 DFF_997_Q_reg ( .D(g26675), .SI(g1785), .SE(n9217), .CLK(n9404), .Q(
        g1783), .QN(n8786) );
  SDFFX1 DFF_998_Q_reg ( .D(n4288), .SI(g1783), .SE(n9217), .CLK(n9404), .Q(
        g1831) );
  SDFFX1 DFF_999_Q_reg ( .D(g1831), .SI(g1831), .SE(n9217), .CLK(n9404), .Q(
        n7988), .QN(DFF_999_n1) );
  SDFFX1 DFF_1000_Q_reg ( .D(n4565), .SI(n7988), .SE(n9217), .CLK(n9404), .Q(
        g1833) );
  SDFFX1 DFF_1001_Q_reg ( .D(g1833), .SI(g1833), .SE(n9217), .CLK(n9404), .Q(
        n7987), .QN(DFF_1001_n1) );
  SDFFX1 DFF_1002_Q_reg ( .D(n4557), .SI(n7987), .SE(n9218), .CLK(n9405), .Q(
        g1835) );
  SDFFX1 DFF_1003_Q_reg ( .D(g1835), .SI(g1835), .SE(n9218), .CLK(n9405), .Q(
        n7986), .QN(DFF_1003_n1) );
  SDFFX1 DFF_1004_Q_reg ( .D(n4326), .SI(n7986), .SE(n9218), .CLK(n9405), .Q(
        g1661) );
  SDFFX1 DFF_1005_Q_reg ( .D(g1661), .SI(g1661), .SE(n9218), .CLK(n9405), .Q(
        n7985), .QN(DFF_1005_n1) );
  SDFFX1 DFF_1006_Q_reg ( .D(n4390), .SI(n7985), .SE(n9218), .CLK(n9405), .Q(
        g1663) );
  SDFFX1 DFF_1007_Q_reg ( .D(g1663), .SI(g1663), .SE(n9218), .CLK(n9405), .Q(
        n7984), .QN(DFF_1007_n1) );
  SDFFX1 DFF_1008_Q_reg ( .D(n4320), .SI(n7984), .SE(n9218), .CLK(n9405), .Q(
        g1665) );
  SDFFX1 DFF_1009_Q_reg ( .D(g1665), .SI(g1665), .SE(n9218), .CLK(n9405), .Q(
        n7983), .QN(DFF_1009_n1) );
  SDFFX1 DFF_1010_Q_reg ( .D(n4374), .SI(n7983), .SE(n9218), .CLK(n9405), .Q(
        g1667) );
  SDFFX1 DFF_1011_Q_reg ( .D(g1667), .SI(g1667), .SE(n9218), .CLK(n9405), .Q(
        test_so61), .QN(DFF_1011_n1) );
  SDFFX1 DFF_1012_Q_reg ( .D(n4378), .SI(test_si62), .SE(n9132), .CLK(n9319), 
        .Q(g1669) );
  SDFFX1 DFF_1013_Q_reg ( .D(g1669), .SI(g1669), .SE(n9132), .CLK(n9319), .Q(
        n7980), .QN(DFF_1013_n1) );
  SDFFX1 DFF_1014_Q_reg ( .D(g2877), .SI(n7980), .SE(n9138), .CLK(n9325), .Q(
        g1671) );
  SDFFX1 DFF_1015_Q_reg ( .D(g1671), .SI(g1671), .SE(n9138), .CLK(n9325), .Q(
        n7979), .QN(n4484) );
  SDFFX1 DFF_1016_Q_reg ( .D(n4284), .SI(n7979), .SE(n9215), .CLK(n9402), .Q(
        g1680), .QN(n4488) );
  SDFFX1 DFF_1017_Q_reg ( .D(n465), .SI(g1680), .SE(n9229), .CLK(n9416), .Q(
        g1686) );
  SDFFX1 DFF_1028_Q_reg ( .D(n4276), .SI(g1686), .SE(n9218), .CLK(n9405), .Q(
        n7978), .QN(n16491) );
  SDFFX1 DFF_1029_Q_reg ( .D(g1735), .SI(n7978), .SE(n9218), .CLK(n9405), .Q(
        g1723) );
  SDFFX1 DFF_1030_Q_reg ( .D(g1723), .SI(g1723), .SE(n9219), .CLK(n9406), .Q(
        g1730) );
  SDFFX1 DFF_1031_Q_reg ( .D(g1724), .SI(g1730), .SE(n9219), .CLK(n9406), .Q(
        g1731) );
  SDFFX1 DFF_1032_Q_reg ( .D(g1731), .SI(g1731), .SE(n9219), .CLK(n9406), .Q(
        g1732) );
  SDFFX1 DFF_1033_Q_reg ( .D(g1727), .SI(g1732), .SE(n9219), .CLK(n9406), .Q(
        g1733) );
  SDFFX1 DFF_1034_Q_reg ( .D(g1733), .SI(g1733), .SE(n9219), .CLK(n9406), .Q(
        g1734) );
  SDFFX1 DFF_1035_Q_reg ( .D(g1750), .SI(g1734), .SE(n9219), .CLK(n9406), .Q(
        g1738) );
  SDFFX1 DFF_1036_Q_reg ( .D(g1738), .SI(g1738), .SE(n9219), .CLK(n9406), .Q(
        g1745) );
  SDFFX1 DFF_1037_Q_reg ( .D(g1739), .SI(g1745), .SE(n9219), .CLK(n9406), .Q(
        test_so62) );
  SDFFX1 DFF_1038_Q_reg ( .D(test_so62), .SI(test_si63), .SE(n9219), .CLK(
        n9406), .Q(g1747) );
  SDFFX1 DFF_1039_Q_reg ( .D(g1742), .SI(g1747), .SE(n9219), .CLK(n9406), .Q(
        g1748) );
  SDFFX1 DFF_1040_Q_reg ( .D(g1748), .SI(g1748), .SE(n9219), .CLK(n9406), .Q(
        g1749) );
  SDFFX1 DFF_1041_Q_reg ( .D(g1765), .SI(g1749), .SE(n9219), .CLK(n9406), .Q(
        g1753) );
  SDFFX1 DFF_1042_Q_reg ( .D(g1753), .SI(g1753), .SE(n9220), .CLK(n9407), .Q(
        g1760) );
  SDFFX1 DFF_1043_Q_reg ( .D(g1754), .SI(g1760), .SE(n9220), .CLK(n9407), .Q(
        g1761) );
  SDFFX1 DFF_1044_Q_reg ( .D(g1761), .SI(g1761), .SE(n9220), .CLK(n9407), .Q(
        g1762) );
  SDFFX1 DFF_1045_Q_reg ( .D(g1757), .SI(g1762), .SE(n9220), .CLK(n9407), .Q(
        g1763) );
  SDFFX1 DFF_1046_Q_reg ( .D(g1763), .SI(g1763), .SE(n9220), .CLK(n9407), .Q(
        g1764) );
  SDFFX1 DFF_1047_Q_reg ( .D(g1779), .SI(g1764), .SE(n9220), .CLK(n9407), .Q(
        g1768) );
  SDFFX1 DFF_1048_Q_reg ( .D(g1768), .SI(g1768), .SE(n9220), .CLK(n9407), .Q(
        g1775) );
  SDFFX1 DFF_1049_Q_reg ( .D(test_so58), .SI(g1775), .SE(n9220), .CLK(n9407), 
        .Q(g1776) );
  SDFFX1 DFF_1050_Q_reg ( .D(g1776), .SI(g1776), .SE(n9220), .CLK(n9407), .Q(
        g1777) );
  SDFFX1 DFF_1051_Q_reg ( .D(g1772), .SI(g1777), .SE(n9220), .CLK(n9407), .Q(
        g1778) );
  SDFFX1 DFF_1052_Q_reg ( .D(g1778), .SI(g1778), .SE(n9220), .CLK(n9407), .Q(
        g1705) );
  SDFFX1 DFF_1053_Q_reg ( .D(n4598), .SI(g1705), .SE(n9220), .CLK(n9407), .Q(
        test_so63) );
  SDFFX1 DFF_1054_Q_reg ( .D(test_so63), .SI(test_si64), .SE(n9221), .CLK(
        n9408), .Q(g5738) );
  SDFFX1 DFF_1055_Q_reg ( .D(g5738), .SI(g5738), .SE(n9221), .CLK(n9408), .Q(
        g1718) );
  SDFFX1 DFF_1056_Q_reg ( .D(n4598), .SI(g1718), .SE(n9221), .CLK(n9408), .Q(
        g7052), .QN(n4296) );
  SDFFX1 DFF_1057_Q_reg ( .D(g7052), .SI(g7052), .SE(n9221), .CLK(n9408), .Q(
        g7194), .QN(n4315) );
  SDFFX1 DFF_1058_Q_reg ( .D(g7194), .SI(g7194), .SE(n9221), .CLK(n9408), .Q(
        g1930), .QN(n4366) );
  SDFFX1 DFF_1059_Q_reg ( .D(g21845), .SI(g1930), .SE(n9221), .CLK(n9408), .Q(
        g1934), .QN(n9051) );
  SDFFX1 DFF_1060_Q_reg ( .D(g18743), .SI(g1934), .SE(n9221), .CLK(n9408), .Q(
        g1937), .QN(n4311) );
  SDFFX1 DFF_1061_Q_reg ( .D(g18794), .SI(g1937), .SE(n9221), .CLK(n9408), .Q(
        g1890), .QN(n4297) );
  SDFFX1 DFF_1062_Q_reg ( .D(n1096), .SI(g1890), .SE(n9222), .CLK(n9409), .Q(
        g1893) );
  SDFFX1 DFF_1063_Q_reg ( .D(g1893), .SI(g1893), .SE(n9222), .CLK(n9409), .Q(
        g1903) );
  SDFFX1 DFF_1064_Q_reg ( .D(g1903), .SI(g1903), .SE(n9222), .CLK(n9409), .Q(
        g1904) );
  SDFFX1 DFF_1065_Q_reg ( .D(g1836), .SI(g1904), .SE(n9222), .CLK(n9409), .Q(
        g1944) );
  SDFFX1 DFF_1066_Q_reg ( .D(g1944), .SI(g1944), .SE(n9223), .CLK(n9410), .Q(
        g1949) );
  SDFFX1 DFF_1067_Q_reg ( .D(test_so65), .SI(g1949), .SE(n9223), .CLK(n9410), 
        .Q(g1950) );
  SDFFX1 DFF_1068_Q_reg ( .D(g1950), .SI(g1950), .SE(n9223), .CLK(n9410), .Q(
        g1951) );
  SDFFX1 DFF_1069_Q_reg ( .D(g1842), .SI(g1951), .SE(n9223), .CLK(n9410), .Q(
        test_so64) );
  SDFFX1 DFF_1070_Q_reg ( .D(test_so64), .SI(test_si65), .SE(n9223), .CLK(
        n9410), .Q(g1953) );
  SDFFX1 DFF_1071_Q_reg ( .D(g1846), .SI(g1953), .SE(n9223), .CLK(n9410), .Q(
        g1954) );
  SDFFX1 DFF_1072_Q_reg ( .D(g1954), .SI(g1954), .SE(n9223), .CLK(n9410), .Q(
        g1945) );
  SDFFX1 DFF_1073_Q_reg ( .D(g1849), .SI(g1945), .SE(n9223), .CLK(n9410), .Q(
        g1946) );
  SDFFX1 DFF_1074_Q_reg ( .D(g1946), .SI(g1946), .SE(n9223), .CLK(n9410), .Q(
        g1947) );
  SDFFX1 DFF_1075_Q_reg ( .D(g1852), .SI(g1947), .SE(n9223), .CLK(n9410), .Q(
        g1948) );
  SDFFX1 DFF_1076_Q_reg ( .D(g1948), .SI(g1948), .SE(n9223), .CLK(n9410), .Q(
        g1870) );
  SDFFX1 DFF_1077_Q_reg ( .D(g2950), .SI(g1870), .SE(n9223), .CLK(n9410), .Q(
        g8012), .QN(n4458) );
  SDFFX1 DFF_1078_Q_reg ( .D(g8012), .SI(g8012), .SE(n9224), .CLK(n9411), .Q(
        g8082), .QN(n4457) );
  SDFFX1 DFF_1079_Q_reg ( .D(g8082), .SI(g8082), .SE(n9224), .CLK(n9411), .Q(
        g1866), .QN(n4464) );
  SDFFX1 DFF_1080_Q_reg ( .D(g23097), .SI(g1866), .SE(n9225), .CLK(n9412), .Q(
        g1867) );
  SDFFX1 DFF_1081_Q_reg ( .D(g23124), .SI(g1867), .SE(n9225), .CLK(n9412), .Q(
        g1868) );
  SDFFX1 DFF_1082_Q_reg ( .D(g23137), .SI(g1868), .SE(n9225), .CLK(n9412), .Q(
        g1869) );
  SDFFX1 DFF_1083_Q_reg ( .D(g23400), .SI(g1869), .SE(n9225), .CLK(n9412), .Q(
        g1836) );
  SDFFX1 DFF_1084_Q_reg ( .D(g23413), .SI(g1836), .SE(n9225), .CLK(n9412), .Q(
        test_so65) );
  SDFFX1 DFF_1085_Q_reg ( .D(g24182), .SI(test_si66), .SE(n9224), .CLK(n9411), 
        .Q(g1842) );
  SDFFX1 DFF_1086_Q_reg ( .D(g24208), .SI(g1842), .SE(n9224), .CLK(n9411), .Q(
        g1858) );
  SDFFX1 DFF_1087_Q_reg ( .D(g24219), .SI(g1858), .SE(n9224), .CLK(n9411), .Q(
        g1859) );
  SDFFX1 DFF_1088_Q_reg ( .D(g24231), .SI(g1859), .SE(n9224), .CLK(n9411), .Q(
        g1860) );
  SDFFX1 DFF_1089_Q_reg ( .D(g23123), .SI(g1860), .SE(n9224), .CLK(n9411), .Q(
        g1861) );
  SDFFX1 DFF_1090_Q_reg ( .D(g23030), .SI(g1861), .SE(n9224), .CLK(n9411), .Q(
        g1865) );
  SDFFX1 DFF_1091_Q_reg ( .D(g23058), .SI(g1865), .SE(n9224), .CLK(n9411), .Q(
        g1845) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24218), .SI(g1845), .SE(n9224), .CLK(n9411), .Q(
        g1846) );
  SDFFX1 DFF_1093_Q_reg ( .D(g24230), .SI(g1846), .SE(n9224), .CLK(n9411), .Q(
        g1849) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24243), .SI(g1849), .SE(n9224), .CLK(n9411), .Q(
        g1852) );
  SDFFX1 DFF_1095_Q_reg ( .D(n1073), .SI(g1852), .SE(n9225), .CLK(n9412), .Q(
        g1908) );
  SDFFX1 DFF_1096_Q_reg ( .D(g1908), .SI(g1908), .SE(n9225), .CLK(n9412), .Q(
        g1915) );
  SDFFX1 DFF_1097_Q_reg ( .D(g1915), .SI(g1915), .SE(n9225), .CLK(n9412), .Q(
        g1922) );
  SDFFX1 DFF_1098_Q_reg ( .D(g13164), .SI(g1922), .SE(n9225), .CLK(n9412), .Q(
        g1923) );
  SDFFX1 DFF_1099_Q_reg ( .D(g1923), .SI(g1923), .SE(n9225), .CLK(n9412), .Q(
        test_so66), .QN(DFF_1099_n1) );
  SDFFX1 DFF_1100_Q_reg ( .D(n490), .SI(test_si67), .SE(n9226), .CLK(n9413), 
        .Q(n7971), .QN(DFF_1100_n1) );
  SDFFX1 DFF_1101_Q_reg ( .D(g13135), .SI(n7971), .SE(n9225), .CLK(n9412), .Q(
        g1929) );
  SDFFX1 DFF_1102_Q_reg ( .D(g1929), .SI(g1929), .SE(n9225), .CLK(n9412), .Q(
        g1880), .QN(n4545) );
  SDFFX1 DFF_1103_Q_reg ( .D(g13182), .SI(g1880), .SE(n9226), .CLK(n9413), .Q(
        g1938) );
  SDFFX1 DFF_1104_Q_reg ( .D(g1938), .SI(g1938), .SE(n9226), .CLK(n9413), .Q(
        g1939) );
  SDFFX1 DFF_1105_Q_reg ( .D(g27290), .SI(g1939), .SE(n9226), .CLK(n9413), .Q(
        g1956), .QN(n8444) );
  SDFFX1 DFF_1106_Q_reg ( .D(g27305), .SI(g1956), .SE(n9226), .CLK(n9413), .Q(
        g1957), .QN(n8446) );
  SDFFX1 DFF_1107_Q_reg ( .D(g27319), .SI(g1957), .SE(n9226), .CLK(n9413), .Q(
        g1955), .QN(n8445) );
  SDFFX1 DFF_1108_Q_reg ( .D(g27306), .SI(g1955), .SE(n9227), .CLK(n9414), .Q(
        g1959), .QN(n8456) );
  SDFFX1 DFF_1109_Q_reg ( .D(g27320), .SI(g1959), .SE(n9227), .CLK(n9414), .Q(
        g1960), .QN(n8458) );
  SDFFX1 DFF_1110_Q_reg ( .D(g27331), .SI(g1960), .SE(n9226), .CLK(n9413), .Q(
        g1958), .QN(n8457) );
  SDFFX1 DFF_1111_Q_reg ( .D(g27321), .SI(g1958), .SE(n9226), .CLK(n9413), .Q(
        g1962), .QN(n8289) );
  SDFFX1 DFF_1112_Q_reg ( .D(g27332), .SI(g1962), .SE(n9226), .CLK(n9413), .Q(
        g1963), .QN(n8291) );
  SDFFX1 DFF_1113_Q_reg ( .D(g27340), .SI(g1963), .SE(n9226), .CLK(n9413), .Q(
        g1961), .QN(n8290) );
  SDFFX1 DFF_1114_Q_reg ( .D(g27333), .SI(g1961), .SE(n9226), .CLK(n9413), .Q(
        test_so67), .QN(n9125) );
  SDFFX1 DFF_1115_Q_reg ( .D(g27341), .SI(test_si68), .SE(n9227), .CLK(n9414), 
        .Q(g1966), .QN(n8468) );
  SDFFX1 DFF_1116_Q_reg ( .D(g27346), .SI(g1966), .SE(n9227), .CLK(n9414), .Q(
        g1964), .QN(n8467) );
  SDFFX1 DFF_1117_Q_reg ( .D(g24513), .SI(g1964), .SE(n9227), .CLK(n9414), .Q(
        g1967) );
  SDFFX1 DFF_1118_Q_reg ( .D(g24524), .SI(g1967), .SE(n9227), .CLK(n9414), .Q(
        g1970) );
  SDFFX1 DFF_1119_Q_reg ( .D(g24534), .SI(g1970), .SE(n9227), .CLK(n9414), .Q(
        g1973) );
  SDFFX1 DFF_1120_Q_reg ( .D(g24525), .SI(g1973), .SE(n9227), .CLK(n9414), .Q(
        g1976) );
  SDFFX1 DFF_1121_Q_reg ( .D(g24535), .SI(g1976), .SE(n9227), .CLK(n9414), .Q(
        g1979) );
  SDFFX1 DFF_1122_Q_reg ( .D(g24545), .SI(g1979), .SE(n9227), .CLK(n9414), .Q(
        g1982) );
  SDFFX1 DFF_1123_Q_reg ( .D(g28357), .SI(g1982), .SE(n9227), .CLK(n9414), .Q(
        g1994) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28362), .SI(g1994), .SE(n9227), .CLK(n9414), .Q(
        g1997) );
  SDFFX1 DFF_1125_Q_reg ( .D(g28366), .SI(g1997), .SE(n9226), .CLK(n9413), .Q(
        g2000) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28352), .SI(g2000), .SE(n9228), .CLK(n9415), .Q(
        g1985) );
  SDFFX1 DFF_1127_Q_reg ( .D(g28356), .SI(g1985), .SE(n9228), .CLK(n9415), .Q(
        g1988) );
  SDFFX1 DFF_1128_Q_reg ( .D(g28361), .SI(g1988), .SE(n9228), .CLK(n9415), .Q(
        g1991) );
  SDFFX1 DFF_1129_Q_reg ( .D(g26559), .SI(g1991), .SE(n9228), .CLK(n9415), .Q(
        test_so68) );
  SDFFX1 DFF_1130_Q_reg ( .D(g26573), .SI(test_si69), .SE(n9228), .CLK(n9415), 
        .Q(g1874) );
  SDFFX1 DFF_1131_Q_reg ( .D(g26592), .SI(g1874), .SE(n9228), .CLK(n9415), .Q(
        g1877) );
  SDFFX1 DFF_1132_Q_reg ( .D(g1880), .SI(g1877), .SE(n9228), .CLK(n9415), .Q(
        g1886), .QN(n4493) );
  SDFFX1 DFF_1133_Q_reg ( .D(g22651), .SI(g1886), .SE(n9228), .CLK(n9415), .Q(
        n7968), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(n515), .SI(n7968), .SE(n9228), .CLK(n9415), .Q(
        g16399), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(g16399), .SI(g16399), .SE(n9228), .CLK(n9415), 
        .Q(g1905), .QN(n8826) );
  SDFFX1 DFF_1144_Q_reg ( .D(DFF_999_n1), .SI(g1905), .SE(n9228), .CLK(n9415), 
        .Q(n7967) );
  SDFFX1 DFF_1145_Q_reg ( .D(DFF_1001_n1), .SI(n7967), .SE(n9228), .CLK(n9415), 
        .Q(n7966) );
  SDFFX1 DFF_1146_Q_reg ( .D(DFF_1003_n1), .SI(n7966), .SE(n9229), .CLK(n9416), 
        .Q(n7965) );
  SDFFX1 DFF_1147_Q_reg ( .D(DFF_1005_n1), .SI(n7965), .SE(n9229), .CLK(n9416), 
        .Q(n7964) );
  SDFFX1 DFF_1148_Q_reg ( .D(DFF_1007_n1), .SI(n7964), .SE(n9229), .CLK(n9416), 
        .Q(n7963) );
  SDFFX1 DFF_1149_Q_reg ( .D(DFF_1009_n1), .SI(n7963), .SE(n9229), .CLK(n9416), 
        .Q(n7962) );
  SDFFX1 DFF_1150_Q_reg ( .D(DFF_1011_n1), .SI(n7962), .SE(n9229), .CLK(n9416), 
        .Q(g1916) );
  SDFFX1 DFF_1151_Q_reg ( .D(DFF_1013_n1), .SI(g1916), .SE(n9229), .CLK(n9416), 
        .Q(g1917) );
  SDFFX1 DFF_1152_Q_reg ( .D(g24083), .SI(g1917), .SE(n9229), .CLK(n9416), .Q(
        test_so69), .QN(n9127) );
  SDFFX1 DFF_1153_Q_reg ( .D(n4484), .SI(test_si70), .SE(n9138), .CLK(n9325), 
        .Q(n7960) );
  SDFFX1 DFF_1155_Q_reg ( .D(g7229), .SI(g7229), .SE(n9138), .CLK(n9325), .Q(
        g7357), .QN(n4357) );
  SDFFX1 DFF_1156_Q_reg ( .D(g7357), .SI(g7357), .SE(n9138), .CLK(n9325), .Q(
        g2009), .QN(n4293) );
  SDFFX1 DFF_1157_Q_reg ( .D(g16692), .SI(g2009), .SE(n9221), .CLK(n9408), .Q(
        g2010), .QN(n9084) );
  SDFFX1 DFF_1158_Q_reg ( .D(g20353), .SI(g2010), .SE(n9221), .CLK(n9408), .Q(
        g2039) );
  SDFFX1 DFF_1159_Q_reg ( .D(g20752), .SI(g2039), .SE(n9221), .CLK(n9408), .Q(
        g2020), .QN(n4400) );
  SDFFX1 DFF_1160_Q_reg ( .D(g21972), .SI(g2020), .SE(n9221), .CLK(n9408), .Q(
        g2013), .QN(n4474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g23339), .SI(g2013), .SE(n9222), .CLK(n9409), .Q(
        g2033), .QN(n4420) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24434), .SI(g2033), .SE(n9222), .CLK(n9409), .Q(
        g2026), .QN(n4410) );
  SDFFX1 DFF_1163_Q_reg ( .D(g25194), .SI(g2026), .SE(n9222), .CLK(n9409), .Q(
        g2040), .QN(n4399) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26671), .SI(g2040), .SE(n9222), .CLK(n9409), .Q(
        g2052), .QN(n4409) );
  SDFFX1 DFF_1165_Q_reg ( .D(g26789), .SI(g2052), .SE(n9222), .CLK(n9409), .Q(
        g2046), .QN(n4468) );
  SDFFX1 DFF_1166_Q_reg ( .D(g27682), .SI(g2046), .SE(n9222), .CLK(n9409), .Q(
        g2059), .QN(n4473) );
  SDFFX1 DFF_1167_Q_reg ( .D(g27722), .SI(g2059), .SE(n9222), .CLK(n9409), .Q(
        test_so70), .QN(n9124) );
  SDFFX1 DFF_1168_Q_reg ( .D(g28325), .SI(test_si71), .SE(n9222), .CLK(n9409), 
        .Q(g2072), .QN(n4416) );
  SDFFX1 DFF_1169_Q_reg ( .D(g20899), .SI(g2072), .SE(n9229), .CLK(n9416), .Q(
        g2079), .QN(n8904) );
  SDFFX1 DFF_1170_Q_reg ( .D(g20915), .SI(g2079), .SE(n9229), .CLK(n9416), .Q(
        g2080), .QN(n8903) );
  SDFFX1 DFF_1171_Q_reg ( .D(g20934), .SI(g2080), .SE(n9231), .CLK(n9418), .Q(
        g2078), .QN(n8958) );
  SDFFX1 DFF_1172_Q_reg ( .D(g20916), .SI(g2078), .SE(n9231), .CLK(n9418), .Q(
        g2082), .QN(n8902) );
  SDFFX1 DFF_1173_Q_reg ( .D(g20935), .SI(g2082), .SE(n9231), .CLK(n9418), .Q(
        g2083), .QN(n8901) );
  SDFFX1 DFF_1174_Q_reg ( .D(g20953), .SI(g2083), .SE(n9231), .CLK(n9418), .Q(
        g2081), .QN(n8957) );
  SDFFX1 DFF_1175_Q_reg ( .D(g20936), .SI(g2081), .SE(n9232), .CLK(n9419), .Q(
        g2085), .QN(n8900) );
  SDFFX1 DFF_1176_Q_reg ( .D(g20954), .SI(g2085), .SE(n9232), .CLK(n9419), .Q(
        g2086), .QN(n8899) );
  SDFFX1 DFF_1177_Q_reg ( .D(g20977), .SI(g2086), .SE(n9232), .CLK(n9419), .Q(
        g2084), .QN(n8956) );
  SDFFX1 DFF_1178_Q_reg ( .D(g20955), .SI(g2084), .SE(n9232), .CLK(n9419), .Q(
        g2088), .QN(n8898) );
  SDFFX1 DFF_1179_Q_reg ( .D(g20978), .SI(g2088), .SE(n9232), .CLK(n9419), .Q(
        g2089), .QN(n8897) );
  SDFFX1 DFF_1180_Q_reg ( .D(g20999), .SI(g2089), .SE(n9232), .CLK(n9419), .Q(
        g2087), .QN(n8955) );
  SDFFX1 DFF_1181_Q_reg ( .D(g20979), .SI(g2087), .SE(n9232), .CLK(n9419), .Q(
        g2091), .QN(n8896) );
  SDFFX1 DFF_1182_Q_reg ( .D(g21000), .SI(g2091), .SE(n9232), .CLK(n9419), .Q(
        test_so71) );
  SDFFX1 DFF_1183_Q_reg ( .D(g21019), .SI(test_si72), .SE(n9229), .CLK(n9416), 
        .Q(g2090), .QN(n8954) );
  SDFFX1 DFF_1184_Q_reg ( .D(g21001), .SI(g2090), .SE(n9229), .CLK(n9416), .Q(
        g2094), .QN(n8895) );
  SDFFX1 DFF_1185_Q_reg ( .D(g21020), .SI(g2094), .SE(n9230), .CLK(n9417), .Q(
        g2095), .QN(n8894) );
  SDFFX1 DFF_1186_Q_reg ( .D(g21039), .SI(g2095), .SE(n9230), .CLK(n9417), .Q(
        g2093), .QN(n8953) );
  SDFFX1 DFF_1187_Q_reg ( .D(g21021), .SI(g2093), .SE(n9230), .CLK(n9417), .Q(
        g2097), .QN(n8893) );
  SDFFX1 DFF_1188_Q_reg ( .D(g21040), .SI(g2097), .SE(n9230), .CLK(n9417), .Q(
        g2098), .QN(n8892) );
  SDFFX1 DFF_1189_Q_reg ( .D(g21054), .SI(g2098), .SE(n9230), .CLK(n9417), .Q(
        g2096), .QN(n8952) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21041), .SI(g2096), .SE(n9230), .CLK(n9417), .Q(
        g2100), .QN(n8891) );
  SDFFX1 DFF_1191_Q_reg ( .D(g21055), .SI(g2100), .SE(n9230), .CLK(n9417), .Q(
        g2101), .QN(n8890) );
  SDFFX1 DFF_1192_Q_reg ( .D(g21071), .SI(g2101), .SE(n9230), .CLK(n9417), .Q(
        g2099), .QN(n8951) );
  SDFFX1 DFF_1193_Q_reg ( .D(g21056), .SI(g2099), .SE(n9230), .CLK(n9417), .Q(
        g2103), .QN(n8889) );
  SDFFX1 DFF_1194_Q_reg ( .D(g21072), .SI(g2103), .SE(n9230), .CLK(n9417), .Q(
        g2104), .QN(n8888) );
  SDFFX1 DFF_1195_Q_reg ( .D(g21080), .SI(g2104), .SE(n9230), .CLK(n9417), .Q(
        g2102), .QN(n8950) );
  SDFFX1 DFF_1196_Q_reg ( .D(g20900), .SI(g2102), .SE(n9230), .CLK(n9417), .Q(
        g2106), .QN(n8887) );
  SDFFX1 DFF_1197_Q_reg ( .D(g20917), .SI(g2106), .SE(n9231), .CLK(n9418), .Q(
        test_so72) );
  SDFFX1 DFF_1198_Q_reg ( .D(g20937), .SI(test_si73), .SE(n9231), .CLK(n9418), 
        .Q(g2105), .QN(n8949) );
  SDFFX1 DFF_1199_Q_reg ( .D(g20980), .SI(g2105), .SE(n9231), .CLK(n9418), .Q(
        g2109), .QN(n8680) );
  SDFFX1 DFF_1200_Q_reg ( .D(g21002), .SI(g2109), .SE(n9231), .CLK(n9418), .Q(
        g2110), .QN(n8672) );
  SDFFX1 DFF_1201_Q_reg ( .D(g21022), .SI(g2110), .SE(n9231), .CLK(n9418), .Q(
        g2108), .QN(n8735) );
  SDFFX1 DFF_1202_Q_reg ( .D(g21003), .SI(g2108), .SE(n9231), .CLK(n9418), .Q(
        g2112), .QN(n8679) );
  SDFFX1 DFF_1203_Q_reg ( .D(g21023), .SI(g2112), .SE(n9231), .CLK(n9418), .Q(
        g2113), .QN(n8671) );
  SDFFX1 DFF_1204_Q_reg ( .D(g21042), .SI(g2113), .SE(n9231), .CLK(n9418), .Q(
        g2111), .QN(n8734) );
  SDFFX1 DFF_1205_Q_reg ( .D(g25268), .SI(g2111), .SE(n9232), .CLK(n9419), .Q(
        g2115) );
  SDFFX1 DFF_1206_Q_reg ( .D(g25271), .SI(g2115), .SE(n9232), .CLK(n9419), .Q(
        g2116) );
  SDFFX1 DFF_1207_Q_reg ( .D(g25279), .SI(g2116), .SE(n9232), .CLK(n9419), .Q(
        g2114) );
  SDFFX1 DFF_1208_Q_reg ( .D(g22249), .SI(g2114), .SE(n9232), .CLK(n9419), .Q(
        g2118) );
  SDFFX1 DFF_1209_Q_reg ( .D(g22267), .SI(g2118), .SE(n9233), .CLK(n9420), .Q(
        g2119) );
  SDFFX1 DFF_1210_Q_reg ( .D(g22280), .SI(g2119), .SE(n9234), .CLK(n9421), .Q(
        g2117) );
  SDFFX1 DFF_1211_Q_reg ( .D(g2950), .SI(g2117), .SE(n9234), .CLK(n9421), .Q(
        g6837), .QN(n4324) );
  SDFFX1 DFF_1212_Q_reg ( .D(g6837), .SI(g6837), .SE(n9234), .CLK(n9421), .Q(
        test_so73), .QN(n9119) );
  SDFFX1 DFF_1213_Q_reg ( .D(test_so73), .SI(test_si74), .SE(n9234), .CLK(
        n9421), .Q(g2241), .QN(n4367) );
  SDFFX1 DFF_1214_Q_reg ( .D(g22170), .SI(g2241), .SE(n9234), .CLK(n9421), .Q(
        g2206), .QN(n8997) );
  SDFFX1 DFF_1215_Q_reg ( .D(g22182), .SI(g2206), .SE(n9238), .CLK(n9425), .Q(
        g2207), .QN(n8996) );
  SDFFX1 DFF_1216_Q_reg ( .D(g22192), .SI(g2207), .SE(n9238), .CLK(n9425), .Q(
        g2205), .QN(n8634) );
  SDFFX1 DFF_1217_Q_reg ( .D(g22183), .SI(g2205), .SE(n9238), .CLK(n9425), .Q(
        g2209), .QN(n8995) );
  SDFFX1 DFF_1218_Q_reg ( .D(g22193), .SI(g2209), .SE(n9238), .CLK(n9425), .Q(
        g2210), .QN(n8994) );
  SDFFX1 DFF_1219_Q_reg ( .D(g22200), .SI(g2210), .SE(n9238), .CLK(n9425), .Q(
        g2208), .QN(n8633) );
  SDFFX1 DFF_1220_Q_reg ( .D(g22045), .SI(g2208), .SE(n9238), .CLK(n9425), .Q(
        g2218), .QN(n8993) );
  SDFFX1 DFF_1221_Q_reg ( .D(g22060), .SI(g2218), .SE(n9238), .CLK(n9425), .Q(
        g2219), .QN(n8992) );
  SDFFX1 DFF_1222_Q_reg ( .D(g22076), .SI(g2219), .SE(n9238), .CLK(n9425), .Q(
        g2217), .QN(n8632) );
  SDFFX1 DFF_1223_Q_reg ( .D(g22061), .SI(g2217), .SE(n9238), .CLK(n9425), .Q(
        g2221), .QN(n8991) );
  SDFFX1 DFF_1224_Q_reg ( .D(g22077), .SI(g2221), .SE(n9238), .CLK(n9425), .Q(
        g2222), .QN(n8990) );
  SDFFX1 DFF_1225_Q_reg ( .D(g22097), .SI(g2222), .SE(n9238), .CLK(n9425), .Q(
        g2220), .QN(n8631) );
  SDFFX1 DFF_1226_Q_reg ( .D(g22078), .SI(g2220), .SE(n9238), .CLK(n9425), .Q(
        g2224), .QN(n8989) );
  SDFFX1 DFF_1227_Q_reg ( .D(g22098), .SI(g2224), .SE(n9239), .CLK(n9426), .Q(
        test_so74) );
  SDFFX1 DFF_1228_Q_reg ( .D(g22115), .SI(test_si75), .SE(n9236), .CLK(n9423), 
        .Q(g2223), .QN(n8630) );
  SDFFX1 DFF_1229_Q_reg ( .D(g22099), .SI(g2223), .SE(n9236), .CLK(n9423), .Q(
        g2227) );
  SDFFX1 DFF_1230_Q_reg ( .D(g22116), .SI(g2227), .SE(n9239), .CLK(n9426), .Q(
        g2228) );
  SDFFX1 DFF_1231_Q_reg ( .D(g22138), .SI(g2228), .SE(n9239), .CLK(n9426), .Q(
        g2226) );
  SDFFX1 DFF_1232_Q_reg ( .D(g22117), .SI(g2226), .SE(n9239), .CLK(n9426), .Q(
        g2230) );
  SDFFX1 DFF_1233_Q_reg ( .D(g22139), .SI(g2230), .SE(n9239), .CLK(n9426), .Q(
        g2231) );
  SDFFX1 DFF_1234_Q_reg ( .D(g22153), .SI(g2231), .SE(n9239), .CLK(n9426), .Q(
        g2229) );
  SDFFX1 DFF_1235_Q_reg ( .D(g22140), .SI(g2229), .SE(n9239), .CLK(n9426), .Q(
        g2233), .QN(n8984) );
  SDFFX1 DFF_1236_Q_reg ( .D(g22154), .SI(g2233), .SE(n9239), .CLK(n9426), .Q(
        g2234), .QN(n8983) );
  SDFFX1 DFF_1237_Q_reg ( .D(g22171), .SI(g2234), .SE(n9239), .CLK(n9426), .Q(
        g2232), .QN(n8627) );
  SDFFX1 DFF_1238_Q_reg ( .D(g22155), .SI(g2232), .SE(n9239), .CLK(n9426), .Q(
        g2236) );
  SDFFX1 DFF_1239_Q_reg ( .D(g22172), .SI(g2236), .SE(n9239), .CLK(n9426), .Q(
        g2237) );
  SDFFX1 DFF_1240_Q_reg ( .D(g22184), .SI(g2237), .SE(n9239), .CLK(n9426), .Q(
        g2235) );
  SDFFX1 DFF_1241_Q_reg ( .D(g22173), .SI(g2235), .SE(n9234), .CLK(n9421), .Q(
        g2239) );
  SDFFX1 DFF_1242_Q_reg ( .D(g22185), .SI(g2239), .SE(n9240), .CLK(n9427), .Q(
        test_so75) );
  SDFFX1 DFF_1243_Q_reg ( .D(g22194), .SI(test_si76), .SE(n9236), .CLK(n9423), 
        .Q(g2238) );
  SDFFX1 DFF_1244_Q_reg ( .D(g25227), .SI(g2238), .SE(n9237), .CLK(n9424), .Q(
        g2245), .QN(n8696) );
  SDFFX1 DFF_1245_Q_reg ( .D(g25236), .SI(g2245), .SE(n9237), .CLK(n9424), .Q(
        g2246), .QN(n8695) );
  SDFFX1 DFF_1246_Q_reg ( .D(g25245), .SI(g2246), .SE(n9237), .CLK(n9424), .Q(
        g2244), .QN(n8694) );
  SDFFX1 DFF_1247_Q_reg ( .D(g25237), .SI(g2244), .SE(n9237), .CLK(n9424), .Q(
        g2248), .QN(n8693) );
  SDFFX1 DFF_1248_Q_reg ( .D(g25246), .SI(g2248), .SE(n9237), .CLK(n9424), .Q(
        g2249), .QN(n8692) );
  SDFFX1 DFF_1249_Q_reg ( .D(g25251), .SI(g2249), .SE(n9237), .CLK(n9424), .Q(
        g2247), .QN(n8691) );
  SDFFX1 DFF_1250_Q_reg ( .D(g25247), .SI(g2247), .SE(n9237), .CLK(n9424), .Q(
        g2251), .QN(n8690) );
  SDFFX1 DFF_1251_Q_reg ( .D(g25252), .SI(g2251), .SE(n9237), .CLK(n9424), .Q(
        g2252), .QN(n8689) );
  SDFFX1 DFF_1252_Q_reg ( .D(g25256), .SI(g2252), .SE(n9237), .CLK(n9424), .Q(
        g2250), .QN(n8688) );
  SDFFX1 DFF_1253_Q_reg ( .D(g25253), .SI(g2250), .SE(n9237), .CLK(n9424), .Q(
        g2254), .QN(n8687) );
  SDFFX1 DFF_1254_Q_reg ( .D(g25257), .SI(g2254), .SE(n9237), .CLK(n9424), .Q(
        g2255), .QN(n8686) );
  SDFFX1 DFF_1255_Q_reg ( .D(g25259), .SI(g2255), .SE(n9237), .CLK(n9424), .Q(
        g2253), .QN(n8685) );
  SDFFX1 DFF_1256_Q_reg ( .D(g30289), .SI(g2253), .SE(n9249), .CLK(n9436), .Q(
        g2261) );
  SDFFX1 DFF_1257_Q_reg ( .D(g30296), .SI(g2261), .SE(n9249), .CLK(n9436), .Q(
        test_so76) );
  SDFFX1 DFF_1258_Q_reg ( .D(g30300), .SI(test_si77), .SE(n9249), .CLK(n9436), 
        .Q(g2267) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30660), .SI(g2267), .SE(n9250), .CLK(n9437), .Q(
        g2306) );
  SDFFX1 DFF_1260_Q_reg ( .D(g30666), .SI(g2306), .SE(n9250), .CLK(n9437), .Q(
        g2309) );
  SDFFX1 DFF_1261_Q_reg ( .D(g30672), .SI(g2309), .SE(n9250), .CLK(n9437), .Q(
        g2312) );
  SDFFX1 DFF_1262_Q_reg ( .D(g30690), .SI(g2312), .SE(n9250), .CLK(n9437), .Q(
        g2270) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30693), .SI(g2270), .SE(n9250), .CLK(n9437), .Q(
        g2273) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30695), .SI(g2273), .SE(n9240), .CLK(n9427), .Q(
        g2276) );
  SDFFX1 DFF_1265_Q_reg ( .D(g30667), .SI(g2276), .SE(n9240), .CLK(n9427), .Q(
        g2315) );
  SDFFX1 DFF_1266_Q_reg ( .D(g30673), .SI(g2315), .SE(n9240), .CLK(n9427), .Q(
        g2318) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30679), .SI(g2318), .SE(n9240), .CLK(n9427), .Q(
        g2321) );
  SDFFX1 DFF_1268_Q_reg ( .D(g30301), .SI(g2321), .SE(n9240), .CLK(n9427), .Q(
        g2279) );
  SDFFX1 DFF_1269_Q_reg ( .D(g30303), .SI(g2279), .SE(n9240), .CLK(n9427), .Q(
        g2282) );
  SDFFX1 DFF_1270_Q_reg ( .D(g30304), .SI(g2282), .SE(n9240), .CLK(n9427), .Q(
        g2285) );
  SDFFX1 DFF_1271_Q_reg ( .D(g30274), .SI(g2285), .SE(n9240), .CLK(n9427), .Q(
        g2324) );
  SDFFX1 DFF_1272_Q_reg ( .D(g30282), .SI(g2324), .SE(n9240), .CLK(n9427), .Q(
        test_so77) );
  SDFFX1 DFF_1273_Q_reg ( .D(g30290), .SI(test_si78), .SE(n9240), .CLK(n9427), 
        .Q(g2330) );
  SDFFX1 DFF_1274_Q_reg ( .D(g30253), .SI(g2330), .SE(n9240), .CLK(n9427), .Q(
        g2288) );
  SDFFX1 DFF_1275_Q_reg ( .D(g30256), .SI(g2288), .SE(n9241), .CLK(n9428), .Q(
        g2291) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30260), .SI(g2291), .SE(n9241), .CLK(n9428), .Q(
        g2294) );
  SDFFX1 DFF_1277_Q_reg ( .D(g30283), .SI(g2294), .SE(n9241), .CLK(n9428), .Q(
        g2333) );
  SDFFX1 DFF_1278_Q_reg ( .D(g30291), .SI(g2333), .SE(n9241), .CLK(n9428), .Q(
        g2336) );
  SDFFX1 DFF_1279_Q_reg ( .D(g30297), .SI(g2336), .SE(n9241), .CLK(n9428), .Q(
        g2339) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30652), .SI(g2339), .SE(n9241), .CLK(n9428), .Q(
        g2297) );
  SDFFX1 DFF_1281_Q_reg ( .D(g30659), .SI(g2297), .SE(n9241), .CLK(n9428), .Q(
        g2300) );
  SDFFX1 DFF_1282_Q_reg ( .D(g30665), .SI(g2300), .SE(n9234), .CLK(n9421), .Q(
        g2303) );
  SDFFX1 DFF_1283_Q_reg ( .D(g30686), .SI(g2303), .SE(n9234), .CLK(n9421), .Q(
        g2342) );
  SDFFX1 DFF_1284_Q_reg ( .D(g30691), .SI(g2342), .SE(n9234), .CLK(n9421), .Q(
        g2345) );
  SDFFX1 DFF_1285_Q_reg ( .D(g30694), .SI(g2345), .SE(n9235), .CLK(n9422), .Q(
        g2348) );
  SDFFX1 DFF_1286_Q_reg ( .D(g25067), .SI(g2348), .SE(n9235), .CLK(n9422), .Q(
        g2160), .QN(n8809) );
  SDFFX1 DFF_1287_Q_reg ( .D(g25940), .SI(g2160), .SE(n9235), .CLK(n9422), .Q(
        test_so78) );
  SDFFX1 DFF_1288_Q_reg ( .D(g26532), .SI(test_si79), .SE(n9235), .CLK(n9422), 
        .Q(g2151), .QN(n8808) );
  SDFFX1 DFF_1289_Q_reg ( .D(g27131), .SI(g2151), .SE(n9235), .CLK(n9422), .Q(
        g2147), .QN(n9116) );
  SDFFX1 DFF_1290_Q_reg ( .D(g27621), .SI(g2147), .SE(n9235), .CLK(n9422), .Q(
        g2142), .QN(n8807) );
  SDFFX1 DFF_1291_Q_reg ( .D(g28148), .SI(g2142), .SE(n9235), .CLK(n9422), .Q(
        g2138), .QN(n9098) );
  SDFFX1 DFF_1292_Q_reg ( .D(g28637), .SI(g2138), .SE(n9235), .CLK(n9422), .Q(
        g2133), .QN(n8806) );
  SDFFX1 DFF_1293_Q_reg ( .D(g29112), .SI(g2133), .SE(n9235), .CLK(n9422), .Q(
        g2129), .QN(n9104) );
  SDFFX1 DFF_1294_Q_reg ( .D(g29357), .SI(g2129), .SE(n9235), .CLK(n9422), .Q(
        g2124), .QN(n8437) );
  SDFFX1 DFF_1295_Q_reg ( .D(g29582), .SI(g2124), .SE(n9235), .CLK(n9422), .Q(
        g2120), .QN(n8283) );
  SDFFX1 DFF_1296_Q_reg ( .D(g13110), .SI(g2120), .SE(n9235), .CLK(n9422), .Q(
        g2256) );
  SDFFX1 DFF_1297_Q_reg ( .D(g2256), .SI(g2256), .SE(n9236), .CLK(n9423), .Q(
        g5637) );
  SDFFX1 DFF_1298_Q_reg ( .D(g5637), .SI(g5637), .SE(n9236), .CLK(n9423), .Q(
        g2257), .QN(n9091) );
  SDFFX1 DFF_1299_Q_reg ( .D(g2950), .SI(g2257), .SE(n9236), .CLK(n9423), .Q(
        g5555), .QN(n4516) );
  SDFFX1 DFF_1302_Q_reg ( .D(g5637), .SI(n4606), .SE(n9236), .CLK(n9423), .Q(
        test_so79), .QN(n9121) );
  SDFFX1 DFF_1303_Q_reg ( .D(g27276), .SI(test_si80), .SE(n9249), .CLK(n9436), 
        .Q(g2429), .QN(n8764) );
  SDFFX1 DFF_1304_Q_reg ( .D(g27291), .SI(g2429), .SE(n9249), .CLK(n9436), .Q(
        g2418), .QN(n8763) );
  SDFFX1 DFF_1305_Q_reg ( .D(g27307), .SI(g2418), .SE(n9249), .CLK(n9436), .Q(
        g2421), .QN(n8762) );
  SDFFX1 DFF_1306_Q_reg ( .D(g27292), .SI(g2421), .SE(n9249), .CLK(n9436), .Q(
        g2444), .QN(n8741) );
  SDFFX1 DFF_1307_Q_reg ( .D(g27308), .SI(g2444), .SE(n9249), .CLK(n9436), .Q(
        g2433), .QN(n8740) );
  SDFFX1 DFF_1308_Q_reg ( .D(g27322), .SI(g2433), .SE(n9248), .CLK(n9435), .Q(
        g2436), .QN(n8739) );
  SDFFX1 DFF_1309_Q_reg ( .D(g27309), .SI(g2436), .SE(n9249), .CLK(n9436), .Q(
        g2459), .QN(n8486) );
  SDFFX1 DFF_1310_Q_reg ( .D(g27323), .SI(g2459), .SE(n9249), .CLK(n9436), .Q(
        g2448), .QN(n8488) );
  SDFFX1 DFF_1311_Q_reg ( .D(g27334), .SI(g2448), .SE(n9248), .CLK(n9435), .Q(
        g2451), .QN(n8487) );
  SDFFX1 DFF_1312_Q_reg ( .D(g27324), .SI(g2451), .SE(n9249), .CLK(n9436), .Q(
        g2473), .QN(n8753) );
  SDFFX1 DFF_1313_Q_reg ( .D(g27335), .SI(g2473), .SE(n9249), .CLK(n9436), .Q(
        g2463), .QN(n8752) );
  SDFFX1 DFF_1314_Q_reg ( .D(g27342), .SI(g2463), .SE(n9241), .CLK(n9428), .Q(
        g2466), .QN(n8751) );
  SDFFX1 DFF_1315_Q_reg ( .D(g28763), .SI(g2466), .SE(n9242), .CLK(n9429), .Q(
        g2483) );
  SDFFX1 DFF_1316_Q_reg ( .D(g28773), .SI(g2483), .SE(n9248), .CLK(n9435), .Q(
        g2486) );
  SDFFX1 DFF_1317_Q_reg ( .D(g28782), .SI(g2486), .SE(n9248), .CLK(n9435), .Q(
        test_so80) );
  SDFFX1 DFF_1318_Q_reg ( .D(g29213), .SI(test_si81), .SE(n9242), .CLK(n9429), 
        .Q(g2492) );
  SDFFX1 DFF_1319_Q_reg ( .D(g29221), .SI(g2492), .SE(n9242), .CLK(n9429), .Q(
        g2495) );
  SDFFX1 DFF_1320_Q_reg ( .D(g29226), .SI(g2495), .SE(n9242), .CLK(n9429), .Q(
        g2498) );
  SDFFX1 DFF_1321_Q_reg ( .D(g28774), .SI(g2498), .SE(n9245), .CLK(n9432), .Q(
        g2502), .QN(n8785) );
  SDFFX1 DFF_1322_Q_reg ( .D(g28783), .SI(g2502), .SE(n9245), .CLK(n9432), .Q(
        g2503), .QN(n8775) );
  SDFFX1 DFF_1323_Q_reg ( .D(g28788), .SI(g2503), .SE(n9245), .CLK(n9432), .Q(
        g2501), .QN(n8784) );
  SDFFX1 DFF_1324_Q_reg ( .D(g26817), .SI(g2501), .SE(n9245), .CLK(n9432), .Q(
        g2504) );
  SDFFX1 DFF_1325_Q_reg ( .D(g26822), .SI(g2504), .SE(n9245), .CLK(n9432), .Q(
        g2507) );
  SDFFX1 DFF_1326_Q_reg ( .D(g26825), .SI(g2507), .SE(n9245), .CLK(n9432), .Q(
        g2510) );
  SDFFX1 DFF_1327_Q_reg ( .D(g26823), .SI(g2510), .SE(n9246), .CLK(n9433), .Q(
        g2513) );
  SDFFX1 DFF_1328_Q_reg ( .D(g26826), .SI(g2513), .SE(n9246), .CLK(n9433), .Q(
        g2516) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26827), .SI(g2516), .SE(n9246), .CLK(n9433), .Q(
        g2519) );
  SDFFX1 DFF_1330_Q_reg ( .D(g27767), .SI(g2519), .SE(n9246), .CLK(n9433), .Q(
        g2523), .QN(n8783) );
  SDFFX1 DFF_1331_Q_reg ( .D(g27769), .SI(g2523), .SE(n9246), .CLK(n9433), .Q(
        g2524), .QN(n8774) );
  SDFFX1 DFF_1332_Q_reg ( .D(g27771), .SI(g2524), .SE(n9246), .CLK(n9433), .Q(
        test_so81) );
  SDFFX1 DFF_1333_Q_reg ( .D(g29618), .SI(test_si82), .SE(n9241), .CLK(n9428), 
        .Q(g2387), .QN(n8388) );
  SDFFX1 DFF_1334_Q_reg ( .D(g29621), .SI(g2387), .SE(n9241), .CLK(n9428), .Q(
        g2388), .QN(n8376) );
  SDFFX1 DFF_1335_Q_reg ( .D(g29623), .SI(g2388), .SE(n9241), .CLK(n9428), .Q(
        g2389), .QN(n8387) );
  SDFFX1 DFF_1336_Q_reg ( .D(g30707), .SI(g2389), .SE(n9241), .CLK(n9428), .Q(
        g2390), .QN(n8386) );
  SDFFX1 DFF_1337_Q_reg ( .D(g30709), .SI(g2390), .SE(n9234), .CLK(n9421), .Q(
        g2391), .QN(n8375) );
  SDFFX1 DFF_1338_Q_reg ( .D(g30566), .SI(g2391), .SE(n9236), .CLK(n9423), .Q(
        g2392), .QN(n8385) );
  SDFFX1 DFF_1339_Q_reg ( .D(g30505), .SI(g2392), .SE(n9234), .CLK(n9421), .Q(
        g2393), .QN(n8384) );
  SDFFX1 DFF_1340_Q_reg ( .D(g30341), .SI(g2393), .SE(n9236), .CLK(n9423), .Q(
        g2394), .QN(n8374) );
  SDFFX1 DFF_1341_Q_reg ( .D(g30356), .SI(g2394), .SE(n9236), .CLK(n9423), .Q(
        g2395), .QN(n8383) );
  SDFFX1 DFF_1342_Q_reg ( .D(g29182), .SI(g2395), .SE(n9250), .CLK(n9437), .Q(
        g2397) );
  SDFFX1 DFF_1343_Q_reg ( .D(g29185), .SI(g2397), .SE(n9250), .CLK(n9437), .Q(
        g2398) );
  SDFFX1 DFF_1344_Q_reg ( .D(g29187), .SI(g2398), .SE(n9250), .CLK(n9437), .Q(
        g2396) );
  SDFFX1 DFF_1345_Q_reg ( .D(g26672), .SI(g2396), .SE(n9250), .CLK(n9437), .Q(
        g2478), .QN(n8782) );
  SDFFX1 DFF_1346_Q_reg ( .D(g26676), .SI(g2478), .SE(n9250), .CLK(n9437), .Q(
        g2479), .QN(n8773) );
  SDFFX1 DFF_1347_Q_reg ( .D(g26025), .SI(g2479), .SE(n9250), .CLK(n9437), .Q(
        test_so82) );
  SDFFX1 DFF_1348_Q_reg ( .D(n4287), .SI(test_si83), .SE(n9143), .CLK(n9330), 
        .Q(g2525) );
  SDFFX1 DFF_1349_Q_reg ( .D(g2525), .SI(g2525), .SE(n9143), .CLK(n9330), .Q(
        n7946), .QN(DFF_1349_n1) );
  SDFFX1 DFF_1350_Q_reg ( .D(n4563), .SI(n7946), .SE(n9143), .CLK(n9330), .Q(
        g2527) );
  SDFFX1 DFF_1351_Q_reg ( .D(g2527), .SI(g2527), .SE(n9143), .CLK(n9330), .Q(
        n7945), .QN(DFF_1351_n1) );
  SDFFX1 DFF_1352_Q_reg ( .D(n4555), .SI(n7945), .SE(n9143), .CLK(n9330), .Q(
        g2529) );
  SDFFX1 DFF_1353_Q_reg ( .D(g2529), .SI(g2529), .SE(n9143), .CLK(n9330), .Q(
        n7944), .QN(DFF_1353_n1) );
  SDFFX1 DFF_1354_Q_reg ( .D(n4325), .SI(n7944), .SE(n9143), .CLK(n9330), .Q(
        g2355) );
  SDFFX1 DFF_1355_Q_reg ( .D(g2355), .SI(g2355), .SE(n9143), .CLK(n9330), .Q(
        n7943), .QN(DFF_1355_n1) );
  SDFFX1 DFF_1356_Q_reg ( .D(n4389), .SI(n7943), .SE(n9144), .CLK(n9331), .Q(
        g2357) );
  SDFFX1 DFF_1357_Q_reg ( .D(g2357), .SI(g2357), .SE(n9144), .CLK(n9331), .Q(
        n7942), .QN(DFF_1357_n1) );
  SDFFX1 DFF_1358_Q_reg ( .D(n4319), .SI(n7942), .SE(n9144), .CLK(n9331), .Q(
        g2359) );
  SDFFX1 DFF_1359_Q_reg ( .D(g2359), .SI(g2359), .SE(n9144), .CLK(n9331), .Q(
        n7941), .QN(DFF_1359_n1) );
  SDFFX1 DFF_1360_Q_reg ( .D(n4373), .SI(n7941), .SE(n9144), .CLK(n9331), .Q(
        g2361) );
  SDFFX1 DFF_1361_Q_reg ( .D(g2361), .SI(g2361), .SE(n9144), .CLK(n9331), .Q(
        n7940), .QN(DFF_1361_n1) );
  SDFFX1 DFF_1362_Q_reg ( .D(n4377), .SI(n7940), .SE(n9144), .CLK(n9331), .Q(
        test_so83) );
  SDFFX1 DFF_1363_Q_reg ( .D(test_so83), .SI(test_si84), .SE(n9144), .CLK(
        n9331), .Q(n7938), .QN(DFF_1363_n1) );
  SDFFX1 DFF_1364_Q_reg ( .D(g2878), .SI(n7938), .SE(n9149), .CLK(n9336), .Q(
        g2365) );
  SDFFX1 DFF_1365_Q_reg ( .D(g2365), .SI(g2365), .SE(n9149), .CLK(n9336), .Q(
        n7937), .QN(n4483) );
  SDFFX1 DFF_1366_Q_reg ( .D(n4285), .SI(n7937), .SE(n9248), .CLK(n9435), .Q(
        g2374), .QN(n4487) );
  SDFFX1 DFF_1367_Q_reg ( .D(g30055), .SI(g2374), .SE(n9253), .CLK(n9440), .Q(
        g2380) );
  SDFFX1 DFF_1378_Q_reg ( .D(n4275), .SI(g2380), .SE(n9250), .CLK(n9437), .Q(
        n7936), .QN(DFF_1378_n1) );
  SDFFX1 DFF_1379_Q_reg ( .D(g2429), .SI(n7936), .SE(n9251), .CLK(n9438), .Q(
        g2417) );
  SDFFX1 DFF_1380_Q_reg ( .D(g2417), .SI(g2417), .SE(n9251), .CLK(n9438), .Q(
        g2424) );
  SDFFX1 DFF_1381_Q_reg ( .D(g2418), .SI(g2424), .SE(n9251), .CLK(n9438), .Q(
        g2425) );
  SDFFX1 DFF_1382_Q_reg ( .D(g2425), .SI(g2425), .SE(n9251), .CLK(n9438), .Q(
        g2426) );
  SDFFX1 DFF_1383_Q_reg ( .D(g2421), .SI(g2426), .SE(n9251), .CLK(n9438), .Q(
        g2427) );
  SDFFX1 DFF_1384_Q_reg ( .D(g2427), .SI(g2427), .SE(n9251), .CLK(n9438), .Q(
        g2428) );
  SDFFX1 DFF_1385_Q_reg ( .D(g2444), .SI(g2428), .SE(n9251), .CLK(n9438), .Q(
        g2432) );
  SDFFX1 DFF_1386_Q_reg ( .D(g2432), .SI(g2432), .SE(n9251), .CLK(n9438), .Q(
        g2439) );
  SDFFX1 DFF_1387_Q_reg ( .D(g2433), .SI(g2439), .SE(n9251), .CLK(n9438), .Q(
        test_so84) );
  SDFFX1 DFF_1388_Q_reg ( .D(test_so84), .SI(test_si85), .SE(n9251), .CLK(
        n9438), .Q(g2441) );
  SDFFX1 DFF_1389_Q_reg ( .D(g2436), .SI(g2441), .SE(n9251), .CLK(n9438), .Q(
        g2442) );
  SDFFX1 DFF_1390_Q_reg ( .D(g2442), .SI(g2442), .SE(n9251), .CLK(n9438), .Q(
        g2443) );
  SDFFX1 DFF_1391_Q_reg ( .D(g2459), .SI(g2443), .SE(n9252), .CLK(n9439), .Q(
        g2447) );
  SDFFX1 DFF_1392_Q_reg ( .D(g2447), .SI(g2447), .SE(n9252), .CLK(n9439), .Q(
        g2454) );
  SDFFX1 DFF_1393_Q_reg ( .D(g2448), .SI(g2454), .SE(n9252), .CLK(n9439), .Q(
        g2455) );
  SDFFX1 DFF_1394_Q_reg ( .D(g2455), .SI(g2455), .SE(n9252), .CLK(n9439), .Q(
        g2456) );
  SDFFX1 DFF_1395_Q_reg ( .D(g2451), .SI(g2456), .SE(n9252), .CLK(n9439), .Q(
        g2457) );
  SDFFX1 DFF_1396_Q_reg ( .D(g2457), .SI(g2457), .SE(n9252), .CLK(n9439), .Q(
        g2458) );
  SDFFX1 DFF_1397_Q_reg ( .D(g2473), .SI(g2458), .SE(n9252), .CLK(n9439), .Q(
        g2462) );
  SDFFX1 DFF_1398_Q_reg ( .D(g2462), .SI(g2462), .SE(n9252), .CLK(n9439), .Q(
        g2469) );
  SDFFX1 DFF_1399_Q_reg ( .D(g2463), .SI(g2469), .SE(n9252), .CLK(n9439), .Q(
        g2470) );
  SDFFX1 DFF_1400_Q_reg ( .D(g2470), .SI(g2470), .SE(n9252), .CLK(n9439), .Q(
        g2471) );
  SDFFX1 DFF_1401_Q_reg ( .D(g2466), .SI(g2471), .SE(n9252), .CLK(n9439), .Q(
        g2472) );
  SDFFX1 DFF_1402_Q_reg ( .D(g2472), .SI(g2472), .SE(n9252), .CLK(n9439), .Q(
        test_so85) );
  SDFFX1 DFF_1403_Q_reg ( .D(n4598), .SI(test_si86), .SE(n9129), .CLK(n9316), 
        .Q(g5747) );
  SDFFX1 DFF_1404_Q_reg ( .D(g5747), .SI(g5747), .SE(n9129), .CLK(n9316), .Q(
        g5796) );
  SDFFX1 DFF_1405_Q_reg ( .D(g5796), .SI(g5796), .SE(n9129), .CLK(n9316), .Q(
        g2412) );
  SDFFX1 DFF_1406_Q_reg ( .D(n4598), .SI(g2412), .SE(n9129), .CLK(n9316), .Q(
        g7302), .QN(n4314) );
  SDFFX1 DFF_1407_Q_reg ( .D(g7302), .SI(g7302), .SE(n9129), .CLK(n9316), .Q(
        g7390), .QN(n4370) );
  SDFFX1 DFF_1408_Q_reg ( .D(g7390), .SI(g7390), .SE(n9129), .CLK(n9316), .Q(
        g2624), .QN(n4299) );
  SDFFX1 DFF_1409_Q_reg ( .D(g21847), .SI(g2624), .SE(n9152), .CLK(n9339), .Q(
        g2628), .QN(n9050) );
  SDFFX1 DFF_1410_Q_reg ( .D(g18780), .SI(g2628), .SE(n9152), .CLK(n9339), .Q(
        g2631), .QN(n4352) );
  SDFFX1 DFF_1411_Q_reg ( .D(g18820), .SI(g2631), .SE(n9152), .CLK(n9339), .Q(
        g2584), .QN(n4303) );
  SDFFX1 DFF_1412_Q_reg ( .D(n1386), .SI(g2584), .SE(n9244), .CLK(n9431), .Q(
        g2587) );
  SDFFX1 DFF_1413_Q_reg ( .D(g2587), .SI(g2587), .SE(n9244), .CLK(n9431), .Q(
        g2597) );
  SDFFX1 DFF_1414_Q_reg ( .D(g2597), .SI(g2597), .SE(n9244), .CLK(n9431), .Q(
        g2598) );
  SDFFX1 DFF_1415_Q_reg ( .D(g2530), .SI(g2598), .SE(n9244), .CLK(n9431), .Q(
        g2638) );
  SDFFX1 DFF_1416_Q_reg ( .D(g2638), .SI(g2638), .SE(n9244), .CLK(n9431), .Q(
        g2643) );
  SDFFX1 DFF_1417_Q_reg ( .D(g2533), .SI(g2643), .SE(n9244), .CLK(n9431), .Q(
        test_so86) );
  SDFFX1 DFF_1418_Q_reg ( .D(test_so86), .SI(test_si87), .SE(n9244), .CLK(
        n9431), .Q(g2645) );
  SDFFX1 DFF_1419_Q_reg ( .D(g2536), .SI(g2645), .SE(n9244), .CLK(n9431), .Q(
        g2646) );
  SDFFX1 DFF_1420_Q_reg ( .D(g2646), .SI(g2646), .SE(n9244), .CLK(n9431), .Q(
        g2647) );
  SDFFX1 DFF_1421_Q_reg ( .D(g2540), .SI(g2647), .SE(n9242), .CLK(n9429), .Q(
        g2648) );
  SDFFX1 DFF_1422_Q_reg ( .D(g2648), .SI(g2648), .SE(n9242), .CLK(n9429), .Q(
        g2639) );
  SDFFX1 DFF_1423_Q_reg ( .D(g2543), .SI(g2639), .SE(n9242), .CLK(n9429), .Q(
        g2640) );
  SDFFX1 DFF_1424_Q_reg ( .D(g2640), .SI(g2640), .SE(n9242), .CLK(n9429), .Q(
        g2641) );
  SDFFX1 DFF_1425_Q_reg ( .D(g2546), .SI(g2641), .SE(n9243), .CLK(n9430), .Q(
        g2642) );
  SDFFX1 DFF_1426_Q_reg ( .D(g2642), .SI(g2642), .SE(n9243), .CLK(n9430), .Q(
        g2564) );
  SDFFX1 DFF_1427_Q_reg ( .D(g2950), .SI(g2564), .SE(n9243), .CLK(n9430), .Q(
        g8087), .QN(n4456) );
  SDFFX1 DFF_1428_Q_reg ( .D(g8087), .SI(g8087), .SE(n9243), .CLK(n9430), .Q(
        g8167), .QN(n4455) );
  SDFFX1 DFF_1429_Q_reg ( .D(g8167), .SI(g8167), .SE(n9243), .CLK(n9430), .Q(
        g2560), .QN(n4463) );
  SDFFX1 DFF_1430_Q_reg ( .D(g23114), .SI(g2560), .SE(n9246), .CLK(n9433), .Q(
        g2561) );
  SDFFX1 DFF_1431_Q_reg ( .D(g23133), .SI(g2561), .SE(n9246), .CLK(n9433), .Q(
        g2562) );
  SDFFX1 DFF_1432_Q_reg ( .D(g21970), .SI(g2562), .SE(n9246), .CLK(n9433), .Q(
        test_so87) );
  SDFFX1 DFF_1433_Q_reg ( .D(g23407), .SI(test_si88), .SE(n9243), .CLK(n9430), 
        .Q(g2530) );
  SDFFX1 DFF_1434_Q_reg ( .D(g23418), .SI(g2530), .SE(n9243), .CLK(n9430), .Q(
        g2533) );
  SDFFX1 DFF_1435_Q_reg ( .D(g24209), .SI(g2533), .SE(n9244), .CLK(n9431), .Q(
        g2536) );
  SDFFX1 DFF_1436_Q_reg ( .D(g24214), .SI(g2536), .SE(n9244), .CLK(n9431), .Q(
        g2552) );
  SDFFX1 DFF_1437_Q_reg ( .D(g24226), .SI(g2552), .SE(n9244), .CLK(n9431), .Q(
        g2553) );
  SDFFX1 DFF_1438_Q_reg ( .D(g24238), .SI(g2553), .SE(n9245), .CLK(n9432), .Q(
        g2554) );
  SDFFX1 DFF_1439_Q_reg ( .D(g23132), .SI(g2554), .SE(n9242), .CLK(n9429), .Q(
        g2555) );
  SDFFX1 DFF_1440_Q_reg ( .D(g23047), .SI(g2555), .SE(n9242), .CLK(n9429), .Q(
        g2559) );
  SDFFX1 DFF_1441_Q_reg ( .D(g23076), .SI(g2559), .SE(n9242), .CLK(n9429), .Q(
        g2539) );
  SDFFX1 DFF_1442_Q_reg ( .D(g24225), .SI(g2539), .SE(n9242), .CLK(n9429), .Q(
        g2540) );
  SDFFX1 DFF_1443_Q_reg ( .D(g24237), .SI(g2540), .SE(n9243), .CLK(n9430), .Q(
        g2543) );
  SDFFX1 DFF_1444_Q_reg ( .D(g24250), .SI(g2543), .SE(n9243), .CLK(n9430), .Q(
        g2546) );
  SDFFX1 DFF_1445_Q_reg ( .D(n1359), .SI(g2546), .SE(n9243), .CLK(n9430), .Q(
        g2602) );
  SDFFX1 DFF_1446_Q_reg ( .D(g2602), .SI(g2602), .SE(n9243), .CLK(n9430), .Q(
        g2609) );
  SDFFX1 DFF_1447_Q_reg ( .D(g2609), .SI(g2609), .SE(n9243), .CLK(n9430), .Q(
        test_so88) );
  SDFFX1 DFF_1448_Q_reg ( .D(g13175), .SI(test_si89), .SE(n9245), .CLK(n9432), 
        .Q(g2617) );
  SDFFX1 DFF_1449_Q_reg ( .D(g2617), .SI(g2617), .SE(n9245), .CLK(n9432), .Q(
        n7930) );
  SDFFX1 DFF_1450_Q_reg ( .D(g30072), .SI(n7930), .SE(n9245), .CLK(n9432), .Q(
        n7929) );
  SDFFX1 DFF_1451_Q_reg ( .D(g13143), .SI(n7929), .SE(n9245), .CLK(n9432), .Q(
        g2623) );
  SDFFX1 DFF_1452_Q_reg ( .D(g2623), .SI(g2623), .SE(n9245), .CLK(n9432), .Q(
        g2574), .QN(n4543) );
  SDFFX1 DFF_1453_Q_reg ( .D(g13194), .SI(g2574), .SE(n9246), .CLK(n9433), .Q(
        g2632) );
  SDFFX1 DFF_1454_Q_reg ( .D(g2632), .SI(g2632), .SE(n9246), .CLK(n9433), .Q(
        g2633) );
  SDFFX1 DFF_1455_Q_reg ( .D(g27310), .SI(g2633), .SE(n9246), .CLK(n9433), .Q(
        g2650), .QN(n8441) );
  SDFFX1 DFF_1456_Q_reg ( .D(g27325), .SI(g2650), .SE(n9248), .CLK(n9435), .Q(
        g2651), .QN(n8443) );
  SDFFX1 DFF_1457_Q_reg ( .D(g27336), .SI(g2651), .SE(n9248), .CLK(n9435), .Q(
        g2649), .QN(n8442) );
  SDFFX1 DFF_1458_Q_reg ( .D(g27326), .SI(g2649), .SE(n9248), .CLK(n9435), .Q(
        g2653), .QN(n8453) );
  SDFFX1 DFF_1459_Q_reg ( .D(g27337), .SI(g2653), .SE(n9248), .CLK(n9435), .Q(
        g2654), .QN(n8455) );
  SDFFX1 DFF_1460_Q_reg ( .D(g27343), .SI(g2654), .SE(n9248), .CLK(n9435), .Q(
        g2652), .QN(n8454) );
  SDFFX1 DFF_1461_Q_reg ( .D(g27338), .SI(g2652), .SE(n9248), .CLK(n9435), .Q(
        g2656), .QN(n8287) );
  SDFFX1 DFF_1462_Q_reg ( .D(g27344), .SI(g2656), .SE(n9248), .CLK(n9435), .Q(
        test_so89) );
  SDFFX1 DFF_1463_Q_reg ( .D(g27347), .SI(test_si90), .SE(n9247), .CLK(n9434), 
        .Q(g2655), .QN(n8288) );
  SDFFX1 DFF_1464_Q_reg ( .D(g27345), .SI(g2655), .SE(n9247), .CLK(n9434), .Q(
        g2659), .QN(n8464) );
  SDFFX1 DFF_1465_Q_reg ( .D(g27348), .SI(g2659), .SE(n9247), .CLK(n9434), .Q(
        g2660), .QN(n8466) );
  SDFFX1 DFF_1466_Q_reg ( .D(g27354), .SI(g2660), .SE(n9247), .CLK(n9434), .Q(
        g2658), .QN(n8465) );
  SDFFX1 DFF_1467_Q_reg ( .D(g24527), .SI(g2658), .SE(n9247), .CLK(n9434), .Q(
        g2661) );
  SDFFX1 DFF_1468_Q_reg ( .D(g24537), .SI(g2661), .SE(n9247), .CLK(n9434), .Q(
        g2664) );
  SDFFX1 DFF_1469_Q_reg ( .D(g24547), .SI(g2664), .SE(n9247), .CLK(n9434), .Q(
        g2667) );
  SDFFX1 DFF_1470_Q_reg ( .D(g24538), .SI(g2667), .SE(n9247), .CLK(n9434), .Q(
        g2670) );
  SDFFX1 DFF_1471_Q_reg ( .D(g24548), .SI(g2670), .SE(n9247), .CLK(n9434), .Q(
        g2673) );
  SDFFX1 DFF_1472_Q_reg ( .D(g24557), .SI(g2673), .SE(n9247), .CLK(n9434), .Q(
        g2676) );
  SDFFX1 DFF_1473_Q_reg ( .D(g28364), .SI(g2676), .SE(n9247), .CLK(n9434), .Q(
        g2688) );
  SDFFX1 DFF_1474_Q_reg ( .D(g28368), .SI(g2688), .SE(n9247), .CLK(n9434), .Q(
        g2691) );
  SDFFX1 DFF_1475_Q_reg ( .D(g28371), .SI(g2691), .SE(n9153), .CLK(n9340), .Q(
        g2694) );
  SDFFX1 DFF_1476_Q_reg ( .D(g28358), .SI(g2694), .SE(n9253), .CLK(n9440), .Q(
        g2679) );
  SDFFX1 DFF_1477_Q_reg ( .D(g28363), .SI(g2679), .SE(n9253), .CLK(n9440), .Q(
        test_so90) );
  SDFFX1 DFF_1478_Q_reg ( .D(g28367), .SI(test_si91), .SE(n9253), .CLK(n9440), 
        .Q(g2685) );
  SDFFX1 DFF_1479_Q_reg ( .D(g26575), .SI(g2685), .SE(n9253), .CLK(n9440), .Q(
        g2565) );
  SDFFX1 DFF_1480_Q_reg ( .D(g26596), .SI(g2565), .SE(n9253), .CLK(n9440), .Q(
        g2568) );
  SDFFX1 DFF_1481_Q_reg ( .D(g26616), .SI(g2568), .SE(n9253), .CLK(n9440), .Q(
        g2571) );
  SDFFX1 DFF_1482_Q_reg ( .D(g2574), .SI(g2571), .SE(n9253), .CLK(n9440), .Q(
        g2580), .QN(n8602) );
  SDFFX1 DFF_1483_Q_reg ( .D(g22687), .SI(g2580), .SE(n9153), .CLK(n9340), .Q(
        n7926) );
  SDFFX1 DFF_1492_Q_reg ( .D(g30061), .SI(n7926), .SE(n9153), .CLK(n9340), .Q(
        g16437) );
  SDFFX1 DFF_1493_Q_reg ( .D(g16437), .SI(g16437), .SE(n9154), .CLK(n9341), 
        .Q(g2599), .QN(n8825) );
  SDFFX1 DFF_1494_Q_reg ( .D(DFF_1349_n1), .SI(g2599), .SE(n9154), .CLK(n9341), 
        .Q(n7925) );
  SDFFX1 DFF_1495_Q_reg ( .D(DFF_1351_n1), .SI(n7925), .SE(n9154), .CLK(n9341), 
        .Q(n7924) );
  SDFFX1 DFF_1496_Q_reg ( .D(DFF_1353_n1), .SI(n7924), .SE(n9154), .CLK(n9341), 
        .Q(n7923) );
  SDFFX1 DFF_1497_Q_reg ( .D(DFF_1355_n1), .SI(n7923), .SE(n9154), .CLK(n9341), 
        .Q(n7922) );
  SDFFX1 DFF_1498_Q_reg ( .D(DFF_1357_n1), .SI(n7922), .SE(n9154), .CLK(n9341), 
        .Q(n7921) );
  SDFFX1 DFF_1499_Q_reg ( .D(DFF_1359_n1), .SI(n7921), .SE(n9154), .CLK(n9341), 
        .Q(n7920) );
  SDFFX1 DFF_1500_Q_reg ( .D(DFF_1361_n1), .SI(n7920), .SE(n9154), .CLK(n9341), 
        .Q(test_so91) );
  SDFFX1 DFF_1501_Q_reg ( .D(DFF_1363_n1), .SI(test_si92), .SE(n9144), .CLK(
        n9331), .Q(g2611) );
  SDFFX1 DFF_1502_Q_reg ( .D(g24092), .SI(g2611), .SE(n9254), .CLK(n9441), .Q(
        g2612), .QN(n4490) );
  SDFFX1 DFF_1503_Q_reg ( .D(n4483), .SI(g2612), .SE(n9149), .CLK(n9336), .Q(
        n7918) );
  SDFFX1 DFF_1505_Q_reg ( .D(g7425), .SI(g7425), .SE(n9150), .CLK(n9337), .Q(
        g7487), .QN(n4356) );
  SDFFX1 DFF_1506_Q_reg ( .D(g7487), .SI(g7487), .SE(n9150), .CLK(n9337), .Q(
        g2703), .QN(n4292) );
  SDFFX1 DFF_1507_Q_reg ( .D(g16718), .SI(g2703), .SE(n9152), .CLK(n9339), .Q(
        g2704), .QN(n9085) );
  SDFFX1 DFF_1508_Q_reg ( .D(g20375), .SI(g2704), .SE(n9152), .CLK(n9339), .Q(
        g2733) );
  SDFFX1 DFF_1509_Q_reg ( .D(g20789), .SI(g2733), .SE(n9152), .CLK(n9339), .Q(
        g2714), .QN(n4398) );
  SDFFX1 DFF_1510_Q_reg ( .D(g21974), .SI(g2714), .SE(n9152), .CLK(n9339), .Q(
        g2707), .QN(n4472) );
  SDFFX1 DFF_1511_Q_reg ( .D(g23348), .SI(g2707), .SE(n9152), .CLK(n9339), .Q(
        g2727), .QN(n4419) );
  SDFFX1 DFF_1512_Q_reg ( .D(g24438), .SI(g2727), .SE(n9152), .CLK(n9339), .Q(
        g2720), .QN(n4408) );
  SDFFX1 DFF_1513_Q_reg ( .D(g25197), .SI(g2720), .SE(n9153), .CLK(n9340), .Q(
        g2734), .QN(n4397) );
  SDFFX1 DFF_1514_Q_reg ( .D(g26677), .SI(g2734), .SE(n9153), .CLK(n9340), .Q(
        g2746), .QN(n4407) );
  SDFFX1 DFF_1515_Q_reg ( .D(g26795), .SI(g2746), .SE(n9153), .CLK(n9340), .Q(
        test_so92), .QN(n9122) );
  SDFFX1 DFF_1516_Q_reg ( .D(g27243), .SI(test_si93), .SE(n9153), .CLK(n9340), 
        .Q(g2753), .QN(n4471) );
  SDFFX1 DFF_1517_Q_reg ( .D(g27724), .SI(g2753), .SE(n9153), .CLK(n9340), .Q(
        g2760), .QN(n4393) );
  SDFFX1 DFF_1518_Q_reg ( .D(g28328), .SI(g2760), .SE(n9153), .CLK(n9340), .Q(
        g2766), .QN(n4415) );
  SDFFX1 DFF_1519_Q_reg ( .D(g20918), .SI(g2766), .SE(n9153), .CLK(n9340), .Q(
        g2773), .QN(n8886) );
  SDFFX1 DFF_1520_Q_reg ( .D(g20939), .SI(g2773), .SE(n9154), .CLK(n9341), .Q(
        g2774), .QN(n8885) );
  SDFFX1 DFF_1521_Q_reg ( .D(g20962), .SI(g2774), .SE(n9154), .CLK(n9341), .Q(
        g2772), .QN(n8948) );
  SDFFX1 DFF_1522_Q_reg ( .D(g20940), .SI(g2772), .SE(n9155), .CLK(n9342), .Q(
        g2776), .QN(n8884) );
  SDFFX1 DFF_1523_Q_reg ( .D(g20963), .SI(g2776), .SE(n9155), .CLK(n9342), .Q(
        g2777), .QN(n8883) );
  SDFFX1 DFF_1524_Q_reg ( .D(g20981), .SI(g2777), .SE(n9155), .CLK(n9342), .Q(
        g2775), .QN(n8947) );
  SDFFX1 DFF_1525_Q_reg ( .D(g20964), .SI(g2775), .SE(n9155), .CLK(n9342), .Q(
        g2779), .QN(n8882) );
  SDFFX1 DFF_1526_Q_reg ( .D(g20982), .SI(g2779), .SE(n9155), .CLK(n9342), .Q(
        g2780), .QN(n8881) );
  SDFFX1 DFF_1527_Q_reg ( .D(g21004), .SI(g2780), .SE(n9155), .CLK(n9342), .Q(
        g2778), .QN(n8946) );
  SDFFX1 DFF_1528_Q_reg ( .D(g20983), .SI(g2778), .SE(n9155), .CLK(n9342), .Q(
        g2782), .QN(n8880) );
  SDFFX1 DFF_1529_Q_reg ( .D(g21005), .SI(g2782), .SE(n9155), .CLK(n9342), .Q(
        g2783), .QN(n8879) );
  SDFFX1 DFF_1530_Q_reg ( .D(g21025), .SI(g2783), .SE(n9157), .CLK(n9344), .Q(
        test_so93) );
  SDFFX1 DFF_1531_Q_reg ( .D(g21006), .SI(test_si94), .SE(n9153), .CLK(n9340), 
        .Q(g2785), .QN(n8878) );
  SDFFX1 DFF_1532_Q_reg ( .D(g21026), .SI(g2785), .SE(n9154), .CLK(n9341), .Q(
        g2786), .QN(n8877) );
  SDFFX1 DFF_1533_Q_reg ( .D(g21043), .SI(g2786), .SE(n9156), .CLK(n9343), .Q(
        g2784), .QN(n8945) );
  SDFFX1 DFF_1534_Q_reg ( .D(g21027), .SI(g2784), .SE(n9156), .CLK(n9343), .Q(
        g2788), .QN(n8876) );
  SDFFX1 DFF_1535_Q_reg ( .D(g21044), .SI(g2788), .SE(n9156), .CLK(n9343), .Q(
        g2789), .QN(n8875) );
  SDFFX1 DFF_1536_Q_reg ( .D(g21060), .SI(g2789), .SE(n9156), .CLK(n9343), .Q(
        g2787), .QN(n8944) );
  SDFFX1 DFF_1537_Q_reg ( .D(g21045), .SI(g2787), .SE(n9156), .CLK(n9343), .Q(
        g2791), .QN(n8874) );
  SDFFX1 DFF_1538_Q_reg ( .D(g21061), .SI(g2791), .SE(n9156), .CLK(n9343), .Q(
        g2792), .QN(n8873) );
  SDFFX1 DFF_1539_Q_reg ( .D(g21073), .SI(g2792), .SE(n9156), .CLK(n9343), .Q(
        g2790), .QN(n8943) );
  SDFFX1 DFF_1540_Q_reg ( .D(g21062), .SI(g2790), .SE(n9156), .CLK(n9343), .Q(
        g2794), .QN(n8872) );
  SDFFX1 DFF_1541_Q_reg ( .D(g21074), .SI(g2794), .SE(n9156), .CLK(n9343), .Q(
        g2795), .QN(n8871) );
  SDFFX1 DFF_1542_Q_reg ( .D(g21081), .SI(g2795), .SE(n9156), .CLK(n9343), .Q(
        g2793), .QN(n8942) );
  SDFFX1 DFF_1543_Q_reg ( .D(g21075), .SI(g2793), .SE(n9156), .CLK(n9343), .Q(
        g2797), .QN(n8870) );
  SDFFX1 DFF_1544_Q_reg ( .D(g21082), .SI(g2797), .SE(n9156), .CLK(n9343), .Q(
        g2798), .QN(n8869) );
  SDFFX1 DFF_1545_Q_reg ( .D(g21094), .SI(g2798), .SE(n9157), .CLK(n9344), .Q(
        test_so94) );
  SDFFX1 DFF_1546_Q_reg ( .D(g20919), .SI(test_si95), .SE(n9153), .CLK(n9340), 
        .Q(g2800), .QN(n8868) );
  SDFFX1 DFF_1547_Q_reg ( .D(g20941), .SI(g2800), .SE(n9154), .CLK(n9341), .Q(
        g2801), .QN(n8867) );
  SDFFX1 DFF_1548_Q_reg ( .D(g20965), .SI(g2801), .SE(n9155), .CLK(n9342), .Q(
        g2799), .QN(n8941) );
  SDFFX1 DFF_1549_Q_reg ( .D(g21007), .SI(g2799), .SE(n9155), .CLK(n9342), .Q(
        g2803), .QN(n8678) );
  SDFFX1 DFF_1550_Q_reg ( .D(g21028), .SI(g2803), .SE(n9155), .CLK(n9342), .Q(
        g2804), .QN(n8670) );
  SDFFX1 DFF_1551_Q_reg ( .D(g21046), .SI(g2804), .SE(n9155), .CLK(n9342), .Q(
        g2802), .QN(n8733) );
  SDFFX1 DFF_1552_Q_reg ( .D(g21029), .SI(g2802), .SE(n9253), .CLK(n9440), .Q(
        g2806), .QN(n8677) );
  SDFFX1 DFF_1553_Q_reg ( .D(g21047), .SI(g2806), .SE(n9253), .CLK(n9440), .Q(
        g2807), .QN(n8669) );
  SDFFX1 DFF_1554_Q_reg ( .D(g21063), .SI(g2807), .SE(n9253), .CLK(n9440), .Q(
        g2805), .QN(n8732) );
  SDFFX1 DFF_1555_Q_reg ( .D(g25272), .SI(g2805), .SE(n9150), .CLK(n9337), .Q(
        g2809) );
  SDFFX1 DFF_1556_Q_reg ( .D(g25280), .SI(g2809), .SE(n9253), .CLK(n9440), .Q(
        g2810) );
  SDFFX1 DFF_1557_Q_reg ( .D(g25288), .SI(g2810), .SE(n9157), .CLK(n9344), .Q(
        g2808) );
  SDFFX1 DFF_1558_Q_reg ( .D(g22269), .SI(g2808), .SE(n9157), .CLK(n9344), .Q(
        g2812) );
  SDFFX1 DFF_1559_Q_reg ( .D(g22284), .SI(g2812), .SE(n9157), .CLK(n9344), .Q(
        g2813) );
  SDFFX1 DFF_1560_Q_reg ( .D(g22299), .SI(g2813), .SE(n9157), .CLK(n9344), .Q(
        test_so95) );
  SDFFX1 DFF_1561_Q_reg ( .D(g20877), .SI(test_si96), .SE(n9129), .CLK(n9316), 
        .Q(n7913) );
  SDFFX1 DFF_1562_Q_reg ( .D(g20884), .SI(n7913), .SE(n9129), .CLK(n9316), .Q(
        n7912) );
  SDFFX1 DFF_1563_Q_reg ( .D(n4263), .SI(n7912), .SE(n9129), .CLK(n9316), .Q(
        n4598), .QN(n9094) );
  SDFFX1 DFF_1564_Q_reg ( .D(n4269), .SI(n4598), .SE(n9134), .CLK(n9321), .Q(
        g3043) );
  SDFFX1 DFF_1565_Q_reg ( .D(n4268), .SI(g3043), .SE(n9134), .CLK(n9321), .Q(
        g3044) );
  SDFFX1 DFF_1566_Q_reg ( .D(n4267), .SI(g3044), .SE(n9134), .CLK(n9321), .Q(
        g3045) );
  SDFFX1 DFF_1567_Q_reg ( .D(n4266), .SI(g3045), .SE(n9134), .CLK(n9321), .Q(
        g3046) );
  SDFFX1 DFF_1568_Q_reg ( .D(n4265), .SI(g3046), .SE(n9134), .CLK(n9321), .Q(
        g3047) );
  SDFFX1 DFF_1569_Q_reg ( .D(n4272), .SI(g3047), .SE(n9135), .CLK(n9322), .Q(
        g3048) );
  SDFFX1 DFF_1570_Q_reg ( .D(n4271), .SI(g3048), .SE(n9135), .CLK(n9322), .Q(
        g3049) );
  SDFFX1 DFF_1571_Q_reg ( .D(n4270), .SI(g3049), .SE(n9135), .CLK(n9322), .Q(
        g3050) );
  SDFFX1 DFF_1572_Q_reg ( .D(n4259), .SI(g3050), .SE(n9135), .CLK(n9322), .Q(
        g3051) );
  SDFFX1 DFF_1573_Q_reg ( .D(n4236), .SI(g3051), .SE(n9135), .CLK(n9322), .Q(
        g3052) );
  SDFFX1 DFF_1574_Q_reg ( .D(n4239), .SI(g3052), .SE(n9135), .CLK(n9322), .Q(
        g3053) );
  SDFFX1 DFF_1575_Q_reg ( .D(n4237), .SI(g3053), .SE(n9135), .CLK(n9322), .Q(
        test_so96) );
  SDFFX1 DFF_1576_Q_reg ( .D(n4234), .SI(test_si97), .SE(n9233), .CLK(n9420), 
        .Q(g3056) );
  SDFFX1 DFF_1577_Q_reg ( .D(n4233), .SI(g3056), .SE(n9233), .CLK(n9420), .Q(
        g3057) );
  SDFFX1 DFF_1578_Q_reg ( .D(n4238), .SI(g3057), .SE(n9233), .CLK(n9420), .Q(
        g3058) );
  SDFFX1 DFF_1579_Q_reg ( .D(n4235), .SI(g3058), .SE(n9233), .CLK(n9420), .Q(
        g3059) );
  SDFFX1 DFF_1580_Q_reg ( .D(n4240), .SI(g3059), .SE(n9233), .CLK(n9420), .Q(
        g3060) );
  SDFFX1 DFF_1581_Q_reg ( .D(n4232), .SI(g3060), .SE(n9233), .CLK(n9420), .Q(
        g3061) );
  SDFFX1 DFF_1582_Q_reg ( .D(n4245), .SI(g3061), .SE(n9254), .CLK(n9441), .Q(
        g3062) );
  SDFFX1 DFF_1583_Q_reg ( .D(n4248), .SI(g3062), .SE(n9254), .CLK(n9441), .Q(
        g3063) );
  SDFFX1 DFF_1584_Q_reg ( .D(n4246), .SI(g3063), .SE(n9254), .CLK(n9441), .Q(
        g3064) );
  SDFFX1 DFF_1585_Q_reg ( .D(n4243), .SI(g3064), .SE(n9254), .CLK(n9441), .Q(
        g3065) );
  SDFFX1 DFF_1586_Q_reg ( .D(n4242), .SI(g3065), .SE(n9254), .CLK(n9441), .Q(
        g3066) );
  SDFFX1 DFF_1587_Q_reg ( .D(n4247), .SI(g3066), .SE(n9254), .CLK(n9441), .Q(
        g3067) );
  SDFFX1 DFF_1588_Q_reg ( .D(n4244), .SI(g3067), .SE(n9255), .CLK(n9442), .Q(
        g3068) );
  SDFFX1 DFF_1589_Q_reg ( .D(n4249), .SI(g3068), .SE(n9255), .CLK(n9442), .Q(
        g3069) );
  SDFFX1 DFF_1590_Q_reg ( .D(n4241), .SI(g3069), .SE(n9255), .CLK(n9442), .Q(
        test_so97) );
  SDFFX1 DFF_1591_Q_reg ( .D(n4254), .SI(test_si98), .SE(n9150), .CLK(n9337), 
        .Q(g3071) );
  SDFFX1 DFF_1592_Q_reg ( .D(n4257), .SI(g3071), .SE(n9150), .CLK(n9337), .Q(
        g3072) );
  SDFFX1 DFF_1593_Q_reg ( .D(n4255), .SI(g3072), .SE(n9150), .CLK(n9337), .Q(
        g3073) );
  SDFFX1 DFF_1594_Q_reg ( .D(n4252), .SI(g3073), .SE(n9150), .CLK(n9337), .Q(
        g3074) );
  SDFFX1 DFF_1595_Q_reg ( .D(n4251), .SI(g3074), .SE(n9150), .CLK(n9337), .Q(
        g3075) );
  SDFFX1 DFF_1596_Q_reg ( .D(n4256), .SI(g3075), .SE(n9150), .CLK(n9337), .Q(
        g3076) );
  SDFFX1 DFF_1597_Q_reg ( .D(n4253), .SI(g3076), .SE(n9150), .CLK(n9337), .Q(
        g3077) );
  SDFFX1 DFF_1598_Q_reg ( .D(n4258), .SI(g3077), .SE(n9150), .CLK(n9337), .Q(
        g3078) );
  SDFFX1 DFF_1599_Q_reg ( .D(n4250), .SI(g3078), .SE(n9151), .CLK(n9338), .Q(
        g2997) );
  SDFFX1 DFF_1600_Q_reg ( .D(g25265), .SI(g2997), .SE(n9151), .CLK(n9338), .Q(
        g2993), .QN(n9095) );
  SDFFX1 DFF_1601_Q_reg ( .D(g26048), .SI(g2993), .SE(n9151), .CLK(n9338), .Q(
        n7909), .QN(n16493) );
  SDFFX1 DFF_1602_Q_reg ( .D(g23330), .SI(n7909), .SE(n9151), .CLK(n9338), .Q(
        g3006), .QN(n9093) );
  SDFFX1 DFF_1603_Q_reg ( .D(g24445), .SI(g3006), .SE(n9151), .CLK(n9338), .Q(
        g3002), .QN(n8282) );
  SDFFX1 DFF_1604_Q_reg ( .D(g25191), .SI(g3002), .SE(n9151), .CLK(n9338), .Q(
        g3013), .QN(n9092) );
  SDFFX1 DFF_1605_Q_reg ( .D(g26031), .SI(g3013), .SE(n9151), .CLK(n9338), .Q(
        test_so98) );
  SDFFX1 DFF_1606_Q_reg ( .D(g26786), .SI(test_si99), .SE(n9151), .CLK(n9338), 
        .Q(g3024), .QN(n8281) );
  SDFFX1 DFF_1607_Q_reg ( .D(n4262), .SI(g3024), .SE(n9151), .CLK(n9338), .Q(
        g3018), .QN(n4481) );
  SDFFX1 DFF_1608_Q_reg ( .D(g23359), .SI(g3018), .SE(n9152), .CLK(n9339), .Q(
        g3028), .QN(n4350) );
  SDFFX1 DFF_1609_Q_reg ( .D(g24446), .SI(g3028), .SE(n9152), .CLK(n9339), .Q(
        g3036), .QN(n4480) );
  SDFFX1 DFF_1610_Q_reg ( .D(g25202), .SI(g3036), .SE(n9151), .CLK(n9338), .Q(
        g3032), .QN(n9086) );
  SDFFX1 DFF_1611_Q_reg ( .D(g3234), .SI(g3032), .SE(n9151), .CLK(n9338), .Q(
        g5388) );
  SDFFX1 DFF_1612_Q_reg ( .D(g5388), .SI(g5388), .SE(n9151), .CLK(n9338), .Q(
        n7907), .QN(DFF_1612_n1) );
  SDFFX1 DFF_1613_Q_reg ( .D(g16496), .SI(n7907), .SE(n9152), .CLK(n9339), .Q(
        g2987), .QN(n4365) );
  SDFFX1 DFF_1614_Q_reg ( .D(g16824), .SI(g2987), .SE(n9254), .CLK(n9441), .Q(
        g8275), .QN(n9074) );
  SDFFX1 DFF_1615_Q_reg ( .D(g16844), .SI(g8275), .SE(n9254), .CLK(n9441), .Q(
        g8274), .QN(n9076) );
  SDFFX1 DFF_1616_Q_reg ( .D(g16853), .SI(g8274), .SE(n9254), .CLK(n9441), .Q(
        g8273), .QN(n16495) );
  SDFFX1 DFF_1617_Q_reg ( .D(g16860), .SI(g8273), .SE(n9254), .CLK(n9441), .Q(
        g8272), .QN(n16496) );
  SDFFX1 DFF_1618_Q_reg ( .D(g16803), .SI(g8272), .SE(n9254), .CLK(n9441), .Q(
        g8268), .QN(DFF_1618_n1) );
  SDFFX1 DFF_1619_Q_reg ( .D(g16835), .SI(g8268), .SE(n9255), .CLK(n9442), .Q(
        g8269), .QN(n9077) );
  SDFFX1 DFF_1620_Q_reg ( .D(g16851), .SI(g8269), .SE(n9255), .CLK(n9442), .Q(
        test_so99) );
  SDFFX1 DFF_1621_Q_reg ( .D(g16857), .SI(test_si100), .SE(n9255), .CLK(n9442), 
        .Q(g8271), .QN(n9075) );
  SDFFX1 DFF_1622_Q_reg ( .D(g16866), .SI(g8271), .SE(n9255), .CLK(n9442), .Q(
        g3083), .QN(n9080) );
  SDFFX1 DFF_1623_Q_reg ( .D(n4261), .SI(g3083), .SE(n9255), .CLK(n9442), .Q(
        g8267) );
  SDFFX1 DFF_1624_Q_reg ( .D(N995), .SI(g8267), .SE(n9255), .CLK(n9442), .Q(
        n4577) );
  SDFFX1 DFF_1625_Q_reg ( .D(g16845), .SI(n4577), .SE(n9255), .CLK(n9442), .Q(
        g8266), .QN(n16497) );
  SDFFX1 DFF_1626_Q_reg ( .D(g16854), .SI(g8266), .SE(n9255), .CLK(n9442), .Q(
        g8265), .QN(n16498) );
  SDFFX1 DFF_1627_Q_reg ( .D(g16861), .SI(g8265), .SE(n9135), .CLK(n9322), .Q(
        g8264), .QN(n9057) );
  SDFFX1 DFF_1628_Q_reg ( .D(g16880), .SI(g8264), .SE(n9233), .CLK(n9420), .Q(
        g8262), .QN(DFF_1628_n1) );
  SDFFX1 DFF_1629_Q_reg ( .D(g18755), .SI(g8262), .SE(n9233), .CLK(n9420), .Q(
        g8263), .QN(n9058) );
  SDFFX1 DFF_1630_Q_reg ( .D(g18804), .SI(g8263), .SE(n9233), .CLK(n9420), .Q(
        g8260), .QN(n9054) );
  SDFFX1 DFF_1631_Q_reg ( .D(g18837), .SI(g8260), .SE(n9233), .CLK(n9420), .Q(
        g8261), .QN(n9055) );
  SDFFX1 DFF_1632_Q_reg ( .D(g18868), .SI(g8261), .SE(n9233), .CLK(n9420), .Q(
        g8259), .QN(n9056) );
  SDFFX1 DFF_1633_Q_reg ( .D(g18907), .SI(g8259), .SE(n9234), .CLK(n9421), .Q(
        g2990), .QN(n9078) );
  SDFFX1 DFF_1634_Q_reg ( .D(N690), .SI(g2990), .SE(n9135), .CLK(n9322), .Q(
        n4578) );
  SDFFX1 DFF_1635_Q_reg ( .D(n4260), .SI(n4578), .SE(n9259), .CLK(n9446), .Q(
        test_so100) );
  SDFFX1 DFF_454_Q_reg ( .D(n4598), .SI(n8040), .SE(n9147), .CLK(n9334), .Q(
        g6677), .QN(n4309) );
  SDFFX1 DFF_804_Q_reg ( .D(n4598), .SI(test_si49), .SE(n9129), .CLK(n9316), 
        .Q(g6979), .QN(n4308) );
  SDFFX1 DFF_1154_Q_reg ( .D(n4598), .SI(n7960), .SE(n9138), .CLK(n9325), .Q(
        g7229), .QN(n4307) );
  SDFFX1 DFF_1504_Q_reg ( .D(n4598), .SI(n7918), .SE(n9150), .CLK(n9337), .Q(
        g7425), .QN(n4306) );
  SDFFX1 DFF_1300_Q_reg ( .D(g5555), .SI(g5555), .SE(n9236), .CLK(n9423), .Q(
        g7264), .QN(n4524) );
  SDFFX1 DFF_950_Q_reg ( .D(g5511), .SI(g5511), .SE(n9208), .CLK(n9395), .Q(
        g7014), .QN(n4525) );
  SDFFX1 DFF_951_Q_reg ( .D(g7014), .SI(g7014), .SE(n9208), .CLK(n9395), .Q(
        n4618), .QN(n4511) );
  SDFFX1 DFF_1301_Q_reg ( .D(g7264), .SI(g7264), .SE(n9236), .CLK(n9423), .Q(
        n4606), .QN(n4509) );
  SDFFX1 DFF_250_Q_reg ( .D(g5437), .SI(g5437), .SE(n9133), .CLK(n9320), .Q(
        g6447), .QN(n4499) );
  SDFFX1 DFF_249_Q_reg ( .D(g2950), .SI(g181), .SE(n9133), .CLK(n9320), .Q(
        g5437), .QN(n4520) );
  NOR2X0 Trojan1 ( .IN1(n2459), .IN2(n2309), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(n2237), .IN2(n2279), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(n2381), .IN2(n2207), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(n2542), .IN2(n2489), .QN(Tj_OUT4) );
  AND4X1 Trojan1234 ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  OR2X1 Trojan5 ( .IN1(n3260), .IN2(n3301), .Q(Tj_OUT5) );
  OR2X1 Trojan6 ( .IN1(n3380), .IN2(n3341), .Q(Tj_OUT6) );
  OR2X1 Trojan7 ( .IN1(n3374), .IN2(n3293), .Q(Tj_OUT7) );
  OR2X1 Trojan8 ( .IN1(n3334), .IN2(n9117), .Q(Tj_OUT8) );
  AND4X1 Trojan5678 ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND2X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .Q(Tj_Trigger)
         );
  OR2X1 Trojan_Payload_1 ( .IN1(Tj_Trigger), .IN2(n4149), .Q(n4149_Tj_Payload)
         );
  OR2X1 Trojan_Payload_2 ( .IN1(Tj_Trigger), .IN2(n590), .Q(n4161_Tj_Payload)
         );
  OR2X1 Trojan_Payload_3 ( .IN1(Tj_Trigger), .IN2(n869), .Q(n4160_Tj_Payload)
         );
  OR2X1 Trojan_Payload_4 ( .IN1(Tj_Trigger), .IN2(n4122), .Q(n4122_Tj_Payload)
         );
  NBUFFX2 U9017 ( .INP(n9303), .Z(n9129) );
  NBUFFX2 U9018 ( .INP(n9303), .Z(n9130) );
  NBUFFX2 U9019 ( .INP(n9296), .Z(n9151) );
  NBUFFX2 U9020 ( .INP(n9294), .Z(n9156) );
  NBUFFX2 U9021 ( .INP(n9294), .Z(n9155) );
  NBUFFX2 U9022 ( .INP(n9296), .Z(n9150) );
  NBUFFX2 U9023 ( .INP(n9261), .Z(n9254) );
  NBUFFX2 U9024 ( .INP(n9295), .Z(n9154) );
  NBUFFX2 U9025 ( .INP(n9295), .Z(n9153) );
  NBUFFX2 U9026 ( .INP(n9264), .Z(n9247) );
  NBUFFX2 U9027 ( .INP(n9265), .Z(n9243) );
  NBUFFX2 U9028 ( .INP(n9265), .Z(n9244) );
  NBUFFX2 U9029 ( .INP(n9295), .Z(n9152) );
  NBUFFX2 U9030 ( .INP(n9262), .Z(n9252) );
  NBUFFX2 U9031 ( .INP(n9262), .Z(n9251) );
  NBUFFX2 U9032 ( .INP(n9262), .Z(n9253) );
  NBUFFX2 U9033 ( .INP(n9264), .Z(n9246) );
  NBUFFX2 U9034 ( .INP(n9264), .Z(n9245) );
  NBUFFX2 U9035 ( .INP(n9265), .Z(n9242) );
  NBUFFX2 U9036 ( .INP(n9263), .Z(n9248) );
  NBUFFX2 U9037 ( .INP(n9268), .Z(n9235) );
  NBUFFX2 U9038 ( .INP(n9266), .Z(n9241) );
  NBUFFX2 U9039 ( .INP(n9263), .Z(n9250) );
  NBUFFX2 U9040 ( .INP(n9263), .Z(n9249) );
  NBUFFX2 U9041 ( .INP(n9267), .Z(n9237) );
  NBUFFX2 U9042 ( .INP(n9266), .Z(n9240) );
  NBUFFX2 U9043 ( .INP(n9267), .Z(n9236) );
  NBUFFX2 U9044 ( .INP(n9266), .Z(n9239) );
  NBUFFX2 U9045 ( .INP(n9267), .Z(n9238) );
  NBUFFX2 U9046 ( .INP(n9268), .Z(n9234) );
  NBUFFX2 U9047 ( .INP(n9268), .Z(n9233) );
  NBUFFX2 U9048 ( .INP(n9269), .Z(n9230) );
  NBUFFX2 U9049 ( .INP(n9269), .Z(n9232) );
  NBUFFX2 U9050 ( .INP(n9269), .Z(n9231) );
  NBUFFX2 U9051 ( .INP(n9270), .Z(n9228) );
  NBUFFX2 U9052 ( .INP(n9270), .Z(n9227) );
  NBUFFX2 U9053 ( .INP(n9271), .Z(n9226) );
  NBUFFX2 U9054 ( .INP(n9271), .Z(n9225) );
  NBUFFX2 U9055 ( .INP(n9271), .Z(n9224) );
  NBUFFX2 U9056 ( .INP(n9272), .Z(n9223) );
  NBUFFX2 U9057 ( .INP(n9272), .Z(n9222) );
  NBUFFX2 U9058 ( .INP(n9272), .Z(n9221) );
  NBUFFX2 U9059 ( .INP(n9273), .Z(n9220) );
  NBUFFX2 U9060 ( .INP(n9273), .Z(n9219) );
  NBUFFX2 U9061 ( .INP(n9270), .Z(n9229) );
  NBUFFX2 U9062 ( .INP(n9273), .Z(n9218) );
  NBUFFX2 U9063 ( .INP(n9275), .Z(n9214) );
  NBUFFX2 U9064 ( .INP(n9274), .Z(n9215) );
  NBUFFX2 U9065 ( .INP(n9277), .Z(n9208) );
  NBUFFX2 U9066 ( .INP(n9275), .Z(n9213) );
  NBUFFX2 U9067 ( .INP(n9275), .Z(n9212) );
  NBUFFX2 U9068 ( .INP(n9274), .Z(n9217) );
  NBUFFX2 U9069 ( .INP(n9274), .Z(n9216) );
  NBUFFX2 U9070 ( .INP(n9276), .Z(n9211) );
  NBUFFX2 U9071 ( .INP(n9276), .Z(n9210) );
  NBUFFX2 U9072 ( .INP(n9277), .Z(n9207) );
  NBUFFX2 U9073 ( .INP(n9276), .Z(n9209) );
  NBUFFX2 U9074 ( .INP(n9277), .Z(n9206) );
  NBUFFX2 U9075 ( .INP(n9278), .Z(n9205) );
  NBUFFX2 U9076 ( .INP(n9278), .Z(n9204) );
  NBUFFX2 U9077 ( .INP(n9278), .Z(n9203) );
  NBUFFX2 U9078 ( .INP(n9279), .Z(n9202) );
  NBUFFX2 U9079 ( .INP(n9279), .Z(n9201) );
  NBUFFX2 U9080 ( .INP(n9279), .Z(n9200) );
  NBUFFX2 U9081 ( .INP(n9280), .Z(n9199) );
  NBUFFX2 U9082 ( .INP(n9280), .Z(n9198) );
  NBUFFX2 U9083 ( .INP(n9280), .Z(n9197) );
  NBUFFX2 U9084 ( .INP(n9281), .Z(n9196) );
  NBUFFX2 U9085 ( .INP(n9281), .Z(n9195) );
  NBUFFX2 U9086 ( .INP(n9281), .Z(n9194) );
  NBUFFX2 U9087 ( .INP(n9282), .Z(n9193) );
  NBUFFX2 U9088 ( .INP(n9282), .Z(n9192) );
  NBUFFX2 U9089 ( .INP(n9282), .Z(n9191) );
  NBUFFX2 U9090 ( .INP(n9283), .Z(n9188) );
  NBUFFX2 U9091 ( .INP(n9285), .Z(n9183) );
  NBUFFX2 U9092 ( .INP(n9285), .Z(n9182) );
  NBUFFX2 U9093 ( .INP(n9286), .Z(n9181) );
  NBUFFX2 U9094 ( .INP(n9283), .Z(n9190) );
  NBUFFX2 U9095 ( .INP(n9283), .Z(n9189) );
  NBUFFX2 U9096 ( .INP(n9284), .Z(n9187) );
  NBUFFX2 U9097 ( .INP(n9284), .Z(n9186) );
  NBUFFX2 U9098 ( .INP(n9284), .Z(n9185) );
  NBUFFX2 U9099 ( .INP(n9285), .Z(n9184) );
  NBUFFX2 U9100 ( .INP(n9286), .Z(n9180) );
  NBUFFX2 U9101 ( .INP(n9289), .Z(n9171) );
  NBUFFX2 U9102 ( .INP(n9289), .Z(n9170) );
  NBUFFX2 U9103 ( .INP(n9290), .Z(n9169) );
  NBUFFX2 U9104 ( .INP(n9286), .Z(n9179) );
  NBUFFX2 U9105 ( .INP(n9287), .Z(n9178) );
  NBUFFX2 U9106 ( .INP(n9287), .Z(n9177) );
  NBUFFX2 U9107 ( .INP(n9287), .Z(n9176) );
  NBUFFX2 U9108 ( .INP(n9288), .Z(n9175) );
  NBUFFX2 U9109 ( .INP(n9288), .Z(n9174) );
  NBUFFX2 U9110 ( .INP(n9288), .Z(n9173) );
  NBUFFX2 U9111 ( .INP(n9289), .Z(n9172) );
  NBUFFX2 U9112 ( .INP(n9290), .Z(n9168) );
  NBUFFX2 U9113 ( .INP(n9297), .Z(n9146) );
  NBUFFX2 U9114 ( .INP(n9292), .Z(n9163) );
  NBUFFX2 U9115 ( .INP(n9290), .Z(n9167) );
  NBUFFX2 U9116 ( .INP(n9291), .Z(n9166) );
  NBUFFX2 U9117 ( .INP(n9291), .Z(n9164) );
  NBUFFX2 U9118 ( .INP(n9291), .Z(n9165) );
  NBUFFX2 U9119 ( .INP(n9292), .Z(n9162) );
  NBUFFX2 U9120 ( .INP(n9292), .Z(n9161) );
  NBUFFX2 U9121 ( .INP(n9293), .Z(n9160) );
  NBUFFX2 U9122 ( .INP(n9301), .Z(n9134) );
  NBUFFX2 U9123 ( .INP(n9293), .Z(n9159) );
  NBUFFX2 U9124 ( .INP(n9297), .Z(n9148) );
  NBUFFX2 U9125 ( .INP(n9297), .Z(n9147) );
  NBUFFX2 U9126 ( .INP(n9298), .Z(n9145) );
  NBUFFX2 U9127 ( .INP(n9298), .Z(n9144) );
  NBUFFX2 U9128 ( .INP(n9301), .Z(n9135) );
  NBUFFX2 U9129 ( .INP(n9300), .Z(n9137) );
  NBUFFX2 U9130 ( .INP(n9301), .Z(n9136) );
  NBUFFX2 U9131 ( .INP(n9260), .Z(n9258) );
  NBUFFX2 U9132 ( .INP(n9260), .Z(n9257) );
  NBUFFX2 U9133 ( .INP(n9261), .Z(n9256) );
  NBUFFX2 U9134 ( .INP(n9261), .Z(n9255) );
  NBUFFX2 U9135 ( .INP(n9296), .Z(n9149) );
  NBUFFX2 U9136 ( .INP(n9298), .Z(n9143) );
  NBUFFX2 U9137 ( .INP(n9299), .Z(n9142) );
  NBUFFX2 U9138 ( .INP(n9299), .Z(n9141) );
  NBUFFX2 U9139 ( .INP(n9299), .Z(n9140) );
  NBUFFX2 U9140 ( .INP(n9300), .Z(n9139) );
  NBUFFX2 U9141 ( .INP(n9300), .Z(n9138) );
  NBUFFX2 U9142 ( .INP(n9302), .Z(n9131) );
  NBUFFX2 U9143 ( .INP(n9293), .Z(n9158) );
  NBUFFX2 U9144 ( .INP(n9294), .Z(n9157) );
  NBUFFX2 U9145 ( .INP(n9302), .Z(n9133) );
  NBUFFX2 U9146 ( .INP(n9302), .Z(n9132) );
  NBUFFX2 U9147 ( .INP(n9490), .Z(n9316) );
  NBUFFX2 U9148 ( .INP(n9490), .Z(n9317) );
  NBUFFX2 U9149 ( .INP(n9483), .Z(n9338) );
  NBUFFX2 U9150 ( .INP(n9481), .Z(n9343) );
  NBUFFX2 U9151 ( .INP(n9481), .Z(n9342) );
  NBUFFX2 U9152 ( .INP(n9483), .Z(n9337) );
  NBUFFX2 U9153 ( .INP(n9448), .Z(n9441) );
  NBUFFX2 U9154 ( .INP(n9482), .Z(n9341) );
  NBUFFX2 U9155 ( .INP(n9482), .Z(n9340) );
  NBUFFX2 U9156 ( .INP(n9451), .Z(n9434) );
  NBUFFX2 U9157 ( .INP(n9452), .Z(n9430) );
  NBUFFX2 U9158 ( .INP(n9452), .Z(n9431) );
  NBUFFX2 U9159 ( .INP(n9482), .Z(n9339) );
  NBUFFX2 U9160 ( .INP(n9449), .Z(n9439) );
  NBUFFX2 U9161 ( .INP(n9449), .Z(n9438) );
  NBUFFX2 U9162 ( .INP(n9449), .Z(n9440) );
  NBUFFX2 U9163 ( .INP(n9451), .Z(n9433) );
  NBUFFX2 U9164 ( .INP(n9451), .Z(n9432) );
  NBUFFX2 U9165 ( .INP(n9452), .Z(n9429) );
  NBUFFX2 U9166 ( .INP(n9450), .Z(n9435) );
  NBUFFX2 U9167 ( .INP(n9455), .Z(n9422) );
  NBUFFX2 U9168 ( .INP(n9453), .Z(n9428) );
  NBUFFX2 U9169 ( .INP(n9450), .Z(n9437) );
  NBUFFX2 U9170 ( .INP(n9450), .Z(n9436) );
  NBUFFX2 U9171 ( .INP(n9454), .Z(n9424) );
  NBUFFX2 U9172 ( .INP(n9453), .Z(n9427) );
  NBUFFX2 U9173 ( .INP(n9454), .Z(n9423) );
  NBUFFX2 U9174 ( .INP(n9453), .Z(n9426) );
  NBUFFX2 U9175 ( .INP(n9454), .Z(n9425) );
  NBUFFX2 U9176 ( .INP(n9455), .Z(n9421) );
  NBUFFX2 U9177 ( .INP(n9455), .Z(n9420) );
  NBUFFX2 U9178 ( .INP(n9456), .Z(n9417) );
  NBUFFX2 U9179 ( .INP(n9456), .Z(n9419) );
  NBUFFX2 U9180 ( .INP(n9456), .Z(n9418) );
  NBUFFX2 U9181 ( .INP(n9457), .Z(n9415) );
  NBUFFX2 U9182 ( .INP(n9457), .Z(n9414) );
  NBUFFX2 U9183 ( .INP(n9458), .Z(n9413) );
  NBUFFX2 U9184 ( .INP(n9458), .Z(n9412) );
  NBUFFX2 U9185 ( .INP(n9458), .Z(n9411) );
  NBUFFX2 U9186 ( .INP(n9459), .Z(n9410) );
  NBUFFX2 U9187 ( .INP(n9459), .Z(n9409) );
  NBUFFX2 U9188 ( .INP(n9459), .Z(n9408) );
  NBUFFX2 U9189 ( .INP(n9460), .Z(n9407) );
  NBUFFX2 U9190 ( .INP(n9460), .Z(n9406) );
  NBUFFX2 U9191 ( .INP(n9457), .Z(n9416) );
  NBUFFX2 U9192 ( .INP(n9460), .Z(n9405) );
  NBUFFX2 U9193 ( .INP(n9462), .Z(n9401) );
  NBUFFX2 U9194 ( .INP(n9461), .Z(n9402) );
  NBUFFX2 U9195 ( .INP(n9464), .Z(n9395) );
  NBUFFX2 U9196 ( .INP(n9462), .Z(n9400) );
  NBUFFX2 U9197 ( .INP(n9462), .Z(n9399) );
  NBUFFX2 U9198 ( .INP(n9461), .Z(n9404) );
  NBUFFX2 U9199 ( .INP(n9461), .Z(n9403) );
  NBUFFX2 U9200 ( .INP(n9463), .Z(n9398) );
  NBUFFX2 U9201 ( .INP(n9463), .Z(n9397) );
  NBUFFX2 U9202 ( .INP(n9464), .Z(n9394) );
  NBUFFX2 U9203 ( .INP(n9463), .Z(n9396) );
  NBUFFX2 U9204 ( .INP(n9464), .Z(n9393) );
  NBUFFX2 U9205 ( .INP(n9465), .Z(n9392) );
  NBUFFX2 U9206 ( .INP(n9465), .Z(n9391) );
  NBUFFX2 U9207 ( .INP(n9465), .Z(n9390) );
  NBUFFX2 U9208 ( .INP(n9466), .Z(n9389) );
  NBUFFX2 U9209 ( .INP(n9466), .Z(n9388) );
  NBUFFX2 U9210 ( .INP(n9466), .Z(n9387) );
  NBUFFX2 U9211 ( .INP(n9467), .Z(n9386) );
  NBUFFX2 U9212 ( .INP(n9467), .Z(n9385) );
  NBUFFX2 U9213 ( .INP(n9467), .Z(n9384) );
  NBUFFX2 U9214 ( .INP(n9468), .Z(n9383) );
  NBUFFX2 U9215 ( .INP(n9468), .Z(n9382) );
  NBUFFX2 U9216 ( .INP(n9468), .Z(n9381) );
  NBUFFX2 U9217 ( .INP(n9469), .Z(n9380) );
  NBUFFX2 U9218 ( .INP(n9469), .Z(n9379) );
  NBUFFX2 U9219 ( .INP(n9469), .Z(n9378) );
  NBUFFX2 U9220 ( .INP(n9470), .Z(n9375) );
  NBUFFX2 U9221 ( .INP(n9472), .Z(n9370) );
  NBUFFX2 U9222 ( .INP(n9472), .Z(n9369) );
  NBUFFX2 U9223 ( .INP(n9473), .Z(n9368) );
  NBUFFX2 U9224 ( .INP(n9470), .Z(n9377) );
  NBUFFX2 U9225 ( .INP(n9470), .Z(n9376) );
  NBUFFX2 U9226 ( .INP(n9471), .Z(n9374) );
  NBUFFX2 U9227 ( .INP(n9471), .Z(n9373) );
  NBUFFX2 U9228 ( .INP(n9471), .Z(n9372) );
  NBUFFX2 U9229 ( .INP(n9472), .Z(n9371) );
  NBUFFX2 U9230 ( .INP(n9473), .Z(n9367) );
  NBUFFX2 U9231 ( .INP(n9476), .Z(n9358) );
  NBUFFX2 U9232 ( .INP(n9476), .Z(n9357) );
  NBUFFX2 U9233 ( .INP(n9477), .Z(n9356) );
  NBUFFX2 U9234 ( .INP(n9473), .Z(n9366) );
  NBUFFX2 U9235 ( .INP(n9474), .Z(n9365) );
  NBUFFX2 U9236 ( .INP(n9474), .Z(n9364) );
  NBUFFX2 U9237 ( .INP(n9474), .Z(n9363) );
  NBUFFX2 U9238 ( .INP(n9475), .Z(n9362) );
  NBUFFX2 U9239 ( .INP(n9475), .Z(n9361) );
  NBUFFX2 U9240 ( .INP(n9475), .Z(n9360) );
  NBUFFX2 U9241 ( .INP(n9476), .Z(n9359) );
  NBUFFX2 U9242 ( .INP(n9477), .Z(n9355) );
  NBUFFX2 U9243 ( .INP(n9484), .Z(n9333) );
  NBUFFX2 U9244 ( .INP(n9479), .Z(n9350) );
  NBUFFX2 U9245 ( .INP(n9477), .Z(n9354) );
  NBUFFX2 U9246 ( .INP(n9478), .Z(n9353) );
  NBUFFX2 U9247 ( .INP(n9478), .Z(n9351) );
  NBUFFX2 U9248 ( .INP(n9478), .Z(n9352) );
  NBUFFX2 U9249 ( .INP(n9479), .Z(n9349) );
  NBUFFX2 U9250 ( .INP(n9479), .Z(n9348) );
  NBUFFX2 U9251 ( .INP(n9480), .Z(n9347) );
  NBUFFX2 U9252 ( .INP(n9488), .Z(n9321) );
  NBUFFX2 U9253 ( .INP(n9480), .Z(n9346) );
  NBUFFX2 U9254 ( .INP(n9484), .Z(n9335) );
  NBUFFX2 U9255 ( .INP(n9484), .Z(n9334) );
  NBUFFX2 U9256 ( .INP(n9485), .Z(n9332) );
  NBUFFX2 U9257 ( .INP(n9485), .Z(n9331) );
  NBUFFX2 U9258 ( .INP(n9488), .Z(n9322) );
  NBUFFX2 U9259 ( .INP(n9487), .Z(n9324) );
  NBUFFX2 U9260 ( .INP(n9488), .Z(n9323) );
  NBUFFX2 U9261 ( .INP(n9447), .Z(n9445) );
  NBUFFX2 U9262 ( .INP(n9447), .Z(n9444) );
  NBUFFX2 U9263 ( .INP(n9448), .Z(n9443) );
  NBUFFX2 U9264 ( .INP(n9448), .Z(n9442) );
  NBUFFX2 U9265 ( .INP(n9483), .Z(n9336) );
  NBUFFX2 U9266 ( .INP(n9485), .Z(n9330) );
  NBUFFX2 U9267 ( .INP(n9486), .Z(n9329) );
  NBUFFX2 U9268 ( .INP(n9486), .Z(n9328) );
  NBUFFX2 U9269 ( .INP(n9486), .Z(n9327) );
  NBUFFX2 U9270 ( .INP(n9487), .Z(n9326) );
  NBUFFX2 U9271 ( .INP(n9487), .Z(n9325) );
  NBUFFX2 U9272 ( .INP(n9489), .Z(n9318) );
  NBUFFX2 U9273 ( .INP(n9480), .Z(n9345) );
  NBUFFX2 U9274 ( .INP(n9481), .Z(n9344) );
  NBUFFX2 U9275 ( .INP(n9489), .Z(n9320) );
  NBUFFX2 U9276 ( .INP(n9489), .Z(n9319) );
  NBUFFX2 U9277 ( .INP(n9260), .Z(n9259) );
  NBUFFX2 U9278 ( .INP(n9447), .Z(n9446) );
  NBUFFX2 U9279 ( .INP(n9499), .Z(n9449) );
  NBUFFX2 U9280 ( .INP(n9312), .Z(n9262) );
  NBUFFX2 U9281 ( .INP(n9499), .Z(n9450) );
  NBUFFX2 U9282 ( .INP(n9312), .Z(n9263) );
  NBUFFX2 U9283 ( .INP(n9499), .Z(n9447) );
  NBUFFX2 U9284 ( .INP(n9312), .Z(n9260) );
  NBUFFX2 U9285 ( .INP(n9499), .Z(n9448) );
  NBUFFX2 U9286 ( .INP(n9312), .Z(n9261) );
  NBUFFX2 U9287 ( .INP(n9492), .Z(n9482) );
  NBUFFX2 U9288 ( .INP(n9305), .Z(n9295) );
  NBUFFX2 U9289 ( .INP(n9498), .Z(n9451) );
  NBUFFX2 U9290 ( .INP(n9311), .Z(n9264) );
  NBUFFX2 U9291 ( .INP(n9498), .Z(n9452) );
  NBUFFX2 U9292 ( .INP(n9311), .Z(n9265) );
  NBUFFX2 U9293 ( .INP(n9498), .Z(n9453) );
  NBUFFX2 U9294 ( .INP(n9311), .Z(n9266) );
  NBUFFX2 U9295 ( .INP(n9498), .Z(n9454) );
  NBUFFX2 U9296 ( .INP(n9311), .Z(n9267) );
  NBUFFX2 U9297 ( .INP(n9498), .Z(n9455) );
  NBUFFX2 U9298 ( .INP(n9311), .Z(n9268) );
  NBUFFX2 U9299 ( .INP(n9497), .Z(n9456) );
  NBUFFX2 U9300 ( .INP(n9310), .Z(n9269) );
  NBUFFX2 U9301 ( .INP(n9497), .Z(n9458) );
  NBUFFX2 U9302 ( .INP(n9310), .Z(n9271) );
  NBUFFX2 U9303 ( .INP(n9497), .Z(n9459) );
  NBUFFX2 U9304 ( .INP(n9310), .Z(n9272) );
  NBUFFX2 U9305 ( .INP(n9497), .Z(n9457) );
  NBUFFX2 U9306 ( .INP(n9310), .Z(n9270) );
  NBUFFX2 U9307 ( .INP(n9497), .Z(n9460) );
  NBUFFX2 U9308 ( .INP(n9310), .Z(n9273) );
  NBUFFX2 U9309 ( .INP(n9496), .Z(n9462) );
  NBUFFX2 U9310 ( .INP(n9309), .Z(n9275) );
  NBUFFX2 U9311 ( .INP(n9496), .Z(n9461) );
  NBUFFX2 U9312 ( .INP(n9309), .Z(n9274) );
  NBUFFX2 U9313 ( .INP(n9496), .Z(n9463) );
  NBUFFX2 U9314 ( .INP(n9309), .Z(n9276) );
  NBUFFX2 U9315 ( .INP(n9496), .Z(n9464) );
  NBUFFX2 U9316 ( .INP(n9309), .Z(n9277) );
  NBUFFX2 U9317 ( .INP(n9496), .Z(n9465) );
  NBUFFX2 U9318 ( .INP(n9309), .Z(n9278) );
  NBUFFX2 U9319 ( .INP(n9495), .Z(n9466) );
  NBUFFX2 U9320 ( .INP(n9308), .Z(n9279) );
  NBUFFX2 U9321 ( .INP(n9495), .Z(n9467) );
  NBUFFX2 U9322 ( .INP(n9308), .Z(n9280) );
  NBUFFX2 U9323 ( .INP(n9495), .Z(n9468) );
  NBUFFX2 U9324 ( .INP(n9308), .Z(n9281) );
  NBUFFX2 U9325 ( .INP(n9495), .Z(n9469) );
  NBUFFX2 U9326 ( .INP(n9308), .Z(n9282) );
  NBUFFX2 U9327 ( .INP(n9495), .Z(n9470) );
  NBUFFX2 U9328 ( .INP(n9308), .Z(n9283) );
  NBUFFX2 U9329 ( .INP(n9494), .Z(n9471) );
  NBUFFX2 U9330 ( .INP(n9307), .Z(n9284) );
  NBUFFX2 U9331 ( .INP(n9494), .Z(n9472) );
  NBUFFX2 U9332 ( .INP(n9307), .Z(n9285) );
  NBUFFX2 U9333 ( .INP(n9494), .Z(n9473) );
  NBUFFX2 U9334 ( .INP(n9307), .Z(n9286) );
  NBUFFX2 U9335 ( .INP(n9494), .Z(n9474) );
  NBUFFX2 U9336 ( .INP(n9307), .Z(n9287) );
  NBUFFX2 U9337 ( .INP(n9494), .Z(n9475) );
  NBUFFX2 U9338 ( .INP(n9307), .Z(n9288) );
  NBUFFX2 U9339 ( .INP(n9493), .Z(n9476) );
  NBUFFX2 U9340 ( .INP(n9306), .Z(n9289) );
  NBUFFX2 U9341 ( .INP(n9493), .Z(n9477) );
  NBUFFX2 U9342 ( .INP(n9306), .Z(n9290) );
  NBUFFX2 U9343 ( .INP(n9493), .Z(n9478) );
  NBUFFX2 U9344 ( .INP(n9306), .Z(n9291) );
  NBUFFX2 U9345 ( .INP(n9493), .Z(n9479) );
  NBUFFX2 U9346 ( .INP(n9306), .Z(n9292) );
  NBUFFX2 U9347 ( .INP(n9492), .Z(n9484) );
  NBUFFX2 U9348 ( .INP(n9305), .Z(n9297) );
  NBUFFX2 U9349 ( .INP(n9491), .Z(n9488) );
  NBUFFX2 U9350 ( .INP(n9304), .Z(n9301) );
  NBUFFX2 U9351 ( .INP(n9492), .Z(n9483) );
  NBUFFX2 U9352 ( .INP(n9305), .Z(n9296) );
  NBUFFX2 U9353 ( .INP(n9492), .Z(n9485) );
  NBUFFX2 U9354 ( .INP(n9305), .Z(n9298) );
  NBUFFX2 U9355 ( .INP(n9491), .Z(n9486) );
  NBUFFX2 U9356 ( .INP(n9304), .Z(n9299) );
  NBUFFX2 U9357 ( .INP(n9491), .Z(n9487) );
  NBUFFX2 U9358 ( .INP(n9304), .Z(n9300) );
  NBUFFX2 U9359 ( .INP(n9493), .Z(n9480) );
  NBUFFX2 U9360 ( .INP(n9306), .Z(n9293) );
  NBUFFX2 U9361 ( .INP(n9492), .Z(n9481) );
  NBUFFX2 U9362 ( .INP(n9305), .Z(n9294) );
  NBUFFX2 U9363 ( .INP(n9491), .Z(n9489) );
  NBUFFX2 U9364 ( .INP(n9304), .Z(n9302) );
  NBUFFX2 U9365 ( .INP(n9491), .Z(n9490) );
  NBUFFX2 U9366 ( .INP(n9304), .Z(n9303) );
  NBUFFX2 U9367 ( .INP(n9315), .Z(n9304) );
  NBUFFX2 U9368 ( .INP(n9315), .Z(n9305) );
  NBUFFX2 U9369 ( .INP(n9315), .Z(n9306) );
  NBUFFX2 U9370 ( .INP(n9314), .Z(n9307) );
  NBUFFX2 U9371 ( .INP(n9314), .Z(n9308) );
  NBUFFX2 U9372 ( .INP(n9314), .Z(n9309) );
  NBUFFX2 U9373 ( .INP(n9313), .Z(n9310) );
  NBUFFX2 U9374 ( .INP(n9313), .Z(n9311) );
  NBUFFX2 U9375 ( .INP(n9313), .Z(n9312) );
  NBUFFX2 U9376 ( .INP(test_se), .Z(n9313) );
  NBUFFX2 U9377 ( .INP(test_se), .Z(n9314) );
  NBUFFX2 U9378 ( .INP(test_se), .Z(n9315) );
  NBUFFX2 U9379 ( .INP(n9502), .Z(n9491) );
  NBUFFX2 U9380 ( .INP(n9502), .Z(n9492) );
  NBUFFX2 U9381 ( .INP(n9502), .Z(n9493) );
  NBUFFX2 U9382 ( .INP(n9501), .Z(n9494) );
  NBUFFX2 U9383 ( .INP(n9501), .Z(n9495) );
  NBUFFX2 U9384 ( .INP(n9501), .Z(n9496) );
  NBUFFX2 U9385 ( .INP(n9500), .Z(n9497) );
  NBUFFX2 U9386 ( .INP(n9500), .Z(n9498) );
  NBUFFX2 U9387 ( .INP(n9500), .Z(n9499) );
  NBUFFX2 U9388 ( .INP(CK), .Z(n9500) );
  NBUFFX2 U9389 ( .INP(CK), .Z(n9501) );
  NBUFFX2 U9390 ( .INP(CK), .Z(n9502) );
  INVX0 U9391 ( .INP(n9503), .ZN(n932) );
  INVX0 U9392 ( .INP(n9504), .ZN(n811) );
  INVX0 U9393 ( .INP(n9505), .ZN(n8) );
  AND2X1 U9394 ( .IN1(n9506), .IN2(n9507), .Q(n9505) );
  OR2X1 U9395 ( .IN1(n9508), .IN2(n9509), .Q(n9506) );
  AND2X1 U9396 ( .IN1(n9510), .IN2(n4482), .Q(n9508) );
  INVX0 U9397 ( .INP(n9511), .ZN(n785) );
  INVX0 U9398 ( .INP(n9512), .ZN(n640) );
  INVX0 U9399 ( .INP(n9513), .ZN(n519) );
  INVX0 U9400 ( .INP(n9514), .ZN(n516) );
  INVX0 U9401 ( .INP(n9515), .ZN(n492) );
  INVX0 U9402 ( .INP(n9516), .ZN(n488) );
  INVX0 U9403 ( .INP(n9517), .ZN(n484) );
  XOR2X1 U9404 ( .IN1(n9079), .IN2(n9518), .Q(n4281) );
  XOR2X1 U9405 ( .IN1(g2934), .IN2(n9519), .Q(n4280) );
  OR2X1 U9406 ( .IN1(n9520), .IN2(n4351), .Q(n4279) );
  AND2X1 U9407 ( .IN1(DFF_18_n1), .IN2(g8021), .Q(n9520) );
  AND2X1 U9408 ( .IN1(n9521), .IN2(n9522), .Q(n4278) );
  OR2X1 U9409 ( .IN1(n9523), .IN2(n9524), .Q(n9522) );
  OR2X1 U9410 ( .IN1(n9525), .IN2(n9526), .Q(n9524) );
  OR2X1 U9411 ( .IN1(n9527), .IN2(n9528), .Q(n9526) );
  OR2X1 U9412 ( .IN1(n9529), .IN2(n9530), .Q(n9528) );
  XNOR2X1 U9413 ( .IN1(n9113), .IN2(n9531), .Q(n9530) );
  XNOR2X1 U9414 ( .IN1(n9096), .IN2(n9532), .Q(n9529) );
  XNOR2X1 U9415 ( .IN1(n9105), .IN2(n9533), .Q(n9527) );
  OR2X1 U9416 ( .IN1(n9534), .IN2(n9535), .Q(n9525) );
  OR2X1 U9417 ( .IN1(n9536), .IN2(n9537), .Q(n9535) );
  XNOR2X1 U9418 ( .IN1(n8818), .IN2(n9538), .Q(n9537) );
  XNOR2X1 U9419 ( .IN1(n8286), .IN2(n9539), .Q(n9536) );
  XNOR2X1 U9420 ( .IN1(n8440), .IN2(n9540), .Q(n9534) );
  OR2X1 U9421 ( .IN1(n9541), .IN2(n9542), .Q(n9523) );
  OR2X1 U9422 ( .IN1(n9543), .IN2(n9544), .Q(n9542) );
  OR2X1 U9423 ( .IN1(n9545), .IN2(n9546), .Q(n9544) );
  XNOR2X1 U9424 ( .IN1(n8821), .IN2(n9547), .Q(n9546) );
  XNOR2X1 U9425 ( .IN1(n8820), .IN2(n9548), .Q(n9545) );
  XNOR2X1 U9426 ( .IN1(n8819), .IN2(n9549), .Q(n9543) );
  OR2X1 U9427 ( .IN1(n9550), .IN2(n9551), .Q(n9541) );
  OR2X1 U9428 ( .IN1(n9552), .IN2(n9553), .Q(n9551) );
  XOR2X1 U9429 ( .IN1(test_so15), .IN2(n9554), .Q(n9550) );
  OR2X1 U9430 ( .IN1(n9555), .IN2(n9556), .Q(n9521) );
  AND2X1 U9431 ( .IN1(n9557), .IN2(n9558), .Q(n4277) );
  OR2X1 U9432 ( .IN1(n9559), .IN2(n9560), .Q(n9558) );
  OR2X1 U9433 ( .IN1(n9561), .IN2(n9562), .Q(n9560) );
  OR2X1 U9434 ( .IN1(n9563), .IN2(n9564), .Q(n9562) );
  OR2X1 U9435 ( .IN1(n9565), .IN2(n9566), .Q(n9564) );
  XNOR2X1 U9436 ( .IN1(n9100), .IN2(n9567), .Q(n9566) );
  XNOR2X1 U9437 ( .IN1(n9099), .IN2(n9568), .Q(n9565) );
  XNOR2X1 U9438 ( .IN1(n9101), .IN2(n9569), .Q(n9563) );
  OR2X1 U9439 ( .IN1(n9570), .IN2(n9571), .Q(n9561) );
  OR2X1 U9440 ( .IN1(n9572), .IN2(n9573), .Q(n9571) );
  XNOR2X1 U9441 ( .IN1(n8814), .IN2(n9574), .Q(n9573) );
  XOR2X1 U9442 ( .IN1(n8285), .IN2(n9575), .Q(n9572) );
  XNOR2X1 U9443 ( .IN1(n8817), .IN2(n9576), .Q(n9570) );
  OR2X1 U9444 ( .IN1(n9577), .IN2(n9578), .Q(n9559) );
  OR2X1 U9445 ( .IN1(n9579), .IN2(n9580), .Q(n9578) );
  OR2X1 U9446 ( .IN1(n9581), .IN2(n9582), .Q(n9580) );
  XNOR2X1 U9447 ( .IN1(n8815), .IN2(n9583), .Q(n9582) );
  XNOR2X1 U9448 ( .IN1(n8439), .IN2(n9584), .Q(n9581) );
  XNOR2X1 U9449 ( .IN1(n8816), .IN2(n9585), .Q(n9579) );
  OR2X1 U9450 ( .IN1(n9586), .IN2(n9587), .Q(n9577) );
  OR2X1 U9451 ( .IN1(n9552), .IN2(n9588), .Q(n9587) );
  XOR2X1 U9452 ( .IN1(test_so36), .IN2(n9589), .Q(n9586) );
  OR2X1 U9453 ( .IN1(n2542), .IN2(n9590), .Q(n9557) );
  AND2X1 U9454 ( .IN1(n9591), .IN2(n9592), .Q(n4276) );
  OR2X1 U9455 ( .IN1(n9593), .IN2(n9594), .Q(n9592) );
  OR2X1 U9456 ( .IN1(n9595), .IN2(n9596), .Q(n9594) );
  OR2X1 U9457 ( .IN1(n9597), .IN2(n9598), .Q(n9596) );
  OR2X1 U9458 ( .IN1(n9599), .IN2(n9600), .Q(n9598) );
  XNOR2X1 U9459 ( .IN1(n9114), .IN2(n9601), .Q(n9600) );
  XNOR2X1 U9460 ( .IN1(n9097), .IN2(n9602), .Q(n9599) );
  XNOR2X1 U9461 ( .IN1(n9103), .IN2(n9603), .Q(n9597) );
  OR2X1 U9462 ( .IN1(n9604), .IN2(n9605), .Q(n9595) );
  OR2X1 U9463 ( .IN1(n9606), .IN2(n9607), .Q(n9605) );
  XNOR2X1 U9464 ( .IN1(n8813), .IN2(n9608), .Q(n9607) );
  XNOR2X1 U9465 ( .IN1(n8284), .IN2(n9609), .Q(n9606) );
  XNOR2X1 U9466 ( .IN1(n9115), .IN2(n9610), .Q(n9604) );
  OR2X1 U9467 ( .IN1(n9611), .IN2(n9612), .Q(n9593) );
  OR2X1 U9468 ( .IN1(n9613), .IN2(n9614), .Q(n9612) );
  OR2X1 U9469 ( .IN1(n9615), .IN2(n9616), .Q(n9614) );
  XNOR2X1 U9470 ( .IN1(n8812), .IN2(n9617), .Q(n9616) );
  XNOR2X1 U9471 ( .IN1(n8438), .IN2(n9618), .Q(n9615) );
  XNOR2X1 U9472 ( .IN1(n8810), .IN2(n9619), .Q(n9613) );
  OR2X1 U9473 ( .IN1(n9620), .IN2(n9621), .Q(n9611) );
  OR2X1 U9474 ( .IN1(n9552), .IN2(n9622), .Q(n9621) );
  XNOR2X1 U9475 ( .IN1(n8811), .IN2(n9623), .Q(n9620) );
  OR2X1 U9476 ( .IN1(n9624), .IN2(n9625), .Q(n9591) );
  AND2X1 U9477 ( .IN1(n9626), .IN2(n9627), .Q(n4275) );
  OR2X1 U9478 ( .IN1(n9628), .IN2(n9629), .Q(n9627) );
  OR2X1 U9479 ( .IN1(n9630), .IN2(n9631), .Q(n9629) );
  OR2X1 U9480 ( .IN1(n9632), .IN2(n9633), .Q(n9631) );
  OR2X1 U9481 ( .IN1(n9634), .IN2(n9635), .Q(n9633) );
  XNOR2X1 U9482 ( .IN1(n8283), .IN2(n9636), .Q(n9635) );
  XNOR2X1 U9483 ( .IN1(n9098), .IN2(n9637), .Q(n9634) );
  XNOR2X1 U9484 ( .IN1(n9104), .IN2(n9638), .Q(n9632) );
  OR2X1 U9485 ( .IN1(n9639), .IN2(n9640), .Q(n9630) );
  OR2X1 U9486 ( .IN1(n9641), .IN2(n9642), .Q(n9640) );
  XNOR2X1 U9487 ( .IN1(n8437), .IN2(n9643), .Q(n9642) );
  XNOR2X1 U9488 ( .IN1(n9116), .IN2(n9644), .Q(n9641) );
  XNOR2X1 U9489 ( .IN1(n8809), .IN2(n9645), .Q(n9639) );
  OR2X1 U9490 ( .IN1(n9646), .IN2(n9647), .Q(n9628) );
  OR2X1 U9491 ( .IN1(n9648), .IN2(n9649), .Q(n9647) );
  OR2X1 U9492 ( .IN1(n9650), .IN2(n9651), .Q(n9649) );
  XNOR2X1 U9493 ( .IN1(n8807), .IN2(n9652), .Q(n9651) );
  XNOR2X1 U9494 ( .IN1(n8806), .IN2(n9653), .Q(n9650) );
  XNOR2X1 U9495 ( .IN1(n8808), .IN2(n9654), .Q(n9648) );
  OR2X1 U9496 ( .IN1(n9655), .IN2(n9656), .Q(n9646) );
  OR2X1 U9497 ( .IN1(n9552), .IN2(n9657), .Q(n9656) );
  XNOR2X1 U9498 ( .IN1(test_so78), .IN2(n9658), .Q(n9655) );
  OR2X1 U9499 ( .IN1(n2489), .IN2(n9659), .Q(n9626) );
  OR2X1 U9500 ( .IN1(n9660), .IN2(n9661), .Q(n4274) );
  INVX0 U9501 ( .INP(n9662), .ZN(n9661) );
  AND2X1 U9502 ( .IN1(n9663), .IN2(n9664), .Q(n9660) );
  INVX0 U9503 ( .INP(n9665), .ZN(n9663) );
  AND2X1 U9504 ( .IN1(n4330), .IN2(n4423), .Q(n9665) );
  OR2X1 U9505 ( .IN1(n9666), .IN2(n9667), .Q(n4272) );
  OR2X1 U9506 ( .IN1(n9668), .IN2(n9669), .Q(n9667) );
  AND2X1 U9507 ( .IN1(test_so27), .IN2(n9670), .Q(n9669) );
  AND2X1 U9508 ( .IN1(n9671), .IN2(n9672), .Q(n9668) );
  OR2X1 U9509 ( .IN1(n9673), .IN2(n9674), .Q(n4271) );
  OR2X1 U9510 ( .IN1(n9675), .IN2(n9676), .Q(n9674) );
  AND2X1 U9511 ( .IN1(n9670), .IN2(g536), .Q(n9676) );
  AND2X1 U9512 ( .IN1(n9671), .IN2(n9677), .Q(n9675) );
  AND2X1 U9513 ( .IN1(n2446), .IN2(n9678), .Q(n9673) );
  OR2X1 U9514 ( .IN1(n9679), .IN2(n9680), .Q(n4270) );
  OR2X1 U9515 ( .IN1(n9681), .IN2(n9682), .Q(n9680) );
  AND2X1 U9516 ( .IN1(n9670), .IN2(g537), .Q(n9682) );
  AND2X1 U9517 ( .IN1(n9671), .IN2(n9683), .Q(n9681) );
  AND2X1 U9518 ( .IN1(n2446), .IN2(n9684), .Q(n9679) );
  OR2X1 U9519 ( .IN1(n9685), .IN2(n9686), .Q(n4269) );
  OR2X1 U9520 ( .IN1(n9687), .IN2(n9688), .Q(n9686) );
  AND2X1 U9521 ( .IN1(n9670), .IN2(n8047), .Q(n9688) );
  AND2X1 U9522 ( .IN1(n9689), .IN2(n9690), .Q(n9687) );
  AND2X1 U9523 ( .IN1(n9691), .IN2(n9692), .Q(n9689) );
  OR2X1 U9524 ( .IN1(n9693), .IN2(n9694), .Q(n4268) );
  OR2X1 U9525 ( .IN1(n9695), .IN2(n9696), .Q(n9693) );
  AND2X1 U9526 ( .IN1(n9670), .IN2(n8046), .Q(n9696) );
  AND2X1 U9527 ( .IN1(n9697), .IN2(n9690), .Q(n9695) );
  AND2X1 U9528 ( .IN1(n9698), .IN2(n9692), .Q(n9697) );
  OR2X1 U9529 ( .IN1(n9699), .IN2(n9694), .Q(n4267) );
  OR2X1 U9530 ( .IN1(n9666), .IN2(n9700), .Q(n9694) );
  INVX0 U9531 ( .INP(n2440), .ZN(n9700) );
  OR2X1 U9532 ( .IN1(n9701), .IN2(n9702), .Q(n9699) );
  AND2X1 U9533 ( .IN1(n9670), .IN2(n8045), .Q(n9702) );
  AND2X1 U9534 ( .IN1(n9703), .IN2(n9690), .Q(n9701) );
  AND2X1 U9535 ( .IN1(n9704), .IN2(n9692), .Q(n9703) );
  OR2X1 U9536 ( .IN1(n9685), .IN2(n9705), .Q(n4266) );
  OR2X1 U9537 ( .IN1(n9706), .IN2(n9707), .Q(n9705) );
  AND2X1 U9538 ( .IN1(n9670), .IN2(n8044), .Q(n9707) );
  AND2X1 U9539 ( .IN1(n9708), .IN2(n9690), .Q(n9706) );
  AND2X1 U9540 ( .IN1(n9709), .IN2(n9692), .Q(n9708) );
  OR2X1 U9541 ( .IN1(n9710), .IN2(n9666), .Q(n9685) );
  AND2X1 U9542 ( .IN1(n2446), .IN2(n2445), .Q(n9710) );
  OR2X1 U9543 ( .IN1(n9666), .IN2(n9711), .Q(n4265) );
  OR2X1 U9544 ( .IN1(n9712), .IN2(n9713), .Q(n9711) );
  AND2X1 U9545 ( .IN1(n9670), .IN2(n8043), .Q(n9713) );
  AND2X1 U9546 ( .IN1(n9714), .IN2(n9690), .Q(n9670) );
  AND2X1 U9547 ( .IN1(n9671), .IN2(n9715), .Q(n9712) );
  AND2X1 U9548 ( .IN1(n9692), .IN2(n9690), .Q(n9671) );
  INVX0 U9549 ( .INP(n9716), .ZN(n9690) );
  INVX0 U9550 ( .INP(n2426), .ZN(n9666) );
  OR2X1 U9551 ( .IN1(g3234), .IN2(n7912), .Q(n4263) );
  INVX0 U9552 ( .INP(n9717), .ZN(n4262) );
  AND2X1 U9553 ( .IN1(n9718), .IN2(n9719), .Q(n9717) );
  OR2X1 U9554 ( .IN1(n9720), .IN2(n9721), .Q(n9718) );
  AND2X1 U9555 ( .IN1(n9722), .IN2(n4481), .Q(n9720) );
  XOR2X1 U9556 ( .IN1(n9723), .IN2(n9724), .Q(n4261) );
  XOR2X1 U9557 ( .IN1(n9725), .IN2(n9723), .Q(n4260) );
  OR2X1 U9558 ( .IN1(n16492), .IN2(g3231), .Q(n9723) );
  OR2X1 U9559 ( .IN1(n9726), .IN2(n9727), .Q(n4259) );
  OR2X1 U9560 ( .IN1(n9728), .IN2(n9729), .Q(n9727) );
  AND2X1 U9561 ( .IN1(n9730), .IN2(g557), .Q(n9729) );
  XOR2X1 U9562 ( .IN1(n9678), .IN2(n9684), .Q(n9730) );
  OR2X1 U9563 ( .IN1(n9731), .IN2(n9732), .Q(n9684) );
  OR2X1 U9564 ( .IN1(n9733), .IN2(n9734), .Q(n9731) );
  AND2X1 U9565 ( .IN1(n9735), .IN2(n9736), .Q(n9734) );
  AND2X1 U9566 ( .IN1(n9737), .IN2(n9738), .Q(n9733) );
  OR2X1 U9567 ( .IN1(n9739), .IN2(n9740), .Q(n9678) );
  OR2X1 U9568 ( .IN1(n9741), .IN2(n9742), .Q(n9740) );
  AND2X1 U9569 ( .IN1(n9743), .IN2(n9744), .Q(n9742) );
  AND2X1 U9570 ( .IN1(n9745), .IN2(n9746), .Q(n9741) );
  AND2X1 U9571 ( .IN1(n9747), .IN2(n9748), .Q(n9728) );
  AND2X1 U9572 ( .IN1(n9749), .IN2(n9750), .Q(n9748) );
  OR2X1 U9573 ( .IN1(g3229), .IN2(n8040), .Q(n9750) );
  INVX0 U9574 ( .INP(n9751), .ZN(n9749) );
  AND2X1 U9575 ( .IN1(g3229), .IN2(n4492), .Q(n9751) );
  INVX0 U9576 ( .INP(n9752), .ZN(n9747) );
  OR2X1 U9577 ( .IN1(n9692), .IN2(n9716), .Q(n9752) );
  OR2X1 U9578 ( .IN1(n9517), .IN2(n9753), .Q(n9692) );
  AND2X1 U9579 ( .IN1(test_so22), .IN2(n9754), .Q(n9726) );
  XOR2X1 U9580 ( .IN1(n9755), .IN2(n9756), .Q(n9754) );
  XOR2X1 U9581 ( .IN1(n9757), .IN2(n9758), .Q(n9756) );
  XNOR2X1 U9582 ( .IN1(n9715), .IN2(n9709), .Q(n9758) );
  OR2X1 U9583 ( .IN1(n9759), .IN2(n9760), .Q(n9709) );
  OR2X1 U9584 ( .IN1(n9761), .IN2(n9762), .Q(n9760) );
  AND2X1 U9585 ( .IN1(n9735), .IN2(n9763), .Q(n9762) );
  AND2X1 U9586 ( .IN1(n9764), .IN2(n9738), .Q(n9761) );
  INVX0 U9587 ( .INP(n9763), .ZN(n9764) );
  OR2X1 U9588 ( .IN1(n9739), .IN2(n9765), .Q(n9715) );
  OR2X1 U9589 ( .IN1(n9766), .IN2(n9767), .Q(n9765) );
  AND2X1 U9590 ( .IN1(n9768), .IN2(n9744), .Q(n9767) );
  AND2X1 U9591 ( .IN1(n9745), .IN2(n9769), .Q(n9766) );
  XNOR2X1 U9592 ( .IN1(n9704), .IN2(n9698), .Q(n9757) );
  OR2X1 U9593 ( .IN1(n9759), .IN2(n9770), .Q(n9698) );
  OR2X1 U9594 ( .IN1(n9771), .IN2(n9772), .Q(n9770) );
  AND2X1 U9595 ( .IN1(n9735), .IN2(n9773), .Q(n9772) );
  AND2X1 U9596 ( .IN1(n9774), .IN2(n9738), .Q(n9771) );
  OR2X1 U9597 ( .IN1(n9759), .IN2(n9775), .Q(n9704) );
  OR2X1 U9598 ( .IN1(n9776), .IN2(n9777), .Q(n9775) );
  AND2X1 U9599 ( .IN1(n9778), .IN2(n9744), .Q(n9777) );
  INVX0 U9600 ( .INP(n9779), .ZN(n9778) );
  AND2X1 U9601 ( .IN1(n9745), .IN2(n9779), .Q(n9776) );
  XOR2X1 U9602 ( .IN1(n9780), .IN2(n9781), .Q(n9755) );
  XNOR2X1 U9603 ( .IN1(n9691), .IN2(n9683), .Q(n9781) );
  OR2X1 U9604 ( .IN1(n9759), .IN2(n9782), .Q(n9683) );
  OR2X1 U9605 ( .IN1(n9783), .IN2(n9784), .Q(n9782) );
  AND2X1 U9606 ( .IN1(n9735), .IN2(n9785), .Q(n9784) );
  AND2X1 U9607 ( .IN1(n9786), .IN2(n9738), .Q(n9783) );
  INVX0 U9608 ( .INP(n9785), .ZN(n9786) );
  OR2X1 U9609 ( .IN1(n9759), .IN2(n9787), .Q(n9691) );
  OR2X1 U9610 ( .IN1(n9788), .IN2(n9789), .Q(n9787) );
  AND2X1 U9611 ( .IN1(n9790), .IN2(n9744), .Q(n9789) );
  INVX0 U9612 ( .INP(n9791), .ZN(n9790) );
  AND2X1 U9613 ( .IN1(n9745), .IN2(n9791), .Q(n9788) );
  XNOR2X1 U9614 ( .IN1(n9677), .IN2(n9672), .Q(n9780) );
  OR2X1 U9615 ( .IN1(n9792), .IN2(n9732), .Q(n9672) );
  OR2X1 U9616 ( .IN1(n9793), .IN2(n9759), .Q(n9732) );
  INVX0 U9617 ( .INP(n2459), .ZN(n9793) );
  OR2X1 U9618 ( .IN1(n9794), .IN2(n9795), .Q(n9792) );
  AND2X1 U9619 ( .IN1(n9735), .IN2(n9796), .Q(n9795) );
  AND2X1 U9620 ( .IN1(n9797), .IN2(n9798), .Q(n9735) );
  AND2X1 U9621 ( .IN1(n9799), .IN2(n9738), .Q(n9794) );
  OR2X1 U9622 ( .IN1(n9739), .IN2(n9800), .Q(n9677) );
  OR2X1 U9623 ( .IN1(n9801), .IN2(n9802), .Q(n9800) );
  AND2X1 U9624 ( .IN1(n9803), .IN2(n9744), .Q(n9802) );
  AND2X1 U9625 ( .IN1(n9745), .IN2(n9804), .Q(n9801) );
  AND2X1 U9626 ( .IN1(n9797), .IN2(n9805), .Q(n9745) );
  OR2X1 U9627 ( .IN1(n9806), .IN2(n9759), .Q(n9739) );
  OR2X1 U9628 ( .IN1(n4541), .IN2(n9517), .Q(n9759) );
  OR2X1 U9629 ( .IN1(n9807), .IN2(n9808), .Q(n9517) );
  OR2X1 U9630 ( .IN1(g559), .IN2(g21851), .Q(n9808) );
  OR2X1 U9631 ( .IN1(g563), .IN2(n9809), .Q(n9807) );
  AND2X1 U9632 ( .IN1(n4541), .IN2(n9810), .Q(n9809) );
  INVX0 U9633 ( .INP(n9811), .ZN(n9806) );
  OR2X1 U9634 ( .IN1(n9797), .IN2(n9805), .Q(n9811) );
  OR2X1 U9635 ( .IN1(n9812), .IN2(n9813), .Q(n4258) );
  OR2X1 U9636 ( .IN1(n9814), .IN2(n9815), .Q(n9813) );
  AND2X1 U9637 ( .IN1(n9816), .IN2(g2611), .Q(n9815) );
  AND2X1 U9638 ( .IN1(n9817), .IN2(n9818), .Q(n9814) );
  AND2X1 U9639 ( .IN1(n2361), .IN2(n9819), .Q(n9812) );
  OR2X1 U9640 ( .IN1(n9820), .IN2(n9821), .Q(n4257) );
  OR2X1 U9641 ( .IN1(n9822), .IN2(n9823), .Q(n9821) );
  AND2X1 U9642 ( .IN1(n9816), .IN2(n7924), .Q(n9822) );
  OR2X1 U9643 ( .IN1(n9824), .IN2(n9825), .Q(n9820) );
  AND2X1 U9644 ( .IN1(n9826), .IN2(n9827), .Q(n9825) );
  AND2X1 U9645 ( .IN1(n9828), .IN2(n9829), .Q(n9826) );
  OR2X1 U9646 ( .IN1(n9830), .IN2(n9831), .Q(n4256) );
  OR2X1 U9647 ( .IN1(n9824), .IN2(n9832), .Q(n9831) );
  AND2X1 U9648 ( .IN1(n9817), .IN2(n9833), .Q(n9832) );
  AND2X1 U9649 ( .IN1(n9816), .IN2(n7920), .Q(n9830) );
  OR2X1 U9650 ( .IN1(n9834), .IN2(n9835), .Q(n4255) );
  OR2X1 U9651 ( .IN1(n9836), .IN2(n9823), .Q(n9835) );
  INVX0 U9652 ( .INP(n2375), .ZN(n9823) );
  AND2X1 U9653 ( .IN1(n9816), .IN2(n7923), .Q(n9836) );
  OR2X1 U9654 ( .IN1(n9824), .IN2(n9837), .Q(n9834) );
  AND2X1 U9655 ( .IN1(n9838), .IN2(n9827), .Q(n9837) );
  AND2X1 U9656 ( .IN1(n9839), .IN2(n9829), .Q(n9838) );
  OR2X1 U9657 ( .IN1(n9840), .IN2(n9841), .Q(n4254) );
  OR2X1 U9658 ( .IN1(n9842), .IN2(n9843), .Q(n9841) );
  AND2X1 U9659 ( .IN1(n9816), .IN2(n7925), .Q(n9843) );
  AND2X1 U9660 ( .IN1(n9844), .IN2(n9827), .Q(n9842) );
  AND2X1 U9661 ( .IN1(n9845), .IN2(n9829), .Q(n9844) );
  OR2X1 U9662 ( .IN1(n9846), .IN2(n9847), .Q(n4253) );
  OR2X1 U9663 ( .IN1(n9848), .IN2(n9849), .Q(n9847) );
  AND2X1 U9664 ( .IN1(test_so91), .IN2(n9816), .Q(n9849) );
  AND2X1 U9665 ( .IN1(n9817), .IN2(n9850), .Q(n9848) );
  AND2X1 U9666 ( .IN1(n2361), .IN2(n9851), .Q(n9846) );
  OR2X1 U9667 ( .IN1(n9840), .IN2(n9852), .Q(n4252) );
  OR2X1 U9668 ( .IN1(n9853), .IN2(n9854), .Q(n9852) );
  AND2X1 U9669 ( .IN1(n9816), .IN2(n7922), .Q(n9854) );
  AND2X1 U9670 ( .IN1(n9855), .IN2(n9827), .Q(n9853) );
  AND2X1 U9671 ( .IN1(n9856), .IN2(n9829), .Q(n9855) );
  OR2X1 U9672 ( .IN1(n9824), .IN2(n9857), .Q(n9840) );
  AND2X1 U9673 ( .IN1(n2361), .IN2(n2374), .Q(n9857) );
  OR2X1 U9674 ( .IN1(n9858), .IN2(n9859), .Q(n4251) );
  OR2X1 U9675 ( .IN1(n9824), .IN2(n9860), .Q(n9859) );
  AND2X1 U9676 ( .IN1(n9817), .IN2(n9861), .Q(n9860) );
  AND2X1 U9677 ( .IN1(n9829), .IN2(n9827), .Q(n9817) );
  AND2X1 U9678 ( .IN1(n9862), .IN2(n2361), .Q(n9824) );
  AND2X1 U9679 ( .IN1(n9816), .IN2(n7921), .Q(n9858) );
  AND2X1 U9680 ( .IN1(n9863), .IN2(n9827), .Q(n9816) );
  INVX0 U9681 ( .INP(n9864), .ZN(n9827) );
  OR2X1 U9682 ( .IN1(n9865), .IN2(n9866), .Q(n4250) );
  OR2X1 U9683 ( .IN1(n9867), .IN2(n9868), .Q(n9866) );
  AND2X1 U9684 ( .IN1(n9869), .IN2(g2584), .Q(n9868) );
  XOR2X1 U9685 ( .IN1(n9870), .IN2(n9871), .Q(n9869) );
  XOR2X1 U9686 ( .IN1(n9872), .IN2(n9873), .Q(n9871) );
  XOR2X1 U9687 ( .IN1(n9856), .IN2(n9861), .Q(n9873) );
  OR2X1 U9688 ( .IN1(n9874), .IN2(n9875), .Q(n9861) );
  OR2X1 U9689 ( .IN1(n9876), .IN2(n9877), .Q(n9875) );
  AND2X1 U9690 ( .IN1(n9878), .IN2(n9879), .Q(n9877) );
  AND2X1 U9691 ( .IN1(n9880), .IN2(n9881), .Q(n9876) );
  OR2X1 U9692 ( .IN1(n9882), .IN2(n9883), .Q(n9856) );
  OR2X1 U9693 ( .IN1(n9884), .IN2(n9885), .Q(n9883) );
  AND2X1 U9694 ( .IN1(n9886), .IN2(n9887), .Q(n9885) );
  AND2X1 U9695 ( .IN1(n9888), .IN2(n9889), .Q(n9884) );
  INVX0 U9696 ( .INP(n9887), .ZN(n9888) );
  XOR2X1 U9697 ( .IN1(n9845), .IN2(n9850), .Q(n9872) );
  OR2X1 U9698 ( .IN1(n9874), .IN2(n9890), .Q(n9850) );
  OR2X1 U9699 ( .IN1(n9891), .IN2(n9892), .Q(n9890) );
  AND2X1 U9700 ( .IN1(n9893), .IN2(n9879), .Q(n9892) );
  AND2X1 U9701 ( .IN1(n9880), .IN2(n9894), .Q(n9891) );
  OR2X1 U9702 ( .IN1(n9882), .IN2(n9895), .Q(n9845) );
  OR2X1 U9703 ( .IN1(n9896), .IN2(n9897), .Q(n9895) );
  AND2X1 U9704 ( .IN1(n9898), .IN2(n9879), .Q(n9897) );
  INVX0 U9705 ( .INP(n9899), .ZN(n9898) );
  AND2X1 U9706 ( .IN1(n9880), .IN2(n9899), .Q(n9896) );
  XOR2X1 U9707 ( .IN1(n9900), .IN2(n9901), .Q(n9870) );
  XOR2X1 U9708 ( .IN1(n9833), .IN2(n9839), .Q(n9901) );
  OR2X1 U9709 ( .IN1(n9882), .IN2(n9902), .Q(n9839) );
  OR2X1 U9710 ( .IN1(n9903), .IN2(n9904), .Q(n9902) );
  AND2X1 U9711 ( .IN1(n9905), .IN2(n9879), .Q(n9904) );
  INVX0 U9712 ( .INP(n9906), .ZN(n9905) );
  AND2X1 U9713 ( .IN1(n9880), .IN2(n9906), .Q(n9903) );
  OR2X1 U9714 ( .IN1(n9907), .IN2(n9908), .Q(n9833) );
  OR2X1 U9715 ( .IN1(n9909), .IN2(n9910), .Q(n9907) );
  AND2X1 U9716 ( .IN1(n9886), .IN2(n9911), .Q(n9910) );
  AND2X1 U9717 ( .IN1(n9912), .IN2(n9889), .Q(n9909) );
  XOR2X1 U9718 ( .IN1(n9818), .IN2(n9828), .Q(n9900) );
  OR2X1 U9719 ( .IN1(n9882), .IN2(n9913), .Q(n9828) );
  OR2X1 U9720 ( .IN1(n9914), .IN2(n9915), .Q(n9913) );
  AND2X1 U9721 ( .IN1(n9886), .IN2(n9916), .Q(n9915) );
  AND2X1 U9722 ( .IN1(n9917), .IN2(n9889), .Q(n9914) );
  OR2X1 U9723 ( .IN1(n9882), .IN2(n9918), .Q(n9818) );
  OR2X1 U9724 ( .IN1(n9919), .IN2(n9920), .Q(n9918) );
  AND2X1 U9725 ( .IN1(n9886), .IN2(n9921), .Q(n9920) );
  AND2X1 U9726 ( .IN1(n9922), .IN2(n9889), .Q(n9919) );
  INVX0 U9727 ( .INP(n9921), .ZN(n9922) );
  AND2X1 U9728 ( .IN1(n9923), .IN2(n9924), .Q(n9867) );
  AND2X1 U9729 ( .IN1(n9925), .IN2(n9926), .Q(n9924) );
  OR2X1 U9730 ( .IN1(g3229), .IN2(n7918), .Q(n9926) );
  INVX0 U9731 ( .INP(n9927), .ZN(n9925) );
  AND2X1 U9732 ( .IN1(g3229), .IN2(n4490), .Q(n9927) );
  INVX0 U9733 ( .INP(n9928), .ZN(n9923) );
  OR2X1 U9734 ( .IN1(n9829), .IN2(n9864), .Q(n9928) );
  OR2X1 U9735 ( .IN1(n9862), .IN2(n9929), .Q(n9829) );
  AND2X1 U9736 ( .IN1(n9930), .IN2(g2631), .Q(n9865) );
  XOR2X1 U9737 ( .IN1(n9819), .IN2(n9851), .Q(n9930) );
  OR2X1 U9738 ( .IN1(n9874), .IN2(n9931), .Q(n9851) );
  OR2X1 U9739 ( .IN1(n9932), .IN2(n9933), .Q(n9931) );
  AND2X1 U9740 ( .IN1(n9934), .IN2(n9879), .Q(n9933) );
  AND2X1 U9741 ( .IN1(n9880), .IN2(n9935), .Q(n9932) );
  AND2X1 U9742 ( .IN1(n9936), .IN2(n9937), .Q(n9880) );
  OR2X1 U9743 ( .IN1(n9938), .IN2(n9882), .Q(n9874) );
  INVX0 U9744 ( .INP(n9939), .ZN(n9938) );
  OR2X1 U9745 ( .IN1(n9936), .IN2(n9937), .Q(n9939) );
  OR2X1 U9746 ( .IN1(n9940), .IN2(n9908), .Q(n9819) );
  OR2X1 U9747 ( .IN1(n9941), .IN2(n9882), .Q(n9908) );
  OR2X1 U9748 ( .IN1(n4543), .IN2(n9862), .Q(n9882) );
  OR2X1 U9749 ( .IN1(g2633), .IN2(n9942), .Q(n9862) );
  OR2X1 U9750 ( .IN1(g2637), .IN2(g30072), .Q(n9942) );
  INVX0 U9751 ( .INP(n2381), .ZN(n9941) );
  OR2X1 U9752 ( .IN1(n9943), .IN2(n9944), .Q(n9940) );
  AND2X1 U9753 ( .IN1(n9886), .IN2(n9945), .Q(n9944) );
  AND2X1 U9754 ( .IN1(n9936), .IN2(n9946), .Q(n9886) );
  AND2X1 U9755 ( .IN1(n9947), .IN2(n9889), .Q(n9943) );
  OR2X1 U9756 ( .IN1(n9948), .IN2(n9949), .Q(n4249) );
  OR2X1 U9757 ( .IN1(n9950), .IN2(n9951), .Q(n9949) );
  AND2X1 U9758 ( .IN1(n9952), .IN2(g1917), .Q(n9951) );
  AND2X1 U9759 ( .IN1(n9953), .IN2(n9954), .Q(n9950) );
  AND2X1 U9760 ( .IN1(n2289), .IN2(n9955), .Q(n9948) );
  OR2X1 U9761 ( .IN1(n9956), .IN2(n9957), .Q(n4248) );
  OR2X1 U9762 ( .IN1(n9958), .IN2(n9959), .Q(n9956) );
  AND2X1 U9763 ( .IN1(n9952), .IN2(n7966), .Q(n9959) );
  AND2X1 U9764 ( .IN1(n9960), .IN2(n9961), .Q(n9958) );
  AND2X1 U9765 ( .IN1(n9962), .IN2(n9963), .Q(n9960) );
  OR2X1 U9766 ( .IN1(n9964), .IN2(n9965), .Q(n4247) );
  OR2X1 U9767 ( .IN1(n9966), .IN2(n9967), .Q(n9965) );
  AND2X1 U9768 ( .IN1(n9952), .IN2(n7962), .Q(n9967) );
  AND2X1 U9769 ( .IN1(n9953), .IN2(n9968), .Q(n9966) );
  OR2X1 U9770 ( .IN1(n9969), .IN2(n9957), .Q(n4246) );
  OR2X1 U9771 ( .IN1(n9964), .IN2(n9970), .Q(n9957) );
  INVX0 U9772 ( .INP(n2303), .ZN(n9970) );
  OR2X1 U9773 ( .IN1(n9971), .IN2(n9972), .Q(n9969) );
  AND2X1 U9774 ( .IN1(n9952), .IN2(n7965), .Q(n9972) );
  AND2X1 U9775 ( .IN1(n9973), .IN2(n9961), .Q(n9971) );
  AND2X1 U9776 ( .IN1(n9974), .IN2(n9963), .Q(n9973) );
  OR2X1 U9777 ( .IN1(n9975), .IN2(n9976), .Q(n4245) );
  OR2X1 U9778 ( .IN1(n9977), .IN2(n9978), .Q(n9976) );
  AND2X1 U9779 ( .IN1(n9952), .IN2(n7967), .Q(n9978) );
  AND2X1 U9780 ( .IN1(n9979), .IN2(n9961), .Q(n9977) );
  AND2X1 U9781 ( .IN1(n9980), .IN2(n9963), .Q(n9979) );
  OR2X1 U9782 ( .IN1(n9981), .IN2(n9982), .Q(n4244) );
  OR2X1 U9783 ( .IN1(n9983), .IN2(n9984), .Q(n9982) );
  AND2X1 U9784 ( .IN1(n9952), .IN2(g1916), .Q(n9984) );
  AND2X1 U9785 ( .IN1(n9953), .IN2(n9985), .Q(n9983) );
  AND2X1 U9786 ( .IN1(n2289), .IN2(n9986), .Q(n9981) );
  OR2X1 U9787 ( .IN1(n9975), .IN2(n9987), .Q(n4243) );
  OR2X1 U9788 ( .IN1(n9988), .IN2(n9989), .Q(n9987) );
  AND2X1 U9789 ( .IN1(n9952), .IN2(n7964), .Q(n9989) );
  AND2X1 U9790 ( .IN1(n9990), .IN2(n9961), .Q(n9988) );
  AND2X1 U9791 ( .IN1(n9991), .IN2(n9963), .Q(n9990) );
  OR2X1 U9792 ( .IN1(n9992), .IN2(n9964), .Q(n9975) );
  AND2X1 U9793 ( .IN1(n2289), .IN2(n2302), .Q(n9992) );
  OR2X1 U9794 ( .IN1(n9964), .IN2(n9993), .Q(n4242) );
  OR2X1 U9795 ( .IN1(n9994), .IN2(n9995), .Q(n9993) );
  AND2X1 U9796 ( .IN1(n9952), .IN2(n7963), .Q(n9995) );
  AND2X1 U9797 ( .IN1(n9996), .IN2(n9961), .Q(n9952) );
  AND2X1 U9798 ( .IN1(n9953), .IN2(n9997), .Q(n9994) );
  AND2X1 U9799 ( .IN1(n9963), .IN2(n9961), .Q(n9953) );
  INVX0 U9800 ( .INP(n9998), .ZN(n9961) );
  INVX0 U9801 ( .INP(n2275), .ZN(n9964) );
  OR2X1 U9802 ( .IN1(n9999), .IN2(n10000), .Q(n4241) );
  OR2X1 U9803 ( .IN1(n10001), .IN2(n10002), .Q(n10000) );
  AND2X1 U9804 ( .IN1(n10003), .IN2(g1890), .Q(n10002) );
  XOR2X1 U9805 ( .IN1(n10004), .IN2(n10005), .Q(n10003) );
  XOR2X1 U9806 ( .IN1(n10006), .IN2(n10007), .Q(n10005) );
  XOR2X1 U9807 ( .IN1(n9991), .IN2(n9997), .Q(n10007) );
  OR2X1 U9808 ( .IN1(n10008), .IN2(n10009), .Q(n9997) );
  OR2X1 U9809 ( .IN1(n10010), .IN2(n10011), .Q(n10009) );
  AND2X1 U9810 ( .IN1(n10012), .IN2(n10013), .Q(n10011) );
  AND2X1 U9811 ( .IN1(n10014), .IN2(n10015), .Q(n10010) );
  OR2X1 U9812 ( .IN1(n10016), .IN2(n10017), .Q(n9991) );
  OR2X1 U9813 ( .IN1(n10018), .IN2(n10019), .Q(n10017) );
  AND2X1 U9814 ( .IN1(n10020), .IN2(n10021), .Q(n10019) );
  AND2X1 U9815 ( .IN1(n10022), .IN2(n10023), .Q(n10018) );
  XOR2X1 U9816 ( .IN1(n9980), .IN2(n9985), .Q(n10006) );
  OR2X1 U9817 ( .IN1(n10008), .IN2(n10024), .Q(n9985) );
  OR2X1 U9818 ( .IN1(n10025), .IN2(n10026), .Q(n10024) );
  AND2X1 U9819 ( .IN1(n10027), .IN2(n10013), .Q(n10026) );
  AND2X1 U9820 ( .IN1(n10014), .IN2(n10028), .Q(n10025) );
  OR2X1 U9821 ( .IN1(n10016), .IN2(n10029), .Q(n9980) );
  OR2X1 U9822 ( .IN1(n10030), .IN2(n10031), .Q(n10029) );
  AND2X1 U9823 ( .IN1(n10032), .IN2(n10013), .Q(n10031) );
  INVX0 U9824 ( .INP(n10033), .ZN(n10032) );
  AND2X1 U9825 ( .IN1(n10014), .IN2(n10033), .Q(n10030) );
  XOR2X1 U9826 ( .IN1(n10034), .IN2(n10035), .Q(n10004) );
  XOR2X1 U9827 ( .IN1(n9968), .IN2(n9974), .Q(n10035) );
  OR2X1 U9828 ( .IN1(n10016), .IN2(n10036), .Q(n9974) );
  OR2X1 U9829 ( .IN1(n10037), .IN2(n10038), .Q(n10036) );
  AND2X1 U9830 ( .IN1(n10039), .IN2(n10013), .Q(n10038) );
  INVX0 U9831 ( .INP(n10040), .ZN(n10039) );
  AND2X1 U9832 ( .IN1(n10014), .IN2(n10040), .Q(n10037) );
  OR2X1 U9833 ( .IN1(n10041), .IN2(n10042), .Q(n9968) );
  OR2X1 U9834 ( .IN1(n10043), .IN2(n10044), .Q(n10041) );
  AND2X1 U9835 ( .IN1(n10020), .IN2(n10045), .Q(n10044) );
  AND2X1 U9836 ( .IN1(n10046), .IN2(n10023), .Q(n10043) );
  XOR2X1 U9837 ( .IN1(n9954), .IN2(n9962), .Q(n10034) );
  OR2X1 U9838 ( .IN1(n10016), .IN2(n10047), .Q(n9962) );
  OR2X1 U9839 ( .IN1(n10048), .IN2(n10049), .Q(n10047) );
  AND2X1 U9840 ( .IN1(n10020), .IN2(n10050), .Q(n10049) );
  AND2X1 U9841 ( .IN1(n10051), .IN2(n10023), .Q(n10048) );
  INVX0 U9842 ( .INP(n10050), .ZN(n10051) );
  OR2X1 U9843 ( .IN1(n10016), .IN2(n10052), .Q(n9954) );
  OR2X1 U9844 ( .IN1(n10053), .IN2(n10054), .Q(n10052) );
  AND2X1 U9845 ( .IN1(n10020), .IN2(n10055), .Q(n10054) );
  AND2X1 U9846 ( .IN1(n10056), .IN2(n10023), .Q(n10053) );
  INVX0 U9847 ( .INP(n10055), .ZN(n10056) );
  AND2X1 U9848 ( .IN1(n10057), .IN2(n10058), .Q(n10001) );
  AND2X1 U9849 ( .IN1(n10059), .IN2(n10060), .Q(n10058) );
  OR2X1 U9850 ( .IN1(test_so69), .IN2(n10061), .Q(n10060) );
  OR2X1 U9851 ( .IN1(g3229), .IN2(n7960), .Q(n10059) );
  INVX0 U9852 ( .INP(n10062), .ZN(n10057) );
  OR2X1 U9853 ( .IN1(n9963), .IN2(n9998), .Q(n10062) );
  OR2X1 U9854 ( .IN1(n10063), .IN2(n9516), .Q(n9963) );
  AND2X1 U9855 ( .IN1(n10064), .IN2(g1937), .Q(n9999) );
  XOR2X1 U9856 ( .IN1(n9955), .IN2(n9986), .Q(n10064) );
  OR2X1 U9857 ( .IN1(n10008), .IN2(n10065), .Q(n9986) );
  OR2X1 U9858 ( .IN1(n10066), .IN2(n10067), .Q(n10065) );
  AND2X1 U9859 ( .IN1(n10068), .IN2(n10013), .Q(n10067) );
  AND2X1 U9860 ( .IN1(n10014), .IN2(n10069), .Q(n10066) );
  AND2X1 U9861 ( .IN1(n10070), .IN2(n10071), .Q(n10014) );
  OR2X1 U9862 ( .IN1(n10072), .IN2(n10016), .Q(n10008) );
  INVX0 U9863 ( .INP(n2279), .ZN(n10072) );
  OR2X1 U9864 ( .IN1(n10073), .IN2(n10042), .Q(n9955) );
  OR2X1 U9865 ( .IN1(n10074), .IN2(n10016), .Q(n10042) );
  OR2X1 U9866 ( .IN1(n4545), .IN2(n9516), .Q(n10016) );
  OR2X1 U9867 ( .IN1(g1939), .IN2(n10075), .Q(n9516) );
  OR2X1 U9868 ( .IN1(g1943), .IN2(n490), .Q(n10075) );
  INVX0 U9869 ( .INP(n2309), .ZN(n10074) );
  OR2X1 U9870 ( .IN1(n10076), .IN2(n10077), .Q(n10073) );
  AND2X1 U9871 ( .IN1(n10020), .IN2(n10078), .Q(n10077) );
  AND2X1 U9872 ( .IN1(n10070), .IN2(n10079), .Q(n10020) );
  AND2X1 U9873 ( .IN1(n10080), .IN2(n10023), .Q(n10076) );
  OR2X1 U9874 ( .IN1(n10081), .IN2(n10082), .Q(n4240) );
  OR2X1 U9875 ( .IN1(n10083), .IN2(n10084), .Q(n10082) );
  AND2X1 U9876 ( .IN1(n10085), .IN2(g1223), .Q(n10084) );
  AND2X1 U9877 ( .IN1(n10086), .IN2(n10087), .Q(n10083) );
  AND2X1 U9878 ( .IN1(n2217), .IN2(n10088), .Q(n10081) );
  OR2X1 U9879 ( .IN1(n10089), .IN2(n10090), .Q(n4239) );
  OR2X1 U9880 ( .IN1(n10091), .IN2(n10092), .Q(n10090) );
  AND2X1 U9881 ( .IN1(n10085), .IN2(n8007), .Q(n10091) );
  OR2X1 U9882 ( .IN1(n10093), .IN2(n10094), .Q(n10089) );
  AND2X1 U9883 ( .IN1(n10095), .IN2(n10096), .Q(n10094) );
  AND2X1 U9884 ( .IN1(n10097), .IN2(n10098), .Q(n10095) );
  OR2X1 U9885 ( .IN1(n10099), .IN2(n10100), .Q(n4238) );
  OR2X1 U9886 ( .IN1(n10093), .IN2(n10101), .Q(n10100) );
  AND2X1 U9887 ( .IN1(n10086), .IN2(n10102), .Q(n10101) );
  AND2X1 U9888 ( .IN1(n10085), .IN2(n8003), .Q(n10099) );
  OR2X1 U9889 ( .IN1(n10103), .IN2(n10104), .Q(n4237) );
  OR2X1 U9890 ( .IN1(n10105), .IN2(n10092), .Q(n10104) );
  INVX0 U9891 ( .INP(n2231), .ZN(n10092) );
  AND2X1 U9892 ( .IN1(n10085), .IN2(n8006), .Q(n10105) );
  OR2X1 U9893 ( .IN1(n10093), .IN2(n10106), .Q(n10103) );
  AND2X1 U9894 ( .IN1(n10107), .IN2(n10096), .Q(n10106) );
  AND2X1 U9895 ( .IN1(n10108), .IN2(n10098), .Q(n10107) );
  OR2X1 U9896 ( .IN1(n10109), .IN2(n10110), .Q(n4236) );
  OR2X1 U9897 ( .IN1(n10111), .IN2(n10112), .Q(n10110) );
  AND2X1 U9898 ( .IN1(n10085), .IN2(n8008), .Q(n10112) );
  AND2X1 U9899 ( .IN1(n10113), .IN2(n10096), .Q(n10111) );
  AND2X1 U9900 ( .IN1(n10114), .IN2(n10098), .Q(n10113) );
  OR2X1 U9901 ( .IN1(n10115), .IN2(n10116), .Q(n4235) );
  OR2X1 U9902 ( .IN1(n10117), .IN2(n10118), .Q(n10116) );
  AND2X1 U9903 ( .IN1(n10085), .IN2(g1222), .Q(n10118) );
  AND2X1 U9904 ( .IN1(n10086), .IN2(n10119), .Q(n10117) );
  AND2X1 U9905 ( .IN1(n2217), .IN2(n10120), .Q(n10115) );
  OR2X1 U9906 ( .IN1(n10109), .IN2(n10121), .Q(n4234) );
  OR2X1 U9907 ( .IN1(n10122), .IN2(n10123), .Q(n10121) );
  AND2X1 U9908 ( .IN1(n10085), .IN2(n8005), .Q(n10123) );
  AND2X1 U9909 ( .IN1(n10124), .IN2(n10096), .Q(n10122) );
  AND2X1 U9910 ( .IN1(n10125), .IN2(n10098), .Q(n10124) );
  OR2X1 U9911 ( .IN1(n10093), .IN2(n10126), .Q(n10109) );
  AND2X1 U9912 ( .IN1(n2217), .IN2(n2230), .Q(n10126) );
  OR2X1 U9913 ( .IN1(n10127), .IN2(n10128), .Q(n4233) );
  OR2X1 U9914 ( .IN1(n10093), .IN2(n10129), .Q(n10128) );
  AND2X1 U9915 ( .IN1(n10086), .IN2(n10130), .Q(n10129) );
  AND2X1 U9916 ( .IN1(n10098), .IN2(n10096), .Q(n10086) );
  AND2X1 U9917 ( .IN1(n10131), .IN2(n2217), .Q(n10093) );
  AND2X1 U9918 ( .IN1(n10085), .IN2(n8004), .Q(n10127) );
  AND2X1 U9919 ( .IN1(n10132), .IN2(n10096), .Q(n10085) );
  INVX0 U9920 ( .INP(n10133), .ZN(n10096) );
  OR2X1 U9921 ( .IN1(n10134), .IN2(n10135), .Q(n4232) );
  OR2X1 U9922 ( .IN1(n10136), .IN2(n10137), .Q(n10135) );
  AND2X1 U9923 ( .IN1(n10138), .IN2(g1196), .Q(n10137) );
  XOR2X1 U9924 ( .IN1(n10139), .IN2(n10140), .Q(n10138) );
  XOR2X1 U9925 ( .IN1(n10141), .IN2(n10142), .Q(n10140) );
  XOR2X1 U9926 ( .IN1(n10125), .IN2(n10130), .Q(n10142) );
  OR2X1 U9927 ( .IN1(n10143), .IN2(n10144), .Q(n10130) );
  OR2X1 U9928 ( .IN1(n10145), .IN2(n10146), .Q(n10144) );
  AND2X1 U9929 ( .IN1(n10147), .IN2(n10148), .Q(n10146) );
  AND2X1 U9930 ( .IN1(n10149), .IN2(n10150), .Q(n10145) );
  OR2X1 U9931 ( .IN1(n10151), .IN2(n10152), .Q(n10125) );
  OR2X1 U9932 ( .IN1(n10153), .IN2(n10154), .Q(n10152) );
  AND2X1 U9933 ( .IN1(n10155), .IN2(n10156), .Q(n10154) );
  AND2X1 U9934 ( .IN1(n10157), .IN2(n10158), .Q(n10153) );
  INVX0 U9935 ( .INP(n10156), .ZN(n10157) );
  XOR2X1 U9936 ( .IN1(n10114), .IN2(n10119), .Q(n10141) );
  OR2X1 U9937 ( .IN1(n10143), .IN2(n10159), .Q(n10119) );
  OR2X1 U9938 ( .IN1(n10160), .IN2(n10161), .Q(n10159) );
  AND2X1 U9939 ( .IN1(n10162), .IN2(n10148), .Q(n10161) );
  AND2X1 U9940 ( .IN1(n10149), .IN2(n10163), .Q(n10160) );
  OR2X1 U9941 ( .IN1(n10151), .IN2(n10164), .Q(n10114) );
  OR2X1 U9942 ( .IN1(n10165), .IN2(n10166), .Q(n10164) );
  AND2X1 U9943 ( .IN1(n10167), .IN2(n10148), .Q(n10166) );
  INVX0 U9944 ( .INP(n10168), .ZN(n10167) );
  AND2X1 U9945 ( .IN1(n10149), .IN2(n10168), .Q(n10165) );
  XOR2X1 U9946 ( .IN1(n10169), .IN2(n10170), .Q(n10139) );
  XOR2X1 U9947 ( .IN1(n10102), .IN2(n10108), .Q(n10170) );
  OR2X1 U9948 ( .IN1(n10151), .IN2(n10171), .Q(n10108) );
  OR2X1 U9949 ( .IN1(n10172), .IN2(n10173), .Q(n10171) );
  AND2X1 U9950 ( .IN1(n10174), .IN2(n10148), .Q(n10173) );
  AND2X1 U9951 ( .IN1(n10149), .IN2(n10175), .Q(n10172) );
  OR2X1 U9952 ( .IN1(n10176), .IN2(n10177), .Q(n10102) );
  OR2X1 U9953 ( .IN1(n10178), .IN2(n10179), .Q(n10176) );
  AND2X1 U9954 ( .IN1(n10155), .IN2(n10180), .Q(n10179) );
  AND2X1 U9955 ( .IN1(n10181), .IN2(n10158), .Q(n10178) );
  XOR2X1 U9956 ( .IN1(n10087), .IN2(n10097), .Q(n10169) );
  OR2X1 U9957 ( .IN1(n10151), .IN2(n10182), .Q(n10097) );
  OR2X1 U9958 ( .IN1(n10183), .IN2(n10184), .Q(n10182) );
  AND2X1 U9959 ( .IN1(n10155), .IN2(n10185), .Q(n10184) );
  AND2X1 U9960 ( .IN1(n10186), .IN2(n10158), .Q(n10183) );
  INVX0 U9961 ( .INP(n10185), .ZN(n10186) );
  OR2X1 U9962 ( .IN1(n10151), .IN2(n10187), .Q(n10087) );
  OR2X1 U9963 ( .IN1(n10188), .IN2(n10189), .Q(n10187) );
  AND2X1 U9964 ( .IN1(n10155), .IN2(n10190), .Q(n10189) );
  AND2X1 U9965 ( .IN1(n10191), .IN2(n10158), .Q(n10188) );
  INVX0 U9966 ( .INP(n10190), .ZN(n10191) );
  AND2X1 U9967 ( .IN1(n10192), .IN2(n10193), .Q(n10136) );
  AND2X1 U9968 ( .IN1(n10194), .IN2(n10195), .Q(n10193) );
  INVX0 U9969 ( .INP(n10196), .ZN(n10195) );
  AND2X1 U9970 ( .IN1(g3229), .IN2(n4489), .Q(n10196) );
  OR2X1 U9971 ( .IN1(test_so48), .IN2(g3229), .Q(n10194) );
  INVX0 U9972 ( .INP(n10197), .ZN(n10192) );
  OR2X1 U9973 ( .IN1(n10098), .IN2(n10133), .Q(n10197) );
  OR2X1 U9974 ( .IN1(n10131), .IN2(n10198), .Q(n10098) );
  AND2X1 U9975 ( .IN1(n10199), .IN2(g1243), .Q(n10134) );
  XOR2X1 U9976 ( .IN1(n10088), .IN2(n10120), .Q(n10199) );
  OR2X1 U9977 ( .IN1(n10143), .IN2(n10200), .Q(n10120) );
  OR2X1 U9978 ( .IN1(n10201), .IN2(n10202), .Q(n10200) );
  AND2X1 U9979 ( .IN1(n10203), .IN2(n10148), .Q(n10202) );
  AND2X1 U9980 ( .IN1(n10149), .IN2(n10204), .Q(n10201) );
  AND2X1 U9981 ( .IN1(n10205), .IN2(n10206), .Q(n10149) );
  OR2X1 U9982 ( .IN1(n10207), .IN2(n10151), .Q(n10143) );
  INVX0 U9983 ( .INP(n2207), .ZN(n10207) );
  OR2X1 U9984 ( .IN1(n10208), .IN2(n10177), .Q(n10088) );
  OR2X1 U9985 ( .IN1(n10209), .IN2(n10151), .Q(n10177) );
  OR2X1 U9986 ( .IN1(n4548), .IN2(n10131), .Q(n10151) );
  OR2X1 U9987 ( .IN1(g1245), .IN2(n10210), .Q(n10131) );
  OR2X1 U9988 ( .IN1(g1249), .IN2(n486), .Q(n10210) );
  INVX0 U9989 ( .INP(n2237), .ZN(n10209) );
  OR2X1 U9990 ( .IN1(n10211), .IN2(n10212), .Q(n10208) );
  AND2X1 U9991 ( .IN1(n10155), .IN2(n10213), .Q(n10212) );
  AND2X1 U9992 ( .IN1(n10205), .IN2(n10214), .Q(n10155) );
  AND2X1 U9993 ( .IN1(n10215), .IN2(n10158), .Q(n10211) );
  INVX0 U9994 ( .INP(n10216), .ZN(n4521) );
  AND2X1 U9995 ( .IN1(test_so15), .IN2(n3692), .Q(n10216) );
  OR2X1 U9996 ( .IN1(n9113), .IN2(n10217), .Q(n4528) );
  OR2X1 U9997 ( .IN1(n9114), .IN2(n10218), .Q(n4527) );
  OR2X1 U9998 ( .IN1(n9115), .IN2(n10219), .Q(n4523) );
  OR2X1 U9999 ( .IN1(n9116), .IN2(n10220), .Q(n4522) );
  INVX0 U10000 ( .INP(n10221), .ZN(n338) );
  OR2X1 U10001 ( .IN1(n10222), .IN2(n10223), .Q(n3254) );
  INVX0 U10002 ( .INP(n10224), .ZN(n10223) );
  OR2X1 U10003 ( .IN1(n10225), .IN2(n10226), .Q(n10224) );
  INVX0 U10004 ( .INP(g24734), .ZN(n312) );
  INVX0 U10005 ( .INP(g25435), .ZN(n308) );
  INVX0 U10006 ( .INP(g26135), .ZN(n282) );
  OR2X1 U10007 ( .IN1(n10227), .IN2(n10228), .Q(n2800) );
  AND2X1 U10008 ( .IN1(n10229), .IN2(n10230), .Q(n10228) );
  AND2X1 U10009 ( .IN1(n10231), .IN2(n10232), .Q(n10229) );
  INVX0 U10010 ( .INP(n10233), .ZN(n10227) );
  OR2X1 U10011 ( .IN1(n10231), .IN2(n10230), .Q(n10233) );
  OR2X1 U10012 ( .IN1(n10234), .IN2(n10235), .Q(n10231) );
  OR2X1 U10013 ( .IN1(n10236), .IN2(n10237), .Q(n10235) );
  AND2X1 U10014 ( .IN1(n10238), .IN2(n10239), .Q(n10237) );
  OR2X1 U10015 ( .IN1(n10240), .IN2(n10241), .Q(n10234) );
  AND2X1 U10016 ( .IN1(n10242), .IN2(n10243), .Q(n10241) );
  AND2X1 U10017 ( .IN1(n10244), .IN2(n10245), .Q(n10242) );
  OR2X1 U10018 ( .IN1(n10246), .IN2(n10247), .Q(n10244) );
  AND2X1 U10019 ( .IN1(n10230), .IN2(n10248), .Q(n10246) );
  AND2X1 U10020 ( .IN1(n10249), .IN2(n10250), .Q(n10240) );
  OR2X1 U10021 ( .IN1(n4387), .IN2(n10251), .Q(n10250) );
  XNOR2X1 U10022 ( .IN1(n9540), .IN2(n10252), .Q(n2719) );
  XNOR2X1 U10023 ( .IN1(n9618), .IN2(n4530), .Q(n2686) );
  XNOR2X1 U10024 ( .IN1(n9643), .IN2(n4529), .Q(n2671) );
  INVX0 U10025 ( .INP(n10253), .ZN(n2617) );
  XNOR2X1 U10026 ( .IN1(n10249), .IN2(n10254), .Q(n2616) );
  OR2X1 U10027 ( .IN1(n10255), .IN2(n10256), .Q(n10254) );
  OR2X1 U10028 ( .IN1(n10257), .IN2(n10258), .Q(n10256) );
  AND2X1 U10029 ( .IN1(n10259), .IN2(n10249), .Q(n10258) );
  AND2X1 U10030 ( .IN1(n10260), .IN2(n10245), .Q(n10259) );
  AND2X1 U10031 ( .IN1(n10261), .IN2(n10262), .Q(n10260) );
  OR2X1 U10032 ( .IN1(n10230), .IN2(n10263), .Q(n10262) );
  OR2X1 U10033 ( .IN1(n10264), .IN2(n10239), .Q(n10261) );
  AND2X1 U10034 ( .IN1(n10265), .IN2(n10266), .Q(n10264) );
  AND2X1 U10035 ( .IN1(n10267), .IN2(n10232), .Q(n10266) );
  AND2X1 U10036 ( .IN1(n10268), .IN2(n10269), .Q(n10265) );
  OR2X1 U10037 ( .IN1(n10247), .IN2(n10248), .Q(n10269) );
  INVX0 U10038 ( .INP(n10270), .ZN(n10248) );
  AND2X1 U10039 ( .IN1(n10271), .IN2(n10243), .Q(n10257) );
  OR2X1 U10040 ( .IN1(n10272), .IN2(n10247), .Q(n10271) );
  AND2X1 U10041 ( .IN1(n10273), .IN2(n10274), .Q(n10272) );
  INVX0 U10042 ( .INP(n10275), .ZN(n10274) );
  AND2X1 U10043 ( .IN1(n10276), .IN2(n10277), .Q(n10273) );
  INVX0 U10044 ( .INP(n10278), .ZN(n10277) );
  OR2X1 U10045 ( .IN1(n10239), .IN2(n10279), .Q(n10276) );
  OR2X1 U10046 ( .IN1(n10270), .IN2(n10280), .Q(n10279) );
  AND2X1 U10047 ( .IN1(n10236), .IN2(n10281), .Q(n10255) );
  OR2X1 U10048 ( .IN1(n9798), .IN2(n9797), .Q(n2459) );
  AND2X1 U10049 ( .IN1(n9716), .IN2(n9714), .Q(n2446) );
  INVX0 U10050 ( .INP(n9753), .ZN(n9714) );
  OR2X1 U10051 ( .IN1(test_so22), .IN2(n10282), .Q(n9753) );
  AND2X1 U10052 ( .IN1(n8828), .IN2(n4360), .Q(n10282) );
  OR2X1 U10053 ( .IN1(n10283), .IN2(g557), .Q(n9716) );
  AND2X1 U10054 ( .IN1(n8828), .IN2(n9126), .Q(n10283) );
  OR2X1 U10055 ( .IN1(n10284), .IN2(n4541), .Q(n2445) );
  AND2X1 U10056 ( .IN1(n10285), .IN2(n10286), .Q(n10284) );
  AND2X1 U10057 ( .IN1(n10287), .IN2(n9797), .Q(n10286) );
  OR2X1 U10058 ( .IN1(n10288), .IN2(n10289), .Q(n9797) );
  OR2X1 U10059 ( .IN1(n10290), .IN2(n10291), .Q(n10289) );
  OR2X1 U10060 ( .IN1(n9791), .IN2(n10292), .Q(n10291) );
  OR2X1 U10061 ( .IN1(n9763), .IN2(n9785), .Q(n10292) );
  OR2X1 U10062 ( .IN1(n9779), .IN2(n10293), .Q(n10290) );
  OR2X1 U10063 ( .IN1(n10294), .IN2(n9773), .Q(n10293) );
  AND2X1 U10064 ( .IN1(n10295), .IN2(n10296), .Q(n10294) );
  OR2X1 U10065 ( .IN1(n4295), .IN2(g737), .Q(n10296) );
  AND2X1 U10066 ( .IN1(n10297), .IN2(n10298), .Q(n10295) );
  OR2X1 U10067 ( .IN1(n4359), .IN2(g739), .Q(n10298) );
  OR2X1 U10068 ( .IN1(n4309), .IN2(g738), .Q(n10297) );
  OR2X1 U10069 ( .IN1(n10299), .IN2(n10300), .Q(n10288) );
  OR2X1 U10070 ( .IN1(n10301), .IN2(n10302), .Q(n10300) );
  OR2X1 U10071 ( .IN1(n9743), .IN2(n9737), .Q(n10302) );
  INVX0 U10072 ( .INP(n10303), .ZN(n10301) );
  OR2X1 U10073 ( .IN1(n9768), .IN2(n10304), .Q(n10299) );
  OR2X1 U10074 ( .IN1(n9799), .IN2(n9803), .Q(n10304) );
  OR2X1 U10075 ( .IN1(n4359), .IN2(g736), .Q(n10287) );
  AND2X1 U10076 ( .IN1(n10305), .IN2(n10306), .Q(n10285) );
  OR2X1 U10077 ( .IN1(n4309), .IN2(g735), .Q(n10306) );
  OR2X1 U10078 ( .IN1(n4295), .IN2(g734), .Q(n10305) );
  OR2X1 U10079 ( .IN1(n9946), .IN2(n9936), .Q(n2381) );
  OR2X1 U10080 ( .IN1(n10307), .IN2(n4543), .Q(n2374) );
  AND2X1 U10081 ( .IN1(n10308), .IN2(n10309), .Q(n10307) );
  AND2X1 U10082 ( .IN1(n10310), .IN2(n9936), .Q(n10309) );
  OR2X1 U10083 ( .IN1(n10311), .IN2(n10312), .Q(n9936) );
  OR2X1 U10084 ( .IN1(n10313), .IN2(n10314), .Q(n10312) );
  OR2X1 U10085 ( .IN1(n9921), .IN2(n10315), .Q(n10314) );
  OR2X1 U10086 ( .IN1(n9887), .IN2(n9899), .Q(n10315) );
  OR2X1 U10087 ( .IN1(n9906), .IN2(n10316), .Q(n10313) );
  OR2X1 U10088 ( .IN1(n10317), .IN2(n9916), .Q(n10316) );
  AND2X1 U10089 ( .IN1(n10318), .IN2(n10319), .Q(n10317) );
  OR2X1 U10090 ( .IN1(n4292), .IN2(test_so95), .Q(n10319) );
  AND2X1 U10091 ( .IN1(n10320), .IN2(n10321), .Q(n10318) );
  OR2X1 U10092 ( .IN1(n4356), .IN2(g2813), .Q(n10321) );
  OR2X1 U10093 ( .IN1(n4306), .IN2(g2812), .Q(n10320) );
  OR2X1 U10094 ( .IN1(n10322), .IN2(n10323), .Q(n10311) );
  OR2X1 U10095 ( .IN1(n10324), .IN2(n10325), .Q(n10323) );
  OR2X1 U10096 ( .IN1(n9934), .IN2(n9947), .Q(n10325) );
  INVX0 U10097 ( .INP(n10326), .ZN(n10324) );
  OR2X1 U10098 ( .IN1(n9878), .IN2(n10327), .Q(n10322) );
  OR2X1 U10099 ( .IN1(n9912), .IN2(n9893), .Q(n10327) );
  OR2X1 U10100 ( .IN1(n4356), .IN2(g2810), .Q(n10310) );
  AND2X1 U10101 ( .IN1(n10328), .IN2(n10329), .Q(n10308) );
  OR2X1 U10102 ( .IN1(n4306), .IN2(g2809), .Q(n10329) );
  OR2X1 U10103 ( .IN1(n4292), .IN2(g2808), .Q(n10328) );
  AND2X1 U10104 ( .IN1(n9864), .IN2(n9863), .Q(n2361) );
  INVX0 U10105 ( .INP(n9929), .ZN(n9863) );
  OR2X1 U10106 ( .IN1(n10330), .IN2(g2584), .Q(n9929) );
  AND2X1 U10107 ( .IN1(n4352), .IN2(n8825), .Q(n10330) );
  OR2X1 U10108 ( .IN1(n10331), .IN2(g2631), .Q(n9864) );
  AND2X1 U10109 ( .IN1(n8825), .IN2(n4303), .Q(n10331) );
  OR2X1 U10110 ( .IN1(n10079), .IN2(n10070), .Q(n2309) );
  OR2X1 U10111 ( .IN1(n10332), .IN2(n4545), .Q(n2302) );
  AND2X1 U10112 ( .IN1(n10333), .IN2(n10334), .Q(n10332) );
  AND2X1 U10113 ( .IN1(n10335), .IN2(n10070), .Q(n10334) );
  OR2X1 U10114 ( .IN1(n4357), .IN2(g2116), .Q(n10335) );
  AND2X1 U10115 ( .IN1(n10336), .IN2(n10337), .Q(n10333) );
  OR2X1 U10116 ( .IN1(n4307), .IN2(g2115), .Q(n10337) );
  OR2X1 U10117 ( .IN1(n4293), .IN2(g2114), .Q(n10336) );
  AND2X1 U10118 ( .IN1(n9998), .IN2(n9996), .Q(n2289) );
  INVX0 U10119 ( .INP(n10063), .ZN(n9996) );
  OR2X1 U10120 ( .IN1(n10338), .IN2(g1890), .Q(n10063) );
  AND2X1 U10121 ( .IN1(n8826), .IN2(n4311), .Q(n10338) );
  OR2X1 U10122 ( .IN1(n10339), .IN2(g1937), .Q(n9998) );
  AND2X1 U10123 ( .IN1(n4297), .IN2(n8826), .Q(n10339) );
  OR2X1 U10124 ( .IN1(n10071), .IN2(n10070), .Q(n2279) );
  OR2X1 U10125 ( .IN1(n10340), .IN2(n10341), .Q(n10070) );
  OR2X1 U10126 ( .IN1(n10342), .IN2(n10343), .Q(n10341) );
  OR2X1 U10127 ( .IN1(n10055), .IN2(n10344), .Q(n10343) );
  OR2X1 U10128 ( .IN1(n10033), .IN2(n10021), .Q(n10344) );
  INVX0 U10129 ( .INP(n10022), .ZN(n10021) );
  OR2X1 U10130 ( .IN1(n10050), .IN2(n10345), .Q(n10342) );
  OR2X1 U10131 ( .IN1(n10346), .IN2(n10040), .Q(n10345) );
  AND2X1 U10132 ( .IN1(n10347), .IN2(n10348), .Q(n10346) );
  OR2X1 U10133 ( .IN1(n4293), .IN2(g2117), .Q(n10348) );
  AND2X1 U10134 ( .IN1(n10349), .IN2(n10350), .Q(n10347) );
  OR2X1 U10135 ( .IN1(n4357), .IN2(g2119), .Q(n10350) );
  OR2X1 U10136 ( .IN1(n4307), .IN2(g2118), .Q(n10349) );
  OR2X1 U10137 ( .IN1(n10351), .IN2(n10352), .Q(n10340) );
  OR2X1 U10138 ( .IN1(n10353), .IN2(n10354), .Q(n10352) );
  OR2X1 U10139 ( .IN1(n10068), .IN2(n10080), .Q(n10354) );
  INVX0 U10140 ( .INP(n10355), .ZN(n10353) );
  OR2X1 U10141 ( .IN1(n10012), .IN2(n10356), .Q(n10351) );
  OR2X1 U10142 ( .IN1(n10046), .IN2(n10027), .Q(n10356) );
  OR2X1 U10143 ( .IN1(n10214), .IN2(n10205), .Q(n2237) );
  OR2X1 U10144 ( .IN1(n10357), .IN2(n4548), .Q(n2230) );
  AND2X1 U10145 ( .IN1(n10358), .IN2(n10359), .Q(n10357) );
  AND2X1 U10146 ( .IN1(n10360), .IN2(n10205), .Q(n10359) );
  OR2X1 U10147 ( .IN1(n4358), .IN2(g1422), .Q(n10360) );
  AND2X1 U10148 ( .IN1(n10361), .IN2(n10362), .Q(n10358) );
  OR2X1 U10149 ( .IN1(n4308), .IN2(g1421), .Q(n10362) );
  OR2X1 U10150 ( .IN1(n4294), .IN2(g1420), .Q(n10361) );
  AND2X1 U10151 ( .IN1(n10133), .IN2(n10132), .Q(n2217) );
  INVX0 U10152 ( .INP(n10198), .ZN(n10132) );
  OR2X1 U10153 ( .IN1(n10363), .IN2(g1196), .Q(n10198) );
  AND2X1 U10154 ( .IN1(n4353), .IN2(n8827), .Q(n10363) );
  OR2X1 U10155 ( .IN1(n10364), .IN2(g1243), .Q(n10133) );
  AND2X1 U10156 ( .IN1(n8827), .IN2(n4304), .Q(n10364) );
  OR2X1 U10157 ( .IN1(n10206), .IN2(n10205), .Q(n2207) );
  OR2X1 U10158 ( .IN1(n10365), .IN2(n10366), .Q(n10205) );
  OR2X1 U10159 ( .IN1(n10367), .IN2(n10368), .Q(n10366) );
  OR2X1 U10160 ( .IN1(n10190), .IN2(n10369), .Q(n10368) );
  OR2X1 U10161 ( .IN1(n10168), .IN2(n10156), .Q(n10369) );
  OR2X1 U10162 ( .IN1(n10185), .IN2(n10370), .Q(n10367) );
  OR2X1 U10163 ( .IN1(n10371), .IN2(n10175), .Q(n10370) );
  INVX0 U10164 ( .INP(n10174), .ZN(n10175) );
  AND2X1 U10165 ( .IN1(n10372), .IN2(n10373), .Q(n10371) );
  OR2X1 U10166 ( .IN1(n4294), .IN2(g1423), .Q(n10373) );
  AND2X1 U10167 ( .IN1(n10374), .IN2(n10375), .Q(n10372) );
  OR2X1 U10168 ( .IN1(n4358), .IN2(g1425), .Q(n10375) );
  OR2X1 U10169 ( .IN1(n4308), .IN2(g1424), .Q(n10374) );
  OR2X1 U10170 ( .IN1(n10376), .IN2(n10377), .Q(n10365) );
  OR2X1 U10171 ( .IN1(n10378), .IN2(n10379), .Q(n10377) );
  OR2X1 U10172 ( .IN1(n10215), .IN2(n10203), .Q(n10379) );
  INVX0 U10173 ( .INP(n10380), .ZN(n10378) );
  OR2X1 U10174 ( .IN1(n10147), .IN2(n10381), .Q(n10376) );
  OR2X1 U10175 ( .IN1(n10181), .IN2(n10162), .Q(n10381) );
  INVX0 U10176 ( .INP(n10382), .ZN(n1386) );
  INVX0 U10177 ( .INP(n10383), .ZN(n1359) );
  INVX0 U10178 ( .INP(n10384), .ZN(n1348) );
  INVX0 U10179 ( .INP(n10385), .ZN(n4526) );
  AND2X1 U10180 ( .IN1(test_so78), .IN2(n3887), .Q(n10385) );
  INVX0 U10181 ( .INP(n10386), .ZN(n1221) );
  INVX0 U10182 ( .INP(g27380), .ZN(n122) );
  INVX0 U10183 ( .INP(n10387), .ZN(n1096) );
  INVX0 U10184 ( .INP(n10388), .ZN(n1073) );
  OR2X1 U10185 ( .IN1(n10389), .IN2(n10390), .Q(g30801) );
  AND2X1 U10186 ( .IN1(g30072), .IN2(g3109), .Q(n10390) );
  AND2X1 U10187 ( .IN1(n4494), .IN2(g3108), .Q(n10389) );
  OR2X1 U10188 ( .IN1(n10391), .IN2(n10392), .Q(g30798) );
  AND2X1 U10189 ( .IN1(g30072), .IN2(g8030), .Q(n10392) );
  AND2X1 U10190 ( .IN1(n4383), .IN2(g3107), .Q(n10391) );
  OR2X1 U10191 ( .IN1(n10393), .IN2(n10394), .Q(g30796) );
  AND2X1 U10192 ( .IN1(g30072), .IN2(g8106), .Q(n10394) );
  AND2X1 U10193 ( .IN1(n4382), .IN2(g3106), .Q(n10393) );
  OR2X1 U10194 ( .IN1(n10395), .IN2(n10396), .Q(g30709) );
  INVX0 U10195 ( .INP(n10397), .ZN(n10396) );
  OR2X1 U10196 ( .IN1(n10398), .IN2(n8375), .Q(n10397) );
  AND2X1 U10197 ( .IN1(n10399), .IN2(g7264), .Q(n10395) );
  OR2X1 U10198 ( .IN1(n10400), .IN2(n10401), .Q(g30708) );
  INVX0 U10199 ( .INP(n10402), .ZN(n10401) );
  OR2X1 U10200 ( .IN1(n10403), .IN2(n8391), .Q(n10402) );
  AND2X1 U10201 ( .IN1(n10404), .IN2(n4618), .Q(n10400) );
  OR2X1 U10202 ( .IN1(n10405), .IN2(n10406), .Q(g30707) );
  INVX0 U10203 ( .INP(n10407), .ZN(n10406) );
  OR2X1 U10204 ( .IN1(n10408), .IN2(n8386), .Q(n10407) );
  AND2X1 U10205 ( .IN1(n10399), .IN2(g5555), .Q(n10405) );
  OR2X1 U10206 ( .IN1(n10409), .IN2(n10410), .Q(g30706) );
  INVX0 U10207 ( .INP(n10411), .ZN(n10410) );
  OR2X1 U10208 ( .IN1(n10412), .IN2(n8378), .Q(n10411) );
  AND2X1 U10209 ( .IN1(n10404), .IN2(g7014), .Q(n10409) );
  OR2X1 U10210 ( .IN1(n10413), .IN2(n10414), .Q(g30705) );
  AND2X1 U10211 ( .IN1(n2594), .IN2(g1088), .Q(n10414) );
  INVX0 U10212 ( .INP(n10415), .ZN(n10413) );
  OR2X1 U10213 ( .IN1(g1088), .IN2(n8396), .Q(n10415) );
  OR2X1 U10214 ( .IN1(n10416), .IN2(n10417), .Q(g30704) );
  INVX0 U10215 ( .INP(n10418), .ZN(n10417) );
  OR2X1 U10216 ( .IN1(n10419), .IN2(n8392), .Q(n10418) );
  AND2X1 U10217 ( .IN1(n10404), .IN2(g5511), .Q(n10416) );
  AND2X1 U10218 ( .IN1(n10420), .IN2(n10421), .Q(n10404) );
  XNOR2X1 U10219 ( .IN1(n10422), .IN2(n10423), .Q(n10421) );
  OR2X1 U10220 ( .IN1(n10424), .IN2(n10425), .Q(n10422) );
  OR2X1 U10221 ( .IN1(n10426), .IN2(n10427), .Q(n10425) );
  AND2X1 U10222 ( .IN1(n10428), .IN2(n10423), .Q(n10427) );
  AND2X1 U10223 ( .IN1(n10429), .IN2(n10430), .Q(n10428) );
  AND2X1 U10224 ( .IN1(n10431), .IN2(n10432), .Q(n10429) );
  OR2X1 U10225 ( .IN1(n10433), .IN2(n10434), .Q(n10432) );
  OR2X1 U10226 ( .IN1(n10435), .IN2(n10436), .Q(n10431) );
  AND2X1 U10227 ( .IN1(n10437), .IN2(n10438), .Q(n10435) );
  AND2X1 U10228 ( .IN1(n10439), .IN2(n10440), .Q(n10438) );
  AND2X1 U10229 ( .IN1(n10441), .IN2(n10442), .Q(n10437) );
  OR2X1 U10230 ( .IN1(n10443), .IN2(n10444), .Q(n10442) );
  AND2X1 U10231 ( .IN1(n10445), .IN2(n10446), .Q(n10426) );
  OR2X1 U10232 ( .IN1(n10447), .IN2(n10443), .Q(n10445) );
  AND2X1 U10233 ( .IN1(n10448), .IN2(n10449), .Q(n10447) );
  INVX0 U10234 ( .INP(n10450), .ZN(n10449) );
  AND2X1 U10235 ( .IN1(n10451), .IN2(n10452), .Q(n10448) );
  INVX0 U10236 ( .INP(n10453), .ZN(n10452) );
  OR2X1 U10237 ( .IN1(n10436), .IN2(n10454), .Q(n10451) );
  OR2X1 U10238 ( .IN1(n10455), .IN2(n10456), .Q(n10454) );
  AND2X1 U10239 ( .IN1(n10457), .IN2(n10458), .Q(n10424) );
  OR2X1 U10240 ( .IN1(n10459), .IN2(n10460), .Q(g30703) );
  AND2X1 U10241 ( .IN1(n2594), .IN2(g6712), .Q(n10460) );
  INVX0 U10242 ( .INP(n10461), .ZN(n10459) );
  OR2X1 U10243 ( .IN1(g6712), .IN2(n8381), .Q(n10461) );
  OR2X1 U10244 ( .IN1(n10462), .IN2(n10463), .Q(g30702) );
  INVX0 U10245 ( .INP(n10464), .ZN(n10463) );
  OR2X1 U10246 ( .IN1(n10465), .IN2(n8403), .Q(n10464) );
  AND2X1 U10247 ( .IN1(n10466), .IN2(n4640), .Q(n10462) );
  OR2X1 U10248 ( .IN1(n10467), .IN2(n10468), .Q(g30701) );
  AND2X1 U10249 ( .IN1(n2594), .IN2(g5472), .Q(n10468) );
  INVX0 U10250 ( .INP(n10469), .ZN(n10467) );
  OR2X1 U10251 ( .IN1(g5472), .IN2(n8397), .Q(n10469) );
  OR2X1 U10252 ( .IN1(n10470), .IN2(n10471), .Q(g30700) );
  AND2X1 U10253 ( .IN1(test_so18), .IN2(n4499), .Q(n10471) );
  AND2X1 U10254 ( .IN1(n10466), .IN2(g6447), .Q(n10470) );
  OR2X1 U10255 ( .IN1(n10472), .IN2(n10473), .Q(g30699) );
  INVX0 U10256 ( .INP(n10474), .ZN(n10473) );
  OR2X1 U10257 ( .IN1(n10475), .IN2(n8404), .Q(n10474) );
  AND2X1 U10258 ( .IN1(n10466), .IN2(g5437), .Q(n10472) );
  AND2X1 U10259 ( .IN1(n10476), .IN2(n10477), .Q(n10466) );
  XNOR2X1 U10260 ( .IN1(n10478), .IN2(n10479), .Q(n10477) );
  OR2X1 U10261 ( .IN1(n10480), .IN2(n10481), .Q(n10478) );
  OR2X1 U10262 ( .IN1(n10482), .IN2(n10483), .Q(n10481) );
  AND2X1 U10263 ( .IN1(n10484), .IN2(n10479), .Q(n10483) );
  AND2X1 U10264 ( .IN1(n10485), .IN2(n10486), .Q(n10484) );
  AND2X1 U10265 ( .IN1(n10487), .IN2(n10488), .Q(n10485) );
  OR2X1 U10266 ( .IN1(n10489), .IN2(n10490), .Q(n10488) );
  OR2X1 U10267 ( .IN1(n10491), .IN2(n10492), .Q(n10487) );
  AND2X1 U10268 ( .IN1(n10493), .IN2(n10494), .Q(n10491) );
  AND2X1 U10269 ( .IN1(n10495), .IN2(n10496), .Q(n10494) );
  AND2X1 U10270 ( .IN1(n10497), .IN2(n10498), .Q(n10493) );
  OR2X1 U10271 ( .IN1(n10499), .IN2(n10500), .Q(n10498) );
  AND2X1 U10272 ( .IN1(n10501), .IN2(n10502), .Q(n10482) );
  OR2X1 U10273 ( .IN1(n10503), .IN2(n10499), .Q(n10501) );
  AND2X1 U10274 ( .IN1(n10504), .IN2(n10505), .Q(n10503) );
  INVX0 U10275 ( .INP(n10506), .ZN(n10505) );
  AND2X1 U10276 ( .IN1(n10507), .IN2(n10508), .Q(n10504) );
  INVX0 U10277 ( .INP(n10509), .ZN(n10508) );
  OR2X1 U10278 ( .IN1(n10492), .IN2(n10510), .Q(n10507) );
  OR2X1 U10279 ( .IN1(n10511), .IN2(n10512), .Q(n10510) );
  AND2X1 U10280 ( .IN1(n10513), .IN2(n10514), .Q(n10480) );
  OR2X1 U10281 ( .IN1(n10515), .IN2(n10516), .Q(g30695) );
  AND2X1 U10282 ( .IN1(n10517), .IN2(g2241), .Q(n10516) );
  AND2X1 U10283 ( .IN1(n4367), .IN2(g2276), .Q(n10515) );
  OR2X1 U10284 ( .IN1(n10518), .IN2(n10519), .Q(g30694) );
  AND2X1 U10285 ( .IN1(n10520), .IN2(g2241), .Q(n10519) );
  AND2X1 U10286 ( .IN1(n4367), .IN2(g2348), .Q(n10518) );
  OR2X1 U10287 ( .IN1(n10521), .IN2(n10522), .Q(g30693) );
  AND2X1 U10288 ( .IN1(test_so73), .IN2(n10517), .Q(n10522) );
  AND2X1 U10289 ( .IN1(g2273), .IN2(n9119), .Q(n10521) );
  OR2X1 U10290 ( .IN1(n10523), .IN2(n10524), .Q(g30692) );
  AND2X1 U10291 ( .IN1(n10525), .IN2(g1547), .Q(n10524) );
  AND2X1 U10292 ( .IN1(n4368), .IN2(g1582), .Q(n10523) );
  OR2X1 U10293 ( .IN1(n10526), .IN2(n10527), .Q(g30691) );
  AND2X1 U10294 ( .IN1(n10520), .IN2(test_so73), .Q(n10527) );
  AND2X1 U10295 ( .IN1(g2345), .IN2(n9119), .Q(n10526) );
  OR2X1 U10296 ( .IN1(n10528), .IN2(n10529), .Q(g30690) );
  AND2X1 U10297 ( .IN1(n10517), .IN2(g6837), .Q(n10529) );
  OR2X1 U10298 ( .IN1(n10530), .IN2(n10531), .Q(n10517) );
  OR2X1 U10299 ( .IN1(n10532), .IN2(n10533), .Q(n10531) );
  AND2X1 U10300 ( .IN1(n10534), .IN2(g2175), .Q(n10533) );
  AND2X1 U10301 ( .IN1(n10535), .IN2(n10536), .Q(n10532) );
  XNOR2X1 U10302 ( .IN1(n10537), .IN2(n10538), .Q(n10535) );
  AND2X1 U10303 ( .IN1(n4324), .IN2(g2270), .Q(n10528) );
  OR2X1 U10304 ( .IN1(n10539), .IN2(n10540), .Q(g30689) );
  AND2X1 U10305 ( .IN1(n10541), .IN2(g1547), .Q(n10540) );
  AND2X1 U10306 ( .IN1(n4368), .IN2(g1654), .Q(n10539) );
  OR2X1 U10307 ( .IN1(n10542), .IN2(n10543), .Q(g30688) );
  AND2X1 U10308 ( .IN1(n10525), .IN2(g6782), .Q(n10543) );
  AND2X1 U10309 ( .IN1(n4515), .IN2(g1579), .Q(n10542) );
  OR2X1 U10310 ( .IN1(n10544), .IN2(n10545), .Q(g30687) );
  AND2X1 U10311 ( .IN1(test_so31), .IN2(n10546), .Q(n10545) );
  AND2X1 U10312 ( .IN1(g888), .IN2(n9118), .Q(n10544) );
  OR2X1 U10313 ( .IN1(n10547), .IN2(n10548), .Q(g30686) );
  AND2X1 U10314 ( .IN1(n10520), .IN2(g6837), .Q(n10548) );
  INVX0 U10315 ( .INP(n10549), .ZN(n10520) );
  OR2X1 U10316 ( .IN1(n10550), .IN2(n10551), .Q(n10549) );
  OR2X1 U10317 ( .IN1(n10552), .IN2(n10553), .Q(n10551) );
  AND2X1 U10318 ( .IN1(n10554), .IN2(n10536), .Q(n10553) );
  XOR2X1 U10319 ( .IN1(n9636), .IN2(n2669), .Q(n10554) );
  AND2X1 U10320 ( .IN1(n10534), .IN2(n10555), .Q(n10550) );
  AND2X1 U10321 ( .IN1(n4324), .IN2(g2342), .Q(n10547) );
  OR2X1 U10322 ( .IN1(n10556), .IN2(n10557), .Q(g30684) );
  AND2X1 U10323 ( .IN1(n10541), .IN2(g6782), .Q(n10557) );
  AND2X1 U10324 ( .IN1(n4515), .IN2(g1651), .Q(n10556) );
  OR2X1 U10325 ( .IN1(n10558), .IN2(n10559), .Q(g30683) );
  AND2X1 U10326 ( .IN1(n10525), .IN2(g6573), .Q(n10559) );
  OR2X1 U10327 ( .IN1(n10560), .IN2(n10561), .Q(n10525) );
  OR2X1 U10328 ( .IN1(n10562), .IN2(n10563), .Q(n10561) );
  AND2X1 U10329 ( .IN1(n10564), .IN2(g1481), .Q(n10563) );
  AND2X1 U10330 ( .IN1(n10565), .IN2(n10566), .Q(n10562) );
  XNOR2X1 U10331 ( .IN1(n10567), .IN2(n10568), .Q(n10565) );
  AND2X1 U10332 ( .IN1(n4317), .IN2(g1576), .Q(n10558) );
  OR2X1 U10333 ( .IN1(n10569), .IN2(n10570), .Q(g30682) );
  AND2X1 U10334 ( .IN1(n10571), .IN2(test_so31), .Q(n10570) );
  AND2X1 U10335 ( .IN1(g960), .IN2(n9118), .Q(n10569) );
  OR2X1 U10336 ( .IN1(n10572), .IN2(n10573), .Q(g30681) );
  AND2X1 U10337 ( .IN1(n10546), .IN2(g6518), .Q(n10573) );
  AND2X1 U10338 ( .IN1(n4312), .IN2(g885), .Q(n10572) );
  OR2X1 U10339 ( .IN1(n10574), .IN2(n10575), .Q(g30680) );
  AND2X1 U10340 ( .IN1(n10576), .IN2(g165), .Q(n10575) );
  AND2X1 U10341 ( .IN1(n4369), .IN2(g201), .Q(n10574) );
  OR2X1 U10342 ( .IN1(n10577), .IN2(n10578), .Q(g30679) );
  AND2X1 U10343 ( .IN1(n10579), .IN2(g2241), .Q(n10578) );
  AND2X1 U10344 ( .IN1(n4367), .IN2(g2321), .Q(n10577) );
  OR2X1 U10345 ( .IN1(n10580), .IN2(n10581), .Q(g30678) );
  AND2X1 U10346 ( .IN1(n10541), .IN2(g6573), .Q(n10581) );
  INVX0 U10347 ( .INP(n10582), .ZN(n10541) );
  OR2X1 U10348 ( .IN1(n10583), .IN2(n10584), .Q(n10582) );
  OR2X1 U10349 ( .IN1(n10585), .IN2(n10586), .Q(n10584) );
  AND2X1 U10350 ( .IN1(n10587), .IN2(n10566), .Q(n10586) );
  XNOR2X1 U10351 ( .IN1(n10588), .IN2(n2684), .Q(n10587) );
  AND2X1 U10352 ( .IN1(n10564), .IN2(n10589), .Q(n10583) );
  AND2X1 U10353 ( .IN1(n4317), .IN2(g1648), .Q(n10580) );
  OR2X1 U10354 ( .IN1(n10590), .IN2(n10591), .Q(g30677) );
  AND2X1 U10355 ( .IN1(n10571), .IN2(g6518), .Q(n10591) );
  AND2X1 U10356 ( .IN1(n4312), .IN2(g957), .Q(n10590) );
  OR2X1 U10357 ( .IN1(n10592), .IN2(n10593), .Q(g30676) );
  AND2X1 U10358 ( .IN1(n10546), .IN2(g6368), .Q(n10593) );
  OR2X1 U10359 ( .IN1(n10594), .IN2(n10595), .Q(n10546) );
  OR2X1 U10360 ( .IN1(n10596), .IN2(n10597), .Q(n10595) );
  AND2X1 U10361 ( .IN1(n10598), .IN2(g793), .Q(n10597) );
  AND2X1 U10362 ( .IN1(n10599), .IN2(n10600), .Q(n10596) );
  XNOR2X1 U10363 ( .IN1(n10601), .IN2(n9585), .Q(n10599) );
  AND2X1 U10364 ( .IN1(n4323), .IN2(g882), .Q(n10592) );
  OR2X1 U10365 ( .IN1(n10602), .IN2(n10603), .Q(g30675) );
  AND2X1 U10366 ( .IN1(n10604), .IN2(g165), .Q(n10603) );
  AND2X1 U10367 ( .IN1(n4369), .IN2(g273), .Q(n10602) );
  OR2X1 U10368 ( .IN1(n10605), .IN2(n10606), .Q(g30674) );
  AND2X1 U10369 ( .IN1(n10576), .IN2(g6313), .Q(n10606) );
  AND2X1 U10370 ( .IN1(n4512), .IN2(g198), .Q(n10605) );
  OR2X1 U10371 ( .IN1(n10607), .IN2(n10608), .Q(g30673) );
  AND2X1 U10372 ( .IN1(n10579), .IN2(test_so73), .Q(n10608) );
  AND2X1 U10373 ( .IN1(g2318), .IN2(n9119), .Q(n10607) );
  OR2X1 U10374 ( .IN1(n10609), .IN2(n10610), .Q(g30672) );
  AND2X1 U10375 ( .IN1(n10611), .IN2(g2241), .Q(n10610) );
  AND2X1 U10376 ( .IN1(n4367), .IN2(g2312), .Q(n10609) );
  OR2X1 U10377 ( .IN1(n10612), .IN2(n10613), .Q(g30671) );
  AND2X1 U10378 ( .IN1(n10614), .IN2(g1547), .Q(n10613) );
  AND2X1 U10379 ( .IN1(n4368), .IN2(g1627), .Q(n10612) );
  OR2X1 U10380 ( .IN1(n10615), .IN2(n10616), .Q(g30670) );
  AND2X1 U10381 ( .IN1(n10571), .IN2(g6368), .Q(n10616) );
  INVX0 U10382 ( .INP(n10617), .ZN(n10571) );
  OR2X1 U10383 ( .IN1(n10618), .IN2(n10619), .Q(n10617) );
  OR2X1 U10384 ( .IN1(n10620), .IN2(n10621), .Q(n10619) );
  AND2X1 U10385 ( .IN1(n10600), .IN2(n10622), .Q(n10621) );
  XOR2X1 U10386 ( .IN1(n10623), .IN2(n10624), .Q(n10622) );
  OR2X1 U10387 ( .IN1(n10625), .IN2(n10626), .Q(n10624) );
  XNOR2X1 U10388 ( .IN1(n10627), .IN2(n10628), .Q(n10625) );
  AND2X1 U10389 ( .IN1(n10598), .IN2(n10629), .Q(n10618) );
  AND2X1 U10390 ( .IN1(n4323), .IN2(g954), .Q(n10615) );
  OR2X1 U10391 ( .IN1(n10630), .IN2(n10631), .Q(g30669) );
  AND2X1 U10392 ( .IN1(n10604), .IN2(g6313), .Q(n10631) );
  AND2X1 U10393 ( .IN1(n4512), .IN2(g270), .Q(n10630) );
  OR2X1 U10394 ( .IN1(n10632), .IN2(n10633), .Q(g30668) );
  AND2X1 U10395 ( .IN1(n10576), .IN2(g6231), .Q(n10633) );
  OR2X1 U10396 ( .IN1(n10634), .IN2(n10635), .Q(n10576) );
  OR2X1 U10397 ( .IN1(n10636), .IN2(n10637), .Q(n10635) );
  AND2X1 U10398 ( .IN1(n10638), .IN2(g105), .Q(n10637) );
  AND2X1 U10399 ( .IN1(n10639), .IN2(n10640), .Q(n10636) );
  XNOR2X1 U10400 ( .IN1(n10641), .IN2(n10642), .Q(n10639) );
  AND2X1 U10401 ( .IN1(n4318), .IN2(g195), .Q(n10632) );
  OR2X1 U10402 ( .IN1(n10643), .IN2(n10644), .Q(g30667) );
  AND2X1 U10403 ( .IN1(n10579), .IN2(g6837), .Q(n10644) );
  INVX0 U10404 ( .INP(n10645), .ZN(n10579) );
  OR2X1 U10405 ( .IN1(n10646), .IN2(n10647), .Q(n10645) );
  OR2X1 U10406 ( .IN1(n10552), .IN2(n10648), .Q(n10647) );
  AND2X1 U10407 ( .IN1(n10536), .IN2(n10649), .Q(n10648) );
  XNOR2X1 U10408 ( .IN1(n10650), .IN2(n9644), .Q(n10649) );
  AND2X1 U10409 ( .IN1(n10537), .IN2(n10651), .Q(n10650) );
  XNOR2X1 U10410 ( .IN1(n9654), .IN2(n4529), .Q(n10651) );
  INVX0 U10411 ( .INP(n10652), .ZN(n10537) );
  AND2X1 U10412 ( .IN1(n10534), .IN2(n4389), .Q(n10646) );
  AND2X1 U10413 ( .IN1(n4324), .IN2(g2315), .Q(n10643) );
  OR2X1 U10414 ( .IN1(n10653), .IN2(n10654), .Q(g30666) );
  AND2X1 U10415 ( .IN1(n10611), .IN2(test_so73), .Q(n10654) );
  AND2X1 U10416 ( .IN1(g2309), .IN2(n9119), .Q(n10653) );
  OR2X1 U10417 ( .IN1(n10655), .IN2(n10656), .Q(g30665) );
  AND2X1 U10418 ( .IN1(n10657), .IN2(g2241), .Q(n10656) );
  AND2X1 U10419 ( .IN1(n4367), .IN2(g2303), .Q(n10655) );
  OR2X1 U10420 ( .IN1(n10658), .IN2(n10659), .Q(g30664) );
  AND2X1 U10421 ( .IN1(n10614), .IN2(g6782), .Q(n10659) );
  AND2X1 U10422 ( .IN1(n4515), .IN2(g1624), .Q(n10658) );
  OR2X1 U10423 ( .IN1(n10660), .IN2(n10661), .Q(g30663) );
  AND2X1 U10424 ( .IN1(n10662), .IN2(g1547), .Q(n10661) );
  AND2X1 U10425 ( .IN1(n4368), .IN2(g1618), .Q(n10660) );
  OR2X1 U10426 ( .IN1(n10663), .IN2(n10664), .Q(g30662) );
  AND2X1 U10427 ( .IN1(n10665), .IN2(test_so31), .Q(n10664) );
  AND2X1 U10428 ( .IN1(g933), .IN2(n9118), .Q(n10663) );
  OR2X1 U10429 ( .IN1(n10666), .IN2(n10667), .Q(g30661) );
  AND2X1 U10430 ( .IN1(n10604), .IN2(g6231), .Q(n10667) );
  INVX0 U10431 ( .INP(n10668), .ZN(n10604) );
  OR2X1 U10432 ( .IN1(n10669), .IN2(n10670), .Q(n10668) );
  OR2X1 U10433 ( .IN1(n10671), .IN2(n10672), .Q(n10670) );
  AND2X1 U10434 ( .IN1(n10673), .IN2(n10640), .Q(n10672) );
  XOR2X1 U10435 ( .IN1(n9539), .IN2(n2717), .Q(n10673) );
  AND2X1 U10436 ( .IN1(n10638), .IN2(n10674), .Q(n10669) );
  AND2X1 U10437 ( .IN1(n4318), .IN2(g267), .Q(n10666) );
  OR2X1 U10438 ( .IN1(n10675), .IN2(n10676), .Q(g30660) );
  AND2X1 U10439 ( .IN1(n10611), .IN2(g6837), .Q(n10676) );
  INVX0 U10440 ( .INP(n10677), .ZN(n10611) );
  OR2X1 U10441 ( .IN1(n10678), .IN2(n10679), .Q(n10677) );
  OR2X1 U10442 ( .IN1(n10552), .IN2(n10680), .Q(n10679) );
  AND2X1 U10443 ( .IN1(n10536), .IN2(n10681), .Q(n10680) );
  XNOR2X1 U10444 ( .IN1(n10682), .IN2(n9658), .Q(n10681) );
  AND2X1 U10445 ( .IN1(n4529), .IN2(n10683), .Q(n10552) );
  AND2X1 U10446 ( .IN1(n10534), .IN2(n4373), .Q(n10678) );
  AND2X1 U10447 ( .IN1(n4324), .IN2(g2306), .Q(n10675) );
  OR2X1 U10448 ( .IN1(n10684), .IN2(n10685), .Q(g30659) );
  AND2X1 U10449 ( .IN1(test_so73), .IN2(n10657), .Q(n10685) );
  AND2X1 U10450 ( .IN1(g2300), .IN2(n9119), .Q(n10684) );
  OR2X1 U10451 ( .IN1(n10686), .IN2(n10687), .Q(g30658) );
  AND2X1 U10452 ( .IN1(test_so55), .IN2(n4317), .Q(n10687) );
  AND2X1 U10453 ( .IN1(n10614), .IN2(g6573), .Q(n10686) );
  INVX0 U10454 ( .INP(n10688), .ZN(n10614) );
  OR2X1 U10455 ( .IN1(n10689), .IN2(n10690), .Q(n10688) );
  OR2X1 U10456 ( .IN1(n10585), .IN2(n10691), .Q(n10690) );
  AND2X1 U10457 ( .IN1(n10566), .IN2(n10692), .Q(n10691) );
  XNOR2X1 U10458 ( .IN1(n10693), .IN2(n9610), .Q(n10692) );
  AND2X1 U10459 ( .IN1(n10567), .IN2(n10694), .Q(n10693) );
  XNOR2X1 U10460 ( .IN1(n9617), .IN2(n4530), .Q(n10694) );
  INVX0 U10461 ( .INP(n10695), .ZN(n10567) );
  AND2X1 U10462 ( .IN1(n10564), .IN2(n4390), .Q(n10689) );
  OR2X1 U10463 ( .IN1(n10696), .IN2(n10697), .Q(g30657) );
  AND2X1 U10464 ( .IN1(n10662), .IN2(g6782), .Q(n10697) );
  AND2X1 U10465 ( .IN1(n4515), .IN2(g1615), .Q(n10696) );
  OR2X1 U10466 ( .IN1(n10698), .IN2(n10699), .Q(g30656) );
  AND2X1 U10467 ( .IN1(n10700), .IN2(g1547), .Q(n10699) );
  AND2X1 U10468 ( .IN1(n4368), .IN2(g1609), .Q(n10698) );
  OR2X1 U10469 ( .IN1(n10701), .IN2(n10702), .Q(g30655) );
  AND2X1 U10470 ( .IN1(n10665), .IN2(g6518), .Q(n10702) );
  AND2X1 U10471 ( .IN1(n4312), .IN2(g930), .Q(n10701) );
  OR2X1 U10472 ( .IN1(n10703), .IN2(n10704), .Q(g30654) );
  AND2X1 U10473 ( .IN1(n10705), .IN2(test_so31), .Q(n10704) );
  AND2X1 U10474 ( .IN1(test_so34), .IN2(n9118), .Q(n10703) );
  OR2X1 U10475 ( .IN1(n10706), .IN2(n10707), .Q(g30653) );
  AND2X1 U10476 ( .IN1(n10708), .IN2(g165), .Q(n10707) );
  AND2X1 U10477 ( .IN1(n4369), .IN2(g246), .Q(n10706) );
  OR2X1 U10478 ( .IN1(n10709), .IN2(n10710), .Q(g30652) );
  AND2X1 U10479 ( .IN1(n10657), .IN2(g6837), .Q(n10710) );
  OR2X1 U10480 ( .IN1(n10530), .IN2(n10711), .Q(n10657) );
  OR2X1 U10481 ( .IN1(n10712), .IN2(n10713), .Q(n10711) );
  AND2X1 U10482 ( .IN1(n10534), .IN2(n10714), .Q(n10713) );
  AND2X1 U10483 ( .IN1(n10715), .IN2(n10536), .Q(n10712) );
  XNOR2X1 U10484 ( .IN1(n9643), .IN2(n2670), .Q(n10715) );
  OR2X1 U10485 ( .IN1(n10716), .IN2(n10717), .Q(n2670) );
  XNOR2X1 U10486 ( .IN1(n10718), .IN2(n9638), .Q(n10716) );
  AND2X1 U10487 ( .IN1(n10683), .IN2(n10719), .Q(n10530) );
  INVX0 U10488 ( .INP(n10720), .ZN(n10683) );
  AND2X1 U10489 ( .IN1(n4324), .IN2(g2297), .Q(n10709) );
  OR2X1 U10490 ( .IN1(n10721), .IN2(n10722), .Q(g30651) );
  AND2X1 U10491 ( .IN1(n10662), .IN2(g6573), .Q(n10722) );
  INVX0 U10492 ( .INP(n10723), .ZN(n10662) );
  OR2X1 U10493 ( .IN1(n10724), .IN2(n10725), .Q(n10723) );
  OR2X1 U10494 ( .IN1(n10585), .IN2(n10726), .Q(n10725) );
  AND2X1 U10495 ( .IN1(n10566), .IN2(n10727), .Q(n10726) );
  XNOR2X1 U10496 ( .IN1(n10728), .IN2(n10729), .Q(n10727) );
  AND2X1 U10497 ( .IN1(n4530), .IN2(n10730), .Q(n10585) );
  AND2X1 U10498 ( .IN1(n10564), .IN2(n4374), .Q(n10724) );
  AND2X1 U10499 ( .IN1(n4317), .IN2(g1612), .Q(n10721) );
  OR2X1 U10500 ( .IN1(n10731), .IN2(n10732), .Q(g30650) );
  AND2X1 U10501 ( .IN1(n10700), .IN2(g6782), .Q(n10732) );
  AND2X1 U10502 ( .IN1(test_so56), .IN2(n4515), .Q(n10731) );
  OR2X1 U10503 ( .IN1(n10733), .IN2(n10734), .Q(g30649) );
  AND2X1 U10504 ( .IN1(n10665), .IN2(g6368), .Q(n10734) );
  INVX0 U10505 ( .INP(n10735), .ZN(n10665) );
  OR2X1 U10506 ( .IN1(n10736), .IN2(n10737), .Q(n10735) );
  OR2X1 U10507 ( .IN1(n10620), .IN2(n10738), .Q(n10737) );
  AND2X1 U10508 ( .IN1(n10600), .IN2(n10739), .Q(n10738) );
  XNOR2X1 U10509 ( .IN1(n9567), .IN2(n10740), .Q(n10739) );
  AND2X1 U10510 ( .IN1(n10741), .IN2(n10742), .Q(n10740) );
  OR2X1 U10511 ( .IN1(n9585), .IN2(n10743), .Q(n10742) );
  INVX0 U10512 ( .INP(n10744), .ZN(n10741) );
  AND2X1 U10513 ( .IN1(n10598), .IN2(n4391), .Q(n10736) );
  AND2X1 U10514 ( .IN1(n4323), .IN2(g927), .Q(n10733) );
  OR2X1 U10515 ( .IN1(n10745), .IN2(n10746), .Q(g30648) );
  AND2X1 U10516 ( .IN1(n10705), .IN2(g6518), .Q(n10746) );
  AND2X1 U10517 ( .IN1(n4312), .IN2(g921), .Q(n10745) );
  OR2X1 U10518 ( .IN1(n10747), .IN2(n10748), .Q(g30647) );
  AND2X1 U10519 ( .IN1(test_so31), .IN2(n10749), .Q(n10748) );
  AND2X1 U10520 ( .IN1(g915), .IN2(n9118), .Q(n10747) );
  OR2X1 U10521 ( .IN1(n10750), .IN2(n10751), .Q(g30646) );
  AND2X1 U10522 ( .IN1(n10708), .IN2(g6313), .Q(n10751) );
  AND2X1 U10523 ( .IN1(n4512), .IN2(g243), .Q(n10750) );
  OR2X1 U10524 ( .IN1(n10752), .IN2(n10753), .Q(g30645) );
  AND2X1 U10525 ( .IN1(n10754), .IN2(g165), .Q(n10753) );
  AND2X1 U10526 ( .IN1(n4369), .IN2(g237), .Q(n10752) );
  OR2X1 U10527 ( .IN1(n10755), .IN2(n10756), .Q(g30644) );
  AND2X1 U10528 ( .IN1(n10700), .IN2(g6573), .Q(n10756) );
  OR2X1 U10529 ( .IN1(n10560), .IN2(n10757), .Q(n10700) );
  OR2X1 U10530 ( .IN1(n10758), .IN2(n10759), .Q(n10757) );
  AND2X1 U10531 ( .IN1(n10564), .IN2(n10760), .Q(n10759) );
  AND2X1 U10532 ( .IN1(n10761), .IN2(n10566), .Q(n10758) );
  XOR2X1 U10533 ( .IN1(n10762), .IN2(n2685), .Q(n10761) );
  OR2X1 U10534 ( .IN1(n10763), .IN2(n10764), .Q(n2685) );
  XNOR2X1 U10535 ( .IN1(n10765), .IN2(n9603), .Q(n10763) );
  AND2X1 U10536 ( .IN1(n10730), .IN2(n10766), .Q(n10560) );
  INVX0 U10537 ( .INP(n10767), .ZN(n10730) );
  AND2X1 U10538 ( .IN1(n4317), .IN2(g1603), .Q(n10755) );
  OR2X1 U10539 ( .IN1(n10768), .IN2(n10769), .Q(g30643) );
  AND2X1 U10540 ( .IN1(n10705), .IN2(g6368), .Q(n10769) );
  INVX0 U10541 ( .INP(n10770), .ZN(n10705) );
  OR2X1 U10542 ( .IN1(n10771), .IN2(n10772), .Q(n10770) );
  OR2X1 U10543 ( .IN1(n10620), .IN2(n10773), .Q(n10772) );
  AND2X1 U10544 ( .IN1(n10600), .IN2(n10774), .Q(n10773) );
  XNOR2X1 U10545 ( .IN1(n10775), .IN2(n10776), .Q(n10774) );
  AND2X1 U10546 ( .IN1(n10627), .IN2(n10777), .Q(n10620) );
  AND2X1 U10547 ( .IN1(n10598), .IN2(n4375), .Q(n10771) );
  AND2X1 U10548 ( .IN1(n4323), .IN2(g918), .Q(n10768) );
  OR2X1 U10549 ( .IN1(n10778), .IN2(n10779), .Q(g30642) );
  AND2X1 U10550 ( .IN1(n10749), .IN2(g6518), .Q(n10779) );
  AND2X1 U10551 ( .IN1(n4312), .IN2(g912), .Q(n10778) );
  OR2X1 U10552 ( .IN1(n10780), .IN2(n10781), .Q(g30641) );
  AND2X1 U10553 ( .IN1(n10708), .IN2(g6231), .Q(n10781) );
  INVX0 U10554 ( .INP(n10782), .ZN(n10708) );
  OR2X1 U10555 ( .IN1(n10783), .IN2(n10784), .Q(n10782) );
  OR2X1 U10556 ( .IN1(n10671), .IN2(n10785), .Q(n10784) );
  AND2X1 U10557 ( .IN1(n10640), .IN2(n10786), .Q(n10785) );
  XNOR2X1 U10558 ( .IN1(n10787), .IN2(n9554), .Q(n10786) );
  AND2X1 U10559 ( .IN1(n10641), .IN2(n10788), .Q(n10787) );
  XNOR2X1 U10560 ( .IN1(n9548), .IN2(n10252), .Q(n10788) );
  INVX0 U10561 ( .INP(n10789), .ZN(n10641) );
  AND2X1 U10562 ( .IN1(n10638), .IN2(n4392), .Q(n10783) );
  AND2X1 U10563 ( .IN1(n4318), .IN2(g240), .Q(n10780) );
  OR2X1 U10564 ( .IN1(n10790), .IN2(n10791), .Q(g30640) );
  AND2X1 U10565 ( .IN1(n10754), .IN2(g6313), .Q(n10791) );
  AND2X1 U10566 ( .IN1(n4512), .IN2(g234), .Q(n10790) );
  OR2X1 U10567 ( .IN1(n10792), .IN2(n10793), .Q(g30639) );
  AND2X1 U10568 ( .IN1(n10794), .IN2(g165), .Q(n10793) );
  AND2X1 U10569 ( .IN1(n4369), .IN2(g228), .Q(n10792) );
  OR2X1 U10570 ( .IN1(n10795), .IN2(n10796), .Q(g30638) );
  AND2X1 U10571 ( .IN1(n10749), .IN2(g6368), .Q(n10796) );
  OR2X1 U10572 ( .IN1(n10594), .IN2(n10797), .Q(n10749) );
  OR2X1 U10573 ( .IN1(n10798), .IN2(n10799), .Q(n10797) );
  AND2X1 U10574 ( .IN1(n10598), .IN2(n10800), .Q(n10799) );
  AND2X1 U10575 ( .IN1(n10801), .IN2(n10600), .Q(n10798) );
  XNOR2X1 U10576 ( .IN1(n10626), .IN2(n9584), .Q(n10801) );
  OR2X1 U10577 ( .IN1(n10802), .IN2(n10803), .Q(n10626) );
  OR2X1 U10578 ( .IN1(n10804), .IN2(n10805), .Q(n10803) );
  INVX0 U10579 ( .INP(n10806), .ZN(n10805) );
  OR2X1 U10580 ( .IN1(n10743), .IN2(n9589), .Q(n10806) );
  AND2X1 U10581 ( .IN1(n10807), .IN2(n9589), .Q(n10804) );
  AND2X1 U10582 ( .IN1(n10777), .IN2(n10743), .Q(n10594) );
  AND2X1 U10583 ( .IN1(n4323), .IN2(g909), .Q(n10795) );
  OR2X1 U10584 ( .IN1(n10808), .IN2(n10809), .Q(g30637) );
  AND2X1 U10585 ( .IN1(n10754), .IN2(g6231), .Q(n10809) );
  INVX0 U10586 ( .INP(n10810), .ZN(n10754) );
  OR2X1 U10587 ( .IN1(n10811), .IN2(n10812), .Q(n10810) );
  OR2X1 U10588 ( .IN1(n10671), .IN2(n10813), .Q(n10812) );
  AND2X1 U10589 ( .IN1(n10640), .IN2(n10814), .Q(n10813) );
  XOR2X1 U10590 ( .IN1(n10815), .IN2(n9531), .Q(n10814) );
  AND2X1 U10591 ( .IN1(n10252), .IN2(n10816), .Q(n10671) );
  AND2X1 U10592 ( .IN1(n10638), .IN2(n4376), .Q(n10811) );
  AND2X1 U10593 ( .IN1(n4318), .IN2(g231), .Q(n10808) );
  OR2X1 U10594 ( .IN1(n10817), .IN2(n10818), .Q(g30636) );
  AND2X1 U10595 ( .IN1(n10794), .IN2(g6313), .Q(n10818) );
  AND2X1 U10596 ( .IN1(n4512), .IN2(g225), .Q(n10817) );
  OR2X1 U10597 ( .IN1(n10819), .IN2(n10820), .Q(g30635) );
  AND2X1 U10598 ( .IN1(n10794), .IN2(g6231), .Q(n10820) );
  OR2X1 U10599 ( .IN1(n10634), .IN2(n10821), .Q(n10794) );
  OR2X1 U10600 ( .IN1(n10822), .IN2(n10823), .Q(n10821) );
  AND2X1 U10601 ( .IN1(n10638), .IN2(n10824), .Q(n10823) );
  AND2X1 U10602 ( .IN1(n10825), .IN2(n10640), .Q(n10822) );
  XNOR2X1 U10603 ( .IN1(n9540), .IN2(n2718), .Q(n10825) );
  OR2X1 U10604 ( .IN1(n10826), .IN2(n10827), .Q(n2718) );
  XNOR2X1 U10605 ( .IN1(n10252), .IN2(n10828), .Q(n10826) );
  AND2X1 U10606 ( .IN1(n10816), .IN2(n10829), .Q(n10634) );
  AND2X1 U10607 ( .IN1(n4318), .IN2(g222), .Q(n10819) );
  OR2X1 U10608 ( .IN1(n10830), .IN2(n10831), .Q(g30566) );
  INVX0 U10609 ( .INP(n10832), .ZN(n10831) );
  OR2X1 U10610 ( .IN1(n10833), .IN2(n8385), .Q(n10832) );
  AND2X1 U10611 ( .IN1(n10399), .IN2(n4606), .Q(n10830) );
  AND2X1 U10612 ( .IN1(n10834), .IN2(n10835), .Q(n10399) );
  XNOR2X1 U10613 ( .IN1(n10836), .IN2(n10837), .Q(n10835) );
  OR2X1 U10614 ( .IN1(n10838), .IN2(n10839), .Q(n10836) );
  OR2X1 U10615 ( .IN1(n10840), .IN2(n10841), .Q(n10839) );
  AND2X1 U10616 ( .IN1(n10842), .IN2(n10837), .Q(n10841) );
  AND2X1 U10617 ( .IN1(n10843), .IN2(n10844), .Q(n10842) );
  AND2X1 U10618 ( .IN1(n10845), .IN2(n10846), .Q(n10843) );
  OR2X1 U10619 ( .IN1(n10847), .IN2(n10848), .Q(n10846) );
  OR2X1 U10620 ( .IN1(n10849), .IN2(n10850), .Q(n10845) );
  AND2X1 U10621 ( .IN1(n10851), .IN2(n10852), .Q(n10849) );
  AND2X1 U10622 ( .IN1(n10853), .IN2(n10854), .Q(n10852) );
  AND2X1 U10623 ( .IN1(n10855), .IN2(n10856), .Q(n10851) );
  OR2X1 U10624 ( .IN1(n10857), .IN2(n10858), .Q(n10856) );
  AND2X1 U10625 ( .IN1(n10859), .IN2(n10860), .Q(n10840) );
  OR2X1 U10626 ( .IN1(n10861), .IN2(n10857), .Q(n10859) );
  AND2X1 U10627 ( .IN1(n10862), .IN2(n10863), .Q(n10861) );
  INVX0 U10628 ( .INP(n10864), .ZN(n10863) );
  AND2X1 U10629 ( .IN1(n10865), .IN2(n10866), .Q(n10862) );
  INVX0 U10630 ( .INP(n10867), .ZN(n10866) );
  OR2X1 U10631 ( .IN1(n10850), .IN2(n10868), .Q(n10865) );
  OR2X1 U10632 ( .IN1(n10869), .IN2(n10870), .Q(n10868) );
  AND2X1 U10633 ( .IN1(n10871), .IN2(n10872), .Q(n10838) );
  OR2X1 U10634 ( .IN1(n10873), .IN2(n10874), .Q(g30505) );
  INVX0 U10635 ( .INP(n10875), .ZN(n10874) );
  OR2X1 U10636 ( .IN1(n10408), .IN2(n8384), .Q(n10875) );
  AND2X1 U10637 ( .IN1(n10876), .IN2(g5555), .Q(n10873) );
  OR2X1 U10638 ( .IN1(n10877), .IN2(n10878), .Q(g30503) );
  INVX0 U10639 ( .INP(n10879), .ZN(n10878) );
  OR2X1 U10640 ( .IN1(n10412), .IN2(n8377), .Q(n10879) );
  AND2X1 U10641 ( .IN1(n10880), .IN2(g7014), .Q(n10877) );
  OR2X1 U10642 ( .IN1(n10881), .IN2(n10882), .Q(g30500) );
  AND2X1 U10643 ( .IN1(test_so39), .IN2(n4381), .Q(n10882) );
  AND2X1 U10644 ( .IN1(n2798), .IN2(g1088), .Q(n10881) );
  OR2X1 U10645 ( .IN1(n10883), .IN2(n10884), .Q(g30487) );
  INVX0 U10646 ( .INP(n10885), .ZN(n10884) );
  OR2X1 U10647 ( .IN1(n10419), .IN2(n8390), .Q(n10885) );
  AND2X1 U10648 ( .IN1(n10880), .IN2(g5511), .Q(n10883) );
  OR2X1 U10649 ( .IN1(n10886), .IN2(n10887), .Q(g30485) );
  AND2X1 U10650 ( .IN1(n2798), .IN2(g6712), .Q(n10887) );
  INVX0 U10651 ( .INP(n10888), .ZN(n10886) );
  OR2X1 U10652 ( .IN1(g6712), .IN2(n8380), .Q(n10888) );
  OR2X1 U10653 ( .IN1(n10889), .IN2(n10890), .Q(g30482) );
  INVX0 U10654 ( .INP(n10891), .ZN(n10890) );
  OR2X1 U10655 ( .IN1(n10465), .IN2(n8400), .Q(n10891) );
  AND2X1 U10656 ( .IN1(n10892), .IN2(n4640), .Q(n10889) );
  OR2X1 U10657 ( .IN1(n10893), .IN2(n10894), .Q(g30470) );
  AND2X1 U10658 ( .IN1(n2798), .IN2(g5472), .Q(n10894) );
  INVX0 U10659 ( .INP(n10895), .ZN(n10893) );
  OR2X1 U10660 ( .IN1(g5472), .IN2(n8395), .Q(n10895) );
  OR2X1 U10661 ( .IN1(n10896), .IN2(n10897), .Q(g30468) );
  INVX0 U10662 ( .INP(n10898), .ZN(n10897) );
  OR2X1 U10663 ( .IN1(n10899), .IN2(n8401), .Q(n10898) );
  AND2X1 U10664 ( .IN1(n10892), .IN2(g6447), .Q(n10896) );
  OR2X1 U10665 ( .IN1(n10900), .IN2(n10901), .Q(g30455) );
  INVX0 U10666 ( .INP(n10902), .ZN(n10901) );
  OR2X1 U10667 ( .IN1(n10475), .IN2(n8402), .Q(n10902) );
  AND2X1 U10668 ( .IN1(n10892), .IN2(g5437), .Q(n10900) );
  AND2X1 U10669 ( .IN1(n10476), .IN2(n10903), .Q(n10892) );
  AND2X1 U10670 ( .IN1(n10904), .IN2(n10905), .Q(n10903) );
  INVX0 U10671 ( .INP(n10906), .ZN(n10905) );
  AND2X1 U10672 ( .IN1(n10907), .IN2(n10908), .Q(n10906) );
  OR2X1 U10673 ( .IN1(n10513), .IN2(n10492), .Q(n10907) );
  OR2X1 U10674 ( .IN1(n10908), .IN2(n10492), .Q(n10904) );
  OR2X1 U10675 ( .IN1(n10909), .IN2(n10910), .Q(n10908) );
  OR2X1 U10676 ( .IN1(n10513), .IN2(n10911), .Q(n10910) );
  AND2X1 U10677 ( .IN1(n10912), .IN2(n10492), .Q(n10911) );
  OR2X1 U10678 ( .IN1(n10913), .IN2(n10914), .Q(n10909) );
  AND2X1 U10679 ( .IN1(n10915), .IN2(n10502), .Q(n10914) );
  AND2X1 U10680 ( .IN1(n10916), .IN2(n10486), .Q(n10915) );
  OR2X1 U10681 ( .IN1(n10917), .IN2(n10499), .Q(n10916) );
  AND2X1 U10682 ( .IN1(n10489), .IN2(n10500), .Q(n10917) );
  INVX0 U10683 ( .INP(n10511), .ZN(n10500) );
  AND2X1 U10684 ( .IN1(n10479), .IN2(n10918), .Q(n10913) );
  OR2X1 U10685 ( .IN1(n4388), .IN2(n10919), .Q(n10918) );
  OR2X1 U10686 ( .IN1(n10920), .IN2(n10921), .Q(g30356) );
  INVX0 U10687 ( .INP(n10922), .ZN(n10921) );
  OR2X1 U10688 ( .IN1(n10833), .IN2(n8383), .Q(n10922) );
  AND2X1 U10689 ( .IN1(n10876), .IN2(n4606), .Q(n10920) );
  OR2X1 U10690 ( .IN1(n10923), .IN2(n10924), .Q(g30341) );
  INVX0 U10691 ( .INP(n10925), .ZN(n10924) );
  OR2X1 U10692 ( .IN1(n10398), .IN2(n8374), .Q(n10925) );
  AND2X1 U10693 ( .IN1(n10876), .IN2(g7264), .Q(n10923) );
  AND2X1 U10694 ( .IN1(n10834), .IN2(n10926), .Q(n10876) );
  AND2X1 U10695 ( .IN1(n10927), .IN2(n10928), .Q(n10926) );
  INVX0 U10696 ( .INP(n10929), .ZN(n10928) );
  AND2X1 U10697 ( .IN1(n10930), .IN2(n10931), .Q(n10929) );
  OR2X1 U10698 ( .IN1(n10871), .IN2(n10850), .Q(n10930) );
  OR2X1 U10699 ( .IN1(n10931), .IN2(n10850), .Q(n10927) );
  OR2X1 U10700 ( .IN1(n10932), .IN2(n10933), .Q(n10931) );
  OR2X1 U10701 ( .IN1(n10871), .IN2(n10934), .Q(n10933) );
  AND2X1 U10702 ( .IN1(n10935), .IN2(n10850), .Q(n10934) );
  OR2X1 U10703 ( .IN1(n10936), .IN2(n10937), .Q(n10932) );
  AND2X1 U10704 ( .IN1(n10938), .IN2(n10860), .Q(n10937) );
  AND2X1 U10705 ( .IN1(n10939), .IN2(n10844), .Q(n10938) );
  OR2X1 U10706 ( .IN1(n10940), .IN2(n10857), .Q(n10939) );
  AND2X1 U10707 ( .IN1(n10847), .IN2(n10858), .Q(n10940) );
  INVX0 U10708 ( .INP(n10870), .ZN(n10858) );
  AND2X1 U10709 ( .IN1(n10837), .IN2(n10941), .Q(n10936) );
  OR2X1 U10710 ( .IN1(n10942), .IN2(n9121), .Q(n10941) );
  OR2X1 U10711 ( .IN1(n10943), .IN2(n10944), .Q(g30338) );
  INVX0 U10712 ( .INP(n10945), .ZN(n10944) );
  OR2X1 U10713 ( .IN1(n10403), .IN2(n8389), .Q(n10945) );
  AND2X1 U10714 ( .IN1(n10880), .IN2(n4618), .Q(n10943) );
  AND2X1 U10715 ( .IN1(n10420), .IN2(n10946), .Q(n10880) );
  AND2X1 U10716 ( .IN1(n10947), .IN2(n10948), .Q(n10946) );
  INVX0 U10717 ( .INP(n10949), .ZN(n10948) );
  AND2X1 U10718 ( .IN1(n10950), .IN2(n10951), .Q(n10949) );
  OR2X1 U10719 ( .IN1(n10457), .IN2(n10436), .Q(n10950) );
  OR2X1 U10720 ( .IN1(n10951), .IN2(n10436), .Q(n10947) );
  OR2X1 U10721 ( .IN1(n10952), .IN2(n10953), .Q(n10951) );
  OR2X1 U10722 ( .IN1(n10457), .IN2(n10954), .Q(n10953) );
  AND2X1 U10723 ( .IN1(n10955), .IN2(n10436), .Q(n10954) );
  OR2X1 U10724 ( .IN1(n10956), .IN2(n10957), .Q(n10952) );
  AND2X1 U10725 ( .IN1(n10958), .IN2(n10446), .Q(n10957) );
  AND2X1 U10726 ( .IN1(n10959), .IN2(n10430), .Q(n10958) );
  OR2X1 U10727 ( .IN1(n10960), .IN2(n10443), .Q(n10959) );
  AND2X1 U10728 ( .IN1(n10433), .IN2(n10444), .Q(n10960) );
  AND2X1 U10729 ( .IN1(n10423), .IN2(n10961), .Q(n10956) );
  OR2X1 U10730 ( .IN1(n4386), .IN2(n10962), .Q(n10961) );
  OR2X1 U10731 ( .IN1(n10963), .IN2(n10964), .Q(g30304) );
  AND2X1 U10732 ( .IN1(n10965), .IN2(g2241), .Q(n10964) );
  AND2X1 U10733 ( .IN1(n4367), .IN2(g2285), .Q(n10963) );
  OR2X1 U10734 ( .IN1(n10966), .IN2(n10967), .Q(g30303) );
  AND2X1 U10735 ( .IN1(test_so73), .IN2(n10965), .Q(n10967) );
  AND2X1 U10736 ( .IN1(g2282), .IN2(n9119), .Q(n10966) );
  OR2X1 U10737 ( .IN1(n10968), .IN2(n10969), .Q(g30302) );
  AND2X1 U10738 ( .IN1(n10970), .IN2(g1547), .Q(n10969) );
  AND2X1 U10739 ( .IN1(n4368), .IN2(g1591), .Q(n10968) );
  OR2X1 U10740 ( .IN1(n10971), .IN2(n10972), .Q(g30301) );
  AND2X1 U10741 ( .IN1(n10965), .IN2(g6837), .Q(n10972) );
  OR2X1 U10742 ( .IN1(n10973), .IN2(n10974), .Q(n10965) );
  AND2X1 U10743 ( .IN1(n10534), .IN2(g2185), .Q(n10974) );
  AND2X1 U10744 ( .IN1(n10975), .IN2(n10536), .Q(n10973) );
  XNOR2X1 U10745 ( .IN1(n9652), .IN2(n10976), .Q(n10975) );
  AND2X1 U10746 ( .IN1(n4324), .IN2(g2279), .Q(n10971) );
  OR2X1 U10747 ( .IN1(n10977), .IN2(n10978), .Q(g30300) );
  AND2X1 U10748 ( .IN1(n10979), .IN2(g2241), .Q(n10978) );
  AND2X1 U10749 ( .IN1(n4367), .IN2(g2267), .Q(n10977) );
  OR2X1 U10750 ( .IN1(n10980), .IN2(n10981), .Q(g30299) );
  AND2X1 U10751 ( .IN1(n10970), .IN2(g6782), .Q(n10981) );
  AND2X1 U10752 ( .IN1(n4515), .IN2(g1588), .Q(n10980) );
  OR2X1 U10753 ( .IN1(n10982), .IN2(n10983), .Q(g30298) );
  AND2X1 U10754 ( .IN1(test_so31), .IN2(n10984), .Q(n10983) );
  AND2X1 U10755 ( .IN1(g897), .IN2(n9118), .Q(n10982) );
  OR2X1 U10756 ( .IN1(n10985), .IN2(n10986), .Q(g30297) );
  AND2X1 U10757 ( .IN1(n10987), .IN2(g2241), .Q(n10986) );
  AND2X1 U10758 ( .IN1(n4367), .IN2(g2339), .Q(n10985) );
  OR2X1 U10759 ( .IN1(n10988), .IN2(n10989), .Q(g30296) );
  AND2X1 U10760 ( .IN1(test_so73), .IN2(n10979), .Q(n10989) );
  AND2X1 U10761 ( .IN1(test_so76), .IN2(n9119), .Q(n10988) );
  OR2X1 U10762 ( .IN1(n10990), .IN2(n10991), .Q(g30295) );
  AND2X1 U10763 ( .IN1(n10970), .IN2(g6573), .Q(n10991) );
  OR2X1 U10764 ( .IN1(n10992), .IN2(n10993), .Q(n10970) );
  AND2X1 U10765 ( .IN1(n10564), .IN2(g1491), .Q(n10993) );
  AND2X1 U10766 ( .IN1(n10994), .IN2(n10566), .Q(n10992) );
  XNOR2X1 U10767 ( .IN1(n9623), .IN2(n10995), .Q(n10994) );
  AND2X1 U10768 ( .IN1(n4317), .IN2(g1585), .Q(n10990) );
  OR2X1 U10769 ( .IN1(n10996), .IN2(n10997), .Q(g30294) );
  AND2X1 U10770 ( .IN1(n10998), .IN2(g1547), .Q(n10997) );
  AND2X1 U10771 ( .IN1(n4368), .IN2(g1573), .Q(n10996) );
  OR2X1 U10772 ( .IN1(n10999), .IN2(n11000), .Q(g30293) );
  AND2X1 U10773 ( .IN1(n10984), .IN2(g6518), .Q(n11000) );
  AND2X1 U10774 ( .IN1(n4312), .IN2(g894), .Q(n10999) );
  OR2X1 U10775 ( .IN1(n11001), .IN2(n11002), .Q(g30292) );
  AND2X1 U10776 ( .IN1(n11003), .IN2(g165), .Q(n11002) );
  AND2X1 U10777 ( .IN1(n4369), .IN2(g210), .Q(n11001) );
  OR2X1 U10778 ( .IN1(n11004), .IN2(n11005), .Q(g30291) );
  AND2X1 U10779 ( .IN1(test_so73), .IN2(n10987), .Q(n11005) );
  AND2X1 U10780 ( .IN1(g2336), .IN2(n9119), .Q(n11004) );
  OR2X1 U10781 ( .IN1(n11006), .IN2(n11007), .Q(g30290) );
  AND2X1 U10782 ( .IN1(n11008), .IN2(g2241), .Q(n11007) );
  AND2X1 U10783 ( .IN1(n4367), .IN2(g2330), .Q(n11006) );
  OR2X1 U10784 ( .IN1(n11009), .IN2(n11010), .Q(g30289) );
  AND2X1 U10785 ( .IN1(n10979), .IN2(g6837), .Q(n11010) );
  OR2X1 U10786 ( .IN1(n11011), .IN2(n11012), .Q(n10979) );
  AND2X1 U10787 ( .IN1(n10534), .IN2(g2165), .Q(n11012) );
  AND2X1 U10788 ( .IN1(n10536), .IN2(n11013), .Q(n11011) );
  XNOR2X1 U10789 ( .IN1(n11014), .IN2(n9645), .Q(n11013) );
  AND2X1 U10790 ( .IN1(n4324), .IN2(g2261), .Q(n11009) );
  OR2X1 U10791 ( .IN1(n11015), .IN2(n11016), .Q(g30288) );
  AND2X1 U10792 ( .IN1(n11017), .IN2(g1547), .Q(n11016) );
  AND2X1 U10793 ( .IN1(n4368), .IN2(g1645), .Q(n11015) );
  OR2X1 U10794 ( .IN1(n11018), .IN2(n11019), .Q(g30287) );
  AND2X1 U10795 ( .IN1(n10998), .IN2(g6782), .Q(n11019) );
  AND2X1 U10796 ( .IN1(n4515), .IN2(g1570), .Q(n11018) );
  OR2X1 U10797 ( .IN1(n11020), .IN2(n11021), .Q(g30286) );
  AND2X1 U10798 ( .IN1(n10984), .IN2(g6368), .Q(n11021) );
  OR2X1 U10799 ( .IN1(n11022), .IN2(n11023), .Q(n10984) );
  AND2X1 U10800 ( .IN1(n10598), .IN2(g801), .Q(n11023) );
  AND2X1 U10801 ( .IN1(n11024), .IN2(n10600), .Q(n11022) );
  XNOR2X1 U10802 ( .IN1(n11025), .IN2(n9583), .Q(n11024) );
  AND2X1 U10803 ( .IN1(n4323), .IN2(g891), .Q(n11020) );
  OR2X1 U10804 ( .IN1(n11026), .IN2(n11027), .Q(g30285) );
  AND2X1 U10805 ( .IN1(test_so31), .IN2(n11028), .Q(n11027) );
  AND2X1 U10806 ( .IN1(g879), .IN2(n9118), .Q(n11026) );
  OR2X1 U10807 ( .IN1(n11029), .IN2(n11030), .Q(g30284) );
  AND2X1 U10808 ( .IN1(n11003), .IN2(g6313), .Q(n11030) );
  AND2X1 U10809 ( .IN1(n4512), .IN2(g207), .Q(n11029) );
  OR2X1 U10810 ( .IN1(n11031), .IN2(n11032), .Q(g30283) );
  AND2X1 U10811 ( .IN1(n10987), .IN2(g6837), .Q(n11032) );
  OR2X1 U10812 ( .IN1(n11033), .IN2(n11034), .Q(n10987) );
  AND2X1 U10813 ( .IN1(n10534), .IN2(g2200), .Q(n11034) );
  AND2X1 U10814 ( .IN1(n11035), .IN2(n11036), .Q(n11033) );
  XNOR2X1 U10815 ( .IN1(n10717), .IN2(n9638), .Q(n11036) );
  OR2X1 U10816 ( .IN1(n11037), .IN2(n11038), .Q(n10717) );
  XNOR2X1 U10817 ( .IN1(n4529), .IN2(n11039), .Q(n11037) );
  INVX0 U10818 ( .INP(n9653), .ZN(n11039) );
  AND2X1 U10819 ( .IN1(n4324), .IN2(g2333), .Q(n11031) );
  OR2X1 U10820 ( .IN1(n11040), .IN2(n11041), .Q(g30282) );
  AND2X1 U10821 ( .IN1(test_so73), .IN2(n11008), .Q(n11041) );
  AND2X1 U10822 ( .IN1(test_so77), .IN2(n9119), .Q(n11040) );
  OR2X1 U10823 ( .IN1(n11042), .IN2(n11043), .Q(g30281) );
  AND2X1 U10824 ( .IN1(n11017), .IN2(g6782), .Q(n11043) );
  AND2X1 U10825 ( .IN1(n4515), .IN2(g1642), .Q(n11042) );
  OR2X1 U10826 ( .IN1(n11044), .IN2(n11045), .Q(g30280) );
  AND2X1 U10827 ( .IN1(n11046), .IN2(g1547), .Q(n11045) );
  AND2X1 U10828 ( .IN1(n4368), .IN2(g1636), .Q(n11044) );
  OR2X1 U10829 ( .IN1(n11047), .IN2(n11048), .Q(g30279) );
  AND2X1 U10830 ( .IN1(n10998), .IN2(g6573), .Q(n11048) );
  OR2X1 U10831 ( .IN1(n11049), .IN2(n11050), .Q(n10998) );
  AND2X1 U10832 ( .IN1(n10564), .IN2(g1471), .Q(n11050) );
  AND2X1 U10833 ( .IN1(n10566), .IN2(n11051), .Q(n11049) );
  XNOR2X1 U10834 ( .IN1(n11052), .IN2(n9608), .Q(n11051) );
  AND2X1 U10835 ( .IN1(n4317), .IN2(g1567), .Q(n11047) );
  OR2X1 U10836 ( .IN1(n11053), .IN2(n11054), .Q(g30278) );
  AND2X1 U10837 ( .IN1(test_so31), .IN2(n11055), .Q(n11054) );
  AND2X1 U10838 ( .IN1(g951), .IN2(n9118), .Q(n11053) );
  OR2X1 U10839 ( .IN1(n11056), .IN2(n11057), .Q(g30277) );
  AND2X1 U10840 ( .IN1(n11028), .IN2(g6518), .Q(n11057) );
  AND2X1 U10841 ( .IN1(n4312), .IN2(g876), .Q(n11056) );
  OR2X1 U10842 ( .IN1(n11058), .IN2(n11059), .Q(g30276) );
  AND2X1 U10843 ( .IN1(n11003), .IN2(g6231), .Q(n11059) );
  OR2X1 U10844 ( .IN1(n11060), .IN2(n11061), .Q(n11003) );
  AND2X1 U10845 ( .IN1(n10638), .IN2(g113), .Q(n11061) );
  AND2X1 U10846 ( .IN1(n11062), .IN2(n10640), .Q(n11060) );
  XNOR2X1 U10847 ( .IN1(n9549), .IN2(n11063), .Q(n11062) );
  AND2X1 U10848 ( .IN1(n4318), .IN2(g204), .Q(n11058) );
  OR2X1 U10849 ( .IN1(n11064), .IN2(n11065), .Q(g30275) );
  AND2X1 U10850 ( .IN1(n11066), .IN2(g165), .Q(n11065) );
  AND2X1 U10851 ( .IN1(n4369), .IN2(g192), .Q(n11064) );
  OR2X1 U10852 ( .IN1(n11067), .IN2(n11068), .Q(g30274) );
  AND2X1 U10853 ( .IN1(n11008), .IN2(g6837), .Q(n11068) );
  OR2X1 U10854 ( .IN1(n11069), .IN2(n11070), .Q(n11008) );
  AND2X1 U10855 ( .IN1(n10534), .IN2(g2190), .Q(n11070) );
  AND2X1 U10856 ( .IN1(n11035), .IN2(n11071), .Q(n11069) );
  XNOR2X1 U10857 ( .IN1(n11072), .IN2(n11073), .Q(n11071) );
  AND2X1 U10858 ( .IN1(n11074), .IN2(n11075), .Q(n11073) );
  OR2X1 U10859 ( .IN1(n9652), .IN2(n10718), .Q(n11075) );
  INVX0 U10860 ( .INP(n11076), .ZN(n11074) );
  AND2X1 U10861 ( .IN1(n10536), .IN2(n10720), .Q(n11035) );
  AND2X1 U10862 ( .IN1(n4324), .IN2(g2324), .Q(n11067) );
  OR2X1 U10863 ( .IN1(n11077), .IN2(n11078), .Q(g30273) );
  AND2X1 U10864 ( .IN1(n11017), .IN2(g6573), .Q(n11078) );
  OR2X1 U10865 ( .IN1(n11079), .IN2(n11080), .Q(n11017) );
  AND2X1 U10866 ( .IN1(n10564), .IN2(g1506), .Q(n11080) );
  AND2X1 U10867 ( .IN1(n11081), .IN2(n11082), .Q(n11079) );
  XNOR2X1 U10868 ( .IN1(n10764), .IN2(n9603), .Q(n11082) );
  OR2X1 U10869 ( .IN1(n11083), .IN2(n11084), .Q(n10764) );
  XNOR2X1 U10870 ( .IN1(n4530), .IN2(n11085), .Q(n11083) );
  INVX0 U10871 ( .INP(n9619), .ZN(n11085) );
  AND2X1 U10872 ( .IN1(n4317), .IN2(g1639), .Q(n11077) );
  OR2X1 U10873 ( .IN1(n11086), .IN2(n11087), .Q(g30272) );
  AND2X1 U10874 ( .IN1(n11046), .IN2(g6782), .Q(n11087) );
  AND2X1 U10875 ( .IN1(n4515), .IN2(g1633), .Q(n11086) );
  OR2X1 U10876 ( .IN1(n11088), .IN2(n11089), .Q(g30271) );
  AND2X1 U10877 ( .IN1(n11055), .IN2(g6518), .Q(n11089) );
  AND2X1 U10878 ( .IN1(n4312), .IN2(g948), .Q(n11088) );
  OR2X1 U10879 ( .IN1(n11090), .IN2(n11091), .Q(g30270) );
  AND2X1 U10880 ( .IN1(test_so31), .IN2(n11092), .Q(n11091) );
  AND2X1 U10881 ( .IN1(g942), .IN2(n9118), .Q(n11090) );
  OR2X1 U10882 ( .IN1(n11093), .IN2(n11094), .Q(g30269) );
  AND2X1 U10883 ( .IN1(n11028), .IN2(g6368), .Q(n11094) );
  OR2X1 U10884 ( .IN1(n11095), .IN2(n11096), .Q(n11028) );
  AND2X1 U10885 ( .IN1(n10598), .IN2(g785), .Q(n11096) );
  AND2X1 U10886 ( .IN1(n10600), .IN2(n11097), .Q(n11095) );
  XNOR2X1 U10887 ( .IN1(n11098), .IN2(n9576), .Q(n11097) );
  AND2X1 U10888 ( .IN1(n4323), .IN2(g873), .Q(n11093) );
  OR2X1 U10889 ( .IN1(n11099), .IN2(n11100), .Q(g30268) );
  AND2X1 U10890 ( .IN1(n11101), .IN2(g165), .Q(n11100) );
  AND2X1 U10891 ( .IN1(n4369), .IN2(g264), .Q(n11099) );
  OR2X1 U10892 ( .IN1(n11102), .IN2(n11103), .Q(g30267) );
  AND2X1 U10893 ( .IN1(n11066), .IN2(g6313), .Q(n11103) );
  AND2X1 U10894 ( .IN1(test_so13), .IN2(n4512), .Q(n11102) );
  OR2X1 U10895 ( .IN1(n11104), .IN2(n11105), .Q(g30266) );
  AND2X1 U10896 ( .IN1(n11046), .IN2(g6573), .Q(n11105) );
  OR2X1 U10897 ( .IN1(n11106), .IN2(n11107), .Q(n11046) );
  AND2X1 U10898 ( .IN1(n10564), .IN2(g1496), .Q(n11107) );
  AND2X1 U10899 ( .IN1(n11081), .IN2(n11108), .Q(n11106) );
  XNOR2X1 U10900 ( .IN1(n11109), .IN2(n11110), .Q(n11108) );
  AND2X1 U10901 ( .IN1(n11111), .IN2(n11112), .Q(n11110) );
  OR2X1 U10902 ( .IN1(n9623), .IN2(n10765), .Q(n11112) );
  INVX0 U10903 ( .INP(n11113), .ZN(n11111) );
  AND2X1 U10904 ( .IN1(n10566), .IN2(n10767), .Q(n11081) );
  AND2X1 U10905 ( .IN1(n4317), .IN2(g1630), .Q(n11104) );
  OR2X1 U10906 ( .IN1(n11114), .IN2(n11115), .Q(g30265) );
  AND2X1 U10907 ( .IN1(n11055), .IN2(g6368), .Q(n11115) );
  OR2X1 U10908 ( .IN1(n11116), .IN2(n11117), .Q(n11055) );
  AND2X1 U10909 ( .IN1(n10598), .IN2(g813), .Q(n11117) );
  AND2X1 U10910 ( .IN1(n11118), .IN2(n10600), .Q(n11116) );
  XNOR2X1 U10911 ( .IN1(n11119), .IN2(n9589), .Q(n11118) );
  OR2X1 U10912 ( .IN1(n11120), .IN2(n10802), .Q(n11119) );
  OR2X1 U10913 ( .IN1(n11121), .IN2(n11122), .Q(n10802) );
  AND2X1 U10914 ( .IN1(n10743), .IN2(n9574), .Q(n11121) );
  AND2X1 U10915 ( .IN1(n10627), .IN2(n10807), .Q(n11120) );
  INVX0 U10916 ( .INP(n9574), .ZN(n10807) );
  AND2X1 U10917 ( .IN1(test_so35), .IN2(n4323), .Q(n11114) );
  OR2X1 U10918 ( .IN1(n11123), .IN2(n11124), .Q(g30264) );
  AND2X1 U10919 ( .IN1(n11092), .IN2(g6518), .Q(n11124) );
  AND2X1 U10920 ( .IN1(n4312), .IN2(g939), .Q(n11123) );
  OR2X1 U10921 ( .IN1(n11125), .IN2(n11126), .Q(g30263) );
  AND2X1 U10922 ( .IN1(n11101), .IN2(g6313), .Q(n11126) );
  AND2X1 U10923 ( .IN1(n4512), .IN2(g261), .Q(n11125) );
  OR2X1 U10924 ( .IN1(n11127), .IN2(n11128), .Q(g30262) );
  AND2X1 U10925 ( .IN1(n11129), .IN2(g165), .Q(n11128) );
  AND2X1 U10926 ( .IN1(n4369), .IN2(test_so14), .Q(n11127) );
  OR2X1 U10927 ( .IN1(n11130), .IN2(n11131), .Q(g30261) );
  AND2X1 U10928 ( .IN1(n11066), .IN2(g6231), .Q(n11131) );
  OR2X1 U10929 ( .IN1(n11132), .IN2(n11133), .Q(n11066) );
  AND2X1 U10930 ( .IN1(n10638), .IN2(g97), .Q(n11133) );
  AND2X1 U10931 ( .IN1(n10640), .IN2(n11134), .Q(n11132) );
  XNOR2X1 U10932 ( .IN1(n11135), .IN2(n9547), .Q(n11134) );
  AND2X1 U10933 ( .IN1(n4318), .IN2(g186), .Q(n11130) );
  OR2X1 U10934 ( .IN1(n11136), .IN2(n11137), .Q(g30260) );
  AND2X1 U10935 ( .IN1(n11138), .IN2(g2241), .Q(n11137) );
  AND2X1 U10936 ( .IN1(n4367), .IN2(g2294), .Q(n11136) );
  OR2X1 U10937 ( .IN1(n11139), .IN2(n11140), .Q(g30259) );
  AND2X1 U10938 ( .IN1(n11092), .IN2(g6368), .Q(n11140) );
  OR2X1 U10939 ( .IN1(n11141), .IN2(n11142), .Q(n11092) );
  AND2X1 U10940 ( .IN1(n10598), .IN2(g805), .Q(n11142) );
  AND2X1 U10941 ( .IN1(n11143), .IN2(n10600), .Q(n11141) );
  XNOR2X1 U10942 ( .IN1(n11144), .IN2(n9568), .Q(n11143) );
  OR2X1 U10943 ( .IN1(n11145), .IN2(n11146), .Q(n11144) );
  AND2X1 U10944 ( .IN1(n10627), .IN2(n11147), .Q(n11145) );
  AND2X1 U10945 ( .IN1(n4323), .IN2(g936), .Q(n11139) );
  OR2X1 U10946 ( .IN1(n11148), .IN2(n11149), .Q(g30258) );
  AND2X1 U10947 ( .IN1(n11101), .IN2(g6231), .Q(n11149) );
  OR2X1 U10948 ( .IN1(n11150), .IN2(n11151), .Q(n11101) );
  AND2X1 U10949 ( .IN1(n10638), .IN2(g125), .Q(n11151) );
  AND2X1 U10950 ( .IN1(n11152), .IN2(n10640), .Q(n11150) );
  XNOR2X1 U10951 ( .IN1(n10827), .IN2(n9533), .Q(n11152) );
  OR2X1 U10952 ( .IN1(n11153), .IN2(n11154), .Q(n10827) );
  XNOR2X1 U10953 ( .IN1(n10252), .IN2(n11155), .Q(n11153) );
  INVX0 U10954 ( .INP(n9538), .ZN(n11155) );
  AND2X1 U10955 ( .IN1(n4318), .IN2(g258), .Q(n11148) );
  OR2X1 U10956 ( .IN1(n11156), .IN2(n11157), .Q(g30257) );
  AND2X1 U10957 ( .IN1(n11129), .IN2(g6313), .Q(n11157) );
  AND2X1 U10958 ( .IN1(n4512), .IN2(g252), .Q(n11156) );
  OR2X1 U10959 ( .IN1(n11158), .IN2(n11159), .Q(g30256) );
  AND2X1 U10960 ( .IN1(test_so73), .IN2(n11138), .Q(n11159) );
  AND2X1 U10961 ( .IN1(g2291), .IN2(n9119), .Q(n11158) );
  OR2X1 U10962 ( .IN1(n11160), .IN2(n11161), .Q(g30255) );
  AND2X1 U10963 ( .IN1(n11162), .IN2(g1547), .Q(n11161) );
  AND2X1 U10964 ( .IN1(n4368), .IN2(g1600), .Q(n11160) );
  OR2X1 U10965 ( .IN1(n11163), .IN2(n11164), .Q(g30254) );
  AND2X1 U10966 ( .IN1(n11129), .IN2(g6231), .Q(n11164) );
  OR2X1 U10967 ( .IN1(n11165), .IN2(n11166), .Q(n11129) );
  AND2X1 U10968 ( .IN1(n10638), .IN2(g117), .Q(n11166) );
  AND2X1 U10969 ( .IN1(n11167), .IN2(n10640), .Q(n11165) );
  XNOR2X1 U10970 ( .IN1(n11168), .IN2(n11169), .Q(n11167) );
  AND2X1 U10971 ( .IN1(n11170), .IN2(n11171), .Q(n11169) );
  OR2X1 U10972 ( .IN1(n9549), .IN2(n10829), .Q(n11171) );
  INVX0 U10973 ( .INP(n11172), .ZN(n11170) );
  AND2X1 U10974 ( .IN1(n4318), .IN2(g249), .Q(n11163) );
  OR2X1 U10975 ( .IN1(n11173), .IN2(n11174), .Q(g30253) );
  AND2X1 U10976 ( .IN1(n11138), .IN2(g6837), .Q(n11174) );
  OR2X1 U10977 ( .IN1(n11175), .IN2(n11176), .Q(n11138) );
  AND2X1 U10978 ( .IN1(n10534), .IN2(g2195), .Q(n11176) );
  AND2X1 U10979 ( .IN1(n10720), .IN2(n11177), .Q(n10534) );
  INVX0 U10980 ( .INP(n10536), .ZN(n11177) );
  OR2X1 U10981 ( .IN1(n11178), .IN2(n11179), .Q(n10720) );
  INVX0 U10982 ( .INP(n11180), .ZN(n11179) );
  AND2X1 U10983 ( .IN1(n11181), .IN2(n10536), .Q(n11175) );
  AND2X1 U10984 ( .IN1(n11182), .IN2(n11180), .Q(n10536) );
  AND2X1 U10985 ( .IN1(n11183), .IN2(n11184), .Q(n11180) );
  AND2X1 U10986 ( .IN1(n10834), .IN2(n11185), .Q(n11184) );
  OR2X1 U10987 ( .IN1(n11186), .IN2(n10871), .Q(n11185) );
  AND2X1 U10988 ( .IN1(n11187), .IN2(n10844), .Q(n11186) );
  OR2X1 U10989 ( .IN1(n10855), .IN2(n10860), .Q(n11187) );
  OR2X1 U10990 ( .IN1(n10848), .IN2(n11188), .Q(n10855) );
  OR2X1 U10991 ( .IN1(n11189), .IN2(n10848), .Q(n11183) );
  OR2X1 U10992 ( .IN1(n11190), .IN2(n11191), .Q(n10848) );
  AND2X1 U10993 ( .IN1(n11192), .IN2(n11193), .Q(n11190) );
  OR2X1 U10994 ( .IN1(n4524), .IN2(g2398), .Q(n11193) );
  AND2X1 U10995 ( .IN1(n11194), .IN2(n11195), .Q(n11192) );
  OR2X1 U10996 ( .IN1(n4516), .IN2(g2397), .Q(n11195) );
  OR2X1 U10997 ( .IN1(n4509), .IN2(g2396), .Q(n11194) );
  OR2X1 U10998 ( .IN1(n11178), .IN2(n11196), .Q(n11182) );
  AND2X1 U10999 ( .IN1(n11197), .IN2(n4529), .Q(n11196) );
  OR2X1 U11000 ( .IN1(n11198), .IN2(n11014), .Q(n11178) );
  AND2X1 U11001 ( .IN1(n11197), .IN2(n2489), .Q(n11198) );
  OR2X1 U11002 ( .IN1(n11199), .IN2(n11200), .Q(n2489) );
  OR2X1 U11003 ( .IN1(n11201), .IN2(n11202), .Q(n11200) );
  OR2X1 U11004 ( .IN1(n9643), .IN2(n9636), .Q(n11202) );
  OR2X1 U11005 ( .IN1(n9644), .IN2(n11203), .Q(n11199) );
  OR2X1 U11006 ( .IN1(n11204), .IN2(n9654), .Q(n11203) );
  OR2X1 U11007 ( .IN1(n11205), .IN2(n11206), .Q(n11197) );
  OR2X1 U11008 ( .IN1(n10719), .IN2(n11207), .Q(n11206) );
  OR2X1 U11009 ( .IN1(n10538), .IN2(n11201), .Q(n11207) );
  OR2X1 U11010 ( .IN1(n11208), .IN2(n11209), .Q(n11201) );
  OR2X1 U11011 ( .IN1(n9637), .IN2(n9638), .Q(n11209) );
  OR2X1 U11012 ( .IN1(n9645), .IN2(n11210), .Q(n11208) );
  OR2X1 U11013 ( .IN1(n9653), .IN2(n9652), .Q(n11210) );
  INVX0 U11014 ( .INP(n4529), .ZN(n10719) );
  INVX0 U11015 ( .INP(n11211), .ZN(n11205) );
  AND2X1 U11016 ( .IN1(n11212), .IN2(n11213), .Q(n11211) );
  AND2X1 U11017 ( .IN1(n9644), .IN2(n9643), .Q(n11213) );
  AND2X1 U11018 ( .IN1(n11204), .IN2(n9636), .Q(n11212) );
  XNOR2X1 U11019 ( .IN1(n11038), .IN2(n9653), .Q(n11181) );
  OR2X1 U11020 ( .IN1(n11076), .IN2(n11214), .Q(n11038) );
  OR2X1 U11021 ( .IN1(n11215), .IN2(n11216), .Q(n11214) );
  AND2X1 U11022 ( .IN1(n4529), .IN2(n11072), .Q(n11216) );
  INVX0 U11023 ( .INP(n9637), .ZN(n11072) );
  AND2X1 U11024 ( .IN1(n11217), .IN2(n9637), .Q(n11215) );
  INVX0 U11025 ( .INP(n9652), .ZN(n11217) );
  OR2X1 U11026 ( .IN1(n11218), .IN2(n10976), .Q(n11076) );
  OR2X1 U11027 ( .IN1(n11219), .IN2(n11220), .Q(n10976) );
  OR2X1 U11028 ( .IN1(n11221), .IN2(n10652), .Q(n11220) );
  OR2X1 U11029 ( .IN1(n11222), .IN2(n10682), .Q(n10652) );
  OR2X1 U11030 ( .IN1(n11014), .IN2(n11223), .Q(n10682) );
  XNOR2X1 U11031 ( .IN1(n4529), .IN2(n11224), .Q(n11223) );
  INVX0 U11032 ( .INP(n9645), .ZN(n11224) );
  AND2X1 U11033 ( .IN1(n9659), .IN2(n10718), .Q(n11014) );
  XNOR2X1 U11034 ( .IN1(n4529), .IN2(n9658), .Q(n11222) );
  AND2X1 U11035 ( .IN1(n4529), .IN2(n11225), .Q(n11221) );
  OR2X1 U11036 ( .IN1(n11226), .IN2(n11227), .Q(n11219) );
  AND2X1 U11037 ( .IN1(n10538), .IN2(n9644), .Q(n11227) );
  INVX0 U11038 ( .INP(n9654), .ZN(n10538) );
  AND2X1 U11039 ( .IN1(n10718), .IN2(n9654), .Q(n11226) );
  AND2X1 U11040 ( .IN1(n10718), .IN2(n9652), .Q(n11218) );
  AND2X1 U11041 ( .IN1(n4324), .IN2(g2288), .Q(n11173) );
  OR2X1 U11042 ( .IN1(n11228), .IN2(n11229), .Q(g30252) );
  AND2X1 U11043 ( .IN1(n11162), .IN2(g6782), .Q(n11229) );
  AND2X1 U11044 ( .IN1(n4515), .IN2(g1597), .Q(n11228) );
  OR2X1 U11045 ( .IN1(n11230), .IN2(n11231), .Q(g30251) );
  AND2X1 U11046 ( .IN1(test_so31), .IN2(n11232), .Q(n11231) );
  AND2X1 U11047 ( .IN1(g906), .IN2(n9118), .Q(n11230) );
  OR2X1 U11048 ( .IN1(n11233), .IN2(n11234), .Q(g30250) );
  AND2X1 U11049 ( .IN1(n11162), .IN2(g6573), .Q(n11234) );
  OR2X1 U11050 ( .IN1(n11235), .IN2(n11236), .Q(n11162) );
  AND2X1 U11051 ( .IN1(n10564), .IN2(g1501), .Q(n11236) );
  AND2X1 U11052 ( .IN1(n10767), .IN2(n11237), .Q(n10564) );
  INVX0 U11053 ( .INP(n10566), .ZN(n11237) );
  OR2X1 U11054 ( .IN1(n11238), .IN2(n11239), .Q(n10767) );
  INVX0 U11055 ( .INP(n11240), .ZN(n11239) );
  AND2X1 U11056 ( .IN1(n11241), .IN2(n10566), .Q(n11235) );
  AND2X1 U11057 ( .IN1(n11242), .IN2(n11240), .Q(n10566) );
  AND2X1 U11058 ( .IN1(n11243), .IN2(n11244), .Q(n11240) );
  AND2X1 U11059 ( .IN1(n10420), .IN2(n11245), .Q(n11244) );
  OR2X1 U11060 ( .IN1(n11246), .IN2(n10457), .Q(n11245) );
  AND2X1 U11061 ( .IN1(n11247), .IN2(n10430), .Q(n11246) );
  OR2X1 U11062 ( .IN1(n10441), .IN2(n10446), .Q(n11247) );
  OR2X1 U11063 ( .IN1(n10434), .IN2(n11248), .Q(n10441) );
  OR2X1 U11064 ( .IN1(n11249), .IN2(n10434), .Q(n11243) );
  OR2X1 U11065 ( .IN1(n11250), .IN2(n11251), .Q(n10434) );
  AND2X1 U11066 ( .IN1(n11252), .IN2(n11253), .Q(n11250) );
  OR2X1 U11067 ( .IN1(n4525), .IN2(g1704), .Q(n11253) );
  AND2X1 U11068 ( .IN1(n11254), .IN2(n11255), .Q(n11252) );
  OR2X1 U11069 ( .IN1(n4518), .IN2(g1703), .Q(n11255) );
  OR2X1 U11070 ( .IN1(n4511), .IN2(g1702), .Q(n11254) );
  OR2X1 U11071 ( .IN1(n11238), .IN2(n11256), .Q(n11242) );
  AND2X1 U11072 ( .IN1(n11257), .IN2(n4530), .Q(n11256) );
  OR2X1 U11073 ( .IN1(n11258), .IN2(n11052), .Q(n11238) );
  AND2X1 U11074 ( .IN1(n11257), .IN2(n9624), .Q(n11258) );
  OR2X1 U11075 ( .IN1(n11259), .IN2(n11260), .Q(n9624) );
  OR2X1 U11076 ( .IN1(n11261), .IN2(n11262), .Q(n11260) );
  OR2X1 U11077 ( .IN1(n9610), .IN2(n9601), .Q(n11262) );
  OR2X1 U11078 ( .IN1(n9609), .IN2(n11263), .Q(n11259) );
  OR2X1 U11079 ( .IN1(n9618), .IN2(n9617), .Q(n11263) );
  OR2X1 U11080 ( .IN1(n11264), .IN2(n11265), .Q(n11257) );
  OR2X1 U11081 ( .IN1(n10766), .IN2(n11266), .Q(n11265) );
  OR2X1 U11082 ( .IN1(n10568), .IN2(n11261), .Q(n11266) );
  OR2X1 U11083 ( .IN1(n11267), .IN2(n11268), .Q(n11261) );
  OR2X1 U11084 ( .IN1(n9602), .IN2(n9603), .Q(n11268) );
  OR2X1 U11085 ( .IN1(n9608), .IN2(n11269), .Q(n11267) );
  OR2X1 U11086 ( .IN1(n9623), .IN2(n9619), .Q(n11269) );
  INVX0 U11087 ( .INP(n4530), .ZN(n10766) );
  OR2X1 U11088 ( .IN1(n11270), .IN2(n11271), .Q(n11264) );
  OR2X1 U11089 ( .IN1(n11272), .IN2(n10762), .Q(n11271) );
  INVX0 U11090 ( .INP(n9618), .ZN(n10762) );
  OR2X1 U11091 ( .IN1(n10729), .IN2(n10588), .Q(n11270) );
  XNOR2X1 U11092 ( .IN1(n11084), .IN2(n9619), .Q(n11241) );
  OR2X1 U11093 ( .IN1(n11113), .IN2(n11273), .Q(n11084) );
  OR2X1 U11094 ( .IN1(n11274), .IN2(n11275), .Q(n11273) );
  AND2X1 U11095 ( .IN1(n4530), .IN2(n11109), .Q(n11275) );
  INVX0 U11096 ( .INP(n9602), .ZN(n11109) );
  AND2X1 U11097 ( .IN1(n11276), .IN2(n9602), .Q(n11274) );
  INVX0 U11098 ( .INP(n9623), .ZN(n11276) );
  OR2X1 U11099 ( .IN1(n11277), .IN2(n10995), .Q(n11113) );
  OR2X1 U11100 ( .IN1(n11278), .IN2(n11279), .Q(n10995) );
  OR2X1 U11101 ( .IN1(n11280), .IN2(n10695), .Q(n11279) );
  OR2X1 U11102 ( .IN1(n11281), .IN2(n10728), .Q(n10695) );
  OR2X1 U11103 ( .IN1(n11052), .IN2(n11282), .Q(n10728) );
  XNOR2X1 U11104 ( .IN1(n4530), .IN2(n11283), .Q(n11282) );
  INVX0 U11105 ( .INP(n9608), .ZN(n11283) );
  AND2X1 U11106 ( .IN1(n9625), .IN2(n10765), .Q(n11052) );
  XNOR2X1 U11107 ( .IN1(n4530), .IN2(n10729), .Q(n11281) );
  INVX0 U11108 ( .INP(n9601), .ZN(n10729) );
  AND2X1 U11109 ( .IN1(n4530), .IN2(n11272), .Q(n11280) );
  INVX0 U11110 ( .INP(n9610), .ZN(n11272) );
  OR2X1 U11111 ( .IN1(n11284), .IN2(n11285), .Q(n11278) );
  AND2X1 U11112 ( .IN1(n10568), .IN2(n9610), .Q(n11285) );
  INVX0 U11113 ( .INP(n9617), .ZN(n10568) );
  AND2X1 U11114 ( .IN1(n10765), .IN2(n9617), .Q(n11284) );
  AND2X1 U11115 ( .IN1(n10765), .IN2(n9623), .Q(n11277) );
  AND2X1 U11116 ( .IN1(n4317), .IN2(g1594), .Q(n11233) );
  OR2X1 U11117 ( .IN1(n11286), .IN2(n11287), .Q(g30249) );
  AND2X1 U11118 ( .IN1(n11232), .IN2(g6518), .Q(n11287) );
  AND2X1 U11119 ( .IN1(n4312), .IN2(g903), .Q(n11286) );
  OR2X1 U11120 ( .IN1(n11288), .IN2(n11289), .Q(g30248) );
  AND2X1 U11121 ( .IN1(n11290), .IN2(g165), .Q(n11289) );
  AND2X1 U11122 ( .IN1(n4369), .IN2(g219), .Q(n11288) );
  OR2X1 U11123 ( .IN1(n11291), .IN2(n11292), .Q(g30247) );
  AND2X1 U11124 ( .IN1(n11232), .IN2(g6368), .Q(n11292) );
  OR2X1 U11125 ( .IN1(n11293), .IN2(n11294), .Q(n11232) );
  AND2X1 U11126 ( .IN1(n10598), .IN2(g809), .Q(n11294) );
  INVX0 U11127 ( .INP(n11295), .ZN(n10598) );
  OR2X1 U11128 ( .IN1(n10777), .IN2(n10600), .Q(n11295) );
  AND2X1 U11129 ( .IN1(n11296), .IN2(n11297), .Q(n10777) );
  INVX0 U11130 ( .INP(n11298), .ZN(n11297) );
  OR2X1 U11131 ( .IN1(n11098), .IN2(n11299), .Q(n11298) );
  AND2X1 U11132 ( .IN1(n2542), .IN2(n11300), .Q(n11299) );
  AND2X1 U11133 ( .IN1(n11301), .IN2(n10600), .Q(n11293) );
  AND2X1 U11134 ( .IN1(n11302), .IN2(n11296), .Q(n10600) );
  AND2X1 U11135 ( .IN1(n11303), .IN2(n11304), .Q(n11296) );
  AND2X1 U11136 ( .IN1(n10253), .IN2(n11305), .Q(n11304) );
  OR2X1 U11137 ( .IN1(n11306), .IN2(n10236), .Q(n11305) );
  AND2X1 U11138 ( .IN1(n11307), .IN2(n10245), .Q(n11306) );
  OR2X1 U11139 ( .IN1(n10268), .IN2(n10243), .Q(n11307) );
  OR2X1 U11140 ( .IN1(n11308), .IN2(n10263), .Q(n10268) );
  OR2X1 U11141 ( .IN1(n11309), .IN2(n10263), .Q(n11303) );
  OR2X1 U11142 ( .IN1(n11310), .IN2(n11311), .Q(n10263) );
  AND2X1 U11143 ( .IN1(n11312), .IN2(n11313), .Q(n11310) );
  OR2X1 U11144 ( .IN1(n4364), .IN2(g1010), .Q(n11313) );
  AND2X1 U11145 ( .IN1(n11314), .IN2(n11315), .Q(n11312) );
  OR2X1 U11146 ( .IN1(n4363), .IN2(g1009), .Q(n11315) );
  OR2X1 U11147 ( .IN1(n4381), .IN2(g1008), .Q(n11314) );
  OR2X1 U11148 ( .IN1(n11098), .IN2(n11316), .Q(n11302) );
  AND2X1 U11149 ( .IN1(n11300), .IN2(n11317), .Q(n11316) );
  OR2X1 U11150 ( .IN1(n10627), .IN2(n2542), .Q(n11317) );
  OR2X1 U11151 ( .IN1(n11318), .IN2(n11319), .Q(n2542) );
  OR2X1 U11152 ( .IN1(n11320), .IN2(n11321), .Q(n11319) );
  OR2X1 U11153 ( .IN1(n9567), .IN2(n9569), .Q(n11321) );
  OR2X1 U11154 ( .IN1(n10623), .IN2(n11322), .Q(n11318) );
  OR2X1 U11155 ( .IN1(n9584), .IN2(n9585), .Q(n11322) );
  OR2X1 U11156 ( .IN1(n11323), .IN2(n11324), .Q(n11300) );
  OR2X1 U11157 ( .IN1(n10743), .IN2(n11325), .Q(n11324) );
  OR2X1 U11158 ( .IN1(n11326), .IN2(n11320), .Q(n11325) );
  OR2X1 U11159 ( .IN1(n11327), .IN2(n11328), .Q(n11320) );
  OR2X1 U11160 ( .IN1(n9576), .IN2(n9568), .Q(n11328) );
  OR2X1 U11161 ( .IN1(n9574), .IN2(n11329), .Q(n11327) );
  OR2X1 U11162 ( .IN1(n9589), .IN2(n9583), .Q(n11329) );
  OR2X1 U11163 ( .IN1(n11330), .IN2(n11331), .Q(n11323) );
  OR2X1 U11164 ( .IN1(n9575), .IN2(n10628), .Q(n11331) );
  INVX0 U11165 ( .INP(n9584), .ZN(n10628) );
  OR2X1 U11166 ( .IN1(n10776), .IN2(n11332), .Q(n11330) );
  XNOR2X1 U11167 ( .IN1(n11122), .IN2(n9574), .Q(n11301) );
  OR2X1 U11168 ( .IN1(n11146), .IN2(n11333), .Q(n11122) );
  OR2X1 U11169 ( .IN1(n11334), .IN2(n11335), .Q(n11333) );
  INVX0 U11170 ( .INP(n11336), .ZN(n11335) );
  OR2X1 U11171 ( .IN1(n10743), .IN2(n9568), .Q(n11336) );
  AND2X1 U11172 ( .IN1(n11147), .IN2(n9568), .Q(n11334) );
  OR2X1 U11173 ( .IN1(n11337), .IN2(n11025), .Q(n11146) );
  OR2X1 U11174 ( .IN1(n10744), .IN2(n11338), .Q(n11025) );
  OR2X1 U11175 ( .IN1(n11339), .IN2(n11340), .Q(n11338) );
  AND2X1 U11176 ( .IN1(n10627), .IN2(n11332), .Q(n11340) );
  INVX0 U11177 ( .INP(n9567), .ZN(n11332) );
  AND2X1 U11178 ( .IN1(n11326), .IN2(n9567), .Q(n11339) );
  OR2X1 U11179 ( .IN1(n11341), .IN2(n10601), .Q(n10744) );
  OR2X1 U11180 ( .IN1(n11342), .IN2(n10775), .Q(n10601) );
  OR2X1 U11181 ( .IN1(n11098), .IN2(n11343), .Q(n10775) );
  XNOR2X1 U11182 ( .IN1(n10627), .IN2(n11344), .Q(n11343) );
  AND2X1 U11183 ( .IN1(n9590), .IN2(n10743), .Q(n11098) );
  XNOR2X1 U11184 ( .IN1(n10627), .IN2(n10776), .Q(n11342) );
  INVX0 U11185 ( .INP(n9569), .ZN(n10776) );
  AND2X1 U11186 ( .IN1(n10743), .IN2(n9585), .Q(n11341) );
  AND2X1 U11187 ( .IN1(n10743), .IN2(n9583), .Q(n11337) );
  AND2X1 U11188 ( .IN1(n4323), .IN2(g900), .Q(n11291) );
  OR2X1 U11189 ( .IN1(n11345), .IN2(n11346), .Q(g30246) );
  AND2X1 U11190 ( .IN1(n11290), .IN2(g6313), .Q(n11346) );
  AND2X1 U11191 ( .IN1(n4512), .IN2(g216), .Q(n11345) );
  OR2X1 U11192 ( .IN1(n11347), .IN2(n11348), .Q(g30245) );
  AND2X1 U11193 ( .IN1(n11290), .IN2(g6231), .Q(n11348) );
  OR2X1 U11194 ( .IN1(n11349), .IN2(n11350), .Q(n11290) );
  AND2X1 U11195 ( .IN1(n10638), .IN2(g121), .Q(n11350) );
  INVX0 U11196 ( .INP(n11351), .ZN(n10638) );
  OR2X1 U11197 ( .IN1(n10816), .IN2(n10640), .Q(n11351) );
  AND2X1 U11198 ( .IN1(n11352), .IN2(n11353), .Q(n10816) );
  INVX0 U11199 ( .INP(n11354), .ZN(n11352) );
  AND2X1 U11200 ( .IN1(n11355), .IN2(n10640), .Q(n11349) );
  AND2X1 U11201 ( .IN1(n11356), .IN2(n11353), .Q(n10640) );
  AND2X1 U11202 ( .IN1(n11357), .IN2(n11358), .Q(n11353) );
  AND2X1 U11203 ( .IN1(n10476), .IN2(n11359), .Q(n11358) );
  OR2X1 U11204 ( .IN1(n11360), .IN2(n10513), .Q(n11359) );
  AND2X1 U11205 ( .IN1(n11361), .IN2(n10486), .Q(n11360) );
  OR2X1 U11206 ( .IN1(n10497), .IN2(n10502), .Q(n11361) );
  OR2X1 U11207 ( .IN1(n10490), .IN2(n11362), .Q(n10497) );
  OR2X1 U11208 ( .IN1(n11363), .IN2(n10490), .Q(n11357) );
  OR2X1 U11209 ( .IN1(n11364), .IN2(n11365), .Q(n10490) );
  AND2X1 U11210 ( .IN1(n11366), .IN2(n11367), .Q(n11364) );
  OR2X1 U11211 ( .IN1(n4499), .IN2(g323), .Q(n11367) );
  AND2X1 U11212 ( .IN1(n11368), .IN2(n11369), .Q(n11366) );
  OR2X1 U11213 ( .IN1(n4520), .IN2(g322), .Q(n11369) );
  OR2X1 U11214 ( .IN1(n4506), .IN2(g321), .Q(n11368) );
  OR2X1 U11215 ( .IN1(n11354), .IN2(n11370), .Q(n11356) );
  AND2X1 U11216 ( .IN1(n11371), .IN2(n10252), .Q(n11370) );
  OR2X1 U11217 ( .IN1(n11372), .IN2(n11135), .Q(n11354) );
  AND2X1 U11218 ( .IN1(n11371), .IN2(n9555), .Q(n11372) );
  OR2X1 U11219 ( .IN1(n11373), .IN2(n11374), .Q(n9555) );
  OR2X1 U11220 ( .IN1(n11375), .IN2(n11376), .Q(n11374) );
  OR2X1 U11221 ( .IN1(n9540), .IN2(n9531), .Q(n11376) );
  OR2X1 U11222 ( .IN1(n9539), .IN2(n11377), .Q(n11373) );
  OR2X1 U11223 ( .IN1(n9554), .IN2(n9548), .Q(n11377) );
  OR2X1 U11224 ( .IN1(n11378), .IN2(n11379), .Q(n11371) );
  OR2X1 U11225 ( .IN1(n10829), .IN2(n11380), .Q(n11379) );
  OR2X1 U11226 ( .IN1(n10642), .IN2(n11375), .Q(n11380) );
  OR2X1 U11227 ( .IN1(n11381), .IN2(n11382), .Q(n11375) );
  INVX0 U11228 ( .INP(n11383), .ZN(n11382) );
  AND2X1 U11229 ( .IN1(n10828), .IN2(n4513), .Q(n11383) );
  INVX0 U11230 ( .INP(n9533), .ZN(n10828) );
  OR2X1 U11231 ( .IN1(n9532), .IN2(n11384), .Q(n11381) );
  OR2X1 U11232 ( .IN1(n9549), .IN2(n9538), .Q(n11384) );
  INVX0 U11233 ( .INP(n11385), .ZN(n11378) );
  AND2X1 U11234 ( .IN1(n11386), .IN2(n11387), .Q(n11385) );
  AND2X1 U11235 ( .IN1(n9554), .IN2(n9540), .Q(n11387) );
  AND2X1 U11236 ( .IN1(n9531), .IN2(n9539), .Q(n11386) );
  XNOR2X1 U11237 ( .IN1(n11154), .IN2(n9538), .Q(n11355) );
  OR2X1 U11238 ( .IN1(n11172), .IN2(n11388), .Q(n11154) );
  OR2X1 U11239 ( .IN1(n11389), .IN2(n11390), .Q(n11388) );
  AND2X1 U11240 ( .IN1(n10252), .IN2(n11168), .Q(n11390) );
  INVX0 U11241 ( .INP(n9532), .ZN(n11168) );
  AND2X1 U11242 ( .IN1(n11391), .IN2(n9532), .Q(n11389) );
  INVX0 U11243 ( .INP(n9549), .ZN(n11391) );
  OR2X1 U11244 ( .IN1(n11392), .IN2(n11063), .Q(n11172) );
  OR2X1 U11245 ( .IN1(n11393), .IN2(n11394), .Q(n11063) );
  OR2X1 U11246 ( .IN1(n11395), .IN2(n10789), .Q(n11394) );
  OR2X1 U11247 ( .IN1(n11396), .IN2(n10815), .Q(n10789) );
  OR2X1 U11248 ( .IN1(n11135), .IN2(n11397), .Q(n10815) );
  XNOR2X1 U11249 ( .IN1(n10252), .IN2(n4513), .Q(n11397) );
  INVX0 U11250 ( .INP(n9547), .ZN(n4513) );
  OR2X1 U11251 ( .IN1(n11398), .IN2(n11399), .Q(n9547) );
  OR2X1 U11252 ( .IN1(n11400), .IN2(n11401), .Q(n11399) );
  AND2X1 U11253 ( .IN1(g165), .IN2(g192), .Q(n11401) );
  AND2X1 U11254 ( .IN1(g6231), .IN2(g186), .Q(n11400) );
  AND2X1 U11255 ( .IN1(test_so13), .IN2(g6313), .Q(n11398) );
  AND2X1 U11256 ( .IN1(n9556), .IN2(n10829), .Q(n11135) );
  XNOR2X1 U11257 ( .IN1(n10829), .IN2(n9531), .Q(n11396) );
  INVX0 U11258 ( .INP(n11402), .ZN(n11395) );
  OR2X1 U11259 ( .IN1(n10829), .IN2(n9554), .Q(n11402) );
  OR2X1 U11260 ( .IN1(n11403), .IN2(n11404), .Q(n11393) );
  AND2X1 U11261 ( .IN1(n10642), .IN2(n9554), .Q(n11404) );
  INVX0 U11262 ( .INP(n9548), .ZN(n10642) );
  AND2X1 U11263 ( .IN1(n10829), .IN2(n9548), .Q(n11403) );
  AND2X1 U11264 ( .IN1(n10829), .IN2(n9549), .Q(n11392) );
  AND2X1 U11265 ( .IN1(n4318), .IN2(g213), .Q(n11347) );
  OR2X1 U11266 ( .IN1(n11405), .IN2(n11406), .Q(g30072) );
  AND2X1 U11267 ( .IN1(n4543), .IN2(n11407), .Q(n11406) );
  OR2X1 U11268 ( .IN1(n11408), .IN2(n11409), .Q(n11407) );
  AND2X1 U11269 ( .IN1(n11410), .IN2(n7929), .Q(n11409) );
  INVX0 U11270 ( .INP(g7302), .ZN(n11410) );
  AND2X1 U11271 ( .IN1(n490), .IN2(n11411), .Q(n11408) );
  AND2X1 U11272 ( .IN1(g2574), .IN2(n7930), .Q(n11405) );
  OR2X1 U11273 ( .IN1(n11412), .IN2(n11413), .Q(g30061) );
  AND2X1 U11274 ( .IN1(n8602), .IN2(n11414), .Q(n11413) );
  OR2X1 U11275 ( .IN1(n11415), .IN2(n11416), .Q(n11414) );
  AND2X1 U11276 ( .IN1(n515), .IN2(g7390), .Q(n11416) );
  INVX0 U11277 ( .INP(n11417), .ZN(n515) );
  OR2X1 U11278 ( .IN1(n11418), .IN2(n11419), .Q(n11417) );
  AND2X1 U11279 ( .IN1(n4493), .IN2(n11420), .Q(n11419) );
  OR2X1 U11280 ( .IN1(n11421), .IN2(n11422), .Q(n11420) );
  AND2X1 U11281 ( .IN1(n9514), .IN2(g7194), .Q(n11422) );
  OR2X1 U11282 ( .IN1(n11423), .IN2(n11424), .Q(n9514) );
  AND2X1 U11283 ( .IN1(n4454), .IN2(n11425), .Q(n11424) );
  OR2X1 U11284 ( .IN1(n11426), .IN2(n11427), .Q(n11425) );
  INVX0 U11285 ( .INP(n11428), .ZN(n11427) );
  OR2X1 U11286 ( .IN1(n517), .IN2(n4316), .Q(n11428) );
  OR2X1 U11287 ( .IN1(n11429), .IN2(n11430), .Q(n517) );
  AND2X1 U11288 ( .IN1(n4570), .IN2(n11431), .Q(n11430) );
  OR2X1 U11289 ( .IN1(g6642), .IN2(g16297), .Q(n11431) );
  AND2X1 U11290 ( .IN1(g506), .IN2(n4571), .Q(n11429) );
  AND2X1 U11291 ( .IN1(n4316), .IN2(DFF_792_n1), .Q(n11426) );
  AND2X1 U11292 ( .IN1(g1192), .IN2(DFF_783_n1), .Q(n11423) );
  AND2X1 U11293 ( .IN1(n4315), .IN2(DFF_1142_n1), .Q(n11421) );
  AND2X1 U11294 ( .IN1(g1886), .IN2(DFF_1133_n1), .Q(n11418) );
  AND2X1 U11295 ( .IN1(n4370), .IN2(g16437), .Q(n11415) );
  AND2X1 U11296 ( .IN1(g2580), .IN2(n7926), .Q(n11412) );
  OR2X1 U11297 ( .IN1(n11432), .IN2(n11433), .Q(g30055) );
  AND2X1 U11298 ( .IN1(n11434), .IN2(g2374), .Q(n11433) );
  OR2X1 U11299 ( .IN1(n11435), .IN2(n11436), .Q(n11434) );
  AND2X1 U11300 ( .IN1(n4524), .IN2(g2380), .Q(n11436) );
  AND2X1 U11301 ( .IN1(g7264), .IN2(n465), .Q(n11435) );
  OR2X1 U11302 ( .IN1(n11437), .IN2(n11438), .Q(n465) );
  AND2X1 U11303 ( .IN1(n11439), .IN2(g1680), .Q(n11438) );
  OR2X1 U11304 ( .IN1(n11440), .IN2(n11441), .Q(n11439) );
  AND2X1 U11305 ( .IN1(n4525), .IN2(g1686), .Q(n11441) );
  AND2X1 U11306 ( .IN1(g7014), .IN2(n467), .Q(n11440) );
  INVX0 U11307 ( .INP(n11442), .ZN(n467) );
  OR2X1 U11308 ( .IN1(n11443), .IN2(n11444), .Q(n11442) );
  AND2X1 U11309 ( .IN1(n11445), .IN2(g986), .Q(n11444) );
  OR2X1 U11310 ( .IN1(n11446), .IN2(n11447), .Q(n11445) );
  AND2X1 U11311 ( .IN1(n11448), .IN2(g6712), .Q(n11447) );
  INVX0 U11312 ( .INP(g21346), .ZN(n11448) );
  AND2X1 U11313 ( .IN1(n4364), .IN2(n8824), .Q(n11446) );
  AND2X1 U11314 ( .IN1(n4432), .IN2(n8017), .Q(n11443) );
  AND2X1 U11315 ( .IN1(n16491), .IN2(n4488), .Q(n11437) );
  AND2X1 U11316 ( .IN1(n4487), .IN2(DFF_1378_n1), .Q(n11432) );
  OR2X1 U11317 ( .IN1(n11449), .IN2(n11450), .Q(g29941) );
  AND2X1 U11318 ( .IN1(n490), .IN2(g3109), .Q(n11450) );
  AND2X1 U11319 ( .IN1(n4494), .IN2(g3105), .Q(n11449) );
  OR2X1 U11320 ( .IN1(n11451), .IN2(n11452), .Q(g29939) );
  AND2X1 U11321 ( .IN1(n490), .IN2(g8030), .Q(n11452) );
  AND2X1 U11322 ( .IN1(n4383), .IN2(g3104), .Q(n11451) );
  OR2X1 U11323 ( .IN1(n11453), .IN2(n11454), .Q(g29936) );
  AND2X1 U11324 ( .IN1(n490), .IN2(g8106), .Q(n11454) );
  INVX0 U11325 ( .INP(n11455), .ZN(n490) );
  OR2X1 U11326 ( .IN1(n11456), .IN2(n11457), .Q(n11455) );
  AND2X1 U11327 ( .IN1(n11458), .IN2(n4545), .Q(n11457) );
  AND2X1 U11328 ( .IN1(n11459), .IN2(n11460), .Q(n11458) );
  OR2X1 U11329 ( .IN1(n4296), .IN2(n11461), .Q(n11460) );
  OR2X1 U11330 ( .IN1(g7052), .IN2(DFF_1100_n1), .Q(n11459) );
  AND2X1 U11331 ( .IN1(g1880), .IN2(DFF_1099_n1), .Q(n11456) );
  AND2X1 U11332 ( .IN1(n4382), .IN2(g3103), .Q(n11453) );
  OR2X1 U11333 ( .IN1(n11462), .IN2(n11463), .Q(g29623) );
  INVX0 U11334 ( .INP(n11464), .ZN(n11463) );
  OR2X1 U11335 ( .IN1(n10833), .IN2(n8387), .Q(n11464) );
  AND2X1 U11336 ( .IN1(n11465), .IN2(n4606), .Q(n11462) );
  OR2X1 U11337 ( .IN1(n11466), .IN2(n11467), .Q(g29621) );
  INVX0 U11338 ( .INP(n11468), .ZN(n11467) );
  OR2X1 U11339 ( .IN1(n10398), .IN2(n8376), .Q(n11468) );
  AND2X1 U11340 ( .IN1(n11465), .IN2(g7264), .Q(n11466) );
  OR2X1 U11341 ( .IN1(n11469), .IN2(n11470), .Q(g29620) );
  INVX0 U11342 ( .INP(n11471), .ZN(n11470) );
  OR2X1 U11343 ( .IN1(n10403), .IN2(n8393), .Q(n11471) );
  AND2X1 U11344 ( .IN1(n11472), .IN2(n4618), .Q(n11469) );
  OR2X1 U11345 ( .IN1(n11473), .IN2(n11474), .Q(g29618) );
  INVX0 U11346 ( .INP(n11475), .ZN(n11474) );
  OR2X1 U11347 ( .IN1(n10408), .IN2(n8388), .Q(n11475) );
  AND2X1 U11348 ( .IN1(n11465), .IN2(g5555), .Q(n11473) );
  AND2X1 U11349 ( .IN1(n11476), .IN2(n10834), .Q(n11465) );
  OR2X1 U11350 ( .IN1(n11477), .IN2(n11191), .Q(n10834) );
  INVX0 U11351 ( .INP(n11478), .ZN(n11477) );
  OR2X1 U11352 ( .IN1(n11479), .IN2(n4529), .Q(n11476) );
  INVX0 U11353 ( .INP(n10718), .ZN(n4529) );
  OR2X1 U11354 ( .IN1(n10850), .IN2(n11480), .Q(n10718) );
  OR2X1 U11355 ( .IN1(n10837), .IN2(n10854), .Q(n11480) );
  INVX0 U11356 ( .INP(n10860), .ZN(n10837) );
  AND2X1 U11357 ( .IN1(n11189), .IN2(n11481), .Q(n11479) );
  AND2X1 U11358 ( .IN1(n11188), .IN2(n10854), .Q(n11481) );
  OR2X1 U11359 ( .IN1(n11482), .IN2(n11483), .Q(g29617) );
  INVX0 U11360 ( .INP(n11484), .ZN(n11483) );
  OR2X1 U11361 ( .IN1(n10412), .IN2(n8379), .Q(n11484) );
  AND2X1 U11362 ( .IN1(n11472), .IN2(g7014), .Q(n11482) );
  OR2X1 U11363 ( .IN1(n11485), .IN2(n11486), .Q(g29616) );
  AND2X1 U11364 ( .IN1(n11487), .IN2(g1088), .Q(n11486) );
  INVX0 U11365 ( .INP(n11488), .ZN(n11485) );
  OR2X1 U11366 ( .IN1(g1088), .IN2(n8398), .Q(n11488) );
  OR2X1 U11367 ( .IN1(n11489), .IN2(n11490), .Q(g29613) );
  INVX0 U11368 ( .INP(n11491), .ZN(n11490) );
  OR2X1 U11369 ( .IN1(n10419), .IN2(n8394), .Q(n11491) );
  AND2X1 U11370 ( .IN1(n11472), .IN2(g5511), .Q(n11489) );
  AND2X1 U11371 ( .IN1(n11492), .IN2(n10420), .Q(n11472) );
  OR2X1 U11372 ( .IN1(n11493), .IN2(n11251), .Q(n10420) );
  INVX0 U11373 ( .INP(n11494), .ZN(n11493) );
  OR2X1 U11374 ( .IN1(n11495), .IN2(n4530), .Q(n11492) );
  INVX0 U11375 ( .INP(n10765), .ZN(n4530) );
  OR2X1 U11376 ( .IN1(n10436), .IN2(n11496), .Q(n10765) );
  OR2X1 U11377 ( .IN1(n10423), .IN2(n10440), .Q(n11496) );
  INVX0 U11378 ( .INP(n10446), .ZN(n10423) );
  AND2X1 U11379 ( .IN1(n11249), .IN2(n11497), .Q(n11495) );
  AND2X1 U11380 ( .IN1(n11248), .IN2(n10440), .Q(n11497) );
  OR2X1 U11381 ( .IN1(n11498), .IN2(n11499), .Q(g29612) );
  AND2X1 U11382 ( .IN1(n11487), .IN2(g6712), .Q(n11499) );
  INVX0 U11383 ( .INP(n11500), .ZN(n11498) );
  OR2X1 U11384 ( .IN1(g6712), .IN2(n8382), .Q(n11500) );
  OR2X1 U11385 ( .IN1(n11501), .IN2(n11502), .Q(g29611) );
  INVX0 U11386 ( .INP(n11503), .ZN(n11502) );
  OR2X1 U11387 ( .IN1(n10465), .IN2(n8405), .Q(n11503) );
  AND2X1 U11388 ( .IN1(n11504), .IN2(n4640), .Q(n11501) );
  OR2X1 U11389 ( .IN1(n11505), .IN2(n11506), .Q(g29609) );
  AND2X1 U11390 ( .IN1(n11487), .IN2(g5472), .Q(n11506) );
  AND2X1 U11391 ( .IN1(n11507), .IN2(n10253), .Q(n11487) );
  OR2X1 U11392 ( .IN1(n11508), .IN2(n11311), .Q(n10253) );
  INVX0 U11393 ( .INP(n11509), .ZN(n11508) );
  OR2X1 U11394 ( .IN1(n11510), .IN2(n10627), .Q(n11507) );
  INVX0 U11395 ( .INP(n10743), .ZN(n10627) );
  OR2X1 U11396 ( .IN1(n10239), .IN2(n11511), .Q(n10743) );
  OR2X1 U11397 ( .IN1(n10249), .IN2(n10232), .Q(n11511) );
  INVX0 U11398 ( .INP(n10243), .ZN(n10249) );
  AND2X1 U11399 ( .IN1(n11309), .IN2(n11512), .Q(n11510) );
  AND2X1 U11400 ( .IN1(n11308), .IN2(n10232), .Q(n11512) );
  INVX0 U11401 ( .INP(n11513), .ZN(n11505) );
  OR2X1 U11402 ( .IN1(g5472), .IN2(n8399), .Q(n11513) );
  OR2X1 U11403 ( .IN1(n11514), .IN2(n11515), .Q(g29608) );
  INVX0 U11404 ( .INP(n11516), .ZN(n11515) );
  OR2X1 U11405 ( .IN1(n10899), .IN2(n8406), .Q(n11516) );
  AND2X1 U11406 ( .IN1(n11504), .IN2(g6447), .Q(n11514) );
  OR2X1 U11407 ( .IN1(n11517), .IN2(n11518), .Q(g29606) );
  INVX0 U11408 ( .INP(n11519), .ZN(n11518) );
  OR2X1 U11409 ( .IN1(n10475), .IN2(n8407), .Q(n11519) );
  AND2X1 U11410 ( .IN1(n11504), .IN2(g5437), .Q(n11517) );
  AND2X1 U11411 ( .IN1(n11520), .IN2(n10476), .Q(n11504) );
  OR2X1 U11412 ( .IN1(n11521), .IN2(n11365), .Q(n10476) );
  INVX0 U11413 ( .INP(n11522), .ZN(n11521) );
  OR2X1 U11414 ( .IN1(n11523), .IN2(n10252), .Q(n11520) );
  INVX0 U11415 ( .INP(n10829), .ZN(n10252) );
  OR2X1 U11416 ( .IN1(n10492), .IN2(n11524), .Q(n10829) );
  OR2X1 U11417 ( .IN1(n10479), .IN2(n10496), .Q(n11524) );
  INVX0 U11418 ( .INP(n10502), .ZN(n10479) );
  AND2X1 U11419 ( .IN1(n11363), .IN2(n11525), .Q(n11523) );
  AND2X1 U11420 ( .IN1(n11362), .IN2(n10496), .Q(n11525) );
  AND2X1 U11421 ( .IN1(n11526), .IN2(n11527), .Q(g29582) );
  XOR2X1 U11422 ( .IN1(n8283), .IN2(n2981), .Q(n11526) );
  AND2X1 U11423 ( .IN1(n11528), .IN2(n11529), .Q(g29581) );
  XOR2X1 U11424 ( .IN1(n8284), .IN2(n2984), .Q(n11528) );
  AND2X1 U11425 ( .IN1(n11530), .IN2(n11531), .Q(g29580) );
  XOR2X1 U11426 ( .IN1(n8285), .IN2(n2987), .Q(n11530) );
  AND2X1 U11427 ( .IN1(n11532), .IN2(n11533), .Q(g29579) );
  XOR2X1 U11428 ( .IN1(n8286), .IN2(n2990), .Q(n11532) );
  AND2X1 U11429 ( .IN1(n11534), .IN2(n11527), .Q(g29357) );
  XNOR2X1 U11430 ( .IN1(n11535), .IN2(n8437), .Q(n11534) );
  AND2X1 U11431 ( .IN1(n11536), .IN2(n11529), .Q(g29355) );
  XNOR2X1 U11432 ( .IN1(n11537), .IN2(n8438), .Q(n11536) );
  AND2X1 U11433 ( .IN1(n11538), .IN2(n11531), .Q(g29354) );
  XNOR2X1 U11434 ( .IN1(n8439), .IN2(n11539), .Q(n11538) );
  AND2X1 U11435 ( .IN1(n11540), .IN2(n11533), .Q(g29353) );
  XNOR2X1 U11436 ( .IN1(n11541), .IN2(n8440), .Q(n11540) );
  OR2X1 U11437 ( .IN1(n11542), .IN2(n11543), .Q(g29226) );
  AND2X1 U11438 ( .IN1(n4509), .IN2(g2498), .Q(n11543) );
  AND2X1 U11439 ( .IN1(n11544), .IN2(n4606), .Q(n11542) );
  OR2X1 U11440 ( .IN1(n11545), .IN2(n11546), .Q(g29221) );
  AND2X1 U11441 ( .IN1(n4524), .IN2(g2495), .Q(n11546) );
  AND2X1 U11442 ( .IN1(n11544), .IN2(g7264), .Q(n11545) );
  OR2X1 U11443 ( .IN1(n11547), .IN2(n11548), .Q(g29218) );
  AND2X1 U11444 ( .IN1(n4511), .IN2(g1804), .Q(n11548) );
  AND2X1 U11445 ( .IN1(n4618), .IN2(n11549), .Q(n11547) );
  OR2X1 U11446 ( .IN1(n11550), .IN2(n11551), .Q(g29213) );
  AND2X1 U11447 ( .IN1(n4516), .IN2(g2492), .Q(n11551) );
  AND2X1 U11448 ( .IN1(n11544), .IN2(g5555), .Q(n11550) );
  XNOR2X1 U11449 ( .IN1(n11552), .IN2(n11553), .Q(n11544) );
  AND2X1 U11450 ( .IN1(n11554), .IN2(test_so79), .Q(n11553) );
  AND2X1 U11451 ( .IN1(n11555), .IN2(n11556), .Q(n11554) );
  OR2X1 U11452 ( .IN1(n11552), .IN2(n11557), .Q(n11556) );
  AND2X1 U11453 ( .IN1(n11558), .IN2(n11559), .Q(n11557) );
  AND2X1 U11454 ( .IN1(n11560), .IN2(n11561), .Q(n11558) );
  OR2X1 U11455 ( .IN1(n4285), .IN2(n11562), .Q(n11555) );
  AND2X1 U11456 ( .IN1(n11563), .IN2(n11564), .Q(n11562) );
  OR2X1 U11457 ( .IN1(n11565), .IN2(n11566), .Q(n11564) );
  INVX0 U11458 ( .INP(n10844), .ZN(n11566) );
  AND2X1 U11459 ( .IN1(n11559), .IN2(n11561), .Q(n11565) );
  OR2X1 U11460 ( .IN1(n11567), .IN2(n11568), .Q(g29212) );
  AND2X1 U11461 ( .IN1(n4525), .IN2(g1801), .Q(n11568) );
  AND2X1 U11462 ( .IN1(g7014), .IN2(n11549), .Q(n11567) );
  OR2X1 U11463 ( .IN1(n11569), .IN2(n11570), .Q(g29209) );
  AND2X1 U11464 ( .IN1(n11571), .IN2(g1088), .Q(n11570) );
  AND2X1 U11465 ( .IN1(n4381), .IN2(g1110), .Q(n11569) );
  OR2X1 U11466 ( .IN1(n11572), .IN2(n11573), .Q(g29205) );
  AND2X1 U11467 ( .IN1(n4518), .IN2(g1798), .Q(n11573) );
  AND2X1 U11468 ( .IN1(g5511), .IN2(n11549), .Q(n11572) );
  XNOR2X1 U11469 ( .IN1(n4284), .IN2(n11574), .Q(n11549) );
  AND2X1 U11470 ( .IN1(n11575), .IN2(n11576), .Q(n11574) );
  OR2X1 U11471 ( .IN1(n11577), .IN2(n11578), .Q(n11576) );
  OR2X1 U11472 ( .IN1(n11579), .IN2(n10430), .Q(n11578) );
  OR2X1 U11473 ( .IN1(n4386), .IN2(n4284), .Q(n11577) );
  OR2X1 U11474 ( .IN1(n11580), .IN2(n11581), .Q(n11575) );
  OR2X1 U11475 ( .IN1(n11582), .IN2(n11583), .Q(n11581) );
  XNOR2X1 U11476 ( .IN1(n11584), .IN2(n11579), .Q(n11583) );
  OR2X1 U11477 ( .IN1(n4386), .IN2(n11585), .Q(n11580) );
  OR2X1 U11478 ( .IN1(n11586), .IN2(n11587), .Q(g29204) );
  AND2X1 U11479 ( .IN1(n11571), .IN2(g6712), .Q(n11587) );
  AND2X1 U11480 ( .IN1(n4364), .IN2(g1107), .Q(n11586) );
  OR2X1 U11481 ( .IN1(n11588), .IN2(n11589), .Q(g29201) );
  AND2X1 U11482 ( .IN1(n4506), .IN2(g423), .Q(n11589) );
  AND2X1 U11483 ( .IN1(n4640), .IN2(n11590), .Q(n11588) );
  OR2X1 U11484 ( .IN1(n11591), .IN2(n11592), .Q(g29198) );
  AND2X1 U11485 ( .IN1(n11571), .IN2(g5472), .Q(n11592) );
  XNOR2X1 U11486 ( .IN1(n11593), .IN2(n11594), .Q(n11571) );
  AND2X1 U11487 ( .IN1(n11595), .IN2(g996), .Q(n11594) );
  AND2X1 U11488 ( .IN1(n11596), .IN2(n11597), .Q(n11595) );
  OR2X1 U11489 ( .IN1(n11593), .IN2(n11598), .Q(n11597) );
  AND2X1 U11490 ( .IN1(n11599), .IN2(n11600), .Q(n11598) );
  AND2X1 U11491 ( .IN1(n11601), .IN2(n11602), .Q(n11599) );
  OR2X1 U11492 ( .IN1(n4283), .IN2(n11603), .Q(n11596) );
  AND2X1 U11493 ( .IN1(n11604), .IN2(n11605), .Q(n11603) );
  OR2X1 U11494 ( .IN1(n11606), .IN2(n11607), .Q(n11605) );
  INVX0 U11495 ( .INP(n10245), .ZN(n11607) );
  AND2X1 U11496 ( .IN1(n11600), .IN2(n11602), .Q(n11606) );
  AND2X1 U11497 ( .IN1(n4363), .IN2(g1104), .Q(n11591) );
  OR2X1 U11498 ( .IN1(n11608), .IN2(n11609), .Q(g29197) );
  AND2X1 U11499 ( .IN1(n4499), .IN2(g420), .Q(n11609) );
  AND2X1 U11500 ( .IN1(g6447), .IN2(n11590), .Q(n11608) );
  OR2X1 U11501 ( .IN1(n11610), .IN2(n11611), .Q(g29194) );
  AND2X1 U11502 ( .IN1(n4520), .IN2(g417), .Q(n11611) );
  AND2X1 U11503 ( .IN1(g5437), .IN2(n11590), .Q(n11610) );
  XNOR2X1 U11504 ( .IN1(n4282), .IN2(n11612), .Q(n11590) );
  AND2X1 U11505 ( .IN1(n11613), .IN2(n11614), .Q(n11612) );
  OR2X1 U11506 ( .IN1(n11615), .IN2(n11616), .Q(n11614) );
  OR2X1 U11507 ( .IN1(n11617), .IN2(n10486), .Q(n11616) );
  OR2X1 U11508 ( .IN1(n4388), .IN2(n4282), .Q(n11615) );
  OR2X1 U11509 ( .IN1(n11618), .IN2(n11619), .Q(n11613) );
  OR2X1 U11510 ( .IN1(n11620), .IN2(n11621), .Q(n11619) );
  XNOR2X1 U11511 ( .IN1(n11622), .IN2(n11617), .Q(n11621) );
  OR2X1 U11512 ( .IN1(n4388), .IN2(n11623), .Q(n11618) );
  OR2X1 U11513 ( .IN1(n11624), .IN2(n11625), .Q(g29187) );
  AND2X1 U11514 ( .IN1(n11626), .IN2(n10833), .Q(n11625) );
  AND2X1 U11515 ( .IN1(n11627), .IN2(g2396), .Q(n11624) );
  OR2X1 U11516 ( .IN1(n4509), .IN2(n11628), .Q(n11627) );
  OR2X1 U11517 ( .IN1(n11629), .IN2(n11630), .Q(g29185) );
  AND2X1 U11518 ( .IN1(n11626), .IN2(n10398), .Q(n11630) );
  AND2X1 U11519 ( .IN1(n11631), .IN2(g2398), .Q(n11629) );
  OR2X1 U11520 ( .IN1(n4524), .IN2(n11628), .Q(n11631) );
  OR2X1 U11521 ( .IN1(n11632), .IN2(n11633), .Q(g29184) );
  AND2X1 U11522 ( .IN1(n11634), .IN2(n10403), .Q(n11633) );
  AND2X1 U11523 ( .IN1(n11635), .IN2(g1702), .Q(n11632) );
  OR2X1 U11524 ( .IN1(n4511), .IN2(n11636), .Q(n11635) );
  OR2X1 U11525 ( .IN1(n11637), .IN2(n11638), .Q(g29182) );
  AND2X1 U11526 ( .IN1(n11626), .IN2(n10408), .Q(n11638) );
  AND2X1 U11527 ( .IN1(n11628), .IN2(n11639), .Q(n11626) );
  INVX0 U11528 ( .INP(n11640), .ZN(n11639) );
  OR2X1 U11529 ( .IN1(n11641), .IN2(n11642), .Q(n11640) );
  AND2X1 U11530 ( .IN1(n10935), .IN2(n11189), .Q(n11642) );
  AND2X1 U11531 ( .IN1(n11643), .IN2(g2397), .Q(n11637) );
  OR2X1 U11532 ( .IN1(n4516), .IN2(n11628), .Q(n11643) );
  OR2X1 U11533 ( .IN1(n11191), .IN2(n11644), .Q(n11628) );
  OR2X1 U11534 ( .IN1(n11641), .IN2(n11645), .Q(n11644) );
  AND2X1 U11535 ( .IN1(n11646), .IN2(n11189), .Q(n11645) );
  OR2X1 U11536 ( .IN1(n10935), .IN2(n11647), .Q(n11646) );
  OR2X1 U11537 ( .IN1(n10871), .IN2(n10942), .Q(n11647) );
  OR2X1 U11538 ( .IN1(n10850), .IN2(n11188), .Q(n10942) );
  OR2X1 U11539 ( .IN1(n10869), .IN2(n11648), .Q(n11188) );
  AND2X1 U11540 ( .IN1(n3038), .IN2(n11649), .Q(n11648) );
  OR2X1 U11541 ( .IN1(n10867), .IN2(n10864), .Q(n11649) );
  OR2X1 U11542 ( .IN1(n11650), .IN2(n11651), .Q(n10864) );
  AND2X1 U11543 ( .IN1(n11652), .IN2(n11653), .Q(n11651) );
  AND2X1 U11544 ( .IN1(n11654), .IN2(n11655), .Q(n11652) );
  OR2X1 U11545 ( .IN1(n11656), .IN2(n11657), .Q(n11655) );
  OR2X1 U11546 ( .IN1(n11658), .IN2(n11659), .Q(n11654) );
  AND2X1 U11547 ( .IN1(n11660), .IN2(n11657), .Q(n11650) );
  AND2X1 U11548 ( .IN1(n11661), .IN2(n11662), .Q(n11660) );
  OR2X1 U11549 ( .IN1(n11653), .IN2(n11659), .Q(n11662) );
  AND2X1 U11550 ( .IN1(n11658), .IN2(n11663), .Q(n10867) );
  AND2X1 U11551 ( .IN1(n11664), .IN2(n11665), .Q(n11663) );
  OR2X1 U11552 ( .IN1(n11653), .IN2(n11656), .Q(n11664) );
  INVX0 U11553 ( .INP(n10853), .ZN(n10869) );
  OR2X1 U11554 ( .IN1(n11666), .IN2(n10857), .Q(n10853) );
  AND2X1 U11555 ( .IN1(n11667), .IN2(n11668), .Q(n11666) );
  OR2X1 U11556 ( .IN1(n11669), .IN2(n11670), .Q(n11668) );
  OR2X1 U11557 ( .IN1(n11671), .IN2(n11672), .Q(n11670) );
  AND2X1 U11558 ( .IN1(n11673), .IN2(n11674), .Q(n11672) );
  AND2X1 U11559 ( .IN1(n11675), .IN2(n11676), .Q(n11671) );
  AND2X1 U11560 ( .IN1(n11677), .IN2(n11678), .Q(n11667) );
  OR2X1 U11561 ( .IN1(n11675), .IN2(n11679), .Q(n11678) );
  OR2X1 U11562 ( .IN1(n11680), .IN2(n11681), .Q(n11679) );
  AND2X1 U11563 ( .IN1(n11669), .IN2(n11673), .Q(n11681) );
  OR2X1 U11564 ( .IN1(n11674), .IN2(n11682), .Q(n11677) );
  OR2X1 U11565 ( .IN1(n11683), .IN2(n11684), .Q(n11682) );
  AND2X1 U11566 ( .IN1(n11675), .IN2(n11673), .Q(n11684) );
  AND2X1 U11567 ( .IN1(n11669), .IN2(n11676), .Q(n11683) );
  OR2X1 U11568 ( .IN1(n10870), .IN2(n10857), .Q(n10935) );
  AND2X1 U11569 ( .IN1(n11685), .IN2(n11686), .Q(n10870) );
  INVX0 U11570 ( .INP(n11687), .ZN(n11686) );
  OR2X1 U11571 ( .IN1(n11688), .IN2(n11665), .Q(n11687) );
  OR2X1 U11572 ( .IN1(n11657), .IN2(n11659), .Q(n11665) );
  XNOR2X1 U11573 ( .IN1(n4563), .IN2(n9653), .Q(n11659) );
  OR2X1 U11574 ( .IN1(n11689), .IN2(n11690), .Q(n9653) );
  OR2X1 U11575 ( .IN1(n11691), .IN2(n11692), .Q(n11690) );
  AND2X1 U11576 ( .IN1(g2241), .IN2(g2294), .Q(n11692) );
  AND2X1 U11577 ( .IN1(g6837), .IN2(g2288), .Q(n11691) );
  AND2X1 U11578 ( .IN1(test_so73), .IN2(g2291), .Q(n11689) );
  XNOR2X1 U11579 ( .IN1(n11693), .IN2(n9643), .Q(n11657) );
  OR2X1 U11580 ( .IN1(n11694), .IN2(n11695), .Q(n9643) );
  OR2X1 U11581 ( .IN1(n11696), .IN2(n11697), .Q(n11695) );
  AND2X1 U11582 ( .IN1(g2241), .IN2(g2303), .Q(n11697) );
  AND2X1 U11583 ( .IN1(g6837), .IN2(g2297), .Q(n11696) );
  AND2X1 U11584 ( .IN1(test_so73), .IN2(g2300), .Q(n11694) );
  OR2X1 U11585 ( .IN1(n11653), .IN2(n11661), .Q(n11688) );
  OR2X1 U11586 ( .IN1(n11658), .IN2(n11656), .Q(n11661) );
  XNOR2X1 U11587 ( .IN1(n4319), .IN2(n9654), .Q(n11656) );
  OR2X1 U11588 ( .IN1(n11698), .IN2(n11699), .Q(n9654) );
  OR2X1 U11589 ( .IN1(n11700), .IN2(n11701), .Q(n11699) );
  AND2X1 U11590 ( .IN1(g2241), .IN2(g2276), .Q(n11701) );
  AND2X1 U11591 ( .IN1(g6837), .IN2(g2270), .Q(n11700) );
  AND2X1 U11592 ( .IN1(test_so73), .IN2(g2273), .Q(n11698) );
  XNOR2X1 U11593 ( .IN1(n4377), .IN2(n9645), .Q(n11658) );
  OR2X1 U11594 ( .IN1(n11702), .IN2(n11703), .Q(n9645) );
  OR2X1 U11595 ( .IN1(n11704), .IN2(n11705), .Q(n11703) );
  AND2X1 U11596 ( .IN1(g2241), .IN2(g2267), .Q(n11705) );
  AND2X1 U11597 ( .IN1(g6837), .IN2(g2261), .Q(n11704) );
  AND2X1 U11598 ( .IN1(test_so76), .IN2(test_so73), .Q(n11702) );
  XNOR2X1 U11599 ( .IN1(n4325), .IN2(n9652), .Q(n11653) );
  OR2X1 U11600 ( .IN1(n11706), .IN2(n11707), .Q(n9652) );
  OR2X1 U11601 ( .IN1(n11708), .IN2(n11709), .Q(n11707) );
  AND2X1 U11602 ( .IN1(g2241), .IN2(g2285), .Q(n11709) );
  AND2X1 U11603 ( .IN1(g6837), .IN2(g2279), .Q(n11708) );
  AND2X1 U11604 ( .IN1(test_so73), .IN2(g2282), .Q(n11706) );
  AND2X1 U11605 ( .IN1(n11710), .IN2(n11711), .Q(n11685) );
  AND2X1 U11606 ( .IN1(n11669), .IN2(n11675), .Q(n11711) );
  XOR2X1 U11607 ( .IN1(n10555), .IN2(n9636), .Q(n11675) );
  OR2X1 U11608 ( .IN1(n11712), .IN2(n11713), .Q(n9636) );
  OR2X1 U11609 ( .IN1(n11714), .IN2(n11715), .Q(n11713) );
  AND2X1 U11610 ( .IN1(g2241), .IN2(g2348), .Q(n11715) );
  AND2X1 U11611 ( .IN1(g6837), .IN2(g2342), .Q(n11714) );
  AND2X1 U11612 ( .IN1(test_so73), .IN2(g2345), .Q(n11712) );
  XNOR2X1 U11613 ( .IN1(g2190), .IN2(n9637), .Q(n11669) );
  OR2X1 U11614 ( .IN1(n11716), .IN2(n11717), .Q(n9637) );
  OR2X1 U11615 ( .IN1(n11718), .IN2(n11719), .Q(n11717) );
  AND2X1 U11616 ( .IN1(g2241), .IN2(g2330), .Q(n11719) );
  AND2X1 U11617 ( .IN1(g6837), .IN2(g2324), .Q(n11718) );
  AND2X1 U11618 ( .IN1(test_so77), .IN2(test_so73), .Q(n11716) );
  AND2X1 U11619 ( .IN1(n11673), .IN2(n11680), .Q(n11710) );
  AND2X1 U11620 ( .IN1(n11674), .IN2(n11676), .Q(n11680) );
  XNOR2X1 U11621 ( .IN1(n4389), .IN2(n11225), .Q(n11676) );
  INVX0 U11622 ( .INP(n9644), .ZN(n11225) );
  OR2X1 U11623 ( .IN1(n11720), .IN2(n11721), .Q(n9644) );
  OR2X1 U11624 ( .IN1(n11722), .IN2(n11723), .Q(n11721) );
  AND2X1 U11625 ( .IN1(g2241), .IN2(g2321), .Q(n11723) );
  AND2X1 U11626 ( .IN1(g6837), .IN2(g2315), .Q(n11722) );
  AND2X1 U11627 ( .IN1(test_so73), .IN2(g2318), .Q(n11720) );
  XNOR2X1 U11628 ( .IN1(n4373), .IN2(n9658), .Q(n11674) );
  INVX0 U11629 ( .INP(n11204), .ZN(n9658) );
  OR2X1 U11630 ( .IN1(n11724), .IN2(n11725), .Q(n11204) );
  OR2X1 U11631 ( .IN1(n11726), .IN2(n11727), .Q(n11725) );
  AND2X1 U11632 ( .IN1(g2241), .IN2(g2312), .Q(n11727) );
  AND2X1 U11633 ( .IN1(g6837), .IN2(g2306), .Q(n11726) );
  AND2X1 U11634 ( .IN1(test_so73), .IN2(g2309), .Q(n11724) );
  XNOR2X1 U11635 ( .IN1(g2200), .IN2(n9638), .Q(n11673) );
  OR2X1 U11636 ( .IN1(n11728), .IN2(n11729), .Q(n9638) );
  OR2X1 U11637 ( .IN1(n11730), .IN2(n11731), .Q(n11729) );
  AND2X1 U11638 ( .IN1(g2241), .IN2(g2339), .Q(n11731) );
  AND2X1 U11639 ( .IN1(g6837), .IN2(g2333), .Q(n11730) );
  AND2X1 U11640 ( .IN1(test_so73), .IN2(g2336), .Q(n11728) );
  AND2X1 U11641 ( .IN1(n11732), .IN2(n9121), .Q(n11641) );
  OR2X1 U11642 ( .IN1(n11733), .IN2(n11734), .Q(g29181) );
  AND2X1 U11643 ( .IN1(n11634), .IN2(n10412), .Q(n11734) );
  AND2X1 U11644 ( .IN1(n11735), .IN2(g1704), .Q(n11733) );
  OR2X1 U11645 ( .IN1(n4525), .IN2(n11636), .Q(n11735) );
  OR2X1 U11646 ( .IN1(n11736), .IN2(n11737), .Q(g29179) );
  AND2X1 U11647 ( .IN1(n11738), .IN2(g1088), .Q(n11737) );
  AND2X1 U11648 ( .IN1(n11739), .IN2(g1008), .Q(n11736) );
  OR2X1 U11649 ( .IN1(n4381), .IN2(n11740), .Q(n11739) );
  OR2X1 U11650 ( .IN1(n11741), .IN2(n11742), .Q(g29178) );
  AND2X1 U11651 ( .IN1(n11634), .IN2(n10419), .Q(n11742) );
  AND2X1 U11652 ( .IN1(n11636), .IN2(n11743), .Q(n11634) );
  INVX0 U11653 ( .INP(n11744), .ZN(n11743) );
  OR2X1 U11654 ( .IN1(n11745), .IN2(n11746), .Q(n11744) );
  AND2X1 U11655 ( .IN1(n10955), .IN2(n11249), .Q(n11746) );
  AND2X1 U11656 ( .IN1(n11747), .IN2(g1703), .Q(n11741) );
  OR2X1 U11657 ( .IN1(n4518), .IN2(n11636), .Q(n11747) );
  OR2X1 U11658 ( .IN1(n11251), .IN2(n11748), .Q(n11636) );
  OR2X1 U11659 ( .IN1(n11745), .IN2(n11749), .Q(n11748) );
  AND2X1 U11660 ( .IN1(n11750), .IN2(n11249), .Q(n11749) );
  OR2X1 U11661 ( .IN1(n10955), .IN2(n11751), .Q(n11750) );
  OR2X1 U11662 ( .IN1(n10457), .IN2(n10962), .Q(n11751) );
  OR2X1 U11663 ( .IN1(n10436), .IN2(n11248), .Q(n10962) );
  OR2X1 U11664 ( .IN1(n10455), .IN2(n11752), .Q(n11248) );
  AND2X1 U11665 ( .IN1(n3070), .IN2(n11753), .Q(n11752) );
  OR2X1 U11666 ( .IN1(n10453), .IN2(n10450), .Q(n11753) );
  OR2X1 U11667 ( .IN1(n11754), .IN2(n11755), .Q(n10450) );
  AND2X1 U11668 ( .IN1(n11756), .IN2(n11757), .Q(n11755) );
  AND2X1 U11669 ( .IN1(n11758), .IN2(n11759), .Q(n11756) );
  OR2X1 U11670 ( .IN1(n11760), .IN2(n11761), .Q(n11759) );
  OR2X1 U11671 ( .IN1(n11762), .IN2(n11763), .Q(n11758) );
  AND2X1 U11672 ( .IN1(n11764), .IN2(n11761), .Q(n11754) );
  AND2X1 U11673 ( .IN1(n11765), .IN2(n11766), .Q(n11764) );
  OR2X1 U11674 ( .IN1(n11757), .IN2(n11763), .Q(n11766) );
  AND2X1 U11675 ( .IN1(n11762), .IN2(n11767), .Q(n10453) );
  AND2X1 U11676 ( .IN1(n11768), .IN2(n11769), .Q(n11767) );
  OR2X1 U11677 ( .IN1(n11757), .IN2(n11760), .Q(n11768) );
  INVX0 U11678 ( .INP(n10439), .ZN(n10455) );
  OR2X1 U11679 ( .IN1(n11770), .IN2(n10443), .Q(n10439) );
  AND2X1 U11680 ( .IN1(n11771), .IN2(n11772), .Q(n11770) );
  OR2X1 U11681 ( .IN1(n11773), .IN2(n11774), .Q(n11772) );
  OR2X1 U11682 ( .IN1(n11775), .IN2(n11776), .Q(n11774) );
  AND2X1 U11683 ( .IN1(n11777), .IN2(n11778), .Q(n11776) );
  AND2X1 U11684 ( .IN1(n11779), .IN2(n11780), .Q(n11775) );
  AND2X1 U11685 ( .IN1(n11781), .IN2(n11782), .Q(n11771) );
  OR2X1 U11686 ( .IN1(n11779), .IN2(n11783), .Q(n11782) );
  OR2X1 U11687 ( .IN1(n11784), .IN2(n11785), .Q(n11783) );
  AND2X1 U11688 ( .IN1(n11773), .IN2(n11777), .Q(n11785) );
  AND2X1 U11689 ( .IN1(n11780), .IN2(n11778), .Q(n11784) );
  OR2X1 U11690 ( .IN1(n11778), .IN2(n11786), .Q(n11781) );
  OR2X1 U11691 ( .IN1(n11787), .IN2(n11788), .Q(n11786) );
  AND2X1 U11692 ( .IN1(n11779), .IN2(n11777), .Q(n11788) );
  INVX0 U11693 ( .INP(n11789), .ZN(n11779) );
  AND2X1 U11694 ( .IN1(n11773), .IN2(n11780), .Q(n11787) );
  INVX0 U11695 ( .INP(n11790), .ZN(n11780) );
  INVX0 U11696 ( .INP(n11791), .ZN(n11773) );
  INVX0 U11697 ( .INP(n11792), .ZN(n11778) );
  OR2X1 U11698 ( .IN1(n10456), .IN2(n10443), .Q(n10955) );
  INVX0 U11699 ( .INP(n10444), .ZN(n10456) );
  OR2X1 U11700 ( .IN1(n11793), .IN2(n11794), .Q(n10444) );
  OR2X1 U11701 ( .IN1(n11795), .IN2(n11769), .Q(n11794) );
  OR2X1 U11702 ( .IN1(n11761), .IN2(n11763), .Q(n11769) );
  XNOR2X1 U11703 ( .IN1(n4565), .IN2(n9619), .Q(n11763) );
  OR2X1 U11704 ( .IN1(n11796), .IN2(n11797), .Q(n9619) );
  OR2X1 U11705 ( .IN1(n11798), .IN2(n11799), .Q(n11797) );
  AND2X1 U11706 ( .IN1(g1547), .IN2(g1600), .Q(n11799) );
  AND2X1 U11707 ( .IN1(g6573), .IN2(g1594), .Q(n11798) );
  AND2X1 U11708 ( .IN1(g6782), .IN2(g1597), .Q(n11796) );
  XNOR2X1 U11709 ( .IN1(n11800), .IN2(n9618), .Q(n11761) );
  OR2X1 U11710 ( .IN1(n11801), .IN2(n11802), .Q(n9618) );
  OR2X1 U11711 ( .IN1(n11803), .IN2(n11804), .Q(n11802) );
  AND2X1 U11712 ( .IN1(g1547), .IN2(g1609), .Q(n11804) );
  AND2X1 U11713 ( .IN1(g6573), .IN2(g1603), .Q(n11803) );
  AND2X1 U11714 ( .IN1(test_so56), .IN2(g6782), .Q(n11801) );
  OR2X1 U11715 ( .IN1(n11757), .IN2(n11765), .Q(n11795) );
  OR2X1 U11716 ( .IN1(n11762), .IN2(n11760), .Q(n11765) );
  XNOR2X1 U11717 ( .IN1(n4320), .IN2(n9617), .Q(n11760) );
  OR2X1 U11718 ( .IN1(n11805), .IN2(n11806), .Q(n9617) );
  OR2X1 U11719 ( .IN1(n11807), .IN2(n11808), .Q(n11806) );
  AND2X1 U11720 ( .IN1(g1547), .IN2(g1582), .Q(n11808) );
  AND2X1 U11721 ( .IN1(g6573), .IN2(g1576), .Q(n11807) );
  AND2X1 U11722 ( .IN1(g6782), .IN2(g1579), .Q(n11805) );
  XNOR2X1 U11723 ( .IN1(n4378), .IN2(n9608), .Q(n11762) );
  OR2X1 U11724 ( .IN1(n11809), .IN2(n11810), .Q(n9608) );
  OR2X1 U11725 ( .IN1(n11811), .IN2(n11812), .Q(n11810) );
  AND2X1 U11726 ( .IN1(g1547), .IN2(g1573), .Q(n11812) );
  AND2X1 U11727 ( .IN1(g6573), .IN2(g1567), .Q(n11811) );
  AND2X1 U11728 ( .IN1(g6782), .IN2(g1570), .Q(n11809) );
  XNOR2X1 U11729 ( .IN1(n4326), .IN2(n9623), .Q(n11757) );
  OR2X1 U11730 ( .IN1(n11813), .IN2(n11814), .Q(n9623) );
  OR2X1 U11731 ( .IN1(n11815), .IN2(n11816), .Q(n11814) );
  AND2X1 U11732 ( .IN1(g1547), .IN2(g1591), .Q(n11816) );
  AND2X1 U11733 ( .IN1(g6573), .IN2(g1585), .Q(n11815) );
  AND2X1 U11734 ( .IN1(g6782), .IN2(g1588), .Q(n11813) );
  OR2X1 U11735 ( .IN1(n11817), .IN2(n11818), .Q(n11793) );
  OR2X1 U11736 ( .IN1(n11791), .IN2(n11789), .Q(n11818) );
  XNOR2X1 U11737 ( .IN1(n10588), .IN2(n11819), .Q(n11789) );
  INVX0 U11738 ( .INP(n9609), .ZN(n10588) );
  OR2X1 U11739 ( .IN1(n11820), .IN2(n11821), .Q(n9609) );
  OR2X1 U11740 ( .IN1(n11822), .IN2(n11823), .Q(n11821) );
  AND2X1 U11741 ( .IN1(g1547), .IN2(g1654), .Q(n11823) );
  AND2X1 U11742 ( .IN1(g6573), .IN2(g1648), .Q(n11822) );
  AND2X1 U11743 ( .IN1(g6782), .IN2(g1651), .Q(n11820) );
  XNOR2X1 U11744 ( .IN1(n4557), .IN2(n9602), .Q(n11791) );
  OR2X1 U11745 ( .IN1(n11824), .IN2(n11825), .Q(n9602) );
  OR2X1 U11746 ( .IN1(n11826), .IN2(n11827), .Q(n11825) );
  AND2X1 U11747 ( .IN1(g1547), .IN2(g1636), .Q(n11827) );
  AND2X1 U11748 ( .IN1(g6573), .IN2(g1630), .Q(n11826) );
  AND2X1 U11749 ( .IN1(g6782), .IN2(g1633), .Q(n11824) );
  OR2X1 U11750 ( .IN1(n11828), .IN2(n11829), .Q(n11817) );
  OR2X1 U11751 ( .IN1(n11792), .IN2(n11790), .Q(n11829) );
  XNOR2X1 U11752 ( .IN1(n4390), .IN2(n9610), .Q(n11790) );
  OR2X1 U11753 ( .IN1(n11830), .IN2(n11831), .Q(n9610) );
  OR2X1 U11754 ( .IN1(n11832), .IN2(n11833), .Q(n11831) );
  AND2X1 U11755 ( .IN1(g1547), .IN2(g1627), .Q(n11833) );
  AND2X1 U11756 ( .IN1(test_so55), .IN2(g6573), .Q(n11832) );
  AND2X1 U11757 ( .IN1(g6782), .IN2(g1624), .Q(n11830) );
  XNOR2X1 U11758 ( .IN1(n4374), .IN2(n9601), .Q(n11792) );
  OR2X1 U11759 ( .IN1(n11834), .IN2(n11835), .Q(n9601) );
  OR2X1 U11760 ( .IN1(n11836), .IN2(n11837), .Q(n11835) );
  AND2X1 U11761 ( .IN1(g1547), .IN2(g1618), .Q(n11837) );
  AND2X1 U11762 ( .IN1(g6573), .IN2(g1612), .Q(n11836) );
  AND2X1 U11763 ( .IN1(g6782), .IN2(g1615), .Q(n11834) );
  INVX0 U11764 ( .INP(n11777), .ZN(n11828) );
  XOR2X1 U11765 ( .IN1(n4288), .IN2(n9603), .Q(n11777) );
  OR2X1 U11766 ( .IN1(n11838), .IN2(n11839), .Q(n9603) );
  OR2X1 U11767 ( .IN1(n11840), .IN2(n11841), .Q(n11839) );
  AND2X1 U11768 ( .IN1(g1547), .IN2(g1645), .Q(n11841) );
  AND2X1 U11769 ( .IN1(g6573), .IN2(g1639), .Q(n11840) );
  AND2X1 U11770 ( .IN1(g6782), .IN2(g1642), .Q(n11838) );
  AND2X1 U11771 ( .IN1(n4386), .IN2(n11842), .Q(n11745) );
  OR2X1 U11772 ( .IN1(n11843), .IN2(n11844), .Q(g29173) );
  AND2X1 U11773 ( .IN1(n11738), .IN2(g6712), .Q(n11844) );
  AND2X1 U11774 ( .IN1(n11845), .IN2(g1010), .Q(n11843) );
  OR2X1 U11775 ( .IN1(n4364), .IN2(n11740), .Q(n11845) );
  OR2X1 U11776 ( .IN1(n11846), .IN2(n11847), .Q(g29172) );
  AND2X1 U11777 ( .IN1(n11848), .IN2(n10465), .Q(n11847) );
  AND2X1 U11778 ( .IN1(n11849), .IN2(g321), .Q(n11846) );
  OR2X1 U11779 ( .IN1(n4506), .IN2(n11850), .Q(n11849) );
  OR2X1 U11780 ( .IN1(n11851), .IN2(n11852), .Q(g29170) );
  AND2X1 U11781 ( .IN1(n11738), .IN2(g5472), .Q(n11852) );
  AND2X1 U11782 ( .IN1(n11740), .IN2(n11853), .Q(n11738) );
  INVX0 U11783 ( .INP(n11854), .ZN(n11853) );
  OR2X1 U11784 ( .IN1(n11855), .IN2(n11856), .Q(n11854) );
  AND2X1 U11785 ( .IN1(n11309), .IN2(n10238), .Q(n11856) );
  AND2X1 U11786 ( .IN1(n11857), .IN2(g1009), .Q(n11851) );
  OR2X1 U11787 ( .IN1(n4363), .IN2(n11740), .Q(n11857) );
  OR2X1 U11788 ( .IN1(n11311), .IN2(n11858), .Q(n11740) );
  OR2X1 U11789 ( .IN1(n11855), .IN2(n11859), .Q(n11858) );
  AND2X1 U11790 ( .IN1(n11860), .IN2(n11309), .Q(n11859) );
  OR2X1 U11791 ( .IN1(n10238), .IN2(n11861), .Q(n11860) );
  OR2X1 U11792 ( .IN1(n10236), .IN2(n10251), .Q(n11861) );
  OR2X1 U11793 ( .IN1(n10239), .IN2(n11308), .Q(n10251) );
  OR2X1 U11794 ( .IN1(n10280), .IN2(n11862), .Q(n11308) );
  AND2X1 U11795 ( .IN1(n3102), .IN2(n11863), .Q(n11862) );
  OR2X1 U11796 ( .IN1(n10278), .IN2(n10275), .Q(n11863) );
  OR2X1 U11797 ( .IN1(n11864), .IN2(n11865), .Q(n10275) );
  AND2X1 U11798 ( .IN1(n11866), .IN2(n11867), .Q(n11865) );
  AND2X1 U11799 ( .IN1(n11868), .IN2(n11869), .Q(n11866) );
  OR2X1 U11800 ( .IN1(n11870), .IN2(n11871), .Q(n11869) );
  OR2X1 U11801 ( .IN1(n11872), .IN2(n11873), .Q(n11868) );
  AND2X1 U11802 ( .IN1(n11874), .IN2(n11871), .Q(n11864) );
  AND2X1 U11803 ( .IN1(n11875), .IN2(n11876), .Q(n11874) );
  OR2X1 U11804 ( .IN1(n11867), .IN2(n11873), .Q(n11876) );
  AND2X1 U11805 ( .IN1(n11872), .IN2(n11877), .Q(n10278) );
  AND2X1 U11806 ( .IN1(n11878), .IN2(n11879), .Q(n11877) );
  OR2X1 U11807 ( .IN1(n11867), .IN2(n11870), .Q(n11878) );
  INVX0 U11808 ( .INP(n10267), .ZN(n10280) );
  OR2X1 U11809 ( .IN1(n11880), .IN2(n10247), .Q(n10267) );
  AND2X1 U11810 ( .IN1(n11881), .IN2(n11882), .Q(n11880) );
  OR2X1 U11811 ( .IN1(n11883), .IN2(n11884), .Q(n11882) );
  OR2X1 U11812 ( .IN1(n11885), .IN2(n11886), .Q(n11884) );
  AND2X1 U11813 ( .IN1(n11887), .IN2(n11888), .Q(n11885) );
  AND2X1 U11814 ( .IN1(n11889), .IN2(n11890), .Q(n11881) );
  OR2X1 U11815 ( .IN1(n11888), .IN2(n11891), .Q(n11890) );
  OR2X1 U11816 ( .IN1(n11892), .IN2(n11893), .Q(n11891) );
  AND2X1 U11817 ( .IN1(n11883), .IN2(n11894), .Q(n11893) );
  AND2X1 U11818 ( .IN1(n11887), .IN2(n11895), .Q(n11892) );
  OR2X1 U11819 ( .IN1(n11895), .IN2(n11896), .Q(n11889) );
  OR2X1 U11820 ( .IN1(n11897), .IN2(n11898), .Q(n11896) );
  AND2X1 U11821 ( .IN1(n11888), .IN2(n11894), .Q(n11897) );
  OR2X1 U11822 ( .IN1(n10270), .IN2(n10247), .Q(n10238) );
  AND2X1 U11823 ( .IN1(n11899), .IN2(n11900), .Q(n10270) );
  AND2X1 U11824 ( .IN1(n11901), .IN2(n11898), .Q(n11900) );
  AND2X1 U11825 ( .IN1(n11887), .IN2(n11883), .Q(n11898) );
  XNOR2X1 U11826 ( .IN1(g805), .IN2(n9568), .Q(n11883) );
  OR2X1 U11827 ( .IN1(n11902), .IN2(n11903), .Q(n9568) );
  OR2X1 U11828 ( .IN1(n11904), .IN2(n11905), .Q(n11903) );
  AND2X1 U11829 ( .IN1(g6368), .IN2(g936), .Q(n11905) );
  AND2X1 U11830 ( .IN1(g6518), .IN2(g939), .Q(n11904) );
  AND2X1 U11831 ( .IN1(test_so31), .IN2(g942), .Q(n11902) );
  XOR2X1 U11832 ( .IN1(n4391), .IN2(n9567), .Q(n11887) );
  OR2X1 U11833 ( .IN1(n11906), .IN2(n11907), .Q(n9567) );
  OR2X1 U11834 ( .IN1(n11908), .IN2(n11909), .Q(n11907) );
  AND2X1 U11835 ( .IN1(g6368), .IN2(g927), .Q(n11909) );
  AND2X1 U11836 ( .IN1(g6518), .IN2(g930), .Q(n11908) );
  AND2X1 U11837 ( .IN1(test_so31), .IN2(g933), .Q(n11906) );
  AND2X1 U11838 ( .IN1(n11888), .IN2(n11886), .Q(n11901) );
  AND2X1 U11839 ( .IN1(n11894), .IN2(n11895), .Q(n11886) );
  XOR2X1 U11840 ( .IN1(n4375), .IN2(n9569), .Q(n11895) );
  OR2X1 U11841 ( .IN1(n11910), .IN2(n11911), .Q(n9569) );
  OR2X1 U11842 ( .IN1(n11912), .IN2(n11913), .Q(n11911) );
  AND2X1 U11843 ( .IN1(g6368), .IN2(g918), .Q(n11913) );
  AND2X1 U11844 ( .IN1(g6518), .IN2(g921), .Q(n11912) );
  AND2X1 U11845 ( .IN1(test_so34), .IN2(test_so31), .Q(n11910) );
  XNOR2X1 U11846 ( .IN1(g813), .IN2(n9589), .Q(n11894) );
  OR2X1 U11847 ( .IN1(n11914), .IN2(n11915), .Q(n9589) );
  OR2X1 U11848 ( .IN1(n11916), .IN2(n11917), .Q(n11915) );
  AND2X1 U11849 ( .IN1(test_so35), .IN2(g6368), .Q(n11917) );
  AND2X1 U11850 ( .IN1(g6518), .IN2(g948), .Q(n11916) );
  AND2X1 U11851 ( .IN1(test_so31), .IN2(g951), .Q(n11914) );
  XNOR2X1 U11852 ( .IN1(n10629), .IN2(n9575), .Q(n11888) );
  INVX0 U11853 ( .INP(n10623), .ZN(n9575) );
  OR2X1 U11854 ( .IN1(n11918), .IN2(n11919), .Q(n10623) );
  OR2X1 U11855 ( .IN1(n11920), .IN2(n11921), .Q(n11919) );
  AND2X1 U11856 ( .IN1(g6368), .IN2(g954), .Q(n11921) );
  AND2X1 U11857 ( .IN1(g6518), .IN2(g957), .Q(n11920) );
  AND2X1 U11858 ( .IN1(test_so31), .IN2(g960), .Q(n11918) );
  INVX0 U11859 ( .INP(n11922), .ZN(n11899) );
  OR2X1 U11860 ( .IN1(n11923), .IN2(n11879), .Q(n11922) );
  OR2X1 U11861 ( .IN1(n11873), .IN2(n11871), .Q(n11879) );
  XNOR2X1 U11862 ( .IN1(n11924), .IN2(n9584), .Q(n11871) );
  OR2X1 U11863 ( .IN1(n11925), .IN2(n11926), .Q(n9584) );
  OR2X1 U11864 ( .IN1(n11927), .IN2(n11928), .Q(n11926) );
  AND2X1 U11865 ( .IN1(g6368), .IN2(g909), .Q(n11928) );
  AND2X1 U11866 ( .IN1(g6518), .IN2(g912), .Q(n11927) );
  AND2X1 U11867 ( .IN1(test_so31), .IN2(g915), .Q(n11925) );
  XNOR2X1 U11868 ( .IN1(n4567), .IN2(n9574), .Q(n11873) );
  OR2X1 U11869 ( .IN1(n11929), .IN2(n11930), .Q(n9574) );
  OR2X1 U11870 ( .IN1(n11931), .IN2(n11932), .Q(n11930) );
  AND2X1 U11871 ( .IN1(g6368), .IN2(g900), .Q(n11932) );
  AND2X1 U11872 ( .IN1(g6518), .IN2(g903), .Q(n11931) );
  AND2X1 U11873 ( .IN1(test_so31), .IN2(g906), .Q(n11929) );
  OR2X1 U11874 ( .IN1(n11867), .IN2(n11875), .Q(n11923) );
  OR2X1 U11875 ( .IN1(n11870), .IN2(n11872), .Q(n11875) );
  XNOR2X1 U11876 ( .IN1(g785), .IN2(n11344), .Q(n11872) );
  INVX0 U11877 ( .INP(n9576), .ZN(n11344) );
  OR2X1 U11878 ( .IN1(n11933), .IN2(n11934), .Q(n9576) );
  OR2X1 U11879 ( .IN1(n11935), .IN2(n11936), .Q(n11934) );
  AND2X1 U11880 ( .IN1(g6368), .IN2(g873), .Q(n11936) );
  AND2X1 U11881 ( .IN1(g6518), .IN2(g876), .Q(n11935) );
  AND2X1 U11882 ( .IN1(test_so31), .IN2(g879), .Q(n11933) );
  XNOR2X1 U11883 ( .IN1(g793), .IN2(n11326), .Q(n11870) );
  INVX0 U11884 ( .INP(n9585), .ZN(n11326) );
  OR2X1 U11885 ( .IN1(n11937), .IN2(n11938), .Q(n9585) );
  OR2X1 U11886 ( .IN1(n11939), .IN2(n11940), .Q(n11938) );
  AND2X1 U11887 ( .IN1(g6368), .IN2(g882), .Q(n11940) );
  AND2X1 U11888 ( .IN1(g6518), .IN2(g885), .Q(n11939) );
  AND2X1 U11889 ( .IN1(test_so31), .IN2(g888), .Q(n11937) );
  XNOR2X1 U11890 ( .IN1(g801), .IN2(n11147), .Q(n11867) );
  INVX0 U11891 ( .INP(n9583), .ZN(n11147) );
  OR2X1 U11892 ( .IN1(n11941), .IN2(n11942), .Q(n9583) );
  OR2X1 U11893 ( .IN1(n11943), .IN2(n11944), .Q(n11942) );
  AND2X1 U11894 ( .IN1(g6368), .IN2(g891), .Q(n11944) );
  AND2X1 U11895 ( .IN1(g6518), .IN2(g894), .Q(n11943) );
  AND2X1 U11896 ( .IN1(test_so31), .IN2(g897), .Q(n11941) );
  AND2X1 U11897 ( .IN1(n4387), .IN2(n11945), .Q(n11855) );
  OR2X1 U11898 ( .IN1(n11946), .IN2(n11947), .Q(g29169) );
  AND2X1 U11899 ( .IN1(n11848), .IN2(n10899), .Q(n11947) );
  AND2X1 U11900 ( .IN1(n11948), .IN2(g323), .Q(n11946) );
  OR2X1 U11901 ( .IN1(n4499), .IN2(n11850), .Q(n11948) );
  OR2X1 U11902 ( .IN1(n11949), .IN2(n11950), .Q(g29167) );
  AND2X1 U11903 ( .IN1(n11848), .IN2(n10475), .Q(n11950) );
  AND2X1 U11904 ( .IN1(n11850), .IN2(n11951), .Q(n11848) );
  INVX0 U11905 ( .INP(n11952), .ZN(n11951) );
  OR2X1 U11906 ( .IN1(n11953), .IN2(n11954), .Q(n11952) );
  AND2X1 U11907 ( .IN1(n10912), .IN2(n11363), .Q(n11954) );
  AND2X1 U11908 ( .IN1(n11955), .IN2(g322), .Q(n11949) );
  OR2X1 U11909 ( .IN1(n4520), .IN2(n11850), .Q(n11955) );
  OR2X1 U11910 ( .IN1(n11365), .IN2(n11956), .Q(n11850) );
  OR2X1 U11911 ( .IN1(n11953), .IN2(n11957), .Q(n11956) );
  AND2X1 U11912 ( .IN1(n11958), .IN2(n11363), .Q(n11957) );
  OR2X1 U11913 ( .IN1(n10912), .IN2(n11959), .Q(n11958) );
  OR2X1 U11914 ( .IN1(n10513), .IN2(n10919), .Q(n11959) );
  OR2X1 U11915 ( .IN1(n10492), .IN2(n11362), .Q(n10919) );
  OR2X1 U11916 ( .IN1(n10512), .IN2(n11960), .Q(n11362) );
  AND2X1 U11917 ( .IN1(n3130), .IN2(n11961), .Q(n11960) );
  OR2X1 U11918 ( .IN1(n10509), .IN2(n10506), .Q(n11961) );
  OR2X1 U11919 ( .IN1(n11962), .IN2(n11963), .Q(n10506) );
  AND2X1 U11920 ( .IN1(n11964), .IN2(n11965), .Q(n11963) );
  AND2X1 U11921 ( .IN1(n11966), .IN2(n11967), .Q(n11964) );
  OR2X1 U11922 ( .IN1(n11968), .IN2(n11969), .Q(n11967) );
  OR2X1 U11923 ( .IN1(n11970), .IN2(n11971), .Q(n11966) );
  AND2X1 U11924 ( .IN1(n11972), .IN2(n11969), .Q(n11962) );
  AND2X1 U11925 ( .IN1(n11973), .IN2(n11974), .Q(n11972) );
  OR2X1 U11926 ( .IN1(n11965), .IN2(n11971), .Q(n11974) );
  AND2X1 U11927 ( .IN1(n11970), .IN2(n11975), .Q(n10509) );
  AND2X1 U11928 ( .IN1(n11976), .IN2(n11977), .Q(n11975) );
  OR2X1 U11929 ( .IN1(n11965), .IN2(n11968), .Q(n11976) );
  INVX0 U11930 ( .INP(n10495), .ZN(n10512) );
  OR2X1 U11931 ( .IN1(n11978), .IN2(n10499), .Q(n10495) );
  AND2X1 U11932 ( .IN1(n11979), .IN2(n11980), .Q(n11978) );
  OR2X1 U11933 ( .IN1(n11981), .IN2(n11982), .Q(n11980) );
  OR2X1 U11934 ( .IN1(n11983), .IN2(n11984), .Q(n11982) );
  AND2X1 U11935 ( .IN1(n11985), .IN2(n11986), .Q(n11984) );
  AND2X1 U11936 ( .IN1(n11987), .IN2(n11988), .Q(n11983) );
  AND2X1 U11937 ( .IN1(n11989), .IN2(n11990), .Q(n11979) );
  OR2X1 U11938 ( .IN1(n11987), .IN2(n11991), .Q(n11990) );
  OR2X1 U11939 ( .IN1(n11992), .IN2(n11993), .Q(n11991) );
  AND2X1 U11940 ( .IN1(n11981), .IN2(n11985), .Q(n11993) );
  OR2X1 U11941 ( .IN1(n11986), .IN2(n11994), .Q(n11989) );
  OR2X1 U11942 ( .IN1(n11995), .IN2(n11996), .Q(n11994) );
  AND2X1 U11943 ( .IN1(n11987), .IN2(n11985), .Q(n11996) );
  AND2X1 U11944 ( .IN1(n11981), .IN2(n11988), .Q(n11995) );
  OR2X1 U11945 ( .IN1(n10511), .IN2(n10499), .Q(n10912) );
  AND2X1 U11946 ( .IN1(n11997), .IN2(n11998), .Q(n10511) );
  INVX0 U11947 ( .INP(n11999), .ZN(n11998) );
  OR2X1 U11948 ( .IN1(n12000), .IN2(n11977), .Q(n11999) );
  OR2X1 U11949 ( .IN1(n11969), .IN2(n11971), .Q(n11977) );
  XNOR2X1 U11950 ( .IN1(n4569), .IN2(n9538), .Q(n11971) );
  OR2X1 U11951 ( .IN1(n12001), .IN2(n12002), .Q(n9538) );
  OR2X1 U11952 ( .IN1(n12003), .IN2(n12004), .Q(n12002) );
  AND2X1 U11953 ( .IN1(g165), .IN2(g219), .Q(n12004) );
  AND2X1 U11954 ( .IN1(g6231), .IN2(g213), .Q(n12003) );
  AND2X1 U11955 ( .IN1(g6313), .IN2(g216), .Q(n12001) );
  XNOR2X1 U11956 ( .IN1(n12005), .IN2(n9540), .Q(n11969) );
  OR2X1 U11957 ( .IN1(n12006), .IN2(n12007), .Q(n9540) );
  OR2X1 U11958 ( .IN1(n12008), .IN2(n12009), .Q(n12007) );
  AND2X1 U11959 ( .IN1(g165), .IN2(g228), .Q(n12009) );
  AND2X1 U11960 ( .IN1(g6231), .IN2(g222), .Q(n12008) );
  AND2X1 U11961 ( .IN1(g6313), .IN2(g225), .Q(n12006) );
  OR2X1 U11962 ( .IN1(n11965), .IN2(n11973), .Q(n12000) );
  OR2X1 U11963 ( .IN1(n11968), .IN2(n11970), .Q(n11973) );
  XOR2X1 U11964 ( .IN1(n4513), .IN2(n4380), .Q(n11970) );
  XNOR2X1 U11965 ( .IN1(n4322), .IN2(n9548), .Q(n11968) );
  OR2X1 U11966 ( .IN1(n12010), .IN2(n12011), .Q(n9548) );
  OR2X1 U11967 ( .IN1(n12012), .IN2(n12013), .Q(n12011) );
  AND2X1 U11968 ( .IN1(g165), .IN2(g201), .Q(n12013) );
  AND2X1 U11969 ( .IN1(g6231), .IN2(g195), .Q(n12012) );
  AND2X1 U11970 ( .IN1(g6313), .IN2(g198), .Q(n12010) );
  XNOR2X1 U11971 ( .IN1(n4328), .IN2(n9549), .Q(n11965) );
  OR2X1 U11972 ( .IN1(n12014), .IN2(n12015), .Q(n9549) );
  OR2X1 U11973 ( .IN1(n12016), .IN2(n12017), .Q(n12015) );
  AND2X1 U11974 ( .IN1(g165), .IN2(g210), .Q(n12017) );
  AND2X1 U11975 ( .IN1(g6231), .IN2(g204), .Q(n12016) );
  AND2X1 U11976 ( .IN1(g6313), .IN2(g207), .Q(n12014) );
  AND2X1 U11977 ( .IN1(n12018), .IN2(n12019), .Q(n11997) );
  AND2X1 U11978 ( .IN1(n11981), .IN2(n11987), .Q(n12019) );
  XOR2X1 U11979 ( .IN1(n10674), .IN2(n9539), .Q(n11987) );
  OR2X1 U11980 ( .IN1(n12020), .IN2(n12021), .Q(n9539) );
  OR2X1 U11981 ( .IN1(n12022), .IN2(n12023), .Q(n12021) );
  AND2X1 U11982 ( .IN1(g165), .IN2(g273), .Q(n12023) );
  AND2X1 U11983 ( .IN1(g6231), .IN2(g267), .Q(n12022) );
  AND2X1 U11984 ( .IN1(g6313), .IN2(g270), .Q(n12020) );
  XNOR2X1 U11985 ( .IN1(g117), .IN2(n9532), .Q(n11981) );
  OR2X1 U11986 ( .IN1(n12024), .IN2(n12025), .Q(n9532) );
  OR2X1 U11987 ( .IN1(n12026), .IN2(n12027), .Q(n12025) );
  AND2X1 U11988 ( .IN1(test_so14), .IN2(g165), .Q(n12027) );
  AND2X1 U11989 ( .IN1(g6231), .IN2(g249), .Q(n12026) );
  AND2X1 U11990 ( .IN1(g6313), .IN2(g252), .Q(n12024) );
  AND2X1 U11991 ( .IN1(n11985), .IN2(n11992), .Q(n12018) );
  AND2X1 U11992 ( .IN1(n11986), .IN2(n11988), .Q(n11992) );
  XOR2X1 U11993 ( .IN1(n4392), .IN2(n9554), .Q(n11988) );
  OR2X1 U11994 ( .IN1(n12028), .IN2(n12029), .Q(n9554) );
  OR2X1 U11995 ( .IN1(n12030), .IN2(n12031), .Q(n12029) );
  AND2X1 U11996 ( .IN1(g165), .IN2(g246), .Q(n12031) );
  AND2X1 U11997 ( .IN1(g6231), .IN2(g240), .Q(n12030) );
  AND2X1 U11998 ( .IN1(g6313), .IN2(g243), .Q(n12028) );
  XOR2X1 U11999 ( .IN1(n4376), .IN2(n9531), .Q(n11986) );
  OR2X1 U12000 ( .IN1(n12032), .IN2(n12033), .Q(n9531) );
  OR2X1 U12001 ( .IN1(n12034), .IN2(n12035), .Q(n12033) );
  AND2X1 U12002 ( .IN1(g165), .IN2(g237), .Q(n12035) );
  AND2X1 U12003 ( .IN1(g6231), .IN2(g231), .Q(n12034) );
  AND2X1 U12004 ( .IN1(g6313), .IN2(g234), .Q(n12032) );
  XOR2X1 U12005 ( .IN1(n4290), .IN2(n9533), .Q(n11985) );
  OR2X1 U12006 ( .IN1(n12036), .IN2(n12037), .Q(n9533) );
  OR2X1 U12007 ( .IN1(n12038), .IN2(n12039), .Q(n12037) );
  AND2X1 U12008 ( .IN1(g165), .IN2(g264), .Q(n12039) );
  AND2X1 U12009 ( .IN1(g6231), .IN2(g258), .Q(n12038) );
  AND2X1 U12010 ( .IN1(g6313), .IN2(g261), .Q(n12036) );
  AND2X1 U12011 ( .IN1(n4388), .IN2(n12040), .Q(n11953) );
  AND2X1 U12012 ( .IN1(n12041), .IN2(n12042), .Q(g29112) );
  OR2X1 U12013 ( .IN1(n3159), .IN2(g2129), .Q(n12042) );
  AND2X1 U12014 ( .IN1(n11527), .IN2(n1291), .Q(n12041) );
  INVX0 U12015 ( .INP(n11535), .ZN(n1291) );
  AND2X1 U12016 ( .IN1(g2129), .IN2(n3159), .Q(n11535) );
  AND2X1 U12017 ( .IN1(n12043), .IN2(n12044), .Q(g29111) );
  OR2X1 U12018 ( .IN1(n3163), .IN2(g1435), .Q(n12044) );
  AND2X1 U12019 ( .IN1(n11529), .IN2(n1005), .Q(n12043) );
  INVX0 U12020 ( .INP(n11537), .ZN(n1005) );
  AND2X1 U12021 ( .IN1(g1435), .IN2(n3163), .Q(n11537) );
  AND2X1 U12022 ( .IN1(n12045), .IN2(n12046), .Q(g29110) );
  OR2X1 U12023 ( .IN1(n3167), .IN2(test_so36), .Q(n12046) );
  AND2X1 U12024 ( .IN1(n11531), .IN2(n716), .Q(n12045) );
  INVX0 U12025 ( .INP(n11539), .ZN(n716) );
  AND2X1 U12026 ( .IN1(n3167), .IN2(test_so36), .Q(n11539) );
  AND2X1 U12027 ( .IN1(n12047), .IN2(n12048), .Q(g29109) );
  OR2X1 U12028 ( .IN1(n3171), .IN2(g61), .Q(n12048) );
  AND2X1 U12029 ( .IN1(n11533), .IN2(n407), .Q(n12047) );
  INVX0 U12030 ( .INP(n11541), .ZN(n407) );
  AND2X1 U12031 ( .IN1(g61), .IN2(n3171), .Q(n11541) );
  OR2X1 U12032 ( .IN1(n12049), .IN2(n12050), .Q(g28788) );
  AND2X1 U12033 ( .IN1(n12051), .IN2(n10833), .Q(n12050) );
  AND2X1 U12034 ( .IN1(n12052), .IN2(g2501), .Q(n12049) );
  OR2X1 U12035 ( .IN1(n4509), .IN2(n12053), .Q(n12052) );
  OR2X1 U12036 ( .IN1(n12054), .IN2(n12055), .Q(g28783) );
  AND2X1 U12037 ( .IN1(n12051), .IN2(n10398), .Q(n12055) );
  AND2X1 U12038 ( .IN1(n12056), .IN2(g2503), .Q(n12054) );
  OR2X1 U12039 ( .IN1(n4524), .IN2(n12053), .Q(n12056) );
  OR2X1 U12040 ( .IN1(n12057), .IN2(n12058), .Q(g28782) );
  AND2X1 U12041 ( .IN1(test_so80), .IN2(n4509), .Q(n12058) );
  AND2X1 U12042 ( .IN1(n4606), .IN2(n12059), .Q(n12057) );
  OR2X1 U12043 ( .IN1(n12060), .IN2(n12061), .Q(g28778) );
  AND2X1 U12044 ( .IN1(n12062), .IN2(n10403), .Q(n12061) );
  AND2X1 U12045 ( .IN1(n12063), .IN2(g1807), .Q(n12060) );
  OR2X1 U12046 ( .IN1(n4511), .IN2(n12064), .Q(n12063) );
  OR2X1 U12047 ( .IN1(n12065), .IN2(n12066), .Q(g28774) );
  AND2X1 U12048 ( .IN1(n12051), .IN2(n10408), .Q(n12066) );
  AND2X1 U12049 ( .IN1(n12067), .IN2(g2502), .Q(n12065) );
  OR2X1 U12050 ( .IN1(n4516), .IN2(n12053), .Q(n12067) );
  OR2X1 U12051 ( .IN1(n11559), .IN2(n12068), .Q(n12053) );
  OR2X1 U12052 ( .IN1(n12069), .IN2(n12070), .Q(g28773) );
  AND2X1 U12053 ( .IN1(n4524), .IN2(g2486), .Q(n12070) );
  AND2X1 U12054 ( .IN1(g7264), .IN2(n12059), .Q(n12069) );
  OR2X1 U12055 ( .IN1(n12071), .IN2(n12072), .Q(g28772) );
  AND2X1 U12056 ( .IN1(n12062), .IN2(n10412), .Q(n12072) );
  AND2X1 U12057 ( .IN1(n12073), .IN2(g1809), .Q(n12071) );
  OR2X1 U12058 ( .IN1(n4525), .IN2(n12064), .Q(n12073) );
  OR2X1 U12059 ( .IN1(n12074), .IN2(n12075), .Q(g28771) );
  AND2X1 U12060 ( .IN1(n4511), .IN2(g1795), .Q(n12075) );
  AND2X1 U12061 ( .IN1(n4618), .IN2(n12076), .Q(n12074) );
  OR2X1 U12062 ( .IN1(n12077), .IN2(n12078), .Q(g28767) );
  AND2X1 U12063 ( .IN1(n12079), .IN2(g1088), .Q(n12078) );
  AND2X1 U12064 ( .IN1(n12080), .IN2(g1113), .Q(n12077) );
  OR2X1 U12065 ( .IN1(n4381), .IN2(n12081), .Q(n12080) );
  OR2X1 U12066 ( .IN1(n12082), .IN2(n12083), .Q(g28763) );
  AND2X1 U12067 ( .IN1(n4516), .IN2(g2483), .Q(n12083) );
  AND2X1 U12068 ( .IN1(g5555), .IN2(n12059), .Q(n12082) );
  OR2X1 U12069 ( .IN1(n12084), .IN2(n12051), .Q(n12059) );
  INVX0 U12070 ( .INP(n12085), .ZN(n12051) );
  OR2X1 U12071 ( .IN1(n11561), .IN2(n12068), .Q(n12085) );
  OR2X1 U12072 ( .IN1(n12086), .IN2(n9121), .Q(n12068) );
  AND2X1 U12073 ( .IN1(n12087), .IN2(n11561), .Q(n12084) );
  OR2X1 U12074 ( .IN1(n12088), .IN2(n12089), .Q(n11561) );
  OR2X1 U12075 ( .IN1(n12090), .IN2(n12091), .Q(n12089) );
  AND2X1 U12076 ( .IN1(g7264), .IN2(g2486), .Q(n12091) );
  AND2X1 U12077 ( .IN1(test_so80), .IN2(n4606), .Q(n12090) );
  AND2X1 U12078 ( .IN1(g5555), .IN2(g2483), .Q(n12088) );
  OR2X1 U12079 ( .IN1(n12092), .IN2(n9121), .Q(n12087) );
  INVX0 U12080 ( .INP(n12093), .ZN(n12092) );
  OR2X1 U12081 ( .IN1(n11559), .IN2(n12086), .Q(n12093) );
  INVX0 U12082 ( .INP(n12094), .ZN(n12086) );
  OR2X1 U12083 ( .IN1(n12095), .IN2(n12096), .Q(n12094) );
  AND2X1 U12084 ( .IN1(n12097), .IN2(n11552), .Q(n12096) );
  AND2X1 U12085 ( .IN1(n11563), .IN2(n10844), .Q(n12097) );
  OR2X1 U12086 ( .IN1(n9091), .IN2(n10386), .Q(n10844) );
  OR2X1 U12087 ( .IN1(n12098), .IN2(n12099), .Q(n10386) );
  OR2X1 U12088 ( .IN1(n12100), .IN2(n12101), .Q(n12099) );
  AND2X1 U12089 ( .IN1(n8694), .IN2(g2241), .Q(n12101) );
  AND2X1 U12090 ( .IN1(n8696), .IN2(g6837), .Q(n12100) );
  AND2X1 U12091 ( .IN1(n8695), .IN2(test_so73), .Q(n12098) );
  INVX0 U12092 ( .INP(n11560), .ZN(n11563) );
  AND2X1 U12093 ( .IN1(n11560), .IN2(n4285), .Q(n12095) );
  OR2X1 U12094 ( .IN1(n12102), .IN2(n12103), .Q(n11560) );
  OR2X1 U12095 ( .IN1(n11693), .IN2(n10555), .Q(n12103) );
  OR2X1 U12096 ( .IN1(n12104), .IN2(n12105), .Q(n11559) );
  OR2X1 U12097 ( .IN1(n12106), .IN2(n12107), .Q(n12105) );
  AND2X1 U12098 ( .IN1(n8785), .IN2(n10408), .Q(n12107) );
  AND2X1 U12099 ( .IN1(n8784), .IN2(n10833), .Q(n12106) );
  AND2X1 U12100 ( .IN1(n8775), .IN2(n10398), .Q(n12104) );
  OR2X1 U12101 ( .IN1(n12108), .IN2(n12109), .Q(g28761) );
  AND2X1 U12102 ( .IN1(n12062), .IN2(n10419), .Q(n12109) );
  AND2X1 U12103 ( .IN1(n12110), .IN2(g1808), .Q(n12108) );
  OR2X1 U12104 ( .IN1(n4518), .IN2(n12064), .Q(n12110) );
  INVX0 U12105 ( .INP(n12111), .ZN(n12064) );
  AND2X1 U12106 ( .IN1(n11582), .IN2(n12112), .Q(n12111) );
  OR2X1 U12107 ( .IN1(n12113), .IN2(n12114), .Q(g28760) );
  AND2X1 U12108 ( .IN1(n4525), .IN2(g1792), .Q(n12114) );
  AND2X1 U12109 ( .IN1(g7014), .IN2(n12076), .Q(n12113) );
  OR2X1 U12110 ( .IN1(n12115), .IN2(n12116), .Q(g28759) );
  AND2X1 U12111 ( .IN1(n12079), .IN2(g6712), .Q(n12116) );
  AND2X1 U12112 ( .IN1(n12117), .IN2(g1115), .Q(n12115) );
  OR2X1 U12113 ( .IN1(n4364), .IN2(n12081), .Q(n12117) );
  OR2X1 U12114 ( .IN1(n12118), .IN2(n12119), .Q(g28758) );
  AND2X1 U12115 ( .IN1(n12120), .IN2(g1088), .Q(n12119) );
  AND2X1 U12116 ( .IN1(n4381), .IN2(g1101), .Q(n12118) );
  OR2X1 U12117 ( .IN1(n12121), .IN2(n12122), .Q(g28754) );
  AND2X1 U12118 ( .IN1(n12123), .IN2(n10465), .Q(n12122) );
  AND2X1 U12119 ( .IN1(n12124), .IN2(g426), .Q(n12121) );
  OR2X1 U12120 ( .IN1(n4506), .IN2(n12125), .Q(n12124) );
  OR2X1 U12121 ( .IN1(n12126), .IN2(n12127), .Q(g28749) );
  AND2X1 U12122 ( .IN1(n4518), .IN2(g1789), .Q(n12127) );
  AND2X1 U12123 ( .IN1(g5511), .IN2(n12076), .Q(n12126) );
  OR2X1 U12124 ( .IN1(n12128), .IN2(n12062), .Q(n12076) );
  AND2X1 U12125 ( .IN1(n11585), .IN2(n12112), .Q(n12062) );
  AND2X1 U12126 ( .IN1(g1690), .IN2(n12129), .Q(n12112) );
  INVX0 U12127 ( .INP(n12130), .ZN(n11585) );
  AND2X1 U12128 ( .IN1(n12131), .IN2(n12130), .Q(n12128) );
  OR2X1 U12129 ( .IN1(n12132), .IN2(n12133), .Q(n12130) );
  OR2X1 U12130 ( .IN1(n12134), .IN2(n12135), .Q(n12133) );
  AND2X1 U12131 ( .IN1(g7014), .IN2(g1792), .Q(n12135) );
  AND2X1 U12132 ( .IN1(n4618), .IN2(g1795), .Q(n12134) );
  AND2X1 U12133 ( .IN1(g5511), .IN2(g1789), .Q(n12132) );
  OR2X1 U12134 ( .IN1(n12136), .IN2(n4386), .Q(n12131) );
  AND2X1 U12135 ( .IN1(n11582), .IN2(n12129), .Q(n12136) );
  OR2X1 U12136 ( .IN1(n12137), .IN2(n12138), .Q(n12129) );
  AND2X1 U12137 ( .IN1(n12139), .IN2(n11584), .Q(n12138) );
  AND2X1 U12138 ( .IN1(n12140), .IN2(n10430), .Q(n12139) );
  OR2X1 U12139 ( .IN1(n9090), .IN2(n9503), .Q(n10430) );
  OR2X1 U12140 ( .IN1(n12141), .IN2(n12142), .Q(n9503) );
  OR2X1 U12141 ( .IN1(n12143), .IN2(n12144), .Q(n12142) );
  AND2X1 U12142 ( .IN1(n8705), .IN2(g1547), .Q(n12144) );
  AND2X1 U12143 ( .IN1(n8707), .IN2(g6573), .Q(n12143) );
  AND2X1 U12144 ( .IN1(n8706), .IN2(g6782), .Q(n12141) );
  INVX0 U12145 ( .INP(n11579), .ZN(n12140) );
  AND2X1 U12146 ( .IN1(n11579), .IN2(n4284), .Q(n12137) );
  OR2X1 U12147 ( .IN1(n12145), .IN2(n12146), .Q(n11579) );
  OR2X1 U12148 ( .IN1(n11800), .IN2(n10589), .Q(n12146) );
  INVX0 U12149 ( .INP(n12147), .ZN(n11582) );
  OR2X1 U12150 ( .IN1(n12148), .IN2(n12149), .Q(n12147) );
  OR2X1 U12151 ( .IN1(n12150), .IN2(n12151), .Q(n12149) );
  AND2X1 U12152 ( .IN1(n8790), .IN2(n10419), .Q(n12151) );
  AND2X1 U12153 ( .IN1(n8789), .IN2(n10403), .Q(n12150) );
  AND2X1 U12154 ( .IN1(n8778), .IN2(n10412), .Q(n12148) );
  OR2X1 U12155 ( .IN1(n12152), .IN2(n12153), .Q(g28747) );
  AND2X1 U12156 ( .IN1(n12079), .IN2(g5472), .Q(n12153) );
  AND2X1 U12157 ( .IN1(n12154), .IN2(g1114), .Q(n12152) );
  OR2X1 U12158 ( .IN1(n4363), .IN2(n12081), .Q(n12154) );
  OR2X1 U12159 ( .IN1(n11600), .IN2(n12155), .Q(n12081) );
  OR2X1 U12160 ( .IN1(n12156), .IN2(n12157), .Q(g28746) );
  AND2X1 U12161 ( .IN1(n12120), .IN2(g6712), .Q(n12157) );
  AND2X1 U12162 ( .IN1(n4364), .IN2(g1098), .Q(n12156) );
  OR2X1 U12163 ( .IN1(n12158), .IN2(n12159), .Q(g28745) );
  AND2X1 U12164 ( .IN1(n12123), .IN2(n10899), .Q(n12159) );
  AND2X1 U12165 ( .IN1(n12160), .IN2(g428), .Q(n12158) );
  OR2X1 U12166 ( .IN1(n4499), .IN2(n12125), .Q(n12160) );
  OR2X1 U12167 ( .IN1(n12161), .IN2(n12162), .Q(g28744) );
  AND2X1 U12168 ( .IN1(n4506), .IN2(g414), .Q(n12162) );
  AND2X1 U12169 ( .IN1(n4640), .IN2(n12163), .Q(n12161) );
  OR2X1 U12170 ( .IN1(n12164), .IN2(n12165), .Q(g28738) );
  AND2X1 U12171 ( .IN1(n12120), .IN2(g5472), .Q(n12165) );
  OR2X1 U12172 ( .IN1(n12166), .IN2(n12079), .Q(n12120) );
  INVX0 U12173 ( .INP(n12167), .ZN(n12079) );
  OR2X1 U12174 ( .IN1(n11602), .IN2(n12155), .Q(n12167) );
  OR2X1 U12175 ( .IN1(n4387), .IN2(n12168), .Q(n12155) );
  AND2X1 U12176 ( .IN1(n12169), .IN2(n11602), .Q(n12166) );
  OR2X1 U12177 ( .IN1(n12170), .IN2(n12171), .Q(n11602) );
  OR2X1 U12178 ( .IN1(n12172), .IN2(n12173), .Q(n12171) );
  AND2X1 U12179 ( .IN1(g6712), .IN2(g1098), .Q(n12173) );
  AND2X1 U12180 ( .IN1(g5472), .IN2(g1095), .Q(n12172) );
  AND2X1 U12181 ( .IN1(g1088), .IN2(g1101), .Q(n12170) );
  OR2X1 U12182 ( .IN1(n12174), .IN2(n4387), .Q(n12169) );
  INVX0 U12183 ( .INP(n12175), .ZN(n12174) );
  OR2X1 U12184 ( .IN1(n11600), .IN2(n12168), .Q(n12175) );
  INVX0 U12185 ( .INP(n12176), .ZN(n12168) );
  OR2X1 U12186 ( .IN1(n12177), .IN2(n12178), .Q(n12176) );
  AND2X1 U12187 ( .IN1(n12179), .IN2(n11593), .Q(n12178) );
  AND2X1 U12188 ( .IN1(n11604), .IN2(n10245), .Q(n12179) );
  OR2X1 U12189 ( .IN1(n9089), .IN2(n9512), .Q(n10245) );
  OR2X1 U12190 ( .IN1(n12180), .IN2(n12181), .Q(n9512) );
  OR2X1 U12191 ( .IN1(n12182), .IN2(n12183), .Q(n12181) );
  AND2X1 U12192 ( .IN1(n8718), .IN2(g6368), .Q(n12183) );
  INVX0 U12193 ( .INP(n12184), .ZN(n12182) );
  OR2X1 U12194 ( .IN1(n4312), .IN2(test_so33), .Q(n12184) );
  AND2X1 U12195 ( .IN1(test_so31), .IN2(n8717), .Q(n12180) );
  INVX0 U12196 ( .INP(n11601), .ZN(n11604) );
  AND2X1 U12197 ( .IN1(n11601), .IN2(n4283), .Q(n12177) );
  OR2X1 U12198 ( .IN1(n12185), .IN2(n12186), .Q(n11601) );
  OR2X1 U12199 ( .IN1(n10629), .IN2(n11924), .Q(n12186) );
  OR2X1 U12200 ( .IN1(n12187), .IN2(n12188), .Q(n11600) );
  OR2X1 U12201 ( .IN1(n12189), .IN2(n12190), .Q(n12188) );
  AND2X1 U12202 ( .IN1(n8781), .IN2(g6712), .Q(n12190) );
  AND2X1 U12203 ( .IN1(n8796), .IN2(g5472), .Q(n12189) );
  AND2X1 U12204 ( .IN1(n8795), .IN2(g1088), .Q(n12187) );
  AND2X1 U12205 ( .IN1(n4363), .IN2(g1095), .Q(n12164) );
  OR2X1 U12206 ( .IN1(n12191), .IN2(n12192), .Q(g28736) );
  AND2X1 U12207 ( .IN1(n12123), .IN2(n10475), .Q(n12192) );
  AND2X1 U12208 ( .IN1(test_so17), .IN2(n12193), .Q(n12191) );
  OR2X1 U12209 ( .IN1(n4520), .IN2(n12125), .Q(n12193) );
  INVX0 U12210 ( .INP(n12194), .ZN(n12125) );
  AND2X1 U12211 ( .IN1(n11620), .IN2(n12195), .Q(n12194) );
  OR2X1 U12212 ( .IN1(n12196), .IN2(n12197), .Q(g28735) );
  AND2X1 U12213 ( .IN1(n4499), .IN2(g411), .Q(n12197) );
  AND2X1 U12214 ( .IN1(g6447), .IN2(n12163), .Q(n12196) );
  OR2X1 U12215 ( .IN1(n12198), .IN2(n12199), .Q(g28732) );
  AND2X1 U12216 ( .IN1(n4520), .IN2(g408), .Q(n12199) );
  AND2X1 U12217 ( .IN1(g5437), .IN2(n12163), .Q(n12198) );
  OR2X1 U12218 ( .IN1(n12200), .IN2(n12123), .Q(n12163) );
  AND2X1 U12219 ( .IN1(n11623), .IN2(n12195), .Q(n12123) );
  AND2X1 U12220 ( .IN1(g309), .IN2(n12201), .Q(n12195) );
  INVX0 U12221 ( .INP(n12202), .ZN(n11623) );
  AND2X1 U12222 ( .IN1(n12203), .IN2(n12202), .Q(n12200) );
  OR2X1 U12223 ( .IN1(n12204), .IN2(n12205), .Q(n12202) );
  OR2X1 U12224 ( .IN1(n12206), .IN2(n12207), .Q(n12205) );
  AND2X1 U12225 ( .IN1(g6447), .IN2(g411), .Q(n12207) );
  AND2X1 U12226 ( .IN1(n4640), .IN2(g414), .Q(n12206) );
  AND2X1 U12227 ( .IN1(g5437), .IN2(g408), .Q(n12204) );
  OR2X1 U12228 ( .IN1(n12208), .IN2(n4388), .Q(n12203) );
  AND2X1 U12229 ( .IN1(n11620), .IN2(n12201), .Q(n12208) );
  OR2X1 U12230 ( .IN1(n12209), .IN2(n12210), .Q(n12201) );
  AND2X1 U12231 ( .IN1(n12211), .IN2(n11622), .Q(n12210) );
  AND2X1 U12232 ( .IN1(n12212), .IN2(n10486), .Q(n12211) );
  OR2X1 U12233 ( .IN1(n9088), .IN2(n10221), .Q(n10486) );
  OR2X1 U12234 ( .IN1(n12213), .IN2(n12214), .Q(n10221) );
  OR2X1 U12235 ( .IN1(n12215), .IN2(n12216), .Q(n12214) );
  AND2X1 U12236 ( .IN1(n8728), .IN2(g165), .Q(n12216) );
  AND2X1 U12237 ( .IN1(n8730), .IN2(g6231), .Q(n12215) );
  AND2X1 U12238 ( .IN1(n8729), .IN2(g6313), .Q(n12213) );
  INVX0 U12239 ( .INP(n11617), .ZN(n12212) );
  AND2X1 U12240 ( .IN1(n11617), .IN2(n4282), .Q(n12209) );
  OR2X1 U12241 ( .IN1(n12217), .IN2(n12218), .Q(n11617) );
  OR2X1 U12242 ( .IN1(n12005), .IN2(n10674), .Q(n12218) );
  INVX0 U12243 ( .INP(n12219), .ZN(n11620) );
  OR2X1 U12244 ( .IN1(n12220), .IN2(n12221), .Q(n12219) );
  OR2X1 U12245 ( .IN1(n12222), .IN2(n12223), .Q(n12221) );
  AND2X1 U12246 ( .IN1(n8803), .IN2(n10465), .Q(n12223) );
  AND2X1 U12247 ( .IN1(n8804), .IN2(n10899), .Q(n12222) );
  INVX0 U12248 ( .INP(n12224), .ZN(n12220) );
  OR2X1 U12249 ( .IN1(n4520), .IN2(test_so17), .Q(n12224) );
  AND2X1 U12250 ( .IN1(n12225), .IN2(n12226), .Q(g28668) );
  XOR2X1 U12251 ( .IN1(n12227), .IN2(n4418), .Q(n12225) );
  OR2X1 U12252 ( .IN1(n4396), .IN2(n12228), .Q(n12227) );
  AND2X1 U12253 ( .IN1(n12229), .IN2(n11527), .Q(g28637) );
  XNOR2X1 U12254 ( .IN1(n12230), .IN2(n8806), .Q(n12229) );
  AND2X1 U12255 ( .IN1(n12231), .IN2(n11529), .Q(g28636) );
  XNOR2X1 U12256 ( .IN1(n12232), .IN2(n8810), .Q(n12231) );
  AND2X1 U12257 ( .IN1(n12233), .IN2(n11531), .Q(g28635) );
  XNOR2X1 U12258 ( .IN1(n12234), .IN2(n8814), .Q(n12233) );
  AND2X1 U12259 ( .IN1(n12235), .IN2(n11533), .Q(g28634) );
  XNOR2X1 U12260 ( .IN1(n12236), .IN2(n8818), .Q(n12235) );
  OR2X1 U12261 ( .IN1(n12237), .IN2(n12238), .Q(g28425) );
  AND2X1 U12262 ( .IN1(n486), .IN2(g3109), .Q(n12238) );
  AND2X1 U12263 ( .IN1(n4494), .IN2(g3102), .Q(n12237) );
  OR2X1 U12264 ( .IN1(n12239), .IN2(n12240), .Q(g28421) );
  AND2X1 U12265 ( .IN1(n486), .IN2(g8030), .Q(n12240) );
  AND2X1 U12266 ( .IN1(n4383), .IN2(test_so7), .Q(n12239) );
  OR2X1 U12267 ( .IN1(n12241), .IN2(n12242), .Q(g28420) );
  AND2X1 U12268 ( .IN1(n486), .IN2(g8106), .Q(n12242) );
  INVX0 U12269 ( .INP(n11461), .ZN(n486) );
  OR2X1 U12270 ( .IN1(n12243), .IN2(n12244), .Q(n11461) );
  AND2X1 U12271 ( .IN1(n12245), .IN2(n4548), .Q(n12244) );
  AND2X1 U12272 ( .IN1(n12246), .IN2(n12247), .Q(n12245) );
  INVX0 U12273 ( .INP(n12248), .ZN(n12247) );
  AND2X1 U12274 ( .IN1(g21851), .IN2(g6750), .Q(n12248) );
  OR2X1 U12275 ( .IN1(n8269), .IN2(n12249), .Q(n12246) );
  AND2X1 U12276 ( .IN1(n8268), .IN2(g1186), .Q(n12243) );
  AND2X1 U12277 ( .IN1(n4382), .IN2(g3100), .Q(n12241) );
  OR2X1 U12278 ( .IN1(n12250), .IN2(n12251), .Q(g28371) );
  AND2X1 U12279 ( .IN1(n12252), .IN2(g2624), .Q(n12251) );
  AND2X1 U12280 ( .IN1(n4299), .IN2(g2694), .Q(n12250) );
  OR2X1 U12281 ( .IN1(n12253), .IN2(n12254), .Q(g28368) );
  AND2X1 U12282 ( .IN1(n12252), .IN2(g7390), .Q(n12254) );
  AND2X1 U12283 ( .IN1(n4370), .IN2(g2691), .Q(n12253) );
  OR2X1 U12284 ( .IN1(n12255), .IN2(n12256), .Q(g28367) );
  AND2X1 U12285 ( .IN1(n12257), .IN2(g2624), .Q(n12256) );
  AND2X1 U12286 ( .IN1(n4299), .IN2(g2685), .Q(n12255) );
  OR2X1 U12287 ( .IN1(n12258), .IN2(n12259), .Q(g28366) );
  AND2X1 U12288 ( .IN1(n12260), .IN2(g1930), .Q(n12259) );
  AND2X1 U12289 ( .IN1(n4366), .IN2(g2000), .Q(n12258) );
  OR2X1 U12290 ( .IN1(n12261), .IN2(n12262), .Q(g28364) );
  AND2X1 U12291 ( .IN1(n12252), .IN2(n11411), .Q(n12262) );
  OR2X1 U12292 ( .IN1(n12263), .IN2(n12264), .Q(n12252) );
  AND2X1 U12293 ( .IN1(n9889), .IN2(n12265), .Q(n12264) );
  AND2X1 U12294 ( .IN1(n3252), .IN2(n12266), .Q(n12263) );
  AND2X1 U12295 ( .IN1(n4314), .IN2(g2688), .Q(n12261) );
  OR2X1 U12296 ( .IN1(n12267), .IN2(n12268), .Q(g28363) );
  AND2X1 U12297 ( .IN1(n12257), .IN2(g7390), .Q(n12268) );
  AND2X1 U12298 ( .IN1(n4370), .IN2(test_so90), .Q(n12267) );
  OR2X1 U12299 ( .IN1(n12269), .IN2(n12270), .Q(g28362) );
  AND2X1 U12300 ( .IN1(n12260), .IN2(g7194), .Q(n12270) );
  AND2X1 U12301 ( .IN1(n4315), .IN2(g1997), .Q(n12269) );
  OR2X1 U12302 ( .IN1(n12271), .IN2(n12272), .Q(g28361) );
  AND2X1 U12303 ( .IN1(n12273), .IN2(g1930), .Q(n12272) );
  AND2X1 U12304 ( .IN1(n4366), .IN2(g1991), .Q(n12271) );
  OR2X1 U12305 ( .IN1(n12274), .IN2(n12275), .Q(g28360) );
  AND2X1 U12306 ( .IN1(n12276), .IN2(g1236), .Q(n12275) );
  AND2X1 U12307 ( .IN1(n4300), .IN2(g1306), .Q(n12274) );
  OR2X1 U12308 ( .IN1(n12277), .IN2(n12278), .Q(g28358) );
  AND2X1 U12309 ( .IN1(n4314), .IN2(g2679), .Q(n12278) );
  AND2X1 U12310 ( .IN1(g7302), .IN2(n12257), .Q(n12277) );
  OR2X1 U12311 ( .IN1(n12279), .IN2(n12280), .Q(n12257) );
  AND2X1 U12312 ( .IN1(n9879), .IN2(n12265), .Q(n12280) );
  AND2X1 U12313 ( .IN1(n3260), .IN2(n12281), .Q(n12279) );
  INVX0 U12314 ( .INP(n10226), .ZN(n12281) );
  OR2X1 U12315 ( .IN1(n12282), .IN2(n12283), .Q(n10226) );
  OR2X1 U12316 ( .IN1(n12284), .IN2(n12285), .Q(n12283) );
  AND2X1 U12317 ( .IN1(n12286), .IN2(n12287), .Q(n12285) );
  AND2X1 U12318 ( .IN1(n12288), .IN2(n12289), .Q(n12286) );
  OR2X1 U12319 ( .IN1(n12290), .IN2(n12291), .Q(n12288) );
  AND2X1 U12320 ( .IN1(n12292), .IN2(n12293), .Q(n12290) );
  OR2X1 U12321 ( .IN1(n12294), .IN2(n12295), .Q(n12293) );
  AND2X1 U12322 ( .IN1(n12296), .IN2(n12297), .Q(n12284) );
  OR2X1 U12323 ( .IN1(n12298), .IN2(n12299), .Q(n12297) );
  AND2X1 U12324 ( .IN1(n12300), .IN2(n12301), .Q(n12299) );
  OR2X1 U12325 ( .IN1(n12302), .IN2(n12292), .Q(n12300) );
  AND2X1 U12326 ( .IN1(n12303), .IN2(n12304), .Q(n12302) );
  AND2X1 U12327 ( .IN1(n12305), .IN2(n12306), .Q(n12298) );
  AND2X1 U12328 ( .IN1(n12294), .IN2(n12295), .Q(n12306) );
  AND2X1 U12329 ( .IN1(n12292), .IN2(n12307), .Q(n12305) );
  OR2X1 U12330 ( .IN1(n12308), .IN2(n12309), .Q(n12282) );
  AND2X1 U12331 ( .IN1(n12310), .IN2(n12304), .Q(n12309) );
  AND2X1 U12332 ( .IN1(n12311), .IN2(n12312), .Q(n12310) );
  OR2X1 U12333 ( .IN1(n12313), .IN2(n12314), .Q(n12312) );
  AND2X1 U12334 ( .IN1(n12315), .IN2(n12316), .Q(n12313) );
  AND2X1 U12335 ( .IN1(n12317), .IN2(n12318), .Q(n12308) );
  OR2X1 U12336 ( .IN1(n12319), .IN2(n12320), .Q(n12318) );
  AND2X1 U12337 ( .IN1(n12321), .IN2(n12315), .Q(n12320) );
  OR2X1 U12338 ( .IN1(n12322), .IN2(n12323), .Q(n12315) );
  AND2X1 U12339 ( .IN1(n12324), .IN2(n12287), .Q(n12322) );
  AND2X1 U12340 ( .IN1(n12325), .IN2(n12314), .Q(n12319) );
  OR2X1 U12341 ( .IN1(n12326), .IN2(n12327), .Q(n12314) );
  AND2X1 U12342 ( .IN1(n12323), .IN2(n12287), .Q(n12327) );
  AND2X1 U12343 ( .IN1(n12307), .IN2(n12296), .Q(n12326) );
  AND2X1 U12344 ( .IN1(n12266), .IN2(n12328), .Q(n3260) );
  INVX0 U12345 ( .INP(n12329), .ZN(n12328) );
  OR2X1 U12346 ( .IN1(n10222), .IN2(n12330), .Q(n12329) );
  INVX0 U12347 ( .INP(n12331), .ZN(n12330) );
  OR2X1 U12348 ( .IN1(n10384), .IN2(n12332), .Q(n12331) );
  OR2X1 U12349 ( .IN1(n12333), .IN2(n12334), .Q(n10384) );
  OR2X1 U12350 ( .IN1(n12335), .IN2(n12336), .Q(n12334) );
  AND2X1 U12351 ( .IN1(n12337), .IN2(n12287), .Q(n12336) );
  OR2X1 U12352 ( .IN1(n12338), .IN2(n12339), .Q(n12337) );
  AND2X1 U12353 ( .IN1(n12317), .IN2(n12340), .Q(n12339) );
  OR2X1 U12354 ( .IN1(n12341), .IN2(n12342), .Q(n12340) );
  OR2X1 U12355 ( .IN1(n12343), .IN2(n12344), .Q(n12342) );
  AND2X1 U12356 ( .IN1(n12291), .IN2(n12307), .Q(n12344) );
  AND2X1 U12357 ( .IN1(n12294), .IN2(n12345), .Q(n12291) );
  AND2X1 U12358 ( .IN1(n12295), .IN2(n12303), .Q(n12345) );
  AND2X1 U12359 ( .IN1(n12346), .IN2(n12292), .Q(n12343) );
  AND2X1 U12360 ( .IN1(n12311), .IN2(n12323), .Q(n12341) );
  AND2X1 U12361 ( .IN1(n12325), .IN2(n12301), .Q(n12338) );
  AND2X1 U12362 ( .IN1(n12347), .IN2(n12311), .Q(n12335) );
  INVX0 U12363 ( .INP(n12295), .ZN(n12311) );
  AND2X1 U12364 ( .IN1(n12348), .IN2(n12289), .Q(n12347) );
  OR2X1 U12365 ( .IN1(n12349), .IN2(n12350), .Q(n12348) );
  AND2X1 U12366 ( .IN1(n12317), .IN2(n12316), .Q(n12350) );
  AND2X1 U12367 ( .IN1(n12296), .IN2(n12294), .Q(n12349) );
  AND2X1 U12368 ( .IN1(n12351), .IN2(n12304), .Q(n12333) );
  OR2X1 U12369 ( .IN1(n12352), .IN2(n12353), .Q(n12351) );
  AND2X1 U12370 ( .IN1(n12296), .IN2(n12354), .Q(n12353) );
  OR2X1 U12371 ( .IN1(n12355), .IN2(n12356), .Q(n12354) );
  OR2X1 U12372 ( .IN1(n12357), .IN2(n12358), .Q(n12356) );
  AND2X1 U12373 ( .IN1(n12346), .IN2(n12325), .Q(n12358) );
  AND2X1 U12374 ( .IN1(n12295), .IN2(n12316), .Q(n12325) );
  AND2X1 U12375 ( .IN1(n12359), .IN2(n12303), .Q(n12357) );
  AND2X1 U12376 ( .IN1(n12323), .IN2(n12295), .Q(n12359) );
  OR2X1 U12377 ( .IN1(n12360), .IN2(n12361), .Q(n12295) );
  OR2X1 U12378 ( .IN1(n12362), .IN2(n12363), .Q(n12361) );
  AND2X1 U12379 ( .IN1(g2412), .IN2(g2443), .Q(n12363) );
  AND2X1 U12380 ( .IN1(g5747), .IN2(g2439), .Q(n12362) );
  AND2X1 U12381 ( .IN1(g5796), .IN2(g2441), .Q(n12360) );
  AND2X1 U12382 ( .IN1(n12292), .IN2(n12289), .Q(n12355) );
  INVX0 U12383 ( .INP(n12316), .ZN(n12292) );
  OR2X1 U12384 ( .IN1(n12364), .IN2(n12365), .Q(n12316) );
  OR2X1 U12385 ( .IN1(n12366), .IN2(n12367), .Q(n12365) );
  AND2X1 U12386 ( .IN1(g2412), .IN2(g2458), .Q(n12367) );
  AND2X1 U12387 ( .IN1(g5747), .IN2(g2454), .Q(n12366) );
  AND2X1 U12388 ( .IN1(g5796), .IN2(g2456), .Q(n12364) );
  INVX0 U12389 ( .INP(n12287), .ZN(n12296) );
  OR2X1 U12390 ( .IN1(n12368), .IN2(n12369), .Q(n12287) );
  OR2X1 U12391 ( .IN1(n12370), .IN2(n12371), .Q(n12369) );
  AND2X1 U12392 ( .IN1(g2412), .IN2(g2428), .Q(n12371) );
  AND2X1 U12393 ( .IN1(g5747), .IN2(g2424), .Q(n12370) );
  AND2X1 U12394 ( .IN1(g5796), .IN2(g2426), .Q(n12368) );
  AND2X1 U12395 ( .IN1(n12372), .IN2(n12321), .Q(n12352) );
  INVX0 U12396 ( .INP(n12303), .ZN(n12321) );
  OR2X1 U12397 ( .IN1(n12373), .IN2(n12374), .Q(n12303) );
  OR2X1 U12398 ( .IN1(n12375), .IN2(n12376), .Q(n12374) );
  AND2X1 U12399 ( .IN1(test_so85), .IN2(g2412), .Q(n12376) );
  AND2X1 U12400 ( .IN1(g5747), .IN2(g2469), .Q(n12375) );
  AND2X1 U12401 ( .IN1(g5796), .IN2(g2471), .Q(n12373) );
  AND2X1 U12402 ( .IN1(n12307), .IN2(n12294), .Q(n12372) );
  AND2X1 U12403 ( .IN1(n10225), .IN2(n12332), .Q(n10222) );
  OR2X1 U12404 ( .IN1(n12377), .IN2(n12378), .Q(g28357) );
  AND2X1 U12405 ( .IN1(n12260), .IN2(n12379), .Q(n12378) );
  OR2X1 U12406 ( .IN1(n12380), .IN2(n12381), .Q(n12260) );
  AND2X1 U12407 ( .IN1(n10023), .IN2(n12265), .Q(n12381) );
  AND2X1 U12408 ( .IN1(n3293), .IN2(n12382), .Q(n12380) );
  INVX0 U12409 ( .INP(n12383), .ZN(n12382) );
  AND2X1 U12410 ( .IN1(n12266), .IN2(n12384), .Q(n3293) );
  INVX0 U12411 ( .INP(n12385), .ZN(n12384) );
  OR2X1 U12412 ( .IN1(n12386), .IN2(n12387), .Q(n12385) );
  INVX0 U12413 ( .INP(n12388), .ZN(n12387) );
  OR2X1 U12414 ( .IN1(n12389), .IN2(n12390), .Q(n12388) );
  AND2X1 U12415 ( .IN1(n4296), .IN2(g1994), .Q(n12377) );
  OR2X1 U12416 ( .IN1(n12391), .IN2(n12392), .Q(g28356) );
  AND2X1 U12417 ( .IN1(n12273), .IN2(g7194), .Q(n12392) );
  AND2X1 U12418 ( .IN1(n4315), .IN2(g1988), .Q(n12391) );
  OR2X1 U12419 ( .IN1(n12393), .IN2(n12394), .Q(g28355) );
  AND2X1 U12420 ( .IN1(n12276), .IN2(g6944), .Q(n12394) );
  AND2X1 U12421 ( .IN1(n4316), .IN2(g1303), .Q(n12393) );
  OR2X1 U12422 ( .IN1(n12395), .IN2(n12396), .Q(g28354) );
  AND2X1 U12423 ( .IN1(n12397), .IN2(g1236), .Q(n12396) );
  AND2X1 U12424 ( .IN1(n4300), .IN2(g1297), .Q(n12395) );
  OR2X1 U12425 ( .IN1(n12398), .IN2(n12399), .Q(g28353) );
  AND2X1 U12426 ( .IN1(n12400), .IN2(g550), .Q(n12399) );
  AND2X1 U12427 ( .IN1(n4313), .IN2(test_so26), .Q(n12398) );
  OR2X1 U12428 ( .IN1(n12401), .IN2(n12402), .Q(g28352) );
  AND2X1 U12429 ( .IN1(n4296), .IN2(g1985), .Q(n12402) );
  AND2X1 U12430 ( .IN1(g7052), .IN2(n12273), .Q(n12401) );
  OR2X1 U12431 ( .IN1(n12403), .IN2(n12404), .Q(n12273) );
  AND2X1 U12432 ( .IN1(n10013), .IN2(n12265), .Q(n12404) );
  AND2X1 U12433 ( .IN1(n3301), .IN2(n12405), .Q(n12403) );
  INVX0 U12434 ( .INP(n12390), .ZN(n12405) );
  OR2X1 U12435 ( .IN1(n12406), .IN2(n12407), .Q(n12390) );
  OR2X1 U12436 ( .IN1(n12408), .IN2(n12409), .Q(n12407) );
  AND2X1 U12437 ( .IN1(n12410), .IN2(n12411), .Q(n12409) );
  AND2X1 U12438 ( .IN1(n12412), .IN2(n12413), .Q(n12410) );
  OR2X1 U12439 ( .IN1(n12414), .IN2(n12415), .Q(n12412) );
  AND2X1 U12440 ( .IN1(n12416), .IN2(n12417), .Q(n12414) );
  OR2X1 U12441 ( .IN1(n12418), .IN2(n12419), .Q(n12417) );
  AND2X1 U12442 ( .IN1(n12420), .IN2(n12421), .Q(n12408) );
  OR2X1 U12443 ( .IN1(n12422), .IN2(n12423), .Q(n12421) );
  AND2X1 U12444 ( .IN1(n12424), .IN2(n12425), .Q(n12423) );
  OR2X1 U12445 ( .IN1(n12426), .IN2(n12416), .Q(n12424) );
  AND2X1 U12446 ( .IN1(n12427), .IN2(n12428), .Q(n12426) );
  AND2X1 U12447 ( .IN1(n12429), .IN2(n12430), .Q(n12422) );
  AND2X1 U12448 ( .IN1(n12418), .IN2(n12419), .Q(n12430) );
  AND2X1 U12449 ( .IN1(n12416), .IN2(n12431), .Q(n12429) );
  OR2X1 U12450 ( .IN1(n12432), .IN2(n12433), .Q(n12406) );
  AND2X1 U12451 ( .IN1(n12434), .IN2(n12428), .Q(n12433) );
  AND2X1 U12452 ( .IN1(n12435), .IN2(n12436), .Q(n12434) );
  OR2X1 U12453 ( .IN1(n12437), .IN2(n12438), .Q(n12436) );
  AND2X1 U12454 ( .IN1(n12439), .IN2(n12440), .Q(n12437) );
  AND2X1 U12455 ( .IN1(n12441), .IN2(n12442), .Q(n12432) );
  OR2X1 U12456 ( .IN1(n12443), .IN2(n12444), .Q(n12442) );
  AND2X1 U12457 ( .IN1(n12445), .IN2(n12439), .Q(n12444) );
  OR2X1 U12458 ( .IN1(n12446), .IN2(n12447), .Q(n12439) );
  AND2X1 U12459 ( .IN1(n12448), .IN2(n12411), .Q(n12446) );
  AND2X1 U12460 ( .IN1(n12449), .IN2(n12438), .Q(n12443) );
  OR2X1 U12461 ( .IN1(n12450), .IN2(n12451), .Q(n12438) );
  AND2X1 U12462 ( .IN1(n12447), .IN2(n12411), .Q(n12451) );
  AND2X1 U12463 ( .IN1(n12431), .IN2(n12420), .Q(n12450) );
  AND2X1 U12464 ( .IN1(n12266), .IN2(n12452), .Q(n3301) );
  INVX0 U12465 ( .INP(n12453), .ZN(n12452) );
  OR2X1 U12466 ( .IN1(n12386), .IN2(n12454), .Q(n12453) );
  INVX0 U12467 ( .INP(n12455), .ZN(n12454) );
  OR2X1 U12468 ( .IN1(n12456), .IN2(n12383), .Q(n12455) );
  OR2X1 U12469 ( .IN1(n12457), .IN2(n12458), .Q(n12383) );
  OR2X1 U12470 ( .IN1(n12459), .IN2(n12460), .Q(n12458) );
  AND2X1 U12471 ( .IN1(n12461), .IN2(n12411), .Q(n12460) );
  OR2X1 U12472 ( .IN1(n12462), .IN2(n12463), .Q(n12461) );
  AND2X1 U12473 ( .IN1(n12441), .IN2(n12464), .Q(n12463) );
  OR2X1 U12474 ( .IN1(n12465), .IN2(n12466), .Q(n12464) );
  OR2X1 U12475 ( .IN1(n12467), .IN2(n12468), .Q(n12466) );
  AND2X1 U12476 ( .IN1(n12415), .IN2(n12431), .Q(n12468) );
  AND2X1 U12477 ( .IN1(n12418), .IN2(n12469), .Q(n12415) );
  AND2X1 U12478 ( .IN1(n12419), .IN2(n12427), .Q(n12469) );
  AND2X1 U12479 ( .IN1(n12470), .IN2(n12416), .Q(n12467) );
  AND2X1 U12480 ( .IN1(n12435), .IN2(n12447), .Q(n12465) );
  AND2X1 U12481 ( .IN1(n12449), .IN2(n12425), .Q(n12462) );
  AND2X1 U12482 ( .IN1(n12471), .IN2(n12435), .Q(n12459) );
  INVX0 U12483 ( .INP(n12419), .ZN(n12435) );
  AND2X1 U12484 ( .IN1(n12472), .IN2(n12413), .Q(n12471) );
  OR2X1 U12485 ( .IN1(n12473), .IN2(n12474), .Q(n12472) );
  AND2X1 U12486 ( .IN1(n12441), .IN2(n12440), .Q(n12474) );
  AND2X1 U12487 ( .IN1(n12420), .IN2(n12418), .Q(n12473) );
  AND2X1 U12488 ( .IN1(n12475), .IN2(n12428), .Q(n12457) );
  OR2X1 U12489 ( .IN1(n12476), .IN2(n12477), .Q(n12475) );
  AND2X1 U12490 ( .IN1(n12420), .IN2(n12478), .Q(n12477) );
  OR2X1 U12491 ( .IN1(n12479), .IN2(n12480), .Q(n12478) );
  OR2X1 U12492 ( .IN1(n12481), .IN2(n12482), .Q(n12480) );
  AND2X1 U12493 ( .IN1(n12470), .IN2(n12449), .Q(n12482) );
  AND2X1 U12494 ( .IN1(n12419), .IN2(n12440), .Q(n12449) );
  AND2X1 U12495 ( .IN1(n12483), .IN2(n12427), .Q(n12481) );
  AND2X1 U12496 ( .IN1(n12447), .IN2(n12419), .Q(n12483) );
  OR2X1 U12497 ( .IN1(n12484), .IN2(n12485), .Q(n12419) );
  OR2X1 U12498 ( .IN1(n12486), .IN2(n12487), .Q(n12485) );
  AND2X1 U12499 ( .IN1(g5738), .IN2(g1747), .Q(n12487) );
  AND2X1 U12500 ( .IN1(g1718), .IN2(g1749), .Q(n12486) );
  AND2X1 U12501 ( .IN1(test_so63), .IN2(g1745), .Q(n12484) );
  AND2X1 U12502 ( .IN1(n12416), .IN2(n12413), .Q(n12479) );
  INVX0 U12503 ( .INP(n12440), .ZN(n12416) );
  OR2X1 U12504 ( .IN1(n12488), .IN2(n12489), .Q(n12440) );
  OR2X1 U12505 ( .IN1(n12490), .IN2(n12491), .Q(n12489) );
  AND2X1 U12506 ( .IN1(g5738), .IN2(g1762), .Q(n12491) );
  AND2X1 U12507 ( .IN1(g1718), .IN2(g1764), .Q(n12490) );
  AND2X1 U12508 ( .IN1(test_so63), .IN2(g1760), .Q(n12488) );
  INVX0 U12509 ( .INP(n12411), .ZN(n12420) );
  OR2X1 U12510 ( .IN1(n12492), .IN2(n12493), .Q(n12411) );
  OR2X1 U12511 ( .IN1(n12494), .IN2(n12495), .Q(n12493) );
  AND2X1 U12512 ( .IN1(g5738), .IN2(g1732), .Q(n12495) );
  AND2X1 U12513 ( .IN1(g1718), .IN2(g1734), .Q(n12494) );
  AND2X1 U12514 ( .IN1(test_so63), .IN2(g1730), .Q(n12492) );
  AND2X1 U12515 ( .IN1(n12496), .IN2(n12445), .Q(n12476) );
  INVX0 U12516 ( .INP(n12427), .ZN(n12445) );
  OR2X1 U12517 ( .IN1(n12497), .IN2(n12498), .Q(n12427) );
  OR2X1 U12518 ( .IN1(n12499), .IN2(n12500), .Q(n12498) );
  AND2X1 U12519 ( .IN1(g5738), .IN2(g1777), .Q(n12500) );
  AND2X1 U12520 ( .IN1(g1718), .IN2(g1705), .Q(n12499) );
  AND2X1 U12521 ( .IN1(test_so63), .IN2(g1775), .Q(n12497) );
  AND2X1 U12522 ( .IN1(n12431), .IN2(n12418), .Q(n12496) );
  AND2X1 U12523 ( .IN1(n12389), .IN2(n12456), .Q(n12386) );
  OR2X1 U12524 ( .IN1(n12501), .IN2(n12502), .Q(g28351) );
  AND2X1 U12525 ( .IN1(n12276), .IN2(n12249), .Q(n12502) );
  OR2X1 U12526 ( .IN1(n12503), .IN2(n12504), .Q(n12276) );
  AND2X1 U12527 ( .IN1(n10158), .IN2(n12265), .Q(n12504) );
  AND2X1 U12528 ( .IN1(n3334), .IN2(n12505), .Q(n12503) );
  INVX0 U12529 ( .INP(n12506), .ZN(n12505) );
  AND2X1 U12530 ( .IN1(n12266), .IN2(n12507), .Q(n3334) );
  INVX0 U12531 ( .INP(n12508), .ZN(n12507) );
  OR2X1 U12532 ( .IN1(n12509), .IN2(n12510), .Q(n12508) );
  INVX0 U12533 ( .INP(n12511), .ZN(n12510) );
  OR2X1 U12534 ( .IN1(n12512), .IN2(n12513), .Q(n12511) );
  AND2X1 U12535 ( .IN1(n4371), .IN2(g1300), .Q(n12501) );
  OR2X1 U12536 ( .IN1(n12514), .IN2(n12515), .Q(g28350) );
  AND2X1 U12537 ( .IN1(n12397), .IN2(g6944), .Q(n12515) );
  AND2X1 U12538 ( .IN1(n4316), .IN2(g1294), .Q(n12514) );
  OR2X1 U12539 ( .IN1(n12516), .IN2(n12517), .Q(g28349) );
  AND2X1 U12540 ( .IN1(n12400), .IN2(g6642), .Q(n12517) );
  AND2X1 U12541 ( .IN1(n4372), .IN2(g617), .Q(n12516) );
  OR2X1 U12542 ( .IN1(n12518), .IN2(n12519), .Q(g28348) );
  AND2X1 U12543 ( .IN1(n12520), .IN2(g550), .Q(n12519) );
  AND2X1 U12544 ( .IN1(n4313), .IN2(g611), .Q(n12518) );
  OR2X1 U12545 ( .IN1(n12521), .IN2(n12522), .Q(g28346) );
  AND2X1 U12546 ( .IN1(n4371), .IN2(g1291), .Q(n12522) );
  AND2X1 U12547 ( .IN1(g6750), .IN2(n12397), .Q(n12521) );
  OR2X1 U12548 ( .IN1(n12523), .IN2(n12524), .Q(n12397) );
  AND2X1 U12549 ( .IN1(n10148), .IN2(n12265), .Q(n12524) );
  AND2X1 U12550 ( .IN1(n3341), .IN2(n12525), .Q(n12523) );
  INVX0 U12551 ( .INP(n12513), .ZN(n12525) );
  OR2X1 U12552 ( .IN1(n12526), .IN2(n12527), .Q(n12513) );
  OR2X1 U12553 ( .IN1(n12528), .IN2(n12529), .Q(n12527) );
  AND2X1 U12554 ( .IN1(n12530), .IN2(n12531), .Q(n12529) );
  AND2X1 U12555 ( .IN1(n12532), .IN2(n12533), .Q(n12530) );
  OR2X1 U12556 ( .IN1(n12534), .IN2(n12535), .Q(n12532) );
  AND2X1 U12557 ( .IN1(n12536), .IN2(n12537), .Q(n12534) );
  OR2X1 U12558 ( .IN1(n12538), .IN2(n12539), .Q(n12537) );
  AND2X1 U12559 ( .IN1(n12540), .IN2(n12541), .Q(n12528) );
  OR2X1 U12560 ( .IN1(n12542), .IN2(n12543), .Q(n12541) );
  AND2X1 U12561 ( .IN1(n12544), .IN2(n12545), .Q(n12543) );
  OR2X1 U12562 ( .IN1(n12546), .IN2(n12536), .Q(n12544) );
  AND2X1 U12563 ( .IN1(n12547), .IN2(n12548), .Q(n12546) );
  AND2X1 U12564 ( .IN1(n12549), .IN2(n12550), .Q(n12542) );
  AND2X1 U12565 ( .IN1(n12538), .IN2(n12539), .Q(n12550) );
  AND2X1 U12566 ( .IN1(n12536), .IN2(n12551), .Q(n12549) );
  OR2X1 U12567 ( .IN1(n12552), .IN2(n12553), .Q(n12526) );
  AND2X1 U12568 ( .IN1(n12554), .IN2(n12548), .Q(n12553) );
  AND2X1 U12569 ( .IN1(n12555), .IN2(n12556), .Q(n12554) );
  OR2X1 U12570 ( .IN1(n12557), .IN2(n12558), .Q(n12556) );
  AND2X1 U12571 ( .IN1(n12559), .IN2(n12560), .Q(n12557) );
  AND2X1 U12572 ( .IN1(n12561), .IN2(n12562), .Q(n12552) );
  OR2X1 U12573 ( .IN1(n12563), .IN2(n12564), .Q(n12562) );
  AND2X1 U12574 ( .IN1(n12565), .IN2(n12559), .Q(n12564) );
  OR2X1 U12575 ( .IN1(n12566), .IN2(n12567), .Q(n12559) );
  AND2X1 U12576 ( .IN1(n12568), .IN2(n12531), .Q(n12566) );
  AND2X1 U12577 ( .IN1(n12569), .IN2(n12558), .Q(n12563) );
  OR2X1 U12578 ( .IN1(n12570), .IN2(n12571), .Q(n12558) );
  AND2X1 U12579 ( .IN1(n12567), .IN2(n12531), .Q(n12571) );
  AND2X1 U12580 ( .IN1(n12551), .IN2(n12540), .Q(n12570) );
  AND2X1 U12581 ( .IN1(n12266), .IN2(n12572), .Q(n3341) );
  INVX0 U12582 ( .INP(n12573), .ZN(n12572) );
  OR2X1 U12583 ( .IN1(n12509), .IN2(n12574), .Q(n12573) );
  INVX0 U12584 ( .INP(n12575), .ZN(n12574) );
  OR2X1 U12585 ( .IN1(n12576), .IN2(n12506), .Q(n12575) );
  OR2X1 U12586 ( .IN1(n12577), .IN2(n12578), .Q(n12506) );
  OR2X1 U12587 ( .IN1(n12579), .IN2(n12580), .Q(n12578) );
  AND2X1 U12588 ( .IN1(n12581), .IN2(n12531), .Q(n12580) );
  OR2X1 U12589 ( .IN1(n12582), .IN2(n12583), .Q(n12581) );
  AND2X1 U12590 ( .IN1(n12561), .IN2(n12584), .Q(n12583) );
  OR2X1 U12591 ( .IN1(n12585), .IN2(n12586), .Q(n12584) );
  OR2X1 U12592 ( .IN1(n12587), .IN2(n12588), .Q(n12586) );
  AND2X1 U12593 ( .IN1(n12535), .IN2(n12551), .Q(n12588) );
  AND2X1 U12594 ( .IN1(n12538), .IN2(n12589), .Q(n12535) );
  AND2X1 U12595 ( .IN1(n12539), .IN2(n12547), .Q(n12589) );
  AND2X1 U12596 ( .IN1(n12590), .IN2(n12536), .Q(n12587) );
  AND2X1 U12597 ( .IN1(n12555), .IN2(n12567), .Q(n12585) );
  AND2X1 U12598 ( .IN1(n12569), .IN2(n12545), .Q(n12582) );
  AND2X1 U12599 ( .IN1(n12591), .IN2(n12555), .Q(n12579) );
  INVX0 U12600 ( .INP(n12539), .ZN(n12555) );
  AND2X1 U12601 ( .IN1(n12592), .IN2(n12533), .Q(n12591) );
  OR2X1 U12602 ( .IN1(n12593), .IN2(n12594), .Q(n12592) );
  AND2X1 U12603 ( .IN1(n12561), .IN2(n12560), .Q(n12594) );
  AND2X1 U12604 ( .IN1(n12540), .IN2(n12538), .Q(n12593) );
  AND2X1 U12605 ( .IN1(n12595), .IN2(n12548), .Q(n12577) );
  OR2X1 U12606 ( .IN1(n12596), .IN2(n12597), .Q(n12595) );
  AND2X1 U12607 ( .IN1(n12540), .IN2(n12598), .Q(n12597) );
  OR2X1 U12608 ( .IN1(n12599), .IN2(n12600), .Q(n12598) );
  OR2X1 U12609 ( .IN1(n12601), .IN2(n12602), .Q(n12600) );
  AND2X1 U12610 ( .IN1(n12590), .IN2(n12569), .Q(n12602) );
  AND2X1 U12611 ( .IN1(n12539), .IN2(n12560), .Q(n12569) );
  AND2X1 U12612 ( .IN1(n12603), .IN2(n12547), .Q(n12601) );
  AND2X1 U12613 ( .IN1(n12567), .IN2(n12539), .Q(n12603) );
  OR2X1 U12614 ( .IN1(n12604), .IN2(n12605), .Q(n12539) );
  OR2X1 U12615 ( .IN1(n12606), .IN2(n12607), .Q(n12605) );
  AND2X1 U12616 ( .IN1(g1024), .IN2(g1055), .Q(n12607) );
  AND2X1 U12617 ( .IN1(g5657), .IN2(g1051), .Q(n12606) );
  AND2X1 U12618 ( .IN1(g5686), .IN2(g1053), .Q(n12604) );
  AND2X1 U12619 ( .IN1(n12536), .IN2(n12533), .Q(n12599) );
  INVX0 U12620 ( .INP(n12560), .ZN(n12536) );
  OR2X1 U12621 ( .IN1(n12608), .IN2(n12609), .Q(n12560) );
  OR2X1 U12622 ( .IN1(n12610), .IN2(n12611), .Q(n12609) );
  AND2X1 U12623 ( .IN1(g1024), .IN2(g1070), .Q(n12611) );
  AND2X1 U12624 ( .IN1(g5657), .IN2(g1066), .Q(n12610) );
  AND2X1 U12625 ( .IN1(g5686), .IN2(g1068), .Q(n12608) );
  INVX0 U12626 ( .INP(n12531), .ZN(n12540) );
  OR2X1 U12627 ( .IN1(n12612), .IN2(n12613), .Q(n12531) );
  OR2X1 U12628 ( .IN1(n12614), .IN2(n12615), .Q(n12613) );
  AND2X1 U12629 ( .IN1(g1024), .IN2(g1040), .Q(n12615) );
  AND2X1 U12630 ( .IN1(g5657), .IN2(g1036), .Q(n12614) );
  AND2X1 U12631 ( .IN1(g5686), .IN2(g1038), .Q(n12612) );
  AND2X1 U12632 ( .IN1(n12616), .IN2(n12565), .Q(n12596) );
  INVX0 U12633 ( .INP(n12547), .ZN(n12565) );
  OR2X1 U12634 ( .IN1(n12617), .IN2(n12618), .Q(n12547) );
  OR2X1 U12635 ( .IN1(n12619), .IN2(n12620), .Q(n12618) );
  AND2X1 U12636 ( .IN1(g1024), .IN2(g1011), .Q(n12620) );
  AND2X1 U12637 ( .IN1(g5657), .IN2(g1081), .Q(n12619) );
  AND2X1 U12638 ( .IN1(g5686), .IN2(g1083), .Q(n12617) );
  AND2X1 U12639 ( .IN1(n12551), .IN2(n12538), .Q(n12616) );
  AND2X1 U12640 ( .IN1(n12512), .IN2(n12576), .Q(n12509) );
  OR2X1 U12641 ( .IN1(n12621), .IN2(n12622), .Q(g28345) );
  AND2X1 U12642 ( .IN1(n12400), .IN2(n9810), .Q(n12622) );
  OR2X1 U12643 ( .IN1(n12623), .IN2(n12624), .Q(n12400) );
  AND2X1 U12644 ( .IN1(n9738), .IN2(n12265), .Q(n12624) );
  AND2X1 U12645 ( .IN1(n3374), .IN2(n12625), .Q(n12623) );
  INVX0 U12646 ( .INP(n12626), .ZN(n12625) );
  AND2X1 U12647 ( .IN1(n12266), .IN2(n12627), .Q(n3374) );
  INVX0 U12648 ( .INP(n12628), .ZN(n12627) );
  OR2X1 U12649 ( .IN1(n12629), .IN2(n12630), .Q(n12628) );
  INVX0 U12650 ( .INP(n12631), .ZN(n12630) );
  OR2X1 U12651 ( .IN1(n12632), .IN2(n12633), .Q(n12631) );
  AND2X1 U12652 ( .IN1(n4298), .IN2(g614), .Q(n12621) );
  OR2X1 U12653 ( .IN1(n12634), .IN2(n12635), .Q(g28344) );
  AND2X1 U12654 ( .IN1(n12520), .IN2(g6642), .Q(n12635) );
  AND2X1 U12655 ( .IN1(n4372), .IN2(g608), .Q(n12634) );
  OR2X1 U12656 ( .IN1(n12636), .IN2(n12637), .Q(g28342) );
  AND2X1 U12657 ( .IN1(n4298), .IN2(g605), .Q(n12637) );
  AND2X1 U12658 ( .IN1(g6485), .IN2(n12520), .Q(n12636) );
  OR2X1 U12659 ( .IN1(n12638), .IN2(n12639), .Q(n12520) );
  AND2X1 U12660 ( .IN1(n9744), .IN2(n12265), .Q(n12639) );
  AND2X1 U12661 ( .IN1(n3380), .IN2(n12640), .Q(n12638) );
  INVX0 U12662 ( .INP(n12633), .ZN(n12640) );
  OR2X1 U12663 ( .IN1(n12641), .IN2(n12642), .Q(n12633) );
  OR2X1 U12664 ( .IN1(n12643), .IN2(n12644), .Q(n12642) );
  AND2X1 U12665 ( .IN1(n12645), .IN2(n12646), .Q(n12644) );
  AND2X1 U12666 ( .IN1(n12647), .IN2(n12648), .Q(n12645) );
  OR2X1 U12667 ( .IN1(n12649), .IN2(n12650), .Q(n12647) );
  AND2X1 U12668 ( .IN1(n12651), .IN2(n12652), .Q(n12649) );
  OR2X1 U12669 ( .IN1(n12653), .IN2(n12654), .Q(n12652) );
  AND2X1 U12670 ( .IN1(n12655), .IN2(n12656), .Q(n12643) );
  OR2X1 U12671 ( .IN1(n12657), .IN2(n12658), .Q(n12656) );
  AND2X1 U12672 ( .IN1(n12659), .IN2(n12660), .Q(n12658) );
  OR2X1 U12673 ( .IN1(n12661), .IN2(n12651), .Q(n12659) );
  AND2X1 U12674 ( .IN1(n12662), .IN2(n12663), .Q(n12661) );
  AND2X1 U12675 ( .IN1(n12664), .IN2(n12665), .Q(n12657) );
  AND2X1 U12676 ( .IN1(n12653), .IN2(n12654), .Q(n12665) );
  AND2X1 U12677 ( .IN1(n12651), .IN2(n12666), .Q(n12664) );
  OR2X1 U12678 ( .IN1(n12667), .IN2(n12668), .Q(n12641) );
  AND2X1 U12679 ( .IN1(n12669), .IN2(n12663), .Q(n12668) );
  AND2X1 U12680 ( .IN1(n12670), .IN2(n12671), .Q(n12669) );
  OR2X1 U12681 ( .IN1(n12672), .IN2(n12673), .Q(n12671) );
  AND2X1 U12682 ( .IN1(n12674), .IN2(n12675), .Q(n12672) );
  AND2X1 U12683 ( .IN1(n12676), .IN2(n12677), .Q(n12667) );
  OR2X1 U12684 ( .IN1(n12678), .IN2(n12679), .Q(n12677) );
  AND2X1 U12685 ( .IN1(n12680), .IN2(n12674), .Q(n12679) );
  OR2X1 U12686 ( .IN1(n12681), .IN2(n12682), .Q(n12674) );
  AND2X1 U12687 ( .IN1(n12683), .IN2(n12646), .Q(n12681) );
  AND2X1 U12688 ( .IN1(n12684), .IN2(n12673), .Q(n12678) );
  OR2X1 U12689 ( .IN1(n12685), .IN2(n12686), .Q(n12673) );
  AND2X1 U12690 ( .IN1(n12682), .IN2(n12646), .Q(n12686) );
  AND2X1 U12691 ( .IN1(n12666), .IN2(n12655), .Q(n12685) );
  AND2X1 U12692 ( .IN1(n12266), .IN2(n12687), .Q(n3380) );
  INVX0 U12693 ( .INP(n12688), .ZN(n12687) );
  OR2X1 U12694 ( .IN1(n12629), .IN2(n12689), .Q(n12688) );
  INVX0 U12695 ( .INP(n12690), .ZN(n12689) );
  OR2X1 U12696 ( .IN1(n12691), .IN2(n12626), .Q(n12690) );
  OR2X1 U12697 ( .IN1(n12692), .IN2(n12693), .Q(n12626) );
  OR2X1 U12698 ( .IN1(n12694), .IN2(n12695), .Q(n12693) );
  AND2X1 U12699 ( .IN1(n12696), .IN2(n12646), .Q(n12695) );
  OR2X1 U12700 ( .IN1(n12697), .IN2(n12698), .Q(n12696) );
  AND2X1 U12701 ( .IN1(n12676), .IN2(n12699), .Q(n12698) );
  OR2X1 U12702 ( .IN1(n12700), .IN2(n12701), .Q(n12699) );
  OR2X1 U12703 ( .IN1(n12702), .IN2(n12703), .Q(n12701) );
  AND2X1 U12704 ( .IN1(n12650), .IN2(n12666), .Q(n12703) );
  AND2X1 U12705 ( .IN1(n12653), .IN2(n12704), .Q(n12650) );
  AND2X1 U12706 ( .IN1(n12654), .IN2(n12662), .Q(n12704) );
  AND2X1 U12707 ( .IN1(n12705), .IN2(n12651), .Q(n12702) );
  AND2X1 U12708 ( .IN1(n12670), .IN2(n12682), .Q(n12700) );
  AND2X1 U12709 ( .IN1(n12684), .IN2(n12660), .Q(n12697) );
  AND2X1 U12710 ( .IN1(n12706), .IN2(n12670), .Q(n12694) );
  INVX0 U12711 ( .INP(n12654), .ZN(n12670) );
  AND2X1 U12712 ( .IN1(n12707), .IN2(n12648), .Q(n12706) );
  OR2X1 U12713 ( .IN1(n12708), .IN2(n12709), .Q(n12707) );
  AND2X1 U12714 ( .IN1(n12676), .IN2(n12675), .Q(n12709) );
  AND2X1 U12715 ( .IN1(n12655), .IN2(n12653), .Q(n12708) );
  AND2X1 U12716 ( .IN1(n12710), .IN2(n12663), .Q(n12692) );
  OR2X1 U12717 ( .IN1(n12711), .IN2(n12712), .Q(n12710) );
  AND2X1 U12718 ( .IN1(n12655), .IN2(n12713), .Q(n12712) );
  OR2X1 U12719 ( .IN1(n12714), .IN2(n12715), .Q(n12713) );
  OR2X1 U12720 ( .IN1(n12716), .IN2(n12717), .Q(n12715) );
  AND2X1 U12721 ( .IN1(n12705), .IN2(n12684), .Q(n12717) );
  AND2X1 U12722 ( .IN1(n12654), .IN2(n12675), .Q(n12684) );
  AND2X1 U12723 ( .IN1(n12718), .IN2(n12662), .Q(n12716) );
  AND2X1 U12724 ( .IN1(n12682), .IN2(n12654), .Q(n12718) );
  OR2X1 U12725 ( .IN1(n12719), .IN2(n12720), .Q(n12654) );
  OR2X1 U12726 ( .IN1(n12721), .IN2(n12722), .Q(n12720) );
  AND2X1 U12727 ( .IN1(g337), .IN2(g368), .Q(n12722) );
  AND2X1 U12728 ( .IN1(g5629), .IN2(g364), .Q(n12721) );
  AND2X1 U12729 ( .IN1(g5648), .IN2(g366), .Q(n12719) );
  AND2X1 U12730 ( .IN1(n12651), .IN2(n12648), .Q(n12714) );
  INVX0 U12731 ( .INP(n12675), .ZN(n12651) );
  OR2X1 U12732 ( .IN1(n12723), .IN2(n12724), .Q(n12675) );
  OR2X1 U12733 ( .IN1(n12725), .IN2(n12726), .Q(n12724) );
  AND2X1 U12734 ( .IN1(g337), .IN2(g383), .Q(n12726) );
  AND2X1 U12735 ( .IN1(g5629), .IN2(g379), .Q(n12725) );
  AND2X1 U12736 ( .IN1(g5648), .IN2(g381), .Q(n12723) );
  INVX0 U12737 ( .INP(n12646), .ZN(n12655) );
  OR2X1 U12738 ( .IN1(n12727), .IN2(n12728), .Q(n12646) );
  OR2X1 U12739 ( .IN1(n12729), .IN2(n12730), .Q(n12728) );
  AND2X1 U12740 ( .IN1(g337), .IN2(g353), .Q(n12730) );
  AND2X1 U12741 ( .IN1(g5629), .IN2(g349), .Q(n12729) );
  AND2X1 U12742 ( .IN1(g5648), .IN2(g351), .Q(n12727) );
  AND2X1 U12743 ( .IN1(n12731), .IN2(n12680), .Q(n12711) );
  INVX0 U12744 ( .INP(n12662), .ZN(n12680) );
  OR2X1 U12745 ( .IN1(n12732), .IN2(n12733), .Q(n12662) );
  OR2X1 U12746 ( .IN1(n12734), .IN2(n12735), .Q(n12733) );
  AND2X1 U12747 ( .IN1(g337), .IN2(g324), .Q(n12735) );
  AND2X1 U12748 ( .IN1(g5629), .IN2(g394), .Q(n12734) );
  AND2X1 U12749 ( .IN1(g5648), .IN2(g396), .Q(n12732) );
  AND2X1 U12750 ( .IN1(n12666), .IN2(n12653), .Q(n12731) );
  AND2X1 U12751 ( .IN1(n12632), .IN2(n12691), .Q(n12629) );
  INVX0 U12752 ( .INP(n12265), .ZN(n12266) );
  AND2X1 U12753 ( .IN1(n12736), .IN2(n12737), .Q(g28328) );
  XOR2X1 U12754 ( .IN1(n12738), .IN2(n4415), .Q(n12736) );
  OR2X1 U12755 ( .IN1(n4393), .IN2(n12739), .Q(n12738) );
  AND2X1 U12756 ( .IN1(n12740), .IN2(n12741), .Q(g28325) );
  XOR2X1 U12757 ( .IN1(n12742), .IN2(n4416), .Q(n12740) );
  OR2X1 U12758 ( .IN1(n12743), .IN2(n9124), .Q(n12742) );
  AND2X1 U12759 ( .IN1(n12744), .IN2(n12745), .Q(g28321) );
  XOR2X1 U12760 ( .IN1(n12746), .IN2(n4417), .Q(n12744) );
  OR2X1 U12761 ( .IN1(n4395), .IN2(n12747), .Q(n12746) );
  AND2X1 U12762 ( .IN1(n12748), .IN2(n12226), .Q(g28199) );
  XOR2X1 U12763 ( .IN1(n12228), .IN2(n4396), .Q(n12748) );
  AND2X1 U12764 ( .IN1(n12749), .IN2(n12750), .Q(g28148) );
  OR2X1 U12765 ( .IN1(n3424), .IN2(g2138), .Q(n12750) );
  AND2X1 U12766 ( .IN1(n11527), .IN2(n1289), .Q(n12749) );
  INVX0 U12767 ( .INP(n12230), .ZN(n1289) );
  AND2X1 U12768 ( .IN1(g2138), .IN2(n3424), .Q(n12230) );
  AND2X1 U12769 ( .IN1(n12751), .IN2(n12752), .Q(g28147) );
  OR2X1 U12770 ( .IN1(n3427), .IN2(g1444), .Q(n12752) );
  AND2X1 U12771 ( .IN1(n11529), .IN2(n1003), .Q(n12751) );
  INVX0 U12772 ( .INP(n12232), .ZN(n1003) );
  AND2X1 U12773 ( .IN1(g1444), .IN2(n3427), .Q(n12232) );
  AND2X1 U12774 ( .IN1(n12753), .IN2(n12754), .Q(g28146) );
  OR2X1 U12775 ( .IN1(n3430), .IN2(g758), .Q(n12754) );
  AND2X1 U12776 ( .IN1(n11531), .IN2(n714), .Q(n12753) );
  INVX0 U12777 ( .INP(n12234), .ZN(n714) );
  AND2X1 U12778 ( .IN1(g758), .IN2(n3430), .Q(n12234) );
  AND2X1 U12779 ( .IN1(n12755), .IN2(n12756), .Q(g28145) );
  OR2X1 U12780 ( .IN1(n3433), .IN2(g70), .Q(n12756) );
  AND2X1 U12781 ( .IN1(n11533), .IN2(n405), .Q(n12755) );
  INVX0 U12782 ( .INP(n12236), .ZN(n405) );
  AND2X1 U12783 ( .IN1(g70), .IN2(n3433), .Q(n12236) );
  OR2X1 U12784 ( .IN1(n12757), .IN2(n12758), .Q(g27771) );
  AND2X1 U12785 ( .IN1(n12759), .IN2(n10833), .Q(n12758) );
  AND2X1 U12786 ( .IN1(test_so81), .IN2(n12760), .Q(n12757) );
  OR2X1 U12787 ( .IN1(n4509), .IN2(n12761), .Q(n12760) );
  OR2X1 U12788 ( .IN1(n12762), .IN2(n12763), .Q(g27769) );
  AND2X1 U12789 ( .IN1(n12759), .IN2(n10398), .Q(n12763) );
  AND2X1 U12790 ( .IN1(n12764), .IN2(g2524), .Q(n12762) );
  OR2X1 U12791 ( .IN1(n4524), .IN2(n12761), .Q(n12764) );
  OR2X1 U12792 ( .IN1(n12765), .IN2(n12766), .Q(g27768) );
  AND2X1 U12793 ( .IN1(n12767), .IN2(n10403), .Q(n12766) );
  AND2X1 U12794 ( .IN1(n12768), .IN2(g1828), .Q(n12765) );
  OR2X1 U12795 ( .IN1(n4511), .IN2(n12769), .Q(n12768) );
  OR2X1 U12796 ( .IN1(n12770), .IN2(n12771), .Q(g27767) );
  AND2X1 U12797 ( .IN1(n12759), .IN2(n10408), .Q(n12771) );
  AND2X1 U12798 ( .IN1(test_so79), .IN2(n12772), .Q(n12759) );
  INVX0 U12799 ( .INP(n12773), .ZN(n12772) );
  OR2X1 U12800 ( .IN1(n12774), .IN2(n12775), .Q(n12773) );
  AND2X1 U12801 ( .IN1(n12776), .IN2(n12777), .Q(n12775) );
  OR2X1 U12802 ( .IN1(n12778), .IN2(n12779), .Q(n12776) );
  AND2X1 U12803 ( .IN1(n12780), .IN2(n12781), .Q(n12774) );
  OR2X1 U12804 ( .IN1(n12782), .IN2(n12783), .Q(n12781) );
  AND2X1 U12805 ( .IN1(n12784), .IN2(g2523), .Q(n12770) );
  OR2X1 U12806 ( .IN1(n4516), .IN2(n12761), .Q(n12784) );
  OR2X1 U12807 ( .IN1(n12785), .IN2(n12786), .Q(n12761) );
  OR2X1 U12808 ( .IN1(n12787), .IN2(n12788), .Q(n12786) );
  INVX0 U12809 ( .INP(n12789), .ZN(n12787) );
  OR2X1 U12810 ( .IN1(n12790), .IN2(n12791), .Q(g27766) );
  AND2X1 U12811 ( .IN1(n12767), .IN2(n10412), .Q(n12791) );
  AND2X1 U12812 ( .IN1(n12792), .IN2(g1830), .Q(n12790) );
  OR2X1 U12813 ( .IN1(n4525), .IN2(n12769), .Q(n12792) );
  OR2X1 U12814 ( .IN1(n12793), .IN2(n12794), .Q(g27765) );
  AND2X1 U12815 ( .IN1(n12795), .IN2(g1088), .Q(n12794) );
  AND2X1 U12816 ( .IN1(n12796), .IN2(g1134), .Q(n12793) );
  OR2X1 U12817 ( .IN1(n4381), .IN2(n12797), .Q(n12796) );
  OR2X1 U12818 ( .IN1(n12798), .IN2(n12799), .Q(g27764) );
  AND2X1 U12819 ( .IN1(n12767), .IN2(n10419), .Q(n12799) );
  AND2X1 U12820 ( .IN1(g1690), .IN2(n12800), .Q(n12767) );
  INVX0 U12821 ( .INP(n12801), .ZN(n12800) );
  OR2X1 U12822 ( .IN1(n12802), .IN2(n12803), .Q(n12801) );
  AND2X1 U12823 ( .IN1(n12804), .IN2(n12805), .Q(n12803) );
  OR2X1 U12824 ( .IN1(n12806), .IN2(n12807), .Q(n12804) );
  AND2X1 U12825 ( .IN1(n12808), .IN2(n12809), .Q(n12802) );
  OR2X1 U12826 ( .IN1(n12810), .IN2(n12811), .Q(n12809) );
  AND2X1 U12827 ( .IN1(n12812), .IN2(g1829), .Q(n12798) );
  OR2X1 U12828 ( .IN1(n4518), .IN2(n12769), .Q(n12812) );
  OR2X1 U12829 ( .IN1(n12813), .IN2(n12814), .Q(n12769) );
  OR2X1 U12830 ( .IN1(n12815), .IN2(n12816), .Q(n12814) );
  AND2X1 U12831 ( .IN1(n8777), .IN2(n10412), .Q(n12815) );
  OR2X1 U12832 ( .IN1(n12817), .IN2(n12818), .Q(g27763) );
  AND2X1 U12833 ( .IN1(n12795), .IN2(g6712), .Q(n12818) );
  AND2X1 U12834 ( .IN1(n12819), .IN2(g1136), .Q(n12817) );
  OR2X1 U12835 ( .IN1(n4364), .IN2(n12797), .Q(n12819) );
  OR2X1 U12836 ( .IN1(n12820), .IN2(n12821), .Q(g27762) );
  AND2X1 U12837 ( .IN1(n12822), .IN2(n10465), .Q(n12821) );
  AND2X1 U12838 ( .IN1(n12823), .IN2(g447), .Q(n12820) );
  OR2X1 U12839 ( .IN1(n4506), .IN2(n12824), .Q(n12823) );
  OR2X1 U12840 ( .IN1(n12825), .IN2(n12826), .Q(g27761) );
  AND2X1 U12841 ( .IN1(n12795), .IN2(g5472), .Q(n12826) );
  AND2X1 U12842 ( .IN1(g996), .IN2(n12827), .Q(n12795) );
  INVX0 U12843 ( .INP(n12828), .ZN(n12827) );
  OR2X1 U12844 ( .IN1(n12829), .IN2(n12830), .Q(n12828) );
  AND2X1 U12845 ( .IN1(n12831), .IN2(n12832), .Q(n12830) );
  OR2X1 U12846 ( .IN1(n12833), .IN2(n12834), .Q(n12831) );
  AND2X1 U12847 ( .IN1(n12835), .IN2(n12836), .Q(n12829) );
  OR2X1 U12848 ( .IN1(n12837), .IN2(n12838), .Q(n12836) );
  AND2X1 U12849 ( .IN1(n12839), .IN2(g1135), .Q(n12825) );
  OR2X1 U12850 ( .IN1(n4363), .IN2(n12797), .Q(n12839) );
  OR2X1 U12851 ( .IN1(n12840), .IN2(n12841), .Q(n12797) );
  OR2X1 U12852 ( .IN1(n12842), .IN2(n12843), .Q(n12841) );
  AND2X1 U12853 ( .IN1(n8780), .IN2(g6712), .Q(n12842) );
  OR2X1 U12854 ( .IN1(n12844), .IN2(n12845), .Q(g27760) );
  AND2X1 U12855 ( .IN1(n12822), .IN2(n10899), .Q(n12845) );
  AND2X1 U12856 ( .IN1(n12846), .IN2(g449), .Q(n12844) );
  OR2X1 U12857 ( .IN1(n4499), .IN2(n12824), .Q(n12846) );
  OR2X1 U12858 ( .IN1(n12847), .IN2(n12848), .Q(g27759) );
  AND2X1 U12859 ( .IN1(n12822), .IN2(n10475), .Q(n12848) );
  AND2X1 U12860 ( .IN1(g309), .IN2(n12849), .Q(n12822) );
  INVX0 U12861 ( .INP(n12850), .ZN(n12849) );
  OR2X1 U12862 ( .IN1(n12851), .IN2(n12852), .Q(n12850) );
  AND2X1 U12863 ( .IN1(n12853), .IN2(n12854), .Q(n12852) );
  OR2X1 U12864 ( .IN1(n12855), .IN2(n12856), .Q(n12853) );
  AND2X1 U12865 ( .IN1(n12857), .IN2(n12858), .Q(n12851) );
  OR2X1 U12866 ( .IN1(n12859), .IN2(n12860), .Q(n12858) );
  AND2X1 U12867 ( .IN1(n12861), .IN2(g448), .Q(n12847) );
  OR2X1 U12868 ( .IN1(n4520), .IN2(n12824), .Q(n12861) );
  OR2X1 U12869 ( .IN1(n12862), .IN2(n12863), .Q(n12824) );
  OR2X1 U12870 ( .IN1(n12864), .IN2(n12865), .Q(n12863) );
  AND2X1 U12871 ( .IN1(n8800), .IN2(n10465), .Q(n12864) );
  AND2X1 U12872 ( .IN1(n12866), .IN2(n12737), .Q(g27724) );
  XOR2X1 U12873 ( .IN1(n12739), .IN2(n4393), .Q(n12866) );
  AND2X1 U12874 ( .IN1(n12867), .IN2(n12741), .Q(g27722) );
  XNOR2X1 U12875 ( .IN1(test_so70), .IN2(n12743), .Q(n12867) );
  AND2X1 U12876 ( .IN1(n12868), .IN2(n12745), .Q(g27718) );
  XOR2X1 U12877 ( .IN1(n12747), .IN2(n4395), .Q(n12868) );
  AND2X1 U12878 ( .IN1(n12869), .IN2(n12870), .Q(g27682) );
  INVX0 U12879 ( .INP(n12871), .ZN(n12870) );
  AND2X1 U12880 ( .IN1(n12872), .IN2(n4473), .Q(n12871) );
  OR2X1 U12881 ( .IN1(n12873), .IN2(n4468), .Q(n12872) );
  AND2X1 U12882 ( .IN1(n12743), .IN2(n12741), .Q(n12869) );
  OR2X1 U12883 ( .IN1(n12873), .IN2(n12874), .Q(n12743) );
  OR2X1 U12884 ( .IN1(n4473), .IN2(n4468), .Q(n12874) );
  AND2X1 U12885 ( .IN1(n12875), .IN2(n12876), .Q(g27678) );
  INVX0 U12886 ( .INP(n12877), .ZN(n12876) );
  AND2X1 U12887 ( .IN1(n12878), .IN2(n4475), .Q(n12877) );
  OR2X1 U12888 ( .IN1(n12879), .IN2(n4469), .Q(n12878) );
  AND2X1 U12889 ( .IN1(n12747), .IN2(n12745), .Q(n12875) );
  OR2X1 U12890 ( .IN1(n12879), .IN2(n12880), .Q(n12747) );
  OR2X1 U12891 ( .IN1(n4475), .IN2(n4469), .Q(n12880) );
  AND2X1 U12892 ( .IN1(n12881), .IN2(n12882), .Q(g27672) );
  INVX0 U12893 ( .INP(n12883), .ZN(n12882) );
  AND2X1 U12894 ( .IN1(n12884), .IN2(n4477), .Q(n12883) );
  OR2X1 U12895 ( .IN1(n9123), .IN2(n12885), .Q(n12884) );
  AND2X1 U12896 ( .IN1(n12228), .IN2(n12226), .Q(n12881) );
  OR2X1 U12897 ( .IN1(n9123), .IN2(n12886), .Q(n12228) );
  OR2X1 U12898 ( .IN1(n4477), .IN2(n12885), .Q(n12886) );
  AND2X1 U12899 ( .IN1(n12887), .IN2(n11527), .Q(g27621) );
  XOR2X1 U12900 ( .IN1(n8807), .IN2(n4522), .Q(n12887) );
  AND2X1 U12901 ( .IN1(n12888), .IN2(n11529), .Q(g27612) );
  XOR2X1 U12902 ( .IN1(n8811), .IN2(n4523), .Q(n12888) );
  AND2X1 U12903 ( .IN1(n12889), .IN2(n11531), .Q(g27603) );
  XNOR2X1 U12904 ( .IN1(n12890), .IN2(n8815), .Q(n12889) );
  AND2X1 U12905 ( .IN1(n12891), .IN2(n11533), .Q(g27594) );
  XOR2X1 U12906 ( .IN1(n8819), .IN2(n4521), .Q(n12891) );
  OR2X1 U12907 ( .IN1(n12892), .IN2(n12893), .Q(g27380) );
  OR2X1 U12908 ( .IN1(n12894), .IN2(n12895), .Q(n12893) );
  OR2X1 U12909 ( .IN1(n12896), .IN2(n12897), .Q(n12895) );
  AND2X1 U12910 ( .IN1(n8545), .IN2(n12898), .Q(n12897) );
  AND2X1 U12911 ( .IN1(n12899), .IN2(n8079), .Q(n12896) );
  OR2X1 U12912 ( .IN1(n12900), .IN2(n12901), .Q(n12892) );
  OR2X1 U12913 ( .IN1(n12902), .IN2(n12903), .Q(n12901) );
  AND2X1 U12914 ( .IN1(n12904), .IN2(g3151), .Q(n12903) );
  AND2X1 U12915 ( .IN1(n12905), .IN2(n12906), .Q(n12902) );
  OR2X1 U12916 ( .IN1(n12907), .IN2(n3705), .Q(n12906) );
  AND2X1 U12917 ( .IN1(n4384), .IN2(n12908), .Q(n12907) );
  OR2X1 U12918 ( .IN1(n12909), .IN2(n12910), .Q(n12900) );
  AND2X1 U12919 ( .IN1(n12911), .IN2(n12912), .Q(n12910) );
  INVX0 U12920 ( .INP(n12913), .ZN(n12912) );
  OR2X1 U12921 ( .IN1(n12914), .IN2(n12915), .Q(n12913) );
  AND2X1 U12922 ( .IN1(n8081), .IN2(n12916), .Q(n12915) );
  AND2X1 U12923 ( .IN1(n8082), .IN2(n12917), .Q(n12914) );
  AND2X1 U12924 ( .IN1(n12918), .IN2(n12919), .Q(n12911) );
  OR2X1 U12925 ( .IN1(n12920), .IN2(n12921), .Q(g27354) );
  AND2X1 U12926 ( .IN1(n12922), .IN2(n12923), .Q(n12921) );
  INVX0 U12927 ( .INP(n12924), .ZN(n12920) );
  OR2X1 U12928 ( .IN1(n12922), .IN2(n8465), .Q(n12924) );
  OR2X1 U12929 ( .IN1(n12925), .IN2(n12926), .Q(g27348) );
  AND2X1 U12930 ( .IN1(n12927), .IN2(n12923), .Q(n12926) );
  INVX0 U12931 ( .INP(n12928), .ZN(n12925) );
  OR2X1 U12932 ( .IN1(n12927), .IN2(n8466), .Q(n12928) );
  OR2X1 U12933 ( .IN1(n12929), .IN2(n12930), .Q(g27347) );
  AND2X1 U12934 ( .IN1(n12922), .IN2(n12931), .Q(n12930) );
  INVX0 U12935 ( .INP(n12932), .ZN(n12929) );
  OR2X1 U12936 ( .IN1(n12922), .IN2(n8288), .Q(n12932) );
  OR2X1 U12937 ( .IN1(n12933), .IN2(n12934), .Q(g27346) );
  AND2X1 U12938 ( .IN1(n12935), .IN2(n12936), .Q(n12934) );
  INVX0 U12939 ( .INP(n12937), .ZN(n12933) );
  OR2X1 U12940 ( .IN1(n12935), .IN2(n8467), .Q(n12937) );
  OR2X1 U12941 ( .IN1(n12938), .IN2(n12939), .Q(g27345) );
  AND2X1 U12942 ( .IN1(n12940), .IN2(n12923), .Q(n12939) );
  OR2X1 U12943 ( .IN1(n12941), .IN2(n12942), .Q(n12923) );
  OR2X1 U12944 ( .IN1(n12323), .IN2(n12289), .Q(n12942) );
  INVX0 U12945 ( .INP(n12943), .ZN(n12938) );
  OR2X1 U12946 ( .IN1(n12940), .IN2(n8464), .Q(n12943) );
  OR2X1 U12947 ( .IN1(n12944), .IN2(n12945), .Q(g27344) );
  AND2X1 U12948 ( .IN1(n12927), .IN2(n12931), .Q(n12945) );
  AND2X1 U12949 ( .IN1(test_so89), .IN2(n12946), .Q(n12944) );
  INVX0 U12950 ( .INP(n12927), .ZN(n12946) );
  OR2X1 U12951 ( .IN1(n12947), .IN2(n12948), .Q(g27343) );
  AND2X1 U12952 ( .IN1(n12949), .IN2(n12922), .Q(n12948) );
  INVX0 U12953 ( .INP(n12950), .ZN(n12947) );
  OR2X1 U12954 ( .IN1(n12922), .IN2(n8454), .Q(n12950) );
  OR2X1 U12955 ( .IN1(n12951), .IN2(n12952), .Q(g27342) );
  AND2X1 U12956 ( .IN1(n12953), .IN2(n12954), .Q(n12952) );
  INVX0 U12957 ( .INP(n12955), .ZN(n12951) );
  OR2X1 U12958 ( .IN1(n12953), .IN2(n8751), .Q(n12955) );
  OR2X1 U12959 ( .IN1(n12956), .IN2(n12957), .Q(g27341) );
  AND2X1 U12960 ( .IN1(n12958), .IN2(n12936), .Q(n12957) );
  INVX0 U12961 ( .INP(n12959), .ZN(n12956) );
  OR2X1 U12962 ( .IN1(n12958), .IN2(n8468), .Q(n12959) );
  OR2X1 U12963 ( .IN1(n12960), .IN2(n12961), .Q(g27340) );
  AND2X1 U12964 ( .IN1(n12935), .IN2(n12962), .Q(n12961) );
  INVX0 U12965 ( .INP(n12963), .ZN(n12960) );
  OR2X1 U12966 ( .IN1(n12935), .IN2(n8290), .Q(n12963) );
  OR2X1 U12967 ( .IN1(n12964), .IN2(n12965), .Q(g27339) );
  AND2X1 U12968 ( .IN1(n12966), .IN2(n12967), .Q(n12965) );
  INVX0 U12969 ( .INP(n12968), .ZN(n12964) );
  OR2X1 U12970 ( .IN1(n12966), .IN2(n8470), .Q(n12968) );
  OR2X1 U12971 ( .IN1(n12969), .IN2(n12970), .Q(g27338) );
  AND2X1 U12972 ( .IN1(n12940), .IN2(n12931), .Q(n12970) );
  AND2X1 U12973 ( .IN1(n12971), .IN2(n12972), .Q(n12931) );
  OR2X1 U12974 ( .IN1(n12941), .IN2(n12307), .Q(n12972) );
  INVX0 U12975 ( .INP(n12973), .ZN(n12971) );
  AND2X1 U12976 ( .IN1(n12346), .IN2(n12941), .Q(n12973) );
  INVX0 U12977 ( .INP(n12974), .ZN(n12941) );
  AND2X1 U12978 ( .IN1(n12324), .IN2(n12307), .Q(n12346) );
  INVX0 U12979 ( .INP(n12975), .ZN(n12969) );
  OR2X1 U12980 ( .IN1(n12940), .IN2(n8287), .Q(n12975) );
  OR2X1 U12981 ( .IN1(n12976), .IN2(n12977), .Q(g27337) );
  AND2X1 U12982 ( .IN1(n12949), .IN2(n12927), .Q(n12977) );
  INVX0 U12983 ( .INP(n12978), .ZN(n12976) );
  OR2X1 U12984 ( .IN1(n12927), .IN2(n8455), .Q(n12978) );
  OR2X1 U12985 ( .IN1(n12979), .IN2(n12980), .Q(g27336) );
  AND2X1 U12986 ( .IN1(n12981), .IN2(n12922), .Q(n12980) );
  INVX0 U12987 ( .INP(n12982), .ZN(n12979) );
  OR2X1 U12988 ( .IN1(n12922), .IN2(n8442), .Q(n12982) );
  AND2X1 U12989 ( .IN1(g2624), .IN2(g22687), .Q(n12922) );
  OR2X1 U12990 ( .IN1(n12983), .IN2(n12984), .Q(g27335) );
  AND2X1 U12991 ( .IN1(n12985), .IN2(n12954), .Q(n12984) );
  INVX0 U12992 ( .INP(n12986), .ZN(n12983) );
  OR2X1 U12993 ( .IN1(n12985), .IN2(n8752), .Q(n12986) );
  OR2X1 U12994 ( .IN1(n12987), .IN2(n12988), .Q(g27334) );
  AND2X1 U12995 ( .IN1(n12953), .IN2(n12989), .Q(n12988) );
  INVX0 U12996 ( .INP(n12990), .ZN(n12987) );
  OR2X1 U12997 ( .IN1(n12953), .IN2(n8487), .Q(n12990) );
  OR2X1 U12998 ( .IN1(n12991), .IN2(n12992), .Q(g27333) );
  AND2X1 U12999 ( .IN1(n12993), .IN2(n12936), .Q(n12992) );
  OR2X1 U13000 ( .IN1(n12994), .IN2(n12995), .Q(n12936) );
  OR2X1 U13001 ( .IN1(n12447), .IN2(n12413), .Q(n12995) );
  INVX0 U13002 ( .INP(n12996), .ZN(n12991) );
  OR2X1 U13003 ( .IN1(n9125), .IN2(n12993), .Q(n12996) );
  OR2X1 U13004 ( .IN1(n12997), .IN2(n12998), .Q(g27332) );
  AND2X1 U13005 ( .IN1(n12958), .IN2(n12962), .Q(n12998) );
  INVX0 U13006 ( .INP(n12999), .ZN(n12997) );
  OR2X1 U13007 ( .IN1(n12958), .IN2(n8291), .Q(n12999) );
  OR2X1 U13008 ( .IN1(n13000), .IN2(n13001), .Q(g27331) );
  AND2X1 U13009 ( .IN1(n13002), .IN2(n12935), .Q(n13001) );
  INVX0 U13010 ( .INP(n13003), .ZN(n13000) );
  OR2X1 U13011 ( .IN1(n12935), .IN2(n8457), .Q(n13003) );
  OR2X1 U13012 ( .IN1(n13004), .IN2(n13005), .Q(g27330) );
  AND2X1 U13013 ( .IN1(n13006), .IN2(n13007), .Q(n13005) );
  INVX0 U13014 ( .INP(n13008), .ZN(n13004) );
  OR2X1 U13015 ( .IN1(n13006), .IN2(n8754), .Q(n13008) );
  OR2X1 U13016 ( .IN1(n13009), .IN2(n13010), .Q(g27329) );
  AND2X1 U13017 ( .IN1(n13011), .IN2(n12967), .Q(n13010) );
  INVX0 U13018 ( .INP(n13012), .ZN(n13009) );
  OR2X1 U13019 ( .IN1(n13011), .IN2(n8471), .Q(n13012) );
  OR2X1 U13020 ( .IN1(n13013), .IN2(n13014), .Q(g27328) );
  AND2X1 U13021 ( .IN1(n12966), .IN2(n13015), .Q(n13014) );
  AND2X1 U13022 ( .IN1(test_so46), .IN2(n13016), .Q(n13013) );
  INVX0 U13023 ( .INP(n12966), .ZN(n13016) );
  OR2X1 U13024 ( .IN1(n13017), .IN2(n13018), .Q(g27327) );
  AND2X1 U13025 ( .IN1(n13019), .IN2(n13020), .Q(n13018) );
  INVX0 U13026 ( .INP(n13021), .ZN(n13017) );
  OR2X1 U13027 ( .IN1(n13019), .IN2(n8473), .Q(n13021) );
  OR2X1 U13028 ( .IN1(n13022), .IN2(n13023), .Q(g27326) );
  AND2X1 U13029 ( .IN1(n12949), .IN2(n12940), .Q(n13023) );
  AND2X1 U13030 ( .IN1(n13024), .IN2(n13025), .Q(n12949) );
  OR2X1 U13031 ( .IN1(n12974), .IN2(n12294), .Q(n13024) );
  INVX0 U13032 ( .INP(n12323), .ZN(n12294) );
  XNOR2X1 U13033 ( .IN1(g3229), .IN2(n12317), .Q(n12974) );
  INVX0 U13034 ( .INP(n12304), .ZN(n12317) );
  INVX0 U13035 ( .INP(n13026), .ZN(n13022) );
  OR2X1 U13036 ( .IN1(n12940), .IN2(n8453), .Q(n13026) );
  OR2X1 U13037 ( .IN1(n13027), .IN2(n13028), .Q(g27325) );
  AND2X1 U13038 ( .IN1(n12981), .IN2(n12927), .Q(n13028) );
  INVX0 U13039 ( .INP(n13029), .ZN(n13027) );
  OR2X1 U13040 ( .IN1(n12927), .IN2(n8443), .Q(n13029) );
  AND2X1 U13041 ( .IN1(g7390), .IN2(g22687), .Q(n12927) );
  OR2X1 U13042 ( .IN1(n13030), .IN2(n13031), .Q(g27324) );
  AND2X1 U13043 ( .IN1(n13032), .IN2(n12954), .Q(n13031) );
  OR2X1 U13044 ( .IN1(n13033), .IN2(n13034), .Q(n12954) );
  OR2X1 U13045 ( .IN1(n13035), .IN2(n13036), .Q(n13034) );
  INVX0 U13046 ( .INP(n13037), .ZN(n13030) );
  OR2X1 U13047 ( .IN1(n13032), .IN2(n8753), .Q(n13037) );
  OR2X1 U13048 ( .IN1(n13038), .IN2(n13039), .Q(g27323) );
  AND2X1 U13049 ( .IN1(n12985), .IN2(n12989), .Q(n13039) );
  INVX0 U13050 ( .INP(n13040), .ZN(n13038) );
  OR2X1 U13051 ( .IN1(n12985), .IN2(n8488), .Q(n13040) );
  OR2X1 U13052 ( .IN1(n13041), .IN2(n13042), .Q(g27322) );
  AND2X1 U13053 ( .IN1(n13043), .IN2(n12953), .Q(n13042) );
  INVX0 U13054 ( .INP(n13044), .ZN(n13041) );
  OR2X1 U13055 ( .IN1(n12953), .IN2(n8739), .Q(n13044) );
  OR2X1 U13056 ( .IN1(n13045), .IN2(n13046), .Q(g27321) );
  AND2X1 U13057 ( .IN1(n12993), .IN2(n12962), .Q(n13046) );
  AND2X1 U13058 ( .IN1(n13047), .IN2(n13048), .Q(n12962) );
  OR2X1 U13059 ( .IN1(n12994), .IN2(n12431), .Q(n13048) );
  INVX0 U13060 ( .INP(n13049), .ZN(n13047) );
  AND2X1 U13061 ( .IN1(n12470), .IN2(n12994), .Q(n13049) );
  INVX0 U13062 ( .INP(n13050), .ZN(n12994) );
  AND2X1 U13063 ( .IN1(n12448), .IN2(n12431), .Q(n12470) );
  INVX0 U13064 ( .INP(n13051), .ZN(n13045) );
  OR2X1 U13065 ( .IN1(n12993), .IN2(n8289), .Q(n13051) );
  OR2X1 U13066 ( .IN1(n13052), .IN2(n13053), .Q(g27320) );
  AND2X1 U13067 ( .IN1(n13002), .IN2(n12958), .Q(n13053) );
  INVX0 U13068 ( .INP(n13054), .ZN(n13052) );
  OR2X1 U13069 ( .IN1(n12958), .IN2(n8458), .Q(n13054) );
  OR2X1 U13070 ( .IN1(n13055), .IN2(n13056), .Q(g27319) );
  AND2X1 U13071 ( .IN1(n13057), .IN2(n12935), .Q(n13056) );
  INVX0 U13072 ( .INP(n13058), .ZN(n13055) );
  OR2X1 U13073 ( .IN1(n12935), .IN2(n8445), .Q(n13058) );
  AND2X1 U13074 ( .IN1(g1930), .IN2(g22651), .Q(n12935) );
  OR2X1 U13075 ( .IN1(n13059), .IN2(n13060), .Q(g27318) );
  AND2X1 U13076 ( .IN1(n13061), .IN2(n13007), .Q(n13060) );
  AND2X1 U13077 ( .IN1(test_so58), .IN2(n13062), .Q(n13059) );
  INVX0 U13078 ( .INP(n13061), .ZN(n13062) );
  OR2X1 U13079 ( .IN1(n13063), .IN2(n13064), .Q(g27317) );
  AND2X1 U13080 ( .IN1(n13006), .IN2(n13065), .Q(n13064) );
  INVX0 U13081 ( .INP(n13066), .ZN(n13063) );
  OR2X1 U13082 ( .IN1(n13006), .IN2(n8490), .Q(n13066) );
  OR2X1 U13083 ( .IN1(n13067), .IN2(n13068), .Q(g27316) );
  AND2X1 U13084 ( .IN1(n13069), .IN2(n12967), .Q(n13068) );
  OR2X1 U13085 ( .IN1(n13070), .IN2(n13071), .Q(n12967) );
  OR2X1 U13086 ( .IN1(n12567), .IN2(n12533), .Q(n13071) );
  INVX0 U13087 ( .INP(n13072), .ZN(n13067) );
  OR2X1 U13088 ( .IN1(n13069), .IN2(n8469), .Q(n13072) );
  OR2X1 U13089 ( .IN1(n13073), .IN2(n13074), .Q(g27315) );
  AND2X1 U13090 ( .IN1(n13011), .IN2(n13015), .Q(n13074) );
  INVX0 U13091 ( .INP(n13075), .ZN(n13073) );
  OR2X1 U13092 ( .IN1(n13011), .IN2(n8293), .Q(n13075) );
  OR2X1 U13093 ( .IN1(n13076), .IN2(n13077), .Q(g27314) );
  AND2X1 U13094 ( .IN1(n13078), .IN2(n12966), .Q(n13077) );
  INVX0 U13095 ( .INP(n13079), .ZN(n13076) );
  OR2X1 U13096 ( .IN1(n12966), .IN2(n8460), .Q(n13079) );
  OR2X1 U13097 ( .IN1(n13080), .IN2(n13081), .Q(g27313) );
  AND2X1 U13098 ( .IN1(n13082), .IN2(n13083), .Q(n13081) );
  INVX0 U13099 ( .INP(n13084), .ZN(n13080) );
  OR2X1 U13100 ( .IN1(n13082), .IN2(n8756), .Q(n13084) );
  OR2X1 U13101 ( .IN1(n13085), .IN2(n13086), .Q(g27312) );
  AND2X1 U13102 ( .IN1(n13087), .IN2(n13020), .Q(n13086) );
  INVX0 U13103 ( .INP(n13088), .ZN(n13085) );
  OR2X1 U13104 ( .IN1(n13087), .IN2(n8474), .Q(n13088) );
  OR2X1 U13105 ( .IN1(n13089), .IN2(n13090), .Q(g27311) );
  AND2X1 U13106 ( .IN1(n13019), .IN2(n13091), .Q(n13090) );
  INVX0 U13107 ( .INP(n13092), .ZN(n13089) );
  OR2X1 U13108 ( .IN1(n13019), .IN2(n8295), .Q(n13092) );
  OR2X1 U13109 ( .IN1(n13093), .IN2(n13094), .Q(g27310) );
  AND2X1 U13110 ( .IN1(n12981), .IN2(n12940), .Q(n13094) );
  INVX0 U13111 ( .INP(n13095), .ZN(n12981) );
  OR2X1 U13112 ( .IN1(n13096), .IN2(n13097), .Q(n13095) );
  OR2X1 U13113 ( .IN1(n13098), .IN2(n13099), .Q(n13097) );
  AND2X1 U13114 ( .IN1(n13100), .IN2(n13025), .Q(n13099) );
  AND2X1 U13115 ( .IN1(n12324), .IN2(n12304), .Q(n13100) );
  OR2X1 U13116 ( .IN1(n13101), .IN2(n13102), .Q(n12304) );
  OR2X1 U13117 ( .IN1(n13103), .IN2(n13104), .Q(n13102) );
  AND2X1 U13118 ( .IN1(n8441), .IN2(n11411), .Q(n13104) );
  AND2X1 U13119 ( .IN1(n8442), .IN2(g2624), .Q(n13103) );
  AND2X1 U13120 ( .IN1(n8443), .IN2(g7390), .Q(n13101) );
  INVX0 U13121 ( .INP(n12301), .ZN(n12324) );
  INVX0 U13122 ( .INP(n13105), .ZN(n13098) );
  OR2X1 U13123 ( .IN1(n13025), .IN2(g3229), .Q(n13105) );
  OR2X1 U13124 ( .IN1(n12307), .IN2(n12323), .Q(n13025) );
  OR2X1 U13125 ( .IN1(n13106), .IN2(n13107), .Q(n12323) );
  OR2X1 U13126 ( .IN1(n13108), .IN2(n13109), .Q(n13107) );
  AND2X1 U13127 ( .IN1(n8287), .IN2(n11411), .Q(n13109) );
  AND2X1 U13128 ( .IN1(n8288), .IN2(g2624), .Q(n13108) );
  INVX0 U13129 ( .INP(n13110), .ZN(n13106) );
  OR2X1 U13130 ( .IN1(n4370), .IN2(test_so89), .Q(n13110) );
  INVX0 U13131 ( .INP(n12289), .ZN(n12307) );
  OR2X1 U13132 ( .IN1(n13111), .IN2(n13112), .Q(n12289) );
  OR2X1 U13133 ( .IN1(n13113), .IN2(n13114), .Q(n13112) );
  AND2X1 U13134 ( .IN1(n8453), .IN2(n11411), .Q(n13114) );
  AND2X1 U13135 ( .IN1(n8454), .IN2(g2624), .Q(n13113) );
  AND2X1 U13136 ( .IN1(n8455), .IN2(g7390), .Q(n13111) );
  AND2X1 U13137 ( .IN1(g3229), .IN2(n12301), .Q(n13096) );
  OR2X1 U13138 ( .IN1(n13115), .IN2(n13116), .Q(n12301) );
  OR2X1 U13139 ( .IN1(n13117), .IN2(n13118), .Q(n13116) );
  AND2X1 U13140 ( .IN1(n8464), .IN2(n11411), .Q(n13118) );
  AND2X1 U13141 ( .IN1(n8465), .IN2(g2624), .Q(n13117) );
  AND2X1 U13142 ( .IN1(n8466), .IN2(g7390), .Q(n13115) );
  INVX0 U13143 ( .INP(n13119), .ZN(n13093) );
  OR2X1 U13144 ( .IN1(n12940), .IN2(n8441), .Q(n13119) );
  AND2X1 U13145 ( .IN1(g22687), .IN2(g7302), .Q(n12940) );
  OR2X1 U13146 ( .IN1(n13120), .IN2(n13121), .Q(g27309) );
  AND2X1 U13147 ( .IN1(n13032), .IN2(n12989), .Q(n13121) );
  AND2X1 U13148 ( .IN1(n13122), .IN2(n13123), .Q(n12989) );
  OR2X1 U13149 ( .IN1(n13124), .IN2(n13033), .Q(n13123) );
  OR2X1 U13150 ( .IN1(n13125), .IN2(n13126), .Q(n13124) );
  OR2X1 U13151 ( .IN1(n13036), .IN2(n13127), .Q(n13122) );
  INVX0 U13152 ( .INP(n13128), .ZN(n13120) );
  OR2X1 U13153 ( .IN1(n13032), .IN2(n8486), .Q(n13128) );
  OR2X1 U13154 ( .IN1(n13129), .IN2(n13130), .Q(g27308) );
  AND2X1 U13155 ( .IN1(n13043), .IN2(n12985), .Q(n13130) );
  INVX0 U13156 ( .INP(n13131), .ZN(n13129) );
  OR2X1 U13157 ( .IN1(n12985), .IN2(n8740), .Q(n13131) );
  OR2X1 U13158 ( .IN1(n13132), .IN2(n13133), .Q(g27307) );
  AND2X1 U13159 ( .IN1(n13134), .IN2(n12953), .Q(n13133) );
  INVX0 U13160 ( .INP(n13135), .ZN(n13132) );
  OR2X1 U13161 ( .IN1(n12953), .IN2(n8762), .Q(n13135) );
  AND2X1 U13162 ( .IN1(n10833), .IN2(n13136), .Q(n12953) );
  OR2X1 U13163 ( .IN1(n13137), .IN2(n13138), .Q(g27306) );
  AND2X1 U13164 ( .IN1(n13002), .IN2(n12993), .Q(n13138) );
  AND2X1 U13165 ( .IN1(n13139), .IN2(n13140), .Q(n13002) );
  OR2X1 U13166 ( .IN1(n13050), .IN2(n12418), .Q(n13139) );
  INVX0 U13167 ( .INP(n12447), .ZN(n12418) );
  XNOR2X1 U13168 ( .IN1(g3229), .IN2(n12441), .Q(n13050) );
  INVX0 U13169 ( .INP(n12428), .ZN(n12441) );
  INVX0 U13170 ( .INP(n13141), .ZN(n13137) );
  OR2X1 U13171 ( .IN1(n12993), .IN2(n8456), .Q(n13141) );
  OR2X1 U13172 ( .IN1(n13142), .IN2(n13143), .Q(g27305) );
  AND2X1 U13173 ( .IN1(n13057), .IN2(n12958), .Q(n13143) );
  INVX0 U13174 ( .INP(n13144), .ZN(n13142) );
  OR2X1 U13175 ( .IN1(n12958), .IN2(n8446), .Q(n13144) );
  AND2X1 U13176 ( .IN1(g7194), .IN2(g22651), .Q(n12958) );
  OR2X1 U13177 ( .IN1(n13145), .IN2(n13146), .Q(g27304) );
  AND2X1 U13178 ( .IN1(n13147), .IN2(n13007), .Q(n13146) );
  OR2X1 U13179 ( .IN1(n13148), .IN2(n13149), .Q(n13007) );
  OR2X1 U13180 ( .IN1(n13150), .IN2(n13151), .Q(n13149) );
  INVX0 U13181 ( .INP(n13152), .ZN(n13145) );
  OR2X1 U13182 ( .IN1(n13147), .IN2(n8755), .Q(n13152) );
  OR2X1 U13183 ( .IN1(n13153), .IN2(n13154), .Q(g27303) );
  AND2X1 U13184 ( .IN1(n13061), .IN2(n13065), .Q(n13154) );
  INVX0 U13185 ( .INP(n13155), .ZN(n13153) );
  OR2X1 U13186 ( .IN1(n13061), .IN2(n8491), .Q(n13155) );
  OR2X1 U13187 ( .IN1(n13156), .IN2(n13157), .Q(g27302) );
  AND2X1 U13188 ( .IN1(n13158), .IN2(n13006), .Q(n13157) );
  INVX0 U13189 ( .INP(n13159), .ZN(n13156) );
  OR2X1 U13190 ( .IN1(n13006), .IN2(n8742), .Q(n13159) );
  OR2X1 U13191 ( .IN1(n13160), .IN2(n13161), .Q(g27301) );
  AND2X1 U13192 ( .IN1(n13069), .IN2(n13015), .Q(n13161) );
  AND2X1 U13193 ( .IN1(n13162), .IN2(n13163), .Q(n13015) );
  OR2X1 U13194 ( .IN1(n13070), .IN2(n12551), .Q(n13163) );
  INVX0 U13195 ( .INP(n13164), .ZN(n13162) );
  AND2X1 U13196 ( .IN1(n12590), .IN2(n13070), .Q(n13164) );
  INVX0 U13197 ( .INP(n13165), .ZN(n13070) );
  AND2X1 U13198 ( .IN1(n12568), .IN2(n12551), .Q(n12590) );
  INVX0 U13199 ( .INP(n13166), .ZN(n13160) );
  OR2X1 U13200 ( .IN1(n13069), .IN2(n8292), .Q(n13166) );
  OR2X1 U13201 ( .IN1(n13167), .IN2(n13168), .Q(g27300) );
  AND2X1 U13202 ( .IN1(n13078), .IN2(n13011), .Q(n13168) );
  INVX0 U13203 ( .INP(n13169), .ZN(n13167) );
  OR2X1 U13204 ( .IN1(n13011), .IN2(n8461), .Q(n13169) );
  OR2X1 U13205 ( .IN1(n13170), .IN2(n13171), .Q(g27299) );
  AND2X1 U13206 ( .IN1(n13172), .IN2(n12966), .Q(n13171) );
  INVX0 U13207 ( .INP(n13173), .ZN(n13170) );
  OR2X1 U13208 ( .IN1(n12966), .IN2(n8448), .Q(n13173) );
  AND2X1 U13209 ( .IN1(g1236), .IN2(g22615), .Q(n12966) );
  OR2X1 U13210 ( .IN1(n13174), .IN2(n13175), .Q(g27298) );
  AND2X1 U13211 ( .IN1(n13176), .IN2(n13083), .Q(n13175) );
  INVX0 U13212 ( .INP(n13177), .ZN(n13174) );
  OR2X1 U13213 ( .IN1(n13176), .IN2(n8757), .Q(n13177) );
  OR2X1 U13214 ( .IN1(n13178), .IN2(n13179), .Q(g27297) );
  AND2X1 U13215 ( .IN1(n13082), .IN2(n13180), .Q(n13179) );
  INVX0 U13216 ( .INP(n13181), .ZN(n13178) );
  OR2X1 U13217 ( .IN1(n13082), .IN2(n8493), .Q(n13181) );
  OR2X1 U13218 ( .IN1(n13182), .IN2(n13183), .Q(g27296) );
  AND2X1 U13219 ( .IN1(n13184), .IN2(n13020), .Q(n13183) );
  OR2X1 U13220 ( .IN1(n13185), .IN2(n13186), .Q(n13020) );
  OR2X1 U13221 ( .IN1(n12682), .IN2(n12648), .Q(n13186) );
  INVX0 U13222 ( .INP(n13187), .ZN(n13182) );
  OR2X1 U13223 ( .IN1(n13184), .IN2(n8472), .Q(n13187) );
  OR2X1 U13224 ( .IN1(n13188), .IN2(n13189), .Q(g27295) );
  AND2X1 U13225 ( .IN1(n13087), .IN2(n13091), .Q(n13189) );
  INVX0 U13226 ( .INP(n13190), .ZN(n13188) );
  OR2X1 U13227 ( .IN1(n13087), .IN2(n8296), .Q(n13190) );
  OR2X1 U13228 ( .IN1(n13191), .IN2(n13192), .Q(g27294) );
  AND2X1 U13229 ( .IN1(n13193), .IN2(n13019), .Q(n13192) );
  INVX0 U13230 ( .INP(n13194), .ZN(n13191) );
  OR2X1 U13231 ( .IN1(n13019), .IN2(n8463), .Q(n13194) );
  OR2X1 U13232 ( .IN1(n13195), .IN2(n13196), .Q(g27293) );
  AND2X1 U13233 ( .IN1(n13197), .IN2(n13198), .Q(n13196) );
  INVX0 U13234 ( .INP(n13199), .ZN(n13195) );
  OR2X1 U13235 ( .IN1(n13197), .IN2(n8759), .Q(n13199) );
  OR2X1 U13236 ( .IN1(n13200), .IN2(n13201), .Q(g27292) );
  AND2X1 U13237 ( .IN1(n13043), .IN2(n13032), .Q(n13201) );
  INVX0 U13238 ( .INP(n13202), .ZN(n13043) );
  OR2X1 U13239 ( .IN1(n13203), .IN2(n13204), .Q(n13202) );
  AND2X1 U13240 ( .IN1(n13036), .IN2(n13035), .Q(n13203) );
  INVX0 U13241 ( .INP(n13126), .ZN(n13036) );
  XOR2X1 U13242 ( .IN1(g3229), .IN2(n13205), .Q(n13126) );
  INVX0 U13243 ( .INP(n13206), .ZN(n13200) );
  OR2X1 U13244 ( .IN1(n13032), .IN2(n8741), .Q(n13206) );
  OR2X1 U13245 ( .IN1(n13207), .IN2(n13208), .Q(g27291) );
  AND2X1 U13246 ( .IN1(n13134), .IN2(n12985), .Q(n13208) );
  INVX0 U13247 ( .INP(n13209), .ZN(n13207) );
  OR2X1 U13248 ( .IN1(n12985), .IN2(n8763), .Q(n13209) );
  AND2X1 U13249 ( .IN1(g7264), .IN2(n13136), .Q(n12985) );
  OR2X1 U13250 ( .IN1(n13210), .IN2(n13211), .Q(g27290) );
  AND2X1 U13251 ( .IN1(n13057), .IN2(n12993), .Q(n13211) );
  INVX0 U13252 ( .INP(n13212), .ZN(n13057) );
  OR2X1 U13253 ( .IN1(n13213), .IN2(n13214), .Q(n13212) );
  OR2X1 U13254 ( .IN1(n13215), .IN2(n13216), .Q(n13214) );
  AND2X1 U13255 ( .IN1(n13217), .IN2(n13140), .Q(n13216) );
  AND2X1 U13256 ( .IN1(n12448), .IN2(n12428), .Q(n13217) );
  OR2X1 U13257 ( .IN1(n13218), .IN2(n13219), .Q(n12428) );
  OR2X1 U13258 ( .IN1(n13220), .IN2(n13221), .Q(n13219) );
  AND2X1 U13259 ( .IN1(n8446), .IN2(g7194), .Q(n13221) );
  AND2X1 U13260 ( .IN1(n8444), .IN2(n12379), .Q(n13220) );
  AND2X1 U13261 ( .IN1(n8445), .IN2(g1930), .Q(n13218) );
  INVX0 U13262 ( .INP(n12425), .ZN(n12448) );
  INVX0 U13263 ( .INP(n13222), .ZN(n13215) );
  OR2X1 U13264 ( .IN1(n13140), .IN2(g3229), .Q(n13222) );
  OR2X1 U13265 ( .IN1(n12431), .IN2(n12447), .Q(n13140) );
  OR2X1 U13266 ( .IN1(n13223), .IN2(n13224), .Q(n12447) );
  OR2X1 U13267 ( .IN1(n13225), .IN2(n13226), .Q(n13224) );
  AND2X1 U13268 ( .IN1(n8291), .IN2(g7194), .Q(n13226) );
  AND2X1 U13269 ( .IN1(n8289), .IN2(n12379), .Q(n13225) );
  AND2X1 U13270 ( .IN1(n8290), .IN2(g1930), .Q(n13223) );
  INVX0 U13271 ( .INP(n12413), .ZN(n12431) );
  OR2X1 U13272 ( .IN1(n13227), .IN2(n13228), .Q(n12413) );
  OR2X1 U13273 ( .IN1(n13229), .IN2(n13230), .Q(n13228) );
  AND2X1 U13274 ( .IN1(n8458), .IN2(g7194), .Q(n13230) );
  AND2X1 U13275 ( .IN1(n8456), .IN2(n12379), .Q(n13229) );
  AND2X1 U13276 ( .IN1(n8457), .IN2(g1930), .Q(n13227) );
  AND2X1 U13277 ( .IN1(g3229), .IN2(n12425), .Q(n13213) );
  OR2X1 U13278 ( .IN1(n13231), .IN2(n13232), .Q(n12425) );
  OR2X1 U13279 ( .IN1(n13233), .IN2(n13234), .Q(n13232) );
  AND2X1 U13280 ( .IN1(n8468), .IN2(g7194), .Q(n13234) );
  AND2X1 U13281 ( .IN1(n12379), .IN2(n9125), .Q(n13233) );
  AND2X1 U13282 ( .IN1(n8467), .IN2(g1930), .Q(n13231) );
  INVX0 U13283 ( .INP(n13235), .ZN(n13210) );
  OR2X1 U13284 ( .IN1(n12993), .IN2(n8444), .Q(n13235) );
  AND2X1 U13285 ( .IN1(g22651), .IN2(g7052), .Q(n12993) );
  OR2X1 U13286 ( .IN1(n13236), .IN2(n13237), .Q(g27289) );
  AND2X1 U13287 ( .IN1(n13147), .IN2(n13065), .Q(n13237) );
  AND2X1 U13288 ( .IN1(n13238), .IN2(n13239), .Q(n13065) );
  INVX0 U13289 ( .INP(n13240), .ZN(n13239) );
  AND2X1 U13290 ( .IN1(n13241), .IN2(n13242), .Q(n13240) );
  AND2X1 U13291 ( .IN1(n13243), .IN2(n13151), .Q(n13241) );
  OR2X1 U13292 ( .IN1(n13151), .IN2(n13242), .Q(n13238) );
  INVX0 U13293 ( .INP(n13244), .ZN(n13236) );
  OR2X1 U13294 ( .IN1(n13147), .IN2(n8489), .Q(n13244) );
  OR2X1 U13295 ( .IN1(n13245), .IN2(n13246), .Q(g27288) );
  AND2X1 U13296 ( .IN1(n13158), .IN2(n13061), .Q(n13246) );
  INVX0 U13297 ( .INP(n13247), .ZN(n13245) );
  OR2X1 U13298 ( .IN1(n13061), .IN2(n8743), .Q(n13247) );
  OR2X1 U13299 ( .IN1(n13248), .IN2(n13249), .Q(g27287) );
  AND2X1 U13300 ( .IN1(n13250), .IN2(n13006), .Q(n13249) );
  INVX0 U13301 ( .INP(n13251), .ZN(n13248) );
  OR2X1 U13302 ( .IN1(n13006), .IN2(n8765), .Q(n13251) );
  AND2X1 U13303 ( .IN1(n10403), .IN2(n13252), .Q(n13006) );
  OR2X1 U13304 ( .IN1(n13253), .IN2(n13254), .Q(g27286) );
  AND2X1 U13305 ( .IN1(n13078), .IN2(n13069), .Q(n13254) );
  AND2X1 U13306 ( .IN1(n13255), .IN2(n13256), .Q(n13078) );
  OR2X1 U13307 ( .IN1(n13165), .IN2(n12538), .Q(n13255) );
  INVX0 U13308 ( .INP(n12567), .ZN(n12538) );
  XNOR2X1 U13309 ( .IN1(g3229), .IN2(n12561), .Q(n13165) );
  INVX0 U13310 ( .INP(n12548), .ZN(n12561) );
  INVX0 U13311 ( .INP(n13257), .ZN(n13253) );
  OR2X1 U13312 ( .IN1(n13069), .IN2(n8459), .Q(n13257) );
  OR2X1 U13313 ( .IN1(n13258), .IN2(n13259), .Q(g27285) );
  AND2X1 U13314 ( .IN1(n13172), .IN2(n13011), .Q(n13259) );
  INVX0 U13315 ( .INP(n13260), .ZN(n13258) );
  OR2X1 U13316 ( .IN1(n13011), .IN2(n8449), .Q(n13260) );
  AND2X1 U13317 ( .IN1(g6944), .IN2(g22615), .Q(n13011) );
  OR2X1 U13318 ( .IN1(n13261), .IN2(n13262), .Q(g27284) );
  INVX0 U13319 ( .INP(n13263), .ZN(n13262) );
  OR2X1 U13320 ( .IN1(n13264), .IN2(n8758), .Q(n13263) );
  AND2X1 U13321 ( .IN1(n13264), .IN2(n13083), .Q(n13261) );
  OR2X1 U13322 ( .IN1(n13265), .IN2(n13266), .Q(n13083) );
  OR2X1 U13323 ( .IN1(n13267), .IN2(n13268), .Q(n13266) );
  OR2X1 U13324 ( .IN1(n13269), .IN2(n13270), .Q(g27283) );
  AND2X1 U13325 ( .IN1(n13176), .IN2(n13180), .Q(n13270) );
  INVX0 U13326 ( .INP(n13271), .ZN(n13269) );
  OR2X1 U13327 ( .IN1(n13176), .IN2(n8492), .Q(n13271) );
  OR2X1 U13328 ( .IN1(n13272), .IN2(n13273), .Q(g27282) );
  AND2X1 U13329 ( .IN1(n13274), .IN2(n13082), .Q(n13273) );
  INVX0 U13330 ( .INP(n13275), .ZN(n13272) );
  OR2X1 U13331 ( .IN1(n13082), .IN2(n8745), .Q(n13275) );
  OR2X1 U13332 ( .IN1(n13276), .IN2(n13277), .Q(g27281) );
  AND2X1 U13333 ( .IN1(n13184), .IN2(n13091), .Q(n13277) );
  AND2X1 U13334 ( .IN1(n13278), .IN2(n13279), .Q(n13091) );
  OR2X1 U13335 ( .IN1(n13185), .IN2(n12666), .Q(n13279) );
  INVX0 U13336 ( .INP(n13280), .ZN(n13278) );
  AND2X1 U13337 ( .IN1(n12705), .IN2(n13185), .Q(n13280) );
  INVX0 U13338 ( .INP(n13281), .ZN(n13185) );
  AND2X1 U13339 ( .IN1(n12683), .IN2(n12666), .Q(n12705) );
  INVX0 U13340 ( .INP(n13282), .ZN(n13276) );
  OR2X1 U13341 ( .IN1(n13184), .IN2(n8294), .Q(n13282) );
  OR2X1 U13342 ( .IN1(n13283), .IN2(n13284), .Q(g27280) );
  AND2X1 U13343 ( .IN1(n13193), .IN2(n13087), .Q(n13284) );
  AND2X1 U13344 ( .IN1(test_so25), .IN2(n13285), .Q(n13283) );
  INVX0 U13345 ( .INP(n13087), .ZN(n13285) );
  OR2X1 U13346 ( .IN1(n13286), .IN2(n13287), .Q(g27279) );
  AND2X1 U13347 ( .IN1(n13288), .IN2(n13019), .Q(n13287) );
  INVX0 U13348 ( .INP(n13289), .ZN(n13286) );
  OR2X1 U13349 ( .IN1(n13019), .IN2(n8451), .Q(n13289) );
  AND2X1 U13350 ( .IN1(g550), .IN2(g22578), .Q(n13019) );
  OR2X1 U13351 ( .IN1(n13290), .IN2(n13291), .Q(g27278) );
  AND2X1 U13352 ( .IN1(n13292), .IN2(n13198), .Q(n13291) );
  INVX0 U13353 ( .INP(n13293), .ZN(n13290) );
  OR2X1 U13354 ( .IN1(n13292), .IN2(n8760), .Q(n13293) );
  OR2X1 U13355 ( .IN1(n13294), .IN2(n13295), .Q(g27277) );
  AND2X1 U13356 ( .IN1(n13197), .IN2(n13296), .Q(n13295) );
  INVX0 U13357 ( .INP(n13297), .ZN(n13294) );
  OR2X1 U13358 ( .IN1(n13197), .IN2(n8495), .Q(n13297) );
  OR2X1 U13359 ( .IN1(n13298), .IN2(n13299), .Q(g27276) );
  AND2X1 U13360 ( .IN1(n13134), .IN2(n13032), .Q(n13299) );
  INVX0 U13361 ( .INP(n13300), .ZN(n13134) );
  OR2X1 U13362 ( .IN1(n13301), .IN2(n13302), .Q(n13300) );
  OR2X1 U13363 ( .IN1(n13303), .IN2(n13304), .Q(n13302) );
  AND2X1 U13364 ( .IN1(n13305), .IN2(n13306), .Q(n13304) );
  AND2X1 U13365 ( .IN1(n13307), .IN2(n13205), .Q(n13305) );
  OR2X1 U13366 ( .IN1(n13308), .IN2(n13309), .Q(n13205) );
  OR2X1 U13367 ( .IN1(n13310), .IN2(n13311), .Q(n13309) );
  AND2X1 U13368 ( .IN1(n8764), .IN2(n10408), .Q(n13311) );
  AND2X1 U13369 ( .IN1(n8762), .IN2(n10833), .Q(n13310) );
  AND2X1 U13370 ( .IN1(n8763), .IN2(n10398), .Q(n13308) );
  INVX0 U13371 ( .INP(n13125), .ZN(n13307) );
  AND2X1 U13372 ( .IN1(n13204), .IN2(n10061), .Q(n13303) );
  INVX0 U13373 ( .INP(n13306), .ZN(n13204) );
  OR2X1 U13374 ( .IN1(n13127), .IN2(n13035), .Q(n13306) );
  OR2X1 U13375 ( .IN1(n13312), .IN2(n13313), .Q(n13035) );
  OR2X1 U13376 ( .IN1(n13314), .IN2(n13315), .Q(n13313) );
  AND2X1 U13377 ( .IN1(n8486), .IN2(n10408), .Q(n13315) );
  AND2X1 U13378 ( .IN1(n8487), .IN2(n10833), .Q(n13314) );
  AND2X1 U13379 ( .IN1(n8488), .IN2(n10398), .Q(n13312) );
  INVX0 U13380 ( .INP(n13033), .ZN(n13127) );
  OR2X1 U13381 ( .IN1(n13316), .IN2(n13317), .Q(n13033) );
  OR2X1 U13382 ( .IN1(n13318), .IN2(n13319), .Q(n13317) );
  AND2X1 U13383 ( .IN1(n8741), .IN2(n10408), .Q(n13319) );
  AND2X1 U13384 ( .IN1(n8739), .IN2(n10833), .Q(n13318) );
  AND2X1 U13385 ( .IN1(n8740), .IN2(n10398), .Q(n13316) );
  AND2X1 U13386 ( .IN1(g3229), .IN2(n13125), .Q(n13301) );
  OR2X1 U13387 ( .IN1(n13320), .IN2(n13321), .Q(n13125) );
  OR2X1 U13388 ( .IN1(n13322), .IN2(n13323), .Q(n13321) );
  AND2X1 U13389 ( .IN1(n8753), .IN2(n10408), .Q(n13323) );
  AND2X1 U13390 ( .IN1(n8751), .IN2(n10833), .Q(n13322) );
  AND2X1 U13391 ( .IN1(n8752), .IN2(n10398), .Q(n13320) );
  INVX0 U13392 ( .INP(n13324), .ZN(n13298) );
  OR2X1 U13393 ( .IN1(n13032), .IN2(n8764), .Q(n13324) );
  AND2X1 U13394 ( .IN1(g5555), .IN2(n13136), .Q(n13032) );
  INVX0 U13395 ( .INP(n13325), .ZN(n13136) );
  OR2X1 U13396 ( .IN1(n13326), .IN2(n9657), .Q(n13325) );
  AND2X1 U13397 ( .IN1(n9552), .IN2(n9659), .Q(n13326) );
  OR2X1 U13398 ( .IN1(n13327), .IN2(n13328), .Q(g27275) );
  AND2X1 U13399 ( .IN1(n13158), .IN2(n13147), .Q(n13328) );
  AND2X1 U13400 ( .IN1(n13329), .IN2(n13330), .Q(n13158) );
  INVX0 U13401 ( .INP(n13331), .ZN(n13329) );
  AND2X1 U13402 ( .IN1(n13151), .IN2(n13150), .Q(n13331) );
  XNOR2X1 U13403 ( .IN1(g3229), .IN2(n13332), .Q(n13151) );
  INVX0 U13404 ( .INP(n13333), .ZN(n13327) );
  OR2X1 U13405 ( .IN1(n13147), .IN2(n8744), .Q(n13333) );
  OR2X1 U13406 ( .IN1(n13334), .IN2(n13335), .Q(g27274) );
  AND2X1 U13407 ( .IN1(n13250), .IN2(n13061), .Q(n13335) );
  INVX0 U13408 ( .INP(n13336), .ZN(n13334) );
  OR2X1 U13409 ( .IN1(n13061), .IN2(n8766), .Q(n13336) );
  AND2X1 U13410 ( .IN1(g7014), .IN2(n13252), .Q(n13061) );
  OR2X1 U13411 ( .IN1(n13337), .IN2(n13338), .Q(g27273) );
  AND2X1 U13412 ( .IN1(n13172), .IN2(n13069), .Q(n13338) );
  INVX0 U13413 ( .INP(n13339), .ZN(n13172) );
  OR2X1 U13414 ( .IN1(n13340), .IN2(n13341), .Q(n13339) );
  OR2X1 U13415 ( .IN1(n13342), .IN2(n13343), .Q(n13341) );
  AND2X1 U13416 ( .IN1(n13344), .IN2(n13256), .Q(n13343) );
  AND2X1 U13417 ( .IN1(n12568), .IN2(n12548), .Q(n13344) );
  OR2X1 U13418 ( .IN1(n13345), .IN2(n13346), .Q(n12548) );
  OR2X1 U13419 ( .IN1(n13347), .IN2(n13348), .Q(n13346) );
  AND2X1 U13420 ( .IN1(n8449), .IN2(g6944), .Q(n13348) );
  AND2X1 U13421 ( .IN1(n8448), .IN2(g1236), .Q(n13347) );
  AND2X1 U13422 ( .IN1(n8447), .IN2(n12249), .Q(n13345) );
  INVX0 U13423 ( .INP(n12545), .ZN(n12568) );
  INVX0 U13424 ( .INP(n13349), .ZN(n13342) );
  OR2X1 U13425 ( .IN1(n13256), .IN2(g3229), .Q(n13349) );
  OR2X1 U13426 ( .IN1(n12551), .IN2(n12567), .Q(n13256) );
  OR2X1 U13427 ( .IN1(n13350), .IN2(n13351), .Q(n12567) );
  OR2X1 U13428 ( .IN1(n13352), .IN2(n13353), .Q(n13351) );
  AND2X1 U13429 ( .IN1(n8293), .IN2(g6944), .Q(n13353) );
  INVX0 U13430 ( .INP(n13354), .ZN(n13352) );
  OR2X1 U13431 ( .IN1(n4300), .IN2(test_so46), .Q(n13354) );
  AND2X1 U13432 ( .IN1(n8292), .IN2(n12249), .Q(n13350) );
  INVX0 U13433 ( .INP(n12533), .ZN(n12551) );
  OR2X1 U13434 ( .IN1(n13355), .IN2(n13356), .Q(n12533) );
  OR2X1 U13435 ( .IN1(n13357), .IN2(n13358), .Q(n13356) );
  AND2X1 U13436 ( .IN1(n8461), .IN2(g6944), .Q(n13358) );
  AND2X1 U13437 ( .IN1(n8460), .IN2(g1236), .Q(n13357) );
  AND2X1 U13438 ( .IN1(n8459), .IN2(n12249), .Q(n13355) );
  AND2X1 U13439 ( .IN1(g3229), .IN2(n12545), .Q(n13340) );
  OR2X1 U13440 ( .IN1(n13359), .IN2(n13360), .Q(n12545) );
  OR2X1 U13441 ( .IN1(n13361), .IN2(n13362), .Q(n13360) );
  AND2X1 U13442 ( .IN1(n8471), .IN2(g6944), .Q(n13362) );
  AND2X1 U13443 ( .IN1(n8470), .IN2(g1236), .Q(n13361) );
  AND2X1 U13444 ( .IN1(n8469), .IN2(n12249), .Q(n13359) );
  INVX0 U13445 ( .INP(n13363), .ZN(n13337) );
  OR2X1 U13446 ( .IN1(n13069), .IN2(n8447), .Q(n13363) );
  AND2X1 U13447 ( .IN1(g22615), .IN2(g6750), .Q(n13069) );
  OR2X1 U13448 ( .IN1(n13364), .IN2(n13365), .Q(g27272) );
  AND2X1 U13449 ( .IN1(n13264), .IN2(n13180), .Q(n13365) );
  AND2X1 U13450 ( .IN1(n13366), .IN2(n13367), .Q(n13180) );
  OR2X1 U13451 ( .IN1(n13368), .IN2(n13265), .Q(n13367) );
  OR2X1 U13452 ( .IN1(n13369), .IN2(n13370), .Q(n13368) );
  OR2X1 U13453 ( .IN1(n13268), .IN2(n13371), .Q(n13366) );
  AND2X1 U13454 ( .IN1(test_so37), .IN2(n13372), .Q(n13364) );
  OR2X1 U13455 ( .IN1(n13373), .IN2(n13374), .Q(g27271) );
  AND2X1 U13456 ( .IN1(n13274), .IN2(n13176), .Q(n13374) );
  INVX0 U13457 ( .INP(n13375), .ZN(n13373) );
  OR2X1 U13458 ( .IN1(n13176), .IN2(n8746), .Q(n13375) );
  OR2X1 U13459 ( .IN1(n13376), .IN2(n13377), .Q(g27270) );
  AND2X1 U13460 ( .IN1(n13378), .IN2(n13082), .Q(n13377) );
  INVX0 U13461 ( .INP(n13379), .ZN(n13376) );
  OR2X1 U13462 ( .IN1(n13082), .IN2(n8768), .Q(n13379) );
  AND2X1 U13463 ( .IN1(g1088), .IN2(n13380), .Q(n13082) );
  OR2X1 U13464 ( .IN1(n13381), .IN2(n13382), .Q(g27269) );
  AND2X1 U13465 ( .IN1(n13193), .IN2(n13184), .Q(n13382) );
  AND2X1 U13466 ( .IN1(n13383), .IN2(n13384), .Q(n13193) );
  OR2X1 U13467 ( .IN1(n13281), .IN2(n12653), .Q(n13383) );
  INVX0 U13468 ( .INP(n12682), .ZN(n12653) );
  XNOR2X1 U13469 ( .IN1(g3229), .IN2(n12676), .Q(n13281) );
  INVX0 U13470 ( .INP(n12663), .ZN(n12676) );
  INVX0 U13471 ( .INP(n13385), .ZN(n13381) );
  OR2X1 U13472 ( .IN1(n13184), .IN2(n8462), .Q(n13385) );
  OR2X1 U13473 ( .IN1(n13386), .IN2(n13387), .Q(g27268) );
  AND2X1 U13474 ( .IN1(n13288), .IN2(n13087), .Q(n13387) );
  INVX0 U13475 ( .INP(n13388), .ZN(n13386) );
  OR2X1 U13476 ( .IN1(n13087), .IN2(n8452), .Q(n13388) );
  AND2X1 U13477 ( .IN1(g6642), .IN2(g22578), .Q(n13087) );
  OR2X1 U13478 ( .IN1(n13389), .IN2(n13390), .Q(g27267) );
  AND2X1 U13479 ( .IN1(n13391), .IN2(n13198), .Q(n13390) );
  OR2X1 U13480 ( .IN1(n13392), .IN2(n13393), .Q(n13198) );
  OR2X1 U13481 ( .IN1(n13394), .IN2(n13395), .Q(n13393) );
  INVX0 U13482 ( .INP(n13396), .ZN(n13389) );
  OR2X1 U13483 ( .IN1(n13391), .IN2(n8761), .Q(n13396) );
  OR2X1 U13484 ( .IN1(n13397), .IN2(n13398), .Q(g27266) );
  AND2X1 U13485 ( .IN1(n13292), .IN2(n13296), .Q(n13398) );
  INVX0 U13486 ( .INP(n13399), .ZN(n13397) );
  OR2X1 U13487 ( .IN1(n13292), .IN2(n8496), .Q(n13399) );
  OR2X1 U13488 ( .IN1(n13400), .IN2(n13401), .Q(g27265) );
  AND2X1 U13489 ( .IN1(n13402), .IN2(n13197), .Q(n13401) );
  INVX0 U13490 ( .INP(n13403), .ZN(n13400) );
  OR2X1 U13491 ( .IN1(n13197), .IN2(n8748), .Q(n13403) );
  OR2X1 U13492 ( .IN1(n13404), .IN2(n13405), .Q(g27264) );
  AND2X1 U13493 ( .IN1(n13250), .IN2(n13147), .Q(n13405) );
  AND2X1 U13494 ( .IN1(n13406), .IN2(n13407), .Q(n13250) );
  AND2X1 U13495 ( .IN1(n13408), .IN2(n13409), .Q(n13407) );
  INVX0 U13496 ( .INP(n13410), .ZN(n13409) );
  AND2X1 U13497 ( .IN1(n13411), .IN2(n13330), .Q(n13410) );
  AND2X1 U13498 ( .IN1(n13243), .IN2(n13332), .Q(n13411) );
  OR2X1 U13499 ( .IN1(n13412), .IN2(n13413), .Q(n13332) );
  OR2X1 U13500 ( .IN1(n13414), .IN2(n13415), .Q(n13413) );
  AND2X1 U13501 ( .IN1(n8767), .IN2(n10419), .Q(n13415) );
  AND2X1 U13502 ( .IN1(n8765), .IN2(n10403), .Q(n13414) );
  AND2X1 U13503 ( .IN1(n8766), .IN2(n10412), .Q(n13412) );
  OR2X1 U13504 ( .IN1(n13330), .IN2(g3229), .Q(n13408) );
  OR2X1 U13505 ( .IN1(n13242), .IN2(n13150), .Q(n13330) );
  OR2X1 U13506 ( .IN1(n13416), .IN2(n13417), .Q(n13150) );
  OR2X1 U13507 ( .IN1(n13418), .IN2(n13419), .Q(n13417) );
  AND2X1 U13508 ( .IN1(n8489), .IN2(n10419), .Q(n13419) );
  AND2X1 U13509 ( .IN1(n8490), .IN2(n10403), .Q(n13418) );
  AND2X1 U13510 ( .IN1(n8491), .IN2(n10412), .Q(n13416) );
  INVX0 U13511 ( .INP(n13148), .ZN(n13242) );
  OR2X1 U13512 ( .IN1(n13420), .IN2(n13421), .Q(n13148) );
  OR2X1 U13513 ( .IN1(n13422), .IN2(n13423), .Q(n13421) );
  AND2X1 U13514 ( .IN1(n8744), .IN2(n10419), .Q(n13423) );
  AND2X1 U13515 ( .IN1(n8742), .IN2(n10403), .Q(n13422) );
  AND2X1 U13516 ( .IN1(n8743), .IN2(n10412), .Q(n13420) );
  OR2X1 U13517 ( .IN1(n10061), .IN2(n13243), .Q(n13406) );
  AND2X1 U13518 ( .IN1(n13424), .IN2(n13425), .Q(n13243) );
  INVX0 U13519 ( .INP(n13426), .ZN(n13425) );
  OR2X1 U13520 ( .IN1(n13427), .IN2(n13428), .Q(n13426) );
  AND2X1 U13521 ( .IN1(n8755), .IN2(n10419), .Q(n13428) );
  AND2X1 U13522 ( .IN1(n8754), .IN2(n10403), .Q(n13427) );
  OR2X1 U13523 ( .IN1(n4525), .IN2(test_so58), .Q(n13424) );
  INVX0 U13524 ( .INP(n13429), .ZN(n13404) );
  OR2X1 U13525 ( .IN1(n13147), .IN2(n8767), .Q(n13429) );
  AND2X1 U13526 ( .IN1(g5511), .IN2(n13252), .Q(n13147) );
  INVX0 U13527 ( .INP(n13430), .ZN(n13252) );
  OR2X1 U13528 ( .IN1(n13431), .IN2(n9622), .Q(n13430) );
  AND2X1 U13529 ( .IN1(n9552), .IN2(n9625), .Q(n13431) );
  OR2X1 U13530 ( .IN1(n13432), .IN2(n13433), .Q(g27263) );
  AND2X1 U13531 ( .IN1(n13274), .IN2(n13264), .Q(n13433) );
  INVX0 U13532 ( .INP(n13434), .ZN(n13274) );
  OR2X1 U13533 ( .IN1(n13435), .IN2(n13436), .Q(n13434) );
  AND2X1 U13534 ( .IN1(n13268), .IN2(n13267), .Q(n13435) );
  INVX0 U13535 ( .INP(n13370), .ZN(n13268) );
  XOR2X1 U13536 ( .IN1(g3229), .IN2(n13437), .Q(n13370) );
  INVX0 U13537 ( .INP(n13438), .ZN(n13432) );
  OR2X1 U13538 ( .IN1(n13264), .IN2(n8747), .Q(n13438) );
  OR2X1 U13539 ( .IN1(n13439), .IN2(n13440), .Q(g27262) );
  AND2X1 U13540 ( .IN1(n13378), .IN2(n13176), .Q(n13440) );
  INVX0 U13541 ( .INP(n13441), .ZN(n13439) );
  OR2X1 U13542 ( .IN1(n13176), .IN2(n8769), .Q(n13441) );
  AND2X1 U13543 ( .IN1(g6712), .IN2(n13380), .Q(n13176) );
  INVX0 U13544 ( .INP(n13442), .ZN(n13380) );
  OR2X1 U13545 ( .IN1(n13443), .IN2(n13444), .Q(g27261) );
  AND2X1 U13546 ( .IN1(n13288), .IN2(n13184), .Q(n13444) );
  INVX0 U13547 ( .INP(n13445), .ZN(n13288) );
  OR2X1 U13548 ( .IN1(n13446), .IN2(n13447), .Q(n13445) );
  OR2X1 U13549 ( .IN1(n13448), .IN2(n13449), .Q(n13447) );
  AND2X1 U13550 ( .IN1(n13450), .IN2(n13384), .Q(n13449) );
  AND2X1 U13551 ( .IN1(n12683), .IN2(n12663), .Q(n13450) );
  OR2X1 U13552 ( .IN1(n13451), .IN2(n13452), .Q(n12663) );
  OR2X1 U13553 ( .IN1(n13453), .IN2(n13454), .Q(n13452) );
  AND2X1 U13554 ( .IN1(n8451), .IN2(g550), .Q(n13454) );
  AND2X1 U13555 ( .IN1(n8450), .IN2(n9810), .Q(n13453) );
  AND2X1 U13556 ( .IN1(n8452), .IN2(g6642), .Q(n13451) );
  INVX0 U13557 ( .INP(n12660), .ZN(n12683) );
  INVX0 U13558 ( .INP(n13455), .ZN(n13448) );
  OR2X1 U13559 ( .IN1(n13384), .IN2(g3229), .Q(n13455) );
  OR2X1 U13560 ( .IN1(n12666), .IN2(n12682), .Q(n13384) );
  OR2X1 U13561 ( .IN1(n13456), .IN2(n13457), .Q(n12682) );
  OR2X1 U13562 ( .IN1(n13458), .IN2(n13459), .Q(n13457) );
  AND2X1 U13563 ( .IN1(n8295), .IN2(g550), .Q(n13459) );
  AND2X1 U13564 ( .IN1(n8294), .IN2(n9810), .Q(n13458) );
  AND2X1 U13565 ( .IN1(n8296), .IN2(g6642), .Q(n13456) );
  INVX0 U13566 ( .INP(n12648), .ZN(n12666) );
  OR2X1 U13567 ( .IN1(n13460), .IN2(n13461), .Q(n12648) );
  OR2X1 U13568 ( .IN1(n13462), .IN2(n13463), .Q(n13461) );
  AND2X1 U13569 ( .IN1(n8463), .IN2(g550), .Q(n13463) );
  AND2X1 U13570 ( .IN1(n8462), .IN2(n9810), .Q(n13462) );
  INVX0 U13571 ( .INP(n13464), .ZN(n13460) );
  OR2X1 U13572 ( .IN1(n4372), .IN2(test_so25), .Q(n13464) );
  AND2X1 U13573 ( .IN1(g3229), .IN2(n12660), .Q(n13446) );
  OR2X1 U13574 ( .IN1(n13465), .IN2(n13466), .Q(n12660) );
  OR2X1 U13575 ( .IN1(n13467), .IN2(n13468), .Q(n13466) );
  AND2X1 U13576 ( .IN1(n8473), .IN2(g550), .Q(n13468) );
  AND2X1 U13577 ( .IN1(n8472), .IN2(n9810), .Q(n13467) );
  AND2X1 U13578 ( .IN1(n8474), .IN2(g6642), .Q(n13465) );
  INVX0 U13579 ( .INP(n13469), .ZN(n13443) );
  OR2X1 U13580 ( .IN1(n13184), .IN2(n8450), .Q(n13469) );
  AND2X1 U13581 ( .IN1(g22578), .IN2(g6485), .Q(n13184) );
  OR2X1 U13582 ( .IN1(n13470), .IN2(n13471), .Q(g27260) );
  AND2X1 U13583 ( .IN1(n13391), .IN2(n13296), .Q(n13471) );
  AND2X1 U13584 ( .IN1(n13472), .IN2(n13473), .Q(n13296) );
  OR2X1 U13585 ( .IN1(n13474), .IN2(n13392), .Q(n13473) );
  OR2X1 U13586 ( .IN1(n13475), .IN2(n13476), .Q(n13474) );
  OR2X1 U13587 ( .IN1(n13395), .IN2(n13477), .Q(n13472) );
  INVX0 U13588 ( .INP(n13478), .ZN(n13470) );
  OR2X1 U13589 ( .IN1(n13391), .IN2(n8494), .Q(n13478) );
  OR2X1 U13590 ( .IN1(n13479), .IN2(n13480), .Q(g27259) );
  AND2X1 U13591 ( .IN1(n13402), .IN2(n13292), .Q(n13480) );
  INVX0 U13592 ( .INP(n13481), .ZN(n13479) );
  OR2X1 U13593 ( .IN1(n13292), .IN2(n8749), .Q(n13481) );
  OR2X1 U13594 ( .IN1(n13482), .IN2(n13483), .Q(g27258) );
  AND2X1 U13595 ( .IN1(n13484), .IN2(n13197), .Q(n13483) );
  INVX0 U13596 ( .INP(n13485), .ZN(n13197) );
  AND2X1 U13597 ( .IN1(test_so16), .IN2(n13485), .Q(n13482) );
  OR2X1 U13598 ( .IN1(n4506), .IN2(n13486), .Q(n13485) );
  OR2X1 U13599 ( .IN1(n13487), .IN2(n13488), .Q(g27257) );
  AND2X1 U13600 ( .IN1(n13378), .IN2(n13264), .Q(n13488) );
  INVX0 U13601 ( .INP(n13489), .ZN(n13378) );
  OR2X1 U13602 ( .IN1(n13490), .IN2(n13491), .Q(n13489) );
  OR2X1 U13603 ( .IN1(n13492), .IN2(n13493), .Q(n13491) );
  AND2X1 U13604 ( .IN1(n13494), .IN2(n13495), .Q(n13493) );
  AND2X1 U13605 ( .IN1(n13496), .IN2(n13437), .Q(n13494) );
  OR2X1 U13606 ( .IN1(n13497), .IN2(n13498), .Q(n13437) );
  OR2X1 U13607 ( .IN1(n13499), .IN2(n13500), .Q(n13498) );
  AND2X1 U13608 ( .IN1(n8769), .IN2(g6712), .Q(n13500) );
  AND2X1 U13609 ( .IN1(n8770), .IN2(g5472), .Q(n13499) );
  AND2X1 U13610 ( .IN1(n8768), .IN2(g1088), .Q(n13497) );
  INVX0 U13611 ( .INP(n13369), .ZN(n13496) );
  AND2X1 U13612 ( .IN1(n13436), .IN2(n10061), .Q(n13492) );
  INVX0 U13613 ( .INP(n13495), .ZN(n13436) );
  OR2X1 U13614 ( .IN1(n13371), .IN2(n13267), .Q(n13495) );
  OR2X1 U13615 ( .IN1(n13501), .IN2(n13502), .Q(n13267) );
  OR2X1 U13616 ( .IN1(n13503), .IN2(n13504), .Q(n13502) );
  AND2X1 U13617 ( .IN1(n8492), .IN2(g6712), .Q(n13504) );
  INVX0 U13618 ( .INP(n13505), .ZN(n13503) );
  OR2X1 U13619 ( .IN1(n4363), .IN2(test_so37), .Q(n13505) );
  AND2X1 U13620 ( .IN1(n8493), .IN2(g1088), .Q(n13501) );
  INVX0 U13621 ( .INP(n13265), .ZN(n13371) );
  OR2X1 U13622 ( .IN1(n13506), .IN2(n13507), .Q(n13265) );
  OR2X1 U13623 ( .IN1(n13508), .IN2(n13509), .Q(n13507) );
  AND2X1 U13624 ( .IN1(n8746), .IN2(g6712), .Q(n13509) );
  AND2X1 U13625 ( .IN1(n8747), .IN2(g5472), .Q(n13508) );
  AND2X1 U13626 ( .IN1(n8745), .IN2(g1088), .Q(n13506) );
  AND2X1 U13627 ( .IN1(g3229), .IN2(n13369), .Q(n13490) );
  OR2X1 U13628 ( .IN1(n13510), .IN2(n13511), .Q(n13369) );
  OR2X1 U13629 ( .IN1(n13512), .IN2(n13513), .Q(n13511) );
  AND2X1 U13630 ( .IN1(n8757), .IN2(g6712), .Q(n13513) );
  AND2X1 U13631 ( .IN1(n8758), .IN2(g5472), .Q(n13512) );
  AND2X1 U13632 ( .IN1(n8756), .IN2(g1088), .Q(n13510) );
  INVX0 U13633 ( .INP(n13514), .ZN(n13487) );
  OR2X1 U13634 ( .IN1(n13264), .IN2(n8770), .Q(n13514) );
  INVX0 U13635 ( .INP(n13372), .ZN(n13264) );
  OR2X1 U13636 ( .IN1(n4363), .IN2(n13442), .Q(n13372) );
  OR2X1 U13637 ( .IN1(n13515), .IN2(n9588), .Q(n13442) );
  AND2X1 U13638 ( .IN1(n9552), .IN2(n9590), .Q(n13515) );
  OR2X1 U13639 ( .IN1(n13516), .IN2(n13517), .Q(g27256) );
  AND2X1 U13640 ( .IN1(n13402), .IN2(n13391), .Q(n13517) );
  INVX0 U13641 ( .INP(n13518), .ZN(n13402) );
  OR2X1 U13642 ( .IN1(n13519), .IN2(n13520), .Q(n13518) );
  AND2X1 U13643 ( .IN1(n13395), .IN2(n13394), .Q(n13519) );
  INVX0 U13644 ( .INP(n13476), .ZN(n13395) );
  XOR2X1 U13645 ( .IN1(g3229), .IN2(n13521), .Q(n13476) );
  INVX0 U13646 ( .INP(n13522), .ZN(n13516) );
  OR2X1 U13647 ( .IN1(n13391), .IN2(n8750), .Q(n13522) );
  OR2X1 U13648 ( .IN1(n13523), .IN2(n13524), .Q(g27255) );
  AND2X1 U13649 ( .IN1(n13484), .IN2(n13292), .Q(n13524) );
  INVX0 U13650 ( .INP(n13525), .ZN(n13523) );
  OR2X1 U13651 ( .IN1(n13292), .IN2(n8771), .Q(n13525) );
  AND2X1 U13652 ( .IN1(g6447), .IN2(n13526), .Q(n13292) );
  OR2X1 U13653 ( .IN1(n13527), .IN2(n13528), .Q(g27253) );
  AND2X1 U13654 ( .IN1(n13484), .IN2(n13391), .Q(n13528) );
  INVX0 U13655 ( .INP(n13529), .ZN(n13484) );
  OR2X1 U13656 ( .IN1(n13530), .IN2(n13531), .Q(n13529) );
  OR2X1 U13657 ( .IN1(n13532), .IN2(n13533), .Q(n13531) );
  AND2X1 U13658 ( .IN1(n13534), .IN2(n13535), .Q(n13533) );
  AND2X1 U13659 ( .IN1(n13536), .IN2(n13521), .Q(n13534) );
  OR2X1 U13660 ( .IN1(n13537), .IN2(n13538), .Q(n13521) );
  OR2X1 U13661 ( .IN1(n13539), .IN2(n13540), .Q(n13538) );
  INVX0 U13662 ( .INP(n13541), .ZN(n13540) );
  OR2X1 U13663 ( .IN1(n4506), .IN2(test_so16), .Q(n13541) );
  AND2X1 U13664 ( .IN1(n8771), .IN2(n10899), .Q(n13539) );
  AND2X1 U13665 ( .IN1(n8772), .IN2(n10475), .Q(n13537) );
  INVX0 U13666 ( .INP(n13475), .ZN(n13536) );
  AND2X1 U13667 ( .IN1(n13520), .IN2(n10061), .Q(n13532) );
  INVX0 U13668 ( .INP(n13535), .ZN(n13520) );
  OR2X1 U13669 ( .IN1(n13477), .IN2(n13394), .Q(n13535) );
  OR2X1 U13670 ( .IN1(n13542), .IN2(n13543), .Q(n13394) );
  OR2X1 U13671 ( .IN1(n13544), .IN2(n13545), .Q(n13543) );
  AND2X1 U13672 ( .IN1(n8495), .IN2(n10465), .Q(n13545) );
  AND2X1 U13673 ( .IN1(n8496), .IN2(n10899), .Q(n13544) );
  AND2X1 U13674 ( .IN1(n8494), .IN2(n10475), .Q(n13542) );
  INVX0 U13675 ( .INP(n13392), .ZN(n13477) );
  OR2X1 U13676 ( .IN1(n13546), .IN2(n13547), .Q(n13392) );
  OR2X1 U13677 ( .IN1(n13548), .IN2(n13549), .Q(n13547) );
  AND2X1 U13678 ( .IN1(n8748), .IN2(n10465), .Q(n13549) );
  AND2X1 U13679 ( .IN1(n8749), .IN2(n10899), .Q(n13548) );
  AND2X1 U13680 ( .IN1(n8750), .IN2(n10475), .Q(n13546) );
  AND2X1 U13681 ( .IN1(g3229), .IN2(n13475), .Q(n13530) );
  OR2X1 U13682 ( .IN1(n13550), .IN2(n13551), .Q(n13475) );
  OR2X1 U13683 ( .IN1(n13552), .IN2(n13553), .Q(n13551) );
  AND2X1 U13684 ( .IN1(n8759), .IN2(n10465), .Q(n13553) );
  AND2X1 U13685 ( .IN1(n8760), .IN2(n10899), .Q(n13552) );
  AND2X1 U13686 ( .IN1(n8761), .IN2(n10475), .Q(n13550) );
  INVX0 U13687 ( .INP(n13554), .ZN(n13527) );
  OR2X1 U13688 ( .IN1(n13391), .IN2(n8772), .Q(n13554) );
  AND2X1 U13689 ( .IN1(g5437), .IN2(n13526), .Q(n13391) );
  INVX0 U13690 ( .INP(n13486), .ZN(n13526) );
  OR2X1 U13691 ( .IN1(n13555), .IN2(n9553), .Q(n13486) );
  AND2X1 U13692 ( .IN1(n9552), .IN2(n9556), .Q(n13555) );
  AND2X1 U13693 ( .IN1(n13556), .IN2(n13557), .Q(g27243) );
  INVX0 U13694 ( .INP(n13558), .ZN(n13557) );
  AND2X1 U13695 ( .IN1(n13559), .IN2(n4471), .Q(n13558) );
  OR2X1 U13696 ( .IN1(n9122), .IN2(n13560), .Q(n13559) );
  AND2X1 U13697 ( .IN1(n12739), .IN2(n12737), .Q(n13556) );
  OR2X1 U13698 ( .IN1(n9122), .IN2(n13561), .Q(n12739) );
  OR2X1 U13699 ( .IN1(n4471), .IN2(n13560), .Q(n13561) );
  AND2X1 U13700 ( .IN1(n13562), .IN2(n4522), .Q(g27131) );
  AND2X1 U13701 ( .IN1(n13563), .IN2(n11527), .Q(n13562) );
  INVX0 U13702 ( .INP(n13564), .ZN(n13563) );
  AND2X1 U13703 ( .IN1(n10220), .IN2(n9116), .Q(n13564) );
  INVX0 U13704 ( .INP(n3683), .ZN(n10220) );
  AND2X1 U13705 ( .IN1(n13565), .IN2(n4523), .Q(g27129) );
  AND2X1 U13706 ( .IN1(n13566), .IN2(n11529), .Q(n13565) );
  INVX0 U13707 ( .INP(n13567), .ZN(n13566) );
  AND2X1 U13708 ( .IN1(n10219), .IN2(n9115), .Q(n13567) );
  INVX0 U13709 ( .INP(n3686), .ZN(n10219) );
  AND2X1 U13710 ( .IN1(n13568), .IN2(n13569), .Q(g27123) );
  OR2X1 U13711 ( .IN1(n3689), .IN2(g767), .Q(n13569) );
  AND2X1 U13712 ( .IN1(n11531), .IN2(n712), .Q(n13568) );
  INVX0 U13713 ( .INP(n12890), .ZN(n712) );
  AND2X1 U13714 ( .IN1(g767), .IN2(n3689), .Q(n12890) );
  AND2X1 U13715 ( .IN1(n13570), .IN2(n4521), .Q(g27120) );
  AND2X1 U13716 ( .IN1(n13571), .IN2(n11533), .Q(n13570) );
  OR2X1 U13717 ( .IN1(n3692), .IN2(test_so15), .Q(n13571) );
  OR2X1 U13718 ( .IN1(n13572), .IN2(n13573), .Q(g26827) );
  AND2X1 U13719 ( .IN1(n4509), .IN2(g2519), .Q(n13573) );
  AND2X1 U13720 ( .IN1(n13574), .IN2(n4606), .Q(n13572) );
  OR2X1 U13721 ( .IN1(n13575), .IN2(n13576), .Q(g26826) );
  AND2X1 U13722 ( .IN1(n4524), .IN2(g2516), .Q(n13576) );
  AND2X1 U13723 ( .IN1(n13574), .IN2(g7264), .Q(n13575) );
  OR2X1 U13724 ( .IN1(n13577), .IN2(n13578), .Q(g26825) );
  AND2X1 U13725 ( .IN1(n4509), .IN2(g2510), .Q(n13578) );
  AND2X1 U13726 ( .IN1(n4606), .IN2(n13579), .Q(n13577) );
  OR2X1 U13727 ( .IN1(n13580), .IN2(n13581), .Q(g26824) );
  AND2X1 U13728 ( .IN1(test_so59), .IN2(n4511), .Q(n13581) );
  AND2X1 U13729 ( .IN1(n13582), .IN2(n4618), .Q(n13580) );
  OR2X1 U13730 ( .IN1(n13583), .IN2(n13584), .Q(g26823) );
  AND2X1 U13731 ( .IN1(n4516), .IN2(g2513), .Q(n13584) );
  AND2X1 U13732 ( .IN1(n13574), .IN2(g5555), .Q(n13583) );
  XNOR2X1 U13733 ( .IN1(n13585), .IN2(n12782), .Q(n13574) );
  OR2X1 U13734 ( .IN1(n13586), .IN2(n12788), .Q(n13585) );
  OR2X1 U13735 ( .IN1(n9121), .IN2(n13587), .Q(n12788) );
  OR2X1 U13736 ( .IN1(n13588), .IN2(n13589), .Q(n13587) );
  AND2X1 U13737 ( .IN1(n13590), .IN2(n12783), .Q(n13589) );
  OR2X1 U13738 ( .IN1(n12782), .IN2(n12777), .Q(n13590) );
  INVX0 U13739 ( .INP(n12780), .ZN(n12777) );
  AND2X1 U13740 ( .IN1(n12779), .IN2(n13591), .Q(n13588) );
  OR2X1 U13741 ( .IN1(n12780), .IN2(n12778), .Q(n13591) );
  INVX0 U13742 ( .INP(n12782), .ZN(n12778) );
  INVX0 U13743 ( .INP(n12783), .ZN(n12779) );
  AND2X1 U13744 ( .IN1(n13592), .IN2(n12789), .Q(n13586) );
  OR2X1 U13745 ( .IN1(n4509), .IN2(test_so81), .Q(n12789) );
  INVX0 U13746 ( .INP(n12785), .ZN(n13592) );
  OR2X1 U13747 ( .IN1(n13593), .IN2(n13594), .Q(n12785) );
  AND2X1 U13748 ( .IN1(n8774), .IN2(n10398), .Q(n13594) );
  AND2X1 U13749 ( .IN1(n8783), .IN2(n10408), .Q(n13593) );
  OR2X1 U13750 ( .IN1(n13595), .IN2(n13596), .Q(g26822) );
  AND2X1 U13751 ( .IN1(n4524), .IN2(g2507), .Q(n13596) );
  AND2X1 U13752 ( .IN1(g7264), .IN2(n13579), .Q(n13595) );
  OR2X1 U13753 ( .IN1(n13597), .IN2(n13598), .Q(g26821) );
  AND2X1 U13754 ( .IN1(n4525), .IN2(g1822), .Q(n13598) );
  AND2X1 U13755 ( .IN1(n13582), .IN2(g7014), .Q(n13597) );
  OR2X1 U13756 ( .IN1(n13599), .IN2(n13600), .Q(g26820) );
  AND2X1 U13757 ( .IN1(n4511), .IN2(g1816), .Q(n13600) );
  AND2X1 U13758 ( .IN1(n4618), .IN2(n13601), .Q(n13599) );
  OR2X1 U13759 ( .IN1(n13602), .IN2(n13603), .Q(g26818) );
  AND2X1 U13760 ( .IN1(n13604), .IN2(g1088), .Q(n13603) );
  AND2X1 U13761 ( .IN1(n4381), .IN2(g1131), .Q(n13602) );
  OR2X1 U13762 ( .IN1(n13605), .IN2(n13606), .Q(g26817) );
  AND2X1 U13763 ( .IN1(n4516), .IN2(g2504), .Q(n13606) );
  AND2X1 U13764 ( .IN1(g5555), .IN2(n13579), .Q(n13605) );
  OR2X1 U13765 ( .IN1(n13607), .IN2(n13608), .Q(n13579) );
  AND2X1 U13766 ( .IN1(n12783), .IN2(n9121), .Q(n13608) );
  OR2X1 U13767 ( .IN1(n13609), .IN2(n13610), .Q(n12783) );
  OR2X1 U13768 ( .IN1(n13611), .IN2(n13612), .Q(n13610) );
  AND2X1 U13769 ( .IN1(g7264), .IN2(g2507), .Q(n13612) );
  AND2X1 U13770 ( .IN1(n4606), .IN2(g2510), .Q(n13611) );
  AND2X1 U13771 ( .IN1(g5555), .IN2(g2504), .Q(n13609) );
  AND2X1 U13772 ( .IN1(n12780), .IN2(test_so79), .Q(n13607) );
  AND2X1 U13773 ( .IN1(n13613), .IN2(n13614), .Q(n12780) );
  INVX0 U13774 ( .INP(n12102), .ZN(n13614) );
  OR2X1 U13775 ( .IN1(n13615), .IN2(n13616), .Q(n13613) );
  AND2X1 U13776 ( .IN1(test_so73), .IN2(n8686), .Q(n13616) );
  OR2X1 U13777 ( .IN1(n13617), .IN2(n13618), .Q(n13615) );
  AND2X1 U13778 ( .IN1(g6837), .IN2(n8687), .Q(n13618) );
  AND2X1 U13779 ( .IN1(g2241), .IN2(n8685), .Q(n13617) );
  OR2X1 U13780 ( .IN1(n13619), .IN2(n13620), .Q(g26816) );
  AND2X1 U13781 ( .IN1(n4518), .IN2(g1819), .Q(n13620) );
  AND2X1 U13782 ( .IN1(n13582), .IN2(g5511), .Q(n13619) );
  XNOR2X1 U13783 ( .IN1(n13621), .IN2(n12805), .Q(n13582) );
  OR2X1 U13784 ( .IN1(n13622), .IN2(n12816), .Q(n13621) );
  OR2X1 U13785 ( .IN1(n4386), .IN2(n13623), .Q(n12816) );
  OR2X1 U13786 ( .IN1(n13624), .IN2(n13625), .Q(n13623) );
  AND2X1 U13787 ( .IN1(n13626), .IN2(n12811), .Q(n13625) );
  OR2X1 U13788 ( .IN1(n12810), .IN2(n12805), .Q(n13626) );
  AND2X1 U13789 ( .IN1(n12807), .IN2(n13627), .Q(n13624) );
  OR2X1 U13790 ( .IN1(n12808), .IN2(n12806), .Q(n13627) );
  INVX0 U13791 ( .INP(n12805), .ZN(n12808) );
  INVX0 U13792 ( .INP(n12811), .ZN(n12807) );
  AND2X1 U13793 ( .IN1(n13628), .IN2(n13629), .Q(n13622) );
  OR2X1 U13794 ( .IN1(n4525), .IN2(g1830), .Q(n13629) );
  INVX0 U13795 ( .INP(n12813), .ZN(n13628) );
  OR2X1 U13796 ( .IN1(n13630), .IN2(n13631), .Q(n12813) );
  AND2X1 U13797 ( .IN1(n8788), .IN2(n10419), .Q(n13631) );
  AND2X1 U13798 ( .IN1(n8787), .IN2(n10403), .Q(n13630) );
  OR2X1 U13799 ( .IN1(n13632), .IN2(n13633), .Q(g26815) );
  AND2X1 U13800 ( .IN1(n4525), .IN2(g1813), .Q(n13633) );
  AND2X1 U13801 ( .IN1(g7014), .IN2(n13601), .Q(n13632) );
  OR2X1 U13802 ( .IN1(n13634), .IN2(n13635), .Q(g26814) );
  AND2X1 U13803 ( .IN1(n13604), .IN2(g6712), .Q(n13635) );
  AND2X1 U13804 ( .IN1(n4364), .IN2(g1128), .Q(n13634) );
  OR2X1 U13805 ( .IN1(n13636), .IN2(n13637), .Q(g26813) );
  AND2X1 U13806 ( .IN1(n13638), .IN2(g1088), .Q(n13637) );
  AND2X1 U13807 ( .IN1(n4381), .IN2(g1122), .Q(n13636) );
  OR2X1 U13808 ( .IN1(n13639), .IN2(n13640), .Q(g26812) );
  AND2X1 U13809 ( .IN1(n4506), .IN2(g444), .Q(n13640) );
  AND2X1 U13810 ( .IN1(n13641), .IN2(n4640), .Q(n13639) );
  OR2X1 U13811 ( .IN1(n13642), .IN2(n13643), .Q(g26811) );
  AND2X1 U13812 ( .IN1(n4518), .IN2(g1810), .Q(n13643) );
  AND2X1 U13813 ( .IN1(g5511), .IN2(n13601), .Q(n13642) );
  OR2X1 U13814 ( .IN1(n13644), .IN2(n13645), .Q(n13601) );
  AND2X1 U13815 ( .IN1(n4386), .IN2(n12811), .Q(n13645) );
  OR2X1 U13816 ( .IN1(n13646), .IN2(n13647), .Q(n12811) );
  OR2X1 U13817 ( .IN1(n13648), .IN2(n13649), .Q(n13647) );
  AND2X1 U13818 ( .IN1(g7014), .IN2(g1813), .Q(n13649) );
  AND2X1 U13819 ( .IN1(n4618), .IN2(g1816), .Q(n13648) );
  AND2X1 U13820 ( .IN1(g5511), .IN2(g1810), .Q(n13646) );
  AND2X1 U13821 ( .IN1(n12806), .IN2(g1690), .Q(n13644) );
  INVX0 U13822 ( .INP(n12810), .ZN(n12806) );
  OR2X1 U13823 ( .IN1(n13650), .IN2(n12145), .Q(n12810) );
  AND2X1 U13824 ( .IN1(n13651), .IN2(n13652), .Q(n13650) );
  INVX0 U13825 ( .INP(n13653), .ZN(n13652) );
  AND2X1 U13826 ( .IN1(g6573), .IN2(n8699), .Q(n13653) );
  AND2X1 U13827 ( .IN1(n13654), .IN2(n13655), .Q(n13651) );
  INVX0 U13828 ( .INP(n13656), .ZN(n13655) );
  AND2X1 U13829 ( .IN1(g6782), .IN2(n8698), .Q(n13656) );
  OR2X1 U13830 ( .IN1(n4368), .IN2(g1559), .Q(n13654) );
  OR2X1 U13831 ( .IN1(n13657), .IN2(n13658), .Q(g26810) );
  AND2X1 U13832 ( .IN1(n13604), .IN2(g5472), .Q(n13658) );
  XNOR2X1 U13833 ( .IN1(n13659), .IN2(n12832), .Q(n13604) );
  OR2X1 U13834 ( .IN1(n13660), .IN2(n12843), .Q(n13659) );
  OR2X1 U13835 ( .IN1(n4387), .IN2(n13661), .Q(n12843) );
  OR2X1 U13836 ( .IN1(n13662), .IN2(n13663), .Q(n13661) );
  AND2X1 U13837 ( .IN1(n13664), .IN2(n12838), .Q(n13663) );
  OR2X1 U13838 ( .IN1(n12837), .IN2(n12832), .Q(n13664) );
  AND2X1 U13839 ( .IN1(n12834), .IN2(n13665), .Q(n13662) );
  OR2X1 U13840 ( .IN1(n12835), .IN2(n12833), .Q(n13665) );
  INVX0 U13841 ( .INP(n12832), .ZN(n12835) );
  INVX0 U13842 ( .INP(n12838), .ZN(n12834) );
  AND2X1 U13843 ( .IN1(n13666), .IN2(n13667), .Q(n13660) );
  OR2X1 U13844 ( .IN1(n4364), .IN2(g1136), .Q(n13667) );
  INVX0 U13845 ( .INP(n12840), .ZN(n13666) );
  OR2X1 U13846 ( .IN1(n13668), .IN2(n13669), .Q(n12840) );
  AND2X1 U13847 ( .IN1(n8793), .IN2(g1088), .Q(n13669) );
  AND2X1 U13848 ( .IN1(n8794), .IN2(g5472), .Q(n13668) );
  AND2X1 U13849 ( .IN1(n4363), .IN2(g1125), .Q(n13657) );
  OR2X1 U13850 ( .IN1(n13670), .IN2(n13671), .Q(g26809) );
  AND2X1 U13851 ( .IN1(n4364), .IN2(test_so38), .Q(n13671) );
  AND2X1 U13852 ( .IN1(n13638), .IN2(g6712), .Q(n13670) );
  OR2X1 U13853 ( .IN1(n13672), .IN2(n13673), .Q(g26808) );
  AND2X1 U13854 ( .IN1(n4499), .IN2(g441), .Q(n13673) );
  AND2X1 U13855 ( .IN1(n13641), .IN2(g6447), .Q(n13672) );
  OR2X1 U13856 ( .IN1(n13674), .IN2(n13675), .Q(g26807) );
  AND2X1 U13857 ( .IN1(n4506), .IN2(g435), .Q(n13675) );
  AND2X1 U13858 ( .IN1(n4640), .IN2(n13676), .Q(n13674) );
  OR2X1 U13859 ( .IN1(n13677), .IN2(n13678), .Q(g26806) );
  AND2X1 U13860 ( .IN1(n13638), .IN2(g5472), .Q(n13678) );
  OR2X1 U13861 ( .IN1(n13679), .IN2(n13680), .Q(n13638) );
  AND2X1 U13862 ( .IN1(n4387), .IN2(n12838), .Q(n13680) );
  OR2X1 U13863 ( .IN1(n13681), .IN2(n13682), .Q(n12838) );
  OR2X1 U13864 ( .IN1(n13683), .IN2(n13684), .Q(n13682) );
  AND2X1 U13865 ( .IN1(test_so38), .IN2(g6712), .Q(n13684) );
  AND2X1 U13866 ( .IN1(g5472), .IN2(g1116), .Q(n13683) );
  AND2X1 U13867 ( .IN1(g1088), .IN2(g1122), .Q(n13681) );
  AND2X1 U13868 ( .IN1(n12833), .IN2(g996), .Q(n13679) );
  INVX0 U13869 ( .INP(n12837), .ZN(n12833) );
  OR2X1 U13870 ( .IN1(n13685), .IN2(n12185), .Q(n12837) );
  AND2X1 U13871 ( .IN1(n13686), .IN2(n13687), .Q(n13685) );
  OR2X1 U13872 ( .IN1(n4312), .IN2(g867), .Q(n13687) );
  INVX0 U13873 ( .INP(n13688), .ZN(n13686) );
  OR2X1 U13874 ( .IN1(n13689), .IN2(n13690), .Q(n13688) );
  AND2X1 U13875 ( .IN1(test_so31), .IN2(n8708), .Q(n13690) );
  AND2X1 U13876 ( .IN1(g6368), .IN2(n8710), .Q(n13689) );
  AND2X1 U13877 ( .IN1(n4363), .IN2(g1116), .Q(n13677) );
  OR2X1 U13878 ( .IN1(n13691), .IN2(n13692), .Q(g26805) );
  AND2X1 U13879 ( .IN1(n4520), .IN2(g438), .Q(n13692) );
  AND2X1 U13880 ( .IN1(n13641), .IN2(g5437), .Q(n13691) );
  XNOR2X1 U13881 ( .IN1(n13693), .IN2(n12859), .Q(n13641) );
  OR2X1 U13882 ( .IN1(n13694), .IN2(n12865), .Q(n13693) );
  OR2X1 U13883 ( .IN1(n4388), .IN2(n13695), .Q(n12865) );
  OR2X1 U13884 ( .IN1(n13696), .IN2(n13697), .Q(n13695) );
  AND2X1 U13885 ( .IN1(n13698), .IN2(n12860), .Q(n13697) );
  OR2X1 U13886 ( .IN1(n12859), .IN2(n12854), .Q(n13698) );
  INVX0 U13887 ( .INP(n12857), .ZN(n12854) );
  AND2X1 U13888 ( .IN1(n12856), .IN2(n13699), .Q(n13696) );
  OR2X1 U13889 ( .IN1(n12857), .IN2(n12855), .Q(n13699) );
  INVX0 U13890 ( .INP(n12859), .ZN(n12855) );
  INVX0 U13891 ( .INP(n12860), .ZN(n12856) );
  AND2X1 U13892 ( .IN1(n13700), .IN2(n13701), .Q(n13694) );
  OR2X1 U13893 ( .IN1(n4506), .IN2(g447), .Q(n13701) );
  INVX0 U13894 ( .INP(n12862), .ZN(n13700) );
  OR2X1 U13895 ( .IN1(n13702), .IN2(n13703), .Q(n12862) );
  AND2X1 U13896 ( .IN1(n8802), .IN2(n10475), .Q(n13703) );
  AND2X1 U13897 ( .IN1(n8801), .IN2(n10899), .Q(n13702) );
  OR2X1 U13898 ( .IN1(n13704), .IN2(n13705), .Q(g26804) );
  AND2X1 U13899 ( .IN1(n4499), .IN2(g432), .Q(n13705) );
  AND2X1 U13900 ( .IN1(g6447), .IN2(n13676), .Q(n13704) );
  OR2X1 U13901 ( .IN1(n13706), .IN2(n13707), .Q(g26803) );
  AND2X1 U13902 ( .IN1(n4520), .IN2(g429), .Q(n13707) );
  AND2X1 U13903 ( .IN1(g5437), .IN2(n13676), .Q(n13706) );
  OR2X1 U13904 ( .IN1(n13708), .IN2(n13709), .Q(n13676) );
  AND2X1 U13905 ( .IN1(n4388), .IN2(n12860), .Q(n13709) );
  OR2X1 U13906 ( .IN1(n13710), .IN2(n13711), .Q(n12860) );
  OR2X1 U13907 ( .IN1(n13712), .IN2(n13713), .Q(n13711) );
  AND2X1 U13908 ( .IN1(g6447), .IN2(g432), .Q(n13713) );
  AND2X1 U13909 ( .IN1(n4640), .IN2(g435), .Q(n13712) );
  AND2X1 U13910 ( .IN1(g5437), .IN2(g429), .Q(n13710) );
  AND2X1 U13911 ( .IN1(n12857), .IN2(g309), .Q(n13708) );
  AND2X1 U13912 ( .IN1(n13714), .IN2(n13715), .Q(n12857) );
  INVX0 U13913 ( .INP(n12217), .ZN(n13715) );
  OR2X1 U13914 ( .IN1(n13716), .IN2(n13717), .Q(n13714) );
  AND2X1 U13915 ( .IN1(g6313), .IN2(n8720), .Q(n13717) );
  OR2X1 U13916 ( .IN1(n13718), .IN2(n13719), .Q(n13716) );
  AND2X1 U13917 ( .IN1(g6231), .IN2(n8721), .Q(n13719) );
  AND2X1 U13918 ( .IN1(g165), .IN2(n8719), .Q(n13718) );
  AND2X1 U13919 ( .IN1(n13720), .IN2(n9662), .Q(g26798) );
  XOR2X1 U13920 ( .IN1(n13721), .IN2(n4355), .Q(n13720) );
  AND2X1 U13921 ( .IN1(n13722), .IN2(n12737), .Q(g26795) );
  XNOR2X1 U13922 ( .IN1(test_so92), .IN2(n13560), .Q(n13722) );
  AND2X1 U13923 ( .IN1(n13723), .IN2(n12741), .Q(g26789) );
  XOR2X1 U13924 ( .IN1(n12873), .IN2(n4468), .Q(n13723) );
  AND2X1 U13925 ( .IN1(n13724), .IN2(n13725), .Q(g26786) );
  XOR2X1 U13926 ( .IN1(n8281), .IN2(n3741), .Q(n13725) );
  AND2X1 U13927 ( .IN1(n13726), .IN2(n12745), .Q(g26781) );
  XOR2X1 U13928 ( .IN1(n12879), .IN2(n4469), .Q(n13726) );
  AND2X1 U13929 ( .IN1(n13727), .IN2(n12226), .Q(g26776) );
  XNOR2X1 U13930 ( .IN1(test_so28), .IN2(n12885), .Q(n13727) );
  AND2X1 U13931 ( .IN1(n13728), .IN2(n13729), .Q(g26677) );
  INVX0 U13932 ( .INP(n13730), .ZN(n13729) );
  AND2X1 U13933 ( .IN1(n13731), .IN2(n4407), .Q(n13730) );
  OR2X1 U13934 ( .IN1(n13732), .IN2(n4397), .Q(n13731) );
  AND2X1 U13935 ( .IN1(n13560), .IN2(n12737), .Q(n13728) );
  OR2X1 U13936 ( .IN1(n13732), .IN2(n13733), .Q(n13560) );
  OR2X1 U13937 ( .IN1(n4407), .IN2(n4397), .Q(n13733) );
  OR2X1 U13938 ( .IN1(n13734), .IN2(n13735), .Q(g26676) );
  AND2X1 U13939 ( .IN1(n13736), .IN2(n10398), .Q(n13735) );
  AND2X1 U13940 ( .IN1(n13737), .IN2(g2479), .Q(n13734) );
  OR2X1 U13941 ( .IN1(n4524), .IN2(n13738), .Q(n13737) );
  OR2X1 U13942 ( .IN1(n13739), .IN2(n13740), .Q(g26675) );
  AND2X1 U13943 ( .IN1(n13741), .IN2(n10403), .Q(n13740) );
  AND2X1 U13944 ( .IN1(n13742), .IN2(g1783), .Q(n13739) );
  OR2X1 U13945 ( .IN1(n4511), .IN2(n13743), .Q(n13742) );
  OR2X1 U13946 ( .IN1(n13744), .IN2(n13745), .Q(g26672) );
  AND2X1 U13947 ( .IN1(n13736), .IN2(n10408), .Q(n13745) );
  AND2X1 U13948 ( .IN1(n13746), .IN2(g2478), .Q(n13744) );
  OR2X1 U13949 ( .IN1(n4516), .IN2(n13738), .Q(n13746) );
  AND2X1 U13950 ( .IN1(n13747), .IN2(n13748), .Q(g26671) );
  INVX0 U13951 ( .INP(n13749), .ZN(n13748) );
  AND2X1 U13952 ( .IN1(n13750), .IN2(n4409), .Q(n13749) );
  OR2X1 U13953 ( .IN1(n13751), .IN2(n4399), .Q(n13750) );
  AND2X1 U13954 ( .IN1(n12873), .IN2(n12741), .Q(n13747) );
  OR2X1 U13955 ( .IN1(n13751), .IN2(n13752), .Q(n12873) );
  OR2X1 U13956 ( .IN1(n4409), .IN2(n4399), .Q(n13752) );
  OR2X1 U13957 ( .IN1(n13753), .IN2(n13754), .Q(g26670) );
  AND2X1 U13958 ( .IN1(n13741), .IN2(n10412), .Q(n13754) );
  AND2X1 U13959 ( .IN1(n13755), .IN2(g1785), .Q(n13753) );
  OR2X1 U13960 ( .IN1(n4525), .IN2(n13743), .Q(n13755) );
  OR2X1 U13961 ( .IN1(n13756), .IN2(n13757), .Q(g26669) );
  AND2X1 U13962 ( .IN1(n13758), .IN2(g1088), .Q(n13757) );
  AND2X1 U13963 ( .IN1(n13759), .IN2(g1089), .Q(n13756) );
  OR2X1 U13964 ( .IN1(n4381), .IN2(n13760), .Q(n13759) );
  OR2X1 U13965 ( .IN1(n13761), .IN2(n13762), .Q(g26667) );
  AND2X1 U13966 ( .IN1(n13741), .IN2(n10419), .Q(n13762) );
  AND2X1 U13967 ( .IN1(g1690), .IN2(n13743), .Q(n13741) );
  AND2X1 U13968 ( .IN1(test_so60), .IN2(n13763), .Q(n13761) );
  OR2X1 U13969 ( .IN1(n4518), .IN2(n13743), .Q(n13763) );
  OR2X1 U13970 ( .IN1(n11494), .IN2(n13764), .Q(n13743) );
  OR2X1 U13971 ( .IN1(n4386), .IN2(n11251), .Q(n13764) );
  OR2X1 U13972 ( .IN1(n13765), .IN2(n13766), .Q(n11251) );
  OR2X1 U13973 ( .IN1(n13767), .IN2(n13768), .Q(n13766) );
  OR2X1 U13974 ( .IN1(n13769), .IN2(n13770), .Q(n13768) );
  XNOR2X1 U13975 ( .IN1(n13771), .IN2(n10760), .Q(n13770) );
  AND2X1 U13976 ( .IN1(n13772), .IN2(n13773), .Q(n13771) );
  OR2X1 U13977 ( .IN1(n4368), .IN2(g1541), .Q(n13773) );
  AND2X1 U13978 ( .IN1(n13774), .IN2(n13775), .Q(n13772) );
  OR2X1 U13979 ( .IN1(n4317), .IN2(g1542), .Q(n13775) );
  OR2X1 U13980 ( .IN1(n4515), .IN2(g1543), .Q(n13774) );
  XNOR2X1 U13981 ( .IN1(g1481), .IN2(n13776), .Q(n13769) );
  AND2X1 U13982 ( .IN1(n13777), .IN2(n13778), .Q(n13776) );
  OR2X1 U13983 ( .IN1(n4368), .IN2(g1523), .Q(n13778) );
  AND2X1 U13984 ( .IN1(n13779), .IN2(n13780), .Q(n13777) );
  OR2X1 U13985 ( .IN1(n4515), .IN2(g1525), .Q(n13780) );
  OR2X1 U13986 ( .IN1(n4317), .IN2(g1524), .Q(n13779) );
  OR2X1 U13987 ( .IN1(n13781), .IN2(n13782), .Q(n13767) );
  OR2X1 U13988 ( .IN1(n13783), .IN2(n13784), .Q(n13782) );
  XNOR2X1 U13989 ( .IN1(g1471), .IN2(n13785), .Q(n13784) );
  AND2X1 U13990 ( .IN1(n13786), .IN2(n13787), .Q(n13785) );
  OR2X1 U13991 ( .IN1(n4368), .IN2(g1511), .Q(n13787) );
  AND2X1 U13992 ( .IN1(n13788), .IN2(n13789), .Q(n13786) );
  OR2X1 U13993 ( .IN1(n4515), .IN2(g1513), .Q(n13789) );
  OR2X1 U13994 ( .IN1(n4317), .IN2(g1512), .Q(n13788) );
  XNOR2X1 U13995 ( .IN1(g1476), .IN2(n13790), .Q(n13783) );
  AND2X1 U13996 ( .IN1(n13791), .IN2(n13792), .Q(n13790) );
  OR2X1 U13997 ( .IN1(n4368), .IN2(g1514), .Q(n13792) );
  AND2X1 U13998 ( .IN1(n13793), .IN2(n13794), .Q(n13791) );
  OR2X1 U13999 ( .IN1(n4515), .IN2(g1516), .Q(n13794) );
  OR2X1 U14000 ( .IN1(n4317), .IN2(test_so52), .Q(n13793) );
  XNOR2X1 U14001 ( .IN1(n13795), .IN2(n11819), .Q(n13781) );
  AND2X1 U14002 ( .IN1(n13796), .IN2(n13797), .Q(n13795) );
  OR2X1 U14003 ( .IN1(n4368), .IN2(g1544), .Q(n13797) );
  AND2X1 U14004 ( .IN1(n13798), .IN2(n13799), .Q(n13796) );
  OR2X1 U14005 ( .IN1(n4317), .IN2(g1545), .Q(n13799) );
  OR2X1 U14006 ( .IN1(n4515), .IN2(g1546), .Q(n13798) );
  OR2X1 U14007 ( .IN1(n13800), .IN2(n13801), .Q(n13765) );
  OR2X1 U14008 ( .IN1(n13802), .IN2(n13803), .Q(n13801) );
  OR2X1 U14009 ( .IN1(n13804), .IN2(n13805), .Q(n13803) );
  XNOR2X1 U14010 ( .IN1(g1501), .IN2(n13806), .Q(n13805) );
  AND2X1 U14011 ( .IN1(n13807), .IN2(n13808), .Q(n13806) );
  OR2X1 U14012 ( .IN1(n4368), .IN2(g1535), .Q(n13808) );
  AND2X1 U14013 ( .IN1(n13809), .IN2(n13810), .Q(n13807) );
  OR2X1 U14014 ( .IN1(n4317), .IN2(g1536), .Q(n13810) );
  OR2X1 U14015 ( .IN1(n4515), .IN2(test_so53), .Q(n13809) );
  XNOR2X1 U14016 ( .IN1(g1496), .IN2(n13811), .Q(n13804) );
  AND2X1 U14017 ( .IN1(n13812), .IN2(n13813), .Q(n13811) );
  OR2X1 U14018 ( .IN1(n4368), .IN2(g1532), .Q(n13813) );
  AND2X1 U14019 ( .IN1(n13814), .IN2(n13815), .Q(n13812) );
  OR2X1 U14020 ( .IN1(n4317), .IN2(g1533), .Q(n13815) );
  OR2X1 U14021 ( .IN1(n4515), .IN2(g1534), .Q(n13814) );
  XNOR2X1 U14022 ( .IN1(g1486), .IN2(n13816), .Q(n13802) );
  AND2X1 U14023 ( .IN1(n13817), .IN2(n13818), .Q(n13816) );
  OR2X1 U14024 ( .IN1(n4368), .IN2(g1526), .Q(n13818) );
  AND2X1 U14025 ( .IN1(n13819), .IN2(n13820), .Q(n13817) );
  OR2X1 U14026 ( .IN1(n4515), .IN2(g1528), .Q(n13820) );
  OR2X1 U14027 ( .IN1(n4317), .IN2(g1527), .Q(n13819) );
  OR2X1 U14028 ( .IN1(n13821), .IN2(n13822), .Q(n13800) );
  OR2X1 U14029 ( .IN1(n10443), .IN2(n13823), .Q(n13822) );
  XNOR2X1 U14030 ( .IN1(g1506), .IN2(n13824), .Q(n13823) );
  AND2X1 U14031 ( .IN1(n13825), .IN2(n13826), .Q(n13824) );
  OR2X1 U14032 ( .IN1(n4368), .IN2(g1538), .Q(n13826) );
  AND2X1 U14033 ( .IN1(n13827), .IN2(n13828), .Q(n13825) );
  OR2X1 U14034 ( .IN1(n4515), .IN2(g1540), .Q(n13828) );
  OR2X1 U14035 ( .IN1(n4317), .IN2(g1539), .Q(n13827) );
  INVX0 U14036 ( .INP(n3070), .ZN(n10443) );
  XNOR2X1 U14037 ( .IN1(g1491), .IN2(n13829), .Q(n13821) );
  AND2X1 U14038 ( .IN1(n13830), .IN2(n13831), .Q(n13829) );
  OR2X1 U14039 ( .IN1(n4368), .IN2(g1529), .Q(n13831) );
  AND2X1 U14040 ( .IN1(n13832), .IN2(n13833), .Q(n13830) );
  OR2X1 U14041 ( .IN1(n4515), .IN2(g1531), .Q(n13833) );
  OR2X1 U14042 ( .IN1(n4317), .IN2(g1530), .Q(n13832) );
  OR2X1 U14043 ( .IN1(n13834), .IN2(n13835), .Q(n11494) );
  OR2X1 U14044 ( .IN1(n13836), .IN2(n13837), .Q(n13835) );
  INVX0 U14045 ( .INP(n13838), .ZN(n13837) );
  OR2X1 U14046 ( .IN1(n4518), .IN2(test_so60), .Q(n13838) );
  AND2X1 U14047 ( .IN1(n8786), .IN2(n10403), .Q(n13836) );
  AND2X1 U14048 ( .IN1(n8776), .IN2(n10412), .Q(n13834) );
  AND2X1 U14049 ( .IN1(n13839), .IN2(n13840), .Q(g26666) );
  INVX0 U14050 ( .INP(n13841), .ZN(n13840) );
  AND2X1 U14051 ( .IN1(n13842), .IN2(n4411), .Q(n13841) );
  OR2X1 U14052 ( .IN1(n13843), .IN2(n4401), .Q(n13842) );
  AND2X1 U14053 ( .IN1(n12879), .IN2(n12745), .Q(n13839) );
  OR2X1 U14054 ( .IN1(n13843), .IN2(n13844), .Q(n12879) );
  OR2X1 U14055 ( .IN1(n4411), .IN2(n4401), .Q(n13844) );
  OR2X1 U14056 ( .IN1(n13845), .IN2(n13846), .Q(g26665) );
  AND2X1 U14057 ( .IN1(n13758), .IN2(g6712), .Q(n13846) );
  AND2X1 U14058 ( .IN1(n13847), .IN2(g1091), .Q(n13845) );
  OR2X1 U14059 ( .IN1(n4364), .IN2(n13760), .Q(n13847) );
  OR2X1 U14060 ( .IN1(n13848), .IN2(n13849), .Q(g26664) );
  AND2X1 U14061 ( .IN1(n13850), .IN2(n10465), .Q(n13849) );
  AND2X1 U14062 ( .IN1(n13851), .IN2(g402), .Q(n13848) );
  OR2X1 U14063 ( .IN1(n4506), .IN2(n13852), .Q(n13851) );
  OR2X1 U14064 ( .IN1(n13853), .IN2(n13854), .Q(g26661) );
  AND2X1 U14065 ( .IN1(n13758), .IN2(g5472), .Q(n13854) );
  AND2X1 U14066 ( .IN1(g996), .IN2(n13760), .Q(n13758) );
  AND2X1 U14067 ( .IN1(n13855), .IN2(g1090), .Q(n13853) );
  OR2X1 U14068 ( .IN1(n4363), .IN2(n13760), .Q(n13855) );
  OR2X1 U14069 ( .IN1(n11509), .IN2(n13856), .Q(n13760) );
  OR2X1 U14070 ( .IN1(n4387), .IN2(n11311), .Q(n13856) );
  OR2X1 U14071 ( .IN1(n13857), .IN2(n13858), .Q(n11311) );
  OR2X1 U14072 ( .IN1(n13859), .IN2(n13860), .Q(n13858) );
  OR2X1 U14073 ( .IN1(n13861), .IN2(n13862), .Q(n13860) );
  XNOR2X1 U14074 ( .IN1(n10800), .IN2(n13863), .Q(n13862) );
  AND2X1 U14075 ( .IN1(n13864), .IN2(n13865), .Q(n13863) );
  OR2X1 U14076 ( .IN1(n9118), .IN2(g847), .Q(n13865) );
  AND2X1 U14077 ( .IN1(n13866), .IN2(n13867), .Q(n13864) );
  OR2X1 U14078 ( .IN1(n4312), .IN2(g849), .Q(n13867) );
  OR2X1 U14079 ( .IN1(n4323), .IN2(g848), .Q(n13866) );
  XNOR2X1 U14080 ( .IN1(n13868), .IN2(n13869), .Q(n13861) );
  AND2X1 U14081 ( .IN1(n13870), .IN2(n13871), .Q(n13869) );
  OR2X1 U14082 ( .IN1(n9118), .IN2(g850), .Q(n13871) );
  AND2X1 U14083 ( .IN1(n13872), .IN2(n13873), .Q(n13870) );
  OR2X1 U14084 ( .IN1(n4312), .IN2(g852), .Q(n13873) );
  OR2X1 U14085 ( .IN1(n4323), .IN2(g851), .Q(n13872) );
  OR2X1 U14086 ( .IN1(n13874), .IN2(n13875), .Q(n13859) );
  OR2X1 U14087 ( .IN1(n13876), .IN2(n13877), .Q(n13875) );
  XOR2X1 U14088 ( .IN1(g793), .IN2(n13878), .Q(n13877) );
  OR2X1 U14089 ( .IN1(n13879), .IN2(n13880), .Q(n13878) );
  OR2X1 U14090 ( .IN1(n13881), .IN2(n13882), .Q(n13880) );
  AND2X1 U14091 ( .IN1(n9022), .IN2(g6368), .Q(n13882) );
  AND2X1 U14092 ( .IN1(n8657), .IN2(test_so31), .Q(n13881) );
  AND2X1 U14093 ( .IN1(n9021), .IN2(g6518), .Q(n13879) );
  XOR2X1 U14094 ( .IN1(g785), .IN2(n13883), .Q(n13876) );
  OR2X1 U14095 ( .IN1(n13884), .IN2(n13885), .Q(n13883) );
  OR2X1 U14096 ( .IN1(n13886), .IN2(n13887), .Q(n13885) );
  AND2X1 U14097 ( .IN1(n9026), .IN2(g6368), .Q(n13887) );
  AND2X1 U14098 ( .IN1(n8659), .IN2(test_so31), .Q(n13886) );
  AND2X1 U14099 ( .IN1(n9025), .IN2(g6518), .Q(n13884) );
  XNOR2X1 U14100 ( .IN1(n4375), .IN2(n13888), .Q(n13874) );
  OR2X1 U14101 ( .IN1(n13889), .IN2(n13890), .Q(n13888) );
  OR2X1 U14102 ( .IN1(n13891), .IN2(n13892), .Q(n13890) );
  AND2X1 U14103 ( .IN1(n9024), .IN2(g6368), .Q(n13892) );
  AND2X1 U14104 ( .IN1(n8658), .IN2(test_so31), .Q(n13891) );
  AND2X1 U14105 ( .IN1(n9023), .IN2(g6518), .Q(n13889) );
  OR2X1 U14106 ( .IN1(n13893), .IN2(n13894), .Q(n13857) );
  OR2X1 U14107 ( .IN1(n13895), .IN2(n13896), .Q(n13894) );
  OR2X1 U14108 ( .IN1(n13897), .IN2(n13898), .Q(n13896) );
  XNOR2X1 U14109 ( .IN1(g809), .IN2(n13899), .Q(n13898) );
  AND2X1 U14110 ( .IN1(n13900), .IN2(n13901), .Q(n13899) );
  OR2X1 U14111 ( .IN1(n9118), .IN2(g841), .Q(n13901) );
  AND2X1 U14112 ( .IN1(n13902), .IN2(n13903), .Q(n13900) );
  OR2X1 U14113 ( .IN1(n4312), .IN2(g843), .Q(n13903) );
  OR2X1 U14114 ( .IN1(n4323), .IN2(g842), .Q(n13902) );
  XNOR2X1 U14115 ( .IN1(g805), .IN2(n13904), .Q(n13897) );
  AND2X1 U14116 ( .IN1(n13905), .IN2(n13906), .Q(n13904) );
  OR2X1 U14117 ( .IN1(n9118), .IN2(g838), .Q(n13906) );
  AND2X1 U14118 ( .IN1(n13907), .IN2(n13908), .Q(n13905) );
  OR2X1 U14119 ( .IN1(n4312), .IN2(g840), .Q(n13908) );
  OR2X1 U14120 ( .IN1(test_so32), .IN2(n4323), .Q(n13907) );
  XNOR2X1 U14121 ( .IN1(n4391), .IN2(n13909), .Q(n13895) );
  OR2X1 U14122 ( .IN1(n13910), .IN2(n13911), .Q(n13909) );
  OR2X1 U14123 ( .IN1(n13912), .IN2(n13913), .Q(n13911) );
  AND2X1 U14124 ( .IN1(n9020), .IN2(g6368), .Q(n13913) );
  AND2X1 U14125 ( .IN1(n8656), .IN2(test_so31), .Q(n13912) );
  AND2X1 U14126 ( .IN1(n9019), .IN2(g6518), .Q(n13910) );
  OR2X1 U14127 ( .IN1(n13914), .IN2(n13915), .Q(n13893) );
  OR2X1 U14128 ( .IN1(n10247), .IN2(n13916), .Q(n13915) );
  XOR2X1 U14129 ( .IN1(g813), .IN2(n13917), .Q(n13916) );
  OR2X1 U14130 ( .IN1(n13918), .IN2(n13919), .Q(n13917) );
  OR2X1 U14131 ( .IN1(n13920), .IN2(n13921), .Q(n13919) );
  AND2X1 U14132 ( .IN1(n9013), .IN2(g6368), .Q(n13921) );
  AND2X1 U14133 ( .IN1(n8652), .IN2(test_so31), .Q(n13920) );
  AND2X1 U14134 ( .IN1(n9012), .IN2(g6518), .Q(n13918) );
  INVX0 U14135 ( .INP(n3102), .ZN(n10247) );
  XOR2X1 U14136 ( .IN1(g801), .IN2(n13922), .Q(n13914) );
  OR2X1 U14137 ( .IN1(n13923), .IN2(n13924), .Q(n13922) );
  OR2X1 U14138 ( .IN1(n13925), .IN2(n13926), .Q(n13924) );
  AND2X1 U14139 ( .IN1(n9018), .IN2(g6368), .Q(n13926) );
  AND2X1 U14140 ( .IN1(n8655), .IN2(test_so31), .Q(n13925) );
  AND2X1 U14141 ( .IN1(n9017), .IN2(g6518), .Q(n13923) );
  OR2X1 U14142 ( .IN1(n13927), .IN2(n13928), .Q(n11509) );
  OR2X1 U14143 ( .IN1(n13929), .IN2(n13930), .Q(n13928) );
  AND2X1 U14144 ( .IN1(n8779), .IN2(g6712), .Q(n13930) );
  AND2X1 U14145 ( .IN1(n8792), .IN2(g5472), .Q(n13929) );
  AND2X1 U14146 ( .IN1(n8791), .IN2(g1088), .Q(n13927) );
  AND2X1 U14147 ( .IN1(n13931), .IN2(n13932), .Q(g26660) );
  INVX0 U14148 ( .INP(n13933), .ZN(n13932) );
  AND2X1 U14149 ( .IN1(n13934), .IN2(n4413), .Q(n13933) );
  OR2X1 U14150 ( .IN1(n13935), .IN2(n4403), .Q(n13934) );
  AND2X1 U14151 ( .IN1(n12885), .IN2(n12226), .Q(n13931) );
  OR2X1 U14152 ( .IN1(n13935), .IN2(n13936), .Q(n12885) );
  OR2X1 U14153 ( .IN1(n4413), .IN2(n4403), .Q(n13936) );
  OR2X1 U14154 ( .IN1(n13937), .IN2(n13938), .Q(g26659) );
  AND2X1 U14155 ( .IN1(n13850), .IN2(n10899), .Q(n13938) );
  AND2X1 U14156 ( .IN1(n13939), .IN2(g404), .Q(n13937) );
  OR2X1 U14157 ( .IN1(n4499), .IN2(n13852), .Q(n13939) );
  OR2X1 U14158 ( .IN1(n13940), .IN2(n13941), .Q(g26655) );
  AND2X1 U14159 ( .IN1(n13850), .IN2(n10475), .Q(n13941) );
  AND2X1 U14160 ( .IN1(g309), .IN2(n13852), .Q(n13850) );
  AND2X1 U14161 ( .IN1(n13942), .IN2(g403), .Q(n13940) );
  OR2X1 U14162 ( .IN1(n4520), .IN2(n13852), .Q(n13942) );
  OR2X1 U14163 ( .IN1(n11522), .IN2(n13943), .Q(n13852) );
  OR2X1 U14164 ( .IN1(n4388), .IN2(n11365), .Q(n13943) );
  OR2X1 U14165 ( .IN1(n13944), .IN2(n13945), .Q(n11365) );
  OR2X1 U14166 ( .IN1(n13946), .IN2(n13947), .Q(n13945) );
  OR2X1 U14167 ( .IN1(n13948), .IN2(n13949), .Q(n13947) );
  XNOR2X1 U14168 ( .IN1(n13950), .IN2(n10824), .Q(n13949) );
  AND2X1 U14169 ( .IN1(n13951), .IN2(n13952), .Q(n13950) );
  OR2X1 U14170 ( .IN1(n4369), .IN2(g159), .Q(n13952) );
  AND2X1 U14171 ( .IN1(n13953), .IN2(n13954), .Q(n13951) );
  OR2X1 U14172 ( .IN1(n4318), .IN2(g160), .Q(n13954) );
  OR2X1 U14173 ( .IN1(n4512), .IN2(g161), .Q(n13953) );
  XNOR2X1 U14174 ( .IN1(g105), .IN2(n13955), .Q(n13948) );
  AND2X1 U14175 ( .IN1(n13956), .IN2(n13957), .Q(n13955) );
  OR2X1 U14176 ( .IN1(n4369), .IN2(g141), .Q(n13957) );
  AND2X1 U14177 ( .IN1(n13958), .IN2(n13959), .Q(n13956) );
  OR2X1 U14178 ( .IN1(n4512), .IN2(g143), .Q(n13959) );
  OR2X1 U14179 ( .IN1(n4318), .IN2(g142), .Q(n13958) );
  OR2X1 U14180 ( .IN1(n13960), .IN2(n13961), .Q(n13946) );
  OR2X1 U14181 ( .IN1(n13962), .IN2(n13963), .Q(n13961) );
  XOR2X1 U14182 ( .IN1(n4380), .IN2(n13964), .Q(n13963) );
  AND2X1 U14183 ( .IN1(n13965), .IN2(n13966), .Q(n13964) );
  OR2X1 U14184 ( .IN1(n4369), .IN2(g129), .Q(n13966) );
  AND2X1 U14185 ( .IN1(n13967), .IN2(n13968), .Q(n13965) );
  OR2X1 U14186 ( .IN1(n4512), .IN2(g131), .Q(n13968) );
  OR2X1 U14187 ( .IN1(n4318), .IN2(g130), .Q(n13967) );
  XOR2X1 U14188 ( .IN1(n4376), .IN2(n13969), .Q(n13962) );
  AND2X1 U14189 ( .IN1(n13970), .IN2(n13971), .Q(n13969) );
  OR2X1 U14190 ( .IN1(n4369), .IN2(g132), .Q(n13971) );
  AND2X1 U14191 ( .IN1(n13972), .IN2(n13973), .Q(n13970) );
  OR2X1 U14192 ( .IN1(n4512), .IN2(g134), .Q(n13973) );
  OR2X1 U14193 ( .IN1(n4318), .IN2(g133), .Q(n13972) );
  XNOR2X1 U14194 ( .IN1(n13974), .IN2(n13975), .Q(n13960) );
  AND2X1 U14195 ( .IN1(n13976), .IN2(n13977), .Q(n13974) );
  OR2X1 U14196 ( .IN1(n4369), .IN2(g162), .Q(n13977) );
  AND2X1 U14197 ( .IN1(n13978), .IN2(n13979), .Q(n13976) );
  OR2X1 U14198 ( .IN1(n4512), .IN2(g164), .Q(n13979) );
  OR2X1 U14199 ( .IN1(n4318), .IN2(test_so12), .Q(n13978) );
  OR2X1 U14200 ( .IN1(n13980), .IN2(n13981), .Q(n13944) );
  OR2X1 U14201 ( .IN1(n13982), .IN2(n13983), .Q(n13981) );
  OR2X1 U14202 ( .IN1(n13984), .IN2(n13985), .Q(n13983) );
  XNOR2X1 U14203 ( .IN1(g121), .IN2(n13986), .Q(n13985) );
  AND2X1 U14204 ( .IN1(n13987), .IN2(n13988), .Q(n13986) );
  OR2X1 U14205 ( .IN1(n4369), .IN2(g153), .Q(n13988) );
  AND2X1 U14206 ( .IN1(n13989), .IN2(n13990), .Q(n13987) );
  OR2X1 U14207 ( .IN1(n4318), .IN2(g154), .Q(n13990) );
  OR2X1 U14208 ( .IN1(n4512), .IN2(g155), .Q(n13989) );
  XNOR2X1 U14209 ( .IN1(g117), .IN2(n13991), .Q(n13984) );
  AND2X1 U14210 ( .IN1(n13992), .IN2(n13993), .Q(n13991) );
  OR2X1 U14211 ( .IN1(n4369), .IN2(g150), .Q(n13993) );
  AND2X1 U14212 ( .IN1(n13994), .IN2(n13995), .Q(n13992) );
  OR2X1 U14213 ( .IN1(n4318), .IN2(g151), .Q(n13995) );
  OR2X1 U14214 ( .IN1(n4512), .IN2(g152), .Q(n13994) );
  XOR2X1 U14215 ( .IN1(n4392), .IN2(n13996), .Q(n13982) );
  AND2X1 U14216 ( .IN1(n13997), .IN2(n13998), .Q(n13996) );
  OR2X1 U14217 ( .IN1(n4318), .IN2(g145), .Q(n13998) );
  AND2X1 U14218 ( .IN1(n13999), .IN2(n14000), .Q(n13997) );
  OR2X1 U14219 ( .IN1(n4512), .IN2(g146), .Q(n14000) );
  OR2X1 U14220 ( .IN1(n4369), .IN2(test_so11), .Q(n13999) );
  OR2X1 U14221 ( .IN1(n14001), .IN2(n14002), .Q(n13980) );
  OR2X1 U14222 ( .IN1(n10499), .IN2(n14003), .Q(n14002) );
  XOR2X1 U14223 ( .IN1(n4290), .IN2(n14004), .Q(n14003) );
  AND2X1 U14224 ( .IN1(n14005), .IN2(n14006), .Q(n14004) );
  OR2X1 U14225 ( .IN1(n4369), .IN2(g156), .Q(n14006) );
  AND2X1 U14226 ( .IN1(n14007), .IN2(n14008), .Q(n14005) );
  OR2X1 U14227 ( .IN1(n4512), .IN2(g158), .Q(n14008) );
  OR2X1 U14228 ( .IN1(n4318), .IN2(g157), .Q(n14007) );
  INVX0 U14229 ( .INP(n3130), .ZN(n10499) );
  XNOR2X1 U14230 ( .IN1(g113), .IN2(n14009), .Q(n14001) );
  AND2X1 U14231 ( .IN1(n14010), .IN2(n14011), .Q(n14009) );
  OR2X1 U14232 ( .IN1(n4369), .IN2(g147), .Q(n14011) );
  AND2X1 U14233 ( .IN1(n14012), .IN2(n14013), .Q(n14010) );
  OR2X1 U14234 ( .IN1(n4512), .IN2(g149), .Q(n14013) );
  OR2X1 U14235 ( .IN1(n4318), .IN2(g148), .Q(n14012) );
  OR2X1 U14236 ( .IN1(n14014), .IN2(n14015), .Q(n11522) );
  OR2X1 U14237 ( .IN1(n14016), .IN2(n14017), .Q(n14015) );
  AND2X1 U14238 ( .IN1(n8797), .IN2(n10465), .Q(n14017) );
  AND2X1 U14239 ( .IN1(n8798), .IN2(n10899), .Q(n14016) );
  AND2X1 U14240 ( .IN1(n8799), .IN2(n10475), .Q(n14014) );
  OR2X1 U14241 ( .IN1(n14018), .IN2(n14019), .Q(g26616) );
  AND2X1 U14242 ( .IN1(n14020), .IN2(g2624), .Q(n14019) );
  AND2X1 U14243 ( .IN1(n4299), .IN2(g2571), .Q(n14018) );
  OR2X1 U14244 ( .IN1(n14021), .IN2(n14022), .Q(g26596) );
  AND2X1 U14245 ( .IN1(n14020), .IN2(g7390), .Q(n14022) );
  AND2X1 U14246 ( .IN1(n4370), .IN2(g2568), .Q(n14021) );
  OR2X1 U14247 ( .IN1(n14023), .IN2(n14024), .Q(g26592) );
  AND2X1 U14248 ( .IN1(n14025), .IN2(g1930), .Q(n14024) );
  AND2X1 U14249 ( .IN1(n4366), .IN2(g1877), .Q(n14023) );
  OR2X1 U14250 ( .IN1(n14026), .IN2(n14027), .Q(g26575) );
  AND2X1 U14251 ( .IN1(n14020), .IN2(n11411), .Q(n14027) );
  AND2X1 U14252 ( .IN1(n14028), .IN2(n14029), .Q(n14020) );
  AND2X1 U14253 ( .IN1(g2584), .IN2(n9946), .Q(n14029) );
  AND2X1 U14254 ( .IN1(n4314), .IN2(g2565), .Q(n14026) );
  OR2X1 U14255 ( .IN1(n14030), .IN2(n14031), .Q(g26573) );
  AND2X1 U14256 ( .IN1(n14025), .IN2(g7194), .Q(n14031) );
  AND2X1 U14257 ( .IN1(n4315), .IN2(g1874), .Q(n14030) );
  OR2X1 U14258 ( .IN1(n14032), .IN2(n14033), .Q(g26569) );
  AND2X1 U14259 ( .IN1(n14034), .IN2(g1236), .Q(n14033) );
  AND2X1 U14260 ( .IN1(n4300), .IN2(g1183), .Q(n14032) );
  OR2X1 U14261 ( .IN1(n14035), .IN2(n14036), .Q(g26559) );
  AND2X1 U14262 ( .IN1(test_so68), .IN2(n4296), .Q(n14036) );
  AND2X1 U14263 ( .IN1(n14025), .IN2(n12379), .Q(n14035) );
  AND2X1 U14264 ( .IN1(n14037), .IN2(n14038), .Q(n14025) );
  AND2X1 U14265 ( .IN1(g1890), .IN2(n10079), .Q(n14038) );
  OR2X1 U14266 ( .IN1(n14039), .IN2(n14040), .Q(g26557) );
  AND2X1 U14267 ( .IN1(n14034), .IN2(g6944), .Q(n14040) );
  AND2X1 U14268 ( .IN1(n4316), .IN2(g1180), .Q(n14039) );
  OR2X1 U14269 ( .IN1(n14041), .IN2(n14042), .Q(g26553) );
  AND2X1 U14270 ( .IN1(n14043), .IN2(g550), .Q(n14042) );
  AND2X1 U14271 ( .IN1(n4313), .IN2(g496), .Q(n14041) );
  OR2X1 U14272 ( .IN1(n14044), .IN2(n14045), .Q(g26547) );
  AND2X1 U14273 ( .IN1(test_so47), .IN2(n4371), .Q(n14045) );
  AND2X1 U14274 ( .IN1(n14034), .IN2(n12249), .Q(n14044) );
  AND2X1 U14275 ( .IN1(n14046), .IN2(n14047), .Q(n14034) );
  AND2X1 U14276 ( .IN1(g1196), .IN2(n10214), .Q(n14047) );
  OR2X1 U14277 ( .IN1(n14048), .IN2(n14049), .Q(g26545) );
  AND2X1 U14278 ( .IN1(n14043), .IN2(g6642), .Q(n14049) );
  AND2X1 U14279 ( .IN1(n4372), .IN2(g493), .Q(n14048) );
  OR2X1 U14280 ( .IN1(n14050), .IN2(n14051), .Q(g26541) );
  AND2X1 U14281 ( .IN1(n14043), .IN2(n9810), .Q(n14051) );
  AND2X1 U14282 ( .IN1(n14052), .IN2(n14053), .Q(n14043) );
  AND2X1 U14283 ( .IN1(n9798), .IN2(test_so22), .Q(n14053) );
  AND2X1 U14284 ( .IN1(n4298), .IN2(g490), .Q(n14050) );
  AND2X1 U14285 ( .IN1(n14054), .IN2(n11527), .Q(g26532) );
  XOR2X1 U14286 ( .IN1(n8808), .IN2(n4526), .Q(n14054) );
  AND2X1 U14287 ( .IN1(n14055), .IN2(n11529), .Q(g26531) );
  XOR2X1 U14288 ( .IN1(n8812), .IN2(n4527), .Q(n14055) );
  AND2X1 U14289 ( .IN1(n14056), .IN2(n11531), .Q(g26530) );
  XNOR2X1 U14290 ( .IN1(n14057), .IN2(n8816), .Q(n14056) );
  AND2X1 U14291 ( .IN1(n14058), .IN2(n11533), .Q(g26529) );
  XOR2X1 U14292 ( .IN1(n8820), .IN2(n4528), .Q(n14058) );
  OR2X1 U14293 ( .IN1(n14059), .IN2(n14060), .Q(g26149) );
  OR2X1 U14294 ( .IN1(n14061), .IN2(n14062), .Q(n14060) );
  OR2X1 U14295 ( .IN1(n14063), .IN2(n12894), .Q(n14062) );
  AND2X1 U14296 ( .IN1(n12898), .IN2(n8086), .Q(n14063) );
  OR2X1 U14297 ( .IN1(n14064), .IN2(n14065), .Q(n14061) );
  OR2X1 U14298 ( .IN1(n14066), .IN2(n14067), .Q(n14065) );
  AND2X1 U14299 ( .IN1(n14068), .IN2(g3170), .Q(n14067) );
  AND2X1 U14300 ( .IN1(n14069), .IN2(g3173), .Q(n14066) );
  AND2X1 U14301 ( .IN1(n14070), .IN2(n8080), .Q(n14064) );
  OR2X1 U14302 ( .IN1(n14071), .IN2(n14072), .Q(n14059) );
  OR2X1 U14303 ( .IN1(n14073), .IN2(n14074), .Q(n14072) );
  OR2X1 U14304 ( .IN1(n14075), .IN2(n14076), .Q(n14074) );
  AND2X1 U14305 ( .IN1(n14077), .IN2(g3176), .Q(n14076) );
  AND2X1 U14306 ( .IN1(n12899), .IN2(n8076), .Q(n14075) );
  AND2X1 U14307 ( .IN1(n14078), .IN2(g3161), .Q(n14073) );
  OR2X1 U14308 ( .IN1(n14079), .IN2(n14080), .Q(n14071) );
  OR2X1 U14309 ( .IN1(n14081), .IN2(n14082), .Q(n14080) );
  AND2X1 U14310 ( .IN1(n3939), .IN2(n14083), .Q(n14082) );
  OR2X1 U14311 ( .IN1(n14084), .IN2(n14085), .Q(n14083) );
  OR2X1 U14312 ( .IN1(n14086), .IN2(n14087), .Q(n14085) );
  AND2X1 U14313 ( .IN1(n14088), .IN2(g3155), .Q(n14087) );
  AND2X1 U14314 ( .IN1(test_so8), .IN2(n12918), .Q(n14086) );
  AND2X1 U14315 ( .IN1(n3940), .IN2(g3185), .Q(n14084) );
  AND2X1 U14316 ( .IN1(n14089), .IN2(g3167), .Q(n14081) );
  AND2X1 U14317 ( .IN1(n3936), .IN2(n14090), .Q(n14079) );
  OR2X1 U14318 ( .IN1(n14091), .IN2(n14092), .Q(n14090) );
  OR2X1 U14319 ( .IN1(n14093), .IN2(n14094), .Q(n14092) );
  AND2X1 U14320 ( .IN1(n12905), .IN2(g3182), .Q(n14094) );
  AND2X1 U14321 ( .IN1(n14095), .IN2(g3158), .Q(n14093) );
  OR2X1 U14322 ( .IN1(n14096), .IN2(n14097), .Q(n14091) );
  AND2X1 U14323 ( .IN1(n14098), .IN2(g3164), .Q(n14097) );
  AND2X1 U14324 ( .IN1(n14099), .IN2(g3088), .Q(n14096) );
  OR2X1 U14325 ( .IN1(n14100), .IN2(n14101), .Q(g26135) );
  OR2X1 U14326 ( .IN1(n14102), .IN2(n14103), .Q(n14101) );
  OR2X1 U14327 ( .IN1(n12894), .IN2(n14104), .Q(n14103) );
  OR2X1 U14328 ( .IN1(n14105), .IN2(n14106), .Q(n14104) );
  AND2X1 U14329 ( .IN1(n8731), .IN2(n12898), .Q(n14106) );
  AND2X1 U14330 ( .IN1(n14070), .IN2(n8081), .Q(n14105) );
  OR2X1 U14331 ( .IN1(n14107), .IN2(n14108), .Q(n14102) );
  OR2X1 U14332 ( .IN1(n14109), .IN2(n14110), .Q(n14108) );
  AND2X1 U14333 ( .IN1(n14069), .IN2(g3103), .Q(n14110) );
  AND2X1 U14334 ( .IN1(n14078), .IN2(g3099), .Q(n14109) );
  AND2X1 U14335 ( .IN1(n14068), .IN2(g3102), .Q(n14107) );
  OR2X1 U14336 ( .IN1(n14111), .IN2(n14112), .Q(n14100) );
  OR2X1 U14337 ( .IN1(n14113), .IN2(n14114), .Q(n14112) );
  OR2X1 U14338 ( .IN1(n14115), .IN2(n14116), .Q(n14114) );
  AND2X1 U14339 ( .IN1(n12899), .IN2(n8077), .Q(n14116) );
  AND2X1 U14340 ( .IN1(n3936), .IN2(n14117), .Q(n14115) );
  OR2X1 U14341 ( .IN1(n14118), .IN2(n14119), .Q(n14117) );
  OR2X1 U14342 ( .IN1(n14120), .IN2(n14121), .Q(n14119) );
  AND2X1 U14343 ( .IN1(n12905), .IN2(g3106), .Q(n14121) );
  AND2X1 U14344 ( .IN1(n14095), .IN2(g3098), .Q(n14120) );
  OR2X1 U14345 ( .IN1(n14122), .IN2(n14123), .Q(n14118) );
  AND2X1 U14346 ( .IN1(n14098), .IN2(g3100), .Q(n14123) );
  AND2X1 U14347 ( .IN1(n14099), .IN2(g3108), .Q(n14122) );
  AND2X1 U14348 ( .IN1(n14077), .IN2(g3104), .Q(n14113) );
  OR2X1 U14349 ( .IN1(n14124), .IN2(n14125), .Q(n14111) );
  OR2X1 U14350 ( .IN1(n14126), .IN2(n14127), .Q(n14125) );
  AND2X1 U14351 ( .IN1(n3939), .IN2(n14128), .Q(n14127) );
  OR2X1 U14352 ( .IN1(n14129), .IN2(n14130), .Q(n14128) );
  OR2X1 U14353 ( .IN1(n14131), .IN2(n14132), .Q(n14130) );
  AND2X1 U14354 ( .IN1(n14088), .IN2(g3097), .Q(n14132) );
  AND2X1 U14355 ( .IN1(n12918), .IN2(g3105), .Q(n14131) );
  AND2X1 U14356 ( .IN1(n3940), .IN2(g3107), .Q(n14129) );
  AND2X1 U14357 ( .IN1(test_so10), .IN2(n12904), .Q(n14126) );
  OR2X1 U14358 ( .IN1(n14133), .IN2(n14134), .Q(n14124) );
  AND2X1 U14359 ( .IN1(n12909), .IN2(n12916), .Q(n14134) );
  AND2X1 U14360 ( .IN1(test_so7), .IN2(n14089), .Q(n14133) );
  OR2X1 U14361 ( .IN1(n14135), .IN2(n14136), .Q(g26104) );
  OR2X1 U14362 ( .IN1(n14137), .IN2(n14138), .Q(n14136) );
  OR2X1 U14363 ( .IN1(n12894), .IN2(n14139), .Q(n14138) );
  OR2X1 U14364 ( .IN1(n14140), .IN2(n14141), .Q(n14139) );
  AND2X1 U14365 ( .IN1(n12898), .IN2(n8087), .Q(n14141) );
  AND2X1 U14366 ( .IN1(n14070), .IN2(n8082), .Q(n14140) );
  OR2X1 U14367 ( .IN1(n14142), .IN2(n14143), .Q(n14137) );
  OR2X1 U14368 ( .IN1(n14144), .IN2(n14145), .Q(n14143) );
  AND2X1 U14369 ( .IN1(n14069), .IN2(g3091), .Q(n14145) );
  AND2X1 U14370 ( .IN1(n3933), .IN2(n14146), .Q(n14069) );
  AND2X1 U14371 ( .IN1(n4406), .IN2(n12919), .Q(n14146) );
  AND2X1 U14372 ( .IN1(n14078), .IN2(g3084), .Q(n14144) );
  AND2X1 U14373 ( .IN1(n3933), .IN2(n14147), .Q(n14078) );
  AND2X1 U14374 ( .IN1(n4406), .IN2(n3939), .Q(n14147) );
  AND2X1 U14375 ( .IN1(g3207), .IN2(n4405), .Q(n3933) );
  AND2X1 U14376 ( .IN1(n14068), .IN2(g3087), .Q(n14142) );
  AND2X1 U14377 ( .IN1(n14095), .IN2(n12908), .Q(n14068) );
  OR2X1 U14378 ( .IN1(n14148), .IN2(n14149), .Q(n14135) );
  OR2X1 U14379 ( .IN1(n14150), .IN2(n14151), .Q(n14149) );
  OR2X1 U14380 ( .IN1(n14152), .IN2(n14153), .Q(n14151) );
  AND2X1 U14381 ( .IN1(n12899), .IN2(n8078), .Q(n14153) );
  AND2X1 U14382 ( .IN1(n14154), .IN2(n12918), .Q(n12899) );
  AND2X1 U14383 ( .IN1(n3936), .IN2(n14155), .Q(n14152) );
  OR2X1 U14384 ( .IN1(n14156), .IN2(n14157), .Q(n14155) );
  OR2X1 U14385 ( .IN1(n14158), .IN2(n14159), .Q(n14157) );
  AND2X1 U14386 ( .IN1(n12905), .IN2(g3094), .Q(n14159) );
  AND2X1 U14387 ( .IN1(n14095), .IN2(g3211), .Q(n14158) );
  OR2X1 U14388 ( .IN1(n14160), .IN2(n14161), .Q(n14156) );
  AND2X1 U14389 ( .IN1(n14098), .IN2(g3085), .Q(n14161) );
  AND2X1 U14390 ( .IN1(n14099), .IN2(g3096), .Q(n14160) );
  AND2X1 U14391 ( .IN1(g3201), .IN2(g3207), .Q(n14099) );
  AND2X1 U14392 ( .IN1(n14077), .IN2(g3092), .Q(n14150) );
  AND2X1 U14393 ( .IN1(n14098), .IN2(n12908), .Q(n14077) );
  AND2X1 U14394 ( .IN1(g3188), .IN2(n12919), .Q(n12908) );
  AND2X1 U14395 ( .IN1(g3207), .IN2(n4406), .Q(n14098) );
  OR2X1 U14396 ( .IN1(n14162), .IN2(n14163), .Q(n14148) );
  OR2X1 U14397 ( .IN1(n14164), .IN2(n14165), .Q(n14163) );
  AND2X1 U14398 ( .IN1(n3939), .IN2(n14166), .Q(n14165) );
  OR2X1 U14399 ( .IN1(n14167), .IN2(n14168), .Q(n14166) );
  OR2X1 U14400 ( .IN1(n14169), .IN2(n14170), .Q(n14168) );
  AND2X1 U14401 ( .IN1(test_so6), .IN2(n14088), .Q(n14170) );
  AND2X1 U14402 ( .IN1(n12918), .IN2(g3093), .Q(n14169) );
  AND2X1 U14403 ( .IN1(n4405), .IN2(n12905), .Q(n12918) );
  AND2X1 U14404 ( .IN1(g3201), .IN2(n4329), .Q(n12905) );
  AND2X1 U14405 ( .IN1(n3940), .IN2(g3095), .Q(n14167) );
  AND2X1 U14406 ( .IN1(n12904), .IN2(g3142), .Q(n14164) );
  AND2X1 U14407 ( .IN1(n3940), .IN2(n14154), .Q(n12904) );
  OR2X1 U14408 ( .IN1(n14171), .IN2(n14172), .Q(n14162) );
  AND2X1 U14409 ( .IN1(n12909), .IN2(n12917), .Q(n14172) );
  AND2X1 U14410 ( .IN1(n3705), .IN2(n14088), .Q(n12909) );
  AND2X1 U14411 ( .IN1(n14089), .IN2(g3086), .Q(n14171) );
  AND2X1 U14412 ( .IN1(n14088), .IN2(n12919), .Q(n14089) );
  AND2X1 U14413 ( .IN1(g3204), .IN2(n305), .Q(n12919) );
  AND2X1 U14414 ( .IN1(g3197), .IN2(n306), .Q(n305) );
  INVX0 U14415 ( .INP(n14173), .ZN(n306) );
  OR2X1 U14416 ( .IN1(n8088), .IN2(n14174), .Q(n14173) );
  OR2X1 U14417 ( .IN1(n8090), .IN2(n8089), .Q(n14174) );
  OR2X1 U14418 ( .IN1(g3234), .IN2(n14175), .Q(g26048) );
  AND2X1 U14419 ( .IN1(n14176), .IN2(n13724), .Q(n14175) );
  XOR2X1 U14420 ( .IN1(n14177), .IN2(n16493), .Q(n14176) );
  AND2X1 U14421 ( .IN1(n14178), .IN2(n9662), .Q(g26037) );
  AND2X1 U14422 ( .IN1(n14179), .IN2(n13721), .Q(n14178) );
  OR2X1 U14423 ( .IN1(n4291), .IN2(n14180), .Q(n13721) );
  OR2X1 U14424 ( .IN1(n14181), .IN2(g2900), .Q(n14179) );
  AND2X1 U14425 ( .IN1(n13724), .IN2(n14182), .Q(g26031) );
  XNOR2X1 U14426 ( .IN1(test_so98), .IN2(n3742), .Q(n14182) );
  OR2X1 U14427 ( .IN1(n14183), .IN2(n14184), .Q(g26025) );
  AND2X1 U14428 ( .IN1(n13736), .IN2(n10833), .Q(n14184) );
  AND2X1 U14429 ( .IN1(n13738), .IN2(test_so79), .Q(n13736) );
  AND2X1 U14430 ( .IN1(test_so82), .IN2(n14185), .Q(n14183) );
  OR2X1 U14431 ( .IN1(n4509), .IN2(n13738), .Q(n14185) );
  OR2X1 U14432 ( .IN1(n11478), .IN2(n14186), .Q(n13738) );
  OR2X1 U14433 ( .IN1(n11191), .IN2(n9121), .Q(n14186) );
  OR2X1 U14434 ( .IN1(n14187), .IN2(n14188), .Q(n11191) );
  OR2X1 U14435 ( .IN1(n14189), .IN2(n14190), .Q(n14188) );
  OR2X1 U14436 ( .IN1(n14191), .IN2(n14192), .Q(n14190) );
  XNOR2X1 U14437 ( .IN1(n10714), .IN2(n14193), .Q(n14192) );
  AND2X1 U14438 ( .IN1(n14194), .IN2(n14195), .Q(n14193) );
  OR2X1 U14439 ( .IN1(n9119), .IN2(g2237), .Q(n14195) );
  AND2X1 U14440 ( .IN1(n14196), .IN2(n14197), .Q(n14194) );
  OR2X1 U14441 ( .IN1(n4324), .IN2(g2236), .Q(n14197) );
  OR2X1 U14442 ( .IN1(n4367), .IN2(g2235), .Q(n14196) );
  XNOR2X1 U14443 ( .IN1(n4319), .IN2(n14198), .Q(n14191) );
  OR2X1 U14444 ( .IN1(n14199), .IN2(n14200), .Q(n14198) );
  OR2X1 U14445 ( .IN1(n14201), .IN2(n14202), .Q(n14200) );
  AND2X1 U14446 ( .IN1(n8993), .IN2(g6837), .Q(n14202) );
  AND2X1 U14447 ( .IN1(n8992), .IN2(test_so73), .Q(n14201) );
  AND2X1 U14448 ( .IN1(n8632), .IN2(g2241), .Q(n14199) );
  OR2X1 U14449 ( .IN1(n14203), .IN2(n14204), .Q(n14189) );
  OR2X1 U14450 ( .IN1(n14205), .IN2(n14206), .Q(n14204) );
  XNOR2X1 U14451 ( .IN1(n4377), .IN2(n14207), .Q(n14206) );
  OR2X1 U14452 ( .IN1(n14208), .IN2(n14209), .Q(n14207) );
  OR2X1 U14453 ( .IN1(n14210), .IN2(n14211), .Q(n14209) );
  AND2X1 U14454 ( .IN1(n8997), .IN2(g6837), .Q(n14211) );
  AND2X1 U14455 ( .IN1(n8996), .IN2(test_so73), .Q(n14210) );
  AND2X1 U14456 ( .IN1(n8634), .IN2(g2241), .Q(n14208) );
  XNOR2X1 U14457 ( .IN1(n4373), .IN2(n14212), .Q(n14205) );
  OR2X1 U14458 ( .IN1(n14213), .IN2(n14214), .Q(n14212) );
  OR2X1 U14459 ( .IN1(n14215), .IN2(n14216), .Q(n14214) );
  AND2X1 U14460 ( .IN1(n8995), .IN2(g6837), .Q(n14216) );
  AND2X1 U14461 ( .IN1(n8994), .IN2(test_so73), .Q(n14215) );
  AND2X1 U14462 ( .IN1(n8633), .IN2(g2241), .Q(n14213) );
  XNOR2X1 U14463 ( .IN1(n14217), .IN2(n14218), .Q(n14203) );
  AND2X1 U14464 ( .IN1(n14219), .IN2(n14220), .Q(n14218) );
  OR2X1 U14465 ( .IN1(test_so75), .IN2(n9119), .Q(n14220) );
  AND2X1 U14466 ( .IN1(n14221), .IN2(n14222), .Q(n14219) );
  OR2X1 U14467 ( .IN1(n4324), .IN2(g2239), .Q(n14222) );
  OR2X1 U14468 ( .IN1(n4367), .IN2(g2238), .Q(n14221) );
  OR2X1 U14469 ( .IN1(n14223), .IN2(n14224), .Q(n14187) );
  OR2X1 U14470 ( .IN1(n14225), .IN2(n14226), .Q(n14224) );
  OR2X1 U14471 ( .IN1(n14227), .IN2(n14228), .Q(n14226) );
  XNOR2X1 U14472 ( .IN1(g2195), .IN2(n14229), .Q(n14228) );
  AND2X1 U14473 ( .IN1(n14230), .IN2(n14231), .Q(n14229) );
  OR2X1 U14474 ( .IN1(n9119), .IN2(g2231), .Q(n14231) );
  AND2X1 U14475 ( .IN1(n14232), .IN2(n14233), .Q(n14230) );
  OR2X1 U14476 ( .IN1(n4324), .IN2(g2230), .Q(n14233) );
  OR2X1 U14477 ( .IN1(n4367), .IN2(g2229), .Q(n14232) );
  XNOR2X1 U14478 ( .IN1(g2190), .IN2(n14234), .Q(n14227) );
  AND2X1 U14479 ( .IN1(n14235), .IN2(n14236), .Q(n14234) );
  OR2X1 U14480 ( .IN1(n9119), .IN2(g2228), .Q(n14236) );
  AND2X1 U14481 ( .IN1(n14237), .IN2(n14238), .Q(n14235) );
  OR2X1 U14482 ( .IN1(n4324), .IN2(g2227), .Q(n14238) );
  OR2X1 U14483 ( .IN1(n4367), .IN2(g2226), .Q(n14237) );
  XNOR2X1 U14484 ( .IN1(n4389), .IN2(n14239), .Q(n14225) );
  OR2X1 U14485 ( .IN1(n14240), .IN2(n14241), .Q(n14239) );
  OR2X1 U14486 ( .IN1(n14242), .IN2(n14243), .Q(n14241) );
  AND2X1 U14487 ( .IN1(n8991), .IN2(g6837), .Q(n14243) );
  AND2X1 U14488 ( .IN1(n8990), .IN2(test_so73), .Q(n14242) );
  AND2X1 U14489 ( .IN1(n8631), .IN2(g2241), .Q(n14240) );
  OR2X1 U14490 ( .IN1(n14244), .IN2(n14245), .Q(n14223) );
  OR2X1 U14491 ( .IN1(n10857), .IN2(n14246), .Q(n14245) );
  XNOR2X1 U14492 ( .IN1(n4287), .IN2(n14247), .Q(n14246) );
  OR2X1 U14493 ( .IN1(n14248), .IN2(n14249), .Q(n14247) );
  OR2X1 U14494 ( .IN1(n14250), .IN2(n14251), .Q(n14249) );
  AND2X1 U14495 ( .IN1(n8984), .IN2(g6837), .Q(n14251) );
  AND2X1 U14496 ( .IN1(n8983), .IN2(test_so73), .Q(n14250) );
  AND2X1 U14497 ( .IN1(n8627), .IN2(g2241), .Q(n14248) );
  INVX0 U14498 ( .INP(n3038), .ZN(n10857) );
  XNOR2X1 U14499 ( .IN1(n4325), .IN2(n14252), .Q(n14244) );
  OR2X1 U14500 ( .IN1(n14253), .IN2(n14254), .Q(n14252) );
  OR2X1 U14501 ( .IN1(n14255), .IN2(n14256), .Q(n14254) );
  AND2X1 U14502 ( .IN1(n8989), .IN2(g6837), .Q(n14256) );
  INVX0 U14503 ( .INP(n14257), .ZN(n14255) );
  OR2X1 U14504 ( .IN1(n9119), .IN2(test_so74), .Q(n14257) );
  AND2X1 U14505 ( .IN1(n8630), .IN2(g2241), .Q(n14253) );
  OR2X1 U14506 ( .IN1(n14258), .IN2(n14259), .Q(n11478) );
  OR2X1 U14507 ( .IN1(n14260), .IN2(n14261), .Q(n14259) );
  AND2X1 U14508 ( .IN1(n8782), .IN2(n10408), .Q(n14261) );
  INVX0 U14509 ( .INP(n14262), .ZN(n14260) );
  OR2X1 U14510 ( .IN1(n4509), .IN2(test_so82), .Q(n14262) );
  AND2X1 U14511 ( .IN1(n8773), .IN2(n10398), .Q(n14258) );
  AND2X1 U14512 ( .IN1(n14263), .IN2(n4526), .Q(g25940) );
  AND2X1 U14513 ( .IN1(n14264), .IN2(n11527), .Q(n14263) );
  OR2X1 U14514 ( .IN1(n3887), .IN2(test_so78), .Q(n14264) );
  AND2X1 U14515 ( .IN1(n14265), .IN2(n4527), .Q(g25938) );
  AND2X1 U14516 ( .IN1(n14266), .IN2(n11529), .Q(n14265) );
  INVX0 U14517 ( .INP(n14267), .ZN(n14266) );
  AND2X1 U14518 ( .IN1(n10218), .IN2(n9114), .Q(n14267) );
  INVX0 U14519 ( .INP(n3890), .ZN(n10218) );
  AND2X1 U14520 ( .IN1(n14268), .IN2(n14269), .Q(g25935) );
  OR2X1 U14521 ( .IN1(n3893), .IN2(g776), .Q(n14269) );
  AND2X1 U14522 ( .IN1(n11531), .IN2(n710), .Q(n14268) );
  INVX0 U14523 ( .INP(n14057), .ZN(n710) );
  AND2X1 U14524 ( .IN1(g776), .IN2(n3893), .Q(n14057) );
  AND2X1 U14525 ( .IN1(n14270), .IN2(n4528), .Q(g25932) );
  AND2X1 U14526 ( .IN1(n14271), .IN2(n11533), .Q(n14270) );
  INVX0 U14527 ( .INP(n14272), .ZN(n14271) );
  AND2X1 U14528 ( .IN1(n10217), .IN2(n9113), .Q(n14272) );
  INVX0 U14529 ( .INP(n3896), .ZN(n10217) );
  OR2X1 U14530 ( .IN1(n14273), .IN2(n14274), .Q(g25489) );
  AND2X1 U14531 ( .IN1(n14275), .IN2(test_so10), .Q(n14274) );
  AND2X1 U14532 ( .IN1(n14276), .IN2(g3142), .Q(n14275) );
  AND2X1 U14533 ( .IN1(g3151), .IN2(g3097), .Q(n14276) );
  AND2X1 U14534 ( .IN1(n14277), .IN2(n9128), .Q(n14273) );
  OR2X1 U14535 ( .IN1(n14278), .IN2(n14279), .Q(n14277) );
  AND2X1 U14536 ( .IN1(n4301), .IN2(n12917), .Q(n14279) );
  OR2X1 U14537 ( .IN1(test_so1), .IN2(n8099), .Q(n12917) );
  AND2X1 U14538 ( .IN1(n4424), .IN2(n14280), .Q(n14278) );
  OR2X1 U14539 ( .IN1(n4301), .IN2(n12916), .Q(n14280) );
  OR2X1 U14540 ( .IN1(n4577), .IN2(n4578), .Q(n12916) );
  OR2X1 U14541 ( .IN1(n14281), .IN2(n14282), .Q(g25452) );
  AND2X1 U14542 ( .IN1(g21851), .IN2(g3109), .Q(n14282) );
  AND2X1 U14543 ( .IN1(n4494), .IN2(g3099), .Q(n14281) );
  OR2X1 U14544 ( .IN1(n14283), .IN2(n14284), .Q(g25451) );
  AND2X1 U14545 ( .IN1(g21851), .IN2(g8030), .Q(n14284) );
  AND2X1 U14546 ( .IN1(n4383), .IN2(g3098), .Q(n14283) );
  OR2X1 U14547 ( .IN1(n14285), .IN2(n14286), .Q(g25450) );
  AND2X1 U14548 ( .IN1(g21851), .IN2(g8106), .Q(n14286) );
  AND2X1 U14549 ( .IN1(n4382), .IN2(g3097), .Q(n14285) );
  OR2X1 U14550 ( .IN1(n12894), .IN2(n14287), .Q(g25442) );
  OR2X1 U14551 ( .IN1(n14288), .IN2(n14289), .Q(n14287) );
  AND2X1 U14552 ( .IN1(n12898), .IN2(g3124), .Q(n14289) );
  AND2X1 U14553 ( .IN1(n14070), .IN2(g3111), .Q(n14288) );
  OR2X1 U14554 ( .IN1(n12894), .IN2(n14290), .Q(g25435) );
  OR2X1 U14555 ( .IN1(n14291), .IN2(n14292), .Q(n14290) );
  AND2X1 U14556 ( .IN1(n12898), .IN2(DFF_144_n1), .Q(n14292) );
  AND2X1 U14557 ( .IN1(n14070), .IN2(g3110), .Q(n14291) );
  OR2X1 U14558 ( .IN1(n12894), .IN2(n14293), .Q(g25420) );
  OR2X1 U14559 ( .IN1(n14294), .IN2(n14295), .Q(n14293) );
  AND2X1 U14560 ( .IN1(test_so9), .IN2(n12898), .Q(n14295) );
  AND2X1 U14561 ( .IN1(n14070), .IN2(g3112), .Q(n14294) );
  AND2X1 U14562 ( .IN1(n14154), .IN2(n14088), .Q(n14070) );
  AND2X1 U14563 ( .IN1(n4405), .IN2(n14095), .Q(n14088) );
  AND2X1 U14564 ( .IN1(n4329), .IN2(n4406), .Q(n14095) );
  AND2X1 U14565 ( .IN1(g3204), .IN2(n4073), .Q(n14154) );
  OR2X1 U14566 ( .IN1(n14296), .IN2(n14297), .Q(g25288) );
  AND2X1 U14567 ( .IN1(n14298), .IN2(n14299), .Q(n14297) );
  AND2X1 U14568 ( .IN1(n14300), .IN2(g2808), .Q(n14296) );
  OR2X1 U14569 ( .IN1(n14301), .IN2(n14302), .Q(g25280) );
  AND2X1 U14570 ( .IN1(n14303), .IN2(g2810), .Q(n14302) );
  AND2X1 U14571 ( .IN1(n14304), .IN2(n14298), .Q(n14301) );
  OR2X1 U14572 ( .IN1(n14305), .IN2(n14306), .Q(g25279) );
  AND2X1 U14573 ( .IN1(n14307), .IN2(n4149), .Q(n14306) );
  AND2X1 U14574 ( .IN1(n14308), .IN2(g2114), .Q(n14305) );
  OR2X1 U14575 ( .IN1(n14309), .IN2(n14310), .Q(g25272) );
  AND2X1 U14576 ( .IN1(n14311), .IN2(g2809), .Q(n14310) );
  AND2X1 U14577 ( .IN1(n14312), .IN2(n14298), .Q(n14309) );
  INVX0 U14578 ( .INP(n14313), .ZN(n14298) );
  OR2X1 U14579 ( .IN1(n14314), .IN2(n14315), .Q(n14313) );
  OR2X1 U14580 ( .IN1(n14316), .IN2(n10326), .Q(n14315) );
  OR2X1 U14581 ( .IN1(n14317), .IN2(n14318), .Q(n10326) );
  OR2X1 U14582 ( .IN1(n14319), .IN2(n14320), .Q(n14318) );
  AND2X1 U14583 ( .IN1(n8677), .IN2(g7425), .Q(n14320) );
  AND2X1 U14584 ( .IN1(n8732), .IN2(g2703), .Q(n14319) );
  AND2X1 U14585 ( .IN1(n8669), .IN2(g7487), .Q(n14317) );
  AND2X1 U14586 ( .IN1(n8670), .IN2(g7487), .Q(n14316) );
  OR2X1 U14587 ( .IN1(n14321), .IN2(n14322), .Q(n14314) );
  OR2X1 U14588 ( .IN1(n14323), .IN2(n14324), .Q(n14322) );
  AND2X1 U14589 ( .IN1(n8733), .IN2(g2703), .Q(n14324) );
  AND2X1 U14590 ( .IN1(n14325), .IN2(n14326), .Q(n14323) );
  AND2X1 U14591 ( .IN1(n14327), .IN2(n14328), .Q(n14326) );
  AND2X1 U14592 ( .IN1(n14329), .IN2(n14330), .Q(n14328) );
  XNOR2X1 U14593 ( .IN1(n4472), .IN2(n9893), .Q(n14330) );
  INVX0 U14594 ( .INP(n9894), .ZN(n9893) );
  OR2X1 U14595 ( .IN1(n14331), .IN2(n14332), .Q(n9894) );
  OR2X1 U14596 ( .IN1(n14333), .IN2(n14334), .Q(n14332) );
  AND2X1 U14597 ( .IN1(n8884), .IN2(g7425), .Q(n14334) );
  AND2X1 U14598 ( .IN1(n8947), .IN2(g2703), .Q(n14333) );
  AND2X1 U14599 ( .IN1(n8883), .IN2(g7487), .Q(n14331) );
  AND2X1 U14600 ( .IN1(n14335), .IN2(n14336), .Q(n14329) );
  XNOR2X1 U14601 ( .IN1(n9122), .IN2(n9917), .Q(n14336) );
  INVX0 U14602 ( .INP(n9916), .ZN(n9917) );
  OR2X1 U14603 ( .IN1(n14337), .IN2(n14338), .Q(n9916) );
  OR2X1 U14604 ( .IN1(n14339), .IN2(n14340), .Q(n14338) );
  AND2X1 U14605 ( .IN1(n8874), .IN2(g7425), .Q(n14340) );
  AND2X1 U14606 ( .IN1(n8943), .IN2(g2703), .Q(n14339) );
  AND2X1 U14607 ( .IN1(n8873), .IN2(g7487), .Q(n14337) );
  XOR2X1 U14608 ( .IN1(n4398), .IN2(n9921), .Q(n14335) );
  OR2X1 U14609 ( .IN1(n14341), .IN2(n14342), .Q(n9921) );
  OR2X1 U14610 ( .IN1(n14343), .IN2(n14344), .Q(n14342) );
  AND2X1 U14611 ( .IN1(n8886), .IN2(g7425), .Q(n14344) );
  AND2X1 U14612 ( .IN1(n8948), .IN2(g2703), .Q(n14343) );
  AND2X1 U14613 ( .IN1(n8885), .IN2(g7487), .Q(n14341) );
  AND2X1 U14614 ( .IN1(n14345), .IN2(n14346), .Q(n14327) );
  XOR2X1 U14615 ( .IN1(n4397), .IN2(n9887), .Q(n14346) );
  OR2X1 U14616 ( .IN1(n14347), .IN2(n14348), .Q(n9887) );
  OR2X1 U14617 ( .IN1(n14349), .IN2(n14350), .Q(n14348) );
  AND2X1 U14618 ( .IN1(n8878), .IN2(g7425), .Q(n14350) );
  AND2X1 U14619 ( .IN1(n8945), .IN2(g2703), .Q(n14349) );
  AND2X1 U14620 ( .IN1(n8877), .IN2(g7487), .Q(n14347) );
  XOR2X1 U14621 ( .IN1(n4407), .IN2(n9906), .Q(n14345) );
  OR2X1 U14622 ( .IN1(n14351), .IN2(n14352), .Q(n9906) );
  OR2X1 U14623 ( .IN1(n14353), .IN2(n14354), .Q(n14352) );
  AND2X1 U14624 ( .IN1(n8876), .IN2(g7425), .Q(n14354) );
  AND2X1 U14625 ( .IN1(n8944), .IN2(g2703), .Q(n14353) );
  AND2X1 U14626 ( .IN1(n8875), .IN2(g7487), .Q(n14351) );
  AND2X1 U14627 ( .IN1(n14355), .IN2(n14356), .Q(n14325) );
  AND2X1 U14628 ( .IN1(n14357), .IN2(n14358), .Q(n14356) );
  XOR2X1 U14629 ( .IN1(n4471), .IN2(n9899), .Q(n14358) );
  OR2X1 U14630 ( .IN1(n14359), .IN2(n14360), .Q(n9899) );
  OR2X1 U14631 ( .IN1(n14361), .IN2(n14362), .Q(n14360) );
  AND2X1 U14632 ( .IN1(n8872), .IN2(g7425), .Q(n14362) );
  AND2X1 U14633 ( .IN1(n8942), .IN2(g2703), .Q(n14361) );
  AND2X1 U14634 ( .IN1(n8871), .IN2(g7487), .Q(n14359) );
  AND2X1 U14635 ( .IN1(n14363), .IN2(n14364), .Q(n14357) );
  XNOR2X1 U14636 ( .IN1(n4415), .IN2(n9934), .Q(n14364) );
  INVX0 U14637 ( .INP(n9935), .ZN(n9934) );
  OR2X1 U14638 ( .IN1(n14365), .IN2(n14366), .Q(n9935) );
  OR2X1 U14639 ( .IN1(n14367), .IN2(n14368), .Q(n14366) );
  AND2X1 U14640 ( .IN1(n8868), .IN2(g7425), .Q(n14368) );
  AND2X1 U14641 ( .IN1(n8941), .IN2(g2703), .Q(n14367) );
  AND2X1 U14642 ( .IN1(n8867), .IN2(g7487), .Q(n14365) );
  XNOR2X1 U14643 ( .IN1(n4393), .IN2(n9947), .Q(n14363) );
  INVX0 U14644 ( .INP(n9945), .ZN(n9947) );
  OR2X1 U14645 ( .IN1(n14369), .IN2(n14370), .Q(n9945) );
  OR2X1 U14646 ( .IN1(n14371), .IN2(n14372), .Q(n14370) );
  AND2X1 U14647 ( .IN1(n8870), .IN2(g7425), .Q(n14372) );
  INVX0 U14648 ( .INP(n14373), .ZN(n14371) );
  OR2X1 U14649 ( .IN1(n4292), .IN2(test_so94), .Q(n14373) );
  AND2X1 U14650 ( .IN1(n8869), .IN2(g7487), .Q(n14369) );
  AND2X1 U14651 ( .IN1(n14374), .IN2(n14375), .Q(n14355) );
  XNOR2X1 U14652 ( .IN1(n4408), .IN2(n9878), .Q(n14375) );
  INVX0 U14653 ( .INP(n9881), .ZN(n9878) );
  OR2X1 U14654 ( .IN1(n14376), .IN2(n14377), .Q(n9881) );
  OR2X1 U14655 ( .IN1(n14378), .IN2(n14379), .Q(n14377) );
  AND2X1 U14656 ( .IN1(n8880), .IN2(g7425), .Q(n14379) );
  INVX0 U14657 ( .INP(n14380), .ZN(n14378) );
  OR2X1 U14658 ( .IN1(n4292), .IN2(test_so93), .Q(n14380) );
  AND2X1 U14659 ( .IN1(n8879), .IN2(g7487), .Q(n14376) );
  XNOR2X1 U14660 ( .IN1(n4419), .IN2(n9912), .Q(n14374) );
  INVX0 U14661 ( .INP(n9911), .ZN(n9912) );
  OR2X1 U14662 ( .IN1(n14381), .IN2(n14382), .Q(n9911) );
  OR2X1 U14663 ( .IN1(n14383), .IN2(n14384), .Q(n14382) );
  AND2X1 U14664 ( .IN1(n8882), .IN2(g7425), .Q(n14384) );
  AND2X1 U14665 ( .IN1(n8946), .IN2(g2703), .Q(n14383) );
  AND2X1 U14666 ( .IN1(n8881), .IN2(g7487), .Q(n14381) );
  AND2X1 U14667 ( .IN1(n8678), .IN2(g7425), .Q(n14321) );
  OR2X1 U14668 ( .IN1(n14385), .IN2(n14386), .Q(g25271) );
  AND2X1 U14669 ( .IN1(n14387), .IN2(n14307), .Q(n14386) );
  AND2X1 U14670 ( .IN1(n14388), .IN2(g2116), .Q(n14385) );
  OR2X1 U14671 ( .IN1(n14389), .IN2(n14390), .Q(g25270) );
  AND2X1 U14672 ( .IN1(n14391), .IN2(n14392), .Q(n14390) );
  AND2X1 U14673 ( .IN1(n14393), .IN2(g1420), .Q(n14389) );
  OR2X1 U14674 ( .IN1(n14394), .IN2(n14395), .Q(g25268) );
  AND2X1 U14675 ( .IN1(n14396), .IN2(n14307), .Q(n14395) );
  INVX0 U14676 ( .INP(n14397), .ZN(n14307) );
  OR2X1 U14677 ( .IN1(n14398), .IN2(n14399), .Q(n14397) );
  OR2X1 U14678 ( .IN1(n14400), .IN2(n10355), .Q(n14399) );
  OR2X1 U14679 ( .IN1(n14401), .IN2(n14402), .Q(n10355) );
  OR2X1 U14680 ( .IN1(n14403), .IN2(n14404), .Q(n14402) );
  AND2X1 U14681 ( .IN1(n8679), .IN2(g7229), .Q(n14404) );
  AND2X1 U14682 ( .IN1(n8734), .IN2(g2009), .Q(n14403) );
  AND2X1 U14683 ( .IN1(n8671), .IN2(g7357), .Q(n14401) );
  AND2X1 U14684 ( .IN1(n8672), .IN2(g7357), .Q(n14400) );
  OR2X1 U14685 ( .IN1(n14405), .IN2(n14406), .Q(n14398) );
  OR2X1 U14686 ( .IN1(n14407), .IN2(n14408), .Q(n14406) );
  AND2X1 U14687 ( .IN1(n8735), .IN2(g2009), .Q(n14408) );
  AND2X1 U14688 ( .IN1(n14409), .IN2(n14410), .Q(n14407) );
  AND2X1 U14689 ( .IN1(n14411), .IN2(n14412), .Q(n14410) );
  AND2X1 U14690 ( .IN1(n14413), .IN2(n14414), .Q(n14412) );
  XNOR2X1 U14691 ( .IN1(n4474), .IN2(n10027), .Q(n14414) );
  INVX0 U14692 ( .INP(n10028), .ZN(n10027) );
  OR2X1 U14693 ( .IN1(n14415), .IN2(n14416), .Q(n10028) );
  OR2X1 U14694 ( .IN1(n14417), .IN2(n14418), .Q(n14416) );
  AND2X1 U14695 ( .IN1(n8902), .IN2(g7229), .Q(n14418) );
  AND2X1 U14696 ( .IN1(n8957), .IN2(g2009), .Q(n14417) );
  AND2X1 U14697 ( .IN1(n8901), .IN2(g7357), .Q(n14415) );
  AND2X1 U14698 ( .IN1(n14419), .IN2(n14420), .Q(n14413) );
  XNOR2X1 U14699 ( .IN1(n9124), .IN2(n10080), .Q(n14420) );
  INVX0 U14700 ( .INP(n10078), .ZN(n10080) );
  OR2X1 U14701 ( .IN1(n14421), .IN2(n14422), .Q(n10078) );
  OR2X1 U14702 ( .IN1(n14423), .IN2(n14424), .Q(n14422) );
  AND2X1 U14703 ( .IN1(n8889), .IN2(g7229), .Q(n14424) );
  AND2X1 U14704 ( .IN1(n8950), .IN2(g2009), .Q(n14423) );
  AND2X1 U14705 ( .IN1(n8888), .IN2(g7357), .Q(n14421) );
  XOR2X1 U14706 ( .IN1(n4473), .IN2(n10033), .Q(n14419) );
  OR2X1 U14707 ( .IN1(n14425), .IN2(n14426), .Q(n10033) );
  OR2X1 U14708 ( .IN1(n14427), .IN2(n14428), .Q(n14426) );
  AND2X1 U14709 ( .IN1(n8891), .IN2(g7229), .Q(n14428) );
  AND2X1 U14710 ( .IN1(n8951), .IN2(g2009), .Q(n14427) );
  AND2X1 U14711 ( .IN1(n8890), .IN2(g7357), .Q(n14425) );
  AND2X1 U14712 ( .IN1(n14429), .IN2(n14430), .Q(n14411) );
  XOR2X1 U14713 ( .IN1(n4468), .IN2(n10050), .Q(n14430) );
  OR2X1 U14714 ( .IN1(n14431), .IN2(n14432), .Q(n10050) );
  OR2X1 U14715 ( .IN1(n14433), .IN2(n14434), .Q(n14432) );
  AND2X1 U14716 ( .IN1(n8893), .IN2(g7229), .Q(n14434) );
  AND2X1 U14717 ( .IN1(n8952), .IN2(g2009), .Q(n14433) );
  AND2X1 U14718 ( .IN1(n8892), .IN2(g7357), .Q(n14431) );
  XNOR2X1 U14719 ( .IN1(n4410), .IN2(n10012), .Q(n14429) );
  INVX0 U14720 ( .INP(n10015), .ZN(n10012) );
  OR2X1 U14721 ( .IN1(n14435), .IN2(n14436), .Q(n10015) );
  OR2X1 U14722 ( .IN1(n14437), .IN2(n14438), .Q(n14436) );
  AND2X1 U14723 ( .IN1(n8898), .IN2(g7229), .Q(n14438) );
  AND2X1 U14724 ( .IN1(n8955), .IN2(g2009), .Q(n14437) );
  AND2X1 U14725 ( .IN1(n8897), .IN2(g7357), .Q(n14435) );
  AND2X1 U14726 ( .IN1(n14439), .IN2(n14440), .Q(n14409) );
  AND2X1 U14727 ( .IN1(n14441), .IN2(n14442), .Q(n14440) );
  XNOR2X1 U14728 ( .IN1(n4399), .IN2(n10022), .Q(n14442) );
  AND2X1 U14729 ( .IN1(n14443), .IN2(n14444), .Q(n10022) );
  INVX0 U14730 ( .INP(n14445), .ZN(n14444) );
  OR2X1 U14731 ( .IN1(n14446), .IN2(n14447), .Q(n14445) );
  AND2X1 U14732 ( .IN1(n8896), .IN2(g7229), .Q(n14447) );
  AND2X1 U14733 ( .IN1(n8954), .IN2(g2009), .Q(n14446) );
  OR2X1 U14734 ( .IN1(n4357), .IN2(test_so71), .Q(n14443) );
  AND2X1 U14735 ( .IN1(n14448), .IN2(n14449), .Q(n14441) );
  XNOR2X1 U14736 ( .IN1(n4416), .IN2(n10068), .Q(n14449) );
  INVX0 U14737 ( .INP(n10069), .ZN(n10068) );
  OR2X1 U14738 ( .IN1(n14450), .IN2(n14451), .Q(n10069) );
  OR2X1 U14739 ( .IN1(n14452), .IN2(n14453), .Q(n14451) );
  AND2X1 U14740 ( .IN1(n8887), .IN2(g7229), .Q(n14453) );
  AND2X1 U14741 ( .IN1(n8949), .IN2(g2009), .Q(n14452) );
  INVX0 U14742 ( .INP(n14454), .ZN(n14450) );
  OR2X1 U14743 ( .IN1(n4357), .IN2(test_so72), .Q(n14454) );
  XOR2X1 U14744 ( .IN1(n4409), .IN2(n10040), .Q(n14448) );
  OR2X1 U14745 ( .IN1(n14455), .IN2(n14456), .Q(n10040) );
  OR2X1 U14746 ( .IN1(n14457), .IN2(n14458), .Q(n14456) );
  AND2X1 U14747 ( .IN1(n8895), .IN2(g7229), .Q(n14458) );
  AND2X1 U14748 ( .IN1(n8953), .IN2(g2009), .Q(n14457) );
  AND2X1 U14749 ( .IN1(n8894), .IN2(g7357), .Q(n14455) );
  AND2X1 U14750 ( .IN1(n14459), .IN2(n14460), .Q(n14439) );
  XOR2X1 U14751 ( .IN1(n4400), .IN2(n10055), .Q(n14460) );
  OR2X1 U14752 ( .IN1(n14461), .IN2(n14462), .Q(n10055) );
  OR2X1 U14753 ( .IN1(n14463), .IN2(n14464), .Q(n14462) );
  AND2X1 U14754 ( .IN1(n8904), .IN2(g7229), .Q(n14464) );
  AND2X1 U14755 ( .IN1(n8958), .IN2(g2009), .Q(n14463) );
  AND2X1 U14756 ( .IN1(n8903), .IN2(g7357), .Q(n14461) );
  XNOR2X1 U14757 ( .IN1(n4420), .IN2(n10046), .Q(n14459) );
  INVX0 U14758 ( .INP(n10045), .ZN(n10046) );
  OR2X1 U14759 ( .IN1(n14465), .IN2(n14466), .Q(n10045) );
  OR2X1 U14760 ( .IN1(n14467), .IN2(n14468), .Q(n14466) );
  AND2X1 U14761 ( .IN1(n8900), .IN2(g7229), .Q(n14468) );
  AND2X1 U14762 ( .IN1(n8956), .IN2(g2009), .Q(n14467) );
  AND2X1 U14763 ( .IN1(n8899), .IN2(g7357), .Q(n14465) );
  AND2X1 U14764 ( .IN1(n8680), .IN2(g7229), .Q(n14405) );
  AND2X1 U14765 ( .IN1(n14469), .IN2(g2115), .Q(n14394) );
  OR2X1 U14766 ( .IN1(n14470), .IN2(n14471), .Q(g25267) );
  AND2X1 U14767 ( .IN1(n869), .IN2(n14391), .Q(n14471) );
  AND2X1 U14768 ( .IN1(n14472), .IN2(g1422), .Q(n14470) );
  OR2X1 U14769 ( .IN1(n14473), .IN2(n14474), .Q(g25266) );
  AND2X1 U14770 ( .IN1(n14475), .IN2(n590), .Q(n14474) );
  AND2X1 U14771 ( .IN1(n14476), .IN2(g734), .Q(n14473) );
  OR2X1 U14772 ( .IN1(n14477), .IN2(n14478), .Q(g25265) );
  AND2X1 U14773 ( .IN1(n14479), .IN2(n13724), .Q(n14478) );
  XNOR2X1 U14774 ( .IN1(g2993), .IN2(n9094), .Q(n14479) );
  INVX0 U14775 ( .INP(n14480), .ZN(n14477) );
  OR2X1 U14776 ( .IN1(n13724), .IN2(g3234), .Q(n14480) );
  OR2X1 U14777 ( .IN1(n14481), .IN2(n14482), .Q(g25263) );
  AND2X1 U14778 ( .IN1(n14483), .IN2(g1421), .Q(n14482) );
  AND2X1 U14779 ( .IN1(n14484), .IN2(n14391), .Q(n14481) );
  INVX0 U14780 ( .INP(n14485), .ZN(n14391) );
  OR2X1 U14781 ( .IN1(n14486), .IN2(n14487), .Q(n14485) );
  OR2X1 U14782 ( .IN1(n14488), .IN2(n10380), .Q(n14487) );
  OR2X1 U14783 ( .IN1(n14489), .IN2(n14490), .Q(n10380) );
  OR2X1 U14784 ( .IN1(n14491), .IN2(n14492), .Q(n14490) );
  AND2X1 U14785 ( .IN1(n8681), .IN2(g6979), .Q(n14492) );
  AND2X1 U14786 ( .IN1(n8736), .IN2(g1315), .Q(n14491) );
  AND2X1 U14787 ( .IN1(n8673), .IN2(g7161), .Q(n14489) );
  AND2X1 U14788 ( .IN1(n8674), .IN2(g7161), .Q(n14488) );
  OR2X1 U14789 ( .IN1(n14493), .IN2(n14494), .Q(n14486) );
  OR2X1 U14790 ( .IN1(n14495), .IN2(n14496), .Q(n14494) );
  INVX0 U14791 ( .INP(n14497), .ZN(n14496) );
  OR2X1 U14792 ( .IN1(n4294), .IN2(test_so51), .Q(n14497) );
  AND2X1 U14793 ( .IN1(n14498), .IN2(n14499), .Q(n14495) );
  AND2X1 U14794 ( .IN1(n14500), .IN2(n14501), .Q(n14499) );
  AND2X1 U14795 ( .IN1(n14502), .IN2(n14503), .Q(n14501) );
  XOR2X1 U14796 ( .IN1(n4475), .IN2(n10168), .Q(n14503) );
  OR2X1 U14797 ( .IN1(n14504), .IN2(n14505), .Q(n10168) );
  OR2X1 U14798 ( .IN1(n14506), .IN2(n14507), .Q(n14505) );
  AND2X1 U14799 ( .IN1(n8910), .IN2(g6979), .Q(n14507) );
  AND2X1 U14800 ( .IN1(n8961), .IN2(g1315), .Q(n14506) );
  AND2X1 U14801 ( .IN1(n8909), .IN2(g7161), .Q(n14504) );
  AND2X1 U14802 ( .IN1(n14508), .IN2(n14509), .Q(n14502) );
  XOR2X1 U14803 ( .IN1(n4469), .IN2(n10185), .Q(n14509) );
  OR2X1 U14804 ( .IN1(n14510), .IN2(n14511), .Q(n10185) );
  OR2X1 U14805 ( .IN1(n14512), .IN2(n14513), .Q(n14511) );
  AND2X1 U14806 ( .IN1(n8912), .IN2(g6979), .Q(n14513) );
  AND2X1 U14807 ( .IN1(n8962), .IN2(g1315), .Q(n14512) );
  AND2X1 U14808 ( .IN1(n8911), .IN2(g7161), .Q(n14510) );
  XNOR2X1 U14809 ( .IN1(n4476), .IN2(n10162), .Q(n14508) );
  INVX0 U14810 ( .INP(n10163), .ZN(n10162) );
  OR2X1 U14811 ( .IN1(n14514), .IN2(n14515), .Q(n10163) );
  OR2X1 U14812 ( .IN1(n14516), .IN2(n14517), .Q(n14515) );
  AND2X1 U14813 ( .IN1(n8921), .IN2(g6979), .Q(n14517) );
  AND2X1 U14814 ( .IN1(n8967), .IN2(g1315), .Q(n14516) );
  AND2X1 U14815 ( .IN1(n8920), .IN2(g7161), .Q(n14514) );
  AND2X1 U14816 ( .IN1(n14518), .IN2(n14519), .Q(n14500) );
  XNOR2X1 U14817 ( .IN1(n4412), .IN2(n10147), .Q(n14519) );
  INVX0 U14818 ( .INP(n10150), .ZN(n10147) );
  OR2X1 U14819 ( .IN1(n14520), .IN2(n14521), .Q(n10150) );
  OR2X1 U14820 ( .IN1(n14522), .IN2(n14523), .Q(n14521) );
  AND2X1 U14821 ( .IN1(n8917), .IN2(g6979), .Q(n14523) );
  AND2X1 U14822 ( .IN1(n8965), .IN2(g1315), .Q(n14522) );
  AND2X1 U14823 ( .IN1(n8916), .IN2(g7161), .Q(n14520) );
  XNOR2X1 U14824 ( .IN1(n4417), .IN2(n10203), .Q(n14518) );
  INVX0 U14825 ( .INP(n10204), .ZN(n10203) );
  OR2X1 U14826 ( .IN1(n14524), .IN2(n14525), .Q(n10204) );
  OR2X1 U14827 ( .IN1(n14526), .IN2(n14527), .Q(n14525) );
  AND2X1 U14828 ( .IN1(n8906), .IN2(g6979), .Q(n14527) );
  AND2X1 U14829 ( .IN1(n8959), .IN2(g1315), .Q(n14526) );
  AND2X1 U14830 ( .IN1(n8905), .IN2(g7161), .Q(n14524) );
  AND2X1 U14831 ( .IN1(n14528), .IN2(n14529), .Q(n14498) );
  AND2X1 U14832 ( .IN1(n14530), .IN2(n14531), .Q(n14529) );
  XOR2X1 U14833 ( .IN1(n4401), .IN2(n10156), .Q(n14531) );
  OR2X1 U14834 ( .IN1(n14532), .IN2(n14533), .Q(n10156) );
  OR2X1 U14835 ( .IN1(n14534), .IN2(n14535), .Q(n14533) );
  AND2X1 U14836 ( .IN1(n8915), .IN2(g6979), .Q(n14535) );
  AND2X1 U14837 ( .IN1(n8964), .IN2(g1315), .Q(n14534) );
  AND2X1 U14838 ( .IN1(n8914), .IN2(g7161), .Q(n14532) );
  AND2X1 U14839 ( .IN1(n14536), .IN2(n14537), .Q(n14530) );
  XNOR2X1 U14840 ( .IN1(n4395), .IN2(n10215), .Q(n14537) );
  INVX0 U14841 ( .INP(n10213), .ZN(n10215) );
  OR2X1 U14842 ( .IN1(n14538), .IN2(n14539), .Q(n10213) );
  OR2X1 U14843 ( .IN1(n14540), .IN2(n14541), .Q(n14539) );
  AND2X1 U14844 ( .IN1(n8908), .IN2(g6979), .Q(n14541) );
  AND2X1 U14845 ( .IN1(n8960), .IN2(g1315), .Q(n14540) );
  AND2X1 U14846 ( .IN1(n8907), .IN2(g7161), .Q(n14538) );
  XNOR2X1 U14847 ( .IN1(n4411), .IN2(n10174), .Q(n14536) );
  AND2X1 U14848 ( .IN1(n14542), .IN2(n14543), .Q(n10174) );
  INVX0 U14849 ( .INP(n14544), .ZN(n14543) );
  OR2X1 U14850 ( .IN1(n14545), .IN2(n14546), .Q(n14544) );
  AND2X1 U14851 ( .IN1(n8913), .IN2(g6979), .Q(n14546) );
  AND2X1 U14852 ( .IN1(n8963), .IN2(g1315), .Q(n14545) );
  OR2X1 U14853 ( .IN1(n4358), .IN2(test_so50), .Q(n14542) );
  AND2X1 U14854 ( .IN1(n14547), .IN2(n14548), .Q(n14528) );
  XOR2X1 U14855 ( .IN1(n4402), .IN2(n10190), .Q(n14548) );
  OR2X1 U14856 ( .IN1(n14549), .IN2(n14550), .Q(n10190) );
  OR2X1 U14857 ( .IN1(n14551), .IN2(n14552), .Q(n14550) );
  INVX0 U14858 ( .INP(n14553), .ZN(n14552) );
  OR2X1 U14859 ( .IN1(n4308), .IN2(test_so49), .Q(n14553) );
  AND2X1 U14860 ( .IN1(n8968), .IN2(g1315), .Q(n14551) );
  AND2X1 U14861 ( .IN1(n8922), .IN2(g7161), .Q(n14549) );
  XNOR2X1 U14862 ( .IN1(n4421), .IN2(n10181), .Q(n14547) );
  INVX0 U14863 ( .INP(n10180), .ZN(n10181) );
  OR2X1 U14864 ( .IN1(n14554), .IN2(n14555), .Q(n10180) );
  OR2X1 U14865 ( .IN1(n14556), .IN2(n14557), .Q(n14555) );
  AND2X1 U14866 ( .IN1(n8919), .IN2(g6979), .Q(n14557) );
  AND2X1 U14867 ( .IN1(n8966), .IN2(g1315), .Q(n14556) );
  AND2X1 U14868 ( .IN1(n8918), .IN2(g7161), .Q(n14554) );
  AND2X1 U14869 ( .IN1(n8682), .IN2(g6979), .Q(n14493) );
  OR2X1 U14870 ( .IN1(n14558), .IN2(n14559), .Q(g25262) );
  AND2X1 U14871 ( .IN1(n14560), .IN2(g736), .Q(n14559) );
  AND2X1 U14872 ( .IN1(n14561), .IN2(n14475), .Q(n14558) );
  OR2X1 U14873 ( .IN1(n14562), .IN2(n14563), .Q(g25260) );
  AND2X1 U14874 ( .IN1(n14564), .IN2(g735), .Q(n14563) );
  AND2X1 U14875 ( .IN1(n14565), .IN2(n14475), .Q(n14562) );
  INVX0 U14876 ( .INP(n14566), .ZN(n14475) );
  OR2X1 U14877 ( .IN1(n14567), .IN2(n14568), .Q(n14566) );
  OR2X1 U14878 ( .IN1(n14569), .IN2(n10303), .Q(n14568) );
  OR2X1 U14879 ( .IN1(n14570), .IN2(n14571), .Q(n10303) );
  OR2X1 U14880 ( .IN1(n14572), .IN2(n14573), .Q(n14571) );
  AND2X1 U14881 ( .IN1(n8683), .IN2(g6677), .Q(n14573) );
  AND2X1 U14882 ( .IN1(n8737), .IN2(g629), .Q(n14572) );
  AND2X1 U14883 ( .IN1(n8675), .IN2(g6911), .Q(n14570) );
  AND2X1 U14884 ( .IN1(n8676), .IN2(g6911), .Q(n14569) );
  OR2X1 U14885 ( .IN1(n14574), .IN2(n14575), .Q(n14567) );
  OR2X1 U14886 ( .IN1(n14576), .IN2(n14577), .Q(n14575) );
  AND2X1 U14887 ( .IN1(n8738), .IN2(g629), .Q(n14577) );
  AND2X1 U14888 ( .IN1(n14578), .IN2(n14579), .Q(n14576) );
  AND2X1 U14889 ( .IN1(n14580), .IN2(n14581), .Q(n14579) );
  AND2X1 U14890 ( .IN1(n14582), .IN2(n14583), .Q(n14581) );
  XNOR2X1 U14891 ( .IN1(n4478), .IN2(n9803), .Q(n14583) );
  INVX0 U14892 ( .INP(n9804), .ZN(n9803) );
  OR2X1 U14893 ( .IN1(n14584), .IN2(n14585), .Q(n9804) );
  OR2X1 U14894 ( .IN1(n14586), .IN2(n14587), .Q(n14585) );
  AND2X1 U14895 ( .IN1(n8938), .IN2(g6677), .Q(n14587) );
  AND2X1 U14896 ( .IN1(n8977), .IN2(g629), .Q(n14586) );
  AND2X1 U14897 ( .IN1(n8937), .IN2(g6911), .Q(n14584) );
  AND2X1 U14898 ( .IN1(n14588), .IN2(n14589), .Q(n14582) );
  XNOR2X1 U14899 ( .IN1(n9123), .IN2(n9774), .Q(n14589) );
  INVX0 U14900 ( .INP(n9773), .ZN(n9774) );
  OR2X1 U14901 ( .IN1(n14590), .IN2(n14591), .Q(n9773) );
  OR2X1 U14902 ( .IN1(n14592), .IN2(n14593), .Q(n14591) );
  AND2X1 U14903 ( .IN1(n8929), .IN2(g6677), .Q(n14593) );
  AND2X1 U14904 ( .IN1(n8972), .IN2(g629), .Q(n14592) );
  AND2X1 U14905 ( .IN1(n8928), .IN2(g6911), .Q(n14590) );
  XOR2X1 U14906 ( .IN1(n4404), .IN2(n9785), .Q(n14588) );
  OR2X1 U14907 ( .IN1(n14594), .IN2(n14595), .Q(n9785) );
  OR2X1 U14908 ( .IN1(n14596), .IN2(n14597), .Q(n14595) );
  AND2X1 U14909 ( .IN1(n8940), .IN2(g6677), .Q(n14597) );
  AND2X1 U14910 ( .IN1(n8978), .IN2(g629), .Q(n14596) );
  AND2X1 U14911 ( .IN1(n8939), .IN2(g6911), .Q(n14594) );
  AND2X1 U14912 ( .IN1(n14598), .IN2(n14599), .Q(n14580) );
  XOR2X1 U14913 ( .IN1(n4403), .IN2(n9763), .Q(n14599) );
  OR2X1 U14914 ( .IN1(n14600), .IN2(n14601), .Q(n9763) );
  OR2X1 U14915 ( .IN1(n14602), .IN2(n14603), .Q(n14601) );
  INVX0 U14916 ( .INP(n14604), .ZN(n14603) );
  OR2X1 U14917 ( .IN1(n4309), .IN2(test_so29), .Q(n14604) );
  AND2X1 U14918 ( .IN1(n8974), .IN2(g629), .Q(n14602) );
  AND2X1 U14919 ( .IN1(n8932), .IN2(g6911), .Q(n14600) );
  XOR2X1 U14920 ( .IN1(n4413), .IN2(n9779), .Q(n14598) );
  OR2X1 U14921 ( .IN1(n14605), .IN2(n14606), .Q(n9779) );
  OR2X1 U14922 ( .IN1(n14607), .IN2(n14608), .Q(n14606) );
  AND2X1 U14923 ( .IN1(n8931), .IN2(g6677), .Q(n14608) );
  AND2X1 U14924 ( .IN1(n8973), .IN2(g629), .Q(n14607) );
  AND2X1 U14925 ( .IN1(n8930), .IN2(g6911), .Q(n14605) );
  AND2X1 U14926 ( .IN1(n14609), .IN2(n14610), .Q(n14578) );
  AND2X1 U14927 ( .IN1(n14611), .IN2(n14612), .Q(n14610) );
  XOR2X1 U14928 ( .IN1(n4477), .IN2(n9791), .Q(n14612) );
  OR2X1 U14929 ( .IN1(n14613), .IN2(n14614), .Q(n9791) );
  OR2X1 U14930 ( .IN1(n14615), .IN2(n14616), .Q(n14614) );
  AND2X1 U14931 ( .IN1(n8927), .IN2(g6677), .Q(n14616) );
  AND2X1 U14932 ( .IN1(n8971), .IN2(g629), .Q(n14615) );
  AND2X1 U14933 ( .IN1(n8926), .IN2(g6911), .Q(n14613) );
  AND2X1 U14934 ( .IN1(n14617), .IN2(n14618), .Q(n14611) );
  XNOR2X1 U14935 ( .IN1(n4418), .IN2(n9743), .Q(n14618) );
  INVX0 U14936 ( .INP(n9746), .ZN(n9743) );
  OR2X1 U14937 ( .IN1(n14619), .IN2(n14620), .Q(n9746) );
  OR2X1 U14938 ( .IN1(n14621), .IN2(n14622), .Q(n14620) );
  AND2X1 U14939 ( .IN1(n8923), .IN2(g6677), .Q(n14622) );
  AND2X1 U14940 ( .IN1(n8969), .IN2(g629), .Q(n14621) );
  INVX0 U14941 ( .INP(n14623), .ZN(n14619) );
  OR2X1 U14942 ( .IN1(n4359), .IN2(test_so30), .Q(n14623) );
  XNOR2X1 U14943 ( .IN1(n4396), .IN2(n9737), .Q(n14617) );
  INVX0 U14944 ( .INP(n9736), .ZN(n9737) );
  OR2X1 U14945 ( .IN1(n14624), .IN2(n14625), .Q(n9736) );
  OR2X1 U14946 ( .IN1(n14626), .IN2(n14627), .Q(n14625) );
  AND2X1 U14947 ( .IN1(n8925), .IN2(g6677), .Q(n14627) );
  AND2X1 U14948 ( .IN1(n8970), .IN2(g629), .Q(n14626) );
  AND2X1 U14949 ( .IN1(n8924), .IN2(g6911), .Q(n14624) );
  AND2X1 U14950 ( .IN1(n14628), .IN2(n14629), .Q(n14609) );
  XNOR2X1 U14951 ( .IN1(n4414), .IN2(n9768), .Q(n14629) );
  INVX0 U14952 ( .INP(n9769), .ZN(n9768) );
  OR2X1 U14953 ( .IN1(n14630), .IN2(n14631), .Q(n9769) );
  OR2X1 U14954 ( .IN1(n14632), .IN2(n14633), .Q(n14631) );
  AND2X1 U14955 ( .IN1(n8934), .IN2(g6677), .Q(n14633) );
  AND2X1 U14956 ( .IN1(n8975), .IN2(g629), .Q(n14632) );
  AND2X1 U14957 ( .IN1(n8933), .IN2(g6911), .Q(n14630) );
  XNOR2X1 U14958 ( .IN1(n4422), .IN2(n9799), .Q(n14628) );
  INVX0 U14959 ( .INP(n9796), .ZN(n9799) );
  OR2X1 U14960 ( .IN1(n14634), .IN2(n14635), .Q(n9796) );
  OR2X1 U14961 ( .IN1(n14636), .IN2(n14637), .Q(n14635) );
  AND2X1 U14962 ( .IN1(n8936), .IN2(g6677), .Q(n14637) );
  AND2X1 U14963 ( .IN1(n8976), .IN2(g629), .Q(n14636) );
  AND2X1 U14964 ( .IN1(n8935), .IN2(g6911), .Q(n14634) );
  AND2X1 U14965 ( .IN1(n8684), .IN2(g6677), .Q(n14574) );
  OR2X1 U14966 ( .IN1(n14638), .IN2(n14639), .Q(g25259) );
  AND2X1 U14967 ( .IN1(n14640), .IN2(n12102), .Q(n14639) );
  INVX0 U14968 ( .INP(n14641), .ZN(n14638) );
  OR2X1 U14969 ( .IN1(n14640), .IN2(n8685), .Q(n14641) );
  OR2X1 U14970 ( .IN1(n14642), .IN2(n14643), .Q(g25257) );
  AND2X1 U14971 ( .IN1(n9117), .IN2(n12102), .Q(n14643) );
  INVX0 U14972 ( .INP(n14644), .ZN(n14642) );
  OR2X1 U14973 ( .IN1(n9117), .IN2(n8686), .Q(n14644) );
  OR2X1 U14974 ( .IN1(n14645), .IN2(n14646), .Q(g25256) );
  INVX0 U14975 ( .INP(n14647), .ZN(n14646) );
  OR2X1 U14976 ( .IN1(n14640), .IN2(n8688), .Q(n14647) );
  AND2X1 U14977 ( .IN1(n14640), .IN2(n4377), .Q(n14645) );
  OR2X1 U14978 ( .IN1(n14648), .IN2(n14649), .Q(g25255) );
  AND2X1 U14979 ( .IN1(n14650), .IN2(n12145), .Q(n14649) );
  AND2X1 U14980 ( .IN1(n14651), .IN2(g1559), .Q(n14648) );
  OR2X1 U14981 ( .IN1(n14652), .IN2(n14653), .Q(g25253) );
  AND2X1 U14982 ( .IN1(n14654), .IN2(n12102), .Q(n14653) );
  OR2X1 U14983 ( .IN1(n14655), .IN2(n14656), .Q(n12102) );
  OR2X1 U14984 ( .IN1(n14657), .IN2(n14658), .Q(n14656) );
  OR2X1 U14985 ( .IN1(n4319), .IN2(n4287), .Q(n14658) );
  OR2X1 U14986 ( .IN1(n4373), .IN2(n4325), .Q(n14657) );
  OR2X1 U14987 ( .IN1(n14659), .IN2(n14660), .Q(n14655) );
  OR2X1 U14988 ( .IN1(n4389), .IN2(n4377), .Q(n14660) );
  OR2X1 U14989 ( .IN1(n4563), .IN2(n4555), .Q(n14659) );
  INVX0 U14990 ( .INP(n14661), .ZN(n14652) );
  OR2X1 U14991 ( .IN1(n14654), .IN2(n8687), .Q(n14661) );
  OR2X1 U14992 ( .IN1(n14662), .IN2(n14663), .Q(g25252) );
  INVX0 U14993 ( .INP(n14664), .ZN(n14663) );
  OR2X1 U14994 ( .IN1(n9117), .IN2(n8689), .Q(n14664) );
  AND2X1 U14995 ( .IN1(n9117), .IN2(n4377), .Q(n14662) );
  OR2X1 U14996 ( .IN1(n14665), .IN2(n14666), .Q(g25251) );
  INVX0 U14997 ( .INP(n14667), .ZN(n14666) );
  OR2X1 U14998 ( .IN1(n14640), .IN2(n8691), .Q(n14667) );
  AND2X1 U14999 ( .IN1(n14640), .IN2(n4373), .Q(n14665) );
  OR2X1 U15000 ( .IN1(n14668), .IN2(n14669), .Q(g25250) );
  AND2X1 U15001 ( .IN1(n14670), .IN2(n12145), .Q(n14669) );
  INVX0 U15002 ( .INP(n14671), .ZN(n14668) );
  OR2X1 U15003 ( .IN1(n14670), .IN2(n8698), .Q(n14671) );
  OR2X1 U15004 ( .IN1(n14672), .IN2(n14673), .Q(g25249) );
  INVX0 U15005 ( .INP(n14674), .ZN(n14673) );
  OR2X1 U15006 ( .IN1(n14650), .IN2(n8700), .Q(n14674) );
  AND2X1 U15007 ( .IN1(n14650), .IN2(n4378), .Q(n14672) );
  OR2X1 U15008 ( .IN1(n14675), .IN2(n14676), .Q(g25248) );
  AND2X1 U15009 ( .IN1(n14677), .IN2(n12185), .Q(n14676) );
  INVX0 U15010 ( .INP(n14678), .ZN(n14675) );
  OR2X1 U15011 ( .IN1(n14677), .IN2(n8708), .Q(n14678) );
  OR2X1 U15012 ( .IN1(n14679), .IN2(n14680), .Q(g25247) );
  INVX0 U15013 ( .INP(n14681), .ZN(n14680) );
  OR2X1 U15014 ( .IN1(n14654), .IN2(n8690), .Q(n14681) );
  AND2X1 U15015 ( .IN1(n14654), .IN2(n4377), .Q(n14679) );
  OR2X1 U15016 ( .IN1(n14682), .IN2(n14683), .Q(g25246) );
  INVX0 U15017 ( .INP(n14684), .ZN(n14683) );
  OR2X1 U15018 ( .IN1(n9117), .IN2(n8692), .Q(n14684) );
  AND2X1 U15019 ( .IN1(n9117), .IN2(n4373), .Q(n14682) );
  OR2X1 U15020 ( .IN1(n14685), .IN2(n14686), .Q(g25245) );
  AND2X1 U15021 ( .IN1(n14687), .IN2(n14640), .Q(n14686) );
  INVX0 U15022 ( .INP(n14688), .ZN(n14685) );
  OR2X1 U15023 ( .IN1(n14640), .IN2(n8694), .Q(n14688) );
  AND2X1 U15024 ( .IN1(g2241), .IN2(g13110), .Q(n14640) );
  OR2X1 U15025 ( .IN1(n14689), .IN2(n14690), .Q(g25244) );
  AND2X1 U15026 ( .IN1(n14691), .IN2(n12145), .Q(n14690) );
  OR2X1 U15027 ( .IN1(n14692), .IN2(n14693), .Q(n12145) );
  OR2X1 U15028 ( .IN1(n14694), .IN2(n14695), .Q(n14693) );
  OR2X1 U15029 ( .IN1(n4320), .IN2(n4288), .Q(n14695) );
  OR2X1 U15030 ( .IN1(n4374), .IN2(n4326), .Q(n14694) );
  OR2X1 U15031 ( .IN1(n14696), .IN2(n14697), .Q(n14692) );
  OR2X1 U15032 ( .IN1(n4390), .IN2(n4378), .Q(n14697) );
  OR2X1 U15033 ( .IN1(n4565), .IN2(n4557), .Q(n14696) );
  INVX0 U15034 ( .INP(n14698), .ZN(n14689) );
  OR2X1 U15035 ( .IN1(n14691), .IN2(n8699), .Q(n14698) );
  OR2X1 U15036 ( .IN1(n14699), .IN2(n14700), .Q(g25243) );
  INVX0 U15037 ( .INP(n14701), .ZN(n14700) );
  OR2X1 U15038 ( .IN1(n14670), .IN2(n8701), .Q(n14701) );
  AND2X1 U15039 ( .IN1(n14670), .IN2(n4378), .Q(n14699) );
  OR2X1 U15040 ( .IN1(n14702), .IN2(n14703), .Q(g25242) );
  AND2X1 U15041 ( .IN1(n14650), .IN2(n4374), .Q(n14703) );
  AND2X1 U15042 ( .IN1(test_so54), .IN2(n14651), .Q(n14702) );
  INVX0 U15043 ( .INP(n14650), .ZN(n14651) );
  OR2X1 U15044 ( .IN1(n14704), .IN2(n14705), .Q(g25241) );
  AND2X1 U15045 ( .IN1(n14706), .IN2(n12185), .Q(n14705) );
  AND2X1 U15046 ( .IN1(n14707), .IN2(g867), .Q(n14704) );
  OR2X1 U15047 ( .IN1(n14708), .IN2(n14709), .Q(g25240) );
  INVX0 U15048 ( .INP(n14710), .ZN(n14709) );
  OR2X1 U15049 ( .IN1(n14677), .IN2(n8711), .Q(n14710) );
  AND2X1 U15050 ( .IN1(n4379), .IN2(n14677), .Q(n14708) );
  OR2X1 U15051 ( .IN1(n14711), .IN2(n14712), .Q(g25239) );
  AND2X1 U15052 ( .IN1(n14713), .IN2(n12217), .Q(n14712) );
  INVX0 U15053 ( .INP(n14714), .ZN(n14711) );
  OR2X1 U15054 ( .IN1(n14713), .IN2(n8719), .Q(n14714) );
  OR2X1 U15055 ( .IN1(n14715), .IN2(n14716), .Q(g25237) );
  INVX0 U15056 ( .INP(n14717), .ZN(n14716) );
  OR2X1 U15057 ( .IN1(n14654), .IN2(n8693), .Q(n14717) );
  AND2X1 U15058 ( .IN1(n14654), .IN2(n4373), .Q(n14715) );
  OR2X1 U15059 ( .IN1(n14718), .IN2(n14719), .Q(g25236) );
  AND2X1 U15060 ( .IN1(n14687), .IN2(n9117), .Q(n14719) );
  INVX0 U15061 ( .INP(n14720), .ZN(n14718) );
  OR2X1 U15062 ( .IN1(n9117), .IN2(n8695), .Q(n14720) );
  AND2X1 U15063 ( .IN1(g13110), .IN2(test_so73), .Q(n9117) );
  OR2X1 U15064 ( .IN1(n14721), .IN2(n14722), .Q(g25235) );
  INVX0 U15065 ( .INP(n14723), .ZN(n14722) );
  OR2X1 U15066 ( .IN1(n14691), .IN2(n8702), .Q(n14723) );
  AND2X1 U15067 ( .IN1(n14691), .IN2(n4378), .Q(n14721) );
  OR2X1 U15068 ( .IN1(n14724), .IN2(n14725), .Q(g25234) );
  INVX0 U15069 ( .INP(n14726), .ZN(n14725) );
  OR2X1 U15070 ( .IN1(n14670), .IN2(n8703), .Q(n14726) );
  AND2X1 U15071 ( .IN1(n14670), .IN2(n4374), .Q(n14724) );
  OR2X1 U15072 ( .IN1(n14727), .IN2(n14728), .Q(g25233) );
  AND2X1 U15073 ( .IN1(n14729), .IN2(n14650), .Q(n14728) );
  INVX0 U15074 ( .INP(n14730), .ZN(n14727) );
  OR2X1 U15075 ( .IN1(n14650), .IN2(n8705), .Q(n14730) );
  AND2X1 U15076 ( .IN1(g1547), .IN2(g13110), .Q(n14650) );
  OR2X1 U15077 ( .IN1(n14731), .IN2(n14732), .Q(g25232) );
  AND2X1 U15078 ( .IN1(n14733), .IN2(n12185), .Q(n14732) );
  OR2X1 U15079 ( .IN1(n14734), .IN2(n14735), .Q(n12185) );
  OR2X1 U15080 ( .IN1(n14736), .IN2(n14737), .Q(n14735) );
  OR2X1 U15081 ( .IN1(n4321), .IN2(n4289), .Q(n14737) );
  OR2X1 U15082 ( .IN1(n4375), .IN2(n4327), .Q(n14736) );
  OR2X1 U15083 ( .IN1(n14738), .IN2(n14739), .Q(n14734) );
  OR2X1 U15084 ( .IN1(n4391), .IN2(n4379), .Q(n14739) );
  OR2X1 U15085 ( .IN1(n4567), .IN2(n4559), .Q(n14738) );
  INVX0 U15086 ( .INP(n14740), .ZN(n14731) );
  OR2X1 U15087 ( .IN1(n14733), .IN2(n8710), .Q(n14740) );
  OR2X1 U15088 ( .IN1(n14741), .IN2(n14742), .Q(g25231) );
  INVX0 U15089 ( .INP(n14743), .ZN(n14742) );
  OR2X1 U15090 ( .IN1(n14706), .IN2(n8712), .Q(n14743) );
  AND2X1 U15091 ( .IN1(n4379), .IN2(n14706), .Q(n14741) );
  OR2X1 U15092 ( .IN1(n14744), .IN2(n14745), .Q(g25230) );
  INVX0 U15093 ( .INP(n14746), .ZN(n14745) );
  OR2X1 U15094 ( .IN1(n14677), .IN2(n8714), .Q(n14746) );
  AND2X1 U15095 ( .IN1(n14677), .IN2(n4375), .Q(n14744) );
  OR2X1 U15096 ( .IN1(n14747), .IN2(n14748), .Q(g25229) );
  AND2X1 U15097 ( .IN1(n14749), .IN2(n12217), .Q(n14748) );
  INVX0 U15098 ( .INP(n14750), .ZN(n14747) );
  OR2X1 U15099 ( .IN1(n14749), .IN2(n8720), .Q(n14750) );
  OR2X1 U15100 ( .IN1(n14751), .IN2(n14752), .Q(g25228) );
  INVX0 U15101 ( .INP(n14753), .ZN(n14752) );
  OR2X1 U15102 ( .IN1(n14713), .IN2(n8722), .Q(n14753) );
  AND2X1 U15103 ( .IN1(n4380), .IN2(n14713), .Q(n14751) );
  OR2X1 U15104 ( .IN1(n14754), .IN2(n14755), .Q(g25227) );
  AND2X1 U15105 ( .IN1(n14687), .IN2(n14654), .Q(n14755) );
  INVX0 U15106 ( .INP(n14756), .ZN(n14687) );
  OR2X1 U15107 ( .IN1(n14757), .IN2(n14758), .Q(n14756) );
  OR2X1 U15108 ( .IN1(g2190), .IN2(g2195), .Q(n14758) );
  OR2X1 U15109 ( .IN1(n4325), .IN2(n4287), .Q(n14757) );
  INVX0 U15110 ( .INP(n14759), .ZN(n14754) );
  OR2X1 U15111 ( .IN1(n14654), .IN2(n8696), .Q(n14759) );
  AND2X1 U15112 ( .IN1(g6837), .IN2(g13110), .Q(n14654) );
  OR2X1 U15113 ( .IN1(n14760), .IN2(n14761), .Q(g25225) );
  INVX0 U15114 ( .INP(n14762), .ZN(n14761) );
  OR2X1 U15115 ( .IN1(n14691), .IN2(n8704), .Q(n14762) );
  AND2X1 U15116 ( .IN1(n14691), .IN2(n4374), .Q(n14760) );
  OR2X1 U15117 ( .IN1(n14763), .IN2(n14764), .Q(g25224) );
  AND2X1 U15118 ( .IN1(n14729), .IN2(n14670), .Q(n14764) );
  INVX0 U15119 ( .INP(n14765), .ZN(n14763) );
  OR2X1 U15120 ( .IN1(n14670), .IN2(n8706), .Q(n14765) );
  AND2X1 U15121 ( .IN1(g6782), .IN2(g13110), .Q(n14670) );
  OR2X1 U15122 ( .IN1(n14766), .IN2(n14767), .Q(g25223) );
  INVX0 U15123 ( .INP(n14768), .ZN(n14767) );
  OR2X1 U15124 ( .IN1(n14733), .IN2(n8713), .Q(n14768) );
  AND2X1 U15125 ( .IN1(n14733), .IN2(n4379), .Q(n14766) );
  OR2X1 U15126 ( .IN1(n14769), .IN2(n14770), .Q(g25222) );
  INVX0 U15127 ( .INP(n14771), .ZN(n14770) );
  OR2X1 U15128 ( .IN1(n14706), .IN2(n8715), .Q(n14771) );
  AND2X1 U15129 ( .IN1(n14706), .IN2(n4375), .Q(n14769) );
  OR2X1 U15130 ( .IN1(n14772), .IN2(n14773), .Q(g25221) );
  AND2X1 U15131 ( .IN1(n14774), .IN2(n14677), .Q(n14773) );
  INVX0 U15132 ( .INP(n14775), .ZN(n14772) );
  OR2X1 U15133 ( .IN1(n14677), .IN2(n8717), .Q(n14775) );
  AND2X1 U15134 ( .IN1(g13110), .IN2(test_so31), .Q(n14677) );
  OR2X1 U15135 ( .IN1(n14776), .IN2(n14777), .Q(g25220) );
  AND2X1 U15136 ( .IN1(n14778), .IN2(n12217), .Q(n14777) );
  OR2X1 U15137 ( .IN1(n14779), .IN2(n14780), .Q(n12217) );
  OR2X1 U15138 ( .IN1(n14781), .IN2(n14782), .Q(n14780) );
  OR2X1 U15139 ( .IN1(n4322), .IN2(n4290), .Q(n14782) );
  OR2X1 U15140 ( .IN1(n4376), .IN2(n4328), .Q(n14781) );
  OR2X1 U15141 ( .IN1(n14783), .IN2(n14784), .Q(n14779) );
  OR2X1 U15142 ( .IN1(n4392), .IN2(n4380), .Q(n14784) );
  OR2X1 U15143 ( .IN1(n4569), .IN2(n4561), .Q(n14783) );
  INVX0 U15144 ( .INP(n14785), .ZN(n14776) );
  OR2X1 U15145 ( .IN1(n14778), .IN2(n8721), .Q(n14785) );
  OR2X1 U15146 ( .IN1(n14786), .IN2(n14787), .Q(g25219) );
  INVX0 U15147 ( .INP(n14788), .ZN(n14787) );
  OR2X1 U15148 ( .IN1(n14749), .IN2(n8723), .Q(n14788) );
  AND2X1 U15149 ( .IN1(n4380), .IN2(n14749), .Q(n14786) );
  OR2X1 U15150 ( .IN1(n14789), .IN2(n14790), .Q(g25218) );
  INVX0 U15151 ( .INP(n14791), .ZN(n14790) );
  OR2X1 U15152 ( .IN1(n14713), .IN2(n8725), .Q(n14791) );
  AND2X1 U15153 ( .IN1(n14713), .IN2(n4376), .Q(n14789) );
  OR2X1 U15154 ( .IN1(n14792), .IN2(n14793), .Q(g25217) );
  AND2X1 U15155 ( .IN1(n14729), .IN2(n14691), .Q(n14793) );
  INVX0 U15156 ( .INP(n14794), .ZN(n14729) );
  OR2X1 U15157 ( .IN1(n14795), .IN2(n14796), .Q(n14794) );
  OR2X1 U15158 ( .IN1(g1496), .IN2(g1501), .Q(n14796) );
  OR2X1 U15159 ( .IN1(n4326), .IN2(n4288), .Q(n14795) );
  INVX0 U15160 ( .INP(n14797), .ZN(n14792) );
  OR2X1 U15161 ( .IN1(n14691), .IN2(n8707), .Q(n14797) );
  AND2X1 U15162 ( .IN1(g6573), .IN2(g13110), .Q(n14691) );
  OR2X1 U15163 ( .IN1(n14798), .IN2(n14799), .Q(g25215) );
  INVX0 U15164 ( .INP(n14800), .ZN(n14799) );
  OR2X1 U15165 ( .IN1(n14733), .IN2(n8716), .Q(n14800) );
  AND2X1 U15166 ( .IN1(n14733), .IN2(n4375), .Q(n14798) );
  OR2X1 U15167 ( .IN1(n14801), .IN2(n14802), .Q(g25214) );
  AND2X1 U15168 ( .IN1(n14774), .IN2(n14706), .Q(n14802) );
  AND2X1 U15169 ( .IN1(test_so33), .IN2(n14707), .Q(n14801) );
  INVX0 U15170 ( .INP(n14706), .ZN(n14707) );
  AND2X1 U15171 ( .IN1(g6518), .IN2(g13110), .Q(n14706) );
  OR2X1 U15172 ( .IN1(n14803), .IN2(n14804), .Q(g25213) );
  INVX0 U15173 ( .INP(n14805), .ZN(n14804) );
  OR2X1 U15174 ( .IN1(n14778), .IN2(n8724), .Q(n14805) );
  AND2X1 U15175 ( .IN1(n14778), .IN2(n4380), .Q(n14803) );
  OR2X1 U15176 ( .IN1(n14806), .IN2(n14807), .Q(g25212) );
  INVX0 U15177 ( .INP(n14808), .ZN(n14807) );
  OR2X1 U15178 ( .IN1(n14749), .IN2(n8726), .Q(n14808) );
  AND2X1 U15179 ( .IN1(n14749), .IN2(n4376), .Q(n14806) );
  OR2X1 U15180 ( .IN1(n14809), .IN2(n14810), .Q(g25211) );
  AND2X1 U15181 ( .IN1(n14811), .IN2(n14713), .Q(n14810) );
  INVX0 U15182 ( .INP(n14812), .ZN(n14809) );
  OR2X1 U15183 ( .IN1(n14713), .IN2(n8728), .Q(n14812) );
  AND2X1 U15184 ( .IN1(g165), .IN2(g13110), .Q(n14713) );
  OR2X1 U15185 ( .IN1(n14813), .IN2(n14814), .Q(g25209) );
  AND2X1 U15186 ( .IN1(n14774), .IN2(n14733), .Q(n14814) );
  INVX0 U15187 ( .INP(n14815), .ZN(n14774) );
  OR2X1 U15188 ( .IN1(n14816), .IN2(n14817), .Q(n14815) );
  OR2X1 U15189 ( .IN1(g805), .IN2(g809), .Q(n14817) );
  OR2X1 U15190 ( .IN1(n4327), .IN2(n4289), .Q(n14816) );
  INVX0 U15191 ( .INP(n14818), .ZN(n14813) );
  OR2X1 U15192 ( .IN1(n14733), .IN2(n8718), .Q(n14818) );
  AND2X1 U15193 ( .IN1(g6368), .IN2(g13110), .Q(n14733) );
  OR2X1 U15194 ( .IN1(n14819), .IN2(n14820), .Q(g25207) );
  INVX0 U15195 ( .INP(n14821), .ZN(n14820) );
  OR2X1 U15196 ( .IN1(n14778), .IN2(n8727), .Q(n14821) );
  AND2X1 U15197 ( .IN1(n14778), .IN2(n4376), .Q(n14819) );
  OR2X1 U15198 ( .IN1(n14822), .IN2(n14823), .Q(g25206) );
  AND2X1 U15199 ( .IN1(n14811), .IN2(n14749), .Q(n14823) );
  INVX0 U15200 ( .INP(n14824), .ZN(n14822) );
  OR2X1 U15201 ( .IN1(n14749), .IN2(n8729), .Q(n14824) );
  AND2X1 U15202 ( .IN1(g6313), .IN2(g13110), .Q(n14749) );
  OR2X1 U15203 ( .IN1(n14825), .IN2(n14826), .Q(g25204) );
  AND2X1 U15204 ( .IN1(n14811), .IN2(n14778), .Q(n14826) );
  INVX0 U15205 ( .INP(n14827), .ZN(n14811) );
  OR2X1 U15206 ( .IN1(n14828), .IN2(n14829), .Q(n14827) );
  OR2X1 U15207 ( .IN1(g117), .IN2(g121), .Q(n14829) );
  OR2X1 U15208 ( .IN1(n4328), .IN2(n4290), .Q(n14828) );
  INVX0 U15209 ( .INP(n14830), .ZN(n14825) );
  OR2X1 U15210 ( .IN1(n14778), .IN2(n8730), .Q(n14830) );
  AND2X1 U15211 ( .IN1(g6231), .IN2(g13110), .Q(n14778) );
  AND2X1 U15212 ( .IN1(n14831), .IN2(n9719), .Q(g25202) );
  XOR2X1 U15213 ( .IN1(n9086), .IN2(n14832), .Q(n14831) );
  AND2X1 U15214 ( .IN1(n14833), .IN2(n9662), .Q(g25201) );
  INVX0 U15215 ( .INP(n14834), .ZN(n14833) );
  OR2X1 U15216 ( .IN1(n14181), .IN2(n4057), .Q(n14834) );
  INVX0 U15217 ( .INP(n14180), .ZN(n14181) );
  OR2X1 U15218 ( .IN1(n4305), .IN2(n4058), .Q(n14180) );
  OR2X1 U15219 ( .IN1(n9102), .IN2(n14835), .Q(n4058) );
  AND2X1 U15220 ( .IN1(n14836), .IN2(n9507), .Q(g25199) );
  XOR2X1 U15221 ( .IN1(n14837), .IN2(n8822), .Q(n14836) );
  AND2X1 U15222 ( .IN1(n14838), .IN2(n12737), .Q(g25197) );
  XOR2X1 U15223 ( .IN1(n13732), .IN2(n4397), .Q(n14838) );
  AND2X1 U15224 ( .IN1(n14839), .IN2(n12741), .Q(g25194) );
  XOR2X1 U15225 ( .IN1(n13751), .IN2(n4399), .Q(n14839) );
  AND2X1 U15226 ( .IN1(n14840), .IN2(n13724), .Q(g25191) );
  AND2X1 U15227 ( .IN1(n14841), .IN2(n3742), .Q(n14840) );
  OR2X1 U15228 ( .IN1(n9092), .IN2(n14842), .Q(n3742) );
  INVX0 U15229 ( .INP(n14843), .ZN(n14841) );
  AND2X1 U15230 ( .IN1(n14842), .IN2(n9092), .Q(n14843) );
  INVX0 U15231 ( .INP(n4065), .ZN(n14842) );
  AND2X1 U15232 ( .IN1(n14844), .IN2(n12745), .Q(g25189) );
  XOR2X1 U15233 ( .IN1(n13843), .IN2(n4401), .Q(n14844) );
  AND2X1 U15234 ( .IN1(n14845), .IN2(n12226), .Q(g25185) );
  XOR2X1 U15235 ( .IN1(n13935), .IN2(n4403), .Q(n14845) );
  AND2X1 U15236 ( .IN1(n14846), .IN2(n11527), .Q(g25067) );
  OR2X1 U15237 ( .IN1(n14847), .IN2(n14848), .Q(n11527) );
  XOR2X1 U15238 ( .IN1(n3888), .IN2(n8809), .Q(n14846) );
  OR2X1 U15239 ( .IN1(n9552), .IN2(n4367), .Q(n3888) );
  AND2X1 U15240 ( .IN1(n14849), .IN2(n11529), .Q(g25056) );
  OR2X1 U15241 ( .IN1(n14847), .IN2(n14850), .Q(n11529) );
  XOR2X1 U15242 ( .IN1(n3891), .IN2(n8813), .Q(n14849) );
  OR2X1 U15243 ( .IN1(n9552), .IN2(n4368), .Q(n3891) );
  AND2X1 U15244 ( .IN1(n14851), .IN2(n11531), .Q(g25042) );
  OR2X1 U15245 ( .IN1(n14847), .IN2(n14852), .Q(n11531) );
  XOR2X1 U15246 ( .IN1(n8817), .IN2(n3894), .Q(n14851) );
  OR2X1 U15247 ( .IN1(n9552), .IN2(n9118), .Q(n3894) );
  AND2X1 U15248 ( .IN1(n14853), .IN2(n11533), .Q(g25027) );
  OR2X1 U15249 ( .IN1(n14847), .IN2(n14854), .Q(n11533) );
  XOR2X1 U15250 ( .IN1(n3897), .IN2(n8821), .Q(n14853) );
  OR2X1 U15251 ( .IN1(n9552), .IN2(n4369), .Q(n3897) );
  OR2X1 U15252 ( .IN1(n14855), .IN2(n12894), .Q(g24734) );
  INVX0 U15253 ( .INP(n3700), .ZN(n12894) );
  AND2X1 U15254 ( .IN1(n12898), .IN2(DFF_146_n1), .Q(n14855) );
  AND2X1 U15255 ( .IN1(n3705), .IN2(n3940), .Q(n12898) );
  OR2X1 U15256 ( .IN1(n14856), .IN2(n14857), .Q(g24557) );
  AND2X1 U15257 ( .IN1(n4299), .IN2(g2676), .Q(n14857) );
  AND2X1 U15258 ( .IN1(n14858), .IN2(n10225), .Q(n14856) );
  OR2X1 U15259 ( .IN1(n14859), .IN2(n14860), .Q(g24548) );
  AND2X1 U15260 ( .IN1(n14861), .IN2(g7390), .Q(n14860) );
  AND2X1 U15261 ( .IN1(n4370), .IN2(g2673), .Q(n14859) );
  OR2X1 U15262 ( .IN1(n14862), .IN2(n14863), .Q(g24547) );
  AND2X1 U15263 ( .IN1(n4299), .IN2(g2667), .Q(n14863) );
  AND2X1 U15264 ( .IN1(n14858), .IN2(n12332), .Q(n14862) );
  OR2X1 U15265 ( .IN1(n14864), .IN2(n14865), .Q(g24545) );
  AND2X1 U15266 ( .IN1(n4366), .IN2(g1982), .Q(n14865) );
  AND2X1 U15267 ( .IN1(n14866), .IN2(n12389), .Q(n14864) );
  OR2X1 U15268 ( .IN1(n14867), .IN2(n14868), .Q(g24538) );
  AND2X1 U15269 ( .IN1(n4314), .IN2(g2670), .Q(n14868) );
  AND2X1 U15270 ( .IN1(n14861), .IN2(g7302), .Q(n14867) );
  AND2X1 U15271 ( .IN1(n10225), .IN2(n12265), .Q(n14861) );
  OR2X1 U15272 ( .IN1(n14869), .IN2(n14870), .Q(n10225) );
  OR2X1 U15273 ( .IN1(n14871), .IN2(n14872), .Q(n14870) );
  AND2X1 U15274 ( .IN1(g7390), .IN2(g2673), .Q(n14872) );
  AND2X1 U15275 ( .IN1(n11411), .IN2(g2670), .Q(n14871) );
  OR2X1 U15276 ( .IN1(n14873), .IN2(n14874), .Q(n14869) );
  AND2X1 U15277 ( .IN1(g2624), .IN2(g2676), .Q(n14874) );
  AND2X1 U15278 ( .IN1(n14875), .IN2(test_so88), .Q(n14873) );
  AND2X1 U15279 ( .IN1(n10383), .IN2(g185), .Q(n14875) );
  OR2X1 U15280 ( .IN1(n14876), .IN2(n14877), .Q(n10383) );
  OR2X1 U15281 ( .IN1(n14878), .IN2(n14879), .Q(n14877) );
  AND2X1 U15282 ( .IN1(n11411), .IN2(g2639), .Q(n14879) );
  AND2X1 U15283 ( .IN1(g2624), .IN2(g2564), .Q(n14878) );
  AND2X1 U15284 ( .IN1(g7390), .IN2(g2641), .Q(n14876) );
  OR2X1 U15285 ( .IN1(n14880), .IN2(n14881), .Q(g24537) );
  AND2X1 U15286 ( .IN1(n14882), .IN2(g7390), .Q(n14881) );
  AND2X1 U15287 ( .IN1(n4370), .IN2(g2664), .Q(n14880) );
  OR2X1 U15288 ( .IN1(n14883), .IN2(n14884), .Q(g24535) );
  AND2X1 U15289 ( .IN1(n14885), .IN2(g7194), .Q(n14884) );
  AND2X1 U15290 ( .IN1(n4315), .IN2(g1979), .Q(n14883) );
  OR2X1 U15291 ( .IN1(n14886), .IN2(n14887), .Q(g24534) );
  AND2X1 U15292 ( .IN1(n4366), .IN2(g1973), .Q(n14887) );
  AND2X1 U15293 ( .IN1(n14866), .IN2(n12456), .Q(n14886) );
  OR2X1 U15294 ( .IN1(n14888), .IN2(n14889), .Q(g24532) );
  AND2X1 U15295 ( .IN1(n4300), .IN2(g1288), .Q(n14889) );
  AND2X1 U15296 ( .IN1(n14890), .IN2(n12512), .Q(n14888) );
  OR2X1 U15297 ( .IN1(n14891), .IN2(n14892), .Q(g24527) );
  AND2X1 U15298 ( .IN1(n14882), .IN2(n11411), .Q(n14892) );
  AND2X1 U15299 ( .IN1(n12332), .IN2(n12265), .Q(n14882) );
  OR2X1 U15300 ( .IN1(n14893), .IN2(n14894), .Q(n12332) );
  OR2X1 U15301 ( .IN1(n14895), .IN2(n14896), .Q(n14894) );
  AND2X1 U15302 ( .IN1(g7390), .IN2(g2664), .Q(n14896) );
  AND2X1 U15303 ( .IN1(g2624), .IN2(g2667), .Q(n14895) );
  OR2X1 U15304 ( .IN1(n14897), .IN2(n14898), .Q(n14893) );
  AND2X1 U15305 ( .IN1(g7302), .IN2(g2661), .Q(n14898) );
  AND2X1 U15306 ( .IN1(n14899), .IN2(n10382), .Q(n14897) );
  OR2X1 U15307 ( .IN1(n14900), .IN2(n14901), .Q(n10382) );
  OR2X1 U15308 ( .IN1(n14902), .IN2(n14903), .Q(n14901) );
  AND2X1 U15309 ( .IN1(g2624), .IN2(g2647), .Q(n14903) );
  AND2X1 U15310 ( .IN1(g7302), .IN2(g2643), .Q(n14902) );
  AND2X1 U15311 ( .IN1(g7390), .IN2(g2645), .Q(n14900) );
  AND2X1 U15312 ( .IN1(g185), .IN2(g2598), .Q(n14899) );
  AND2X1 U15313 ( .IN1(n4314), .IN2(g2661), .Q(n14891) );
  OR2X1 U15314 ( .IN1(n14904), .IN2(n14905), .Q(g24525) );
  AND2X1 U15315 ( .IN1(n4296), .IN2(g1976), .Q(n14905) );
  AND2X1 U15316 ( .IN1(n14885), .IN2(g7052), .Q(n14904) );
  AND2X1 U15317 ( .IN1(n12389), .IN2(n12265), .Q(n14885) );
  OR2X1 U15318 ( .IN1(n14906), .IN2(n14907), .Q(n12389) );
  OR2X1 U15319 ( .IN1(n14908), .IN2(n14909), .Q(n14907) );
  AND2X1 U15320 ( .IN1(g1930), .IN2(g1982), .Q(n14909) );
  AND2X1 U15321 ( .IN1(g7194), .IN2(g1979), .Q(n14908) );
  OR2X1 U15322 ( .IN1(n14910), .IN2(n14911), .Q(n14906) );
  AND2X1 U15323 ( .IN1(n12379), .IN2(g1976), .Q(n14911) );
  AND2X1 U15324 ( .IN1(n14912), .IN2(n10388), .Q(n14910) );
  OR2X1 U15325 ( .IN1(n14913), .IN2(n14914), .Q(n10388) );
  OR2X1 U15326 ( .IN1(n14915), .IN2(n14916), .Q(n14914) );
  AND2X1 U15327 ( .IN1(g7194), .IN2(g1947), .Q(n14916) );
  AND2X1 U15328 ( .IN1(n12379), .IN2(g1945), .Q(n14915) );
  AND2X1 U15329 ( .IN1(g1930), .IN2(g1870), .Q(n14913) );
  AND2X1 U15330 ( .IN1(g185), .IN2(g1922), .Q(n14912) );
  OR2X1 U15331 ( .IN1(n14917), .IN2(n14918), .Q(g24524) );
  AND2X1 U15332 ( .IN1(n14919), .IN2(g7194), .Q(n14918) );
  AND2X1 U15333 ( .IN1(n4315), .IN2(g1970), .Q(n14917) );
  OR2X1 U15334 ( .IN1(n14920), .IN2(n14921), .Q(g24522) );
  AND2X1 U15335 ( .IN1(n14922), .IN2(g6944), .Q(n14921) );
  AND2X1 U15336 ( .IN1(n4316), .IN2(g1285), .Q(n14920) );
  OR2X1 U15337 ( .IN1(n14923), .IN2(n14924), .Q(g24521) );
  AND2X1 U15338 ( .IN1(n4300), .IN2(g1279), .Q(n14924) );
  AND2X1 U15339 ( .IN1(n14890), .IN2(n12576), .Q(n14923) );
  OR2X1 U15340 ( .IN1(n14925), .IN2(n14926), .Q(g24519) );
  AND2X1 U15341 ( .IN1(n4313), .IN2(g602), .Q(n14926) );
  AND2X1 U15342 ( .IN1(n14927), .IN2(n12632), .Q(n14925) );
  OR2X1 U15343 ( .IN1(n14928), .IN2(n14929), .Q(g24513) );
  AND2X1 U15344 ( .IN1(n14919), .IN2(n12379), .Q(n14929) );
  AND2X1 U15345 ( .IN1(n12456), .IN2(n12265), .Q(n14919) );
  OR2X1 U15346 ( .IN1(n14930), .IN2(n14931), .Q(n12456) );
  OR2X1 U15347 ( .IN1(n14932), .IN2(n14933), .Q(n14931) );
  AND2X1 U15348 ( .IN1(g1930), .IN2(g1973), .Q(n14933) );
  AND2X1 U15349 ( .IN1(g7194), .IN2(g1970), .Q(n14932) );
  OR2X1 U15350 ( .IN1(n14934), .IN2(n14935), .Q(n14930) );
  AND2X1 U15351 ( .IN1(g7052), .IN2(g1967), .Q(n14935) );
  AND2X1 U15352 ( .IN1(n14936), .IN2(n10387), .Q(n14934) );
  OR2X1 U15353 ( .IN1(n14937), .IN2(n14938), .Q(n10387) );
  OR2X1 U15354 ( .IN1(n14939), .IN2(n14940), .Q(n14938) );
  AND2X1 U15355 ( .IN1(g7194), .IN2(g1951), .Q(n14940) );
  AND2X1 U15356 ( .IN1(g7052), .IN2(g1949), .Q(n14939) );
  AND2X1 U15357 ( .IN1(g1930), .IN2(g1953), .Q(n14937) );
  AND2X1 U15358 ( .IN1(g185), .IN2(g1904), .Q(n14936) );
  AND2X1 U15359 ( .IN1(n4296), .IN2(g1967), .Q(n14928) );
  OR2X1 U15360 ( .IN1(n14941), .IN2(n14942), .Q(g24511) );
  AND2X1 U15361 ( .IN1(n4371), .IN2(g1282), .Q(n14942) );
  AND2X1 U15362 ( .IN1(n14922), .IN2(g6750), .Q(n14941) );
  AND2X1 U15363 ( .IN1(n12512), .IN2(n12265), .Q(n14922) );
  OR2X1 U15364 ( .IN1(n14943), .IN2(n14944), .Q(n12512) );
  OR2X1 U15365 ( .IN1(n14945), .IN2(n14946), .Q(n14944) );
  AND2X1 U15366 ( .IN1(n12249), .IN2(g1282), .Q(n14946) );
  AND2X1 U15367 ( .IN1(g6944), .IN2(g1285), .Q(n14945) );
  OR2X1 U15368 ( .IN1(n14947), .IN2(n14948), .Q(n14943) );
  AND2X1 U15369 ( .IN1(g1236), .IN2(g1288), .Q(n14948) );
  AND2X1 U15370 ( .IN1(n14949), .IN2(test_so45), .Q(n14947) );
  AND2X1 U15371 ( .IN1(n9504), .IN2(g185), .Q(n14949) );
  OR2X1 U15372 ( .IN1(n14950), .IN2(n14951), .Q(n9504) );
  OR2X1 U15373 ( .IN1(n14952), .IN2(n14953), .Q(n14951) );
  AND2X1 U15374 ( .IN1(g1236), .IN2(g1176), .Q(n14953) );
  AND2X1 U15375 ( .IN1(g6750), .IN2(g1251), .Q(n14952) );
  AND2X1 U15376 ( .IN1(g6944), .IN2(g1253), .Q(n14950) );
  OR2X1 U15377 ( .IN1(n14954), .IN2(n14955), .Q(g24510) );
  AND2X1 U15378 ( .IN1(n14956), .IN2(g6944), .Q(n14955) );
  AND2X1 U15379 ( .IN1(n4316), .IN2(g1276), .Q(n14954) );
  OR2X1 U15380 ( .IN1(n14957), .IN2(n14958), .Q(g24508) );
  AND2X1 U15381 ( .IN1(n14959), .IN2(g6642), .Q(n14958) );
  AND2X1 U15382 ( .IN1(n4372), .IN2(g599), .Q(n14957) );
  OR2X1 U15383 ( .IN1(n14960), .IN2(n14961), .Q(g24507) );
  AND2X1 U15384 ( .IN1(n4313), .IN2(g593), .Q(n14961) );
  AND2X1 U15385 ( .IN1(n14927), .IN2(n12691), .Q(n14960) );
  OR2X1 U15386 ( .IN1(n14962), .IN2(n14963), .Q(g24501) );
  AND2X1 U15387 ( .IN1(n14956), .IN2(n12249), .Q(n14963) );
  AND2X1 U15388 ( .IN1(n12576), .IN2(n12265), .Q(n14956) );
  OR2X1 U15389 ( .IN1(n14964), .IN2(n14965), .Q(n12576) );
  OR2X1 U15390 ( .IN1(n14966), .IN2(n14967), .Q(n14965) );
  AND2X1 U15391 ( .IN1(g6944), .IN2(g1276), .Q(n14967) );
  AND2X1 U15392 ( .IN1(g1236), .IN2(g1279), .Q(n14966) );
  OR2X1 U15393 ( .IN1(n14968), .IN2(n14969), .Q(n14964) );
  AND2X1 U15394 ( .IN1(g6750), .IN2(g1273), .Q(n14969) );
  AND2X1 U15395 ( .IN1(n14970), .IN2(n9511), .Q(n14968) );
  OR2X1 U15396 ( .IN1(n14971), .IN2(n14972), .Q(n9511) );
  OR2X1 U15397 ( .IN1(n14973), .IN2(n14974), .Q(n14972) );
  AND2X1 U15398 ( .IN1(g6944), .IN2(g1257), .Q(n14974) );
  AND2X1 U15399 ( .IN1(g1236), .IN2(g1259), .Q(n14973) );
  AND2X1 U15400 ( .IN1(n12249), .IN2(g1255), .Q(n14971) );
  AND2X1 U15401 ( .IN1(g185), .IN2(g1210), .Q(n14970) );
  AND2X1 U15402 ( .IN1(n4371), .IN2(g1273), .Q(n14962) );
  OR2X1 U15403 ( .IN1(n14975), .IN2(n14976), .Q(g24499) );
  AND2X1 U15404 ( .IN1(n4298), .IN2(g596), .Q(n14976) );
  AND2X1 U15405 ( .IN1(n14959), .IN2(g6485), .Q(n14975) );
  AND2X1 U15406 ( .IN1(n12632), .IN2(n12265), .Q(n14959) );
  OR2X1 U15407 ( .IN1(n14977), .IN2(n14978), .Q(n12632) );
  OR2X1 U15408 ( .IN1(n14979), .IN2(n14980), .Q(n14978) );
  AND2X1 U15409 ( .IN1(g6642), .IN2(g599), .Q(n14980) );
  AND2X1 U15410 ( .IN1(g550), .IN2(g602), .Q(n14979) );
  OR2X1 U15411 ( .IN1(n14981), .IN2(n14982), .Q(n14977) );
  AND2X1 U15412 ( .IN1(g6485), .IN2(g596), .Q(n14982) );
  AND2X1 U15413 ( .IN1(n14983), .IN2(n9515), .Q(n14981) );
  OR2X1 U15414 ( .IN1(n14984), .IN2(n14985), .Q(n9515) );
  OR2X1 U15415 ( .IN1(n14986), .IN2(n14987), .Q(n14985) );
  AND2X1 U15416 ( .IN1(g550), .IN2(g489), .Q(n14987) );
  AND2X1 U15417 ( .IN1(n9810), .IN2(g565), .Q(n14986) );
  AND2X1 U15418 ( .IN1(g6642), .IN2(g567), .Q(n14984) );
  AND2X1 U15419 ( .IN1(g185), .IN2(g542), .Q(n14983) );
  OR2X1 U15420 ( .IN1(n14988), .IN2(n14989), .Q(g24498) );
  AND2X1 U15421 ( .IN1(n14990), .IN2(g6642), .Q(n14989) );
  AND2X1 U15422 ( .IN1(n4372), .IN2(g590), .Q(n14988) );
  OR2X1 U15423 ( .IN1(n14991), .IN2(n14992), .Q(g24491) );
  AND2X1 U15424 ( .IN1(n14990), .IN2(n9810), .Q(n14992) );
  AND2X1 U15425 ( .IN1(n12691), .IN2(n12265), .Q(n14990) );
  OR2X1 U15426 ( .IN1(n14993), .IN2(n14994), .Q(n12691) );
  OR2X1 U15427 ( .IN1(n14995), .IN2(n14996), .Q(n14994) );
  AND2X1 U15428 ( .IN1(g6642), .IN2(g590), .Q(n14996) );
  AND2X1 U15429 ( .IN1(g550), .IN2(g593), .Q(n14995) );
  OR2X1 U15430 ( .IN1(n14997), .IN2(n14998), .Q(n14993) );
  AND2X1 U15431 ( .IN1(n9810), .IN2(g587), .Q(n14998) );
  AND2X1 U15432 ( .IN1(n14999), .IN2(n9513), .Q(n14997) );
  OR2X1 U15433 ( .IN1(n15000), .IN2(n15001), .Q(n9513) );
  OR2X1 U15434 ( .IN1(n15002), .IN2(n15003), .Q(n15001) );
  AND2X1 U15435 ( .IN1(g550), .IN2(g573), .Q(n15003) );
  AND2X1 U15436 ( .IN1(g6485), .IN2(g569), .Q(n15002) );
  AND2X1 U15437 ( .IN1(g6642), .IN2(g571), .Q(n15000) );
  AND2X1 U15438 ( .IN1(g185), .IN2(g524), .Q(n14999) );
  AND2X1 U15439 ( .IN1(n4298), .IN2(g587), .Q(n14991) );
  AND2X1 U15440 ( .IN1(n15004), .IN2(n15005), .Q(g24476) );
  OR2X1 U15441 ( .IN1(n15006), .IN2(g2924), .Q(n15005) );
  AND2X1 U15442 ( .IN1(n9509), .IN2(g2917), .Q(n15006) );
  AND2X1 U15443 ( .IN1(n14837), .IN2(n9507), .Q(n15004) );
  OR2X1 U15444 ( .IN1(n15007), .IN2(n15008), .Q(n14837) );
  OR2X1 U15445 ( .IN1(n4479), .IN2(n4349), .Q(n15008) );
  AND2X1 U15446 ( .IN1(n15009), .IN2(n9662), .Q(g24473) );
  XOR2X1 U15447 ( .IN1(n14835), .IN2(n9102), .Q(n15009) );
  AND2X1 U15448 ( .IN1(n15010), .IN2(n14832), .Q(g24446) );
  OR2X1 U15449 ( .IN1(n4480), .IN2(n4102), .Q(n14832) );
  OR2X1 U15450 ( .IN1(n4350), .IN2(n15011), .Q(n4102) );
  AND2X1 U15451 ( .IN1(n9719), .IN2(n15012), .Q(n15010) );
  INVX0 U15452 ( .INP(n4101), .ZN(n15012) );
  AND2X1 U15453 ( .IN1(n15013), .IN2(n13724), .Q(g24445) );
  XOR2X1 U15454 ( .IN1(n4066), .IN2(n8282), .Q(n15013) );
  AND2X1 U15455 ( .IN1(n15014), .IN2(n15015), .Q(g24438) );
  INVX0 U15456 ( .INP(n15016), .ZN(n15015) );
  AND2X1 U15457 ( .IN1(n15017), .IN2(n4408), .Q(n15016) );
  OR2X1 U15458 ( .IN1(n15018), .IN2(n4419), .Q(n15017) );
  AND2X1 U15459 ( .IN1(n13732), .IN2(n12737), .Q(n15014) );
  OR2X1 U15460 ( .IN1(n15018), .IN2(n15019), .Q(n13732) );
  OR2X1 U15461 ( .IN1(n4419), .IN2(n4408), .Q(n15019) );
  AND2X1 U15462 ( .IN1(n15020), .IN2(n15021), .Q(g24434) );
  INVX0 U15463 ( .INP(n15022), .ZN(n15021) );
  AND2X1 U15464 ( .IN1(n15023), .IN2(n4410), .Q(n15022) );
  OR2X1 U15465 ( .IN1(n15024), .IN2(n4420), .Q(n15023) );
  AND2X1 U15466 ( .IN1(n13751), .IN2(n12741), .Q(n15020) );
  OR2X1 U15467 ( .IN1(n15024), .IN2(n15025), .Q(n13751) );
  OR2X1 U15468 ( .IN1(n4420), .IN2(n4410), .Q(n15025) );
  AND2X1 U15469 ( .IN1(n15026), .IN2(n15027), .Q(g24430) );
  INVX0 U15470 ( .INP(n15028), .ZN(n15027) );
  AND2X1 U15471 ( .IN1(n15029), .IN2(n4412), .Q(n15028) );
  OR2X1 U15472 ( .IN1(n15030), .IN2(n4421), .Q(n15029) );
  AND2X1 U15473 ( .IN1(n13843), .IN2(n12745), .Q(n15026) );
  OR2X1 U15474 ( .IN1(n15030), .IN2(n15031), .Q(n13843) );
  OR2X1 U15475 ( .IN1(n4421), .IN2(n4412), .Q(n15031) );
  AND2X1 U15476 ( .IN1(n15032), .IN2(n15033), .Q(g24426) );
  INVX0 U15477 ( .INP(n15034), .ZN(n15033) );
  AND2X1 U15478 ( .IN1(n15035), .IN2(n4414), .Q(n15034) );
  OR2X1 U15479 ( .IN1(n15036), .IN2(n4422), .Q(n15035) );
  AND2X1 U15480 ( .IN1(n13935), .IN2(n12226), .Q(n15032) );
  OR2X1 U15481 ( .IN1(n15036), .IN2(n15037), .Q(n13935) );
  OR2X1 U15482 ( .IN1(n4422), .IN2(n4414), .Q(n15037) );
  OR2X1 U15483 ( .IN1(n15038), .IN2(n15039), .Q(g24250) );
  AND2X1 U15484 ( .IN1(n15040), .IN2(g2560), .Q(n15039) );
  AND2X1 U15485 ( .IN1(n4463), .IN2(g2546), .Q(n15038) );
  OR2X1 U15486 ( .IN1(n15041), .IN2(n15042), .Q(g24243) );
  AND2X1 U15487 ( .IN1(n15043), .IN2(g1866), .Q(n15042) );
  AND2X1 U15488 ( .IN1(n4464), .IN2(g1852), .Q(n15041) );
  OR2X1 U15489 ( .IN1(n15044), .IN2(n15045), .Q(g24238) );
  AND2X1 U15490 ( .IN1(n11732), .IN2(g2560), .Q(n15045) );
  AND2X1 U15491 ( .IN1(n4463), .IN2(g2554), .Q(n15044) );
  OR2X1 U15492 ( .IN1(n15046), .IN2(n15047), .Q(g24237) );
  AND2X1 U15493 ( .IN1(n15040), .IN2(g8167), .Q(n15047) );
  AND2X1 U15494 ( .IN1(n4455), .IN2(g2543), .Q(n15046) );
  OR2X1 U15495 ( .IN1(n15048), .IN2(n15049), .Q(g24235) );
  AND2X1 U15496 ( .IN1(n15050), .IN2(g1172), .Q(n15049) );
  AND2X1 U15497 ( .IN1(n4465), .IN2(g1158), .Q(n15048) );
  OR2X1 U15498 ( .IN1(n15051), .IN2(n15052), .Q(g24231) );
  AND2X1 U15499 ( .IN1(n11842), .IN2(g1866), .Q(n15052) );
  AND2X1 U15500 ( .IN1(n4464), .IN2(g1860), .Q(n15051) );
  OR2X1 U15501 ( .IN1(n15053), .IN2(n15054), .Q(g24230) );
  AND2X1 U15502 ( .IN1(n15043), .IN2(g8082), .Q(n15054) );
  AND2X1 U15503 ( .IN1(n4457), .IN2(g1849), .Q(n15053) );
  OR2X1 U15504 ( .IN1(n15055), .IN2(n15056), .Q(g24228) );
  AND2X1 U15505 ( .IN1(n15057), .IN2(g485), .Q(n15056) );
  AND2X1 U15506 ( .IN1(n4466), .IN2(g471), .Q(n15055) );
  OR2X1 U15507 ( .IN1(n15058), .IN2(n15059), .Q(g24226) );
  AND2X1 U15508 ( .IN1(n11732), .IN2(g8167), .Q(n15059) );
  AND2X1 U15509 ( .IN1(n4455), .IN2(g2553), .Q(n15058) );
  OR2X1 U15510 ( .IN1(n15060), .IN2(n15061), .Q(g24225) );
  AND2X1 U15511 ( .IN1(n15040), .IN2(g8087), .Q(n15061) );
  INVX0 U15512 ( .INP(n9659), .ZN(n15040) );
  OR2X1 U15513 ( .IN1(n10854), .IN2(n10872), .Q(n9659) );
  OR2X1 U15514 ( .IN1(n10850), .IN2(n10860), .Q(n10872) );
  AND2X1 U15515 ( .IN1(n4456), .IN2(g2540), .Q(n15060) );
  OR2X1 U15516 ( .IN1(n15062), .IN2(n15063), .Q(g24223) );
  AND2X1 U15517 ( .IN1(n11945), .IN2(g1172), .Q(n15063) );
  AND2X1 U15518 ( .IN1(n4465), .IN2(g1166), .Q(n15062) );
  OR2X1 U15519 ( .IN1(n15064), .IN2(n15065), .Q(g24222) );
  AND2X1 U15520 ( .IN1(n15050), .IN2(g8007), .Q(n15065) );
  AND2X1 U15521 ( .IN1(n4459), .IN2(g1155), .Q(n15064) );
  OR2X1 U15522 ( .IN1(n15066), .IN2(n15067), .Q(g24219) );
  AND2X1 U15523 ( .IN1(n11842), .IN2(g8082), .Q(n15067) );
  AND2X1 U15524 ( .IN1(n4457), .IN2(g1859), .Q(n15066) );
  OR2X1 U15525 ( .IN1(n15068), .IN2(n15069), .Q(g24218) );
  AND2X1 U15526 ( .IN1(n15043), .IN2(g8012), .Q(n15069) );
  INVX0 U15527 ( .INP(n9625), .ZN(n15043) );
  OR2X1 U15528 ( .IN1(n10440), .IN2(n10458), .Q(n9625) );
  OR2X1 U15529 ( .IN1(n10436), .IN2(n10446), .Q(n10458) );
  AND2X1 U15530 ( .IN1(n4458), .IN2(g1846), .Q(n15068) );
  OR2X1 U15531 ( .IN1(n15070), .IN2(n15071), .Q(g24216) );
  AND2X1 U15532 ( .IN1(n12040), .IN2(g485), .Q(n15071) );
  AND2X1 U15533 ( .IN1(n4466), .IN2(g479), .Q(n15070) );
  OR2X1 U15534 ( .IN1(n15072), .IN2(n15073), .Q(g24215) );
  AND2X1 U15535 ( .IN1(test_so24), .IN2(n4461), .Q(n15073) );
  AND2X1 U15536 ( .IN1(n15057), .IN2(g7956), .Q(n15072) );
  OR2X1 U15537 ( .IN1(n15074), .IN2(n15075), .Q(g24214) );
  AND2X1 U15538 ( .IN1(n11732), .IN2(g8087), .Q(n15075) );
  INVX0 U15539 ( .INP(n11189), .ZN(n11732) );
  OR2X1 U15540 ( .IN1(n10860), .IN2(n15076), .Q(n11189) );
  OR2X1 U15541 ( .IN1(n10871), .IN2(n10847), .Q(n15076) );
  INVX0 U15542 ( .INP(n10850), .ZN(n10847) );
  AND2X1 U15543 ( .IN1(n4456), .IN2(g2552), .Q(n15074) );
  OR2X1 U15544 ( .IN1(n15077), .IN2(n15078), .Q(g24213) );
  AND2X1 U15545 ( .IN1(n11945), .IN2(g8007), .Q(n15078) );
  AND2X1 U15546 ( .IN1(n4459), .IN2(g1165), .Q(n15077) );
  OR2X1 U15547 ( .IN1(n15079), .IN2(n15080), .Q(g24212) );
  AND2X1 U15548 ( .IN1(n15050), .IN2(g7961), .Q(n15080) );
  INVX0 U15549 ( .INP(n9590), .ZN(n15050) );
  OR2X1 U15550 ( .IN1(n10232), .IN2(n10281), .Q(n9590) );
  OR2X1 U15551 ( .IN1(n10239), .IN2(n10243), .Q(n10281) );
  AND2X1 U15552 ( .IN1(n4460), .IN2(g1152), .Q(n15079) );
  OR2X1 U15553 ( .IN1(n15081), .IN2(n15082), .Q(g24209) );
  AND2X1 U15554 ( .IN1(n9657), .IN2(g2560), .Q(n15082) );
  AND2X1 U15555 ( .IN1(n4463), .IN2(g2536), .Q(n15081) );
  OR2X1 U15556 ( .IN1(n15083), .IN2(n15084), .Q(g24208) );
  AND2X1 U15557 ( .IN1(n11842), .IN2(g8012), .Q(n15084) );
  INVX0 U15558 ( .INP(n11249), .ZN(n11842) );
  OR2X1 U15559 ( .IN1(n10446), .IN2(n15085), .Q(n11249) );
  OR2X1 U15560 ( .IN1(n10457), .IN2(n10433), .Q(n15085) );
  INVX0 U15561 ( .INP(n10436), .ZN(n10433) );
  AND2X1 U15562 ( .IN1(n4458), .IN2(g1858), .Q(n15083) );
  OR2X1 U15563 ( .IN1(n15086), .IN2(n15087), .Q(g24207) );
  AND2X1 U15564 ( .IN1(n12040), .IN2(g7956), .Q(n15087) );
  AND2X1 U15565 ( .IN1(n4461), .IN2(g478), .Q(n15086) );
  OR2X1 U15566 ( .IN1(n15088), .IN2(n15089), .Q(g24206) );
  AND2X1 U15567 ( .IN1(test_so23), .IN2(n15057), .Q(n15089) );
  INVX0 U15568 ( .INP(n9556), .ZN(n15057) );
  OR2X1 U15569 ( .IN1(n10496), .IN2(n10514), .Q(n9556) );
  OR2X1 U15570 ( .IN1(n10492), .IN2(n10502), .Q(n10514) );
  AND2X1 U15571 ( .IN1(g465), .IN2(n9120), .Q(n15088) );
  OR2X1 U15572 ( .IN1(n15090), .IN2(n15091), .Q(g24182) );
  AND2X1 U15573 ( .IN1(n9622), .IN2(g1866), .Q(n15091) );
  AND2X1 U15574 ( .IN1(n4464), .IN2(g1842), .Q(n15090) );
  OR2X1 U15575 ( .IN1(n15092), .IN2(n15093), .Q(g24181) );
  AND2X1 U15576 ( .IN1(n11945), .IN2(g7961), .Q(n15093) );
  INVX0 U15577 ( .INP(n11309), .ZN(n11945) );
  OR2X1 U15578 ( .IN1(n10243), .IN2(n15094), .Q(n11309) );
  OR2X1 U15579 ( .IN1(n10236), .IN2(n10230), .Q(n15094) );
  INVX0 U15580 ( .INP(n10239), .ZN(n10230) );
  AND2X1 U15581 ( .IN1(n4460), .IN2(g1164), .Q(n15092) );
  OR2X1 U15582 ( .IN1(n15095), .IN2(n15096), .Q(g24179) );
  AND2X1 U15583 ( .IN1(n9588), .IN2(g1172), .Q(n15096) );
  AND2X1 U15584 ( .IN1(n4465), .IN2(g1148), .Q(n15095) );
  OR2X1 U15585 ( .IN1(n15097), .IN2(n15098), .Q(g24178) );
  AND2X1 U15586 ( .IN1(test_so23), .IN2(n12040), .Q(n15098) );
  INVX0 U15587 ( .INP(n11363), .ZN(n12040) );
  OR2X1 U15588 ( .IN1(n10502), .IN2(n15099), .Q(n11363) );
  OR2X1 U15589 ( .IN1(n10513), .IN2(n10489), .Q(n15099) );
  INVX0 U15590 ( .INP(n10492), .ZN(n10489) );
  AND2X1 U15591 ( .IN1(g477), .IN2(n9120), .Q(n15097) );
  OR2X1 U15592 ( .IN1(n15100), .IN2(n15101), .Q(g24174) );
  AND2X1 U15593 ( .IN1(n9553), .IN2(g485), .Q(n15101) );
  AND2X1 U15594 ( .IN1(n4466), .IN2(g461), .Q(n15100) );
  OR2X1 U15595 ( .IN1(n15102), .IN2(n15103), .Q(g24092) );
  AND2X1 U15596 ( .IN1(n10061), .IN2(g2380), .Q(n15103) );
  AND2X1 U15597 ( .IN1(g3229), .IN2(n4483), .Q(n15102) );
  OR2X1 U15598 ( .IN1(n15104), .IN2(n15105), .Q(g24083) );
  AND2X1 U15599 ( .IN1(n10061), .IN2(g1686), .Q(n15105) );
  INVX0 U15600 ( .INP(g3229), .ZN(n10061) );
  AND2X1 U15601 ( .IN1(g3229), .IN2(n4484), .Q(n15104) );
  OR2X1 U15602 ( .IN1(n15106), .IN2(n15107), .Q(g24072) );
  INVX0 U15603 ( .INP(n15108), .ZN(n15107) );
  OR2X1 U15604 ( .IN1(g3229), .IN2(n8824), .Q(n15108) );
  AND2X1 U15605 ( .IN1(g3229), .IN2(n4486), .Q(n15106) );
  OR2X1 U15606 ( .IN1(n15109), .IN2(n15110), .Q(g24059) );
  INVX0 U15607 ( .INP(n15111), .ZN(n15110) );
  OR2X1 U15608 ( .IN1(g3229), .IN2(n8546), .Q(n15111) );
  AND2X1 U15609 ( .IN1(g3229), .IN2(n4485), .Q(n15109) );
  OR2X1 U15610 ( .IN1(n15112), .IN2(n15113), .Q(g23418) );
  AND2X1 U15611 ( .IN1(n9657), .IN2(g8167), .Q(n15113) );
  AND2X1 U15612 ( .IN1(n4455), .IN2(g2533), .Q(n15112) );
  OR2X1 U15613 ( .IN1(n15114), .IN2(n15115), .Q(g23413) );
  AND2X1 U15614 ( .IN1(test_so65), .IN2(n4457), .Q(n15115) );
  AND2X1 U15615 ( .IN1(n9622), .IN2(g8082), .Q(n15114) );
  OR2X1 U15616 ( .IN1(n15116), .IN2(n15117), .Q(g23407) );
  AND2X1 U15617 ( .IN1(n9657), .IN2(g8087), .Q(n15117) );
  AND2X1 U15618 ( .IN1(n10871), .IN2(n15118), .Q(n9657) );
  AND2X1 U15619 ( .IN1(n10860), .IN2(n10850), .Q(n15118) );
  OR2X1 U15620 ( .IN1(n15119), .IN2(n15120), .Q(n10850) );
  OR2X1 U15621 ( .IN1(n15121), .IN2(n15122), .Q(n15120) );
  AND2X1 U15622 ( .IN1(n8384), .IN2(n10408), .Q(n15122) );
  AND2X1 U15623 ( .IN1(n8383), .IN2(n10833), .Q(n15121) );
  AND2X1 U15624 ( .IN1(n8374), .IN2(n10398), .Q(n15119) );
  OR2X1 U15625 ( .IN1(n15123), .IN2(n15124), .Q(n10860) );
  OR2X1 U15626 ( .IN1(n15125), .IN2(n15126), .Q(n15124) );
  AND2X1 U15627 ( .IN1(n8386), .IN2(n10408), .Q(n15126) );
  AND2X1 U15628 ( .IN1(n8385), .IN2(n10833), .Q(n15125) );
  AND2X1 U15629 ( .IN1(n8375), .IN2(n10398), .Q(n15123) );
  INVX0 U15630 ( .INP(n10854), .ZN(n10871) );
  OR2X1 U15631 ( .IN1(n15127), .IN2(n15128), .Q(n10854) );
  OR2X1 U15632 ( .IN1(n15129), .IN2(n15130), .Q(n15128) );
  AND2X1 U15633 ( .IN1(n8388), .IN2(n10408), .Q(n15130) );
  INVX0 U15634 ( .INP(n4516), .ZN(n10408) );
  AND2X1 U15635 ( .IN1(n8387), .IN2(n10833), .Q(n15129) );
  INVX0 U15636 ( .INP(n4509), .ZN(n10833) );
  AND2X1 U15637 ( .IN1(n8376), .IN2(n10398), .Q(n15127) );
  INVX0 U15638 ( .INP(n4524), .ZN(n10398) );
  AND2X1 U15639 ( .IN1(n4456), .IN2(g2530), .Q(n15116) );
  OR2X1 U15640 ( .IN1(n15131), .IN2(n15132), .Q(g23406) );
  AND2X1 U15641 ( .IN1(n9588), .IN2(g8007), .Q(n15132) );
  AND2X1 U15642 ( .IN1(n4459), .IN2(g1145), .Q(n15131) );
  OR2X1 U15643 ( .IN1(n15133), .IN2(n15134), .Q(g23400) );
  AND2X1 U15644 ( .IN1(n9622), .IN2(g8012), .Q(n15134) );
  AND2X1 U15645 ( .IN1(n10457), .IN2(n15135), .Q(n9622) );
  AND2X1 U15646 ( .IN1(n10446), .IN2(n10436), .Q(n15135) );
  OR2X1 U15647 ( .IN1(n15136), .IN2(n15137), .Q(n10436) );
  OR2X1 U15648 ( .IN1(n15138), .IN2(n15139), .Q(n15137) );
  AND2X1 U15649 ( .IN1(n8390), .IN2(n10419), .Q(n15139) );
  AND2X1 U15650 ( .IN1(n8389), .IN2(n10403), .Q(n15138) );
  AND2X1 U15651 ( .IN1(n8377), .IN2(n10412), .Q(n15136) );
  OR2X1 U15652 ( .IN1(n15140), .IN2(n15141), .Q(n10446) );
  OR2X1 U15653 ( .IN1(n15142), .IN2(n15143), .Q(n15141) );
  AND2X1 U15654 ( .IN1(n8392), .IN2(n10419), .Q(n15143) );
  AND2X1 U15655 ( .IN1(n8391), .IN2(n10403), .Q(n15142) );
  AND2X1 U15656 ( .IN1(n8378), .IN2(n10412), .Q(n15140) );
  INVX0 U15657 ( .INP(n10440), .ZN(n10457) );
  OR2X1 U15658 ( .IN1(n15144), .IN2(n15145), .Q(n10440) );
  OR2X1 U15659 ( .IN1(n15146), .IN2(n15147), .Q(n15145) );
  AND2X1 U15660 ( .IN1(n8394), .IN2(n10419), .Q(n15147) );
  INVX0 U15661 ( .INP(n4518), .ZN(n10419) );
  AND2X1 U15662 ( .IN1(n8393), .IN2(n10403), .Q(n15146) );
  INVX0 U15663 ( .INP(n4511), .ZN(n10403) );
  AND2X1 U15664 ( .IN1(n8379), .IN2(n10412), .Q(n15144) );
  INVX0 U15665 ( .INP(n4525), .ZN(n10412) );
  AND2X1 U15666 ( .IN1(n4458), .IN2(g1836), .Q(n15133) );
  OR2X1 U15667 ( .IN1(n15148), .IN2(n15149), .Q(g23399) );
  AND2X1 U15668 ( .IN1(n9553), .IN2(g7956), .Q(n15149) );
  AND2X1 U15669 ( .IN1(n4461), .IN2(g458), .Q(n15148) );
  OR2X1 U15670 ( .IN1(n15150), .IN2(n15151), .Q(g23392) );
  AND2X1 U15671 ( .IN1(n9588), .IN2(g7961), .Q(n15151) );
  AND2X1 U15672 ( .IN1(n10236), .IN2(n15152), .Q(n9588) );
  AND2X1 U15673 ( .IN1(n10243), .IN2(n10239), .Q(n15152) );
  OR2X1 U15674 ( .IN1(n15153), .IN2(n15154), .Q(n10239) );
  OR2X1 U15675 ( .IN1(n15155), .IN2(n15156), .Q(n15154) );
  AND2X1 U15676 ( .IN1(n8380), .IN2(g6712), .Q(n15156) );
  AND2X1 U15677 ( .IN1(n8395), .IN2(g5472), .Q(n15155) );
  INVX0 U15678 ( .INP(n15157), .ZN(n15153) );
  OR2X1 U15679 ( .IN1(n4381), .IN2(test_so39), .Q(n15157) );
  OR2X1 U15680 ( .IN1(n15158), .IN2(n15159), .Q(n10243) );
  OR2X1 U15681 ( .IN1(n15160), .IN2(n15161), .Q(n15159) );
  AND2X1 U15682 ( .IN1(n8381), .IN2(g6712), .Q(n15161) );
  AND2X1 U15683 ( .IN1(n8397), .IN2(g5472), .Q(n15160) );
  AND2X1 U15684 ( .IN1(n8396), .IN2(g1088), .Q(n15158) );
  INVX0 U15685 ( .INP(n10232), .ZN(n10236) );
  OR2X1 U15686 ( .IN1(n15162), .IN2(n15163), .Q(n10232) );
  OR2X1 U15687 ( .IN1(n15164), .IN2(n15165), .Q(n15163) );
  AND2X1 U15688 ( .IN1(n8382), .IN2(g6712), .Q(n15165) );
  AND2X1 U15689 ( .IN1(n8399), .IN2(g5472), .Q(n15164) );
  AND2X1 U15690 ( .IN1(n8398), .IN2(g1088), .Q(n15162) );
  AND2X1 U15691 ( .IN1(n4460), .IN2(g1142), .Q(n15150) );
  OR2X1 U15692 ( .IN1(n15166), .IN2(n15167), .Q(g23385) );
  AND2X1 U15693 ( .IN1(n9553), .IN2(test_so23), .Q(n15167) );
  AND2X1 U15694 ( .IN1(n10513), .IN2(n15168), .Q(n9553) );
  AND2X1 U15695 ( .IN1(n10502), .IN2(n10492), .Q(n15168) );
  OR2X1 U15696 ( .IN1(n15169), .IN2(n15170), .Q(n10492) );
  OR2X1 U15697 ( .IN1(n15171), .IN2(n15172), .Q(n15170) );
  AND2X1 U15698 ( .IN1(n8400), .IN2(n10465), .Q(n15172) );
  AND2X1 U15699 ( .IN1(n8401), .IN2(n10899), .Q(n15171) );
  AND2X1 U15700 ( .IN1(n8402), .IN2(n10475), .Q(n15169) );
  OR2X1 U15701 ( .IN1(n15173), .IN2(n15174), .Q(n10502) );
  OR2X1 U15702 ( .IN1(n15175), .IN2(n15176), .Q(n15174) );
  AND2X1 U15703 ( .IN1(n8403), .IN2(n10465), .Q(n15176) );
  INVX0 U15704 ( .INP(n15177), .ZN(n15175) );
  OR2X1 U15705 ( .IN1(n4499), .IN2(test_so18), .Q(n15177) );
  AND2X1 U15706 ( .IN1(n8404), .IN2(n10475), .Q(n15173) );
  INVX0 U15707 ( .INP(n10496), .ZN(n10513) );
  OR2X1 U15708 ( .IN1(n15178), .IN2(n15179), .Q(n10496) );
  OR2X1 U15709 ( .IN1(n15180), .IN2(n15181), .Q(n15179) );
  AND2X1 U15710 ( .IN1(n8405), .IN2(n10465), .Q(n15181) );
  INVX0 U15711 ( .INP(n4506), .ZN(n10465) );
  AND2X1 U15712 ( .IN1(n8406), .IN2(n10899), .Q(n15180) );
  INVX0 U15713 ( .INP(n4499), .ZN(n10899) );
  AND2X1 U15714 ( .IN1(n8407), .IN2(n10475), .Q(n15178) );
  INVX0 U15715 ( .INP(n4520), .ZN(n10475) );
  AND2X1 U15716 ( .IN1(g455), .IN2(n9120), .Q(n15166) );
  AND2X1 U15717 ( .IN1(n15182), .IN2(n9719), .Q(g23359) );
  OR2X1 U15718 ( .IN1(n15183), .IN2(n13724), .Q(n9719) );
  AND2X1 U15719 ( .IN1(n15184), .IN2(n15185), .Q(n15183) );
  OR2X1 U15720 ( .IN1(n15186), .IN2(n15187), .Q(n15184) );
  INVX0 U15721 ( .INP(n15188), .ZN(n15187) );
  AND2X1 U15722 ( .IN1(n4350), .IN2(n4480), .Q(n15188) );
  OR2X1 U15723 ( .IN1(n9086), .IN2(n4481), .Q(n15186) );
  XNOR2X1 U15724 ( .IN1(n4350), .IN2(n9721), .Q(n15182) );
  INVX0 U15725 ( .INP(n15011), .ZN(n9721) );
  OR2X1 U15726 ( .IN1(n4481), .IN2(n9722), .Q(n15011) );
  AND2X1 U15727 ( .IN1(n15189), .IN2(n9662), .Q(g23358) );
  AND2X1 U15728 ( .IN1(n14835), .IN2(n15190), .Q(n15189) );
  INVX0 U15729 ( .INP(n4122_Tj_Payload), .ZN(n15190) );
  OR2X1 U15730 ( .IN1(n4431), .IN2(n4123), .Q(n14835) );
  OR2X1 U15731 ( .IN1(n9081), .IN2(n9664), .Q(n4123) );
  AND2X1 U15732 ( .IN1(n15191), .IN2(n9507), .Q(g23357) );
  OR2X1 U15733 ( .IN1(n15192), .IN2(n9662), .Q(n9507) );
  AND2X1 U15734 ( .IN1(n16489), .IN2(n15193), .Q(n15192) );
  OR2X1 U15735 ( .IN1(n15194), .IN2(n15195), .Q(n15193) );
  OR2X1 U15736 ( .IN1(g2917), .IN2(g2924), .Q(n15195) );
  OR2X1 U15737 ( .IN1(n8822), .IN2(n4482), .Q(n15194) );
  XNOR2X1 U15738 ( .IN1(n9509), .IN2(n4479), .Q(n15191) );
  INVX0 U15739 ( .INP(n15007), .ZN(n9509) );
  OR2X1 U15740 ( .IN1(n4482), .IN2(n9510), .Q(n15007) );
  AND2X1 U15741 ( .IN1(n15196), .IN2(n12737), .Q(g23348) );
  XOR2X1 U15742 ( .IN1(n15018), .IN2(n4419), .Q(n15196) );
  AND2X1 U15743 ( .IN1(n15197), .IN2(n12741), .Q(g23339) );
  XOR2X1 U15744 ( .IN1(n15024), .IN2(n4420), .Q(n15197) );
  AND2X1 U15745 ( .IN1(n15198), .IN2(n13724), .Q(g23330) );
  AND2X1 U15746 ( .IN1(n9722), .IN2(n15185), .Q(n13724) );
  OR2X1 U15747 ( .IN1(n9094), .IN2(n15199), .Q(n9722) );
  AND2X1 U15748 ( .IN1(n15200), .IN2(n4066), .Q(n15198) );
  OR2X1 U15749 ( .IN1(n14177), .IN2(n15201), .Q(n4066) );
  OR2X1 U15750 ( .IN1(n16493), .IN2(n9093), .Q(n15201) );
  INVX0 U15751 ( .INP(n15202), .ZN(n15200) );
  AND2X1 U15752 ( .IN1(n15203), .IN2(n9093), .Q(n15202) );
  OR2X1 U15753 ( .IN1(n14177), .IN2(n16493), .Q(n15203) );
  OR2X1 U15754 ( .IN1(n9094), .IN2(n9095), .Q(n14177) );
  AND2X1 U15755 ( .IN1(n15204), .IN2(n12745), .Q(g23329) );
  XOR2X1 U15756 ( .IN1(n15030), .IN2(n4421), .Q(n15204) );
  AND2X1 U15757 ( .IN1(n15205), .IN2(n12226), .Q(g23324) );
  XOR2X1 U15758 ( .IN1(n15036), .IN2(n4422), .Q(n15205) );
  OR2X1 U15759 ( .IN1(n15206), .IN2(n15207), .Q(g23137) );
  AND2X1 U15760 ( .IN1(n12805), .IN2(g1866), .Q(n15207) );
  AND2X1 U15761 ( .IN1(n4464), .IN2(g1869), .Q(n15206) );
  AND2X1 U15762 ( .IN1(n15208), .IN2(n15209), .Q(g23136) );
  INVX0 U15763 ( .INP(n15210), .ZN(n15209) );
  AND2X1 U15764 ( .IN1(n15211), .IN2(n4478), .Q(n15210) );
  OR2X1 U15765 ( .IN1(n15212), .IN2(n4404), .Q(n15211) );
  AND2X1 U15766 ( .IN1(n15036), .IN2(n12226), .Q(n15208) );
  OR2X1 U15767 ( .IN1(n15212), .IN2(n15213), .Q(n15036) );
  OR2X1 U15768 ( .IN1(n4478), .IN2(n4404), .Q(n15213) );
  OR2X1 U15769 ( .IN1(n15214), .IN2(n15215), .Q(g23133) );
  AND2X1 U15770 ( .IN1(n12782), .IN2(g8167), .Q(n15215) );
  AND2X1 U15771 ( .IN1(n4455), .IN2(g2562), .Q(n15214) );
  OR2X1 U15772 ( .IN1(n15216), .IN2(n15217), .Q(g23132) );
  AND2X1 U15773 ( .IN1(n11552), .IN2(g8087), .Q(n15217) );
  AND2X1 U15774 ( .IN1(n4456), .IN2(g2555), .Q(n15216) );
  OR2X1 U15775 ( .IN1(n15218), .IN2(n15219), .Q(g23126) );
  AND2X1 U15776 ( .IN1(n12832), .IN2(g1172), .Q(n15219) );
  AND2X1 U15777 ( .IN1(n4465), .IN2(g1175), .Q(n15218) );
  OR2X1 U15778 ( .IN1(n15220), .IN2(n15221), .Q(g23124) );
  AND2X1 U15779 ( .IN1(n12805), .IN2(g8082), .Q(n15221) );
  AND2X1 U15780 ( .IN1(n4457), .IN2(g1868), .Q(n15220) );
  OR2X1 U15781 ( .IN1(n15222), .IN2(n15223), .Q(g23123) );
  AND2X1 U15782 ( .IN1(n11584), .IN2(g8012), .Q(n15223) );
  AND2X1 U15783 ( .IN1(n4458), .IN2(g1861), .Q(n15222) );
  OR2X1 U15784 ( .IN1(n15224), .IN2(n15225), .Q(g23117) );
  AND2X1 U15785 ( .IN1(n12859), .IN2(g485), .Q(n15225) );
  AND2X1 U15786 ( .IN1(n4466), .IN2(g488), .Q(n15224) );
  OR2X1 U15787 ( .IN1(n15226), .IN2(n15227), .Q(g23114) );
  AND2X1 U15788 ( .IN1(n12782), .IN2(g8087), .Q(n15227) );
  AND2X1 U15789 ( .IN1(n4456), .IN2(g2561), .Q(n15226) );
  OR2X1 U15790 ( .IN1(n15228), .IN2(n15229), .Q(g23111) );
  AND2X1 U15791 ( .IN1(n12832), .IN2(g8007), .Q(n15229) );
  AND2X1 U15792 ( .IN1(test_so44), .IN2(n4459), .Q(n15228) );
  OR2X1 U15793 ( .IN1(n15230), .IN2(n15231), .Q(g23110) );
  AND2X1 U15794 ( .IN1(n11593), .IN2(g7961), .Q(n15231) );
  AND2X1 U15795 ( .IN1(n4460), .IN2(g1167), .Q(n15230) );
  OR2X1 U15796 ( .IN1(n15232), .IN2(n15233), .Q(g23097) );
  AND2X1 U15797 ( .IN1(n12805), .IN2(g8012), .Q(n15233) );
  OR2X1 U15798 ( .IN1(n15234), .IN2(n15235), .Q(n12805) );
  OR2X1 U15799 ( .IN1(n15236), .IN2(n15237), .Q(n15235) );
  AND2X1 U15800 ( .IN1(g7014), .IN2(g1822), .Q(n15237) );
  AND2X1 U15801 ( .IN1(test_so59), .IN2(n4618), .Q(n15236) );
  AND2X1 U15802 ( .IN1(g5511), .IN2(g1819), .Q(n15234) );
  AND2X1 U15803 ( .IN1(n4458), .IN2(g1867), .Q(n15232) );
  OR2X1 U15804 ( .IN1(n15238), .IN2(n15239), .Q(g23093) );
  AND2X1 U15805 ( .IN1(n12859), .IN2(g7956), .Q(n15239) );
  AND2X1 U15806 ( .IN1(n4461), .IN2(g487), .Q(n15238) );
  OR2X1 U15807 ( .IN1(n15240), .IN2(n15241), .Q(g23092) );
  AND2X1 U15808 ( .IN1(test_so23), .IN2(n11622), .Q(n15241) );
  AND2X1 U15809 ( .IN1(g480), .IN2(n9120), .Q(n15240) );
  OR2X1 U15810 ( .IN1(n15242), .IN2(n15243), .Q(g23081) );
  AND2X1 U15811 ( .IN1(n12832), .IN2(g7961), .Q(n15243) );
  OR2X1 U15812 ( .IN1(n15244), .IN2(n15245), .Q(n12832) );
  OR2X1 U15813 ( .IN1(n15246), .IN2(n15247), .Q(n15245) );
  AND2X1 U15814 ( .IN1(g6712), .IN2(g1128), .Q(n15247) );
  AND2X1 U15815 ( .IN1(g5472), .IN2(g1125), .Q(n15246) );
  AND2X1 U15816 ( .IN1(g1088), .IN2(g1131), .Q(n15244) );
  AND2X1 U15817 ( .IN1(n4460), .IN2(g1173), .Q(n15242) );
  OR2X1 U15818 ( .IN1(n15248), .IN2(n15249), .Q(g23076) );
  AND2X1 U15819 ( .IN1(n11552), .IN2(g2560), .Q(n15249) );
  AND2X1 U15820 ( .IN1(n4463), .IN2(g2539), .Q(n15248) );
  OR2X1 U15821 ( .IN1(n15250), .IN2(n15251), .Q(g23067) );
  AND2X1 U15822 ( .IN1(test_so23), .IN2(n12859), .Q(n15251) );
  OR2X1 U15823 ( .IN1(n15252), .IN2(n15253), .Q(n12859) );
  OR2X1 U15824 ( .IN1(n15254), .IN2(n15255), .Q(n15253) );
  AND2X1 U15825 ( .IN1(g6447), .IN2(g441), .Q(n15255) );
  AND2X1 U15826 ( .IN1(n4640), .IN2(g444), .Q(n15254) );
  AND2X1 U15827 ( .IN1(g5437), .IN2(g438), .Q(n15252) );
  AND2X1 U15828 ( .IN1(g486), .IN2(n9120), .Q(n15250) );
  OR2X1 U15829 ( .IN1(n15256), .IN2(n15257), .Q(g23058) );
  AND2X1 U15830 ( .IN1(n11584), .IN2(g1866), .Q(n15257) );
  AND2X1 U15831 ( .IN1(n4464), .IN2(g1845), .Q(n15256) );
  OR2X1 U15832 ( .IN1(n15258), .IN2(n15259), .Q(g23047) );
  AND2X1 U15833 ( .IN1(n11552), .IN2(g8167), .Q(n15259) );
  INVX0 U15834 ( .INP(n4285), .ZN(n11552) );
  OR2X1 U15835 ( .IN1(n15260), .IN2(n15261), .Q(n4285) );
  OR2X1 U15836 ( .IN1(n15262), .IN2(n15263), .Q(n15261) );
  AND2X1 U15837 ( .IN1(g7264), .IN2(g2495), .Q(n15263) );
  AND2X1 U15838 ( .IN1(n4606), .IN2(g2498), .Q(n15262) );
  AND2X1 U15839 ( .IN1(g5555), .IN2(g2492), .Q(n15260) );
  AND2X1 U15840 ( .IN1(n4455), .IN2(g2559), .Q(n15258) );
  OR2X1 U15841 ( .IN1(n15264), .IN2(n15265), .Q(g23039) );
  AND2X1 U15842 ( .IN1(n11593), .IN2(g1172), .Q(n15265) );
  AND2X1 U15843 ( .IN1(n4465), .IN2(g1151), .Q(n15264) );
  OR2X1 U15844 ( .IN1(n15266), .IN2(n15267), .Q(g23030) );
  AND2X1 U15845 ( .IN1(n11584), .IN2(g8082), .Q(n15267) );
  INVX0 U15846 ( .INP(n4284), .ZN(n11584) );
  OR2X1 U15847 ( .IN1(n15268), .IN2(n15269), .Q(n4284) );
  OR2X1 U15848 ( .IN1(n15270), .IN2(n15271), .Q(n15269) );
  AND2X1 U15849 ( .IN1(g7014), .IN2(g1801), .Q(n15271) );
  AND2X1 U15850 ( .IN1(n4618), .IN2(g1804), .Q(n15270) );
  AND2X1 U15851 ( .IN1(g5511), .IN2(g1798), .Q(n15268) );
  AND2X1 U15852 ( .IN1(n4457), .IN2(g1865), .Q(n15266) );
  OR2X1 U15853 ( .IN1(n15272), .IN2(n15273), .Q(g23022) );
  AND2X1 U15854 ( .IN1(n11622), .IN2(g485), .Q(n15273) );
  AND2X1 U15855 ( .IN1(n4466), .IN2(g464), .Q(n15272) );
  OR2X1 U15856 ( .IN1(n15274), .IN2(n15275), .Q(g23014) );
  AND2X1 U15857 ( .IN1(n11593), .IN2(g8007), .Q(n15275) );
  INVX0 U15858 ( .INP(n4283), .ZN(n11593) );
  OR2X1 U15859 ( .IN1(n15276), .IN2(n15277), .Q(n4283) );
  OR2X1 U15860 ( .IN1(n15278), .IN2(n15279), .Q(n15277) );
  AND2X1 U15861 ( .IN1(g6712), .IN2(g1107), .Q(n15279) );
  AND2X1 U15862 ( .IN1(g5472), .IN2(g1104), .Q(n15278) );
  AND2X1 U15863 ( .IN1(g1088), .IN2(g1110), .Q(n15276) );
  AND2X1 U15864 ( .IN1(n4459), .IN2(g1171), .Q(n15274) );
  OR2X1 U15865 ( .IN1(n15280), .IN2(n15281), .Q(g23000) );
  AND2X1 U15866 ( .IN1(n11622), .IN2(g7956), .Q(n15281) );
  INVX0 U15867 ( .INP(n4282), .ZN(n11622) );
  OR2X1 U15868 ( .IN1(n15282), .IN2(n15283), .Q(n4282) );
  OR2X1 U15869 ( .IN1(n15284), .IN2(n15285), .Q(n15283) );
  AND2X1 U15870 ( .IN1(g6447), .IN2(g420), .Q(n15285) );
  AND2X1 U15871 ( .IN1(n4640), .IN2(g423), .Q(n15284) );
  AND2X1 U15872 ( .IN1(g5437), .IN2(g417), .Q(n15282) );
  AND2X1 U15873 ( .IN1(n4461), .IN2(g484), .Q(n15280) );
  OR2X1 U15874 ( .IN1(n15286), .IN2(n15287), .Q(g22687) );
  AND2X1 U15875 ( .IN1(n15288), .IN2(n15289), .Q(n15287) );
  OR2X1 U15876 ( .IN1(n14028), .IN2(n9937), .Q(n15288) );
  AND2X1 U15877 ( .IN1(n15290), .IN2(n14028), .Q(n15286) );
  INVX0 U15878 ( .INP(n15291), .ZN(n14028) );
  OR2X1 U15879 ( .IN1(n15292), .IN2(n15293), .Q(n15291) );
  OR2X1 U15880 ( .IN1(n15294), .IN2(n15295), .Q(n15293) );
  AND2X1 U15881 ( .IN1(n11411), .IN2(g2565), .Q(n15295) );
  AND2X1 U15882 ( .IN1(g2624), .IN2(g2571), .Q(n15294) );
  AND2X1 U15883 ( .IN1(g7390), .IN2(g2568), .Q(n15292) );
  AND2X1 U15884 ( .IN1(n9889), .IN2(g2584), .Q(n15290) );
  OR2X1 U15885 ( .IN1(n15296), .IN2(n15297), .Q(g22651) );
  AND2X1 U15886 ( .IN1(n15298), .IN2(n15289), .Q(n15297) );
  OR2X1 U15887 ( .IN1(n14037), .IN2(n10071), .Q(n15298) );
  AND2X1 U15888 ( .IN1(n15299), .IN2(n14037), .Q(n15296) );
  INVX0 U15889 ( .INP(n15300), .ZN(n14037) );
  OR2X1 U15890 ( .IN1(n15301), .IN2(n15302), .Q(n15300) );
  OR2X1 U15891 ( .IN1(n15303), .IN2(n15304), .Q(n15302) );
  AND2X1 U15892 ( .IN1(g7194), .IN2(g1874), .Q(n15304) );
  AND2X1 U15893 ( .IN1(test_so68), .IN2(n12379), .Q(n15303) );
  AND2X1 U15894 ( .IN1(g1930), .IN2(g1877), .Q(n15301) );
  AND2X1 U15895 ( .IN1(n10023), .IN2(g1890), .Q(n15299) );
  OR2X1 U15896 ( .IN1(n15305), .IN2(n15306), .Q(g22615) );
  AND2X1 U15897 ( .IN1(n15307), .IN2(n15289), .Q(n15306) );
  OR2X1 U15898 ( .IN1(n14046), .IN2(n10206), .Q(n15307) );
  AND2X1 U15899 ( .IN1(n15308), .IN2(n14046), .Q(n15305) );
  INVX0 U15900 ( .INP(n15309), .ZN(n14046) );
  OR2X1 U15901 ( .IN1(n15310), .IN2(n15311), .Q(n15309) );
  OR2X1 U15902 ( .IN1(n15312), .IN2(n15313), .Q(n15311) );
  AND2X1 U15903 ( .IN1(g6944), .IN2(g1180), .Q(n15313) );
  AND2X1 U15904 ( .IN1(g1236), .IN2(g1183), .Q(n15312) );
  AND2X1 U15905 ( .IN1(test_so47), .IN2(n12249), .Q(n15310) );
  AND2X1 U15906 ( .IN1(n10158), .IN2(g1196), .Q(n15308) );
  OR2X1 U15907 ( .IN1(n15314), .IN2(n15315), .Q(g22578) );
  AND2X1 U15908 ( .IN1(n15316), .IN2(n15289), .Q(n15315) );
  INVX0 U15909 ( .INP(n15317), .ZN(n15289) );
  OR2X1 U15910 ( .IN1(n14052), .IN2(n9805), .Q(n15316) );
  AND2X1 U15911 ( .IN1(n15318), .IN2(n14052), .Q(n15314) );
  INVX0 U15912 ( .INP(n15319), .ZN(n14052) );
  OR2X1 U15913 ( .IN1(n15320), .IN2(n15321), .Q(n15319) );
  OR2X1 U15914 ( .IN1(n15322), .IN2(n15323), .Q(n15321) );
  AND2X1 U15915 ( .IN1(g550), .IN2(g496), .Q(n15323) );
  AND2X1 U15916 ( .IN1(g6485), .IN2(g490), .Q(n15322) );
  AND2X1 U15917 ( .IN1(g6642), .IN2(g493), .Q(n15320) );
  AND2X1 U15918 ( .IN1(test_so22), .IN2(n9738), .Q(n15318) );
  AND2X1 U15919 ( .IN1(n15324), .IN2(n15325), .Q(g22299) );
  OR2X1 U15920 ( .IN1(n14299), .IN2(test_so95), .Q(n15324) );
  AND2X1 U15921 ( .IN1(n15326), .IN2(n12737), .Q(g22284) );
  OR2X1 U15922 ( .IN1(n14304), .IN2(g2813), .Q(n15326) );
  AND2X1 U15923 ( .IN1(n15327), .IN2(n15328), .Q(g22280) );
  OR2X1 U15924 ( .IN1(n4149_Tj_Payload), .IN2(g2117), .Q(n15327) );
  AND2X1 U15925 ( .IN1(n15329), .IN2(n15330), .Q(g22269) );
  OR2X1 U15926 ( .IN1(n14312), .IN2(g2812), .Q(n15329) );
  AND2X1 U15927 ( .IN1(n15331), .IN2(n12741), .Q(g22267) );
  OR2X1 U15928 ( .IN1(n14387), .IN2(g2119), .Q(n15331) );
  AND2X1 U15929 ( .IN1(n15332), .IN2(n15333), .Q(g22263) );
  OR2X1 U15930 ( .IN1(n14392), .IN2(g1423), .Q(n15332) );
  AND2X1 U15931 ( .IN1(n15334), .IN2(n15335), .Q(g22249) );
  OR2X1 U15932 ( .IN1(n14396), .IN2(g2118), .Q(n15334) );
  AND2X1 U15933 ( .IN1(n15336), .IN2(n12745), .Q(g22247) );
  OR2X1 U15934 ( .IN1(n4160_Tj_Payload), .IN2(g1425), .Q(n15336) );
  AND2X1 U15935 ( .IN1(n15337), .IN2(n15338), .Q(g22242) );
  OR2X1 U15936 ( .IN1(n4161_Tj_Payload), .IN2(g737), .Q(n15337) );
  AND2X1 U15937 ( .IN1(n15339), .IN2(n15340), .Q(g22234) );
  OR2X1 U15938 ( .IN1(n14484), .IN2(g1424), .Q(n15339) );
  AND2X1 U15939 ( .IN1(n15341), .IN2(n12226), .Q(g22231) );
  OR2X1 U15940 ( .IN1(n14561), .IN2(g739), .Q(n15341) );
  AND2X1 U15941 ( .IN1(n15342), .IN2(n15343), .Q(g22218) );
  OR2X1 U15942 ( .IN1(n14565), .IN2(g738), .Q(n15342) );
  OR2X1 U15943 ( .IN1(n15344), .IN2(n15345), .Q(g22200) );
  INVX0 U15944 ( .INP(n15346), .ZN(n15345) );
  OR2X1 U15945 ( .IN1(n15347), .IN2(n8633), .Q(n15346) );
  AND2X1 U15946 ( .IN1(n15347), .IN2(n4373), .Q(n15344) );
  OR2X1 U15947 ( .IN1(n15348), .IN2(n15349), .Q(g22194) );
  AND2X1 U15948 ( .IN1(n14848), .IN2(g2238), .Q(n15349) );
  AND2X1 U15949 ( .IN1(n15347), .IN2(n10555), .Q(n15348) );
  OR2X1 U15950 ( .IN1(n15350), .IN2(n15351), .Q(g22193) );
  INVX0 U15951 ( .INP(n15352), .ZN(n15351) );
  OR2X1 U15952 ( .IN1(n15353), .IN2(n8994), .Q(n15352) );
  AND2X1 U15953 ( .IN1(n15353), .IN2(n4373), .Q(n15350) );
  OR2X1 U15954 ( .IN1(n15354), .IN2(n15355), .Q(g22192) );
  INVX0 U15955 ( .INP(n15356), .ZN(n15355) );
  OR2X1 U15956 ( .IN1(n15347), .IN2(n8634), .Q(n15356) );
  AND2X1 U15957 ( .IN1(n15347), .IN2(n4377), .Q(n15354) );
  OR2X1 U15958 ( .IN1(n15357), .IN2(n15358), .Q(g22191) );
  AND2X1 U15959 ( .IN1(n14850), .IN2(g1514), .Q(n15358) );
  AND2X1 U15960 ( .IN1(n15359), .IN2(n4374), .Q(n15357) );
  OR2X1 U15961 ( .IN1(n15360), .IN2(n15361), .Q(g22185) );
  AND2X1 U15962 ( .IN1(n15353), .IN2(n10555), .Q(n15361) );
  AND2X1 U15963 ( .IN1(test_so75), .IN2(n15362), .Q(n15360) );
  OR2X1 U15964 ( .IN1(n15363), .IN2(n15364), .Q(g22184) );
  AND2X1 U15965 ( .IN1(n14848), .IN2(g2235), .Q(n15364) );
  AND2X1 U15966 ( .IN1(n11693), .IN2(n15347), .Q(n15363) );
  OR2X1 U15967 ( .IN1(n15365), .IN2(n15366), .Q(g22183) );
  INVX0 U15968 ( .INP(n15367), .ZN(n15366) );
  OR2X1 U15969 ( .IN1(n15368), .IN2(n8995), .Q(n15367) );
  AND2X1 U15970 ( .IN1(n15368), .IN2(n4373), .Q(n15365) );
  OR2X1 U15971 ( .IN1(n15369), .IN2(n15370), .Q(g22182) );
  INVX0 U15972 ( .INP(n15371), .ZN(n15370) );
  OR2X1 U15973 ( .IN1(n15353), .IN2(n8996), .Q(n15371) );
  AND2X1 U15974 ( .IN1(n15353), .IN2(n4377), .Q(n15369) );
  OR2X1 U15975 ( .IN1(n15372), .IN2(n15373), .Q(g22180) );
  AND2X1 U15976 ( .IN1(n14850), .IN2(g1544), .Q(n15373) );
  AND2X1 U15977 ( .IN1(n15359), .IN2(n10589), .Q(n15372) );
  OR2X1 U15978 ( .IN1(n15374), .IN2(n15375), .Q(g22179) );
  AND2X1 U15979 ( .IN1(n15376), .IN2(g1516), .Q(n15375) );
  AND2X1 U15980 ( .IN1(n15377), .IN2(n4374), .Q(n15374) );
  OR2X1 U15981 ( .IN1(n15378), .IN2(n15379), .Q(g22178) );
  AND2X1 U15982 ( .IN1(n14850), .IN2(g1511), .Q(n15379) );
  AND2X1 U15983 ( .IN1(n15359), .IN2(n4378), .Q(n15378) );
  OR2X1 U15984 ( .IN1(n15380), .IN2(n15381), .Q(g22177) );
  INVX0 U15985 ( .INP(n15382), .ZN(n15381) );
  OR2X1 U15986 ( .IN1(n15383), .IN2(n8658), .Q(n15382) );
  AND2X1 U15987 ( .IN1(n15383), .IN2(n4375), .Q(n15380) );
  OR2X1 U15988 ( .IN1(n15384), .IN2(n15385), .Q(g22173) );
  AND2X1 U15989 ( .IN1(n15386), .IN2(g2239), .Q(n15385) );
  AND2X1 U15990 ( .IN1(n15368), .IN2(n10555), .Q(n15384) );
  INVX0 U15991 ( .INP(n14217), .ZN(n10555) );
  OR2X1 U15992 ( .IN1(n15387), .IN2(n15388), .Q(n14217) );
  OR2X1 U15993 ( .IN1(n15389), .IN2(n15390), .Q(n15388) );
  AND2X1 U15994 ( .IN1(n8691), .IN2(g2241), .Q(n15390) );
  AND2X1 U15995 ( .IN1(n8693), .IN2(g6837), .Q(n15389) );
  AND2X1 U15996 ( .IN1(n8692), .IN2(test_so73), .Q(n15387) );
  OR2X1 U15997 ( .IN1(n15391), .IN2(n15392), .Q(g22172) );
  AND2X1 U15998 ( .IN1(n15362), .IN2(g2237), .Q(n15392) );
  AND2X1 U15999 ( .IN1(n11693), .IN2(n15353), .Q(n15391) );
  OR2X1 U16000 ( .IN1(n15393), .IN2(n15394), .Q(g22171) );
  INVX0 U16001 ( .INP(n15395), .ZN(n15394) );
  OR2X1 U16002 ( .IN1(n15347), .IN2(n8627), .Q(n15395) );
  AND2X1 U16003 ( .IN1(n15347), .IN2(n4287), .Q(n15393) );
  OR2X1 U16004 ( .IN1(n15396), .IN2(n15397), .Q(g22170) );
  INVX0 U16005 ( .INP(n15398), .ZN(n15397) );
  OR2X1 U16006 ( .IN1(n15368), .IN2(n8997), .Q(n15398) );
  AND2X1 U16007 ( .IN1(n15368), .IN2(n4377), .Q(n15396) );
  OR2X1 U16008 ( .IN1(n15399), .IN2(n15400), .Q(g22169) );
  AND2X1 U16009 ( .IN1(n15376), .IN2(g1546), .Q(n15400) );
  AND2X1 U16010 ( .IN1(n15377), .IN2(n10589), .Q(n15399) );
  OR2X1 U16011 ( .IN1(n15401), .IN2(n15402), .Q(g22168) );
  AND2X1 U16012 ( .IN1(n14850), .IN2(g1541), .Q(n15402) );
  AND2X1 U16013 ( .IN1(n11800), .IN2(n15359), .Q(n15401) );
  OR2X1 U16014 ( .IN1(n15403), .IN2(n15404), .Q(g22167) );
  AND2X1 U16015 ( .IN1(n15405), .IN2(n4374), .Q(n15404) );
  AND2X1 U16016 ( .IN1(test_so52), .IN2(n15406), .Q(n15403) );
  OR2X1 U16017 ( .IN1(n15407), .IN2(n15408), .Q(g22166) );
  AND2X1 U16018 ( .IN1(n15376), .IN2(g1513), .Q(n15408) );
  AND2X1 U16019 ( .IN1(n15377), .IN2(n4378), .Q(n15407) );
  OR2X1 U16020 ( .IN1(n15409), .IN2(n15410), .Q(g22164) );
  AND2X1 U16021 ( .IN1(n14852), .IN2(g850), .Q(n15410) );
  AND2X1 U16022 ( .IN1(n15383), .IN2(n10629), .Q(n15409) );
  OR2X1 U16023 ( .IN1(n15411), .IN2(n15412), .Q(g22163) );
  INVX0 U16024 ( .INP(n15413), .ZN(n15412) );
  OR2X1 U16025 ( .IN1(n15414), .IN2(n9023), .Q(n15413) );
  AND2X1 U16026 ( .IN1(n15414), .IN2(n4375), .Q(n15411) );
  OR2X1 U16027 ( .IN1(n15415), .IN2(n15416), .Q(g22162) );
  INVX0 U16028 ( .INP(n15417), .ZN(n15416) );
  OR2X1 U16029 ( .IN1(n15383), .IN2(n8659), .Q(n15417) );
  AND2X1 U16030 ( .IN1(n4379), .IN2(n15383), .Q(n15415) );
  OR2X1 U16031 ( .IN1(n15418), .IN2(n15419), .Q(g22161) );
  AND2X1 U16032 ( .IN1(n14854), .IN2(g132), .Q(n15419) );
  AND2X1 U16033 ( .IN1(n15420), .IN2(n4376), .Q(n15418) );
  OR2X1 U16034 ( .IN1(n15421), .IN2(n15422), .Q(g22155) );
  AND2X1 U16035 ( .IN1(n15386), .IN2(g2236), .Q(n15422) );
  AND2X1 U16036 ( .IN1(n15368), .IN2(n11693), .Q(n15421) );
  INVX0 U16037 ( .INP(n10714), .ZN(n11693) );
  OR2X1 U16038 ( .IN1(n15423), .IN2(n15424), .Q(n10714) );
  OR2X1 U16039 ( .IN1(n15425), .IN2(n15426), .Q(n15424) );
  AND2X1 U16040 ( .IN1(n8688), .IN2(g2241), .Q(n15426) );
  AND2X1 U16041 ( .IN1(n8690), .IN2(g6837), .Q(n15425) );
  AND2X1 U16042 ( .IN1(n8689), .IN2(test_so73), .Q(n15423) );
  OR2X1 U16043 ( .IN1(n15427), .IN2(n15428), .Q(g22154) );
  INVX0 U16044 ( .INP(n15429), .ZN(n15428) );
  OR2X1 U16045 ( .IN1(n15353), .IN2(n8983), .Q(n15429) );
  AND2X1 U16046 ( .IN1(n15353), .IN2(n4287), .Q(n15427) );
  OR2X1 U16047 ( .IN1(n15430), .IN2(n15431), .Q(g22153) );
  AND2X1 U16048 ( .IN1(n14848), .IN2(g2229), .Q(n15431) );
  AND2X1 U16049 ( .IN1(n15347), .IN2(n4563), .Q(n15430) );
  OR2X1 U16050 ( .IN1(n15432), .IN2(n15433), .Q(g22152) );
  AND2X1 U16051 ( .IN1(n15406), .IN2(g1545), .Q(n15433) );
  AND2X1 U16052 ( .IN1(n15405), .IN2(n10589), .Q(n15432) );
  INVX0 U16053 ( .INP(n11819), .ZN(n10589) );
  OR2X1 U16054 ( .IN1(n15434), .IN2(n15435), .Q(n11819) );
  OR2X1 U16055 ( .IN1(n15436), .IN2(n15437), .Q(n15435) );
  INVX0 U16056 ( .INP(n15438), .ZN(n15437) );
  OR2X1 U16057 ( .IN1(n4368), .IN2(test_so54), .Q(n15438) );
  AND2X1 U16058 ( .IN1(n8704), .IN2(g6573), .Q(n15436) );
  AND2X1 U16059 ( .IN1(n8703), .IN2(g6782), .Q(n15434) );
  OR2X1 U16060 ( .IN1(n15439), .IN2(n15440), .Q(g22151) );
  AND2X1 U16061 ( .IN1(n15376), .IN2(g1543), .Q(n15440) );
  AND2X1 U16062 ( .IN1(n11800), .IN2(n15377), .Q(n15439) );
  OR2X1 U16063 ( .IN1(n15441), .IN2(n15442), .Q(g22150) );
  AND2X1 U16064 ( .IN1(n14850), .IN2(g1538), .Q(n15442) );
  AND2X1 U16065 ( .IN1(n15359), .IN2(n4288), .Q(n15441) );
  OR2X1 U16066 ( .IN1(n15443), .IN2(n15444), .Q(g22149) );
  AND2X1 U16067 ( .IN1(n15406), .IN2(g1512), .Q(n15444) );
  AND2X1 U16068 ( .IN1(n15405), .IN2(n4378), .Q(n15443) );
  OR2X1 U16069 ( .IN1(n15445), .IN2(n15446), .Q(g22148) );
  AND2X1 U16070 ( .IN1(n15447), .IN2(g852), .Q(n15446) );
  AND2X1 U16071 ( .IN1(n15414), .IN2(n10629), .Q(n15445) );
  OR2X1 U16072 ( .IN1(n15448), .IN2(n15449), .Q(g22147) );
  AND2X1 U16073 ( .IN1(n14852), .IN2(g847), .Q(n15449) );
  AND2X1 U16074 ( .IN1(n11924), .IN2(n15383), .Q(n15448) );
  OR2X1 U16075 ( .IN1(n15450), .IN2(n15451), .Q(g22146) );
  INVX0 U16076 ( .INP(n15452), .ZN(n15451) );
  OR2X1 U16077 ( .IN1(n15453), .IN2(n9024), .Q(n15452) );
  AND2X1 U16078 ( .IN1(n15453), .IN2(n4375), .Q(n15450) );
  OR2X1 U16079 ( .IN1(n15454), .IN2(n15455), .Q(g22145) );
  INVX0 U16080 ( .INP(n15456), .ZN(n15455) );
  OR2X1 U16081 ( .IN1(n15414), .IN2(n9025), .Q(n15456) );
  AND2X1 U16082 ( .IN1(n15414), .IN2(n4379), .Q(n15454) );
  OR2X1 U16083 ( .IN1(n15457), .IN2(n15458), .Q(g22143) );
  AND2X1 U16084 ( .IN1(n14854), .IN2(g162), .Q(n15458) );
  AND2X1 U16085 ( .IN1(n15420), .IN2(n10674), .Q(n15457) );
  OR2X1 U16086 ( .IN1(n15459), .IN2(n15460), .Q(g22142) );
  AND2X1 U16087 ( .IN1(n15461), .IN2(g134), .Q(n15460) );
  AND2X1 U16088 ( .IN1(n15462), .IN2(n4376), .Q(n15459) );
  OR2X1 U16089 ( .IN1(n15463), .IN2(n15464), .Q(g22141) );
  AND2X1 U16090 ( .IN1(n14854), .IN2(g129), .Q(n15464) );
  AND2X1 U16091 ( .IN1(n4380), .IN2(n15420), .Q(n15463) );
  OR2X1 U16092 ( .IN1(n15465), .IN2(n15466), .Q(g22140) );
  INVX0 U16093 ( .INP(n15467), .ZN(n15466) );
  OR2X1 U16094 ( .IN1(n15368), .IN2(n8984), .Q(n15467) );
  AND2X1 U16095 ( .IN1(n15368), .IN2(n4287), .Q(n15465) );
  OR2X1 U16096 ( .IN1(n15468), .IN2(n15469), .Q(g22139) );
  AND2X1 U16097 ( .IN1(n15362), .IN2(g2231), .Q(n15469) );
  AND2X1 U16098 ( .IN1(n15353), .IN2(n4563), .Q(n15468) );
  OR2X1 U16099 ( .IN1(n15470), .IN2(n15471), .Q(g22138) );
  AND2X1 U16100 ( .IN1(n14848), .IN2(g2226), .Q(n15471) );
  AND2X1 U16101 ( .IN1(n15347), .IN2(n4555), .Q(n15470) );
  OR2X1 U16102 ( .IN1(n15472), .IN2(n15473), .Q(g22132) );
  AND2X1 U16103 ( .IN1(n15406), .IN2(g1542), .Q(n15473) );
  AND2X1 U16104 ( .IN1(n15405), .IN2(n11800), .Q(n15472) );
  INVX0 U16105 ( .INP(n10760), .ZN(n11800) );
  OR2X1 U16106 ( .IN1(n15474), .IN2(n15475), .Q(n10760) );
  OR2X1 U16107 ( .IN1(n15476), .IN2(n15477), .Q(n15475) );
  AND2X1 U16108 ( .IN1(n8700), .IN2(g1547), .Q(n15477) );
  AND2X1 U16109 ( .IN1(n8702), .IN2(g6573), .Q(n15476) );
  AND2X1 U16110 ( .IN1(n8701), .IN2(g6782), .Q(n15474) );
  OR2X1 U16111 ( .IN1(n15478), .IN2(n15479), .Q(g22131) );
  AND2X1 U16112 ( .IN1(n15376), .IN2(g1540), .Q(n15479) );
  AND2X1 U16113 ( .IN1(n15377), .IN2(n4288), .Q(n15478) );
  OR2X1 U16114 ( .IN1(n15480), .IN2(n15481), .Q(g22130) );
  AND2X1 U16115 ( .IN1(n14850), .IN2(g1535), .Q(n15481) );
  AND2X1 U16116 ( .IN1(n15359), .IN2(n4565), .Q(n15480) );
  OR2X1 U16117 ( .IN1(n15482), .IN2(n15483), .Q(g22129) );
  AND2X1 U16118 ( .IN1(n15484), .IN2(g851), .Q(n15483) );
  AND2X1 U16119 ( .IN1(n15453), .IN2(n10629), .Q(n15482) );
  INVX0 U16120 ( .INP(n13868), .ZN(n10629) );
  OR2X1 U16121 ( .IN1(n15485), .IN2(n15486), .Q(n13868) );
  OR2X1 U16122 ( .IN1(n15487), .IN2(n15488), .Q(n15486) );
  AND2X1 U16123 ( .IN1(n8716), .IN2(g6368), .Q(n15488) );
  AND2X1 U16124 ( .IN1(n8715), .IN2(g6518), .Q(n15487) );
  AND2X1 U16125 ( .IN1(n8714), .IN2(test_so31), .Q(n15485) );
  OR2X1 U16126 ( .IN1(n15489), .IN2(n15490), .Q(g22128) );
  AND2X1 U16127 ( .IN1(n15447), .IN2(g849), .Q(n15490) );
  AND2X1 U16128 ( .IN1(n11924), .IN2(n15414), .Q(n15489) );
  OR2X1 U16129 ( .IN1(n15491), .IN2(n15492), .Q(g22127) );
  INVX0 U16130 ( .INP(n15493), .ZN(n15492) );
  OR2X1 U16131 ( .IN1(n15383), .IN2(n8652), .Q(n15493) );
  AND2X1 U16132 ( .IN1(n4289), .IN2(n15383), .Q(n15491) );
  OR2X1 U16133 ( .IN1(n15494), .IN2(n15495), .Q(g22126) );
  INVX0 U16134 ( .INP(n15496), .ZN(n15495) );
  OR2X1 U16135 ( .IN1(n15453), .IN2(n9026), .Q(n15496) );
  AND2X1 U16136 ( .IN1(n15453), .IN2(n4379), .Q(n15494) );
  OR2X1 U16137 ( .IN1(n15497), .IN2(n15498), .Q(g22125) );
  AND2X1 U16138 ( .IN1(n15461), .IN2(g164), .Q(n15498) );
  AND2X1 U16139 ( .IN1(n15462), .IN2(n10674), .Q(n15497) );
  OR2X1 U16140 ( .IN1(n15499), .IN2(n15500), .Q(g22124) );
  AND2X1 U16141 ( .IN1(n14854), .IN2(g159), .Q(n15500) );
  AND2X1 U16142 ( .IN1(n12005), .IN2(n15420), .Q(n15499) );
  OR2X1 U16143 ( .IN1(n15501), .IN2(n15502), .Q(g22123) );
  AND2X1 U16144 ( .IN1(n15503), .IN2(g133), .Q(n15502) );
  AND2X1 U16145 ( .IN1(n15504), .IN2(n4376), .Q(n15501) );
  OR2X1 U16146 ( .IN1(n15505), .IN2(n15506), .Q(g22122) );
  AND2X1 U16147 ( .IN1(n15461), .IN2(g131), .Q(n15506) );
  AND2X1 U16148 ( .IN1(n15462), .IN2(n4380), .Q(n15505) );
  OR2X1 U16149 ( .IN1(n15507), .IN2(n15508), .Q(g22117) );
  AND2X1 U16150 ( .IN1(n15386), .IN2(g2230), .Q(n15508) );
  AND2X1 U16151 ( .IN1(n15368), .IN2(n4563), .Q(n15507) );
  OR2X1 U16152 ( .IN1(n15509), .IN2(n15510), .Q(g22116) );
  AND2X1 U16153 ( .IN1(n15362), .IN2(g2228), .Q(n15510) );
  AND2X1 U16154 ( .IN1(n15353), .IN2(n4555), .Q(n15509) );
  OR2X1 U16155 ( .IN1(n15511), .IN2(n15512), .Q(g22115) );
  INVX0 U16156 ( .INP(n15513), .ZN(n15512) );
  OR2X1 U16157 ( .IN1(n15347), .IN2(n8630), .Q(n15513) );
  AND2X1 U16158 ( .IN1(n15347), .IN2(n4325), .Q(n15511) );
  OR2X1 U16159 ( .IN1(n15514), .IN2(n15515), .Q(g22114) );
  AND2X1 U16160 ( .IN1(n15406), .IN2(g1539), .Q(n15515) );
  AND2X1 U16161 ( .IN1(n15405), .IN2(n4288), .Q(n15514) );
  OR2X1 U16162 ( .IN1(n15516), .IN2(n15517), .Q(g22113) );
  AND2X1 U16163 ( .IN1(n15377), .IN2(n4565), .Q(n15517) );
  AND2X1 U16164 ( .IN1(test_so53), .IN2(n15376), .Q(n15516) );
  OR2X1 U16165 ( .IN1(n15518), .IN2(n15519), .Q(g22112) );
  AND2X1 U16166 ( .IN1(n14850), .IN2(g1532), .Q(n15519) );
  AND2X1 U16167 ( .IN1(n15359), .IN2(n4557), .Q(n15518) );
  OR2X1 U16168 ( .IN1(n15520), .IN2(n15521), .Q(g22106) );
  AND2X1 U16169 ( .IN1(n15484), .IN2(g848), .Q(n15521) );
  AND2X1 U16170 ( .IN1(n15453), .IN2(n11924), .Q(n15520) );
  INVX0 U16171 ( .INP(n10800), .ZN(n11924) );
  OR2X1 U16172 ( .IN1(n15522), .IN2(n15523), .Q(n10800) );
  OR2X1 U16173 ( .IN1(n15524), .IN2(n15525), .Q(n15523) );
  AND2X1 U16174 ( .IN1(n8713), .IN2(g6368), .Q(n15525) );
  AND2X1 U16175 ( .IN1(n8712), .IN2(g6518), .Q(n15524) );
  AND2X1 U16176 ( .IN1(n8711), .IN2(test_so31), .Q(n15522) );
  OR2X1 U16177 ( .IN1(n15526), .IN2(n15527), .Q(g22105) );
  INVX0 U16178 ( .INP(n15528), .ZN(n15527) );
  OR2X1 U16179 ( .IN1(n15414), .IN2(n9012), .Q(n15528) );
  AND2X1 U16180 ( .IN1(n4289), .IN2(n15414), .Q(n15526) );
  OR2X1 U16181 ( .IN1(n15529), .IN2(n15530), .Q(g22104) );
  AND2X1 U16182 ( .IN1(n14852), .IN2(g841), .Q(n15530) );
  AND2X1 U16183 ( .IN1(n15383), .IN2(n4567), .Q(n15529) );
  OR2X1 U16184 ( .IN1(n15531), .IN2(n15532), .Q(g22103) );
  AND2X1 U16185 ( .IN1(n15504), .IN2(n10674), .Q(n15532) );
  INVX0 U16186 ( .INP(n13975), .ZN(n10674) );
  OR2X1 U16187 ( .IN1(n15533), .IN2(n15534), .Q(n13975) );
  OR2X1 U16188 ( .IN1(n15535), .IN2(n15536), .Q(n15534) );
  AND2X1 U16189 ( .IN1(n8725), .IN2(g165), .Q(n15536) );
  AND2X1 U16190 ( .IN1(n8727), .IN2(g6231), .Q(n15535) );
  AND2X1 U16191 ( .IN1(n8726), .IN2(g6313), .Q(n15533) );
  AND2X1 U16192 ( .IN1(test_so12), .IN2(n15503), .Q(n15531) );
  OR2X1 U16193 ( .IN1(n15537), .IN2(n15538), .Q(g22102) );
  AND2X1 U16194 ( .IN1(n15461), .IN2(g161), .Q(n15538) );
  AND2X1 U16195 ( .IN1(n12005), .IN2(n15462), .Q(n15537) );
  OR2X1 U16196 ( .IN1(n15539), .IN2(n15540), .Q(g22101) );
  AND2X1 U16197 ( .IN1(n14854), .IN2(g156), .Q(n15540) );
  AND2X1 U16198 ( .IN1(n4290), .IN2(n15420), .Q(n15539) );
  OR2X1 U16199 ( .IN1(n15541), .IN2(n15542), .Q(g22100) );
  AND2X1 U16200 ( .IN1(n15503), .IN2(g130), .Q(n15542) );
  AND2X1 U16201 ( .IN1(n15504), .IN2(n4380), .Q(n15541) );
  OR2X1 U16202 ( .IN1(n15543), .IN2(n15544), .Q(g22099) );
  AND2X1 U16203 ( .IN1(n15386), .IN2(g2227), .Q(n15544) );
  AND2X1 U16204 ( .IN1(n15368), .IN2(n4555), .Q(n15543) );
  OR2X1 U16205 ( .IN1(n15545), .IN2(n15546), .Q(g22098) );
  AND2X1 U16206 ( .IN1(n15353), .IN2(n4325), .Q(n15546) );
  AND2X1 U16207 ( .IN1(test_so74), .IN2(n15362), .Q(n15545) );
  OR2X1 U16208 ( .IN1(n15547), .IN2(n15548), .Q(g22097) );
  INVX0 U16209 ( .INP(n15549), .ZN(n15548) );
  OR2X1 U16210 ( .IN1(n15347), .IN2(n8631), .Q(n15549) );
  AND2X1 U16211 ( .IN1(n15347), .IN2(n4389), .Q(n15547) );
  OR2X1 U16212 ( .IN1(n15550), .IN2(n15551), .Q(g22092) );
  AND2X1 U16213 ( .IN1(n15406), .IN2(g1536), .Q(n15551) );
  AND2X1 U16214 ( .IN1(n15405), .IN2(n4565), .Q(n15550) );
  OR2X1 U16215 ( .IN1(n15552), .IN2(n15553), .Q(g22091) );
  AND2X1 U16216 ( .IN1(n15376), .IN2(g1534), .Q(n15553) );
  AND2X1 U16217 ( .IN1(n15377), .IN2(n4557), .Q(n15552) );
  OR2X1 U16218 ( .IN1(n15554), .IN2(n15555), .Q(g22090) );
  AND2X1 U16219 ( .IN1(n14850), .IN2(g1529), .Q(n15555) );
  AND2X1 U16220 ( .IN1(n15359), .IN2(n4326), .Q(n15554) );
  OR2X1 U16221 ( .IN1(n15556), .IN2(n15557), .Q(g22089) );
  INVX0 U16222 ( .INP(n15558), .ZN(n15557) );
  OR2X1 U16223 ( .IN1(n15453), .IN2(n9013), .Q(n15558) );
  AND2X1 U16224 ( .IN1(n4289), .IN2(n15453), .Q(n15556) );
  OR2X1 U16225 ( .IN1(n15559), .IN2(n15560), .Q(g22088) );
  AND2X1 U16226 ( .IN1(n15447), .IN2(g843), .Q(n15560) );
  AND2X1 U16227 ( .IN1(n15414), .IN2(n4567), .Q(n15559) );
  OR2X1 U16228 ( .IN1(n15561), .IN2(n15562), .Q(g22087) );
  AND2X1 U16229 ( .IN1(n14852), .IN2(g838), .Q(n15562) );
  AND2X1 U16230 ( .IN1(n15383), .IN2(n4559), .Q(n15561) );
  OR2X1 U16231 ( .IN1(n15563), .IN2(n15564), .Q(g22081) );
  AND2X1 U16232 ( .IN1(n15503), .IN2(g160), .Q(n15564) );
  AND2X1 U16233 ( .IN1(n15504), .IN2(n12005), .Q(n15563) );
  INVX0 U16234 ( .INP(n10824), .ZN(n12005) );
  OR2X1 U16235 ( .IN1(n15565), .IN2(n15566), .Q(n10824) );
  OR2X1 U16236 ( .IN1(n15567), .IN2(n15568), .Q(n15566) );
  AND2X1 U16237 ( .IN1(n8722), .IN2(g165), .Q(n15568) );
  AND2X1 U16238 ( .IN1(n8724), .IN2(g6231), .Q(n15567) );
  AND2X1 U16239 ( .IN1(n8723), .IN2(g6313), .Q(n15565) );
  OR2X1 U16240 ( .IN1(n15569), .IN2(n15570), .Q(g22080) );
  AND2X1 U16241 ( .IN1(n15461), .IN2(g158), .Q(n15570) );
  AND2X1 U16242 ( .IN1(n4290), .IN2(n15462), .Q(n15569) );
  OR2X1 U16243 ( .IN1(n15571), .IN2(n15572), .Q(g22079) );
  AND2X1 U16244 ( .IN1(n14854), .IN2(g153), .Q(n15572) );
  AND2X1 U16245 ( .IN1(n15420), .IN2(n4569), .Q(n15571) );
  OR2X1 U16246 ( .IN1(n15573), .IN2(n15574), .Q(g22078) );
  INVX0 U16247 ( .INP(n15575), .ZN(n15574) );
  OR2X1 U16248 ( .IN1(n15368), .IN2(n8989), .Q(n15575) );
  AND2X1 U16249 ( .IN1(n15368), .IN2(n4325), .Q(n15573) );
  OR2X1 U16250 ( .IN1(n15576), .IN2(n15577), .Q(g22077) );
  INVX0 U16251 ( .INP(n15578), .ZN(n15577) );
  OR2X1 U16252 ( .IN1(n15353), .IN2(n8990), .Q(n15578) );
  AND2X1 U16253 ( .IN1(n15353), .IN2(n4389), .Q(n15576) );
  OR2X1 U16254 ( .IN1(n15579), .IN2(n15580), .Q(g22076) );
  INVX0 U16255 ( .INP(n15581), .ZN(n15580) );
  OR2X1 U16256 ( .IN1(n15347), .IN2(n8632), .Q(n15581) );
  AND2X1 U16257 ( .IN1(n15347), .IN2(n4319), .Q(n15579) );
  INVX0 U16258 ( .INP(n14848), .ZN(n15347) );
  OR2X1 U16259 ( .IN1(n4367), .IN2(n9091), .Q(n14848) );
  OR2X1 U16260 ( .IN1(n15582), .IN2(n15583), .Q(g22075) );
  AND2X1 U16261 ( .IN1(n15406), .IN2(g1533), .Q(n15583) );
  AND2X1 U16262 ( .IN1(n15405), .IN2(n4557), .Q(n15582) );
  OR2X1 U16263 ( .IN1(n15584), .IN2(n15585), .Q(g22074) );
  AND2X1 U16264 ( .IN1(n15376), .IN2(g1531), .Q(n15585) );
  AND2X1 U16265 ( .IN1(n15377), .IN2(n4326), .Q(n15584) );
  OR2X1 U16266 ( .IN1(n15586), .IN2(n15587), .Q(g22073) );
  AND2X1 U16267 ( .IN1(n14850), .IN2(g1526), .Q(n15587) );
  AND2X1 U16268 ( .IN1(n15359), .IN2(n4390), .Q(n15586) );
  OR2X1 U16269 ( .IN1(n15588), .IN2(n15589), .Q(g22068) );
  AND2X1 U16270 ( .IN1(n15484), .IN2(g842), .Q(n15589) );
  AND2X1 U16271 ( .IN1(n15453), .IN2(n4567), .Q(n15588) );
  OR2X1 U16272 ( .IN1(n15590), .IN2(n15591), .Q(g22067) );
  AND2X1 U16273 ( .IN1(n15447), .IN2(g840), .Q(n15591) );
  AND2X1 U16274 ( .IN1(n15414), .IN2(n4559), .Q(n15590) );
  OR2X1 U16275 ( .IN1(n15592), .IN2(n15593), .Q(g22066) );
  INVX0 U16276 ( .INP(n15594), .ZN(n15593) );
  OR2X1 U16277 ( .IN1(n15383), .IN2(n8655), .Q(n15594) );
  AND2X1 U16278 ( .IN1(n4327), .IN2(n15383), .Q(n15592) );
  OR2X1 U16279 ( .IN1(n15595), .IN2(n15596), .Q(g22065) );
  AND2X1 U16280 ( .IN1(n15503), .IN2(g157), .Q(n15596) );
  AND2X1 U16281 ( .IN1(n4290), .IN2(n15504), .Q(n15595) );
  OR2X1 U16282 ( .IN1(n15597), .IN2(n15598), .Q(g22064) );
  AND2X1 U16283 ( .IN1(n15461), .IN2(g155), .Q(n15598) );
  AND2X1 U16284 ( .IN1(n15462), .IN2(n4569), .Q(n15597) );
  OR2X1 U16285 ( .IN1(n15599), .IN2(n15600), .Q(g22063) );
  AND2X1 U16286 ( .IN1(n14854), .IN2(g150), .Q(n15600) );
  AND2X1 U16287 ( .IN1(n15420), .IN2(n4561), .Q(n15599) );
  OR2X1 U16288 ( .IN1(n15601), .IN2(n15602), .Q(g22061) );
  INVX0 U16289 ( .INP(n15603), .ZN(n15602) );
  OR2X1 U16290 ( .IN1(n15368), .IN2(n8991), .Q(n15603) );
  AND2X1 U16291 ( .IN1(n15368), .IN2(n4389), .Q(n15601) );
  OR2X1 U16292 ( .IN1(n15604), .IN2(n15605), .Q(g22060) );
  INVX0 U16293 ( .INP(n15606), .ZN(n15605) );
  OR2X1 U16294 ( .IN1(n15353), .IN2(n8992), .Q(n15606) );
  AND2X1 U16295 ( .IN1(n15353), .IN2(n4319), .Q(n15604) );
  INVX0 U16296 ( .INP(n15362), .ZN(n15353) );
  OR2X1 U16297 ( .IN1(n9091), .IN2(n9119), .Q(n15362) );
  OR2X1 U16298 ( .IN1(n15607), .IN2(n15608), .Q(g22059) );
  AND2X1 U16299 ( .IN1(n15406), .IN2(g1530), .Q(n15608) );
  AND2X1 U16300 ( .IN1(n15405), .IN2(n4326), .Q(n15607) );
  OR2X1 U16301 ( .IN1(n15609), .IN2(n15610), .Q(g22058) );
  AND2X1 U16302 ( .IN1(n15376), .IN2(g1528), .Q(n15610) );
  AND2X1 U16303 ( .IN1(n15377), .IN2(n4390), .Q(n15609) );
  OR2X1 U16304 ( .IN1(n15611), .IN2(n15612), .Q(g22057) );
  AND2X1 U16305 ( .IN1(n14850), .IN2(g1523), .Q(n15612) );
  AND2X1 U16306 ( .IN1(n15359), .IN2(n4320), .Q(n15611) );
  INVX0 U16307 ( .INP(n14850), .ZN(n15359) );
  OR2X1 U16308 ( .IN1(n4368), .IN2(n9090), .Q(n14850) );
  OR2X1 U16309 ( .IN1(n15613), .IN2(n15614), .Q(g22056) );
  AND2X1 U16310 ( .IN1(n15453), .IN2(n4559), .Q(n15614) );
  AND2X1 U16311 ( .IN1(test_so32), .IN2(n15484), .Q(n15613) );
  OR2X1 U16312 ( .IN1(n15615), .IN2(n15616), .Q(g22055) );
  INVX0 U16313 ( .INP(n15617), .ZN(n15616) );
  OR2X1 U16314 ( .IN1(n15414), .IN2(n9017), .Q(n15617) );
  AND2X1 U16315 ( .IN1(n4327), .IN2(n15414), .Q(n15615) );
  OR2X1 U16316 ( .IN1(n15618), .IN2(n15619), .Q(g22054) );
  INVX0 U16317 ( .INP(n15620), .ZN(n15619) );
  OR2X1 U16318 ( .IN1(n15383), .IN2(n8656), .Q(n15620) );
  AND2X1 U16319 ( .IN1(n15383), .IN2(n4391), .Q(n15618) );
  OR2X1 U16320 ( .IN1(n15621), .IN2(n15622), .Q(g22049) );
  AND2X1 U16321 ( .IN1(n15503), .IN2(g154), .Q(n15622) );
  AND2X1 U16322 ( .IN1(n15504), .IN2(n4569), .Q(n15621) );
  OR2X1 U16323 ( .IN1(n15623), .IN2(n15624), .Q(g22048) );
  AND2X1 U16324 ( .IN1(n15461), .IN2(g152), .Q(n15624) );
  AND2X1 U16325 ( .IN1(n15462), .IN2(n4561), .Q(n15623) );
  OR2X1 U16326 ( .IN1(n15625), .IN2(n15626), .Q(g22047) );
  AND2X1 U16327 ( .IN1(n14854), .IN2(g147), .Q(n15626) );
  AND2X1 U16328 ( .IN1(n4328), .IN2(n15420), .Q(n15625) );
  OR2X1 U16329 ( .IN1(n15627), .IN2(n15628), .Q(g22045) );
  INVX0 U16330 ( .INP(n15629), .ZN(n15628) );
  OR2X1 U16331 ( .IN1(n15368), .IN2(n8993), .Q(n15629) );
  AND2X1 U16332 ( .IN1(n15368), .IN2(n4319), .Q(n15627) );
  INVX0 U16333 ( .INP(n15386), .ZN(n15368) );
  OR2X1 U16334 ( .IN1(n4324), .IN2(n9091), .Q(n15386) );
  OR2X1 U16335 ( .IN1(n15630), .IN2(n15631), .Q(g22044) );
  AND2X1 U16336 ( .IN1(n15406), .IN2(g1527), .Q(n15631) );
  AND2X1 U16337 ( .IN1(n15405), .IN2(n4390), .Q(n15630) );
  OR2X1 U16338 ( .IN1(n15632), .IN2(n15633), .Q(g22043) );
  AND2X1 U16339 ( .IN1(n15376), .IN2(g1525), .Q(n15633) );
  AND2X1 U16340 ( .IN1(n15377), .IN2(n4320), .Q(n15632) );
  INVX0 U16341 ( .INP(n15376), .ZN(n15377) );
  OR2X1 U16342 ( .IN1(n4515), .IN2(n9090), .Q(n15376) );
  OR2X1 U16343 ( .IN1(n15634), .IN2(n15635), .Q(g22042) );
  INVX0 U16344 ( .INP(n15636), .ZN(n15635) );
  OR2X1 U16345 ( .IN1(n15453), .IN2(n9018), .Q(n15636) );
  AND2X1 U16346 ( .IN1(n4327), .IN2(n15453), .Q(n15634) );
  OR2X1 U16347 ( .IN1(n15637), .IN2(n15638), .Q(g22041) );
  INVX0 U16348 ( .INP(n15639), .ZN(n15638) );
  OR2X1 U16349 ( .IN1(n15414), .IN2(n9019), .Q(n15639) );
  AND2X1 U16350 ( .IN1(n15414), .IN2(n4391), .Q(n15637) );
  OR2X1 U16351 ( .IN1(n15640), .IN2(n15641), .Q(g22040) );
  INVX0 U16352 ( .INP(n15642), .ZN(n15641) );
  OR2X1 U16353 ( .IN1(n15383), .IN2(n8657), .Q(n15642) );
  AND2X1 U16354 ( .IN1(n4321), .IN2(n15383), .Q(n15640) );
  INVX0 U16355 ( .INP(n14852), .ZN(n15383) );
  OR2X1 U16356 ( .IN1(n9089), .IN2(n9118), .Q(n14852) );
  OR2X1 U16357 ( .IN1(n15643), .IN2(n15644), .Q(g22039) );
  AND2X1 U16358 ( .IN1(n15503), .IN2(g151), .Q(n15644) );
  AND2X1 U16359 ( .IN1(n15504), .IN2(n4561), .Q(n15643) );
  OR2X1 U16360 ( .IN1(n15645), .IN2(n15646), .Q(g22038) );
  AND2X1 U16361 ( .IN1(n15461), .IN2(g149), .Q(n15646) );
  AND2X1 U16362 ( .IN1(n4328), .IN2(n15462), .Q(n15645) );
  OR2X1 U16363 ( .IN1(n15647), .IN2(n15648), .Q(g22037) );
  AND2X1 U16364 ( .IN1(n15420), .IN2(n4392), .Q(n15648) );
  AND2X1 U16365 ( .IN1(test_so11), .IN2(n14854), .Q(n15647) );
  OR2X1 U16366 ( .IN1(n15649), .IN2(n15650), .Q(g22035) );
  AND2X1 U16367 ( .IN1(n15406), .IN2(g1524), .Q(n15650) );
  AND2X1 U16368 ( .IN1(n15405), .IN2(n4320), .Q(n15649) );
  INVX0 U16369 ( .INP(n15406), .ZN(n15405) );
  OR2X1 U16370 ( .IN1(n4317), .IN2(n9090), .Q(n15406) );
  OR2X1 U16371 ( .IN1(n15651), .IN2(n15652), .Q(g22034) );
  INVX0 U16372 ( .INP(n15653), .ZN(n15652) );
  OR2X1 U16373 ( .IN1(n15453), .IN2(n9020), .Q(n15653) );
  AND2X1 U16374 ( .IN1(n15453), .IN2(n4391), .Q(n15651) );
  OR2X1 U16375 ( .IN1(n15654), .IN2(n15655), .Q(g22033) );
  INVX0 U16376 ( .INP(n15656), .ZN(n15655) );
  OR2X1 U16377 ( .IN1(n15414), .IN2(n9021), .Q(n15656) );
  AND2X1 U16378 ( .IN1(n4321), .IN2(n15414), .Q(n15654) );
  INVX0 U16379 ( .INP(n15447), .ZN(n15414) );
  OR2X1 U16380 ( .IN1(n4312), .IN2(n9089), .Q(n15447) );
  OR2X1 U16381 ( .IN1(n15657), .IN2(n15658), .Q(g22032) );
  AND2X1 U16382 ( .IN1(n15503), .IN2(g148), .Q(n15658) );
  AND2X1 U16383 ( .IN1(n4328), .IN2(n15504), .Q(n15657) );
  OR2X1 U16384 ( .IN1(n15659), .IN2(n15660), .Q(g22031) );
  AND2X1 U16385 ( .IN1(n15461), .IN2(g146), .Q(n15660) );
  AND2X1 U16386 ( .IN1(n15462), .IN2(n4392), .Q(n15659) );
  OR2X1 U16387 ( .IN1(n15661), .IN2(n15662), .Q(g22030) );
  AND2X1 U16388 ( .IN1(n14854), .IN2(g141), .Q(n15662) );
  AND2X1 U16389 ( .IN1(n4322), .IN2(n15420), .Q(n15661) );
  INVX0 U16390 ( .INP(n14854), .ZN(n15420) );
  OR2X1 U16391 ( .IN1(n4369), .IN2(n9088), .Q(n14854) );
  OR2X1 U16392 ( .IN1(n15663), .IN2(n15664), .Q(g22029) );
  INVX0 U16393 ( .INP(n15665), .ZN(n15664) );
  OR2X1 U16394 ( .IN1(n15453), .IN2(n9022), .Q(n15665) );
  AND2X1 U16395 ( .IN1(n4321), .IN2(n15453), .Q(n15663) );
  INVX0 U16396 ( .INP(n15484), .ZN(n15453) );
  OR2X1 U16397 ( .IN1(n4323), .IN2(n9089), .Q(n15484) );
  OR2X1 U16398 ( .IN1(n15666), .IN2(n15667), .Q(g22028) );
  AND2X1 U16399 ( .IN1(n15503), .IN2(g145), .Q(n15667) );
  AND2X1 U16400 ( .IN1(n15504), .IN2(n4392), .Q(n15666) );
  OR2X1 U16401 ( .IN1(n15668), .IN2(n15669), .Q(g22027) );
  AND2X1 U16402 ( .IN1(n15461), .IN2(g143), .Q(n15669) );
  AND2X1 U16403 ( .IN1(n4322), .IN2(n15462), .Q(n15668) );
  INVX0 U16404 ( .INP(n15461), .ZN(n15462) );
  OR2X1 U16405 ( .IN1(n4512), .IN2(n9088), .Q(n15461) );
  AND2X1 U16406 ( .IN1(n15670), .IN2(n9662), .Q(g22026) );
  AND2X1 U16407 ( .IN1(n9510), .IN2(n16489), .Q(n9662) );
  OR2X1 U16408 ( .IN1(n15671), .IN2(n15672), .Q(n9510) );
  INVX0 U16409 ( .INP(n15673), .ZN(n15672) );
  AND2X1 U16410 ( .IN1(n15674), .IN2(n4330), .Q(n15673) );
  AND2X1 U16411 ( .IN1(n4182), .IN2(n4431), .Q(n15674) );
  OR2X1 U16412 ( .IN1(n15675), .IN2(n15676), .Q(n15671) );
  OR2X1 U16413 ( .IN1(n4355), .IN2(g2900), .Q(n15676) );
  OR2X1 U16414 ( .IN1(n9081), .IN2(n4423), .Q(n15675) );
  XOR2X1 U16415 ( .IN1(n9664), .IN2(n9081), .Q(n15670) );
  OR2X1 U16416 ( .IN1(n4330), .IN2(n4423), .Q(n9664) );
  OR2X1 U16417 ( .IN1(n15677), .IN2(n15678), .Q(g22025) );
  AND2X1 U16418 ( .IN1(n15503), .IN2(g142), .Q(n15678) );
  AND2X1 U16419 ( .IN1(n4322), .IN2(n15504), .Q(n15677) );
  INVX0 U16420 ( .INP(n15503), .ZN(n15504) );
  OR2X1 U16421 ( .IN1(n4318), .IN2(n9088), .Q(n15503) );
  AND2X1 U16422 ( .IN1(n15679), .IN2(n15680), .Q(g21974) );
  INVX0 U16423 ( .INP(n15681), .ZN(n15680) );
  AND2X1 U16424 ( .IN1(n15682), .IN2(n4472), .Q(n15681) );
  OR2X1 U16425 ( .IN1(n15683), .IN2(n4398), .Q(n15682) );
  AND2X1 U16426 ( .IN1(n15018), .IN2(n12737), .Q(n15679) );
  OR2X1 U16427 ( .IN1(n15683), .IN2(n15684), .Q(n15018) );
  OR2X1 U16428 ( .IN1(n4472), .IN2(n4398), .Q(n15684) );
  AND2X1 U16429 ( .IN1(n15685), .IN2(n15686), .Q(g21972) );
  INVX0 U16430 ( .INP(n15687), .ZN(n15686) );
  AND2X1 U16431 ( .IN1(n15688), .IN2(n4474), .Q(n15687) );
  OR2X1 U16432 ( .IN1(n15689), .IN2(n4400), .Q(n15688) );
  AND2X1 U16433 ( .IN1(n15024), .IN2(n12741), .Q(n15685) );
  OR2X1 U16434 ( .IN1(n15689), .IN2(n15690), .Q(n15024) );
  OR2X1 U16435 ( .IN1(n4474), .IN2(n4400), .Q(n15690) );
  OR2X1 U16436 ( .IN1(n15691), .IN2(n15692), .Q(g21970) );
  AND2X1 U16437 ( .IN1(n12782), .IN2(g2560), .Q(n15692) );
  OR2X1 U16438 ( .IN1(n15693), .IN2(n15694), .Q(n12782) );
  OR2X1 U16439 ( .IN1(n15695), .IN2(n15696), .Q(n15694) );
  AND2X1 U16440 ( .IN1(g7264), .IN2(g2516), .Q(n15696) );
  AND2X1 U16441 ( .IN1(n4606), .IN2(g2519), .Q(n15695) );
  AND2X1 U16442 ( .IN1(g5555), .IN2(g2513), .Q(n15693) );
  AND2X1 U16443 ( .IN1(test_so87), .IN2(n4463), .Q(n15691) );
  AND2X1 U16444 ( .IN1(n15697), .IN2(n15698), .Q(g21969) );
  INVX0 U16445 ( .INP(n15699), .ZN(n15698) );
  AND2X1 U16446 ( .IN1(n15700), .IN2(n4476), .Q(n15699) );
  OR2X1 U16447 ( .IN1(n15701), .IN2(n4402), .Q(n15700) );
  AND2X1 U16448 ( .IN1(n15030), .IN2(n12745), .Q(n15697) );
  OR2X1 U16449 ( .IN1(n15701), .IN2(n15702), .Q(n15030) );
  OR2X1 U16450 ( .IN1(n4476), .IN2(n4402), .Q(n15702) );
  OR2X1 U16451 ( .IN1(n15703), .IN2(n15704), .Q(g21882) );
  AND2X1 U16452 ( .IN1(n15705), .IN2(g2879), .Q(n15704) );
  AND2X1 U16453 ( .IN1(n4351), .IN2(g2878), .Q(n15703) );
  OR2X1 U16454 ( .IN1(n15706), .IN2(n15707), .Q(g21880) );
  AND2X1 U16455 ( .IN1(n15708), .IN2(g2879), .Q(n15707) );
  AND2X1 U16456 ( .IN1(n4351), .IN2(g2877), .Q(n15706) );
  OR2X1 U16457 ( .IN1(n15709), .IN2(n15710), .Q(g21878) );
  AND2X1 U16458 ( .IN1(n15705), .IN2(n4351), .Q(n15710) );
  XNOR2X1 U16459 ( .IN1(n15711), .IN2(n9518), .Q(n15705) );
  XNOR2X1 U16460 ( .IN1(n15712), .IN2(n15713), .Q(n9518) );
  XOR2X1 U16461 ( .IN1(n15714), .IN2(n15715), .Q(n15713) );
  XNOR2X1 U16462 ( .IN1(g2969), .IN2(n9071), .Q(n15715) );
  XNOR2X1 U16463 ( .IN1(test_so2), .IN2(g2981), .Q(n15714) );
  XOR2X1 U16464 ( .IN1(n15716), .IN2(n15717), .Q(n15712) );
  XNOR2X1 U16465 ( .IN1(g2972), .IN2(n9069), .Q(n15717) );
  XNOR2X1 U16466 ( .IN1(n9067), .IN2(n9068), .Q(n15716) );
  AND2X1 U16467 ( .IN1(test_so4), .IN2(g2879), .Q(n15709) );
  OR2X1 U16468 ( .IN1(n15718), .IN2(n15719), .Q(g21851) );
  AND2X1 U16469 ( .IN1(n15720), .IN2(n4541), .Q(n15719) );
  AND2X1 U16470 ( .IN1(n4298), .IN2(g548), .Q(n15720) );
  AND2X1 U16471 ( .IN1(g499), .IN2(g544), .Q(n15718) );
  OR2X1 U16472 ( .IN1(n15721), .IN2(n14858), .Q(g21847) );
  AND2X1 U16473 ( .IN1(g2624), .IN2(n12265), .Q(n14858) );
  INVX0 U16474 ( .INP(n15722), .ZN(n15721) );
  OR2X1 U16475 ( .IN1(g2624), .IN2(n9050), .Q(n15722) );
  OR2X1 U16476 ( .IN1(n15723), .IN2(n14866), .Q(g21845) );
  AND2X1 U16477 ( .IN1(g1930), .IN2(n12265), .Q(n14866) );
  INVX0 U16478 ( .INP(n15724), .ZN(n15723) );
  OR2X1 U16479 ( .IN1(g1930), .IN2(n9051), .Q(n15724) );
  OR2X1 U16480 ( .IN1(n15725), .IN2(n14890), .Q(g21843) );
  AND2X1 U16481 ( .IN1(g1236), .IN2(n12265), .Q(n14890) );
  INVX0 U16482 ( .INP(n15726), .ZN(n15725) );
  OR2X1 U16483 ( .IN1(g1236), .IN2(n9052), .Q(n15726) );
  OR2X1 U16484 ( .IN1(n15727), .IN2(n14927), .Q(g21842) );
  AND2X1 U16485 ( .IN1(g550), .IN2(n12265), .Q(n14927) );
  OR2X1 U16486 ( .IN1(n15728), .IN2(n15729), .Q(n12265) );
  INVX0 U16487 ( .INP(n15730), .ZN(n15729) );
  AND2X1 U16488 ( .IN1(n4480), .IN2(n9086), .Q(n15730) );
  OR2X1 U16489 ( .IN1(n15199), .IN2(n15731), .Q(n15728) );
  OR2X1 U16490 ( .IN1(n4481), .IN2(n4350), .Q(n15731) );
  OR2X1 U16491 ( .IN1(n15732), .IN2(n15733), .Q(n15199) );
  OR2X1 U16492 ( .IN1(g2993), .IN2(n15734), .Q(n15733) );
  OR2X1 U16493 ( .IN1(n8281), .IN2(g3006), .Q(n15734) );
  OR2X1 U16494 ( .IN1(n15735), .IN2(n15736), .Q(n15732) );
  OR2X1 U16495 ( .IN1(n9092), .IN2(n8282), .Q(n15736) );
  OR2X1 U16496 ( .IN1(test_so98), .IN2(n16493), .Q(n15735) );
  INVX0 U16497 ( .INP(n15737), .ZN(n15727) );
  OR2X1 U16498 ( .IN1(g550), .IN2(n9053), .Q(n15737) );
  OR2X1 U16499 ( .IN1(n15738), .IN2(n15739), .Q(g21346) );
  INVX0 U16500 ( .INP(n15740), .ZN(n15739) );
  OR2X1 U16501 ( .IN1(n15741), .IN2(n16490), .Q(n15740) );
  OR2X1 U16502 ( .IN1(g6447), .IN2(n8546), .Q(n15741) );
  AND2X1 U16503 ( .IN1(n16490), .IN2(DFF_328_n1), .Q(n15738) );
  OR2X1 U16504 ( .IN1(n15742), .IN2(n15743), .Q(g21094) );
  AND2X1 U16505 ( .IN1(n4393), .IN2(n14299), .Q(n15743) );
  AND2X1 U16506 ( .IN1(test_so94), .IN2(n14300), .Q(n15742) );
  OR2X1 U16507 ( .IN1(n15744), .IN2(n15745), .Q(g21082) );
  INVX0 U16508 ( .INP(n15746), .ZN(n15745) );
  OR2X1 U16509 ( .IN1(n14304), .IN2(n8869), .Q(n15746) );
  AND2X1 U16510 ( .IN1(n4393), .IN2(n14304), .Q(n15744) );
  OR2X1 U16511 ( .IN1(n15747), .IN2(n15748), .Q(g21081) );
  INVX0 U16512 ( .INP(n15749), .ZN(n15748) );
  OR2X1 U16513 ( .IN1(n14299), .IN2(n8942), .Q(n15749) );
  AND2X1 U16514 ( .IN1(n14299), .IN2(n4471), .Q(n15747) );
  OR2X1 U16515 ( .IN1(n15750), .IN2(n15751), .Q(g21080) );
  INVX0 U16516 ( .INP(n15752), .ZN(n15751) );
  OR2X1 U16517 ( .IN1(n4149), .IN2(n8950), .Q(n15752) );
  AND2X1 U16518 ( .IN1(n4149), .IN2(n9124), .Q(n15750) );
  OR2X1 U16519 ( .IN1(n15753), .IN2(n15754), .Q(g21075) );
  INVX0 U16520 ( .INP(n15755), .ZN(n15754) );
  OR2X1 U16521 ( .IN1(n14312), .IN2(n8870), .Q(n15755) );
  AND2X1 U16522 ( .IN1(n4393), .IN2(n14312), .Q(n15753) );
  OR2X1 U16523 ( .IN1(n15756), .IN2(n15757), .Q(g21074) );
  INVX0 U16524 ( .INP(n15758), .ZN(n15757) );
  OR2X1 U16525 ( .IN1(n14304), .IN2(n8871), .Q(n15758) );
  AND2X1 U16526 ( .IN1(n14304), .IN2(n4471), .Q(n15756) );
  OR2X1 U16527 ( .IN1(n15759), .IN2(n15760), .Q(g21073) );
  INVX0 U16528 ( .INP(n15761), .ZN(n15760) );
  OR2X1 U16529 ( .IN1(n14299), .IN2(n8943), .Q(n15761) );
  AND2X1 U16530 ( .IN1(n14299), .IN2(n9122), .Q(n15759) );
  OR2X1 U16531 ( .IN1(n15762), .IN2(n15763), .Q(g21072) );
  INVX0 U16532 ( .INP(n15764), .ZN(n15763) );
  OR2X1 U16533 ( .IN1(n14387), .IN2(n8888), .Q(n15764) );
  AND2X1 U16534 ( .IN1(n14387), .IN2(n9124), .Q(n15762) );
  OR2X1 U16535 ( .IN1(n15765), .IN2(n15766), .Q(g21071) );
  INVX0 U16536 ( .INP(n15767), .ZN(n15766) );
  OR2X1 U16537 ( .IN1(n4149), .IN2(n8951), .Q(n15767) );
  AND2X1 U16538 ( .IN1(n4149), .IN2(n4473), .Q(n15765) );
  OR2X1 U16539 ( .IN1(n15768), .IN2(n15769), .Q(g21070) );
  INVX0 U16540 ( .INP(n15770), .ZN(n15769) );
  OR2X1 U16541 ( .IN1(n14392), .IN2(n8960), .Q(n15770) );
  AND2X1 U16542 ( .IN1(n4395), .IN2(n14392), .Q(n15768) );
  OR2X1 U16543 ( .IN1(n15771), .IN2(n15772), .Q(g21063) );
  INVX0 U16544 ( .INP(n15773), .ZN(n15772) );
  OR2X1 U16545 ( .IN1(n15774), .IN2(n8732), .Q(n15773) );
  AND2X1 U16546 ( .IN1(n15774), .IN2(n9937), .Q(n15771) );
  OR2X1 U16547 ( .IN1(n15775), .IN2(n15776), .Q(g21062) );
  INVX0 U16548 ( .INP(n15777), .ZN(n15776) );
  OR2X1 U16549 ( .IN1(n14312), .IN2(n8872), .Q(n15777) );
  AND2X1 U16550 ( .IN1(n14312), .IN2(n4471), .Q(n15775) );
  OR2X1 U16551 ( .IN1(n15778), .IN2(n15779), .Q(g21061) );
  INVX0 U16552 ( .INP(n15780), .ZN(n15779) );
  OR2X1 U16553 ( .IN1(n14304), .IN2(n8873), .Q(n15780) );
  AND2X1 U16554 ( .IN1(n14304), .IN2(n9122), .Q(n15778) );
  OR2X1 U16555 ( .IN1(n15781), .IN2(n15782), .Q(g21060) );
  INVX0 U16556 ( .INP(n15783), .ZN(n15782) );
  OR2X1 U16557 ( .IN1(n14299), .IN2(n8944), .Q(n15783) );
  AND2X1 U16558 ( .IN1(n14299), .IN2(n4407), .Q(n15781) );
  OR2X1 U16559 ( .IN1(n15784), .IN2(n15785), .Q(g21056) );
  INVX0 U16560 ( .INP(n15786), .ZN(n15785) );
  OR2X1 U16561 ( .IN1(n14396), .IN2(n8889), .Q(n15786) );
  AND2X1 U16562 ( .IN1(n14396), .IN2(n9124), .Q(n15784) );
  OR2X1 U16563 ( .IN1(n15787), .IN2(n15788), .Q(g21055) );
  INVX0 U16564 ( .INP(n15789), .ZN(n15788) );
  OR2X1 U16565 ( .IN1(n14387), .IN2(n8890), .Q(n15789) );
  AND2X1 U16566 ( .IN1(n14387), .IN2(n4473), .Q(n15787) );
  OR2X1 U16567 ( .IN1(n15790), .IN2(n15791), .Q(g21054) );
  INVX0 U16568 ( .INP(n15792), .ZN(n15791) );
  OR2X1 U16569 ( .IN1(n4149), .IN2(n8952), .Q(n15792) );
  AND2X1 U16570 ( .IN1(n4468), .IN2(n4149), .Q(n15790) );
  OR2X1 U16571 ( .IN1(n15793), .IN2(n15794), .Q(g21053) );
  INVX0 U16572 ( .INP(n15795), .ZN(n15794) );
  OR2X1 U16573 ( .IN1(n869), .IN2(n8907), .Q(n15795) );
  AND2X1 U16574 ( .IN1(n4395), .IN2(n869), .Q(n15793) );
  OR2X1 U16575 ( .IN1(n15796), .IN2(n15797), .Q(g21052) );
  INVX0 U16576 ( .INP(n15798), .ZN(n15797) );
  OR2X1 U16577 ( .IN1(n14392), .IN2(n8961), .Q(n15798) );
  AND2X1 U16578 ( .IN1(n14392), .IN2(n4475), .Q(n15796) );
  OR2X1 U16579 ( .IN1(n15799), .IN2(n15800), .Q(g21051) );
  INVX0 U16580 ( .INP(n15801), .ZN(n15800) );
  OR2X1 U16581 ( .IN1(n590), .IN2(n8970), .Q(n15801) );
  AND2X1 U16582 ( .IN1(n4396), .IN2(n590), .Q(n15799) );
  OR2X1 U16583 ( .IN1(n15802), .IN2(n15803), .Q(g21047) );
  INVX0 U16584 ( .INP(n15804), .ZN(n15803) );
  OR2X1 U16585 ( .IN1(n15805), .IN2(n8669), .Q(n15804) );
  AND2X1 U16586 ( .IN1(n15805), .IN2(n9937), .Q(n15802) );
  OR2X1 U16587 ( .IN1(n15806), .IN2(n15807), .Q(g21046) );
  INVX0 U16588 ( .INP(n15808), .ZN(n15807) );
  OR2X1 U16589 ( .IN1(n15774), .IN2(n8733), .Q(n15808) );
  AND2X1 U16590 ( .IN1(n15774), .IN2(n9946), .Q(n15806) );
  INVX0 U16591 ( .INP(n15325), .ZN(n15774) );
  OR2X1 U16592 ( .IN1(n4292), .IN2(n9085), .Q(n15325) );
  OR2X1 U16593 ( .IN1(n15809), .IN2(n15810), .Q(g21045) );
  INVX0 U16594 ( .INP(n15811), .ZN(n15810) );
  OR2X1 U16595 ( .IN1(n14312), .IN2(n8874), .Q(n15811) );
  AND2X1 U16596 ( .IN1(n14312), .IN2(n9122), .Q(n15809) );
  OR2X1 U16597 ( .IN1(n15812), .IN2(n15813), .Q(g21044) );
  INVX0 U16598 ( .INP(n15814), .ZN(n15813) );
  OR2X1 U16599 ( .IN1(n14304), .IN2(n8875), .Q(n15814) );
  AND2X1 U16600 ( .IN1(n14304), .IN2(n4407), .Q(n15812) );
  OR2X1 U16601 ( .IN1(n15815), .IN2(n15816), .Q(g21043) );
  INVX0 U16602 ( .INP(n15817), .ZN(n15816) );
  OR2X1 U16603 ( .IN1(n14299), .IN2(n8945), .Q(n15817) );
  AND2X1 U16604 ( .IN1(n4397), .IN2(n14299), .Q(n15815) );
  OR2X1 U16605 ( .IN1(n15818), .IN2(n15819), .Q(g21042) );
  INVX0 U16606 ( .INP(n15820), .ZN(n15819) );
  OR2X1 U16607 ( .IN1(n15821), .IN2(n8734), .Q(n15820) );
  AND2X1 U16608 ( .IN1(n15821), .IN2(n10071), .Q(n15818) );
  OR2X1 U16609 ( .IN1(n15822), .IN2(n15823), .Q(g21041) );
  INVX0 U16610 ( .INP(n15824), .ZN(n15823) );
  OR2X1 U16611 ( .IN1(n14396), .IN2(n8891), .Q(n15824) );
  AND2X1 U16612 ( .IN1(n14396), .IN2(n4473), .Q(n15822) );
  OR2X1 U16613 ( .IN1(n15825), .IN2(n15826), .Q(g21040) );
  INVX0 U16614 ( .INP(n15827), .ZN(n15826) );
  OR2X1 U16615 ( .IN1(n14387), .IN2(n8892), .Q(n15827) );
  AND2X1 U16616 ( .IN1(n4468), .IN2(n14387), .Q(n15825) );
  OR2X1 U16617 ( .IN1(n15828), .IN2(n15829), .Q(g21039) );
  INVX0 U16618 ( .INP(n15830), .ZN(n15829) );
  OR2X1 U16619 ( .IN1(n4149), .IN2(n8953), .Q(n15830) );
  AND2X1 U16620 ( .IN1(n4149), .IN2(n4409), .Q(n15828) );
  OR2X1 U16621 ( .IN1(n15831), .IN2(n15832), .Q(g21035) );
  INVX0 U16622 ( .INP(n15833), .ZN(n15832) );
  OR2X1 U16623 ( .IN1(n14484), .IN2(n8908), .Q(n15833) );
  AND2X1 U16624 ( .IN1(n4395), .IN2(n14484), .Q(n15831) );
  OR2X1 U16625 ( .IN1(n15834), .IN2(n15835), .Q(g21034) );
  INVX0 U16626 ( .INP(n15836), .ZN(n15835) );
  OR2X1 U16627 ( .IN1(n869), .IN2(n8909), .Q(n15836) );
  AND2X1 U16628 ( .IN1(n869), .IN2(n4475), .Q(n15834) );
  OR2X1 U16629 ( .IN1(n15837), .IN2(n15838), .Q(g21033) );
  INVX0 U16630 ( .INP(n15839), .ZN(n15838) );
  OR2X1 U16631 ( .IN1(n14392), .IN2(n8962), .Q(n15839) );
  AND2X1 U16632 ( .IN1(n4469), .IN2(n14392), .Q(n15837) );
  OR2X1 U16633 ( .IN1(n15840), .IN2(n15841), .Q(g21032) );
  INVX0 U16634 ( .INP(n15842), .ZN(n15841) );
  OR2X1 U16635 ( .IN1(n14561), .IN2(n8924), .Q(n15842) );
  AND2X1 U16636 ( .IN1(n4396), .IN2(n14561), .Q(n15840) );
  OR2X1 U16637 ( .IN1(n15843), .IN2(n15844), .Q(g21031) );
  INVX0 U16638 ( .INP(n15845), .ZN(n15844) );
  OR2X1 U16639 ( .IN1(n590), .IN2(n8971), .Q(n15845) );
  AND2X1 U16640 ( .IN1(n590), .IN2(n4477), .Q(n15843) );
  OR2X1 U16641 ( .IN1(n15846), .IN2(n15847), .Q(g21029) );
  INVX0 U16642 ( .INP(n15848), .ZN(n15847) );
  OR2X1 U16643 ( .IN1(n15849), .IN2(n8677), .Q(n15848) );
  AND2X1 U16644 ( .IN1(n15849), .IN2(n9937), .Q(n15846) );
  INVX0 U16645 ( .INP(n9879), .ZN(n9937) );
  OR2X1 U16646 ( .IN1(n15850), .IN2(n15851), .Q(n9879) );
  OR2X1 U16647 ( .IN1(n15852), .IN2(n15853), .Q(n15851) );
  AND2X1 U16648 ( .IN1(g2624), .IN2(g2685), .Q(n15853) );
  AND2X1 U16649 ( .IN1(g7302), .IN2(g2679), .Q(n15852) );
  AND2X1 U16650 ( .IN1(test_so90), .IN2(g7390), .Q(n15850) );
  OR2X1 U16651 ( .IN1(n15854), .IN2(n15855), .Q(g21028) );
  INVX0 U16652 ( .INP(n15856), .ZN(n15855) );
  OR2X1 U16653 ( .IN1(n15805), .IN2(n8670), .Q(n15856) );
  AND2X1 U16654 ( .IN1(n15805), .IN2(n9946), .Q(n15854) );
  INVX0 U16655 ( .INP(n12737), .ZN(n15805) );
  OR2X1 U16656 ( .IN1(n15857), .IN2(n15858), .Q(g21027) );
  INVX0 U16657 ( .INP(n15859), .ZN(n15858) );
  OR2X1 U16658 ( .IN1(n14312), .IN2(n8876), .Q(n15859) );
  AND2X1 U16659 ( .IN1(n14312), .IN2(n4407), .Q(n15857) );
  OR2X1 U16660 ( .IN1(n15860), .IN2(n15861), .Q(g21026) );
  INVX0 U16661 ( .INP(n15862), .ZN(n15861) );
  OR2X1 U16662 ( .IN1(n14304), .IN2(n8877), .Q(n15862) );
  AND2X1 U16663 ( .IN1(n4397), .IN2(n14304), .Q(n15860) );
  OR2X1 U16664 ( .IN1(n15863), .IN2(n15864), .Q(g21025) );
  AND2X1 U16665 ( .IN1(n14299), .IN2(n4408), .Q(n15864) );
  AND2X1 U16666 ( .IN1(test_so93), .IN2(n14300), .Q(n15863) );
  OR2X1 U16667 ( .IN1(n15865), .IN2(n15866), .Q(g21023) );
  INVX0 U16668 ( .INP(n15867), .ZN(n15866) );
  OR2X1 U16669 ( .IN1(n15868), .IN2(n8671), .Q(n15867) );
  AND2X1 U16670 ( .IN1(n15868), .IN2(n10071), .Q(n15865) );
  OR2X1 U16671 ( .IN1(n15869), .IN2(n15870), .Q(g21022) );
  INVX0 U16672 ( .INP(n15871), .ZN(n15870) );
  OR2X1 U16673 ( .IN1(n15821), .IN2(n8735), .Q(n15871) );
  AND2X1 U16674 ( .IN1(n15821), .IN2(n10079), .Q(n15869) );
  INVX0 U16675 ( .INP(n15328), .ZN(n15821) );
  OR2X1 U16676 ( .IN1(n4293), .IN2(n9084), .Q(n15328) );
  OR2X1 U16677 ( .IN1(n15872), .IN2(n15873), .Q(g21021) );
  INVX0 U16678 ( .INP(n15874), .ZN(n15873) );
  OR2X1 U16679 ( .IN1(n14396), .IN2(n8893), .Q(n15874) );
  AND2X1 U16680 ( .IN1(n4468), .IN2(n14396), .Q(n15872) );
  OR2X1 U16681 ( .IN1(n15875), .IN2(n15876), .Q(g21020) );
  INVX0 U16682 ( .INP(n15877), .ZN(n15876) );
  OR2X1 U16683 ( .IN1(n14387), .IN2(n8894), .Q(n15877) );
  AND2X1 U16684 ( .IN1(n14387), .IN2(n4409), .Q(n15875) );
  OR2X1 U16685 ( .IN1(n15878), .IN2(n15879), .Q(g21019) );
  INVX0 U16686 ( .INP(n15880), .ZN(n15879) );
  OR2X1 U16687 ( .IN1(n4149), .IN2(n8954), .Q(n15880) );
  AND2X1 U16688 ( .IN1(n4399), .IN2(n4149), .Q(n15878) );
  OR2X1 U16689 ( .IN1(n15881), .IN2(n15882), .Q(g21018) );
  INVX0 U16690 ( .INP(n15883), .ZN(n15882) );
  OR2X1 U16691 ( .IN1(n15884), .IN2(n8736), .Q(n15883) );
  AND2X1 U16692 ( .IN1(n15884), .IN2(n10206), .Q(n15881) );
  OR2X1 U16693 ( .IN1(n15885), .IN2(n15886), .Q(g21017) );
  INVX0 U16694 ( .INP(n15887), .ZN(n15886) );
  OR2X1 U16695 ( .IN1(n14484), .IN2(n8910), .Q(n15887) );
  AND2X1 U16696 ( .IN1(n14484), .IN2(n4475), .Q(n15885) );
  OR2X1 U16697 ( .IN1(n15888), .IN2(n15889), .Q(g21016) );
  INVX0 U16698 ( .INP(n15890), .ZN(n15889) );
  OR2X1 U16699 ( .IN1(n869), .IN2(n8911), .Q(n15890) );
  AND2X1 U16700 ( .IN1(n4469), .IN2(n869), .Q(n15888) );
  OR2X1 U16701 ( .IN1(n15891), .IN2(n15892), .Q(g21015) );
  INVX0 U16702 ( .INP(n15893), .ZN(n15892) );
  OR2X1 U16703 ( .IN1(n14392), .IN2(n8963), .Q(n15893) );
  AND2X1 U16704 ( .IN1(n14392), .IN2(n4411), .Q(n15891) );
  OR2X1 U16705 ( .IN1(n15894), .IN2(n15895), .Q(g21011) );
  INVX0 U16706 ( .INP(n15896), .ZN(n15895) );
  OR2X1 U16707 ( .IN1(n14565), .IN2(n8925), .Q(n15896) );
  AND2X1 U16708 ( .IN1(n4396), .IN2(n14565), .Q(n15894) );
  OR2X1 U16709 ( .IN1(n15897), .IN2(n15898), .Q(g21010) );
  INVX0 U16710 ( .INP(n15899), .ZN(n15898) );
  OR2X1 U16711 ( .IN1(n14561), .IN2(n8926), .Q(n15899) );
  AND2X1 U16712 ( .IN1(n14561), .IN2(n4477), .Q(n15897) );
  OR2X1 U16713 ( .IN1(n15900), .IN2(n15901), .Q(g21009) );
  INVX0 U16714 ( .INP(n15902), .ZN(n15901) );
  OR2X1 U16715 ( .IN1(n590), .IN2(n8972), .Q(n15902) );
  AND2X1 U16716 ( .IN1(n590), .IN2(n9123), .Q(n15900) );
  OR2X1 U16717 ( .IN1(n15903), .IN2(n15904), .Q(g21007) );
  INVX0 U16718 ( .INP(n15905), .ZN(n15904) );
  OR2X1 U16719 ( .IN1(n15849), .IN2(n8678), .Q(n15905) );
  AND2X1 U16720 ( .IN1(n15849), .IN2(n9946), .Q(n15903) );
  INVX0 U16721 ( .INP(n9889), .ZN(n9946) );
  OR2X1 U16722 ( .IN1(n15906), .IN2(n15907), .Q(n9889) );
  OR2X1 U16723 ( .IN1(n15908), .IN2(n15909), .Q(n15907) );
  AND2X1 U16724 ( .IN1(n11411), .IN2(g2688), .Q(n15909) );
  INVX0 U16725 ( .INP(n4314), .ZN(n11411) );
  AND2X1 U16726 ( .IN1(g2624), .IN2(g2694), .Q(n15908) );
  AND2X1 U16727 ( .IN1(g7390), .IN2(g2691), .Q(n15906) );
  INVX0 U16728 ( .INP(n15330), .ZN(n15849) );
  OR2X1 U16729 ( .IN1(n4306), .IN2(n9085), .Q(n15330) );
  OR2X1 U16730 ( .IN1(n15910), .IN2(n15911), .Q(g21006) );
  INVX0 U16731 ( .INP(n15912), .ZN(n15911) );
  OR2X1 U16732 ( .IN1(n14312), .IN2(n8878), .Q(n15912) );
  AND2X1 U16733 ( .IN1(n4397), .IN2(n14312), .Q(n15910) );
  OR2X1 U16734 ( .IN1(n15913), .IN2(n15914), .Q(g21005) );
  INVX0 U16735 ( .INP(n15915), .ZN(n15914) );
  OR2X1 U16736 ( .IN1(n14304), .IN2(n8879), .Q(n15915) );
  AND2X1 U16737 ( .IN1(n14304), .IN2(n4408), .Q(n15913) );
  OR2X1 U16738 ( .IN1(n15916), .IN2(n15917), .Q(g21004) );
  INVX0 U16739 ( .INP(n15918), .ZN(n15917) );
  OR2X1 U16740 ( .IN1(n14299), .IN2(n8946), .Q(n15918) );
  AND2X1 U16741 ( .IN1(n4419), .IN2(n14299), .Q(n15916) );
  OR2X1 U16742 ( .IN1(n15919), .IN2(n15920), .Q(g21003) );
  INVX0 U16743 ( .INP(n15921), .ZN(n15920) );
  OR2X1 U16744 ( .IN1(n15922), .IN2(n8679), .Q(n15921) );
  AND2X1 U16745 ( .IN1(n15922), .IN2(n10071), .Q(n15919) );
  INVX0 U16746 ( .INP(n10013), .ZN(n10071) );
  OR2X1 U16747 ( .IN1(n15923), .IN2(n15924), .Q(n10013) );
  OR2X1 U16748 ( .IN1(n15925), .IN2(n15926), .Q(n15924) );
  AND2X1 U16749 ( .IN1(g7194), .IN2(g1988), .Q(n15926) );
  AND2X1 U16750 ( .IN1(g7052), .IN2(g1985), .Q(n15925) );
  AND2X1 U16751 ( .IN1(g1930), .IN2(g1991), .Q(n15923) );
  OR2X1 U16752 ( .IN1(n15927), .IN2(n15928), .Q(g21002) );
  INVX0 U16753 ( .INP(n15929), .ZN(n15928) );
  OR2X1 U16754 ( .IN1(n15868), .IN2(n8672), .Q(n15929) );
  AND2X1 U16755 ( .IN1(n15868), .IN2(n10079), .Q(n15927) );
  INVX0 U16756 ( .INP(n12741), .ZN(n15868) );
  OR2X1 U16757 ( .IN1(n15930), .IN2(n15931), .Q(g21001) );
  INVX0 U16758 ( .INP(n15932), .ZN(n15931) );
  OR2X1 U16759 ( .IN1(n14396), .IN2(n8895), .Q(n15932) );
  AND2X1 U16760 ( .IN1(n14396), .IN2(n4409), .Q(n15930) );
  OR2X1 U16761 ( .IN1(n15933), .IN2(n15934), .Q(g21000) );
  AND2X1 U16762 ( .IN1(n4399), .IN2(n14387), .Q(n15934) );
  AND2X1 U16763 ( .IN1(test_so71), .IN2(n14388), .Q(n15933) );
  OR2X1 U16764 ( .IN1(n15935), .IN2(n15936), .Q(g20999) );
  INVX0 U16765 ( .INP(n15937), .ZN(n15936) );
  OR2X1 U16766 ( .IN1(n4149), .IN2(n8955), .Q(n15937) );
  AND2X1 U16767 ( .IN1(n4149), .IN2(n4410), .Q(n15935) );
  OR2X1 U16768 ( .IN1(n15938), .IN2(n15939), .Q(g20997) );
  INVX0 U16769 ( .INP(n15940), .ZN(n15939) );
  OR2X1 U16770 ( .IN1(n15941), .IN2(n8673), .Q(n15940) );
  AND2X1 U16771 ( .IN1(n15941), .IN2(n10206), .Q(n15938) );
  OR2X1 U16772 ( .IN1(n15942), .IN2(n15943), .Q(g20996) );
  AND2X1 U16773 ( .IN1(n15884), .IN2(n10214), .Q(n15943) );
  INVX0 U16774 ( .INP(n15333), .ZN(n15884) );
  AND2X1 U16775 ( .IN1(test_so51), .IN2(n15333), .Q(n15942) );
  OR2X1 U16776 ( .IN1(n4294), .IN2(n9083), .Q(n15333) );
  OR2X1 U16777 ( .IN1(n15944), .IN2(n15945), .Q(g20995) );
  INVX0 U16778 ( .INP(n15946), .ZN(n15945) );
  OR2X1 U16779 ( .IN1(n14484), .IN2(n8912), .Q(n15946) );
  AND2X1 U16780 ( .IN1(n4469), .IN2(n14484), .Q(n15944) );
  OR2X1 U16781 ( .IN1(n15947), .IN2(n15948), .Q(g20994) );
  AND2X1 U16782 ( .IN1(n869), .IN2(n4411), .Q(n15948) );
  AND2X1 U16783 ( .IN1(test_so50), .IN2(n14472), .Q(n15947) );
  OR2X1 U16784 ( .IN1(n15949), .IN2(n15950), .Q(g20993) );
  INVX0 U16785 ( .INP(n15951), .ZN(n15950) );
  OR2X1 U16786 ( .IN1(n14392), .IN2(n8964), .Q(n15951) );
  AND2X1 U16787 ( .IN1(n4401), .IN2(n14392), .Q(n15949) );
  OR2X1 U16788 ( .IN1(n15952), .IN2(n15953), .Q(g20992) );
  INVX0 U16789 ( .INP(n15954), .ZN(n15953) );
  OR2X1 U16790 ( .IN1(n15955), .IN2(n8737), .Q(n15954) );
  AND2X1 U16791 ( .IN1(n15955), .IN2(n9805), .Q(n15952) );
  OR2X1 U16792 ( .IN1(n15956), .IN2(n15957), .Q(g20991) );
  INVX0 U16793 ( .INP(n15958), .ZN(n15957) );
  OR2X1 U16794 ( .IN1(n14565), .IN2(n8927), .Q(n15958) );
  AND2X1 U16795 ( .IN1(n14565), .IN2(n4477), .Q(n15956) );
  OR2X1 U16796 ( .IN1(n15959), .IN2(n15960), .Q(g20990) );
  INVX0 U16797 ( .INP(n15961), .ZN(n15960) );
  OR2X1 U16798 ( .IN1(n14561), .IN2(n8928), .Q(n15961) );
  AND2X1 U16799 ( .IN1(n14561), .IN2(n9123), .Q(n15959) );
  OR2X1 U16800 ( .IN1(n15962), .IN2(n15963), .Q(g20989) );
  INVX0 U16801 ( .INP(n15964), .ZN(n15963) );
  OR2X1 U16802 ( .IN1(n590), .IN2(n8973), .Q(n15964) );
  AND2X1 U16803 ( .IN1(n590), .IN2(n4413), .Q(n15962) );
  OR2X1 U16804 ( .IN1(n15965), .IN2(n15966), .Q(g20983) );
  INVX0 U16805 ( .INP(n15967), .ZN(n15966) );
  OR2X1 U16806 ( .IN1(n14312), .IN2(n8880), .Q(n15967) );
  AND2X1 U16807 ( .IN1(n14312), .IN2(n4408), .Q(n15965) );
  OR2X1 U16808 ( .IN1(n15968), .IN2(n15969), .Q(g20982) );
  INVX0 U16809 ( .INP(n15970), .ZN(n15969) );
  OR2X1 U16810 ( .IN1(n14304), .IN2(n8881), .Q(n15970) );
  AND2X1 U16811 ( .IN1(n4419), .IN2(n14304), .Q(n15968) );
  OR2X1 U16812 ( .IN1(n15971), .IN2(n15972), .Q(g20981) );
  INVX0 U16813 ( .INP(n15973), .ZN(n15972) );
  OR2X1 U16814 ( .IN1(n14299), .IN2(n8947), .Q(n15973) );
  AND2X1 U16815 ( .IN1(n14299), .IN2(n4472), .Q(n15971) );
  OR2X1 U16816 ( .IN1(n15974), .IN2(n15975), .Q(g20980) );
  INVX0 U16817 ( .INP(n15976), .ZN(n15975) );
  OR2X1 U16818 ( .IN1(n15922), .IN2(n8680), .Q(n15976) );
  AND2X1 U16819 ( .IN1(n15922), .IN2(n10079), .Q(n15974) );
  INVX0 U16820 ( .INP(n10023), .ZN(n10079) );
  OR2X1 U16821 ( .IN1(n15977), .IN2(n15978), .Q(n10023) );
  OR2X1 U16822 ( .IN1(n15979), .IN2(n15980), .Q(n15978) );
  AND2X1 U16823 ( .IN1(g7194), .IN2(g1997), .Q(n15980) );
  AND2X1 U16824 ( .IN1(n12379), .IN2(g1994), .Q(n15979) );
  INVX0 U16825 ( .INP(n4296), .ZN(n12379) );
  AND2X1 U16826 ( .IN1(g1930), .IN2(g2000), .Q(n15977) );
  INVX0 U16827 ( .INP(n15335), .ZN(n15922) );
  OR2X1 U16828 ( .IN1(n4307), .IN2(n9084), .Q(n15335) );
  OR2X1 U16829 ( .IN1(n15981), .IN2(n15982), .Q(g20979) );
  INVX0 U16830 ( .INP(n15983), .ZN(n15982) );
  OR2X1 U16831 ( .IN1(n14396), .IN2(n8896), .Q(n15983) );
  AND2X1 U16832 ( .IN1(n4399), .IN2(n14396), .Q(n15981) );
  OR2X1 U16833 ( .IN1(n15984), .IN2(n15985), .Q(g20978) );
  INVX0 U16834 ( .INP(n15986), .ZN(n15985) );
  OR2X1 U16835 ( .IN1(n14387), .IN2(n8897), .Q(n15986) );
  AND2X1 U16836 ( .IN1(n14387), .IN2(n4410), .Q(n15984) );
  OR2X1 U16837 ( .IN1(n15987), .IN2(n15988), .Q(g20977) );
  INVX0 U16838 ( .INP(n15989), .ZN(n15988) );
  OR2X1 U16839 ( .IN1(n4149), .IN2(n8956), .Q(n15989) );
  AND2X1 U16840 ( .IN1(n4420), .IN2(n4149), .Q(n15987) );
  OR2X1 U16841 ( .IN1(n15990), .IN2(n15991), .Q(g20976) );
  INVX0 U16842 ( .INP(n15992), .ZN(n15991) );
  OR2X1 U16843 ( .IN1(n15993), .IN2(n8681), .Q(n15992) );
  AND2X1 U16844 ( .IN1(n15993), .IN2(n10206), .Q(n15990) );
  INVX0 U16845 ( .INP(n10148), .ZN(n10206) );
  OR2X1 U16846 ( .IN1(n15994), .IN2(n15995), .Q(n10148) );
  OR2X1 U16847 ( .IN1(n15996), .IN2(n15997), .Q(n15995) );
  AND2X1 U16848 ( .IN1(g1236), .IN2(g1297), .Q(n15997) );
  AND2X1 U16849 ( .IN1(g6750), .IN2(g1291), .Q(n15996) );
  AND2X1 U16850 ( .IN1(g6944), .IN2(g1294), .Q(n15994) );
  OR2X1 U16851 ( .IN1(n15998), .IN2(n15999), .Q(g20975) );
  INVX0 U16852 ( .INP(n16000), .ZN(n15999) );
  OR2X1 U16853 ( .IN1(n15941), .IN2(n8674), .Q(n16000) );
  AND2X1 U16854 ( .IN1(n15941), .IN2(n10214), .Q(n15998) );
  INVX0 U16855 ( .INP(n12745), .ZN(n15941) );
  OR2X1 U16856 ( .IN1(n16001), .IN2(n16002), .Q(g20974) );
  INVX0 U16857 ( .INP(n16003), .ZN(n16002) );
  OR2X1 U16858 ( .IN1(n14484), .IN2(n8913), .Q(n16003) );
  AND2X1 U16859 ( .IN1(n14484), .IN2(n4411), .Q(n16001) );
  OR2X1 U16860 ( .IN1(n16004), .IN2(n16005), .Q(g20973) );
  INVX0 U16861 ( .INP(n16006), .ZN(n16005) );
  OR2X1 U16862 ( .IN1(n869), .IN2(n8914), .Q(n16006) );
  AND2X1 U16863 ( .IN1(n4401), .IN2(n869), .Q(n16004) );
  OR2X1 U16864 ( .IN1(n16007), .IN2(n16008), .Q(g20972) );
  INVX0 U16865 ( .INP(n16009), .ZN(n16008) );
  OR2X1 U16866 ( .IN1(n14392), .IN2(n8965), .Q(n16009) );
  AND2X1 U16867 ( .IN1(n14392), .IN2(n4412), .Q(n16007) );
  OR2X1 U16868 ( .IN1(n16010), .IN2(n16011), .Q(g20970) );
  INVX0 U16869 ( .INP(n16012), .ZN(n16011) );
  OR2X1 U16870 ( .IN1(n16013), .IN2(n8675), .Q(n16012) );
  AND2X1 U16871 ( .IN1(n16013), .IN2(n9805), .Q(n16010) );
  OR2X1 U16872 ( .IN1(n16014), .IN2(n16015), .Q(g20969) );
  INVX0 U16873 ( .INP(n16016), .ZN(n16015) );
  OR2X1 U16874 ( .IN1(n15955), .IN2(n8738), .Q(n16016) );
  AND2X1 U16875 ( .IN1(n15955), .IN2(n9798), .Q(n16014) );
  INVX0 U16876 ( .INP(n15338), .ZN(n15955) );
  OR2X1 U16877 ( .IN1(n4295), .IN2(n9082), .Q(n15338) );
  OR2X1 U16878 ( .IN1(n16017), .IN2(n16018), .Q(g20968) );
  INVX0 U16879 ( .INP(n16019), .ZN(n16018) );
  OR2X1 U16880 ( .IN1(n14565), .IN2(n8929), .Q(n16019) );
  AND2X1 U16881 ( .IN1(n14565), .IN2(n9123), .Q(n16017) );
  OR2X1 U16882 ( .IN1(n16020), .IN2(n16021), .Q(g20967) );
  INVX0 U16883 ( .INP(n16022), .ZN(n16021) );
  OR2X1 U16884 ( .IN1(n14561), .IN2(n8930), .Q(n16022) );
  AND2X1 U16885 ( .IN1(n14561), .IN2(n4413), .Q(n16020) );
  OR2X1 U16886 ( .IN1(n16023), .IN2(n16024), .Q(g20966) );
  INVX0 U16887 ( .INP(n16025), .ZN(n16024) );
  OR2X1 U16888 ( .IN1(n590), .IN2(n8974), .Q(n16025) );
  AND2X1 U16889 ( .IN1(n4403), .IN2(n590), .Q(n16023) );
  OR2X1 U16890 ( .IN1(n16026), .IN2(n16027), .Q(g20965) );
  INVX0 U16891 ( .INP(n16028), .ZN(n16027) );
  OR2X1 U16892 ( .IN1(n14299), .IN2(n8941), .Q(n16028) );
  AND2X1 U16893 ( .IN1(n4415), .IN2(n14299), .Q(n16026) );
  OR2X1 U16894 ( .IN1(n16029), .IN2(n16030), .Q(g20964) );
  INVX0 U16895 ( .INP(n16031), .ZN(n16030) );
  OR2X1 U16896 ( .IN1(n14312), .IN2(n8882), .Q(n16031) );
  AND2X1 U16897 ( .IN1(n4419), .IN2(n14312), .Q(n16029) );
  OR2X1 U16898 ( .IN1(n16032), .IN2(n16033), .Q(g20963) );
  INVX0 U16899 ( .INP(n16034), .ZN(n16033) );
  OR2X1 U16900 ( .IN1(n14304), .IN2(n8883), .Q(n16034) );
  AND2X1 U16901 ( .IN1(n14304), .IN2(n4472), .Q(n16032) );
  OR2X1 U16902 ( .IN1(n16035), .IN2(n16036), .Q(g20962) );
  INVX0 U16903 ( .INP(n16037), .ZN(n16036) );
  OR2X1 U16904 ( .IN1(n14299), .IN2(n8948), .Q(n16037) );
  AND2X1 U16905 ( .IN1(n4398), .IN2(n14299), .Q(n16035) );
  INVX0 U16906 ( .INP(n14300), .ZN(n14299) );
  OR2X1 U16907 ( .IN1(n15683), .IN2(n16038), .Q(n14300) );
  OR2X1 U16908 ( .IN1(n16039), .IN2(n16040), .Q(g20955) );
  INVX0 U16909 ( .INP(n16041), .ZN(n16040) );
  OR2X1 U16910 ( .IN1(n14396), .IN2(n8898), .Q(n16041) );
  AND2X1 U16911 ( .IN1(n14396), .IN2(n4410), .Q(n16039) );
  OR2X1 U16912 ( .IN1(n16042), .IN2(n16043), .Q(g20954) );
  INVX0 U16913 ( .INP(n16044), .ZN(n16043) );
  OR2X1 U16914 ( .IN1(n14387), .IN2(n8899), .Q(n16044) );
  AND2X1 U16915 ( .IN1(n4420), .IN2(n14387), .Q(n16042) );
  OR2X1 U16916 ( .IN1(n16045), .IN2(n16046), .Q(g20953) );
  INVX0 U16917 ( .INP(n16047), .ZN(n16046) );
  OR2X1 U16918 ( .IN1(n4149), .IN2(n8957), .Q(n16047) );
  AND2X1 U16919 ( .IN1(n4149), .IN2(n4474), .Q(n16045) );
  OR2X1 U16920 ( .IN1(n16048), .IN2(n16049), .Q(g20952) );
  INVX0 U16921 ( .INP(n16050), .ZN(n16049) );
  OR2X1 U16922 ( .IN1(n15993), .IN2(n8682), .Q(n16050) );
  AND2X1 U16923 ( .IN1(n15993), .IN2(n10214), .Q(n16048) );
  INVX0 U16924 ( .INP(n10158), .ZN(n10214) );
  OR2X1 U16925 ( .IN1(n16051), .IN2(n16052), .Q(n10158) );
  OR2X1 U16926 ( .IN1(n16053), .IN2(n16054), .Q(n16052) );
  AND2X1 U16927 ( .IN1(g6944), .IN2(g1303), .Q(n16054) );
  AND2X1 U16928 ( .IN1(g1236), .IN2(g1306), .Q(n16053) );
  AND2X1 U16929 ( .IN1(n12249), .IN2(g1300), .Q(n16051) );
  INVX0 U16930 ( .INP(n4371), .ZN(n12249) );
  INVX0 U16931 ( .INP(n15340), .ZN(n15993) );
  OR2X1 U16932 ( .IN1(n4308), .IN2(n9083), .Q(n15340) );
  OR2X1 U16933 ( .IN1(n16055), .IN2(n16056), .Q(g20951) );
  INVX0 U16934 ( .INP(n16057), .ZN(n16056) );
  OR2X1 U16935 ( .IN1(n14484), .IN2(n8915), .Q(n16057) );
  AND2X1 U16936 ( .IN1(n4401), .IN2(n14484), .Q(n16055) );
  OR2X1 U16937 ( .IN1(n16058), .IN2(n16059), .Q(g20950) );
  INVX0 U16938 ( .INP(n16060), .ZN(n16059) );
  OR2X1 U16939 ( .IN1(n869), .IN2(n8916), .Q(n16060) );
  AND2X1 U16940 ( .IN1(n869), .IN2(n4412), .Q(n16058) );
  OR2X1 U16941 ( .IN1(n16061), .IN2(n16062), .Q(g20949) );
  INVX0 U16942 ( .INP(n16063), .ZN(n16062) );
  OR2X1 U16943 ( .IN1(n14392), .IN2(n8966), .Q(n16063) );
  AND2X1 U16944 ( .IN1(n4421), .IN2(n14392), .Q(n16061) );
  OR2X1 U16945 ( .IN1(n16064), .IN2(n16065), .Q(g20948) );
  INVX0 U16946 ( .INP(n16066), .ZN(n16065) );
  OR2X1 U16947 ( .IN1(n16067), .IN2(n8683), .Q(n16066) );
  AND2X1 U16948 ( .IN1(n16067), .IN2(n9805), .Q(n16064) );
  INVX0 U16949 ( .INP(n9744), .ZN(n9805) );
  OR2X1 U16950 ( .IN1(n16068), .IN2(n16069), .Q(n9744) );
  OR2X1 U16951 ( .IN1(n16070), .IN2(n16071), .Q(n16069) );
  AND2X1 U16952 ( .IN1(g550), .IN2(g611), .Q(n16071) );
  AND2X1 U16953 ( .IN1(n9810), .IN2(g605), .Q(n16070) );
  INVX0 U16954 ( .INP(n4298), .ZN(n9810) );
  AND2X1 U16955 ( .IN1(g6642), .IN2(g608), .Q(n16068) );
  OR2X1 U16956 ( .IN1(n16072), .IN2(n16073), .Q(g20947) );
  INVX0 U16957 ( .INP(n16074), .ZN(n16073) );
  OR2X1 U16958 ( .IN1(n16013), .IN2(n8676), .Q(n16074) );
  AND2X1 U16959 ( .IN1(n16013), .IN2(n9798), .Q(n16072) );
  INVX0 U16960 ( .INP(n12226), .ZN(n16013) );
  OR2X1 U16961 ( .IN1(n16075), .IN2(n16076), .Q(g20946) );
  INVX0 U16962 ( .INP(n16077), .ZN(n16076) );
  OR2X1 U16963 ( .IN1(n14565), .IN2(n8931), .Q(n16077) );
  AND2X1 U16964 ( .IN1(n14565), .IN2(n4413), .Q(n16075) );
  OR2X1 U16965 ( .IN1(n16078), .IN2(n16079), .Q(g20945) );
  INVX0 U16966 ( .INP(n16080), .ZN(n16079) );
  OR2X1 U16967 ( .IN1(n14561), .IN2(n8932), .Q(n16080) );
  AND2X1 U16968 ( .IN1(n4403), .IN2(n14561), .Q(n16078) );
  OR2X1 U16969 ( .IN1(n16081), .IN2(n16082), .Q(g20944) );
  INVX0 U16970 ( .INP(n16083), .ZN(n16082) );
  OR2X1 U16971 ( .IN1(n590), .IN2(n8975), .Q(n16083) );
  AND2X1 U16972 ( .IN1(n590), .IN2(n4414), .Q(n16081) );
  OR2X1 U16973 ( .IN1(n16084), .IN2(n16085), .Q(g20941) );
  INVX0 U16974 ( .INP(n16086), .ZN(n16085) );
  OR2X1 U16975 ( .IN1(n14304), .IN2(n8867), .Q(n16086) );
  AND2X1 U16976 ( .IN1(n4415), .IN2(n14304), .Q(n16084) );
  OR2X1 U16977 ( .IN1(n16087), .IN2(n16088), .Q(g20940) );
  INVX0 U16978 ( .INP(n16089), .ZN(n16088) );
  OR2X1 U16979 ( .IN1(n14312), .IN2(n8884), .Q(n16089) );
  AND2X1 U16980 ( .IN1(n14312), .IN2(n4472), .Q(n16087) );
  OR2X1 U16981 ( .IN1(n16090), .IN2(n16091), .Q(g20939) );
  INVX0 U16982 ( .INP(n16092), .ZN(n16091) );
  OR2X1 U16983 ( .IN1(n14304), .IN2(n8885), .Q(n16092) );
  AND2X1 U16984 ( .IN1(n4398), .IN2(n14304), .Q(n16090) );
  INVX0 U16985 ( .INP(n14303), .ZN(n14304) );
  OR2X1 U16986 ( .IN1(n4356), .IN2(n16093), .Q(n14303) );
  OR2X1 U16987 ( .IN1(n16094), .IN2(n16095), .Q(g20937) );
  INVX0 U16988 ( .INP(n16096), .ZN(n16095) );
  OR2X1 U16989 ( .IN1(n4149), .IN2(n8949), .Q(n16096) );
  AND2X1 U16990 ( .IN1(n4416), .IN2(n4149), .Q(n16094) );
  OR2X1 U16991 ( .IN1(n16097), .IN2(n16098), .Q(g20936) );
  INVX0 U16992 ( .INP(n16099), .ZN(n16098) );
  OR2X1 U16993 ( .IN1(n14396), .IN2(n8900), .Q(n16099) );
  AND2X1 U16994 ( .IN1(n4420), .IN2(n14396), .Q(n16097) );
  OR2X1 U16995 ( .IN1(n16100), .IN2(n16101), .Q(g20935) );
  INVX0 U16996 ( .INP(n16102), .ZN(n16101) );
  OR2X1 U16997 ( .IN1(n14387), .IN2(n8901), .Q(n16102) );
  AND2X1 U16998 ( .IN1(n14387), .IN2(n4474), .Q(n16100) );
  OR2X1 U16999 ( .IN1(n16103), .IN2(n16104), .Q(g20934) );
  INVX0 U17000 ( .INP(n16105), .ZN(n16104) );
  OR2X1 U17001 ( .IN1(n4149), .IN2(n8958), .Q(n16105) );
  AND2X1 U17002 ( .IN1(n4400), .IN2(n4149), .Q(n16103) );
  INVX0 U17003 ( .INP(n14308), .ZN(n4149) );
  OR2X1 U17004 ( .IN1(n15689), .IN2(n16106), .Q(n14308) );
  OR2X1 U17005 ( .IN1(n16107), .IN2(n16108), .Q(g20927) );
  INVX0 U17006 ( .INP(n16109), .ZN(n16108) );
  OR2X1 U17007 ( .IN1(n14484), .IN2(n8917), .Q(n16109) );
  AND2X1 U17008 ( .IN1(n14484), .IN2(n4412), .Q(n16107) );
  OR2X1 U17009 ( .IN1(n16110), .IN2(n16111), .Q(g20926) );
  INVX0 U17010 ( .INP(n16112), .ZN(n16111) );
  OR2X1 U17011 ( .IN1(n869), .IN2(n8918), .Q(n16112) );
  AND2X1 U17012 ( .IN1(n4421), .IN2(n869), .Q(n16110) );
  OR2X1 U17013 ( .IN1(n16113), .IN2(n16114), .Q(g20925) );
  INVX0 U17014 ( .INP(n16115), .ZN(n16114) );
  OR2X1 U17015 ( .IN1(n14392), .IN2(n8967), .Q(n16115) );
  AND2X1 U17016 ( .IN1(n14392), .IN2(n4476), .Q(n16113) );
  OR2X1 U17017 ( .IN1(n16116), .IN2(n16117), .Q(g20924) );
  INVX0 U17018 ( .INP(n16118), .ZN(n16117) );
  OR2X1 U17019 ( .IN1(n16067), .IN2(n8684), .Q(n16118) );
  AND2X1 U17020 ( .IN1(n16067), .IN2(n9798), .Q(n16116) );
  INVX0 U17021 ( .INP(n9738), .ZN(n9798) );
  OR2X1 U17022 ( .IN1(n16119), .IN2(n16120), .Q(n9738) );
  OR2X1 U17023 ( .IN1(n16121), .IN2(n16122), .Q(n16120) );
  AND2X1 U17024 ( .IN1(test_so26), .IN2(g550), .Q(n16122) );
  AND2X1 U17025 ( .IN1(g6485), .IN2(g614), .Q(n16121) );
  AND2X1 U17026 ( .IN1(g6642), .IN2(g617), .Q(n16119) );
  INVX0 U17027 ( .INP(n15343), .ZN(n16067) );
  OR2X1 U17028 ( .IN1(n4309), .IN2(n9082), .Q(n15343) );
  OR2X1 U17029 ( .IN1(n16123), .IN2(n16124), .Q(g20923) );
  AND2X1 U17030 ( .IN1(n4403), .IN2(n14565), .Q(n16124) );
  AND2X1 U17031 ( .IN1(test_so29), .IN2(n14564), .Q(n16123) );
  OR2X1 U17032 ( .IN1(n16125), .IN2(n16126), .Q(g20922) );
  INVX0 U17033 ( .INP(n16127), .ZN(n16126) );
  OR2X1 U17034 ( .IN1(n14561), .IN2(n8933), .Q(n16127) );
  AND2X1 U17035 ( .IN1(n14561), .IN2(n4414), .Q(n16125) );
  OR2X1 U17036 ( .IN1(n16128), .IN2(n16129), .Q(g20921) );
  INVX0 U17037 ( .INP(n16130), .ZN(n16129) );
  OR2X1 U17038 ( .IN1(n590), .IN2(n8976), .Q(n16130) );
  AND2X1 U17039 ( .IN1(n4422), .IN2(n590), .Q(n16128) );
  OR2X1 U17040 ( .IN1(n16131), .IN2(n16132), .Q(g20919) );
  INVX0 U17041 ( .INP(n16133), .ZN(n16132) );
  OR2X1 U17042 ( .IN1(n14312), .IN2(n8868), .Q(n16133) );
  AND2X1 U17043 ( .IN1(n4415), .IN2(n14312), .Q(n16131) );
  OR2X1 U17044 ( .IN1(n16134), .IN2(n16135), .Q(g20918) );
  INVX0 U17045 ( .INP(n16136), .ZN(n16135) );
  OR2X1 U17046 ( .IN1(n14312), .IN2(n8886), .Q(n16136) );
  AND2X1 U17047 ( .IN1(n4398), .IN2(n14312), .Q(n16134) );
  INVX0 U17048 ( .INP(n14311), .ZN(n14312) );
  OR2X1 U17049 ( .IN1(n4306), .IN2(n16093), .Q(n14311) );
  OR2X1 U17050 ( .IN1(g2733), .IN2(n16038), .Q(n16093) );
  OR2X1 U17051 ( .IN1(n8825), .IN2(n4490), .Q(n16038) );
  OR2X1 U17052 ( .IN1(n16137), .IN2(n16138), .Q(g20917) );
  AND2X1 U17053 ( .IN1(n4416), .IN2(n14387), .Q(n16138) );
  AND2X1 U17054 ( .IN1(test_so72), .IN2(n14388), .Q(n16137) );
  OR2X1 U17055 ( .IN1(n16139), .IN2(n16140), .Q(g20916) );
  INVX0 U17056 ( .INP(n16141), .ZN(n16140) );
  OR2X1 U17057 ( .IN1(n14396), .IN2(n8902), .Q(n16141) );
  AND2X1 U17058 ( .IN1(n14396), .IN2(n4474), .Q(n16139) );
  OR2X1 U17059 ( .IN1(n16142), .IN2(n16143), .Q(g20915) );
  INVX0 U17060 ( .INP(n16144), .ZN(n16143) );
  OR2X1 U17061 ( .IN1(n14387), .IN2(n8903), .Q(n16144) );
  AND2X1 U17062 ( .IN1(n4400), .IN2(n14387), .Q(n16142) );
  INVX0 U17063 ( .INP(n14388), .ZN(n14387) );
  OR2X1 U17064 ( .IN1(n16106), .IN2(n16145), .Q(n14388) );
  OR2X1 U17065 ( .IN1(n4357), .IN2(g2039), .Q(n16145) );
  OR2X1 U17066 ( .IN1(n16146), .IN2(n16147), .Q(g20913) );
  INVX0 U17067 ( .INP(n16148), .ZN(n16147) );
  OR2X1 U17068 ( .IN1(n14392), .IN2(n8959), .Q(n16148) );
  AND2X1 U17069 ( .IN1(n4417), .IN2(n14392), .Q(n16146) );
  OR2X1 U17070 ( .IN1(n16149), .IN2(n16150), .Q(g20912) );
  INVX0 U17071 ( .INP(n16151), .ZN(n16150) );
  OR2X1 U17072 ( .IN1(n14484), .IN2(n8919), .Q(n16151) );
  AND2X1 U17073 ( .IN1(n4421), .IN2(n14484), .Q(n16149) );
  OR2X1 U17074 ( .IN1(n16152), .IN2(n16153), .Q(g20911) );
  INVX0 U17075 ( .INP(n16154), .ZN(n16153) );
  OR2X1 U17076 ( .IN1(n869), .IN2(n8920), .Q(n16154) );
  AND2X1 U17077 ( .IN1(n869), .IN2(n4476), .Q(n16152) );
  OR2X1 U17078 ( .IN1(n16155), .IN2(n16156), .Q(g20910) );
  INVX0 U17079 ( .INP(n16157), .ZN(n16156) );
  OR2X1 U17080 ( .IN1(n14392), .IN2(n8968), .Q(n16157) );
  AND2X1 U17081 ( .IN1(n4402), .IN2(n14392), .Q(n16155) );
  INVX0 U17082 ( .INP(n14393), .ZN(n14392) );
  OR2X1 U17083 ( .IN1(n15701), .IN2(n16158), .Q(n14393) );
  OR2X1 U17084 ( .IN1(n16159), .IN2(n16160), .Q(g20903) );
  INVX0 U17085 ( .INP(n16161), .ZN(n16160) );
  OR2X1 U17086 ( .IN1(n14565), .IN2(n8934), .Q(n16161) );
  AND2X1 U17087 ( .IN1(n14565), .IN2(n4414), .Q(n16159) );
  OR2X1 U17088 ( .IN1(n16162), .IN2(n16163), .Q(g20902) );
  INVX0 U17089 ( .INP(n16164), .ZN(n16163) );
  OR2X1 U17090 ( .IN1(n14561), .IN2(n8935), .Q(n16164) );
  AND2X1 U17091 ( .IN1(n4422), .IN2(n14561), .Q(n16162) );
  OR2X1 U17092 ( .IN1(n16165), .IN2(n16166), .Q(g20901) );
  INVX0 U17093 ( .INP(n16167), .ZN(n16166) );
  OR2X1 U17094 ( .IN1(n590), .IN2(n8977), .Q(n16167) );
  AND2X1 U17095 ( .IN1(n590), .IN2(n4478), .Q(n16165) );
  OR2X1 U17096 ( .IN1(n16168), .IN2(n16169), .Q(g20900) );
  INVX0 U17097 ( .INP(n16170), .ZN(n16169) );
  OR2X1 U17098 ( .IN1(n14396), .IN2(n8887), .Q(n16170) );
  AND2X1 U17099 ( .IN1(n4416), .IN2(n14396), .Q(n16168) );
  OR2X1 U17100 ( .IN1(n16171), .IN2(n16172), .Q(g20899) );
  INVX0 U17101 ( .INP(n16173), .ZN(n16172) );
  OR2X1 U17102 ( .IN1(n14396), .IN2(n8904), .Q(n16173) );
  AND2X1 U17103 ( .IN1(n4400), .IN2(n14396), .Q(n16171) );
  INVX0 U17104 ( .INP(n14469), .ZN(n14396) );
  OR2X1 U17105 ( .IN1(n16106), .IN2(n16174), .Q(n14469) );
  OR2X1 U17106 ( .IN1(n4307), .IN2(g2039), .Q(n16174) );
  OR2X1 U17107 ( .IN1(n8826), .IN2(n9127), .Q(n16106) );
  OR2X1 U17108 ( .IN1(n16175), .IN2(n16176), .Q(g20898) );
  INVX0 U17109 ( .INP(n16177), .ZN(n16176) );
  OR2X1 U17110 ( .IN1(n869), .IN2(n8905), .Q(n16177) );
  AND2X1 U17111 ( .IN1(n4417), .IN2(n869), .Q(n16175) );
  OR2X1 U17112 ( .IN1(n16178), .IN2(n16179), .Q(g20897) );
  INVX0 U17113 ( .INP(n16180), .ZN(n16179) );
  OR2X1 U17114 ( .IN1(n14484), .IN2(n8921), .Q(n16180) );
  AND2X1 U17115 ( .IN1(n14484), .IN2(n4476), .Q(n16178) );
  OR2X1 U17116 ( .IN1(n16181), .IN2(n16182), .Q(g20896) );
  INVX0 U17117 ( .INP(n16183), .ZN(n16182) );
  OR2X1 U17118 ( .IN1(n869), .IN2(n8922), .Q(n16183) );
  AND2X1 U17119 ( .IN1(n4402), .IN2(n869), .Q(n16181) );
  INVX0 U17120 ( .INP(n14472), .ZN(n869) );
  OR2X1 U17121 ( .IN1(n4358), .IN2(n16184), .Q(n14472) );
  OR2X1 U17122 ( .IN1(n16185), .IN2(n16186), .Q(g20894) );
  INVX0 U17123 ( .INP(n16187), .ZN(n16186) );
  OR2X1 U17124 ( .IN1(n590), .IN2(n8969), .Q(n16187) );
  AND2X1 U17125 ( .IN1(n4418), .IN2(n590), .Q(n16185) );
  OR2X1 U17126 ( .IN1(n16188), .IN2(n16189), .Q(g20893) );
  INVX0 U17127 ( .INP(n16190), .ZN(n16189) );
  OR2X1 U17128 ( .IN1(n14565), .IN2(n8936), .Q(n16190) );
  AND2X1 U17129 ( .IN1(n4422), .IN2(n14565), .Q(n16188) );
  OR2X1 U17130 ( .IN1(n16191), .IN2(n16192), .Q(g20892) );
  INVX0 U17131 ( .INP(n16193), .ZN(n16192) );
  OR2X1 U17132 ( .IN1(n14561), .IN2(n8937), .Q(n16193) );
  AND2X1 U17133 ( .IN1(n14561), .IN2(n4478), .Q(n16191) );
  OR2X1 U17134 ( .IN1(n16194), .IN2(n16195), .Q(g20891) );
  INVX0 U17135 ( .INP(n16196), .ZN(n16195) );
  OR2X1 U17136 ( .IN1(n590), .IN2(n8978), .Q(n16196) );
  AND2X1 U17137 ( .IN1(n4404), .IN2(n590), .Q(n16194) );
  INVX0 U17138 ( .INP(n14476), .ZN(n590) );
  OR2X1 U17139 ( .IN1(n15212), .IN2(n16197), .Q(n14476) );
  AND2X1 U17140 ( .IN1(n15185), .IN2(n7913), .Q(g20884) );
  INVX0 U17141 ( .INP(g3234), .ZN(n15185) );
  OR2X1 U17142 ( .IN1(n16198), .IN2(n16199), .Q(g20883) );
  INVX0 U17143 ( .INP(n16200), .ZN(n16199) );
  OR2X1 U17144 ( .IN1(n14484), .IN2(n8906), .Q(n16200) );
  AND2X1 U17145 ( .IN1(n4417), .IN2(n14484), .Q(n16198) );
  OR2X1 U17146 ( .IN1(n16201), .IN2(n16202), .Q(g20882) );
  AND2X1 U17147 ( .IN1(n4402), .IN2(n14484), .Q(n16202) );
  INVX0 U17148 ( .INP(n14483), .ZN(n14484) );
  AND2X1 U17149 ( .IN1(test_so49), .IN2(n14483), .Q(n16201) );
  OR2X1 U17150 ( .IN1(n4308), .IN2(n16184), .Q(n14483) );
  OR2X1 U17151 ( .IN1(g1345), .IN2(n16158), .Q(n16184) );
  OR2X1 U17152 ( .IN1(n8827), .IN2(n4489), .Q(n16158) );
  OR2X1 U17153 ( .IN1(n16203), .IN2(n16204), .Q(g20881) );
  AND2X1 U17154 ( .IN1(n4418), .IN2(n14561), .Q(n16204) );
  AND2X1 U17155 ( .IN1(test_so30), .IN2(n14560), .Q(n16203) );
  OR2X1 U17156 ( .IN1(n16205), .IN2(n16206), .Q(g20880) );
  INVX0 U17157 ( .INP(n16207), .ZN(n16206) );
  OR2X1 U17158 ( .IN1(n14565), .IN2(n8938), .Q(n16207) );
  AND2X1 U17159 ( .IN1(n14565), .IN2(n4478), .Q(n16205) );
  OR2X1 U17160 ( .IN1(n16208), .IN2(n16209), .Q(g20879) );
  INVX0 U17161 ( .INP(n16210), .ZN(n16209) );
  OR2X1 U17162 ( .IN1(n14561), .IN2(n8939), .Q(n16210) );
  AND2X1 U17163 ( .IN1(n4404), .IN2(n14561), .Q(n16208) );
  INVX0 U17164 ( .INP(n14560), .ZN(n14561) );
  OR2X1 U17165 ( .IN1(n4359), .IN2(n16211), .Q(n14560) );
  OR2X1 U17166 ( .IN1(n16212), .IN2(n16213), .Q(g20876) );
  INVX0 U17167 ( .INP(n16214), .ZN(n16213) );
  OR2X1 U17168 ( .IN1(n14565), .IN2(n8923), .Q(n16214) );
  AND2X1 U17169 ( .IN1(n4418), .IN2(n14565), .Q(n16212) );
  OR2X1 U17170 ( .IN1(n16215), .IN2(n16216), .Q(g20875) );
  INVX0 U17171 ( .INP(n16217), .ZN(n16216) );
  OR2X1 U17172 ( .IN1(n14565), .IN2(n8940), .Q(n16217) );
  AND2X1 U17173 ( .IN1(n4404), .IN2(n14565), .Q(n16215) );
  INVX0 U17174 ( .INP(n14564), .ZN(n14565) );
  OR2X1 U17175 ( .IN1(n4309), .IN2(n16211), .Q(n14564) );
  OR2X1 U17176 ( .IN1(g659), .IN2(n16197), .Q(n16211) );
  OR2X1 U17177 ( .IN1(n8828), .IN2(n4492), .Q(n16197) );
  OR2X1 U17178 ( .IN1(n16218), .IN2(n16219), .Q(g20874) );
  AND2X1 U17179 ( .IN1(n4351), .IN2(n15708), .Q(n16219) );
  XOR2X1 U17180 ( .IN1(n15711), .IN2(n9519), .Q(n15708) );
  XNOR2X1 U17181 ( .IN1(n16220), .IN2(n16221), .Q(n9519) );
  XOR2X1 U17182 ( .IN1(n16222), .IN2(n16223), .Q(n16221) );
  XNOR2X1 U17183 ( .IN1(g2953), .IN2(n9063), .Q(n16223) );
  XNOR2X1 U17184 ( .IN1(g2956), .IN2(n9065), .Q(n16222) );
  XOR2X1 U17185 ( .IN1(n16224), .IN2(n16225), .Q(n16220) );
  XNOR2X1 U17186 ( .IN1(g2938), .IN2(n9061), .Q(n16225) );
  XNOR2X1 U17187 ( .IN1(n9059), .IN2(n9060), .Q(n16224) );
  OR2X1 U17188 ( .IN1(n16494), .IN2(g3231), .Q(n15711) );
  AND2X1 U17189 ( .IN1(g2879), .IN2(g8096), .Q(n16218) );
  AND2X1 U17190 ( .IN1(n16226), .IN2(n12737), .Q(g20789) );
  OR2X1 U17191 ( .IN1(n4356), .IN2(n9085), .Q(n12737) );
  XOR2X1 U17192 ( .IN1(n15683), .IN2(n4398), .Q(n16226) );
  OR2X1 U17193 ( .IN1(n4292), .IN2(g2733), .Q(n15683) );
  AND2X1 U17194 ( .IN1(n16227), .IN2(n12741), .Q(g20752) );
  OR2X1 U17195 ( .IN1(n4357), .IN2(n9084), .Q(n12741) );
  XOR2X1 U17196 ( .IN1(n15689), .IN2(n4400), .Q(n16227) );
  OR2X1 U17197 ( .IN1(n4293), .IN2(g2039), .Q(n15689) );
  AND2X1 U17198 ( .IN1(n16228), .IN2(n12745), .Q(g20717) );
  OR2X1 U17199 ( .IN1(n4358), .IN2(n9083), .Q(n12745) );
  XOR2X1 U17200 ( .IN1(n15701), .IN2(n4402), .Q(n16228) );
  OR2X1 U17201 ( .IN1(n4294), .IN2(g1345), .Q(n15701) );
  AND2X1 U17202 ( .IN1(n16229), .IN2(n12226), .Q(g20682) );
  OR2X1 U17203 ( .IN1(n4359), .IN2(n9082), .Q(n12226) );
  XOR2X1 U17204 ( .IN1(n15212), .IN2(n4404), .Q(n16229) );
  OR2X1 U17205 ( .IN1(n4295), .IN2(g659), .Q(n15212) );
  OR2X1 U17206 ( .IN1(n16230), .IN2(n16231), .Q(g20417) );
  AND2X1 U17207 ( .IN1(g2879), .IN2(g7334), .Q(n16231) );
  AND2X1 U17208 ( .IN1(n4351), .IN2(g2963), .Q(n16230) );
  OR2X1 U17209 ( .IN1(n16232), .IN2(n16233), .Q(g20376) );
  AND2X1 U17210 ( .IN1(g2879), .IN2(g6895), .Q(n16233) );
  AND2X1 U17211 ( .IN1(test_so2), .IN2(n4351), .Q(n16232) );
  OR2X1 U17212 ( .IN1(n16234), .IN2(n16235), .Q(g20375) );
  AND2X1 U17213 ( .IN1(n15317), .IN2(g2703), .Q(n16235) );
  AND2X1 U17214 ( .IN1(n4292), .IN2(g2733), .Q(n16234) );
  OR2X1 U17215 ( .IN1(n16236), .IN2(n16237), .Q(g20353) );
  AND2X1 U17216 ( .IN1(n15317), .IN2(g2009), .Q(n16237) );
  AND2X1 U17217 ( .IN1(n4293), .IN2(g2039), .Q(n16236) );
  OR2X1 U17218 ( .IN1(n16238), .IN2(n16239), .Q(g20343) );
  AND2X1 U17219 ( .IN1(g2879), .IN2(g6442), .Q(n16239) );
  AND2X1 U17220 ( .IN1(n4351), .IN2(g2969), .Q(n16238) );
  OR2X1 U17221 ( .IN1(n16240), .IN2(n16241), .Q(g20333) );
  AND2X1 U17222 ( .IN1(n15317), .IN2(g1315), .Q(n16241) );
  AND2X1 U17223 ( .IN1(n4294), .IN2(g1345), .Q(n16240) );
  OR2X1 U17224 ( .IN1(n16242), .IN2(n16243), .Q(g20314) );
  AND2X1 U17225 ( .IN1(n15317), .IN2(g629), .Q(n16243) );
  AND2X1 U17226 ( .IN1(n16244), .IN2(n16245), .Q(n15317) );
  AND2X1 U17227 ( .IN1(n8282), .IN2(n9092), .Q(n16245) );
  AND2X1 U17228 ( .IN1(n8281), .IN2(n16246), .Q(n16244) );
  INVX0 U17229 ( .INP(n16247), .ZN(n16246) );
  OR2X1 U17230 ( .IN1(test_so98), .IN2(g3006), .Q(n16247) );
  AND2X1 U17231 ( .IN1(n4295), .IN2(g659), .Q(n16242) );
  OR2X1 U17232 ( .IN1(n16248), .IN2(n16249), .Q(g20310) );
  AND2X1 U17233 ( .IN1(g2879), .IN2(g6225), .Q(n16249) );
  AND2X1 U17234 ( .IN1(n4351), .IN2(g2972), .Q(n16248) );
  OR2X1 U17235 ( .IN1(n16250), .IN2(n16251), .Q(g19184) );
  AND2X1 U17236 ( .IN1(g2879), .IN2(g4590), .Q(n16251) );
  AND2X1 U17237 ( .IN1(n4351), .IN2(g2975), .Q(n16250) );
  OR2X1 U17238 ( .IN1(n16252), .IN2(n16253), .Q(g19178) );
  AND2X1 U17239 ( .IN1(test_so5), .IN2(g2879), .Q(n16253) );
  AND2X1 U17240 ( .IN1(n4351), .IN2(g2935), .Q(n16252) );
  OR2X1 U17241 ( .IN1(n16254), .IN2(n16255), .Q(g19173) );
  AND2X1 U17242 ( .IN1(g2879), .IN2(g4323), .Q(n16255) );
  AND2X1 U17243 ( .IN1(n4351), .IN2(g2978), .Q(n16254) );
  OR2X1 U17244 ( .IN1(n16256), .IN2(n16257), .Q(g19172) );
  AND2X1 U17245 ( .IN1(g2879), .IN2(g4321), .Q(n16257) );
  AND2X1 U17246 ( .IN1(n4351), .IN2(g2953), .Q(n16256) );
  OR2X1 U17247 ( .IN1(n16258), .IN2(n16259), .Q(g19167) );
  AND2X1 U17248 ( .IN1(g2879), .IN2(g4200), .Q(n16259) );
  AND2X1 U17249 ( .IN1(n4351), .IN2(g2938), .Q(n16258) );
  OR2X1 U17250 ( .IN1(n16260), .IN2(n16261), .Q(g19163) );
  AND2X1 U17251 ( .IN1(g2879), .IN2(g4090), .Q(n16261) );
  AND2X1 U17252 ( .IN1(n4351), .IN2(g2981), .Q(n16260) );
  OR2X1 U17253 ( .IN1(n16262), .IN2(n16263), .Q(g19162) );
  AND2X1 U17254 ( .IN1(g2879), .IN2(g4088), .Q(n16263) );
  AND2X1 U17255 ( .IN1(n4351), .IN2(g2956), .Q(n16262) );
  OR2X1 U17256 ( .IN1(n16264), .IN2(n16265), .Q(g19157) );
  AND2X1 U17257 ( .IN1(g2879), .IN2(g3993), .Q(n16265) );
  AND2X1 U17258 ( .IN1(n4351), .IN2(g2941), .Q(n16264) );
  OR2X1 U17259 ( .IN1(n16266), .IN2(n16267), .Q(g19154) );
  AND2X1 U17260 ( .IN1(test_so3), .IN2(g2879), .Q(n16267) );
  AND2X1 U17261 ( .IN1(n4351), .IN2(g2874), .Q(n16266) );
  OR2X1 U17262 ( .IN1(n16268), .IN2(n16269), .Q(g19153) );
  AND2X1 U17263 ( .IN1(g2879), .IN2(g8249), .Q(n16269) );
  AND2X1 U17264 ( .IN1(n4351), .IN2(g2959), .Q(n16268) );
  OR2X1 U17265 ( .IN1(n16270), .IN2(n16271), .Q(g19149) );
  AND2X1 U17266 ( .IN1(g2879), .IN2(g8175), .Q(n16271) );
  AND2X1 U17267 ( .IN1(n4351), .IN2(g2944), .Q(n16270) );
  OR2X1 U17268 ( .IN1(n16272), .IN2(n16273), .Q(g19144) );
  AND2X1 U17269 ( .IN1(g2879), .IN2(g8023), .Q(n16273) );
  AND2X1 U17270 ( .IN1(n4351), .IN2(g2947), .Q(n16272) );
  OR2X1 U17271 ( .IN1(n16274), .IN2(n16275), .Q(g18975) );
  AND2X1 U17272 ( .IN1(g2879), .IN2(g2981), .Q(n16275) );
  AND2X1 U17273 ( .IN1(n4351), .IN2(g2195), .Q(n16274) );
  OR2X1 U17274 ( .IN1(n16276), .IN2(n16277), .Q(g18968) );
  AND2X1 U17275 ( .IN1(g2879), .IN2(g2978), .Q(n16277) );
  AND2X1 U17276 ( .IN1(n4351), .IN2(g2190), .Q(n16276) );
  OR2X1 U17277 ( .IN1(n16278), .IN2(n16279), .Q(g18957) );
  AND2X1 U17278 ( .IN1(g2879), .IN2(g2963), .Q(n16279) );
  AND2X1 U17279 ( .IN1(n4351), .IN2(g2165), .Q(n16278) );
  OR2X1 U17280 ( .IN1(n16280), .IN2(n16281), .Q(g18942) );
  AND2X1 U17281 ( .IN1(n4351), .IN2(g2185), .Q(n16281) );
  AND2X1 U17282 ( .IN1(g2879), .IN2(g2975), .Q(n16280) );
  OR2X1 U17283 ( .IN1(n16282), .IN2(n16283), .Q(g18907) );
  AND2X1 U17284 ( .IN1(g2987), .IN2(g2997), .Q(n16283) );
  AND2X1 U17285 ( .IN1(n4365), .IN2(g3061), .Q(n16282) );
  OR2X1 U17286 ( .IN1(n16284), .IN2(n16285), .Q(g18906) );
  AND2X1 U17287 ( .IN1(g2879), .IN2(g2972), .Q(n16285) );
  AND2X1 U17288 ( .IN1(n4351), .IN2(g2180), .Q(n16284) );
  OR2X1 U17289 ( .IN1(n16286), .IN2(n16287), .Q(g18885) );
  AND2X1 U17290 ( .IN1(n4351), .IN2(g2200), .Q(n16287) );
  AND2X1 U17291 ( .IN1(g2879), .IN2(g2874), .Q(n16286) );
  OR2X1 U17292 ( .IN1(n16288), .IN2(n16289), .Q(g18883) );
  AND2X1 U17293 ( .IN1(g2879), .IN2(g2935), .Q(n16289) );
  AND2X1 U17294 ( .IN1(n4351), .IN2(g1471), .Q(n16288) );
  OR2X1 U17295 ( .IN1(n16290), .IN2(n16291), .Q(g18868) );
  AND2X1 U17296 ( .IN1(g2987), .IN2(g3078), .Q(n16291) );
  AND2X1 U17297 ( .IN1(n4365), .IN2(g3060), .Q(n16290) );
  OR2X1 U17298 ( .IN1(n16292), .IN2(n16293), .Q(g18867) );
  AND2X1 U17299 ( .IN1(n4351), .IN2(g2175), .Q(n16293) );
  AND2X1 U17300 ( .IN1(g2879), .IN2(g2969), .Q(n16292) );
  OR2X1 U17301 ( .IN1(n16294), .IN2(n16295), .Q(g18866) );
  AND2X1 U17302 ( .IN1(g2879), .IN2(g2938), .Q(n16295) );
  AND2X1 U17303 ( .IN1(n4351), .IN2(g1476), .Q(n16294) );
  OR2X1 U17304 ( .IN1(n16296), .IN2(n16297), .Q(g18852) );
  AND2X1 U17305 ( .IN1(n4351), .IN2(g1481), .Q(n16297) );
  AND2X1 U17306 ( .IN1(g2879), .IN2(g2941), .Q(n16296) );
  OR2X1 U17307 ( .IN1(n16298), .IN2(n16299), .Q(g18837) );
  AND2X1 U17308 ( .IN1(g2987), .IN2(g3077), .Q(n16299) );
  AND2X1 U17309 ( .IN1(n4365), .IN2(g3059), .Q(n16298) );
  OR2X1 U17310 ( .IN1(n16300), .IN2(n16301), .Q(g18836) );
  AND2X1 U17311 ( .IN1(test_so2), .IN2(g2879), .Q(n16301) );
  AND2X1 U17312 ( .IN1(n4351), .IN2(g2170), .Q(n16300) );
  OR2X1 U17313 ( .IN1(n16302), .IN2(n16303), .Q(g18835) );
  AND2X1 U17314 ( .IN1(g2879), .IN2(g2944), .Q(n16303) );
  AND2X1 U17315 ( .IN1(n4351), .IN2(g1486), .Q(n16302) );
  OR2X1 U17316 ( .IN1(n16304), .IN2(n16305), .Q(g18821) );
  AND2X1 U17317 ( .IN1(n4351), .IN2(g1491), .Q(n16305) );
  AND2X1 U17318 ( .IN1(g2879), .IN2(g2947), .Q(n16304) );
  OR2X1 U17319 ( .IN1(n16306), .IN2(n16307), .Q(g18820) );
  AND2X1 U17320 ( .IN1(g2624), .IN2(g2631), .Q(n16307) );
  AND2X1 U17321 ( .IN1(n4299), .IN2(g2584), .Q(n16306) );
  OR2X1 U17322 ( .IN1(n16308), .IN2(n16309), .Q(g18804) );
  AND2X1 U17323 ( .IN1(g2987), .IN2(g3076), .Q(n16309) );
  AND2X1 U17324 ( .IN1(n4365), .IN2(g3058), .Q(n16308) );
  OR2X1 U17325 ( .IN1(n16310), .IN2(n16311), .Q(g18803) );
  AND2X1 U17326 ( .IN1(g2879), .IN2(g2953), .Q(n16311) );
  AND2X1 U17327 ( .IN1(n4351), .IN2(g1496), .Q(n16310) );
  OR2X1 U17328 ( .IN1(n16312), .IN2(n16313), .Q(g18794) );
  AND2X1 U17329 ( .IN1(n4366), .IN2(g1890), .Q(n16313) );
  AND2X1 U17330 ( .IN1(g1937), .IN2(g1930), .Q(n16312) );
  OR2X1 U17331 ( .IN1(n16314), .IN2(n16315), .Q(g18782) );
  AND2X1 U17332 ( .IN1(n4494), .IN2(g3084), .Q(n16315) );
  AND2X1 U17333 ( .IN1(g3109), .IN2(g559), .Q(n16314) );
  OR2X1 U17334 ( .IN1(n16316), .IN2(n16317), .Q(g18781) );
  AND2X1 U17335 ( .IN1(g2879), .IN2(g2956), .Q(n16317) );
  AND2X1 U17336 ( .IN1(n4351), .IN2(g1501), .Q(n16316) );
  OR2X1 U17337 ( .IN1(n16318), .IN2(n16319), .Q(g18780) );
  AND2X1 U17338 ( .IN1(n9050), .IN2(g2624), .Q(n16319) );
  AND2X1 U17339 ( .IN1(n4299), .IN2(g2631), .Q(n16318) );
  OR2X1 U17340 ( .IN1(n16320), .IN2(n16321), .Q(g18763) );
  AND2X1 U17341 ( .IN1(g1236), .IN2(g1243), .Q(n16321) );
  AND2X1 U17342 ( .IN1(n4300), .IN2(g1196), .Q(n16320) );
  OR2X1 U17343 ( .IN1(n16322), .IN2(n16323), .Q(g18755) );
  AND2X1 U17344 ( .IN1(g2987), .IN2(g3075), .Q(n16323) );
  AND2X1 U17345 ( .IN1(n4365), .IN2(g3057), .Q(n16322) );
  OR2X1 U17346 ( .IN1(n16324), .IN2(n16325), .Q(g18754) );
  AND2X1 U17347 ( .IN1(n4351), .IN2(g1506), .Q(n16325) );
  AND2X1 U17348 ( .IN1(g2879), .IN2(g2959), .Q(n16324) );
  OR2X1 U17349 ( .IN1(n16326), .IN2(n16327), .Q(g18743) );
  AND2X1 U17350 ( .IN1(n4366), .IN2(g1937), .Q(n16327) );
  AND2X1 U17351 ( .IN1(n9051), .IN2(g1930), .Q(n16326) );
  OR2X1 U17352 ( .IN1(n16328), .IN2(n16329), .Q(g18726) );
  AND2X1 U17353 ( .IN1(g550), .IN2(g557), .Q(n16329) );
  AND2X1 U17354 ( .IN1(n4313), .IN2(test_so22), .Q(n16328) );
  OR2X1 U17355 ( .IN1(n16330), .IN2(n16331), .Q(g18719) );
  AND2X1 U17356 ( .IN1(g8030), .IN2(g559), .Q(n16331) );
  AND2X1 U17357 ( .IN1(n4383), .IN2(g3211), .Q(n16330) );
  OR2X1 U17358 ( .IN1(n16332), .IN2(n16333), .Q(g18707) );
  AND2X1 U17359 ( .IN1(n9052), .IN2(g1236), .Q(n16333) );
  AND2X1 U17360 ( .IN1(n4300), .IN2(g1243), .Q(n16332) );
  OR2X1 U17361 ( .IN1(n16334), .IN2(n16335), .Q(g18678) );
  AND2X1 U17362 ( .IN1(n9053), .IN2(g550), .Q(n16335) );
  AND2X1 U17363 ( .IN1(n4313), .IN2(g557), .Q(n16334) );
  OR2X1 U17364 ( .IN1(n16336), .IN2(n16337), .Q(g18669) );
  AND2X1 U17365 ( .IN1(g8106), .IN2(g559), .Q(n16337) );
  AND2X1 U17366 ( .IN1(n4382), .IN2(test_so6), .Q(n16336) );
  OR2X1 U17367 ( .IN1(n16338), .IN2(n16339), .Q(g17429) );
  AND2X1 U17368 ( .IN1(n4494), .IN2(g3088), .Q(n16339) );
  AND2X1 U17369 ( .IN1(g3109), .IN2(g2574), .Q(n16338) );
  OR2X1 U17370 ( .IN1(n16340), .IN2(n16341), .Q(g17383) );
  AND2X1 U17371 ( .IN1(g3109), .IN2(g1880), .Q(n16341) );
  AND2X1 U17372 ( .IN1(n4494), .IN2(test_so8), .Q(n16340) );
  OR2X1 U17373 ( .IN1(n16342), .IN2(n16343), .Q(g17341) );
  AND2X1 U17374 ( .IN1(g8030), .IN2(g2574), .Q(n16343) );
  AND2X1 U17375 ( .IN1(n4383), .IN2(g3185), .Q(n16342) );
  OR2X1 U17376 ( .IN1(n16344), .IN2(n16345), .Q(g17340) );
  AND2X1 U17377 ( .IN1(n4494), .IN2(g3170), .Q(n16345) );
  AND2X1 U17378 ( .IN1(g3109), .IN2(g1186), .Q(n16344) );
  OR2X1 U17379 ( .IN1(n16346), .IN2(n16347), .Q(g17303) );
  AND2X1 U17380 ( .IN1(g8030), .IN2(g1880), .Q(n16347) );
  AND2X1 U17381 ( .IN1(n4383), .IN2(g3176), .Q(n16346) );
  OR2X1 U17382 ( .IN1(n16348), .IN2(n16349), .Q(g17302) );
  AND2X1 U17383 ( .IN1(n4494), .IN2(g3161), .Q(n16349) );
  AND2X1 U17384 ( .IN1(g3109), .IN2(g499), .Q(n16348) );
  OR2X1 U17385 ( .IN1(n16350), .IN2(n16351), .Q(g17271) );
  AND2X1 U17386 ( .IN1(g8106), .IN2(g2574), .Q(n16351) );
  AND2X1 U17387 ( .IN1(n4382), .IN2(g3182), .Q(n16350) );
  OR2X1 U17388 ( .IN1(n16352), .IN2(n16353), .Q(g17270) );
  AND2X1 U17389 ( .IN1(n4383), .IN2(g3167), .Q(n16353) );
  AND2X1 U17390 ( .IN1(g8030), .IN2(g1186), .Q(n16352) );
  OR2X1 U17391 ( .IN1(n16354), .IN2(n16355), .Q(g17269) );
  AND2X1 U17392 ( .IN1(n4494), .IN2(g3096), .Q(n16355) );
  AND2X1 U17393 ( .IN1(g3109), .IN2(g2633), .Q(n16354) );
  OR2X1 U17394 ( .IN1(n16356), .IN2(n16357), .Q(g17248) );
  AND2X1 U17395 ( .IN1(n4382), .IN2(g3173), .Q(n16357) );
  AND2X1 U17396 ( .IN1(g8106), .IN2(g1880), .Q(n16356) );
  OR2X1 U17397 ( .IN1(n16358), .IN2(n16359), .Q(g17247) );
  AND2X1 U17398 ( .IN1(g8030), .IN2(g499), .Q(n16359) );
  AND2X1 U17399 ( .IN1(n4383), .IN2(g3158), .Q(n16358) );
  OR2X1 U17400 ( .IN1(n16360), .IN2(n16361), .Q(g17246) );
  AND2X1 U17401 ( .IN1(n4494), .IN2(g3093), .Q(n16361) );
  AND2X1 U17402 ( .IN1(g3109), .IN2(g1939), .Q(n16360) );
  OR2X1 U17403 ( .IN1(n16362), .IN2(n16363), .Q(g17236) );
  AND2X1 U17404 ( .IN1(n4382), .IN2(g3164), .Q(n16363) );
  AND2X1 U17405 ( .IN1(g8106), .IN2(g1186), .Q(n16362) );
  OR2X1 U17406 ( .IN1(n16364), .IN2(n16365), .Q(g17235) );
  AND2X1 U17407 ( .IN1(g8030), .IN2(g2633), .Q(n16365) );
  AND2X1 U17408 ( .IN1(n4383), .IN2(g3095), .Q(n16364) );
  OR2X1 U17409 ( .IN1(n16366), .IN2(n16367), .Q(g17234) );
  AND2X1 U17410 ( .IN1(n4494), .IN2(g3087), .Q(n16367) );
  AND2X1 U17411 ( .IN1(g3109), .IN2(g1245), .Q(n16366) );
  OR2X1 U17412 ( .IN1(n16368), .IN2(n16369), .Q(g17229) );
  AND2X1 U17413 ( .IN1(g8106), .IN2(g499), .Q(n16369) );
  AND2X1 U17414 ( .IN1(n4382), .IN2(g3155), .Q(n16368) );
  OR2X1 U17415 ( .IN1(n16370), .IN2(n16371), .Q(g17228) );
  AND2X1 U17416 ( .IN1(g8030), .IN2(g1939), .Q(n16371) );
  AND2X1 U17417 ( .IN1(n4383), .IN2(g3092), .Q(n16370) );
  OR2X1 U17418 ( .IN1(n16372), .IN2(n16373), .Q(g17226) );
  AND2X1 U17419 ( .IN1(g8106), .IN2(g2633), .Q(n16373) );
  AND2X1 U17420 ( .IN1(n4382), .IN2(g3094), .Q(n16372) );
  OR2X1 U17421 ( .IN1(n16374), .IN2(n16375), .Q(g17225) );
  AND2X1 U17422 ( .IN1(n4383), .IN2(g3086), .Q(n16375) );
  AND2X1 U17423 ( .IN1(g8030), .IN2(g1245), .Q(n16374) );
  OR2X1 U17424 ( .IN1(n16376), .IN2(n16377), .Q(g17224) );
  AND2X1 U17425 ( .IN1(g8106), .IN2(g1939), .Q(n16377) );
  AND2X1 U17426 ( .IN1(n4382), .IN2(g3091), .Q(n16376) );
  OR2X1 U17427 ( .IN1(n16378), .IN2(n16379), .Q(g17222) );
  AND2X1 U17428 ( .IN1(n4382), .IN2(g3085), .Q(n16379) );
  AND2X1 U17429 ( .IN1(g8106), .IN2(g1245), .Q(n16378) );
  OR2X1 U17430 ( .IN1(n16380), .IN2(n16381), .Q(g16880) );
  AND2X1 U17431 ( .IN1(g2987), .IN2(g3074), .Q(n16381) );
  AND2X1 U17432 ( .IN1(n4365), .IN2(g3056), .Q(n16380) );
  OR2X1 U17433 ( .IN1(n16382), .IN2(n16383), .Q(g16866) );
  AND2X1 U17434 ( .IN1(test_so97), .IN2(g2987), .Q(n16383) );
  AND2X1 U17435 ( .IN1(n4365), .IN2(g3051), .Q(n16382) );
  OR2X1 U17436 ( .IN1(n16384), .IN2(n16385), .Q(g16861) );
  AND2X1 U17437 ( .IN1(g2987), .IN2(g3073), .Q(n16385) );
  AND2X1 U17438 ( .IN1(test_so96), .IN2(n4365), .Q(n16384) );
  OR2X1 U17439 ( .IN1(n16386), .IN2(n16387), .Q(g16860) );
  AND2X1 U17440 ( .IN1(g2987), .IN2(g3065), .Q(n16387) );
  AND2X1 U17441 ( .IN1(n4365), .IN2(g3046), .Q(n16386) );
  OR2X1 U17442 ( .IN1(n16388), .IN2(n16389), .Q(g16857) );
  AND2X1 U17443 ( .IN1(g2987), .IN2(g3069), .Q(n16389) );
  AND2X1 U17444 ( .IN1(n4365), .IN2(g3050), .Q(n16388) );
  OR2X1 U17445 ( .IN1(n16390), .IN2(n16391), .Q(g16854) );
  AND2X1 U17446 ( .IN1(g2987), .IN2(g3072), .Q(n16391) );
  AND2X1 U17447 ( .IN1(n4365), .IN2(g3053), .Q(n16390) );
  OR2X1 U17448 ( .IN1(n16392), .IN2(n16393), .Q(g16853) );
  AND2X1 U17449 ( .IN1(g2987), .IN2(g3064), .Q(n16393) );
  AND2X1 U17450 ( .IN1(n4365), .IN2(g3045), .Q(n16392) );
  OR2X1 U17451 ( .IN1(n16394), .IN2(n16395), .Q(g16851) );
  AND2X1 U17452 ( .IN1(g2987), .IN2(g3068), .Q(n16395) );
  AND2X1 U17453 ( .IN1(n4365), .IN2(g3049), .Q(n16394) );
  OR2X1 U17454 ( .IN1(n16396), .IN2(n16397), .Q(g16845) );
  AND2X1 U17455 ( .IN1(g2987), .IN2(g3071), .Q(n16397) );
  AND2X1 U17456 ( .IN1(n4365), .IN2(g3052), .Q(n16396) );
  OR2X1 U17457 ( .IN1(n16398), .IN2(n16399), .Q(g16844) );
  AND2X1 U17458 ( .IN1(g2987), .IN2(g3063), .Q(n16399) );
  AND2X1 U17459 ( .IN1(n4365), .IN2(g3044), .Q(n16398) );
  OR2X1 U17460 ( .IN1(n16400), .IN2(n16401), .Q(g16835) );
  AND2X1 U17461 ( .IN1(g2987), .IN2(g3067), .Q(n16401) );
  AND2X1 U17462 ( .IN1(n4365), .IN2(g3048), .Q(n16400) );
  OR2X1 U17463 ( .IN1(n16402), .IN2(n16403), .Q(g16824) );
  AND2X1 U17464 ( .IN1(g2987), .IN2(g3062), .Q(n16403) );
  AND2X1 U17465 ( .IN1(n4365), .IN2(g3043), .Q(n16402) );
  AND2X1 U17466 ( .IN1(n16404), .IN2(n8103), .Q(g16823) );
  OR2X1 U17467 ( .IN1(n16405), .IN2(n16406), .Q(g16803) );
  AND2X1 U17468 ( .IN1(g2987), .IN2(g3066), .Q(n16406) );
  AND2X1 U17469 ( .IN1(n4365), .IN2(g3047), .Q(n16405) );
  AND2X1 U17470 ( .IN1(n16404), .IN2(g2950), .Q(g16802) );
  INVX0 U17471 ( .INP(g51), .ZN(n16404) );
  OR2X1 U17472 ( .IN1(n16407), .IN2(n16408), .Q(g16718) );
  AND2X1 U17473 ( .IN1(g2703), .IN2(g2584), .Q(n16408) );
  INVX0 U17474 ( .INP(n16409), .ZN(n16407) );
  OR2X1 U17475 ( .IN1(g2703), .IN2(n9085), .Q(n16409) );
  OR2X1 U17476 ( .IN1(n16410), .IN2(n16411), .Q(g16692) );
  AND2X1 U17477 ( .IN1(g2009), .IN2(g1890), .Q(n16411) );
  INVX0 U17478 ( .INP(n16412), .ZN(n16410) );
  OR2X1 U17479 ( .IN1(g2009), .IN2(n9084), .Q(n16412) );
  OR2X1 U17480 ( .IN1(n16413), .IN2(n16414), .Q(g16671) );
  AND2X1 U17481 ( .IN1(g1315), .IN2(g1196), .Q(n16414) );
  INVX0 U17482 ( .INP(n16415), .ZN(n16413) );
  OR2X1 U17483 ( .IN1(g1315), .IN2(n9083), .Q(n16415) );
  OR2X1 U17484 ( .IN1(n16416), .IN2(n16417), .Q(g16654) );
  AND2X1 U17485 ( .IN1(test_so22), .IN2(g629), .Q(n16417) );
  INVX0 U17486 ( .INP(n16418), .ZN(n16416) );
  OR2X1 U17487 ( .IN1(g629), .IN2(n9082), .Q(n16418) );
  OR2X1 U17488 ( .IN1(n4365), .IN2(n16419), .Q(g16496) );
  AND2X1 U17489 ( .IN1(DFF_1612_n1), .IN2(g5388), .Q(n16419) );
  AND2X1 U17490 ( .IN1(n16420), .IN2(n16421), .Q(g13194) );
  OR2X1 U17491 ( .IN1(n4370), .IN2(g2561), .Q(n16421) );
  AND2X1 U17492 ( .IN1(n16422), .IN2(n16423), .Q(n16420) );
  OR2X1 U17493 ( .IN1(n4299), .IN2(g2562), .Q(n16423) );
  OR2X1 U17494 ( .IN1(n4314), .IN2(test_so87), .Q(n16422) );
  AND2X1 U17495 ( .IN1(n16424), .IN2(n16425), .Q(g13182) );
  OR2X1 U17496 ( .IN1(n4315), .IN2(g1867), .Q(n16425) );
  AND2X1 U17497 ( .IN1(n16426), .IN2(n16427), .Q(n16424) );
  OR2X1 U17498 ( .IN1(n4366), .IN2(g1868), .Q(n16427) );
  OR2X1 U17499 ( .IN1(n4296), .IN2(g1869), .Q(n16426) );
  AND2X1 U17500 ( .IN1(n16428), .IN2(n16429), .Q(g13175) );
  OR2X1 U17501 ( .IN1(n4370), .IN2(g2552), .Q(n16429) );
  AND2X1 U17502 ( .IN1(n16430), .IN2(n16431), .Q(n16428) );
  OR2X1 U17503 ( .IN1(n4299), .IN2(g2553), .Q(n16431) );
  OR2X1 U17504 ( .IN1(n4314), .IN2(g2554), .Q(n16430) );
  AND2X1 U17505 ( .IN1(n16432), .IN2(n16433), .Q(g13171) );
  OR2X1 U17506 ( .IN1(n4316), .IN2(g1173), .Q(n16433) );
  AND2X1 U17507 ( .IN1(n16434), .IN2(n16435), .Q(n16432) );
  OR2X1 U17508 ( .IN1(n4371), .IN2(g1175), .Q(n16435) );
  OR2X1 U17509 ( .IN1(n4300), .IN2(test_so44), .Q(n16434) );
  AND2X1 U17510 ( .IN1(n16436), .IN2(n16437), .Q(g13164) );
  OR2X1 U17511 ( .IN1(n4315), .IN2(g1858), .Q(n16437) );
  AND2X1 U17512 ( .IN1(n16438), .IN2(n16439), .Q(n16436) );
  OR2X1 U17513 ( .IN1(n4366), .IN2(g1859), .Q(n16439) );
  OR2X1 U17514 ( .IN1(n4296), .IN2(g1860), .Q(n16438) );
  AND2X1 U17515 ( .IN1(n16440), .IN2(n16441), .Q(g13160) );
  OR2X1 U17516 ( .IN1(n4372), .IN2(g486), .Q(n16441) );
  AND2X1 U17517 ( .IN1(n16442), .IN2(n16443), .Q(n16440) );
  OR2X1 U17518 ( .IN1(n4313), .IN2(g487), .Q(n16443) );
  OR2X1 U17519 ( .IN1(n4298), .IN2(g488), .Q(n16442) );
  AND2X1 U17520 ( .IN1(n16444), .IN2(n16445), .Q(g13155) );
  OR2X1 U17521 ( .IN1(n4316), .IN2(g1164), .Q(n16445) );
  AND2X1 U17522 ( .IN1(n16446), .IN2(n16447), .Q(n16444) );
  OR2X1 U17523 ( .IN1(n4300), .IN2(g1165), .Q(n16447) );
  OR2X1 U17524 ( .IN1(n4371), .IN2(g1166), .Q(n16446) );
  AND2X1 U17525 ( .IN1(n16448), .IN2(n16449), .Q(g13149) );
  OR2X1 U17526 ( .IN1(n4372), .IN2(g477), .Q(n16449) );
  AND2X1 U17527 ( .IN1(n16450), .IN2(n16451), .Q(n16448) );
  OR2X1 U17528 ( .IN1(n4313), .IN2(g478), .Q(n16451) );
  OR2X1 U17529 ( .IN1(n4298), .IN2(g479), .Q(n16450) );
  AND2X1 U17530 ( .IN1(n16452), .IN2(n16453), .Q(g13143) );
  OR2X1 U17531 ( .IN1(n4370), .IN2(g2555), .Q(n16453) );
  AND2X1 U17532 ( .IN1(n16454), .IN2(n16455), .Q(n16452) );
  OR2X1 U17533 ( .IN1(n4299), .IN2(g2559), .Q(n16455) );
  OR2X1 U17534 ( .IN1(n4314), .IN2(g2539), .Q(n16454) );
  AND2X1 U17535 ( .IN1(n16456), .IN2(n16457), .Q(g13135) );
  OR2X1 U17536 ( .IN1(n4315), .IN2(g1861), .Q(n16457) );
  AND2X1 U17537 ( .IN1(n16458), .IN2(n16459), .Q(n16456) );
  OR2X1 U17538 ( .IN1(n4366), .IN2(g1865), .Q(n16459) );
  OR2X1 U17539 ( .IN1(n4296), .IN2(g1845), .Q(n16458) );
  AND2X1 U17540 ( .IN1(n16460), .IN2(n16461), .Q(g13124) );
  OR2X1 U17541 ( .IN1(n4316), .IN2(g1167), .Q(n16461) );
  AND2X1 U17542 ( .IN1(n16462), .IN2(n16463), .Q(n16460) );
  OR2X1 U17543 ( .IN1(n4300), .IN2(g1171), .Q(n16463) );
  OR2X1 U17544 ( .IN1(n4371), .IN2(g1151), .Q(n16462) );
  AND2X1 U17545 ( .IN1(n16464), .IN2(n16465), .Q(g13111) );
  OR2X1 U17546 ( .IN1(n4372), .IN2(g480), .Q(n16465) );
  AND2X1 U17547 ( .IN1(n16466), .IN2(n16467), .Q(n16464) );
  OR2X1 U17548 ( .IN1(n4313), .IN2(g484), .Q(n16467) );
  OR2X1 U17549 ( .IN1(n4298), .IN2(g464), .Q(n16466) );
  AND2X1 U17550 ( .IN1(n16468), .IN2(n16469), .Q(g13110) );
  AND2X1 U17551 ( .IN1(n9081), .IN2(n16470), .Q(n16469) );
  AND2X1 U17552 ( .IN1(n4482), .IN2(n8822), .Q(n16470) );
  INVX0 U17553 ( .INP(n16471), .ZN(n16468) );
  OR2X1 U17554 ( .IN1(n16472), .IN2(n16473), .Q(n16471) );
  OR2X1 U17555 ( .IN1(n14847), .IN2(g2917), .Q(n16473) );
  INVX0 U17556 ( .INP(n9552), .ZN(n14847) );
  AND2X1 U17557 ( .IN1(n16474), .IN2(n16475), .Q(n9552) );
  AND2X1 U17558 ( .IN1(n4431), .IN2(n9102), .Q(n16475) );
  AND2X1 U17559 ( .IN1(n4355), .IN2(n16476), .Q(n16474) );
  AND2X1 U17560 ( .IN1(n4291), .IN2(n4305), .Q(n16476) );
  OR2X1 U17561 ( .IN1(n4349), .IN2(n4330), .Q(n16472) );
  XOR2X1 U17562 ( .IN1(n9724), .IN2(n9080), .Q(N995) );
  XOR2X1 U17563 ( .IN1(n16477), .IN2(n16478), .Q(n9724) );
  XOR2X1 U17564 ( .IN1(n16479), .IN2(n16480), .Q(n16478) );
  XOR2X1 U17565 ( .IN1(n16496), .IN2(n9077), .Q(n16480) );
  XOR2X1 U17566 ( .IN1(test_so99), .IN2(n16495), .Q(n16479) );
  XOR2X1 U17567 ( .IN1(n16481), .IN2(n16482), .Q(n16477) );
  XOR2X1 U17568 ( .IN1(n9076), .IN2(n9075), .Q(n16482) );
  XOR2X1 U17569 ( .IN1(DFF_1618_n1), .IN2(n9074), .Q(n16481) );
  XOR2X1 U17570 ( .IN1(n9078), .IN2(n9725), .Q(N690) );
  XNOR2X1 U17571 ( .IN1(n16483), .IN2(n16484), .Q(n9725) );
  XOR2X1 U17572 ( .IN1(n16485), .IN2(n16486), .Q(n16484) );
  XOR2X1 U17573 ( .IN1(n9058), .IN2(n9057), .Q(n16486) );
  XOR2X1 U17574 ( .IN1(n16497), .IN2(n16498), .Q(n16485) );
  XOR2X1 U17575 ( .IN1(n16487), .IN2(n16488), .Q(n16483) );
  XOR2X1 U17576 ( .IN1(n9056), .IN2(n9055), .Q(n16488) );
  XOR2X1 U17577 ( .IN1(DFF_1628_n1), .IN2(n9054), .Q(n16487) );
  OR2X1 U3772_U1 ( .IN1(n2230), .IN2(n2217), .Q(n2231) );
  OR2X1 U3776_U1 ( .IN1(n2374), .IN2(n2361), .Q(n2375) );
  OR2X1 U3777_U1 ( .IN1(g51), .IN2(DFF_2_n1), .Q(n4264) );
  OR2X1 U3778_U1 ( .IN1(n2445), .IN2(n2446), .Q(n2440) );
  OR2X1 U3779_U1 ( .IN1(n484), .IN2(n2446), .Q(n2426) );
  OR2X1 U3780_U1 ( .IN1(n2670), .IN2(n2671), .Q(n2669) );
  OR2X1 U3781_U1 ( .IN1(n2685), .IN2(n2686), .Q(n2684) );
  OR2X1 U3782_U1 ( .IN1(n2718), .IN2(n2719), .Q(n2717) );
  OR2X1 U3783_U1 ( .IN1(n1291), .IN2(g2124), .Q(n2981) );
  OR2X1 U3784_U1 ( .IN1(n1005), .IN2(g1430), .Q(n2984) );
  OR2X1 U3785_U1 ( .IN1(n716), .IN2(g744), .Q(n2987) );
  OR2X1 U3786_U1 ( .IN1(n407), .IN2(g56), .Q(n2990) );
  OR2X1 U3787_U1 ( .IN1(n3742), .IN2(test_so98), .Q(n3741) );
  OR2X1 U3901_U1 ( .IN1(n2302), .IN2(n2289), .Q(n2303) );
  OR2X1 U3902_U1 ( .IN1(n488), .IN2(n2289), .Q(n2275) );
  INVX0 U4467_U2 ( .INP(n3254), .ZN(U4467_n1) );
  AND2X1 U4467_U1 ( .IN1(n1348), .IN2(U4467_n1), .Q(n3252) );
  INVX0 U4904_U2 ( .INP(n2617), .ZN(U4904_n1) );
  AND2X1 U4904_U1 ( .IN1(n2800), .IN2(U4904_n1), .Q(n2798) );
  INVX0 U4930_U2 ( .INP(n2617), .ZN(U4930_n1) );
  AND2X1 U4930_U1 ( .IN1(n2616), .IN2(U4930_n1), .Q(n2594) );
  INVX0 U5128_U2 ( .INP(n4406), .ZN(U5128_n1) );
  AND2X1 U5128_U1 ( .IN1(n3933), .IN2(U5128_n1), .Q(n3940) );
  INVX0 U5141_U2 ( .INP(n4405), .ZN(U5141_n1) );
  AND2X1 U5141_U1 ( .IN1(n3939), .IN2(U5141_n1), .Q(n3936) );
  INVX0 U5749_U2 ( .INP(n1289), .ZN(U5749_n1) );
  AND2X1 U5749_U1 ( .IN1(g2133), .IN2(U5749_n1), .Q(n3159) );
  INVX0 U5750_U2 ( .INP(n1003), .ZN(U5750_n1) );
  AND2X1 U5750_U1 ( .IN1(g1439), .IN2(U5750_n1), .Q(n3163) );
  INVX0 U5751_U2 ( .INP(n714), .ZN(U5751_n1) );
  AND2X1 U5751_U1 ( .IN1(g753), .IN2(U5751_n1), .Q(n3167) );
  INVX0 U5752_U2 ( .INP(n405), .ZN(U5752_n1) );
  AND2X1 U5752_U1 ( .IN1(g65), .IN2(U5752_n1), .Q(n3171) );
  INVX0 U5753_U2 ( .INP(n4522), .ZN(U5753_n1) );
  AND2X1 U5753_U1 ( .IN1(g2142), .IN2(U5753_n1), .Q(n3424) );
  INVX0 U5754_U2 ( .INP(n4526), .ZN(U5754_n1) );
  AND2X1 U5754_U1 ( .IN1(g2151), .IN2(U5754_n1), .Q(n3683) );
  INVX0 U5755_U2 ( .INP(n3888), .ZN(U5755_n1) );
  AND2X1 U5755_U1 ( .IN1(g2160), .IN2(U5755_n1), .Q(n3887) );
  INVX0 U5756_U2 ( .INP(n4523), .ZN(U5756_n1) );
  AND2X1 U5756_U1 ( .IN1(g1448), .IN2(U5756_n1), .Q(n3427) );
  INVX0 U5757_U2 ( .INP(n4527), .ZN(U5757_n1) );
  AND2X1 U5757_U1 ( .IN1(g1457), .IN2(U5757_n1), .Q(n3686) );
  INVX0 U5758_U2 ( .INP(n3891), .ZN(U5758_n1) );
  AND2X1 U5758_U1 ( .IN1(g1466), .IN2(U5758_n1), .Q(n3890) );
  INVX0 U5759_U2 ( .INP(n712), .ZN(U5759_n1) );
  AND2X1 U5759_U1 ( .IN1(g762), .IN2(U5759_n1), .Q(n3430) );
  INVX0 U5760_U2 ( .INP(n710), .ZN(U5760_n1) );
  AND2X1 U5760_U1 ( .IN1(g771), .IN2(U5760_n1), .Q(n3689) );
  INVX0 U5761_U2 ( .INP(n3894), .ZN(U5761_n1) );
  AND2X1 U5761_U1 ( .IN1(g780), .IN2(U5761_n1), .Q(n3893) );
  INVX0 U5762_U2 ( .INP(n4521), .ZN(U5762_n1) );
  AND2X1 U5762_U1 ( .IN1(g74), .IN2(U5762_n1), .Q(n3433) );
  INVX0 U5763_U2 ( .INP(n4528), .ZN(U5763_n1) );
  AND2X1 U5763_U1 ( .IN1(g83), .IN2(U5763_n1), .Q(n3692) );
  INVX0 U5764_U2 ( .INP(n3897), .ZN(U5764_n1) );
  AND2X1 U5764_U1 ( .IN1(g92), .IN2(U5764_n1), .Q(n3896) );
  INVX0 U5882_U2 ( .INP(g3036), .ZN(U5882_n1) );
  AND2X1 U5882_U1 ( .IN1(n4102), .IN2(U5882_n1), .Q(n4101) );
  INVX0 U5939_U2 ( .INP(n1221), .ZN(U5939_n1) );
  AND2X1 U5939_U1 ( .IN1(g2257), .IN2(U5939_n1), .Q(n3038) );
  INVX0 U5940_U2 ( .INP(n932), .ZN(U5940_n1) );
  AND2X1 U5940_U1 ( .IN1(g1563), .IN2(U5940_n1), .Q(n3070) );
  INVX0 U5941_U2 ( .INP(n640), .ZN(U5941_n1) );
  AND2X1 U5941_U1 ( .IN1(g869), .IN2(U5941_n1), .Q(n3102) );
  INVX0 U5942_U2 ( .INP(n338), .ZN(U5942_n1) );
  AND2X1 U5942_U1 ( .IN1(g181), .IN2(U5942_n1), .Q(n3130) );
  INVX0 U6140_U2 ( .INP(n4066), .ZN(U6140_n1) );
  AND2X1 U6140_U1 ( .IN1(g3002), .IN2(U6140_n1), .Q(n4065) );
  INVX0 U6460_U2 ( .INP(g3230), .ZN(U6460_n1) );
  AND2X1 U6460_U1 ( .IN1(g3233), .IN2(U6460_n1), .Q(n3700) );
  INVX0 U6470_U2 ( .INP(n4305), .ZN(U6470_n1) );
  AND2X1 U6470_U1 ( .IN1(g2892), .IN2(U6470_n1), .Q(n4182) );
  INVX0 U6562_U2 ( .INP(g3204), .ZN(U6562_n1) );
  AND2X1 U6562_U1 ( .IN1(n305), .IN2(U6562_n1), .Q(n3939) );
  INVX0 U6563_U2 ( .INP(g3204), .ZN(U6563_n1) );
  AND2X1 U6563_U1 ( .IN1(n4073), .IN2(U6563_n1), .Q(n3705) );
  INVX0 U6718_U2 ( .INP(g3197), .ZN(U6718_n1) );
  AND2X1 U6718_U1 ( .IN1(n306), .IN2(U6718_n1), .Q(n4073) );
  INVX0 U7116_U2 ( .INP(g2903), .ZN(U7116_n1) );
  AND2X1 U7116_U1 ( .IN1(n4058), .IN2(U7116_n1), .Q(n4057) );
  INVX0 U7118_U2 ( .INP(g2896), .ZN(U7118_n1) );
  AND2X1 U7118_U1 ( .IN1(n4123), .IN2(U7118_n1), .Q(n4122) );
  INVX0 U7293_U2 ( .INP(g3234), .ZN(U7293_n1) );
  AND2X1 U7293_U1 ( .IN1(n4598), .IN2(U7293_n1), .Q(g20877) );
endmodule

