module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n1233_, new_n1215_, new_n1105_, new_n1249_, new_n955_, new_n608_, new_n888_, new_n847_, new_n1157_, new_n501_, new_n798_, new_n1180_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n779_, new_n1232_, new_n1025_, new_n566_, new_n641_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n1176_, new_n1207_, new_n1211_, new_n514_, new_n601_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n1125_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n821_, new_n542_, new_n669_, new_n1237_, new_n1172_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n1210_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n1213_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n1188_, new_n344_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n1221_, new_n1167_, new_n1264_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n1238_, new_n792_, new_n1058_, new_n953_, new_n1162_, new_n481_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n1250_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n1151_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1203_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n1083_, new_n655_, new_n759_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n829_, new_n1257_, new_n988_, new_n478_, new_n694_, new_n461_, new_n1228_, new_n710_, new_n971_, new_n565_, new_n361_, new_n764_, new_n906_, new_n683_, new_n1196_, new_n511_, new_n463_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n517_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1216_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n1170_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n420_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n1182_, new_n1200_, new_n650_, new_n708_, new_n750_, new_n1217_, new_n887_, new_n429_, new_n355_, new_n926_, new_n353_, new_n1222_, new_n432_, new_n734_, new_n912_, new_n1062_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1226_, new_n778_, new_n452_, new_n1198_, new_n1219_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n1168_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n1007_, new_n935_, new_n1241_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1159_, new_n1020_, new_n363_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n1133_, new_n398_, new_n1177_, new_n646_, new_n1132_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1026_, new_n1106_, new_n473_, new_n1147_, new_n1229_, new_n790_, new_n1081_, new_n587_, new_n1247_, new_n465_, new_n739_, new_n783_, new_n969_, new_n835_, new_n1234_, new_n996_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n943_, new_n874_, new_n1245_, new_n663_, new_n579_, new_n1209_, new_n347_, new_n659_, new_n1254_, new_n700_, new_n921_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n1218_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n1201_, new_n948_, new_n1231_, new_n762_, new_n1055_, new_n1193_, new_n838_, new_n923_, new_n1187_, new_n469_, new_n1205_, new_n1154_, new_n437_, new_n1085_, new_n1253_, new_n1256_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n1128_, new_n1002_, new_n834_, new_n1169_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n1171_, new_n688_, new_n1255_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1124_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n494_, new_n672_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n1160_, new_n362_, new_n1166_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n1104_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n1175_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1251_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n1095_, new_n1252_, new_n998_, new_n1056_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n963_, new_n586_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n1191_, new_n824_, new_n520_, new_n1001_, new_n717_, new_n403_, new_n475_, new_n868_, new_n1242_, new_n825_, new_n858_, new_n557_, new_n936_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n558_, new_n382_, new_n583_, new_n617_, new_n1080_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n1186_, new_n612_, new_n919_, new_n1015_, new_n755_, new_n1261_, new_n1040_, new_n1246_, new_n922_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n1179_, new_n499_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n1185_, new_n1240_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n1174_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n1195_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n1227_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n1248_, new_n751_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n1244_, new_n1181_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n1072_, new_n769_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n1164_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n732_, new_n687_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n1220_, new_n989_, new_n1204_, new_n1117_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n1096_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n1206_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1008_, new_n640_, new_n684_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n905_, new_n539_, new_n1258_, new_n803_, new_n727_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1173_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1189_, new_n1153_, new_n357_, new_n1197_, new_n780_, new_n984_, new_n643_, new_n474_, new_n1223_, new_n1129_, new_n467_, new_n1013_, new_n1194_, new_n1243_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n1230_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n1165_, new_n1259_, new_n425_, new_n896_, new_n802_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n1236_, new_n709_, new_n373_, new_n866_, new_n1235_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1225_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n889_, new_n536_, new_n464_, new_n1089_, new_n1192_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n343_, N75 );
nand g001 ( new_n344_, N29, N42 );
nor g002 ( new_n345_, new_n344_, new_n343_ );
xor g003 ( N388, new_n345_, keyIn_0_5 );
not g004 ( new_n347_, N80 );
nand g005 ( new_n348_, N29, N36 );
nor g006 ( new_n349_, new_n348_, new_n347_ );
xor g007 ( N389, new_n349_, keyIn_0_6 );
not g008 ( new_n351_, N42 );
nor g009 ( N390, new_n348_, new_n351_ );
nand g010 ( new_n353_, N85, N86 );
xnor g011 ( N391, new_n353_, keyIn_0_11 );
not g012 ( new_n355_, N13 );
nand g013 ( new_n356_, N1, N8 );
nor g014 ( new_n357_, new_n356_, new_n355_ );
nand g015 ( new_n358_, new_n357_, N17 );
xnor g016 ( new_n359_, new_n358_, keyIn_0_0 );
xor g017 ( N418, new_n359_, keyIn_0_40 );
nand g018 ( new_n361_, N1, N26 );
nand g019 ( new_n362_, N13, N17 );
nor g020 ( new_n363_, new_n361_, new_n362_ );
xnor g021 ( new_n364_, new_n363_, keyIn_0_1 );
xnor g022 ( new_n365_, N390, keyIn_0_2 );
nand g023 ( N419, new_n364_, new_n365_ );
nand g024 ( new_n367_, N59, N75 );
nor g025 ( new_n368_, new_n367_, new_n347_ );
xor g026 ( new_n369_, new_n368_, keyIn_0_7 );
xnor g027 ( N420, new_n369_, keyIn_0_46 );
nand g028 ( new_n371_, N36, N59 );
nor g029 ( new_n372_, new_n371_, new_n347_ );
xnor g030 ( new_n373_, new_n372_, keyIn_0_9 );
xnor g031 ( N421, new_n373_, keyIn_0_47 );
nor g032 ( new_n375_, new_n371_, new_n351_ );
xnor g033 ( new_n376_, new_n375_, keyIn_0_10 );
xnor g034 ( N422, new_n376_, keyIn_0_48 );
nor g035 ( new_n378_, N87, N88 );
xor g036 ( new_n379_, new_n378_, keyIn_0_12 );
nand g037 ( new_n380_, new_n379_, N90 );
xnor g038 ( N423, new_n380_, keyIn_0_50 );
not g039 ( new_n382_, new_n365_ );
nor g040 ( new_n383_, new_n382_, keyIn_0_41 );
nand g041 ( new_n384_, new_n382_, keyIn_0_41 );
nand g042 ( new_n385_, new_n384_, new_n364_ );
nor g043 ( new_n386_, new_n385_, new_n383_ );
xnor g044 ( N446, new_n386_, keyIn_0_58 );
not g045 ( new_n388_, N51 );
nor g046 ( new_n389_, new_n361_, new_n388_ );
xor g047 ( new_n390_, new_n389_, keyIn_0_43 );
xnor g048 ( N447, new_n390_, keyIn_0_60 );
nand g049 ( new_n392_, new_n357_, N55 );
nand g050 ( new_n393_, N29, N68 );
nor g051 ( new_n394_, new_n392_, new_n393_ );
xor g052 ( N448, new_n394_, keyIn_0_62 );
not g053 ( new_n396_, new_n392_ );
not g054 ( new_n397_, N74 );
nand g055 ( new_n398_, N59, N68 );
nor g056 ( new_n399_, new_n398_, new_n397_ );
nand g057 ( new_n400_, new_n396_, new_n399_ );
xnor g058 ( new_n401_, new_n400_, keyIn_0_45 );
xnor g059 ( N449, new_n401_, keyIn_0_63 );
nand g060 ( new_n403_, new_n379_, N89 );
xor g061 ( N450, new_n403_, keyIn_0_49 );
not g062 ( new_n405_, N130 );
nor g063 ( new_n406_, N91, N96 );
xnor g064 ( new_n407_, new_n406_, keyIn_0_14 );
nand g065 ( new_n408_, N91, N96 );
xnor g066 ( new_n409_, new_n408_, keyIn_0_13 );
nand g067 ( new_n410_, new_n407_, new_n409_ );
xor g068 ( new_n411_, new_n410_, keyIn_0_51 );
nand g069 ( new_n412_, new_n411_, keyIn_0_64 );
not g070 ( new_n413_, N106 );
nor g071 ( new_n414_, keyIn_0_15, N101 );
nand g072 ( new_n415_, new_n414_, new_n413_ );
nand g073 ( new_n416_, N101, N106 );
not g074 ( new_n417_, new_n416_ );
not g075 ( new_n418_, keyIn_0_15 );
nor g076 ( new_n419_, N101, N106 );
nor g077 ( new_n420_, new_n419_, new_n418_ );
nor g078 ( new_n421_, new_n420_, new_n417_ );
nand g079 ( new_n422_, new_n421_, new_n415_ );
xnor g080 ( new_n423_, new_n422_, keyIn_0_65 );
nor g081 ( new_n424_, new_n411_, keyIn_0_64 );
nor g082 ( new_n425_, new_n424_, new_n423_ );
nand g083 ( new_n426_, new_n425_, new_n412_ );
nor g084 ( new_n427_, new_n426_, keyIn_0_77 );
nand g085 ( new_n428_, new_n426_, keyIn_0_77 );
nand g086 ( new_n429_, new_n411_, new_n422_ );
xor g087 ( new_n430_, new_n429_, keyIn_0_66 );
nand g088 ( new_n431_, new_n428_, new_n430_ );
nor g089 ( new_n432_, new_n431_, new_n427_ );
xor g090 ( new_n433_, new_n432_, keyIn_0_86 );
nor g091 ( new_n434_, new_n433_, new_n405_ );
xnor g092 ( new_n435_, new_n434_, keyIn_0_102 );
nand g093 ( new_n436_, new_n433_, new_n405_ );
xnor g094 ( new_n437_, new_n436_, keyIn_0_103 );
nand g095 ( new_n438_, new_n435_, new_n437_ );
xor g096 ( new_n439_, new_n438_, keyIn_0_122 );
xnor g097 ( new_n440_, new_n439_, keyIn_0_128 );
not g098 ( new_n441_, N135 );
nor g099 ( new_n442_, N111, N116 );
xor g100 ( new_n443_, new_n442_, keyIn_0_17 );
nand g101 ( new_n444_, N111, N116 );
xor g102 ( new_n445_, new_n444_, keyIn_0_16 );
nand g103 ( new_n446_, new_n443_, new_n445_ );
xnor g104 ( new_n447_, new_n446_, keyIn_0_52 );
nand g105 ( new_n448_, new_n447_, keyIn_0_67 );
nor g106 ( new_n449_, new_n447_, keyIn_0_67 );
nor g107 ( new_n450_, keyIn_0_18, N126 );
xor g108 ( new_n451_, new_n450_, keyIn_0_53 );
not g109 ( new_n452_, N121 );
nand g110 ( new_n453_, keyIn_0_18, N126 );
nand g111 ( new_n454_, new_n453_, new_n452_ );
xnor g112 ( new_n455_, new_n451_, new_n454_ );
xnor g113 ( new_n456_, new_n455_, keyIn_0_68 );
nor g114 ( new_n457_, new_n456_, new_n449_ );
nand g115 ( new_n458_, new_n457_, new_n448_ );
nor g116 ( new_n459_, new_n458_, keyIn_0_78 );
nand g117 ( new_n460_, new_n447_, new_n455_ );
xnor g118 ( new_n461_, new_n460_, keyIn_0_69 );
nand g119 ( new_n462_, new_n458_, keyIn_0_78 );
nand g120 ( new_n463_, new_n462_, new_n461_ );
nor g121 ( new_n464_, new_n463_, new_n459_ );
xnor g122 ( new_n465_, new_n464_, keyIn_0_87 );
nand g123 ( new_n466_, new_n465_, new_n441_ );
xnor g124 ( new_n467_, new_n466_, keyIn_0_105 );
nor g125 ( new_n468_, new_n465_, new_n441_ );
xnor g126 ( new_n469_, new_n468_, keyIn_0_104 );
nand g127 ( new_n470_, new_n469_, new_n467_ );
xor g128 ( new_n471_, new_n470_, keyIn_0_123 );
xnor g129 ( new_n472_, new_n471_, keyIn_0_129 );
nor g130 ( new_n473_, new_n440_, new_n472_ );
nand g131 ( new_n474_, new_n473_, keyIn_0_138 );
nor g132 ( new_n475_, new_n439_, new_n471_ );
nor g133 ( new_n476_, new_n473_, keyIn_0_138 );
nor g134 ( new_n477_, new_n476_, new_n475_ );
nand g135 ( new_n478_, new_n477_, new_n474_ );
xor g136 ( N767, new_n478_, keyIn_0_156 );
nor g137 ( new_n480_, N159, N165 );
xnor g138 ( new_n481_, new_n480_, keyIn_0_26 );
nand g139 ( new_n482_, N159, N165 );
xnor g140 ( new_n483_, new_n482_, keyIn_0_25 );
nand g141 ( new_n484_, new_n481_, new_n483_ );
xnor g142 ( new_n485_, new_n484_, keyIn_0_71 );
nor g143 ( new_n486_, N171, N177 );
xor g144 ( new_n487_, new_n486_, keyIn_0_28 );
nand g145 ( new_n488_, N171, N177 );
xor g146 ( new_n489_, new_n488_, keyIn_0_27 );
nand g147 ( new_n490_, new_n487_, new_n489_ );
xnor g148 ( new_n491_, new_n490_, keyIn_0_72 );
nor g149 ( new_n492_, new_n491_, new_n485_ );
xnor g150 ( new_n493_, new_n492_, keyIn_0_84 );
nand g151 ( new_n494_, new_n490_, new_n484_ );
nand g152 ( new_n495_, new_n493_, new_n494_ );
xnor g153 ( new_n496_, new_n495_, keyIn_0_101 );
nor g154 ( new_n497_, new_n496_, N130 );
xnor g155 ( new_n498_, new_n497_, keyIn_0_115 );
nand g156 ( new_n499_, new_n496_, N130 );
xnor g157 ( new_n500_, new_n499_, keyIn_0_114 );
nand g158 ( new_n501_, new_n498_, new_n500_ );
nor g159 ( new_n502_, new_n501_, keyIn_0_136 );
not g160 ( new_n503_, keyIn_0_116 );
not g161 ( new_n504_, N207 );
nor g162 ( new_n505_, N195, N201 );
xnor g163 ( new_n506_, new_n505_, keyIn_0_31 );
nand g164 ( new_n507_, N195, N201 );
xnor g165 ( new_n508_, new_n507_, keyIn_0_30 );
nand g166 ( new_n509_, new_n506_, new_n508_ );
xor g167 ( new_n510_, new_n509_, keyIn_0_57 );
nor g168 ( new_n511_, new_n510_, keyIn_0_73 );
nor g169 ( new_n512_, keyIn_0_29, N189 );
xnor g170 ( new_n513_, new_n512_, keyIn_0_56 );
not g171 ( new_n514_, N183 );
nand g172 ( new_n515_, keyIn_0_29, N189 );
nand g173 ( new_n516_, new_n515_, new_n514_ );
xnor g174 ( new_n517_, new_n513_, new_n516_ );
nand g175 ( new_n518_, new_n510_, keyIn_0_73 );
not g176 ( new_n519_, new_n518_ );
nor g177 ( new_n520_, new_n519_, new_n517_ );
not g178 ( new_n521_, new_n520_ );
nor g179 ( new_n522_, new_n521_, new_n511_ );
not g180 ( new_n523_, new_n522_ );
nor g181 ( new_n524_, new_n523_, keyIn_0_85 );
nand g182 ( new_n525_, new_n523_, keyIn_0_85 );
not g183 ( new_n526_, new_n510_ );
nand g184 ( new_n527_, new_n526_, new_n517_ );
xnor g185 ( new_n528_, new_n527_, keyIn_0_74 );
nand g186 ( new_n529_, new_n525_, new_n528_ );
nor g187 ( new_n530_, new_n529_, new_n524_ );
not g188 ( new_n531_, new_n530_ );
nor g189 ( new_n532_, new_n531_, new_n504_ );
nor g190 ( new_n533_, new_n532_, new_n503_ );
nand g191 ( new_n534_, new_n532_, new_n503_ );
not g192 ( new_n535_, new_n534_ );
nor g193 ( new_n536_, new_n530_, N207 );
nor g194 ( new_n537_, new_n535_, new_n536_ );
not g195 ( new_n538_, new_n537_ );
nor g196 ( new_n539_, new_n538_, new_n533_ );
nand g197 ( new_n540_, new_n501_, keyIn_0_136 );
nand g198 ( new_n541_, new_n539_, new_n540_ );
nor g199 ( new_n542_, new_n541_, new_n502_ );
xnor g200 ( new_n543_, new_n542_, keyIn_0_139 );
not g201 ( new_n544_, new_n539_ );
nand g202 ( new_n545_, new_n544_, new_n501_ );
xnor g203 ( new_n546_, new_n545_, keyIn_0_137 );
nand g204 ( new_n547_, new_n543_, new_n546_ );
xor g205 ( N768, new_n547_, keyIn_0_157 );
not g206 ( new_n549_, keyIn_0_215 );
not g207 ( new_n550_, keyIn_0_192 );
not g208 ( new_n551_, N261 );
not g209 ( new_n552_, keyIn_0_135 );
not g210 ( new_n553_, keyIn_0_127 );
not g211 ( new_n554_, keyIn_0_59 );
not g212 ( new_n555_, keyIn_0_42 );
xnor g213 ( new_n556_, new_n389_, new_n555_ );
xnor g214 ( new_n557_, new_n556_, new_n554_ );
not g215 ( new_n558_, keyIn_0_55 );
nor g216 ( new_n559_, N17, N42 );
xnor g217 ( new_n560_, new_n559_, keyIn_0_23 );
nand g218 ( new_n561_, N17, N42 );
xnor g219 ( new_n562_, new_n561_, keyIn_0_24 );
nor g220 ( new_n563_, new_n560_, new_n562_ );
nor g221 ( new_n564_, new_n563_, new_n558_ );
not g222 ( new_n565_, new_n564_ );
nand g223 ( new_n566_, N59, N156 );
not g224 ( new_n567_, N17 );
nand g225 ( new_n568_, new_n567_, new_n351_ );
nand g226 ( new_n569_, new_n568_, keyIn_0_23 );
not g227 ( new_n570_, keyIn_0_23 );
nand g228 ( new_n571_, new_n559_, new_n570_ );
nand g229 ( new_n572_, new_n569_, new_n571_ );
not g230 ( new_n573_, keyIn_0_24 );
xnor g231 ( new_n574_, new_n561_, new_n573_ );
nand g232 ( new_n575_, new_n572_, new_n574_ );
nor g233 ( new_n576_, new_n575_, keyIn_0_55 );
nor g234 ( new_n577_, new_n576_, new_n566_ );
nand g235 ( new_n578_, new_n577_, new_n565_ );
nor g236 ( new_n579_, new_n578_, new_n557_ );
nand g237 ( new_n580_, new_n579_, keyIn_0_82 );
not g238 ( new_n581_, keyIn_0_82 );
nand g239 ( new_n582_, new_n556_, keyIn_0_59 );
xnor g240 ( new_n583_, new_n389_, keyIn_0_42 );
nand g241 ( new_n584_, new_n583_, new_n554_ );
nand g242 ( new_n585_, new_n582_, new_n584_ );
not g243 ( new_n586_, new_n566_ );
nand g244 ( new_n587_, new_n563_, new_n558_ );
nand g245 ( new_n588_, new_n587_, new_n586_ );
nor g246 ( new_n589_, new_n588_, new_n564_ );
nand g247 ( new_n590_, new_n589_, new_n585_ );
nand g248 ( new_n591_, new_n590_, new_n581_ );
nand g249 ( new_n592_, new_n580_, new_n591_ );
nand g250 ( new_n593_, N17, N51 );
nor g251 ( new_n594_, new_n356_, new_n593_ );
xnor g252 ( new_n595_, new_n594_, keyIn_0_3 );
nand g253 ( new_n596_, N42, N59 );
nor g254 ( new_n597_, new_n596_, new_n343_ );
xnor g255 ( new_n598_, new_n597_, keyIn_0_8 );
nor g256 ( new_n599_, new_n595_, new_n598_ );
xnor g257 ( new_n600_, new_n599_, keyIn_0_70 );
nand g258 ( new_n601_, new_n592_, new_n600_ );
xnor g259 ( new_n602_, new_n601_, keyIn_0_88 );
nand g260 ( new_n603_, new_n602_, N126 );
xnor g261 ( new_n604_, new_n566_, keyIn_0_22 );
nand g262 ( new_n605_, new_n585_, N17 );
nor g263 ( new_n606_, new_n605_, new_n604_ );
nand g264 ( new_n607_, new_n606_, keyIn_0_83 );
not g265 ( new_n608_, new_n607_ );
not g266 ( new_n609_, keyIn_0_83 );
not g267 ( new_n610_, new_n604_ );
not g268 ( new_n611_, new_n605_ );
nand g269 ( new_n612_, new_n611_, new_n610_ );
nand g270 ( new_n613_, new_n612_, new_n609_ );
nand g271 ( new_n614_, new_n613_, N1 );
nor g272 ( new_n615_, new_n614_, new_n608_ );
nand g273 ( new_n616_, new_n615_, keyIn_0_97 );
not g274 ( new_n617_, keyIn_0_97 );
not g275 ( new_n618_, N1 );
nor g276 ( new_n619_, new_n606_, keyIn_0_83 );
nor g277 ( new_n620_, new_n619_, new_n618_ );
nand g278 ( new_n621_, new_n620_, new_n607_ );
nand g279 ( new_n622_, new_n621_, new_n617_ );
nand g280 ( new_n623_, new_n616_, new_n622_ );
nand g281 ( new_n624_, new_n623_, N153 );
nand g282 ( new_n625_, new_n603_, new_n624_ );
nor g283 ( new_n626_, new_n625_, new_n553_ );
nand g284 ( new_n627_, N29, N75 );
not g285 ( new_n628_, new_n627_ );
nand g286 ( new_n629_, new_n628_, N80 );
nand g287 ( new_n630_, new_n585_, N55 );
nor g288 ( new_n631_, new_n630_, new_n629_ );
nand g289 ( new_n632_, new_n631_, keyIn_0_81 );
nor g290 ( new_n633_, new_n631_, keyIn_0_81 );
xor g291 ( new_n634_, keyIn_0_19, N268 );
xnor g292 ( new_n635_, new_n634_, keyIn_0_54 );
nor g293 ( new_n636_, new_n633_, new_n635_ );
nand g294 ( new_n637_, new_n636_, new_n632_ );
nand g295 ( new_n638_, new_n625_, new_n553_ );
nand g296 ( new_n639_, new_n638_, new_n637_ );
nor g297 ( new_n640_, new_n639_, new_n626_ );
nand g298 ( new_n641_, new_n640_, new_n552_ );
not g299 ( new_n642_, new_n626_ );
not g300 ( new_n643_, new_n639_ );
nand g301 ( new_n644_, new_n643_, new_n642_ );
nand g302 ( new_n645_, new_n644_, keyIn_0_135 );
nand g303 ( new_n646_, new_n645_, new_n641_ );
nand g304 ( new_n647_, new_n626_, keyIn_0_135 );
not g305 ( new_n648_, new_n647_ );
nor g306 ( new_n649_, new_n646_, new_n648_ );
nand g307 ( new_n650_, new_n649_, N201 );
xnor g308 ( new_n651_, new_n640_, keyIn_0_135 );
nor g309 ( new_n652_, new_n651_, N201 );
xnor g310 ( new_n653_, new_n652_, keyIn_0_154 );
nand g311 ( new_n654_, new_n653_, new_n650_ );
nor g312 ( new_n655_, new_n654_, new_n551_ );
nand g313 ( new_n656_, new_n655_, new_n550_ );
nor g314 ( new_n657_, new_n655_, new_n550_ );
not g315 ( new_n658_, new_n654_ );
nor g316 ( new_n659_, new_n658_, N261 );
nor g317 ( new_n660_, new_n657_, new_n659_ );
nand g318 ( new_n661_, new_n660_, new_n656_ );
nor g319 ( new_n662_, new_n661_, keyIn_0_209 );
nand g320 ( new_n663_, new_n661_, keyIn_0_209 );
nand g321 ( new_n664_, new_n663_, N219 );
nor g322 ( new_n665_, new_n664_, new_n662_ );
nor g323 ( new_n666_, new_n665_, new_n549_ );
nand g324 ( new_n667_, new_n665_, new_n549_ );
not g325 ( new_n668_, keyIn_0_172 );
not g326 ( new_n669_, N201 );
nand g327 ( new_n670_, new_n651_, new_n647_ );
nor g328 ( new_n671_, new_n670_, new_n669_ );
nand g329 ( new_n672_, new_n671_, new_n668_ );
nand g330 ( new_n673_, new_n650_, keyIn_0_172 );
nand g331 ( new_n674_, new_n672_, new_n673_ );
nand g332 ( new_n675_, new_n674_, N237 );
xnor g333 ( new_n676_, new_n675_, keyIn_0_194 );
not g334 ( new_n677_, N228 );
nor g335 ( new_n678_, new_n654_, new_n677_ );
xnor g336 ( new_n679_, new_n678_, keyIn_0_193 );
nand g337 ( new_n680_, new_n679_, new_n676_ );
xor g338 ( new_n681_, new_n680_, keyIn_0_210 );
not g339 ( new_n682_, keyIn_0_155 );
nand g340 ( new_n683_, new_n649_, N246 );
nand g341 ( new_n684_, new_n683_, new_n682_ );
nand g342 ( new_n685_, N255, N267 );
xnor g343 ( new_n686_, new_n685_, keyIn_0_39 );
nand g344 ( new_n687_, keyIn_0_155, N246 );
nor g345 ( new_n688_, new_n646_, new_n687_ );
nor g346 ( new_n689_, new_n688_, new_n686_ );
nand g347 ( new_n690_, new_n684_, new_n689_ );
nand g348 ( new_n691_, new_n690_, keyIn_0_173 );
nor g349 ( new_n692_, new_n690_, keyIn_0_173 );
nand g350 ( new_n693_, N68, N72 );
nor g351 ( new_n694_, new_n596_, new_n693_ );
xor g352 ( new_n695_, new_n694_, keyIn_0_4 );
nand g353 ( new_n696_, new_n695_, new_n396_ );
xnor g354 ( new_n697_, new_n696_, keyIn_0_44 );
nand g355 ( new_n698_, new_n697_, N73 );
xor g356 ( new_n699_, new_n698_, keyIn_0_61 );
xnor g357 ( new_n700_, new_n699_, keyIn_0_76 );
nand g358 ( new_n701_, new_n700_, N201 );
nand g359 ( new_n702_, N121, N210 );
xor g360 ( new_n703_, new_n702_, keyIn_0_38 );
nand g361 ( new_n704_, new_n701_, new_n703_ );
nor g362 ( new_n705_, new_n692_, new_n704_ );
nand g363 ( new_n706_, new_n705_, new_n691_ );
nor g364 ( new_n707_, new_n681_, new_n706_ );
nand g365 ( new_n708_, new_n707_, new_n667_ );
nor g366 ( new_n709_, new_n708_, new_n666_ );
xnor g367 ( new_n710_, new_n709_, keyIn_0_223 );
xor g368 ( new_n711_, new_n710_, keyIn_0_229 );
xnor g369 ( N850, new_n711_, keyIn_0_234 );
not g370 ( new_n713_, keyIn_0_216 );
not g371 ( new_n714_, keyIn_0_111 );
nand g372 ( new_n715_, new_n602_, N111 );
nor g373 ( new_n716_, new_n715_, new_n714_ );
nand g374 ( new_n717_, new_n623_, N143 );
nand g375 ( new_n718_, new_n715_, new_n714_ );
nand g376 ( new_n719_, new_n718_, new_n717_ );
nor g377 ( new_n720_, new_n719_, new_n716_ );
xor g378 ( new_n721_, new_n720_, keyIn_0_126 );
xor g379 ( new_n722_, new_n637_, keyIn_0_98 );
nand g380 ( new_n723_, new_n721_, new_n722_ );
xor g381 ( new_n724_, new_n723_, keyIn_0_132 );
nand g382 ( new_n725_, new_n724_, N183 );
xnor g383 ( new_n726_, new_n725_, keyIn_0_149 );
not g384 ( new_n727_, new_n724_ );
nand g385 ( new_n728_, new_n727_, new_n514_ );
xnor g386 ( new_n729_, new_n728_, keyIn_0_150 );
not g387 ( new_n730_, new_n729_ );
nor g388 ( new_n731_, new_n730_, new_n726_ );
xnor g389 ( new_n732_, new_n731_, keyIn_0_165 );
not g390 ( new_n733_, new_n732_ );
not g391 ( new_n734_, N189 );
nand g392 ( new_n735_, new_n623_, N146 );
not g393 ( new_n736_, N116 );
not g394 ( new_n737_, keyIn_0_88 );
xnor g395 ( new_n738_, new_n601_, new_n737_ );
nor g396 ( new_n739_, new_n738_, new_n736_ );
xnor g397 ( new_n740_, new_n637_, keyIn_0_99 );
nor g398 ( new_n741_, new_n739_, new_n740_ );
nand g399 ( new_n742_, new_n741_, new_n735_ );
xnor g400 ( new_n743_, new_n742_, keyIn_0_133 );
nand g401 ( new_n744_, new_n743_, new_n734_ );
not g402 ( new_n745_, N195 );
nand g403 ( new_n746_, new_n623_, N149 );
not g404 ( new_n747_, new_n746_ );
nand g405 ( new_n748_, new_n747_, keyIn_0_112 );
not g406 ( new_n749_, keyIn_0_113 );
nand g407 ( new_n750_, new_n749_, N121 );
nor g408 ( new_n751_, new_n738_, new_n750_ );
xor g409 ( new_n752_, new_n637_, keyIn_0_100 );
nor g410 ( new_n753_, new_n751_, new_n752_ );
nand g411 ( new_n754_, new_n748_, new_n753_ );
not g412 ( new_n755_, keyIn_0_112 );
nand g413 ( new_n756_, new_n746_, new_n755_ );
nand g414 ( new_n757_, new_n602_, N121 );
nand g415 ( new_n758_, new_n757_, keyIn_0_113 );
nand g416 ( new_n759_, new_n758_, new_n756_ );
nor g417 ( new_n760_, new_n754_, new_n759_ );
xnor g418 ( new_n761_, new_n760_, keyIn_0_134 );
nand g419 ( new_n762_, new_n761_, new_n745_ );
xnor g420 ( new_n763_, new_n762_, keyIn_0_152 );
not g421 ( new_n764_, new_n763_ );
nand g422 ( new_n765_, new_n653_, N261 );
nor g423 ( new_n766_, new_n765_, new_n764_ );
nand g424 ( new_n767_, new_n766_, new_n744_ );
xnor g425 ( new_n768_, new_n767_, keyIn_0_176 );
xnor g426 ( new_n769_, new_n650_, new_n668_ );
nor g427 ( new_n770_, new_n769_, new_n764_ );
nand g428 ( new_n771_, new_n770_, new_n744_ );
nor g429 ( new_n772_, new_n771_, keyIn_0_197 );
not g430 ( new_n773_, new_n772_ );
not g431 ( new_n774_, keyIn_0_197 );
not g432 ( new_n775_, new_n744_ );
nand g433 ( new_n776_, new_n674_, new_n763_ );
nor g434 ( new_n777_, new_n776_, new_n775_ );
nor g435 ( new_n778_, new_n777_, new_n774_ );
nor g436 ( new_n779_, new_n761_, new_n745_ );
nand g437 ( new_n780_, new_n779_, keyIn_0_169 );
not g438 ( new_n781_, keyIn_0_169 );
not g439 ( new_n782_, keyIn_0_134 );
xnor g440 ( new_n783_, new_n760_, new_n782_ );
nand g441 ( new_n784_, new_n783_, N195 );
nand g442 ( new_n785_, new_n784_, new_n781_ );
nand g443 ( new_n786_, new_n780_, new_n785_ );
nand g444 ( new_n787_, new_n786_, new_n744_ );
xnor g445 ( new_n788_, new_n787_, keyIn_0_196 );
nor g446 ( new_n789_, new_n743_, new_n734_ );
not g447 ( new_n790_, new_n789_ );
nand g448 ( new_n791_, new_n788_, new_n790_ );
nor g449 ( new_n792_, new_n778_, new_n791_ );
nand g450 ( new_n793_, new_n792_, new_n773_ );
nor g451 ( new_n794_, new_n793_, new_n768_ );
nand g452 ( new_n795_, new_n794_, keyIn_0_204 );
not g453 ( new_n796_, keyIn_0_204 );
not g454 ( new_n797_, keyIn_0_176 );
xnor g455 ( new_n798_, new_n767_, new_n797_ );
nand g456 ( new_n799_, new_n771_, keyIn_0_197 );
not g457 ( new_n800_, keyIn_0_196 );
xnor g458 ( new_n801_, new_n787_, new_n800_ );
nor g459 ( new_n802_, new_n801_, new_n789_ );
nand g460 ( new_n803_, new_n799_, new_n802_ );
nor g461 ( new_n804_, new_n803_, new_n772_ );
nand g462 ( new_n805_, new_n804_, new_n798_ );
nand g463 ( new_n806_, new_n805_, new_n796_ );
nand g464 ( new_n807_, new_n795_, new_n806_ );
nor g465 ( new_n808_, new_n733_, new_n807_ );
nor g466 ( new_n809_, new_n808_, keyIn_0_211 );
nand g467 ( new_n810_, new_n733_, new_n807_ );
nand g468 ( new_n811_, new_n808_, keyIn_0_211 );
nand g469 ( new_n812_, new_n811_, new_n810_ );
nor g470 ( new_n813_, new_n812_, new_n809_ );
nand g471 ( new_n814_, new_n813_, new_n713_ );
not g472 ( new_n815_, N219 );
nor g473 ( new_n816_, new_n813_, new_n713_ );
nor g474 ( new_n817_, new_n816_, new_n815_ );
nand g475 ( new_n818_, new_n817_, new_n814_ );
xor g476 ( new_n819_, new_n818_, keyIn_0_220 );
nand g477 ( new_n820_, N106, N210 );
xor g478 ( new_n821_, new_n820_, keyIn_0_34 );
nand g479 ( new_n822_, new_n819_, new_n821_ );
nor g480 ( new_n823_, new_n822_, keyIn_0_226 );
nand g481 ( new_n824_, new_n822_, keyIn_0_226 );
nand g482 ( new_n825_, new_n733_, N228 );
nand g483 ( new_n826_, new_n726_, N237 );
xnor g484 ( new_n827_, new_n826_, keyIn_0_186 );
nand g485 ( new_n828_, new_n825_, new_n827_ );
nor g486 ( new_n829_, new_n828_, keyIn_0_205 );
nand g487 ( new_n830_, new_n828_, keyIn_0_205 );
nand g488 ( new_n831_, new_n724_, N246 );
nand g489 ( new_n832_, new_n700_, N183 );
xnor g490 ( new_n833_, new_n832_, keyIn_0_121 );
nand g491 ( new_n834_, new_n831_, new_n833_ );
xnor g492 ( new_n835_, new_n834_, keyIn_0_166 );
nand g493 ( new_n836_, new_n830_, new_n835_ );
nor g494 ( new_n837_, new_n836_, new_n829_ );
nand g495 ( new_n838_, new_n824_, new_n837_ );
nor g496 ( new_n839_, new_n838_, new_n823_ );
xnor g497 ( new_n840_, new_n839_, keyIn_0_233 );
xnor g498 ( new_n841_, new_n840_, keyIn_0_238 );
xor g499 ( N863, new_n841_, keyIn_0_245 );
not g500 ( new_n843_, keyIn_0_212 );
xor g501 ( new_n844_, new_n766_, keyIn_0_175 );
not g502 ( new_n845_, keyIn_0_195 );
nor g503 ( new_n846_, new_n776_, new_n845_ );
xor g504 ( new_n847_, new_n786_, keyIn_0_189 );
nand g505 ( new_n848_, new_n776_, new_n845_ );
nand g506 ( new_n849_, new_n848_, new_n847_ );
nor g507 ( new_n850_, new_n849_, new_n846_ );
nand g508 ( new_n851_, new_n844_, new_n850_ );
xnor g509 ( new_n852_, new_n851_, keyIn_0_206 );
nand g510 ( new_n853_, new_n790_, new_n744_ );
xnor g511 ( new_n854_, new_n853_, keyIn_0_167 );
nand g512 ( new_n855_, new_n852_, new_n854_ );
nor g513 ( new_n856_, new_n855_, new_n843_ );
nand g514 ( new_n857_, new_n855_, new_n843_ );
nor g515 ( new_n858_, new_n852_, new_n854_ );
nor g516 ( new_n859_, new_n858_, new_n815_ );
nand g517 ( new_n860_, new_n859_, new_n857_ );
nor g518 ( new_n861_, new_n860_, new_n856_ );
nor g519 ( new_n862_, new_n861_, keyIn_0_221 );
nand g520 ( new_n863_, new_n861_, keyIn_0_221 );
nand g521 ( new_n864_, N111, N210 );
xor g522 ( new_n865_, new_n864_, keyIn_0_35 );
nand g523 ( new_n866_, new_n863_, new_n865_ );
nor g524 ( new_n867_, new_n866_, new_n862_ );
xor g525 ( new_n868_, new_n867_, keyIn_0_227 );
nand g526 ( new_n869_, new_n854_, N228 );
xor g527 ( new_n870_, new_n869_, keyIn_0_187 );
not g528 ( new_n871_, keyIn_0_151 );
not g529 ( new_n872_, N246 );
nor g530 ( new_n873_, new_n743_, new_n872_ );
not g531 ( new_n874_, new_n873_ );
nand g532 ( new_n875_, new_n874_, new_n871_ );
not g533 ( new_n876_, new_n875_ );
nand g534 ( new_n877_, new_n873_, keyIn_0_151 );
nand g535 ( new_n878_, N255, N259 );
xnor g536 ( new_n879_, new_n878_, keyIn_0_36 );
nand g537 ( new_n880_, new_n877_, new_n879_ );
nor g538 ( new_n881_, new_n876_, new_n880_ );
nand g539 ( new_n882_, new_n881_, keyIn_0_168 );
nor g540 ( new_n883_, new_n881_, keyIn_0_168 );
not g541 ( new_n884_, N237 );
nor g542 ( new_n885_, new_n790_, new_n884_ );
nand g543 ( new_n886_, new_n885_, keyIn_0_188 );
not g544 ( new_n887_, new_n700_ );
nor g545 ( new_n888_, new_n887_, new_n734_ );
nor g546 ( new_n889_, new_n885_, keyIn_0_188 );
nor g547 ( new_n890_, new_n889_, new_n888_ );
nand g548 ( new_n891_, new_n890_, new_n886_ );
nor g549 ( new_n892_, new_n891_, new_n883_ );
nand g550 ( new_n893_, new_n892_, new_n882_ );
nor g551 ( new_n894_, new_n870_, new_n893_ );
nand g552 ( new_n895_, new_n868_, new_n894_ );
xnor g553 ( new_n896_, new_n895_, keyIn_0_239 );
xor g554 ( N864, new_n896_, keyIn_0_246 );
not g555 ( new_n898_, keyIn_0_228 );
nand g556 ( new_n899_, new_n763_, new_n784_ );
xor g557 ( new_n900_, new_n899_, keyIn_0_170 );
not g558 ( new_n901_, new_n900_ );
nor g559 ( new_n902_, new_n765_, keyIn_0_174 );
nand g560 ( new_n903_, new_n765_, keyIn_0_174 );
nand g561 ( new_n904_, new_n903_, new_n769_ );
nor g562 ( new_n905_, new_n904_, new_n902_ );
xnor g563 ( new_n906_, new_n905_, keyIn_0_207 );
nor g564 ( new_n907_, new_n906_, new_n901_ );
xor g565 ( new_n908_, new_n907_, keyIn_0_213 );
nand g566 ( new_n909_, new_n906_, new_n901_ );
xnor g567 ( new_n910_, new_n909_, keyIn_0_214 );
nor g568 ( new_n911_, new_n908_, new_n910_ );
nor g569 ( new_n912_, new_n911_, keyIn_0_217 );
nand g570 ( new_n913_, new_n911_, keyIn_0_217 );
nand g571 ( new_n914_, new_n913_, N219 );
nor g572 ( new_n915_, new_n914_, new_n912_ );
nand g573 ( new_n916_, new_n915_, keyIn_0_222 );
nand g574 ( new_n917_, N116, N210 );
not g575 ( new_n918_, new_n917_ );
nor g576 ( new_n919_, new_n915_, keyIn_0_222 );
nor g577 ( new_n920_, new_n919_, new_n918_ );
nand g578 ( new_n921_, new_n920_, new_n916_ );
nor g579 ( new_n922_, new_n921_, new_n898_ );
nand g580 ( new_n923_, new_n921_, new_n898_ );
nand g581 ( new_n924_, new_n901_, N228 );
nor g582 ( new_n925_, new_n924_, keyIn_0_190 );
nand g583 ( new_n926_, new_n786_, N237 );
xnor g584 ( new_n927_, new_n926_, keyIn_0_191 );
nand g585 ( new_n928_, new_n924_, keyIn_0_190 );
nand g586 ( new_n929_, new_n928_, new_n927_ );
nor g587 ( new_n930_, new_n929_, new_n925_ );
nor g588 ( new_n931_, new_n930_, keyIn_0_208 );
nand g589 ( new_n932_, new_n930_, keyIn_0_208 );
not g590 ( new_n933_, keyIn_0_153 );
nand g591 ( new_n934_, new_n783_, N246 );
nand g592 ( new_n935_, new_n934_, new_n933_ );
nor g593 ( new_n936_, new_n934_, new_n933_ );
nand g594 ( new_n937_, N255, N260 );
xnor g595 ( new_n938_, new_n937_, keyIn_0_37 );
nor g596 ( new_n939_, new_n936_, new_n938_ );
nand g597 ( new_n940_, new_n939_, new_n935_ );
nor g598 ( new_n941_, new_n940_, keyIn_0_171 );
nand g599 ( new_n942_, new_n700_, N195 );
nand g600 ( new_n943_, new_n940_, keyIn_0_171 );
nand g601 ( new_n944_, new_n943_, new_n942_ );
nor g602 ( new_n945_, new_n944_, new_n941_ );
nand g603 ( new_n946_, new_n932_, new_n945_ );
nor g604 ( new_n947_, new_n946_, new_n931_ );
nand g605 ( new_n948_, new_n923_, new_n947_ );
nor g606 ( new_n949_, new_n948_, new_n922_ );
xnor g607 ( new_n950_, new_n949_, keyIn_0_240 );
xnor g608 ( N865, new_n950_, keyIn_0_247 );
not g609 ( new_n952_, keyIn_0_235 );
not g610 ( new_n953_, keyIn_0_225 );
nor g611 ( new_n954_, new_n630_, new_n604_ );
xnor g612 ( new_n955_, new_n954_, keyIn_0_79 );
nand g613 ( new_n956_, new_n955_, N146 );
xnor g614 ( new_n957_, new_n956_, keyIn_0_91 );
not g615 ( new_n958_, keyIn_0_80 );
nor g616 ( new_n959_, new_n605_, new_n629_ );
nand g617 ( new_n960_, new_n959_, new_n958_ );
nor g618 ( new_n961_, new_n959_, new_n958_ );
nor g619 ( new_n962_, new_n961_, new_n634_ );
nand g620 ( new_n963_, new_n962_, new_n960_ );
xor g621 ( new_n964_, new_n963_, keyIn_0_92 );
nand g622 ( new_n965_, new_n964_, new_n957_ );
xnor g623 ( new_n966_, new_n965_, keyIn_0_107 );
nand g624 ( new_n967_, new_n602_, N96 );
nor g625 ( new_n968_, new_n967_, keyIn_0_106 );
nand g626 ( new_n969_, N51, N138 );
xnor g627 ( new_n970_, new_n969_, keyIn_0_20 );
nand g628 ( new_n971_, new_n967_, keyIn_0_106 );
nand g629 ( new_n972_, new_n971_, new_n970_ );
nor g630 ( new_n973_, new_n972_, new_n968_ );
nand g631 ( new_n974_, new_n966_, new_n973_ );
xnor g632 ( new_n975_, new_n974_, keyIn_0_130 );
nor g633 ( new_n976_, new_n975_, N165 );
xnor g634 ( new_n977_, new_n976_, keyIn_0_144 );
not g635 ( new_n978_, new_n977_ );
not g636 ( new_n979_, N171 );
nand g637 ( new_n980_, new_n602_, N101 );
nand g638 ( new_n981_, N17, N138 );
xor g639 ( new_n982_, new_n981_, keyIn_0_21 );
nand g640 ( new_n983_, new_n980_, new_n982_ );
xnor g641 ( new_n984_, new_n983_, keyIn_0_124 );
nand g642 ( new_n985_, new_n955_, N149 );
xor g643 ( new_n986_, new_n985_, keyIn_0_93 );
xnor g644 ( new_n987_, new_n963_, keyIn_0_94 );
nor g645 ( new_n988_, new_n986_, new_n987_ );
xnor g646 ( new_n989_, new_n988_, keyIn_0_108 );
nand g647 ( new_n990_, new_n989_, new_n984_ );
xnor g648 ( new_n991_, new_n990_, keyIn_0_131 );
nand g649 ( new_n992_, new_n991_, new_n979_ );
xnor g650 ( new_n993_, new_n992_, keyIn_0_145 );
not g651 ( new_n994_, new_n993_ );
nor g652 ( new_n995_, new_n994_, new_n978_ );
not g653 ( new_n996_, new_n995_ );
nand g654 ( new_n997_, new_n807_, new_n729_ );
xnor g655 ( new_n998_, new_n726_, keyIn_0_185 );
nand g656 ( new_n999_, new_n997_, new_n998_ );
nand g657 ( new_n1000_, new_n602_, N106 );
nor g658 ( new_n1001_, new_n1000_, keyIn_0_109 );
nand g659 ( new_n1002_, N138, N152 );
nand g660 ( new_n1003_, new_n1000_, keyIn_0_109 );
nand g661 ( new_n1004_, new_n1003_, new_n1002_ );
nor g662 ( new_n1005_, new_n1004_, new_n1001_ );
nand g663 ( new_n1006_, new_n1005_, keyIn_0_125 );
nor g664 ( new_n1007_, new_n1005_, keyIn_0_125 );
nand g665 ( new_n1008_, new_n955_, N153 );
xnor g666 ( new_n1009_, new_n1008_, keyIn_0_95 );
xnor g667 ( new_n1010_, new_n963_, keyIn_0_96 );
nand g668 ( new_n1011_, new_n1009_, new_n1010_ );
xor g669 ( new_n1012_, new_n1011_, keyIn_0_110 );
nor g670 ( new_n1013_, new_n1007_, new_n1012_ );
nand g671 ( new_n1014_, new_n1013_, new_n1006_ );
nor g672 ( new_n1015_, new_n1014_, N177 );
xor g673 ( new_n1016_, new_n1015_, keyIn_0_147 );
nand g674 ( new_n1017_, new_n999_, new_n1016_ );
nor g675 ( new_n1018_, new_n1017_, new_n996_ );
nand g676 ( new_n1019_, new_n1018_, new_n953_ );
nor g677 ( new_n1020_, new_n1018_, new_n953_ );
not g678 ( new_n1021_, keyIn_0_200 );
nand g679 ( new_n1022_, new_n1014_, N177 );
xor g680 ( new_n1023_, new_n1022_, keyIn_0_146 );
xor g681 ( new_n1024_, new_n1023_, keyIn_0_162 );
not g682 ( new_n1025_, new_n1024_ );
nor g683 ( new_n1026_, new_n1025_, new_n996_ );
nor g684 ( new_n1027_, new_n1026_, new_n1021_ );
nand g685 ( new_n1028_, new_n1026_, new_n1021_ );
nor g686 ( new_n1029_, new_n991_, new_n979_ );
not g687 ( new_n1030_, new_n1029_ );
nor g688 ( new_n1031_, new_n978_, new_n1030_ );
not g689 ( new_n1032_, new_n1031_ );
nor g690 ( new_n1033_, new_n1032_, keyIn_0_199 );
nand g691 ( new_n1034_, new_n1032_, keyIn_0_199 );
nand g692 ( new_n1035_, new_n975_, N165 );
xnor g693 ( new_n1036_, new_n1035_, keyIn_0_143 );
xnor g694 ( new_n1037_, new_n1036_, keyIn_0_179 );
nand g695 ( new_n1038_, new_n1034_, new_n1037_ );
nor g696 ( new_n1039_, new_n1038_, new_n1033_ );
nand g697 ( new_n1040_, new_n1028_, new_n1039_ );
nor g698 ( new_n1041_, new_n1040_, new_n1027_ );
not g699 ( new_n1042_, new_n1041_ );
nor g700 ( new_n1043_, new_n1020_, new_n1042_ );
nand g701 ( new_n1044_, new_n1043_, new_n1019_ );
not g702 ( new_n1045_, N159 );
nand g703 ( new_n1046_, new_n602_, N91 );
xor g704 ( new_n1047_, new_n963_, keyIn_0_90 );
not g705 ( new_n1048_, keyIn_0_89 );
nand g706 ( new_n1049_, new_n955_, N143 );
not g707 ( new_n1050_, new_n1049_ );
nor g708 ( new_n1051_, new_n1050_, new_n1048_ );
nand g709 ( new_n1052_, N8, N138 );
not g710 ( new_n1053_, new_n1052_ );
nor g711 ( new_n1054_, new_n1049_, keyIn_0_89 );
nor g712 ( new_n1055_, new_n1054_, new_n1053_ );
not g713 ( new_n1056_, new_n1055_ );
nor g714 ( new_n1057_, new_n1056_, new_n1051_ );
not g715 ( new_n1058_, new_n1057_ );
nor g716 ( new_n1059_, new_n1058_, new_n1047_ );
nand g717 ( new_n1060_, new_n1059_, new_n1046_ );
not g718 ( new_n1061_, new_n1060_ );
nand g719 ( new_n1062_, new_n1061_, new_n1045_ );
xor g720 ( new_n1063_, new_n1062_, keyIn_0_141 );
nand g721 ( new_n1064_, new_n1044_, new_n1063_ );
nor g722 ( new_n1065_, new_n1064_, new_n952_ );
nand g723 ( new_n1066_, new_n1064_, new_n952_ );
nand g724 ( new_n1067_, new_n1060_, N159 );
xor g725 ( new_n1068_, new_n1067_, keyIn_0_140 );
xnor g726 ( new_n1069_, new_n1068_, keyIn_0_177 );
nand g727 ( new_n1070_, new_n1066_, new_n1069_ );
nor g728 ( new_n1071_, new_n1070_, new_n1065_ );
xnor g729 ( new_n1072_, new_n1071_, keyIn_0_241 );
xnor g730 ( N866, new_n1072_, keyIn_0_248 );
not g731 ( new_n1074_, new_n1016_ );
nor g732 ( new_n1075_, new_n1074_, new_n1023_ );
xor g733 ( new_n1076_, new_n1075_, keyIn_0_163 );
not g734 ( new_n1077_, new_n1076_ );
nand g735 ( new_n1078_, new_n999_, new_n1077_ );
xor g736 ( new_n1079_, new_n1078_, keyIn_0_219 );
not g737 ( new_n1080_, keyIn_0_218 );
not g738 ( new_n1081_, new_n999_ );
nand g739 ( new_n1082_, new_n1081_, new_n1076_ );
nor g740 ( new_n1083_, new_n1082_, new_n1080_ );
nand g741 ( new_n1084_, new_n1082_, new_n1080_ );
nand g742 ( new_n1085_, new_n1084_, N219 );
nor g743 ( new_n1086_, new_n1085_, new_n1083_ );
nand g744 ( new_n1087_, new_n1086_, new_n1079_ );
not g745 ( new_n1088_, keyIn_0_184 );
nand g746 ( new_n1089_, new_n1077_, N228 );
nor g747 ( new_n1090_, new_n1089_, new_n1088_ );
nand g748 ( new_n1091_, new_n1089_, new_n1088_ );
nor g749 ( new_n1092_, new_n1025_, new_n884_ );
not g750 ( new_n1093_, keyIn_0_148 );
nand g751 ( new_n1094_, new_n1014_, N246 );
nor g752 ( new_n1095_, new_n1094_, new_n1093_ );
nand g753 ( new_n1096_, new_n1094_, new_n1093_ );
nand g754 ( new_n1097_, new_n700_, N177 );
xnor g755 ( new_n1098_, new_n1097_, keyIn_0_120 );
nand g756 ( new_n1099_, new_n1096_, new_n1098_ );
nor g757 ( new_n1100_, new_n1099_, new_n1095_ );
nand g758 ( new_n1101_, new_n1100_, keyIn_0_164 );
nor g759 ( new_n1102_, new_n1100_, keyIn_0_164 );
nand g760 ( new_n1103_, N101, N210 );
not g761 ( new_n1104_, new_n1103_ );
nor g762 ( new_n1105_, new_n1102_, new_n1104_ );
nand g763 ( new_n1106_, new_n1105_, new_n1101_ );
nor g764 ( new_n1107_, new_n1092_, new_n1106_ );
nand g765 ( new_n1108_, new_n1091_, new_n1107_ );
nor g766 ( new_n1109_, new_n1108_, new_n1090_ );
nand g767 ( new_n1110_, new_n1087_, new_n1109_ );
xnor g768 ( new_n1111_, new_n1110_, keyIn_0_244 );
xnor g769 ( N874, new_n1111_, keyIn_0_253 );
not g770 ( new_n1113_, keyIn_0_249 );
not g771 ( new_n1114_, new_n1063_ );
not g772 ( new_n1115_, new_n1068_ );
nor g773 ( new_n1116_, new_n1114_, new_n1115_ );
xor g774 ( new_n1117_, new_n1116_, keyIn_0_158 );
not g775 ( new_n1118_, new_n1117_ );
nand g776 ( new_n1119_, new_n1044_, new_n1118_ );
nand g777 ( new_n1120_, new_n1119_, keyIn_0_230 );
not g778 ( new_n1121_, keyIn_0_230 );
not g779 ( new_n1122_, new_n1019_ );
not g780 ( new_n1123_, new_n1017_ );
nand g781 ( new_n1124_, new_n1123_, new_n995_ );
nand g782 ( new_n1125_, new_n1124_, keyIn_0_225 );
nand g783 ( new_n1126_, new_n1125_, new_n1041_ );
nor g784 ( new_n1127_, new_n1126_, new_n1122_ );
nor g785 ( new_n1128_, new_n1127_, new_n1117_ );
nand g786 ( new_n1129_, new_n1128_, new_n1121_ );
nand g787 ( new_n1130_, new_n1129_, new_n1120_ );
nor g788 ( new_n1131_, new_n1044_, new_n1118_ );
not g789 ( new_n1132_, new_n1131_ );
nand g790 ( new_n1133_, new_n1130_, new_n1132_ );
nor g791 ( new_n1134_, new_n1133_, keyIn_0_236 );
nand g792 ( new_n1135_, new_n1133_, keyIn_0_236 );
nand g793 ( new_n1136_, new_n1135_, N219 );
nor g794 ( new_n1137_, new_n1136_, new_n1134_ );
not g795 ( new_n1138_, N210 );
not g796 ( new_n1139_, new_n635_ );
nor g797 ( new_n1140_, new_n1139_, new_n1138_ );
xor g798 ( new_n1141_, new_n1140_, keyIn_0_75 );
not g799 ( new_n1142_, new_n1141_ );
nor g800 ( new_n1143_, new_n1137_, new_n1142_ );
xnor g801 ( new_n1144_, new_n1143_, new_n1113_ );
not g802 ( new_n1145_, keyIn_0_201 );
nor g803 ( new_n1146_, new_n1117_, new_n677_ );
not g804 ( new_n1147_, new_n1146_ );
nand g805 ( new_n1148_, new_n1147_, keyIn_0_178 );
nor g806 ( new_n1149_, new_n1147_, keyIn_0_178 );
nor g807 ( new_n1150_, new_n1068_, new_n884_ );
nor g808 ( new_n1151_, new_n1149_, new_n1150_ );
nand g809 ( new_n1152_, new_n1151_, new_n1148_ );
nor g810 ( new_n1153_, new_n1152_, new_n1145_ );
nand g811 ( new_n1154_, new_n1152_, new_n1145_ );
not g812 ( new_n1155_, keyIn_0_142 );
nand g813 ( new_n1156_, new_n1060_, N246 );
nor g814 ( new_n1157_, new_n1156_, new_n1155_ );
nand g815 ( new_n1158_, new_n700_, N159 );
xnor g816 ( new_n1159_, new_n1158_, keyIn_0_117 );
nand g817 ( new_n1160_, new_n1156_, new_n1155_ );
nand g818 ( new_n1161_, new_n1160_, new_n1159_ );
nor g819 ( new_n1162_, new_n1161_, new_n1157_ );
nand g820 ( new_n1163_, new_n1154_, new_n1162_ );
nor g821 ( new_n1164_, new_n1163_, new_n1153_ );
not g822 ( new_n1165_, new_n1164_ );
nor g823 ( new_n1166_, new_n1144_, new_n1165_ );
nand g824 ( new_n1167_, new_n1166_, keyIn_0_251 );
not g825 ( new_n1168_, keyIn_0_251 );
not g826 ( new_n1169_, new_n1134_ );
not g827 ( new_n1170_, new_n1136_ );
nand g828 ( new_n1171_, new_n1170_, new_n1169_ );
nand g829 ( new_n1172_, new_n1171_, new_n1141_ );
nand g830 ( new_n1173_, new_n1172_, new_n1113_ );
nand g831 ( new_n1174_, new_n1143_, keyIn_0_249 );
nand g832 ( new_n1175_, new_n1173_, new_n1174_ );
nand g833 ( new_n1176_, new_n1175_, new_n1164_ );
nand g834 ( new_n1177_, new_n1176_, new_n1168_ );
nand g835 ( new_n1178_, new_n1167_, new_n1177_ );
nand g836 ( new_n1179_, new_n1178_, keyIn_0_254 );
not g837 ( new_n1180_, keyIn_0_254 );
xnor g838 ( new_n1181_, new_n1176_, keyIn_0_251 );
nand g839 ( new_n1182_, new_n1181_, new_n1180_ );
nand g840 ( N878, new_n1182_, new_n1179_ );
nor g841 ( new_n1184_, new_n1017_, new_n994_ );
nor g842 ( new_n1185_, new_n1184_, keyIn_0_224 );
nand g843 ( new_n1186_, new_n1184_, keyIn_0_224 );
nand g844 ( new_n1187_, new_n1024_, new_n993_ );
nor g845 ( new_n1188_, new_n1187_, keyIn_0_198 );
xor g846 ( new_n1189_, new_n1029_, keyIn_0_181 );
nand g847 ( new_n1190_, new_n1187_, keyIn_0_198 );
nand g848 ( new_n1191_, new_n1190_, new_n1189_ );
nor g849 ( new_n1192_, new_n1191_, new_n1188_ );
nand g850 ( new_n1193_, new_n1186_, new_n1192_ );
nor g851 ( new_n1194_, new_n1193_, new_n1185_ );
nor g852 ( new_n1195_, new_n978_, new_n1036_ );
xnor g853 ( new_n1196_, new_n1195_, keyIn_0_159 );
nand g854 ( new_n1197_, new_n1194_, new_n1196_ );
nor g855 ( new_n1198_, new_n1194_, new_n1196_ );
nor g856 ( new_n1199_, new_n1198_, new_n815_ );
nand g857 ( new_n1200_, new_n1199_, new_n1197_ );
xnor g858 ( new_n1201_, new_n1200_, keyIn_0_242 );
nand g859 ( new_n1202_, N91, N210 );
xor g860 ( new_n1203_, new_n1202_, keyIn_0_32 );
nand g861 ( new_n1204_, new_n1201_, new_n1203_ );
xor g862 ( new_n1205_, new_n1204_, keyIn_0_250 );
not g863 ( new_n1206_, keyIn_0_180 );
not g864 ( new_n1207_, new_n1196_ );
nand g865 ( new_n1208_, new_n1207_, N228 );
nor g866 ( new_n1209_, new_n1208_, new_n1206_ );
nand g867 ( new_n1210_, new_n1036_, N237 );
nand g868 ( new_n1211_, new_n1208_, new_n1206_ );
nand g869 ( new_n1212_, new_n1211_, new_n1210_ );
nor g870 ( new_n1213_, new_n1212_, new_n1209_ );
nor g871 ( new_n1214_, new_n1213_, keyIn_0_202 );
nand g872 ( new_n1215_, new_n1213_, keyIn_0_202 );
not g873 ( new_n1216_, new_n975_ );
nor g874 ( new_n1217_, new_n1216_, new_n872_ );
nand g875 ( new_n1218_, new_n700_, N165 );
xor g876 ( new_n1219_, new_n1218_, keyIn_0_118 );
nor g877 ( new_n1220_, new_n1217_, new_n1219_ );
nand g878 ( new_n1221_, new_n1215_, new_n1220_ );
nor g879 ( new_n1222_, new_n1221_, new_n1214_ );
nand g880 ( new_n1223_, new_n1205_, new_n1222_ );
xor g881 ( N879, new_n1223_, keyIn_0_255 );
nand g882 ( new_n1225_, new_n993_, new_n1030_ );
xor g883 ( new_n1226_, new_n1225_, keyIn_0_160 );
xnor g884 ( new_n1227_, new_n1024_, keyIn_0_183 );
nand g885 ( new_n1228_, new_n1017_, new_n1227_ );
nor g886 ( new_n1229_, new_n1228_, new_n1226_ );
xnor g887 ( new_n1230_, new_n1229_, keyIn_0_231 );
nand g888 ( new_n1231_, new_n1228_, new_n1226_ );
xnor g889 ( new_n1232_, new_n1231_, keyIn_0_232 );
nor g890 ( new_n1233_, new_n1230_, new_n1232_ );
nand g891 ( new_n1234_, new_n1233_, keyIn_0_237 );
nor g892 ( new_n1235_, new_n1233_, keyIn_0_237 );
nor g893 ( new_n1236_, new_n1235_, new_n815_ );
nand g894 ( new_n1237_, new_n1236_, new_n1234_ );
nor g895 ( new_n1238_, new_n1237_, keyIn_0_243 );
nand g896 ( new_n1239_, new_n1237_, keyIn_0_243 );
not g897 ( new_n1240_, keyIn_0_203 );
nand g898 ( new_n1241_, new_n1226_, N228 );
nand g899 ( new_n1242_, new_n1029_, N237 );
xnor g900 ( new_n1243_, new_n1242_, keyIn_0_182 );
nand g901 ( new_n1244_, new_n1241_, new_n1243_ );
nand g902 ( new_n1245_, new_n1244_, new_n1240_ );
not g903 ( new_n1246_, new_n1245_ );
not g904 ( new_n1247_, new_n1244_ );
nand g905 ( new_n1248_, new_n1247_, keyIn_0_203 );
not g906 ( new_n1249_, keyIn_0_161 );
not g907 ( new_n1250_, new_n991_ );
nand g908 ( new_n1251_, new_n1250_, N246 );
nand g909 ( new_n1252_, new_n700_, N171 );
xnor g910 ( new_n1253_, new_n1252_, keyIn_0_119 );
nand g911 ( new_n1254_, new_n1251_, new_n1253_ );
nor g912 ( new_n1255_, new_n1254_, new_n1249_ );
nand g913 ( new_n1256_, new_n1254_, new_n1249_ );
nand g914 ( new_n1257_, N96, N210 );
xor g915 ( new_n1258_, new_n1257_, keyIn_0_33 );
nand g916 ( new_n1259_, new_n1256_, new_n1258_ );
nor g917 ( new_n1260_, new_n1259_, new_n1255_ );
nand g918 ( new_n1261_, new_n1248_, new_n1260_ );
nor g919 ( new_n1262_, new_n1261_, new_n1246_ );
nand g920 ( new_n1263_, new_n1239_, new_n1262_ );
nor g921 ( new_n1264_, new_n1263_, new_n1238_ );
xor g922 ( N880, new_n1264_, keyIn_0_252 );
endmodule