module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n1009_, new_n479_, new_n955_, new_n608_, new_n888_, new_n847_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n1073_, new_n902_, new_n364_, new_n449_, new_n639_, new_n484_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n845_, new_n768_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n1062_, new_n925_, new_n875_, new_n680_, new_n506_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1026_, new_n267_, new_n473_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n1061_, new_n668_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n313_, new_n382_, new_n583_, new_n239_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n337_, new_n623_, new_n446_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n978_, new_n408_, new_n470_, new_n1072_, new_n769_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n697_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n573_, new_n765_, new_n405_;

nand g000 ( new_n215_, N29, N42, N75 );
not g001 ( N388, new_n215_ );
nand g002 ( new_n217_, N29, N36, N80 );
not g003 ( N389, new_n217_ );
nand g004 ( new_n219_, N29, N36, N42 );
not g005 ( N390, new_n219_ );
nand g006 ( new_n221_, N85, N86 );
not g007 ( N391, new_n221_ );
nand g008 ( new_n223_, N1, N8 );
not g009 ( new_n224_, new_n223_ );
nand g010 ( new_n225_, new_n224_, N13, N17 );
not g011 ( N418, new_n225_ );
not g012 ( new_n227_, N13 );
not g013 ( new_n228_, N17 );
nand g014 ( new_n229_, N1, N26 );
nor g015 ( new_n230_, new_n229_, new_n227_, new_n228_ );
nand g016 ( N419, new_n230_, new_n219_ );
nand g017 ( N420, N59, N75, N80 );
nand g018 ( N421, N36, N59, N80 );
nand g019 ( N422, N36, N42, N59 );
not g020 ( new_n235_, N90 );
nor g021 ( new_n236_, N87, N88 );
nor g022 ( N423, new_n236_, new_n235_ );
nand g023 ( N446, new_n230_, N390 );
nand g024 ( new_n239_, N1, N26, N51 );
nand g025 ( new_n240_, new_n239_, keyIn_0_0 );
not g026 ( new_n241_, keyIn_0_0 );
nand g027 ( new_n242_, new_n241_, N1, N26, N51 );
nand g028 ( N447, new_n240_, new_n242_ );
nand g029 ( new_n244_, new_n224_, N13, N55 );
nand g030 ( new_n245_, N29, N68 );
nor g031 ( N448, new_n244_, new_n245_ );
not g032 ( new_n247_, N74 );
not g033 ( new_n248_, new_n244_ );
nand g034 ( new_n249_, new_n248_, N59, N68 );
nor g035 ( N449, new_n249_, new_n247_ );
not g036 ( new_n251_, N89 );
nor g037 ( N450, new_n236_, new_n251_ );
not g038 ( new_n253_, N126 );
nand g039 ( new_n254_, new_n253_, N121 );
not g040 ( new_n255_, N121 );
nand g041 ( new_n256_, new_n255_, N126 );
nand g042 ( new_n257_, new_n254_, new_n256_ );
nand g043 ( new_n258_, new_n257_, keyIn_0_15 );
not g044 ( new_n259_, keyIn_0_15 );
nand g045 ( new_n260_, new_n254_, new_n256_, new_n259_ );
nand g046 ( new_n261_, new_n258_, new_n260_ );
not g047 ( new_n262_, new_n261_ );
not g048 ( new_n263_, N111 );
not g049 ( new_n264_, N116 );
nand g050 ( new_n265_, new_n263_, new_n264_ );
nand g051 ( new_n266_, N111, N116 );
nand g052 ( new_n267_, new_n265_, new_n266_ );
nand g053 ( new_n268_, new_n267_, keyIn_0_14 );
not g054 ( new_n269_, keyIn_0_14 );
nand g055 ( new_n270_, new_n265_, new_n269_, new_n266_ );
nand g056 ( new_n271_, new_n268_, new_n270_ );
nor g057 ( new_n272_, new_n262_, new_n271_ );
not g058 ( new_n273_, new_n272_ );
nand g059 ( new_n274_, new_n273_, keyIn_0_24 );
not g060 ( new_n275_, keyIn_0_24 );
nand g061 ( new_n276_, new_n272_, new_n275_ );
nand g062 ( new_n277_, new_n274_, new_n276_ );
nand g063 ( new_n278_, new_n262_, new_n271_ );
nand g064 ( new_n279_, new_n278_, keyIn_0_29 );
not g065 ( new_n280_, keyIn_0_29 );
nand g066 ( new_n281_, new_n262_, new_n280_, new_n271_ );
nand g067 ( new_n282_, new_n279_, new_n281_ );
nand g068 ( new_n283_, new_n277_, new_n282_ );
nand g069 ( new_n284_, new_n283_, keyIn_0_38 );
not g070 ( new_n285_, keyIn_0_38 );
nand g071 ( new_n286_, new_n277_, new_n285_, new_n282_ );
nand g072 ( new_n287_, new_n284_, new_n286_ );
nand g073 ( new_n288_, new_n287_, N135 );
not g074 ( new_n289_, N135 );
nand g075 ( new_n290_, new_n284_, new_n289_, new_n286_ );
nand g076 ( new_n291_, new_n288_, new_n290_ );
not g077 ( new_n292_, keyIn_0_23 );
not g078 ( new_n293_, N96 );
nand g079 ( new_n294_, new_n293_, N91 );
not g080 ( new_n295_, N91 );
nand g081 ( new_n296_, new_n295_, N96 );
nand g082 ( new_n297_, new_n294_, new_n296_ );
nand g083 ( new_n298_, new_n297_, keyIn_0_12 );
not g084 ( new_n299_, keyIn_0_12 );
nand g085 ( new_n300_, new_n294_, new_n296_, new_n299_ );
nand g086 ( new_n301_, new_n298_, new_n300_ );
not g087 ( new_n302_, new_n301_ );
not g088 ( new_n303_, N101 );
not g089 ( new_n304_, N106 );
nand g090 ( new_n305_, new_n303_, new_n304_ );
nand g091 ( new_n306_, N101, N106 );
nand g092 ( new_n307_, new_n305_, new_n306_ );
nand g093 ( new_n308_, new_n307_, keyIn_0_13 );
not g094 ( new_n309_, keyIn_0_13 );
nand g095 ( new_n310_, new_n305_, new_n309_, new_n306_ );
nand g096 ( new_n311_, new_n308_, new_n310_ );
nor g097 ( new_n312_, new_n302_, new_n311_ );
not g098 ( new_n313_, new_n312_ );
nand g099 ( new_n314_, new_n313_, new_n292_ );
nand g100 ( new_n315_, new_n312_, keyIn_0_23 );
nand g101 ( new_n316_, new_n314_, new_n315_ );
not g102 ( new_n317_, keyIn_0_28 );
nand g103 ( new_n318_, new_n302_, new_n311_ );
nand g104 ( new_n319_, new_n318_, new_n317_ );
nand g105 ( new_n320_, new_n302_, keyIn_0_28, new_n311_ );
nand g106 ( new_n321_, new_n319_, new_n320_ );
nand g107 ( new_n322_, new_n316_, new_n321_ );
nand g108 ( new_n323_, new_n322_, keyIn_0_37 );
not g109 ( new_n324_, keyIn_0_37 );
nand g110 ( new_n325_, new_n316_, new_n324_, new_n321_ );
nand g111 ( new_n326_, new_n323_, new_n325_ );
nand g112 ( new_n327_, new_n326_, N130 );
not g113 ( new_n328_, N130 );
nand g114 ( new_n329_, new_n323_, new_n328_, new_n325_ );
nand g115 ( new_n330_, new_n327_, new_n329_ );
nand g116 ( new_n331_, new_n291_, new_n330_ );
nand g117 ( new_n332_, new_n288_, new_n327_, new_n290_, new_n329_ );
nand g118 ( N767, new_n331_, new_n332_ );
not g119 ( new_n334_, keyIn_0_26 );
nand g120 ( new_n335_, N159, N165 );
not g121 ( new_n336_, new_n335_ );
nor g122 ( new_n337_, N159, N165 );
nor g123 ( new_n338_, new_n336_, new_n337_ );
not g124 ( new_n339_, new_n338_ );
nor g125 ( new_n340_, new_n339_, keyIn_0_18 );
nand g126 ( new_n341_, new_n339_, keyIn_0_18 );
not g127 ( new_n342_, new_n341_ );
nor g128 ( new_n343_, new_n342_, new_n340_ );
not g129 ( new_n344_, new_n343_ );
not g130 ( new_n345_, N177 );
nand g131 ( new_n346_, new_n345_, N171 );
not g132 ( new_n347_, N171 );
nand g133 ( new_n348_, new_n347_, N177 );
nand g134 ( new_n349_, new_n346_, new_n348_ );
nand g135 ( new_n350_, new_n349_, keyIn_0_19 );
not g136 ( new_n351_, keyIn_0_19 );
nand g137 ( new_n352_, new_n346_, new_n348_, new_n351_ );
nand g138 ( new_n353_, new_n350_, new_n352_ );
nand g139 ( new_n354_, new_n344_, new_n353_ );
nand g140 ( new_n355_, new_n354_, new_n334_ );
nand g141 ( new_n356_, new_n344_, keyIn_0_26, new_n353_ );
nand g142 ( new_n357_, new_n355_, new_n356_ );
not g143 ( new_n358_, keyIn_0_35 );
not g144 ( new_n359_, new_n353_ );
nand g145 ( new_n360_, new_n343_, new_n359_ );
nand g146 ( new_n361_, new_n360_, new_n358_ );
nand g147 ( new_n362_, new_n343_, keyIn_0_35, new_n359_ );
nand g148 ( new_n363_, new_n361_, new_n362_ );
nand g149 ( new_n364_, new_n357_, new_n363_ );
nand g150 ( new_n365_, new_n364_, keyIn_0_49 );
not g151 ( new_n366_, keyIn_0_49 );
nand g152 ( new_n367_, new_n357_, new_n366_, new_n363_ );
nand g153 ( new_n368_, new_n365_, new_n367_ );
nand g154 ( new_n369_, new_n368_, new_n328_ );
nand g155 ( new_n370_, new_n365_, N130, new_n367_ );
nand g156 ( new_n371_, new_n369_, new_n370_ );
not g157 ( new_n372_, keyIn_0_36 );
nand g158 ( new_n373_, N195, N201 );
not g159 ( new_n374_, new_n373_ );
nor g160 ( new_n375_, N195, N201 );
nor g161 ( new_n376_, new_n374_, new_n375_ );
not g162 ( new_n377_, new_n376_ );
nor g163 ( new_n378_, new_n377_, keyIn_0_21 );
nand g164 ( new_n379_, new_n377_, keyIn_0_21 );
not g165 ( new_n380_, new_n379_ );
nor g166 ( new_n381_, new_n380_, new_n378_ );
not g167 ( new_n382_, new_n381_ );
not g168 ( new_n383_, N189 );
nand g169 ( new_n384_, new_n383_, N183 );
not g170 ( new_n385_, N183 );
nand g171 ( new_n386_, new_n385_, N189 );
nand g172 ( new_n387_, new_n384_, new_n386_ );
nand g173 ( new_n388_, new_n387_, keyIn_0_20 );
not g174 ( new_n389_, keyIn_0_20 );
nand g175 ( new_n390_, new_n384_, new_n386_, new_n389_ );
nand g176 ( new_n391_, new_n388_, new_n390_ );
nand g177 ( new_n392_, new_n382_, new_n391_ );
nand g178 ( new_n393_, new_n392_, new_n372_ );
nand g179 ( new_n394_, new_n382_, keyIn_0_36, new_n391_ );
nand g180 ( new_n395_, new_n393_, new_n394_ );
not g181 ( new_n396_, new_n391_ );
nand g182 ( new_n397_, new_n381_, new_n396_ );
nand g183 ( new_n398_, new_n397_, keyIn_0_27 );
not g184 ( new_n399_, keyIn_0_27 );
nand g185 ( new_n400_, new_n381_, new_n399_, new_n396_ );
nand g186 ( new_n401_, new_n398_, new_n400_ );
nand g187 ( new_n402_, new_n395_, new_n401_ );
nand g188 ( new_n403_, new_n402_, keyIn_0_50 );
not g189 ( new_n404_, keyIn_0_50 );
nand g190 ( new_n405_, new_n395_, new_n404_, new_n401_ );
nand g191 ( new_n406_, new_n403_, new_n405_ );
nand g192 ( new_n407_, new_n406_, N207 );
not g193 ( new_n408_, N207 );
nand g194 ( new_n409_, new_n403_, new_n408_, new_n405_ );
nand g195 ( new_n410_, new_n407_, new_n409_ );
nand g196 ( new_n411_, new_n371_, new_n410_ );
nand g197 ( new_n412_, new_n369_, new_n407_, new_n370_, new_n409_ );
nand g198 ( N768, new_n411_, new_n412_ );
not g199 ( new_n414_, keyIn_0_112 );
not g200 ( new_n415_, N261 );
not g201 ( new_n416_, keyIn_0_94 );
not g202 ( new_n417_, keyIn_0_62 );
not g203 ( new_n418_, keyIn_0_22 );
not g204 ( new_n419_, keyIn_0_8 );
nand g205 ( new_n420_, N447, new_n419_ );
nand g206 ( new_n421_, new_n240_, keyIn_0_8, new_n242_ );
nand g207 ( new_n422_, new_n420_, new_n421_ );
nand g208 ( new_n423_, new_n422_, new_n418_ );
nand g209 ( new_n424_, new_n420_, keyIn_0_22, new_n421_ );
nand g210 ( new_n425_, new_n423_, new_n424_ );
nand g211 ( new_n426_, N59, N156 );
not g212 ( new_n427_, new_n426_ );
not g213 ( new_n428_, N42 );
nand g214 ( new_n429_, new_n228_, new_n428_ );
nand g215 ( new_n430_, new_n429_, keyIn_0_6 );
not g216 ( new_n431_, keyIn_0_6 );
nand g217 ( new_n432_, new_n431_, new_n228_, new_n428_ );
nand g218 ( new_n433_, new_n430_, new_n432_ );
not g219 ( new_n434_, keyIn_0_7 );
nand g220 ( new_n435_, N17, N42 );
nand g221 ( new_n436_, new_n435_, new_n434_ );
nand g222 ( new_n437_, keyIn_0_7, N17, N42 );
nand g223 ( new_n438_, new_n436_, new_n437_ );
nand g224 ( new_n439_, new_n433_, new_n438_ );
nand g225 ( new_n440_, new_n439_, keyIn_0_17 );
not g226 ( new_n441_, keyIn_0_17 );
nand g227 ( new_n442_, new_n433_, new_n441_, new_n438_ );
nand g228 ( new_n443_, new_n440_, new_n442_ );
nand g229 ( new_n444_, new_n425_, keyIn_0_33, new_n427_, new_n443_ );
not g230 ( new_n445_, keyIn_0_33 );
nand g231 ( new_n446_, new_n425_, new_n427_, new_n443_ );
nand g232 ( new_n447_, new_n446_, new_n445_ );
nand g233 ( new_n448_, N1, N8, N17, N51 );
nand g234 ( new_n449_, new_n448_, keyIn_0_1 );
not g235 ( new_n450_, keyIn_0_1 );
nand g236 ( new_n451_, new_n224_, new_n450_, N17, N51 );
nand g237 ( new_n452_, new_n451_, new_n449_ );
nand g238 ( new_n453_, new_n452_, keyIn_0_9 );
not g239 ( new_n454_, keyIn_0_9 );
nand g240 ( new_n455_, new_n451_, new_n454_, new_n449_ );
nand g241 ( new_n456_, new_n453_, new_n455_ );
not g242 ( new_n457_, keyIn_0_11 );
not g243 ( new_n458_, keyIn_0_3 );
nand g244 ( new_n459_, N42, N59, N75 );
nand g245 ( new_n460_, new_n459_, new_n458_ );
nand g246 ( new_n461_, keyIn_0_3, N42, N59, N75 );
nand g247 ( new_n462_, new_n460_, new_n461_ );
nand g248 ( new_n463_, new_n462_, new_n457_ );
nand g249 ( new_n464_, new_n460_, keyIn_0_11, new_n461_ );
nand g250 ( new_n465_, new_n463_, new_n464_ );
nand g251 ( new_n466_, new_n456_, new_n465_ );
nand g252 ( new_n467_, new_n466_, keyIn_0_25 );
not g253 ( new_n468_, keyIn_0_25 );
nand g254 ( new_n469_, new_n456_, new_n465_, new_n468_ );
nand g255 ( new_n470_, new_n447_, new_n444_, new_n467_, new_n469_ );
nand g256 ( new_n471_, new_n470_, keyIn_0_39 );
not g257 ( new_n472_, keyIn_0_39 );
nand g258 ( new_n473_, new_n467_, new_n469_ );
not g259 ( new_n474_, new_n473_ );
nand g260 ( new_n475_, new_n474_, new_n472_, new_n444_, new_n447_ );
nand g261 ( new_n476_, new_n471_, new_n475_ );
nand g262 ( new_n477_, new_n476_, N126 );
nand g263 ( new_n478_, new_n477_, new_n417_ );
nand g264 ( new_n479_, new_n476_, keyIn_0_62, N126 );
nand g265 ( new_n480_, new_n478_, new_n479_ );
nand g266 ( new_n481_, new_n427_, keyIn_0_5 );
not g267 ( new_n482_, keyIn_0_5 );
nand g268 ( new_n483_, new_n426_, new_n482_ );
nand g269 ( new_n484_, new_n481_, new_n483_ );
not g270 ( new_n485_, new_n484_ );
nand g271 ( new_n486_, new_n425_, N17, new_n485_ );
nand g272 ( new_n487_, new_n486_, keyIn_0_34 );
not g273 ( new_n488_, keyIn_0_34 );
nand g274 ( new_n489_, new_n425_, new_n488_, N17, new_n485_ );
nand g275 ( new_n490_, new_n487_, new_n489_ );
nand g276 ( new_n491_, new_n490_, N1 );
nand g277 ( new_n492_, new_n491_, keyIn_0_44 );
not g278 ( new_n493_, keyIn_0_44 );
nand g279 ( new_n494_, new_n490_, new_n493_, N1 );
nand g280 ( new_n495_, new_n492_, N153, new_n494_ );
nand g281 ( new_n496_, new_n495_, keyIn_0_61 );
not g282 ( new_n497_, keyIn_0_61 );
nand g283 ( new_n498_, new_n492_, new_n494_ );
not g284 ( new_n499_, new_n498_ );
nand g285 ( new_n500_, new_n499_, new_n497_, N153 );
nand g286 ( new_n501_, new_n480_, new_n496_, new_n500_ );
nand g287 ( new_n502_, new_n501_, keyIn_0_70 );
not g288 ( new_n503_, keyIn_0_70 );
nand g289 ( new_n504_, new_n480_, new_n503_, new_n496_, new_n500_ );
nand g290 ( new_n505_, new_n502_, new_n504_ );
not g291 ( new_n506_, keyIn_0_48 );
nand g292 ( new_n507_, N29, N75, N80 );
nand g293 ( new_n508_, new_n507_, keyIn_0_2 );
not g294 ( new_n509_, keyIn_0_2 );
nand g295 ( new_n510_, new_n509_, N29, N75, N80 );
nand g296 ( new_n511_, new_n425_, new_n508_, new_n510_ );
not g297 ( new_n512_, new_n511_ );
nand g298 ( new_n513_, new_n512_, N55 );
nand g299 ( new_n514_, new_n513_, keyIn_0_32 );
not g300 ( new_n515_, keyIn_0_32 );
nand g301 ( new_n516_, new_n512_, new_n515_, N55 );
nand g302 ( new_n517_, new_n514_, new_n516_ );
nand g303 ( new_n518_, keyIn_0_4, N268 );
not g304 ( new_n519_, new_n518_ );
nor g305 ( new_n520_, keyIn_0_4, N268 );
nor g306 ( new_n521_, new_n519_, new_n520_ );
not g307 ( new_n522_, new_n521_ );
nor g308 ( new_n523_, new_n522_, keyIn_0_16 );
nand g309 ( new_n524_, new_n522_, keyIn_0_16 );
not g310 ( new_n525_, new_n524_ );
nor g311 ( new_n526_, new_n525_, new_n523_ );
nand g312 ( new_n527_, new_n517_, new_n526_ );
not g313 ( new_n528_, new_n527_ );
nand g314 ( new_n529_, new_n528_, new_n506_ );
nand g315 ( new_n530_, new_n527_, keyIn_0_48 );
nand g316 ( new_n531_, new_n529_, new_n530_ );
nand g317 ( new_n532_, new_n505_, new_n531_ );
nand g318 ( new_n533_, new_n532_, keyIn_0_78 );
not g319 ( new_n534_, keyIn_0_78 );
nand g320 ( new_n535_, new_n505_, new_n534_, new_n531_ );
nand g321 ( new_n536_, new_n533_, new_n535_ );
nand g322 ( new_n537_, new_n536_, N201 );
nand g323 ( new_n538_, new_n537_, keyIn_0_83 );
not g324 ( new_n539_, keyIn_0_83 );
nand g325 ( new_n540_, new_n536_, new_n539_, N201 );
nand g326 ( new_n541_, new_n538_, new_n540_ );
not g327 ( new_n542_, keyIn_0_84 );
not g328 ( new_n543_, N201 );
nand g329 ( new_n544_, new_n533_, new_n543_, new_n535_ );
nand g330 ( new_n545_, new_n544_, new_n542_ );
nand g331 ( new_n546_, new_n533_, keyIn_0_84, new_n543_, new_n535_ );
nand g332 ( new_n547_, new_n545_, new_n546_ );
not g333 ( new_n548_, new_n547_ );
nand g334 ( new_n549_, new_n548_, new_n541_ );
nand g335 ( new_n550_, new_n549_, new_n416_ );
nand g336 ( new_n551_, new_n548_, new_n541_, keyIn_0_94 );
nand g337 ( new_n552_, new_n550_, new_n415_, new_n551_ );
nand g338 ( new_n553_, new_n550_, new_n551_ );
nand g339 ( new_n554_, new_n553_, N261 );
nand g340 ( new_n555_, new_n554_, N219, new_n552_ );
nand g341 ( new_n556_, new_n553_, N228 );
not g342 ( new_n557_, keyIn_0_93 );
nand g343 ( new_n558_, new_n541_, new_n557_ );
nand g344 ( new_n559_, new_n538_, keyIn_0_93, new_n540_ );
nand g345 ( new_n560_, new_n558_, new_n559_ );
nand g346 ( new_n561_, new_n560_, N237 );
nand g347 ( new_n562_, new_n536_, N246 );
not g348 ( new_n563_, keyIn_0_10 );
not g349 ( new_n564_, N72 );
nor g350 ( new_n565_, new_n249_, new_n428_, new_n564_ );
nor g351 ( new_n566_, new_n565_, new_n563_ );
nand g352 ( new_n567_, new_n565_, new_n563_ );
nand g353 ( new_n568_, new_n567_, N73 );
nor g354 ( new_n569_, new_n568_, new_n566_ );
nand g355 ( new_n570_, new_n569_, N201 );
nand g356 ( new_n571_, N255, N267 );
nand g357 ( new_n572_, N121, N210 );
nand g358 ( new_n573_, new_n570_, new_n571_, new_n572_ );
not g359 ( new_n574_, new_n573_ );
nand g360 ( new_n575_, new_n561_, new_n562_, new_n574_ );
not g361 ( new_n576_, new_n575_ );
nand g362 ( new_n577_, new_n555_, new_n556_, new_n576_ );
nand g363 ( new_n578_, new_n577_, new_n414_ );
nand g364 ( new_n579_, new_n555_, keyIn_0_112, new_n556_, new_n576_ );
nand g365 ( N850, new_n578_, new_n579_ );
not g366 ( new_n581_, keyIn_0_121 );
not g367 ( new_n582_, keyIn_0_89 );
not g368 ( new_n583_, keyIn_0_75 );
not g369 ( new_n584_, keyIn_0_67 );
nand g370 ( new_n585_, new_n499_, N143 );
nand g371 ( new_n586_, new_n585_, keyIn_0_55 );
not g372 ( new_n587_, keyIn_0_56 );
nand g373 ( new_n588_, new_n476_, N111 );
nand g374 ( new_n589_, new_n588_, new_n587_ );
nand g375 ( new_n590_, new_n476_, keyIn_0_56, N111 );
not g376 ( new_n591_, keyIn_0_55 );
nand g377 ( new_n592_, new_n499_, new_n591_, N143 );
nand g378 ( new_n593_, new_n586_, new_n589_, new_n590_, new_n592_ );
nand g379 ( new_n594_, new_n593_, new_n584_ );
not g380 ( new_n595_, keyIn_0_45 );
nand g381 ( new_n596_, new_n528_, new_n595_ );
nand g382 ( new_n597_, new_n527_, keyIn_0_45 );
nand g383 ( new_n598_, new_n596_, new_n597_ );
not g384 ( new_n599_, new_n593_ );
nand g385 ( new_n600_, new_n599_, keyIn_0_67 );
nand g386 ( new_n601_, new_n600_, new_n594_, new_n598_ );
nand g387 ( new_n602_, new_n601_, new_n583_ );
nand g388 ( new_n603_, new_n600_, keyIn_0_75, new_n594_, new_n598_ );
nand g389 ( new_n604_, new_n602_, new_n603_ );
nand g390 ( new_n605_, new_n604_, N183 );
nand g391 ( new_n606_, new_n602_, new_n385_, new_n603_ );
nand g392 ( new_n607_, new_n605_, new_n606_ );
nand g393 ( new_n608_, new_n607_, new_n582_ );
nand g394 ( new_n609_, new_n605_, keyIn_0_89, new_n606_ );
nand g395 ( new_n610_, new_n608_, new_n609_ );
not g396 ( new_n611_, keyIn_0_103 );
not g397 ( new_n612_, keyIn_0_99 );
not g398 ( new_n613_, keyIn_0_76 );
nand g399 ( new_n614_, new_n476_, N116 );
nand g400 ( new_n615_, new_n614_, keyIn_0_58 );
not g401 ( new_n616_, keyIn_0_58 );
nand g402 ( new_n617_, new_n476_, new_n616_, N116 );
nand g403 ( new_n618_, new_n615_, new_n617_ );
nand g404 ( new_n619_, new_n492_, N146, new_n494_ );
nand g405 ( new_n620_, new_n619_, keyIn_0_57 );
not g406 ( new_n621_, keyIn_0_57 );
nand g407 ( new_n622_, new_n499_, new_n621_, N146 );
nand g408 ( new_n623_, new_n618_, keyIn_0_68, new_n620_, new_n622_ );
not g409 ( new_n624_, keyIn_0_68 );
nand g410 ( new_n625_, new_n618_, new_n620_, new_n622_ );
nand g411 ( new_n626_, new_n625_, new_n624_ );
not g412 ( new_n627_, keyIn_0_46 );
nand g413 ( new_n628_, new_n528_, new_n627_ );
nand g414 ( new_n629_, new_n527_, keyIn_0_46 );
nand g415 ( new_n630_, new_n628_, new_n629_ );
not g416 ( new_n631_, new_n630_ );
nand g417 ( new_n632_, new_n626_, new_n623_, new_n631_ );
nand g418 ( new_n633_, new_n632_, new_n613_ );
nand g419 ( new_n634_, new_n626_, keyIn_0_76, new_n623_, new_n631_ );
nand g420 ( new_n635_, new_n633_, new_n634_ );
nand g421 ( new_n636_, new_n635_, new_n383_ );
nand g422 ( new_n637_, new_n636_, keyIn_0_80 );
not g423 ( new_n638_, keyIn_0_80 );
nand g424 ( new_n639_, new_n635_, new_n638_, new_n383_ );
nand g425 ( new_n640_, new_n637_, new_n639_ );
not g426 ( new_n641_, new_n640_ );
not g427 ( new_n642_, N195 );
not g428 ( new_n643_, keyIn_0_77 );
not g429 ( new_n644_, keyIn_0_69 );
nand g430 ( new_n645_, new_n476_, N121 );
nand g431 ( new_n646_, new_n645_, keyIn_0_60 );
not g432 ( new_n647_, keyIn_0_60 );
nand g433 ( new_n648_, new_n476_, new_n647_, N121 );
nand g434 ( new_n649_, new_n646_, new_n648_ );
nand g435 ( new_n650_, new_n492_, N149, new_n494_ );
nand g436 ( new_n651_, new_n650_, keyIn_0_59 );
not g437 ( new_n652_, keyIn_0_59 );
nand g438 ( new_n653_, new_n492_, new_n652_, N149, new_n494_ );
nand g439 ( new_n654_, new_n651_, new_n653_ );
nand g440 ( new_n655_, new_n649_, new_n644_, new_n654_ );
nand g441 ( new_n656_, new_n649_, new_n654_ );
nand g442 ( new_n657_, new_n656_, keyIn_0_69 );
not g443 ( new_n658_, keyIn_0_47 );
nand g444 ( new_n659_, new_n528_, new_n658_ );
nand g445 ( new_n660_, new_n527_, keyIn_0_47 );
nand g446 ( new_n661_, new_n659_, new_n660_ );
not g447 ( new_n662_, new_n661_ );
nand g448 ( new_n663_, new_n657_, new_n655_, new_n662_ );
nand g449 ( new_n664_, new_n663_, new_n643_ );
nand g450 ( new_n665_, new_n657_, keyIn_0_77, new_n655_, new_n662_ );
nand g451 ( new_n666_, new_n664_, new_n665_ );
nand g452 ( new_n667_, new_n666_, new_n642_ );
nand g453 ( new_n668_, new_n667_, keyIn_0_82 );
not g454 ( new_n669_, keyIn_0_82 );
nand g455 ( new_n670_, new_n666_, new_n669_, new_n642_ );
nand g456 ( new_n671_, new_n668_, new_n670_ );
nand g457 ( new_n672_, new_n560_, new_n641_, new_n671_ );
nand g458 ( new_n673_, new_n672_, new_n612_ );
nand g459 ( new_n674_, new_n560_, keyIn_0_99, new_n641_, new_n671_ );
nand g460 ( new_n675_, new_n673_, new_n674_ );
not g461 ( new_n676_, keyIn_0_96 );
not g462 ( new_n677_, new_n671_ );
nand g463 ( new_n678_, new_n545_, N261, new_n546_ );
nor g464 ( new_n679_, new_n677_, new_n678_, new_n640_ );
nor g465 ( new_n680_, new_n679_, new_n676_ );
nand g466 ( new_n681_, new_n671_, N261, new_n545_, new_n546_ );
nor g467 ( new_n682_, new_n681_, keyIn_0_96, new_n640_ );
nor g468 ( new_n683_, new_n680_, new_n682_ );
not g469 ( new_n684_, keyIn_0_91 );
nand g470 ( new_n685_, new_n664_, N195, new_n665_ );
nand g471 ( new_n686_, new_n685_, keyIn_0_81 );
not g472 ( new_n687_, keyIn_0_81 );
nand g473 ( new_n688_, new_n664_, new_n687_, N195, new_n665_ );
nand g474 ( new_n689_, new_n686_, new_n688_ );
nand g475 ( new_n690_, new_n689_, new_n684_ );
nand g476 ( new_n691_, new_n686_, keyIn_0_91, new_n688_ );
nand g477 ( new_n692_, new_n690_, new_n691_ );
nand g478 ( new_n693_, new_n692_, new_n641_ );
nand g479 ( new_n694_, new_n693_, keyIn_0_98 );
not g480 ( new_n695_, keyIn_0_98 );
nand g481 ( new_n696_, new_n692_, new_n695_, new_n641_ );
nand g482 ( new_n697_, new_n694_, new_n696_ );
not g483 ( new_n698_, new_n635_ );
nand g484 ( new_n699_, new_n698_, N189 );
nand g485 ( new_n700_, new_n699_, keyIn_0_79 );
not g486 ( new_n701_, keyIn_0_79 );
nand g487 ( new_n702_, new_n698_, new_n701_, N189 );
nand g488 ( new_n703_, new_n700_, new_n702_ );
not g489 ( new_n704_, new_n703_ );
nand g490 ( new_n705_, new_n697_, new_n704_ );
nor g491 ( new_n706_, new_n705_, new_n683_ );
nand g492 ( new_n707_, new_n706_, new_n675_ );
nand g493 ( new_n708_, new_n707_, new_n611_ );
nand g494 ( new_n709_, new_n706_, keyIn_0_103, new_n675_ );
nand g495 ( new_n710_, new_n708_, new_n709_ );
not g496 ( new_n711_, new_n710_ );
nand g497 ( new_n712_, new_n711_, keyIn_0_106, new_n610_ );
not g498 ( new_n713_, keyIn_0_106 );
nand g499 ( new_n714_, new_n711_, new_n610_ );
nand g500 ( new_n715_, new_n714_, new_n713_ );
nand g501 ( new_n716_, new_n710_, new_n608_, new_n609_ );
nand g502 ( new_n717_, new_n715_, N219, new_n712_, new_n716_ );
nand g503 ( new_n718_, new_n610_, N228 );
nand g504 ( new_n719_, new_n604_, N183, N237 );
nand g505 ( new_n720_, new_n604_, N246 );
nand g506 ( new_n721_, N106, N210 );
nand g507 ( new_n722_, new_n569_, N183 );
nand g508 ( new_n723_, new_n720_, new_n721_, new_n722_ );
not g509 ( new_n724_, new_n723_ );
nand g510 ( new_n725_, new_n718_, new_n719_, new_n724_ );
not g511 ( new_n726_, new_n725_ );
nand g512 ( new_n727_, new_n717_, new_n726_ );
nand g513 ( new_n728_, new_n727_, new_n581_ );
nand g514 ( new_n729_, new_n717_, keyIn_0_121, new_n726_ );
nand g515 ( N863, new_n728_, new_n729_ );
not g516 ( new_n731_, keyIn_0_107 );
nand g517 ( new_n732_, new_n560_, new_n671_ );
nand g518 ( new_n733_, new_n732_, keyIn_0_97 );
not g519 ( new_n734_, keyIn_0_97 );
nand g520 ( new_n735_, new_n560_, new_n734_, new_n671_ );
nand g521 ( new_n736_, new_n733_, new_n735_ );
not g522 ( new_n737_, keyIn_0_95 );
nand g523 ( new_n738_, new_n548_, new_n737_, N261, new_n671_ );
nand g524 ( new_n739_, new_n681_, keyIn_0_95 );
nand g525 ( new_n740_, new_n738_, new_n739_, new_n690_, new_n691_ );
not g526 ( new_n741_, new_n740_ );
nand g527 ( new_n742_, new_n736_, new_n741_ );
nand g528 ( new_n743_, new_n742_, keyIn_0_104 );
not g529 ( new_n744_, keyIn_0_104 );
nand g530 ( new_n745_, new_n736_, new_n744_, new_n741_ );
nand g531 ( new_n746_, new_n743_, new_n745_ );
not g532 ( new_n747_, keyIn_0_90 );
nor g533 ( new_n748_, new_n703_, new_n640_ );
not g534 ( new_n749_, new_n748_ );
nand g535 ( new_n750_, new_n749_, new_n747_ );
nand g536 ( new_n751_, new_n748_, keyIn_0_90 );
nand g537 ( new_n752_, new_n750_, new_n751_ );
not g538 ( new_n753_, new_n752_ );
nand g539 ( new_n754_, new_n746_, new_n731_, new_n753_ );
nand g540 ( new_n755_, new_n746_, new_n753_ );
nand g541 ( new_n756_, new_n755_, keyIn_0_107 );
nand g542 ( new_n757_, new_n743_, new_n745_, new_n752_ );
nand g543 ( new_n758_, new_n756_, N219, new_n754_, new_n757_ );
nand g544 ( new_n759_, new_n753_, N228 );
nand g545 ( new_n760_, new_n703_, N237 );
nand g546 ( new_n761_, new_n698_, N246 );
nand g547 ( new_n762_, new_n569_, N189 );
nand g548 ( new_n763_, N255, N259 );
nand g549 ( new_n764_, N111, N210 );
nand g550 ( new_n765_, new_n761_, new_n762_, new_n763_, new_n764_ );
not g551 ( new_n766_, new_n765_ );
nand g552 ( new_n767_, new_n759_, new_n760_, new_n766_ );
not g553 ( new_n768_, new_n767_ );
nand g554 ( new_n769_, new_n758_, new_n768_ );
nand g555 ( new_n770_, new_n769_, keyIn_0_122 );
not g556 ( new_n771_, keyIn_0_122 );
nand g557 ( new_n772_, new_n758_, new_n771_, new_n768_ );
nand g558 ( N864, new_n770_, new_n772_ );
not g559 ( new_n774_, new_n560_ );
nand g560 ( new_n775_, new_n774_, new_n678_ );
nand g561 ( new_n776_, new_n775_, keyIn_0_105 );
not g562 ( new_n777_, keyIn_0_105 );
nand g563 ( new_n778_, new_n774_, new_n777_, new_n678_ );
nand g564 ( new_n779_, new_n776_, new_n778_ );
not g565 ( new_n780_, new_n779_ );
nand g566 ( new_n781_, new_n671_, new_n689_ );
nand g567 ( new_n782_, new_n781_, keyIn_0_92 );
not g568 ( new_n783_, keyIn_0_92 );
nand g569 ( new_n784_, new_n671_, new_n783_, new_n689_ );
nand g570 ( new_n785_, new_n782_, new_n784_ );
not g571 ( new_n786_, new_n785_ );
nand g572 ( new_n787_, new_n780_, keyIn_0_108, new_n786_ );
not g573 ( new_n788_, keyIn_0_108 );
nand g574 ( new_n789_, new_n780_, new_n786_ );
nand g575 ( new_n790_, new_n789_, new_n788_ );
nand g576 ( new_n791_, new_n779_, new_n785_ );
nand g577 ( new_n792_, new_n790_, N219, new_n787_, new_n791_ );
nand g578 ( new_n793_, new_n786_, N228 );
not g579 ( new_n794_, new_n793_ );
nand g580 ( new_n795_, new_n692_, N237 );
not g581 ( new_n796_, new_n795_ );
nand g582 ( new_n797_, new_n664_, N246, new_n665_ );
nand g583 ( new_n798_, new_n569_, N195 );
nand g584 ( new_n799_, N255, N260 );
nand g585 ( new_n800_, N116, N210 );
nand g586 ( new_n801_, new_n797_, new_n798_, new_n799_, new_n800_ );
nor g587 ( new_n802_, new_n794_, new_n796_, new_n801_ );
nand g588 ( new_n803_, new_n792_, new_n802_ );
nand g589 ( new_n804_, new_n803_, keyIn_0_123 );
not g590 ( new_n805_, keyIn_0_123 );
nand g591 ( new_n806_, new_n792_, new_n805_, new_n802_ );
nand g592 ( N865, new_n804_, new_n806_ );
not g593 ( new_n808_, keyIn_0_116 );
not g594 ( new_n809_, N165 );
not g595 ( new_n810_, keyIn_0_72 );
not g596 ( new_n811_, keyIn_0_31 );
nand g597 ( new_n812_, new_n512_, N17 );
nand g598 ( new_n813_, new_n812_, new_n811_ );
nand g599 ( new_n814_, new_n512_, keyIn_0_31, N17 );
nand g600 ( new_n815_, new_n813_, new_n814_ );
nand g601 ( new_n816_, new_n815_, new_n521_ );
not g602 ( new_n817_, new_n816_ );
nand g603 ( new_n818_, new_n817_, keyIn_0_41 );
not g604 ( new_n819_, keyIn_0_41 );
nand g605 ( new_n820_, new_n816_, new_n819_ );
nand g606 ( new_n821_, new_n818_, new_n820_ );
not g607 ( new_n822_, keyIn_0_30 );
nand g608 ( new_n823_, new_n425_, N55, new_n485_ );
nand g609 ( new_n824_, new_n823_, new_n822_ );
nand g610 ( new_n825_, new_n425_, keyIn_0_30, N55, new_n485_ );
nand g611 ( new_n826_, new_n824_, new_n825_ );
nand g612 ( new_n827_, new_n826_, N146 );
nand g613 ( new_n828_, new_n821_, new_n827_ );
nand g614 ( new_n829_, new_n828_, keyIn_0_52 );
not g615 ( new_n830_, keyIn_0_52 );
nand g616 ( new_n831_, new_n821_, new_n830_, new_n827_ );
nand g617 ( new_n832_, new_n829_, new_n831_ );
not g618 ( new_n833_, keyIn_0_64 );
nand g619 ( new_n834_, new_n476_, N96 );
nand g620 ( new_n835_, N51, N138 );
nand g621 ( new_n836_, new_n834_, new_n835_ );
nand g622 ( new_n837_, new_n836_, new_n833_ );
nand g623 ( new_n838_, new_n834_, keyIn_0_64, new_n835_ );
nand g624 ( new_n839_, new_n837_, new_n838_ );
nand g625 ( new_n840_, new_n832_, new_n839_ );
nand g626 ( new_n841_, new_n840_, new_n810_ );
nand g627 ( new_n842_, new_n832_, keyIn_0_72, new_n839_ );
nand g628 ( new_n843_, new_n841_, new_n809_, new_n842_ );
not g629 ( new_n844_, keyIn_0_53 );
not g630 ( new_n845_, keyIn_0_42 );
nand g631 ( new_n846_, new_n817_, new_n845_ );
nand g632 ( new_n847_, new_n816_, keyIn_0_42 );
nand g633 ( new_n848_, new_n846_, new_n847_ );
nand g634 ( new_n849_, new_n826_, N149 );
nand g635 ( new_n850_, new_n848_, new_n849_ );
nand g636 ( new_n851_, new_n850_, new_n844_ );
nand g637 ( new_n852_, new_n848_, keyIn_0_53, new_n849_ );
nand g638 ( new_n853_, new_n851_, new_n852_ );
nand g639 ( new_n854_, new_n476_, N101 );
nand g640 ( new_n855_, N17, N138 );
nand g641 ( new_n856_, new_n854_, new_n855_ );
nand g642 ( new_n857_, new_n856_, keyIn_0_65 );
not g643 ( new_n858_, keyIn_0_65 );
nand g644 ( new_n859_, new_n854_, new_n858_, new_n855_ );
nand g645 ( new_n860_, new_n857_, new_n859_ );
nand g646 ( new_n861_, new_n853_, new_n860_ );
nand g647 ( new_n862_, new_n861_, keyIn_0_73 );
not g648 ( new_n863_, keyIn_0_73 );
nand g649 ( new_n864_, new_n853_, new_n863_, new_n860_ );
nand g650 ( new_n865_, new_n862_, new_n864_ );
nand g651 ( new_n866_, new_n865_, new_n347_ );
not g652 ( new_n867_, keyIn_0_109 );
nand g653 ( new_n868_, new_n708_, new_n606_, new_n709_ );
nand g654 ( new_n869_, new_n868_, new_n867_ );
nand g655 ( new_n870_, new_n708_, keyIn_0_109, new_n606_, new_n709_ );
nand g656 ( new_n871_, new_n869_, new_n870_ );
nand g657 ( new_n872_, new_n871_, new_n605_ );
nand g658 ( new_n873_, new_n872_, keyIn_0_110 );
not g659 ( new_n874_, keyIn_0_110 );
nand g660 ( new_n875_, new_n871_, new_n874_, new_n605_ );
nand g661 ( new_n876_, new_n873_, new_n875_ );
not g662 ( new_n877_, keyIn_0_74 );
not g663 ( new_n878_, keyIn_0_54 );
not g664 ( new_n879_, keyIn_0_43 );
nand g665 ( new_n880_, new_n817_, new_n879_ );
nand g666 ( new_n881_, new_n816_, keyIn_0_43 );
nand g667 ( new_n882_, new_n880_, new_n881_ );
nand g668 ( new_n883_, new_n826_, N153 );
nand g669 ( new_n884_, new_n882_, new_n883_ );
nand g670 ( new_n885_, new_n884_, new_n878_ );
nand g671 ( new_n886_, new_n882_, keyIn_0_54, new_n883_ );
nand g672 ( new_n887_, new_n885_, new_n886_ );
nand g673 ( new_n888_, new_n476_, N106 );
nand g674 ( new_n889_, N138, N152 );
nand g675 ( new_n890_, new_n888_, new_n889_ );
nand g676 ( new_n891_, new_n890_, keyIn_0_66 );
not g677 ( new_n892_, keyIn_0_66 );
nand g678 ( new_n893_, new_n888_, new_n892_, new_n889_ );
nand g679 ( new_n894_, new_n891_, new_n893_ );
nand g680 ( new_n895_, new_n887_, new_n894_ );
nand g681 ( new_n896_, new_n895_, new_n877_ );
nand g682 ( new_n897_, new_n887_, keyIn_0_74, new_n894_ );
nand g683 ( new_n898_, new_n896_, new_n345_, new_n897_ );
nand g684 ( new_n899_, new_n876_, new_n843_, new_n866_, new_n898_ );
not g685 ( new_n900_, new_n899_ );
nand g686 ( new_n901_, new_n900_, keyIn_0_115 );
not g687 ( new_n902_, keyIn_0_115 );
nand g688 ( new_n903_, new_n899_, new_n902_ );
nand g689 ( new_n904_, new_n901_, new_n903_ );
not g690 ( new_n905_, new_n865_ );
nand g691 ( new_n906_, new_n905_, N171 );
not g692 ( new_n907_, new_n906_ );
nand g693 ( new_n908_, new_n907_, new_n843_ );
nand g694 ( new_n909_, new_n908_, keyIn_0_101 );
nor g695 ( new_n910_, new_n908_, keyIn_0_101 );
nand g696 ( new_n911_, new_n841_, new_n842_ );
nand g697 ( new_n912_, new_n911_, N165 );
not g698 ( new_n913_, new_n912_ );
nor g699 ( new_n914_, new_n910_, new_n913_ );
nand g700 ( new_n915_, new_n914_, new_n909_ );
not g701 ( new_n916_, keyIn_0_102 );
nand g702 ( new_n917_, new_n896_, new_n897_ );
nand g703 ( new_n918_, new_n917_, N177 );
not g704 ( new_n919_, new_n918_ );
nand g705 ( new_n920_, new_n919_, new_n866_ );
not g706 ( new_n921_, new_n920_ );
nand g707 ( new_n922_, new_n921_, new_n843_ );
nand g708 ( new_n923_, new_n922_, new_n916_ );
not g709 ( new_n924_, new_n923_ );
nor g710 ( new_n925_, new_n922_, new_n916_ );
nor g711 ( new_n926_, new_n915_, new_n924_, new_n925_ );
nand g712 ( new_n927_, new_n904_, new_n926_ );
nand g713 ( new_n928_, new_n927_, new_n808_ );
nand g714 ( new_n929_, new_n904_, keyIn_0_116, new_n926_ );
nand g715 ( new_n930_, new_n928_, new_n929_ );
not g716 ( new_n931_, N159 );
nand g717 ( new_n932_, new_n817_, keyIn_0_40 );
not g718 ( new_n933_, keyIn_0_40 );
nand g719 ( new_n934_, new_n816_, new_n933_ );
nand g720 ( new_n935_, new_n932_, new_n934_ );
nand g721 ( new_n936_, new_n826_, N143 );
nand g722 ( new_n937_, new_n935_, new_n936_ );
nand g723 ( new_n938_, new_n937_, keyIn_0_51 );
not g724 ( new_n939_, keyIn_0_51 );
nand g725 ( new_n940_, new_n935_, new_n939_, new_n936_ );
nand g726 ( new_n941_, new_n938_, new_n940_ );
not g727 ( new_n942_, keyIn_0_63 );
nand g728 ( new_n943_, new_n476_, N91 );
nand g729 ( new_n944_, N8, N138 );
nand g730 ( new_n945_, new_n943_, new_n944_ );
nand g731 ( new_n946_, new_n945_, new_n942_ );
nand g732 ( new_n947_, new_n943_, keyIn_0_63, new_n944_ );
nand g733 ( new_n948_, new_n946_, new_n947_ );
nand g734 ( new_n949_, new_n941_, new_n948_ );
nand g735 ( new_n950_, new_n949_, keyIn_0_71 );
not g736 ( new_n951_, keyIn_0_71 );
nand g737 ( new_n952_, new_n941_, new_n951_, new_n948_ );
nand g738 ( new_n953_, new_n950_, new_n931_, new_n952_ );
nand g739 ( new_n954_, new_n930_, new_n953_ );
nand g740 ( new_n955_, new_n950_, new_n952_ );
nand g741 ( new_n956_, new_n955_, N159 );
nand g742 ( N866, new_n954_, new_n956_ );
not g743 ( new_n958_, keyIn_0_124 );
not g744 ( new_n959_, keyIn_0_111 );
not g745 ( new_n960_, keyIn_0_88 );
nand g746 ( new_n961_, new_n918_, new_n898_ );
nand g747 ( new_n962_, new_n961_, new_n960_ );
nand g748 ( new_n963_, new_n918_, keyIn_0_88, new_n898_ );
nand g749 ( new_n964_, new_n962_, new_n963_ );
not g750 ( new_n965_, new_n964_ );
nand g751 ( new_n966_, new_n876_, new_n965_ );
nand g752 ( new_n967_, new_n966_, new_n959_ );
nand g753 ( new_n968_, new_n876_, keyIn_0_111, new_n965_ );
nand g754 ( new_n969_, new_n967_, new_n968_ );
nand g755 ( new_n970_, new_n873_, new_n875_, new_n964_ );
nand g756 ( new_n971_, new_n969_, N219, new_n970_ );
nand g757 ( new_n972_, new_n965_, N228 );
nand g758 ( new_n973_, new_n919_, N237 );
nand g759 ( new_n974_, new_n917_, N246 );
nand g760 ( new_n975_, N101, N210 );
nand g761 ( new_n976_, new_n569_, N177 );
nand g762 ( new_n977_, new_n974_, new_n975_, new_n976_ );
not g763 ( new_n978_, new_n977_ );
nand g764 ( new_n979_, new_n972_, new_n973_, new_n978_ );
not g765 ( new_n980_, new_n979_ );
nand g766 ( new_n981_, new_n971_, new_n980_ );
nand g767 ( new_n982_, new_n981_, new_n958_ );
nand g768 ( new_n983_, new_n971_, keyIn_0_124, new_n980_ );
nand g769 ( N874, new_n982_, new_n983_ );
nand g770 ( new_n985_, new_n956_, new_n953_ );
nand g771 ( new_n986_, new_n985_, keyIn_0_85 );
not g772 ( new_n987_, keyIn_0_85 );
nand g773 ( new_n988_, new_n956_, new_n987_, new_n953_ );
nand g774 ( new_n989_, new_n986_, new_n988_ );
not g775 ( new_n990_, new_n989_ );
nand g776 ( new_n991_, new_n930_, new_n990_ );
nand g777 ( new_n992_, new_n928_, new_n929_, new_n989_ );
nand g778 ( new_n993_, new_n991_, N219, new_n992_ );
nand g779 ( new_n994_, new_n990_, N228 );
nand g780 ( new_n995_, new_n955_, N159, N237 );
nand g781 ( new_n996_, new_n955_, N246 );
not g782 ( new_n997_, new_n526_ );
nand g783 ( new_n998_, new_n997_, N210 );
nand g784 ( new_n999_, new_n569_, N159 );
nand g785 ( new_n1000_, new_n996_, new_n998_, new_n999_ );
not g786 ( new_n1001_, new_n1000_ );
nand g787 ( new_n1002_, new_n994_, new_n995_, new_n1001_ );
not g788 ( new_n1003_, new_n1002_ );
nand g789 ( new_n1004_, new_n993_, new_n1003_ );
nand g790 ( new_n1005_, new_n1004_, keyIn_0_125 );
not g791 ( new_n1006_, keyIn_0_125 );
nand g792 ( new_n1007_, new_n993_, new_n1006_, new_n1003_ );
nand g793 ( N878, new_n1005_, new_n1007_ );
not g794 ( new_n1009_, keyIn_0_126 );
nand g795 ( new_n1010_, new_n912_, new_n843_ );
nand g796 ( new_n1011_, new_n1010_, keyIn_0_86 );
not g797 ( new_n1012_, keyIn_0_86 );
nand g798 ( new_n1013_, new_n912_, new_n1012_, new_n843_ );
nand g799 ( new_n1014_, new_n1011_, new_n1013_ );
not g800 ( new_n1015_, new_n1014_ );
not g801 ( new_n1016_, keyIn_0_117 );
nand g802 ( new_n1017_, new_n876_, new_n898_ );
not g803 ( new_n1018_, new_n1017_ );
nand g804 ( new_n1019_, new_n1018_, keyIn_0_114, new_n866_ );
not g805 ( new_n1020_, keyIn_0_114 );
nand g806 ( new_n1021_, new_n876_, new_n866_, new_n898_ );
nand g807 ( new_n1022_, new_n1021_, new_n1020_ );
not g808 ( new_n1023_, keyIn_0_100 );
nand g809 ( new_n1024_, new_n921_, new_n1023_ );
nand g810 ( new_n1025_, new_n920_, keyIn_0_100 );
nand g811 ( new_n1026_, new_n1024_, new_n906_, new_n1025_ );
not g812 ( new_n1027_, new_n1026_ );
nand g813 ( new_n1028_, new_n1019_, new_n1022_, new_n1027_ );
nand g814 ( new_n1029_, new_n1028_, new_n1016_ );
nand g815 ( new_n1030_, new_n1019_, keyIn_0_117, new_n1022_, new_n1027_ );
nand g816 ( new_n1031_, new_n1029_, keyIn_0_119, new_n1015_, new_n1030_ );
not g817 ( new_n1032_, keyIn_0_119 );
nand g818 ( new_n1033_, new_n1029_, new_n1015_, new_n1030_ );
nand g819 ( new_n1034_, new_n1033_, new_n1032_ );
nand g820 ( new_n1035_, new_n1029_, new_n1030_ );
nand g821 ( new_n1036_, new_n1035_, new_n1014_ );
nand g822 ( new_n1037_, new_n1034_, new_n1036_, N219, new_n1031_ );
nand g823 ( new_n1038_, new_n1015_, N228 );
nand g824 ( new_n1039_, new_n913_, N237 );
nand g825 ( new_n1040_, new_n911_, N246 );
nand g826 ( new_n1041_, N91, N210 );
nand g827 ( new_n1042_, new_n569_, N165 );
nand g828 ( new_n1043_, new_n1040_, new_n1041_, new_n1042_ );
not g829 ( new_n1044_, new_n1043_ );
nand g830 ( new_n1045_, new_n1038_, new_n1039_, new_n1044_ );
not g831 ( new_n1046_, new_n1045_ );
nand g832 ( new_n1047_, new_n1037_, new_n1046_ );
nand g833 ( new_n1048_, new_n1047_, new_n1009_ );
nand g834 ( new_n1049_, new_n1037_, keyIn_0_126, new_n1046_ );
nand g835 ( N879, new_n1048_, new_n1049_ );
not g836 ( new_n1051_, keyIn_0_127 );
not g837 ( new_n1052_, keyIn_0_120 );
nand g838 ( new_n1053_, new_n906_, new_n866_ );
nand g839 ( new_n1054_, new_n1053_, keyIn_0_87 );
not g840 ( new_n1055_, keyIn_0_87 );
nand g841 ( new_n1056_, new_n906_, new_n1055_, new_n866_ );
nand g842 ( new_n1057_, new_n1054_, new_n1056_ );
not g843 ( new_n1058_, new_n1057_ );
not g844 ( new_n1059_, keyIn_0_118 );
nand g845 ( new_n1060_, new_n1018_, keyIn_0_113 );
not g846 ( new_n1061_, keyIn_0_113 );
nand g847 ( new_n1062_, new_n1017_, new_n1061_ );
nand g848 ( new_n1063_, new_n1060_, new_n918_, new_n1062_ );
nand g849 ( new_n1064_, new_n1063_, new_n1059_ );
nand g850 ( new_n1065_, new_n1060_, keyIn_0_118, new_n918_, new_n1062_ );
nand g851 ( new_n1066_, new_n1064_, new_n1052_, new_n1058_, new_n1065_ );
nand g852 ( new_n1067_, new_n1064_, new_n1058_, new_n1065_ );
nand g853 ( new_n1068_, new_n1067_, keyIn_0_120 );
nand g854 ( new_n1069_, new_n1064_, new_n1065_ );
nand g855 ( new_n1070_, new_n1069_, new_n1057_ );
nand g856 ( new_n1071_, new_n1068_, new_n1070_, N219, new_n1066_ );
nand g857 ( new_n1072_, new_n1058_, N228 );
nand g858 ( new_n1073_, new_n907_, N237 );
nand g859 ( new_n1074_, new_n905_, N246 );
nand g860 ( new_n1075_, N96, N210 );
nand g861 ( new_n1076_, new_n569_, N171 );
nand g862 ( new_n1077_, new_n1074_, new_n1075_, new_n1076_ );
not g863 ( new_n1078_, new_n1077_ );
nand g864 ( new_n1079_, new_n1072_, new_n1073_, new_n1078_ );
not g865 ( new_n1080_, new_n1079_ );
nand g866 ( new_n1081_, new_n1071_, new_n1080_ );
nand g867 ( new_n1082_, new_n1081_, new_n1051_ );
nand g868 ( new_n1083_, new_n1071_, keyIn_0_127, new_n1080_ );
nand g869 ( N880, new_n1082_, new_n1083_ );
endmodule