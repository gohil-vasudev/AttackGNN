module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX547, WX644, WX645, n3529, WX647, n3527, WX649, n3525, WX653,
         n3521, WX655, n3519, WX657, n3517, WX659, n3515, WX661, n3513, WX663,
         n3511, WX665, n3509, WX667, n3507, WX669, n3505, WX671, n3503, WX673,
         n3501, WX675, n3499, WX677, n3497, WX679, n3495, WX681, n3493, WX683,
         n3491, WX685, n3489, WX689, n3485, WX691, n3483, WX693, n3481, WX695,
         n3479, WX697, n3477, WX699, n3475, WX701, n3473, WX703, n3471, WX705,
         n3469, WX707, n3467, WX708, WX709, WX710, WX711, WX712, WX713, WX714,
         WX715, WX716, WX717, WX718, WX719, WX720, WX721, WX722, WX724, WX725,
         WX726, WX727, WX728, WX729, WX730, WX731, WX732, WX733, WX734, WX735,
         WX736, WX737, WX738, WX739, WX740, WX741, WX742, WX743, WX744, WX745,
         WX746, WX747, WX748, WX749, WX750, WX751, WX752, WX753, WX754, WX755,
         WX756, WX757, WX758, WX760, WX761, WX762, WX763, WX764, WX765, WX766,
         WX767, WX768, WX769, WX770, WX771, WX772, WX773, WX774, WX775, WX776,
         WX777, WX778, WX779, WX780, WX781, WX782, WX783, WX784, WX785, WX786,
         WX787, WX788, WX789, WX790, WX791, WX792, WX793, WX794, WX796, WX797,
         WX798, WX799, WX800, WX801, WX802, WX803, WX804, WX805, WX806, WX807,
         WX808, WX809, WX810, WX811, WX812, WX813, WX814, WX815, WX816, WX817,
         WX818, WX819, WX820, WX821, WX822, WX823, WX824, WX825, WX826, WX827,
         WX828, WX829, WX830, WX832, WX833, WX834, WX835, WX836, WX837, WX838,
         WX839, WX840, WX841, WX842, WX843, WX844, WX845, WX846, WX847, WX848,
         WX849, WX850, WX851, WX852, WX853, WX854, WX855, WX856, WX857, WX858,
         WX859, WX860, WX861, WX862, WX863, WX864, WX865, WX866, WX868, WX869,
         WX870, WX871, WX872, WX873, WX874, WX875, WX876, WX877, WX878, WX879,
         WX880, WX881, WX882, WX883, WX884, WX885, WX886, WX887, WX888, WX889,
         WX890, WX891, WX892, WX893, WX894, WX895, WX896, WX897, WX898, WX899,
         WX1264, DFF_160_n1, WX1266, WX1268, DFF_162_n1, WX1270, WX1272,
         DFF_164_n1, WX1274, DFF_165_n1, WX1276, DFF_166_n1, WX1278,
         DFF_167_n1, WX1280, DFF_168_n1, WX1282, DFF_169_n1, WX1284, WX1286,
         DFF_171_n1, WX1288, DFF_172_n1, WX1290, DFF_173_n1, WX1292,
         DFF_174_n1, WX1294, WX1296, DFF_176_n1, WX1298, DFF_177_n1, WX1300,
         DFF_178_n1, WX1302, WX1304, DFF_180_n1, WX1306, DFF_181_n1, WX1308,
         DFF_182_n1, WX1310, DFF_183_n1, WX1312, DFF_184_n1, WX1314,
         DFF_185_n1, WX1316, DFF_186_n1, WX1318, DFF_187_n1, WX1320,
         DFF_188_n1, WX1322, DFF_189_n1, WX1324, DFF_190_n1, WX1326,
         DFF_191_n1, WX1778, n8702, n8701, n8700, n8699, n8696, n8695, n8694,
         n8693, n8692, n8691, n8690, n8689, n8688, n8687, n8686, n8685, n8684,
         n8683, n8682, n8681, n8680, n8677, n8676, n8675, n8674, n8673, n8672,
         n8671, WX1839, n8670, WX1937, n8669, WX1939, n8668, WX1941, n8667,
         WX1943, n8666, WX1945, n8665, WX1947, n8664, WX1949, n8663, WX1951,
         n8662, WX1953, n8661, WX1955, WX1957, n8658, WX1959, n8657, WX1961,
         n8656, WX1963, n8655, WX1965, n8654, WX1967, n8653, WX1969, WX1970,
         WX1971, WX1972, WX1973, WX1974, WX1975, WX1976, WX1977, WX1978,
         WX1979, WX1980, WX1981, WX1982, WX1983, WX1984, WX1985, WX1986,
         WX1987, WX1988, WX1989, WX1990, WX1991, WX1993, WX1994, WX1995,
         WX1996, WX1997, WX1998, WX1999, WX2000, WX2001, WX2002, WX2003,
         WX2004, WX2005, WX2006, WX2007, WX2008, WX2009, WX2010, WX2011,
         WX2012, WX2013, WX2014, WX2015, WX2016, WX2017, WX2018, WX2019,
         WX2020, WX2021, WX2022, WX2023, WX2024, WX2025, WX2026, WX2027,
         WX2029, WX2030, WX2031, WX2032, WX2033, WX2034, WX2035, WX2036,
         WX2037, WX2038, WX2039, WX2040, WX2041, WX2042, WX2043, WX2044,
         WX2045, WX2046, WX2047, WX2048, WX2049, WX2050, WX2051, WX2052,
         WX2053, WX2054, WX2055, WX2056, WX2057, WX2058, WX2059, WX2060,
         WX2061, WX2062, WX2063, WX2065, WX2066, WX2067, WX2068, WX2069,
         WX2070, WX2071, WX2072, WX2073, WX2074, WX2075, WX2076, WX2077,
         WX2078, WX2079, WX2080, WX2081, WX2082, WX2083, WX2084, WX2085,
         WX2086, WX2087, WX2088, WX2089, WX2090, WX2091, WX2092, WX2093,
         WX2094, WX2095, WX2096, WX2097, WX2098, WX2099, WX2101, WX2102,
         WX2103, WX2104, WX2105, WX2106, WX2107, WX2108, WX2109, WX2110,
         WX2111, WX2112, WX2113, WX2114, WX2115, WX2116, WX2117, WX2118,
         WX2119, WX2120, WX2121, WX2122, WX2123, WX2124, WX2125, WX2126,
         WX2127, WX2128, WX2129, WX2130, WX2131, WX2132, WX2133, WX2134,
         WX2135, WX2137, WX2138, WX2139, WX2140, WX2141, WX2142, WX2143,
         WX2144, WX2145, WX2146, WX2147, WX2148, WX2149, WX2150, WX2151,
         WX2152, WX2153, WX2154, WX2155, WX2156, WX2157, WX2158, WX2159,
         WX2160, WX2161, WX2162, WX2163, WX2164, WX2165, WX2166, WX2167,
         WX2168, WX2169, WX2170, WX2171, WX2173, WX2174, WX2175, WX2176,
         WX2177, WX2178, WX2179, WX2180, WX2181, WX2182, WX2183, WX2184,
         WX2185, WX2186, WX2187, WX2188, WX2189, WX2190, WX2191, WX2192,
         WX2557, DFF_352_n1, WX2559, DFF_353_n1, WX2561, DFF_354_n1, WX2563,
         DFF_355_n1, WX2565, DFF_356_n1, WX2567, DFF_357_n1, WX2569,
         DFF_358_n1, WX2571, WX2573, DFF_360_n1, WX2575, DFF_361_n1, WX2577,
         DFF_362_n1, WX2579, DFF_363_n1, WX2581, DFF_364_n1, WX2583,
         DFF_365_n1, WX2585, DFF_366_n1, WX2587, DFF_367_n1, WX2589,
         DFF_368_n1, WX2591, DFF_369_n1, WX2593, DFF_370_n1, WX2595,
         DFF_371_n1, WX2597, DFF_372_n1, WX2599, DFF_373_n1, WX2601,
         DFF_374_n1, WX2603, DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609,
         DFF_378_n1, WX2611, DFF_379_n1, WX2613, DFF_380_n1, WX2615,
         DFF_381_n1, WX2617, DFF_382_n1, WX2619, DFF_383_n1, WX3071, n8644,
         n8643, n8642, n8641, n8640, n8639, n8638, n8637, n8636, n8635, n8632,
         n8631, n8630, n8629, n8628, n8627, n8626, n8625, n8624, n8623, n8622,
         n8621, n8620, n8619, n8618, n8617, n8616, n8613, WX3132, n8612,
         WX3230, n8611, WX3232, n8610, WX3234, n8609, WX3236, n8608, WX3238,
         n8607, WX3240, n8606, WX3242, n8605, WX3244, n8604, WX3246, n8603,
         WX3248, n8602, WX3250, n8601, WX3252, n8600, WX3254, n8599, WX3256,
         n8598, WX3258, n8597, WX3260, WX3262, WX3263, WX3264, WX3265, WX3266,
         WX3267, WX3268, WX3269, WX3270, WX3271, WX3272, WX3273, WX3274,
         WX3275, WX3276, WX3277, WX3278, WX3279, WX3280, WX3281, WX3282,
         WX3283, WX3284, WX3285, WX3286, WX3287, WX3288, WX3289, WX3290,
         WX3291, WX3292, WX3293, WX3294, WX3295, WX3296, WX3298, WX3299,
         WX3300, WX3301, WX3302, WX3303, WX3304, WX3305, WX3306, WX3307,
         WX3308, WX3309, WX3310, WX3311, WX3312, WX3313, WX3314, WX3315,
         WX3316, WX3317, WX3318, WX3319, WX3320, WX3321, WX3322, WX3323,
         WX3324, WX3325, WX3326, WX3327, n3753, WX3328, WX3329, n3751, WX3330,
         WX3331, n3749, WX3332, WX3334, WX3335, n3745, WX3336, WX3337, n3743,
         WX3338, WX3339, n3741, WX3340, WX3341, WX3342, WX3343, n3737, WX3344,
         WX3345, WX3346, WX3347, n3733, WX3348, WX3349, n3731, WX3350, WX3351,
         n3729, WX3352, WX3353, n3727, WX3354, WX3355, n3725, WX3356, WX3357,
         n3723, WX3358, WX3359, WX3360, WX3361, WX3362, WX3363, WX3364, WX3365,
         WX3366, WX3367, WX3368, WX3370, WX3371, WX3372, WX3373, WX3374,
         WX3375, WX3376, WX3377, WX3378, WX3379, WX3380, WX3381, WX3382,
         WX3383, WX3384, WX3385, WX3386, WX3387, WX3388, WX3389, WX3390,
         WX3391, WX3392, WX3393, WX3394, WX3395, WX3396, WX3397, WX3398,
         WX3399, WX3400, WX3401, WX3402, WX3403, WX3404, WX3406, WX3407,
         WX3408, WX3409, WX3410, WX3411, WX3412, WX3413, WX3414, WX3415,
         WX3416, WX3417, WX3418, WX3419, WX3420, WX3421, WX3422, WX3423,
         WX3424, WX3425, WX3426, WX3427, WX3428, WX3429, WX3430, WX3431,
         WX3432, WX3433, WX3434, WX3435, WX3436, WX3437, WX3438, WX3440,
         WX3441, WX3442, WX3443, WX3444, WX3445, WX3446, WX3447, WX3448,
         WX3449, WX3450, WX3451, WX3452, WX3453, WX3454, WX3455, WX3456,
         WX3457, WX3458, WX3459, WX3460, WX3461, WX3462, WX3463, WX3464,
         WX3465, WX3466, WX3467, WX3468, WX3469, WX3470, WX3471, WX3472,
         WX3474, WX3475, WX3476, WX3477, WX3478, WX3479, WX3480, WX3481,
         WX3482, WX3483, WX3484, WX3485, WX3850, DFF_544_n1, WX3852,
         DFF_545_n1, WX3854, DFF_546_n1, WX3856, DFF_547_n1, WX3858,
         DFF_548_n1, WX3860, DFF_549_n1, WX3862, DFF_550_n1, WX3864,
         DFF_551_n1, WX3866, DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872,
         DFF_555_n1, WX3874, DFF_556_n1, WX3876, DFF_557_n1, WX3878,
         DFF_558_n1, WX3880, DFF_559_n1, WX3882, DFF_560_n1, WX3884,
         DFF_561_n1, WX3886, DFF_562_n1, WX3888, DFF_563_n1, WX3890,
         DFF_564_n1, WX3892, DFF_565_n1, WX3894, DFF_566_n1, WX3896,
         DFF_567_n1, WX3898, DFF_568_n1, WX3900, DFF_569_n1, WX3902,
         DFF_570_n1, WX3904, WX3906, DFF_572_n1, WX3908, DFF_573_n1, WX3910,
         DFF_574_n1, WX3912, DFF_575_n1, WX4364, n8586, n8585, n8584, n8583,
         n8582, n8581, n8580, n8579, n8578, n8577, n8576, n8573, n8572, n8571,
         n8570, n8569, n8568, n8567, n8566, n8565, n8564, n8563, n8562, n8561,
         n8560, n8559, n8558, n8555, WX4425, n8554, WX4523, n8553, WX4525,
         n8552, WX4527, n8551, WX4529, n8550, WX4531, n8549, WX4533, n8548,
         WX4535, n8547, WX4537, n8546, WX4539, n8545, WX4541, n8544, WX4543,
         n8543, WX4545, n8542, WX4547, n8541, WX4549, n8540, WX4551, WX4553,
         n8537, WX4555, WX4556, WX4557, WX4558, WX4559, WX4560, WX4561, WX4562,
         WX4563, WX4564, WX4565, WX4566, WX4567, WX4568, WX4569, WX4570,
         WX4571, WX4572, WX4573, WX4574, WX4575, WX4576, WX4577, WX4578,
         WX4579, WX4580, WX4581, WX4582, WX4583, WX4584, WX4585, WX4587,
         WX4588, WX4589, WX4590, WX4591, WX4592, WX4593, WX4594, WX4595,
         WX4596, WX4597, WX4598, WX4599, WX4600, WX4601, WX4602, WX4603,
         WX4604, WX4605, WX4606, WX4607, WX4608, WX4609, WX4610, WX4611,
         WX4612, WX4613, WX4614, WX4615, WX4616, WX4617, WX4618, WX4619,
         WX4621, WX4622, n3719, WX4623, WX4624, WX4625, WX4626, n3715, WX4627,
         WX4628, WX4629, WX4630, n3711, WX4631, WX4632, n3709, WX4633, WX4634,
         n3707, WX4635, WX4636, n3705, WX4637, WX4638, n3703, WX4639, WX4640,
         n3701, WX4641, WX4642, n3699, WX4643, WX4644, n3697, WX4645, WX4646,
         n3695, WX4647, WX4648, n3693, WX4649, WX4650, WX4651, WX4652, WX4653,
         WX4655, WX4656, WX4657, WX4658, WX4659, WX4660, WX4661, WX4662,
         WX4663, WX4664, WX4665, WX4666, WX4667, WX4668, WX4669, WX4670,
         WX4671, WX4672, WX4673, WX4674, WX4675, WX4676, WX4677, WX4678,
         WX4679, WX4680, WX4681, WX4682, WX4683, WX4684, WX4685, WX4686,
         WX4687, WX4689, WX4690, WX4691, WX4692, WX4693, WX4694, WX4695,
         WX4696, WX4697, WX4698, WX4699, WX4700, WX4701, WX4702, WX4703,
         WX4704, WX4705, WX4706, WX4707, WX4708, WX4709, WX4710, WX4711,
         WX4712, WX4713, WX4714, WX4715, WX4716, WX4717, WX4718, WX4719,
         WX4720, WX4721, WX4723, WX4724, WX4725, WX4726, WX4727, WX4728,
         WX4729, WX4730, WX4731, WX4732, WX4733, WX4734, WX4735, WX4736,
         WX4737, WX4738, WX4739, WX4740, WX4741, WX4742, WX4743, WX4744,
         WX4745, WX4746, WX4747, WX4748, WX4749, WX4750, WX4751, WX4752,
         WX4753, WX4754, WX4755, WX4757, WX4758, WX4759, WX4760, WX4761,
         WX4762, WX4763, WX4764, WX4765, WX4766, WX4767, WX4768, WX4769,
         WX4770, WX4771, WX4772, WX4773, WX4774, WX4775, WX4776, WX4777,
         WX4778, WX5143, DFF_736_n1, WX5145, DFF_737_n1, WX5147, DFF_738_n1,
         WX5149, DFF_739_n1, WX5151, DFF_740_n1, WX5153, WX5155, DFF_742_n1,
         WX5157, DFF_743_n1, WX5159, DFF_744_n1, WX5161, DFF_745_n1, WX5163,
         DFF_746_n1, WX5165, DFF_747_n1, WX5167, DFF_748_n1, WX5169,
         DFF_749_n1, WX5171, DFF_750_n1, WX5173, DFF_751_n1, WX5175,
         DFF_752_n1, WX5177, DFF_753_n1, WX5179, DFF_754_n1, WX5181,
         DFF_755_n1, WX5183, DFF_756_n1, WX5185, DFF_757_n1, WX5187, WX5189,
         DFF_759_n1, WX5191, DFF_760_n1, WX5193, DFF_761_n1, WX5195,
         DFF_762_n1, WX5197, DFF_763_n1, WX5199, DFF_764_n1, WX5201,
         DFF_765_n1, WX5203, DFF_766_n1, WX5205, DFF_767_n1, WX5657, n8528,
         n8527, n8526, n8525, n8524, n8523, n8520, n8519, n8518, n8517, n8516,
         n8515, n8514, n8513, n8512, n8511, n8510, n8509, n8508, n8507, n8506,
         n8505, n8502, n8501, n8500, n8499, n8498, n8497, WX5718, n8496,
         WX5816, n8495, WX5818, n8494, WX5820, n8493, WX5822, n8492, WX5824,
         n8491, WX5826, n8490, WX5828, n8489, WX5830, n8488, WX5832, n8487,
         WX5834, WX5836, n8484, WX5838, n8483, WX5840, n8482, WX5842, n8481,
         WX5844, n8480, WX5846, n8479, WX5848, WX5849, WX5850, WX5851, WX5852,
         WX5853, WX5854, WX5855, WX5856, WX5857, WX5858, WX5859, WX5860,
         WX5861, WX5862, WX5863, WX5864, WX5865, WX5866, WX5867, WX5868,
         WX5870, WX5871, WX5872, WX5873, WX5874, WX5875, WX5876, WX5877,
         WX5878, WX5879, WX5880, WX5881, WX5882, WX5883, WX5884, WX5885,
         WX5886, WX5887, WX5888, WX5889, WX5890, WX5891, WX5892, WX5893,
         WX5894, WX5895, WX5896, WX5897, WX5898, WX5899, WX5900, WX5901,
         WX5902, WX5904, WX5905, WX5906, WX5907, WX5908, WX5909, WX5910,
         WX5911, WX5912, WX5913, n3689, WX5914, WX5915, n3687, WX5916, WX5917,
         n3685, WX5918, WX5919, n3683, WX5920, WX5921, n3681, WX5922, WX5923,
         n3679, WX5924, WX5925, n3677, WX5926, WX5927, n3675, WX5928, WX5929,
         n3673, WX5930, WX5931, n3671, WX5932, WX5933, WX5934, WX5935, n3667,
         WX5936, WX5938, WX5939, n3663, WX5940, WX5941, WX5942, WX5943, n3659,
         WX5944, WX5945, WX5946, WX5947, WX5948, WX5949, WX5950, WX5951,
         WX5952, WX5953, WX5954, WX5955, WX5956, WX5957, WX5958, WX5959,
         WX5960, WX5961, WX5962, WX5963, WX5964, WX5965, WX5966, WX5967,
         WX5968, WX5969, WX5970, WX5972, WX5973, WX5974, WX5975, WX5976,
         WX5977, WX5978, WX5979, WX5980, WX5981, WX5982, WX5983, WX5984,
         WX5985, WX5986, WX5987, WX5988, WX5989, WX5990, WX5991, WX5992,
         WX5993, WX5994, WX5995, WX5996, WX5997, WX5998, WX5999, WX6000,
         WX6001, WX6002, WX6003, WX6004, WX6006, WX6007, WX6008, WX6009,
         WX6010, WX6011, WX6012, WX6013, WX6014, WX6015, WX6016, WX6017,
         WX6018, WX6019, WX6020, WX6021, WX6022, WX6023, WX6024, WX6025,
         WX6026, WX6027, WX6028, WX6029, WX6030, WX6031, WX6032, WX6033,
         WX6034, WX6035, WX6036, WX6037, WX6038, WX6040, WX6041, WX6042,
         WX6043, WX6044, WX6045, WX6046, WX6047, WX6048, WX6049, WX6050,
         WX6051, WX6052, WX6053, WX6054, WX6055, WX6056, WX6057, WX6058,
         WX6059, WX6060, WX6061, WX6062, WX6063, WX6064, WX6065, WX6066,
         WX6067, WX6068, WX6069, WX6070, WX6071, WX6436, WX6438, DFF_929_n1,
         WX6440, DFF_930_n1, WX6442, DFF_931_n1, WX6444, DFF_932_n1, WX6446,
         DFF_933_n1, WX6448, DFF_934_n1, WX6450, DFF_935_n1, WX6452,
         DFF_936_n1, WX6454, DFF_937_n1, WX6456, DFF_938_n1, WX6458,
         DFF_939_n1, WX6460, DFF_940_n1, WX6462, DFF_941_n1, WX6464,
         DFF_942_n1, WX6466, DFF_943_n1, WX6468, DFF_944_n1, WX6470, WX6472,
         DFF_946_n1, WX6474, DFF_947_n1, WX6476, DFF_948_n1, WX6478,
         DFF_949_n1, WX6480, DFF_950_n1, WX6482, DFF_951_n1, WX6484,
         DFF_952_n1, WX6486, DFF_953_n1, WX6488, DFF_954_n1, WX6490,
         DFF_955_n1, WX6492, DFF_956_n1, WX6494, DFF_957_n1, WX6496,
         DFF_958_n1, WX6498, DFF_959_n1, WX6950, n8470, n8467, n8466, n8465,
         n8464, n8463, n8462, n8461, n8460, n8459, n8458, n8457, n8456, n8455,
         n8454, n8453, n8452, n8449, n8448, n8447, n8446, n8445, n8444, n8443,
         n8442, n8441, n8440, n8439, WX7011, n8438, WX7109, n8437, WX7111,
         n8436, WX7113, n8435, WX7115, n8434, WX7117, WX7119, n8431, WX7121,
         n8430, WX7123, n8429, WX7125, n8428, WX7127, n8427, WX7129, n8426,
         WX7131, n8425, WX7133, n8424, WX7135, n8423, WX7137, n8422, WX7139,
         n8421, WX7141, WX7142, WX7143, WX7144, WX7145, WX7146, WX7147, WX7148,
         WX7149, WX7150, WX7151, WX7153, WX7154, WX7155, WX7156, WX7157,
         WX7158, WX7159, WX7160, WX7161, WX7162, WX7163, WX7164, WX7165,
         WX7166, WX7167, WX7168, WX7169, WX7170, WX7171, WX7172, WX7173,
         WX7174, WX7175, WX7176, WX7177, WX7178, WX7179, WX7180, WX7181,
         WX7182, WX7183, WX7184, WX7185, WX7187, WX7188, WX7189, WX7190,
         WX7191, WX7192, WX7193, WX7194, WX7195, WX7196, WX7197, WX7198,
         WX7199, WX7200, WX7201, WX7202, WX7203, WX7204, WX7205, WX7206, n3657,
         WX7207, WX7208, n3655, WX7209, WX7210, n3653, WX7211, WX7212, n3651,
         WX7213, WX7214, n3649, WX7215, WX7216, WX7217, WX7218, n3645, WX7219,
         WX7221, WX7222, n3641, WX7223, WX7224, WX7225, WX7226, n3637, WX7227,
         WX7228, WX7229, WX7230, n3633, WX7231, WX7232, n3631, WX7233, WX7234,
         n3629, WX7235, WX7236, n3627, WX7237, WX7238, WX7239, WX7240, WX7241,
         WX7242, WX7243, WX7244, WX7245, WX7246, WX7247, WX7248, WX7249,
         WX7250, WX7251, WX7252, WX7253, WX7255, WX7256, WX7257, WX7258,
         WX7259, WX7260, WX7261, WX7262, WX7263, WX7264, WX7265, WX7266,
         WX7267, WX7268, WX7269, WX7270, WX7271, WX7272, WX7273, WX7274,
         WX7275, WX7276, WX7277, WX7278, WX7279, WX7280, WX7281, WX7282,
         WX7283, WX7284, WX7285, WX7286, WX7287, WX7289, WX7290, WX7291,
         WX7292, WX7293, WX7294, WX7295, WX7296, WX7297, WX7298, WX7299,
         WX7300, WX7301, WX7302, WX7303, WX7304, WX7305, WX7306, WX7307,
         WX7308, WX7309, WX7310, WX7311, WX7312, WX7313, WX7314, WX7315,
         WX7316, WX7317, WX7318, WX7319, WX7320, WX7321, WX7323, WX7324,
         WX7325, WX7326, WX7327, WX7328, WX7329, WX7330, WX7331, WX7332,
         WX7333, WX7334, WX7335, WX7336, WX7337, WX7338, WX7339, WX7340,
         WX7341, WX7342, WX7343, WX7344, WX7345, WX7346, WX7347, WX7348,
         WX7349, WX7350, WX7351, WX7352, WX7353, WX7354, WX7355, WX7357,
         WX7358, WX7359, WX7360, WX7361, WX7362, WX7363, WX7364, WX7729,
         DFF_1120_n1, WX7731, DFF_1121_n1, WX7733, DFF_1122_n1, WX7735,
         DFF_1123_n1, WX7737, DFF_1124_n1, WX7739, DFF_1125_n1, WX7741,
         DFF_1126_n1, WX7743, DFF_1127_n1, WX7745, DFF_1128_n1, WX7747,
         DFF_1129_n1, WX7749, DFF_1130_n1, WX7751, DFF_1131_n1, WX7753, WX7755,
         DFF_1133_n1, WX7757, DFF_1134_n1, WX7759, DFF_1135_n1, WX7761,
         DFF_1136_n1, WX7763, DFF_1137_n1, WX7765, DFF_1138_n1, WX7767,
         DFF_1139_n1, WX7769, DFF_1140_n1, WX7771, DFF_1141_n1, WX7773,
         DFF_1142_n1, WX7775, DFF_1143_n1, WX7777, DFF_1144_n1, WX7779,
         DFF_1145_n1, WX7781, DFF_1146_n1, WX7783, DFF_1147_n1, WX7785,
         DFF_1148_n1, WX7787, WX7789, DFF_1150_n1, WX7791, DFF_1151_n1, WX8243,
         n8411, n8410, n8409, n8408, n8407, n8406, n8405, n8404, n8403, n8402,
         n8401, n8400, n8399, n8396, n8395, n8394, n8393, n8392, n8391, n8390,
         n8389, n8388, n8387, n8386, n8385, n8384, n8383, n8382, n8381, WX8304,
         WX8402, n8378, WX8404, n8377, WX8406, n8376, WX8408, n8375, WX8410,
         n8374, WX8412, n8373, WX8414, n8372, WX8416, n8371, WX8418, n8370,
         WX8420, n8369, WX8422, n8368, WX8424, n8367, WX8426, n8366, WX8428,
         n8365, WX8430, n8364, WX8432, n8363, WX8434, WX8436, WX8437, WX8438,
         WX8439, WX8440, WX8441, WX8442, WX8443, WX8444, WX8445, WX8446,
         WX8447, WX8448, WX8449, WX8450, WX8451, WX8452, WX8453, WX8454,
         WX8455, WX8456, WX8457, WX8458, WX8459, WX8460, WX8461, WX8462,
         WX8463, WX8464, WX8465, WX8466, WX8467, WX8468, WX8470, WX8471,
         WX8472, WX8473, WX8474, WX8475, WX8476, WX8477, WX8478, WX8479,
         WX8480, WX8481, WX8482, WX8483, WX8484, WX8485, WX8486, WX8487,
         WX8488, WX8489, WX8490, WX8491, WX8492, WX8493, WX8494, WX8495,
         WX8496, WX8497, WX8498, WX8499, WX8500, WX8501, n3623, WX8502, WX8504,
         WX8505, n3619, WX8506, WX8507, WX8508, WX8509, n3615, WX8510, WX8511,
         WX8512, WX8513, n3611, WX8514, WX8515, n3609, WX8516, WX8517, n3607,
         WX8518, WX8519, n3605, WX8520, WX8521, n3603, WX8522, WX8523, n3601,
         WX8524, WX8525, n3599, WX8526, WX8527, n3597, WX8528, WX8529, n3595,
         WX8530, WX8531, WX8532, WX8533, WX8534, WX8535, WX8536, WX8538,
         WX8539, WX8540, WX8541, WX8542, WX8543, WX8544, WX8545, WX8546,
         WX8547, WX8548, WX8549, WX8550, WX8551, WX8552, WX8553, WX8554,
         WX8555, WX8556, WX8557, WX8558, WX8559, WX8560, WX8561, WX8562,
         WX8563, WX8564, WX8565, WX8566, WX8567, WX8568, WX8569, WX8570,
         WX8572, WX8573, WX8574, WX8575, WX8576, WX8577, WX8578, WX8579,
         WX8580, WX8581, WX8582, WX8583, WX8584, WX8585, WX8586, WX8587,
         WX8588, WX8589, WX8590, WX8591, WX8592, WX8593, WX8594, WX8595,
         WX8596, WX8597, WX8598, WX8599, WX8600, WX8601, WX8602, WX8603,
         WX8604, WX8606, WX8607, WX8608, WX8609, WX8610, WX8611, WX8612,
         WX8613, WX8614, WX8615, WX8616, WX8617, WX8618, WX8619, WX8620,
         WX8621, WX8622, WX8623, WX8624, WX8625, WX8626, WX8627, WX8628,
         WX8629, WX8630, WX8631, WX8632, WX8633, WX8634, WX8635, WX8636,
         WX8637, WX8638, WX8640, WX8641, WX8642, WX8643, WX8644, WX8645,
         WX8646, WX8647, WX8648, WX8649, WX8650, WX8651, WX8652, WX8653,
         WX8654, WX8655, WX8656, WX8657, WX9022, DFF_1312_n1, WX9024,
         DFF_1313_n1, WX9026, DFF_1314_n1, WX9028, DFF_1315_n1, WX9030,
         DFF_1316_n1, WX9032, DFF_1317_n1, WX9034, DFF_1318_n1, WX9036, WX9038,
         DFF_1320_n1, WX9040, DFF_1321_n1, WX9042, DFF_1322_n1, WX9044,
         DFF_1323_n1, WX9046, DFF_1324_n1, WX9048, DFF_1325_n1, WX9050,
         DFF_1326_n1, WX9052, DFF_1327_n1, WX9054, DFF_1328_n1, WX9056,
         DFF_1329_n1, WX9058, DFF_1330_n1, WX9060, DFF_1331_n1, WX9062,
         DFF_1332_n1, WX9064, DFF_1333_n1, WX9066, DFF_1334_n1, WX9068,
         DFF_1335_n1, WX9070, WX9072, DFF_1337_n1, WX9074, DFF_1338_n1, WX9076,
         DFF_1339_n1, WX9078, DFF_1340_n1, WX9080, DFF_1341_n1, WX9082,
         DFF_1342_n1, WX9084, DFF_1343_n1, WX9536, n8353, n8352, n8351, n8350,
         n8349, n8348, n8347, n8346, n8343, n8342, n8341, n8340, n8339, n8338,
         n8337, n8336, n8335, n8334, n8333, n8332, n8331, n8330, n8329, n8328,
         n8325, n8324, n8323, n8322, WX9597, n8321, WX9695, n8320, WX9697,
         n8319, WX9699, n8318, WX9701, n8317, WX9703, n8316, WX9705, n8315,
         WX9707, n8314, WX9709, n8313, WX9711, n8312, WX9713, n8311, WX9715,
         n8310, WX9717, WX9719, n8307, WX9721, n8306, WX9723, n8305, WX9725,
         n8304, WX9727, WX9728, WX9729, WX9730, WX9731, WX9732, WX9733, WX9734,
         WX9735, WX9736, WX9737, WX9738, WX9739, WX9740, WX9741, WX9742,
         WX9743, WX9744, WX9745, WX9746, WX9747, WX9748, WX9749, WX9750,
         WX9751, WX9753, WX9754, WX9755, WX9756, WX9757, WX9758, WX9759,
         WX9760, WX9761, WX9762, WX9763, WX9764, WX9765, WX9766, WX9767,
         WX9768, WX9769, WX9770, WX9771, WX9772, WX9773, WX9774, WX9775,
         WX9776, WX9777, WX9778, WX9779, WX9780, WX9781, WX9782, WX9783,
         WX9784, WX9785, WX9787, WX9788, WX9789, WX9790, WX9791, WX9792, n3593,
         WX9793, WX9794, WX9795, WX9796, n3589, WX9797, WX9798, n3587, WX9799,
         WX9800, n3585, WX9801, WX9802, n3583, WX9803, WX9804, n3581, WX9805,
         WX9806, n3579, WX9807, WX9808, n3577, WX9809, WX9810, n3575, WX9811,
         WX9812, n3573, WX9813, WX9814, n3571, WX9815, WX9816, WX9817, WX9818,
         n3567, WX9819, WX9821, WX9822, n3563, WX9823, WX9824, WX9825, WX9826,
         WX9827, WX9828, WX9829, WX9830, WX9831, WX9832, WX9833, WX9834,
         WX9835, WX9836, WX9837, WX9838, WX9839, WX9840, WX9841, WX9842,
         WX9843, WX9844, WX9845, WX9846, WX9847, WX9848, WX9849, WX9850,
         WX9851, WX9852, WX9853, WX9855, WX9856, WX9857, WX9858, WX9859,
         WX9860, WX9861, WX9862, WX9863, WX9864, WX9865, WX9866, WX9867,
         WX9868, WX9869, WX9870, WX9871, WX9872, WX9873, WX9874, WX9875,
         WX9876, WX9877, WX9878, WX9879, WX9880, WX9881, WX9882, WX9883,
         WX9884, WX9885, WX9886, WX9887, WX9889, WX9890, WX9891, WX9892,
         WX9893, WX9894, WX9895, WX9896, WX9897, WX9898, WX9899, WX9900,
         WX9901, WX9902, WX9903, WX9904, WX9905, WX9906, WX9907, WX9908,
         WX9909, WX9910, WX9911, WX9912, WX9913, WX9914, WX9915, WX9916,
         WX9917, WX9918, WX9919, WX9920, WX9921, WX9923, WX9924, WX9925,
         WX9926, WX9927, WX9928, WX9929, WX9930, WX9931, WX9932, WX9933,
         WX9934, WX9935, WX9936, WX9937, WX9938, WX9939, WX9940, WX9941,
         WX9942, WX9943, WX9944, WX9945, WX9946, WX9947, WX9948, WX9949,
         WX9950, WX10315, DFF_1504_n1, WX10317, DFF_1505_n1, WX10319, WX10321,
         DFF_1507_n1, WX10323, DFF_1508_n1, WX10325, DFF_1509_n1, WX10327,
         DFF_1510_n1, WX10329, DFF_1511_n1, WX10331, DFF_1512_n1, WX10333,
         DFF_1513_n1, WX10335, DFF_1514_n1, WX10337, DFF_1515_n1, WX10339,
         DFF_1516_n1, WX10341, DFF_1517_n1, WX10343, DFF_1518_n1, WX10345,
         DFF_1519_n1, WX10347, DFF_1520_n1, WX10349, DFF_1521_n1, WX10351,
         DFF_1522_n1, WX10353, WX10355, DFF_1524_n1, WX10357, DFF_1525_n1,
         WX10359, DFF_1526_n1, WX10361, DFF_1527_n1, WX10363, DFF_1528_n1,
         WX10365, DFF_1529_n1, WX10367, DFF_1530_n1, WX10369, DFF_1531_n1,
         WX10371, DFF_1532_n1, WX10373, DFF_1533_n1, WX10375, DFF_1534_n1,
         WX10377, DFF_1535_n1, WX10829, n8295, n8294, n8293, n8290, n8289,
         n8288, n8287, n8286, n8285, n8284, n8283, n8282, n8281, n8280, n8279,
         n8278, n8277, n8276, n8275, n8272, n8271, n8270, n8269, n8268, n8267,
         n8266, n8265, n8264, WX10890, n8263, n8262, n8261, n8260, n8259,
         n8258, n8257, n8254, n8253, n8252, n8251, n8250, n8249, n8248, n8247,
         n8246, WX11021, WX11023, WX11025, WX11027, WX11029, WX11031, WX11033,
         WX11037, WX11039, WX11041, WX11043, WX11045, WX11047, WX11049,
         WX11051, WX11052, WX11053, WX11054, WX11055, WX11056, WX11057,
         WX11058, WX11059, WX11060, WX11061, WX11062, WX11063, WX11064,
         WX11065, WX11066, WX11067, WX11068, WX11070, WX11071, WX11072,
         WX11073, WX11074, WX11075, WX11076, WX11077, WX11078, WX11079,
         WX11080, WX11081, WX11082, WX11083, WX11084, WX11085, WX11086,
         WX11087, WX11088, WX11089, WX11090, WX11091, WX11092, WX11093,
         WX11094, WX11095, WX11096, WX11097, WX11098, WX11099, WX11100,
         WX11101, WX11102, WX11104, WX11105, WX11106, WX11107, WX11108,
         WX11109, WX11110, WX11111, WX11112, WX11113, WX11114, WX11115,
         WX11116, WX11117, WX11118, WX11119, WX11120, WX11121, WX11122,
         WX11123, WX11124, WX11125, WX11126, WX11127, WX11128, WX11129,
         WX11130, WX11131, WX11132, WX11133, WX11134, WX11135, WX11136,
         WX11138, WX11139, WX11140, WX11141, WX11142, WX11143, WX11144,
         WX11145, WX11146, WX11147, WX11148, WX11149, WX11150, WX11151,
         WX11152, WX11153, WX11154, WX11155, WX11156, WX11157, WX11158,
         WX11159, WX11160, WX11161, WX11162, WX11163, WX11164, WX11165,
         WX11166, WX11167, WX11168, WX11169, WX11170, WX11172, WX11173,
         WX11174, WX11175, WX11176, WX11177, WX11178, WX11179, WX11180,
         WX11181, WX11182, WX11183, WX11184, WX11185, WX11186, WX11187,
         WX11188, WX11189, WX11190, WX11191, WX11192, WX11193, WX11194,
         WX11195, WX11196, WX11197, WX11198, WX11199, WX11200, WX11201,
         WX11202, WX11203, WX11204, WX11206, WX11207, WX11208, WX11209,
         WX11210, WX11211, WX11212, WX11213, WX11214, WX11215, WX11216,
         WX11217, WX11218, WX11219, WX11220, WX11221, WX11222, WX11223,
         WX11224, WX11225, WX11226, WX11227, WX11228, WX11229, WX11230,
         WX11231, WX11232, WX11233, WX11234, WX11235, WX11236, WX11237,
         WX11238, WX11240, WX11241, WX11242, WX11243, WX11608, DFF_1696_n1,
         WX11610, DFF_1697_n1, WX11612, DFF_1698_n1, WX11614, WX11616,
         DFF_1700_n1, WX11618, DFF_1701_n1, WX11620, DFF_1702_n1, WX11622,
         DFF_1703_n1, WX11624, DFF_1704_n1, WX11626, DFF_1705_n1, WX11628,
         WX11630, DFF_1707_n1, WX11632, DFF_1708_n1, WX11634, DFF_1709_n1,
         WX11636, WX11638, WX11640, DFF_1712_n1, WX11642, DFF_1713_n1, WX11644,
         DFF_1714_n1, WX11646, DFF_1715_n1, WX11648, DFF_1716_n1, WX11650,
         DFF_1717_n1, WX11652, DFF_1718_n1, WX11654, DFF_1719_n1, WX11656,
         DFF_1720_n1, WX11658, DFF_1721_n1, WX11660, DFF_1722_n1, WX11662,
         DFF_1723_n1, WX11664, DFF_1724_n1, WX11666, DFF_1725_n1, WX11668,
         DFF_1726_n1, WX11670, n2245, n2153, n3278, n2152, Tj_OUT1, Tj_OUT2,
         Tj_OUT3, Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8,
         Tj_OUT5678, Tj_Trigger, Stage4, Stage1_1, Stage1_2, Stage1_3,
         Stage1_4, Stage1, Stage2_i, Stage2_7, Stage2_8, Stage2_9, Stage2_10,
         Stage2, Stage3_i, Stage3_12, Stage3_13, Stage3_14, Stage3_15,
         Stage4_i, Stage4_17, Stage4_18, Stage4_19, Stage4_20, Stage4_21, n1,
         n43, n46, n49, n53, n56, n59, n62, n65, n68, n71, n74, n77, n80, n83,
         n86, n89, n92, n95, n98, n101, n104, n108, n111, n114, n117, n120,
         n123, n126, n129, n132, n135, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n2010, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2339, n2340, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9561, n9563, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9578,
         n9580, n9582, n9592, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9604, n9607, n9609, n9611, n9617, n9618, n9619, n9620,
         n9622, n9624, n9626, n9627, n9628, n9629, n9639, n9641, n9643, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9656, n9657,
         n9659, n9665, n9671, n9673, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9686, n9688, n9690, n9699, n9700, n9701,
         n9703, n9704, n9706, n9707, n9708, n9709, n9710, n9715, n9719, n9723,
         n9730, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, U3558_n1, U3871_n1, U3991_n1, U5716_n1, U5717_n1, U5718_n1,
         U5719_n1, U5720_n1, U5721_n1, U5722_n1, U5723_n1, U5724_n1, U5725_n1,
         U5726_n1, U5727_n1, U5728_n1, U5729_n1, U5730_n1, U5731_n1, U5732_n1,
         U5733_n1, U5734_n1, U5735_n1, U5736_n1, U5737_n1, U5738_n1, U5739_n1,
         U5740_n1, U5741_n1, U5742_n1, U5743_n1, U5744_n1, U5745_n1, U5746_n1,
         U5747_n1, U5748_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1, U5753_n1,
         U5754_n1, U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1, U5760_n1,
         U5761_n1, U5762_n1, U5763_n1, U5764_n1, U5765_n1, U5766_n1, U5767_n1,
         U5768_n1, U5769_n1, U5770_n1, U5771_n1, U5772_n1, U5773_n1, U5774_n1,
         U5775_n1, U5776_n1, U5777_n1, U5778_n1, U5779_n1, U5780_n1, U5781_n1,
         U5782_n1, U5783_n1, U5784_n1, U5785_n1, U5786_n1, U5787_n1, U5788_n1,
         U5789_n1, U5790_n1, U5791_n1, U5792_n1, U5793_n1, U5794_n1, U5795_n1,
         U5796_n1, U5797_n1, U5798_n1, U5799_n1, U5800_n1, U5801_n1, U5802_n1,
         U5803_n1, U5804_n1, U5805_n1, U5806_n1, U5807_n1, U5808_n1, U5809_n1,
         U5810_n1, U5811_n1, U5812_n1, U5813_n1, U5814_n1, U5815_n1, U5816_n1,
         U5817_n1, U5818_n1, U5819_n1, U5820_n1, U5821_n1, U5822_n1, U5823_n1,
         U5824_n1, U5825_n1, U5826_n1, U5827_n1, U5828_n1, U5829_n1, U5830_n1,
         U5831_n1, U5832_n1, U5833_n1, U5834_n1, U5835_n1, U5836_n1, U5837_n1,
         U5838_n1, U5839_n1, U5840_n1, U5841_n1, U5842_n1, U5843_n1, U5844_n1,
         U5845_n1, U5846_n1, U5847_n1, U5848_n1, U5849_n1, U5850_n1, U5851_n1,
         U5852_n1, U5853_n1, U5854_n1, U5855_n1, U5856_n1, U5857_n1, U5858_n1,
         U5859_n1, U5860_n1, U5861_n1, U5862_n1, U5863_n1, U5864_n1, U5865_n1,
         U5866_n1, U5867_n1, U5868_n1, U5869_n1, U5870_n1, U5871_n1, U5872_n1,
         U5873_n1, U5874_n1, U5875_n1, U5876_n1, U5877_n1, U5878_n1, U5879_n1,
         U5880_n1, U5881_n1, U5882_n1, U5883_n1, U5884_n1, U5885_n1, U5886_n1,
         U5887_n1, U5888_n1, U5889_n1, U5890_n1, U5891_n1, U5892_n1, U5893_n1,
         U5894_n1, U5895_n1, U5896_n1, U5897_n1, U5898_n1, U5899_n1, U5900_n1,
         U5901_n1, U5902_n1, U5903_n1, U5904_n1, U5905_n1, U5906_n1, U5907_n1,
         U5908_n1, U5909_n1, U5910_n1, U5911_n1, U5912_n1, U5913_n1, U5914_n1,
         U5915_n1, U5916_n1, U5917_n1, U5918_n1, U5919_n1, U5920_n1, U5921_n1,
         U5922_n1, U5923_n1, U5924_n1, U5925_n1, U5926_n1, U5927_n1, U5928_n1,
         U5929_n1, U5930_n1, U5931_n1, U5932_n1, U5933_n1, U5934_n1, U5935_n1,
         U5936_n1, U5937_n1, U5938_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1,
         U5943_n1, U5944_n1, U5945_n1, U5946_n1, U5947_n1, U5948_n1, U5949_n1,
         U5950_n1, U5951_n1, U5952_n1, U5953_n1, U5954_n1, U5955_n1, U5956_n1,
         U5957_n1, U5958_n1, U5959_n1, U5960_n1, U5961_n1, U5962_n1, U5963_n1,
         U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1, U5969_n1, U5970_n1,
         U5971_n1, U5972_n1, U5973_n1, U5974_n1, U5975_n1, U5976_n1, U5977_n1,
         U5978_n1, U5979_n1, U5980_n1, U5981_n1, U5982_n1, U5983_n1, U5984_n1,
         U5985_n1, U5986_n1, U5987_n1, U5988_n1, U5989_n1, U5990_n1, U5991_n1,
         U5992_n1, U5993_n1, U5994_n1, U5995_n1, U5996_n1, U5997_n1, U5998_n1,
         U5999_n1, U6000_n1, U6001_n1, U6002_n1, U6003_n1, U6004_n1, U6005_n1,
         U6006_n1, U6007_n1, U6008_n1, U6009_n1, U6010_n1, U6011_n1, U6012_n1,
         U6013_n1, U6014_n1, U6015_n1, U6016_n1, U6017_n1, U6018_n1, U6019_n1,
         U6020_n1, U6021_n1, U6022_n1, U6023_n1, U6024_n1, U6025_n1, U6026_n1,
         U6027_n1, U6028_n1, U6029_n1, U6030_n1, U6031_n1, U6032_n1, U6033_n1,
         U6034_n1, U6035_n1, U6036_n1, U6037_n1, U6038_n1, U6039_n1, U6040_n1,
         U6041_n1, U6042_n1, U6043_n1, U6044_n1, U6045_n1, U6046_n1, U6047_n1,
         U6048_n1, U6049_n1, U6050_n1, U6051_n1, U6052_n1, U6053_n1, U6054_n1,
         U6055_n1, U6056_n1, U6057_n1, U6058_n1, U6059_n1, U6060_n1, U6061_n1,
         U6062_n1, U6063_n1, U6064_n1, U6065_n1, U6066_n1, U6067_n1, U6068_n1,
         U6069_n1, U6070_n1, U6071_n1, U6072_n1, U6073_n1, U6074_n1, U6075_n1,
         U6076_n1, U6077_n1, U6078_n1, U6079_n1, U6080_n1, U6081_n1, U6082_n1,
         U6083_n1, U6084_n1, U6085_n1, U6086_n1, U6087_n1, U6088_n1, U6089_n1,
         U6090_n1, U6091_n1, U6092_n1, U6093_n1, U6094_n1, U6095_n1, U6096_n1,
         U6097_n1, U6098_n1, U6099_n1, U6100_n1, U6101_n1, U6102_n1, U6103_n1,
         U6104_n1, U6105_n1, U6106_n1, U6107_n1, U6108_n1, U6109_n1, U6110_n1,
         U6111_n1, U6112_n1, U6113_n1, U6114_n1, U6115_n1, U6116_n1, U6117_n1,
         U6118_n1, U6119_n1, U6120_n1, U6121_n1, U6122_n1, U6123_n1, U6124_n1,
         U6125_n1, U6126_n1, U6127_n1, U6128_n1, U6129_n1, U6130_n1, U6131_n1,
         U6132_n1, U6133_n1, U6134_n1, U6135_n1, U6136_n1, U6137_n1, U6138_n1,
         U6139_n1, U6140_n1, U6141_n1, U6142_n1, U6143_n1, U6144_n1, U6145_n1,
         U6146_n1, U6147_n1, U6148_n1, U6149_n1, U6150_n1, U6151_n1, U6152_n1,
         U6153_n1, U6154_n1, U6155_n1, U6156_n1, U6157_n1, U6158_n1, U6159_n1,
         U6160_n1, U6161_n1, U6162_n1, U6163_n1, U6164_n1, U6165_n1, U6166_n1,
         U6167_n1, U6168_n1, U6169_n1, U6170_n1, U6171_n1, U6172_n1, U6173_n1,
         U6174_n1, U6175_n1, U6176_n1, U6177_n1, U6178_n1, U6179_n1, U6180_n1,
         U6181_n1, U6182_n1, U6183_n1, U6184_n1, U6185_n1, U6186_n1, U6187_n1,
         U6188_n1, U6189_n1, U6190_n1, U6191_n1, U6192_n1, U6193_n1, U6194_n1,
         U6195_n1, U6196_n1, U6197_n1, U6198_n1, U6199_n1, U6200_n1, U6201_n1,
         U6202_n1, U6203_n1, U6204_n1, U6205_n1, U6206_n1, U6207_n1, U6208_n1,
         U6209_n1, U6210_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1,
         U6216_n1, U6217_n1, U6218_n1, U6219_n1, U6220_n1, U6221_n1, U6222_n1,
         U6223_n1, U6224_n1, U6225_n1, U6226_n1, U6227_n1, U6228_n1, U6229_n1,
         U6230_n1, U6231_n1, U6232_n1, U6233_n1, U6234_n1, U6235_n1, U6236_n1,
         U6237_n1, U6238_n1, U6239_n1, U6240_n1, U6241_n1, U6242_n1, U6243_n1,
         U6244_n1, U6245_n1, U6246_n1, U6247_n1, U6248_n1, U6249_n1, U6250_n1,
         U6251_n1, U6252_n1, U6253_n1, U6254_n1, U6255_n1, U6256_n1, U6257_n1,
         U6258_n1, U6259_n1, U6260_n1, U6261_n1, U6262_n1, U6263_n1, U6264_n1,
         U6265_n1, U6266_n1, U6267_n1, U6268_n1, U6269_n1, U6270_n1, U6271_n1,
         U6272_n1, U6273_n1, U6274_n1, U6275_n1, U6276_n1, U6277_n1, U6278_n1,
         U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1,
         U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1,
         U6293_n1, U6294_n1, U6295_n1, U6296_n1, U6297_n1, U6298_n1, U6299_n1,
         U6300_n1, U6301_n1, U6302_n1, U6303_n1, U6304_n1, U6305_n1, U6306_n1,
         U6307_n1, U6308_n1, U6309_n1, U6310_n1, U6311_n1, U6312_n1, U6313_n1,
         U6314_n1, U6315_n1, U6316_n1, U6317_n1, U6318_n1, U6319_n1, U6320_n1,
         U6321_n1, U6322_n1, U6323_n1, U6324_n1, U6325_n1, U6326_n1, U6327_n1,
         U6328_n1, U6329_n1, U6330_n1, U6331_n1, U6332_n1, U6333_n1, U6334_n1,
         U6335_n1, U6336_n1, U6337_n1, U6338_n1, U6339_n1, U6340_n1, U6341_n1,
         U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1,
         U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1,
         U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1,
         U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1,
         U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6376_n1,
         U6377_n1, U6378_n1, U6379_n1, U6380_n1, U6381_n1, U6382_n1, U6383_n1,
         U6384_n1, U6385_n1, U6386_n1, U6387_n1, U6388_n1, U6389_n1, U6390_n1,
         U6391_n1, U6392_n1, U6393_n1, U6394_n1, U6395_n1, U6396_n1, U6397_n1,
         U6398_n1, U6399_n1, U6400_n1, U6401_n1, U6402_n1, U6403_n1, U6404_n1,
         U6405_n1, U6406_n1, U6407_n1, U6408_n1, U6409_n1, U6410_n1, U6411_n1,
         U6412_n1, U6413_n1, U6414_n1, U6415_n1, U6416_n1, U6417_n1, U6418_n1,
         U6419_n1, U6420_n1, U6421_n1, U6422_n1, U6423_n1, U6424_n1, U6425_n1,
         U6426_n1, U6427_n1, U6428_n1, U6429_n1, U6430_n1, U6431_n1, U6432_n1,
         U6433_n1, U6434_n1, U6435_n1, U6436_n1, U6437_n1, U6438_n1, U6439_n1,
         U6440_n1, U6441_n1, U6442_n1, U6443_n1, U6444_n1, U6445_n1, U6446_n1,
         U6447_n1, U6448_n1, U6449_n1, U6450_n1, U6451_n1, U6452_n1, U6453_n1,
         U6454_n1, U6455_n1, U6456_n1, U6457_n1, U6458_n1, U6459_n1, U6460_n1,
         U6461_n1, U6462_n1, U6463_n1, U6464_n1, U6465_n1, U6466_n1, U6467_n1,
         U6468_n1, U6469_n1, U6470_n1, U6471_n1, U6472_n1, U6473_n1, U6474_n1,
         U6475_n1, U6476_n1, U6477_n1, U6478_n1, U6479_n1, U6480_n1, U6481_n1,
         U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n10026), .CLK(n10333), 
        .Q(WX485), .QN(n9487) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n10167), .CLK(n10335), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n10167), .CLK(n10335), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n10167), .CLK(n10335), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n10167), .CLK(n10335), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n10167), .CLK(n10335), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n10167), .CLK(n10335), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n10167), .CLK(n10335), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n10167), .CLK(n10335), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n10025), .CLK(n10334), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n10022), .CLK(n10334), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n10023), .CLK(n10334), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n10026), .CLK(n10334), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n10027), .CLK(n10334), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(test_se), .CLK(n10334), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n10028), .CLK(n10334), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n10024), .CLK(n10334), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n10025), .CLK(n10334), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n10022), .CLK(n10334), 
        .Q(WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n10023), .CLK(n10334), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n10026), .CLK(n10334), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(test_se), .CLK(n10333), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n10028), .CLK(n10333), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n10024), .CLK(n10333), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n10025), .CLK(n10333), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n10022), .CLK(n10333), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n10023), .CLK(n10333), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n10026), .CLK(n10333), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n10024), .CLK(n10333), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n10025), .CLK(n10333), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n10022), .CLK(n10333), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(n1), .SI(WX545), .SE(n10023), .CLK(n10333), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n10167), .CLK(n10335), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(n43), .SI(WX645), .SE(n10167), .CLK(n10335), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(n46), .SI(WX647), .SE(n10167), .CLK(n10335), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(n49), .SI(WX649), .SE(n10167), .CLK(n10335), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(n53), .SI(test_si3), .SE(n10166), .CLK(n10336), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(n56), .SI(WX653), .SE(n10166), .CLK(n10336), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(n59), .SI(WX655), .SE(n10166), .CLK(n10336), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(n62), .SI(WX657), .SE(n10166), .CLK(n10336), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(n65), .SI(WX659), .SE(n10166), .CLK(n10336), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(n68), .SI(WX661), .SE(n10166), .CLK(n10336), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(n71), .SI(WX663), .SE(n10165), .CLK(n10337), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(n74), .SI(WX665), .SE(n10165), .CLK(n10337), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(n77), .SI(WX667), .SE(n10165), .CLK(n10337), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(n80), .SI(WX669), .SE(n10165), .CLK(n10337), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(n83), .SI(WX671), .SE(n10165), .CLK(n10337), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(n86), .SI(WX673), .SE(n10164), .CLK(n10338), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(n89), .SI(WX675), .SE(n10164), .CLK(n10338), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(n92), .SI(WX677), .SE(n10164), .CLK(n10338), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(n95), .SI(WX679), .SE(n10163), .CLK(n10339), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(n98), .SI(WX681), .SE(n10163), .CLK(n10339), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(n101), .SI(WX683), .SE(n10163), .CLK(n10339), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(n104), .SI(WX685), .SE(n10162), .CLK(n10340), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(n108), .SI(test_si4), .SE(n10162), .CLK(n10340), 
        .Q(WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(n111), .SI(WX689), .SE(n10162), .CLK(n10340), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(n114), .SI(WX691), .SE(n10161), .CLK(n10341), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(n117), .SI(WX693), .SE(n10161), .CLK(n10341), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(n120), .SI(WX695), .SE(n10161), .CLK(n10341), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(n123), .SI(WX697), .SE(n10160), .CLK(n10342), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(n126), .SI(WX699), .SE(n10160), .CLK(n10342), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(n129), .SI(WX701), .SE(n10160), .CLK(n10342), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(n132), .SI(WX703), .SE(n10159), .CLK(n10343), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(n135), .SI(WX705), .SE(n10159), .CLK(n10343), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n10159), .CLK(n10343), .Q(
        WX709), .QN(n9811) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n10158), .CLK(n10344), .Q(
        WX711), .QN(n9737) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n10158), .CLK(n10344), .Q(
        WX713), .QN(n9748) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n10166), .CLK(n10336), .Q(
        WX715), .QN(n9757) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n10166), .CLK(n10336), .Q(
        WX717), .QN(n9763) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n10166), .CLK(n10336), .Q(
        WX719), .QN(n9766) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n10166), .CLK(n10336), .Q(
        WX721), .QN(n9775) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n10166), .CLK(n10336), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n10166), .CLK(n10336), 
        .Q(WX725), .QN(n9786) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n10165), .CLK(n10337), .Q(
        WX727), .QN(n9798) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n10165), .CLK(n10337), .Q(
        WX729), .QN(n9804) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n10165), .CLK(n10337), .Q(
        WX731) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n10165), .CLK(n10337), .Q(
        WX733), .QN(n9745) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n10165), .CLK(n10337), .Q(
        WX735), .QN(n9760) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n10164), .CLK(n10338), .Q(
        WX737), .QN(n9772) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n10164), .CLK(n10338), .Q(
        WX739), .QN(n9787) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n10164), .CLK(n10338), .Q(
        WX741), .QN(n9801) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n10164), .CLK(n10338), .Q(
        WX743), .QN(n9816) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n10163), .CLK(n10339), .Q(
        WX745), .QN(n9751) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n10163), .CLK(n10339), .Q(
        WX747), .QN(n9778) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n10163), .CLK(n10339), .Q(
        WX749), .QN(n9824) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n10162), .CLK(n10340), .Q(
        WX751), .QN(n9769) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n10162), .CLK(n10340), .Q(
        WX753), .QN(n9779) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n10162), .CLK(n10340), .Q(
        WX755), .QN(n9791) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n10161), .CLK(n10341), .Q(
        WX757), .QN(n9819) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n10161), .CLK(n10341), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n10161), .CLK(n10341), 
        .Q(WX761), .QN(n9794) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n10160), .CLK(n10342), .Q(
        WX763), .QN(n9797) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n10160), .CLK(n10342), .Q(
        WX765), .QN(n9742) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n10160), .CLK(n10342), .Q(
        WX767), .QN(n9817) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n10159), .CLK(n10343), .Q(
        WX769), .QN(n9753) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n10159), .CLK(n10343), .Q(
        WX771), .QN(n9825) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n10159), .CLK(n10343), .Q(
        WX773), .QN(n9812) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n10158), .CLK(n10344), .Q(
        WX775), .QN(n9738) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n10158), .CLK(n10344), .Q(
        WX777), .QN(n9746) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n10158), .CLK(n10344), .Q(
        WX779), .QN(n9755) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n10158), .CLK(n10344), .Q(
        WX781), .QN(n9761) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n10158), .CLK(n10344), .Q(
        WX783), .QN(n9764) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n10157), .CLK(n10345), .Q(
        WX785), .QN(n9773) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n10157), .CLK(n10345), .Q(
        WX787), .QN(n9782) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n10157), .CLK(n10345), .Q(
        WX789), .QN(n9784) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n10157), .CLK(n10345), .Q(
        WX791), .QN(n9799) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n10157), .CLK(n10345), .Q(
        WX793), .QN(n9805) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n10157), .CLK(n10345), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n10165), .CLK(n10337), 
        .Q(WX797), .QN(n9743) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n10165), .CLK(n10337), .Q(
        WX799), .QN(n9758) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n10164), .CLK(n10338), .Q(
        WX801), .QN(n9770) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n10164), .CLK(n10338), .Q(
        WX803), .QN(n9788) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n10164), .CLK(n10338), .Q(
        WX805), .QN(n9802) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n10164), .CLK(n10338), .Q(
        WX807), .QN(n9814) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n10163), .CLK(n10339), .Q(
        WX809), .QN(n9749) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n10163), .CLK(n10339), .Q(
        WX811), .QN(n9776) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n10163), .CLK(n10339), .Q(
        WX813), .QN(n9822) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n10162), .CLK(n10340), .Q(
        WX815), .QN(n9767) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n10162), .CLK(n10340), .Q(
        WX817), .QN(n9780) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n10162), .CLK(n10340), .Q(
        WX819), .QN(n9789) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n10161), .CLK(n10341), .Q(
        WX821), .QN(n9820) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n10161), .CLK(n10341), .Q(
        WX823), .QN(n9807) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n10161), .CLK(n10341), .Q(
        WX825), .QN(n9792) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n10160), .CLK(n10342), .Q(
        WX827), .QN(n9795) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n10160), .CLK(n10342), .Q(
        WX829), .QN(n9740) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n10160), .CLK(n10342), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n10159), .CLK(n10343), 
        .Q(WX833) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n10159), .CLK(n10343), .Q(
        WX835), .QN(n9826) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n10159), .CLK(n10343), .Q(
        WX837), .QN(n9813) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n10158), .CLK(n10344), .Q(
        WX839), .QN(n9739) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n10158), .CLK(n10344), .Q(
        WX841), .QN(n9747) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n10158), .CLK(n10344), .Q(
        WX843), .QN(n9756) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n10158), .CLK(n10344), .Q(
        WX845), .QN(n9762) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n10158), .CLK(n10344), .Q(
        WX847), .QN(n9765) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n10157), .CLK(n10345), .Q(
        WX849), .QN(n9774) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n10157), .CLK(n10345), .Q(
        WX851), .QN(n9783) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n10157), .CLK(n10345), .Q(
        WX853), .QN(n9785) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n10157), .CLK(n10345), .Q(
        WX855), .QN(n9800) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n10157), .CLK(n10345), .Q(
        WX857), .QN(n9806) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n10157), .CLK(n10345), .Q(
        WX859), .QN(n9809) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n10156), .CLK(n10346), .Q(
        WX861), .QN(n9744) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n10156), .CLK(n10346), .Q(
        WX863), .QN(n9759) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n10156), .CLK(n10346), .Q(
        WX865), .QN(n9771) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n10156), .CLK(n10346), .Q(
        test_so8), .QN(n9851) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n10164), .CLK(n10338), 
        .Q(WX869), .QN(n9803) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n10163), .CLK(n10339), .Q(
        WX871), .QN(n9815) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n10163), .CLK(n10339), .Q(
        WX873), .QN(n9750) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n10163), .CLK(n10339), .Q(
        WX875), .QN(n9777) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n10162), .CLK(n10340), .Q(
        WX877), .QN(n9823) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n10162), .CLK(n10340), .Q(
        WX879), .QN(n9768) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n10162), .CLK(n10340), .Q(
        WX881), .QN(n9781) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n10161), .CLK(n10341), .Q(
        WX883), .QN(n9790) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n10161), .CLK(n10341), .Q(
        WX885), .QN(n9821) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n10161), .CLK(n10341), .Q(
        WX887), .QN(n9808) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n10160), .CLK(n10342), .Q(
        WX889), .QN(n9793) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n10160), .CLK(n10342), .Q(
        WX891), .QN(n9796) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n10160), .CLK(n10342), .Q(
        WX893), .QN(n9741) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n10159), .CLK(n10343), .Q(
        WX895) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n10159), .CLK(n10343), .Q(
        WX897), .QN(n9752) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n10159), .CLK(n10343), .Q(
        WX899), .QN(n9827) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n10030), .CLK(n10475), 
        .Q(CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n10030), .CLK(
        n10475), .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n10030), .CLK(n10475), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n10030), .CLK(
        n10475), .Q(CRC_OUT_9_3) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n10030), .CLK(
        n10475), .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n10030), .CLK(
        n10475), .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n10030), .CLK(
        n10475), .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n10030), .CLK(
        n10475), .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_10) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_15) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n10029), .CLK(
        n10476), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n10029), .CLK(
        n10476), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n10156), .CLK(n10346), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n10156), .CLK(
        n10346), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n10156), .CLK(
        n10346), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n10156), .CLK(
        n10346), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n10156), .CLK(
        n10346), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n10156), .CLK(
        n10346), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n10156), .CLK(
        n10346), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n10156), .CLK(
        n10346), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n10024), .CLK(
        n10347), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n10028), .CLK(
        n10347), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(test_se), .CLK(
        n10347), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n10027), .CLK(
        n10347), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n281), .SI(CRC_OUT_9_31), .SE(n10026), .CLK(n10347), .Q(WX1778), .QN(n9495) );
  SDFFX1 DFF_193_Q_reg ( .D(n282), .SI(WX1778), .SE(n10154), .CLK(n10349), .Q(
        n8702) );
  SDFFX1 DFF_194_Q_reg ( .D(n283), .SI(n8702), .SE(n10154), .CLK(n10349), .Q(
        n8701) );
  SDFFX1 DFF_195_Q_reg ( .D(n284), .SI(n8701), .SE(n10154), .CLK(n10349), .Q(
        n8700) );
  SDFFX1 DFF_196_Q_reg ( .D(n285), .SI(n8700), .SE(n10154), .CLK(n10349), .Q(
        n8699) );
  SDFFX1 DFF_197_Q_reg ( .D(n286), .SI(n8699), .SE(n10154), .CLK(n10349), .Q(
        test_so11) );
  SDFFX1 DFF_198_Q_reg ( .D(n287), .SI(test_si12), .SE(n10154), .CLK(n10349), 
        .Q(n8696) );
  SDFFX1 DFF_199_Q_reg ( .D(n288), .SI(n8696), .SE(n10154), .CLK(n10349), .Q(
        n8695) );
  SDFFX1 DFF_200_Q_reg ( .D(n289), .SI(n8695), .SE(n10154), .CLK(n10349), .Q(
        n8694) );
  SDFFX1 DFF_201_Q_reg ( .D(n290), .SI(n8694), .SE(n10154), .CLK(n10349), .Q(
        n8693) );
  SDFFX1 DFF_202_Q_reg ( .D(n291), .SI(n8693), .SE(n10154), .CLK(n10349), .Q(
        n8692) );
  SDFFX1 DFF_203_Q_reg ( .D(n292), .SI(n8692), .SE(n10154), .CLK(n10349), .Q(
        n8691) );
  SDFFX1 DFF_204_Q_reg ( .D(n293), .SI(n8691), .SE(n10154), .CLK(n10349), .Q(
        n8690) );
  SDFFX1 DFF_205_Q_reg ( .D(n294), .SI(n8690), .SE(n10155), .CLK(n10348), .Q(
        n8689) );
  SDFFX1 DFF_206_Q_reg ( .D(n295), .SI(n8689), .SE(n10155), .CLK(n10348), .Q(
        n8688) );
  SDFFX1 DFF_207_Q_reg ( .D(n296), .SI(n8688), .SE(n10155), .CLK(n10348), .Q(
        n8687) );
  SDFFX1 DFF_208_Q_reg ( .D(n297), .SI(n8687), .SE(n10155), .CLK(n10348), .Q(
        n8686) );
  SDFFX1 DFF_209_Q_reg ( .D(n298), .SI(n8686), .SE(n10155), .CLK(n10348), .Q(
        n8685) );
  SDFFX1 DFF_210_Q_reg ( .D(n299), .SI(n8685), .SE(n10155), .CLK(n10348), .Q(
        n8684) );
  SDFFX1 DFF_211_Q_reg ( .D(n300), .SI(n8684), .SE(n10155), .CLK(n10348), .Q(
        n8683) );
  SDFFX1 DFF_212_Q_reg ( .D(n301), .SI(n8683), .SE(n10155), .CLK(n10348), .Q(
        n8682) );
  SDFFX1 DFF_213_Q_reg ( .D(n302), .SI(n8682), .SE(n10155), .CLK(n10348), .Q(
        n8681) );
  SDFFX1 DFF_214_Q_reg ( .D(n303), .SI(n8681), .SE(n10155), .CLK(n10348), .Q(
        n8680) );
  SDFFX1 DFF_215_Q_reg ( .D(n304), .SI(n8680), .SE(n10155), .CLK(n10348), .Q(
        test_so12) );
  SDFFX1 DFF_216_Q_reg ( .D(n305), .SI(test_si13), .SE(n10155), .CLK(n10348), 
        .Q(n8677) );
  SDFFX1 DFF_217_Q_reg ( .D(n306), .SI(n8677), .SE(n10027), .CLK(n10347), .Q(
        n8676) );
  SDFFX1 DFF_218_Q_reg ( .D(n307), .SI(n8676), .SE(test_se), .CLK(n10347), .Q(
        n8675) );
  SDFFX1 DFF_219_Q_reg ( .D(n308), .SI(n8675), .SE(n10028), .CLK(n10347), .Q(
        n8674) );
  SDFFX1 DFF_220_Q_reg ( .D(n309), .SI(n8674), .SE(n10024), .CLK(n10347), .Q(
        n8673) );
  SDFFX1 DFF_221_Q_reg ( .D(n310), .SI(n8673), .SE(n10025), .CLK(n10347), .Q(
        n8672) );
  SDFFX1 DFF_222_Q_reg ( .D(n311), .SI(n8672), .SE(n10022), .CLK(n10347), .Q(
        n8671) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n10023), .CLK(n10347), 
        .Q(n8670) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n10153), .CLK(n10350), 
        .Q(n8669), .QN(n18352) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n10153), .CLK(n10350), 
        .Q(n8668), .QN(n18353) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n10153), .CLK(n10350), 
        .Q(n8667), .QN(n18354) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n10153), .CLK(n10350), 
        .Q(n8666), .QN(n18355) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n10152), .CLK(n10351), 
        .Q(n8665), .QN(n18356) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n10152), .CLK(n10351), 
        .Q(n8664), .QN(n18357) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n10152), .CLK(n10351), 
        .Q(n8663), .QN(n18358) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n10151), .CLK(n10352), 
        .Q(n8662), .QN(n18359) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n10151), .CLK(n10352), 
        .Q(n8661), .QN(n18360) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n10030), .CLK(n10475), 
        .Q(test_so13), .QN(n9845) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n10150), .CLK(n10353), 
        .Q(n8658), .QN(n18361) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n10150), .CLK(n10353), 
        .Q(n8657), .QN(n18362) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n10150), .CLK(n10353), 
        .Q(n8656), .QN(n18363) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n10150), .CLK(n10353), 
        .Q(n8655), .QN(n18364) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n10149), .CLK(n10354), 
        .Q(n8654), .QN(n18365) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n10149), .CLK(n10354), 
        .Q(n8653), .QN(n18366) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n10149), .CLK(n10354), 
        .Q(WX1970), .QN(n9485) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n10148), .CLK(n10355), 
        .Q(WX1972), .QN(n9484) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n10148), .CLK(n10355), 
        .Q(WX1974), .QN(n9482) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n10148), .CLK(n10355), 
        .Q(WX1976), .QN(n9480) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n10147), .CLK(n10356), 
        .Q(WX1978), .QN(n9478) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n10147), .CLK(n10356), 
        .Q(WX1980), .QN(n9476) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n10147), .CLK(n10356), 
        .Q(WX1982), .QN(n9474) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n10146), .CLK(n10357), 
        .Q(WX1984), .QN(n9472) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n10146), .CLK(n10357), 
        .Q(WX1986), .QN(n9470) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n10146), .CLK(n10357), 
        .Q(WX1988), .QN(n9468) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n10025), .CLK(n10358), 
        .Q(WX1990), .QN(n9466) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n10027), .CLK(n10358), 
        .Q(test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n10145), .CLK(n10359), 
        .Q(WX1994), .QN(n9463) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n10145), .CLK(n10359), 
        .Q(WX1996), .QN(n9461) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n10145), .CLK(n10359), 
        .Q(WX1998), .QN(n9459) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n10145), .CLK(n10359), 
        .Q(WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n10153), .CLK(n10350), 
        .Q(WX2002), .QN(n9017) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n10153), .CLK(n10350), 
        .Q(WX2004), .QN(n9243) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n10153), .CLK(n10350), 
        .Q(WX2006), .QN(n9241) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n10153), .CLK(n10350), 
        .Q(WX2008), .QN(n9239) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n10152), .CLK(n10351), 
        .Q(WX2010), .QN(n9237) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n10152), .CLK(n10351), 
        .Q(WX2012), .QN(n9235) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n10152), .CLK(n10351), 
        .Q(WX2014), .QN(n9233) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n10151), .CLK(n10352), 
        .Q(WX2016), .QN(n9231) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n10151), .CLK(n10352), 
        .Q(WX2018), .QN(n9229) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n10151), .CLK(n10352), 
        .Q(WX2020), .QN(n9227) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n10151), .CLK(n10352), 
        .Q(WX2022), .QN(n9225) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n10150), .CLK(n10353), 
        .Q(WX2024), .QN(n9223) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n10150), .CLK(n10353), 
        .Q(WX2026), .QN(n9221) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n10149), .CLK(n10354), 
        .Q(test_so15), .QN(n9870) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n10149), .CLK(n10354), 
        .Q(WX2030), .QN(n9218) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n10149), .CLK(n10354), 
        .Q(WX2032), .QN(n9216) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n10148), .CLK(n10355), 
        .Q(WX2034) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n10148), .CLK(n10355), 
        .Q(WX2036) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n10148), .CLK(n10355), 
        .Q(WX2038) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n10147), .CLK(n10356), 
        .Q(WX2040) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n10147), .CLK(n10356), 
        .Q(WX2042) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n10147), .CLK(n10356), 
        .Q(WX2044) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n10146), .CLK(n10357), 
        .Q(WX2046) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n10146), .CLK(n10357), 
        .Q(WX2048) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n10146), .CLK(n10357), 
        .Q(WX2050) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n10026), .CLK(n10358), 
        .Q(WX2052) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n10024), .CLK(n10358), 
        .Q(WX2054) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n10026), .CLK(n10358), 
        .Q(WX2056) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n10025), .CLK(n10358), 
        .Q(WX2058) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n10145), .CLK(n10359), 
        .Q(WX2060) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n10145), .CLK(n10359), 
        .Q(WX2062) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n10144), .CLK(n10360), 
        .Q(test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n10153), .CLK(n10350), 
        .Q(WX2066), .QN(n9018) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n10153), .CLK(n10350), 
        .Q(WX2068), .QN(n9244) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n10153), .CLK(n10350), 
        .Q(WX2070), .QN(n9242) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n10153), .CLK(n10350), 
        .Q(WX2072), .QN(n9240) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n10152), .CLK(n10351), 
        .Q(WX2074), .QN(n9238) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n10152), .CLK(n10351), 
        .Q(WX2076), .QN(n9236) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n10152), .CLK(n10351), 
        .Q(WX2078), .QN(n9234) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n10151), .CLK(n10352), 
        .Q(WX2080), .QN(n9232) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n10151), .CLK(n10352), 
        .Q(WX2082), .QN(n9230) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n10151), .CLK(n10352), 
        .Q(WX2084), .QN(n9228) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n10150), .CLK(n10353), 
        .Q(WX2086), .QN(n9226) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n10150), .CLK(n10353), 
        .Q(WX2088), .QN(n9224) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n10150), .CLK(n10353), 
        .Q(WX2090), .QN(n9222) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n10149), .CLK(n10354), 
        .Q(WX2092), .QN(n9220) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n10149), .CLK(n10354), 
        .Q(WX2094), .QN(n9219) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n10149), .CLK(n10354), 
        .Q(WX2096), .QN(n9217) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n10148), .CLK(n10355), 
        .Q(WX2098), .QN(n9486) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n10148), .CLK(n10355), 
        .Q(test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n10148), .CLK(n10355), 
        .Q(WX2102), .QN(n9483) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n10147), .CLK(n10356), 
        .Q(WX2104), .QN(n9481) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n10147), .CLK(n10356), 
        .Q(WX2106), .QN(n9479) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n10147), .CLK(n10356), 
        .Q(WX2108), .QN(n9477) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n10146), .CLK(n10357), 
        .Q(WX2110), .QN(n9475) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n10146), .CLK(n10357), 
        .Q(WX2112), .QN(n9473) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n10146), .CLK(n10357), 
        .Q(WX2114), .QN(n9471) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n10023), .CLK(n10358), 
        .Q(WX2116), .QN(n9469) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n10028), .CLK(n10358), 
        .Q(WX2118), .QN(n9467) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n10023), .CLK(n10358), 
        .Q(WX2120), .QN(n9465) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n10145), .CLK(n10359), 
        .Q(WX2122), .QN(n9464) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n10145), .CLK(n10359), 
        .Q(WX2124), .QN(n9462) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n10145), .CLK(n10359), 
        .Q(WX2126), .QN(n9460) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n10144), .CLK(n10360), 
        .Q(WX2128), .QN(n9458) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n10144), .CLK(n10360), 
        .Q(WX2130) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n10144), .CLK(n10360), 
        .Q(WX2132) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n10144), .CLK(n10360), 
        .Q(WX2134) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n10144), .CLK(n10360), 
        .Q(test_so18), .QN(n9832) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n10152), .CLK(n10351), 
        .Q(WX2138) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n10152), .CLK(n10351), 
        .Q(WX2140), .QN(n9715) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n10152), .CLK(n10351), 
        .Q(WX2142) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n10151), .CLK(n10352), 
        .Q(WX2144) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n10151), .CLK(n10352), 
        .Q(WX2146) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n10151), .CLK(n10352), 
        .Q(WX2148), .QN(n9719) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n10150), .CLK(n10353), 
        .Q(WX2150) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n10150), .CLK(n10353), 
        .Q(WX2152) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n10150), .CLK(n10353), 
        .Q(WX2154) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n10149), .CLK(n10354), 
        .Q(WX2156), .QN(n9723) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n10149), .CLK(n10354), 
        .Q(WX2158) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n10149), .CLK(n10354), 
        .Q(WX2160), .QN(n9514) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n10148), .CLK(n10355), 
        .Q(WX2162) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n10148), .CLK(n10355), 
        .Q(WX2164) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n10148), .CLK(n10355), 
        .Q(WX2166) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n10147), .CLK(n10356), 
        .Q(WX2168) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n10147), .CLK(n10356), 
        .Q(WX2170), .QN(n9515) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n10147), .CLK(n10356), 
        .Q(test_so19), .QN(n9836) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n10146), .CLK(n10357), 
        .Q(WX2174) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n10146), .CLK(n10357), 
        .Q(WX2176), .QN(n9730) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n10146), .CLK(n10357), 
        .Q(WX2178) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n10022), .CLK(n10358), 
        .Q(WX2180) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(test_se), .CLK(n10358), 
        .Q(WX2182) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n10022), .CLK(n10358), 
        .Q(WX2184), .QN(n9516) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n10145), .CLK(n10359), 
        .Q(WX2186) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n10145), .CLK(n10359), 
        .Q(WX2188) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n10145), .CLK(n10359), 
        .Q(WX2190) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n10144), .CLK(n10360), 
        .Q(WX2192), .QN(n9524) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n10033), .CLK(n10472), 
        .Q(CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_8_3), .QN(DFF_355_n1) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n10032), .CLK(
        n10473), .Q(test_so20), .QN(n9861) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n10032), .CLK(n10473), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_10), .QN(DFF_362_n1) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n10032), .CLK(
        n10473), .Q(CRC_OUT_8_15), .QN(DFF_367_n1) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n10031), .CLK(
        n10474), .Q(test_so21), .QN(n9862) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n10031), .CLK(n10474), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n10031), .CLK(
        n10474), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n10030), .CLK(
        n10475), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n10030), .CLK(
        n10475), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n10030), .CLK(
        n10475), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n10144), .CLK(
        n10360), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n568), .SI(CRC_OUT_8_31), .SE(n10144), .CLK(n10360), .Q(WX3071), .QN(n9494) );
  SDFFX1 DFF_385_Q_reg ( .D(n569), .SI(WX3071), .SE(n10141), .CLK(n10363), .Q(
        n8644) );
  SDFFX1 DFF_386_Q_reg ( .D(n570), .SI(n8644), .SE(n10141), .CLK(n10363), .Q(
        n8643) );
  SDFFX1 DFF_387_Q_reg ( .D(n571), .SI(n8643), .SE(n10141), .CLK(n10363), .Q(
        n8642) );
  SDFFX1 DFF_388_Q_reg ( .D(n572), .SI(n8642), .SE(n10141), .CLK(n10363), .Q(
        n8641) );
  SDFFX1 DFF_389_Q_reg ( .D(n573), .SI(n8641), .SE(n10142), .CLK(n10362), .Q(
        n8640) );
  SDFFX1 DFF_390_Q_reg ( .D(n574), .SI(n8640), .SE(n10142), .CLK(n10362), .Q(
        n8639) );
  SDFFX1 DFF_391_Q_reg ( .D(n575), .SI(n8639), .SE(n10142), .CLK(n10362), .Q(
        n8638) );
  SDFFX1 DFF_392_Q_reg ( .D(n576), .SI(n8638), .SE(n10142), .CLK(n10362), .Q(
        n8637) );
  SDFFX1 DFF_393_Q_reg ( .D(n577), .SI(n8637), .SE(n10142), .CLK(n10362), .Q(
        n8636) );
  SDFFX1 DFF_394_Q_reg ( .D(n578), .SI(n8636), .SE(n10142), .CLK(n10362), .Q(
        n8635) );
  SDFFX1 DFF_395_Q_reg ( .D(n579), .SI(n8635), .SE(n10142), .CLK(n10362), .Q(
        test_so22) );
  SDFFX1 DFF_396_Q_reg ( .D(n580), .SI(test_si23), .SE(n10142), .CLK(n10362), 
        .Q(n8632) );
  SDFFX1 DFF_397_Q_reg ( .D(n581), .SI(n8632), .SE(n10142), .CLK(n10362), .Q(
        n8631) );
  SDFFX1 DFF_398_Q_reg ( .D(n582), .SI(n8631), .SE(n10142), .CLK(n10362), .Q(
        n8630) );
  SDFFX1 DFF_399_Q_reg ( .D(n583), .SI(n8630), .SE(n10142), .CLK(n10362), .Q(
        n8629) );
  SDFFX1 DFF_400_Q_reg ( .D(n584), .SI(n8629), .SE(n10142), .CLK(n10362), .Q(
        n8628) );
  SDFFX1 DFF_401_Q_reg ( .D(n585), .SI(n8628), .SE(n10143), .CLK(n10361), .Q(
        n8627) );
  SDFFX1 DFF_402_Q_reg ( .D(n586), .SI(n8627), .SE(n10143), .CLK(n10361), .Q(
        n8626) );
  SDFFX1 DFF_403_Q_reg ( .D(n587), .SI(n8626), .SE(n10143), .CLK(n10361), .Q(
        n8625) );
  SDFFX1 DFF_404_Q_reg ( .D(n588), .SI(n8625), .SE(n10143), .CLK(n10361), .Q(
        n8624) );
  SDFFX1 DFF_405_Q_reg ( .D(n589), .SI(n8624), .SE(n10143), .CLK(n10361), .Q(
        n8623) );
  SDFFX1 DFF_406_Q_reg ( .D(n590), .SI(n8623), .SE(n10143), .CLK(n10361), .Q(
        n8622) );
  SDFFX1 DFF_407_Q_reg ( .D(n591), .SI(n8622), .SE(n10143), .CLK(n10361), .Q(
        n8621) );
  SDFFX1 DFF_408_Q_reg ( .D(n592), .SI(n8621), .SE(n10143), .CLK(n10361), .Q(
        n8620) );
  SDFFX1 DFF_409_Q_reg ( .D(n593), .SI(n8620), .SE(n10143), .CLK(n10361), .Q(
        n8619) );
  SDFFX1 DFF_410_Q_reg ( .D(n594), .SI(n8619), .SE(n10143), .CLK(n10361), .Q(
        n8618) );
  SDFFX1 DFF_411_Q_reg ( .D(n595), .SI(n8618), .SE(n10143), .CLK(n10361), .Q(
        n8617) );
  SDFFX1 DFF_412_Q_reg ( .D(n596), .SI(n8617), .SE(n10143), .CLK(n10361), .Q(
        n8616) );
  SDFFX1 DFF_413_Q_reg ( .D(n597), .SI(n8616), .SE(n10144), .CLK(n10360), .Q(
        test_so23) );
  SDFFX1 DFF_414_Q_reg ( .D(n598), .SI(test_si24), .SE(n10144), .CLK(n10360), 
        .Q(n8613) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n10144), .CLK(n10360), 
        .Q(n8612) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n10141), .CLK(n10363), 
        .Q(n8611), .QN(n18367) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n10141), .CLK(n10363), 
        .Q(n8610), .QN(n18368) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n10141), .CLK(n10363), 
        .Q(n8609), .QN(n18369) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n10141), .CLK(n10363), 
        .Q(n8608), .QN(n18370) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n10140), .CLK(n10364), 
        .Q(n8607), .QN(n18371) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n10140), .CLK(n10364), 
        .Q(n8606), .QN(n18372) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n10140), .CLK(n10364), 
        .Q(n8605), .QN(n18373) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n10140), .CLK(n10364), 
        .Q(n8604), .QN(n18374) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n10140), .CLK(n10364), 
        .Q(n8603), .QN(n18375) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n10139), .CLK(n10365), 
        .Q(n8602), .QN(n18376) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n10139), .CLK(n10365), 
        .Q(n8601), .QN(n18377) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n10138), .CLK(n10366), 
        .Q(n8600), .QN(n18378) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n10138), .CLK(n10366), 
        .Q(n8599), .QN(n18379) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n10138), .CLK(n10366), 
        .Q(n8598), .QN(n18380) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n10138), .CLK(n10366), 
        .Q(n8597), .QN(n18381) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n10033), .CLK(n10472), 
        .Q(test_so24), .QN(n9844) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n10025), .CLK(n10367), 
        .Q(WX3263), .QN(n9455) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n10024), .CLK(n10367), 
        .Q(WX3265), .QN(n9453) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n10137), .CLK(n10368), 
        .Q(WX3267), .QN(n9451) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n10137), .CLK(n10368), 
        .Q(WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n10137), .CLK(n10368), 
        .Q(WX3271), .QN(n9447) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n10136), .CLK(n10369), 
        .Q(WX3273), .QN(n9445) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n10136), .CLK(n10369), 
        .Q(WX3275), .QN(n9443) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n10136), .CLK(n10369), 
        .Q(WX3277), .QN(n9442) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n10135), .CLK(n10370), 
        .Q(WX3279), .QN(n9440) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n10135), .CLK(n10370), 
        .Q(WX3281), .QN(n9438) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n10135), .CLK(n10370), 
        .Q(WX3283), .QN(n9436) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n10134), .CLK(n10371), 
        .Q(WX3285), .QN(n9434) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n10134), .CLK(n10371), 
        .Q(WX3287), .QN(n9432) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n10134), .CLK(n10371), 
        .Q(WX3289), .QN(n9430) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n10133), .CLK(n10372), 
        .Q(WX3291), .QN(n9428) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n10133), .CLK(n10372), 
        .Q(WX3293), .QN(n9426) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n10141), .CLK(n10363), 
        .Q(WX3295), .QN(n9015) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n10141), .CLK(n10363), 
        .Q(test_so25) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n10141), .CLK(n10363), 
        .Q(WX3299), .QN(n9213) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n10141), .CLK(n10363), 
        .Q(WX3301), .QN(n9211) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n10140), .CLK(n10364), 
        .Q(WX3303), .QN(n9209) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n10140), .CLK(n10364), 
        .Q(WX3305), .QN(n9208) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n10140), .CLK(n10364), 
        .Q(WX3307), .QN(n9206) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n10140), .CLK(n10364), 
        .Q(WX3309), .QN(n9204) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n10140), .CLK(n10364), 
        .Q(WX3311), .QN(n9202) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n10139), .CLK(n10365), 
        .Q(WX3313), .QN(n9200) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n10139), .CLK(n10365), 
        .Q(WX3315), .QN(n9198) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n10139), .CLK(n10365), 
        .Q(WX3317), .QN(n9196) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n10138), .CLK(n10366), 
        .Q(WX3319), .QN(n9194) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n10138), .CLK(n10366), 
        .Q(WX3321), .QN(n9192) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n10138), .CLK(n10366), 
        .Q(WX3323), .QN(n9190) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n10028), .CLK(n10367), 
        .Q(WX3325), .QN(n9188) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n10026), .CLK(n10367), 
        .Q(WX3327), .QN(n3753) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n10028), .CLK(n10367), 
        .Q(WX3329), .QN(n3751) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n10137), .CLK(n10368), 
        .Q(WX3331), .QN(n3749) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n10137), .CLK(n10368), 
        .Q(test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n10137), .CLK(n10368), 
        .Q(WX3335), .QN(n3745) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n10136), .CLK(n10369), 
        .Q(WX3337), .QN(n3743) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n10136), .CLK(n10369), 
        .Q(WX3339), .QN(n3741) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n10136), .CLK(n10369), 
        .Q(WX3341) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n10135), .CLK(n10370), 
        .Q(WX3343), .QN(n3737) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n10135), .CLK(n10370), 
        .Q(WX3345) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n10135), .CLK(n10370), 
        .Q(WX3347), .QN(n3733) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n10134), .CLK(n10371), 
        .Q(WX3349), .QN(n3731) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n10134), .CLK(n10371), 
        .Q(WX3351), .QN(n3729) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n10134), .CLK(n10371), 
        .Q(WX3353), .QN(n3727) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n10133), .CLK(n10372), 
        .Q(WX3355), .QN(n3725) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n10133), .CLK(n10372), 
        .Q(WX3357), .QN(n3723) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n10133), .CLK(n10372), 
        .Q(WX3359), .QN(n9016) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n10133), .CLK(n10372), 
        .Q(WX3361), .QN(n9215) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n10132), .CLK(n10373), 
        .Q(WX3363), .QN(n9214) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n10132), .CLK(n10373), 
        .Q(WX3365), .QN(n9212) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n10132), .CLK(n10373), 
        .Q(WX3367), .QN(n9210) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n10132), .CLK(n10373), 
        .Q(test_so27) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n10140), .CLK(n10364), 
        .Q(WX3371), .QN(n9207) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n10140), .CLK(n10364), 
        .Q(WX3373), .QN(n9205) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n10139), .CLK(n10365), 
        .Q(WX3375), .QN(n9203) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n10139), .CLK(n10365), 
        .Q(WX3377), .QN(n9201) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n10139), .CLK(n10365), 
        .Q(WX3379), .QN(n9199) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n10139), .CLK(n10365), 
        .Q(WX3381), .QN(n9197) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n10138), .CLK(n10366), 
        .Q(WX3383), .QN(n9195) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n10138), .CLK(n10366), 
        .Q(WX3385), .QN(n9193) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n10138), .CLK(n10366), 
        .Q(WX3387), .QN(n9191) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(test_se), .CLK(n10367), 
        .Q(WX3389), .QN(n9189) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n10023), .CLK(n10367), 
        .Q(WX3391), .QN(n9456) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(test_se), .CLK(n10367), 
        .Q(WX3393), .QN(n9454) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n10137), .CLK(n10368), 
        .Q(WX3395), .QN(n9452) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n10137), .CLK(n10368), 
        .Q(WX3397), .QN(n9450) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n10137), .CLK(n10368), 
        .Q(WX3399), .QN(n9448) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n10136), .CLK(n10369), 
        .Q(WX3401), .QN(n9446) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n10136), .CLK(n10369), 
        .Q(WX3403), .QN(n9444) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n10136), .CLK(n10369), 
        .Q(test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n10135), .CLK(n10370), 
        .Q(WX3407), .QN(n9441) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n10135), .CLK(n10370), 
        .Q(WX3409), .QN(n9439) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n10135), .CLK(n10370), 
        .Q(WX3411), .QN(n9437) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n10134), .CLK(n10371), 
        .Q(WX3413), .QN(n9435) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n10134), .CLK(n10371), 
        .Q(WX3415), .QN(n9433) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n10134), .CLK(n10371), 
        .Q(WX3417), .QN(n9431) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n10133), .CLK(n10372), 
        .Q(WX3419), .QN(n9429) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n10133), .CLK(n10372), 
        .Q(WX3421), .QN(n9427) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n10133), .CLK(n10372), 
        .Q(WX3423) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n10133), .CLK(n10372), 
        .Q(WX3425), .QN(n9686) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n10132), .CLK(n10373), 
        .Q(WX3427) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n10132), .CLK(n10373), 
        .Q(WX3429), .QN(n9688) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n10132), .CLK(n10373), 
        .Q(WX3431) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n10132), .CLK(n10373), 
        .Q(WX3433), .QN(n9690) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n10132), .CLK(n10373), 
        .Q(WX3435) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n10132), .CLK(n10373), 
        .Q(WX3437) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n10132), .CLK(n10373), 
        .Q(test_so29), .QN(n9831) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n10139), .CLK(n10365), 
        .Q(WX3441) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n10139), .CLK(n10365), 
        .Q(WX3443) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n10139), .CLK(n10365), 
        .Q(WX3445) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n10138), .CLK(n10366), 
        .Q(WX3447) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n10138), .CLK(n10366), 
        .Q(WX3449) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n10024), .CLK(n10367), 
        .Q(WX3451) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n10027), .CLK(n10367), 
        .Q(WX3453), .QN(n9511) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n10022), .CLK(n10367), 
        .Q(WX3455), .QN(n9699) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n10027), .CLK(n10367), 
        .Q(WX3457), .QN(n9700) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n10137), .CLK(n10368), 
        .Q(WX3459), .QN(n9701) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n10137), .CLK(n10368), 
        .Q(WX3461) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n10137), .CLK(n10368), 
        .Q(WX3463), .QN(n9512) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n10136), .CLK(n10369), 
        .Q(WX3465), .QN(n9703) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n10136), .CLK(n10369), 
        .Q(WX3467), .QN(n9704) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n10136), .CLK(n10369), 
        .Q(WX3469) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n10135), .CLK(n10370), 
        .Q(WX3471), .QN(n9706) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n10135), .CLK(n10370), 
        .Q(test_so30), .QN(n9835) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n10135), .CLK(n10370), 
        .Q(WX3475), .QN(n9707) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n10134), .CLK(n10371), 
        .Q(WX3477), .QN(n9513) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n10134), .CLK(n10371), 
        .Q(WX3479), .QN(n9708) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n10134), .CLK(n10371), 
        .Q(WX3481), .QN(n9709) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n10133), .CLK(n10372), 
        .Q(WX3483), .QN(n9710) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n10133), .CLK(n10372), 
        .Q(WX3485), .QN(n9523) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n10035), .CLK(n10470), 
        .Q(CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_7_3), .QN(DFF_547_n1) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n10034), .CLK(
        n10471), .Q(test_so31), .QN(n9871) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n10034), .CLK(n10471), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_15), .QN(DFF_559_n1) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n10034), .CLK(
        n10471), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n10033), .CLK(
        n10472), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n10132), .CLK(
        n10373), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n10131), .CLK(
        n10374), .Q(test_so32), .QN(n9860) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n10131), .CLK(n10374), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n10131), .CLK(
        n10374), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n10131), .CLK(
        n10374), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n10131), .CLK(
        n10374), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n809), .SI(CRC_OUT_7_31), .SE(n10131), .CLK(n10374), .Q(WX4364), .QN(n9493) );
  SDFFX1 DFF_577_Q_reg ( .D(n810), .SI(WX4364), .SE(n10128), .CLK(n10377), .Q(
        n8586) );
  SDFFX1 DFF_578_Q_reg ( .D(n811), .SI(n8586), .SE(n10129), .CLK(n10376), .Q(
        n8585) );
  SDFFX1 DFF_579_Q_reg ( .D(n812), .SI(n8585), .SE(n10129), .CLK(n10376), .Q(
        n8584) );
  SDFFX1 DFF_580_Q_reg ( .D(n813), .SI(n8584), .SE(n10129), .CLK(n10376), .Q(
        n8583) );
  SDFFX1 DFF_581_Q_reg ( .D(n814), .SI(n8583), .SE(n10129), .CLK(n10376), .Q(
        n8582) );
  SDFFX1 DFF_582_Q_reg ( .D(n815), .SI(n8582), .SE(n10129), .CLK(n10376), .Q(
        n8581) );
  SDFFX1 DFF_583_Q_reg ( .D(n816), .SI(n8581), .SE(n10129), .CLK(n10376), .Q(
        n8580) );
  SDFFX1 DFF_584_Q_reg ( .D(n817), .SI(n8580), .SE(n10129), .CLK(n10376), .Q(
        n8579) );
  SDFFX1 DFF_585_Q_reg ( .D(n818), .SI(n8579), .SE(n10129), .CLK(n10376), .Q(
        n8578) );
  SDFFX1 DFF_586_Q_reg ( .D(n819), .SI(n8578), .SE(n10129), .CLK(n10376), .Q(
        n8577) );
  SDFFX1 DFF_587_Q_reg ( .D(n820), .SI(n8577), .SE(n10129), .CLK(n10376), .Q(
        n8576) );
  SDFFX1 DFF_588_Q_reg ( .D(n821), .SI(n8576), .SE(n10129), .CLK(n10376), .Q(
        test_so33) );
  SDFFX1 DFF_589_Q_reg ( .D(n822), .SI(test_si34), .SE(n10129), .CLK(n10376), 
        .Q(n8573) );
  SDFFX1 DFF_590_Q_reg ( .D(n823), .SI(n8573), .SE(n10130), .CLK(n10375), .Q(
        n8572) );
  SDFFX1 DFF_591_Q_reg ( .D(n824), .SI(n8572), .SE(n10130), .CLK(n10375), .Q(
        n8571) );
  SDFFX1 DFF_592_Q_reg ( .D(n825), .SI(n8571), .SE(n10130), .CLK(n10375), .Q(
        n8570) );
  SDFFX1 DFF_593_Q_reg ( .D(n826), .SI(n8570), .SE(n10130), .CLK(n10375), .Q(
        n8569) );
  SDFFX1 DFF_594_Q_reg ( .D(n827), .SI(n8569), .SE(n10130), .CLK(n10375), .Q(
        n8568) );
  SDFFX1 DFF_595_Q_reg ( .D(n828), .SI(n8568), .SE(n10130), .CLK(n10375), .Q(
        n8567) );
  SDFFX1 DFF_596_Q_reg ( .D(n829), .SI(n8567), .SE(n10130), .CLK(n10375), .Q(
        n8566) );
  SDFFX1 DFF_597_Q_reg ( .D(n830), .SI(n8566), .SE(n10130), .CLK(n10375), .Q(
        n8565) );
  SDFFX1 DFF_598_Q_reg ( .D(n831), .SI(n8565), .SE(n10130), .CLK(n10375), .Q(
        n8564) );
  SDFFX1 DFF_599_Q_reg ( .D(n832), .SI(n8564), .SE(n10130), .CLK(n10375), .Q(
        n8563) );
  SDFFX1 DFF_600_Q_reg ( .D(n833), .SI(n8563), .SE(n10130), .CLK(n10375), .Q(
        n8562) );
  SDFFX1 DFF_601_Q_reg ( .D(n834), .SI(n8562), .SE(n10130), .CLK(n10375), .Q(
        n8561) );
  SDFFX1 DFF_602_Q_reg ( .D(n835), .SI(n8561), .SE(n10131), .CLK(n10374), .Q(
        n8560) );
  SDFFX1 DFF_603_Q_reg ( .D(n836), .SI(n8560), .SE(n10131), .CLK(n10374), .Q(
        n8559) );
  SDFFX1 DFF_604_Q_reg ( .D(n837), .SI(n8559), .SE(n10131), .CLK(n10374), .Q(
        n8558) );
  SDFFX1 DFF_605_Q_reg ( .D(n838), .SI(n8558), .SE(n10131), .CLK(n10374), .Q(
        test_so34) );
  SDFFX1 DFF_606_Q_reg ( .D(n839), .SI(test_si35), .SE(n10131), .CLK(n10374), 
        .Q(n8555) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n10131), .CLK(n10374), 
        .Q(n8554) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n10128), .CLK(n10377), 
        .Q(n8553), .QN(n18382) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n10128), .CLK(n10377), 
        .Q(n8552), .QN(n18383) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n10128), .CLK(n10377), 
        .Q(n8551), .QN(n18384) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n10128), .CLK(n10377), 
        .Q(n8550), .QN(n18385) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n10128), .CLK(n10377), 
        .Q(n8549), .QN(n18386) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n10127), .CLK(n10378), 
        .Q(n8548), .QN(n18387) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n10127), .CLK(n10378), 
        .Q(n8547), .QN(n18388) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n10126), .CLK(n10379), 
        .Q(n8546), .QN(n18389) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n10126), .CLK(n10379), 
        .Q(n8545), .QN(n18390) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n10126), .CLK(n10379), 
        .Q(n8544), .QN(n18391) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n10126), .CLK(n10379), 
        .Q(n8543), .QN(n18392) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n10125), .CLK(n10380), 
        .Q(n8542), .QN(n18393) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n10125), .CLK(n10380), 
        .Q(n8541), .QN(n18394) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n10124), .CLK(n10381), 
        .Q(n8540), .QN(n18395) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n10124), .CLK(n10381), 
        .Q(test_so35), .QN(n9843) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n10124), .CLK(n10381), 
        .Q(n8537), .QN(n18396) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n10124), .CLK(n10381), 
        .Q(WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n10123), .CLK(n10382), 
        .Q(WX4558), .QN(n9422) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n10123), .CLK(n10382), 
        .Q(WX4560), .QN(n9421) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n10123), .CLK(n10382), 
        .Q(WX4562), .QN(n9419) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n10122), .CLK(n10383), 
        .Q(WX4564), .QN(n9417) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n10122), .CLK(n10383), 
        .Q(WX4566), .QN(n9415) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n10122), .CLK(n10383), 
        .Q(WX4568), .QN(n9413) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n10121), .CLK(n10384), 
        .Q(WX4570), .QN(n9411) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n10121), .CLK(n10384), 
        .Q(WX4572), .QN(n9409) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n10121), .CLK(n10384), 
        .Q(WX4574), .QN(n9407) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n10120), .CLK(n10385), 
        .Q(WX4576), .QN(n9405) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n10120), .CLK(n10385), 
        .Q(WX4578), .QN(n9403) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n10120), .CLK(n10385), 
        .Q(WX4580), .QN(n9401) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n10119), .CLK(n10386), 
        .Q(WX4582), .QN(n9399) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n10119), .CLK(n10386), 
        .Q(WX4584), .QN(n9397) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n10119), .CLK(n10386), 
        .Q(test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n10128), .CLK(n10377), 
        .Q(WX4588), .QN(n9013) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n10128), .CLK(n10377), 
        .Q(WX4590), .QN(n9187) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n10128), .CLK(n10377), 
        .Q(WX4592), .QN(n9185) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n10128), .CLK(n10377), 
        .Q(WX4594), .QN(n9183) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n10127), .CLK(n10378), 
        .Q(WX4596), .QN(n9181) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n10127), .CLK(n10378), 
        .Q(WX4598), .QN(n9179) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n10127), .CLK(n10378), 
        .Q(WX4600), .QN(n9177) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n10127), .CLK(n10378), 
        .Q(WX4602), .QN(n9175) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n10126), .CLK(n10379), 
        .Q(WX4604), .QN(n9173) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n10126), .CLK(n10379), 
        .Q(WX4606), .QN(n9171) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n10125), .CLK(n10380), 
        .Q(WX4608), .QN(n9169) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n10125), .CLK(n10380), 
        .Q(WX4610), .QN(n9167) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n10125), .CLK(n10380), 
        .Q(WX4612), .QN(n9165) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n10125), .CLK(n10380), 
        .Q(WX4614), .QN(n9163) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n10124), .CLK(n10381), 
        .Q(WX4616), .QN(n9161) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n10124), .CLK(n10381), 
        .Q(WX4618), .QN(n9159) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n10123), .CLK(n10382), 
        .Q(test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n10123), .CLK(n10382), 
        .Q(WX4622), .QN(n3719) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n10123), .CLK(n10382), 
        .Q(WX4624) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n10122), .CLK(n10383), 
        .Q(WX4626), .QN(n3715) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n10122), .CLK(n10383), 
        .Q(WX4628) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n10122), .CLK(n10383), 
        .Q(WX4630), .QN(n3711) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n10121), .CLK(n10384), 
        .Q(WX4632), .QN(n3709) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n10121), .CLK(n10384), 
        .Q(WX4634), .QN(n3707) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n10121), .CLK(n10384), 
        .Q(WX4636), .QN(n3705) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n10120), .CLK(n10385), 
        .Q(WX4638), .QN(n3703) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n10120), .CLK(n10385), 
        .Q(WX4640), .QN(n3701) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n10120), .CLK(n10385), 
        .Q(WX4642), .QN(n3699) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n10119), .CLK(n10386), 
        .Q(WX4644), .QN(n3697) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n10119), .CLK(n10386), 
        .Q(WX4646), .QN(n3695) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n10119), .CLK(n10386), 
        .Q(WX4648), .QN(n3693) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n10118), .CLK(n10387), 
        .Q(WX4650) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n10118), .CLK(n10387), 
        .Q(WX4652), .QN(n9014) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n10118), .CLK(n10387), 
        .Q(test_so38) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n10128), .CLK(n10377), 
        .Q(WX4656), .QN(n9186) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n10128), .CLK(n10377), 
        .Q(WX4658), .QN(n9184) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n10127), .CLK(n10378), 
        .Q(WX4660), .QN(n9182) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n10127), .CLK(n10378), 
        .Q(WX4662), .QN(n9180) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n10127), .CLK(n10378), 
        .Q(WX4664), .QN(n9178) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n10126), .CLK(n10379), 
        .Q(WX4666), .QN(n9176) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n10126), .CLK(n10379), 
        .Q(WX4668), .QN(n9174) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n10126), .CLK(n10379), 
        .Q(WX4670), .QN(n9172) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n10125), .CLK(n10380), 
        .Q(WX4672), .QN(n9170) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n10125), .CLK(n10380), 
        .Q(WX4674), .QN(n9168) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n10125), .CLK(n10380), 
        .Q(WX4676), .QN(n9166) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n10124), .CLK(n10381), 
        .Q(WX4678), .QN(n9164) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n10124), .CLK(n10381), 
        .Q(WX4680), .QN(n9162) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n10124), .CLK(n10381), 
        .Q(WX4682), .QN(n9160) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n10123), .CLK(n10382), 
        .Q(WX4684), .QN(n9425) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n10123), .CLK(n10382), 
        .Q(WX4686), .QN(n9423) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n10123), .CLK(n10382), 
        .Q(test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n10122), .CLK(n10383), 
        .Q(WX4690), .QN(n9420) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n10122), .CLK(n10383), 
        .Q(WX4692), .QN(n9418) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n10122), .CLK(n10383), 
        .Q(WX4694), .QN(n9416) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n10121), .CLK(n10384), 
        .Q(WX4696), .QN(n9414) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n10121), .CLK(n10384), 
        .Q(WX4698), .QN(n9412) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n10121), .CLK(n10384), 
        .Q(WX4700), .QN(n9410) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n10120), .CLK(n10385), 
        .Q(WX4702), .QN(n9408) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n10120), .CLK(n10385), 
        .Q(WX4704), .QN(n9406) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n10120), .CLK(n10385), 
        .Q(WX4706), .QN(n9404) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n10119), .CLK(n10386), 
        .Q(WX4708), .QN(n9402) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n10119), .CLK(n10386), 
        .Q(WX4710), .QN(n9400) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n10119), .CLK(n10386), 
        .Q(WX4712), .QN(n9398) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n10118), .CLK(n10387), 
        .Q(WX4714), .QN(n9396) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n10118), .CLK(n10387), 
        .Q(WX4716) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n10118), .CLK(n10387), 
        .Q(WX4718), .QN(n9659) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n10118), .CLK(n10387), 
        .Q(WX4720) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n10118), .CLK(n10387), 
        .Q(test_so40), .QN(n9830) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n10127), .CLK(n10378), 
        .Q(WX4724) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n10127), .CLK(n10378), 
        .Q(WX4726) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n10127), .CLK(n10378), 
        .Q(WX4728) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n10126), .CLK(n10379), 
        .Q(WX4730) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n10126), .CLK(n10379), 
        .Q(WX4732), .QN(n9665) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n10126), .CLK(n10379), 
        .Q(WX4734) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n10125), .CLK(n10380), 
        .Q(WX4736) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n10125), .CLK(n10380), 
        .Q(WX4738) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n10125), .CLK(n10380), 
        .Q(WX4740) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n10124), .CLK(n10381), 
        .Q(WX4742) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n10124), .CLK(n10381), 
        .Q(WX4744), .QN(n9671) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n10124), .CLK(n10381), 
        .Q(WX4746), .QN(n9509) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n10123), .CLK(n10382), 
        .Q(WX4748) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n10123), .CLK(n10382), 
        .Q(WX4750), .QN(n9673) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n10123), .CLK(n10382), 
        .Q(WX4752) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n10122), .CLK(n10383), 
        .Q(WX4754), .QN(n9675) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n10122), .CLK(n10383), 
        .Q(test_so41), .QN(n9850) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n10122), .CLK(n10383), 
        .Q(WX4758), .QN(n9676) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n10121), .CLK(n10384), 
        .Q(WX4760), .QN(n9677) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n10121), .CLK(n10384), 
        .Q(WX4762), .QN(n9678) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n10121), .CLK(n10384), 
        .Q(WX4764), .QN(n9679) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n10120), .CLK(n10385), 
        .Q(WX4766), .QN(n9680) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n10120), .CLK(n10385), 
        .Q(WX4768), .QN(n9681) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n10120), .CLK(n10385), 
        .Q(WX4770), .QN(n9510) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n10119), .CLK(n10386), 
        .Q(WX4772), .QN(n9682) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n10119), .CLK(n10386), 
        .Q(WX4774), .QN(n9683) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n10119), .CLK(n10386), 
        .Q(WX4776), .QN(n9684) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n10118), .CLK(n10387), 
        .Q(WX4778), .QN(n9522) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n10038), .CLK(n10467), 
        .Q(CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_3), .QN(DFF_739_n1) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n10037), .CLK(
        n10468), .Q(test_so42), .QN(n9858) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n10037), .CLK(n10468), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_10), .QN(DFF_746_n1) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n10037), .CLK(
        n10468), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_15), .QN(DFF_751_n1) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n10036), .CLK(
        n10469), .Q(test_so43), .QN(n9859) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n10036), .CLK(n10469), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n10036), .CLK(
        n10469), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n10035), .CLK(
        n10470), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n10118), .CLK(
        n10387), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n10118), .CLK(
        n10387), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n1049), .SI(CRC_OUT_6_31), .SE(n10118), .CLK(
        n10387), .Q(WX5657), .QN(n9492) );
  SDFFX1 DFF_769_Q_reg ( .D(n1050), .SI(WX5657), .SE(n10115), .CLK(n10390), 
        .Q(n8528) );
  SDFFX1 DFF_770_Q_reg ( .D(n1051), .SI(n8528), .SE(n10115), .CLK(n10390), .Q(
        n8527) );
  SDFFX1 DFF_771_Q_reg ( .D(n1052), .SI(n8527), .SE(n10115), .CLK(n10390), .Q(
        n8526) );
  SDFFX1 DFF_772_Q_reg ( .D(n1053), .SI(n8526), .SE(n10115), .CLK(n10390), .Q(
        n8525) );
  SDFFX1 DFF_773_Q_reg ( .D(n1054), .SI(n8525), .SE(n10115), .CLK(n10390), .Q(
        n8524) );
  SDFFX1 DFF_774_Q_reg ( .D(n1055), .SI(n8524), .SE(n10115), .CLK(n10390), .Q(
        n8523) );
  SDFFX1 DFF_775_Q_reg ( .D(n1056), .SI(n8523), .SE(n10115), .CLK(n10390), .Q(
        test_so44) );
  SDFFX1 DFF_776_Q_reg ( .D(n1057), .SI(test_si45), .SE(n10116), .CLK(n10389), 
        .Q(n8520) );
  SDFFX1 DFF_777_Q_reg ( .D(n1058), .SI(n8520), .SE(n10116), .CLK(n10389), .Q(
        n8519) );
  SDFFX1 DFF_778_Q_reg ( .D(n1059), .SI(n8519), .SE(n10116), .CLK(n10389), .Q(
        n8518) );
  SDFFX1 DFF_779_Q_reg ( .D(n1060), .SI(n8518), .SE(n10116), .CLK(n10389), .Q(
        n8517) );
  SDFFX1 DFF_780_Q_reg ( .D(n1061), .SI(n8517), .SE(n10116), .CLK(n10389), .Q(
        n8516) );
  SDFFX1 DFF_781_Q_reg ( .D(n1062), .SI(n8516), .SE(n10116), .CLK(n10389), .Q(
        n8515) );
  SDFFX1 DFF_782_Q_reg ( .D(n1063), .SI(n8515), .SE(n10116), .CLK(n10389), .Q(
        n8514) );
  SDFFX1 DFF_783_Q_reg ( .D(n1064), .SI(n8514), .SE(n10116), .CLK(n10389), .Q(
        n8513) );
  SDFFX1 DFF_784_Q_reg ( .D(n1065), .SI(n8513), .SE(n10116), .CLK(n10389), .Q(
        n8512) );
  SDFFX1 DFF_785_Q_reg ( .D(n1066), .SI(n8512), .SE(n10116), .CLK(n10389), .Q(
        n8511) );
  SDFFX1 DFF_786_Q_reg ( .D(n1067), .SI(n8511), .SE(n10116), .CLK(n10389), .Q(
        n8510) );
  SDFFX1 DFF_787_Q_reg ( .D(n1068), .SI(n8510), .SE(n10116), .CLK(n10389), .Q(
        n8509) );
  SDFFX1 DFF_788_Q_reg ( .D(n1069), .SI(n8509), .SE(n10117), .CLK(n10388), .Q(
        n8508) );
  SDFFX1 DFF_789_Q_reg ( .D(n1070), .SI(n8508), .SE(n10117), .CLK(n10388), .Q(
        n8507) );
  SDFFX1 DFF_790_Q_reg ( .D(n1071), .SI(n8507), .SE(n10117), .CLK(n10388), .Q(
        n8506) );
  SDFFX1 DFF_791_Q_reg ( .D(n1072), .SI(n8506), .SE(n10117), .CLK(n10388), .Q(
        n8505) );
  SDFFX1 DFF_792_Q_reg ( .D(n1073), .SI(n8505), .SE(n10117), .CLK(n10388), .Q(
        test_so45) );
  SDFFX1 DFF_793_Q_reg ( .D(n1074), .SI(test_si46), .SE(n10117), .CLK(n10388), 
        .Q(n8502) );
  SDFFX1 DFF_794_Q_reg ( .D(n1075), .SI(n8502), .SE(n10117), .CLK(n10388), .Q(
        n8501) );
  SDFFX1 DFF_795_Q_reg ( .D(n1076), .SI(n8501), .SE(n10117), .CLK(n10388), .Q(
        n8500) );
  SDFFX1 DFF_796_Q_reg ( .D(n1077), .SI(n8500), .SE(n10117), .CLK(n10388), .Q(
        n8499) );
  SDFFX1 DFF_797_Q_reg ( .D(n1078), .SI(n8499), .SE(n10117), .CLK(n10388), .Q(
        n8498) );
  SDFFX1 DFF_798_Q_reg ( .D(n1079), .SI(n8498), .SE(n10117), .CLK(n10388), .Q(
        n8497) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n10117), .CLK(n10388), 
        .Q(n8496) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n10115), .CLK(n10390), 
        .Q(n8495), .QN(n18397) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n10115), .CLK(n10390), 
        .Q(n8494), .QN(n18398) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n10115), .CLK(n10390), 
        .Q(n8493), .QN(n18399) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n10114), .CLK(n10391), 
        .Q(n8492), .QN(n18400) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n10114), .CLK(n10391), 
        .Q(n8491), .QN(n18401) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n10114), .CLK(n10391), 
        .Q(n8490), .QN(n18402) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n10114), .CLK(n10391), 
        .Q(n8489), .QN(n18403) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n10114), .CLK(n10391), 
        .Q(n8488), .QN(n18404) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n10114), .CLK(n10391), 
        .Q(n8487), .QN(n18405) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n10038), .CLK(n10467), 
        .Q(test_so46), .QN(n9842) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n10113), .CLK(n10392), 
        .Q(n8484), .QN(n18406) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n10113), .CLK(n10392), 
        .Q(n8483), .QN(n18407) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n10113), .CLK(n10392), 
        .Q(n8482), .QN(n18408) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n10112), .CLK(n10393), 
        .Q(n8481), .QN(n18409) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n10112), .CLK(n10393), 
        .Q(n8480), .QN(n18410) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n10112), .CLK(n10393), 
        .Q(n8479), .QN(n18411) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n10112), .CLK(n10393), 
        .Q(WX5849), .QN(n9394) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n10112), .CLK(n10393), 
        .Q(WX5851), .QN(n9392) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n10111), .CLK(n10394), 
        .Q(WX5853), .QN(n9390) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n10111), .CLK(n10394), 
        .Q(WX5855), .QN(n9388) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n10111), .CLK(n10394), 
        .Q(WX5857), .QN(n9386) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n10110), .CLK(n10395), 
        .Q(WX5859), .QN(n9384) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n10110), .CLK(n10395), 
        .Q(WX5861), .QN(n9382) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n10110), .CLK(n10395), 
        .Q(WX5863), .QN(n9380) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n10109), .CLK(n10396), 
        .Q(WX5865), .QN(n9378) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n10109), .CLK(n10396), 
        .Q(WX5867), .QN(n9376) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n10109), .CLK(n10396), 
        .Q(test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n10108), .CLK(n10397), 
        .Q(WX5871), .QN(n9373) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n10108), .CLK(n10397), 
        .Q(WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n10108), .CLK(n10397), 
        .Q(WX5875), .QN(n9369) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n10107), .CLK(n10398), 
        .Q(WX5877), .QN(n9368) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n10107), .CLK(n10398), 
        .Q(WX5879), .QN(n9366) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n10115), .CLK(n10390), 
        .Q(WX5881), .QN(n9011) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n10115), .CLK(n10390), 
        .Q(WX5883), .QN(n9157) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n10114), .CLK(n10391), 
        .Q(WX5885), .QN(n9155) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n10114), .CLK(n10391), 
        .Q(WX5887), .QN(n9153) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n10114), .CLK(n10391), 
        .Q(WX5889), .QN(n9151) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n10114), .CLK(n10391), 
        .Q(WX5891), .QN(n9149) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n10114), .CLK(n10391), 
        .Q(WX5893), .QN(n9147) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n10114), .CLK(n10391), 
        .Q(WX5895), .QN(n9145) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n10113), .CLK(n10392), 
        .Q(WX5897), .QN(n9143) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n10113), .CLK(n10392), 
        .Q(WX5899), .QN(n9141) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n10113), .CLK(n10392), 
        .Q(WX5901), .QN(n9139) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n10113), .CLK(n10392), 
        .Q(test_so48) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n10113), .CLK(n10392), 
        .Q(WX5905), .QN(n9136) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n10113), .CLK(n10392), 
        .Q(WX5907), .QN(n9135) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n10112), .CLK(n10393), 
        .Q(WX5909), .QN(n9133) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n10112), .CLK(n10393), 
        .Q(WX5911), .QN(n9131) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n10112), .CLK(n10393), 
        .Q(WX5913), .QN(n3689) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n10111), .CLK(n10394), 
        .Q(WX5915), .QN(n3687) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n10111), .CLK(n10394), 
        .Q(WX5917), .QN(n3685) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n10111), .CLK(n10394), 
        .Q(WX5919), .QN(n3683) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n10110), .CLK(n10395), 
        .Q(WX5921), .QN(n3681) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n10110), .CLK(n10395), 
        .Q(WX5923), .QN(n3679) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n10110), .CLK(n10395), 
        .Q(WX5925), .QN(n3677) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n10109), .CLK(n10396), 
        .Q(WX5927), .QN(n3675) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n10109), .CLK(n10396), 
        .Q(WX5929), .QN(n3673) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n10109), .CLK(n10396), 
        .Q(WX5931), .QN(n3671) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n10108), .CLK(n10397), 
        .Q(WX5933) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n10108), .CLK(n10397), 
        .Q(WX5935), .QN(n3667) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n10108), .CLK(n10397), 
        .Q(test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n10107), .CLK(n10398), 
        .Q(WX5939), .QN(n3663) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n10107), .CLK(n10398), 
        .Q(WX5941) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n10107), .CLK(n10398), 
        .Q(WX5943), .QN(n3659) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n10107), .CLK(n10398), 
        .Q(WX5945), .QN(n9012) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n10106), .CLK(n10399), 
        .Q(WX5947), .QN(n9158) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n10106), .CLK(n10399), 
        .Q(WX5949), .QN(n9156) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n10106), .CLK(n10399), 
        .Q(WX5951), .QN(n9154) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n10106), .CLK(n10399), 
        .Q(WX5953), .QN(n9152) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n10106), .CLK(n10399), 
        .Q(WX5955), .QN(n9150) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n10106), .CLK(n10399), 
        .Q(WX5957), .QN(n9148) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n10105), .CLK(n10400), 
        .Q(WX5959), .QN(n9146) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n10105), .CLK(n10400), 
        .Q(WX5961), .QN(n9144) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n10105), .CLK(n10400), 
        .Q(WX5963), .QN(n9142) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n10105), .CLK(n10400), 
        .Q(WX5965), .QN(n9140) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n10113), .CLK(n10392), 
        .Q(WX5967), .QN(n9138) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n10113), .CLK(n10392), 
        .Q(WX5969), .QN(n9137) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n10113), .CLK(n10392), 
        .Q(test_so50), .QN(n9869) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n10112), .CLK(n10393), 
        .Q(WX5973), .QN(n9134) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n10112), .CLK(n10393), 
        .Q(WX5975), .QN(n9132) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n10112), .CLK(n10393), 
        .Q(WX5977), .QN(n9395) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n10111), .CLK(n10394), 
        .Q(WX5979), .QN(n9393) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n10111), .CLK(n10394), 
        .Q(WX5981), .QN(n9391) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n10111), .CLK(n10394), 
        .Q(WX5983), .QN(n9389) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n10110), .CLK(n10395), 
        .Q(WX5985), .QN(n9387) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n10110), .CLK(n10395), 
        .Q(WX5987), .QN(n9385) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n10110), .CLK(n10395), 
        .Q(WX5989), .QN(n9383) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n10109), .CLK(n10396), 
        .Q(WX5991), .QN(n9381) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n10109), .CLK(n10396), 
        .Q(WX5993), .QN(n9379) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n10109), .CLK(n10396), 
        .Q(WX5995), .QN(n9377) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n10108), .CLK(n10397), 
        .Q(WX5997), .QN(n9375) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n10108), .CLK(n10397), 
        .Q(WX5999), .QN(n9374) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n10108), .CLK(n10397), 
        .Q(WX6001), .QN(n9372) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n10107), .CLK(n10398), 
        .Q(WX6003), .QN(n9370) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n10107), .CLK(n10398), 
        .Q(test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n10107), .CLK(n10398), 
        .Q(WX6007), .QN(n9367) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n10106), .CLK(n10399), 
        .Q(WX6009) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n10106), .CLK(n10399), 
        .Q(WX6011) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n10106), .CLK(n10399), 
        .Q(WX6013) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n10106), .CLK(n10399), 
        .Q(WX6015) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n10106), .CLK(n10399), 
        .Q(WX6017) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n10106), .CLK(n10399), 
        .Q(WX6019) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n10105), .CLK(n10400), 
        .Q(WX6021) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n10105), .CLK(n10400), 
        .Q(WX6023) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n10105), .CLK(n10400), 
        .Q(WX6025) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n10105), .CLK(n10400), 
        .Q(WX6027), .QN(n9639) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n10105), .CLK(n10400), 
        .Q(WX6029) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n10105), .CLK(n10400), 
        .Q(WX6031), .QN(n9641) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n10105), .CLK(n10400), 
        .Q(WX6033) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n10105), .CLK(n10400), 
        .Q(WX6035), .QN(n9643) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n10104), .CLK(n10401), 
        .Q(WX6037) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n10104), .CLK(n10401), 
        .Q(test_so52), .QN(n9848) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n10112), .CLK(n10393), 
        .Q(WX6041), .QN(n9645) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n10111), .CLK(n10394), 
        .Q(WX6043), .QN(n9646) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n10111), .CLK(n10394), 
        .Q(WX6045), .QN(n9647) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n10111), .CLK(n10394), 
        .Q(WX6047), .QN(n9648) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n10110), .CLK(n10395), 
        .Q(WX6049), .QN(n9507) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n10110), .CLK(n10395), 
        .Q(WX6051), .QN(n9649) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n10110), .CLK(n10395), 
        .Q(WX6053), .QN(n9650) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n10109), .CLK(n10396), 
        .Q(WX6055), .QN(n9651) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n10109), .CLK(n10396), 
        .Q(WX6057), .QN(n9652) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n10109), .CLK(n10396), 
        .Q(WX6059), .QN(n9653) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n10108), .CLK(n10397), 
        .Q(WX6061) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n10108), .CLK(n10397), 
        .Q(WX6063), .QN(n9508) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n10108), .CLK(n10397), 
        .Q(WX6065) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n10107), .CLK(n10398), 
        .Q(WX6067), .QN(n9656) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n10107), .CLK(n10398), 
        .Q(WX6069), .QN(n9657) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n10107), .CLK(n10398), 
        .Q(WX6071), .QN(n9521) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n10039), .CLK(n10466), 
        .Q(test_so53), .QN(n9856) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n10039), .CLK(n10466), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_3), .QN(DFF_931_n1) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_5_10), .QN(DFF_938_n1) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n10038), .CLK(
        n10467), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n10038), .CLK(
        n10467), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n10038), .CLK(
        n10467), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n10038), .CLK(
        n10467), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n10038), .CLK(
        n10467), .Q(CRC_OUT_5_15), .QN(DFF_943_n1) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n10038), .CLK(
        n10467), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n10038), .CLK(
        n10467), .Q(test_so54), .QN(n9857) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n10038), .CLK(n10467), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n10038), .CLK(
        n10467), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n10038), .CLK(
        n10467), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n10104), .CLK(
        n10401), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n10103), .CLK(
        n10402), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n1290), .SI(CRC_OUT_5_31), .SE(n10103), .CLK(
        n10402), .Q(WX6950), .QN(n9491) );
  SDFFX1 DFF_961_Q_reg ( .D(n1291), .SI(WX6950), .SE(n10101), .CLK(n10404), 
        .Q(n8470) );
  SDFFX1 DFF_962_Q_reg ( .D(n1292), .SI(n8470), .SE(n10101), .CLK(n10404), .Q(
        test_so55) );
  SDFFX1 DFF_963_Q_reg ( .D(n1293), .SI(test_si56), .SE(n10101), .CLK(n10404), 
        .Q(n8467) );
  SDFFX1 DFF_964_Q_reg ( .D(n1294), .SI(n8467), .SE(n10101), .CLK(n10404), .Q(
        n8466) );
  SDFFX1 DFF_965_Q_reg ( .D(n1295), .SI(n8466), .SE(n10101), .CLK(n10404), .Q(
        n8465) );
  SDFFX1 DFF_966_Q_reg ( .D(n1296), .SI(n8465), .SE(n10101), .CLK(n10404), .Q(
        n8464) );
  SDFFX1 DFF_967_Q_reg ( .D(n1297), .SI(n8464), .SE(n10101), .CLK(n10404), .Q(
        n8463) );
  SDFFX1 DFF_968_Q_reg ( .D(n1298), .SI(n8463), .SE(n10101), .CLK(n10404), .Q(
        n8462) );
  SDFFX1 DFF_969_Q_reg ( .D(n1299), .SI(n8462), .SE(n10101), .CLK(n10404), .Q(
        n8461) );
  SDFFX1 DFF_970_Q_reg ( .D(n1300), .SI(n8461), .SE(n10102), .CLK(n10403), .Q(
        n8460) );
  SDFFX1 DFF_971_Q_reg ( .D(n1301), .SI(n8460), .SE(n10102), .CLK(n10403), .Q(
        n8459) );
  SDFFX1 DFF_972_Q_reg ( .D(n1302), .SI(n8459), .SE(n10102), .CLK(n10403), .Q(
        n8458) );
  SDFFX1 DFF_973_Q_reg ( .D(n1303), .SI(n8458), .SE(n10102), .CLK(n10403), .Q(
        n8457) );
  SDFFX1 DFF_974_Q_reg ( .D(n1304), .SI(n8457), .SE(n10102), .CLK(n10403), .Q(
        n8456) );
  SDFFX1 DFF_975_Q_reg ( .D(n1305), .SI(n8456), .SE(n10102), .CLK(n10403), .Q(
        n8455) );
  SDFFX1 DFF_976_Q_reg ( .D(n1306), .SI(n8455), .SE(n10102), .CLK(n10403), .Q(
        n8454) );
  SDFFX1 DFF_977_Q_reg ( .D(n1307), .SI(n8454), .SE(n10102), .CLK(n10403), .Q(
        n8453) );
  SDFFX1 DFF_978_Q_reg ( .D(n1308), .SI(n8453), .SE(n10102), .CLK(n10403), .Q(
        n8452) );
  SDFFX1 DFF_979_Q_reg ( .D(n1309), .SI(n8452), .SE(n10102), .CLK(n10403), .Q(
        test_so56) );
  SDFFX1 DFF_980_Q_reg ( .D(n1310), .SI(test_si57), .SE(n10102), .CLK(n10403), 
        .Q(n8449) );
  SDFFX1 DFF_981_Q_reg ( .D(n1311), .SI(n8449), .SE(n10102), .CLK(n10403), .Q(
        n8448) );
  SDFFX1 DFF_982_Q_reg ( .D(n1312), .SI(n8448), .SE(n10103), .CLK(n10402), .Q(
        n8447) );
  SDFFX1 DFF_983_Q_reg ( .D(n1313), .SI(n8447), .SE(n10103), .CLK(n10402), .Q(
        n8446) );
  SDFFX1 DFF_984_Q_reg ( .D(n1314), .SI(n8446), .SE(n10103), .CLK(n10402), .Q(
        n8445) );
  SDFFX1 DFF_985_Q_reg ( .D(n1315), .SI(n8445), .SE(n10103), .CLK(n10402), .Q(
        n8444) );
  SDFFX1 DFF_986_Q_reg ( .D(n1316), .SI(n8444), .SE(n10103), .CLK(n10402), .Q(
        n8443) );
  SDFFX1 DFF_987_Q_reg ( .D(n1317), .SI(n8443), .SE(n10103), .CLK(n10402), .Q(
        n8442) );
  SDFFX1 DFF_988_Q_reg ( .D(n1318), .SI(n8442), .SE(n10103), .CLK(n10402), .Q(
        n8441) );
  SDFFX1 DFF_989_Q_reg ( .D(n1319), .SI(n8441), .SE(n10103), .CLK(n10402), .Q(
        n8440) );
  SDFFX1 DFF_990_Q_reg ( .D(n1320), .SI(n8440), .SE(n10103), .CLK(n10402), .Q(
        n8439) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n10103), .CLK(n10402), 
        .Q(n8438) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n10101), .CLK(n10404), 
        .Q(n8437), .QN(n18412) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n10100), .CLK(n10405), 
        .Q(n8436), .QN(n18413) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n10100), .CLK(n10405), 
        .Q(n8435), .QN(n18414) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n10100), .CLK(n10405), 
        .Q(n8434), .QN(n18415) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n10100), .CLK(n10405), 
        .Q(test_so57), .QN(n9841) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n10100), .CLK(n10405), 
        .Q(n8431), .QN(n18416) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n10100), .CLK(n10405), 
        .Q(n8430), .QN(n18417) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n10099), .CLK(n10406), 
        .Q(n8429), .QN(n18418) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n10099), .CLK(n10406), 
        .Q(n8428), .QN(n18419) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n10099), .CLK(n10406), 
        .Q(n8427), .QN(n18420) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n10099), .CLK(n10406), 
        .Q(n8426), .QN(n18421) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n10098), .CLK(n10407), 
        .Q(n8425), .QN(n18422) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n10098), .CLK(n10407), 
        .Q(n8424), .QN(n18423) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n10098), .CLK(n10407), 
        .Q(n8423), .QN(n18424) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n10097), .CLK(n10408), 
        .Q(n8422), .QN(n18425) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n10097), .CLK(n10408), 
        .Q(n8421), .QN(n18426) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n10097), .CLK(n10408), 
        .Q(WX7142), .QN(n9364) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n10096), .CLK(n10409), 
        .Q(WX7144), .QN(n9362) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n10096), .CLK(n10409), 
        .Q(WX7146), .QN(n9360) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n10096), .CLK(n10409), 
        .Q(WX7148), .QN(n9358) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n10095), .CLK(n10410), 
        .Q(WX7150), .QN(n9356) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n10095), .CLK(n10410), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n10095), .CLK(n10410), .Q(WX7154), .QN(n9353) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n10094), .CLK(n10411), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n10094), .CLK(n10411), 
        .Q(WX7158), .QN(n9349) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n10094), .CLK(n10411), 
        .Q(WX7160), .QN(n9348) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n10093), .CLK(n10412), 
        .Q(WX7162), .QN(n9346) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n10093), .CLK(n10412), 
        .Q(WX7164), .QN(n9344) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n10093), .CLK(n10412), 
        .Q(WX7166), .QN(n9342) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n10092), .CLK(n10413), 
        .Q(WX7168), .QN(n9340) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n10092), .CLK(n10413), 
        .Q(WX7170), .QN(n9338) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n10092), .CLK(n10413), 
        .Q(WX7172), .QN(n9336) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n10101), .CLK(n10404), 
        .Q(WX7174), .QN(n9009) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n10101), .CLK(n10404), 
        .Q(WX7176), .QN(n9129) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n10100), .CLK(n10405), 
        .Q(WX7178), .QN(n9127) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n10100), .CLK(n10405), 
        .Q(WX7180), .QN(n9125) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n10100), .CLK(n10405), 
        .Q(WX7182), .QN(n9123) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n10100), .CLK(n10405), 
        .Q(WX7184), .QN(n9121) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n10100), .CLK(n10405), 
        .Q(test_so59) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n10099), .CLK(n10406), .Q(WX7188), .QN(n9118) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n10099), .CLK(n10406), 
        .Q(WX7190), .QN(n9117) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n10099), .CLK(n10406), 
        .Q(WX7192), .QN(n9115) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n10099), .CLK(n10406), 
        .Q(WX7194), .QN(n9113) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n10098), .CLK(n10407), 
        .Q(WX7196), .QN(n9111) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n10098), .CLK(n10407), 
        .Q(WX7198), .QN(n9109) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n10098), .CLK(n10407), 
        .Q(WX7200), .QN(n9107) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n10097), .CLK(n10408), 
        .Q(WX7202), .QN(n9105) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n10097), .CLK(n10408), 
        .Q(WX7204), .QN(n9103) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n10097), .CLK(n10408), 
        .Q(WX7206), .QN(n3657) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n10096), .CLK(n10409), 
        .Q(WX7208), .QN(n3655) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n10096), .CLK(n10409), 
        .Q(WX7210), .QN(n3653) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n10096), .CLK(n10409), 
        .Q(WX7212), .QN(n3651) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n10095), .CLK(n10410), 
        .Q(WX7214), .QN(n3649) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n10095), .CLK(n10410), 
        .Q(WX7216) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n10095), .CLK(n10410), 
        .Q(WX7218), .QN(n3645) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n10094), .CLK(n10411), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n10094), .CLK(n10411), .Q(WX7222), .QN(n3641) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n10094), .CLK(n10411), 
        .Q(WX7224) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n10093), .CLK(n10412), 
        .Q(WX7226), .QN(n3637) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n10093), .CLK(n10412), 
        .Q(WX7228) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n10093), .CLK(n10412), 
        .Q(WX7230), .QN(n3633) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n10092), .CLK(n10413), 
        .Q(WX7232), .QN(n3631) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n10092), .CLK(n10413), 
        .Q(WX7234), .QN(n3629) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n10092), .CLK(n10413), 
        .Q(WX7236), .QN(n3627) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n10091), .CLK(n10414), 
        .Q(WX7238), .QN(n9010) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n10091), .CLK(n10414), 
        .Q(WX7240), .QN(n9130) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n10091), .CLK(n10414), 
        .Q(WX7242), .QN(n9128) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n10091), .CLK(n10414), 
        .Q(WX7244), .QN(n9126) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n10091), .CLK(n10414), 
        .Q(WX7246), .QN(n9124) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n10091), .CLK(n10414), 
        .Q(WX7248), .QN(n9122) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n10100), .CLK(n10405), 
        .Q(WX7250), .QN(n9120) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n10099), .CLK(n10406), 
        .Q(WX7252), .QN(n9119) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n10099), .CLK(n10406), 
        .Q(test_so61) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n10099), .CLK(n10406), .Q(WX7256), .QN(n9116) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n10099), .CLK(n10406), 
        .Q(WX7258), .QN(n9114) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n10098), .CLK(n10407), 
        .Q(WX7260), .QN(n9112) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n10098), .CLK(n10407), 
        .Q(WX7262), .QN(n9110) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n10098), .CLK(n10407), 
        .Q(WX7264), .QN(n9108) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n10097), .CLK(n10408), 
        .Q(WX7266), .QN(n9106) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n10097), .CLK(n10408), 
        .Q(WX7268), .QN(n9104) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n10097), .CLK(n10408), 
        .Q(WX7270), .QN(n9365) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n10096), .CLK(n10409), 
        .Q(WX7272), .QN(n9363) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n10096), .CLK(n10409), 
        .Q(WX7274), .QN(n9361) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n10096), .CLK(n10409), 
        .Q(WX7276), .QN(n9359) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n10095), .CLK(n10410), 
        .Q(WX7278), .QN(n9357) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n10095), .CLK(n10410), 
        .Q(WX7280), .QN(n9355) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n10095), .CLK(n10410), 
        .Q(WX7282), .QN(n9354) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n10094), .CLK(n10411), 
        .Q(WX7284), .QN(n9352) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n10094), .CLK(n10411), 
        .Q(WX7286), .QN(n9350) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n10094), .CLK(n10411), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n10093), .CLK(n10412), .Q(WX7290), .QN(n9347) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n10093), .CLK(n10412), 
        .Q(WX7292), .QN(n9345) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n10093), .CLK(n10412), 
        .Q(WX7294), .QN(n9343) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n10092), .CLK(n10413), 
        .Q(WX7296), .QN(n9341) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n10092), .CLK(n10413), 
        .Q(WX7298), .QN(n9339) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n10092), .CLK(n10413), 
        .Q(WX7300), .QN(n9337) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n10091), .CLK(n10414), 
        .Q(WX7302) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n10091), .CLK(n10414), 
        .Q(WX7304), .QN(n9604) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n10091), .CLK(n10414), 
        .Q(WX7306) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n10091), .CLK(n10414), 
        .Q(WX7308) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n10091), .CLK(n10414), 
        .Q(WX7310), .QN(n9607) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n10091), .CLK(n10414), 
        .Q(WX7312) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n10090), .CLK(n10415), 
        .Q(WX7314), .QN(n9609) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n10090), .CLK(n10415), 
        .Q(WX7316) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n10090), .CLK(n10415), 
        .Q(WX7318), .QN(n9611) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n10090), .CLK(n10415), 
        .Q(WX7320) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n10090), .CLK(n10415), 
        .Q(test_so63), .QN(n9829) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n10098), .CLK(n10407), .Q(WX7324) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n10098), .CLK(n10407), 
        .Q(WX7326) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n10098), .CLK(n10407), 
        .Q(WX7328) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n10097), .CLK(n10408), 
        .Q(WX7330) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n10097), .CLK(n10408), 
        .Q(WX7332), .QN(n9505) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n10097), .CLK(n10408), 
        .Q(WX7334), .QN(n9617) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n10096), .CLK(n10409), 
        .Q(WX7336), .QN(n9618) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n10096), .CLK(n10409), 
        .Q(WX7338), .QN(n9619) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n10096), .CLK(n10409), 
        .Q(WX7340), .QN(n9620) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n10095), .CLK(n10410), 
        .Q(WX7342), .QN(n9506) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n10095), .CLK(n10410), 
        .Q(WX7344) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n10095), .CLK(n10410), 
        .Q(WX7346), .QN(n9622) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n10094), .CLK(n10411), 
        .Q(WX7348) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n10094), .CLK(n10411), 
        .Q(WX7350), .QN(n9624) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n10094), .CLK(n10411), 
        .Q(WX7352) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n10093), .CLK(n10412), 
        .Q(WX7354), .QN(n9626) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n10093), .CLK(n10412), 
        .Q(test_so64), .QN(n9849) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n10093), .CLK(n10412), .Q(WX7358), .QN(n9627) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n10092), .CLK(n10413), 
        .Q(WX7360), .QN(n9628) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n10092), .CLK(n10413), 
        .Q(WX7362), .QN(n9629) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n10092), .CLK(n10413), 
        .Q(WX7364), .QN(n9520) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n10042), .CLK(n10463), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_3), .QN(DFF_1123_n1) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_10), .QN(DFF_1130_n1) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n10041), .CLK(
        n10464), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n10041), .CLK(
        n10464), .Q(test_so65), .QN(n9854) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n10040), .CLK(n10465), .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_15), .QN(DFF_1135_n1) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n10040), .CLK(
        n10465), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n10039), .CLK(
        n10466), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n10090), .CLK(
        n10415), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n10090), .CLK(
        n10415), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n10090), .CLK(
        n10415), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n10090), .CLK(
        n10415), .Q(test_so66), .QN(n9855) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n10090), .CLK(n10415), .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n10090), .CLK(
        n10415), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n1530), .SI(CRC_OUT_4_31), .SE(n10090), .CLK(
        n10415), .Q(WX8243), .QN(n9490) );
  SDFFX1 DFF_1153_Q_reg ( .D(n1531), .SI(WX8243), .SE(n10087), .CLK(n10418), 
        .Q(n8411) );
  SDFFX1 DFF_1154_Q_reg ( .D(n1532), .SI(n8411), .SE(n10087), .CLK(n10418), 
        .Q(n8410) );
  SDFFX1 DFF_1155_Q_reg ( .D(n1533), .SI(n8410), .SE(n10087), .CLK(n10418), 
        .Q(n8409) );
  SDFFX1 DFF_1156_Q_reg ( .D(n1534), .SI(n8409), .SE(n10087), .CLK(n10418), 
        .Q(n8408) );
  SDFFX1 DFF_1157_Q_reg ( .D(n1535), .SI(n8408), .SE(n10087), .CLK(n10418), 
        .Q(n8407) );
  SDFFX1 DFF_1158_Q_reg ( .D(n1536), .SI(n8407), .SE(n10087), .CLK(n10418), 
        .Q(n8406) );
  SDFFX1 DFF_1159_Q_reg ( .D(n1537), .SI(n8406), .SE(n10087), .CLK(n10418), 
        .Q(n8405) );
  SDFFX1 DFF_1160_Q_reg ( .D(n1538), .SI(n8405), .SE(n10088), .CLK(n10417), 
        .Q(n8404) );
  SDFFX1 DFF_1161_Q_reg ( .D(n1539), .SI(n8404), .SE(n10088), .CLK(n10417), 
        .Q(n8403) );
  SDFFX1 DFF_1162_Q_reg ( .D(n1540), .SI(n8403), .SE(n10088), .CLK(n10417), 
        .Q(n8402) );
  SDFFX1 DFF_1163_Q_reg ( .D(n1541), .SI(n8402), .SE(n10088), .CLK(n10417), 
        .Q(n8401) );
  SDFFX1 DFF_1164_Q_reg ( .D(n1542), .SI(n8401), .SE(n10088), .CLK(n10417), 
        .Q(n8400) );
  SDFFX1 DFF_1165_Q_reg ( .D(n1543), .SI(n8400), .SE(n10088), .CLK(n10417), 
        .Q(n8399) );
  SDFFX1 DFF_1166_Q_reg ( .D(n1544), .SI(n8399), .SE(n10088), .CLK(n10417), 
        .Q(test_so67) );
  SDFFX1 DFF_1167_Q_reg ( .D(n1545), .SI(test_si68), .SE(n10088), .CLK(n10417), 
        .Q(n8396) );
  SDFFX1 DFF_1168_Q_reg ( .D(n1546), .SI(n8396), .SE(n10088), .CLK(n10417), 
        .Q(n8395) );
  SDFFX1 DFF_1169_Q_reg ( .D(n1547), .SI(n8395), .SE(n10088), .CLK(n10417), 
        .Q(n8394) );
  SDFFX1 DFF_1170_Q_reg ( .D(n1548), .SI(n8394), .SE(n10088), .CLK(n10417), 
        .Q(n8393) );
  SDFFX1 DFF_1171_Q_reg ( .D(n1549), .SI(n8393), .SE(n10088), .CLK(n10417), 
        .Q(n8392) );
  SDFFX1 DFF_1172_Q_reg ( .D(n1550), .SI(n8392), .SE(n10089), .CLK(n10416), 
        .Q(n8391) );
  SDFFX1 DFF_1173_Q_reg ( .D(n1551), .SI(n8391), .SE(n10089), .CLK(n10416), 
        .Q(n8390) );
  SDFFX1 DFF_1174_Q_reg ( .D(n1552), .SI(n8390), .SE(n10089), .CLK(n10416), 
        .Q(n8389) );
  SDFFX1 DFF_1175_Q_reg ( .D(n1553), .SI(n8389), .SE(n10089), .CLK(n10416), 
        .Q(n8388) );
  SDFFX1 DFF_1176_Q_reg ( .D(n1554), .SI(n8388), .SE(n10089), .CLK(n10416), 
        .Q(n8387) );
  SDFFX1 DFF_1177_Q_reg ( .D(n1555), .SI(n8387), .SE(n10089), .CLK(n10416), 
        .Q(n8386) );
  SDFFX1 DFF_1178_Q_reg ( .D(n1556), .SI(n8386), .SE(n10089), .CLK(n10416), 
        .Q(n8385) );
  SDFFX1 DFF_1179_Q_reg ( .D(n1557), .SI(n8385), .SE(n10089), .CLK(n10416), 
        .Q(n8384) );
  SDFFX1 DFF_1180_Q_reg ( .D(n1558), .SI(n8384), .SE(n10089), .CLK(n10416), 
        .Q(n8383) );
  SDFFX1 DFF_1181_Q_reg ( .D(n1559), .SI(n8383), .SE(n10089), .CLK(n10416), 
        .Q(n8382) );
  SDFFX1 DFF_1182_Q_reg ( .D(n1560), .SI(n8382), .SE(n10089), .CLK(n10416), 
        .Q(n8381) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n10089), .CLK(n10416), 
        .Q(test_so68) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n10042), .CLK(n10463), .Q(n8378), .QN(n18427) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n10087), .CLK(n10418), 
        .Q(n8377), .QN(n18428) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n10087), .CLK(n10418), 
        .Q(n8376), .QN(n18429) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n10086), .CLK(n10419), 
        .Q(n8375), .QN(n18430) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n10086), .CLK(n10419), 
        .Q(n8374), .QN(n18431) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n10086), .CLK(n10419), 
        .Q(n8373), .QN(n18432) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n10086), .CLK(n10419), 
        .Q(n8372), .QN(n18433) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n10085), .CLK(n10420), 
        .Q(n8371), .QN(n18434) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n10085), .CLK(n10420), 
        .Q(n8370), .QN(n18435) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n10084), .CLK(n10421), 
        .Q(n8369), .QN(n18436) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n10084), .CLK(n10421), 
        .Q(n8368), .QN(n18437) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n10084), .CLK(n10421), 
        .Q(n8367), .QN(n18438) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n10084), .CLK(n10421), 
        .Q(n8366), .QN(n18439) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n10083), .CLK(n10422), 
        .Q(n8365), .QN(n18440) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n10083), .CLK(n10422), 
        .Q(n8364), .QN(n18441) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n10082), .CLK(n10423), 
        .Q(n8363), .QN(n18442) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n10082), .CLK(n10423), 
        .Q(test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n10082), .CLK(n10423), .Q(WX8437), .QN(n9333) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n10082), .CLK(n10423), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n10081), .CLK(n10424), 
        .Q(WX8441), .QN(n9329) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n10081), .CLK(n10424), 
        .Q(WX8443), .QN(n9328) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n10081), .CLK(n10424), 
        .Q(WX8445), .QN(n9326) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n10080), .CLK(n10425), 
        .Q(WX8447), .QN(n9324) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n10080), .CLK(n10425), 
        .Q(WX8449), .QN(n9322) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n10080), .CLK(n10425), 
        .Q(WX8451), .QN(n9320) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n10079), .CLK(n10426), 
        .Q(WX8453), .QN(n9318) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n10079), .CLK(n10426), 
        .Q(WX8455), .QN(n9316) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n10079), .CLK(n10426), 
        .Q(WX8457), .QN(n9314) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n10078), .CLK(n10427), 
        .Q(WX8459), .QN(n9312) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n10078), .CLK(n10427), 
        .Q(WX8461), .QN(n9310) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n10078), .CLK(n10427), 
        .Q(WX8463), .QN(n9308) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n10077), .CLK(n10428), 
        .Q(WX8465), .QN(n9306) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n10077), .CLK(n10428), 
        .Q(WX8467), .QN(n9007) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n10087), .CLK(n10418), 
        .Q(test_so70) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n10086), .CLK(n10419), .Q(WX8471), .QN(n9100) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n10086), .CLK(n10419), 
        .Q(WX8473), .QN(n9099) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n10086), .CLK(n10419), 
        .Q(WX8475), .QN(n9097) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n10086), .CLK(n10419), 
        .Q(WX8477), .QN(n9095) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n10086), .CLK(n10419), 
        .Q(WX8479), .QN(n9093) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n10085), .CLK(n10420), 
        .Q(WX8481), .QN(n9091) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n10085), .CLK(n10420), 
        .Q(WX8483), .QN(n9089) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n10085), .CLK(n10420), 
        .Q(WX8485), .QN(n9087) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n10084), .CLK(n10421), 
        .Q(WX8487), .QN(n9085) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n10084), .CLK(n10421), 
        .Q(WX8489), .QN(n9083) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n10084), .CLK(n10421), 
        .Q(WX8491), .QN(n9081) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n10083), .CLK(n10422), 
        .Q(WX8493), .QN(n9079) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n10083), .CLK(n10422), 
        .Q(WX8495), .QN(n9077) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n10083), .CLK(n10422), 
        .Q(WX8497), .QN(n9075) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n10082), .CLK(n10423), 
        .Q(WX8499) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n10082), .CLK(n10423), 
        .Q(WX8501), .QN(n3623) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n10082), .CLK(n10423), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n10081), .CLK(n10424), .Q(WX8505), .QN(n3619) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n10081), .CLK(n10424), 
        .Q(WX8507) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n10081), .CLK(n10424), 
        .Q(WX8509), .QN(n3615) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n10080), .CLK(n10425), 
        .Q(WX8511) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n10080), .CLK(n10425), 
        .Q(WX8513), .QN(n3611) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n10080), .CLK(n10425), 
        .Q(WX8515), .QN(n3609) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n10079), .CLK(n10426), 
        .Q(WX8517), .QN(n3607) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n10079), .CLK(n10426), 
        .Q(WX8519), .QN(n3605) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n10079), .CLK(n10426), 
        .Q(WX8521), .QN(n3603) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n10078), .CLK(n10427), 
        .Q(WX8523), .QN(n3601) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n10078), .CLK(n10427), 
        .Q(WX8525), .QN(n3599) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n10078), .CLK(n10427), 
        .Q(WX8527), .QN(n3597) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n10077), .CLK(n10428), 
        .Q(WX8529), .QN(n3595) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n10077), .CLK(n10428), 
        .Q(WX8531), .QN(n9008) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n10087), .CLK(n10418), 
        .Q(WX8533), .QN(n9102) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n10087), .CLK(n10418), 
        .Q(WX8535), .QN(n9101) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n10086), .CLK(n10419), 
        .Q(test_so72) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n10086), .CLK(n10419), .Q(WX8539), .QN(n9098) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n10086), .CLK(n10419), 
        .Q(WX8541), .QN(n9096) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n10085), .CLK(n10420), 
        .Q(WX8543), .QN(n9094) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n10085), .CLK(n10420), 
        .Q(WX8545), .QN(n9092) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n10085), .CLK(n10420), 
        .Q(WX8547), .QN(n9090) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n10085), .CLK(n10420), 
        .Q(WX8549), .QN(n9088) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n10084), .CLK(n10421), 
        .Q(WX8551), .QN(n9086) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n10084), .CLK(n10421), 
        .Q(WX8553), .QN(n9084) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n10083), .CLK(n10422), 
        .Q(WX8555), .QN(n9082) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n10083), .CLK(n10422), 
        .Q(WX8557), .QN(n9080) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n10083), .CLK(n10422), 
        .Q(WX8559), .QN(n9078) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n10083), .CLK(n10422), 
        .Q(WX8561), .QN(n9076) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n10082), .CLK(n10423), 
        .Q(WX8563), .QN(n9335) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n10082), .CLK(n10423), 
        .Q(WX8565), .QN(n9334) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n10081), .CLK(n10424), 
        .Q(WX8567), .QN(n9332) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n10081), .CLK(n10424), 
        .Q(WX8569), .QN(n9330) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n10081), .CLK(n10424), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n10080), .CLK(n10425), .Q(WX8573), .QN(n9327) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n10080), .CLK(n10425), 
        .Q(WX8575), .QN(n9325) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n10080), .CLK(n10425), 
        .Q(WX8577), .QN(n9323) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n10079), .CLK(n10426), 
        .Q(WX8579), .QN(n9321) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n10079), .CLK(n10426), 
        .Q(WX8581), .QN(n9319) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n10079), .CLK(n10426), 
        .Q(WX8583), .QN(n9317) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n10078), .CLK(n10427), 
        .Q(WX8585), .QN(n9315) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n10078), .CLK(n10427), 
        .Q(WX8587), .QN(n9313) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n10078), .CLK(n10427), 
        .Q(WX8589), .QN(n9311) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n10077), .CLK(n10428), 
        .Q(WX8591), .QN(n9309) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n10077), .CLK(n10428), 
        .Q(WX8593), .QN(n9307) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n10077), .CLK(n10428), 
        .Q(WX8595) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n10077), .CLK(n10428), 
        .Q(WX8597), .QN(n9578) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n10077), .CLK(n10428), 
        .Q(WX8599) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n10077), .CLK(n10428), 
        .Q(WX8601), .QN(n9580) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n10076), .CLK(n10429), 
        .Q(WX8603) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n10076), .CLK(n10429), 
        .Q(test_so74), .QN(n9828) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n10085), .CLK(n10420), .Q(WX8607), .QN(n9582) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n10085), .CLK(n10420), 
        .Q(WX8609) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n10085), .CLK(n10420), 
        .Q(WX8611) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n10084), .CLK(n10421), 
        .Q(WX8613) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n10084), .CLK(n10421), 
        .Q(WX8615) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n10084), .CLK(n10421), 
        .Q(WX8617) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n10083), .CLK(n10422), 
        .Q(WX8619) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n10083), .CLK(n10422), 
        .Q(WX8621) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n10083), .CLK(n10422), 
        .Q(WX8623) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n10082), .CLK(n10423), 
        .Q(WX8625), .QN(n9502) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n10082), .CLK(n10423), 
        .Q(WX8627) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n10082), .CLK(n10423), 
        .Q(WX8629), .QN(n9592) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n10081), .CLK(n10424), 
        .Q(WX8631) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n10081), .CLK(n10424), 
        .Q(WX8633), .QN(n9594) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n10081), .CLK(n10424), 
        .Q(WX8635), .QN(n9503) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n10080), .CLK(n10425), 
        .Q(WX8637), .QN(n9595) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n10080), .CLK(n10425), 
        .Q(test_so75), .QN(n9834) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n10080), .CLK(n10425), .Q(WX8641), .QN(n9596) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n10079), .CLK(n10426), 
        .Q(WX8643), .QN(n9597) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n10079), .CLK(n10426), 
        .Q(WX8645), .QN(n9598) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n10079), .CLK(n10426), 
        .Q(WX8647), .QN(n9599) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n10078), .CLK(n10427), 
        .Q(WX8649), .QN(n9504) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n10078), .CLK(n10427), 
        .Q(WX8651), .QN(n9600) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n10078), .CLK(n10427), 
        .Q(WX8653), .QN(n9601) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n10077), .CLK(n10428), 
        .Q(WX8655), .QN(n9602) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n10077), .CLK(n10428), 
        .Q(WX8657), .QN(n9519) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n10044), .CLK(n10461), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n10044), .CLK(
        n10461), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n10044), .CLK(
        n10461), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n10044), .CLK(
        n10461), .Q(CRC_OUT_3_3), .QN(DFF_1315_n1) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n10044), .CLK(
        n10461), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n10044), .CLK(
        n10461), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n10044), .CLK(
        n10461), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n10044), .CLK(
        n10461), .Q(test_so76), .QN(n9852) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n10044), .CLK(n10461), .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_10), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_15), .QN(DFF_1327_n1) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n10043), .CLK(
        n10462), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n10042), .CLK(
        n10463), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n10042), .CLK(
        n10463), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n10042), .CLK(
        n10463), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n10042), .CLK(
        n10463), .Q(test_so77), .QN(n9853) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n10042), .CLK(n10463), .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n10042), .CLK(
        n10463), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n10042), .CLK(
        n10463), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n10042), .CLK(
        n10463), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n10042), .CLK(
        n10463), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n10042), .CLK(
        n10463), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n10076), .CLK(
        n10429), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n1771), .SI(CRC_OUT_3_31), .SE(n10076), .CLK(
        n10429), .Q(WX9536), .QN(n9489) );
  SDFFX1 DFF_1345_Q_reg ( .D(n1772), .SI(WX9536), .SE(n10074), .CLK(n10431), 
        .Q(n8353) );
  SDFFX1 DFF_1346_Q_reg ( .D(n1773), .SI(n8353), .SE(n10074), .CLK(n10431), 
        .Q(n8352) );
  SDFFX1 DFF_1347_Q_reg ( .D(n1774), .SI(n8352), .SE(n10074), .CLK(n10431), 
        .Q(n8351) );
  SDFFX1 DFF_1348_Q_reg ( .D(n1775), .SI(n8351), .SE(n10074), .CLK(n10431), 
        .Q(n8350) );
  SDFFX1 DFF_1349_Q_reg ( .D(n1776), .SI(n8350), .SE(n10074), .CLK(n10431), 
        .Q(n8349) );
  SDFFX1 DFF_1350_Q_reg ( .D(n1777), .SI(n8349), .SE(n10074), .CLK(n10431), 
        .Q(n8348) );
  SDFFX1 DFF_1351_Q_reg ( .D(n1778), .SI(n8348), .SE(n10074), .CLK(n10431), 
        .Q(n8347) );
  SDFFX1 DFF_1352_Q_reg ( .D(n1779), .SI(n8347), .SE(n10074), .CLK(n10431), 
        .Q(n8346) );
  SDFFX1 DFF_1353_Q_reg ( .D(n1780), .SI(n8346), .SE(n10074), .CLK(n10431), 
        .Q(test_so78) );
  SDFFX1 DFF_1354_Q_reg ( .D(n1781), .SI(test_si79), .SE(n10074), .CLK(n10431), 
        .Q(n8343) );
  SDFFX1 DFF_1355_Q_reg ( .D(n1782), .SI(n8343), .SE(n10074), .CLK(n10431), 
        .Q(n8342) );
  SDFFX1 DFF_1356_Q_reg ( .D(n1783), .SI(n8342), .SE(n10075), .CLK(n10430), 
        .Q(n8341) );
  SDFFX1 DFF_1357_Q_reg ( .D(n1784), .SI(n8341), .SE(n10075), .CLK(n10430), 
        .Q(n8340) );
  SDFFX1 DFF_1358_Q_reg ( .D(n1785), .SI(n8340), .SE(n10075), .CLK(n10430), 
        .Q(n8339) );
  SDFFX1 DFF_1359_Q_reg ( .D(n1786), .SI(n8339), .SE(n10075), .CLK(n10430), 
        .Q(n8338) );
  SDFFX1 DFF_1360_Q_reg ( .D(n1787), .SI(n8338), .SE(n10075), .CLK(n10430), 
        .Q(n8337) );
  SDFFX1 DFF_1361_Q_reg ( .D(n1788), .SI(n8337), .SE(n10075), .CLK(n10430), 
        .Q(n8336) );
  SDFFX1 DFF_1362_Q_reg ( .D(n1789), .SI(n8336), .SE(n10075), .CLK(n10430), 
        .Q(n8335) );
  SDFFX1 DFF_1363_Q_reg ( .D(n1790), .SI(n8335), .SE(n10075), .CLK(n10430), 
        .Q(n8334) );
  SDFFX1 DFF_1364_Q_reg ( .D(n1791), .SI(n8334), .SE(n10075), .CLK(n10430), 
        .Q(n8333) );
  SDFFX1 DFF_1365_Q_reg ( .D(n1792), .SI(n8333), .SE(n10075), .CLK(n10430), 
        .Q(n8332) );
  SDFFX1 DFF_1366_Q_reg ( .D(n1793), .SI(n8332), .SE(n10075), .CLK(n10430), 
        .Q(n8331) );
  SDFFX1 DFF_1367_Q_reg ( .D(n1794), .SI(n8331), .SE(n10075), .CLK(n10430), 
        .Q(n8330) );
  SDFFX1 DFF_1368_Q_reg ( .D(n1795), .SI(n8330), .SE(n10076), .CLK(n10429), 
        .Q(n8329) );
  SDFFX1 DFF_1369_Q_reg ( .D(n1796), .SI(n8329), .SE(n10076), .CLK(n10429), 
        .Q(n8328) );
  SDFFX1 DFF_1370_Q_reg ( .D(n1797), .SI(n8328), .SE(n10076), .CLK(n10429), 
        .Q(test_so79) );
  SDFFX1 DFF_1371_Q_reg ( .D(n1798), .SI(test_si80), .SE(n10076), .CLK(n10429), 
        .Q(n8325) );
  SDFFX1 DFF_1372_Q_reg ( .D(n1799), .SI(n8325), .SE(n10076), .CLK(n10429), 
        .Q(n8324) );
  SDFFX1 DFF_1373_Q_reg ( .D(n1800), .SI(n8324), .SE(n10076), .CLK(n10429), 
        .Q(n8323) );
  SDFFX1 DFF_1374_Q_reg ( .D(n1801), .SI(n8323), .SE(n10076), .CLK(n10429), 
        .Q(n8322) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n10076), .CLK(n10429), 
        .Q(n8321) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n10074), .CLK(n10431), 
        .Q(n8320), .QN(n18443) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n10073), .CLK(n10432), 
        .Q(n8319), .QN(n18444) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n10073), .CLK(n10432), 
        .Q(n8318), .QN(n18445) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n10073), .CLK(n10432), 
        .Q(n8317), .QN(n18446) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n10073), .CLK(n10432), 
        .Q(n8316), .QN(n18447) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n10073), .CLK(n10432), 
        .Q(n8315), .QN(n18448) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n10073), .CLK(n10432), 
        .Q(n8314), .QN(n18449) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n10072), .CLK(n10433), 
        .Q(n8313), .QN(n18450) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n10072), .CLK(n10433), 
        .Q(n8312), .QN(n18451) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n10072), .CLK(n10433), 
        .Q(n8311), .QN(n18452) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n10072), .CLK(n10433), 
        .Q(n8310), .QN(n18453) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n10044), .CLK(n10461), 
        .Q(test_so80), .QN(n9840) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n10072), .CLK(n10433), .Q(n8307), .QN(n18454) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n10071), .CLK(n10434), 
        .Q(n8306), .QN(n18455) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n10071), .CLK(n10434), 
        .Q(n8305), .QN(n18456) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n10071), .CLK(n10434), 
        .Q(n8304), .QN(n18457) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n10071), .CLK(n10434), 
        .Q(WX9728), .QN(n9304) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n10070), .CLK(n10435), 
        .Q(WX9730), .QN(n9302) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n10070), .CLK(n10435), 
        .Q(WX9732), .QN(n9300) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n10070), .CLK(n10435), 
        .Q(WX9734), .QN(n9298) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n10070), .CLK(n10435), 
        .Q(WX9736), .QN(n9296) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n10069), .CLK(n10436), 
        .Q(WX9738), .QN(n9294) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n10069), .CLK(n10436), 
        .Q(WX9740), .QN(n9292) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n10069), .CLK(n10436), 
        .Q(WX9742), .QN(n9290) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n10068), .CLK(n10437), 
        .Q(WX9744), .QN(n9288) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n10068), .CLK(n10437), 
        .Q(WX9746), .QN(n9286) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n10068), .CLK(n10437), 
        .Q(WX9748), .QN(n9284) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n10067), .CLK(n10438), 
        .Q(WX9750), .QN(n9282) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n10067), .CLK(n10438), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n10066), .CLK(n10439), .Q(WX9754), .QN(n9279) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n10066), .CLK(n10439), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n10066), .CLK(n10439), 
        .Q(WX9758), .QN(n9275) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n10073), .CLK(n10432), 
        .Q(WX9760), .QN(n9005) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n10073), .CLK(n10432), 
        .Q(WX9762), .QN(n9073) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n10073), .CLK(n10432), 
        .Q(WX9764), .QN(n9071) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n10073), .CLK(n10432), 
        .Q(WX9766), .QN(n9069) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n10073), .CLK(n10432), 
        .Q(WX9768), .QN(n9067) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n10073), .CLK(n10432), 
        .Q(WX9770), .QN(n9065) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n10072), .CLK(n10433), 
        .Q(WX9772), .QN(n9063) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n10072), .CLK(n10433), 
        .Q(WX9774), .QN(n9061) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n10072), .CLK(n10433), 
        .Q(WX9776), .QN(n9059) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n10072), .CLK(n10433), 
        .Q(WX9778), .QN(n9057) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n10072), .CLK(n10433), 
        .Q(WX9780), .QN(n9055) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n10072), .CLK(n10433), 
        .Q(WX9782), .QN(n9053) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n10072), .CLK(n10433), 
        .Q(WX9784), .QN(n9051) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n10071), .CLK(n10434), 
        .Q(test_so82), .QN(n9868) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n10071), .CLK(n10434), .Q(WX9788), .QN(n9048) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n10071), .CLK(n10434), 
        .Q(WX9790), .QN(n9047) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n10071), .CLK(n10434), 
        .Q(WX9792), .QN(n3593) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n10070), .CLK(n10435), 
        .Q(WX9794) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n10070), .CLK(n10435), 
        .Q(WX9796), .QN(n3589) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n10070), .CLK(n10435), 
        .Q(WX9798), .QN(n3587) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n10069), .CLK(n10436), 
        .Q(WX9800), .QN(n3585) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n10069), .CLK(n10436), 
        .Q(WX9802), .QN(n3583) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n10069), .CLK(n10436), 
        .Q(WX9804), .QN(n3581) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n10068), .CLK(n10437), 
        .Q(WX9806), .QN(n3579) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n10068), .CLK(n10437), 
        .Q(WX9808), .QN(n3577) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n10068), .CLK(n10437), 
        .Q(WX9810), .QN(n3575) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n10067), .CLK(n10438), 
        .Q(WX9812), .QN(n3573) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n10067), .CLK(n10438), 
        .Q(WX9814), .QN(n3571) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n10067), .CLK(n10438), 
        .Q(WX9816) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n10067), .CLK(n10438), 
        .Q(WX9818), .QN(n3567) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n10066), .CLK(n10439), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n10066), .CLK(n10439), .Q(WX9822), .QN(n3563) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n10066), .CLK(n10439), 
        .Q(WX9824), .QN(n9006) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n10065), .CLK(n10440), 
        .Q(WX9826), .QN(n9074) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n10065), .CLK(n10440), 
        .Q(WX9828), .QN(n9072) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n10065), .CLK(n10440), 
        .Q(WX9830), .QN(n9070) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n10065), .CLK(n10440), 
        .Q(WX9832), .QN(n9068) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n10065), .CLK(n10440), 
        .Q(WX9834), .QN(n9066) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n10065), .CLK(n10440), 
        .Q(WX9836), .QN(n9064) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n10064), .CLK(n10441), 
        .Q(WX9838), .QN(n9062) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n10064), .CLK(n10441), 
        .Q(WX9840), .QN(n9060) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n10064), .CLK(n10441), 
        .Q(WX9842), .QN(n9058) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n10064), .CLK(n10441), 
        .Q(WX9844), .QN(n9056) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n10064), .CLK(n10441), 
        .Q(WX9846), .QN(n9054) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n10064), .CLK(n10441), 
        .Q(WX9848), .QN(n9052) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n10071), .CLK(n10434), 
        .Q(WX9850), .QN(n9050) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n10071), .CLK(n10434), 
        .Q(WX9852), .QN(n9049) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n10071), .CLK(n10434), 
        .Q(test_so84), .QN(n9867) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n10071), .CLK(n10434), .Q(WX9856), .QN(n9305) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n10070), .CLK(n10435), 
        .Q(WX9858), .QN(n9303) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n10070), .CLK(n10435), 
        .Q(WX9860), .QN(n9301) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n10070), .CLK(n10435), 
        .Q(WX9862), .QN(n9299) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n10069), .CLK(n10436), 
        .Q(WX9864), .QN(n9297) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n10069), .CLK(n10436), 
        .Q(WX9866), .QN(n9295) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n10069), .CLK(n10436), 
        .Q(WX9868), .QN(n9293) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n10068), .CLK(n10437), 
        .Q(WX9870), .QN(n9291) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n10068), .CLK(n10437), 
        .Q(WX9872), .QN(n9289) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n10068), .CLK(n10437), 
        .Q(WX9874), .QN(n9287) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n10067), .CLK(n10438), 
        .Q(WX9876), .QN(n9285) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n10067), .CLK(n10438), 
        .Q(WX9878), .QN(n9283) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n10067), .CLK(n10438), 
        .Q(WX9880), .QN(n9281) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n10066), .CLK(n10439), 
        .Q(WX9882), .QN(n9280) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n10066), .CLK(n10439), 
        .Q(WX9884), .QN(n9278) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n10066), .CLK(n10439), 
        .Q(WX9886), .QN(n9276) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n10065), .CLK(n10440), 
        .Q(test_so85), .QN(n9833) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n10065), .CLK(n10440), .Q(WX9890) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n10065), .CLK(n10440), 
        .Q(WX9892) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n10065), .CLK(n10440), 
        .Q(WX9894) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n10065), .CLK(n10440), 
        .Q(WX9896) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n10065), .CLK(n10440), 
        .Q(WX9898) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n10064), .CLK(n10441), 
        .Q(WX9900) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n10064), .CLK(n10441), 
        .Q(WX9902) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n10064), .CLK(n10441), 
        .Q(WX9904) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n10064), .CLK(n10441), 
        .Q(WX9906) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n10064), .CLK(n10441), 
        .Q(WX9908) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n10064), .CLK(n10441), 
        .Q(WX9910), .QN(n9561) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n10063), .CLK(n10442), 
        .Q(WX9912) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n10063), .CLK(n10442), 
        .Q(WX9914), .QN(n9563) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n10063), .CLK(n10442), 
        .Q(WX9916) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n10063), .CLK(n10442), 
        .Q(WX9918), .QN(n9499) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n10063), .CLK(n10442), 
        .Q(WX9920), .QN(n9565) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n10063), .CLK(n10442), 
        .Q(test_so86), .QN(n9837) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n10070), .CLK(n10435), .Q(WX9924), .QN(n9566) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n10070), .CLK(n10435), 
        .Q(WX9926), .QN(n9567) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n10069), .CLK(n10436), 
        .Q(WX9928), .QN(n9500) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n10069), .CLK(n10436), 
        .Q(WX9930), .QN(n9568) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n10069), .CLK(n10436), 
        .Q(WX9932), .QN(n9569) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n10068), .CLK(n10437), 
        .Q(WX9934), .QN(n9570) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n10068), .CLK(n10437), 
        .Q(WX9936), .QN(n9571) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n10068), .CLK(n10437), 
        .Q(WX9938), .QN(n9572) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n10067), .CLK(n10438), 
        .Q(WX9940), .QN(n9573) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n10067), .CLK(n10438), 
        .Q(WX9942), .QN(n9501) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n10067), .CLK(n10438), 
        .Q(WX9944), .QN(n9574) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n10066), .CLK(n10439), 
        .Q(WX9946), .QN(n9575) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n10066), .CLK(n10439), 
        .Q(WX9948) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n10066), .CLK(n10439), 
        .Q(WX9950), .QN(n9518) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n10046), .CLK(n10459), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n10046), .CLK(
        n10459), .Q(test_so87), .QN(n9864) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_2_3), .QN(DFF_1507_n1) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_10), .QN(DFF_1514_n1) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n10045), .CLK(
        n10460), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n10044), .CLK(
        n10461), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n10044), .CLK(
        n10461), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n10063), .CLK(
        n10442), .Q(test_so88), .QN(n9863) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n10063), .CLK(
        n10442), .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n10063), .CLK(
        n10442), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n10063), .CLK(
        n10442), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n10063), .CLK(
        n10442), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n10063), .CLK(
        n10442), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n10062), .CLK(
        n10443), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n10062), .CLK(
        n10443), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n10062), .CLK(
        n10443), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n10062), .CLK(
        n10443), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n10062), .CLK(
        n10443), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n10062), .CLK(
        n10443), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n10062), .CLK(
        n10443), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n2013), .SI(CRC_OUT_2_31), .SE(n10062), .CLK(
        n10443), .Q(WX10829) );
  SDFFX1 DFF_1537_Q_reg ( .D(n2015), .SI(WX10829), .SE(n10059), .CLK(n10446), 
        .Q(n8295), .QN(n9900) );
  SDFFX1 DFF_1538_Q_reg ( .D(n2017), .SI(n8295), .SE(n10059), .CLK(n10446), 
        .Q(n8294), .QN(n9899) );
  SDFFX1 DFF_1539_Q_reg ( .D(n2019), .SI(n8294), .SE(n10059), .CLK(n10446), 
        .Q(n8293), .QN(n9898) );
  SDFFX1 DFF_1540_Q_reg ( .D(n2021), .SI(n8293), .SE(n10060), .CLK(n10445), 
        .Q(test_so89), .QN(n9902) );
  SDFFX1 DFF_1541_Q_reg ( .D(n2023), .SI(test_si90), .SE(n10060), .CLK(n10445), 
        .Q(n8290), .QN(n9897) );
  SDFFX1 DFF_1542_Q_reg ( .D(n2025), .SI(n8290), .SE(n10060), .CLK(n10445), 
        .Q(n8289), .QN(n9896) );
  SDFFX1 DFF_1543_Q_reg ( .D(n2027), .SI(n8289), .SE(n10060), .CLK(n10445), 
        .Q(n8288), .QN(n9895) );
  SDFFX1 DFF_1544_Q_reg ( .D(n2029), .SI(n8288), .SE(n10060), .CLK(n10445), 
        .Q(n8287), .QN(n9894) );
  SDFFX1 DFF_1545_Q_reg ( .D(n2031), .SI(n8287), .SE(n10060), .CLK(n10445), 
        .Q(n8286), .QN(n9893) );
  SDFFX1 DFF_1546_Q_reg ( .D(n2033), .SI(n8286), .SE(n10060), .CLK(n10445), 
        .Q(n8285), .QN(n9892) );
  SDFFX1 DFF_1547_Q_reg ( .D(n2035), .SI(n8285), .SE(n10060), .CLK(n10445), 
        .Q(n8284), .QN(n9891) );
  SDFFX1 DFF_1548_Q_reg ( .D(n2037), .SI(n8284), .SE(n10060), .CLK(n10445), 
        .Q(n8283), .QN(n9890) );
  SDFFX1 DFF_1549_Q_reg ( .D(n2039), .SI(n8283), .SE(n10060), .CLK(n10445), 
        .Q(n8282), .QN(n9889) );
  SDFFX1 DFF_1550_Q_reg ( .D(n2041), .SI(n8282), .SE(n10060), .CLK(n10445), 
        .Q(n8281), .QN(n9888) );
  SDFFX1 DFF_1551_Q_reg ( .D(n2043), .SI(n8281), .SE(n10060), .CLK(n10445), 
        .Q(n8280), .QN(n9887) );
  SDFFX1 DFF_1552_Q_reg ( .D(n2045), .SI(n8280), .SE(n10061), .CLK(n10444), 
        .Q(n8279), .QN(n9886) );
  SDFFX1 DFF_1553_Q_reg ( .D(n2047), .SI(n8279), .SE(n10061), .CLK(n10444), 
        .Q(n8278), .QN(n9885) );
  SDFFX1 DFF_1554_Q_reg ( .D(n2049), .SI(n8278), .SE(n10061), .CLK(n10444), 
        .Q(n8277), .QN(n9884) );
  SDFFX1 DFF_1555_Q_reg ( .D(n2051), .SI(n8277), .SE(n10061), .CLK(n10444), 
        .Q(n8276), .QN(n9883) );
  SDFFX1 DFF_1556_Q_reg ( .D(n2053), .SI(n8276), .SE(n10061), .CLK(n10444), 
        .Q(n8275), .QN(n9882) );
  SDFFX1 DFF_1557_Q_reg ( .D(n2055), .SI(n8275), .SE(n10061), .CLK(n10444), 
        .Q(test_so90), .QN(n9901) );
  SDFFX1 DFF_1558_Q_reg ( .D(n2057), .SI(test_si91), .SE(n10061), .CLK(n10444), 
        .Q(n8272), .QN(n9881) );
  SDFFX1 DFF_1559_Q_reg ( .D(n2059), .SI(n8272), .SE(n10061), .CLK(n10444), 
        .Q(n8271), .QN(n9880) );
  SDFFX1 DFF_1560_Q_reg ( .D(n2061), .SI(n8271), .SE(n10061), .CLK(n10444), 
        .Q(n8270), .QN(n9879) );
  SDFFX1 DFF_1561_Q_reg ( .D(n2063), .SI(n8270), .SE(n10061), .CLK(n10444), 
        .Q(n8269), .QN(n9878) );
  SDFFX1 DFF_1562_Q_reg ( .D(n2065), .SI(n8269), .SE(n10061), .CLK(n10444), 
        .Q(n8268), .QN(n9877) );
  SDFFX1 DFF_1563_Q_reg ( .D(n2067), .SI(n8268), .SE(n10061), .CLK(n10444), 
        .Q(n8267), .QN(n9876) );
  SDFFX1 DFF_1564_Q_reg ( .D(n2069), .SI(n8267), .SE(n10062), .CLK(n10443), 
        .Q(n8266), .QN(n9875) );
  SDFFX1 DFF_1565_Q_reg ( .D(n2071), .SI(n8266), .SE(n10062), .CLK(n10443), 
        .Q(n8265), .QN(n9874) );
  SDFFX1 DFF_1566_Q_reg ( .D(n2073), .SI(n8265), .SE(n10062), .CLK(n10443), 
        .Q(n8264), .QN(n9873) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n10062), .CLK(n10443), 
        .Q(n8263), .QN(n9872) );
  SDFFX1 DFF_1568_Q_reg ( .D(n2010), .SI(n8263), .SE(n10059), .CLK(n10446), 
        .Q(n8262), .QN(n18458) );
  SDFFX1 DFF_1569_Q_reg ( .D(n2012), .SI(n8262), .SE(n10059), .CLK(n10446), 
        .Q(n8261), .QN(n18459) );
  SDFFX1 DFF_1570_Q_reg ( .D(n2014), .SI(n8261), .SE(n10059), .CLK(n10446), 
        .Q(n8260), .QN(n18460) );
  SDFFX1 DFF_1571_Q_reg ( .D(n2016), .SI(n8260), .SE(n10059), .CLK(n10446), 
        .Q(n8259), .QN(n18461) );
  SDFFX1 DFF_1572_Q_reg ( .D(n2018), .SI(n8259), .SE(n10059), .CLK(n10446), 
        .Q(n8258), .QN(n18462) );
  SDFFX1 DFF_1573_Q_reg ( .D(n2020), .SI(n8258), .SE(n10058), .CLK(n10447), 
        .Q(n8257), .QN(n18463) );
  SDFFX1 DFF_1574_Q_reg ( .D(n2022), .SI(n8257), .SE(n10058), .CLK(n10447), 
        .Q(test_so91), .QN(n9846) );
  SDFFX1 DFF_1575_Q_reg ( .D(n2024), .SI(test_si92), .SE(n10058), .CLK(n10447), 
        .Q(n8254), .QN(n18464) );
  SDFFX1 DFF_1576_Q_reg ( .D(n2026), .SI(n8254), .SE(n10058), .CLK(n10447), 
        .Q(n8253), .QN(n18465) );
  SDFFX1 DFF_1577_Q_reg ( .D(n2028), .SI(n8253), .SE(n10058), .CLK(n10447), 
        .Q(n8252), .QN(n18466) );
  SDFFX1 DFF_1578_Q_reg ( .D(n2030), .SI(n8252), .SE(n10057), .CLK(n10448), 
        .Q(n8251), .QN(n18467) );
  SDFFX1 DFF_1579_Q_reg ( .D(n2032), .SI(n8251), .SE(n10057), .CLK(n10448), 
        .Q(n8250), .QN(n18468) );
  SDFFX1 DFF_1580_Q_reg ( .D(n2034), .SI(n8250), .SE(n10057), .CLK(n10448), 
        .Q(n8249), .QN(n18469) );
  SDFFX1 DFF_1581_Q_reg ( .D(n2036), .SI(n8249), .SE(n10057), .CLK(n10448), 
        .Q(n8248), .QN(n18470) );
  SDFFX1 DFF_1582_Q_reg ( .D(n2038), .SI(n8248), .SE(n10056), .CLK(n10449), 
        .Q(n8247), .QN(n18471) );
  SDFFX1 DFF_1583_Q_reg ( .D(n2040), .SI(n8247), .SE(n10056), .CLK(n10449), 
        .Q(n8246), .QN(n18472) );
  SDFFX1 DFF_1584_Q_reg ( .D(n2042), .SI(n8246), .SE(n10055), .CLK(n10450), 
        .Q(WX11021), .QN(n9273) );
  SDFFX1 DFF_1585_Q_reg ( .D(n2044), .SI(WX11021), .SE(n10055), .CLK(n10450), 
        .Q(WX11023), .QN(n9271) );
  SDFFX1 DFF_1586_Q_reg ( .D(n2046), .SI(WX11023), .SE(n10055), .CLK(n10450), 
        .Q(WX11025), .QN(n9269) );
  SDFFX1 DFF_1587_Q_reg ( .D(n2048), .SI(WX11025), .SE(n10055), .CLK(n10450), 
        .Q(WX11027), .QN(n9267) );
  SDFFX1 DFF_1588_Q_reg ( .D(n2050), .SI(WX11027), .SE(n10054), .CLK(n10451), 
        .Q(WX11029), .QN(n9265) );
  SDFFX1 DFF_1589_Q_reg ( .D(n2052), .SI(WX11029), .SE(n10054), .CLK(n10451), 
        .Q(WX11031), .QN(n9263) );
  SDFFX1 DFF_1590_Q_reg ( .D(n2054), .SI(WX11031), .SE(n10054), .CLK(n10451), 
        .Q(WX11033), .QN(n9261) );
  SDFFX1 DFF_1591_Q_reg ( .D(n2056), .SI(WX11033), .SE(n10053), .CLK(n10452), 
        .Q(test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(n2058), .SI(test_si93), .SE(n10053), .CLK(n10452), 
        .Q(WX11037), .QN(n9258) );
  SDFFX1 DFF_1593_Q_reg ( .D(n2060), .SI(WX11037), .SE(n10053), .CLK(n10452), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(n2062), .SI(WX11039), .SE(n10052), .CLK(n10453), 
        .Q(WX11041), .QN(n9254) );
  SDFFX1 DFF_1595_Q_reg ( .D(n2064), .SI(WX11041), .SE(n10052), .CLK(n10453), 
        .Q(WX11043), .QN(n9253) );
  SDFFX1 DFF_1596_Q_reg ( .D(n2066), .SI(WX11043), .SE(n10052), .CLK(n10453), 
        .Q(WX11045), .QN(n9251) );
  SDFFX1 DFF_1597_Q_reg ( .D(n2068), .SI(WX11045), .SE(n10051), .CLK(n10454), 
        .Q(WX11047), .QN(n9249) );
  SDFFX1 DFF_1598_Q_reg ( .D(n2070), .SI(WX11047), .SE(n10051), .CLK(n10454), 
        .Q(WX11049), .QN(n9247) );
  SDFFX1 DFF_1599_Q_reg ( .D(n2072), .SI(WX11049), .SE(n10051), .CLK(n10454), 
        .Q(WX11051), .QN(n9245) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n10059), .CLK(n10446), 
        .Q(WX11053), .QN(n9003) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n10059), .CLK(n10446), 
        .Q(WX11055), .QN(n9045) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n10059), .CLK(n10446), 
        .Q(WX11057), .QN(n9043) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n10059), .CLK(n10446), 
        .Q(WX11059), .QN(n9041) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n10058), .CLK(n10447), 
        .Q(WX11061), .QN(n9039) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n10058), .CLK(n10447), 
        .Q(WX11063), .QN(n9037) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n10058), .CLK(n10447), 
        .Q(WX11065), .QN(n9035) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n10058), .CLK(n10447), 
        .Q(WX11067), .QN(n9033) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n10058), .CLK(n10447), 
        .Q(test_so93), .QN(n9866) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n10057), .CLK(
        n10448), .Q(WX11071), .QN(n9030) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n10057), .CLK(n10448), 
        .Q(WX11073), .QN(n9029) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n10057), .CLK(n10448), 
        .Q(WX11075), .QN(n9027) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n10057), .CLK(n10448), 
        .Q(WX11077), .QN(n9025) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n10057), .CLK(n10448), 
        .Q(WX11079), .QN(n9023) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n10056), .CLK(n10449), 
        .Q(WX11081), .QN(n9021) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n10056), .CLK(n10449), 
        .Q(WX11083), .QN(n9019) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n10056), .CLK(n10449), 
        .Q(WX11085) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n10055), .CLK(n10450), 
        .Q(WX11087) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n10055), .CLK(n10450), 
        .Q(WX11089) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n10055), .CLK(n10450), 
        .Q(WX11091) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n10054), .CLK(n10451), 
        .Q(WX11093) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n10054), .CLK(n10451), 
        .Q(WX11095) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n10054), .CLK(n10451), 
        .Q(WX11097) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n10053), .CLK(n10452), 
        .Q(WX11099) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n10053), .CLK(n10452), 
        .Q(WX11101) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n10053), .CLK(n10452), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n10052), .CLK(
        n10453), .Q(WX11105) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n10052), .CLK(n10453), 
        .Q(WX11107) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n10052), .CLK(n10453), 
        .Q(WX11109) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n10051), .CLK(n10454), 
        .Q(WX11111) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n10051), .CLK(n10454), 
        .Q(WX11113) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n10051), .CLK(n10454), 
        .Q(WX11115) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n10050), .CLK(n10455), 
        .Q(WX11117), .QN(n9004) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n10050), .CLK(n10455), 
        .Q(WX11119), .QN(n9046) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n10050), .CLK(n10455), 
        .Q(WX11121), .QN(n9044) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n10050), .CLK(n10455), 
        .Q(WX11123), .QN(n9042) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n10050), .CLK(n10455), 
        .Q(WX11125), .QN(n9040) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n10049), .CLK(n10456), 
        .Q(WX11127), .QN(n9038) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n10049), .CLK(n10456), 
        .Q(WX11129), .QN(n9036) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n10049), .CLK(n10456), 
        .Q(WX11131), .QN(n9034) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n10058), .CLK(n10447), 
        .Q(WX11133), .QN(n9032) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n10058), .CLK(n10447), 
        .Q(WX11135), .QN(n9031) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n10057), .CLK(n10448), 
        .Q(test_so95), .QN(n9865) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n10057), .CLK(
        n10448), .Q(WX11139), .QN(n9028) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n10057), .CLK(n10448), 
        .Q(WX11141), .QN(n9026) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n10056), .CLK(n10449), 
        .Q(WX11143), .QN(n9024) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n10056), .CLK(n10449), 
        .Q(WX11145), .QN(n9022) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n10056), .CLK(n10449), 
        .Q(WX11147), .QN(n9020) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n10056), .CLK(n10449), 
        .Q(WX11149), .QN(n9274) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n10055), .CLK(n10450), 
        .Q(WX11151), .QN(n9272) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n10055), .CLK(n10450), 
        .Q(WX11153), .QN(n9270) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n10054), .CLK(n10451), 
        .Q(WX11155), .QN(n9268) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155), .SE(n10054), .CLK(n10451), 
        .Q(WX11157), .QN(n9266) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(n10054), .CLK(n10451), 
        .Q(WX11159), .QN(n9264) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(n10053), .CLK(n10452), 
        .Q(WX11161), .QN(n9262) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(n10053), .CLK(n10452), 
        .Q(WX11163), .QN(n9260) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(n10053), .CLK(n10452), 
        .Q(WX11165), .QN(n9259) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(n10052), .CLK(n10453), 
        .Q(WX11167), .QN(n9257) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(n10052), .CLK(n10453), 
        .Q(WX11169), .QN(n9255) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(n10052), .CLK(n10453), 
        .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n10051), .CLK(
        n10454), .Q(WX11173), .QN(n9252) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n10051), .CLK(n10454), 
        .Q(WX11175), .QN(n9250) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n10051), .CLK(n10454), 
        .Q(WX11177), .QN(n9248) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n10050), .CLK(n10455), 
        .Q(WX11179), .QN(n9246) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n10050), .CLK(n10455), 
        .Q(WX11181), .QN(n9525) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n10050), .CLK(n10455), 
        .Q(WX11183), .QN(n9526) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n10050), .CLK(n10455), 
        .Q(WX11185), .QN(n9527) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n10050), .CLK(n10455), 
        .Q(WX11187), .QN(n9528) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n10050), .CLK(n10455), 
        .Q(WX11189), .QN(n9529) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n10049), .CLK(n10456), 
        .Q(WX11191), .QN(n9530) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n10049), .CLK(n10456), 
        .Q(WX11193), .QN(n9531) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n10049), .CLK(n10456), 
        .Q(WX11195), .QN(n9532) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n10049), .CLK(n10456), 
        .Q(WX11197), .QN(n9533) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n10049), .CLK(n10456), 
        .Q(WX11199), .QN(n9534) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n10049), .CLK(n10456), 
        .Q(WX11201), .QN(n9535) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n10049), .CLK(n10456), 
        .Q(WX11203), .QN(n9536) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n10049), .CLK(n10456), 
        .Q(test_so97), .QN(n9839) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n10056), .CLK(
        n10449), .Q(WX11207), .QN(n9537) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n10056), .CLK(n10449), 
        .Q(WX11209), .QN(n9538) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n10056), .CLK(n10449), 
        .Q(WX11211), .QN(n9496) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n10055), .CLK(n10450), 
        .Q(WX11213) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n10055), .CLK(n10450), 
        .Q(WX11215), .QN(n9540) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n10055), .CLK(n10450), 
        .Q(WX11217), .QN(n9541) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n10054), .CLK(n10451), 
        .Q(WX11219), .QN(n9542) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n10054), .CLK(n10451), 
        .Q(WX11221), .QN(n9497) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n10054), .CLK(n10451), 
        .Q(WX11223), .QN(n9543) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n10053), .CLK(n10452), 
        .Q(WX11225), .QN(n9544) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n10053), .CLK(n10452), 
        .Q(WX11227), .QN(n9545) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n10053), .CLK(n10452), 
        .Q(WX11229), .QN(n9546) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n10052), .CLK(n10453), 
        .Q(WX11231), .QN(n9547) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n10052), .CLK(n10453), 
        .Q(WX11233), .QN(n9548) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n10052), .CLK(n10453), 
        .Q(WX11235), .QN(n9498) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n10051), .CLK(n10454), 
        .Q(WX11237), .QN(n9549) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n10051), .CLK(n10454), 
        .Q(test_so98), .QN(n9847) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n10051), .CLK(
        n10454), .Q(WX11241), .QN(n9550) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n10050), .CLK(n10455), 
        .Q(WX11243), .QN(n9517) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n10048), .CLK(n10457), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_3) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_10) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n10047), .CLK(
        n10458), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_15) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n10047), .CLK(
        n10458), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n10046), .CLK(
        n10459), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n10049), .CLK(
        n10456), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n10048), .CLK(
        n10457), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n10048), .CLK(
        n10457), .Q(test_so100), .QN(n9838) );
  NOR2X0 Trojan1 ( .IN1(WX3442), .IN2(WX5974), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(WX806), .IN2(WX782), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(WX11632), .IN2(n584), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(WX5964), .IN2(WX3324), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(WX8634), .IN2(WX3330), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n596), .IN2(n588), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(WX862), .IN2(WX7227), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(WX11616), .IN2(n2047), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(n10175), 
        .Q(Tj_Trigger) );
  NAND3X4 TrojanPayload1 ( .IN1(WX547), .IN2(Tj_Trigger), .IN3(Stage4), .QN(
        Stage1_1) );
  INVX8 TrojanPayload2 ( .INP(Stage1_1), .ZN(Stage1_2) );
  INVX8 TrojanPayload3 ( .INP(Stage1_2), .ZN(Stage1_3) );
  INVX8 TrojanPayload4 ( .INP(Stage1_3), .ZN(Stage1_4) );
  INVX8 TrojanPayload5 ( .INP(Stage1_4), .ZN(Stage1) );
  MUX21X2 TrojanPayload6 ( .IN1(WX544), .IN2(Stage1), .S(1'b0), .Q(Stage2_i)
         );
  INVX8 TrojanPayload7 ( .INP(Stage2_i), .ZN(Stage2_7) );
  INVX8 TrojanPayload8 ( .INP(Stage2_7), .ZN(Stage2_8) );
  INVX8 TrojanPayload9 ( .INP(Stage2_8), .ZN(Stage2_9) );
  INVX8 TrojanPayload10 ( .INP(Stage2_9), .ZN(Stage2_10) );
  INVX8 TrojanPayload11 ( .INP(Stage2_10), .ZN(Stage2) );
  MUX21X2 TrojanPayload12 ( .IN1(n135), .IN2(Stage2), .S(1'b0), .Q(Stage3_i)
         );
  INVX8 TrojanPayload13 ( .INP(Stage3_i), .ZN(Stage3_12) );
  INVX8 TrojanPayload14 ( .INP(Stage3_12), .ZN(Stage3_13) );
  INVX8 TrojanPayload15 ( .INP(Stage3_13), .ZN(Stage3_14) );
  INVX8 TrojanPayload16 ( .INP(Stage3_14), .ZN(Stage3_15) );
  INVX8 TrojanPayload17 ( .INP(Stage3_15) );
  MUX21X2 TrojanPayload18 ( .IN1(n3467), .IN2(1'b0), .S(1'b0), .Q(Stage4_i) );
  INVX8 TrojanPayload19 ( .INP(Stage4_i), .ZN(Stage4_17) );
  INVX8 TrojanPayload20 ( .INP(Stage4_17), .ZN(Stage4_18) );
  INVX8 TrojanPayload21 ( .INP(Stage4_18), .ZN(Stage4_19) );
  INVX8 TrojanPayload22 ( .INP(Stage4_19), .ZN(Stage4_20) );
  INVX8 TrojanPayload23 ( .INP(Stage4_20), .ZN(Stage4_21) );
  INVX8 TrojanPayload24 ( .INP(Stage4_21), .ZN(Stage4) );
  NBUFFX2 U9948 ( .INP(n9957), .Z(n9975) );
  NBUFFX2 U9949 ( .INP(n9980), .Z(n9998) );
  NBUFFX2 U9950 ( .INP(n9980), .Z(n9997) );
  NBUFFX2 U9951 ( .INP(n9980), .Z(n9996) );
  NBUFFX2 U9952 ( .INP(n9979), .Z(n9995) );
  NBUFFX2 U9953 ( .INP(n9979), .Z(n9994) );
  NBUFFX2 U9954 ( .INP(n9979), .Z(n9993) );
  NBUFFX2 U9955 ( .INP(n9979), .Z(n9992) );
  NBUFFX2 U9956 ( .INP(n9979), .Z(n9991) );
  NBUFFX2 U9957 ( .INP(n9978), .Z(n9990) );
  NBUFFX2 U9958 ( .INP(n9978), .Z(n9989) );
  NBUFFX2 U9959 ( .INP(n9978), .Z(n9988) );
  NBUFFX2 U9960 ( .INP(n9978), .Z(n9987) );
  NBUFFX2 U9961 ( .INP(n9978), .Z(n9986) );
  NBUFFX2 U9962 ( .INP(n9977), .Z(n9985) );
  NBUFFX2 U9963 ( .INP(n9977), .Z(n9984) );
  NBUFFX2 U9964 ( .INP(n9977), .Z(n9983) );
  NBUFFX2 U9965 ( .INP(n9977), .Z(n9982) );
  NBUFFX2 U9966 ( .INP(n9977), .Z(n9981) );
  NBUFFX2 U9967 ( .INP(n9957), .Z(n9974) );
  NBUFFX2 U9968 ( .INP(n9957), .Z(n9973) );
  NBUFFX2 U9969 ( .INP(n9955), .Z(n9966) );
  NBUFFX2 U9970 ( .INP(n9955), .Z(n9965) );
  NBUFFX2 U9971 ( .INP(n9955), .Z(n9964) );
  NBUFFX2 U9972 ( .INP(n9955), .Z(n9963) );
  NBUFFX2 U9973 ( .INP(n9954), .Z(n9961) );
  NBUFFX2 U9974 ( .INP(n9954), .Z(n9960) );
  NBUFFX2 U9975 ( .INP(n9954), .Z(n9962) );
  NBUFFX2 U9976 ( .INP(n9956), .Z(n9972) );
  NBUFFX2 U9977 ( .INP(n9956), .Z(n9970) );
  NBUFFX2 U9978 ( .INP(n9956), .Z(n9969) );
  NBUFFX2 U9979 ( .INP(n9956), .Z(n9968) );
  NBUFFX2 U9980 ( .INP(n9955), .Z(n9967) );
  NBUFFX2 U9981 ( .INP(n9956), .Z(n9971) );
  NBUFFX2 U9982 ( .INP(n9954), .Z(n9958) );
  NBUFFX2 U9983 ( .INP(n9954), .Z(n9959) );
  NBUFFX2 U9984 ( .INP(n9957), .Z(n9976) );
  NBUFFX2 U9985 ( .INP(n10505), .Z(n10336) );
  NBUFFX2 U9986 ( .INP(n10505), .Z(n10334) );
  NBUFFX2 U9987 ( .INP(n10505), .Z(n10335) );
  NBUFFX2 U9988 ( .INP(n10505), .Z(n10333) );
  NBUFFX2 U9989 ( .INP(n10480), .Z(n10458) );
  NBUFFX2 U9990 ( .INP(n10480), .Z(n10457) );
  NBUFFX2 U9991 ( .INP(n10481), .Z(n10456) );
  NBUFFX2 U9992 ( .INP(n10481), .Z(n10455) );
  NBUFFX2 U9993 ( .INP(n10481), .Z(n10454) );
  NBUFFX2 U9994 ( .INP(n10481), .Z(n10453) );
  NBUFFX2 U9995 ( .INP(n10481), .Z(n10452) );
  NBUFFX2 U9996 ( .INP(n10482), .Z(n10451) );
  NBUFFX2 U9997 ( .INP(n10482), .Z(n10450) );
  NBUFFX2 U9998 ( .INP(n10482), .Z(n10449) );
  NBUFFX2 U9999 ( .INP(n10482), .Z(n10448) );
  NBUFFX2 U10000 ( .INP(n10482), .Z(n10447) );
  NBUFFX2 U10001 ( .INP(n10483), .Z(n10444) );
  NBUFFX2 U10002 ( .INP(n10483), .Z(n10445) );
  NBUFFX2 U10003 ( .INP(n10483), .Z(n10446) );
  NBUFFX2 U10004 ( .INP(n10483), .Z(n10443) );
  NBUFFX2 U10005 ( .INP(n10480), .Z(n10460) );
  NBUFFX2 U10006 ( .INP(n10480), .Z(n10459) );
  NBUFFX2 U10007 ( .INP(n10483), .Z(n10442) );
  NBUFFX2 U10008 ( .INP(n10484), .Z(n10441) );
  NBUFFX2 U10009 ( .INP(n10484), .Z(n10440) );
  NBUFFX2 U10010 ( .INP(n10484), .Z(n10439) );
  NBUFFX2 U10011 ( .INP(n10484), .Z(n10438) );
  NBUFFX2 U10012 ( .INP(n10484), .Z(n10437) );
  NBUFFX2 U10013 ( .INP(n10485), .Z(n10436) );
  NBUFFX2 U10014 ( .INP(n10485), .Z(n10435) );
  NBUFFX2 U10015 ( .INP(n10485), .Z(n10434) );
  NBUFFX2 U10016 ( .INP(n10485), .Z(n10433) );
  NBUFFX2 U10017 ( .INP(n10485), .Z(n10432) );
  NBUFFX2 U10018 ( .INP(n10486), .Z(n10430) );
  NBUFFX2 U10019 ( .INP(n10486), .Z(n10431) );
  NBUFFX2 U10020 ( .INP(n10479), .Z(n10462) );
  NBUFFX2 U10021 ( .INP(n10480), .Z(n10461) );
  NBUFFX2 U10022 ( .INP(n10486), .Z(n10429) );
  NBUFFX2 U10023 ( .INP(n10486), .Z(n10428) );
  NBUFFX2 U10024 ( .INP(n10486), .Z(n10427) );
  NBUFFX2 U10025 ( .INP(n10487), .Z(n10426) );
  NBUFFX2 U10026 ( .INP(n10487), .Z(n10425) );
  NBUFFX2 U10027 ( .INP(n10487), .Z(n10424) );
  NBUFFX2 U10028 ( .INP(n10487), .Z(n10423) );
  NBUFFX2 U10029 ( .INP(n10487), .Z(n10422) );
  NBUFFX2 U10030 ( .INP(n10488), .Z(n10421) );
  NBUFFX2 U10031 ( .INP(n10488), .Z(n10420) );
  NBUFFX2 U10032 ( .INP(n10488), .Z(n10419) );
  NBUFFX2 U10033 ( .INP(n10489), .Z(n10416) );
  NBUFFX2 U10034 ( .INP(n10488), .Z(n10417) );
  NBUFFX2 U10035 ( .INP(n10488), .Z(n10418) );
  NBUFFX2 U10036 ( .INP(n10479), .Z(n10465) );
  NBUFFX2 U10037 ( .INP(n10479), .Z(n10464) );
  NBUFFX2 U10038 ( .INP(n10479), .Z(n10463) );
  NBUFFX2 U10039 ( .INP(n10489), .Z(n10415) );
  NBUFFX2 U10040 ( .INP(n10489), .Z(n10414) );
  NBUFFX2 U10041 ( .INP(n10489), .Z(n10413) );
  NBUFFX2 U10042 ( .INP(n10489), .Z(n10412) );
  NBUFFX2 U10043 ( .INP(n10490), .Z(n10411) );
  NBUFFX2 U10044 ( .INP(n10490), .Z(n10410) );
  NBUFFX2 U10045 ( .INP(n10490), .Z(n10409) );
  NBUFFX2 U10046 ( .INP(n10490), .Z(n10408) );
  NBUFFX2 U10047 ( .INP(n10490), .Z(n10407) );
  NBUFFX2 U10048 ( .INP(n10491), .Z(n10406) );
  NBUFFX2 U10049 ( .INP(n10491), .Z(n10405) );
  NBUFFX2 U10050 ( .INP(n10491), .Z(n10403) );
  NBUFFX2 U10051 ( .INP(n10491), .Z(n10404) );
  NBUFFX2 U10052 ( .INP(n10491), .Z(n10402) );
  NBUFFX2 U10053 ( .INP(n10479), .Z(n10466) );
  NBUFFX2 U10054 ( .INP(n10492), .Z(n10401) );
  NBUFFX2 U10055 ( .INP(n10492), .Z(n10400) );
  NBUFFX2 U10056 ( .INP(n10492), .Z(n10399) );
  NBUFFX2 U10057 ( .INP(n10492), .Z(n10398) );
  NBUFFX2 U10058 ( .INP(n10492), .Z(n10397) );
  NBUFFX2 U10059 ( .INP(n10493), .Z(n10396) );
  NBUFFX2 U10060 ( .INP(n10493), .Z(n10395) );
  NBUFFX2 U10061 ( .INP(n10493), .Z(n10394) );
  NBUFFX2 U10062 ( .INP(n10493), .Z(n10393) );
  NBUFFX2 U10063 ( .INP(n10493), .Z(n10392) );
  NBUFFX2 U10064 ( .INP(n10494), .Z(n10391) );
  NBUFFX2 U10065 ( .INP(n10494), .Z(n10388) );
  NBUFFX2 U10066 ( .INP(n10494), .Z(n10389) );
  NBUFFX2 U10067 ( .INP(n10494), .Z(n10390) );
  NBUFFX2 U10068 ( .INP(n10478), .Z(n10469) );
  NBUFFX2 U10069 ( .INP(n10478), .Z(n10468) );
  NBUFFX2 U10070 ( .INP(n10478), .Z(n10467) );
  NBUFFX2 U10071 ( .INP(n10494), .Z(n10387) );
  NBUFFX2 U10072 ( .INP(n10495), .Z(n10386) );
  NBUFFX2 U10073 ( .INP(n10495), .Z(n10385) );
  NBUFFX2 U10074 ( .INP(n10495), .Z(n10384) );
  NBUFFX2 U10075 ( .INP(n10495), .Z(n10383) );
  NBUFFX2 U10076 ( .INP(n10495), .Z(n10382) );
  NBUFFX2 U10077 ( .INP(n10496), .Z(n10381) );
  NBUFFX2 U10078 ( .INP(n10496), .Z(n10380) );
  NBUFFX2 U10079 ( .INP(n10496), .Z(n10379) );
  NBUFFX2 U10080 ( .INP(n10496), .Z(n10378) );
  NBUFFX2 U10081 ( .INP(n10497), .Z(n10375) );
  NBUFFX2 U10082 ( .INP(n10497), .Z(n10376) );
  NBUFFX2 U10083 ( .INP(n10496), .Z(n10377) );
  NBUFFX2 U10084 ( .INP(n10497), .Z(n10374) );
  NBUFFX2 U10085 ( .INP(n10478), .Z(n10471) );
  NBUFFX2 U10086 ( .INP(n10478), .Z(n10470) );
  NBUFFX2 U10087 ( .INP(n10497), .Z(n10373) );
  NBUFFX2 U10088 ( .INP(n10497), .Z(n10372) );
  NBUFFX2 U10089 ( .INP(n10498), .Z(n10371) );
  NBUFFX2 U10090 ( .INP(n10498), .Z(n10370) );
  NBUFFX2 U10091 ( .INP(n10498), .Z(n10369) );
  NBUFFX2 U10092 ( .INP(n10498), .Z(n10368) );
  NBUFFX2 U10093 ( .INP(n10498), .Z(n10367) );
  NBUFFX2 U10094 ( .INP(n10499), .Z(n10366) );
  NBUFFX2 U10095 ( .INP(n10499), .Z(n10365) );
  NBUFFX2 U10096 ( .INP(n10499), .Z(n10364) );
  NBUFFX2 U10097 ( .INP(n10500), .Z(n10361) );
  NBUFFX2 U10098 ( .INP(n10499), .Z(n10362) );
  NBUFFX2 U10099 ( .INP(n10499), .Z(n10363) );
  NBUFFX2 U10100 ( .INP(n10477), .Z(n10474) );
  NBUFFX2 U10101 ( .INP(n10477), .Z(n10473) );
  NBUFFX2 U10102 ( .INP(n10477), .Z(n10472) );
  NBUFFX2 U10103 ( .INP(n10500), .Z(n10360) );
  NBUFFX2 U10104 ( .INP(n10500), .Z(n10359) );
  NBUFFX2 U10105 ( .INP(n10500), .Z(n10358) );
  NBUFFX2 U10106 ( .INP(n10500), .Z(n10357) );
  NBUFFX2 U10107 ( .INP(n10501), .Z(n10356) );
  NBUFFX2 U10108 ( .INP(n10501), .Z(n10355) );
  NBUFFX2 U10109 ( .INP(n10501), .Z(n10354) );
  NBUFFX2 U10110 ( .INP(n10501), .Z(n10353) );
  NBUFFX2 U10111 ( .INP(n10501), .Z(n10352) );
  NBUFFX2 U10112 ( .INP(n10502), .Z(n10351) );
  NBUFFX2 U10113 ( .INP(n10502), .Z(n10350) );
  NBUFFX2 U10114 ( .INP(n10502), .Z(n10348) );
  NBUFFX2 U10115 ( .INP(n10502), .Z(n10349) );
  NBUFFX2 U10116 ( .INP(n10502), .Z(n10347) );
  NBUFFX2 U10117 ( .INP(n10477), .Z(n10476) );
  NBUFFX2 U10118 ( .INP(n10477), .Z(n10475) );
  NBUFFX2 U10119 ( .INP(n10503), .Z(n10346) );
  NBUFFX2 U10120 ( .INP(n10503), .Z(n10345) );
  NBUFFX2 U10121 ( .INP(n10503), .Z(n10344) );
  NBUFFX2 U10122 ( .INP(n10503), .Z(n10343) );
  NBUFFX2 U10123 ( .INP(n10503), .Z(n10342) );
  NBUFFX2 U10124 ( .INP(n10504), .Z(n10341) );
  NBUFFX2 U10125 ( .INP(n10504), .Z(n10340) );
  NBUFFX2 U10126 ( .INP(n10504), .Z(n10339) );
  NBUFFX2 U10127 ( .INP(n10504), .Z(n10338) );
  NBUFFX2 U10128 ( .INP(n10504), .Z(n10337) );
  NBUFFX2 U10129 ( .INP(n9906), .Z(n9924) );
  NBUFFX2 U10130 ( .INP(n9906), .Z(n9925) );
  NBUFFX2 U10131 ( .INP(n9906), .Z(n9922) );
  NBUFFX2 U10132 ( .INP(n9906), .Z(n9923) );
  NBUFFX2 U10133 ( .INP(n9905), .Z(n9921) );
  NBUFFX2 U10134 ( .INP(n9903), .Z(n9908) );
  NBUFFX2 U10135 ( .INP(n9903), .Z(n9909) );
  NBUFFX2 U10136 ( .INP(n9903), .Z(n9910) );
  NBUFFX2 U10137 ( .INP(n9903), .Z(n9911) );
  NBUFFX2 U10138 ( .INP(n9904), .Z(n9912) );
  NBUFFX2 U10139 ( .INP(n9904), .Z(n9914) );
  NBUFFX2 U10140 ( .INP(n9905), .Z(n9920) );
  NBUFFX2 U10141 ( .INP(n9905), .Z(n9919) );
  NBUFFX2 U10142 ( .INP(n9905), .Z(n9918) );
  NBUFFX2 U10143 ( .INP(n9905), .Z(n9917) );
  NBUFFX2 U10144 ( .INP(n9904), .Z(n9916) );
  NBUFFX2 U10145 ( .INP(n9904), .Z(n9915) );
  NBUFFX2 U10146 ( .INP(n9903), .Z(n9907) );
  NBUFFX2 U10147 ( .INP(n9904), .Z(n9913) );
  NBUFFX2 U10148 ( .INP(n9906), .Z(n9926) );
  NBUFFX2 U10149 ( .INP(n9999), .Z(n10004) );
  NBUFFX2 U10150 ( .INP(n9999), .Z(n10005) );
  NBUFFX2 U10151 ( .INP(n9999), .Z(n10006) );
  NBUFFX2 U10152 ( .INP(n9999), .Z(n10007) );
  NBUFFX2 U10153 ( .INP(n10000), .Z(n10008) );
  NBUFFX2 U10154 ( .INP(n10000), .Z(n10009) );
  NBUFFX2 U10155 ( .INP(n10000), .Z(n10012) );
  NBUFFX2 U10156 ( .INP(n10000), .Z(n10011) );
  NBUFFX2 U10157 ( .INP(n10000), .Z(n10010) );
  NBUFFX2 U10158 ( .INP(n9999), .Z(n10003) );
  NBUFFX2 U10159 ( .INP(n10001), .Z(n10013) );
  NBUFFX2 U10160 ( .INP(n10002), .Z(n10018) );
  NBUFFX2 U10161 ( .INP(n10002), .Z(n10019) );
  NBUFFX2 U10162 ( .INP(n10002), .Z(n10020) );
  NBUFFX2 U10163 ( .INP(n10001), .Z(n10015) );
  NBUFFX2 U10164 ( .INP(n10001), .Z(n10017) );
  NBUFFX2 U10165 ( .INP(n10001), .Z(n10014) );
  NBUFFX2 U10166 ( .INP(n10001), .Z(n10016) );
  NBUFFX2 U10167 ( .INP(n10002), .Z(n10021) );
  INVX0 U10168 ( .INP(n10026), .ZN(n10176) );
  INVX0 U10169 ( .INP(n10025), .ZN(n10175) );
  INVX0 U10170 ( .INP(n10025), .ZN(n10174) );
  INVX0 U10171 ( .INP(n10024), .ZN(n10173) );
  INVX0 U10172 ( .INP(n10024), .ZN(n10172) );
  INVX0 U10173 ( .INP(n10023), .ZN(n10171) );
  INVX0 U10174 ( .INP(n10023), .ZN(n10170) );
  INVX0 U10175 ( .INP(n10026), .ZN(n10177) );
  INVX0 U10176 ( .INP(n10022), .ZN(n10169) );
  INVX0 U10177 ( .INP(n10022), .ZN(n10168) );
  NBUFFX2 U10178 ( .INP(n10027), .Z(n10025) );
  NBUFFX2 U10179 ( .INP(n10027), .Z(n10024) );
  NBUFFX2 U10180 ( .INP(n10028), .Z(n10023) );
  NBUFFX2 U10181 ( .INP(n10027), .Z(n10026) );
  NBUFFX2 U10182 ( .INP(n10028), .Z(n10022) );
  INVX0 U10183 ( .INP(n10563), .ZN(n9953) );
  NBUFFX2 U10184 ( .INP(n10525), .Z(n9903) );
  NBUFFX2 U10185 ( .INP(n10525), .Z(n9904) );
  NBUFFX2 U10186 ( .INP(n10525), .Z(n9905) );
  NBUFFX2 U10187 ( .INP(n10525), .Z(n9906) );
  INVX0 U10188 ( .INP(n9948), .ZN(n9927) );
  INVX0 U10189 ( .INP(n9948), .ZN(n9928) );
  INVX0 U10190 ( .INP(n9948), .ZN(n9929) );
  INVX0 U10191 ( .INP(n9948), .ZN(n9930) );
  INVX0 U10192 ( .INP(n9948), .ZN(n9931) );
  INVX0 U10193 ( .INP(n9947), .ZN(n9932) );
  INVX0 U10194 ( .INP(n9947), .ZN(n9933) );
  INVX0 U10195 ( .INP(n9947), .ZN(n9934) );
  INVX0 U10196 ( .INP(n9947), .ZN(n9935) );
  INVX0 U10197 ( .INP(n9947), .ZN(n9936) );
  INVX0 U10198 ( .INP(n9947), .ZN(n9937) );
  INVX0 U10199 ( .INP(n9947), .ZN(n9938) );
  INVX0 U10200 ( .INP(n9947), .ZN(n9939) );
  INVX0 U10201 ( .INP(n9946), .ZN(n9940) );
  INVX0 U10202 ( .INP(n9946), .ZN(n9941) );
  INVX0 U10203 ( .INP(n9946), .ZN(n9942) );
  INVX0 U10204 ( .INP(n9946), .ZN(n9943) );
  INVX0 U10205 ( .INP(n9946), .ZN(n9944) );
  INVX0 U10206 ( .INP(n9946), .ZN(n9945) );
  NBUFFX2 U10207 ( .INP(n9953), .Z(n9946) );
  NBUFFX2 U10208 ( .INP(n9953), .Z(n9947) );
  NBUFFX2 U10209 ( .INP(n9953), .Z(n9948) );
  NBUFFX2 U10210 ( .INP(n9953), .Z(n9949) );
  NBUFFX2 U10211 ( .INP(n9953), .Z(n9950) );
  NBUFFX2 U10212 ( .INP(n9953), .Z(n9951) );
  NBUFFX2 U10213 ( .INP(n9953), .Z(n9952) );
  NBUFFX2 U10214 ( .INP(n11344), .Z(n9954) );
  NBUFFX2 U10215 ( .INP(n11344), .Z(n9955) );
  NBUFFX2 U10216 ( .INP(n11344), .Z(n9956) );
  NBUFFX2 U10217 ( .INP(n11344), .Z(n9957) );
  NBUFFX2 U10218 ( .INP(n11345), .Z(n9977) );
  NBUFFX2 U10219 ( .INP(n11345), .Z(n9978) );
  NBUFFX2 U10220 ( .INP(n11345), .Z(n9979) );
  NBUFFX2 U10221 ( .INP(n11345), .Z(n9980) );
  NBUFFX2 U10222 ( .INP(n11655), .Z(n9999) );
  NBUFFX2 U10223 ( .INP(n11655), .Z(n10000) );
  NBUFFX2 U10224 ( .INP(n11655), .Z(n10001) );
  NBUFFX2 U10225 ( .INP(n11655), .Z(n10002) );
  NBUFFX2 U10226 ( .INP(test_se), .Z(n10027) );
  NBUFFX2 U10227 ( .INP(test_se), .Z(n10028) );
  INVX0 U10228 ( .INP(n10176), .ZN(n10029) );
  INVX0 U10229 ( .INP(n10176), .ZN(n10030) );
  INVX0 U10230 ( .INP(n10171), .ZN(n10031) );
  INVX0 U10231 ( .INP(n10173), .ZN(n10032) );
  INVX0 U10232 ( .INP(n10174), .ZN(n10033) );
  INVX0 U10233 ( .INP(n10175), .ZN(n10034) );
  INVX0 U10234 ( .INP(n10174), .ZN(n10035) );
  INVX0 U10235 ( .INP(n10173), .ZN(n10036) );
  INVX0 U10236 ( .INP(n10172), .ZN(n10037) );
  INVX0 U10237 ( .INP(n10176), .ZN(n10038) );
  INVX0 U10238 ( .INP(n10177), .ZN(n10039) );
  INVX0 U10239 ( .INP(n10173), .ZN(n10040) );
  INVX0 U10240 ( .INP(n10177), .ZN(n10041) );
  INVX0 U10241 ( .INP(n10177), .ZN(n10042) );
  INVX0 U10242 ( .INP(n10177), .ZN(n10043) );
  INVX0 U10243 ( .INP(n10177), .ZN(n10044) );
  INVX0 U10244 ( .INP(n10177), .ZN(n10045) );
  INVX0 U10245 ( .INP(n10177), .ZN(n10046) );
  INVX0 U10246 ( .INP(n10176), .ZN(n10047) );
  INVX0 U10247 ( .INP(n10176), .ZN(n10048) );
  INVX0 U10248 ( .INP(n10176), .ZN(n10049) );
  INVX0 U10249 ( .INP(n10176), .ZN(n10050) );
  INVX0 U10250 ( .INP(n10176), .ZN(n10051) );
  INVX0 U10251 ( .INP(n10176), .ZN(n10052) );
  INVX0 U10252 ( .INP(n10175), .ZN(n10053) );
  INVX0 U10253 ( .INP(n10175), .ZN(n10054) );
  INVX0 U10254 ( .INP(n10175), .ZN(n10055) );
  INVX0 U10255 ( .INP(n10175), .ZN(n10056) );
  INVX0 U10256 ( .INP(n10175), .ZN(n10057) );
  INVX0 U10257 ( .INP(n10175), .ZN(n10058) );
  INVX0 U10258 ( .INP(n10174), .ZN(n10059) );
  INVX0 U10259 ( .INP(n10174), .ZN(n10060) );
  INVX0 U10260 ( .INP(n10174), .ZN(n10061) );
  INVX0 U10261 ( .INP(n10174), .ZN(n10062) );
  INVX0 U10262 ( .INP(n10174), .ZN(n10063) );
  INVX0 U10263 ( .INP(n10174), .ZN(n10064) );
  INVX0 U10264 ( .INP(n10173), .ZN(n10065) );
  INVX0 U10265 ( .INP(n10173), .ZN(n10066) );
  INVX0 U10266 ( .INP(n10173), .ZN(n10067) );
  INVX0 U10267 ( .INP(n10173), .ZN(n10068) );
  INVX0 U10268 ( .INP(n10173), .ZN(n10069) );
  INVX0 U10269 ( .INP(n10173), .ZN(n10070) );
  INVX0 U10270 ( .INP(n10172), .ZN(n10071) );
  INVX0 U10271 ( .INP(n10172), .ZN(n10072) );
  INVX0 U10272 ( .INP(n10172), .ZN(n10073) );
  INVX0 U10273 ( .INP(n10172), .ZN(n10074) );
  INVX0 U10274 ( .INP(n10172), .ZN(n10075) );
  INVX0 U10275 ( .INP(n10172), .ZN(n10076) );
  INVX0 U10276 ( .INP(n10171), .ZN(n10077) );
  INVX0 U10277 ( .INP(n10171), .ZN(n10078) );
  INVX0 U10278 ( .INP(n10171), .ZN(n10079) );
  INVX0 U10279 ( .INP(n10171), .ZN(n10080) );
  INVX0 U10280 ( .INP(n10171), .ZN(n10081) );
  INVX0 U10281 ( .INP(n10171), .ZN(n10082) );
  INVX0 U10282 ( .INP(n10170), .ZN(n10083) );
  INVX0 U10283 ( .INP(n10170), .ZN(n10084) );
  INVX0 U10284 ( .INP(n10170), .ZN(n10085) );
  INVX0 U10285 ( .INP(n10170), .ZN(n10086) );
  INVX0 U10286 ( .INP(n10170), .ZN(n10087) );
  INVX0 U10287 ( .INP(n10170), .ZN(n10088) );
  INVX0 U10288 ( .INP(n10169), .ZN(n10089) );
  INVX0 U10289 ( .INP(n10169), .ZN(n10090) );
  INVX0 U10290 ( .INP(n10169), .ZN(n10091) );
  INVX0 U10291 ( .INP(n10169), .ZN(n10092) );
  INVX0 U10292 ( .INP(n10169), .ZN(n10093) );
  INVX0 U10293 ( .INP(n10169), .ZN(n10094) );
  INVX0 U10294 ( .INP(n10168), .ZN(n10095) );
  INVX0 U10295 ( .INP(n10168), .ZN(n10096) );
  INVX0 U10296 ( .INP(n10168), .ZN(n10097) );
  INVX0 U10297 ( .INP(n10168), .ZN(n10098) );
  INVX0 U10298 ( .INP(n10168), .ZN(n10099) );
  INVX0 U10299 ( .INP(n10168), .ZN(n10100) );
  INVX0 U10300 ( .INP(n10171), .ZN(n10101) );
  INVX0 U10301 ( .INP(n10170), .ZN(n10102) );
  INVX0 U10302 ( .INP(n10169), .ZN(n10103) );
  INVX0 U10303 ( .INP(n10168), .ZN(n10104) );
  INVX0 U10304 ( .INP(n10171), .ZN(n10105) );
  INVX0 U10305 ( .INP(n10175), .ZN(n10106) );
  INVX0 U10306 ( .INP(n10171), .ZN(n10107) );
  INVX0 U10307 ( .INP(n10170), .ZN(n10108) );
  INVX0 U10308 ( .INP(n10169), .ZN(n10109) );
  INVX0 U10309 ( .INP(n10168), .ZN(n10110) );
  INVX0 U10310 ( .INP(n10175), .ZN(n10111) );
  INVX0 U10311 ( .INP(n10170), .ZN(n10112) );
  INVX0 U10312 ( .INP(n10169), .ZN(n10113) );
  INVX0 U10313 ( .INP(n10168), .ZN(n10114) );
  INVX0 U10314 ( .INP(n10174), .ZN(n10115) );
  INVX0 U10315 ( .INP(n10174), .ZN(n10116) );
  INVX0 U10316 ( .INP(n10169), .ZN(n10117) );
  INVX0 U10317 ( .INP(n10175), .ZN(n10118) );
  INVX0 U10318 ( .INP(n10176), .ZN(n10119) );
  INVX0 U10319 ( .INP(n10168), .ZN(n10120) );
  INVX0 U10320 ( .INP(n10175), .ZN(n10121) );
  INVX0 U10321 ( .INP(n10174), .ZN(n10122) );
  INVX0 U10322 ( .INP(n10173), .ZN(n10123) );
  INVX0 U10323 ( .INP(n10172), .ZN(n10124) );
  INVX0 U10324 ( .INP(n10172), .ZN(n10125) );
  INVX0 U10325 ( .INP(n10176), .ZN(n10126) );
  INVX0 U10326 ( .INP(n10177), .ZN(n10127) );
  INVX0 U10327 ( .INP(n10171), .ZN(n10128) );
  INVX0 U10328 ( .INP(n10170), .ZN(n10129) );
  INVX0 U10329 ( .INP(n10169), .ZN(n10130) );
  INVX0 U10330 ( .INP(n10173), .ZN(n10131) );
  INVX0 U10331 ( .INP(n10172), .ZN(n10132) );
  INVX0 U10332 ( .INP(n10176), .ZN(n10133) );
  INVX0 U10333 ( .INP(n10177), .ZN(n10134) );
  INVX0 U10334 ( .INP(n10175), .ZN(n10135) );
  INVX0 U10335 ( .INP(n10174), .ZN(n10136) );
  INVX0 U10336 ( .INP(n10176), .ZN(n10137) );
  INVX0 U10337 ( .INP(n10171), .ZN(n10138) );
  INVX0 U10338 ( .INP(n10170), .ZN(n10139) );
  INVX0 U10339 ( .INP(n10169), .ZN(n10140) );
  INVX0 U10340 ( .INP(n10168), .ZN(n10141) );
  INVX0 U10341 ( .INP(n10169), .ZN(n10142) );
  INVX0 U10342 ( .INP(n10168), .ZN(n10143) );
  INVX0 U10343 ( .INP(n10172), .ZN(n10144) );
  INVX0 U10344 ( .INP(n10172), .ZN(n10145) );
  INVX0 U10345 ( .INP(n10168), .ZN(n10146) );
  INVX0 U10346 ( .INP(n10170), .ZN(n10147) );
  INVX0 U10347 ( .INP(n10172), .ZN(n10148) );
  INVX0 U10348 ( .INP(n10171), .ZN(n10149) );
  INVX0 U10349 ( .INP(n10170), .ZN(n10150) );
  INVX0 U10350 ( .INP(n10169), .ZN(n10151) );
  INVX0 U10351 ( .INP(n10168), .ZN(n10152) );
  INVX0 U10352 ( .INP(n10173), .ZN(n10153) );
  INVX0 U10353 ( .INP(n10172), .ZN(n10154) );
  INVX0 U10354 ( .INP(n10176), .ZN(n10155) );
  INVX0 U10355 ( .INP(n10175), .ZN(n10156) );
  INVX0 U10356 ( .INP(n10171), .ZN(n10157) );
  INVX0 U10357 ( .INP(n10170), .ZN(n10158) );
  INVX0 U10358 ( .INP(n10173), .ZN(n10159) );
  INVX0 U10359 ( .INP(n10173), .ZN(n10160) );
  INVX0 U10360 ( .INP(n10174), .ZN(n10161) );
  INVX0 U10361 ( .INP(n10175), .ZN(n10162) );
  INVX0 U10362 ( .INP(n10174), .ZN(n10163) );
  INVX0 U10363 ( .INP(n10171), .ZN(n10164) );
  INVX0 U10364 ( .INP(n10170), .ZN(n10165) );
  INVX0 U10365 ( .INP(n10169), .ZN(n10166) );
  INVX0 U10366 ( .INP(n10168), .ZN(n10167) );
  NBUFFX2 U10367 ( .INP(n10228), .Z(n10178) );
  NBUFFX2 U10368 ( .INP(n10228), .Z(n10179) );
  NBUFFX2 U10369 ( .INP(n10227), .Z(n10180) );
  NBUFFX2 U10370 ( .INP(n10227), .Z(n10181) );
  NBUFFX2 U10371 ( .INP(n10227), .Z(n10182) );
  NBUFFX2 U10372 ( .INP(n10226), .Z(n10183) );
  NBUFFX2 U10373 ( .INP(n10226), .Z(n10184) );
  NBUFFX2 U10374 ( .INP(n10226), .Z(n10185) );
  NBUFFX2 U10375 ( .INP(n10225), .Z(n10186) );
  NBUFFX2 U10376 ( .INP(n10225), .Z(n10187) );
  NBUFFX2 U10377 ( .INP(n10225), .Z(n10188) );
  NBUFFX2 U10378 ( .INP(n10224), .Z(n10189) );
  NBUFFX2 U10379 ( .INP(n10224), .Z(n10190) );
  NBUFFX2 U10380 ( .INP(n10224), .Z(n10191) );
  NBUFFX2 U10381 ( .INP(n10223), .Z(n10192) );
  NBUFFX2 U10382 ( .INP(n10223), .Z(n10193) );
  NBUFFX2 U10383 ( .INP(n10223), .Z(n10194) );
  NBUFFX2 U10384 ( .INP(n10222), .Z(n10195) );
  NBUFFX2 U10385 ( .INP(n10222), .Z(n10196) );
  NBUFFX2 U10386 ( .INP(n10222), .Z(n10197) );
  NBUFFX2 U10387 ( .INP(n10221), .Z(n10198) );
  NBUFFX2 U10388 ( .INP(n10221), .Z(n10199) );
  NBUFFX2 U10389 ( .INP(n10221), .Z(n10200) );
  NBUFFX2 U10390 ( .INP(n10220), .Z(n10201) );
  NBUFFX2 U10391 ( .INP(n10220), .Z(n10202) );
  NBUFFX2 U10392 ( .INP(n10220), .Z(n10203) );
  NBUFFX2 U10393 ( .INP(n10219), .Z(n10204) );
  NBUFFX2 U10394 ( .INP(n10219), .Z(n10205) );
  NBUFFX2 U10395 ( .INP(n10219), .Z(n10206) );
  NBUFFX2 U10396 ( .INP(n10218), .Z(n10207) );
  NBUFFX2 U10397 ( .INP(n10218), .Z(n10208) );
  NBUFFX2 U10398 ( .INP(n10218), .Z(n10209) );
  NBUFFX2 U10399 ( .INP(n10217), .Z(n10210) );
  NBUFFX2 U10400 ( .INP(n10217), .Z(n10211) );
  NBUFFX2 U10401 ( .INP(n10217), .Z(n10212) );
  NBUFFX2 U10402 ( .INP(n10216), .Z(n10213) );
  NBUFFX2 U10403 ( .INP(n10216), .Z(n10214) );
  NBUFFX2 U10404 ( .INP(n10216), .Z(n10215) );
  NBUFFX2 U10405 ( .INP(n10233), .Z(n10216) );
  NBUFFX2 U10406 ( .INP(n10232), .Z(n10217) );
  NBUFFX2 U10407 ( .INP(n10232), .Z(n10218) );
  NBUFFX2 U10408 ( .INP(n10232), .Z(n10219) );
  NBUFFX2 U10409 ( .INP(n10231), .Z(n10220) );
  NBUFFX2 U10410 ( .INP(n10231), .Z(n10221) );
  NBUFFX2 U10411 ( .INP(n10231), .Z(n10222) );
  NBUFFX2 U10412 ( .INP(n10230), .Z(n10223) );
  NBUFFX2 U10413 ( .INP(n10230), .Z(n10224) );
  NBUFFX2 U10414 ( .INP(n10230), .Z(n10225) );
  NBUFFX2 U10415 ( .INP(n10229), .Z(n10226) );
  NBUFFX2 U10416 ( .INP(n10229), .Z(n10227) );
  NBUFFX2 U10417 ( .INP(n10229), .Z(n10228) );
  NBUFFX2 U10418 ( .INP(RESET), .Z(n10229) );
  NBUFFX2 U10419 ( .INP(RESET), .Z(n10230) );
  NBUFFX2 U10420 ( .INP(RESET), .Z(n10231) );
  NBUFFX2 U10421 ( .INP(RESET), .Z(n10232) );
  NBUFFX2 U10422 ( .INP(RESET), .Z(n10233) );
  INVX0 U10423 ( .INP(n10178), .ZN(n10234) );
  INVX0 U10424 ( .INP(n10178), .ZN(n10235) );
  INVX0 U10425 ( .INP(n10178), .ZN(n10236) );
  INVX0 U10426 ( .INP(n10178), .ZN(n10237) );
  INVX0 U10427 ( .INP(n10178), .ZN(n10238) );
  INVX0 U10428 ( .INP(n10178), .ZN(n10239) );
  INVX0 U10429 ( .INP(n10178), .ZN(n10240) );
  INVX0 U10430 ( .INP(n10178), .ZN(n10241) );
  INVX0 U10431 ( .INP(n10179), .ZN(n10242) );
  INVX0 U10432 ( .INP(n10179), .ZN(n10243) );
  INVX0 U10433 ( .INP(n10179), .ZN(n10244) );
  INVX0 U10434 ( .INP(n10180), .ZN(n10245) );
  INVX0 U10435 ( .INP(n10180), .ZN(n10246) );
  INVX0 U10436 ( .INP(n10180), .ZN(n10247) );
  INVX0 U10437 ( .INP(n10180), .ZN(n10248) );
  INVX0 U10438 ( .INP(n10180), .ZN(n10249) );
  INVX0 U10439 ( .INP(n10180), .ZN(n10250) );
  INVX0 U10440 ( .INP(n10180), .ZN(n10251) );
  INVX0 U10441 ( .INP(n10180), .ZN(n10252) );
  INVX0 U10442 ( .INP(n10181), .ZN(n10253) );
  INVX0 U10443 ( .INP(n10181), .ZN(n10254) );
  INVX0 U10444 ( .INP(n10181), .ZN(n10255) );
  INVX0 U10445 ( .INP(n10181), .ZN(n10256) );
  INVX0 U10446 ( .INP(n10181), .ZN(n10257) );
  INVX0 U10447 ( .INP(n10181), .ZN(n10258) );
  INVX0 U10448 ( .INP(n10181), .ZN(n10259) );
  INVX0 U10449 ( .INP(n10181), .ZN(n10260) );
  INVX0 U10450 ( .INP(n10182), .ZN(n10261) );
  INVX0 U10451 ( .INP(n10182), .ZN(n10262) );
  INVX0 U10452 ( .INP(n10182), .ZN(n10263) );
  INVX0 U10453 ( .INP(n10182), .ZN(n10264) );
  INVX0 U10454 ( .INP(n10182), .ZN(n10265) );
  INVX0 U10455 ( .INP(n10182), .ZN(n10266) );
  INVX0 U10456 ( .INP(n10182), .ZN(n10267) );
  INVX0 U10457 ( .INP(n10183), .ZN(n10268) );
  INVX0 U10458 ( .INP(n10183), .ZN(n10269) );
  INVX0 U10459 ( .INP(n10183), .ZN(n10270) );
  INVX0 U10460 ( .INP(n10183), .ZN(n10271) );
  INVX0 U10461 ( .INP(n10183), .ZN(n10272) );
  INVX0 U10462 ( .INP(n10183), .ZN(n10273) );
  INVX0 U10463 ( .INP(n10183), .ZN(n10274) );
  INVX0 U10464 ( .INP(n10183), .ZN(n10275) );
  INVX0 U10465 ( .INP(n10184), .ZN(n10276) );
  INVX0 U10466 ( .INP(n10184), .ZN(n10277) );
  INVX0 U10467 ( .INP(n10184), .ZN(n10278) );
  INVX0 U10468 ( .INP(n10184), .ZN(n10279) );
  INVX0 U10469 ( .INP(n10184), .ZN(n10280) );
  INVX0 U10470 ( .INP(n10184), .ZN(n10281) );
  INVX0 U10471 ( .INP(n10184), .ZN(n10282) );
  INVX0 U10472 ( .INP(n10185), .ZN(n10283) );
  INVX0 U10473 ( .INP(n10185), .ZN(n10284) );
  INVX0 U10474 ( .INP(n10185), .ZN(n10285) );
  INVX0 U10475 ( .INP(n10185), .ZN(n10286) );
  INVX0 U10476 ( .INP(n10185), .ZN(n10287) );
  INVX0 U10477 ( .INP(n10185), .ZN(n10288) );
  INVX0 U10478 ( .INP(n10185), .ZN(n10289) );
  INVX0 U10479 ( .INP(n10185), .ZN(n10290) );
  INVX0 U10480 ( .INP(n10186), .ZN(n10291) );
  INVX0 U10481 ( .INP(n10186), .ZN(n10292) );
  INVX0 U10482 ( .INP(n10186), .ZN(n10293) );
  INVX0 U10483 ( .INP(n10186), .ZN(n10294) );
  INVX0 U10484 ( .INP(n10186), .ZN(n10295) );
  INVX0 U10485 ( .INP(n10186), .ZN(n10296) );
  INVX0 U10486 ( .INP(n10186), .ZN(n10297) );
  INVX0 U10487 ( .INP(n10186), .ZN(n10298) );
  INVX0 U10488 ( .INP(n10187), .ZN(n10299) );
  INVX0 U10489 ( .INP(n10187), .ZN(n10300) );
  INVX0 U10490 ( .INP(n10187), .ZN(n10301) );
  INVX0 U10491 ( .INP(n10187), .ZN(n10302) );
  INVX0 U10492 ( .INP(n10187), .ZN(n10303) );
  INVX0 U10493 ( .INP(n10187), .ZN(n10304) );
  INVX0 U10494 ( .INP(n10187), .ZN(n10305) );
  INVX0 U10495 ( .INP(n10187), .ZN(n10306) );
  INVX0 U10496 ( .INP(n10188), .ZN(n10307) );
  INVX0 U10497 ( .INP(n10188), .ZN(n10308) );
  INVX0 U10498 ( .INP(n10188), .ZN(n10309) );
  INVX0 U10499 ( .INP(n10188), .ZN(n10310) );
  INVX0 U10500 ( .INP(n10188), .ZN(n10311) );
  INVX0 U10501 ( .INP(n10188), .ZN(n10312) );
  INVX0 U10502 ( .INP(n10188), .ZN(n10313) );
  INVX0 U10503 ( .INP(n10188), .ZN(n10314) );
  INVX0 U10504 ( .INP(n10189), .ZN(n10315) );
  INVX0 U10505 ( .INP(n10189), .ZN(n10316) );
  INVX0 U10506 ( .INP(n10189), .ZN(n10317) );
  INVX0 U10507 ( .INP(n10189), .ZN(n10318) );
  INVX0 U10508 ( .INP(n10189), .ZN(n10319) );
  INVX0 U10509 ( .INP(n10189), .ZN(n10320) );
  INVX0 U10510 ( .INP(n10189), .ZN(n10321) );
  INVX0 U10511 ( .INP(n10189), .ZN(n10322) );
  INVX0 U10512 ( .INP(n10190), .ZN(n10323) );
  INVX0 U10513 ( .INP(n10190), .ZN(n10324) );
  INVX0 U10514 ( .INP(n10190), .ZN(n10325) );
  INVX0 U10515 ( .INP(n10190), .ZN(n10326) );
  INVX0 U10516 ( .INP(n10190), .ZN(n10327) );
  INVX0 U10517 ( .INP(n10190), .ZN(n10328) );
  INVX0 U10518 ( .INP(n10190), .ZN(n10329) );
  INVX0 U10519 ( .INP(n10190), .ZN(n10330) );
  INVX0 U10520 ( .INP(n10191), .ZN(n10331) );
  INVX0 U10521 ( .INP(n10191), .ZN(n10332) );
  NBUFFX2 U10522 ( .INP(n10515), .Z(n10477) );
  NBUFFX2 U10523 ( .INP(n10515), .Z(n10478) );
  NBUFFX2 U10524 ( .INP(n10514), .Z(n10479) );
  NBUFFX2 U10525 ( .INP(n10514), .Z(n10480) );
  NBUFFX2 U10526 ( .INP(n10514), .Z(n10481) );
  NBUFFX2 U10527 ( .INP(n10513), .Z(n10482) );
  NBUFFX2 U10528 ( .INP(n10513), .Z(n10483) );
  NBUFFX2 U10529 ( .INP(n10513), .Z(n10484) );
  NBUFFX2 U10530 ( .INP(n10512), .Z(n10485) );
  NBUFFX2 U10531 ( .INP(n10512), .Z(n10486) );
  NBUFFX2 U10532 ( .INP(n10512), .Z(n10487) );
  NBUFFX2 U10533 ( .INP(n10511), .Z(n10488) );
  NBUFFX2 U10534 ( .INP(n10511), .Z(n10489) );
  NBUFFX2 U10535 ( .INP(n10511), .Z(n10490) );
  NBUFFX2 U10536 ( .INP(n10510), .Z(n10491) );
  NBUFFX2 U10537 ( .INP(n10510), .Z(n10492) );
  NBUFFX2 U10538 ( .INP(n10510), .Z(n10493) );
  NBUFFX2 U10539 ( .INP(n10509), .Z(n10494) );
  NBUFFX2 U10540 ( .INP(n10509), .Z(n10495) );
  NBUFFX2 U10541 ( .INP(n10509), .Z(n10496) );
  NBUFFX2 U10542 ( .INP(n10508), .Z(n10497) );
  NBUFFX2 U10543 ( .INP(n10508), .Z(n10498) );
  NBUFFX2 U10544 ( .INP(n10508), .Z(n10499) );
  NBUFFX2 U10545 ( .INP(n10507), .Z(n10500) );
  NBUFFX2 U10546 ( .INP(n10507), .Z(n10501) );
  NBUFFX2 U10547 ( .INP(n10507), .Z(n10502) );
  NBUFFX2 U10548 ( .INP(n10506), .Z(n10503) );
  NBUFFX2 U10549 ( .INP(n10506), .Z(n10504) );
  NBUFFX2 U10550 ( .INP(n10506), .Z(n10505) );
  NBUFFX2 U10551 ( .INP(CK), .Z(n10506) );
  NBUFFX2 U10552 ( .INP(CK), .Z(n10507) );
  NBUFFX2 U10553 ( .INP(n10515), .Z(n10508) );
  NBUFFX2 U10554 ( .INP(CK), .Z(n10509) );
  NBUFFX2 U10555 ( .INP(n10511), .Z(n10510) );
  NBUFFX2 U10556 ( .INP(CK), .Z(n10511) );
  NBUFFX2 U10557 ( .INP(n10506), .Z(n10512) );
  NBUFFX2 U10558 ( .INP(n10507), .Z(n10513) );
  NBUFFX2 U10559 ( .INP(n10509), .Z(n10514) );
  NBUFFX2 U10560 ( .INP(n10346), .Z(n10515) );
  INVX0 U10561 ( .INP(n10516), .ZN(n98) );
  NOR2X0 U10562 ( .IN1(n10517), .IN2(n10518), .QN(n10516) );
  NAND2X0 U10563 ( .IN1(n10519), .IN2(n10520), .QN(n10518) );
  NAND2X0 U10564 ( .IN1(n9950), .IN2(n10521), .QN(n10520) );
  NAND2X0 U10565 ( .IN1(n2152), .IN2(CRC_OUT_9_12), .QN(n10519) );
  NAND2X0 U10566 ( .IN1(n10522), .IN2(n10523), .QN(n10517) );
  INVX0 U10567 ( .INP(n10524), .ZN(n10523) );
  NOR2X0 U10568 ( .IN1(n9923), .IN2(n10526), .QN(n10524) );
  NAND2X0 U10569 ( .IN1(WX520), .IN2(n2339), .QN(n10522) );
  INVX0 U10570 ( .INP(n10527), .ZN(n95) );
  NOR2X0 U10571 ( .IN1(n10528), .IN2(n10529), .QN(n10527) );
  NAND2X0 U10572 ( .IN1(n10530), .IN2(n10531), .QN(n10529) );
  NAND2X0 U10573 ( .IN1(n9948), .IN2(n10532), .QN(n10531) );
  NAND2X0 U10574 ( .IN1(n2152), .IN2(CRC_OUT_9_13), .QN(n10530) );
  NAND2X0 U10575 ( .IN1(n10533), .IN2(n10534), .QN(n10528) );
  INVX0 U10576 ( .INP(n10535), .ZN(n10534) );
  NOR2X0 U10577 ( .IN1(n9926), .IN2(n10536), .QN(n10535) );
  NAND2X0 U10578 ( .IN1(WX518), .IN2(n2339), .QN(n10533) );
  INVX0 U10579 ( .INP(n10537), .ZN(n92) );
  NOR2X0 U10580 ( .IN1(n10538), .IN2(n10539), .QN(n10537) );
  NAND2X0 U10581 ( .IN1(n10540), .IN2(n10541), .QN(n10539) );
  NAND2X0 U10582 ( .IN1(n9948), .IN2(n10542), .QN(n10541) );
  NAND2X0 U10583 ( .IN1(n2152), .IN2(CRC_OUT_9_14), .QN(n10540) );
  NAND2X0 U10584 ( .IN1(n10543), .IN2(n10544), .QN(n10538) );
  NAND2X0 U10585 ( .IN1(n10545), .IN2(n2153), .QN(n10544) );
  NAND2X0 U10586 ( .IN1(WX516), .IN2(n2339), .QN(n10543) );
  INVX0 U10587 ( .INP(n10546), .ZN(n89) );
  NOR2X0 U10588 ( .IN1(n10547), .IN2(n10548), .QN(n10546) );
  NAND2X0 U10589 ( .IN1(n10549), .IN2(n10550), .QN(n10548) );
  NAND2X0 U10590 ( .IN1(n9948), .IN2(n10551), .QN(n10550) );
  NAND2X0 U10591 ( .IN1(n2152), .IN2(CRC_OUT_9_15), .QN(n10549) );
  NAND2X0 U10592 ( .IN1(n10552), .IN2(n10553), .QN(n10547) );
  INVX0 U10593 ( .INP(n10554), .ZN(n10553) );
  NOR2X0 U10594 ( .IN1(n9926), .IN2(n10555), .QN(n10554) );
  NAND2X0 U10595 ( .IN1(WX514), .IN2(n2339), .QN(n10552) );
  INVX0 U10596 ( .INP(n10556), .ZN(n86) );
  NOR2X0 U10597 ( .IN1(n10557), .IN2(n10558), .QN(n10556) );
  NAND2X0 U10598 ( .IN1(n10559), .IN2(n10560), .QN(n10558) );
  INVX0 U10599 ( .INP(n10561), .ZN(n10560) );
  NOR2X0 U10600 ( .IN1(n10562), .IN2(n9927), .QN(n10561) );
  NAND2X0 U10601 ( .IN1(n2152), .IN2(CRC_OUT_9_16), .QN(n10559) );
  NAND2X0 U10602 ( .IN1(n10564), .IN2(n10565), .QN(n10557) );
  INVX0 U10603 ( .INP(n10566), .ZN(n10565) );
  NOR2X0 U10604 ( .IN1(n9926), .IN2(n10567), .QN(n10566) );
  NAND2X0 U10605 ( .IN1(WX512), .IN2(n2339), .QN(n10564) );
  INVX0 U10606 ( .INP(n10568), .ZN(n839) );
  INVX0 U10607 ( .INP(n10569), .ZN(n838) );
  INVX0 U10608 ( .INP(n10570), .ZN(n837) );
  INVX0 U10609 ( .INP(n10571), .ZN(n836) );
  INVX0 U10610 ( .INP(n10572), .ZN(n835) );
  INVX0 U10611 ( .INP(n10573), .ZN(n834) );
  INVX0 U10612 ( .INP(n10574), .ZN(n833) );
  INVX0 U10613 ( .INP(n10575), .ZN(n832) );
  INVX0 U10614 ( .INP(n10576), .ZN(n831) );
  INVX0 U10615 ( .INP(n10577), .ZN(n830) );
  INVX0 U10616 ( .INP(n10578), .ZN(n83) );
  NOR2X0 U10617 ( .IN1(n10579), .IN2(n10580), .QN(n10578) );
  NAND2X0 U10618 ( .IN1(n10581), .IN2(n10582), .QN(n10580) );
  NAND2X0 U10619 ( .IN1(n9949), .IN2(n10583), .QN(n10582) );
  NAND2X0 U10620 ( .IN1(n2152), .IN2(CRC_OUT_9_17), .QN(n10581) );
  NAND2X0 U10621 ( .IN1(n10584), .IN2(n10585), .QN(n10579) );
  INVX0 U10622 ( .INP(n10586), .ZN(n10585) );
  NOR2X0 U10623 ( .IN1(n9926), .IN2(n10587), .QN(n10586) );
  NAND2X0 U10624 ( .IN1(WX510), .IN2(n2339), .QN(n10584) );
  INVX0 U10625 ( .INP(n10588), .ZN(n829) );
  INVX0 U10626 ( .INP(n10589), .ZN(n828) );
  INVX0 U10627 ( .INP(n10590), .ZN(n827) );
  INVX0 U10628 ( .INP(n10591), .ZN(n826) );
  INVX0 U10629 ( .INP(n10592), .ZN(n825) );
  INVX0 U10630 ( .INP(n10593), .ZN(n824) );
  INVX0 U10631 ( .INP(n10594), .ZN(n823) );
  INVX0 U10632 ( .INP(n10595), .ZN(n822) );
  INVX0 U10633 ( .INP(n10596), .ZN(n821) );
  INVX0 U10634 ( .INP(n10597), .ZN(n820) );
  INVX0 U10635 ( .INP(n10598), .ZN(n819) );
  INVX0 U10636 ( .INP(n10599), .ZN(n818) );
  INVX0 U10637 ( .INP(n10600), .ZN(n817) );
  INVX0 U10638 ( .INP(n10601), .ZN(n816) );
  INVX0 U10639 ( .INP(n10602), .ZN(n815) );
  INVX0 U10640 ( .INP(n10603), .ZN(n814) );
  INVX0 U10641 ( .INP(n10604), .ZN(n813) );
  INVX0 U10642 ( .INP(n10605), .ZN(n812) );
  INVX0 U10643 ( .INP(n10606), .ZN(n811) );
  INVX0 U10644 ( .INP(n10607), .ZN(n810) );
  INVX0 U10645 ( .INP(n10608), .ZN(n809) );
  INVX0 U10646 ( .INP(n10609), .ZN(n80) );
  NOR2X0 U10647 ( .IN1(n10610), .IN2(n10611), .QN(n10609) );
  NAND2X0 U10648 ( .IN1(n10612), .IN2(n10613), .QN(n10611) );
  NAND2X0 U10649 ( .IN1(n9949), .IN2(n10614), .QN(n10613) );
  NAND2X0 U10650 ( .IN1(n2152), .IN2(CRC_OUT_9_18), .QN(n10612) );
  NAND2X0 U10651 ( .IN1(n10615), .IN2(n10616), .QN(n10610) );
  NAND2X0 U10652 ( .IN1(n10617), .IN2(n2153), .QN(n10616) );
  NAND2X0 U10653 ( .IN1(WX508), .IN2(n2339), .QN(n10615) );
  INVX0 U10654 ( .INP(n10618), .ZN(n77) );
  NOR2X0 U10655 ( .IN1(n10619), .IN2(n10620), .QN(n10618) );
  NAND2X0 U10656 ( .IN1(n10621), .IN2(n10622), .QN(n10620) );
  NAND2X0 U10657 ( .IN1(n9949), .IN2(n10623), .QN(n10622) );
  NAND2X0 U10658 ( .IN1(test_so10), .IN2(n2152), .QN(n10621) );
  NAND2X0 U10659 ( .IN1(n10624), .IN2(n10625), .QN(n10619) );
  INVX0 U10660 ( .INP(n10626), .ZN(n10625) );
  NOR2X0 U10661 ( .IN1(n9926), .IN2(n10627), .QN(n10626) );
  NAND2X0 U10662 ( .IN1(WX506), .IN2(n2339), .QN(n10624) );
  INVX0 U10663 ( .INP(n10628), .ZN(n74) );
  NOR2X0 U10664 ( .IN1(n10629), .IN2(n10630), .QN(n10628) );
  NAND2X0 U10665 ( .IN1(n10631), .IN2(n10632), .QN(n10630) );
  INVX0 U10666 ( .INP(n10633), .ZN(n10632) );
  NOR2X0 U10667 ( .IN1(n10634), .IN2(n9927), .QN(n10633) );
  NAND2X0 U10668 ( .IN1(n2152), .IN2(CRC_OUT_9_20), .QN(n10631) );
  NAND2X0 U10669 ( .IN1(n10635), .IN2(n10636), .QN(n10629) );
  INVX0 U10670 ( .INP(n10637), .ZN(n10636) );
  NOR2X0 U10671 ( .IN1(n9926), .IN2(n10638), .QN(n10637) );
  NAND2X0 U10672 ( .IN1(WX504), .IN2(n2339), .QN(n10635) );
  INVX0 U10673 ( .INP(n10639), .ZN(n71) );
  NOR2X0 U10674 ( .IN1(n10640), .IN2(n10641), .QN(n10639) );
  NAND2X0 U10675 ( .IN1(n10642), .IN2(n10643), .QN(n10641) );
  NAND2X0 U10676 ( .IN1(n9949), .IN2(n10644), .QN(n10643) );
  NAND2X0 U10677 ( .IN1(n2152), .IN2(CRC_OUT_9_21), .QN(n10642) );
  NAND2X0 U10678 ( .IN1(n10645), .IN2(n10646), .QN(n10640) );
  INVX0 U10679 ( .INP(n10647), .ZN(n10646) );
  NOR2X0 U10680 ( .IN1(n9926), .IN2(n10648), .QN(n10647) );
  NAND2X0 U10681 ( .IN1(WX502), .IN2(n2339), .QN(n10645) );
  INVX0 U10682 ( .INP(n10649), .ZN(n68) );
  NOR2X0 U10683 ( .IN1(n10650), .IN2(n10651), .QN(n10649) );
  NAND2X0 U10684 ( .IN1(n10652), .IN2(n10653), .QN(n10651) );
  NAND2X0 U10685 ( .IN1(n9949), .IN2(n10654), .QN(n10653) );
  NAND2X0 U10686 ( .IN1(n2152), .IN2(CRC_OUT_9_22), .QN(n10652) );
  NAND2X0 U10687 ( .IN1(n10655), .IN2(n10656), .QN(n10650) );
  NAND2X0 U10688 ( .IN1(n10657), .IN2(n2153), .QN(n10656) );
  NAND2X0 U10689 ( .IN1(WX500), .IN2(n2339), .QN(n10655) );
  INVX0 U10690 ( .INP(n10658), .ZN(n65) );
  NOR2X0 U10691 ( .IN1(n10659), .IN2(n10660), .QN(n10658) );
  NAND2X0 U10692 ( .IN1(n10661), .IN2(n10662), .QN(n10660) );
  NAND2X0 U10693 ( .IN1(n9949), .IN2(n10663), .QN(n10662) );
  NAND2X0 U10694 ( .IN1(n2152), .IN2(CRC_OUT_9_23), .QN(n10661) );
  NAND2X0 U10695 ( .IN1(n10664), .IN2(n10665), .QN(n10659) );
  INVX0 U10696 ( .INP(n10666), .ZN(n10665) );
  NOR2X0 U10697 ( .IN1(n9925), .IN2(n10667), .QN(n10666) );
  NAND2X0 U10698 ( .IN1(WX498), .IN2(n2339), .QN(n10664) );
  INVX0 U10699 ( .INP(n10668), .ZN(n62) );
  NOR2X0 U10700 ( .IN1(n10669), .IN2(n10670), .QN(n10668) );
  NAND2X0 U10701 ( .IN1(n10671), .IN2(n10672), .QN(n10670) );
  INVX0 U10702 ( .INP(n10673), .ZN(n10672) );
  NOR2X0 U10703 ( .IN1(n10674), .IN2(n9927), .QN(n10673) );
  NAND2X0 U10704 ( .IN1(n2152), .IN2(CRC_OUT_9_24), .QN(n10671) );
  NAND2X0 U10705 ( .IN1(n10675), .IN2(n10676), .QN(n10669) );
  INVX0 U10706 ( .INP(n10677), .ZN(n10676) );
  NOR2X0 U10707 ( .IN1(n9925), .IN2(n10678), .QN(n10677) );
  NAND2X0 U10708 ( .IN1(WX496), .IN2(n2339), .QN(n10675) );
  INVX0 U10709 ( .INP(n10679), .ZN(n598) );
  INVX0 U10710 ( .INP(n10680), .ZN(n597) );
  INVX0 U10711 ( .INP(n10681), .ZN(n596) );
  INVX0 U10712 ( .INP(n10682), .ZN(n595) );
  INVX0 U10713 ( .INP(n10683), .ZN(n594) );
  INVX0 U10714 ( .INP(n10684), .ZN(n593) );
  INVX0 U10715 ( .INP(n10685), .ZN(n592) );
  INVX0 U10716 ( .INP(n10686), .ZN(n591) );
  INVX0 U10717 ( .INP(n10687), .ZN(n590) );
  INVX0 U10718 ( .INP(n10688), .ZN(n59) );
  NOR2X0 U10719 ( .IN1(n10689), .IN2(n10690), .QN(n10688) );
  NAND2X0 U10720 ( .IN1(n10691), .IN2(n10692), .QN(n10690) );
  NAND2X0 U10721 ( .IN1(n9949), .IN2(n10693), .QN(n10692) );
  NAND2X0 U10722 ( .IN1(n2152), .IN2(CRC_OUT_9_25), .QN(n10691) );
  NAND2X0 U10723 ( .IN1(n10694), .IN2(n10695), .QN(n10689) );
  INVX0 U10724 ( .INP(n10696), .ZN(n10695) );
  NOR2X0 U10725 ( .IN1(n9925), .IN2(n10697), .QN(n10696) );
  NAND2X0 U10726 ( .IN1(WX494), .IN2(n2339), .QN(n10694) );
  INVX0 U10727 ( .INP(n10698), .ZN(n589) );
  INVX0 U10728 ( .INP(n10699), .ZN(n588) );
  INVX0 U10729 ( .INP(n10700), .ZN(n587) );
  INVX0 U10730 ( .INP(n10701), .ZN(n586) );
  INVX0 U10731 ( .INP(n10702), .ZN(n585) );
  INVX0 U10732 ( .INP(n10703), .ZN(n584) );
  INVX0 U10733 ( .INP(n10704), .ZN(n583) );
  INVX0 U10734 ( .INP(n10705), .ZN(n582) );
  INVX0 U10735 ( .INP(n10706), .ZN(n581) );
  INVX0 U10736 ( .INP(n10707), .ZN(n580) );
  INVX0 U10737 ( .INP(n10708), .ZN(n579) );
  INVX0 U10738 ( .INP(n10709), .ZN(n578) );
  INVX0 U10739 ( .INP(n10710), .ZN(n577) );
  INVX0 U10740 ( .INP(n10711), .ZN(n576) );
  INVX0 U10741 ( .INP(n10712), .ZN(n575) );
  INVX0 U10742 ( .INP(n10713), .ZN(n574) );
  INVX0 U10743 ( .INP(n10714), .ZN(n573) );
  INVX0 U10744 ( .INP(n10715), .ZN(n572) );
  INVX0 U10745 ( .INP(n10716), .ZN(n571) );
  INVX0 U10746 ( .INP(n10717), .ZN(n570) );
  INVX0 U10747 ( .INP(n10718), .ZN(n569) );
  INVX0 U10748 ( .INP(n10719), .ZN(n568) );
  INVX0 U10749 ( .INP(n10720), .ZN(n56) );
  NOR2X0 U10750 ( .IN1(n10721), .IN2(n10722), .QN(n10720) );
  NAND2X0 U10751 ( .IN1(n10723), .IN2(n10724), .QN(n10722) );
  NAND2X0 U10752 ( .IN1(n9949), .IN2(n10725), .QN(n10724) );
  NAND2X0 U10753 ( .IN1(n2152), .IN2(CRC_OUT_9_26), .QN(n10723) );
  NAND2X0 U10754 ( .IN1(n10726), .IN2(n10727), .QN(n10721) );
  INVX0 U10755 ( .INP(n10728), .ZN(n10727) );
  NOR2X0 U10756 ( .IN1(n9925), .IN2(n10729), .QN(n10728) );
  NAND2X0 U10757 ( .IN1(WX492), .IN2(n2339), .QN(n10726) );
  INVX0 U10758 ( .INP(n10730), .ZN(n53) );
  NOR2X0 U10759 ( .IN1(n10731), .IN2(n10732), .QN(n10730) );
  NAND2X0 U10760 ( .IN1(n10733), .IN2(n10734), .QN(n10732) );
  NAND2X0 U10761 ( .IN1(n9949), .IN2(n10735), .QN(n10734) );
  NAND2X0 U10762 ( .IN1(n2152), .IN2(CRC_OUT_9_27), .QN(n10733) );
  NAND2X0 U10763 ( .IN1(n10736), .IN2(n10737), .QN(n10731) );
  INVX0 U10764 ( .INP(n10738), .ZN(n10737) );
  NOR2X0 U10765 ( .IN1(n9925), .IN2(n10739), .QN(n10738) );
  NAND2X0 U10766 ( .IN1(WX490), .IN2(n2339), .QN(n10736) );
  INVX0 U10767 ( .INP(n10740), .ZN(n49) );
  NOR2X0 U10768 ( .IN1(n10741), .IN2(n10742), .QN(n10740) );
  NAND2X0 U10769 ( .IN1(n10743), .IN2(n10744), .QN(n10742) );
  INVX0 U10770 ( .INP(n10745), .ZN(n10744) );
  NOR2X0 U10771 ( .IN1(n10746), .IN2(n9927), .QN(n10745) );
  NAND2X0 U10772 ( .IN1(n2152), .IN2(CRC_OUT_9_28), .QN(n10743) );
  NAND2X0 U10773 ( .IN1(n10747), .IN2(n10748), .QN(n10741) );
  NAND2X0 U10774 ( .IN1(n10749), .IN2(n2153), .QN(n10748) );
  NAND2X0 U10775 ( .IN1(WX488), .IN2(n2339), .QN(n10747) );
  INVX0 U10776 ( .INP(n10750), .ZN(n46) );
  NOR2X0 U10777 ( .IN1(n10751), .IN2(n10752), .QN(n10750) );
  NAND2X0 U10778 ( .IN1(n10753), .IN2(n10754), .QN(n10752) );
  NAND2X0 U10779 ( .IN1(n9950), .IN2(n10755), .QN(n10754) );
  NAND2X0 U10780 ( .IN1(n2152), .IN2(CRC_OUT_9_29), .QN(n10753) );
  NAND2X0 U10781 ( .IN1(n10756), .IN2(n10757), .QN(n10751) );
  INVX0 U10782 ( .INP(n10758), .ZN(n10757) );
  NOR2X0 U10783 ( .IN1(n9925), .IN2(n10759), .QN(n10758) );
  NAND2X0 U10784 ( .IN1(WX486), .IN2(n2339), .QN(n10756) );
  INVX0 U10785 ( .INP(n10760), .ZN(n43) );
  NOR2X0 U10786 ( .IN1(n10761), .IN2(n10762), .QN(n10760) );
  NAND2X0 U10787 ( .IN1(n10763), .IN2(n10764), .QN(n10762) );
  NAND2X0 U10788 ( .IN1(n9950), .IN2(n10765), .QN(n10764) );
  NAND2X0 U10789 ( .IN1(n2152), .IN2(CRC_OUT_9_30), .QN(n10763) );
  NAND2X0 U10790 ( .IN1(n10766), .IN2(n10767), .QN(n10761) );
  INVX0 U10791 ( .INP(n10768), .ZN(n10767) );
  NOR2X0 U10792 ( .IN1(n9925), .IN2(n10769), .QN(n10768) );
  NAND2X0 U10793 ( .IN1(WX484), .IN2(n2339), .QN(n10766) );
  NOR2X0 U10794 ( .IN1(TM1), .IN2(n10234), .QN(n3278) );
  INVX0 U10795 ( .INP(n10770), .ZN(n311) );
  INVX0 U10796 ( .INP(n10771), .ZN(n310) );
  INVX0 U10797 ( .INP(n10772), .ZN(n309) );
  INVX0 U10798 ( .INP(n10773), .ZN(n308) );
  INVX0 U10799 ( .INP(n10774), .ZN(n307) );
  INVX0 U10800 ( .INP(n10775), .ZN(n306) );
  INVX0 U10801 ( .INP(n10776), .ZN(n305) );
  INVX0 U10802 ( .INP(n10777), .ZN(n304) );
  INVX0 U10803 ( .INP(n10778), .ZN(n303) );
  INVX0 U10804 ( .INP(n10779), .ZN(n302) );
  INVX0 U10805 ( .INP(n10780), .ZN(n301) );
  INVX0 U10806 ( .INP(n10781), .ZN(n300) );
  INVX0 U10807 ( .INP(n10782), .ZN(n299) );
  INVX0 U10808 ( .INP(n10783), .ZN(n298) );
  INVX0 U10809 ( .INP(n10784), .ZN(n297) );
  INVX0 U10810 ( .INP(n10785), .ZN(n296) );
  INVX0 U10811 ( .INP(n10786), .ZN(n295) );
  INVX0 U10812 ( .INP(n10787), .ZN(n294) );
  INVX0 U10813 ( .INP(n10788), .ZN(n293) );
  INVX0 U10814 ( .INP(n10789), .ZN(n292) );
  INVX0 U10815 ( .INP(n10790), .ZN(n291) );
  INVX0 U10816 ( .INP(n10791), .ZN(n290) );
  INVX0 U10817 ( .INP(n10792), .ZN(n289) );
  INVX0 U10818 ( .INP(n10793), .ZN(n288) );
  INVX0 U10819 ( .INP(n10794), .ZN(n287) );
  INVX0 U10820 ( .INP(n10795), .ZN(n286) );
  INVX0 U10821 ( .INP(n10796), .ZN(n285) );
  INVX0 U10822 ( .INP(n10797), .ZN(n284) );
  INVX0 U10823 ( .INP(n10798), .ZN(n283) );
  INVX0 U10824 ( .INP(n10799), .ZN(n282) );
  INVX0 U10825 ( .INP(n10800), .ZN(n281) );
  INVX0 U10826 ( .INP(n10801), .ZN(n2072) );
  NOR2X0 U10827 ( .IN1(n10802), .IN2(n10803), .QN(n10801) );
  NAND2X0 U10828 ( .IN1(n10804), .IN2(n10805), .QN(n10803) );
  NAND2X0 U10829 ( .IN1(DATA_0_0), .IN2(n2153), .QN(n10805) );
  NAND2X0 U10830 ( .IN1(n2152), .IN2(CRC_OUT_1_0), .QN(n10804) );
  NAND2X0 U10831 ( .IN1(n10806), .IN2(n10807), .QN(n10802) );
  INVX0 U10832 ( .INP(n10808), .ZN(n10807) );
  NOR2X0 U10833 ( .IN1(n10563), .IN2(n10809), .QN(n10808) );
  NAND2X0 U10834 ( .IN1(n2073), .IN2(n2339), .QN(n10806) );
  NOR2X0 U10835 ( .IN1(n10311), .IN2(n9872), .QN(n2073) );
  INVX0 U10836 ( .INP(n10810), .ZN(n2070) );
  NOR2X0 U10837 ( .IN1(n10811), .IN2(n10812), .QN(n10810) );
  NAND2X0 U10838 ( .IN1(n10813), .IN2(n10814), .QN(n10812) );
  NAND2X0 U10839 ( .IN1(DATA_0_1), .IN2(n2153), .QN(n10814) );
  NAND2X0 U10840 ( .IN1(n2152), .IN2(CRC_OUT_1_1), .QN(n10813) );
  NAND2X0 U10841 ( .IN1(n10815), .IN2(n10816), .QN(n10811) );
  INVX0 U10842 ( .INP(n10817), .ZN(n10816) );
  NOR2X0 U10843 ( .IN1(n9945), .IN2(n10818), .QN(n10817) );
  NAND2X0 U10844 ( .IN1(n2071), .IN2(n2339), .QN(n10815) );
  NOR2X0 U10845 ( .IN1(n10326), .IN2(n9873), .QN(n2071) );
  INVX0 U10846 ( .INP(n10819), .ZN(n2068) );
  NOR2X0 U10847 ( .IN1(n10820), .IN2(n10821), .QN(n10819) );
  NAND2X0 U10848 ( .IN1(n10822), .IN2(n10823), .QN(n10821) );
  NAND2X0 U10849 ( .IN1(DATA_0_2), .IN2(n2153), .QN(n10823) );
  NAND2X0 U10850 ( .IN1(n2152), .IN2(CRC_OUT_1_2), .QN(n10822) );
  NAND2X0 U10851 ( .IN1(n10824), .IN2(n10825), .QN(n10820) );
  NAND2X0 U10852 ( .IN1(n10826), .IN2(n9952), .QN(n10825) );
  NAND2X0 U10853 ( .IN1(n2069), .IN2(n2339), .QN(n10824) );
  NOR2X0 U10854 ( .IN1(n10319), .IN2(n9874), .QN(n2069) );
  INVX0 U10855 ( .INP(n10827), .ZN(n2066) );
  NOR2X0 U10856 ( .IN1(n10828), .IN2(n10829), .QN(n10827) );
  NAND2X0 U10857 ( .IN1(n10830), .IN2(n10831), .QN(n10829) );
  NAND2X0 U10858 ( .IN1(DATA_0_3), .IN2(n2153), .QN(n10831) );
  NAND2X0 U10859 ( .IN1(n2152), .IN2(CRC_OUT_1_3), .QN(n10830) );
  NAND2X0 U10860 ( .IN1(n10832), .IN2(n10833), .QN(n10828) );
  INVX0 U10861 ( .INP(n10834), .ZN(n10833) );
  NOR2X0 U10862 ( .IN1(n9945), .IN2(n10835), .QN(n10834) );
  NAND2X0 U10863 ( .IN1(n2067), .IN2(n2339), .QN(n10832) );
  NOR2X0 U10864 ( .IN1(n10319), .IN2(n9875), .QN(n2067) );
  INVX0 U10865 ( .INP(n10836), .ZN(n2064) );
  NOR2X0 U10866 ( .IN1(n10837), .IN2(n10838), .QN(n10836) );
  NAND2X0 U10867 ( .IN1(n10839), .IN2(n10840), .QN(n10838) );
  NAND2X0 U10868 ( .IN1(DATA_0_4), .IN2(n2153), .QN(n10840) );
  NAND2X0 U10869 ( .IN1(n2152), .IN2(CRC_OUT_1_4), .QN(n10839) );
  NAND2X0 U10870 ( .IN1(n10841), .IN2(n10842), .QN(n10837) );
  NAND2X0 U10871 ( .IN1(n10843), .IN2(n9952), .QN(n10842) );
  NAND2X0 U10872 ( .IN1(n2065), .IN2(n2339), .QN(n10841) );
  NOR2X0 U10873 ( .IN1(n10319), .IN2(n9876), .QN(n2065) );
  INVX0 U10874 ( .INP(n10844), .ZN(n2062) );
  NOR2X0 U10875 ( .IN1(n10845), .IN2(n10846), .QN(n10844) );
  NAND2X0 U10876 ( .IN1(n10847), .IN2(n10848), .QN(n10846) );
  NAND2X0 U10877 ( .IN1(DATA_0_5), .IN2(n2153), .QN(n10848) );
  NAND2X0 U10878 ( .IN1(n2152), .IN2(CRC_OUT_1_5), .QN(n10847) );
  NAND2X0 U10879 ( .IN1(n10849), .IN2(n10850), .QN(n10845) );
  INVX0 U10880 ( .INP(n10851), .ZN(n10850) );
  NOR2X0 U10881 ( .IN1(n9945), .IN2(n10852), .QN(n10851) );
  NAND2X0 U10882 ( .IN1(n2063), .IN2(n2339), .QN(n10849) );
  NOR2X0 U10883 ( .IN1(n10319), .IN2(n9877), .QN(n2063) );
  INVX0 U10884 ( .INP(n10853), .ZN(n2060) );
  NOR2X0 U10885 ( .IN1(n10854), .IN2(n10855), .QN(n10853) );
  NAND2X0 U10886 ( .IN1(n10856), .IN2(n10857), .QN(n10855) );
  NAND2X0 U10887 ( .IN1(DATA_0_6), .IN2(n2153), .QN(n10857) );
  NAND2X0 U10888 ( .IN1(n2152), .IN2(CRC_OUT_1_6), .QN(n10856) );
  NAND2X0 U10889 ( .IN1(n10858), .IN2(n10859), .QN(n10854) );
  NAND2X0 U10890 ( .IN1(n10860), .IN2(n9952), .QN(n10859) );
  NAND2X0 U10891 ( .IN1(n2061), .IN2(n2339), .QN(n10858) );
  NOR2X0 U10892 ( .IN1(n10319), .IN2(n9878), .QN(n2061) );
  INVX0 U10893 ( .INP(n10861), .ZN(n2058) );
  NOR2X0 U10894 ( .IN1(n10862), .IN2(n10863), .QN(n10861) );
  NAND2X0 U10895 ( .IN1(n10864), .IN2(n10865), .QN(n10863) );
  NAND2X0 U10896 ( .IN1(DATA_0_7), .IN2(n2153), .QN(n10865) );
  NAND2X0 U10897 ( .IN1(n2152), .IN2(CRC_OUT_1_7), .QN(n10864) );
  NAND2X0 U10898 ( .IN1(n10866), .IN2(n10867), .QN(n10862) );
  INVX0 U10899 ( .INP(n10868), .ZN(n10867) );
  NOR2X0 U10900 ( .IN1(n9945), .IN2(n10869), .QN(n10868) );
  NAND2X0 U10901 ( .IN1(n2059), .IN2(n2339), .QN(n10866) );
  NOR2X0 U10902 ( .IN1(n10319), .IN2(n9879), .QN(n2059) );
  INVX0 U10903 ( .INP(n10870), .ZN(n2056) );
  NOR2X0 U10904 ( .IN1(n10871), .IN2(n10872), .QN(n10870) );
  NAND2X0 U10905 ( .IN1(n10873), .IN2(n10874), .QN(n10872) );
  NAND2X0 U10906 ( .IN1(DATA_0_8), .IN2(n2153), .QN(n10874) );
  NAND2X0 U10907 ( .IN1(n2152), .IN2(CRC_OUT_1_8), .QN(n10873) );
  NAND2X0 U10908 ( .IN1(n10875), .IN2(n10876), .QN(n10871) );
  NAND2X0 U10909 ( .IN1(n10877), .IN2(n9952), .QN(n10876) );
  NAND2X0 U10910 ( .IN1(n2057), .IN2(n2339), .QN(n10875) );
  NOR2X0 U10911 ( .IN1(n10319), .IN2(n9880), .QN(n2057) );
  INVX0 U10912 ( .INP(n10878), .ZN(n2054) );
  NOR2X0 U10913 ( .IN1(n10879), .IN2(n10880), .QN(n10878) );
  NAND2X0 U10914 ( .IN1(n10881), .IN2(n10882), .QN(n10880) );
  NAND2X0 U10915 ( .IN1(DATA_0_9), .IN2(n2153), .QN(n10882) );
  NAND2X0 U10916 ( .IN1(n2152), .IN2(CRC_OUT_1_9), .QN(n10881) );
  NAND2X0 U10917 ( .IN1(n10883), .IN2(n10884), .QN(n10879) );
  INVX0 U10918 ( .INP(n10885), .ZN(n10884) );
  NOR2X0 U10919 ( .IN1(n9945), .IN2(n10886), .QN(n10885) );
  NAND2X0 U10920 ( .IN1(n2055), .IN2(n2339), .QN(n10883) );
  NOR2X0 U10921 ( .IN1(n10319), .IN2(n9881), .QN(n2055) );
  INVX0 U10922 ( .INP(n10887), .ZN(n2052) );
  NOR2X0 U10923 ( .IN1(n10888), .IN2(n10889), .QN(n10887) );
  NAND2X0 U10924 ( .IN1(n10890), .IN2(n10891), .QN(n10889) );
  NAND2X0 U10925 ( .IN1(DATA_0_10), .IN2(n2153), .QN(n10891) );
  NAND2X0 U10926 ( .IN1(n2152), .IN2(CRC_OUT_1_10), .QN(n10890) );
  NAND2X0 U10927 ( .IN1(n10892), .IN2(n10893), .QN(n10888) );
  INVX0 U10928 ( .INP(n10894), .ZN(n10893) );
  NOR2X0 U10929 ( .IN1(n9945), .IN2(n10895), .QN(n10894) );
  NAND2X0 U10930 ( .IN1(n2053), .IN2(n2339), .QN(n10892) );
  NOR2X0 U10931 ( .IN1(n9901), .IN2(n10234), .QN(n2053) );
  INVX0 U10932 ( .INP(n10896), .ZN(n2050) );
  NOR2X0 U10933 ( .IN1(n10897), .IN2(n10898), .QN(n10896) );
  NAND2X0 U10934 ( .IN1(n10899), .IN2(n10900), .QN(n10898) );
  NAND2X0 U10935 ( .IN1(DATA_0_11), .IN2(n2153), .QN(n10900) );
  NAND2X0 U10936 ( .IN1(n2152), .IN2(CRC_OUT_1_11), .QN(n10899) );
  NAND2X0 U10937 ( .IN1(n10901), .IN2(n10902), .QN(n10897) );
  INVX0 U10938 ( .INP(n10903), .ZN(n10902) );
  NOR2X0 U10939 ( .IN1(n9945), .IN2(n10904), .QN(n10903) );
  NAND2X0 U10940 ( .IN1(n2051), .IN2(n2339), .QN(n10901) );
  NOR2X0 U10941 ( .IN1(n10319), .IN2(n9882), .QN(n2051) );
  INVX0 U10942 ( .INP(n10905), .ZN(n2048) );
  NOR2X0 U10943 ( .IN1(n10906), .IN2(n10907), .QN(n10905) );
  NAND2X0 U10944 ( .IN1(n10908), .IN2(n10909), .QN(n10907) );
  NAND2X0 U10945 ( .IN1(DATA_0_12), .IN2(n2153), .QN(n10909) );
  NAND2X0 U10946 ( .IN1(n2152), .IN2(CRC_OUT_1_12), .QN(n10908) );
  NAND2X0 U10947 ( .IN1(n10910), .IN2(n10911), .QN(n10906) );
  INVX0 U10948 ( .INP(n10912), .ZN(n10911) );
  NOR2X0 U10949 ( .IN1(n9945), .IN2(n10913), .QN(n10912) );
  NAND2X0 U10950 ( .IN1(n2049), .IN2(n2339), .QN(n10910) );
  NOR2X0 U10951 ( .IN1(n10319), .IN2(n9883), .QN(n2049) );
  INVX0 U10952 ( .INP(n10914), .ZN(n2046) );
  NOR2X0 U10953 ( .IN1(n10915), .IN2(n10916), .QN(n10914) );
  NAND2X0 U10954 ( .IN1(n10917), .IN2(n10918), .QN(n10916) );
  NAND2X0 U10955 ( .IN1(DATA_0_13), .IN2(n2153), .QN(n10918) );
  NAND2X0 U10956 ( .IN1(n2152), .IN2(CRC_OUT_1_13), .QN(n10917) );
  NAND2X0 U10957 ( .IN1(n10919), .IN2(n10920), .QN(n10915) );
  INVX0 U10958 ( .INP(n10921), .ZN(n10920) );
  NOR2X0 U10959 ( .IN1(n9945), .IN2(n10922), .QN(n10921) );
  NAND2X0 U10960 ( .IN1(n2047), .IN2(n2339), .QN(n10919) );
  NOR2X0 U10961 ( .IN1(n10319), .IN2(n9884), .QN(n2047) );
  INVX0 U10962 ( .INP(n10923), .ZN(n2044) );
  NOR2X0 U10963 ( .IN1(n10924), .IN2(n10925), .QN(n10923) );
  NAND2X0 U10964 ( .IN1(n10926), .IN2(n10927), .QN(n10925) );
  NAND2X0 U10965 ( .IN1(DATA_0_14), .IN2(n2153), .QN(n10927) );
  NAND2X0 U10966 ( .IN1(test_so99), .IN2(n2152), .QN(n10926) );
  NAND2X0 U10967 ( .IN1(n10928), .IN2(n10929), .QN(n10924) );
  INVX0 U10968 ( .INP(n10930), .ZN(n10929) );
  NOR2X0 U10969 ( .IN1(n9945), .IN2(n10931), .QN(n10930) );
  NAND2X0 U10970 ( .IN1(n2045), .IN2(n2339), .QN(n10928) );
  NOR2X0 U10971 ( .IN1(n10319), .IN2(n9885), .QN(n2045) );
  INVX0 U10972 ( .INP(n10932), .ZN(n2042) );
  NOR2X0 U10973 ( .IN1(n10933), .IN2(n10934), .QN(n10932) );
  NAND2X0 U10974 ( .IN1(n10935), .IN2(n10936), .QN(n10934) );
  NAND2X0 U10975 ( .IN1(DATA_0_15), .IN2(n2153), .QN(n10936) );
  NAND2X0 U10976 ( .IN1(n2152), .IN2(CRC_OUT_1_15), .QN(n10935) );
  NAND2X0 U10977 ( .IN1(n10937), .IN2(n10938), .QN(n10933) );
  INVX0 U10978 ( .INP(n10939), .ZN(n10938) );
  NOR2X0 U10979 ( .IN1(n9945), .IN2(n10940), .QN(n10939) );
  NAND2X0 U10980 ( .IN1(n2043), .IN2(n2339), .QN(n10937) );
  NOR2X0 U10981 ( .IN1(n10320), .IN2(n9886), .QN(n2043) );
  INVX0 U10982 ( .INP(n10941), .ZN(n2040) );
  NOR2X0 U10983 ( .IN1(n10942), .IN2(n10943), .QN(n10941) );
  NAND2X0 U10984 ( .IN1(n10944), .IN2(n10945), .QN(n10943) );
  NAND2X0 U10985 ( .IN1(DATA_0_16), .IN2(n2153), .QN(n10945) );
  NAND2X0 U10986 ( .IN1(n2152), .IN2(CRC_OUT_1_16), .QN(n10944) );
  NAND2X0 U10987 ( .IN1(n10946), .IN2(n10947), .QN(n10942) );
  INVX0 U10988 ( .INP(n10948), .ZN(n10947) );
  NOR2X0 U10989 ( .IN1(n9945), .IN2(n10949), .QN(n10948) );
  NAND2X0 U10990 ( .IN1(n2041), .IN2(n2339), .QN(n10946) );
  NOR2X0 U10991 ( .IN1(n10320), .IN2(n9887), .QN(n2041) );
  INVX0 U10992 ( .INP(n10950), .ZN(n2038) );
  NOR2X0 U10993 ( .IN1(n10951), .IN2(n10952), .QN(n10950) );
  NAND2X0 U10994 ( .IN1(n10953), .IN2(n10954), .QN(n10952) );
  NAND2X0 U10995 ( .IN1(DATA_0_17), .IN2(n2153), .QN(n10954) );
  NAND2X0 U10996 ( .IN1(n2152), .IN2(CRC_OUT_1_17), .QN(n10953) );
  NAND2X0 U10997 ( .IN1(n10955), .IN2(n10956), .QN(n10951) );
  INVX0 U10998 ( .INP(n10957), .ZN(n10956) );
  NOR2X0 U10999 ( .IN1(n9945), .IN2(n10958), .QN(n10957) );
  NAND2X0 U11000 ( .IN1(n2039), .IN2(n2339), .QN(n10955) );
  NOR2X0 U11001 ( .IN1(n10320), .IN2(n9888), .QN(n2039) );
  INVX0 U11002 ( .INP(n10959), .ZN(n2036) );
  NOR2X0 U11003 ( .IN1(n10960), .IN2(n10961), .QN(n10959) );
  NAND2X0 U11004 ( .IN1(n10962), .IN2(n10963), .QN(n10961) );
  NAND2X0 U11005 ( .IN1(DATA_0_18), .IN2(n2153), .QN(n10963) );
  NAND2X0 U11006 ( .IN1(n2152), .IN2(CRC_OUT_1_18), .QN(n10962) );
  NAND2X0 U11007 ( .IN1(n10964), .IN2(n10965), .QN(n10960) );
  INVX0 U11008 ( .INP(n10966), .ZN(n10965) );
  NOR2X0 U11009 ( .IN1(n9944), .IN2(n10967), .QN(n10966) );
  NAND2X0 U11010 ( .IN1(n2037), .IN2(n2339), .QN(n10964) );
  NOR2X0 U11011 ( .IN1(n10320), .IN2(n9889), .QN(n2037) );
  INVX0 U11012 ( .INP(n10968), .ZN(n2034) );
  NOR2X0 U11013 ( .IN1(n10969), .IN2(n10970), .QN(n10968) );
  NAND2X0 U11014 ( .IN1(n10971), .IN2(n10972), .QN(n10970) );
  NAND2X0 U11015 ( .IN1(DATA_0_19), .IN2(n2153), .QN(n10972) );
  NAND2X0 U11016 ( .IN1(n2152), .IN2(CRC_OUT_1_19), .QN(n10971) );
  NAND2X0 U11017 ( .IN1(n10973), .IN2(n10974), .QN(n10969) );
  NAND2X0 U11018 ( .IN1(n10975), .IN2(n9952), .QN(n10974) );
  NAND2X0 U11019 ( .IN1(n2035), .IN2(n2339), .QN(n10973) );
  NOR2X0 U11020 ( .IN1(n10320), .IN2(n9890), .QN(n2035) );
  INVX0 U11021 ( .INP(n10976), .ZN(n2032) );
  NOR2X0 U11022 ( .IN1(n10977), .IN2(n10978), .QN(n10976) );
  NAND2X0 U11023 ( .IN1(n10979), .IN2(n10980), .QN(n10978) );
  NAND2X0 U11024 ( .IN1(DATA_0_20), .IN2(n2153), .QN(n10980) );
  NAND2X0 U11025 ( .IN1(n2152), .IN2(CRC_OUT_1_20), .QN(n10979) );
  NAND2X0 U11026 ( .IN1(n10981), .IN2(n10982), .QN(n10977) );
  INVX0 U11027 ( .INP(n10983), .ZN(n10982) );
  NOR2X0 U11028 ( .IN1(n9944), .IN2(n10984), .QN(n10983) );
  NAND2X0 U11029 ( .IN1(n2033), .IN2(n2339), .QN(n10981) );
  NOR2X0 U11030 ( .IN1(n10320), .IN2(n9891), .QN(n2033) );
  INVX0 U11031 ( .INP(n10985), .ZN(n2030) );
  NOR2X0 U11032 ( .IN1(n10986), .IN2(n10987), .QN(n10985) );
  NAND2X0 U11033 ( .IN1(n10988), .IN2(n10989), .QN(n10987) );
  NAND2X0 U11034 ( .IN1(DATA_0_21), .IN2(n2153), .QN(n10989) );
  NAND2X0 U11035 ( .IN1(n2152), .IN2(CRC_OUT_1_21), .QN(n10988) );
  NAND2X0 U11036 ( .IN1(n10990), .IN2(n10991), .QN(n10986) );
  NAND2X0 U11037 ( .IN1(n10992), .IN2(n9952), .QN(n10991) );
  NAND2X0 U11038 ( .IN1(n2031), .IN2(n2339), .QN(n10990) );
  NOR2X0 U11039 ( .IN1(n10320), .IN2(n9892), .QN(n2031) );
  INVX0 U11040 ( .INP(n10993), .ZN(n2028) );
  NOR2X0 U11041 ( .IN1(n10994), .IN2(n10995), .QN(n10993) );
  NAND2X0 U11042 ( .IN1(n10996), .IN2(n10997), .QN(n10995) );
  NAND2X0 U11043 ( .IN1(DATA_0_22), .IN2(n2153), .QN(n10997) );
  NAND2X0 U11044 ( .IN1(n2152), .IN2(CRC_OUT_1_22), .QN(n10996) );
  NAND2X0 U11045 ( .IN1(n10998), .IN2(n10999), .QN(n10994) );
  INVX0 U11046 ( .INP(n11000), .ZN(n10999) );
  NOR2X0 U11047 ( .IN1(n9944), .IN2(n11001), .QN(n11000) );
  NAND2X0 U11048 ( .IN1(n2029), .IN2(n2339), .QN(n10998) );
  NOR2X0 U11049 ( .IN1(n10320), .IN2(n9893), .QN(n2029) );
  INVX0 U11050 ( .INP(n11002), .ZN(n2026) );
  NOR2X0 U11051 ( .IN1(n11003), .IN2(n11004), .QN(n11002) );
  NAND2X0 U11052 ( .IN1(n11005), .IN2(n11006), .QN(n11004) );
  NAND2X0 U11053 ( .IN1(DATA_0_23), .IN2(n2153), .QN(n11006) );
  NAND2X0 U11054 ( .IN1(n2152), .IN2(CRC_OUT_1_23), .QN(n11005) );
  NAND2X0 U11055 ( .IN1(n11007), .IN2(n11008), .QN(n11003) );
  NAND2X0 U11056 ( .IN1(n11009), .IN2(n9952), .QN(n11008) );
  NAND2X0 U11057 ( .IN1(n2027), .IN2(n2339), .QN(n11007) );
  NOR2X0 U11058 ( .IN1(n10320), .IN2(n9894), .QN(n2027) );
  INVX0 U11059 ( .INP(n11010), .ZN(n2024) );
  NOR2X0 U11060 ( .IN1(n11011), .IN2(n11012), .QN(n11010) );
  NAND2X0 U11061 ( .IN1(n11013), .IN2(n11014), .QN(n11012) );
  NAND2X0 U11062 ( .IN1(DATA_0_24), .IN2(n2153), .QN(n11014) );
  NAND2X0 U11063 ( .IN1(n2152), .IN2(CRC_OUT_1_24), .QN(n11013) );
  NAND2X0 U11064 ( .IN1(n11015), .IN2(n11016), .QN(n11011) );
  INVX0 U11065 ( .INP(n11017), .ZN(n11016) );
  NOR2X0 U11066 ( .IN1(n9944), .IN2(n11018), .QN(n11017) );
  NAND2X0 U11067 ( .IN1(n2025), .IN2(n2339), .QN(n11015) );
  NOR2X0 U11068 ( .IN1(n10320), .IN2(n9895), .QN(n2025) );
  INVX0 U11069 ( .INP(n11019), .ZN(n2022) );
  NOR2X0 U11070 ( .IN1(n11020), .IN2(n11021), .QN(n11019) );
  NAND2X0 U11071 ( .IN1(n11022), .IN2(n11023), .QN(n11021) );
  NAND2X0 U11072 ( .IN1(DATA_0_25), .IN2(n2153), .QN(n11023) );
  NAND2X0 U11073 ( .IN1(n2152), .IN2(CRC_OUT_1_25), .QN(n11022) );
  NAND2X0 U11074 ( .IN1(n11024), .IN2(n11025), .QN(n11020) );
  NAND2X0 U11075 ( .IN1(n11026), .IN2(n9952), .QN(n11025) );
  NAND2X0 U11076 ( .IN1(n2023), .IN2(n2339), .QN(n11024) );
  NOR2X0 U11077 ( .IN1(n10320), .IN2(n9896), .QN(n2023) );
  INVX0 U11078 ( .INP(n11027), .ZN(n2020) );
  NOR2X0 U11079 ( .IN1(n11028), .IN2(n11029), .QN(n11027) );
  NAND2X0 U11080 ( .IN1(n11030), .IN2(n11031), .QN(n11029) );
  NAND2X0 U11081 ( .IN1(DATA_0_26), .IN2(n2153), .QN(n11031) );
  NAND2X0 U11082 ( .IN1(n2152), .IN2(CRC_OUT_1_26), .QN(n11030) );
  NAND2X0 U11083 ( .IN1(n11032), .IN2(n11033), .QN(n11028) );
  INVX0 U11084 ( .INP(n11034), .ZN(n11033) );
  NOR2X0 U11085 ( .IN1(n9944), .IN2(n11035), .QN(n11034) );
  NAND2X0 U11086 ( .IN1(n2021), .IN2(n2339), .QN(n11032) );
  NOR2X0 U11087 ( .IN1(n10320), .IN2(n9897), .QN(n2021) );
  INVX0 U11088 ( .INP(n11036), .ZN(n2018) );
  NOR2X0 U11089 ( .IN1(n11037), .IN2(n11038), .QN(n11036) );
  NAND2X0 U11090 ( .IN1(n11039), .IN2(n11040), .QN(n11038) );
  NAND2X0 U11091 ( .IN1(DATA_0_27), .IN2(n2153), .QN(n11040) );
  NAND2X0 U11092 ( .IN1(n2152), .IN2(CRC_OUT_1_27), .QN(n11039) );
  NAND2X0 U11093 ( .IN1(n11041), .IN2(n11042), .QN(n11037) );
  INVX0 U11094 ( .INP(n11043), .ZN(n11042) );
  NOR2X0 U11095 ( .IN1(n9944), .IN2(n11044), .QN(n11043) );
  NAND2X0 U11096 ( .IN1(n2019), .IN2(n2339), .QN(n11041) );
  NOR2X0 U11097 ( .IN1(n9902), .IN2(n10234), .QN(n2019) );
  INVX0 U11098 ( .INP(n11045), .ZN(n2016) );
  NOR2X0 U11099 ( .IN1(n11046), .IN2(n11047), .QN(n11045) );
  NAND2X0 U11100 ( .IN1(n11048), .IN2(n11049), .QN(n11047) );
  NAND2X0 U11101 ( .IN1(DATA_0_28), .IN2(n2153), .QN(n11049) );
  NAND2X0 U11102 ( .IN1(n2152), .IN2(CRC_OUT_1_28), .QN(n11048) );
  NAND2X0 U11103 ( .IN1(n11050), .IN2(n11051), .QN(n11046) );
  INVX0 U11104 ( .INP(n11052), .ZN(n11051) );
  NOR2X0 U11105 ( .IN1(n9944), .IN2(n11053), .QN(n11052) );
  NAND2X0 U11106 ( .IN1(n2017), .IN2(n2339), .QN(n11050) );
  NOR2X0 U11107 ( .IN1(n10320), .IN2(n9898), .QN(n2017) );
  INVX0 U11108 ( .INP(n11054), .ZN(n2014) );
  NOR2X0 U11109 ( .IN1(n11055), .IN2(n11056), .QN(n11054) );
  NAND2X0 U11110 ( .IN1(n11057), .IN2(n11058), .QN(n11056) );
  NAND2X0 U11111 ( .IN1(DATA_0_29), .IN2(n2153), .QN(n11058) );
  NAND2X0 U11112 ( .IN1(n2152), .IN2(CRC_OUT_1_29), .QN(n11057) );
  NAND2X0 U11113 ( .IN1(n11059), .IN2(n11060), .QN(n11055) );
  INVX0 U11114 ( .INP(n11061), .ZN(n11060) );
  NOR2X0 U11115 ( .IN1(n9944), .IN2(n11062), .QN(n11061) );
  NAND2X0 U11116 ( .IN1(n2015), .IN2(n2339), .QN(n11059) );
  NOR2X0 U11117 ( .IN1(n10321), .IN2(n9899), .QN(n2015) );
  INVX0 U11118 ( .INP(n11063), .ZN(n2012) );
  NOR2X0 U11119 ( .IN1(n11064), .IN2(n11065), .QN(n11063) );
  NAND2X0 U11120 ( .IN1(n11066), .IN2(n11067), .QN(n11065) );
  NAND2X0 U11121 ( .IN1(DATA_0_30), .IN2(n2153), .QN(n11067) );
  NAND2X0 U11122 ( .IN1(n2152), .IN2(CRC_OUT_1_30), .QN(n11066) );
  NAND2X0 U11123 ( .IN1(n11068), .IN2(n11069), .QN(n11064) );
  INVX0 U11124 ( .INP(n11070), .ZN(n11069) );
  NOR2X0 U11125 ( .IN1(n9944), .IN2(n11071), .QN(n11070) );
  NAND2X0 U11126 ( .IN1(n2013), .IN2(n2339), .QN(n11068) );
  NOR2X0 U11127 ( .IN1(n10321), .IN2(n9900), .QN(n2013) );
  INVX0 U11128 ( .INP(n11072), .ZN(n2010) );
  NOR2X0 U11129 ( .IN1(n11073), .IN2(n11074), .QN(n11072) );
  NAND2X0 U11130 ( .IN1(n11075), .IN2(n11076), .QN(n11074) );
  NAND2X0 U11131 ( .IN1(test_so100), .IN2(n2152), .QN(n11076) );
  NAND2X0 U11132 ( .IN1(n2245), .IN2(WX10829), .QN(n11075) );
  NAND2X0 U11133 ( .IN1(n11077), .IN2(n11078), .QN(n11073) );
  INVX0 U11134 ( .INP(n11079), .ZN(n11078) );
  NOR2X0 U11135 ( .IN1(n9944), .IN2(n11080), .QN(n11079) );
  NAND2X0 U11136 ( .IN1(DATA_0_31), .IN2(n2153), .QN(n11077) );
  INVX0 U11137 ( .INP(n11081), .ZN(n1801) );
  INVX0 U11138 ( .INP(n11082), .ZN(n1800) );
  INVX0 U11139 ( .INP(n11083), .ZN(n1799) );
  INVX0 U11140 ( .INP(n11084), .ZN(n1798) );
  INVX0 U11141 ( .INP(n11085), .ZN(n1797) );
  INVX0 U11142 ( .INP(n11086), .ZN(n1796) );
  INVX0 U11143 ( .INP(n11087), .ZN(n1795) );
  INVX0 U11144 ( .INP(n11088), .ZN(n1794) );
  INVX0 U11145 ( .INP(n11089), .ZN(n1793) );
  INVX0 U11146 ( .INP(n11090), .ZN(n1792) );
  INVX0 U11147 ( .INP(n11091), .ZN(n1791) );
  INVX0 U11148 ( .INP(n11092), .ZN(n1790) );
  INVX0 U11149 ( .INP(n11093), .ZN(n1789) );
  INVX0 U11150 ( .INP(n11094), .ZN(n1788) );
  INVX0 U11151 ( .INP(n11095), .ZN(n1787) );
  INVX0 U11152 ( .INP(n11096), .ZN(n1786) );
  INVX0 U11153 ( .INP(n11097), .ZN(n1785) );
  INVX0 U11154 ( .INP(n11098), .ZN(n1784) );
  INVX0 U11155 ( .INP(n11099), .ZN(n1783) );
  INVX0 U11156 ( .INP(n11100), .ZN(n1782) );
  INVX0 U11157 ( .INP(n11101), .ZN(n1781) );
  INVX0 U11158 ( .INP(n11102), .ZN(n1780) );
  INVX0 U11159 ( .INP(n11103), .ZN(n1779) );
  INVX0 U11160 ( .INP(n11104), .ZN(n1778) );
  INVX0 U11161 ( .INP(n11105), .ZN(n1777) );
  INVX0 U11162 ( .INP(n11106), .ZN(n1776) );
  INVX0 U11163 ( .INP(n11107), .ZN(n1775) );
  INVX0 U11164 ( .INP(n11108), .ZN(n1774) );
  INVX0 U11165 ( .INP(n11109), .ZN(n1773) );
  INVX0 U11166 ( .INP(n11110), .ZN(n1772) );
  INVX0 U11167 ( .INP(n11111), .ZN(n1771) );
  INVX0 U11168 ( .INP(n11112), .ZN(n1560) );
  INVX0 U11169 ( .INP(n11113), .ZN(n1559) );
  INVX0 U11170 ( .INP(n11114), .ZN(n1558) );
  INVX0 U11171 ( .INP(n11115), .ZN(n1557) );
  INVX0 U11172 ( .INP(n11116), .ZN(n1556) );
  INVX0 U11173 ( .INP(n11117), .ZN(n1555) );
  INVX0 U11174 ( .INP(n11118), .ZN(n1554) );
  INVX0 U11175 ( .INP(n11119), .ZN(n1553) );
  INVX0 U11176 ( .INP(n11120), .ZN(n1552) );
  INVX0 U11177 ( .INP(n11121), .ZN(n1551) );
  INVX0 U11178 ( .INP(n11122), .ZN(n1550) );
  INVX0 U11179 ( .INP(n11123), .ZN(n1549) );
  INVX0 U11180 ( .INP(n11124), .ZN(n1548) );
  INVX0 U11181 ( .INP(n11125), .ZN(n1547) );
  INVX0 U11182 ( .INP(n11126), .ZN(n1546) );
  INVX0 U11183 ( .INP(n11127), .ZN(n1545) );
  INVX0 U11184 ( .INP(n11128), .ZN(n1544) );
  INVX0 U11185 ( .INP(n11129), .ZN(n1543) );
  INVX0 U11186 ( .INP(n11130), .ZN(n1542) );
  INVX0 U11187 ( .INP(n11131), .ZN(n1541) );
  INVX0 U11188 ( .INP(n11132), .ZN(n1540) );
  INVX0 U11189 ( .INP(n11133), .ZN(n1539) );
  INVX0 U11190 ( .INP(n11134), .ZN(n1538) );
  INVX0 U11191 ( .INP(n11135), .ZN(n1537) );
  INVX0 U11192 ( .INP(n11136), .ZN(n1536) );
  INVX0 U11193 ( .INP(n11137), .ZN(n1535) );
  INVX0 U11194 ( .INP(n11138), .ZN(n1534) );
  INVX0 U11195 ( .INP(n11139), .ZN(n1533) );
  INVX0 U11196 ( .INP(n11140), .ZN(n1532) );
  INVX0 U11197 ( .INP(n11141), .ZN(n1531) );
  INVX0 U11198 ( .INP(n11142), .ZN(n1530) );
  INVX0 U11199 ( .INP(n11143), .ZN(n135) );
  NOR2X0 U11200 ( .IN1(n11144), .IN2(n11145), .QN(n11143) );
  NAND2X0 U11201 ( .IN1(n11146), .IN2(n11147), .QN(n11145) );
  NAND2X0 U11202 ( .IN1(n9950), .IN2(n11148), .QN(n11147) );
  NAND2X0 U11203 ( .IN1(n2152), .IN2(CRC_OUT_9_0), .QN(n11146) );
  NAND2X0 U11204 ( .IN1(n11149), .IN2(n11150), .QN(n11144) );
  NAND2X0 U11205 ( .IN1(n11151), .IN2(n2153), .QN(n11150) );
  NAND2X0 U11206 ( .IN1(WX544), .IN2(n2339), .QN(n11149) );
  INVX0 U11207 ( .INP(n11152), .ZN(n1320) );
  INVX0 U11208 ( .INP(n11153), .ZN(n132) );
  NOR2X0 U11209 ( .IN1(n11154), .IN2(n11155), .QN(n11153) );
  NAND2X0 U11210 ( .IN1(n11156), .IN2(n11157), .QN(n11155) );
  NAND2X0 U11211 ( .IN1(n9950), .IN2(n11158), .QN(n11157) );
  NAND2X0 U11212 ( .IN1(test_so9), .IN2(n2152), .QN(n11156) );
  NAND2X0 U11213 ( .IN1(n11159), .IN2(n11160), .QN(n11154) );
  INVX0 U11214 ( .INP(n11161), .ZN(n11160) );
  NOR2X0 U11215 ( .IN1(n9925), .IN2(n11162), .QN(n11161) );
  NAND2X0 U11216 ( .IN1(WX542), .IN2(n2339), .QN(n11159) );
  INVX0 U11217 ( .INP(n11163), .ZN(n1319) );
  INVX0 U11218 ( .INP(n11164), .ZN(n1318) );
  INVX0 U11219 ( .INP(n11165), .ZN(n1317) );
  INVX0 U11220 ( .INP(n11166), .ZN(n1316) );
  INVX0 U11221 ( .INP(n11167), .ZN(n1315) );
  INVX0 U11222 ( .INP(n11168), .ZN(n1314) );
  INVX0 U11223 ( .INP(n11169), .ZN(n1313) );
  INVX0 U11224 ( .INP(n11170), .ZN(n1312) );
  INVX0 U11225 ( .INP(n11171), .ZN(n1311) );
  INVX0 U11226 ( .INP(n11172), .ZN(n1310) );
  INVX0 U11227 ( .INP(n11173), .ZN(n1309) );
  INVX0 U11228 ( .INP(n11174), .ZN(n1308) );
  INVX0 U11229 ( .INP(n11175), .ZN(n1307) );
  INVX0 U11230 ( .INP(n11176), .ZN(n1306) );
  INVX0 U11231 ( .INP(n11177), .ZN(n1305) );
  INVX0 U11232 ( .INP(n11178), .ZN(n1304) );
  INVX0 U11233 ( .INP(n11179), .ZN(n1303) );
  INVX0 U11234 ( .INP(n11180), .ZN(n1302) );
  INVX0 U11235 ( .INP(n11181), .ZN(n1301) );
  INVX0 U11236 ( .INP(n11182), .ZN(n1300) );
  INVX0 U11237 ( .INP(n11183), .ZN(n1299) );
  INVX0 U11238 ( .INP(n11184), .ZN(n1298) );
  INVX0 U11239 ( .INP(n11185), .ZN(n1297) );
  INVX0 U11240 ( .INP(n11186), .ZN(n1296) );
  INVX0 U11241 ( .INP(n11187), .ZN(n1295) );
  INVX0 U11242 ( .INP(n11188), .ZN(n1294) );
  INVX0 U11243 ( .INP(n11189), .ZN(n1293) );
  INVX0 U11244 ( .INP(n11190), .ZN(n1292) );
  INVX0 U11245 ( .INP(n11191), .ZN(n1291) );
  INVX0 U11246 ( .INP(n11192), .ZN(n1290) );
  INVX0 U11247 ( .INP(n11193), .ZN(n129) );
  NOR2X0 U11248 ( .IN1(n11194), .IN2(n11195), .QN(n11193) );
  NAND2X0 U11249 ( .IN1(n11196), .IN2(n11197), .QN(n11195) );
  INVX0 U11250 ( .INP(n11198), .ZN(n11197) );
  NOR2X0 U11251 ( .IN1(n11199), .IN2(n9927), .QN(n11198) );
  NAND2X0 U11252 ( .IN1(n2152), .IN2(CRC_OUT_9_2), .QN(n11196) );
  NAND2X0 U11253 ( .IN1(n11200), .IN2(n11201), .QN(n11194) );
  INVX0 U11254 ( .INP(n11202), .ZN(n11201) );
  NOR2X0 U11255 ( .IN1(n9925), .IN2(n11203), .QN(n11202) );
  NAND2X0 U11256 ( .IN1(WX540), .IN2(n2339), .QN(n11200) );
  INVX0 U11257 ( .INP(n11204), .ZN(n126) );
  NOR2X0 U11258 ( .IN1(n11205), .IN2(n11206), .QN(n11204) );
  NAND2X0 U11259 ( .IN1(n11207), .IN2(n11208), .QN(n11206) );
  NAND2X0 U11260 ( .IN1(n9950), .IN2(n11209), .QN(n11208) );
  NAND2X0 U11261 ( .IN1(n2152), .IN2(CRC_OUT_9_3), .QN(n11207) );
  NAND2X0 U11262 ( .IN1(n11210), .IN2(n11211), .QN(n11205) );
  INVX0 U11263 ( .INP(n11212), .ZN(n11211) );
  NOR2X0 U11264 ( .IN1(n9925), .IN2(n11213), .QN(n11212) );
  NAND2X0 U11265 ( .IN1(WX538), .IN2(n2339), .QN(n11210) );
  INVX0 U11266 ( .INP(n11214), .ZN(n123) );
  NOR2X0 U11267 ( .IN1(n11215), .IN2(n11216), .QN(n11214) );
  NAND2X0 U11268 ( .IN1(n11217), .IN2(n11218), .QN(n11216) );
  NAND2X0 U11269 ( .IN1(n9950), .IN2(n11219), .QN(n11218) );
  NAND2X0 U11270 ( .IN1(n2152), .IN2(CRC_OUT_9_4), .QN(n11217) );
  NAND2X0 U11271 ( .IN1(n11220), .IN2(n11221), .QN(n11215) );
  NAND2X0 U11272 ( .IN1(n11222), .IN2(n2153), .QN(n11221) );
  NAND2X0 U11273 ( .IN1(WX536), .IN2(n2339), .QN(n11220) );
  INVX0 U11274 ( .INP(n11223), .ZN(n120) );
  NOR2X0 U11275 ( .IN1(n11224), .IN2(n11225), .QN(n11223) );
  NAND2X0 U11276 ( .IN1(n11226), .IN2(n11227), .QN(n11225) );
  NAND2X0 U11277 ( .IN1(n9950), .IN2(n11228), .QN(n11227) );
  NAND2X0 U11278 ( .IN1(n2152), .IN2(CRC_OUT_9_5), .QN(n11226) );
  NAND2X0 U11279 ( .IN1(n11229), .IN2(n11230), .QN(n11224) );
  INVX0 U11280 ( .INP(n11231), .ZN(n11230) );
  NOR2X0 U11281 ( .IN1(n9925), .IN2(n11232), .QN(n11231) );
  NAND2X0 U11282 ( .IN1(WX534), .IN2(n2339), .QN(n11229) );
  INVX0 U11283 ( .INP(n11233), .ZN(n117) );
  NOR2X0 U11284 ( .IN1(n11234), .IN2(n11235), .QN(n11233) );
  NAND2X0 U11285 ( .IN1(n11236), .IN2(n11237), .QN(n11235) );
  INVX0 U11286 ( .INP(n11238), .ZN(n11237) );
  NOR2X0 U11287 ( .IN1(n11239), .IN2(n9927), .QN(n11238) );
  NAND2X0 U11288 ( .IN1(n2152), .IN2(CRC_OUT_9_6), .QN(n11236) );
  NAND2X0 U11289 ( .IN1(n11240), .IN2(n11241), .QN(n11234) );
  INVX0 U11290 ( .INP(n11242), .ZN(n11241) );
  NOR2X0 U11291 ( .IN1(n9925), .IN2(n11243), .QN(n11242) );
  NAND2X0 U11292 ( .IN1(WX532), .IN2(n2339), .QN(n11240) );
  INVX0 U11293 ( .INP(n11244), .ZN(n114) );
  NOR2X0 U11294 ( .IN1(n11245), .IN2(n11246), .QN(n11244) );
  NAND2X0 U11295 ( .IN1(n11247), .IN2(n11248), .QN(n11246) );
  NAND2X0 U11296 ( .IN1(n9951), .IN2(n11249), .QN(n11248) );
  NAND2X0 U11297 ( .IN1(n2152), .IN2(CRC_OUT_9_7), .QN(n11247) );
  NAND2X0 U11298 ( .IN1(n11250), .IN2(n11251), .QN(n11245) );
  INVX0 U11299 ( .INP(n11252), .ZN(n11251) );
  NOR2X0 U11300 ( .IN1(n9925), .IN2(n11253), .QN(n11252) );
  NAND2X0 U11301 ( .IN1(WX530), .IN2(n2339), .QN(n11250) );
  INVX0 U11302 ( .INP(n11254), .ZN(n111) );
  NOR2X0 U11303 ( .IN1(n11255), .IN2(n11256), .QN(n11254) );
  NAND2X0 U11304 ( .IN1(n11257), .IN2(n11258), .QN(n11256) );
  NAND2X0 U11305 ( .IN1(n9950), .IN2(n11259), .QN(n11258) );
  NAND2X0 U11306 ( .IN1(n2152), .IN2(CRC_OUT_9_8), .QN(n11257) );
  NAND2X0 U11307 ( .IN1(n11260), .IN2(n11261), .QN(n11255) );
  INVX0 U11308 ( .INP(n11262), .ZN(n11261) );
  NOR2X0 U11309 ( .IN1(n9924), .IN2(n11263), .QN(n11262) );
  NAND2X0 U11310 ( .IN1(WX528), .IN2(n2339), .QN(n11260) );
  INVX0 U11311 ( .INP(n11264), .ZN(n108) );
  NOR2X0 U11312 ( .IN1(n11265), .IN2(n11266), .QN(n11264) );
  NAND2X0 U11313 ( .IN1(n11267), .IN2(n11268), .QN(n11266) );
  NAND2X0 U11314 ( .IN1(n9951), .IN2(n11269), .QN(n11268) );
  NAND2X0 U11315 ( .IN1(n2152), .IN2(CRC_OUT_9_9), .QN(n11267) );
  NAND2X0 U11316 ( .IN1(n11270), .IN2(n11271), .QN(n11265) );
  INVX0 U11317 ( .INP(n11272), .ZN(n11271) );
  NOR2X0 U11318 ( .IN1(n9924), .IN2(n11273), .QN(n11272) );
  NAND2X0 U11319 ( .IN1(WX526), .IN2(n2339), .QN(n11270) );
  INVX0 U11320 ( .INP(n11274), .ZN(n1079) );
  INVX0 U11321 ( .INP(n11275), .ZN(n1078) );
  INVX0 U11322 ( .INP(n11276), .ZN(n1077) );
  INVX0 U11323 ( .INP(n11277), .ZN(n1076) );
  INVX0 U11324 ( .INP(n11278), .ZN(n1075) );
  INVX0 U11325 ( .INP(n11279), .ZN(n1074) );
  INVX0 U11326 ( .INP(n11280), .ZN(n1073) );
  INVX0 U11327 ( .INP(n11281), .ZN(n1072) );
  INVX0 U11328 ( .INP(n11282), .ZN(n1071) );
  INVX0 U11329 ( .INP(n11283), .ZN(n1070) );
  INVX0 U11330 ( .INP(n11284), .ZN(n1069) );
  INVX0 U11331 ( .INP(n11285), .ZN(n1068) );
  INVX0 U11332 ( .INP(n11286), .ZN(n1067) );
  INVX0 U11333 ( .INP(n11287), .ZN(n1066) );
  INVX0 U11334 ( .INP(n11288), .ZN(n1065) );
  INVX0 U11335 ( .INP(n11289), .ZN(n1064) );
  INVX0 U11336 ( .INP(n11290), .ZN(n1063) );
  INVX0 U11337 ( .INP(n11291), .ZN(n1062) );
  INVX0 U11338 ( .INP(n11292), .ZN(n1061) );
  INVX0 U11339 ( .INP(n11293), .ZN(n1060) );
  INVX0 U11340 ( .INP(n11294), .ZN(n1059) );
  INVX0 U11341 ( .INP(n11295), .ZN(n1058) );
  INVX0 U11342 ( .INP(n11296), .ZN(n1057) );
  INVX0 U11343 ( .INP(n11297), .ZN(n1056) );
  INVX0 U11344 ( .INP(n11298), .ZN(n1055) );
  INVX0 U11345 ( .INP(n11299), .ZN(n1054) );
  INVX0 U11346 ( .INP(n11300), .ZN(n1053) );
  INVX0 U11347 ( .INP(n11301), .ZN(n1052) );
  INVX0 U11348 ( .INP(n11302), .ZN(n1051) );
  INVX0 U11349 ( .INP(n11303), .ZN(n1050) );
  INVX0 U11350 ( .INP(n11304), .ZN(n1049) );
  INVX0 U11351 ( .INP(n11305), .ZN(n104) );
  NOR2X0 U11352 ( .IN1(n11306), .IN2(n11307), .QN(n11305) );
  NAND2X0 U11353 ( .IN1(n11308), .IN2(n11309), .QN(n11307) );
  INVX0 U11354 ( .INP(n11310), .ZN(n11309) );
  NOR2X0 U11355 ( .IN1(n11311), .IN2(n9927), .QN(n11310) );
  NAND2X0 U11356 ( .IN1(n2152), .IN2(CRC_OUT_9_10), .QN(n11308) );
  NAND2X0 U11357 ( .IN1(n11312), .IN2(n11313), .QN(n11306) );
  NAND2X0 U11358 ( .IN1(n11314), .IN2(n2153), .QN(n11313) );
  NAND2X0 U11359 ( .IN1(WX524), .IN2(n2339), .QN(n11312) );
  INVX0 U11360 ( .INP(n11315), .ZN(n101) );
  NOR2X0 U11361 ( .IN1(n11316), .IN2(n11317), .QN(n11315) );
  NAND2X0 U11362 ( .IN1(n11318), .IN2(n11319), .QN(n11317) );
  NAND2X0 U11363 ( .IN1(n9951), .IN2(n11320), .QN(n11319) );
  NAND2X0 U11364 ( .IN1(n2152), .IN2(CRC_OUT_9_11), .QN(n11318) );
  NAND2X0 U11365 ( .IN1(n11321), .IN2(n11322), .QN(n11316) );
  INVX0 U11366 ( .INP(n11323), .ZN(n11322) );
  NOR2X0 U11367 ( .IN1(n9924), .IN2(n11324), .QN(n11323) );
  NAND2X0 U11368 ( .IN1(WX522), .IN2(n2339), .QN(n11321) );
  NOR2X0 U11369 ( .IN1(n10321), .IN2(WX485), .QN(n1) );
  NOR2X0 U11370 ( .IN1(n18457), .IN2(n10234), .QN(WX9789) );
  NOR2X0 U11371 ( .IN1(n18456), .IN2(n10234), .QN(WX9787) );
  NOR2X0 U11372 ( .IN1(n18455), .IN2(n10234), .QN(WX9785) );
  NOR2X0 U11373 ( .IN1(n18454), .IN2(n10234), .QN(WX9783) );
  NOR2X0 U11374 ( .IN1(n10321), .IN2(n9840), .QN(WX9781) );
  NOR2X0 U11375 ( .IN1(n18453), .IN2(n10234), .QN(WX9779) );
  NOR2X0 U11376 ( .IN1(n18452), .IN2(n10234), .QN(WX9777) );
  NOR2X0 U11377 ( .IN1(n18451), .IN2(n10234), .QN(WX9775) );
  NOR2X0 U11378 ( .IN1(n18450), .IN2(n10234), .QN(WX9773) );
  NOR2X0 U11379 ( .IN1(n18449), .IN2(n10234), .QN(WX9771) );
  NOR2X0 U11380 ( .IN1(n18448), .IN2(n10235), .QN(WX9769) );
  NOR2X0 U11381 ( .IN1(n18447), .IN2(n10235), .QN(WX9767) );
  NOR2X0 U11382 ( .IN1(n18446), .IN2(n10235), .QN(WX9765) );
  NOR2X0 U11383 ( .IN1(n18445), .IN2(n10235), .QN(WX9763) );
  NOR2X0 U11384 ( .IN1(n18444), .IN2(n10235), .QN(WX9761) );
  NOR2X0 U11385 ( .IN1(n18443), .IN2(n10235), .QN(WX9759) );
  NAND2X0 U11386 ( .IN1(n11325), .IN2(n11326), .QN(WX9757) );
  NOR2X0 U11387 ( .IN1(n11327), .IN2(n11328), .QN(n11326) );
  NOR2X0 U11388 ( .IN1(n11329), .IN2(n9935), .QN(n11328) );
  NOR2X0 U11389 ( .IN1(n10809), .IN2(n9907), .QN(n11327) );
  NOR2X0 U11390 ( .IN1(n11330), .IN2(n11331), .QN(n10809) );
  INVX0 U11391 ( .INP(n11332), .ZN(n11331) );
  NAND2X0 U11392 ( .IN1(n11333), .IN2(n11334), .QN(n11332) );
  NOR2X0 U11393 ( .IN1(n11334), .IN2(n11333), .QN(n11330) );
  INVX0 U11394 ( .INP(n11335), .ZN(n11333) );
  NOR2X0 U11395 ( .IN1(n11336), .IN2(n11337), .QN(n11335) );
  NOR2X0 U11396 ( .IN1(WX11243), .IN2(n9246), .QN(n11337) );
  INVX0 U11397 ( .INP(n11338), .ZN(n11336) );
  NAND2X0 U11398 ( .IN1(n9246), .IN2(WX11243), .QN(n11338) );
  NOR2X0 U11399 ( .IN1(n11339), .IN2(n11340), .QN(n11334) );
  INVX0 U11400 ( .INP(n11341), .ZN(n11340) );
  NAND2X0 U11401 ( .IN1(n9245), .IN2(WX11115), .QN(n11341) );
  NOR2X0 U11402 ( .IN1(WX11115), .IN2(n9245), .QN(n11339) );
  NOR2X0 U11403 ( .IN1(n11342), .IN2(n11343), .QN(n11325) );
  NOR2X0 U11404 ( .IN1(DFF_1504_n1), .IN2(n9964), .QN(n11343) );
  NOR2X0 U11405 ( .IN1(n11345), .IN2(n11081), .QN(n11342) );
  NAND2X0 U11406 ( .IN1(n10197), .IN2(n8321), .QN(n11081) );
  NAND2X0 U11407 ( .IN1(n11346), .IN2(n11347), .QN(WX9755) );
  NOR2X0 U11408 ( .IN1(n11348), .IN2(n11349), .QN(n11347) );
  NOR2X0 U11409 ( .IN1(n9944), .IN2(n11350), .QN(n11349) );
  NOR2X0 U11410 ( .IN1(n10818), .IN2(n9907), .QN(n11348) );
  NOR2X0 U11411 ( .IN1(n11351), .IN2(n11352), .QN(n10818) );
  INVX0 U11412 ( .INP(n11353), .ZN(n11352) );
  NAND2X0 U11413 ( .IN1(n11354), .IN2(n11355), .QN(n11353) );
  NOR2X0 U11414 ( .IN1(n11355), .IN2(n11354), .QN(n11351) );
  INVX0 U11415 ( .INP(n11356), .ZN(n11354) );
  NOR2X0 U11416 ( .IN1(n11357), .IN2(n11358), .QN(n11356) );
  NOR2X0 U11417 ( .IN1(WX11241), .IN2(n9248), .QN(n11358) );
  INVX0 U11418 ( .INP(n11359), .ZN(n11357) );
  NAND2X0 U11419 ( .IN1(n9248), .IN2(WX11241), .QN(n11359) );
  NOR2X0 U11420 ( .IN1(n11360), .IN2(n11361), .QN(n11355) );
  INVX0 U11421 ( .INP(n11362), .ZN(n11361) );
  NAND2X0 U11422 ( .IN1(n9247), .IN2(WX11113), .QN(n11362) );
  NOR2X0 U11423 ( .IN1(WX11113), .IN2(n9247), .QN(n11360) );
  NOR2X0 U11424 ( .IN1(n11363), .IN2(n11364), .QN(n11346) );
  NOR2X0 U11425 ( .IN1(DFF_1505_n1), .IN2(n9966), .QN(n11364) );
  NOR2X0 U11426 ( .IN1(n9998), .IN2(n11082), .QN(n11363) );
  NAND2X0 U11427 ( .IN1(n10197), .IN2(n8322), .QN(n11082) );
  NAND2X0 U11428 ( .IN1(n11365), .IN2(n11366), .QN(WX9753) );
  NOR2X0 U11429 ( .IN1(n11367), .IN2(n11368), .QN(n11366) );
  NOR2X0 U11430 ( .IN1(n11369), .IN2(n9927), .QN(n11368) );
  INVX0 U11431 ( .INP(n11370), .ZN(n11367) );
  NAND2X0 U11432 ( .IN1(n2153), .IN2(n10826), .QN(n11370) );
  NOR2X0 U11433 ( .IN1(n11371), .IN2(n11372), .QN(n10826) );
  INVX0 U11434 ( .INP(n11373), .ZN(n11372) );
  NAND2X0 U11435 ( .IN1(n11374), .IN2(n11375), .QN(n11373) );
  NOR2X0 U11436 ( .IN1(n11375), .IN2(n11374), .QN(n11371) );
  INVX0 U11437 ( .INP(n11376), .ZN(n11374) );
  NOR2X0 U11438 ( .IN1(n11377), .IN2(n11378), .QN(n11376) );
  NOR2X0 U11439 ( .IN1(n9847), .IN2(n9250), .QN(n11378) );
  INVX0 U11440 ( .INP(n11379), .ZN(n11377) );
  NAND2X0 U11441 ( .IN1(n9250), .IN2(n9847), .QN(n11379) );
  NOR2X0 U11442 ( .IN1(n11380), .IN2(n11381), .QN(n11375) );
  INVX0 U11443 ( .INP(n11382), .ZN(n11381) );
  NAND2X0 U11444 ( .IN1(n9249), .IN2(WX11111), .QN(n11382) );
  NOR2X0 U11445 ( .IN1(WX11111), .IN2(n9249), .QN(n11380) );
  NOR2X0 U11446 ( .IN1(n11383), .IN2(n11384), .QN(n11365) );
  NOR2X0 U11447 ( .IN1(n9976), .IN2(n9864), .QN(n11384) );
  NOR2X0 U11448 ( .IN1(n9998), .IN2(n11083), .QN(n11383) );
  NAND2X0 U11449 ( .IN1(n10197), .IN2(n8323), .QN(n11083) );
  NAND2X0 U11450 ( .IN1(n11385), .IN2(n11386), .QN(WX9751) );
  NOR2X0 U11451 ( .IN1(n11387), .IN2(n11388), .QN(n11386) );
  NOR2X0 U11452 ( .IN1(n9943), .IN2(n11389), .QN(n11388) );
  NOR2X0 U11453 ( .IN1(n10835), .IN2(n9907), .QN(n11387) );
  NOR2X0 U11454 ( .IN1(n11390), .IN2(n11391), .QN(n10835) );
  INVX0 U11455 ( .INP(n11392), .ZN(n11391) );
  NAND2X0 U11456 ( .IN1(n11393), .IN2(n11394), .QN(n11392) );
  NOR2X0 U11457 ( .IN1(n11394), .IN2(n11393), .QN(n11390) );
  INVX0 U11458 ( .INP(n11395), .ZN(n11393) );
  NOR2X0 U11459 ( .IN1(n11396), .IN2(n11397), .QN(n11395) );
  NOR2X0 U11460 ( .IN1(WX11237), .IN2(n9252), .QN(n11397) );
  INVX0 U11461 ( .INP(n11398), .ZN(n11396) );
  NAND2X0 U11462 ( .IN1(n9252), .IN2(WX11237), .QN(n11398) );
  NOR2X0 U11463 ( .IN1(n11399), .IN2(n11400), .QN(n11394) );
  INVX0 U11464 ( .INP(n11401), .ZN(n11400) );
  NAND2X0 U11465 ( .IN1(n9251), .IN2(WX11109), .QN(n11401) );
  NOR2X0 U11466 ( .IN1(WX11109), .IN2(n9251), .QN(n11399) );
  NOR2X0 U11467 ( .IN1(n11402), .IN2(n11403), .QN(n11385) );
  NOR2X0 U11468 ( .IN1(DFF_1507_n1), .IN2(n9966), .QN(n11403) );
  NOR2X0 U11469 ( .IN1(n9998), .IN2(n11084), .QN(n11402) );
  NAND2X0 U11470 ( .IN1(n10197), .IN2(n8324), .QN(n11084) );
  NAND2X0 U11471 ( .IN1(n11404), .IN2(n11405), .QN(WX9749) );
  NOR2X0 U11472 ( .IN1(n11406), .IN2(n11407), .QN(n11405) );
  NOR2X0 U11473 ( .IN1(n11408), .IN2(n9927), .QN(n11407) );
  INVX0 U11474 ( .INP(n11409), .ZN(n11406) );
  NAND2X0 U11475 ( .IN1(n2153), .IN2(n10843), .QN(n11409) );
  NOR2X0 U11476 ( .IN1(n11410), .IN2(n11411), .QN(n10843) );
  INVX0 U11477 ( .INP(n11412), .ZN(n11411) );
  NAND2X0 U11478 ( .IN1(n11413), .IN2(n11414), .QN(n11412) );
  NOR2X0 U11479 ( .IN1(n11414), .IN2(n11413), .QN(n11410) );
  INVX0 U11480 ( .INP(n11415), .ZN(n11413) );
  NOR2X0 U11481 ( .IN1(n11416), .IN2(n11417), .QN(n11415) );
  INVX0 U11482 ( .INP(n11418), .ZN(n11417) );
  NAND2X0 U11483 ( .IN1(test_so96), .IN2(WX11235), .QN(n11418) );
  NOR2X0 U11484 ( .IN1(WX11235), .IN2(test_so96), .QN(n11416) );
  NOR2X0 U11485 ( .IN1(n11419), .IN2(n11420), .QN(n11414) );
  INVX0 U11486 ( .INP(n11421), .ZN(n11420) );
  NAND2X0 U11487 ( .IN1(n9253), .IN2(WX11107), .QN(n11421) );
  NOR2X0 U11488 ( .IN1(WX11107), .IN2(n9253), .QN(n11419) );
  NOR2X0 U11489 ( .IN1(n11422), .IN2(n11423), .QN(n11404) );
  NOR2X0 U11490 ( .IN1(DFF_1508_n1), .IN2(n9966), .QN(n11423) );
  NOR2X0 U11491 ( .IN1(n9998), .IN2(n11085), .QN(n11422) );
  NAND2X0 U11492 ( .IN1(n10197), .IN2(n8325), .QN(n11085) );
  NAND2X0 U11493 ( .IN1(n11424), .IN2(n11425), .QN(WX9747) );
  NOR2X0 U11494 ( .IN1(n11426), .IN2(n11427), .QN(n11425) );
  NOR2X0 U11495 ( .IN1(n11428), .IN2(n9927), .QN(n11427) );
  NOR2X0 U11496 ( .IN1(n10852), .IN2(n9907), .QN(n11426) );
  NOR2X0 U11497 ( .IN1(n11429), .IN2(n11430), .QN(n10852) );
  INVX0 U11498 ( .INP(n11431), .ZN(n11430) );
  NAND2X0 U11499 ( .IN1(n11432), .IN2(n11433), .QN(n11431) );
  NOR2X0 U11500 ( .IN1(n11433), .IN2(n11432), .QN(n11429) );
  INVX0 U11501 ( .INP(n11434), .ZN(n11432) );
  NOR2X0 U11502 ( .IN1(n11435), .IN2(n11436), .QN(n11434) );
  NOR2X0 U11503 ( .IN1(WX11233), .IN2(n9255), .QN(n11436) );
  INVX0 U11504 ( .INP(n11437), .ZN(n11435) );
  NAND2X0 U11505 ( .IN1(n9255), .IN2(WX11233), .QN(n11437) );
  NOR2X0 U11506 ( .IN1(n11438), .IN2(n11439), .QN(n11433) );
  INVX0 U11507 ( .INP(n11440), .ZN(n11439) );
  NAND2X0 U11508 ( .IN1(n9254), .IN2(WX11105), .QN(n11440) );
  NOR2X0 U11509 ( .IN1(WX11105), .IN2(n9254), .QN(n11438) );
  NOR2X0 U11510 ( .IN1(n11441), .IN2(n11442), .QN(n11424) );
  NOR2X0 U11511 ( .IN1(DFF_1509_n1), .IN2(n9966), .QN(n11442) );
  NOR2X0 U11512 ( .IN1(n9998), .IN2(n11086), .QN(n11441) );
  NAND2X0 U11513 ( .IN1(test_so79), .IN2(n10215), .QN(n11086) );
  NAND2X0 U11514 ( .IN1(n11443), .IN2(n11444), .QN(WX9745) );
  NOR2X0 U11515 ( .IN1(n11445), .IN2(n11446), .QN(n11444) );
  NOR2X0 U11516 ( .IN1(n11447), .IN2(n9927), .QN(n11446) );
  INVX0 U11517 ( .INP(n11448), .ZN(n11445) );
  NAND2X0 U11518 ( .IN1(n2153), .IN2(n10860), .QN(n11448) );
  NOR2X0 U11519 ( .IN1(n11449), .IN2(n11450), .QN(n10860) );
  INVX0 U11520 ( .INP(n11451), .ZN(n11450) );
  NAND2X0 U11521 ( .IN1(n11452), .IN2(n11453), .QN(n11451) );
  NOR2X0 U11522 ( .IN1(n11453), .IN2(n11452), .QN(n11449) );
  INVX0 U11523 ( .INP(n11454), .ZN(n11452) );
  NOR2X0 U11524 ( .IN1(n11455), .IN2(n11456), .QN(n11454) );
  INVX0 U11525 ( .INP(n11457), .ZN(n11456) );
  NAND2X0 U11526 ( .IN1(test_so94), .IN2(WX11231), .QN(n11457) );
  NOR2X0 U11527 ( .IN1(WX11231), .IN2(test_so94), .QN(n11455) );
  NOR2X0 U11528 ( .IN1(n11458), .IN2(n11459), .QN(n11453) );
  INVX0 U11529 ( .INP(n11460), .ZN(n11459) );
  NAND2X0 U11530 ( .IN1(n9257), .IN2(WX11039), .QN(n11460) );
  NOR2X0 U11531 ( .IN1(WX11039), .IN2(n9257), .QN(n11458) );
  NOR2X0 U11532 ( .IN1(n11461), .IN2(n11462), .QN(n11443) );
  NOR2X0 U11533 ( .IN1(DFF_1510_n1), .IN2(n9966), .QN(n11462) );
  NOR2X0 U11534 ( .IN1(n9998), .IN2(n11087), .QN(n11461) );
  NAND2X0 U11535 ( .IN1(n10196), .IN2(n8328), .QN(n11087) );
  NAND2X0 U11536 ( .IN1(n11463), .IN2(n11464), .QN(WX9743) );
  NOR2X0 U11537 ( .IN1(n11465), .IN2(n11466), .QN(n11464) );
  NOR2X0 U11538 ( .IN1(n11467), .IN2(n9928), .QN(n11466) );
  NOR2X0 U11539 ( .IN1(n10869), .IN2(n9907), .QN(n11465) );
  NOR2X0 U11540 ( .IN1(n11468), .IN2(n11469), .QN(n10869) );
  INVX0 U11541 ( .INP(n11470), .ZN(n11469) );
  NAND2X0 U11542 ( .IN1(n11471), .IN2(n11472), .QN(n11470) );
  NOR2X0 U11543 ( .IN1(n11472), .IN2(n11471), .QN(n11468) );
  INVX0 U11544 ( .INP(n11473), .ZN(n11471) );
  NOR2X0 U11545 ( .IN1(n11474), .IN2(n11475), .QN(n11473) );
  NOR2X0 U11546 ( .IN1(WX11229), .IN2(n9259), .QN(n11475) );
  INVX0 U11547 ( .INP(n11476), .ZN(n11474) );
  NAND2X0 U11548 ( .IN1(n9259), .IN2(WX11229), .QN(n11476) );
  NOR2X0 U11549 ( .IN1(n11477), .IN2(n11478), .QN(n11472) );
  INVX0 U11550 ( .INP(n11479), .ZN(n11478) );
  NAND2X0 U11551 ( .IN1(n9258), .IN2(WX11101), .QN(n11479) );
  NOR2X0 U11552 ( .IN1(WX11101), .IN2(n9258), .QN(n11477) );
  NOR2X0 U11553 ( .IN1(n11480), .IN2(n11481), .QN(n11463) );
  NOR2X0 U11554 ( .IN1(DFF_1511_n1), .IN2(n9966), .QN(n11481) );
  NOR2X0 U11555 ( .IN1(n9998), .IN2(n11088), .QN(n11480) );
  NAND2X0 U11556 ( .IN1(n10196), .IN2(n8329), .QN(n11088) );
  NAND2X0 U11557 ( .IN1(n11482), .IN2(n11483), .QN(WX9741) );
  NOR2X0 U11558 ( .IN1(n11484), .IN2(n11485), .QN(n11483) );
  NOR2X0 U11559 ( .IN1(n11486), .IN2(n9928), .QN(n11485) );
  INVX0 U11560 ( .INP(n11487), .ZN(n11484) );
  NAND2X0 U11561 ( .IN1(n2153), .IN2(n10877), .QN(n11487) );
  NOR2X0 U11562 ( .IN1(n11488), .IN2(n11489), .QN(n10877) );
  INVX0 U11563 ( .INP(n11490), .ZN(n11489) );
  NAND2X0 U11564 ( .IN1(n11491), .IN2(n11492), .QN(n11490) );
  NOR2X0 U11565 ( .IN1(n11492), .IN2(n11491), .QN(n11488) );
  INVX0 U11566 ( .INP(n11493), .ZN(n11491) );
  NOR2X0 U11567 ( .IN1(n11494), .IN2(n11495), .QN(n11493) );
  INVX0 U11568 ( .INP(n11496), .ZN(n11495) );
  NAND2X0 U11569 ( .IN1(test_so92), .IN2(WX11227), .QN(n11496) );
  NOR2X0 U11570 ( .IN1(WX11227), .IN2(test_so92), .QN(n11494) );
  NOR2X0 U11571 ( .IN1(n11497), .IN2(n11498), .QN(n11492) );
  INVX0 U11572 ( .INP(n11499), .ZN(n11498) );
  NAND2X0 U11573 ( .IN1(n9260), .IN2(WX11099), .QN(n11499) );
  NOR2X0 U11574 ( .IN1(WX11099), .IN2(n9260), .QN(n11497) );
  NOR2X0 U11575 ( .IN1(n11500), .IN2(n11501), .QN(n11482) );
  NOR2X0 U11576 ( .IN1(DFF_1512_n1), .IN2(n9966), .QN(n11501) );
  NOR2X0 U11577 ( .IN1(n9998), .IN2(n11089), .QN(n11500) );
  NAND2X0 U11578 ( .IN1(n10196), .IN2(n8330), .QN(n11089) );
  NAND2X0 U11579 ( .IN1(n11502), .IN2(n11503), .QN(WX9739) );
  NOR2X0 U11580 ( .IN1(n11504), .IN2(n11505), .QN(n11503) );
  NOR2X0 U11581 ( .IN1(n11506), .IN2(n9928), .QN(n11505) );
  NOR2X0 U11582 ( .IN1(n10886), .IN2(n9907), .QN(n11504) );
  NOR2X0 U11583 ( .IN1(n11507), .IN2(n11508), .QN(n10886) );
  INVX0 U11584 ( .INP(n11509), .ZN(n11508) );
  NAND2X0 U11585 ( .IN1(n11510), .IN2(n11511), .QN(n11509) );
  NOR2X0 U11586 ( .IN1(n11511), .IN2(n11510), .QN(n11507) );
  INVX0 U11587 ( .INP(n11512), .ZN(n11510) );
  NOR2X0 U11588 ( .IN1(n11513), .IN2(n11514), .QN(n11512) );
  NOR2X0 U11589 ( .IN1(WX11225), .IN2(n9262), .QN(n11514) );
  INVX0 U11590 ( .INP(n11515), .ZN(n11513) );
  NAND2X0 U11591 ( .IN1(n9262), .IN2(WX11225), .QN(n11515) );
  NOR2X0 U11592 ( .IN1(n11516), .IN2(n11517), .QN(n11511) );
  INVX0 U11593 ( .INP(n11518), .ZN(n11517) );
  NAND2X0 U11594 ( .IN1(n9261), .IN2(WX11097), .QN(n11518) );
  NOR2X0 U11595 ( .IN1(WX11097), .IN2(n9261), .QN(n11516) );
  NOR2X0 U11596 ( .IN1(n11519), .IN2(n11520), .QN(n11502) );
  NOR2X0 U11597 ( .IN1(DFF_1513_n1), .IN2(n9966), .QN(n11520) );
  NOR2X0 U11598 ( .IN1(n9998), .IN2(n11090), .QN(n11519) );
  NAND2X0 U11599 ( .IN1(n10196), .IN2(n8331), .QN(n11090) );
  NAND2X0 U11600 ( .IN1(n11521), .IN2(n11522), .QN(WX9737) );
  NOR2X0 U11601 ( .IN1(n11523), .IN2(n11524), .QN(n11522) );
  NOR2X0 U11602 ( .IN1(n11525), .IN2(n9928), .QN(n11524) );
  NOR2X0 U11603 ( .IN1(n10895), .IN2(n9907), .QN(n11523) );
  NOR2X0 U11604 ( .IN1(n11526), .IN2(n11527), .QN(n10895) );
  INVX0 U11605 ( .INP(n11528), .ZN(n11527) );
  NAND2X0 U11606 ( .IN1(n11529), .IN2(n11530), .QN(n11528) );
  NOR2X0 U11607 ( .IN1(n11530), .IN2(n11529), .QN(n11526) );
  INVX0 U11608 ( .INP(n11531), .ZN(n11529) );
  NOR2X0 U11609 ( .IN1(n11532), .IN2(n11533), .QN(n11531) );
  NOR2X0 U11610 ( .IN1(WX11223), .IN2(n9264), .QN(n11533) );
  INVX0 U11611 ( .INP(n11534), .ZN(n11532) );
  NAND2X0 U11612 ( .IN1(n9264), .IN2(WX11223), .QN(n11534) );
  NOR2X0 U11613 ( .IN1(n11535), .IN2(n11536), .QN(n11530) );
  INVX0 U11614 ( .INP(n11537), .ZN(n11536) );
  NAND2X0 U11615 ( .IN1(n9263), .IN2(WX11095), .QN(n11537) );
  NOR2X0 U11616 ( .IN1(WX11095), .IN2(n9263), .QN(n11535) );
  NOR2X0 U11617 ( .IN1(n11538), .IN2(n11539), .QN(n11521) );
  NOR2X0 U11618 ( .IN1(DFF_1514_n1), .IN2(n9966), .QN(n11539) );
  NOR2X0 U11619 ( .IN1(n9998), .IN2(n11091), .QN(n11538) );
  NAND2X0 U11620 ( .IN1(n10196), .IN2(n8332), .QN(n11091) );
  NAND2X0 U11621 ( .IN1(n11540), .IN2(n11541), .QN(WX9735) );
  NOR2X0 U11622 ( .IN1(n11542), .IN2(n11543), .QN(n11541) );
  NOR2X0 U11623 ( .IN1(n11544), .IN2(n9928), .QN(n11543) );
  NOR2X0 U11624 ( .IN1(n10904), .IN2(n9907), .QN(n11542) );
  NOR2X0 U11625 ( .IN1(n11545), .IN2(n11546), .QN(n10904) );
  INVX0 U11626 ( .INP(n11547), .ZN(n11546) );
  NAND2X0 U11627 ( .IN1(n11548), .IN2(n11549), .QN(n11547) );
  NOR2X0 U11628 ( .IN1(n11549), .IN2(n11548), .QN(n11545) );
  INVX0 U11629 ( .INP(n11550), .ZN(n11548) );
  NOR2X0 U11630 ( .IN1(n11551), .IN2(n11552), .QN(n11550) );
  NOR2X0 U11631 ( .IN1(WX11221), .IN2(n9266), .QN(n11552) );
  INVX0 U11632 ( .INP(n11553), .ZN(n11551) );
  NAND2X0 U11633 ( .IN1(n9266), .IN2(WX11221), .QN(n11553) );
  NOR2X0 U11634 ( .IN1(n11554), .IN2(n11555), .QN(n11549) );
  INVX0 U11635 ( .INP(n11556), .ZN(n11555) );
  NAND2X0 U11636 ( .IN1(n9265), .IN2(WX11093), .QN(n11556) );
  NOR2X0 U11637 ( .IN1(WX11093), .IN2(n9265), .QN(n11554) );
  NOR2X0 U11638 ( .IN1(n11557), .IN2(n11558), .QN(n11540) );
  NOR2X0 U11639 ( .IN1(DFF_1515_n1), .IN2(n9966), .QN(n11558) );
  NOR2X0 U11640 ( .IN1(n9998), .IN2(n11092), .QN(n11557) );
  NAND2X0 U11641 ( .IN1(n10196), .IN2(n8333), .QN(n11092) );
  NAND2X0 U11642 ( .IN1(n11559), .IN2(n11560), .QN(WX9733) );
  NOR2X0 U11643 ( .IN1(n11561), .IN2(n11562), .QN(n11560) );
  NOR2X0 U11644 ( .IN1(n11563), .IN2(n9928), .QN(n11562) );
  NOR2X0 U11645 ( .IN1(n10913), .IN2(n9907), .QN(n11561) );
  NOR2X0 U11646 ( .IN1(n11564), .IN2(n11565), .QN(n10913) );
  INVX0 U11647 ( .INP(n11566), .ZN(n11565) );
  NAND2X0 U11648 ( .IN1(n11567), .IN2(n11568), .QN(n11566) );
  NOR2X0 U11649 ( .IN1(n11568), .IN2(n11567), .QN(n11564) );
  INVX0 U11650 ( .INP(n11569), .ZN(n11567) );
  NOR2X0 U11651 ( .IN1(n11570), .IN2(n11571), .QN(n11569) );
  NOR2X0 U11652 ( .IN1(WX11219), .IN2(n9268), .QN(n11571) );
  INVX0 U11653 ( .INP(n11572), .ZN(n11570) );
  NAND2X0 U11654 ( .IN1(n9268), .IN2(WX11219), .QN(n11572) );
  NOR2X0 U11655 ( .IN1(n11573), .IN2(n11574), .QN(n11568) );
  INVX0 U11656 ( .INP(n11575), .ZN(n11574) );
  NAND2X0 U11657 ( .IN1(n9267), .IN2(WX11091), .QN(n11575) );
  NOR2X0 U11658 ( .IN1(WX11091), .IN2(n9267), .QN(n11573) );
  NOR2X0 U11659 ( .IN1(n11576), .IN2(n11577), .QN(n11559) );
  NOR2X0 U11660 ( .IN1(DFF_1516_n1), .IN2(n9966), .QN(n11577) );
  NOR2X0 U11661 ( .IN1(n9998), .IN2(n11093), .QN(n11576) );
  NAND2X0 U11662 ( .IN1(n10196), .IN2(n8334), .QN(n11093) );
  NAND2X0 U11663 ( .IN1(n11578), .IN2(n11579), .QN(WX9731) );
  NOR2X0 U11664 ( .IN1(n11580), .IN2(n11581), .QN(n11579) );
  NOR2X0 U11665 ( .IN1(n11582), .IN2(n9928), .QN(n11581) );
  NOR2X0 U11666 ( .IN1(n10922), .IN2(n9907), .QN(n11580) );
  NOR2X0 U11667 ( .IN1(n11583), .IN2(n11584), .QN(n10922) );
  INVX0 U11668 ( .INP(n11585), .ZN(n11584) );
  NAND2X0 U11669 ( .IN1(n11586), .IN2(n11587), .QN(n11585) );
  NOR2X0 U11670 ( .IN1(n11587), .IN2(n11586), .QN(n11583) );
  INVX0 U11671 ( .INP(n11588), .ZN(n11586) );
  NOR2X0 U11672 ( .IN1(n11589), .IN2(n11590), .QN(n11588) );
  NOR2X0 U11673 ( .IN1(WX11217), .IN2(n9270), .QN(n11590) );
  INVX0 U11674 ( .INP(n11591), .ZN(n11589) );
  NAND2X0 U11675 ( .IN1(n9270), .IN2(WX11217), .QN(n11591) );
  NOR2X0 U11676 ( .IN1(n11592), .IN2(n11593), .QN(n11587) );
  INVX0 U11677 ( .INP(n11594), .ZN(n11593) );
  NAND2X0 U11678 ( .IN1(n9269), .IN2(WX11089), .QN(n11594) );
  NOR2X0 U11679 ( .IN1(WX11089), .IN2(n9269), .QN(n11592) );
  NOR2X0 U11680 ( .IN1(n11595), .IN2(n11596), .QN(n11578) );
  NOR2X0 U11681 ( .IN1(DFF_1517_n1), .IN2(n9966), .QN(n11596) );
  NOR2X0 U11682 ( .IN1(n9997), .IN2(n11094), .QN(n11595) );
  NAND2X0 U11683 ( .IN1(n10196), .IN2(n8335), .QN(n11094) );
  NAND2X0 U11684 ( .IN1(n11597), .IN2(n11598), .QN(WX9729) );
  NOR2X0 U11685 ( .IN1(n11599), .IN2(n11600), .QN(n11598) );
  NOR2X0 U11686 ( .IN1(n9944), .IN2(n11601), .QN(n11600) );
  NOR2X0 U11687 ( .IN1(n10931), .IN2(n9907), .QN(n11599) );
  NOR2X0 U11688 ( .IN1(n11602), .IN2(n11603), .QN(n10931) );
  INVX0 U11689 ( .INP(n11604), .ZN(n11603) );
  NAND2X0 U11690 ( .IN1(n11605), .IN2(n11606), .QN(n11604) );
  NOR2X0 U11691 ( .IN1(n11606), .IN2(n11605), .QN(n11602) );
  INVX0 U11692 ( .INP(n11607), .ZN(n11605) );
  NOR2X0 U11693 ( .IN1(n11608), .IN2(n11609), .QN(n11607) );
  NOR2X0 U11694 ( .IN1(WX11215), .IN2(n9272), .QN(n11609) );
  INVX0 U11695 ( .INP(n11610), .ZN(n11608) );
  NAND2X0 U11696 ( .IN1(n9272), .IN2(WX11215), .QN(n11610) );
  NOR2X0 U11697 ( .IN1(n11611), .IN2(n11612), .QN(n11606) );
  INVX0 U11698 ( .INP(n11613), .ZN(n11612) );
  NAND2X0 U11699 ( .IN1(n9271), .IN2(WX11087), .QN(n11613) );
  NOR2X0 U11700 ( .IN1(WX11087), .IN2(n9271), .QN(n11611) );
  NOR2X0 U11701 ( .IN1(n11614), .IN2(n11615), .QN(n11597) );
  NOR2X0 U11702 ( .IN1(DFF_1518_n1), .IN2(n9965), .QN(n11615) );
  NOR2X0 U11703 ( .IN1(n9997), .IN2(n11095), .QN(n11614) );
  NAND2X0 U11704 ( .IN1(n10196), .IN2(n8336), .QN(n11095) );
  NAND2X0 U11705 ( .IN1(n11616), .IN2(n11617), .QN(WX9727) );
  NOR2X0 U11706 ( .IN1(n11618), .IN2(n11619), .QN(n11617) );
  NOR2X0 U11707 ( .IN1(n11620), .IN2(n9928), .QN(n11619) );
  NOR2X0 U11708 ( .IN1(n10940), .IN2(n9908), .QN(n11618) );
  NOR2X0 U11709 ( .IN1(n11621), .IN2(n11622), .QN(n10940) );
  INVX0 U11710 ( .INP(n11623), .ZN(n11622) );
  NAND2X0 U11711 ( .IN1(n11624), .IN2(n11625), .QN(n11623) );
  NOR2X0 U11712 ( .IN1(n11625), .IN2(n11624), .QN(n11621) );
  INVX0 U11713 ( .INP(n11626), .ZN(n11624) );
  NOR2X0 U11714 ( .IN1(n11627), .IN2(n11628), .QN(n11626) );
  NOR2X0 U11715 ( .IN1(WX11213), .IN2(n9274), .QN(n11628) );
  INVX0 U11716 ( .INP(n11629), .ZN(n11627) );
  NAND2X0 U11717 ( .IN1(n9274), .IN2(WX11213), .QN(n11629) );
  NOR2X0 U11718 ( .IN1(n11630), .IN2(n11631), .QN(n11625) );
  INVX0 U11719 ( .INP(n11632), .ZN(n11631) );
  NAND2X0 U11720 ( .IN1(n9273), .IN2(WX11085), .QN(n11632) );
  NOR2X0 U11721 ( .IN1(WX11085), .IN2(n9273), .QN(n11630) );
  NOR2X0 U11722 ( .IN1(n11633), .IN2(n11634), .QN(n11616) );
  NOR2X0 U11723 ( .IN1(DFF_1519_n1), .IN2(n9965), .QN(n11634) );
  NOR2X0 U11724 ( .IN1(n9997), .IN2(n11096), .QN(n11633) );
  NAND2X0 U11725 ( .IN1(n10195), .IN2(n8337), .QN(n11096) );
  NAND2X0 U11726 ( .IN1(n11635), .IN2(n11636), .QN(WX9725) );
  NOR2X0 U11727 ( .IN1(n11637), .IN2(n11638), .QN(n11636) );
  NOR2X0 U11728 ( .IN1(n9943), .IN2(n11639), .QN(n11638) );
  NOR2X0 U11729 ( .IN1(n10949), .IN2(n9908), .QN(n11637) );
  NOR2X0 U11730 ( .IN1(n11640), .IN2(n11641), .QN(n10949) );
  INVX0 U11731 ( .INP(n11642), .ZN(n11641) );
  NAND2X0 U11732 ( .IN1(n11643), .IN2(n11644), .QN(n11642) );
  NOR2X0 U11733 ( .IN1(n11644), .IN2(n11643), .QN(n11640) );
  NAND2X0 U11734 ( .IN1(n11645), .IN2(n11646), .QN(n11643) );
  NAND2X0 U11735 ( .IN1(n9020), .IN2(n11647), .QN(n11646) );
  INVX0 U11736 ( .INP(n11648), .ZN(n11645) );
  NOR2X0 U11737 ( .IN1(n11647), .IN2(n9020), .QN(n11648) );
  NOR2X0 U11738 ( .IN1(n11649), .IN2(n11650), .QN(n11647) );
  INVX0 U11739 ( .INP(n11651), .ZN(n11650) );
  NAND2X0 U11740 ( .IN1(n18472), .IN2(WX11211), .QN(n11651) );
  NOR2X0 U11741 ( .IN1(WX11211), .IN2(n18472), .QN(n11649) );
  NOR2X0 U11742 ( .IN1(n11652), .IN2(n11653), .QN(n11644) );
  INVX0 U11743 ( .INP(n11654), .ZN(n11653) );
  NAND2X0 U11744 ( .IN1(n9019), .IN2(n10019), .QN(n11654) );
  NOR2X0 U11745 ( .IN1(n10003), .IN2(n9019), .QN(n11652) );
  NOR2X0 U11746 ( .IN1(n11656), .IN2(n11657), .QN(n11635) );
  NOR2X0 U11747 ( .IN1(DFF_1520_n1), .IN2(n9965), .QN(n11657) );
  NOR2X0 U11748 ( .IN1(n9997), .IN2(n11097), .QN(n11656) );
  NAND2X0 U11749 ( .IN1(n10195), .IN2(n8338), .QN(n11097) );
  NAND2X0 U11750 ( .IN1(n11658), .IN2(n11659), .QN(WX9723) );
  NOR2X0 U11751 ( .IN1(n11660), .IN2(n11661), .QN(n11659) );
  NOR2X0 U11752 ( .IN1(n11662), .IN2(n9928), .QN(n11661) );
  NOR2X0 U11753 ( .IN1(n10958), .IN2(n9908), .QN(n11660) );
  NOR2X0 U11754 ( .IN1(n11663), .IN2(n11664), .QN(n10958) );
  INVX0 U11755 ( .INP(n11665), .ZN(n11664) );
  NAND2X0 U11756 ( .IN1(n11666), .IN2(n11667), .QN(n11665) );
  NOR2X0 U11757 ( .IN1(n11667), .IN2(n11666), .QN(n11663) );
  NAND2X0 U11758 ( .IN1(n11668), .IN2(n11669), .QN(n11666) );
  NAND2X0 U11759 ( .IN1(n9022), .IN2(n11670), .QN(n11669) );
  INVX0 U11760 ( .INP(n11671), .ZN(n11668) );
  NOR2X0 U11761 ( .IN1(n11670), .IN2(n9022), .QN(n11671) );
  NOR2X0 U11762 ( .IN1(n11672), .IN2(n11673), .QN(n11670) );
  INVX0 U11763 ( .INP(n11674), .ZN(n11673) );
  NAND2X0 U11764 ( .IN1(n18471), .IN2(WX11209), .QN(n11674) );
  NOR2X0 U11765 ( .IN1(WX11209), .IN2(n18471), .QN(n11672) );
  NOR2X0 U11766 ( .IN1(n11675), .IN2(n11676), .QN(n11667) );
  INVX0 U11767 ( .INP(n11677), .ZN(n11676) );
  NAND2X0 U11768 ( .IN1(n9021), .IN2(n10016), .QN(n11677) );
  NOR2X0 U11769 ( .IN1(n10003), .IN2(n9021), .QN(n11675) );
  NOR2X0 U11770 ( .IN1(n11678), .IN2(n11679), .QN(n11658) );
  NOR2X0 U11771 ( .IN1(DFF_1521_n1), .IN2(n9965), .QN(n11679) );
  NOR2X0 U11772 ( .IN1(n9997), .IN2(n11098), .QN(n11678) );
  NAND2X0 U11773 ( .IN1(n10195), .IN2(n8339), .QN(n11098) );
  NAND2X0 U11774 ( .IN1(n11680), .IN2(n11681), .QN(WX9721) );
  NOR2X0 U11775 ( .IN1(n11682), .IN2(n11683), .QN(n11681) );
  NOR2X0 U11776 ( .IN1(n9943), .IN2(n11684), .QN(n11683) );
  NOR2X0 U11777 ( .IN1(n10967), .IN2(n9908), .QN(n11682) );
  NOR2X0 U11778 ( .IN1(n11685), .IN2(n11686), .QN(n10967) );
  INVX0 U11779 ( .INP(n11687), .ZN(n11686) );
  NAND2X0 U11780 ( .IN1(n11688), .IN2(n11689), .QN(n11687) );
  NOR2X0 U11781 ( .IN1(n11689), .IN2(n11688), .QN(n11685) );
  NAND2X0 U11782 ( .IN1(n11690), .IN2(n11691), .QN(n11688) );
  NAND2X0 U11783 ( .IN1(n9024), .IN2(n11692), .QN(n11691) );
  INVX0 U11784 ( .INP(n11693), .ZN(n11690) );
  NOR2X0 U11785 ( .IN1(n11692), .IN2(n9024), .QN(n11693) );
  NOR2X0 U11786 ( .IN1(n11694), .IN2(n11695), .QN(n11692) );
  INVX0 U11787 ( .INP(n11696), .ZN(n11695) );
  NAND2X0 U11788 ( .IN1(n18470), .IN2(WX11207), .QN(n11696) );
  NOR2X0 U11789 ( .IN1(WX11207), .IN2(n18470), .QN(n11694) );
  NOR2X0 U11790 ( .IN1(n11697), .IN2(n11698), .QN(n11689) );
  INVX0 U11791 ( .INP(n11699), .ZN(n11698) );
  NAND2X0 U11792 ( .IN1(n9023), .IN2(n10016), .QN(n11699) );
  NOR2X0 U11793 ( .IN1(n10003), .IN2(n9023), .QN(n11697) );
  NOR2X0 U11794 ( .IN1(n11700), .IN2(n11701), .QN(n11680) );
  NOR2X0 U11795 ( .IN1(DFF_1522_n1), .IN2(n9965), .QN(n11701) );
  NOR2X0 U11796 ( .IN1(n9997), .IN2(n11099), .QN(n11700) );
  NAND2X0 U11797 ( .IN1(n10195), .IN2(n8340), .QN(n11099) );
  NAND2X0 U11798 ( .IN1(n11702), .IN2(n11703), .QN(WX9719) );
  NOR2X0 U11799 ( .IN1(n11704), .IN2(n11705), .QN(n11703) );
  NOR2X0 U11800 ( .IN1(n11706), .IN2(n9928), .QN(n11705) );
  INVX0 U11801 ( .INP(n11707), .ZN(n11704) );
  NAND2X0 U11802 ( .IN1(n2153), .IN2(n10975), .QN(n11707) );
  NOR2X0 U11803 ( .IN1(n11708), .IN2(n11709), .QN(n10975) );
  INVX0 U11804 ( .INP(n11710), .ZN(n11709) );
  NAND2X0 U11805 ( .IN1(n11711), .IN2(n11712), .QN(n11710) );
  NOR2X0 U11806 ( .IN1(n11712), .IN2(n11711), .QN(n11708) );
  NAND2X0 U11807 ( .IN1(n11713), .IN2(n11714), .QN(n11711) );
  NAND2X0 U11808 ( .IN1(n11715), .IN2(WX11141), .QN(n11714) );
  NAND2X0 U11809 ( .IN1(n11716), .IN2(n11717), .QN(n11715) );
  NAND2X0 U11810 ( .IN1(test_so97), .IN2(WX11077), .QN(n11717) );
  NAND2X0 U11811 ( .IN1(n9025), .IN2(n9839), .QN(n11716) );
  NAND2X0 U11812 ( .IN1(n9026), .IN2(n11718), .QN(n11713) );
  NOR2X0 U11813 ( .IN1(n11719), .IN2(n11720), .QN(n11718) );
  NOR2X0 U11814 ( .IN1(test_so97), .IN2(WX11077), .QN(n11720) );
  NOR2X0 U11815 ( .IN1(n9025), .IN2(n9839), .QN(n11719) );
  NOR2X0 U11816 ( .IN1(n11721), .IN2(n11722), .QN(n11712) );
  INVX0 U11817 ( .INP(n11723), .ZN(n11722) );
  NAND2X0 U11818 ( .IN1(n18469), .IN2(n10016), .QN(n11723) );
  NOR2X0 U11819 ( .IN1(n10003), .IN2(n18469), .QN(n11721) );
  NOR2X0 U11820 ( .IN1(n11724), .IN2(n11725), .QN(n11702) );
  NOR2X0 U11821 ( .IN1(n9975), .IN2(n9863), .QN(n11725) );
  NOR2X0 U11822 ( .IN1(n9997), .IN2(n11100), .QN(n11724) );
  NAND2X0 U11823 ( .IN1(n10195), .IN2(n8341), .QN(n11100) );
  NAND2X0 U11824 ( .IN1(n11726), .IN2(n11727), .QN(WX9717) );
  NOR2X0 U11825 ( .IN1(n11728), .IN2(n11729), .QN(n11727) );
  NOR2X0 U11826 ( .IN1(n9943), .IN2(n11730), .QN(n11729) );
  NOR2X0 U11827 ( .IN1(n10984), .IN2(n9908), .QN(n11728) );
  NOR2X0 U11828 ( .IN1(n11731), .IN2(n11732), .QN(n10984) );
  INVX0 U11829 ( .INP(n11733), .ZN(n11732) );
  NAND2X0 U11830 ( .IN1(n11734), .IN2(n11735), .QN(n11733) );
  NOR2X0 U11831 ( .IN1(n11735), .IN2(n11734), .QN(n11731) );
  NAND2X0 U11832 ( .IN1(n11736), .IN2(n11737), .QN(n11734) );
  NAND2X0 U11833 ( .IN1(n9028), .IN2(n11738), .QN(n11737) );
  INVX0 U11834 ( .INP(n11739), .ZN(n11736) );
  NOR2X0 U11835 ( .IN1(n11738), .IN2(n9028), .QN(n11739) );
  NOR2X0 U11836 ( .IN1(n11740), .IN2(n11741), .QN(n11738) );
  INVX0 U11837 ( .INP(n11742), .ZN(n11741) );
  NAND2X0 U11838 ( .IN1(n18468), .IN2(WX11203), .QN(n11742) );
  NOR2X0 U11839 ( .IN1(WX11203), .IN2(n18468), .QN(n11740) );
  NOR2X0 U11840 ( .IN1(n11743), .IN2(n11744), .QN(n11735) );
  INVX0 U11841 ( .INP(n11745), .ZN(n11744) );
  NAND2X0 U11842 ( .IN1(n9027), .IN2(n10016), .QN(n11745) );
  NOR2X0 U11843 ( .IN1(n10003), .IN2(n9027), .QN(n11743) );
  NOR2X0 U11844 ( .IN1(n11746), .IN2(n11747), .QN(n11726) );
  NOR2X0 U11845 ( .IN1(DFF_1524_n1), .IN2(n9965), .QN(n11747) );
  NOR2X0 U11846 ( .IN1(n9997), .IN2(n11101), .QN(n11746) );
  NAND2X0 U11847 ( .IN1(n10195), .IN2(n8342), .QN(n11101) );
  NAND2X0 U11848 ( .IN1(n11748), .IN2(n11749), .QN(WX9715) );
  NOR2X0 U11849 ( .IN1(n11750), .IN2(n11751), .QN(n11749) );
  NOR2X0 U11850 ( .IN1(n11752), .IN2(n9928), .QN(n11751) );
  INVX0 U11851 ( .INP(n11753), .ZN(n11750) );
  NAND2X0 U11852 ( .IN1(n2153), .IN2(n10992), .QN(n11753) );
  NOR2X0 U11853 ( .IN1(n11754), .IN2(n11755), .QN(n10992) );
  INVX0 U11854 ( .INP(n11756), .ZN(n11755) );
  NAND2X0 U11855 ( .IN1(n11757), .IN2(n11758), .QN(n11756) );
  NOR2X0 U11856 ( .IN1(n11758), .IN2(n11757), .QN(n11754) );
  NAND2X0 U11857 ( .IN1(n11759), .IN2(n11760), .QN(n11757) );
  NAND2X0 U11858 ( .IN1(n9535), .IN2(n11761), .QN(n11760) );
  INVX0 U11859 ( .INP(n11762), .ZN(n11761) );
  NAND2X0 U11860 ( .IN1(n11762), .IN2(WX11201), .QN(n11759) );
  NAND2X0 U11861 ( .IN1(n11763), .IN2(n11764), .QN(n11762) );
  INVX0 U11862 ( .INP(n11765), .ZN(n11764) );
  NOR2X0 U11863 ( .IN1(n9865), .IN2(n18467), .QN(n11765) );
  NAND2X0 U11864 ( .IN1(n18467), .IN2(n9865), .QN(n11763) );
  NOR2X0 U11865 ( .IN1(n11766), .IN2(n11767), .QN(n11758) );
  INVX0 U11866 ( .INP(n11768), .ZN(n11767) );
  NAND2X0 U11867 ( .IN1(n9029), .IN2(n10016), .QN(n11768) );
  NOR2X0 U11868 ( .IN1(n10004), .IN2(n9029), .QN(n11766) );
  NOR2X0 U11869 ( .IN1(n11769), .IN2(n11770), .QN(n11748) );
  NOR2X0 U11870 ( .IN1(DFF_1525_n1), .IN2(n9965), .QN(n11770) );
  NOR2X0 U11871 ( .IN1(n9997), .IN2(n11102), .QN(n11769) );
  NAND2X0 U11872 ( .IN1(n10195), .IN2(n8343), .QN(n11102) );
  NAND2X0 U11873 ( .IN1(n11771), .IN2(n11772), .QN(WX9713) );
  NOR2X0 U11874 ( .IN1(n11773), .IN2(n11774), .QN(n11772) );
  NOR2X0 U11875 ( .IN1(n11775), .IN2(n9928), .QN(n11774) );
  NOR2X0 U11876 ( .IN1(n11001), .IN2(n9908), .QN(n11773) );
  NOR2X0 U11877 ( .IN1(n11776), .IN2(n11777), .QN(n11001) );
  INVX0 U11878 ( .INP(n11778), .ZN(n11777) );
  NAND2X0 U11879 ( .IN1(n11779), .IN2(n11780), .QN(n11778) );
  NOR2X0 U11880 ( .IN1(n11780), .IN2(n11779), .QN(n11776) );
  NAND2X0 U11881 ( .IN1(n11781), .IN2(n11782), .QN(n11779) );
  NAND2X0 U11882 ( .IN1(n9031), .IN2(n11783), .QN(n11782) );
  INVX0 U11883 ( .INP(n11784), .ZN(n11781) );
  NOR2X0 U11884 ( .IN1(n11783), .IN2(n9031), .QN(n11784) );
  NOR2X0 U11885 ( .IN1(n11785), .IN2(n11786), .QN(n11783) );
  INVX0 U11886 ( .INP(n11787), .ZN(n11786) );
  NAND2X0 U11887 ( .IN1(n18466), .IN2(WX11199), .QN(n11787) );
  NOR2X0 U11888 ( .IN1(WX11199), .IN2(n18466), .QN(n11785) );
  NOR2X0 U11889 ( .IN1(n11788), .IN2(n11789), .QN(n11780) );
  INVX0 U11890 ( .INP(n11790), .ZN(n11789) );
  NAND2X0 U11891 ( .IN1(n9030), .IN2(n10016), .QN(n11790) );
  NOR2X0 U11892 ( .IN1(n10003), .IN2(n9030), .QN(n11788) );
  NOR2X0 U11893 ( .IN1(n11791), .IN2(n11792), .QN(n11771) );
  NOR2X0 U11894 ( .IN1(DFF_1526_n1), .IN2(n9965), .QN(n11792) );
  NOR2X0 U11895 ( .IN1(n9997), .IN2(n11103), .QN(n11791) );
  NAND2X0 U11896 ( .IN1(test_so78), .IN2(n10215), .QN(n11103) );
  NAND2X0 U11897 ( .IN1(n11793), .IN2(n11794), .QN(WX9711) );
  NOR2X0 U11898 ( .IN1(n11795), .IN2(n11796), .QN(n11794) );
  NOR2X0 U11899 ( .IN1(n11797), .IN2(n9929), .QN(n11796) );
  INVX0 U11900 ( .INP(n11798), .ZN(n11795) );
  NAND2X0 U11901 ( .IN1(n2153), .IN2(n11009), .QN(n11798) );
  NOR2X0 U11902 ( .IN1(n11799), .IN2(n11800), .QN(n11009) );
  INVX0 U11903 ( .INP(n11801), .ZN(n11800) );
  NAND2X0 U11904 ( .IN1(n11802), .IN2(n11803), .QN(n11801) );
  NOR2X0 U11905 ( .IN1(n11803), .IN2(n11802), .QN(n11799) );
  NAND2X0 U11906 ( .IN1(n11804), .IN2(n11805), .QN(n11802) );
  NAND2X0 U11907 ( .IN1(n9533), .IN2(n11806), .QN(n11805) );
  INVX0 U11908 ( .INP(n11807), .ZN(n11806) );
  NAND2X0 U11909 ( .IN1(n11807), .IN2(WX11197), .QN(n11804) );
  NAND2X0 U11910 ( .IN1(n11808), .IN2(n11809), .QN(n11807) );
  INVX0 U11911 ( .INP(n11810), .ZN(n11809) );
  NOR2X0 U11912 ( .IN1(n9866), .IN2(n18465), .QN(n11810) );
  NAND2X0 U11913 ( .IN1(n18465), .IN2(n9866), .QN(n11808) );
  NOR2X0 U11914 ( .IN1(n11811), .IN2(n11812), .QN(n11803) );
  INVX0 U11915 ( .INP(n11813), .ZN(n11812) );
  NAND2X0 U11916 ( .IN1(n9032), .IN2(n10016), .QN(n11813) );
  NOR2X0 U11917 ( .IN1(n10003), .IN2(n9032), .QN(n11811) );
  NOR2X0 U11918 ( .IN1(n11814), .IN2(n11815), .QN(n11793) );
  NOR2X0 U11919 ( .IN1(DFF_1527_n1), .IN2(n9965), .QN(n11815) );
  NOR2X0 U11920 ( .IN1(n9997), .IN2(n11104), .QN(n11814) );
  NAND2X0 U11921 ( .IN1(n10195), .IN2(n8346), .QN(n11104) );
  NAND2X0 U11922 ( .IN1(n11816), .IN2(n11817), .QN(WX9709) );
  NOR2X0 U11923 ( .IN1(n11818), .IN2(n11819), .QN(n11817) );
  NOR2X0 U11924 ( .IN1(n11820), .IN2(n9929), .QN(n11819) );
  NOR2X0 U11925 ( .IN1(n11018), .IN2(n9908), .QN(n11818) );
  NOR2X0 U11926 ( .IN1(n11821), .IN2(n11822), .QN(n11018) );
  INVX0 U11927 ( .INP(n11823), .ZN(n11822) );
  NAND2X0 U11928 ( .IN1(n11824), .IN2(n11825), .QN(n11823) );
  NOR2X0 U11929 ( .IN1(n11825), .IN2(n11824), .QN(n11821) );
  NAND2X0 U11930 ( .IN1(n11826), .IN2(n11827), .QN(n11824) );
  NAND2X0 U11931 ( .IN1(n9034), .IN2(n11828), .QN(n11827) );
  INVX0 U11932 ( .INP(n11829), .ZN(n11826) );
  NOR2X0 U11933 ( .IN1(n11828), .IN2(n9034), .QN(n11829) );
  NOR2X0 U11934 ( .IN1(n11830), .IN2(n11831), .QN(n11828) );
  INVX0 U11935 ( .INP(n11832), .ZN(n11831) );
  NAND2X0 U11936 ( .IN1(n18464), .IN2(WX11195), .QN(n11832) );
  NOR2X0 U11937 ( .IN1(WX11195), .IN2(n18464), .QN(n11830) );
  NOR2X0 U11938 ( .IN1(n11833), .IN2(n11834), .QN(n11825) );
  INVX0 U11939 ( .INP(n11835), .ZN(n11834) );
  NAND2X0 U11940 ( .IN1(n9033), .IN2(n10016), .QN(n11835) );
  NOR2X0 U11941 ( .IN1(n10004), .IN2(n9033), .QN(n11833) );
  NOR2X0 U11942 ( .IN1(n11836), .IN2(n11837), .QN(n11816) );
  NOR2X0 U11943 ( .IN1(DFF_1528_n1), .IN2(n9965), .QN(n11837) );
  NOR2X0 U11944 ( .IN1(n9997), .IN2(n11105), .QN(n11836) );
  NAND2X0 U11945 ( .IN1(n10195), .IN2(n8347), .QN(n11105) );
  NAND2X0 U11946 ( .IN1(n11838), .IN2(n11839), .QN(WX9707) );
  NOR2X0 U11947 ( .IN1(n11840), .IN2(n11841), .QN(n11839) );
  NOR2X0 U11948 ( .IN1(n11842), .IN2(n9929), .QN(n11841) );
  INVX0 U11949 ( .INP(n11843), .ZN(n11840) );
  NAND2X0 U11950 ( .IN1(n2153), .IN2(n11026), .QN(n11843) );
  NOR2X0 U11951 ( .IN1(n11844), .IN2(n11845), .QN(n11026) );
  INVX0 U11952 ( .INP(n11846), .ZN(n11845) );
  NAND2X0 U11953 ( .IN1(n11847), .IN2(n11848), .QN(n11846) );
  NOR2X0 U11954 ( .IN1(n11848), .IN2(n11847), .QN(n11844) );
  NAND2X0 U11955 ( .IN1(n11849), .IN2(n11850), .QN(n11847) );
  NAND2X0 U11956 ( .IN1(n11851), .IN2(WX11129), .QN(n11850) );
  NAND2X0 U11957 ( .IN1(n11852), .IN2(n11853), .QN(n11851) );
  NAND2X0 U11958 ( .IN1(test_so91), .IN2(WX11065), .QN(n11853) );
  NAND2X0 U11959 ( .IN1(n9035), .IN2(n9846), .QN(n11852) );
  NAND2X0 U11960 ( .IN1(n9036), .IN2(n11854), .QN(n11849) );
  NOR2X0 U11961 ( .IN1(n11855), .IN2(n11856), .QN(n11854) );
  NOR2X0 U11962 ( .IN1(test_so91), .IN2(WX11065), .QN(n11856) );
  NOR2X0 U11963 ( .IN1(n9035), .IN2(n9846), .QN(n11855) );
  INVX0 U11964 ( .INP(n11857), .ZN(n11848) );
  NAND2X0 U11965 ( .IN1(n11858), .IN2(n11859), .QN(n11857) );
  NAND2X0 U11966 ( .IN1(n9531), .IN2(n10016), .QN(n11859) );
  NAND2X0 U11967 ( .IN1(TM1), .IN2(WX11193), .QN(n11858) );
  NOR2X0 U11968 ( .IN1(n11860), .IN2(n11861), .QN(n11838) );
  NOR2X0 U11969 ( .IN1(DFF_1529_n1), .IN2(n9965), .QN(n11861) );
  NOR2X0 U11970 ( .IN1(n9996), .IN2(n11106), .QN(n11860) );
  NAND2X0 U11971 ( .IN1(n10194), .IN2(n8348), .QN(n11106) );
  NAND2X0 U11972 ( .IN1(n11862), .IN2(n11863), .QN(WX9705) );
  NOR2X0 U11973 ( .IN1(n11864), .IN2(n11865), .QN(n11863) );
  NOR2X0 U11974 ( .IN1(n11866), .IN2(n9929), .QN(n11865) );
  NOR2X0 U11975 ( .IN1(n11035), .IN2(n9908), .QN(n11864) );
  NOR2X0 U11976 ( .IN1(n11867), .IN2(n11868), .QN(n11035) );
  INVX0 U11977 ( .INP(n11869), .ZN(n11868) );
  NAND2X0 U11978 ( .IN1(n11870), .IN2(n11871), .QN(n11869) );
  NOR2X0 U11979 ( .IN1(n11871), .IN2(n11870), .QN(n11867) );
  NAND2X0 U11980 ( .IN1(n11872), .IN2(n11873), .QN(n11870) );
  NAND2X0 U11981 ( .IN1(n9038), .IN2(n11874), .QN(n11873) );
  INVX0 U11982 ( .INP(n11875), .ZN(n11872) );
  NOR2X0 U11983 ( .IN1(n11874), .IN2(n9038), .QN(n11875) );
  NOR2X0 U11984 ( .IN1(n11876), .IN2(n11877), .QN(n11874) );
  INVX0 U11985 ( .INP(n11878), .ZN(n11877) );
  NAND2X0 U11986 ( .IN1(n18463), .IN2(WX11191), .QN(n11878) );
  NOR2X0 U11987 ( .IN1(WX11191), .IN2(n18463), .QN(n11876) );
  NOR2X0 U11988 ( .IN1(n11879), .IN2(n11880), .QN(n11871) );
  INVX0 U11989 ( .INP(n11881), .ZN(n11880) );
  NAND2X0 U11990 ( .IN1(n9037), .IN2(n10016), .QN(n11881) );
  NOR2X0 U11991 ( .IN1(n10003), .IN2(n9037), .QN(n11879) );
  NOR2X0 U11992 ( .IN1(n11882), .IN2(n11883), .QN(n11862) );
  NOR2X0 U11993 ( .IN1(DFF_1530_n1), .IN2(n9965), .QN(n11883) );
  NOR2X0 U11994 ( .IN1(n9996), .IN2(n11107), .QN(n11882) );
  NAND2X0 U11995 ( .IN1(n10194), .IN2(n8349), .QN(n11107) );
  NAND2X0 U11996 ( .IN1(n11884), .IN2(n11885), .QN(WX9703) );
  NOR2X0 U11997 ( .IN1(n11886), .IN2(n11887), .QN(n11885) );
  NOR2X0 U11998 ( .IN1(n11888), .IN2(n9929), .QN(n11887) );
  NOR2X0 U11999 ( .IN1(n11044), .IN2(n9908), .QN(n11886) );
  NOR2X0 U12000 ( .IN1(n11889), .IN2(n11890), .QN(n11044) );
  INVX0 U12001 ( .INP(n11891), .ZN(n11890) );
  NAND2X0 U12002 ( .IN1(n11892), .IN2(n11893), .QN(n11891) );
  NOR2X0 U12003 ( .IN1(n11893), .IN2(n11892), .QN(n11889) );
  NAND2X0 U12004 ( .IN1(n11894), .IN2(n11895), .QN(n11892) );
  NAND2X0 U12005 ( .IN1(n9040), .IN2(n11896), .QN(n11895) );
  INVX0 U12006 ( .INP(n11897), .ZN(n11894) );
  NOR2X0 U12007 ( .IN1(n11896), .IN2(n9040), .QN(n11897) );
  NOR2X0 U12008 ( .IN1(n11898), .IN2(n11899), .QN(n11896) );
  INVX0 U12009 ( .INP(n11900), .ZN(n11899) );
  NAND2X0 U12010 ( .IN1(n18462), .IN2(WX11189), .QN(n11900) );
  NOR2X0 U12011 ( .IN1(WX11189), .IN2(n18462), .QN(n11898) );
  NOR2X0 U12012 ( .IN1(n11901), .IN2(n11902), .QN(n11893) );
  INVX0 U12013 ( .INP(n11903), .ZN(n11902) );
  NAND2X0 U12014 ( .IN1(n9039), .IN2(n10016), .QN(n11903) );
  NOR2X0 U12015 ( .IN1(n10004), .IN2(n9039), .QN(n11901) );
  NOR2X0 U12016 ( .IN1(n11904), .IN2(n11905), .QN(n11884) );
  NOR2X0 U12017 ( .IN1(DFF_1531_n1), .IN2(n9964), .QN(n11905) );
  NOR2X0 U12018 ( .IN1(n9996), .IN2(n11108), .QN(n11904) );
  NAND2X0 U12019 ( .IN1(n10194), .IN2(n8350), .QN(n11108) );
  NAND2X0 U12020 ( .IN1(n11906), .IN2(n11907), .QN(WX9701) );
  NOR2X0 U12021 ( .IN1(n11908), .IN2(n11909), .QN(n11907) );
  NOR2X0 U12022 ( .IN1(n11910), .IN2(n9929), .QN(n11909) );
  NOR2X0 U12023 ( .IN1(n11053), .IN2(n9908), .QN(n11908) );
  NOR2X0 U12024 ( .IN1(n11911), .IN2(n11912), .QN(n11053) );
  INVX0 U12025 ( .INP(n11913), .ZN(n11912) );
  NAND2X0 U12026 ( .IN1(n11914), .IN2(n11915), .QN(n11913) );
  NOR2X0 U12027 ( .IN1(n11915), .IN2(n11914), .QN(n11911) );
  NAND2X0 U12028 ( .IN1(n11916), .IN2(n11917), .QN(n11914) );
  NAND2X0 U12029 ( .IN1(n9042), .IN2(n11918), .QN(n11917) );
  INVX0 U12030 ( .INP(n11919), .ZN(n11916) );
  NOR2X0 U12031 ( .IN1(n11918), .IN2(n9042), .QN(n11919) );
  NOR2X0 U12032 ( .IN1(n11920), .IN2(n11921), .QN(n11918) );
  INVX0 U12033 ( .INP(n11922), .ZN(n11921) );
  NAND2X0 U12034 ( .IN1(n18461), .IN2(WX11187), .QN(n11922) );
  NOR2X0 U12035 ( .IN1(WX11187), .IN2(n18461), .QN(n11920) );
  NOR2X0 U12036 ( .IN1(n11923), .IN2(n11924), .QN(n11915) );
  INVX0 U12037 ( .INP(n11925), .ZN(n11924) );
  NAND2X0 U12038 ( .IN1(n9041), .IN2(n10016), .QN(n11925) );
  NOR2X0 U12039 ( .IN1(n10004), .IN2(n9041), .QN(n11923) );
  NOR2X0 U12040 ( .IN1(n11926), .IN2(n11927), .QN(n11906) );
  NOR2X0 U12041 ( .IN1(DFF_1532_n1), .IN2(n9967), .QN(n11927) );
  NOR2X0 U12042 ( .IN1(n9996), .IN2(n11109), .QN(n11926) );
  NAND2X0 U12043 ( .IN1(n10194), .IN2(n8351), .QN(n11109) );
  NAND2X0 U12044 ( .IN1(n11928), .IN2(n11929), .QN(WX9699) );
  NOR2X0 U12045 ( .IN1(n11930), .IN2(n11931), .QN(n11929) );
  NOR2X0 U12046 ( .IN1(n11932), .IN2(n9929), .QN(n11931) );
  NOR2X0 U12047 ( .IN1(n11062), .IN2(n9908), .QN(n11930) );
  NOR2X0 U12048 ( .IN1(n11933), .IN2(n11934), .QN(n11062) );
  INVX0 U12049 ( .INP(n11935), .ZN(n11934) );
  NAND2X0 U12050 ( .IN1(n11936), .IN2(n11937), .QN(n11935) );
  NOR2X0 U12051 ( .IN1(n11937), .IN2(n11936), .QN(n11933) );
  NAND2X0 U12052 ( .IN1(n11938), .IN2(n11939), .QN(n11936) );
  NAND2X0 U12053 ( .IN1(n9044), .IN2(n11940), .QN(n11939) );
  INVX0 U12054 ( .INP(n11941), .ZN(n11938) );
  NOR2X0 U12055 ( .IN1(n11940), .IN2(n9044), .QN(n11941) );
  NOR2X0 U12056 ( .IN1(n11942), .IN2(n11943), .QN(n11940) );
  INVX0 U12057 ( .INP(n11944), .ZN(n11943) );
  NAND2X0 U12058 ( .IN1(n18460), .IN2(WX11185), .QN(n11944) );
  NOR2X0 U12059 ( .IN1(WX11185), .IN2(n18460), .QN(n11942) );
  NOR2X0 U12060 ( .IN1(n11945), .IN2(n11946), .QN(n11937) );
  INVX0 U12061 ( .INP(n11947), .ZN(n11946) );
  NAND2X0 U12062 ( .IN1(n9043), .IN2(n10015), .QN(n11947) );
  NOR2X0 U12063 ( .IN1(n10004), .IN2(n9043), .QN(n11945) );
  NOR2X0 U12064 ( .IN1(n11948), .IN2(n11949), .QN(n11928) );
  NOR2X0 U12065 ( .IN1(DFF_1533_n1), .IN2(n9964), .QN(n11949) );
  NOR2X0 U12066 ( .IN1(n9996), .IN2(n11110), .QN(n11948) );
  NAND2X0 U12067 ( .IN1(n10194), .IN2(n8352), .QN(n11110) );
  NAND2X0 U12068 ( .IN1(n11950), .IN2(n11951), .QN(WX9697) );
  NOR2X0 U12069 ( .IN1(n11952), .IN2(n11953), .QN(n11951) );
  NOR2X0 U12070 ( .IN1(n11954), .IN2(n9929), .QN(n11953) );
  NOR2X0 U12071 ( .IN1(n11071), .IN2(n9908), .QN(n11952) );
  NOR2X0 U12072 ( .IN1(n11955), .IN2(n11956), .QN(n11071) );
  INVX0 U12073 ( .INP(n11957), .ZN(n11956) );
  NAND2X0 U12074 ( .IN1(n11958), .IN2(n11959), .QN(n11957) );
  NOR2X0 U12075 ( .IN1(n11959), .IN2(n11958), .QN(n11955) );
  NAND2X0 U12076 ( .IN1(n11960), .IN2(n11961), .QN(n11958) );
  NAND2X0 U12077 ( .IN1(n9046), .IN2(n11962), .QN(n11961) );
  INVX0 U12078 ( .INP(n11963), .ZN(n11960) );
  NOR2X0 U12079 ( .IN1(n11962), .IN2(n9046), .QN(n11963) );
  NOR2X0 U12080 ( .IN1(n11964), .IN2(n11965), .QN(n11962) );
  INVX0 U12081 ( .INP(n11966), .ZN(n11965) );
  NAND2X0 U12082 ( .IN1(n18459), .IN2(WX11183), .QN(n11966) );
  NOR2X0 U12083 ( .IN1(WX11183), .IN2(n18459), .QN(n11964) );
  NOR2X0 U12084 ( .IN1(n11967), .IN2(n11968), .QN(n11959) );
  INVX0 U12085 ( .INP(n11969), .ZN(n11968) );
  NAND2X0 U12086 ( .IN1(n9045), .IN2(n10015), .QN(n11969) );
  NOR2X0 U12087 ( .IN1(n10004), .IN2(n9045), .QN(n11967) );
  NOR2X0 U12088 ( .IN1(n11970), .IN2(n11971), .QN(n11950) );
  NOR2X0 U12089 ( .IN1(DFF_1534_n1), .IN2(n9964), .QN(n11971) );
  NOR2X0 U12090 ( .IN1(n9996), .IN2(n11111), .QN(n11970) );
  NAND2X0 U12091 ( .IN1(n10194), .IN2(n8353), .QN(n11111) );
  NAND2X0 U12092 ( .IN1(n11972), .IN2(n11973), .QN(WX9695) );
  NOR2X0 U12093 ( .IN1(n11974), .IN2(n11975), .QN(n11973) );
  NOR2X0 U12094 ( .IN1(n9942), .IN2(n11976), .QN(n11975) );
  NOR2X0 U12095 ( .IN1(n11080), .IN2(n9909), .QN(n11974) );
  NOR2X0 U12096 ( .IN1(n11977), .IN2(n11978), .QN(n11080) );
  INVX0 U12097 ( .INP(n11979), .ZN(n11978) );
  NAND2X0 U12098 ( .IN1(n11980), .IN2(n11981), .QN(n11979) );
  NOR2X0 U12099 ( .IN1(n11981), .IN2(n11980), .QN(n11977) );
  NAND2X0 U12100 ( .IN1(n11982), .IN2(n11983), .QN(n11980) );
  NAND2X0 U12101 ( .IN1(n9004), .IN2(n11984), .QN(n11983) );
  INVX0 U12102 ( .INP(n11985), .ZN(n11982) );
  NOR2X0 U12103 ( .IN1(n11984), .IN2(n9004), .QN(n11985) );
  NOR2X0 U12104 ( .IN1(n11986), .IN2(n11987), .QN(n11984) );
  INVX0 U12105 ( .INP(n11988), .ZN(n11987) );
  NAND2X0 U12106 ( .IN1(n18458), .IN2(WX11181), .QN(n11988) );
  NOR2X0 U12107 ( .IN1(WX11181), .IN2(n18458), .QN(n11986) );
  NOR2X0 U12108 ( .IN1(n11989), .IN2(n11990), .QN(n11981) );
  INVX0 U12109 ( .INP(n11991), .ZN(n11990) );
  NAND2X0 U12110 ( .IN1(n9003), .IN2(n10015), .QN(n11991) );
  NOR2X0 U12111 ( .IN1(n10004), .IN2(n9003), .QN(n11989) );
  NOR2X0 U12112 ( .IN1(n11992), .IN2(n11993), .QN(n11972) );
  NOR2X0 U12113 ( .IN1(n9489), .IN2(n11994), .QN(n11993) );
  NOR2X0 U12114 ( .IN1(DFF_1535_n1), .IN2(n9964), .QN(n11992) );
  INVX0 U12115 ( .INP(n11995), .ZN(WX9597) );
  NAND2X0 U12116 ( .IN1(n10194), .IN2(n9489), .QN(n11995) );
  NOR2X0 U12117 ( .IN1(n10321), .IN2(n11996), .QN(WX9084) );
  NAND2X0 U12118 ( .IN1(n11997), .IN2(n11998), .QN(n11996) );
  INVX0 U12119 ( .INP(n11999), .ZN(n11998) );
  NOR2X0 U12120 ( .IN1(WX8595), .IN2(DFF_1342_n1), .QN(n11999) );
  NAND2X0 U12121 ( .IN1(DFF_1342_n1), .IN2(WX8595), .QN(n11997) );
  NOR2X0 U12122 ( .IN1(n10321), .IN2(n12000), .QN(WX9082) );
  NAND2X0 U12123 ( .IN1(n12001), .IN2(n12002), .QN(n12000) );
  INVX0 U12124 ( .INP(n12003), .ZN(n12002) );
  NOR2X0 U12125 ( .IN1(WX8597), .IN2(DFF_1341_n1), .QN(n12003) );
  NAND2X0 U12126 ( .IN1(DFF_1341_n1), .IN2(WX8597), .QN(n12001) );
  NOR2X0 U12127 ( .IN1(n10321), .IN2(n12004), .QN(WX9080) );
  NAND2X0 U12128 ( .IN1(n12005), .IN2(n12006), .QN(n12004) );
  INVX0 U12129 ( .INP(n12007), .ZN(n12006) );
  NOR2X0 U12130 ( .IN1(WX8599), .IN2(DFF_1340_n1), .QN(n12007) );
  NAND2X0 U12131 ( .IN1(DFF_1340_n1), .IN2(WX8599), .QN(n12005) );
  NOR2X0 U12132 ( .IN1(n10321), .IN2(n12008), .QN(WX9078) );
  NAND2X0 U12133 ( .IN1(n12009), .IN2(n12010), .QN(n12008) );
  INVX0 U12134 ( .INP(n12011), .ZN(n12010) );
  NOR2X0 U12135 ( .IN1(WX8601), .IN2(DFF_1339_n1), .QN(n12011) );
  NAND2X0 U12136 ( .IN1(DFF_1339_n1), .IN2(WX8601), .QN(n12009) );
  NOR2X0 U12137 ( .IN1(n10321), .IN2(n12012), .QN(WX9076) );
  NAND2X0 U12138 ( .IN1(n12013), .IN2(n12014), .QN(n12012) );
  INVX0 U12139 ( .INP(n12015), .ZN(n12014) );
  NOR2X0 U12140 ( .IN1(WX8603), .IN2(DFF_1338_n1), .QN(n12015) );
  NAND2X0 U12141 ( .IN1(DFF_1338_n1), .IN2(WX8603), .QN(n12013) );
  NOR2X0 U12142 ( .IN1(n10321), .IN2(n12016), .QN(WX9074) );
  NOR2X0 U12143 ( .IN1(n12017), .IN2(n12018), .QN(n12016) );
  INVX0 U12144 ( .INP(n12019), .ZN(n12018) );
  NAND2X0 U12145 ( .IN1(n9828), .IN2(DFF_1337_n1), .QN(n12019) );
  NOR2X0 U12146 ( .IN1(DFF_1337_n1), .IN2(n9828), .QN(n12017) );
  NOR2X0 U12147 ( .IN1(n10321), .IN2(n12020), .QN(WX9072) );
  NOR2X0 U12148 ( .IN1(n12021), .IN2(n12022), .QN(n12020) );
  NOR2X0 U12149 ( .IN1(test_so77), .IN2(WX8607), .QN(n12022) );
  NOR2X0 U12150 ( .IN1(n9582), .IN2(n9853), .QN(n12021) );
  NOR2X0 U12151 ( .IN1(n10321), .IN2(n12023), .QN(WX9070) );
  NAND2X0 U12152 ( .IN1(n12024), .IN2(n12025), .QN(n12023) );
  INVX0 U12153 ( .INP(n12026), .ZN(n12025) );
  NOR2X0 U12154 ( .IN1(WX8609), .IN2(DFF_1335_n1), .QN(n12026) );
  NAND2X0 U12155 ( .IN1(DFF_1335_n1), .IN2(WX8609), .QN(n12024) );
  NOR2X0 U12156 ( .IN1(n10321), .IN2(n12027), .QN(WX9068) );
  NAND2X0 U12157 ( .IN1(n12028), .IN2(n12029), .QN(n12027) );
  INVX0 U12158 ( .INP(n12030), .ZN(n12029) );
  NOR2X0 U12159 ( .IN1(WX8611), .IN2(DFF_1334_n1), .QN(n12030) );
  NAND2X0 U12160 ( .IN1(DFF_1334_n1), .IN2(WX8611), .QN(n12028) );
  NOR2X0 U12161 ( .IN1(n10322), .IN2(n12031), .QN(WX9066) );
  NAND2X0 U12162 ( .IN1(n12032), .IN2(n12033), .QN(n12031) );
  INVX0 U12163 ( .INP(n12034), .ZN(n12033) );
  NOR2X0 U12164 ( .IN1(WX8613), .IN2(DFF_1333_n1), .QN(n12034) );
  NAND2X0 U12165 ( .IN1(DFF_1333_n1), .IN2(WX8613), .QN(n12032) );
  NOR2X0 U12166 ( .IN1(n10322), .IN2(n12035), .QN(WX9064) );
  NAND2X0 U12167 ( .IN1(n12036), .IN2(n12037), .QN(n12035) );
  INVX0 U12168 ( .INP(n12038), .ZN(n12037) );
  NOR2X0 U12169 ( .IN1(WX8615), .IN2(DFF_1332_n1), .QN(n12038) );
  NAND2X0 U12170 ( .IN1(DFF_1332_n1), .IN2(WX8615), .QN(n12036) );
  NOR2X0 U12171 ( .IN1(n10322), .IN2(n12039), .QN(WX9062) );
  NAND2X0 U12172 ( .IN1(n12040), .IN2(n12041), .QN(n12039) );
  INVX0 U12173 ( .INP(n12042), .ZN(n12041) );
  NOR2X0 U12174 ( .IN1(WX8617), .IN2(DFF_1331_n1), .QN(n12042) );
  NAND2X0 U12175 ( .IN1(DFF_1331_n1), .IN2(WX8617), .QN(n12040) );
  NOR2X0 U12176 ( .IN1(n10322), .IN2(n12043), .QN(WX9060) );
  NAND2X0 U12177 ( .IN1(n12044), .IN2(n12045), .QN(n12043) );
  INVX0 U12178 ( .INP(n12046), .ZN(n12045) );
  NOR2X0 U12179 ( .IN1(WX8619), .IN2(DFF_1330_n1), .QN(n12046) );
  NAND2X0 U12180 ( .IN1(DFF_1330_n1), .IN2(WX8619), .QN(n12044) );
  NOR2X0 U12181 ( .IN1(n10322), .IN2(n12047), .QN(WX9058) );
  NAND2X0 U12182 ( .IN1(n12048), .IN2(n12049), .QN(n12047) );
  INVX0 U12183 ( .INP(n12050), .ZN(n12049) );
  NOR2X0 U12184 ( .IN1(WX8621), .IN2(DFF_1329_n1), .QN(n12050) );
  NAND2X0 U12185 ( .IN1(DFF_1329_n1), .IN2(WX8621), .QN(n12048) );
  NOR2X0 U12186 ( .IN1(n10322), .IN2(n12051), .QN(WX9056) );
  NAND2X0 U12187 ( .IN1(n12052), .IN2(n12053), .QN(n12051) );
  INVX0 U12188 ( .INP(n12054), .ZN(n12053) );
  NOR2X0 U12189 ( .IN1(WX8623), .IN2(DFF_1328_n1), .QN(n12054) );
  NAND2X0 U12190 ( .IN1(DFF_1328_n1), .IN2(WX8623), .QN(n12052) );
  NOR2X0 U12191 ( .IN1(n10322), .IN2(n12055), .QN(WX9054) );
  NOR2X0 U12192 ( .IN1(n12056), .IN2(n12057), .QN(n12055) );
  INVX0 U12193 ( .INP(n12058), .ZN(n12057) );
  NAND2X0 U12194 ( .IN1(CRC_OUT_3_15), .IN2(n12059), .QN(n12058) );
  NOR2X0 U12195 ( .IN1(n12059), .IN2(CRC_OUT_3_15), .QN(n12056) );
  NAND2X0 U12196 ( .IN1(n12060), .IN2(n12061), .QN(n12059) );
  NAND2X0 U12197 ( .IN1(n9502), .IN2(CRC_OUT_3_31), .QN(n12061) );
  NAND2X0 U12198 ( .IN1(DFF_1343_n1), .IN2(WX8625), .QN(n12060) );
  NOR2X0 U12199 ( .IN1(n10322), .IN2(n12062), .QN(WX9052) );
  NAND2X0 U12200 ( .IN1(n12063), .IN2(n12064), .QN(n12062) );
  INVX0 U12201 ( .INP(n12065), .ZN(n12064) );
  NOR2X0 U12202 ( .IN1(WX8627), .IN2(DFF_1326_n1), .QN(n12065) );
  NAND2X0 U12203 ( .IN1(DFF_1326_n1), .IN2(WX8627), .QN(n12063) );
  NOR2X0 U12204 ( .IN1(n10322), .IN2(n12066), .QN(WX9050) );
  NAND2X0 U12205 ( .IN1(n12067), .IN2(n12068), .QN(n12066) );
  INVX0 U12206 ( .INP(n12069), .ZN(n12068) );
  NOR2X0 U12207 ( .IN1(WX8629), .IN2(DFF_1325_n1), .QN(n12069) );
  NAND2X0 U12208 ( .IN1(DFF_1325_n1), .IN2(WX8629), .QN(n12067) );
  NOR2X0 U12209 ( .IN1(n10322), .IN2(n12070), .QN(WX9048) );
  NAND2X0 U12210 ( .IN1(n12071), .IN2(n12072), .QN(n12070) );
  INVX0 U12211 ( .INP(n12073), .ZN(n12072) );
  NOR2X0 U12212 ( .IN1(WX8631), .IN2(DFF_1324_n1), .QN(n12073) );
  NAND2X0 U12213 ( .IN1(DFF_1324_n1), .IN2(WX8631), .QN(n12071) );
  NOR2X0 U12214 ( .IN1(n10322), .IN2(n12074), .QN(WX9046) );
  NAND2X0 U12215 ( .IN1(n12075), .IN2(n12076), .QN(n12074) );
  INVX0 U12216 ( .INP(n12077), .ZN(n12076) );
  NOR2X0 U12217 ( .IN1(WX8633), .IN2(DFF_1323_n1), .QN(n12077) );
  NAND2X0 U12218 ( .IN1(DFF_1323_n1), .IN2(WX8633), .QN(n12075) );
  NOR2X0 U12219 ( .IN1(n10322), .IN2(n12078), .QN(WX9044) );
  NOR2X0 U12220 ( .IN1(n12079), .IN2(n12080), .QN(n12078) );
  INVX0 U12221 ( .INP(n12081), .ZN(n12080) );
  NAND2X0 U12222 ( .IN1(CRC_OUT_3_10), .IN2(n12082), .QN(n12081) );
  NOR2X0 U12223 ( .IN1(n12082), .IN2(CRC_OUT_3_10), .QN(n12079) );
  NAND2X0 U12224 ( .IN1(n12083), .IN2(n12084), .QN(n12082) );
  NAND2X0 U12225 ( .IN1(n9503), .IN2(CRC_OUT_3_31), .QN(n12084) );
  NAND2X0 U12226 ( .IN1(DFF_1343_n1), .IN2(WX8635), .QN(n12083) );
  NOR2X0 U12227 ( .IN1(n10322), .IN2(n12085), .QN(WX9042) );
  NAND2X0 U12228 ( .IN1(n12086), .IN2(n12087), .QN(n12085) );
  INVX0 U12229 ( .INP(n12088), .ZN(n12087) );
  NOR2X0 U12230 ( .IN1(WX8637), .IN2(DFF_1321_n1), .QN(n12088) );
  NAND2X0 U12231 ( .IN1(DFF_1321_n1), .IN2(WX8637), .QN(n12086) );
  NOR2X0 U12232 ( .IN1(n10323), .IN2(n12089), .QN(WX9040) );
  NOR2X0 U12233 ( .IN1(n12090), .IN2(n12091), .QN(n12089) );
  INVX0 U12234 ( .INP(n12092), .ZN(n12091) );
  NAND2X0 U12235 ( .IN1(n9834), .IN2(DFF_1320_n1), .QN(n12092) );
  NOR2X0 U12236 ( .IN1(DFF_1320_n1), .IN2(n9834), .QN(n12090) );
  NOR2X0 U12237 ( .IN1(n10323), .IN2(n12093), .QN(WX9038) );
  NOR2X0 U12238 ( .IN1(n12094), .IN2(n12095), .QN(n12093) );
  NOR2X0 U12239 ( .IN1(test_so76), .IN2(WX8641), .QN(n12095) );
  NOR2X0 U12240 ( .IN1(n9596), .IN2(n9852), .QN(n12094) );
  NOR2X0 U12241 ( .IN1(n10323), .IN2(n12096), .QN(WX9036) );
  NAND2X0 U12242 ( .IN1(n12097), .IN2(n12098), .QN(n12096) );
  INVX0 U12243 ( .INP(n12099), .ZN(n12098) );
  NOR2X0 U12244 ( .IN1(WX8643), .IN2(DFF_1318_n1), .QN(n12099) );
  NAND2X0 U12245 ( .IN1(DFF_1318_n1), .IN2(WX8643), .QN(n12097) );
  NOR2X0 U12246 ( .IN1(n10323), .IN2(n12100), .QN(WX9034) );
  NAND2X0 U12247 ( .IN1(n12101), .IN2(n12102), .QN(n12100) );
  INVX0 U12248 ( .INP(n12103), .ZN(n12102) );
  NOR2X0 U12249 ( .IN1(WX8645), .IN2(DFF_1317_n1), .QN(n12103) );
  NAND2X0 U12250 ( .IN1(DFF_1317_n1), .IN2(WX8645), .QN(n12101) );
  NOR2X0 U12251 ( .IN1(n10323), .IN2(n12104), .QN(WX9032) );
  NAND2X0 U12252 ( .IN1(n12105), .IN2(n12106), .QN(n12104) );
  INVX0 U12253 ( .INP(n12107), .ZN(n12106) );
  NOR2X0 U12254 ( .IN1(WX8647), .IN2(DFF_1316_n1), .QN(n12107) );
  NAND2X0 U12255 ( .IN1(DFF_1316_n1), .IN2(WX8647), .QN(n12105) );
  NOR2X0 U12256 ( .IN1(n10323), .IN2(n12108), .QN(WX9030) );
  NOR2X0 U12257 ( .IN1(n12109), .IN2(n12110), .QN(n12108) );
  INVX0 U12258 ( .INP(n12111), .ZN(n12110) );
  NAND2X0 U12259 ( .IN1(CRC_OUT_3_3), .IN2(n12112), .QN(n12111) );
  NOR2X0 U12260 ( .IN1(n12112), .IN2(CRC_OUT_3_3), .QN(n12109) );
  NAND2X0 U12261 ( .IN1(n12113), .IN2(n12114), .QN(n12112) );
  NAND2X0 U12262 ( .IN1(n9504), .IN2(CRC_OUT_3_31), .QN(n12114) );
  NAND2X0 U12263 ( .IN1(DFF_1343_n1), .IN2(WX8649), .QN(n12113) );
  NOR2X0 U12264 ( .IN1(n10323), .IN2(n12115), .QN(WX9028) );
  NAND2X0 U12265 ( .IN1(n12116), .IN2(n12117), .QN(n12115) );
  INVX0 U12266 ( .INP(n12118), .ZN(n12117) );
  NOR2X0 U12267 ( .IN1(WX8651), .IN2(DFF_1314_n1), .QN(n12118) );
  NAND2X0 U12268 ( .IN1(DFF_1314_n1), .IN2(WX8651), .QN(n12116) );
  NOR2X0 U12269 ( .IN1(n10323), .IN2(n12119), .QN(WX9026) );
  NAND2X0 U12270 ( .IN1(n12120), .IN2(n12121), .QN(n12119) );
  INVX0 U12271 ( .INP(n12122), .ZN(n12121) );
  NOR2X0 U12272 ( .IN1(WX8653), .IN2(DFF_1313_n1), .QN(n12122) );
  NAND2X0 U12273 ( .IN1(DFF_1313_n1), .IN2(WX8653), .QN(n12120) );
  NOR2X0 U12274 ( .IN1(n10323), .IN2(n12123), .QN(WX9024) );
  NAND2X0 U12275 ( .IN1(n12124), .IN2(n12125), .QN(n12123) );
  INVX0 U12276 ( .INP(n12126), .ZN(n12125) );
  NOR2X0 U12277 ( .IN1(WX8655), .IN2(DFF_1312_n1), .QN(n12126) );
  NAND2X0 U12278 ( .IN1(DFF_1312_n1), .IN2(WX8655), .QN(n12124) );
  NOR2X0 U12279 ( .IN1(n10323), .IN2(n12127), .QN(WX9022) );
  NAND2X0 U12280 ( .IN1(n12128), .IN2(n12129), .QN(n12127) );
  NAND2X0 U12281 ( .IN1(n9519), .IN2(CRC_OUT_3_31), .QN(n12129) );
  NAND2X0 U12282 ( .IN1(DFF_1343_n1), .IN2(WX8657), .QN(n12128) );
  NOR2X0 U12283 ( .IN1(n18442), .IN2(n10235), .QN(WX8496) );
  NOR2X0 U12284 ( .IN1(n18441), .IN2(n10235), .QN(WX8494) );
  NOR2X0 U12285 ( .IN1(n18440), .IN2(n10235), .QN(WX8492) );
  NOR2X0 U12286 ( .IN1(n18439), .IN2(n10235), .QN(WX8490) );
  NOR2X0 U12287 ( .IN1(n18438), .IN2(n10235), .QN(WX8488) );
  NOR2X0 U12288 ( .IN1(n18437), .IN2(n10235), .QN(WX8486) );
  NOR2X0 U12289 ( .IN1(n18436), .IN2(n10236), .QN(WX8484) );
  NOR2X0 U12290 ( .IN1(n18435), .IN2(n10236), .QN(WX8482) );
  NOR2X0 U12291 ( .IN1(n18434), .IN2(n10236), .QN(WX8480) );
  NOR2X0 U12292 ( .IN1(n18433), .IN2(n10236), .QN(WX8478) );
  NOR2X0 U12293 ( .IN1(n18432), .IN2(n10236), .QN(WX8476) );
  NOR2X0 U12294 ( .IN1(n18431), .IN2(n10236), .QN(WX8474) );
  NOR2X0 U12295 ( .IN1(n18430), .IN2(n10236), .QN(WX8472) );
  NOR2X0 U12296 ( .IN1(n18429), .IN2(n10236), .QN(WX8470) );
  NOR2X0 U12297 ( .IN1(n18428), .IN2(n10236), .QN(WX8468) );
  NOR2X0 U12298 ( .IN1(n18427), .IN2(n10236), .QN(WX8466) );
  NAND2X0 U12299 ( .IN1(n12130), .IN2(n12131), .QN(WX8464) );
  NOR2X0 U12300 ( .IN1(n12132), .IN2(n12133), .QN(n12131) );
  NOR2X0 U12301 ( .IN1(n12134), .IN2(n9929), .QN(n12133) );
  NOR2X0 U12302 ( .IN1(n11329), .IN2(n9909), .QN(n12132) );
  INVX0 U12303 ( .INP(n12135), .ZN(n11329) );
  NAND2X0 U12304 ( .IN1(n12136), .IN2(n12137), .QN(n12135) );
  NAND2X0 U12305 ( .IN1(n12138), .IN2(n12139), .QN(n12137) );
  NAND2X0 U12306 ( .IN1(n12140), .IN2(n12141), .QN(n12139) );
  NAND2X0 U12307 ( .IN1(n9276), .IN2(WX9758), .QN(n12141) );
  NAND2X0 U12308 ( .IN1(n9275), .IN2(WX9886), .QN(n12140) );
  NOR2X0 U12309 ( .IN1(n12142), .IN2(n12143), .QN(n12138) );
  NOR2X0 U12310 ( .IN1(n9518), .IN2(WX9822), .QN(n12143) );
  NOR2X0 U12311 ( .IN1(n3563), .IN2(WX9950), .QN(n12142) );
  NAND2X0 U12312 ( .IN1(n12144), .IN2(n12145), .QN(n12136) );
  NAND2X0 U12313 ( .IN1(n12146), .IN2(n12147), .QN(n12145) );
  NAND2X0 U12314 ( .IN1(n9518), .IN2(WX9822), .QN(n12147) );
  NAND2X0 U12315 ( .IN1(n3563), .IN2(WX9950), .QN(n12146) );
  NOR2X0 U12316 ( .IN1(n12148), .IN2(n12149), .QN(n12144) );
  NOR2X0 U12317 ( .IN1(n9276), .IN2(WX9758), .QN(n12149) );
  NOR2X0 U12318 ( .IN1(n9275), .IN2(WX9886), .QN(n12148) );
  NOR2X0 U12319 ( .IN1(n12150), .IN2(n12151), .QN(n12130) );
  NOR2X0 U12320 ( .IN1(DFF_1312_n1), .IN2(n9964), .QN(n12151) );
  NOR2X0 U12321 ( .IN1(n9996), .IN2(n11112), .QN(n12150) );
  NAND2X0 U12322 ( .IN1(test_so68), .IN2(n10215), .QN(n11112) );
  NAND2X0 U12323 ( .IN1(n12152), .IN2(n12153), .QN(WX8462) );
  NOR2X0 U12324 ( .IN1(n12154), .IN2(n12155), .QN(n12153) );
  NOR2X0 U12325 ( .IN1(n12156), .IN2(n9929), .QN(n12155) );
  NOR2X0 U12326 ( .IN1(n9923), .IN2(n11350), .QN(n12154) );
  NAND2X0 U12327 ( .IN1(n12157), .IN2(n12158), .QN(n11350) );
  INVX0 U12328 ( .INP(n12159), .ZN(n12158) );
  NOR2X0 U12329 ( .IN1(n12160), .IN2(n12161), .QN(n12159) );
  NAND2X0 U12330 ( .IN1(n12161), .IN2(n12160), .QN(n12157) );
  NOR2X0 U12331 ( .IN1(n12162), .IN2(n12163), .QN(n12160) );
  INVX0 U12332 ( .INP(n12164), .ZN(n12163) );
  NAND2X0 U12333 ( .IN1(test_so83), .IN2(WX9948), .QN(n12164) );
  NOR2X0 U12334 ( .IN1(WX9948), .IN2(test_so83), .QN(n12162) );
  NAND2X0 U12335 ( .IN1(n12165), .IN2(n12166), .QN(n12161) );
  NAND2X0 U12336 ( .IN1(n9278), .IN2(WX9756), .QN(n12166) );
  INVX0 U12337 ( .INP(n12167), .ZN(n12165) );
  NOR2X0 U12338 ( .IN1(WX9756), .IN2(n9278), .QN(n12167) );
  NOR2X0 U12339 ( .IN1(n12168), .IN2(n12169), .QN(n12152) );
  NOR2X0 U12340 ( .IN1(DFF_1313_n1), .IN2(n9964), .QN(n12169) );
  NOR2X0 U12341 ( .IN1(n9996), .IN2(n11113), .QN(n12168) );
  NAND2X0 U12342 ( .IN1(n10194), .IN2(n8381), .QN(n11113) );
  NAND2X0 U12343 ( .IN1(n12170), .IN2(n12171), .QN(WX8460) );
  NOR2X0 U12344 ( .IN1(n12172), .IN2(n12173), .QN(n12171) );
  NOR2X0 U12345 ( .IN1(n12174), .IN2(n9929), .QN(n12173) );
  NOR2X0 U12346 ( .IN1(n11369), .IN2(n9909), .QN(n12172) );
  INVX0 U12347 ( .INP(n12175), .ZN(n11369) );
  NAND2X0 U12348 ( .IN1(n12176), .IN2(n12177), .QN(n12175) );
  NAND2X0 U12349 ( .IN1(n12178), .IN2(n12179), .QN(n12177) );
  NAND2X0 U12350 ( .IN1(n12180), .IN2(n12181), .QN(n12179) );
  NAND2X0 U12351 ( .IN1(n9280), .IN2(WX9754), .QN(n12181) );
  NAND2X0 U12352 ( .IN1(n9279), .IN2(WX9882), .QN(n12180) );
  NOR2X0 U12353 ( .IN1(n12182), .IN2(n12183), .QN(n12178) );
  NOR2X0 U12354 ( .IN1(n9575), .IN2(WX9818), .QN(n12183) );
  NOR2X0 U12355 ( .IN1(n3567), .IN2(WX9946), .QN(n12182) );
  NAND2X0 U12356 ( .IN1(n12184), .IN2(n12185), .QN(n12176) );
  NAND2X0 U12357 ( .IN1(n12186), .IN2(n12187), .QN(n12185) );
  NAND2X0 U12358 ( .IN1(n9575), .IN2(WX9818), .QN(n12187) );
  NAND2X0 U12359 ( .IN1(n3567), .IN2(WX9946), .QN(n12186) );
  NOR2X0 U12360 ( .IN1(n12188), .IN2(n12189), .QN(n12184) );
  NOR2X0 U12361 ( .IN1(n9280), .IN2(WX9754), .QN(n12189) );
  NOR2X0 U12362 ( .IN1(n9279), .IN2(WX9882), .QN(n12188) );
  NOR2X0 U12363 ( .IN1(n12190), .IN2(n12191), .QN(n12170) );
  NOR2X0 U12364 ( .IN1(DFF_1314_n1), .IN2(n9964), .QN(n12191) );
  NOR2X0 U12365 ( .IN1(n9996), .IN2(n11114), .QN(n12190) );
  NAND2X0 U12366 ( .IN1(n10193), .IN2(n8382), .QN(n11114) );
  NAND2X0 U12367 ( .IN1(n12192), .IN2(n12193), .QN(WX8458) );
  NOR2X0 U12368 ( .IN1(n12194), .IN2(n12195), .QN(n12193) );
  NOR2X0 U12369 ( .IN1(n12196), .IN2(n9929), .QN(n12195) );
  NOR2X0 U12370 ( .IN1(n9923), .IN2(n11389), .QN(n12194) );
  NAND2X0 U12371 ( .IN1(n12197), .IN2(n12198), .QN(n11389) );
  INVX0 U12372 ( .INP(n12199), .ZN(n12198) );
  NOR2X0 U12373 ( .IN1(n12200), .IN2(n12201), .QN(n12199) );
  NAND2X0 U12374 ( .IN1(n12201), .IN2(n12200), .QN(n12197) );
  NOR2X0 U12375 ( .IN1(n12202), .IN2(n12203), .QN(n12200) );
  INVX0 U12376 ( .INP(n12204), .ZN(n12203) );
  NAND2X0 U12377 ( .IN1(test_so81), .IN2(WX9944), .QN(n12204) );
  NOR2X0 U12378 ( .IN1(WX9944), .IN2(test_so81), .QN(n12202) );
  NAND2X0 U12379 ( .IN1(n12205), .IN2(n12206), .QN(n12201) );
  NAND2X0 U12380 ( .IN1(n9281), .IN2(WX9816), .QN(n12206) );
  INVX0 U12381 ( .INP(n12207), .ZN(n12205) );
  NOR2X0 U12382 ( .IN1(WX9816), .IN2(n9281), .QN(n12207) );
  NOR2X0 U12383 ( .IN1(n12208), .IN2(n12209), .QN(n12192) );
  NOR2X0 U12384 ( .IN1(DFF_1315_n1), .IN2(n9964), .QN(n12209) );
  NOR2X0 U12385 ( .IN1(n9996), .IN2(n11115), .QN(n12208) );
  NAND2X0 U12386 ( .IN1(n10193), .IN2(n8383), .QN(n11115) );
  NAND2X0 U12387 ( .IN1(n12210), .IN2(n12211), .QN(WX8456) );
  NOR2X0 U12388 ( .IN1(n12212), .IN2(n12213), .QN(n12211) );
  NOR2X0 U12389 ( .IN1(n12214), .IN2(n9930), .QN(n12213) );
  NOR2X0 U12390 ( .IN1(n11408), .IN2(n9909), .QN(n12212) );
  INVX0 U12391 ( .INP(n12215), .ZN(n11408) );
  NAND2X0 U12392 ( .IN1(n12216), .IN2(n12217), .QN(n12215) );
  NAND2X0 U12393 ( .IN1(n12218), .IN2(n12219), .QN(n12217) );
  NAND2X0 U12394 ( .IN1(n12220), .IN2(n12221), .QN(n12219) );
  NAND2X0 U12395 ( .IN1(n9283), .IN2(WX9750), .QN(n12221) );
  NAND2X0 U12396 ( .IN1(n9282), .IN2(WX9878), .QN(n12220) );
  NOR2X0 U12397 ( .IN1(n12222), .IN2(n12223), .QN(n12218) );
  NOR2X0 U12398 ( .IN1(n9501), .IN2(WX9814), .QN(n12223) );
  NOR2X0 U12399 ( .IN1(n3571), .IN2(WX9942), .QN(n12222) );
  NAND2X0 U12400 ( .IN1(n12224), .IN2(n12225), .QN(n12216) );
  NAND2X0 U12401 ( .IN1(n12226), .IN2(n12227), .QN(n12225) );
  NAND2X0 U12402 ( .IN1(n9501), .IN2(WX9814), .QN(n12227) );
  NAND2X0 U12403 ( .IN1(n3571), .IN2(WX9942), .QN(n12226) );
  NOR2X0 U12404 ( .IN1(n12228), .IN2(n12229), .QN(n12224) );
  NOR2X0 U12405 ( .IN1(n9283), .IN2(WX9750), .QN(n12229) );
  NOR2X0 U12406 ( .IN1(n9282), .IN2(WX9878), .QN(n12228) );
  NOR2X0 U12407 ( .IN1(n12230), .IN2(n12231), .QN(n12210) );
  NOR2X0 U12408 ( .IN1(DFF_1316_n1), .IN2(n9964), .QN(n12231) );
  NOR2X0 U12409 ( .IN1(n9996), .IN2(n11116), .QN(n12230) );
  NAND2X0 U12410 ( .IN1(n10193), .IN2(n8384), .QN(n11116) );
  NAND2X0 U12411 ( .IN1(n12232), .IN2(n12233), .QN(WX8454) );
  NOR2X0 U12412 ( .IN1(n12234), .IN2(n12235), .QN(n12233) );
  NOR2X0 U12413 ( .IN1(n12236), .IN2(n9930), .QN(n12235) );
  NOR2X0 U12414 ( .IN1(n11428), .IN2(n9909), .QN(n12234) );
  INVX0 U12415 ( .INP(n12237), .ZN(n11428) );
  NAND2X0 U12416 ( .IN1(n12238), .IN2(n12239), .QN(n12237) );
  NAND2X0 U12417 ( .IN1(n12240), .IN2(n12241), .QN(n12239) );
  NAND2X0 U12418 ( .IN1(n12242), .IN2(n12243), .QN(n12241) );
  NAND2X0 U12419 ( .IN1(n9285), .IN2(WX9748), .QN(n12243) );
  NAND2X0 U12420 ( .IN1(n9284), .IN2(WX9876), .QN(n12242) );
  NOR2X0 U12421 ( .IN1(n12244), .IN2(n12245), .QN(n12240) );
  NOR2X0 U12422 ( .IN1(n9573), .IN2(WX9812), .QN(n12245) );
  NOR2X0 U12423 ( .IN1(n3573), .IN2(WX9940), .QN(n12244) );
  NAND2X0 U12424 ( .IN1(n12246), .IN2(n12247), .QN(n12238) );
  NAND2X0 U12425 ( .IN1(n12248), .IN2(n12249), .QN(n12247) );
  NAND2X0 U12426 ( .IN1(n9573), .IN2(WX9812), .QN(n12249) );
  NAND2X0 U12427 ( .IN1(n3573), .IN2(WX9940), .QN(n12248) );
  NOR2X0 U12428 ( .IN1(n12250), .IN2(n12251), .QN(n12246) );
  NOR2X0 U12429 ( .IN1(n9285), .IN2(WX9748), .QN(n12251) );
  NOR2X0 U12430 ( .IN1(n9284), .IN2(WX9876), .QN(n12250) );
  NOR2X0 U12431 ( .IN1(n12252), .IN2(n12253), .QN(n12232) );
  NOR2X0 U12432 ( .IN1(DFF_1317_n1), .IN2(n9964), .QN(n12253) );
  NOR2X0 U12433 ( .IN1(n9996), .IN2(n11117), .QN(n12252) );
  NAND2X0 U12434 ( .IN1(n10193), .IN2(n8385), .QN(n11117) );
  NAND2X0 U12435 ( .IN1(n12254), .IN2(n12255), .QN(WX8452) );
  NOR2X0 U12436 ( .IN1(n12256), .IN2(n12257), .QN(n12255) );
  NOR2X0 U12437 ( .IN1(n12258), .IN2(n9930), .QN(n12257) );
  NOR2X0 U12438 ( .IN1(n11447), .IN2(n9909), .QN(n12256) );
  INVX0 U12439 ( .INP(n12259), .ZN(n11447) );
  NAND2X0 U12440 ( .IN1(n12260), .IN2(n12261), .QN(n12259) );
  NAND2X0 U12441 ( .IN1(n12262), .IN2(n12263), .QN(n12261) );
  NAND2X0 U12442 ( .IN1(n12264), .IN2(n12265), .QN(n12263) );
  NAND2X0 U12443 ( .IN1(n9287), .IN2(WX9746), .QN(n12265) );
  NAND2X0 U12444 ( .IN1(n9286), .IN2(WX9874), .QN(n12264) );
  NOR2X0 U12445 ( .IN1(n12266), .IN2(n12267), .QN(n12262) );
  NOR2X0 U12446 ( .IN1(n9572), .IN2(WX9810), .QN(n12267) );
  NOR2X0 U12447 ( .IN1(n3575), .IN2(WX9938), .QN(n12266) );
  NAND2X0 U12448 ( .IN1(n12268), .IN2(n12269), .QN(n12260) );
  NAND2X0 U12449 ( .IN1(n12270), .IN2(n12271), .QN(n12269) );
  NAND2X0 U12450 ( .IN1(n9572), .IN2(WX9810), .QN(n12271) );
  NAND2X0 U12451 ( .IN1(n3575), .IN2(WX9938), .QN(n12270) );
  NOR2X0 U12452 ( .IN1(n12272), .IN2(n12273), .QN(n12268) );
  NOR2X0 U12453 ( .IN1(n9287), .IN2(WX9746), .QN(n12273) );
  NOR2X0 U12454 ( .IN1(n9286), .IN2(WX9874), .QN(n12272) );
  NOR2X0 U12455 ( .IN1(n12274), .IN2(n12275), .QN(n12254) );
  NOR2X0 U12456 ( .IN1(DFF_1318_n1), .IN2(n9964), .QN(n12275) );
  NOR2X0 U12457 ( .IN1(n9995), .IN2(n11118), .QN(n12274) );
  NAND2X0 U12458 ( .IN1(n10193), .IN2(n8386), .QN(n11118) );
  NAND2X0 U12459 ( .IN1(n12276), .IN2(n12277), .QN(WX8450) );
  NOR2X0 U12460 ( .IN1(n12278), .IN2(n12279), .QN(n12277) );
  NOR2X0 U12461 ( .IN1(n12280), .IN2(n9930), .QN(n12279) );
  NOR2X0 U12462 ( .IN1(n11467), .IN2(n9909), .QN(n12278) );
  INVX0 U12463 ( .INP(n12281), .ZN(n11467) );
  NAND2X0 U12464 ( .IN1(n12282), .IN2(n12283), .QN(n12281) );
  NAND2X0 U12465 ( .IN1(n12284), .IN2(n12285), .QN(n12283) );
  NAND2X0 U12466 ( .IN1(n12286), .IN2(n12287), .QN(n12285) );
  NAND2X0 U12467 ( .IN1(n9289), .IN2(WX9744), .QN(n12287) );
  NAND2X0 U12468 ( .IN1(n9288), .IN2(WX9872), .QN(n12286) );
  NOR2X0 U12469 ( .IN1(n12288), .IN2(n12289), .QN(n12284) );
  NOR2X0 U12470 ( .IN1(n9571), .IN2(WX9808), .QN(n12289) );
  NOR2X0 U12471 ( .IN1(n3577), .IN2(WX9936), .QN(n12288) );
  NAND2X0 U12472 ( .IN1(n12290), .IN2(n12291), .QN(n12282) );
  NAND2X0 U12473 ( .IN1(n12292), .IN2(n12293), .QN(n12291) );
  NAND2X0 U12474 ( .IN1(n9571), .IN2(WX9808), .QN(n12293) );
  NAND2X0 U12475 ( .IN1(n3577), .IN2(WX9936), .QN(n12292) );
  NOR2X0 U12476 ( .IN1(n12294), .IN2(n12295), .QN(n12290) );
  NOR2X0 U12477 ( .IN1(n9289), .IN2(WX9744), .QN(n12295) );
  NOR2X0 U12478 ( .IN1(n9288), .IN2(WX9872), .QN(n12294) );
  NOR2X0 U12479 ( .IN1(n12296), .IN2(n12297), .QN(n12276) );
  NOR2X0 U12480 ( .IN1(n9975), .IN2(n9852), .QN(n12297) );
  NOR2X0 U12481 ( .IN1(n9995), .IN2(n11119), .QN(n12296) );
  NAND2X0 U12482 ( .IN1(n10193), .IN2(n8387), .QN(n11119) );
  NAND2X0 U12483 ( .IN1(n12298), .IN2(n12299), .QN(WX8448) );
  NOR2X0 U12484 ( .IN1(n12300), .IN2(n12301), .QN(n12299) );
  NOR2X0 U12485 ( .IN1(n12302), .IN2(n9930), .QN(n12301) );
  NOR2X0 U12486 ( .IN1(n11486), .IN2(n9909), .QN(n12300) );
  INVX0 U12487 ( .INP(n12303), .ZN(n11486) );
  NAND2X0 U12488 ( .IN1(n12304), .IN2(n12305), .QN(n12303) );
  NAND2X0 U12489 ( .IN1(n12306), .IN2(n12307), .QN(n12305) );
  NAND2X0 U12490 ( .IN1(n12308), .IN2(n12309), .QN(n12307) );
  NAND2X0 U12491 ( .IN1(n9291), .IN2(WX9742), .QN(n12309) );
  NAND2X0 U12492 ( .IN1(n9290), .IN2(WX9870), .QN(n12308) );
  NOR2X0 U12493 ( .IN1(n12310), .IN2(n12311), .QN(n12306) );
  NOR2X0 U12494 ( .IN1(n9570), .IN2(WX9806), .QN(n12311) );
  NOR2X0 U12495 ( .IN1(n3579), .IN2(WX9934), .QN(n12310) );
  NAND2X0 U12496 ( .IN1(n12312), .IN2(n12313), .QN(n12304) );
  NAND2X0 U12497 ( .IN1(n12314), .IN2(n12315), .QN(n12313) );
  NAND2X0 U12498 ( .IN1(n9570), .IN2(WX9806), .QN(n12315) );
  NAND2X0 U12499 ( .IN1(n3579), .IN2(WX9934), .QN(n12314) );
  NOR2X0 U12500 ( .IN1(n12316), .IN2(n12317), .QN(n12312) );
  NOR2X0 U12501 ( .IN1(n9291), .IN2(WX9742), .QN(n12317) );
  NOR2X0 U12502 ( .IN1(n9290), .IN2(WX9870), .QN(n12316) );
  NOR2X0 U12503 ( .IN1(n12318), .IN2(n12319), .QN(n12298) );
  NOR2X0 U12504 ( .IN1(DFF_1320_n1), .IN2(n9963), .QN(n12319) );
  NOR2X0 U12505 ( .IN1(n9995), .IN2(n11120), .QN(n12318) );
  NAND2X0 U12506 ( .IN1(n10193), .IN2(n8388), .QN(n11120) );
  NAND2X0 U12507 ( .IN1(n12320), .IN2(n12321), .QN(WX8446) );
  NOR2X0 U12508 ( .IN1(n12322), .IN2(n12323), .QN(n12321) );
  NOR2X0 U12509 ( .IN1(n9943), .IN2(n12324), .QN(n12323) );
  NOR2X0 U12510 ( .IN1(n11506), .IN2(n9909), .QN(n12322) );
  INVX0 U12511 ( .INP(n12325), .ZN(n11506) );
  NAND2X0 U12512 ( .IN1(n12326), .IN2(n12327), .QN(n12325) );
  NAND2X0 U12513 ( .IN1(n12328), .IN2(n12329), .QN(n12327) );
  NAND2X0 U12514 ( .IN1(n12330), .IN2(n12331), .QN(n12329) );
  NAND2X0 U12515 ( .IN1(n9293), .IN2(WX9740), .QN(n12331) );
  NAND2X0 U12516 ( .IN1(n9292), .IN2(WX9868), .QN(n12330) );
  NOR2X0 U12517 ( .IN1(n12332), .IN2(n12333), .QN(n12328) );
  NOR2X0 U12518 ( .IN1(n9569), .IN2(WX9804), .QN(n12333) );
  NOR2X0 U12519 ( .IN1(n3581), .IN2(WX9932), .QN(n12332) );
  NAND2X0 U12520 ( .IN1(n12334), .IN2(n12335), .QN(n12326) );
  NAND2X0 U12521 ( .IN1(n12336), .IN2(n12337), .QN(n12335) );
  NAND2X0 U12522 ( .IN1(n9569), .IN2(WX9804), .QN(n12337) );
  NAND2X0 U12523 ( .IN1(n3581), .IN2(WX9932), .QN(n12336) );
  NOR2X0 U12524 ( .IN1(n12338), .IN2(n12339), .QN(n12334) );
  NOR2X0 U12525 ( .IN1(n9293), .IN2(WX9740), .QN(n12339) );
  NOR2X0 U12526 ( .IN1(n9292), .IN2(WX9868), .QN(n12338) );
  NOR2X0 U12527 ( .IN1(n12340), .IN2(n12341), .QN(n12320) );
  NOR2X0 U12528 ( .IN1(DFF_1321_n1), .IN2(n9963), .QN(n12341) );
  NOR2X0 U12529 ( .IN1(n9995), .IN2(n11121), .QN(n12340) );
  NAND2X0 U12530 ( .IN1(n10193), .IN2(n8389), .QN(n11121) );
  NAND2X0 U12531 ( .IN1(n12342), .IN2(n12343), .QN(WX8444) );
  NOR2X0 U12532 ( .IN1(n12344), .IN2(n12345), .QN(n12343) );
  NOR2X0 U12533 ( .IN1(n12346), .IN2(n9930), .QN(n12345) );
  NOR2X0 U12534 ( .IN1(n11525), .IN2(n9909), .QN(n12344) );
  INVX0 U12535 ( .INP(n12347), .ZN(n11525) );
  NAND2X0 U12536 ( .IN1(n12348), .IN2(n12349), .QN(n12347) );
  NAND2X0 U12537 ( .IN1(n12350), .IN2(n12351), .QN(n12349) );
  NAND2X0 U12538 ( .IN1(n12352), .IN2(n12353), .QN(n12351) );
  NAND2X0 U12539 ( .IN1(n9295), .IN2(WX9738), .QN(n12353) );
  NAND2X0 U12540 ( .IN1(n9294), .IN2(WX9866), .QN(n12352) );
  NOR2X0 U12541 ( .IN1(n12354), .IN2(n12355), .QN(n12350) );
  NOR2X0 U12542 ( .IN1(n9568), .IN2(WX9802), .QN(n12355) );
  NOR2X0 U12543 ( .IN1(n3583), .IN2(WX9930), .QN(n12354) );
  NAND2X0 U12544 ( .IN1(n12356), .IN2(n12357), .QN(n12348) );
  NAND2X0 U12545 ( .IN1(n12358), .IN2(n12359), .QN(n12357) );
  NAND2X0 U12546 ( .IN1(n9568), .IN2(WX9802), .QN(n12359) );
  NAND2X0 U12547 ( .IN1(n3583), .IN2(WX9930), .QN(n12358) );
  NOR2X0 U12548 ( .IN1(n12360), .IN2(n12361), .QN(n12356) );
  NOR2X0 U12549 ( .IN1(n9295), .IN2(WX9738), .QN(n12361) );
  NOR2X0 U12550 ( .IN1(n9294), .IN2(WX9866), .QN(n12360) );
  NOR2X0 U12551 ( .IN1(n12362), .IN2(n12363), .QN(n12342) );
  NOR2X0 U12552 ( .IN1(DFF_1322_n1), .IN2(n9963), .QN(n12363) );
  NOR2X0 U12553 ( .IN1(n9995), .IN2(n11122), .QN(n12362) );
  NAND2X0 U12554 ( .IN1(n10193), .IN2(n8390), .QN(n11122) );
  NAND2X0 U12555 ( .IN1(n12364), .IN2(n12365), .QN(WX8442) );
  NOR2X0 U12556 ( .IN1(n12366), .IN2(n12367), .QN(n12365) );
  NOR2X0 U12557 ( .IN1(n9941), .IN2(n12368), .QN(n12367) );
  NOR2X0 U12558 ( .IN1(n11544), .IN2(n9909), .QN(n12366) );
  INVX0 U12559 ( .INP(n12369), .ZN(n11544) );
  NAND2X0 U12560 ( .IN1(n12370), .IN2(n12371), .QN(n12369) );
  NAND2X0 U12561 ( .IN1(n12372), .IN2(n12373), .QN(n12371) );
  NAND2X0 U12562 ( .IN1(n12374), .IN2(n12375), .QN(n12373) );
  NAND2X0 U12563 ( .IN1(n9297), .IN2(WX9736), .QN(n12375) );
  NAND2X0 U12564 ( .IN1(n9296), .IN2(WX9864), .QN(n12374) );
  NOR2X0 U12565 ( .IN1(n12376), .IN2(n12377), .QN(n12372) );
  NOR2X0 U12566 ( .IN1(n9500), .IN2(WX9800), .QN(n12377) );
  NOR2X0 U12567 ( .IN1(n3585), .IN2(WX9928), .QN(n12376) );
  NAND2X0 U12568 ( .IN1(n12378), .IN2(n12379), .QN(n12370) );
  NAND2X0 U12569 ( .IN1(n12380), .IN2(n12381), .QN(n12379) );
  NAND2X0 U12570 ( .IN1(n9500), .IN2(WX9800), .QN(n12381) );
  NAND2X0 U12571 ( .IN1(n3585), .IN2(WX9928), .QN(n12380) );
  NOR2X0 U12572 ( .IN1(n12382), .IN2(n12383), .QN(n12378) );
  NOR2X0 U12573 ( .IN1(n9297), .IN2(WX9736), .QN(n12383) );
  NOR2X0 U12574 ( .IN1(n9296), .IN2(WX9864), .QN(n12382) );
  NOR2X0 U12575 ( .IN1(n12384), .IN2(n12385), .QN(n12364) );
  NOR2X0 U12576 ( .IN1(DFF_1323_n1), .IN2(n9963), .QN(n12385) );
  NOR2X0 U12577 ( .IN1(n9995), .IN2(n11123), .QN(n12384) );
  NAND2X0 U12578 ( .IN1(n10192), .IN2(n8391), .QN(n11123) );
  NAND2X0 U12579 ( .IN1(n12386), .IN2(n12387), .QN(WX8440) );
  NOR2X0 U12580 ( .IN1(n12388), .IN2(n12389), .QN(n12387) );
  NOR2X0 U12581 ( .IN1(n12390), .IN2(n9930), .QN(n12389) );
  NOR2X0 U12582 ( .IN1(n11563), .IN2(n9919), .QN(n12388) );
  INVX0 U12583 ( .INP(n12391), .ZN(n11563) );
  NAND2X0 U12584 ( .IN1(n12392), .IN2(n12393), .QN(n12391) );
  NAND2X0 U12585 ( .IN1(n12394), .IN2(n12395), .QN(n12393) );
  NAND2X0 U12586 ( .IN1(n12396), .IN2(n12397), .QN(n12395) );
  NAND2X0 U12587 ( .IN1(n9299), .IN2(WX9734), .QN(n12397) );
  NAND2X0 U12588 ( .IN1(n9298), .IN2(WX9862), .QN(n12396) );
  NOR2X0 U12589 ( .IN1(n12398), .IN2(n12399), .QN(n12394) );
  NOR2X0 U12590 ( .IN1(n9567), .IN2(WX9798), .QN(n12399) );
  NOR2X0 U12591 ( .IN1(n3587), .IN2(WX9926), .QN(n12398) );
  NAND2X0 U12592 ( .IN1(n12400), .IN2(n12401), .QN(n12392) );
  NAND2X0 U12593 ( .IN1(n12402), .IN2(n12403), .QN(n12401) );
  NAND2X0 U12594 ( .IN1(n9567), .IN2(WX9798), .QN(n12403) );
  NAND2X0 U12595 ( .IN1(n3587), .IN2(WX9926), .QN(n12402) );
  NOR2X0 U12596 ( .IN1(n12404), .IN2(n12405), .QN(n12400) );
  NOR2X0 U12597 ( .IN1(n9299), .IN2(WX9734), .QN(n12405) );
  NOR2X0 U12598 ( .IN1(n9298), .IN2(WX9862), .QN(n12404) );
  NOR2X0 U12599 ( .IN1(n12406), .IN2(n12407), .QN(n12386) );
  NOR2X0 U12600 ( .IN1(DFF_1324_n1), .IN2(n9963), .QN(n12407) );
  NOR2X0 U12601 ( .IN1(n9995), .IN2(n11124), .QN(n12406) );
  NAND2X0 U12602 ( .IN1(n10192), .IN2(n8392), .QN(n11124) );
  NAND2X0 U12603 ( .IN1(n12408), .IN2(n12409), .QN(WX8438) );
  NOR2X0 U12604 ( .IN1(n12410), .IN2(n12411), .QN(n12409) );
  NOR2X0 U12605 ( .IN1(n9943), .IN2(n12412), .QN(n12411) );
  NOR2X0 U12606 ( .IN1(n11582), .IN2(n9909), .QN(n12410) );
  INVX0 U12607 ( .INP(n12413), .ZN(n11582) );
  NAND2X0 U12608 ( .IN1(n12414), .IN2(n12415), .QN(n12413) );
  NAND2X0 U12609 ( .IN1(n12416), .IN2(n12417), .QN(n12415) );
  NAND2X0 U12610 ( .IN1(n12418), .IN2(n12419), .QN(n12417) );
  NAND2X0 U12611 ( .IN1(n9301), .IN2(WX9732), .QN(n12419) );
  NAND2X0 U12612 ( .IN1(n9300), .IN2(WX9860), .QN(n12418) );
  NOR2X0 U12613 ( .IN1(n12420), .IN2(n12421), .QN(n12416) );
  NOR2X0 U12614 ( .IN1(n9566), .IN2(WX9796), .QN(n12421) );
  NOR2X0 U12615 ( .IN1(n3589), .IN2(WX9924), .QN(n12420) );
  NAND2X0 U12616 ( .IN1(n12422), .IN2(n12423), .QN(n12414) );
  NAND2X0 U12617 ( .IN1(n12424), .IN2(n12425), .QN(n12423) );
  NAND2X0 U12618 ( .IN1(n9566), .IN2(WX9796), .QN(n12425) );
  NAND2X0 U12619 ( .IN1(n3589), .IN2(WX9924), .QN(n12424) );
  NOR2X0 U12620 ( .IN1(n12426), .IN2(n12427), .QN(n12422) );
  NOR2X0 U12621 ( .IN1(n9301), .IN2(WX9732), .QN(n12427) );
  NOR2X0 U12622 ( .IN1(n9300), .IN2(WX9860), .QN(n12426) );
  NOR2X0 U12623 ( .IN1(n12428), .IN2(n12429), .QN(n12408) );
  NOR2X0 U12624 ( .IN1(DFF_1325_n1), .IN2(n9963), .QN(n12429) );
  NOR2X0 U12625 ( .IN1(n9995), .IN2(n11125), .QN(n12428) );
  NAND2X0 U12626 ( .IN1(n10192), .IN2(n8393), .QN(n11125) );
  NAND2X0 U12627 ( .IN1(n12430), .IN2(n12431), .QN(WX8436) );
  NOR2X0 U12628 ( .IN1(n12432), .IN2(n12433), .QN(n12431) );
  NOR2X0 U12629 ( .IN1(n12434), .IN2(n9930), .QN(n12433) );
  NOR2X0 U12630 ( .IN1(n9922), .IN2(n11601), .QN(n12432) );
  NAND2X0 U12631 ( .IN1(n12435), .IN2(n12436), .QN(n11601) );
  INVX0 U12632 ( .INP(n12437), .ZN(n12436) );
  NOR2X0 U12633 ( .IN1(n12438), .IN2(n12439), .QN(n12437) );
  NAND2X0 U12634 ( .IN1(n12439), .IN2(n12438), .QN(n12435) );
  NOR2X0 U12635 ( .IN1(n12440), .IN2(n12441), .QN(n12438) );
  NOR2X0 U12636 ( .IN1(n9837), .IN2(n9303), .QN(n12441) );
  INVX0 U12637 ( .INP(n12442), .ZN(n12440) );
  NAND2X0 U12638 ( .IN1(n9303), .IN2(n9837), .QN(n12442) );
  NAND2X0 U12639 ( .IN1(n12443), .IN2(n12444), .QN(n12439) );
  NAND2X0 U12640 ( .IN1(n9302), .IN2(WX9794), .QN(n12444) );
  INVX0 U12641 ( .INP(n12445), .ZN(n12443) );
  NOR2X0 U12642 ( .IN1(WX9794), .IN2(n9302), .QN(n12445) );
  NOR2X0 U12643 ( .IN1(n12446), .IN2(n12447), .QN(n12430) );
  NOR2X0 U12644 ( .IN1(DFF_1326_n1), .IN2(n9963), .QN(n12447) );
  NOR2X0 U12645 ( .IN1(n9995), .IN2(n11126), .QN(n12446) );
  NAND2X0 U12646 ( .IN1(n10192), .IN2(n8394), .QN(n11126) );
  NAND2X0 U12647 ( .IN1(n12448), .IN2(n12449), .QN(WX8434) );
  NOR2X0 U12648 ( .IN1(n12450), .IN2(n12451), .QN(n12449) );
  NOR2X0 U12649 ( .IN1(n9941), .IN2(n12452), .QN(n12451) );
  NOR2X0 U12650 ( .IN1(n11620), .IN2(n9910), .QN(n12450) );
  INVX0 U12651 ( .INP(n12453), .ZN(n11620) );
  NAND2X0 U12652 ( .IN1(n12454), .IN2(n12455), .QN(n12453) );
  NAND2X0 U12653 ( .IN1(n12456), .IN2(n12457), .QN(n12455) );
  NAND2X0 U12654 ( .IN1(n12458), .IN2(n12459), .QN(n12457) );
  NAND2X0 U12655 ( .IN1(n9305), .IN2(WX9728), .QN(n12459) );
  NAND2X0 U12656 ( .IN1(n9304), .IN2(WX9856), .QN(n12458) );
  NOR2X0 U12657 ( .IN1(n12460), .IN2(n12461), .QN(n12456) );
  NOR2X0 U12658 ( .IN1(n9565), .IN2(WX9792), .QN(n12461) );
  NOR2X0 U12659 ( .IN1(n3593), .IN2(WX9920), .QN(n12460) );
  NAND2X0 U12660 ( .IN1(n12462), .IN2(n12463), .QN(n12454) );
  NAND2X0 U12661 ( .IN1(n12464), .IN2(n12465), .QN(n12463) );
  NAND2X0 U12662 ( .IN1(n9565), .IN2(WX9792), .QN(n12465) );
  NAND2X0 U12663 ( .IN1(n3593), .IN2(WX9920), .QN(n12464) );
  NOR2X0 U12664 ( .IN1(n12466), .IN2(n12467), .QN(n12462) );
  NOR2X0 U12665 ( .IN1(n9305), .IN2(WX9728), .QN(n12467) );
  NOR2X0 U12666 ( .IN1(n9304), .IN2(WX9856), .QN(n12466) );
  NOR2X0 U12667 ( .IN1(n12468), .IN2(n12469), .QN(n12448) );
  NOR2X0 U12668 ( .IN1(DFF_1327_n1), .IN2(n9963), .QN(n12469) );
  NOR2X0 U12669 ( .IN1(n9995), .IN2(n11127), .QN(n12468) );
  NAND2X0 U12670 ( .IN1(n10192), .IN2(n8395), .QN(n11127) );
  NAND2X0 U12671 ( .IN1(n12470), .IN2(n12471), .QN(WX8432) );
  NOR2X0 U12672 ( .IN1(n12472), .IN2(n12473), .QN(n12471) );
  NOR2X0 U12673 ( .IN1(n12474), .IN2(n9930), .QN(n12473) );
  NOR2X0 U12674 ( .IN1(n9924), .IN2(n11639), .QN(n12472) );
  NAND2X0 U12675 ( .IN1(n12475), .IN2(n12476), .QN(n11639) );
  NAND2X0 U12676 ( .IN1(n12477), .IN2(n12478), .QN(n12476) );
  INVX0 U12677 ( .INP(n12479), .ZN(n12475) );
  NOR2X0 U12678 ( .IN1(n12478), .IN2(n12477), .QN(n12479) );
  NAND2X0 U12679 ( .IN1(n12480), .IN2(n12481), .QN(n12477) );
  NAND2X0 U12680 ( .IN1(n9499), .IN2(n12482), .QN(n12481) );
  INVX0 U12681 ( .INP(n12483), .ZN(n12482) );
  NAND2X0 U12682 ( .IN1(n12483), .IN2(WX9918), .QN(n12480) );
  NAND2X0 U12683 ( .IN1(n12484), .IN2(n12485), .QN(n12483) );
  INVX0 U12684 ( .INP(n12486), .ZN(n12485) );
  NOR2X0 U12685 ( .IN1(n9867), .IN2(n18457), .QN(n12486) );
  NAND2X0 U12686 ( .IN1(n18457), .IN2(n9867), .QN(n12484) );
  NOR2X0 U12687 ( .IN1(n12487), .IN2(n12488), .QN(n12478) );
  INVX0 U12688 ( .INP(n12489), .ZN(n12488) );
  NAND2X0 U12689 ( .IN1(n9047), .IN2(n10015), .QN(n12489) );
  NOR2X0 U12690 ( .IN1(n10004), .IN2(n9047), .QN(n12487) );
  NOR2X0 U12691 ( .IN1(n12490), .IN2(n12491), .QN(n12470) );
  NOR2X0 U12692 ( .IN1(DFF_1328_n1), .IN2(n9963), .QN(n12491) );
  NOR2X0 U12693 ( .IN1(n9995), .IN2(n11128), .QN(n12490) );
  NAND2X0 U12694 ( .IN1(n10192), .IN2(n8396), .QN(n11128) );
  NAND2X0 U12695 ( .IN1(n12492), .IN2(n12493), .QN(WX8430) );
  NOR2X0 U12696 ( .IN1(n12494), .IN2(n12495), .QN(n12493) );
  NOR2X0 U12697 ( .IN1(n12496), .IN2(n9930), .QN(n12495) );
  NOR2X0 U12698 ( .IN1(n11662), .IN2(n9910), .QN(n12494) );
  NOR2X0 U12699 ( .IN1(n12497), .IN2(n12498), .QN(n11662) );
  INVX0 U12700 ( .INP(n12499), .ZN(n12498) );
  NAND2X0 U12701 ( .IN1(n12500), .IN2(n12501), .QN(n12499) );
  NOR2X0 U12702 ( .IN1(n12501), .IN2(n12500), .QN(n12497) );
  NAND2X0 U12703 ( .IN1(n12502), .IN2(n12503), .QN(n12500) );
  NAND2X0 U12704 ( .IN1(n9049), .IN2(n12504), .QN(n12503) );
  INVX0 U12705 ( .INP(n12505), .ZN(n12502) );
  NOR2X0 U12706 ( .IN1(n12504), .IN2(n9049), .QN(n12505) );
  NOR2X0 U12707 ( .IN1(n12506), .IN2(n12507), .QN(n12504) );
  INVX0 U12708 ( .INP(n12508), .ZN(n12507) );
  NAND2X0 U12709 ( .IN1(n18456), .IN2(WX9916), .QN(n12508) );
  NOR2X0 U12710 ( .IN1(WX9916), .IN2(n18456), .QN(n12506) );
  NOR2X0 U12711 ( .IN1(n12509), .IN2(n12510), .QN(n12501) );
  INVX0 U12712 ( .INP(n12511), .ZN(n12510) );
  NAND2X0 U12713 ( .IN1(n9048), .IN2(n10015), .QN(n12511) );
  NOR2X0 U12714 ( .IN1(n10004), .IN2(n9048), .QN(n12509) );
  NOR2X0 U12715 ( .IN1(n12512), .IN2(n12513), .QN(n12492) );
  NOR2X0 U12716 ( .IN1(DFF_1329_n1), .IN2(n9963), .QN(n12513) );
  NOR2X0 U12717 ( .IN1(n9995), .IN2(n11129), .QN(n12512) );
  NAND2X0 U12718 ( .IN1(test_so67), .IN2(n10215), .QN(n11129) );
  NAND2X0 U12719 ( .IN1(n12514), .IN2(n12515), .QN(WX8428) );
  NOR2X0 U12720 ( .IN1(n12516), .IN2(n12517), .QN(n12515) );
  NOR2X0 U12721 ( .IN1(n12518), .IN2(n9930), .QN(n12517) );
  NOR2X0 U12722 ( .IN1(n9923), .IN2(n11684), .QN(n12516) );
  NAND2X0 U12723 ( .IN1(n12519), .IN2(n12520), .QN(n11684) );
  NAND2X0 U12724 ( .IN1(n12521), .IN2(n12522), .QN(n12520) );
  INVX0 U12725 ( .INP(n12523), .ZN(n12519) );
  NOR2X0 U12726 ( .IN1(n12522), .IN2(n12521), .QN(n12523) );
  NAND2X0 U12727 ( .IN1(n12524), .IN2(n12525), .QN(n12521) );
  NAND2X0 U12728 ( .IN1(n9563), .IN2(n12526), .QN(n12525) );
  INVX0 U12729 ( .INP(n12527), .ZN(n12526) );
  NAND2X0 U12730 ( .IN1(n12527), .IN2(WX9914), .QN(n12524) );
  NAND2X0 U12731 ( .IN1(n12528), .IN2(n12529), .QN(n12527) );
  INVX0 U12732 ( .INP(n12530), .ZN(n12529) );
  NOR2X0 U12733 ( .IN1(n9868), .IN2(n18455), .QN(n12530) );
  NAND2X0 U12734 ( .IN1(n18455), .IN2(n9868), .QN(n12528) );
  NOR2X0 U12735 ( .IN1(n12531), .IN2(n12532), .QN(n12522) );
  INVX0 U12736 ( .INP(n12533), .ZN(n12532) );
  NAND2X0 U12737 ( .IN1(n9050), .IN2(n10015), .QN(n12533) );
  NOR2X0 U12738 ( .IN1(n10004), .IN2(n9050), .QN(n12531) );
  NOR2X0 U12739 ( .IN1(n12534), .IN2(n12535), .QN(n12514) );
  NOR2X0 U12740 ( .IN1(DFF_1330_n1), .IN2(n9963), .QN(n12535) );
  NOR2X0 U12741 ( .IN1(n9994), .IN2(n11130), .QN(n12534) );
  NAND2X0 U12742 ( .IN1(n10192), .IN2(n8399), .QN(n11130) );
  NAND2X0 U12743 ( .IN1(n12536), .IN2(n12537), .QN(WX8426) );
  NOR2X0 U12744 ( .IN1(n12538), .IN2(n12539), .QN(n12537) );
  NOR2X0 U12745 ( .IN1(n12540), .IN2(n9930), .QN(n12539) );
  NOR2X0 U12746 ( .IN1(n11706), .IN2(n9910), .QN(n12538) );
  NOR2X0 U12747 ( .IN1(n12541), .IN2(n12542), .QN(n11706) );
  INVX0 U12748 ( .INP(n12543), .ZN(n12542) );
  NAND2X0 U12749 ( .IN1(n12544), .IN2(n12545), .QN(n12543) );
  NOR2X0 U12750 ( .IN1(n12545), .IN2(n12544), .QN(n12541) );
  NAND2X0 U12751 ( .IN1(n12546), .IN2(n12547), .QN(n12544) );
  NAND2X0 U12752 ( .IN1(n9052), .IN2(n12548), .QN(n12547) );
  INVX0 U12753 ( .INP(n12549), .ZN(n12546) );
  NOR2X0 U12754 ( .IN1(n12548), .IN2(n9052), .QN(n12549) );
  NOR2X0 U12755 ( .IN1(n12550), .IN2(n12551), .QN(n12548) );
  INVX0 U12756 ( .INP(n12552), .ZN(n12551) );
  NAND2X0 U12757 ( .IN1(n18454), .IN2(WX9912), .QN(n12552) );
  NOR2X0 U12758 ( .IN1(WX9912), .IN2(n18454), .QN(n12550) );
  NOR2X0 U12759 ( .IN1(n12553), .IN2(n12554), .QN(n12545) );
  INVX0 U12760 ( .INP(n12555), .ZN(n12554) );
  NAND2X0 U12761 ( .IN1(n9051), .IN2(n10015), .QN(n12555) );
  NOR2X0 U12762 ( .IN1(n10004), .IN2(n9051), .QN(n12553) );
  NOR2X0 U12763 ( .IN1(n12556), .IN2(n12557), .QN(n12536) );
  NOR2X0 U12764 ( .IN1(DFF_1331_n1), .IN2(n9963), .QN(n12557) );
  NOR2X0 U12765 ( .IN1(n9994), .IN2(n11131), .QN(n12556) );
  NAND2X0 U12766 ( .IN1(n10192), .IN2(n8400), .QN(n11131) );
  NAND2X0 U12767 ( .IN1(n12558), .IN2(n12559), .QN(WX8424) );
  NOR2X0 U12768 ( .IN1(n12560), .IN2(n12561), .QN(n12559) );
  NOR2X0 U12769 ( .IN1(n12562), .IN2(n9931), .QN(n12561) );
  NOR2X0 U12770 ( .IN1(n9922), .IN2(n11730), .QN(n12560) );
  NAND2X0 U12771 ( .IN1(n12563), .IN2(n12564), .QN(n11730) );
  INVX0 U12772 ( .INP(n12565), .ZN(n12564) );
  NOR2X0 U12773 ( .IN1(n12566), .IN2(n12567), .QN(n12565) );
  NAND2X0 U12774 ( .IN1(n12567), .IN2(n12566), .QN(n12563) );
  INVX0 U12775 ( .INP(n12568), .ZN(n12566) );
  NAND2X0 U12776 ( .IN1(n12569), .IN2(n12570), .QN(n12568) );
  NAND2X0 U12777 ( .IN1(n12571), .IN2(WX9846), .QN(n12570) );
  NAND2X0 U12778 ( .IN1(n12572), .IN2(n12573), .QN(n12571) );
  NAND2X0 U12779 ( .IN1(test_so80), .IN2(WX9782), .QN(n12573) );
  NAND2X0 U12780 ( .IN1(n9053), .IN2(n9840), .QN(n12572) );
  NAND2X0 U12781 ( .IN1(n9054), .IN2(n12574), .QN(n12569) );
  NOR2X0 U12782 ( .IN1(n12575), .IN2(n12576), .QN(n12574) );
  NOR2X0 U12783 ( .IN1(test_so80), .IN2(WX9782), .QN(n12576) );
  NOR2X0 U12784 ( .IN1(n9053), .IN2(n9840), .QN(n12575) );
  NAND2X0 U12785 ( .IN1(n12577), .IN2(n12578), .QN(n12567) );
  NAND2X0 U12786 ( .IN1(n9561), .IN2(n10015), .QN(n12578) );
  NAND2X0 U12787 ( .IN1(TM1), .IN2(WX9910), .QN(n12577) );
  NOR2X0 U12788 ( .IN1(n12579), .IN2(n12580), .QN(n12558) );
  NOR2X0 U12789 ( .IN1(DFF_1332_n1), .IN2(n9962), .QN(n12580) );
  NOR2X0 U12790 ( .IN1(n9994), .IN2(n11132), .QN(n12579) );
  NAND2X0 U12791 ( .IN1(n10192), .IN2(n8401), .QN(n11132) );
  NAND2X0 U12792 ( .IN1(n12581), .IN2(n12582), .QN(WX8422) );
  NOR2X0 U12793 ( .IN1(n12583), .IN2(n12584), .QN(n12582) );
  NOR2X0 U12794 ( .IN1(n12585), .IN2(n9931), .QN(n12584) );
  NOR2X0 U12795 ( .IN1(n11752), .IN2(n9910), .QN(n12583) );
  NOR2X0 U12796 ( .IN1(n12586), .IN2(n12587), .QN(n11752) );
  INVX0 U12797 ( .INP(n12588), .ZN(n12587) );
  NAND2X0 U12798 ( .IN1(n12589), .IN2(n12590), .QN(n12588) );
  NOR2X0 U12799 ( .IN1(n12590), .IN2(n12589), .QN(n12586) );
  NAND2X0 U12800 ( .IN1(n12591), .IN2(n12592), .QN(n12589) );
  NAND2X0 U12801 ( .IN1(n9056), .IN2(n12593), .QN(n12592) );
  INVX0 U12802 ( .INP(n12594), .ZN(n12591) );
  NOR2X0 U12803 ( .IN1(n12593), .IN2(n9056), .QN(n12594) );
  NOR2X0 U12804 ( .IN1(n12595), .IN2(n12596), .QN(n12593) );
  INVX0 U12805 ( .INP(n12597), .ZN(n12596) );
  NAND2X0 U12806 ( .IN1(n18453), .IN2(WX9908), .QN(n12597) );
  NOR2X0 U12807 ( .IN1(WX9908), .IN2(n18453), .QN(n12595) );
  NOR2X0 U12808 ( .IN1(n12598), .IN2(n12599), .QN(n12590) );
  INVX0 U12809 ( .INP(n12600), .ZN(n12599) );
  NAND2X0 U12810 ( .IN1(n9055), .IN2(n10015), .QN(n12600) );
  NOR2X0 U12811 ( .IN1(n10005), .IN2(n9055), .QN(n12598) );
  NOR2X0 U12812 ( .IN1(n12601), .IN2(n12602), .QN(n12581) );
  NOR2X0 U12813 ( .IN1(DFF_1333_n1), .IN2(n9962), .QN(n12602) );
  NOR2X0 U12814 ( .IN1(n9994), .IN2(n11133), .QN(n12601) );
  NAND2X0 U12815 ( .IN1(n10191), .IN2(n8402), .QN(n11133) );
  NAND2X0 U12816 ( .IN1(n12603), .IN2(n12604), .QN(WX8420) );
  NOR2X0 U12817 ( .IN1(n12605), .IN2(n12606), .QN(n12604) );
  NOR2X0 U12818 ( .IN1(n12607), .IN2(n9931), .QN(n12606) );
  NOR2X0 U12819 ( .IN1(n11775), .IN2(n9910), .QN(n12605) );
  NOR2X0 U12820 ( .IN1(n12608), .IN2(n12609), .QN(n11775) );
  INVX0 U12821 ( .INP(n12610), .ZN(n12609) );
  NAND2X0 U12822 ( .IN1(n12611), .IN2(n12612), .QN(n12610) );
  NOR2X0 U12823 ( .IN1(n12612), .IN2(n12611), .QN(n12608) );
  NAND2X0 U12824 ( .IN1(n12613), .IN2(n12614), .QN(n12611) );
  NAND2X0 U12825 ( .IN1(n9058), .IN2(n12615), .QN(n12614) );
  INVX0 U12826 ( .INP(n12616), .ZN(n12613) );
  NOR2X0 U12827 ( .IN1(n12615), .IN2(n9058), .QN(n12616) );
  NOR2X0 U12828 ( .IN1(n12617), .IN2(n12618), .QN(n12615) );
  INVX0 U12829 ( .INP(n12619), .ZN(n12618) );
  NAND2X0 U12830 ( .IN1(n18452), .IN2(WX9906), .QN(n12619) );
  NOR2X0 U12831 ( .IN1(WX9906), .IN2(n18452), .QN(n12617) );
  NOR2X0 U12832 ( .IN1(n12620), .IN2(n12621), .QN(n12612) );
  INVX0 U12833 ( .INP(n12622), .ZN(n12621) );
  NAND2X0 U12834 ( .IN1(n9057), .IN2(n10015), .QN(n12622) );
  NOR2X0 U12835 ( .IN1(n10004), .IN2(n9057), .QN(n12620) );
  NOR2X0 U12836 ( .IN1(n12623), .IN2(n12624), .QN(n12603) );
  NOR2X0 U12837 ( .IN1(DFF_1334_n1), .IN2(n9962), .QN(n12624) );
  NOR2X0 U12838 ( .IN1(n9994), .IN2(n11134), .QN(n12623) );
  NAND2X0 U12839 ( .IN1(n10191), .IN2(n8403), .QN(n11134) );
  NAND2X0 U12840 ( .IN1(n12625), .IN2(n12626), .QN(WX8418) );
  NOR2X0 U12841 ( .IN1(n12627), .IN2(n12628), .QN(n12626) );
  NOR2X0 U12842 ( .IN1(n12629), .IN2(n9931), .QN(n12628) );
  NOR2X0 U12843 ( .IN1(n11797), .IN2(n9910), .QN(n12627) );
  NOR2X0 U12844 ( .IN1(n12630), .IN2(n12631), .QN(n11797) );
  INVX0 U12845 ( .INP(n12632), .ZN(n12631) );
  NAND2X0 U12846 ( .IN1(n12633), .IN2(n12634), .QN(n12632) );
  NOR2X0 U12847 ( .IN1(n12634), .IN2(n12633), .QN(n12630) );
  NAND2X0 U12848 ( .IN1(n12635), .IN2(n12636), .QN(n12633) );
  NAND2X0 U12849 ( .IN1(n9060), .IN2(n12637), .QN(n12636) );
  INVX0 U12850 ( .INP(n12638), .ZN(n12635) );
  NOR2X0 U12851 ( .IN1(n12637), .IN2(n9060), .QN(n12638) );
  NOR2X0 U12852 ( .IN1(n12639), .IN2(n12640), .QN(n12637) );
  INVX0 U12853 ( .INP(n12641), .ZN(n12640) );
  NAND2X0 U12854 ( .IN1(n18451), .IN2(WX9904), .QN(n12641) );
  NOR2X0 U12855 ( .IN1(WX9904), .IN2(n18451), .QN(n12639) );
  NOR2X0 U12856 ( .IN1(n12642), .IN2(n12643), .QN(n12634) );
  INVX0 U12857 ( .INP(n12644), .ZN(n12643) );
  NAND2X0 U12858 ( .IN1(n9059), .IN2(n10015), .QN(n12644) );
  NOR2X0 U12859 ( .IN1(n10004), .IN2(n9059), .QN(n12642) );
  NOR2X0 U12860 ( .IN1(n12645), .IN2(n12646), .QN(n12625) );
  NOR2X0 U12861 ( .IN1(DFF_1335_n1), .IN2(n9962), .QN(n12646) );
  NOR2X0 U12862 ( .IN1(n9994), .IN2(n11135), .QN(n12645) );
  NAND2X0 U12863 ( .IN1(n10191), .IN2(n8404), .QN(n11135) );
  NAND2X0 U12864 ( .IN1(n12647), .IN2(n12648), .QN(WX8416) );
  NOR2X0 U12865 ( .IN1(n12649), .IN2(n12650), .QN(n12648) );
  NOR2X0 U12866 ( .IN1(n12651), .IN2(n9931), .QN(n12650) );
  NOR2X0 U12867 ( .IN1(n11820), .IN2(n9910), .QN(n12649) );
  NOR2X0 U12868 ( .IN1(n12652), .IN2(n12653), .QN(n11820) );
  INVX0 U12869 ( .INP(n12654), .ZN(n12653) );
  NAND2X0 U12870 ( .IN1(n12655), .IN2(n12656), .QN(n12654) );
  NOR2X0 U12871 ( .IN1(n12656), .IN2(n12655), .QN(n12652) );
  NAND2X0 U12872 ( .IN1(n12657), .IN2(n12658), .QN(n12655) );
  NAND2X0 U12873 ( .IN1(n9062), .IN2(n12659), .QN(n12658) );
  INVX0 U12874 ( .INP(n12660), .ZN(n12657) );
  NOR2X0 U12875 ( .IN1(n12659), .IN2(n9062), .QN(n12660) );
  NOR2X0 U12876 ( .IN1(n12661), .IN2(n12662), .QN(n12659) );
  INVX0 U12877 ( .INP(n12663), .ZN(n12662) );
  NAND2X0 U12878 ( .IN1(n18450), .IN2(WX9902), .QN(n12663) );
  NOR2X0 U12879 ( .IN1(WX9902), .IN2(n18450), .QN(n12661) );
  NOR2X0 U12880 ( .IN1(n12664), .IN2(n12665), .QN(n12656) );
  INVX0 U12881 ( .INP(n12666), .ZN(n12665) );
  NAND2X0 U12882 ( .IN1(n9061), .IN2(n10015), .QN(n12666) );
  NOR2X0 U12883 ( .IN1(n10005), .IN2(n9061), .QN(n12664) );
  NOR2X0 U12884 ( .IN1(n12667), .IN2(n12668), .QN(n12647) );
  NOR2X0 U12885 ( .IN1(n9976), .IN2(n9853), .QN(n12668) );
  NOR2X0 U12886 ( .IN1(n9994), .IN2(n11136), .QN(n12667) );
  NAND2X0 U12887 ( .IN1(n10191), .IN2(n8405), .QN(n11136) );
  NAND2X0 U12888 ( .IN1(n12669), .IN2(n12670), .QN(WX8414) );
  NOR2X0 U12889 ( .IN1(n12671), .IN2(n12672), .QN(n12670) );
  NOR2X0 U12890 ( .IN1(n12673), .IN2(n9931), .QN(n12672) );
  NOR2X0 U12891 ( .IN1(n11842), .IN2(n9910), .QN(n12671) );
  NOR2X0 U12892 ( .IN1(n12674), .IN2(n12675), .QN(n11842) );
  INVX0 U12893 ( .INP(n12676), .ZN(n12675) );
  NAND2X0 U12894 ( .IN1(n12677), .IN2(n12678), .QN(n12676) );
  NOR2X0 U12895 ( .IN1(n12678), .IN2(n12677), .QN(n12674) );
  NAND2X0 U12896 ( .IN1(n12679), .IN2(n12680), .QN(n12677) );
  NAND2X0 U12897 ( .IN1(n9064), .IN2(n12681), .QN(n12680) );
  INVX0 U12898 ( .INP(n12682), .ZN(n12679) );
  NOR2X0 U12899 ( .IN1(n12681), .IN2(n9064), .QN(n12682) );
  NOR2X0 U12900 ( .IN1(n12683), .IN2(n12684), .QN(n12681) );
  INVX0 U12901 ( .INP(n12685), .ZN(n12684) );
  NAND2X0 U12902 ( .IN1(n18449), .IN2(WX9900), .QN(n12685) );
  NOR2X0 U12903 ( .IN1(WX9900), .IN2(n18449), .QN(n12683) );
  NOR2X0 U12904 ( .IN1(n12686), .IN2(n12687), .QN(n12678) );
  INVX0 U12905 ( .INP(n12688), .ZN(n12687) );
  NAND2X0 U12906 ( .IN1(n9063), .IN2(n10014), .QN(n12688) );
  NOR2X0 U12907 ( .IN1(n10005), .IN2(n9063), .QN(n12686) );
  NOR2X0 U12908 ( .IN1(n12689), .IN2(n12690), .QN(n12669) );
  NOR2X0 U12909 ( .IN1(DFF_1337_n1), .IN2(n9962), .QN(n12690) );
  NOR2X0 U12910 ( .IN1(n9994), .IN2(n11137), .QN(n12689) );
  NAND2X0 U12911 ( .IN1(n10191), .IN2(n8406), .QN(n11137) );
  NAND2X0 U12912 ( .IN1(n12691), .IN2(n12692), .QN(WX8412) );
  NOR2X0 U12913 ( .IN1(n12693), .IN2(n12694), .QN(n12692) );
  NOR2X0 U12914 ( .IN1(n9941), .IN2(n12695), .QN(n12694) );
  NOR2X0 U12915 ( .IN1(n11866), .IN2(n9910), .QN(n12693) );
  NOR2X0 U12916 ( .IN1(n12696), .IN2(n12697), .QN(n11866) );
  INVX0 U12917 ( .INP(n12698), .ZN(n12697) );
  NAND2X0 U12918 ( .IN1(n12699), .IN2(n12700), .QN(n12698) );
  NOR2X0 U12919 ( .IN1(n12700), .IN2(n12699), .QN(n12696) );
  NAND2X0 U12920 ( .IN1(n12701), .IN2(n12702), .QN(n12699) );
  NAND2X0 U12921 ( .IN1(n9066), .IN2(n12703), .QN(n12702) );
  INVX0 U12922 ( .INP(n12704), .ZN(n12701) );
  NOR2X0 U12923 ( .IN1(n12703), .IN2(n9066), .QN(n12704) );
  NOR2X0 U12924 ( .IN1(n12705), .IN2(n12706), .QN(n12703) );
  INVX0 U12925 ( .INP(n12707), .ZN(n12706) );
  NAND2X0 U12926 ( .IN1(n18448), .IN2(WX9898), .QN(n12707) );
  NOR2X0 U12927 ( .IN1(WX9898), .IN2(n18448), .QN(n12705) );
  NOR2X0 U12928 ( .IN1(n12708), .IN2(n12709), .QN(n12700) );
  INVX0 U12929 ( .INP(n12710), .ZN(n12709) );
  NAND2X0 U12930 ( .IN1(n9065), .IN2(n10014), .QN(n12710) );
  NOR2X0 U12931 ( .IN1(n10005), .IN2(n9065), .QN(n12708) );
  NOR2X0 U12932 ( .IN1(n12711), .IN2(n12712), .QN(n12691) );
  NOR2X0 U12933 ( .IN1(DFF_1338_n1), .IN2(n9962), .QN(n12712) );
  NOR2X0 U12934 ( .IN1(n9994), .IN2(n11138), .QN(n12711) );
  NAND2X0 U12935 ( .IN1(n10191), .IN2(n8407), .QN(n11138) );
  NAND2X0 U12936 ( .IN1(n12713), .IN2(n12714), .QN(WX8410) );
  NOR2X0 U12937 ( .IN1(n12715), .IN2(n12716), .QN(n12714) );
  NOR2X0 U12938 ( .IN1(n12717), .IN2(n9931), .QN(n12716) );
  NOR2X0 U12939 ( .IN1(n11888), .IN2(n9910), .QN(n12715) );
  NOR2X0 U12940 ( .IN1(n12718), .IN2(n12719), .QN(n11888) );
  INVX0 U12941 ( .INP(n12720), .ZN(n12719) );
  NAND2X0 U12942 ( .IN1(n12721), .IN2(n12722), .QN(n12720) );
  NOR2X0 U12943 ( .IN1(n12722), .IN2(n12721), .QN(n12718) );
  NAND2X0 U12944 ( .IN1(n12723), .IN2(n12724), .QN(n12721) );
  NAND2X0 U12945 ( .IN1(n9068), .IN2(n12725), .QN(n12724) );
  INVX0 U12946 ( .INP(n12726), .ZN(n12723) );
  NOR2X0 U12947 ( .IN1(n12725), .IN2(n9068), .QN(n12726) );
  NOR2X0 U12948 ( .IN1(n12727), .IN2(n12728), .QN(n12725) );
  INVX0 U12949 ( .INP(n12729), .ZN(n12728) );
  NAND2X0 U12950 ( .IN1(n18447), .IN2(WX9896), .QN(n12729) );
  NOR2X0 U12951 ( .IN1(WX9896), .IN2(n18447), .QN(n12727) );
  NOR2X0 U12952 ( .IN1(n12730), .IN2(n12731), .QN(n12722) );
  INVX0 U12953 ( .INP(n12732), .ZN(n12731) );
  NAND2X0 U12954 ( .IN1(n9067), .IN2(n10014), .QN(n12732) );
  NOR2X0 U12955 ( .IN1(n10005), .IN2(n9067), .QN(n12730) );
  NOR2X0 U12956 ( .IN1(n12733), .IN2(n12734), .QN(n12713) );
  NOR2X0 U12957 ( .IN1(DFF_1339_n1), .IN2(n9962), .QN(n12734) );
  NOR2X0 U12958 ( .IN1(n9994), .IN2(n11139), .QN(n12733) );
  NAND2X0 U12959 ( .IN1(n10194), .IN2(n8408), .QN(n11139) );
  NAND2X0 U12960 ( .IN1(n12735), .IN2(n12736), .QN(WX8408) );
  NOR2X0 U12961 ( .IN1(n12737), .IN2(n12738), .QN(n12736) );
  NOR2X0 U12962 ( .IN1(n9941), .IN2(n12739), .QN(n12738) );
  NOR2X0 U12963 ( .IN1(n11910), .IN2(n9910), .QN(n12737) );
  NOR2X0 U12964 ( .IN1(n12740), .IN2(n12741), .QN(n11910) );
  INVX0 U12965 ( .INP(n12742), .ZN(n12741) );
  NAND2X0 U12966 ( .IN1(n12743), .IN2(n12744), .QN(n12742) );
  NOR2X0 U12967 ( .IN1(n12744), .IN2(n12743), .QN(n12740) );
  NAND2X0 U12968 ( .IN1(n12745), .IN2(n12746), .QN(n12743) );
  NAND2X0 U12969 ( .IN1(n9070), .IN2(n12747), .QN(n12746) );
  INVX0 U12970 ( .INP(n12748), .ZN(n12745) );
  NOR2X0 U12971 ( .IN1(n12747), .IN2(n9070), .QN(n12748) );
  NOR2X0 U12972 ( .IN1(n12749), .IN2(n12750), .QN(n12747) );
  INVX0 U12973 ( .INP(n12751), .ZN(n12750) );
  NAND2X0 U12974 ( .IN1(n18446), .IN2(WX9894), .QN(n12751) );
  NOR2X0 U12975 ( .IN1(WX9894), .IN2(n18446), .QN(n12749) );
  NOR2X0 U12976 ( .IN1(n12752), .IN2(n12753), .QN(n12744) );
  INVX0 U12977 ( .INP(n12754), .ZN(n12753) );
  NAND2X0 U12978 ( .IN1(n9069), .IN2(n10014), .QN(n12754) );
  NOR2X0 U12979 ( .IN1(n10005), .IN2(n9069), .QN(n12752) );
  NOR2X0 U12980 ( .IN1(n12755), .IN2(n12756), .QN(n12735) );
  NOR2X0 U12981 ( .IN1(DFF_1340_n1), .IN2(n9962), .QN(n12756) );
  NOR2X0 U12982 ( .IN1(n9994), .IN2(n11140), .QN(n12755) );
  NAND2X0 U12983 ( .IN1(n10213), .IN2(n8409), .QN(n11140) );
  NAND2X0 U12984 ( .IN1(n12757), .IN2(n12758), .QN(WX8406) );
  NOR2X0 U12985 ( .IN1(n12759), .IN2(n12760), .QN(n12758) );
  NOR2X0 U12986 ( .IN1(n12761), .IN2(n9931), .QN(n12760) );
  NOR2X0 U12987 ( .IN1(n11932), .IN2(n9910), .QN(n12759) );
  NOR2X0 U12988 ( .IN1(n12762), .IN2(n12763), .QN(n11932) );
  INVX0 U12989 ( .INP(n12764), .ZN(n12763) );
  NAND2X0 U12990 ( .IN1(n12765), .IN2(n12766), .QN(n12764) );
  NOR2X0 U12991 ( .IN1(n12766), .IN2(n12765), .QN(n12762) );
  NAND2X0 U12992 ( .IN1(n12767), .IN2(n12768), .QN(n12765) );
  NAND2X0 U12993 ( .IN1(n9072), .IN2(n12769), .QN(n12768) );
  INVX0 U12994 ( .INP(n12770), .ZN(n12767) );
  NOR2X0 U12995 ( .IN1(n12769), .IN2(n9072), .QN(n12770) );
  NOR2X0 U12996 ( .IN1(n12771), .IN2(n12772), .QN(n12769) );
  INVX0 U12997 ( .INP(n12773), .ZN(n12772) );
  NAND2X0 U12998 ( .IN1(n18445), .IN2(WX9892), .QN(n12773) );
  NOR2X0 U12999 ( .IN1(WX9892), .IN2(n18445), .QN(n12771) );
  NOR2X0 U13000 ( .IN1(n12774), .IN2(n12775), .QN(n12766) );
  INVX0 U13001 ( .INP(n12776), .ZN(n12775) );
  NAND2X0 U13002 ( .IN1(n9071), .IN2(n10014), .QN(n12776) );
  NOR2X0 U13003 ( .IN1(n10005), .IN2(n9071), .QN(n12774) );
  NOR2X0 U13004 ( .IN1(n12777), .IN2(n12778), .QN(n12757) );
  NOR2X0 U13005 ( .IN1(DFF_1341_n1), .IN2(n9962), .QN(n12778) );
  NOR2X0 U13006 ( .IN1(n9994), .IN2(n11141), .QN(n12777) );
  NAND2X0 U13007 ( .IN1(n10214), .IN2(n8410), .QN(n11141) );
  NAND2X0 U13008 ( .IN1(n12779), .IN2(n12780), .QN(WX8404) );
  NOR2X0 U13009 ( .IN1(n12781), .IN2(n12782), .QN(n12780) );
  NOR2X0 U13010 ( .IN1(n9941), .IN2(n12783), .QN(n12782) );
  NOR2X0 U13011 ( .IN1(n11954), .IN2(n9911), .QN(n12781) );
  NOR2X0 U13012 ( .IN1(n12784), .IN2(n12785), .QN(n11954) );
  INVX0 U13013 ( .INP(n12786), .ZN(n12785) );
  NAND2X0 U13014 ( .IN1(n12787), .IN2(n12788), .QN(n12786) );
  NOR2X0 U13015 ( .IN1(n12788), .IN2(n12787), .QN(n12784) );
  NAND2X0 U13016 ( .IN1(n12789), .IN2(n12790), .QN(n12787) );
  NAND2X0 U13017 ( .IN1(n9074), .IN2(n12791), .QN(n12790) );
  INVX0 U13018 ( .INP(n12792), .ZN(n12789) );
  NOR2X0 U13019 ( .IN1(n12791), .IN2(n9074), .QN(n12792) );
  NOR2X0 U13020 ( .IN1(n12793), .IN2(n12794), .QN(n12791) );
  INVX0 U13021 ( .INP(n12795), .ZN(n12794) );
  NAND2X0 U13022 ( .IN1(n18444), .IN2(WX9890), .QN(n12795) );
  NOR2X0 U13023 ( .IN1(WX9890), .IN2(n18444), .QN(n12793) );
  NOR2X0 U13024 ( .IN1(n12796), .IN2(n12797), .QN(n12788) );
  INVX0 U13025 ( .INP(n12798), .ZN(n12797) );
  NAND2X0 U13026 ( .IN1(n9073), .IN2(n10014), .QN(n12798) );
  NOR2X0 U13027 ( .IN1(n10005), .IN2(n9073), .QN(n12796) );
  NOR2X0 U13028 ( .IN1(n12799), .IN2(n12800), .QN(n12779) );
  NOR2X0 U13029 ( .IN1(DFF_1342_n1), .IN2(n9962), .QN(n12800) );
  NOR2X0 U13030 ( .IN1(n9993), .IN2(n11142), .QN(n12799) );
  NAND2X0 U13031 ( .IN1(n10214), .IN2(n8411), .QN(n11142) );
  NAND2X0 U13032 ( .IN1(n12801), .IN2(n12802), .QN(WX8402) );
  NOR2X0 U13033 ( .IN1(n12803), .IN2(n12804), .QN(n12802) );
  NOR2X0 U13034 ( .IN1(n12805), .IN2(n9931), .QN(n12804) );
  NOR2X0 U13035 ( .IN1(n9921), .IN2(n11976), .QN(n12803) );
  NAND2X0 U13036 ( .IN1(n12806), .IN2(n12807), .QN(n11976) );
  NAND2X0 U13037 ( .IN1(n12808), .IN2(n12809), .QN(n12807) );
  INVX0 U13038 ( .INP(n12810), .ZN(n12806) );
  NOR2X0 U13039 ( .IN1(n12809), .IN2(n12808), .QN(n12810) );
  NAND2X0 U13040 ( .IN1(n12811), .IN2(n12812), .QN(n12808) );
  NAND2X0 U13041 ( .IN1(n12813), .IN2(WX9824), .QN(n12812) );
  NAND2X0 U13042 ( .IN1(n12814), .IN2(n12815), .QN(n12813) );
  NAND2X0 U13043 ( .IN1(test_so85), .IN2(WX9760), .QN(n12815) );
  NAND2X0 U13044 ( .IN1(n9005), .IN2(n9833), .QN(n12814) );
  NAND2X0 U13045 ( .IN1(n9006), .IN2(n12816), .QN(n12811) );
  NOR2X0 U13046 ( .IN1(n12817), .IN2(n12818), .QN(n12816) );
  NOR2X0 U13047 ( .IN1(test_so85), .IN2(WX9760), .QN(n12818) );
  NOR2X0 U13048 ( .IN1(n9005), .IN2(n9833), .QN(n12817) );
  NOR2X0 U13049 ( .IN1(n12819), .IN2(n12820), .QN(n12809) );
  INVX0 U13050 ( .INP(n12821), .ZN(n12820) );
  NAND2X0 U13051 ( .IN1(n18443), .IN2(n10014), .QN(n12821) );
  NOR2X0 U13052 ( .IN1(n10005), .IN2(n18443), .QN(n12819) );
  NOR2X0 U13053 ( .IN1(n12822), .IN2(n12823), .QN(n12801) );
  NOR2X0 U13054 ( .IN1(n9490), .IN2(n11994), .QN(n12823) );
  NOR2X0 U13055 ( .IN1(DFF_1343_n1), .IN2(n9962), .QN(n12822) );
  INVX0 U13056 ( .INP(n12824), .ZN(WX8304) );
  NAND2X0 U13057 ( .IN1(n10214), .IN2(n9490), .QN(n12824) );
  NOR2X0 U13058 ( .IN1(n10323), .IN2(n12825), .QN(WX7791) );
  NAND2X0 U13059 ( .IN1(n12826), .IN2(n12827), .QN(n12825) );
  INVX0 U13060 ( .INP(n12828), .ZN(n12827) );
  NOR2X0 U13061 ( .IN1(WX7302), .IN2(DFF_1150_n1), .QN(n12828) );
  NAND2X0 U13062 ( .IN1(DFF_1150_n1), .IN2(WX7302), .QN(n12826) );
  NOR2X0 U13063 ( .IN1(n10323), .IN2(n12829), .QN(WX7789) );
  NOR2X0 U13064 ( .IN1(n12830), .IN2(n12831), .QN(n12829) );
  NOR2X0 U13065 ( .IN1(test_so66), .IN2(WX7304), .QN(n12831) );
  NOR2X0 U13066 ( .IN1(n9604), .IN2(n9855), .QN(n12830) );
  NOR2X0 U13067 ( .IN1(n10323), .IN2(n12832), .QN(WX7787) );
  NAND2X0 U13068 ( .IN1(n12833), .IN2(n12834), .QN(n12832) );
  INVX0 U13069 ( .INP(n12835), .ZN(n12834) );
  NOR2X0 U13070 ( .IN1(WX7306), .IN2(DFF_1148_n1), .QN(n12835) );
  NAND2X0 U13071 ( .IN1(DFF_1148_n1), .IN2(WX7306), .QN(n12833) );
  NOR2X0 U13072 ( .IN1(n10324), .IN2(n12836), .QN(WX7785) );
  NAND2X0 U13073 ( .IN1(n12837), .IN2(n12838), .QN(n12836) );
  INVX0 U13074 ( .INP(n12839), .ZN(n12838) );
  NOR2X0 U13075 ( .IN1(WX7308), .IN2(DFF_1147_n1), .QN(n12839) );
  NAND2X0 U13076 ( .IN1(DFF_1147_n1), .IN2(WX7308), .QN(n12837) );
  NOR2X0 U13077 ( .IN1(n10324), .IN2(n12840), .QN(WX7783) );
  NAND2X0 U13078 ( .IN1(n12841), .IN2(n12842), .QN(n12840) );
  INVX0 U13079 ( .INP(n12843), .ZN(n12842) );
  NOR2X0 U13080 ( .IN1(WX7310), .IN2(DFF_1146_n1), .QN(n12843) );
  NAND2X0 U13081 ( .IN1(DFF_1146_n1), .IN2(WX7310), .QN(n12841) );
  NOR2X0 U13082 ( .IN1(n10324), .IN2(n12844), .QN(WX7781) );
  NAND2X0 U13083 ( .IN1(n12845), .IN2(n12846), .QN(n12844) );
  INVX0 U13084 ( .INP(n12847), .ZN(n12846) );
  NOR2X0 U13085 ( .IN1(WX7312), .IN2(DFF_1145_n1), .QN(n12847) );
  NAND2X0 U13086 ( .IN1(DFF_1145_n1), .IN2(WX7312), .QN(n12845) );
  NOR2X0 U13087 ( .IN1(n10324), .IN2(n12848), .QN(WX7779) );
  NAND2X0 U13088 ( .IN1(n12849), .IN2(n12850), .QN(n12848) );
  INVX0 U13089 ( .INP(n12851), .ZN(n12850) );
  NOR2X0 U13090 ( .IN1(WX7314), .IN2(DFF_1144_n1), .QN(n12851) );
  NAND2X0 U13091 ( .IN1(DFF_1144_n1), .IN2(WX7314), .QN(n12849) );
  NOR2X0 U13092 ( .IN1(n10324), .IN2(n12852), .QN(WX7777) );
  NAND2X0 U13093 ( .IN1(n12853), .IN2(n12854), .QN(n12852) );
  INVX0 U13094 ( .INP(n12855), .ZN(n12854) );
  NOR2X0 U13095 ( .IN1(WX7316), .IN2(DFF_1143_n1), .QN(n12855) );
  NAND2X0 U13096 ( .IN1(DFF_1143_n1), .IN2(WX7316), .QN(n12853) );
  NOR2X0 U13097 ( .IN1(n10324), .IN2(n12856), .QN(WX7775) );
  NAND2X0 U13098 ( .IN1(n12857), .IN2(n12858), .QN(n12856) );
  INVX0 U13099 ( .INP(n12859), .ZN(n12858) );
  NOR2X0 U13100 ( .IN1(WX7318), .IN2(DFF_1142_n1), .QN(n12859) );
  NAND2X0 U13101 ( .IN1(DFF_1142_n1), .IN2(WX7318), .QN(n12857) );
  NOR2X0 U13102 ( .IN1(n10324), .IN2(n12860), .QN(WX7773) );
  NAND2X0 U13103 ( .IN1(n12861), .IN2(n12862), .QN(n12860) );
  INVX0 U13104 ( .INP(n12863), .ZN(n12862) );
  NOR2X0 U13105 ( .IN1(WX7320), .IN2(DFF_1141_n1), .QN(n12863) );
  NAND2X0 U13106 ( .IN1(DFF_1141_n1), .IN2(WX7320), .QN(n12861) );
  NOR2X0 U13107 ( .IN1(n10324), .IN2(n12864), .QN(WX7771) );
  NOR2X0 U13108 ( .IN1(n12865), .IN2(n12866), .QN(n12864) );
  INVX0 U13109 ( .INP(n12867), .ZN(n12866) );
  NAND2X0 U13110 ( .IN1(n9829), .IN2(DFF_1140_n1), .QN(n12867) );
  NOR2X0 U13111 ( .IN1(DFF_1140_n1), .IN2(n9829), .QN(n12865) );
  NOR2X0 U13112 ( .IN1(n10324), .IN2(n12868), .QN(WX7769) );
  NAND2X0 U13113 ( .IN1(n12869), .IN2(n12870), .QN(n12868) );
  INVX0 U13114 ( .INP(n12871), .ZN(n12870) );
  NOR2X0 U13115 ( .IN1(WX7324), .IN2(DFF_1139_n1), .QN(n12871) );
  NAND2X0 U13116 ( .IN1(DFF_1139_n1), .IN2(WX7324), .QN(n12869) );
  NOR2X0 U13117 ( .IN1(n10324), .IN2(n12872), .QN(WX7767) );
  NAND2X0 U13118 ( .IN1(n12873), .IN2(n12874), .QN(n12872) );
  INVX0 U13119 ( .INP(n12875), .ZN(n12874) );
  NOR2X0 U13120 ( .IN1(WX7326), .IN2(DFF_1138_n1), .QN(n12875) );
  NAND2X0 U13121 ( .IN1(DFF_1138_n1), .IN2(WX7326), .QN(n12873) );
  NOR2X0 U13122 ( .IN1(n10324), .IN2(n12876), .QN(WX7765) );
  NAND2X0 U13123 ( .IN1(n12877), .IN2(n12878), .QN(n12876) );
  INVX0 U13124 ( .INP(n12879), .ZN(n12878) );
  NOR2X0 U13125 ( .IN1(WX7328), .IN2(DFF_1137_n1), .QN(n12879) );
  NAND2X0 U13126 ( .IN1(DFF_1137_n1), .IN2(WX7328), .QN(n12877) );
  NOR2X0 U13127 ( .IN1(n10324), .IN2(n12880), .QN(WX7763) );
  NAND2X0 U13128 ( .IN1(n12881), .IN2(n12882), .QN(n12880) );
  INVX0 U13129 ( .INP(n12883), .ZN(n12882) );
  NOR2X0 U13130 ( .IN1(WX7330), .IN2(DFF_1136_n1), .QN(n12883) );
  NAND2X0 U13131 ( .IN1(DFF_1136_n1), .IN2(WX7330), .QN(n12881) );
  NOR2X0 U13132 ( .IN1(n10324), .IN2(n12884), .QN(WX7761) );
  NOR2X0 U13133 ( .IN1(n12885), .IN2(n12886), .QN(n12884) );
  INVX0 U13134 ( .INP(n12887), .ZN(n12886) );
  NAND2X0 U13135 ( .IN1(CRC_OUT_4_15), .IN2(n12888), .QN(n12887) );
  NOR2X0 U13136 ( .IN1(n12888), .IN2(CRC_OUT_4_15), .QN(n12885) );
  NAND2X0 U13137 ( .IN1(n12889), .IN2(n12890), .QN(n12888) );
  NAND2X0 U13138 ( .IN1(n9505), .IN2(CRC_OUT_4_31), .QN(n12890) );
  NAND2X0 U13139 ( .IN1(DFF_1151_n1), .IN2(WX7332), .QN(n12889) );
  NOR2X0 U13140 ( .IN1(n10325), .IN2(n12891), .QN(WX7759) );
  NAND2X0 U13141 ( .IN1(n12892), .IN2(n12893), .QN(n12891) );
  INVX0 U13142 ( .INP(n12894), .ZN(n12893) );
  NOR2X0 U13143 ( .IN1(WX7334), .IN2(DFF_1134_n1), .QN(n12894) );
  NAND2X0 U13144 ( .IN1(DFF_1134_n1), .IN2(WX7334), .QN(n12892) );
  NOR2X0 U13145 ( .IN1(n10325), .IN2(n12895), .QN(WX7757) );
  NAND2X0 U13146 ( .IN1(n12896), .IN2(n12897), .QN(n12895) );
  INVX0 U13147 ( .INP(n12898), .ZN(n12897) );
  NOR2X0 U13148 ( .IN1(WX7336), .IN2(DFF_1133_n1), .QN(n12898) );
  NAND2X0 U13149 ( .IN1(DFF_1133_n1), .IN2(WX7336), .QN(n12896) );
  NOR2X0 U13150 ( .IN1(n10325), .IN2(n12899), .QN(WX7755) );
  NOR2X0 U13151 ( .IN1(n12900), .IN2(n12901), .QN(n12899) );
  NOR2X0 U13152 ( .IN1(test_so65), .IN2(WX7338), .QN(n12901) );
  NOR2X0 U13153 ( .IN1(n9619), .IN2(n9854), .QN(n12900) );
  NOR2X0 U13154 ( .IN1(n10325), .IN2(n12902), .QN(WX7753) );
  NAND2X0 U13155 ( .IN1(n12903), .IN2(n12904), .QN(n12902) );
  INVX0 U13156 ( .INP(n12905), .ZN(n12904) );
  NOR2X0 U13157 ( .IN1(WX7340), .IN2(DFF_1131_n1), .QN(n12905) );
  NAND2X0 U13158 ( .IN1(DFF_1131_n1), .IN2(WX7340), .QN(n12903) );
  NOR2X0 U13159 ( .IN1(n10325), .IN2(n12906), .QN(WX7751) );
  NOR2X0 U13160 ( .IN1(n12907), .IN2(n12908), .QN(n12906) );
  INVX0 U13161 ( .INP(n12909), .ZN(n12908) );
  NAND2X0 U13162 ( .IN1(CRC_OUT_4_10), .IN2(n12910), .QN(n12909) );
  NOR2X0 U13163 ( .IN1(n12910), .IN2(CRC_OUT_4_10), .QN(n12907) );
  NAND2X0 U13164 ( .IN1(n12911), .IN2(n12912), .QN(n12910) );
  NAND2X0 U13165 ( .IN1(n9506), .IN2(CRC_OUT_4_31), .QN(n12912) );
  NAND2X0 U13166 ( .IN1(DFF_1151_n1), .IN2(WX7342), .QN(n12911) );
  NOR2X0 U13167 ( .IN1(n10325), .IN2(n12913), .QN(WX7749) );
  NAND2X0 U13168 ( .IN1(n12914), .IN2(n12915), .QN(n12913) );
  INVX0 U13169 ( .INP(n12916), .ZN(n12915) );
  NOR2X0 U13170 ( .IN1(WX7344), .IN2(DFF_1129_n1), .QN(n12916) );
  NAND2X0 U13171 ( .IN1(DFF_1129_n1), .IN2(WX7344), .QN(n12914) );
  NOR2X0 U13172 ( .IN1(n10325), .IN2(n12917), .QN(WX7747) );
  NAND2X0 U13173 ( .IN1(n12918), .IN2(n12919), .QN(n12917) );
  INVX0 U13174 ( .INP(n12920), .ZN(n12919) );
  NOR2X0 U13175 ( .IN1(WX7346), .IN2(DFF_1128_n1), .QN(n12920) );
  NAND2X0 U13176 ( .IN1(DFF_1128_n1), .IN2(WX7346), .QN(n12918) );
  NOR2X0 U13177 ( .IN1(n10325), .IN2(n12921), .QN(WX7745) );
  NAND2X0 U13178 ( .IN1(n12922), .IN2(n12923), .QN(n12921) );
  INVX0 U13179 ( .INP(n12924), .ZN(n12923) );
  NOR2X0 U13180 ( .IN1(WX7348), .IN2(DFF_1127_n1), .QN(n12924) );
  NAND2X0 U13181 ( .IN1(DFF_1127_n1), .IN2(WX7348), .QN(n12922) );
  NOR2X0 U13182 ( .IN1(n10325), .IN2(n12925), .QN(WX7743) );
  NAND2X0 U13183 ( .IN1(n12926), .IN2(n12927), .QN(n12925) );
  INVX0 U13184 ( .INP(n12928), .ZN(n12927) );
  NOR2X0 U13185 ( .IN1(WX7350), .IN2(DFF_1126_n1), .QN(n12928) );
  NAND2X0 U13186 ( .IN1(DFF_1126_n1), .IN2(WX7350), .QN(n12926) );
  NOR2X0 U13187 ( .IN1(n10325), .IN2(n12929), .QN(WX7741) );
  NAND2X0 U13188 ( .IN1(n12930), .IN2(n12931), .QN(n12929) );
  INVX0 U13189 ( .INP(n12932), .ZN(n12931) );
  NOR2X0 U13190 ( .IN1(WX7352), .IN2(DFF_1125_n1), .QN(n12932) );
  NAND2X0 U13191 ( .IN1(DFF_1125_n1), .IN2(WX7352), .QN(n12930) );
  NOR2X0 U13192 ( .IN1(n10325), .IN2(n12933), .QN(WX7739) );
  NAND2X0 U13193 ( .IN1(n12934), .IN2(n12935), .QN(n12933) );
  INVX0 U13194 ( .INP(n12936), .ZN(n12935) );
  NOR2X0 U13195 ( .IN1(WX7354), .IN2(DFF_1124_n1), .QN(n12936) );
  NAND2X0 U13196 ( .IN1(DFF_1124_n1), .IN2(WX7354), .QN(n12934) );
  NOR2X0 U13197 ( .IN1(n10325), .IN2(n12937), .QN(WX7737) );
  NAND2X0 U13198 ( .IN1(n12938), .IN2(n12939), .QN(n12937) );
  INVX0 U13199 ( .INP(n12940), .ZN(n12939) );
  NOR2X0 U13200 ( .IN1(CRC_OUT_4_3), .IN2(n12941), .QN(n12940) );
  NAND2X0 U13201 ( .IN1(n12941), .IN2(CRC_OUT_4_3), .QN(n12938) );
  NAND2X0 U13202 ( .IN1(n12942), .IN2(n12943), .QN(n12941) );
  NAND2X0 U13203 ( .IN1(test_so64), .IN2(CRC_OUT_4_31), .QN(n12943) );
  NAND2X0 U13204 ( .IN1(DFF_1151_n1), .IN2(n9849), .QN(n12942) );
  NOR2X0 U13205 ( .IN1(n10325), .IN2(n12944), .QN(WX7735) );
  NAND2X0 U13206 ( .IN1(n12945), .IN2(n12946), .QN(n12944) );
  INVX0 U13207 ( .INP(n12947), .ZN(n12946) );
  NOR2X0 U13208 ( .IN1(WX7358), .IN2(DFF_1122_n1), .QN(n12947) );
  NAND2X0 U13209 ( .IN1(DFF_1122_n1), .IN2(WX7358), .QN(n12945) );
  NOR2X0 U13210 ( .IN1(n10326), .IN2(n12948), .QN(WX7733) );
  NAND2X0 U13211 ( .IN1(n12949), .IN2(n12950), .QN(n12948) );
  INVX0 U13212 ( .INP(n12951), .ZN(n12950) );
  NOR2X0 U13213 ( .IN1(WX7360), .IN2(DFF_1121_n1), .QN(n12951) );
  NAND2X0 U13214 ( .IN1(DFF_1121_n1), .IN2(WX7360), .QN(n12949) );
  NOR2X0 U13215 ( .IN1(n10326), .IN2(n12952), .QN(WX7731) );
  NAND2X0 U13216 ( .IN1(n12953), .IN2(n12954), .QN(n12952) );
  INVX0 U13217 ( .INP(n12955), .ZN(n12954) );
  NOR2X0 U13218 ( .IN1(WX7362), .IN2(DFF_1120_n1), .QN(n12955) );
  NAND2X0 U13219 ( .IN1(DFF_1120_n1), .IN2(WX7362), .QN(n12953) );
  NOR2X0 U13220 ( .IN1(n10326), .IN2(n12956), .QN(WX7729) );
  NAND2X0 U13221 ( .IN1(n12957), .IN2(n12958), .QN(n12956) );
  NAND2X0 U13222 ( .IN1(n9520), .IN2(CRC_OUT_4_31), .QN(n12958) );
  NAND2X0 U13223 ( .IN1(DFF_1151_n1), .IN2(WX7364), .QN(n12957) );
  NOR2X0 U13224 ( .IN1(n18426), .IN2(n10236), .QN(WX7203) );
  NOR2X0 U13225 ( .IN1(n18425), .IN2(n10236), .QN(WX7201) );
  NOR2X0 U13226 ( .IN1(n18424), .IN2(n10237), .QN(WX7199) );
  NOR2X0 U13227 ( .IN1(n18423), .IN2(n10237), .QN(WX7197) );
  NOR2X0 U13228 ( .IN1(n18422), .IN2(n10237), .QN(WX7195) );
  NOR2X0 U13229 ( .IN1(n18421), .IN2(n10237), .QN(WX7193) );
  NOR2X0 U13230 ( .IN1(n18420), .IN2(n10237), .QN(WX7191) );
  NOR2X0 U13231 ( .IN1(n18419), .IN2(n10237), .QN(WX7189) );
  NOR2X0 U13232 ( .IN1(n18418), .IN2(n10237), .QN(WX7187) );
  NOR2X0 U13233 ( .IN1(n18417), .IN2(n10237), .QN(WX7185) );
  NOR2X0 U13234 ( .IN1(n18416), .IN2(n10237), .QN(WX7183) );
  NOR2X0 U13235 ( .IN1(n10326), .IN2(n9841), .QN(WX7181) );
  NOR2X0 U13236 ( .IN1(n18415), .IN2(n10237), .QN(WX7179) );
  NOR2X0 U13237 ( .IN1(n18414), .IN2(n10237), .QN(WX7177) );
  NOR2X0 U13238 ( .IN1(n18413), .IN2(n10237), .QN(WX7175) );
  NOR2X0 U13239 ( .IN1(n18412), .IN2(n10238), .QN(WX7173) );
  NAND2X0 U13240 ( .IN1(n12959), .IN2(n12960), .QN(WX7171) );
  NOR2X0 U13241 ( .IN1(n12961), .IN2(n12962), .QN(n12960) );
  NOR2X0 U13242 ( .IN1(n12963), .IN2(n9931), .QN(n12962) );
  NOR2X0 U13243 ( .IN1(n12134), .IN2(n9911), .QN(n12961) );
  INVX0 U13244 ( .INP(n12964), .ZN(n12134) );
  NAND2X0 U13245 ( .IN1(n12965), .IN2(n12966), .QN(n12964) );
  NAND2X0 U13246 ( .IN1(n12967), .IN2(n12968), .QN(n12966) );
  NAND2X0 U13247 ( .IN1(n12969), .IN2(n12970), .QN(n12968) );
  NAND2X0 U13248 ( .IN1(n9307), .IN2(WX8465), .QN(n12970) );
  NAND2X0 U13249 ( .IN1(n9306), .IN2(WX8593), .QN(n12969) );
  NOR2X0 U13250 ( .IN1(n12971), .IN2(n12972), .QN(n12967) );
  NOR2X0 U13251 ( .IN1(n9519), .IN2(WX8529), .QN(n12972) );
  NOR2X0 U13252 ( .IN1(n3595), .IN2(WX8657), .QN(n12971) );
  NAND2X0 U13253 ( .IN1(n12973), .IN2(n12974), .QN(n12965) );
  NAND2X0 U13254 ( .IN1(n12975), .IN2(n12976), .QN(n12974) );
  NAND2X0 U13255 ( .IN1(n9519), .IN2(WX8529), .QN(n12976) );
  NAND2X0 U13256 ( .IN1(n3595), .IN2(WX8657), .QN(n12975) );
  NOR2X0 U13257 ( .IN1(n12977), .IN2(n12978), .QN(n12973) );
  NOR2X0 U13258 ( .IN1(n9307), .IN2(WX8465), .QN(n12978) );
  NOR2X0 U13259 ( .IN1(n9306), .IN2(WX8593), .QN(n12977) );
  NOR2X0 U13260 ( .IN1(n12979), .IN2(n12980), .QN(n12959) );
  NOR2X0 U13261 ( .IN1(DFF_1120_n1), .IN2(n9961), .QN(n12980) );
  NOR2X0 U13262 ( .IN1(n9993), .IN2(n11152), .QN(n12979) );
  NAND2X0 U13263 ( .IN1(n10214), .IN2(n8438), .QN(n11152) );
  NAND2X0 U13264 ( .IN1(n12981), .IN2(n12982), .QN(WX7169) );
  NOR2X0 U13265 ( .IN1(n12983), .IN2(n12984), .QN(n12982) );
  NOR2X0 U13266 ( .IN1(n12985), .IN2(n9931), .QN(n12984) );
  NOR2X0 U13267 ( .IN1(n12156), .IN2(n9911), .QN(n12983) );
  INVX0 U13268 ( .INP(n12986), .ZN(n12156) );
  NAND2X0 U13269 ( .IN1(n12987), .IN2(n12988), .QN(n12986) );
  NAND2X0 U13270 ( .IN1(n12989), .IN2(n12990), .QN(n12988) );
  NAND2X0 U13271 ( .IN1(n12991), .IN2(n12992), .QN(n12990) );
  NAND2X0 U13272 ( .IN1(n9309), .IN2(WX8463), .QN(n12992) );
  NAND2X0 U13273 ( .IN1(n9308), .IN2(WX8591), .QN(n12991) );
  NOR2X0 U13274 ( .IN1(n12993), .IN2(n12994), .QN(n12989) );
  NOR2X0 U13275 ( .IN1(n9602), .IN2(WX8527), .QN(n12994) );
  NOR2X0 U13276 ( .IN1(n3597), .IN2(WX8655), .QN(n12993) );
  NAND2X0 U13277 ( .IN1(n12995), .IN2(n12996), .QN(n12987) );
  NAND2X0 U13278 ( .IN1(n12997), .IN2(n12998), .QN(n12996) );
  NAND2X0 U13279 ( .IN1(n9602), .IN2(WX8527), .QN(n12998) );
  NAND2X0 U13280 ( .IN1(n3597), .IN2(WX8655), .QN(n12997) );
  NOR2X0 U13281 ( .IN1(n12999), .IN2(n13000), .QN(n12995) );
  NOR2X0 U13282 ( .IN1(n9309), .IN2(WX8463), .QN(n13000) );
  NOR2X0 U13283 ( .IN1(n9308), .IN2(WX8591), .QN(n12999) );
  NOR2X0 U13284 ( .IN1(n13001), .IN2(n13002), .QN(n12981) );
  NOR2X0 U13285 ( .IN1(DFF_1121_n1), .IN2(n9961), .QN(n13002) );
  NOR2X0 U13286 ( .IN1(n9993), .IN2(n11163), .QN(n13001) );
  NAND2X0 U13287 ( .IN1(n10213), .IN2(n8439), .QN(n11163) );
  NAND2X0 U13288 ( .IN1(n13003), .IN2(n13004), .QN(WX7167) );
  NOR2X0 U13289 ( .IN1(n13005), .IN2(n13006), .QN(n13004) );
  NOR2X0 U13290 ( .IN1(n13007), .IN2(n9931), .QN(n13006) );
  NOR2X0 U13291 ( .IN1(n12174), .IN2(n9911), .QN(n13005) );
  INVX0 U13292 ( .INP(n13008), .ZN(n12174) );
  NAND2X0 U13293 ( .IN1(n13009), .IN2(n13010), .QN(n13008) );
  NAND2X0 U13294 ( .IN1(n13011), .IN2(n13012), .QN(n13010) );
  NAND2X0 U13295 ( .IN1(n13013), .IN2(n13014), .QN(n13012) );
  NAND2X0 U13296 ( .IN1(n9311), .IN2(WX8461), .QN(n13014) );
  NAND2X0 U13297 ( .IN1(n9310), .IN2(WX8589), .QN(n13013) );
  NOR2X0 U13298 ( .IN1(n13015), .IN2(n13016), .QN(n13011) );
  NOR2X0 U13299 ( .IN1(n9601), .IN2(WX8525), .QN(n13016) );
  NOR2X0 U13300 ( .IN1(n3599), .IN2(WX8653), .QN(n13015) );
  NAND2X0 U13301 ( .IN1(n13017), .IN2(n13018), .QN(n13009) );
  NAND2X0 U13302 ( .IN1(n13019), .IN2(n13020), .QN(n13018) );
  NAND2X0 U13303 ( .IN1(n9601), .IN2(WX8525), .QN(n13020) );
  NAND2X0 U13304 ( .IN1(n3599), .IN2(WX8653), .QN(n13019) );
  NOR2X0 U13305 ( .IN1(n13021), .IN2(n13022), .QN(n13017) );
  NOR2X0 U13306 ( .IN1(n9311), .IN2(WX8461), .QN(n13022) );
  NOR2X0 U13307 ( .IN1(n9310), .IN2(WX8589), .QN(n13021) );
  NOR2X0 U13308 ( .IN1(n13023), .IN2(n13024), .QN(n13003) );
  NOR2X0 U13309 ( .IN1(DFF_1122_n1), .IN2(n9961), .QN(n13024) );
  NOR2X0 U13310 ( .IN1(n9993), .IN2(n11164), .QN(n13023) );
  NAND2X0 U13311 ( .IN1(n10212), .IN2(n8440), .QN(n11164) );
  NAND2X0 U13312 ( .IN1(n13025), .IN2(n13026), .QN(WX7165) );
  NOR2X0 U13313 ( .IN1(n13027), .IN2(n13028), .QN(n13026) );
  NOR2X0 U13314 ( .IN1(n13029), .IN2(n9932), .QN(n13028) );
  NOR2X0 U13315 ( .IN1(n12196), .IN2(n9911), .QN(n13027) );
  INVX0 U13316 ( .INP(n13030), .ZN(n12196) );
  NAND2X0 U13317 ( .IN1(n13031), .IN2(n13032), .QN(n13030) );
  NAND2X0 U13318 ( .IN1(n13033), .IN2(n13034), .QN(n13032) );
  NAND2X0 U13319 ( .IN1(n13035), .IN2(n13036), .QN(n13034) );
  NAND2X0 U13320 ( .IN1(n9313), .IN2(WX8459), .QN(n13036) );
  NAND2X0 U13321 ( .IN1(n9312), .IN2(WX8587), .QN(n13035) );
  NOR2X0 U13322 ( .IN1(n13037), .IN2(n13038), .QN(n13033) );
  NOR2X0 U13323 ( .IN1(n9600), .IN2(WX8523), .QN(n13038) );
  NOR2X0 U13324 ( .IN1(n3601), .IN2(WX8651), .QN(n13037) );
  NAND2X0 U13325 ( .IN1(n13039), .IN2(n13040), .QN(n13031) );
  NAND2X0 U13326 ( .IN1(n13041), .IN2(n13042), .QN(n13040) );
  NAND2X0 U13327 ( .IN1(n9600), .IN2(WX8523), .QN(n13042) );
  NAND2X0 U13328 ( .IN1(n3601), .IN2(WX8651), .QN(n13041) );
  NOR2X0 U13329 ( .IN1(n13043), .IN2(n13044), .QN(n13039) );
  NOR2X0 U13330 ( .IN1(n9313), .IN2(WX8459), .QN(n13044) );
  NOR2X0 U13331 ( .IN1(n9312), .IN2(WX8587), .QN(n13043) );
  NOR2X0 U13332 ( .IN1(n13045), .IN2(n13046), .QN(n13025) );
  NOR2X0 U13333 ( .IN1(DFF_1123_n1), .IN2(n9961), .QN(n13046) );
  NOR2X0 U13334 ( .IN1(n9993), .IN2(n11165), .QN(n13045) );
  NAND2X0 U13335 ( .IN1(n10214), .IN2(n8441), .QN(n11165) );
  NAND2X0 U13336 ( .IN1(n13047), .IN2(n13048), .QN(WX7163) );
  NOR2X0 U13337 ( .IN1(n13049), .IN2(n13050), .QN(n13048) );
  NOR2X0 U13338 ( .IN1(n9942), .IN2(n13051), .QN(n13050) );
  NOR2X0 U13339 ( .IN1(n12214), .IN2(n9911), .QN(n13049) );
  INVX0 U13340 ( .INP(n13052), .ZN(n12214) );
  NAND2X0 U13341 ( .IN1(n13053), .IN2(n13054), .QN(n13052) );
  NAND2X0 U13342 ( .IN1(n13055), .IN2(n13056), .QN(n13054) );
  NAND2X0 U13343 ( .IN1(n13057), .IN2(n13058), .QN(n13056) );
  NAND2X0 U13344 ( .IN1(n9315), .IN2(WX8457), .QN(n13058) );
  NAND2X0 U13345 ( .IN1(n9314), .IN2(WX8585), .QN(n13057) );
  NOR2X0 U13346 ( .IN1(n13059), .IN2(n13060), .QN(n13055) );
  NOR2X0 U13347 ( .IN1(n9504), .IN2(WX8521), .QN(n13060) );
  NOR2X0 U13348 ( .IN1(n3603), .IN2(WX8649), .QN(n13059) );
  NAND2X0 U13349 ( .IN1(n13061), .IN2(n13062), .QN(n13053) );
  NAND2X0 U13350 ( .IN1(n13063), .IN2(n13064), .QN(n13062) );
  NAND2X0 U13351 ( .IN1(n9504), .IN2(WX8521), .QN(n13064) );
  NAND2X0 U13352 ( .IN1(n3603), .IN2(WX8649), .QN(n13063) );
  NOR2X0 U13353 ( .IN1(n13065), .IN2(n13066), .QN(n13061) );
  NOR2X0 U13354 ( .IN1(n9315), .IN2(WX8457), .QN(n13066) );
  NOR2X0 U13355 ( .IN1(n9314), .IN2(WX8585), .QN(n13065) );
  NOR2X0 U13356 ( .IN1(n13067), .IN2(n13068), .QN(n13047) );
  NOR2X0 U13357 ( .IN1(DFF_1124_n1), .IN2(n9961), .QN(n13068) );
  NOR2X0 U13358 ( .IN1(n9993), .IN2(n11166), .QN(n13067) );
  NAND2X0 U13359 ( .IN1(n10213), .IN2(n8442), .QN(n11166) );
  NAND2X0 U13360 ( .IN1(n13069), .IN2(n13070), .QN(WX7161) );
  NOR2X0 U13361 ( .IN1(n13071), .IN2(n13072), .QN(n13070) );
  NOR2X0 U13362 ( .IN1(n13073), .IN2(n9932), .QN(n13072) );
  NOR2X0 U13363 ( .IN1(n12236), .IN2(n9911), .QN(n13071) );
  INVX0 U13364 ( .INP(n13074), .ZN(n12236) );
  NAND2X0 U13365 ( .IN1(n13075), .IN2(n13076), .QN(n13074) );
  NAND2X0 U13366 ( .IN1(n13077), .IN2(n13078), .QN(n13076) );
  NAND2X0 U13367 ( .IN1(n13079), .IN2(n13080), .QN(n13078) );
  NAND2X0 U13368 ( .IN1(n9317), .IN2(WX8455), .QN(n13080) );
  NAND2X0 U13369 ( .IN1(n9316), .IN2(WX8583), .QN(n13079) );
  NOR2X0 U13370 ( .IN1(n13081), .IN2(n13082), .QN(n13077) );
  NOR2X0 U13371 ( .IN1(n9599), .IN2(WX8519), .QN(n13082) );
  NOR2X0 U13372 ( .IN1(n3605), .IN2(WX8647), .QN(n13081) );
  NAND2X0 U13373 ( .IN1(n13083), .IN2(n13084), .QN(n13075) );
  NAND2X0 U13374 ( .IN1(n13085), .IN2(n13086), .QN(n13084) );
  NAND2X0 U13375 ( .IN1(n9599), .IN2(WX8519), .QN(n13086) );
  NAND2X0 U13376 ( .IN1(n3605), .IN2(WX8647), .QN(n13085) );
  NOR2X0 U13377 ( .IN1(n13087), .IN2(n13088), .QN(n13083) );
  NOR2X0 U13378 ( .IN1(n9317), .IN2(WX8455), .QN(n13088) );
  NOR2X0 U13379 ( .IN1(n9316), .IN2(WX8583), .QN(n13087) );
  NOR2X0 U13380 ( .IN1(n13089), .IN2(n13090), .QN(n13069) );
  NOR2X0 U13381 ( .IN1(DFF_1125_n1), .IN2(n9961), .QN(n13090) );
  NOR2X0 U13382 ( .IN1(n9993), .IN2(n11167), .QN(n13089) );
  NAND2X0 U13383 ( .IN1(n10213), .IN2(n8443), .QN(n11167) );
  NAND2X0 U13384 ( .IN1(n13091), .IN2(n13092), .QN(WX7159) );
  NOR2X0 U13385 ( .IN1(n13093), .IN2(n13094), .QN(n13092) );
  NOR2X0 U13386 ( .IN1(n9942), .IN2(n13095), .QN(n13094) );
  NOR2X0 U13387 ( .IN1(n12258), .IN2(n9911), .QN(n13093) );
  INVX0 U13388 ( .INP(n13096), .ZN(n12258) );
  NAND2X0 U13389 ( .IN1(n13097), .IN2(n13098), .QN(n13096) );
  NAND2X0 U13390 ( .IN1(n13099), .IN2(n13100), .QN(n13098) );
  NAND2X0 U13391 ( .IN1(n13101), .IN2(n13102), .QN(n13100) );
  NAND2X0 U13392 ( .IN1(n9319), .IN2(WX8453), .QN(n13102) );
  NAND2X0 U13393 ( .IN1(n9318), .IN2(WX8581), .QN(n13101) );
  NOR2X0 U13394 ( .IN1(n13103), .IN2(n13104), .QN(n13099) );
  NOR2X0 U13395 ( .IN1(n9598), .IN2(WX8517), .QN(n13104) );
  NOR2X0 U13396 ( .IN1(n3607), .IN2(WX8645), .QN(n13103) );
  NAND2X0 U13397 ( .IN1(n13105), .IN2(n13106), .QN(n13097) );
  NAND2X0 U13398 ( .IN1(n13107), .IN2(n13108), .QN(n13106) );
  NAND2X0 U13399 ( .IN1(n9598), .IN2(WX8517), .QN(n13108) );
  NAND2X0 U13400 ( .IN1(n3607), .IN2(WX8645), .QN(n13107) );
  NOR2X0 U13401 ( .IN1(n13109), .IN2(n13110), .QN(n13105) );
  NOR2X0 U13402 ( .IN1(n9319), .IN2(WX8453), .QN(n13110) );
  NOR2X0 U13403 ( .IN1(n9318), .IN2(WX8581), .QN(n13109) );
  NOR2X0 U13404 ( .IN1(n13111), .IN2(n13112), .QN(n13091) );
  NOR2X0 U13405 ( .IN1(DFF_1126_n1), .IN2(n9961), .QN(n13112) );
  NOR2X0 U13406 ( .IN1(n9993), .IN2(n11168), .QN(n13111) );
  NAND2X0 U13407 ( .IN1(n10213), .IN2(n8444), .QN(n11168) );
  NAND2X0 U13408 ( .IN1(n13113), .IN2(n13114), .QN(WX7157) );
  NOR2X0 U13409 ( .IN1(n13115), .IN2(n13116), .QN(n13114) );
  NOR2X0 U13410 ( .IN1(n13117), .IN2(n9932), .QN(n13116) );
  NOR2X0 U13411 ( .IN1(n12280), .IN2(n9911), .QN(n13115) );
  INVX0 U13412 ( .INP(n13118), .ZN(n12280) );
  NAND2X0 U13413 ( .IN1(n13119), .IN2(n13120), .QN(n13118) );
  NAND2X0 U13414 ( .IN1(n13121), .IN2(n13122), .QN(n13120) );
  NAND2X0 U13415 ( .IN1(n13123), .IN2(n13124), .QN(n13122) );
  NAND2X0 U13416 ( .IN1(n9321), .IN2(WX8451), .QN(n13124) );
  NAND2X0 U13417 ( .IN1(n9320), .IN2(WX8579), .QN(n13123) );
  NOR2X0 U13418 ( .IN1(n13125), .IN2(n13126), .QN(n13121) );
  NOR2X0 U13419 ( .IN1(n9597), .IN2(WX8515), .QN(n13126) );
  NOR2X0 U13420 ( .IN1(n3609), .IN2(WX8643), .QN(n13125) );
  NAND2X0 U13421 ( .IN1(n13127), .IN2(n13128), .QN(n13119) );
  NAND2X0 U13422 ( .IN1(n13129), .IN2(n13130), .QN(n13128) );
  NAND2X0 U13423 ( .IN1(n9597), .IN2(WX8515), .QN(n13130) );
  NAND2X0 U13424 ( .IN1(n3609), .IN2(WX8643), .QN(n13129) );
  NOR2X0 U13425 ( .IN1(n13131), .IN2(n13132), .QN(n13127) );
  NOR2X0 U13426 ( .IN1(n9321), .IN2(WX8451), .QN(n13132) );
  NOR2X0 U13427 ( .IN1(n9320), .IN2(WX8579), .QN(n13131) );
  NOR2X0 U13428 ( .IN1(n13133), .IN2(n13134), .QN(n13113) );
  NOR2X0 U13429 ( .IN1(DFF_1127_n1), .IN2(n9961), .QN(n13134) );
  NOR2X0 U13430 ( .IN1(n9993), .IN2(n11169), .QN(n13133) );
  NAND2X0 U13431 ( .IN1(n10213), .IN2(n8445), .QN(n11169) );
  NAND2X0 U13432 ( .IN1(n13135), .IN2(n13136), .QN(WX7155) );
  NOR2X0 U13433 ( .IN1(n13137), .IN2(n13138), .QN(n13136) );
  NOR2X0 U13434 ( .IN1(n9942), .IN2(n13139), .QN(n13138) );
  NOR2X0 U13435 ( .IN1(n12302), .IN2(n9911), .QN(n13137) );
  INVX0 U13436 ( .INP(n13140), .ZN(n12302) );
  NAND2X0 U13437 ( .IN1(n13141), .IN2(n13142), .QN(n13140) );
  NAND2X0 U13438 ( .IN1(n13143), .IN2(n13144), .QN(n13142) );
  NAND2X0 U13439 ( .IN1(n13145), .IN2(n13146), .QN(n13144) );
  NAND2X0 U13440 ( .IN1(n9323), .IN2(WX8449), .QN(n13146) );
  NAND2X0 U13441 ( .IN1(n9322), .IN2(WX8577), .QN(n13145) );
  NOR2X0 U13442 ( .IN1(n13147), .IN2(n13148), .QN(n13143) );
  NOR2X0 U13443 ( .IN1(n9596), .IN2(WX8513), .QN(n13148) );
  NOR2X0 U13444 ( .IN1(n3611), .IN2(WX8641), .QN(n13147) );
  NAND2X0 U13445 ( .IN1(n13149), .IN2(n13150), .QN(n13141) );
  NAND2X0 U13446 ( .IN1(n13151), .IN2(n13152), .QN(n13150) );
  NAND2X0 U13447 ( .IN1(n9596), .IN2(WX8513), .QN(n13152) );
  NAND2X0 U13448 ( .IN1(n3611), .IN2(WX8641), .QN(n13151) );
  NOR2X0 U13449 ( .IN1(n13153), .IN2(n13154), .QN(n13149) );
  NOR2X0 U13450 ( .IN1(n9323), .IN2(WX8449), .QN(n13154) );
  NOR2X0 U13451 ( .IN1(n9322), .IN2(WX8577), .QN(n13153) );
  NOR2X0 U13452 ( .IN1(n13155), .IN2(n13156), .QN(n13135) );
  NOR2X0 U13453 ( .IN1(DFF_1128_n1), .IN2(n9961), .QN(n13156) );
  NOR2X0 U13454 ( .IN1(n9993), .IN2(n11170), .QN(n13155) );
  NAND2X0 U13455 ( .IN1(n10212), .IN2(n8446), .QN(n11170) );
  NAND2X0 U13456 ( .IN1(n13157), .IN2(n13158), .QN(WX7153) );
  NOR2X0 U13457 ( .IN1(n13159), .IN2(n13160), .QN(n13158) );
  NOR2X0 U13458 ( .IN1(n13161), .IN2(n9932), .QN(n13160) );
  NOR2X0 U13459 ( .IN1(n9921), .IN2(n12324), .QN(n13159) );
  NAND2X0 U13460 ( .IN1(n13162), .IN2(n13163), .QN(n12324) );
  INVX0 U13461 ( .INP(n13164), .ZN(n13163) );
  NOR2X0 U13462 ( .IN1(n13165), .IN2(n13166), .QN(n13164) );
  NAND2X0 U13463 ( .IN1(n13166), .IN2(n13165), .QN(n13162) );
  NOR2X0 U13464 ( .IN1(n13167), .IN2(n13168), .QN(n13165) );
  NOR2X0 U13465 ( .IN1(n9834), .IN2(n9325), .QN(n13168) );
  INVX0 U13466 ( .INP(n13169), .ZN(n13167) );
  NAND2X0 U13467 ( .IN1(n9325), .IN2(n9834), .QN(n13169) );
  NAND2X0 U13468 ( .IN1(n13170), .IN2(n13171), .QN(n13166) );
  NAND2X0 U13469 ( .IN1(n9324), .IN2(WX8511), .QN(n13171) );
  INVX0 U13470 ( .INP(n13172), .ZN(n13170) );
  NOR2X0 U13471 ( .IN1(WX8511), .IN2(n9324), .QN(n13172) );
  NOR2X0 U13472 ( .IN1(n13173), .IN2(n13174), .QN(n13157) );
  NOR2X0 U13473 ( .IN1(DFF_1129_n1), .IN2(n9961), .QN(n13174) );
  NOR2X0 U13474 ( .IN1(n9993), .IN2(n11171), .QN(n13173) );
  NAND2X0 U13475 ( .IN1(n10212), .IN2(n8447), .QN(n11171) );
  NAND2X0 U13476 ( .IN1(n13175), .IN2(n13176), .QN(WX7151) );
  NOR2X0 U13477 ( .IN1(n13177), .IN2(n13178), .QN(n13176) );
  NOR2X0 U13478 ( .IN1(n9941), .IN2(n13179), .QN(n13178) );
  NOR2X0 U13479 ( .IN1(n12346), .IN2(n9911), .QN(n13177) );
  INVX0 U13480 ( .INP(n13180), .ZN(n12346) );
  NAND2X0 U13481 ( .IN1(n13181), .IN2(n13182), .QN(n13180) );
  NAND2X0 U13482 ( .IN1(n13183), .IN2(n13184), .QN(n13182) );
  NAND2X0 U13483 ( .IN1(n13185), .IN2(n13186), .QN(n13184) );
  NAND2X0 U13484 ( .IN1(n9327), .IN2(WX8445), .QN(n13186) );
  NAND2X0 U13485 ( .IN1(n9326), .IN2(WX8573), .QN(n13185) );
  NOR2X0 U13486 ( .IN1(n13187), .IN2(n13188), .QN(n13183) );
  NOR2X0 U13487 ( .IN1(n9595), .IN2(WX8509), .QN(n13188) );
  NOR2X0 U13488 ( .IN1(n3615), .IN2(WX8637), .QN(n13187) );
  NAND2X0 U13489 ( .IN1(n13189), .IN2(n13190), .QN(n13181) );
  NAND2X0 U13490 ( .IN1(n13191), .IN2(n13192), .QN(n13190) );
  NAND2X0 U13491 ( .IN1(n9595), .IN2(WX8509), .QN(n13192) );
  NAND2X0 U13492 ( .IN1(n3615), .IN2(WX8637), .QN(n13191) );
  NOR2X0 U13493 ( .IN1(n13193), .IN2(n13194), .QN(n13189) );
  NOR2X0 U13494 ( .IN1(n9327), .IN2(WX8445), .QN(n13194) );
  NOR2X0 U13495 ( .IN1(n9326), .IN2(WX8573), .QN(n13193) );
  NOR2X0 U13496 ( .IN1(n13195), .IN2(n13196), .QN(n13175) );
  NOR2X0 U13497 ( .IN1(DFF_1130_n1), .IN2(n9961), .QN(n13196) );
  NOR2X0 U13498 ( .IN1(n9993), .IN2(n11172), .QN(n13195) );
  NAND2X0 U13499 ( .IN1(n10213), .IN2(n8448), .QN(n11172) );
  NAND2X0 U13500 ( .IN1(n13197), .IN2(n13198), .QN(WX7149) );
  NOR2X0 U13501 ( .IN1(n13199), .IN2(n13200), .QN(n13198) );
  NOR2X0 U13502 ( .IN1(n13201), .IN2(n9932), .QN(n13200) );
  NOR2X0 U13503 ( .IN1(n9921), .IN2(n12368), .QN(n13199) );
  NAND2X0 U13504 ( .IN1(n13202), .IN2(n13203), .QN(n12368) );
  INVX0 U13505 ( .INP(n13204), .ZN(n13203) );
  NOR2X0 U13506 ( .IN1(n13205), .IN2(n13206), .QN(n13204) );
  NAND2X0 U13507 ( .IN1(n13206), .IN2(n13205), .QN(n13202) );
  NOR2X0 U13508 ( .IN1(n13207), .IN2(n13208), .QN(n13205) );
  INVX0 U13509 ( .INP(n13209), .ZN(n13208) );
  NAND2X0 U13510 ( .IN1(test_so73), .IN2(WX8635), .QN(n13209) );
  NOR2X0 U13511 ( .IN1(WX8635), .IN2(test_so73), .QN(n13207) );
  NAND2X0 U13512 ( .IN1(n13210), .IN2(n13211), .QN(n13206) );
  NAND2X0 U13513 ( .IN1(n9328), .IN2(WX8507), .QN(n13211) );
  INVX0 U13514 ( .INP(n13212), .ZN(n13210) );
  NOR2X0 U13515 ( .IN1(WX8507), .IN2(n9328), .QN(n13212) );
  NOR2X0 U13516 ( .IN1(n13213), .IN2(n13214), .QN(n13197) );
  NOR2X0 U13517 ( .IN1(DFF_1131_n1), .IN2(n9961), .QN(n13214) );
  NOR2X0 U13518 ( .IN1(n9992), .IN2(n11173), .QN(n13213) );
  NAND2X0 U13519 ( .IN1(n10211), .IN2(n8449), .QN(n11173) );
  NAND2X0 U13520 ( .IN1(n13215), .IN2(n13216), .QN(WX7147) );
  NOR2X0 U13521 ( .IN1(n13217), .IN2(n13218), .QN(n13216) );
  NOR2X0 U13522 ( .IN1(n13219), .IN2(n9932), .QN(n13218) );
  NOR2X0 U13523 ( .IN1(n12390), .IN2(n9911), .QN(n13217) );
  INVX0 U13524 ( .INP(n13220), .ZN(n12390) );
  NAND2X0 U13525 ( .IN1(n13221), .IN2(n13222), .QN(n13220) );
  NAND2X0 U13526 ( .IN1(n13223), .IN2(n13224), .QN(n13222) );
  NAND2X0 U13527 ( .IN1(n13225), .IN2(n13226), .QN(n13224) );
  NAND2X0 U13528 ( .IN1(n9330), .IN2(WX8441), .QN(n13226) );
  NAND2X0 U13529 ( .IN1(n9329), .IN2(WX8569), .QN(n13225) );
  NOR2X0 U13530 ( .IN1(n13227), .IN2(n13228), .QN(n13223) );
  NOR2X0 U13531 ( .IN1(n9594), .IN2(WX8505), .QN(n13228) );
  NOR2X0 U13532 ( .IN1(n3619), .IN2(WX8633), .QN(n13227) );
  NAND2X0 U13533 ( .IN1(n13229), .IN2(n13230), .QN(n13221) );
  NAND2X0 U13534 ( .IN1(n13231), .IN2(n13232), .QN(n13230) );
  NAND2X0 U13535 ( .IN1(n9594), .IN2(WX8505), .QN(n13232) );
  NAND2X0 U13536 ( .IN1(n3619), .IN2(WX8633), .QN(n13231) );
  NOR2X0 U13537 ( .IN1(n13233), .IN2(n13234), .QN(n13229) );
  NOR2X0 U13538 ( .IN1(n9330), .IN2(WX8441), .QN(n13234) );
  NOR2X0 U13539 ( .IN1(n9329), .IN2(WX8569), .QN(n13233) );
  NOR2X0 U13540 ( .IN1(n13235), .IN2(n13236), .QN(n13215) );
  NOR2X0 U13541 ( .IN1(n9976), .IN2(n9854), .QN(n13236) );
  NOR2X0 U13542 ( .IN1(n9992), .IN2(n11174), .QN(n13235) );
  NAND2X0 U13543 ( .IN1(test_so56), .IN2(n10215), .QN(n11174) );
  NAND2X0 U13544 ( .IN1(n13237), .IN2(n13238), .QN(WX7145) );
  NOR2X0 U13545 ( .IN1(n13239), .IN2(n13240), .QN(n13238) );
  NOR2X0 U13546 ( .IN1(n13241), .IN2(n9932), .QN(n13240) );
  NOR2X0 U13547 ( .IN1(n9922), .IN2(n12412), .QN(n13239) );
  NAND2X0 U13548 ( .IN1(n13242), .IN2(n13243), .QN(n12412) );
  INVX0 U13549 ( .INP(n13244), .ZN(n13243) );
  NOR2X0 U13550 ( .IN1(n13245), .IN2(n13246), .QN(n13244) );
  NAND2X0 U13551 ( .IN1(n13246), .IN2(n13245), .QN(n13242) );
  NOR2X0 U13552 ( .IN1(n13247), .IN2(n13248), .QN(n13245) );
  INVX0 U13553 ( .INP(n13249), .ZN(n13248) );
  NAND2X0 U13554 ( .IN1(test_so71), .IN2(WX8631), .QN(n13249) );
  NOR2X0 U13555 ( .IN1(WX8631), .IN2(test_so71), .QN(n13247) );
  NAND2X0 U13556 ( .IN1(n13250), .IN2(n13251), .QN(n13246) );
  NAND2X0 U13557 ( .IN1(n9332), .IN2(WX8439), .QN(n13251) );
  INVX0 U13558 ( .INP(n13252), .ZN(n13250) );
  NOR2X0 U13559 ( .IN1(WX8439), .IN2(n9332), .QN(n13252) );
  NOR2X0 U13560 ( .IN1(n13253), .IN2(n13254), .QN(n13237) );
  NOR2X0 U13561 ( .IN1(DFF_1133_n1), .IN2(n9960), .QN(n13254) );
  NOR2X0 U13562 ( .IN1(n9992), .IN2(n11175), .QN(n13253) );
  NAND2X0 U13563 ( .IN1(n10213), .IN2(n8452), .QN(n11175) );
  NAND2X0 U13564 ( .IN1(n13255), .IN2(n13256), .QN(WX7143) );
  NOR2X0 U13565 ( .IN1(n13257), .IN2(n13258), .QN(n13256) );
  NOR2X0 U13566 ( .IN1(n13259), .IN2(n9932), .QN(n13258) );
  NOR2X0 U13567 ( .IN1(n12434), .IN2(n9912), .QN(n13257) );
  INVX0 U13568 ( .INP(n13260), .ZN(n12434) );
  NAND2X0 U13569 ( .IN1(n13261), .IN2(n13262), .QN(n13260) );
  NAND2X0 U13570 ( .IN1(n13263), .IN2(n13264), .QN(n13262) );
  NAND2X0 U13571 ( .IN1(n13265), .IN2(n13266), .QN(n13264) );
  NAND2X0 U13572 ( .IN1(n9334), .IN2(WX8437), .QN(n13266) );
  NAND2X0 U13573 ( .IN1(n9333), .IN2(WX8565), .QN(n13265) );
  NOR2X0 U13574 ( .IN1(n13267), .IN2(n13268), .QN(n13263) );
  NOR2X0 U13575 ( .IN1(n9592), .IN2(WX8501), .QN(n13268) );
  NOR2X0 U13576 ( .IN1(n3623), .IN2(WX8629), .QN(n13267) );
  NAND2X0 U13577 ( .IN1(n13269), .IN2(n13270), .QN(n13261) );
  NAND2X0 U13578 ( .IN1(n13271), .IN2(n13272), .QN(n13270) );
  NAND2X0 U13579 ( .IN1(n9592), .IN2(WX8501), .QN(n13272) );
  NAND2X0 U13580 ( .IN1(n3623), .IN2(WX8629), .QN(n13271) );
  NOR2X0 U13581 ( .IN1(n13273), .IN2(n13274), .QN(n13269) );
  NOR2X0 U13582 ( .IN1(n9334), .IN2(WX8437), .QN(n13274) );
  NOR2X0 U13583 ( .IN1(n9333), .IN2(WX8565), .QN(n13273) );
  NOR2X0 U13584 ( .IN1(n13275), .IN2(n13276), .QN(n13255) );
  NOR2X0 U13585 ( .IN1(DFF_1134_n1), .IN2(n9960), .QN(n13276) );
  NOR2X0 U13586 ( .IN1(n9992), .IN2(n11176), .QN(n13275) );
  NAND2X0 U13587 ( .IN1(n10213), .IN2(n8453), .QN(n11176) );
  NAND2X0 U13588 ( .IN1(n13277), .IN2(n13278), .QN(WX7141) );
  NOR2X0 U13589 ( .IN1(n13279), .IN2(n13280), .QN(n13278) );
  NOR2X0 U13590 ( .IN1(n13281), .IN2(n9932), .QN(n13280) );
  NOR2X0 U13591 ( .IN1(n9921), .IN2(n12452), .QN(n13279) );
  NAND2X0 U13592 ( .IN1(n13282), .IN2(n13283), .QN(n12452) );
  INVX0 U13593 ( .INP(n13284), .ZN(n13283) );
  NOR2X0 U13594 ( .IN1(n13285), .IN2(n13286), .QN(n13284) );
  NAND2X0 U13595 ( .IN1(n13286), .IN2(n13285), .QN(n13282) );
  NOR2X0 U13596 ( .IN1(n13287), .IN2(n13288), .QN(n13285) );
  INVX0 U13597 ( .INP(n13289), .ZN(n13288) );
  NAND2X0 U13598 ( .IN1(test_so69), .IN2(WX8627), .QN(n13289) );
  NOR2X0 U13599 ( .IN1(WX8627), .IN2(test_so69), .QN(n13287) );
  NAND2X0 U13600 ( .IN1(n13290), .IN2(n13291), .QN(n13286) );
  NAND2X0 U13601 ( .IN1(n9335), .IN2(WX8499), .QN(n13291) );
  INVX0 U13602 ( .INP(n13292), .ZN(n13290) );
  NOR2X0 U13603 ( .IN1(WX8499), .IN2(n9335), .QN(n13292) );
  NOR2X0 U13604 ( .IN1(n13293), .IN2(n13294), .QN(n13277) );
  NOR2X0 U13605 ( .IN1(DFF_1135_n1), .IN2(n9960), .QN(n13294) );
  NOR2X0 U13606 ( .IN1(n9992), .IN2(n11177), .QN(n13293) );
  NAND2X0 U13607 ( .IN1(n10212), .IN2(n8454), .QN(n11177) );
  NAND2X0 U13608 ( .IN1(n13295), .IN2(n13296), .QN(WX7139) );
  NOR2X0 U13609 ( .IN1(n13297), .IN2(n13298), .QN(n13296) );
  NOR2X0 U13610 ( .IN1(n13299), .IN2(n9932), .QN(n13298) );
  NOR2X0 U13611 ( .IN1(n12474), .IN2(n9912), .QN(n13297) );
  NOR2X0 U13612 ( .IN1(n13300), .IN2(n13301), .QN(n12474) );
  INVX0 U13613 ( .INP(n13302), .ZN(n13301) );
  NAND2X0 U13614 ( .IN1(n13303), .IN2(n13304), .QN(n13302) );
  NOR2X0 U13615 ( .IN1(n13304), .IN2(n13303), .QN(n13300) );
  NAND2X0 U13616 ( .IN1(n13305), .IN2(n13306), .QN(n13303) );
  NAND2X0 U13617 ( .IN1(n9076), .IN2(n13307), .QN(n13306) );
  INVX0 U13618 ( .INP(n13308), .ZN(n13305) );
  NOR2X0 U13619 ( .IN1(n13307), .IN2(n9076), .QN(n13308) );
  NOR2X0 U13620 ( .IN1(n13309), .IN2(n13310), .QN(n13307) );
  INVX0 U13621 ( .INP(n13311), .ZN(n13310) );
  NAND2X0 U13622 ( .IN1(n18442), .IN2(WX8625), .QN(n13311) );
  NOR2X0 U13623 ( .IN1(WX8625), .IN2(n18442), .QN(n13309) );
  NOR2X0 U13624 ( .IN1(n13312), .IN2(n13313), .QN(n13304) );
  INVX0 U13625 ( .INP(n13314), .ZN(n13313) );
  NAND2X0 U13626 ( .IN1(n9075), .IN2(n10014), .QN(n13314) );
  NOR2X0 U13627 ( .IN1(n10005), .IN2(n9075), .QN(n13312) );
  NOR2X0 U13628 ( .IN1(n13315), .IN2(n13316), .QN(n13295) );
  NOR2X0 U13629 ( .IN1(DFF_1136_n1), .IN2(n9960), .QN(n13316) );
  NOR2X0 U13630 ( .IN1(n9992), .IN2(n11178), .QN(n13315) );
  NAND2X0 U13631 ( .IN1(n10212), .IN2(n8455), .QN(n11178) );
  NAND2X0 U13632 ( .IN1(n13317), .IN2(n13318), .QN(WX7137) );
  NOR2X0 U13633 ( .IN1(n13319), .IN2(n13320), .QN(n13318) );
  NOR2X0 U13634 ( .IN1(n13321), .IN2(n9932), .QN(n13320) );
  NOR2X0 U13635 ( .IN1(n12496), .IN2(n9912), .QN(n13319) );
  NOR2X0 U13636 ( .IN1(n13322), .IN2(n13323), .QN(n12496) );
  INVX0 U13637 ( .INP(n13324), .ZN(n13323) );
  NAND2X0 U13638 ( .IN1(n13325), .IN2(n13326), .QN(n13324) );
  NOR2X0 U13639 ( .IN1(n13326), .IN2(n13325), .QN(n13322) );
  NAND2X0 U13640 ( .IN1(n13327), .IN2(n13328), .QN(n13325) );
  NAND2X0 U13641 ( .IN1(n9078), .IN2(n13329), .QN(n13328) );
  INVX0 U13642 ( .INP(n13330), .ZN(n13327) );
  NOR2X0 U13643 ( .IN1(n13329), .IN2(n9078), .QN(n13330) );
  NOR2X0 U13644 ( .IN1(n13331), .IN2(n13332), .QN(n13329) );
  INVX0 U13645 ( .INP(n13333), .ZN(n13332) );
  NAND2X0 U13646 ( .IN1(n18441), .IN2(WX8623), .QN(n13333) );
  NOR2X0 U13647 ( .IN1(WX8623), .IN2(n18441), .QN(n13331) );
  NOR2X0 U13648 ( .IN1(n13334), .IN2(n13335), .QN(n13326) );
  INVX0 U13649 ( .INP(n13336), .ZN(n13335) );
  NAND2X0 U13650 ( .IN1(n9077), .IN2(n10013), .QN(n13336) );
  NOR2X0 U13651 ( .IN1(n10005), .IN2(n9077), .QN(n13334) );
  NOR2X0 U13652 ( .IN1(n13337), .IN2(n13338), .QN(n13317) );
  NOR2X0 U13653 ( .IN1(DFF_1137_n1), .IN2(n9960), .QN(n13338) );
  NOR2X0 U13654 ( .IN1(n9992), .IN2(n11179), .QN(n13337) );
  NAND2X0 U13655 ( .IN1(n10212), .IN2(n8456), .QN(n11179) );
  NAND2X0 U13656 ( .IN1(n13339), .IN2(n13340), .QN(WX7135) );
  NOR2X0 U13657 ( .IN1(n13341), .IN2(n13342), .QN(n13340) );
  NOR2X0 U13658 ( .IN1(n13343), .IN2(n9932), .QN(n13342) );
  NOR2X0 U13659 ( .IN1(n12518), .IN2(n9912), .QN(n13341) );
  NOR2X0 U13660 ( .IN1(n13344), .IN2(n13345), .QN(n12518) );
  INVX0 U13661 ( .INP(n13346), .ZN(n13345) );
  NAND2X0 U13662 ( .IN1(n13347), .IN2(n13348), .QN(n13346) );
  NOR2X0 U13663 ( .IN1(n13348), .IN2(n13347), .QN(n13344) );
  NAND2X0 U13664 ( .IN1(n13349), .IN2(n13350), .QN(n13347) );
  NAND2X0 U13665 ( .IN1(n9080), .IN2(n13351), .QN(n13350) );
  INVX0 U13666 ( .INP(n13352), .ZN(n13349) );
  NOR2X0 U13667 ( .IN1(n13351), .IN2(n9080), .QN(n13352) );
  NOR2X0 U13668 ( .IN1(n13353), .IN2(n13354), .QN(n13351) );
  INVX0 U13669 ( .INP(n13355), .ZN(n13354) );
  NAND2X0 U13670 ( .IN1(n18440), .IN2(WX8621), .QN(n13355) );
  NOR2X0 U13671 ( .IN1(WX8621), .IN2(n18440), .QN(n13353) );
  NOR2X0 U13672 ( .IN1(n13356), .IN2(n13357), .QN(n13348) );
  INVX0 U13673 ( .INP(n13358), .ZN(n13357) );
  NAND2X0 U13674 ( .IN1(n9079), .IN2(n10013), .QN(n13358) );
  NOR2X0 U13675 ( .IN1(n10005), .IN2(n9079), .QN(n13356) );
  NOR2X0 U13676 ( .IN1(n13359), .IN2(n13360), .QN(n13339) );
  NOR2X0 U13677 ( .IN1(DFF_1138_n1), .IN2(n9960), .QN(n13360) );
  NOR2X0 U13678 ( .IN1(n9992), .IN2(n11180), .QN(n13359) );
  NAND2X0 U13679 ( .IN1(n10212), .IN2(n8457), .QN(n11180) );
  NAND2X0 U13680 ( .IN1(n13361), .IN2(n13362), .QN(WX7133) );
  NOR2X0 U13681 ( .IN1(n13363), .IN2(n13364), .QN(n13362) );
  NOR2X0 U13682 ( .IN1(n13365), .IN2(n9933), .QN(n13364) );
  NOR2X0 U13683 ( .IN1(n12540), .IN2(n9912), .QN(n13363) );
  NOR2X0 U13684 ( .IN1(n13366), .IN2(n13367), .QN(n12540) );
  INVX0 U13685 ( .INP(n13368), .ZN(n13367) );
  NAND2X0 U13686 ( .IN1(n13369), .IN2(n13370), .QN(n13368) );
  NOR2X0 U13687 ( .IN1(n13370), .IN2(n13369), .QN(n13366) );
  NAND2X0 U13688 ( .IN1(n13371), .IN2(n13372), .QN(n13369) );
  NAND2X0 U13689 ( .IN1(n9082), .IN2(n13373), .QN(n13372) );
  INVX0 U13690 ( .INP(n13374), .ZN(n13371) );
  NOR2X0 U13691 ( .IN1(n13373), .IN2(n9082), .QN(n13374) );
  NOR2X0 U13692 ( .IN1(n13375), .IN2(n13376), .QN(n13373) );
  INVX0 U13693 ( .INP(n13377), .ZN(n13376) );
  NAND2X0 U13694 ( .IN1(n18439), .IN2(WX8619), .QN(n13377) );
  NOR2X0 U13695 ( .IN1(WX8619), .IN2(n18439), .QN(n13375) );
  NOR2X0 U13696 ( .IN1(n13378), .IN2(n13379), .QN(n13370) );
  INVX0 U13697 ( .INP(n13380), .ZN(n13379) );
  NAND2X0 U13698 ( .IN1(n9081), .IN2(n10014), .QN(n13380) );
  NOR2X0 U13699 ( .IN1(n10005), .IN2(n9081), .QN(n13378) );
  NOR2X0 U13700 ( .IN1(n13381), .IN2(n13382), .QN(n13361) );
  NOR2X0 U13701 ( .IN1(DFF_1139_n1), .IN2(n9960), .QN(n13382) );
  NOR2X0 U13702 ( .IN1(n9992), .IN2(n11181), .QN(n13381) );
  NAND2X0 U13703 ( .IN1(n10212), .IN2(n8458), .QN(n11181) );
  NAND2X0 U13704 ( .IN1(n13383), .IN2(n13384), .QN(WX7131) );
  NOR2X0 U13705 ( .IN1(n13385), .IN2(n13386), .QN(n13384) );
  NOR2X0 U13706 ( .IN1(n13387), .IN2(n9933), .QN(n13386) );
  NOR2X0 U13707 ( .IN1(n12562), .IN2(n9912), .QN(n13385) );
  NOR2X0 U13708 ( .IN1(n13388), .IN2(n13389), .QN(n12562) );
  INVX0 U13709 ( .INP(n13390), .ZN(n13389) );
  NAND2X0 U13710 ( .IN1(n13391), .IN2(n13392), .QN(n13390) );
  NOR2X0 U13711 ( .IN1(n13392), .IN2(n13391), .QN(n13388) );
  NAND2X0 U13712 ( .IN1(n13393), .IN2(n13394), .QN(n13391) );
  NAND2X0 U13713 ( .IN1(n9084), .IN2(n13395), .QN(n13394) );
  INVX0 U13714 ( .INP(n13396), .ZN(n13393) );
  NOR2X0 U13715 ( .IN1(n13395), .IN2(n9084), .QN(n13396) );
  NOR2X0 U13716 ( .IN1(n13397), .IN2(n13398), .QN(n13395) );
  INVX0 U13717 ( .INP(n13399), .ZN(n13398) );
  NAND2X0 U13718 ( .IN1(n18438), .IN2(WX8617), .QN(n13399) );
  NOR2X0 U13719 ( .IN1(WX8617), .IN2(n18438), .QN(n13397) );
  NOR2X0 U13720 ( .IN1(n13400), .IN2(n13401), .QN(n13392) );
  INVX0 U13721 ( .INP(n13402), .ZN(n13401) );
  NAND2X0 U13722 ( .IN1(n9083), .IN2(n10014), .QN(n13402) );
  NOR2X0 U13723 ( .IN1(n10006), .IN2(n9083), .QN(n13400) );
  NOR2X0 U13724 ( .IN1(n13403), .IN2(n13404), .QN(n13383) );
  NOR2X0 U13725 ( .IN1(DFF_1140_n1), .IN2(n9960), .QN(n13404) );
  NOR2X0 U13726 ( .IN1(n9992), .IN2(n11182), .QN(n13403) );
  NAND2X0 U13727 ( .IN1(n10211), .IN2(n8459), .QN(n11182) );
  NAND2X0 U13728 ( .IN1(n13405), .IN2(n13406), .QN(WX7129) );
  NOR2X0 U13729 ( .IN1(n13407), .IN2(n13408), .QN(n13406) );
  NOR2X0 U13730 ( .IN1(n9942), .IN2(n13409), .QN(n13408) );
  NOR2X0 U13731 ( .IN1(n12585), .IN2(n9912), .QN(n13407) );
  NOR2X0 U13732 ( .IN1(n13410), .IN2(n13411), .QN(n12585) );
  INVX0 U13733 ( .INP(n13412), .ZN(n13411) );
  NAND2X0 U13734 ( .IN1(n13413), .IN2(n13414), .QN(n13412) );
  NOR2X0 U13735 ( .IN1(n13414), .IN2(n13413), .QN(n13410) );
  NAND2X0 U13736 ( .IN1(n13415), .IN2(n13416), .QN(n13413) );
  NAND2X0 U13737 ( .IN1(n9086), .IN2(n13417), .QN(n13416) );
  INVX0 U13738 ( .INP(n13418), .ZN(n13415) );
  NOR2X0 U13739 ( .IN1(n13417), .IN2(n9086), .QN(n13418) );
  NOR2X0 U13740 ( .IN1(n13419), .IN2(n13420), .QN(n13417) );
  INVX0 U13741 ( .INP(n13421), .ZN(n13420) );
  NAND2X0 U13742 ( .IN1(n18437), .IN2(WX8615), .QN(n13421) );
  NOR2X0 U13743 ( .IN1(WX8615), .IN2(n18437), .QN(n13419) );
  NOR2X0 U13744 ( .IN1(n13422), .IN2(n13423), .QN(n13414) );
  INVX0 U13745 ( .INP(n13424), .ZN(n13423) );
  NAND2X0 U13746 ( .IN1(n9085), .IN2(n10014), .QN(n13424) );
  NOR2X0 U13747 ( .IN1(n10006), .IN2(n9085), .QN(n13422) );
  NOR2X0 U13748 ( .IN1(n13425), .IN2(n13426), .QN(n13405) );
  NOR2X0 U13749 ( .IN1(DFF_1141_n1), .IN2(n9960), .QN(n13426) );
  NOR2X0 U13750 ( .IN1(n9992), .IN2(n11183), .QN(n13425) );
  NAND2X0 U13751 ( .IN1(n10211), .IN2(n8460), .QN(n11183) );
  NAND2X0 U13752 ( .IN1(n13427), .IN2(n13428), .QN(WX7127) );
  NOR2X0 U13753 ( .IN1(n13429), .IN2(n13430), .QN(n13428) );
  NOR2X0 U13754 ( .IN1(n13431), .IN2(n9933), .QN(n13430) );
  NOR2X0 U13755 ( .IN1(n12607), .IN2(n9912), .QN(n13429) );
  NOR2X0 U13756 ( .IN1(n13432), .IN2(n13433), .QN(n12607) );
  INVX0 U13757 ( .INP(n13434), .ZN(n13433) );
  NAND2X0 U13758 ( .IN1(n13435), .IN2(n13436), .QN(n13434) );
  NOR2X0 U13759 ( .IN1(n13436), .IN2(n13435), .QN(n13432) );
  NAND2X0 U13760 ( .IN1(n13437), .IN2(n13438), .QN(n13435) );
  NAND2X0 U13761 ( .IN1(n9088), .IN2(n13439), .QN(n13438) );
  INVX0 U13762 ( .INP(n13440), .ZN(n13437) );
  NOR2X0 U13763 ( .IN1(n13439), .IN2(n9088), .QN(n13440) );
  NOR2X0 U13764 ( .IN1(n13441), .IN2(n13442), .QN(n13439) );
  INVX0 U13765 ( .INP(n13443), .ZN(n13442) );
  NAND2X0 U13766 ( .IN1(n18436), .IN2(WX8613), .QN(n13443) );
  NOR2X0 U13767 ( .IN1(WX8613), .IN2(n18436), .QN(n13441) );
  NOR2X0 U13768 ( .IN1(n13444), .IN2(n13445), .QN(n13436) );
  INVX0 U13769 ( .INP(n13446), .ZN(n13445) );
  NAND2X0 U13770 ( .IN1(n9087), .IN2(n10014), .QN(n13446) );
  NOR2X0 U13771 ( .IN1(n10006), .IN2(n9087), .QN(n13444) );
  NOR2X0 U13772 ( .IN1(n13447), .IN2(n13448), .QN(n13427) );
  NOR2X0 U13773 ( .IN1(DFF_1142_n1), .IN2(n9960), .QN(n13448) );
  NOR2X0 U13774 ( .IN1(n9992), .IN2(n11184), .QN(n13447) );
  NAND2X0 U13775 ( .IN1(n10211), .IN2(n8461), .QN(n11184) );
  NAND2X0 U13776 ( .IN1(n13449), .IN2(n13450), .QN(WX7125) );
  NOR2X0 U13777 ( .IN1(n13451), .IN2(n13452), .QN(n13450) );
  NOR2X0 U13778 ( .IN1(n9942), .IN2(n13453), .QN(n13452) );
  NOR2X0 U13779 ( .IN1(n12629), .IN2(n9912), .QN(n13451) );
  NOR2X0 U13780 ( .IN1(n13454), .IN2(n13455), .QN(n12629) );
  INVX0 U13781 ( .INP(n13456), .ZN(n13455) );
  NAND2X0 U13782 ( .IN1(n13457), .IN2(n13458), .QN(n13456) );
  NOR2X0 U13783 ( .IN1(n13458), .IN2(n13457), .QN(n13454) );
  NAND2X0 U13784 ( .IN1(n13459), .IN2(n13460), .QN(n13457) );
  NAND2X0 U13785 ( .IN1(n9090), .IN2(n13461), .QN(n13460) );
  INVX0 U13786 ( .INP(n13462), .ZN(n13459) );
  NOR2X0 U13787 ( .IN1(n13461), .IN2(n9090), .QN(n13462) );
  NOR2X0 U13788 ( .IN1(n13463), .IN2(n13464), .QN(n13461) );
  INVX0 U13789 ( .INP(n13465), .ZN(n13464) );
  NAND2X0 U13790 ( .IN1(n18435), .IN2(WX8611), .QN(n13465) );
  NOR2X0 U13791 ( .IN1(WX8611), .IN2(n18435), .QN(n13463) );
  NOR2X0 U13792 ( .IN1(n13466), .IN2(n13467), .QN(n13458) );
  INVX0 U13793 ( .INP(n13468), .ZN(n13467) );
  NAND2X0 U13794 ( .IN1(n9089), .IN2(n10013), .QN(n13468) );
  NOR2X0 U13795 ( .IN1(n10006), .IN2(n9089), .QN(n13466) );
  NOR2X0 U13796 ( .IN1(n13469), .IN2(n13470), .QN(n13449) );
  NOR2X0 U13797 ( .IN1(DFF_1143_n1), .IN2(n9960), .QN(n13470) );
  NOR2X0 U13798 ( .IN1(n9991), .IN2(n11185), .QN(n13469) );
  NAND2X0 U13799 ( .IN1(n10212), .IN2(n8462), .QN(n11185) );
  NAND2X0 U13800 ( .IN1(n13471), .IN2(n13472), .QN(WX7123) );
  NOR2X0 U13801 ( .IN1(n13473), .IN2(n13474), .QN(n13472) );
  NOR2X0 U13802 ( .IN1(n13475), .IN2(n9933), .QN(n13474) );
  NOR2X0 U13803 ( .IN1(n12651), .IN2(n9912), .QN(n13473) );
  NOR2X0 U13804 ( .IN1(n13476), .IN2(n13477), .QN(n12651) );
  INVX0 U13805 ( .INP(n13478), .ZN(n13477) );
  NAND2X0 U13806 ( .IN1(n13479), .IN2(n13480), .QN(n13478) );
  NOR2X0 U13807 ( .IN1(n13480), .IN2(n13479), .QN(n13476) );
  NAND2X0 U13808 ( .IN1(n13481), .IN2(n13482), .QN(n13479) );
  NAND2X0 U13809 ( .IN1(n9092), .IN2(n13483), .QN(n13482) );
  INVX0 U13810 ( .INP(n13484), .ZN(n13481) );
  NOR2X0 U13811 ( .IN1(n13483), .IN2(n9092), .QN(n13484) );
  NOR2X0 U13812 ( .IN1(n13485), .IN2(n13486), .QN(n13483) );
  INVX0 U13813 ( .INP(n13487), .ZN(n13486) );
  NAND2X0 U13814 ( .IN1(n18434), .IN2(WX8609), .QN(n13487) );
  NOR2X0 U13815 ( .IN1(WX8609), .IN2(n18434), .QN(n13485) );
  NOR2X0 U13816 ( .IN1(n13488), .IN2(n13489), .QN(n13480) );
  INVX0 U13817 ( .INP(n13490), .ZN(n13489) );
  NAND2X0 U13818 ( .IN1(n9091), .IN2(n10013), .QN(n13490) );
  NOR2X0 U13819 ( .IN1(n10006), .IN2(n9091), .QN(n13488) );
  NOR2X0 U13820 ( .IN1(n13491), .IN2(n13492), .QN(n13471) );
  NOR2X0 U13821 ( .IN1(DFF_1144_n1), .IN2(n9960), .QN(n13492) );
  NOR2X0 U13822 ( .IN1(n9991), .IN2(n11186), .QN(n13491) );
  NAND2X0 U13823 ( .IN1(n10211), .IN2(n8463), .QN(n11186) );
  NAND2X0 U13824 ( .IN1(n13493), .IN2(n13494), .QN(WX7121) );
  NOR2X0 U13825 ( .IN1(n13495), .IN2(n13496), .QN(n13494) );
  NOR2X0 U13826 ( .IN1(n9942), .IN2(n13497), .QN(n13496) );
  NOR2X0 U13827 ( .IN1(n12673), .IN2(n9912), .QN(n13495) );
  NOR2X0 U13828 ( .IN1(n13498), .IN2(n13499), .QN(n12673) );
  INVX0 U13829 ( .INP(n13500), .ZN(n13499) );
  NAND2X0 U13830 ( .IN1(n13501), .IN2(n13502), .QN(n13500) );
  NOR2X0 U13831 ( .IN1(n13502), .IN2(n13501), .QN(n13498) );
  NAND2X0 U13832 ( .IN1(n13503), .IN2(n13504), .QN(n13501) );
  NAND2X0 U13833 ( .IN1(n9094), .IN2(n13505), .QN(n13504) );
  INVX0 U13834 ( .INP(n13506), .ZN(n13503) );
  NOR2X0 U13835 ( .IN1(n13505), .IN2(n9094), .QN(n13506) );
  NOR2X0 U13836 ( .IN1(n13507), .IN2(n13508), .QN(n13505) );
  INVX0 U13837 ( .INP(n13509), .ZN(n13508) );
  NAND2X0 U13838 ( .IN1(n18433), .IN2(WX8607), .QN(n13509) );
  NOR2X0 U13839 ( .IN1(WX8607), .IN2(n18433), .QN(n13507) );
  NOR2X0 U13840 ( .IN1(n13510), .IN2(n13511), .QN(n13502) );
  INVX0 U13841 ( .INP(n13512), .ZN(n13511) );
  NAND2X0 U13842 ( .IN1(n9093), .IN2(n10013), .QN(n13512) );
  NOR2X0 U13843 ( .IN1(n10006), .IN2(n9093), .QN(n13510) );
  NOR2X0 U13844 ( .IN1(n13513), .IN2(n13514), .QN(n13493) );
  NOR2X0 U13845 ( .IN1(DFF_1145_n1), .IN2(n9959), .QN(n13514) );
  NOR2X0 U13846 ( .IN1(n9991), .IN2(n11187), .QN(n13513) );
  NAND2X0 U13847 ( .IN1(n10211), .IN2(n8464), .QN(n11187) );
  NAND2X0 U13848 ( .IN1(n13515), .IN2(n13516), .QN(WX7119) );
  NOR2X0 U13849 ( .IN1(n13517), .IN2(n13518), .QN(n13516) );
  NOR2X0 U13850 ( .IN1(n13519), .IN2(n9933), .QN(n13518) );
  NOR2X0 U13851 ( .IN1(n9921), .IN2(n12695), .QN(n13517) );
  NAND2X0 U13852 ( .IN1(n13520), .IN2(n13521), .QN(n12695) );
  NAND2X0 U13853 ( .IN1(n13522), .IN2(n13523), .QN(n13521) );
  INVX0 U13854 ( .INP(n13524), .ZN(n13520) );
  NOR2X0 U13855 ( .IN1(n13523), .IN2(n13522), .QN(n13524) );
  NAND2X0 U13856 ( .IN1(n13525), .IN2(n13526), .QN(n13522) );
  NAND2X0 U13857 ( .IN1(n13527), .IN2(WX8541), .QN(n13526) );
  NAND2X0 U13858 ( .IN1(n13528), .IN2(n13529), .QN(n13527) );
  NAND2X0 U13859 ( .IN1(test_so74), .IN2(WX8477), .QN(n13529) );
  NAND2X0 U13860 ( .IN1(n9095), .IN2(n9828), .QN(n13528) );
  NAND2X0 U13861 ( .IN1(n9096), .IN2(n13530), .QN(n13525) );
  NOR2X0 U13862 ( .IN1(n13531), .IN2(n13532), .QN(n13530) );
  NOR2X0 U13863 ( .IN1(test_so74), .IN2(WX8477), .QN(n13532) );
  NOR2X0 U13864 ( .IN1(n9095), .IN2(n9828), .QN(n13531) );
  NOR2X0 U13865 ( .IN1(n13533), .IN2(n13534), .QN(n13523) );
  INVX0 U13866 ( .INP(n13535), .ZN(n13534) );
  NAND2X0 U13867 ( .IN1(n18432), .IN2(n10017), .QN(n13535) );
  NOR2X0 U13868 ( .IN1(n10006), .IN2(n18432), .QN(n13533) );
  NOR2X0 U13869 ( .IN1(n13536), .IN2(n13537), .QN(n13515) );
  NOR2X0 U13870 ( .IN1(DFF_1146_n1), .IN2(n9959), .QN(n13537) );
  NOR2X0 U13871 ( .IN1(n9991), .IN2(n11188), .QN(n13536) );
  NAND2X0 U13872 ( .IN1(n10209), .IN2(n8465), .QN(n11188) );
  NAND2X0 U13873 ( .IN1(n13538), .IN2(n13539), .QN(WX7117) );
  NOR2X0 U13874 ( .IN1(n13540), .IN2(n13541), .QN(n13539) );
  NOR2X0 U13875 ( .IN1(n9942), .IN2(n13542), .QN(n13541) );
  NOR2X0 U13876 ( .IN1(n12717), .IN2(n9912), .QN(n13540) );
  NOR2X0 U13877 ( .IN1(n13543), .IN2(n13544), .QN(n12717) );
  INVX0 U13878 ( .INP(n13545), .ZN(n13544) );
  NAND2X0 U13879 ( .IN1(n13546), .IN2(n13547), .QN(n13545) );
  NOR2X0 U13880 ( .IN1(n13547), .IN2(n13546), .QN(n13543) );
  NAND2X0 U13881 ( .IN1(n13548), .IN2(n13549), .QN(n13546) );
  NAND2X0 U13882 ( .IN1(n9098), .IN2(n13550), .QN(n13549) );
  INVX0 U13883 ( .INP(n13551), .ZN(n13548) );
  NOR2X0 U13884 ( .IN1(n13550), .IN2(n9098), .QN(n13551) );
  NOR2X0 U13885 ( .IN1(n13552), .IN2(n13553), .QN(n13550) );
  INVX0 U13886 ( .INP(n13554), .ZN(n13553) );
  NAND2X0 U13887 ( .IN1(n18431), .IN2(WX8603), .QN(n13554) );
  NOR2X0 U13888 ( .IN1(WX8603), .IN2(n18431), .QN(n13552) );
  NOR2X0 U13889 ( .IN1(n13555), .IN2(n13556), .QN(n13547) );
  INVX0 U13890 ( .INP(n13557), .ZN(n13556) );
  NAND2X0 U13891 ( .IN1(n9097), .IN2(n10017), .QN(n13557) );
  NOR2X0 U13892 ( .IN1(n10006), .IN2(n9097), .QN(n13555) );
  NOR2X0 U13893 ( .IN1(n13558), .IN2(n13559), .QN(n13538) );
  NOR2X0 U13894 ( .IN1(DFF_1147_n1), .IN2(n9959), .QN(n13559) );
  NOR2X0 U13895 ( .IN1(n9991), .IN2(n11189), .QN(n13558) );
  NAND2X0 U13896 ( .IN1(n10210), .IN2(n8466), .QN(n11189) );
  NAND2X0 U13897 ( .IN1(n13560), .IN2(n13561), .QN(WX7115) );
  NOR2X0 U13898 ( .IN1(n13562), .IN2(n13563), .QN(n13561) );
  NOR2X0 U13899 ( .IN1(n13564), .IN2(n9933), .QN(n13563) );
  NOR2X0 U13900 ( .IN1(n9922), .IN2(n12739), .QN(n13562) );
  NAND2X0 U13901 ( .IN1(n13565), .IN2(n13566), .QN(n12739) );
  INVX0 U13902 ( .INP(n13567), .ZN(n13566) );
  NOR2X0 U13903 ( .IN1(n13568), .IN2(n13569), .QN(n13567) );
  NAND2X0 U13904 ( .IN1(n13569), .IN2(n13568), .QN(n13565) );
  NOR2X0 U13905 ( .IN1(n13570), .IN2(n13571), .QN(n13568) );
  INVX0 U13906 ( .INP(n13572), .ZN(n13571) );
  NAND2X0 U13907 ( .IN1(n9580), .IN2(n13573), .QN(n13572) );
  NOR2X0 U13908 ( .IN1(n13573), .IN2(n9580), .QN(n13570) );
  NOR2X0 U13909 ( .IN1(n13574), .IN2(n13575), .QN(n13573) );
  INVX0 U13910 ( .INP(n13576), .ZN(n13575) );
  NAND2X0 U13911 ( .IN1(test_so72), .IN2(n8375), .QN(n13576) );
  NOR2X0 U13912 ( .IN1(n8375), .IN2(test_so72), .QN(n13574) );
  NAND2X0 U13913 ( .IN1(n13577), .IN2(n13578), .QN(n13569) );
  NAND2X0 U13914 ( .IN1(n9099), .IN2(n10017), .QN(n13578) );
  INVX0 U13915 ( .INP(n13579), .ZN(n13577) );
  NOR2X0 U13916 ( .IN1(n10006), .IN2(n9099), .QN(n13579) );
  NOR2X0 U13917 ( .IN1(n13580), .IN2(n13581), .QN(n13560) );
  NOR2X0 U13918 ( .IN1(DFF_1148_n1), .IN2(n9959), .QN(n13581) );
  NOR2X0 U13919 ( .IN1(n9991), .IN2(n11190), .QN(n13580) );
  NAND2X0 U13920 ( .IN1(n10211), .IN2(n8467), .QN(n11190) );
  NAND2X0 U13921 ( .IN1(n13582), .IN2(n13583), .QN(WX7113) );
  NOR2X0 U13922 ( .IN1(n13584), .IN2(n13585), .QN(n13583) );
  NOR2X0 U13923 ( .IN1(n13586), .IN2(n9933), .QN(n13585) );
  NOR2X0 U13924 ( .IN1(n12761), .IN2(n9913), .QN(n13584) );
  NOR2X0 U13925 ( .IN1(n13587), .IN2(n13588), .QN(n12761) );
  INVX0 U13926 ( .INP(n13589), .ZN(n13588) );
  NAND2X0 U13927 ( .IN1(n13590), .IN2(n13591), .QN(n13589) );
  NOR2X0 U13928 ( .IN1(n13591), .IN2(n13590), .QN(n13587) );
  NAND2X0 U13929 ( .IN1(n13592), .IN2(n13593), .QN(n13590) );
  NAND2X0 U13930 ( .IN1(n9101), .IN2(n13594), .QN(n13593) );
  INVX0 U13931 ( .INP(n13595), .ZN(n13592) );
  NOR2X0 U13932 ( .IN1(n13594), .IN2(n9101), .QN(n13595) );
  NOR2X0 U13933 ( .IN1(n13596), .IN2(n13597), .QN(n13594) );
  INVX0 U13934 ( .INP(n13598), .ZN(n13597) );
  NAND2X0 U13935 ( .IN1(n18429), .IN2(WX8599), .QN(n13598) );
  NOR2X0 U13936 ( .IN1(WX8599), .IN2(n18429), .QN(n13596) );
  NOR2X0 U13937 ( .IN1(n13599), .IN2(n13600), .QN(n13591) );
  INVX0 U13938 ( .INP(n13601), .ZN(n13600) );
  NAND2X0 U13939 ( .IN1(n9100), .IN2(n10017), .QN(n13601) );
  NOR2X0 U13940 ( .IN1(n10006), .IN2(n9100), .QN(n13599) );
  NOR2X0 U13941 ( .IN1(n13602), .IN2(n13603), .QN(n13582) );
  NOR2X0 U13942 ( .IN1(n9976), .IN2(n9855), .QN(n13603) );
  NOR2X0 U13943 ( .IN1(n9991), .IN2(n11191), .QN(n13602) );
  NAND2X0 U13944 ( .IN1(test_so55), .IN2(n10214), .QN(n11191) );
  NAND2X0 U13945 ( .IN1(n13604), .IN2(n13605), .QN(WX7111) );
  NOR2X0 U13946 ( .IN1(n13606), .IN2(n13607), .QN(n13605) );
  NOR2X0 U13947 ( .IN1(n13608), .IN2(n9933), .QN(n13607) );
  NOR2X0 U13948 ( .IN1(n9922), .IN2(n12783), .QN(n13606) );
  NAND2X0 U13949 ( .IN1(n13609), .IN2(n13610), .QN(n12783) );
  INVX0 U13950 ( .INP(n13611), .ZN(n13610) );
  NOR2X0 U13951 ( .IN1(n13612), .IN2(n13613), .QN(n13611) );
  NAND2X0 U13952 ( .IN1(n13613), .IN2(n13612), .QN(n13609) );
  NOR2X0 U13953 ( .IN1(n13614), .IN2(n13615), .QN(n13612) );
  INVX0 U13954 ( .INP(n13616), .ZN(n13615) );
  NAND2X0 U13955 ( .IN1(n9578), .IN2(n13617), .QN(n13616) );
  NOR2X0 U13956 ( .IN1(n13617), .IN2(n9578), .QN(n13614) );
  NOR2X0 U13957 ( .IN1(n13618), .IN2(n13619), .QN(n13617) );
  INVX0 U13958 ( .INP(n13620), .ZN(n13619) );
  NAND2X0 U13959 ( .IN1(test_so70), .IN2(n8377), .QN(n13620) );
  NOR2X0 U13960 ( .IN1(n8377), .IN2(test_so70), .QN(n13618) );
  NAND2X0 U13961 ( .IN1(n13621), .IN2(n13622), .QN(n13613) );
  NAND2X0 U13962 ( .IN1(n9102), .IN2(n10017), .QN(n13622) );
  INVX0 U13963 ( .INP(n13623), .ZN(n13621) );
  NOR2X0 U13964 ( .IN1(n10006), .IN2(n9102), .QN(n13623) );
  NOR2X0 U13965 ( .IN1(n13624), .IN2(n13625), .QN(n13604) );
  NOR2X0 U13966 ( .IN1(DFF_1150_n1), .IN2(n9959), .QN(n13625) );
  NOR2X0 U13967 ( .IN1(n9991), .IN2(n11192), .QN(n13624) );
  NAND2X0 U13968 ( .IN1(n10211), .IN2(n8470), .QN(n11192) );
  NAND2X0 U13969 ( .IN1(n13626), .IN2(n13627), .QN(WX7109) );
  NOR2X0 U13970 ( .IN1(n13628), .IN2(n13629), .QN(n13627) );
  NOR2X0 U13971 ( .IN1(n13630), .IN2(n9933), .QN(n13629) );
  NOR2X0 U13972 ( .IN1(n12805), .IN2(n9913), .QN(n13628) );
  NOR2X0 U13973 ( .IN1(n13631), .IN2(n13632), .QN(n12805) );
  INVX0 U13974 ( .INP(n13633), .ZN(n13632) );
  NAND2X0 U13975 ( .IN1(n13634), .IN2(n13635), .QN(n13633) );
  NOR2X0 U13976 ( .IN1(n13635), .IN2(n13634), .QN(n13631) );
  NAND2X0 U13977 ( .IN1(n13636), .IN2(n13637), .QN(n13634) );
  NAND2X0 U13978 ( .IN1(n9008), .IN2(n13638), .QN(n13637) );
  INVX0 U13979 ( .INP(n13639), .ZN(n13636) );
  NOR2X0 U13980 ( .IN1(n13638), .IN2(n9008), .QN(n13639) );
  NOR2X0 U13981 ( .IN1(n13640), .IN2(n13641), .QN(n13638) );
  INVX0 U13982 ( .INP(n13642), .ZN(n13641) );
  NAND2X0 U13983 ( .IN1(n18427), .IN2(WX8595), .QN(n13642) );
  NOR2X0 U13984 ( .IN1(WX8595), .IN2(n18427), .QN(n13640) );
  NOR2X0 U13985 ( .IN1(n13643), .IN2(n13644), .QN(n13635) );
  INVX0 U13986 ( .INP(n13645), .ZN(n13644) );
  NAND2X0 U13987 ( .IN1(n9007), .IN2(n10017), .QN(n13645) );
  NOR2X0 U13988 ( .IN1(n10006), .IN2(n9007), .QN(n13643) );
  NOR2X0 U13989 ( .IN1(n13646), .IN2(n13647), .QN(n13626) );
  NOR2X0 U13990 ( .IN1(n9491), .IN2(n11994), .QN(n13647) );
  NOR2X0 U13991 ( .IN1(DFF_1151_n1), .IN2(n9959), .QN(n13646) );
  INVX0 U13992 ( .INP(n13648), .ZN(WX7011) );
  NAND2X0 U13993 ( .IN1(n10211), .IN2(n9491), .QN(n13648) );
  NOR2X0 U13994 ( .IN1(n10326), .IN2(n13649), .QN(WX6498) );
  NAND2X0 U13995 ( .IN1(n13650), .IN2(n13651), .QN(n13649) );
  INVX0 U13996 ( .INP(n13652), .ZN(n13651) );
  NOR2X0 U13997 ( .IN1(WX6009), .IN2(DFF_958_n1), .QN(n13652) );
  NAND2X0 U13998 ( .IN1(DFF_958_n1), .IN2(WX6009), .QN(n13650) );
  NOR2X0 U13999 ( .IN1(n10326), .IN2(n13653), .QN(WX6496) );
  NAND2X0 U14000 ( .IN1(n13654), .IN2(n13655), .QN(n13653) );
  INVX0 U14001 ( .INP(n13656), .ZN(n13655) );
  NOR2X0 U14002 ( .IN1(WX6011), .IN2(DFF_957_n1), .QN(n13656) );
  NAND2X0 U14003 ( .IN1(DFF_957_n1), .IN2(WX6011), .QN(n13654) );
  NOR2X0 U14004 ( .IN1(n10326), .IN2(n13657), .QN(WX6494) );
  NAND2X0 U14005 ( .IN1(n13658), .IN2(n13659), .QN(n13657) );
  INVX0 U14006 ( .INP(n13660), .ZN(n13659) );
  NOR2X0 U14007 ( .IN1(WX6013), .IN2(DFF_956_n1), .QN(n13660) );
  NAND2X0 U14008 ( .IN1(DFF_956_n1), .IN2(WX6013), .QN(n13658) );
  NOR2X0 U14009 ( .IN1(n10326), .IN2(n13661), .QN(WX6492) );
  NAND2X0 U14010 ( .IN1(n13662), .IN2(n13663), .QN(n13661) );
  INVX0 U14011 ( .INP(n13664), .ZN(n13663) );
  NOR2X0 U14012 ( .IN1(WX6015), .IN2(DFF_955_n1), .QN(n13664) );
  NAND2X0 U14013 ( .IN1(DFF_955_n1), .IN2(WX6015), .QN(n13662) );
  NOR2X0 U14014 ( .IN1(n10326), .IN2(n13665), .QN(WX6490) );
  NAND2X0 U14015 ( .IN1(n13666), .IN2(n13667), .QN(n13665) );
  INVX0 U14016 ( .INP(n13668), .ZN(n13667) );
  NOR2X0 U14017 ( .IN1(WX6017), .IN2(DFF_954_n1), .QN(n13668) );
  NAND2X0 U14018 ( .IN1(DFF_954_n1), .IN2(WX6017), .QN(n13666) );
  NOR2X0 U14019 ( .IN1(n10326), .IN2(n13669), .QN(WX6488) );
  NAND2X0 U14020 ( .IN1(n13670), .IN2(n13671), .QN(n13669) );
  INVX0 U14021 ( .INP(n13672), .ZN(n13671) );
  NOR2X0 U14022 ( .IN1(WX6019), .IN2(DFF_953_n1), .QN(n13672) );
  NAND2X0 U14023 ( .IN1(DFF_953_n1), .IN2(WX6019), .QN(n13670) );
  NOR2X0 U14024 ( .IN1(n10326), .IN2(n13673), .QN(WX6486) );
  NAND2X0 U14025 ( .IN1(n13674), .IN2(n13675), .QN(n13673) );
  INVX0 U14026 ( .INP(n13676), .ZN(n13675) );
  NOR2X0 U14027 ( .IN1(WX6021), .IN2(DFF_952_n1), .QN(n13676) );
  NAND2X0 U14028 ( .IN1(DFF_952_n1), .IN2(WX6021), .QN(n13674) );
  NOR2X0 U14029 ( .IN1(n10326), .IN2(n13677), .QN(WX6484) );
  NAND2X0 U14030 ( .IN1(n13678), .IN2(n13679), .QN(n13677) );
  INVX0 U14031 ( .INP(n13680), .ZN(n13679) );
  NOR2X0 U14032 ( .IN1(WX6023), .IN2(DFF_951_n1), .QN(n13680) );
  NAND2X0 U14033 ( .IN1(DFF_951_n1), .IN2(WX6023), .QN(n13678) );
  NOR2X0 U14034 ( .IN1(n10327), .IN2(n13681), .QN(WX6482) );
  NAND2X0 U14035 ( .IN1(n13682), .IN2(n13683), .QN(n13681) );
  INVX0 U14036 ( .INP(n13684), .ZN(n13683) );
  NOR2X0 U14037 ( .IN1(WX6025), .IN2(DFF_950_n1), .QN(n13684) );
  NAND2X0 U14038 ( .IN1(DFF_950_n1), .IN2(WX6025), .QN(n13682) );
  NOR2X0 U14039 ( .IN1(n10327), .IN2(n13685), .QN(WX6480) );
  NAND2X0 U14040 ( .IN1(n13686), .IN2(n13687), .QN(n13685) );
  INVX0 U14041 ( .INP(n13688), .ZN(n13687) );
  NOR2X0 U14042 ( .IN1(WX6027), .IN2(DFF_949_n1), .QN(n13688) );
  NAND2X0 U14043 ( .IN1(DFF_949_n1), .IN2(WX6027), .QN(n13686) );
  NOR2X0 U14044 ( .IN1(n10327), .IN2(n13689), .QN(WX6478) );
  NAND2X0 U14045 ( .IN1(n13690), .IN2(n13691), .QN(n13689) );
  INVX0 U14046 ( .INP(n13692), .ZN(n13691) );
  NOR2X0 U14047 ( .IN1(WX6029), .IN2(DFF_948_n1), .QN(n13692) );
  NAND2X0 U14048 ( .IN1(DFF_948_n1), .IN2(WX6029), .QN(n13690) );
  NOR2X0 U14049 ( .IN1(n10327), .IN2(n13693), .QN(WX6476) );
  NAND2X0 U14050 ( .IN1(n13694), .IN2(n13695), .QN(n13693) );
  INVX0 U14051 ( .INP(n13696), .ZN(n13695) );
  NOR2X0 U14052 ( .IN1(WX6031), .IN2(DFF_947_n1), .QN(n13696) );
  NAND2X0 U14053 ( .IN1(DFF_947_n1), .IN2(WX6031), .QN(n13694) );
  NOR2X0 U14054 ( .IN1(n10327), .IN2(n13697), .QN(WX6474) );
  NAND2X0 U14055 ( .IN1(n13698), .IN2(n13699), .QN(n13697) );
  INVX0 U14056 ( .INP(n13700), .ZN(n13699) );
  NOR2X0 U14057 ( .IN1(WX6033), .IN2(DFF_946_n1), .QN(n13700) );
  NAND2X0 U14058 ( .IN1(DFF_946_n1), .IN2(WX6033), .QN(n13698) );
  NOR2X0 U14059 ( .IN1(n10327), .IN2(n13701), .QN(WX6472) );
  NOR2X0 U14060 ( .IN1(n13702), .IN2(n13703), .QN(n13701) );
  NOR2X0 U14061 ( .IN1(test_so54), .IN2(WX6035), .QN(n13703) );
  NOR2X0 U14062 ( .IN1(n9643), .IN2(n9857), .QN(n13702) );
  NOR2X0 U14063 ( .IN1(n10327), .IN2(n13704), .QN(WX6470) );
  NAND2X0 U14064 ( .IN1(n13705), .IN2(n13706), .QN(n13704) );
  INVX0 U14065 ( .INP(n13707), .ZN(n13706) );
  NOR2X0 U14066 ( .IN1(WX6037), .IN2(DFF_944_n1), .QN(n13707) );
  NAND2X0 U14067 ( .IN1(DFF_944_n1), .IN2(WX6037), .QN(n13705) );
  NOR2X0 U14068 ( .IN1(n10327), .IN2(n13708), .QN(WX6468) );
  NAND2X0 U14069 ( .IN1(n13709), .IN2(n13710), .QN(n13708) );
  INVX0 U14070 ( .INP(n13711), .ZN(n13710) );
  NOR2X0 U14071 ( .IN1(CRC_OUT_5_15), .IN2(n13712), .QN(n13711) );
  NAND2X0 U14072 ( .IN1(n13712), .IN2(CRC_OUT_5_15), .QN(n13709) );
  NAND2X0 U14073 ( .IN1(n13713), .IN2(n13714), .QN(n13712) );
  NAND2X0 U14074 ( .IN1(test_so52), .IN2(CRC_OUT_5_31), .QN(n13714) );
  NAND2X0 U14075 ( .IN1(DFF_959_n1), .IN2(n9848), .QN(n13713) );
  NOR2X0 U14076 ( .IN1(n10327), .IN2(n13715), .QN(WX6466) );
  NAND2X0 U14077 ( .IN1(n13716), .IN2(n13717), .QN(n13715) );
  INVX0 U14078 ( .INP(n13718), .ZN(n13717) );
  NOR2X0 U14079 ( .IN1(WX6041), .IN2(DFF_942_n1), .QN(n13718) );
  NAND2X0 U14080 ( .IN1(DFF_942_n1), .IN2(WX6041), .QN(n13716) );
  NOR2X0 U14081 ( .IN1(n10327), .IN2(n13719), .QN(WX6464) );
  NAND2X0 U14082 ( .IN1(n13720), .IN2(n13721), .QN(n13719) );
  INVX0 U14083 ( .INP(n13722), .ZN(n13721) );
  NOR2X0 U14084 ( .IN1(WX6043), .IN2(DFF_941_n1), .QN(n13722) );
  NAND2X0 U14085 ( .IN1(DFF_941_n1), .IN2(WX6043), .QN(n13720) );
  NOR2X0 U14086 ( .IN1(n10327), .IN2(n13723), .QN(WX6462) );
  NAND2X0 U14087 ( .IN1(n13724), .IN2(n13725), .QN(n13723) );
  INVX0 U14088 ( .INP(n13726), .ZN(n13725) );
  NOR2X0 U14089 ( .IN1(WX6045), .IN2(DFF_940_n1), .QN(n13726) );
  NAND2X0 U14090 ( .IN1(DFF_940_n1), .IN2(WX6045), .QN(n13724) );
  NOR2X0 U14091 ( .IN1(n10327), .IN2(n13727), .QN(WX6460) );
  NAND2X0 U14092 ( .IN1(n13728), .IN2(n13729), .QN(n13727) );
  INVX0 U14093 ( .INP(n13730), .ZN(n13729) );
  NOR2X0 U14094 ( .IN1(WX6047), .IN2(DFF_939_n1), .QN(n13730) );
  NAND2X0 U14095 ( .IN1(DFF_939_n1), .IN2(WX6047), .QN(n13728) );
  NOR2X0 U14096 ( .IN1(n10327), .IN2(n13731), .QN(WX6458) );
  NOR2X0 U14097 ( .IN1(n13732), .IN2(n13733), .QN(n13731) );
  INVX0 U14098 ( .INP(n13734), .ZN(n13733) );
  NAND2X0 U14099 ( .IN1(CRC_OUT_5_10), .IN2(n13735), .QN(n13734) );
  NOR2X0 U14100 ( .IN1(n13735), .IN2(CRC_OUT_5_10), .QN(n13732) );
  NAND2X0 U14101 ( .IN1(n13736), .IN2(n13737), .QN(n13735) );
  NAND2X0 U14102 ( .IN1(n9507), .IN2(CRC_OUT_5_31), .QN(n13737) );
  NAND2X0 U14103 ( .IN1(DFF_959_n1), .IN2(WX6049), .QN(n13736) );
  NOR2X0 U14104 ( .IN1(n10328), .IN2(n13738), .QN(WX6456) );
  NAND2X0 U14105 ( .IN1(n13739), .IN2(n13740), .QN(n13738) );
  INVX0 U14106 ( .INP(n13741), .ZN(n13740) );
  NOR2X0 U14107 ( .IN1(WX6051), .IN2(DFF_937_n1), .QN(n13741) );
  NAND2X0 U14108 ( .IN1(DFF_937_n1), .IN2(WX6051), .QN(n13739) );
  NOR2X0 U14109 ( .IN1(n10328), .IN2(n13742), .QN(WX6454) );
  NAND2X0 U14110 ( .IN1(n13743), .IN2(n13744), .QN(n13742) );
  INVX0 U14111 ( .INP(n13745), .ZN(n13744) );
  NOR2X0 U14112 ( .IN1(WX6053), .IN2(DFF_936_n1), .QN(n13745) );
  NAND2X0 U14113 ( .IN1(DFF_936_n1), .IN2(WX6053), .QN(n13743) );
  NOR2X0 U14114 ( .IN1(n10328), .IN2(n13746), .QN(WX6452) );
  NAND2X0 U14115 ( .IN1(n13747), .IN2(n13748), .QN(n13746) );
  INVX0 U14116 ( .INP(n13749), .ZN(n13748) );
  NOR2X0 U14117 ( .IN1(WX6055), .IN2(DFF_935_n1), .QN(n13749) );
  NAND2X0 U14118 ( .IN1(DFF_935_n1), .IN2(WX6055), .QN(n13747) );
  NOR2X0 U14119 ( .IN1(n10328), .IN2(n13750), .QN(WX6450) );
  NAND2X0 U14120 ( .IN1(n13751), .IN2(n13752), .QN(n13750) );
  INVX0 U14121 ( .INP(n13753), .ZN(n13752) );
  NOR2X0 U14122 ( .IN1(WX6057), .IN2(DFF_934_n1), .QN(n13753) );
  NAND2X0 U14123 ( .IN1(DFF_934_n1), .IN2(WX6057), .QN(n13751) );
  NOR2X0 U14124 ( .IN1(n10328), .IN2(n13754), .QN(WX6448) );
  NAND2X0 U14125 ( .IN1(n13755), .IN2(n13756), .QN(n13754) );
  INVX0 U14126 ( .INP(n13757), .ZN(n13756) );
  NOR2X0 U14127 ( .IN1(WX6059), .IN2(DFF_933_n1), .QN(n13757) );
  NAND2X0 U14128 ( .IN1(DFF_933_n1), .IN2(WX6059), .QN(n13755) );
  NOR2X0 U14129 ( .IN1(n10328), .IN2(n13758), .QN(WX6446) );
  NAND2X0 U14130 ( .IN1(n13759), .IN2(n13760), .QN(n13758) );
  INVX0 U14131 ( .INP(n13761), .ZN(n13760) );
  NOR2X0 U14132 ( .IN1(WX6061), .IN2(DFF_932_n1), .QN(n13761) );
  NAND2X0 U14133 ( .IN1(DFF_932_n1), .IN2(WX6061), .QN(n13759) );
  NOR2X0 U14134 ( .IN1(n10328), .IN2(n13762), .QN(WX6444) );
  NOR2X0 U14135 ( .IN1(n13763), .IN2(n13764), .QN(n13762) );
  INVX0 U14136 ( .INP(n13765), .ZN(n13764) );
  NAND2X0 U14137 ( .IN1(CRC_OUT_5_3), .IN2(n13766), .QN(n13765) );
  NOR2X0 U14138 ( .IN1(n13766), .IN2(CRC_OUT_5_3), .QN(n13763) );
  NAND2X0 U14139 ( .IN1(n13767), .IN2(n13768), .QN(n13766) );
  NAND2X0 U14140 ( .IN1(n9508), .IN2(CRC_OUT_5_31), .QN(n13768) );
  NAND2X0 U14141 ( .IN1(DFF_959_n1), .IN2(WX6063), .QN(n13767) );
  NOR2X0 U14142 ( .IN1(n10328), .IN2(n13769), .QN(WX6442) );
  NAND2X0 U14143 ( .IN1(n13770), .IN2(n13771), .QN(n13769) );
  INVX0 U14144 ( .INP(n13772), .ZN(n13771) );
  NOR2X0 U14145 ( .IN1(WX6065), .IN2(DFF_930_n1), .QN(n13772) );
  NAND2X0 U14146 ( .IN1(DFF_930_n1), .IN2(WX6065), .QN(n13770) );
  NOR2X0 U14147 ( .IN1(n10328), .IN2(n13773), .QN(WX6440) );
  NAND2X0 U14148 ( .IN1(n13774), .IN2(n13775), .QN(n13773) );
  INVX0 U14149 ( .INP(n13776), .ZN(n13775) );
  NOR2X0 U14150 ( .IN1(WX6067), .IN2(DFF_929_n1), .QN(n13776) );
  NAND2X0 U14151 ( .IN1(DFF_929_n1), .IN2(WX6067), .QN(n13774) );
  NAND2X0 U14152 ( .IN1(n13777), .IN2(n13778), .QN(WX644) );
  NOR2X0 U14153 ( .IN1(n13779), .IN2(n13780), .QN(n13778) );
  NOR2X0 U14154 ( .IN1(n13781), .IN2(n9933), .QN(n13780) );
  NOR2X0 U14155 ( .IN1(n13782), .IN2(n9913), .QN(n13779) );
  NOR2X0 U14156 ( .IN1(n13783), .IN2(n13784), .QN(n13777) );
  NOR2X0 U14157 ( .IN1(n9487), .IN2(n11994), .QN(n13784) );
  NOR2X0 U14158 ( .IN1(DFF_191_n1), .IN2(n9959), .QN(n13783) );
  NOR2X0 U14159 ( .IN1(n10328), .IN2(n13785), .QN(WX6438) );
  NOR2X0 U14160 ( .IN1(n13786), .IN2(n13787), .QN(n13785) );
  NOR2X0 U14161 ( .IN1(test_so53), .IN2(WX6069), .QN(n13787) );
  NOR2X0 U14162 ( .IN1(n9657), .IN2(n9856), .QN(n13786) );
  NOR2X0 U14163 ( .IN1(n10328), .IN2(n13788), .QN(WX6436) );
  NAND2X0 U14164 ( .IN1(n13789), .IN2(n13790), .QN(n13788) );
  NAND2X0 U14165 ( .IN1(n9521), .IN2(CRC_OUT_5_31), .QN(n13790) );
  NAND2X0 U14166 ( .IN1(DFF_959_n1), .IN2(WX6071), .QN(n13789) );
  NOR2X0 U14167 ( .IN1(n18411), .IN2(n10238), .QN(WX5910) );
  NOR2X0 U14168 ( .IN1(n18410), .IN2(n10238), .QN(WX5908) );
  NOR2X0 U14169 ( .IN1(n18409), .IN2(n10238), .QN(WX5906) );
  NOR2X0 U14170 ( .IN1(n18408), .IN2(n10238), .QN(WX5904) );
  NOR2X0 U14171 ( .IN1(n18407), .IN2(n10238), .QN(WX5902) );
  NOR2X0 U14172 ( .IN1(n18406), .IN2(n10238), .QN(WX5900) );
  NOR2X0 U14173 ( .IN1(n10328), .IN2(n9842), .QN(WX5898) );
  NOR2X0 U14174 ( .IN1(n18405), .IN2(n10238), .QN(WX5896) );
  NOR2X0 U14175 ( .IN1(n18404), .IN2(n10238), .QN(WX5894) );
  NOR2X0 U14176 ( .IN1(n18403), .IN2(n10238), .QN(WX5892) );
  NOR2X0 U14177 ( .IN1(n18402), .IN2(n10238), .QN(WX5890) );
  NOR2X0 U14178 ( .IN1(n18401), .IN2(n10238), .QN(WX5888) );
  NOR2X0 U14179 ( .IN1(n18400), .IN2(n10239), .QN(WX5886) );
  NOR2X0 U14180 ( .IN1(n18399), .IN2(n10239), .QN(WX5884) );
  NOR2X0 U14181 ( .IN1(n18398), .IN2(n10294), .QN(WX5882) );
  NOR2X0 U14182 ( .IN1(n18397), .IN2(n10293), .QN(WX5880) );
  NAND2X0 U14183 ( .IN1(n13791), .IN2(n13792), .QN(WX5878) );
  NOR2X0 U14184 ( .IN1(n13793), .IN2(n13794), .QN(n13792) );
  NOR2X0 U14185 ( .IN1(n13795), .IN2(n9933), .QN(n13794) );
  NOR2X0 U14186 ( .IN1(n12963), .IN2(n9913), .QN(n13793) );
  INVX0 U14187 ( .INP(n13796), .ZN(n12963) );
  NAND2X0 U14188 ( .IN1(n13797), .IN2(n13798), .QN(n13796) );
  NAND2X0 U14189 ( .IN1(n13799), .IN2(n13800), .QN(n13798) );
  NAND2X0 U14190 ( .IN1(n13801), .IN2(n13802), .QN(n13800) );
  NAND2X0 U14191 ( .IN1(n9337), .IN2(WX7172), .QN(n13802) );
  NAND2X0 U14192 ( .IN1(n9336), .IN2(WX7300), .QN(n13801) );
  NOR2X0 U14193 ( .IN1(n13803), .IN2(n13804), .QN(n13799) );
  NOR2X0 U14194 ( .IN1(n9520), .IN2(WX7236), .QN(n13804) );
  NOR2X0 U14195 ( .IN1(n3627), .IN2(WX7364), .QN(n13803) );
  NAND2X0 U14196 ( .IN1(n13805), .IN2(n13806), .QN(n13797) );
  NAND2X0 U14197 ( .IN1(n13807), .IN2(n13808), .QN(n13806) );
  NAND2X0 U14198 ( .IN1(n9520), .IN2(WX7236), .QN(n13808) );
  NAND2X0 U14199 ( .IN1(n3627), .IN2(WX7364), .QN(n13807) );
  NOR2X0 U14200 ( .IN1(n13809), .IN2(n13810), .QN(n13805) );
  NOR2X0 U14201 ( .IN1(n9337), .IN2(WX7172), .QN(n13810) );
  NOR2X0 U14202 ( .IN1(n9336), .IN2(WX7300), .QN(n13809) );
  NOR2X0 U14203 ( .IN1(n13811), .IN2(n13812), .QN(n13791) );
  NOR2X0 U14204 ( .IN1(n9975), .IN2(n9856), .QN(n13812) );
  NOR2X0 U14205 ( .IN1(n9991), .IN2(n11274), .QN(n13811) );
  NAND2X0 U14206 ( .IN1(n10210), .IN2(n8496), .QN(n11274) );
  NAND2X0 U14207 ( .IN1(n13813), .IN2(n13814), .QN(WX5876) );
  NOR2X0 U14208 ( .IN1(n13815), .IN2(n13816), .QN(n13814) );
  NOR2X0 U14209 ( .IN1(n9943), .IN2(n13817), .QN(n13816) );
  NOR2X0 U14210 ( .IN1(n12985), .IN2(n9913), .QN(n13815) );
  INVX0 U14211 ( .INP(n13818), .ZN(n12985) );
  NAND2X0 U14212 ( .IN1(n13819), .IN2(n13820), .QN(n13818) );
  NAND2X0 U14213 ( .IN1(n13821), .IN2(n13822), .QN(n13820) );
  NAND2X0 U14214 ( .IN1(n13823), .IN2(n13824), .QN(n13822) );
  NAND2X0 U14215 ( .IN1(n9339), .IN2(WX7170), .QN(n13824) );
  NAND2X0 U14216 ( .IN1(n9338), .IN2(WX7298), .QN(n13823) );
  NOR2X0 U14217 ( .IN1(n13825), .IN2(n13826), .QN(n13821) );
  NOR2X0 U14218 ( .IN1(n9629), .IN2(WX7234), .QN(n13826) );
  NOR2X0 U14219 ( .IN1(n3629), .IN2(WX7362), .QN(n13825) );
  NAND2X0 U14220 ( .IN1(n13827), .IN2(n13828), .QN(n13819) );
  NAND2X0 U14221 ( .IN1(n13829), .IN2(n13830), .QN(n13828) );
  NAND2X0 U14222 ( .IN1(n9629), .IN2(WX7234), .QN(n13830) );
  NAND2X0 U14223 ( .IN1(n3629), .IN2(WX7362), .QN(n13829) );
  NOR2X0 U14224 ( .IN1(n13831), .IN2(n13832), .QN(n13827) );
  NOR2X0 U14225 ( .IN1(n9339), .IN2(WX7170), .QN(n13832) );
  NOR2X0 U14226 ( .IN1(n9338), .IN2(WX7298), .QN(n13831) );
  NOR2X0 U14227 ( .IN1(n13833), .IN2(n13834), .QN(n13813) );
  NOR2X0 U14228 ( .IN1(DFF_929_n1), .IN2(n9959), .QN(n13834) );
  NOR2X0 U14229 ( .IN1(n9991), .IN2(n11275), .QN(n13833) );
  NAND2X0 U14230 ( .IN1(n10210), .IN2(n8497), .QN(n11275) );
  NAND2X0 U14231 ( .IN1(n13835), .IN2(n13836), .QN(WX5874) );
  NOR2X0 U14232 ( .IN1(n13837), .IN2(n13838), .QN(n13836) );
  NOR2X0 U14233 ( .IN1(n13839), .IN2(n9933), .QN(n13838) );
  NOR2X0 U14234 ( .IN1(n13007), .IN2(n9913), .QN(n13837) );
  INVX0 U14235 ( .INP(n13840), .ZN(n13007) );
  NAND2X0 U14236 ( .IN1(n13841), .IN2(n13842), .QN(n13840) );
  NAND2X0 U14237 ( .IN1(n13843), .IN2(n13844), .QN(n13842) );
  NAND2X0 U14238 ( .IN1(n13845), .IN2(n13846), .QN(n13844) );
  NAND2X0 U14239 ( .IN1(n9341), .IN2(WX7168), .QN(n13846) );
  NAND2X0 U14240 ( .IN1(n9340), .IN2(WX7296), .QN(n13845) );
  NOR2X0 U14241 ( .IN1(n13847), .IN2(n13848), .QN(n13843) );
  NOR2X0 U14242 ( .IN1(n9628), .IN2(WX7232), .QN(n13848) );
  NOR2X0 U14243 ( .IN1(n3631), .IN2(WX7360), .QN(n13847) );
  NAND2X0 U14244 ( .IN1(n13849), .IN2(n13850), .QN(n13841) );
  NAND2X0 U14245 ( .IN1(n13851), .IN2(n13852), .QN(n13850) );
  NAND2X0 U14246 ( .IN1(n9628), .IN2(WX7232), .QN(n13852) );
  NAND2X0 U14247 ( .IN1(n3631), .IN2(WX7360), .QN(n13851) );
  NOR2X0 U14248 ( .IN1(n13853), .IN2(n13854), .QN(n13849) );
  NOR2X0 U14249 ( .IN1(n9341), .IN2(WX7168), .QN(n13854) );
  NOR2X0 U14250 ( .IN1(n9340), .IN2(WX7296), .QN(n13853) );
  NOR2X0 U14251 ( .IN1(n13855), .IN2(n13856), .QN(n13835) );
  NOR2X0 U14252 ( .IN1(DFF_930_n1), .IN2(n9959), .QN(n13856) );
  NOR2X0 U14253 ( .IN1(n9991), .IN2(n11276), .QN(n13855) );
  NAND2X0 U14254 ( .IN1(n10210), .IN2(n8498), .QN(n11276) );
  NAND2X0 U14255 ( .IN1(n13857), .IN2(n13858), .QN(WX5872) );
  NOR2X0 U14256 ( .IN1(n13859), .IN2(n13860), .QN(n13858) );
  NOR2X0 U14257 ( .IN1(n9943), .IN2(n13861), .QN(n13860) );
  NOR2X0 U14258 ( .IN1(n13029), .IN2(n9913), .QN(n13859) );
  INVX0 U14259 ( .INP(n13862), .ZN(n13029) );
  NAND2X0 U14260 ( .IN1(n13863), .IN2(n13864), .QN(n13862) );
  NAND2X0 U14261 ( .IN1(n13865), .IN2(n13866), .QN(n13864) );
  NAND2X0 U14262 ( .IN1(n13867), .IN2(n13868), .QN(n13866) );
  NAND2X0 U14263 ( .IN1(n9343), .IN2(WX7166), .QN(n13868) );
  NAND2X0 U14264 ( .IN1(n9342), .IN2(WX7294), .QN(n13867) );
  NOR2X0 U14265 ( .IN1(n13869), .IN2(n13870), .QN(n13865) );
  NOR2X0 U14266 ( .IN1(n9627), .IN2(WX7230), .QN(n13870) );
  NOR2X0 U14267 ( .IN1(n3633), .IN2(WX7358), .QN(n13869) );
  NAND2X0 U14268 ( .IN1(n13871), .IN2(n13872), .QN(n13863) );
  NAND2X0 U14269 ( .IN1(n13873), .IN2(n13874), .QN(n13872) );
  NAND2X0 U14270 ( .IN1(n9627), .IN2(WX7230), .QN(n13874) );
  NAND2X0 U14271 ( .IN1(n3633), .IN2(WX7358), .QN(n13873) );
  NOR2X0 U14272 ( .IN1(n13875), .IN2(n13876), .QN(n13871) );
  NOR2X0 U14273 ( .IN1(n9343), .IN2(WX7166), .QN(n13876) );
  NOR2X0 U14274 ( .IN1(n9342), .IN2(WX7294), .QN(n13875) );
  NOR2X0 U14275 ( .IN1(n13877), .IN2(n13878), .QN(n13857) );
  NOR2X0 U14276 ( .IN1(DFF_931_n1), .IN2(n9959), .QN(n13878) );
  NOR2X0 U14277 ( .IN1(n9991), .IN2(n11277), .QN(n13877) );
  NAND2X0 U14278 ( .IN1(n10210), .IN2(n8499), .QN(n11277) );
  NAND2X0 U14279 ( .IN1(n13879), .IN2(n13880), .QN(WX5870) );
  NOR2X0 U14280 ( .IN1(n13881), .IN2(n13882), .QN(n13880) );
  NOR2X0 U14281 ( .IN1(n13883), .IN2(n9934), .QN(n13882) );
  NOR2X0 U14282 ( .IN1(n9922), .IN2(n13051), .QN(n13881) );
  NAND2X0 U14283 ( .IN1(n13884), .IN2(n13885), .QN(n13051) );
  INVX0 U14284 ( .INP(n13886), .ZN(n13885) );
  NOR2X0 U14285 ( .IN1(n13887), .IN2(n13888), .QN(n13886) );
  NAND2X0 U14286 ( .IN1(n13888), .IN2(n13887), .QN(n13884) );
  NOR2X0 U14287 ( .IN1(n13889), .IN2(n13890), .QN(n13887) );
  NOR2X0 U14288 ( .IN1(n9849), .IN2(n9345), .QN(n13890) );
  INVX0 U14289 ( .INP(n13891), .ZN(n13889) );
  NAND2X0 U14290 ( .IN1(n9345), .IN2(n9849), .QN(n13891) );
  NAND2X0 U14291 ( .IN1(n13892), .IN2(n13893), .QN(n13888) );
  NAND2X0 U14292 ( .IN1(n9344), .IN2(WX7228), .QN(n13893) );
  INVX0 U14293 ( .INP(n13894), .ZN(n13892) );
  NOR2X0 U14294 ( .IN1(WX7228), .IN2(n9344), .QN(n13894) );
  NOR2X0 U14295 ( .IN1(n13895), .IN2(n13896), .QN(n13879) );
  NOR2X0 U14296 ( .IN1(DFF_932_n1), .IN2(n9959), .QN(n13896) );
  NOR2X0 U14297 ( .IN1(n9990), .IN2(n11278), .QN(n13895) );
  NAND2X0 U14298 ( .IN1(n10210), .IN2(n8500), .QN(n11278) );
  NAND2X0 U14299 ( .IN1(n13897), .IN2(n13898), .QN(WX5868) );
  NOR2X0 U14300 ( .IN1(n13899), .IN2(n13900), .QN(n13898) );
  NOR2X0 U14301 ( .IN1(n9943), .IN2(n13901), .QN(n13900) );
  NOR2X0 U14302 ( .IN1(n13073), .IN2(n9913), .QN(n13899) );
  INVX0 U14303 ( .INP(n13902), .ZN(n13073) );
  NAND2X0 U14304 ( .IN1(n13903), .IN2(n13904), .QN(n13902) );
  NAND2X0 U14305 ( .IN1(n13905), .IN2(n13906), .QN(n13904) );
  NAND2X0 U14306 ( .IN1(n13907), .IN2(n13908), .QN(n13906) );
  NAND2X0 U14307 ( .IN1(n9347), .IN2(WX7162), .QN(n13908) );
  NAND2X0 U14308 ( .IN1(n9346), .IN2(WX7290), .QN(n13907) );
  NOR2X0 U14309 ( .IN1(n13909), .IN2(n13910), .QN(n13905) );
  NOR2X0 U14310 ( .IN1(n9626), .IN2(WX7226), .QN(n13910) );
  NOR2X0 U14311 ( .IN1(n3637), .IN2(WX7354), .QN(n13909) );
  NAND2X0 U14312 ( .IN1(n13911), .IN2(n13912), .QN(n13903) );
  NAND2X0 U14313 ( .IN1(n13913), .IN2(n13914), .QN(n13912) );
  NAND2X0 U14314 ( .IN1(n9626), .IN2(WX7226), .QN(n13914) );
  NAND2X0 U14315 ( .IN1(n3637), .IN2(WX7354), .QN(n13913) );
  NOR2X0 U14316 ( .IN1(n13915), .IN2(n13916), .QN(n13911) );
  NOR2X0 U14317 ( .IN1(n9347), .IN2(WX7162), .QN(n13916) );
  NOR2X0 U14318 ( .IN1(n9346), .IN2(WX7290), .QN(n13915) );
  NOR2X0 U14319 ( .IN1(n13917), .IN2(n13918), .QN(n13897) );
  NOR2X0 U14320 ( .IN1(DFF_933_n1), .IN2(n9959), .QN(n13918) );
  NOR2X0 U14321 ( .IN1(n9990), .IN2(n11279), .QN(n13917) );
  NAND2X0 U14322 ( .IN1(n10210), .IN2(n8501), .QN(n11279) );
  NAND2X0 U14323 ( .IN1(n13919), .IN2(n13920), .QN(WX5866) );
  NOR2X0 U14324 ( .IN1(n13921), .IN2(n13922), .QN(n13920) );
  NOR2X0 U14325 ( .IN1(n13923), .IN2(n9934), .QN(n13922) );
  NOR2X0 U14326 ( .IN1(n9922), .IN2(n13095), .QN(n13921) );
  NAND2X0 U14327 ( .IN1(n13924), .IN2(n13925), .QN(n13095) );
  INVX0 U14328 ( .INP(n13926), .ZN(n13925) );
  NOR2X0 U14329 ( .IN1(n13927), .IN2(n13928), .QN(n13926) );
  NAND2X0 U14330 ( .IN1(n13928), .IN2(n13927), .QN(n13924) );
  NOR2X0 U14331 ( .IN1(n13929), .IN2(n13930), .QN(n13927) );
  INVX0 U14332 ( .INP(n13931), .ZN(n13930) );
  NAND2X0 U14333 ( .IN1(test_so62), .IN2(WX7352), .QN(n13931) );
  NOR2X0 U14334 ( .IN1(WX7352), .IN2(test_so62), .QN(n13929) );
  NAND2X0 U14335 ( .IN1(n13932), .IN2(n13933), .QN(n13928) );
  NAND2X0 U14336 ( .IN1(n9348), .IN2(WX7224), .QN(n13933) );
  INVX0 U14337 ( .INP(n13934), .ZN(n13932) );
  NOR2X0 U14338 ( .IN1(WX7224), .IN2(n9348), .QN(n13934) );
  NOR2X0 U14339 ( .IN1(n13935), .IN2(n13936), .QN(n13919) );
  NOR2X0 U14340 ( .IN1(DFF_934_n1), .IN2(n9958), .QN(n13936) );
  NOR2X0 U14341 ( .IN1(n9990), .IN2(n11280), .QN(n13935) );
  NAND2X0 U14342 ( .IN1(n10210), .IN2(n8502), .QN(n11280) );
  NAND2X0 U14343 ( .IN1(n13937), .IN2(n13938), .QN(WX5864) );
  NOR2X0 U14344 ( .IN1(n13939), .IN2(n13940), .QN(n13938) );
  NOR2X0 U14345 ( .IN1(n13941), .IN2(n9934), .QN(n13940) );
  NOR2X0 U14346 ( .IN1(n13117), .IN2(n9913), .QN(n13939) );
  INVX0 U14347 ( .INP(n13942), .ZN(n13117) );
  NAND2X0 U14348 ( .IN1(n13943), .IN2(n13944), .QN(n13942) );
  NAND2X0 U14349 ( .IN1(n13945), .IN2(n13946), .QN(n13944) );
  NAND2X0 U14350 ( .IN1(n13947), .IN2(n13948), .QN(n13946) );
  NAND2X0 U14351 ( .IN1(n9350), .IN2(WX7158), .QN(n13948) );
  NAND2X0 U14352 ( .IN1(n9349), .IN2(WX7286), .QN(n13947) );
  NOR2X0 U14353 ( .IN1(n13949), .IN2(n13950), .QN(n13945) );
  NOR2X0 U14354 ( .IN1(n9624), .IN2(WX7222), .QN(n13950) );
  NOR2X0 U14355 ( .IN1(n3641), .IN2(WX7350), .QN(n13949) );
  NAND2X0 U14356 ( .IN1(n13951), .IN2(n13952), .QN(n13943) );
  NAND2X0 U14357 ( .IN1(n13953), .IN2(n13954), .QN(n13952) );
  NAND2X0 U14358 ( .IN1(n9624), .IN2(WX7222), .QN(n13954) );
  NAND2X0 U14359 ( .IN1(n3641), .IN2(WX7350), .QN(n13953) );
  NOR2X0 U14360 ( .IN1(n13955), .IN2(n13956), .QN(n13951) );
  NOR2X0 U14361 ( .IN1(n9350), .IN2(WX7158), .QN(n13956) );
  NOR2X0 U14362 ( .IN1(n9349), .IN2(WX7286), .QN(n13955) );
  NOR2X0 U14363 ( .IN1(n13957), .IN2(n13958), .QN(n13937) );
  NOR2X0 U14364 ( .IN1(DFF_935_n1), .IN2(n9958), .QN(n13958) );
  NOR2X0 U14365 ( .IN1(n9990), .IN2(n11281), .QN(n13957) );
  NAND2X0 U14366 ( .IN1(test_so45), .IN2(n10215), .QN(n11281) );
  NAND2X0 U14367 ( .IN1(n13959), .IN2(n13960), .QN(WX5862) );
  NOR2X0 U14368 ( .IN1(n13961), .IN2(n13962), .QN(n13960) );
  NOR2X0 U14369 ( .IN1(n13963), .IN2(n9934), .QN(n13962) );
  NOR2X0 U14370 ( .IN1(n9922), .IN2(n13139), .QN(n13961) );
  NAND2X0 U14371 ( .IN1(n13964), .IN2(n13965), .QN(n13139) );
  INVX0 U14372 ( .INP(n13966), .ZN(n13965) );
  NOR2X0 U14373 ( .IN1(n13967), .IN2(n13968), .QN(n13966) );
  NAND2X0 U14374 ( .IN1(n13968), .IN2(n13967), .QN(n13964) );
  NOR2X0 U14375 ( .IN1(n13969), .IN2(n13970), .QN(n13967) );
  INVX0 U14376 ( .INP(n13971), .ZN(n13970) );
  NAND2X0 U14377 ( .IN1(test_so60), .IN2(WX7348), .QN(n13971) );
  NOR2X0 U14378 ( .IN1(WX7348), .IN2(test_so60), .QN(n13969) );
  NAND2X0 U14379 ( .IN1(n13972), .IN2(n13973), .QN(n13968) );
  NAND2X0 U14380 ( .IN1(n9352), .IN2(WX7156), .QN(n13973) );
  INVX0 U14381 ( .INP(n13974), .ZN(n13972) );
  NOR2X0 U14382 ( .IN1(WX7156), .IN2(n9352), .QN(n13974) );
  NOR2X0 U14383 ( .IN1(n13975), .IN2(n13976), .QN(n13959) );
  NOR2X0 U14384 ( .IN1(DFF_936_n1), .IN2(n9958), .QN(n13976) );
  NOR2X0 U14385 ( .IN1(n9990), .IN2(n11282), .QN(n13975) );
  NAND2X0 U14386 ( .IN1(n10210), .IN2(n8505), .QN(n11282) );
  NAND2X0 U14387 ( .IN1(n13977), .IN2(n13978), .QN(WX5860) );
  NOR2X0 U14388 ( .IN1(n13979), .IN2(n13980), .QN(n13978) );
  NOR2X0 U14389 ( .IN1(n13981), .IN2(n9934), .QN(n13980) );
  NOR2X0 U14390 ( .IN1(n13161), .IN2(n9913), .QN(n13979) );
  INVX0 U14391 ( .INP(n13982), .ZN(n13161) );
  NAND2X0 U14392 ( .IN1(n13983), .IN2(n13984), .QN(n13982) );
  NAND2X0 U14393 ( .IN1(n13985), .IN2(n13986), .QN(n13984) );
  NAND2X0 U14394 ( .IN1(n13987), .IN2(n13988), .QN(n13986) );
  NAND2X0 U14395 ( .IN1(n9354), .IN2(WX7154), .QN(n13988) );
  NAND2X0 U14396 ( .IN1(n9353), .IN2(WX7282), .QN(n13987) );
  NOR2X0 U14397 ( .IN1(n13989), .IN2(n13990), .QN(n13985) );
  NOR2X0 U14398 ( .IN1(n9622), .IN2(WX7218), .QN(n13990) );
  NOR2X0 U14399 ( .IN1(n3645), .IN2(WX7346), .QN(n13989) );
  NAND2X0 U14400 ( .IN1(n13991), .IN2(n13992), .QN(n13983) );
  NAND2X0 U14401 ( .IN1(n13993), .IN2(n13994), .QN(n13992) );
  NAND2X0 U14402 ( .IN1(n9622), .IN2(WX7218), .QN(n13994) );
  NAND2X0 U14403 ( .IN1(n3645), .IN2(WX7346), .QN(n13993) );
  NOR2X0 U14404 ( .IN1(n13995), .IN2(n13996), .QN(n13991) );
  NOR2X0 U14405 ( .IN1(n9354), .IN2(WX7154), .QN(n13996) );
  NOR2X0 U14406 ( .IN1(n9353), .IN2(WX7282), .QN(n13995) );
  NOR2X0 U14407 ( .IN1(n13997), .IN2(n13998), .QN(n13977) );
  NOR2X0 U14408 ( .IN1(DFF_937_n1), .IN2(n9958), .QN(n13998) );
  NOR2X0 U14409 ( .IN1(n9990), .IN2(n11283), .QN(n13997) );
  NAND2X0 U14410 ( .IN1(n10208), .IN2(n8506), .QN(n11283) );
  NAND2X0 U14411 ( .IN1(n13999), .IN2(n14000), .QN(WX5858) );
  NOR2X0 U14412 ( .IN1(n14001), .IN2(n14002), .QN(n14000) );
  NOR2X0 U14413 ( .IN1(n14003), .IN2(n9934), .QN(n14002) );
  NOR2X0 U14414 ( .IN1(n9923), .IN2(n13179), .QN(n14001) );
  NAND2X0 U14415 ( .IN1(n14004), .IN2(n14005), .QN(n13179) );
  INVX0 U14416 ( .INP(n14006), .ZN(n14005) );
  NOR2X0 U14417 ( .IN1(n14007), .IN2(n14008), .QN(n14006) );
  NAND2X0 U14418 ( .IN1(n14008), .IN2(n14007), .QN(n14004) );
  NOR2X0 U14419 ( .IN1(n14009), .IN2(n14010), .QN(n14007) );
  INVX0 U14420 ( .INP(n14011), .ZN(n14010) );
  NAND2X0 U14421 ( .IN1(test_so58), .IN2(WX7344), .QN(n14011) );
  NOR2X0 U14422 ( .IN1(WX7344), .IN2(test_so58), .QN(n14009) );
  NAND2X0 U14423 ( .IN1(n14012), .IN2(n14013), .QN(n14008) );
  NAND2X0 U14424 ( .IN1(n9355), .IN2(WX7216), .QN(n14013) );
  INVX0 U14425 ( .INP(n14014), .ZN(n14012) );
  NOR2X0 U14426 ( .IN1(WX7216), .IN2(n9355), .QN(n14014) );
  NOR2X0 U14427 ( .IN1(n14015), .IN2(n14016), .QN(n13999) );
  NOR2X0 U14428 ( .IN1(DFF_938_n1), .IN2(n9958), .QN(n14016) );
  NOR2X0 U14429 ( .IN1(n9990), .IN2(n11284), .QN(n14015) );
  NAND2X0 U14430 ( .IN1(n10209), .IN2(n8507), .QN(n11284) );
  NAND2X0 U14431 ( .IN1(n14017), .IN2(n14018), .QN(WX5856) );
  NOR2X0 U14432 ( .IN1(n14019), .IN2(n14020), .QN(n14018) );
  NOR2X0 U14433 ( .IN1(n14021), .IN2(n9934), .QN(n14020) );
  NOR2X0 U14434 ( .IN1(n13201), .IN2(n9913), .QN(n14019) );
  INVX0 U14435 ( .INP(n14022), .ZN(n13201) );
  NAND2X0 U14436 ( .IN1(n14023), .IN2(n14024), .QN(n14022) );
  NAND2X0 U14437 ( .IN1(n14025), .IN2(n14026), .QN(n14024) );
  NAND2X0 U14438 ( .IN1(n14027), .IN2(n14028), .QN(n14026) );
  NAND2X0 U14439 ( .IN1(n9357), .IN2(WX7150), .QN(n14028) );
  NAND2X0 U14440 ( .IN1(n9356), .IN2(WX7278), .QN(n14027) );
  NOR2X0 U14441 ( .IN1(n14029), .IN2(n14030), .QN(n14025) );
  NOR2X0 U14442 ( .IN1(n9506), .IN2(WX7214), .QN(n14030) );
  NOR2X0 U14443 ( .IN1(n3649), .IN2(WX7342), .QN(n14029) );
  NAND2X0 U14444 ( .IN1(n14031), .IN2(n14032), .QN(n14023) );
  NAND2X0 U14445 ( .IN1(n14033), .IN2(n14034), .QN(n14032) );
  NAND2X0 U14446 ( .IN1(n9506), .IN2(WX7214), .QN(n14034) );
  NAND2X0 U14447 ( .IN1(n3649), .IN2(WX7342), .QN(n14033) );
  NOR2X0 U14448 ( .IN1(n14035), .IN2(n14036), .QN(n14031) );
  NOR2X0 U14449 ( .IN1(n9357), .IN2(WX7150), .QN(n14036) );
  NOR2X0 U14450 ( .IN1(n9356), .IN2(WX7278), .QN(n14035) );
  NOR2X0 U14451 ( .IN1(n14037), .IN2(n14038), .QN(n14017) );
  NOR2X0 U14452 ( .IN1(DFF_939_n1), .IN2(n9958), .QN(n14038) );
  NOR2X0 U14453 ( .IN1(n9990), .IN2(n11285), .QN(n14037) );
  NAND2X0 U14454 ( .IN1(n10209), .IN2(n8508), .QN(n11285) );
  NAND2X0 U14455 ( .IN1(n14039), .IN2(n14040), .QN(WX5854) );
  NOR2X0 U14456 ( .IN1(n14041), .IN2(n14042), .QN(n14040) );
  NOR2X0 U14457 ( .IN1(n14043), .IN2(n9934), .QN(n14042) );
  NOR2X0 U14458 ( .IN1(n13219), .IN2(n9913), .QN(n14041) );
  INVX0 U14459 ( .INP(n14044), .ZN(n13219) );
  NAND2X0 U14460 ( .IN1(n14045), .IN2(n14046), .QN(n14044) );
  NAND2X0 U14461 ( .IN1(n14047), .IN2(n14048), .QN(n14046) );
  NAND2X0 U14462 ( .IN1(n14049), .IN2(n14050), .QN(n14048) );
  NAND2X0 U14463 ( .IN1(n9359), .IN2(WX7148), .QN(n14050) );
  NAND2X0 U14464 ( .IN1(n9358), .IN2(WX7276), .QN(n14049) );
  NOR2X0 U14465 ( .IN1(n14051), .IN2(n14052), .QN(n14047) );
  NOR2X0 U14466 ( .IN1(n9620), .IN2(WX7212), .QN(n14052) );
  NOR2X0 U14467 ( .IN1(n3651), .IN2(WX7340), .QN(n14051) );
  NAND2X0 U14468 ( .IN1(n14053), .IN2(n14054), .QN(n14045) );
  NAND2X0 U14469 ( .IN1(n14055), .IN2(n14056), .QN(n14054) );
  NAND2X0 U14470 ( .IN1(n9620), .IN2(WX7212), .QN(n14056) );
  NAND2X0 U14471 ( .IN1(n3651), .IN2(WX7340), .QN(n14055) );
  NOR2X0 U14472 ( .IN1(n14057), .IN2(n14058), .QN(n14053) );
  NOR2X0 U14473 ( .IN1(n9359), .IN2(WX7148), .QN(n14058) );
  NOR2X0 U14474 ( .IN1(n9358), .IN2(WX7276), .QN(n14057) );
  NOR2X0 U14475 ( .IN1(n14059), .IN2(n14060), .QN(n14039) );
  NOR2X0 U14476 ( .IN1(DFF_940_n1), .IN2(n9958), .QN(n14060) );
  NOR2X0 U14477 ( .IN1(n9990), .IN2(n11286), .QN(n14059) );
  NAND2X0 U14478 ( .IN1(n10209), .IN2(n8509), .QN(n11286) );
  NAND2X0 U14479 ( .IN1(n14061), .IN2(n14062), .QN(WX5852) );
  NOR2X0 U14480 ( .IN1(n14063), .IN2(n14064), .QN(n14062) );
  NOR2X0 U14481 ( .IN1(n14065), .IN2(n9934), .QN(n14064) );
  NOR2X0 U14482 ( .IN1(n13241), .IN2(n9914), .QN(n14063) );
  INVX0 U14483 ( .INP(n14066), .ZN(n13241) );
  NAND2X0 U14484 ( .IN1(n14067), .IN2(n14068), .QN(n14066) );
  NAND2X0 U14485 ( .IN1(n14069), .IN2(n14070), .QN(n14068) );
  NAND2X0 U14486 ( .IN1(n14071), .IN2(n14072), .QN(n14070) );
  NAND2X0 U14487 ( .IN1(n9361), .IN2(WX7146), .QN(n14072) );
  NAND2X0 U14488 ( .IN1(n9360), .IN2(WX7274), .QN(n14071) );
  NOR2X0 U14489 ( .IN1(n14073), .IN2(n14074), .QN(n14069) );
  NOR2X0 U14490 ( .IN1(n9619), .IN2(WX7210), .QN(n14074) );
  NOR2X0 U14491 ( .IN1(n3653), .IN2(WX7338), .QN(n14073) );
  NAND2X0 U14492 ( .IN1(n14075), .IN2(n14076), .QN(n14067) );
  NAND2X0 U14493 ( .IN1(n14077), .IN2(n14078), .QN(n14076) );
  NAND2X0 U14494 ( .IN1(n9619), .IN2(WX7210), .QN(n14078) );
  NAND2X0 U14495 ( .IN1(n3653), .IN2(WX7338), .QN(n14077) );
  NOR2X0 U14496 ( .IN1(n14079), .IN2(n14080), .QN(n14075) );
  NOR2X0 U14497 ( .IN1(n9361), .IN2(WX7146), .QN(n14080) );
  NOR2X0 U14498 ( .IN1(n9360), .IN2(WX7274), .QN(n14079) );
  NOR2X0 U14499 ( .IN1(n14081), .IN2(n14082), .QN(n14061) );
  NOR2X0 U14500 ( .IN1(DFF_941_n1), .IN2(n9958), .QN(n14082) );
  NOR2X0 U14501 ( .IN1(n9990), .IN2(n11287), .QN(n14081) );
  NAND2X0 U14502 ( .IN1(n10209), .IN2(n8510), .QN(n11287) );
  NAND2X0 U14503 ( .IN1(n14083), .IN2(n14084), .QN(WX5850) );
  NOR2X0 U14504 ( .IN1(n14085), .IN2(n14086), .QN(n14084) );
  NOR2X0 U14505 ( .IN1(n14087), .IN2(n9934), .QN(n14086) );
  NOR2X0 U14506 ( .IN1(n13259), .IN2(n9914), .QN(n14085) );
  INVX0 U14507 ( .INP(n14088), .ZN(n13259) );
  NAND2X0 U14508 ( .IN1(n14089), .IN2(n14090), .QN(n14088) );
  NAND2X0 U14509 ( .IN1(n14091), .IN2(n14092), .QN(n14090) );
  NAND2X0 U14510 ( .IN1(n14093), .IN2(n14094), .QN(n14092) );
  NAND2X0 U14511 ( .IN1(n9363), .IN2(WX7144), .QN(n14094) );
  NAND2X0 U14512 ( .IN1(n9362), .IN2(WX7272), .QN(n14093) );
  NOR2X0 U14513 ( .IN1(n14095), .IN2(n14096), .QN(n14091) );
  NOR2X0 U14514 ( .IN1(n9618), .IN2(WX7208), .QN(n14096) );
  NOR2X0 U14515 ( .IN1(n3655), .IN2(WX7336), .QN(n14095) );
  NAND2X0 U14516 ( .IN1(n14097), .IN2(n14098), .QN(n14089) );
  NAND2X0 U14517 ( .IN1(n14099), .IN2(n14100), .QN(n14098) );
  NAND2X0 U14518 ( .IN1(n9618), .IN2(WX7208), .QN(n14100) );
  NAND2X0 U14519 ( .IN1(n3655), .IN2(WX7336), .QN(n14099) );
  NOR2X0 U14520 ( .IN1(n14101), .IN2(n14102), .QN(n14097) );
  NOR2X0 U14521 ( .IN1(n9363), .IN2(WX7144), .QN(n14102) );
  NOR2X0 U14522 ( .IN1(n9362), .IN2(WX7272), .QN(n14101) );
  NOR2X0 U14523 ( .IN1(n14103), .IN2(n14104), .QN(n14083) );
  NOR2X0 U14524 ( .IN1(DFF_942_n1), .IN2(n9958), .QN(n14104) );
  NOR2X0 U14525 ( .IN1(n9990), .IN2(n11288), .QN(n14103) );
  NAND2X0 U14526 ( .IN1(n10209), .IN2(n8511), .QN(n11288) );
  NAND2X0 U14527 ( .IN1(n14105), .IN2(n14106), .QN(WX5848) );
  NOR2X0 U14528 ( .IN1(n14107), .IN2(n14108), .QN(n14106) );
  NOR2X0 U14529 ( .IN1(n14109), .IN2(n9934), .QN(n14108) );
  NOR2X0 U14530 ( .IN1(n13281), .IN2(n9914), .QN(n14107) );
  INVX0 U14531 ( .INP(n14110), .ZN(n13281) );
  NAND2X0 U14532 ( .IN1(n14111), .IN2(n14112), .QN(n14110) );
  NAND2X0 U14533 ( .IN1(n14113), .IN2(n14114), .QN(n14112) );
  NAND2X0 U14534 ( .IN1(n14115), .IN2(n14116), .QN(n14114) );
  NAND2X0 U14535 ( .IN1(n9365), .IN2(WX7142), .QN(n14116) );
  NAND2X0 U14536 ( .IN1(n9364), .IN2(WX7270), .QN(n14115) );
  NOR2X0 U14537 ( .IN1(n14117), .IN2(n14118), .QN(n14113) );
  NOR2X0 U14538 ( .IN1(n9617), .IN2(WX7206), .QN(n14118) );
  NOR2X0 U14539 ( .IN1(n3657), .IN2(WX7334), .QN(n14117) );
  NAND2X0 U14540 ( .IN1(n14119), .IN2(n14120), .QN(n14111) );
  NAND2X0 U14541 ( .IN1(n14121), .IN2(n14122), .QN(n14120) );
  NAND2X0 U14542 ( .IN1(n9617), .IN2(WX7206), .QN(n14122) );
  NAND2X0 U14543 ( .IN1(n3657), .IN2(WX7334), .QN(n14121) );
  NOR2X0 U14544 ( .IN1(n14123), .IN2(n14124), .QN(n14119) );
  NOR2X0 U14545 ( .IN1(n9365), .IN2(WX7142), .QN(n14124) );
  NOR2X0 U14546 ( .IN1(n9364), .IN2(WX7270), .QN(n14123) );
  NOR2X0 U14547 ( .IN1(n14125), .IN2(n14126), .QN(n14105) );
  NOR2X0 U14548 ( .IN1(DFF_943_n1), .IN2(n9958), .QN(n14126) );
  NOR2X0 U14549 ( .IN1(n9990), .IN2(n11289), .QN(n14125) );
  NAND2X0 U14550 ( .IN1(n10209), .IN2(n8512), .QN(n11289) );
  NAND2X0 U14551 ( .IN1(n14127), .IN2(n14128), .QN(WX5846) );
  NOR2X0 U14552 ( .IN1(n14129), .IN2(n14130), .QN(n14128) );
  NOR2X0 U14553 ( .IN1(n9944), .IN2(n14131), .QN(n14130) );
  NOR2X0 U14554 ( .IN1(n13299), .IN2(n9914), .QN(n14129) );
  NOR2X0 U14555 ( .IN1(n14132), .IN2(n14133), .QN(n13299) );
  INVX0 U14556 ( .INP(n14134), .ZN(n14133) );
  NAND2X0 U14557 ( .IN1(n14135), .IN2(n14136), .QN(n14134) );
  NOR2X0 U14558 ( .IN1(n14136), .IN2(n14135), .QN(n14132) );
  NAND2X0 U14559 ( .IN1(n14137), .IN2(n14138), .QN(n14135) );
  NAND2X0 U14560 ( .IN1(n9104), .IN2(n14139), .QN(n14138) );
  INVX0 U14561 ( .INP(n14140), .ZN(n14137) );
  NOR2X0 U14562 ( .IN1(n14139), .IN2(n9104), .QN(n14140) );
  NOR2X0 U14563 ( .IN1(n14141), .IN2(n14142), .QN(n14139) );
  INVX0 U14564 ( .INP(n14143), .ZN(n14142) );
  NAND2X0 U14565 ( .IN1(n18426), .IN2(WX7332), .QN(n14143) );
  NOR2X0 U14566 ( .IN1(WX7332), .IN2(n18426), .QN(n14141) );
  NOR2X0 U14567 ( .IN1(n14144), .IN2(n14145), .QN(n14136) );
  INVX0 U14568 ( .INP(n14146), .ZN(n14145) );
  NAND2X0 U14569 ( .IN1(n9103), .IN2(n10017), .QN(n14146) );
  NOR2X0 U14570 ( .IN1(n10006), .IN2(n9103), .QN(n14144) );
  NOR2X0 U14571 ( .IN1(n14147), .IN2(n14148), .QN(n14127) );
  NOR2X0 U14572 ( .IN1(DFF_944_n1), .IN2(n9958), .QN(n14148) );
  NOR2X0 U14573 ( .IN1(n9989), .IN2(n11290), .QN(n14147) );
  NAND2X0 U14574 ( .IN1(n10209), .IN2(n8513), .QN(n11290) );
  NAND2X0 U14575 ( .IN1(n14149), .IN2(n14150), .QN(WX5844) );
  NOR2X0 U14576 ( .IN1(n14151), .IN2(n14152), .QN(n14150) );
  NOR2X0 U14577 ( .IN1(n14153), .IN2(n9934), .QN(n14152) );
  NOR2X0 U14578 ( .IN1(n13321), .IN2(n9914), .QN(n14151) );
  NOR2X0 U14579 ( .IN1(n14154), .IN2(n14155), .QN(n13321) );
  INVX0 U14580 ( .INP(n14156), .ZN(n14155) );
  NAND2X0 U14581 ( .IN1(n14157), .IN2(n14158), .QN(n14156) );
  NOR2X0 U14582 ( .IN1(n14158), .IN2(n14157), .QN(n14154) );
  NAND2X0 U14583 ( .IN1(n14159), .IN2(n14160), .QN(n14157) );
  NAND2X0 U14584 ( .IN1(n9106), .IN2(n14161), .QN(n14160) );
  INVX0 U14585 ( .INP(n14162), .ZN(n14159) );
  NOR2X0 U14586 ( .IN1(n14161), .IN2(n9106), .QN(n14162) );
  NOR2X0 U14587 ( .IN1(n14163), .IN2(n14164), .QN(n14161) );
  INVX0 U14588 ( .INP(n14165), .ZN(n14164) );
  NAND2X0 U14589 ( .IN1(n18425), .IN2(WX7330), .QN(n14165) );
  NOR2X0 U14590 ( .IN1(WX7330), .IN2(n18425), .QN(n14163) );
  NOR2X0 U14591 ( .IN1(n14166), .IN2(n14167), .QN(n14158) );
  INVX0 U14592 ( .INP(n14168), .ZN(n14167) );
  NAND2X0 U14593 ( .IN1(n9105), .IN2(n10017), .QN(n14168) );
  NOR2X0 U14594 ( .IN1(n10007), .IN2(n9105), .QN(n14166) );
  NOR2X0 U14595 ( .IN1(n14169), .IN2(n14170), .QN(n14149) );
  NOR2X0 U14596 ( .IN1(n9976), .IN2(n9857), .QN(n14170) );
  NOR2X0 U14597 ( .IN1(n9989), .IN2(n11291), .QN(n14169) );
  NAND2X0 U14598 ( .IN1(n10209), .IN2(n8514), .QN(n11291) );
  NAND2X0 U14599 ( .IN1(n14171), .IN2(n14172), .QN(WX5842) );
  NOR2X0 U14600 ( .IN1(n14173), .IN2(n14174), .QN(n14172) );
  NOR2X0 U14601 ( .IN1(n10563), .IN2(n14175), .QN(n14174) );
  NOR2X0 U14602 ( .IN1(n13343), .IN2(n9914), .QN(n14173) );
  NOR2X0 U14603 ( .IN1(n14176), .IN2(n14177), .QN(n13343) );
  INVX0 U14604 ( .INP(n14178), .ZN(n14177) );
  NAND2X0 U14605 ( .IN1(n14179), .IN2(n14180), .QN(n14178) );
  NOR2X0 U14606 ( .IN1(n14180), .IN2(n14179), .QN(n14176) );
  NAND2X0 U14607 ( .IN1(n14181), .IN2(n14182), .QN(n14179) );
  NAND2X0 U14608 ( .IN1(n9108), .IN2(n14183), .QN(n14182) );
  INVX0 U14609 ( .INP(n14184), .ZN(n14181) );
  NOR2X0 U14610 ( .IN1(n14183), .IN2(n9108), .QN(n14184) );
  NOR2X0 U14611 ( .IN1(n14185), .IN2(n14186), .QN(n14183) );
  INVX0 U14612 ( .INP(n14187), .ZN(n14186) );
  NAND2X0 U14613 ( .IN1(n18424), .IN2(WX7328), .QN(n14187) );
  NOR2X0 U14614 ( .IN1(WX7328), .IN2(n18424), .QN(n14185) );
  NOR2X0 U14615 ( .IN1(n14188), .IN2(n14189), .QN(n14180) );
  INVX0 U14616 ( .INP(n14190), .ZN(n14189) );
  NAND2X0 U14617 ( .IN1(n9107), .IN2(n10017), .QN(n14190) );
  NOR2X0 U14618 ( .IN1(n10007), .IN2(n9107), .QN(n14188) );
  NOR2X0 U14619 ( .IN1(n14191), .IN2(n14192), .QN(n14171) );
  NOR2X0 U14620 ( .IN1(DFF_946_n1), .IN2(n9962), .QN(n14192) );
  NOR2X0 U14621 ( .IN1(n9989), .IN2(n11292), .QN(n14191) );
  NAND2X0 U14622 ( .IN1(n10208), .IN2(n8515), .QN(n11292) );
  NAND2X0 U14623 ( .IN1(n14193), .IN2(n14194), .QN(WX5840) );
  NOR2X0 U14624 ( .IN1(n14195), .IN2(n14196), .QN(n14194) );
  NOR2X0 U14625 ( .IN1(n14197), .IN2(n9935), .QN(n14196) );
  NOR2X0 U14626 ( .IN1(n13365), .IN2(n9914), .QN(n14195) );
  NOR2X0 U14627 ( .IN1(n14198), .IN2(n14199), .QN(n13365) );
  INVX0 U14628 ( .INP(n14200), .ZN(n14199) );
  NAND2X0 U14629 ( .IN1(n14201), .IN2(n14202), .QN(n14200) );
  NOR2X0 U14630 ( .IN1(n14202), .IN2(n14201), .QN(n14198) );
  NAND2X0 U14631 ( .IN1(n14203), .IN2(n14204), .QN(n14201) );
  NAND2X0 U14632 ( .IN1(n9110), .IN2(n14205), .QN(n14204) );
  INVX0 U14633 ( .INP(n14206), .ZN(n14203) );
  NOR2X0 U14634 ( .IN1(n14205), .IN2(n9110), .QN(n14206) );
  NOR2X0 U14635 ( .IN1(n14207), .IN2(n14208), .QN(n14205) );
  INVX0 U14636 ( .INP(n14209), .ZN(n14208) );
  NAND2X0 U14637 ( .IN1(n18423), .IN2(WX7326), .QN(n14209) );
  NOR2X0 U14638 ( .IN1(WX7326), .IN2(n18423), .QN(n14207) );
  NOR2X0 U14639 ( .IN1(n14210), .IN2(n14211), .QN(n14202) );
  INVX0 U14640 ( .INP(n14212), .ZN(n14211) );
  NAND2X0 U14641 ( .IN1(n9109), .IN2(n10017), .QN(n14212) );
  NOR2X0 U14642 ( .IN1(n10007), .IN2(n9109), .QN(n14210) );
  NOR2X0 U14643 ( .IN1(n14213), .IN2(n14214), .QN(n14193) );
  NOR2X0 U14644 ( .IN1(DFF_947_n1), .IN2(n9974), .QN(n14214) );
  NOR2X0 U14645 ( .IN1(n9989), .IN2(n11293), .QN(n14213) );
  NAND2X0 U14646 ( .IN1(n10208), .IN2(n8516), .QN(n11293) );
  NAND2X0 U14647 ( .IN1(n14215), .IN2(n14216), .QN(WX5838) );
  NOR2X0 U14648 ( .IN1(n14217), .IN2(n14218), .QN(n14216) );
  NOR2X0 U14649 ( .IN1(n10563), .IN2(n14219), .QN(n14218) );
  NOR2X0 U14650 ( .IN1(n13387), .IN2(n9914), .QN(n14217) );
  NOR2X0 U14651 ( .IN1(n14220), .IN2(n14221), .QN(n13387) );
  INVX0 U14652 ( .INP(n14222), .ZN(n14221) );
  NAND2X0 U14653 ( .IN1(n14223), .IN2(n14224), .QN(n14222) );
  NOR2X0 U14654 ( .IN1(n14224), .IN2(n14223), .QN(n14220) );
  NAND2X0 U14655 ( .IN1(n14225), .IN2(n14226), .QN(n14223) );
  NAND2X0 U14656 ( .IN1(n9112), .IN2(n14227), .QN(n14226) );
  INVX0 U14657 ( .INP(n14228), .ZN(n14225) );
  NOR2X0 U14658 ( .IN1(n14227), .IN2(n9112), .QN(n14228) );
  NOR2X0 U14659 ( .IN1(n14229), .IN2(n14230), .QN(n14227) );
  INVX0 U14660 ( .INP(n14231), .ZN(n14230) );
  NAND2X0 U14661 ( .IN1(n18422), .IN2(WX7324), .QN(n14231) );
  NOR2X0 U14662 ( .IN1(WX7324), .IN2(n18422), .QN(n14229) );
  NOR2X0 U14663 ( .IN1(n14232), .IN2(n14233), .QN(n14224) );
  INVX0 U14664 ( .INP(n14234), .ZN(n14233) );
  NAND2X0 U14665 ( .IN1(n9111), .IN2(n10017), .QN(n14234) );
  NOR2X0 U14666 ( .IN1(n10007), .IN2(n9111), .QN(n14232) );
  NOR2X0 U14667 ( .IN1(n14235), .IN2(n14236), .QN(n14215) );
  NOR2X0 U14668 ( .IN1(DFF_948_n1), .IN2(n9975), .QN(n14236) );
  NOR2X0 U14669 ( .IN1(n9989), .IN2(n11294), .QN(n14235) );
  NAND2X0 U14670 ( .IN1(n10208), .IN2(n8517), .QN(n11294) );
  NAND2X0 U14671 ( .IN1(n14237), .IN2(n14238), .QN(WX5836) );
  NOR2X0 U14672 ( .IN1(n14239), .IN2(n14240), .QN(n14238) );
  NOR2X0 U14673 ( .IN1(n14241), .IN2(n9935), .QN(n14240) );
  NOR2X0 U14674 ( .IN1(n9924), .IN2(n13409), .QN(n14239) );
  NAND2X0 U14675 ( .IN1(n14242), .IN2(n14243), .QN(n13409) );
  NAND2X0 U14676 ( .IN1(n14244), .IN2(n14245), .QN(n14243) );
  INVX0 U14677 ( .INP(n14246), .ZN(n14242) );
  NOR2X0 U14678 ( .IN1(n14245), .IN2(n14244), .QN(n14246) );
  NAND2X0 U14679 ( .IN1(n14247), .IN2(n14248), .QN(n14244) );
  NAND2X0 U14680 ( .IN1(n14249), .IN2(WX7258), .QN(n14248) );
  NAND2X0 U14681 ( .IN1(n14250), .IN2(n14251), .QN(n14249) );
  NAND2X0 U14682 ( .IN1(test_so63), .IN2(WX7194), .QN(n14251) );
  NAND2X0 U14683 ( .IN1(n9113), .IN2(n9829), .QN(n14250) );
  NAND2X0 U14684 ( .IN1(n9114), .IN2(n14252), .QN(n14247) );
  NOR2X0 U14685 ( .IN1(n14253), .IN2(n14254), .QN(n14252) );
  NOR2X0 U14686 ( .IN1(test_so63), .IN2(WX7194), .QN(n14254) );
  NOR2X0 U14687 ( .IN1(n9113), .IN2(n9829), .QN(n14253) );
  NOR2X0 U14688 ( .IN1(n14255), .IN2(n14256), .QN(n14245) );
  INVX0 U14689 ( .INP(n14257), .ZN(n14256) );
  NAND2X0 U14690 ( .IN1(n18421), .IN2(n10017), .QN(n14257) );
  NOR2X0 U14691 ( .IN1(n10007), .IN2(n18421), .QN(n14255) );
  NOR2X0 U14692 ( .IN1(n14258), .IN2(n14259), .QN(n14237) );
  NOR2X0 U14693 ( .IN1(DFF_949_n1), .IN2(n9975), .QN(n14259) );
  NOR2X0 U14694 ( .IN1(n9989), .IN2(n11295), .QN(n14258) );
  NAND2X0 U14695 ( .IN1(n10208), .IN2(n8518), .QN(n11295) );
  NAND2X0 U14696 ( .IN1(n14260), .IN2(n14261), .QN(WX5834) );
  NOR2X0 U14697 ( .IN1(n14262), .IN2(n14263), .QN(n14261) );
  NOR2X0 U14698 ( .IN1(n10563), .IN2(n14264), .QN(n14263) );
  NOR2X0 U14699 ( .IN1(n13431), .IN2(n9914), .QN(n14262) );
  NOR2X0 U14700 ( .IN1(n14265), .IN2(n14266), .QN(n13431) );
  INVX0 U14701 ( .INP(n14267), .ZN(n14266) );
  NAND2X0 U14702 ( .IN1(n14268), .IN2(n14269), .QN(n14267) );
  NOR2X0 U14703 ( .IN1(n14269), .IN2(n14268), .QN(n14265) );
  NAND2X0 U14704 ( .IN1(n14270), .IN2(n14271), .QN(n14268) );
  NAND2X0 U14705 ( .IN1(n9116), .IN2(n14272), .QN(n14271) );
  INVX0 U14706 ( .INP(n14273), .ZN(n14270) );
  NOR2X0 U14707 ( .IN1(n14272), .IN2(n9116), .QN(n14273) );
  NOR2X0 U14708 ( .IN1(n14274), .IN2(n14275), .QN(n14272) );
  INVX0 U14709 ( .INP(n14276), .ZN(n14275) );
  NAND2X0 U14710 ( .IN1(n18420), .IN2(WX7320), .QN(n14276) );
  NOR2X0 U14711 ( .IN1(WX7320), .IN2(n18420), .QN(n14274) );
  NOR2X0 U14712 ( .IN1(n14277), .IN2(n14278), .QN(n14269) );
  INVX0 U14713 ( .INP(n14279), .ZN(n14278) );
  NAND2X0 U14714 ( .IN1(n9115), .IN2(n10017), .QN(n14279) );
  NOR2X0 U14715 ( .IN1(n10007), .IN2(n9115), .QN(n14277) );
  NOR2X0 U14716 ( .IN1(n14280), .IN2(n14281), .QN(n14260) );
  NOR2X0 U14717 ( .IN1(DFF_950_n1), .IN2(n9974), .QN(n14281) );
  NOR2X0 U14718 ( .IN1(n9989), .IN2(n11296), .QN(n14280) );
  NAND2X0 U14719 ( .IN1(n10208), .IN2(n8519), .QN(n11296) );
  NAND2X0 U14720 ( .IN1(n14282), .IN2(n14283), .QN(WX5832) );
  NOR2X0 U14721 ( .IN1(n14284), .IN2(n14285), .QN(n14283) );
  NOR2X0 U14722 ( .IN1(n14286), .IN2(n9941), .QN(n14285) );
  NOR2X0 U14723 ( .IN1(n9924), .IN2(n13453), .QN(n14284) );
  NAND2X0 U14724 ( .IN1(n14287), .IN2(n14288), .QN(n13453) );
  INVX0 U14725 ( .INP(n14289), .ZN(n14288) );
  NOR2X0 U14726 ( .IN1(n14290), .IN2(n14291), .QN(n14289) );
  NAND2X0 U14727 ( .IN1(n14291), .IN2(n14290), .QN(n14287) );
  NOR2X0 U14728 ( .IN1(n14292), .IN2(n14293), .QN(n14290) );
  INVX0 U14729 ( .INP(n14294), .ZN(n14293) );
  NAND2X0 U14730 ( .IN1(n9611), .IN2(n14295), .QN(n14294) );
  NOR2X0 U14731 ( .IN1(n14295), .IN2(n9611), .QN(n14292) );
  NOR2X0 U14732 ( .IN1(n14296), .IN2(n14297), .QN(n14295) );
  INVX0 U14733 ( .INP(n14298), .ZN(n14297) );
  NAND2X0 U14734 ( .IN1(test_so61), .IN2(n8428), .QN(n14298) );
  NOR2X0 U14735 ( .IN1(n8428), .IN2(test_so61), .QN(n14296) );
  NAND2X0 U14736 ( .IN1(n14299), .IN2(n14300), .QN(n14291) );
  NAND2X0 U14737 ( .IN1(n9117), .IN2(n10018), .QN(n14300) );
  INVX0 U14738 ( .INP(n14301), .ZN(n14299) );
  NOR2X0 U14739 ( .IN1(n10007), .IN2(n9117), .QN(n14301) );
  NOR2X0 U14740 ( .IN1(n14302), .IN2(n14303), .QN(n14282) );
  NOR2X0 U14741 ( .IN1(DFF_951_n1), .IN2(n9975), .QN(n14303) );
  NOR2X0 U14742 ( .IN1(n9989), .IN2(n11297), .QN(n14302) );
  NAND2X0 U14743 ( .IN1(n10208), .IN2(n8520), .QN(n11297) );
  NAND2X0 U14744 ( .IN1(n14304), .IN2(n14305), .QN(WX5830) );
  NOR2X0 U14745 ( .IN1(n14306), .IN2(n14307), .QN(n14305) );
  NOR2X0 U14746 ( .IN1(n14308), .IN2(n10563), .QN(n14307) );
  NOR2X0 U14747 ( .IN1(n13475), .IN2(n9914), .QN(n14306) );
  NOR2X0 U14748 ( .IN1(n14309), .IN2(n14310), .QN(n13475) );
  INVX0 U14749 ( .INP(n14311), .ZN(n14310) );
  NAND2X0 U14750 ( .IN1(n14312), .IN2(n14313), .QN(n14311) );
  NOR2X0 U14751 ( .IN1(n14313), .IN2(n14312), .QN(n14309) );
  NAND2X0 U14752 ( .IN1(n14314), .IN2(n14315), .QN(n14312) );
  NAND2X0 U14753 ( .IN1(n9119), .IN2(n14316), .QN(n14315) );
  INVX0 U14754 ( .INP(n14317), .ZN(n14314) );
  NOR2X0 U14755 ( .IN1(n14316), .IN2(n9119), .QN(n14317) );
  NOR2X0 U14756 ( .IN1(n14318), .IN2(n14319), .QN(n14316) );
  INVX0 U14757 ( .INP(n14320), .ZN(n14319) );
  NAND2X0 U14758 ( .IN1(n18418), .IN2(WX7316), .QN(n14320) );
  NOR2X0 U14759 ( .IN1(WX7316), .IN2(n18418), .QN(n14318) );
  NOR2X0 U14760 ( .IN1(n14321), .IN2(n14322), .QN(n14313) );
  INVX0 U14761 ( .INP(n14323), .ZN(n14322) );
  NAND2X0 U14762 ( .IN1(n9118), .IN2(n10018), .QN(n14323) );
  NOR2X0 U14763 ( .IN1(n10007), .IN2(n9118), .QN(n14321) );
  NOR2X0 U14764 ( .IN1(n14324), .IN2(n14325), .QN(n14304) );
  NOR2X0 U14765 ( .IN1(DFF_952_n1), .IN2(n9975), .QN(n14325) );
  NOR2X0 U14766 ( .IN1(n9989), .IN2(n11298), .QN(n14324) );
  NAND2X0 U14767 ( .IN1(test_so44), .IN2(n10215), .QN(n11298) );
  NAND2X0 U14768 ( .IN1(n14326), .IN2(n14327), .QN(WX5828) );
  NOR2X0 U14769 ( .IN1(n14328), .IN2(n14329), .QN(n14327) );
  NOR2X0 U14770 ( .IN1(n14330), .IN2(n9941), .QN(n14329) );
  NOR2X0 U14771 ( .IN1(n9924), .IN2(n13497), .QN(n14328) );
  NAND2X0 U14772 ( .IN1(n14331), .IN2(n14332), .QN(n13497) );
  INVX0 U14773 ( .INP(n14333), .ZN(n14332) );
  NOR2X0 U14774 ( .IN1(n14334), .IN2(n14335), .QN(n14333) );
  NAND2X0 U14775 ( .IN1(n14335), .IN2(n14334), .QN(n14331) );
  NOR2X0 U14776 ( .IN1(n14336), .IN2(n14337), .QN(n14334) );
  INVX0 U14777 ( .INP(n14338), .ZN(n14337) );
  NAND2X0 U14778 ( .IN1(n9609), .IN2(n14339), .QN(n14338) );
  NOR2X0 U14779 ( .IN1(n14339), .IN2(n9609), .QN(n14336) );
  NOR2X0 U14780 ( .IN1(n14340), .IN2(n14341), .QN(n14339) );
  INVX0 U14781 ( .INP(n14342), .ZN(n14341) );
  NAND2X0 U14782 ( .IN1(test_so59), .IN2(n8430), .QN(n14342) );
  NOR2X0 U14783 ( .IN1(n8430), .IN2(test_so59), .QN(n14340) );
  NAND2X0 U14784 ( .IN1(n14343), .IN2(n14344), .QN(n14335) );
  NAND2X0 U14785 ( .IN1(n9120), .IN2(n10018), .QN(n14344) );
  INVX0 U14786 ( .INP(n14345), .ZN(n14343) );
  NOR2X0 U14787 ( .IN1(n10007), .IN2(n9120), .QN(n14345) );
  NOR2X0 U14788 ( .IN1(n14346), .IN2(n14347), .QN(n14326) );
  NOR2X0 U14789 ( .IN1(DFF_953_n1), .IN2(n9975), .QN(n14347) );
  NOR2X0 U14790 ( .IN1(n9989), .IN2(n11299), .QN(n14346) );
  NAND2X0 U14791 ( .IN1(n10208), .IN2(n8523), .QN(n11299) );
  NAND2X0 U14792 ( .IN1(n14348), .IN2(n14349), .QN(WX5826) );
  NOR2X0 U14793 ( .IN1(n14350), .IN2(n14351), .QN(n14349) );
  NOR2X0 U14794 ( .IN1(n14352), .IN2(n9940), .QN(n14351) );
  NOR2X0 U14795 ( .IN1(n13519), .IN2(n9914), .QN(n14350) );
  NOR2X0 U14796 ( .IN1(n14353), .IN2(n14354), .QN(n13519) );
  INVX0 U14797 ( .INP(n14355), .ZN(n14354) );
  NAND2X0 U14798 ( .IN1(n14356), .IN2(n14357), .QN(n14355) );
  NOR2X0 U14799 ( .IN1(n14357), .IN2(n14356), .QN(n14353) );
  NAND2X0 U14800 ( .IN1(n14358), .IN2(n14359), .QN(n14356) );
  NAND2X0 U14801 ( .IN1(n9122), .IN2(n14360), .QN(n14359) );
  INVX0 U14802 ( .INP(n14361), .ZN(n14358) );
  NOR2X0 U14803 ( .IN1(n14360), .IN2(n9122), .QN(n14361) );
  NOR2X0 U14804 ( .IN1(n14362), .IN2(n14363), .QN(n14360) );
  INVX0 U14805 ( .INP(n14364), .ZN(n14363) );
  NAND2X0 U14806 ( .IN1(n18416), .IN2(WX7312), .QN(n14364) );
  NOR2X0 U14807 ( .IN1(WX7312), .IN2(n18416), .QN(n14362) );
  NOR2X0 U14808 ( .IN1(n14365), .IN2(n14366), .QN(n14357) );
  INVX0 U14809 ( .INP(n14367), .ZN(n14366) );
  NAND2X0 U14810 ( .IN1(n9121), .IN2(n10018), .QN(n14367) );
  NOR2X0 U14811 ( .IN1(n10007), .IN2(n9121), .QN(n14365) );
  NOR2X0 U14812 ( .IN1(n14368), .IN2(n14369), .QN(n14348) );
  NOR2X0 U14813 ( .IN1(DFF_954_n1), .IN2(n9974), .QN(n14369) );
  NOR2X0 U14814 ( .IN1(n9989), .IN2(n11300), .QN(n14368) );
  NAND2X0 U14815 ( .IN1(n10208), .IN2(n8524), .QN(n11300) );
  NAND2X0 U14816 ( .IN1(n14370), .IN2(n14371), .QN(WX5824) );
  NOR2X0 U14817 ( .IN1(n14372), .IN2(n14373), .QN(n14371) );
  NOR2X0 U14818 ( .IN1(n14374), .IN2(n9940), .QN(n14373) );
  NOR2X0 U14819 ( .IN1(n9924), .IN2(n13542), .QN(n14372) );
  NAND2X0 U14820 ( .IN1(n14375), .IN2(n14376), .QN(n13542) );
  INVX0 U14821 ( .INP(n14377), .ZN(n14376) );
  NOR2X0 U14822 ( .IN1(n14378), .IN2(n14379), .QN(n14377) );
  NAND2X0 U14823 ( .IN1(n14379), .IN2(n14378), .QN(n14375) );
  INVX0 U14824 ( .INP(n14380), .ZN(n14378) );
  NAND2X0 U14825 ( .IN1(n14381), .IN2(n14382), .QN(n14380) );
  NAND2X0 U14826 ( .IN1(n14383), .IN2(WX7246), .QN(n14382) );
  NAND2X0 U14827 ( .IN1(n14384), .IN2(n14385), .QN(n14383) );
  NAND2X0 U14828 ( .IN1(test_so57), .IN2(WX7182), .QN(n14385) );
  NAND2X0 U14829 ( .IN1(n9123), .IN2(n9841), .QN(n14384) );
  NAND2X0 U14830 ( .IN1(n9124), .IN2(n14386), .QN(n14381) );
  NOR2X0 U14831 ( .IN1(n14387), .IN2(n14388), .QN(n14386) );
  NOR2X0 U14832 ( .IN1(test_so57), .IN2(WX7182), .QN(n14388) );
  NOR2X0 U14833 ( .IN1(n9123), .IN2(n9841), .QN(n14387) );
  NAND2X0 U14834 ( .IN1(n14389), .IN2(n14390), .QN(n14379) );
  NAND2X0 U14835 ( .IN1(n9607), .IN2(n10018), .QN(n14390) );
  NAND2X0 U14836 ( .IN1(TM1), .IN2(WX7310), .QN(n14389) );
  NOR2X0 U14837 ( .IN1(n14391), .IN2(n14392), .QN(n14370) );
  NOR2X0 U14838 ( .IN1(DFF_955_n1), .IN2(n9975), .QN(n14392) );
  NOR2X0 U14839 ( .IN1(n9989), .IN2(n11301), .QN(n14391) );
  NAND2X0 U14840 ( .IN1(n10207), .IN2(n8525), .QN(n11301) );
  NAND2X0 U14841 ( .IN1(n14393), .IN2(n14394), .QN(WX5822) );
  NOR2X0 U14842 ( .IN1(n14395), .IN2(n14396), .QN(n14394) );
  NOR2X0 U14843 ( .IN1(n14397), .IN2(n9940), .QN(n14396) );
  NOR2X0 U14844 ( .IN1(n13564), .IN2(n9914), .QN(n14395) );
  NOR2X0 U14845 ( .IN1(n14398), .IN2(n14399), .QN(n13564) );
  INVX0 U14846 ( .INP(n14400), .ZN(n14399) );
  NAND2X0 U14847 ( .IN1(n14401), .IN2(n14402), .QN(n14400) );
  NOR2X0 U14848 ( .IN1(n14402), .IN2(n14401), .QN(n14398) );
  NAND2X0 U14849 ( .IN1(n14403), .IN2(n14404), .QN(n14401) );
  NAND2X0 U14850 ( .IN1(n9126), .IN2(n14405), .QN(n14404) );
  INVX0 U14851 ( .INP(n14406), .ZN(n14403) );
  NOR2X0 U14852 ( .IN1(n14405), .IN2(n9126), .QN(n14406) );
  NOR2X0 U14853 ( .IN1(n14407), .IN2(n14408), .QN(n14405) );
  INVX0 U14854 ( .INP(n14409), .ZN(n14408) );
  NAND2X0 U14855 ( .IN1(n18415), .IN2(WX7308), .QN(n14409) );
  NOR2X0 U14856 ( .IN1(WX7308), .IN2(n18415), .QN(n14407) );
  NOR2X0 U14857 ( .IN1(n14410), .IN2(n14411), .QN(n14402) );
  INVX0 U14858 ( .INP(n14412), .ZN(n14411) );
  NAND2X0 U14859 ( .IN1(n9125), .IN2(n10018), .QN(n14412) );
  NOR2X0 U14860 ( .IN1(n10007), .IN2(n9125), .QN(n14410) );
  NOR2X0 U14861 ( .IN1(n14413), .IN2(n14414), .QN(n14393) );
  NOR2X0 U14862 ( .IN1(DFF_956_n1), .IN2(n9974), .QN(n14414) );
  NOR2X0 U14863 ( .IN1(n9988), .IN2(n11302), .QN(n14413) );
  NAND2X0 U14864 ( .IN1(n10207), .IN2(n8526), .QN(n11302) );
  NAND2X0 U14865 ( .IN1(n14415), .IN2(n14416), .QN(WX5820) );
  NOR2X0 U14866 ( .IN1(n14417), .IN2(n14418), .QN(n14416) );
  NOR2X0 U14867 ( .IN1(n14419), .IN2(n9940), .QN(n14418) );
  NOR2X0 U14868 ( .IN1(n13586), .IN2(n9915), .QN(n14417) );
  NOR2X0 U14869 ( .IN1(n14420), .IN2(n14421), .QN(n13586) );
  INVX0 U14870 ( .INP(n14422), .ZN(n14421) );
  NAND2X0 U14871 ( .IN1(n14423), .IN2(n14424), .QN(n14422) );
  NOR2X0 U14872 ( .IN1(n14424), .IN2(n14423), .QN(n14420) );
  NAND2X0 U14873 ( .IN1(n14425), .IN2(n14426), .QN(n14423) );
  NAND2X0 U14874 ( .IN1(n9128), .IN2(n14427), .QN(n14426) );
  INVX0 U14875 ( .INP(n14428), .ZN(n14425) );
  NOR2X0 U14876 ( .IN1(n14427), .IN2(n9128), .QN(n14428) );
  NOR2X0 U14877 ( .IN1(n14429), .IN2(n14430), .QN(n14427) );
  INVX0 U14878 ( .INP(n14431), .ZN(n14430) );
  NAND2X0 U14879 ( .IN1(n18414), .IN2(WX7306), .QN(n14431) );
  NOR2X0 U14880 ( .IN1(WX7306), .IN2(n18414), .QN(n14429) );
  NOR2X0 U14881 ( .IN1(n14432), .IN2(n14433), .QN(n14424) );
  INVX0 U14882 ( .INP(n14434), .ZN(n14433) );
  NAND2X0 U14883 ( .IN1(n9127), .IN2(n10018), .QN(n14434) );
  NOR2X0 U14884 ( .IN1(n10007), .IN2(n9127), .QN(n14432) );
  NOR2X0 U14885 ( .IN1(n14435), .IN2(n14436), .QN(n14415) );
  NOR2X0 U14886 ( .IN1(DFF_957_n1), .IN2(n9975), .QN(n14436) );
  NOR2X0 U14887 ( .IN1(n9988), .IN2(n11303), .QN(n14435) );
  NAND2X0 U14888 ( .IN1(n10207), .IN2(n8527), .QN(n11303) );
  NAND2X0 U14889 ( .IN1(n14437), .IN2(n14438), .QN(WX5818) );
  NOR2X0 U14890 ( .IN1(n14439), .IN2(n14440), .QN(n14438) );
  NOR2X0 U14891 ( .IN1(n14441), .IN2(n9940), .QN(n14440) );
  NOR2X0 U14892 ( .IN1(n13608), .IN2(n9920), .QN(n14439) );
  NOR2X0 U14893 ( .IN1(n14442), .IN2(n14443), .QN(n13608) );
  INVX0 U14894 ( .INP(n14444), .ZN(n14443) );
  NAND2X0 U14895 ( .IN1(n14445), .IN2(n14446), .QN(n14444) );
  NOR2X0 U14896 ( .IN1(n14446), .IN2(n14445), .QN(n14442) );
  NAND2X0 U14897 ( .IN1(n14447), .IN2(n14448), .QN(n14445) );
  NAND2X0 U14898 ( .IN1(n9130), .IN2(n14449), .QN(n14448) );
  INVX0 U14899 ( .INP(n14450), .ZN(n14447) );
  NOR2X0 U14900 ( .IN1(n14449), .IN2(n9130), .QN(n14450) );
  NOR2X0 U14901 ( .IN1(n14451), .IN2(n14452), .QN(n14449) );
  INVX0 U14902 ( .INP(n14453), .ZN(n14452) );
  NAND2X0 U14903 ( .IN1(n18413), .IN2(WX7304), .QN(n14453) );
  NOR2X0 U14904 ( .IN1(WX7304), .IN2(n18413), .QN(n14451) );
  NOR2X0 U14905 ( .IN1(n14454), .IN2(n14455), .QN(n14446) );
  INVX0 U14906 ( .INP(n14456), .ZN(n14455) );
  NAND2X0 U14907 ( .IN1(n9129), .IN2(n10018), .QN(n14456) );
  NOR2X0 U14908 ( .IN1(n10007), .IN2(n9129), .QN(n14454) );
  NOR2X0 U14909 ( .IN1(n14457), .IN2(n14458), .QN(n14437) );
  NOR2X0 U14910 ( .IN1(DFF_958_n1), .IN2(n9974), .QN(n14458) );
  NOR2X0 U14911 ( .IN1(n9988), .IN2(n11304), .QN(n14457) );
  NAND2X0 U14912 ( .IN1(n10207), .IN2(n8528), .QN(n11304) );
  NAND2X0 U14913 ( .IN1(n14459), .IN2(n14460), .QN(WX5816) );
  NOR2X0 U14914 ( .IN1(n14461), .IN2(n14462), .QN(n14460) );
  NOR2X0 U14915 ( .IN1(n14463), .IN2(n9940), .QN(n14462) );
  NOR2X0 U14916 ( .IN1(n13630), .IN2(n9921), .QN(n14461) );
  NOR2X0 U14917 ( .IN1(n14464), .IN2(n14465), .QN(n13630) );
  INVX0 U14918 ( .INP(n14466), .ZN(n14465) );
  NAND2X0 U14919 ( .IN1(n14467), .IN2(n14468), .QN(n14466) );
  NOR2X0 U14920 ( .IN1(n14468), .IN2(n14467), .QN(n14464) );
  NAND2X0 U14921 ( .IN1(n14469), .IN2(n14470), .QN(n14467) );
  NAND2X0 U14922 ( .IN1(n9010), .IN2(n14471), .QN(n14470) );
  INVX0 U14923 ( .INP(n14472), .ZN(n14469) );
  NOR2X0 U14924 ( .IN1(n14471), .IN2(n9010), .QN(n14472) );
  NOR2X0 U14925 ( .IN1(n14473), .IN2(n14474), .QN(n14471) );
  INVX0 U14926 ( .INP(n14475), .ZN(n14474) );
  NAND2X0 U14927 ( .IN1(n18412), .IN2(WX7302), .QN(n14475) );
  NOR2X0 U14928 ( .IN1(WX7302), .IN2(n18412), .QN(n14473) );
  NOR2X0 U14929 ( .IN1(n14476), .IN2(n14477), .QN(n14468) );
  INVX0 U14930 ( .INP(n14478), .ZN(n14477) );
  NAND2X0 U14931 ( .IN1(n9009), .IN2(n10018), .QN(n14478) );
  NOR2X0 U14932 ( .IN1(n10008), .IN2(n9009), .QN(n14476) );
  NOR2X0 U14933 ( .IN1(n14479), .IN2(n14480), .QN(n14459) );
  NOR2X0 U14934 ( .IN1(n9492), .IN2(n11994), .QN(n14480) );
  NOR2X0 U14935 ( .IN1(DFF_959_n1), .IN2(n9973), .QN(n14479) );
  INVX0 U14936 ( .INP(n14481), .ZN(WX5718) );
  NAND2X0 U14937 ( .IN1(n10207), .IN2(n9492), .QN(n14481) );
  NOR2X0 U14938 ( .IN1(n10328), .IN2(n14482), .QN(WX5205) );
  NAND2X0 U14939 ( .IN1(n14483), .IN2(n14484), .QN(n14482) );
  INVX0 U14940 ( .INP(n14485), .ZN(n14484) );
  NOR2X0 U14941 ( .IN1(WX4716), .IN2(DFF_766_n1), .QN(n14485) );
  NAND2X0 U14942 ( .IN1(DFF_766_n1), .IN2(WX4716), .QN(n14483) );
  NOR2X0 U14943 ( .IN1(n10329), .IN2(n14486), .QN(WX5203) );
  NAND2X0 U14944 ( .IN1(n14487), .IN2(n14488), .QN(n14486) );
  INVX0 U14945 ( .INP(n14489), .ZN(n14488) );
  NOR2X0 U14946 ( .IN1(WX4718), .IN2(DFF_765_n1), .QN(n14489) );
  NAND2X0 U14947 ( .IN1(DFF_765_n1), .IN2(WX4718), .QN(n14487) );
  NOR2X0 U14948 ( .IN1(n10329), .IN2(n14490), .QN(WX5201) );
  NAND2X0 U14949 ( .IN1(n14491), .IN2(n14492), .QN(n14490) );
  INVX0 U14950 ( .INP(n14493), .ZN(n14492) );
  NOR2X0 U14951 ( .IN1(WX4720), .IN2(DFF_764_n1), .QN(n14493) );
  NAND2X0 U14952 ( .IN1(DFF_764_n1), .IN2(WX4720), .QN(n14491) );
  NOR2X0 U14953 ( .IN1(n10329), .IN2(n14494), .QN(WX5199) );
  NOR2X0 U14954 ( .IN1(n14495), .IN2(n14496), .QN(n14494) );
  INVX0 U14955 ( .INP(n14497), .ZN(n14496) );
  NAND2X0 U14956 ( .IN1(n9830), .IN2(DFF_763_n1), .QN(n14497) );
  NOR2X0 U14957 ( .IN1(DFF_763_n1), .IN2(n9830), .QN(n14495) );
  NOR2X0 U14958 ( .IN1(n10329), .IN2(n14498), .QN(WX5197) );
  NAND2X0 U14959 ( .IN1(n14499), .IN2(n14500), .QN(n14498) );
  INVX0 U14960 ( .INP(n14501), .ZN(n14500) );
  NOR2X0 U14961 ( .IN1(WX4724), .IN2(DFF_762_n1), .QN(n14501) );
  NAND2X0 U14962 ( .IN1(DFF_762_n1), .IN2(WX4724), .QN(n14499) );
  NOR2X0 U14963 ( .IN1(n10329), .IN2(n14502), .QN(WX5195) );
  NAND2X0 U14964 ( .IN1(n14503), .IN2(n14504), .QN(n14502) );
  INVX0 U14965 ( .INP(n14505), .ZN(n14504) );
  NOR2X0 U14966 ( .IN1(WX4726), .IN2(DFF_761_n1), .QN(n14505) );
  NAND2X0 U14967 ( .IN1(DFF_761_n1), .IN2(WX4726), .QN(n14503) );
  NOR2X0 U14968 ( .IN1(n10329), .IN2(n14506), .QN(WX5193) );
  NAND2X0 U14969 ( .IN1(n14507), .IN2(n14508), .QN(n14506) );
  INVX0 U14970 ( .INP(n14509), .ZN(n14508) );
  NOR2X0 U14971 ( .IN1(WX4728), .IN2(DFF_760_n1), .QN(n14509) );
  NAND2X0 U14972 ( .IN1(DFF_760_n1), .IN2(WX4728), .QN(n14507) );
  NOR2X0 U14973 ( .IN1(n10329), .IN2(n14510), .QN(WX5191) );
  NAND2X0 U14974 ( .IN1(n14511), .IN2(n14512), .QN(n14510) );
  INVX0 U14975 ( .INP(n14513), .ZN(n14512) );
  NOR2X0 U14976 ( .IN1(WX4730), .IN2(DFF_759_n1), .QN(n14513) );
  NAND2X0 U14977 ( .IN1(DFF_759_n1), .IN2(WX4730), .QN(n14511) );
  NOR2X0 U14978 ( .IN1(n10329), .IN2(n14514), .QN(WX5189) );
  NOR2X0 U14979 ( .IN1(n14515), .IN2(n14516), .QN(n14514) );
  NOR2X0 U14980 ( .IN1(test_so43), .IN2(WX4732), .QN(n14516) );
  NOR2X0 U14981 ( .IN1(n9665), .IN2(n9859), .QN(n14515) );
  NOR2X0 U14982 ( .IN1(n10329), .IN2(n14517), .QN(WX5187) );
  NAND2X0 U14983 ( .IN1(n14518), .IN2(n14519), .QN(n14517) );
  INVX0 U14984 ( .INP(n14520), .ZN(n14519) );
  NOR2X0 U14985 ( .IN1(WX4734), .IN2(DFF_757_n1), .QN(n14520) );
  NAND2X0 U14986 ( .IN1(DFF_757_n1), .IN2(WX4734), .QN(n14518) );
  NOR2X0 U14987 ( .IN1(n10329), .IN2(n14521), .QN(WX5185) );
  NAND2X0 U14988 ( .IN1(n14522), .IN2(n14523), .QN(n14521) );
  INVX0 U14989 ( .INP(n14524), .ZN(n14523) );
  NOR2X0 U14990 ( .IN1(WX4736), .IN2(DFF_756_n1), .QN(n14524) );
  NAND2X0 U14991 ( .IN1(DFF_756_n1), .IN2(WX4736), .QN(n14522) );
  NOR2X0 U14992 ( .IN1(n10329), .IN2(n14525), .QN(WX5183) );
  NAND2X0 U14993 ( .IN1(n14526), .IN2(n14527), .QN(n14525) );
  INVX0 U14994 ( .INP(n14528), .ZN(n14527) );
  NOR2X0 U14995 ( .IN1(WX4738), .IN2(DFF_755_n1), .QN(n14528) );
  NAND2X0 U14996 ( .IN1(DFF_755_n1), .IN2(WX4738), .QN(n14526) );
  NOR2X0 U14997 ( .IN1(n10329), .IN2(n14529), .QN(WX5181) );
  NAND2X0 U14998 ( .IN1(n14530), .IN2(n14531), .QN(n14529) );
  INVX0 U14999 ( .INP(n14532), .ZN(n14531) );
  NOR2X0 U15000 ( .IN1(WX4740), .IN2(DFF_754_n1), .QN(n14532) );
  NAND2X0 U15001 ( .IN1(DFF_754_n1), .IN2(WX4740), .QN(n14530) );
  NOR2X0 U15002 ( .IN1(n10329), .IN2(n14533), .QN(WX5179) );
  NAND2X0 U15003 ( .IN1(n14534), .IN2(n14535), .QN(n14533) );
  INVX0 U15004 ( .INP(n14536), .ZN(n14535) );
  NOR2X0 U15005 ( .IN1(WX4742), .IN2(DFF_753_n1), .QN(n14536) );
  NAND2X0 U15006 ( .IN1(DFF_753_n1), .IN2(WX4742), .QN(n14534) );
  NOR2X0 U15007 ( .IN1(n10330), .IN2(n14537), .QN(WX5177) );
  NAND2X0 U15008 ( .IN1(n14538), .IN2(n14539), .QN(n14537) );
  INVX0 U15009 ( .INP(n14540), .ZN(n14539) );
  NOR2X0 U15010 ( .IN1(WX4744), .IN2(DFF_752_n1), .QN(n14540) );
  NAND2X0 U15011 ( .IN1(DFF_752_n1), .IN2(WX4744), .QN(n14538) );
  NOR2X0 U15012 ( .IN1(n10330), .IN2(n14541), .QN(WX5175) );
  NOR2X0 U15013 ( .IN1(n14542), .IN2(n14543), .QN(n14541) );
  INVX0 U15014 ( .INP(n14544), .ZN(n14543) );
  NAND2X0 U15015 ( .IN1(CRC_OUT_6_15), .IN2(n14545), .QN(n14544) );
  NOR2X0 U15016 ( .IN1(n14545), .IN2(CRC_OUT_6_15), .QN(n14542) );
  NAND2X0 U15017 ( .IN1(n14546), .IN2(n14547), .QN(n14545) );
  NAND2X0 U15018 ( .IN1(n9509), .IN2(CRC_OUT_6_31), .QN(n14547) );
  NAND2X0 U15019 ( .IN1(DFF_767_n1), .IN2(WX4746), .QN(n14546) );
  NOR2X0 U15020 ( .IN1(n10330), .IN2(n14548), .QN(WX5173) );
  NAND2X0 U15021 ( .IN1(n14549), .IN2(n14550), .QN(n14548) );
  INVX0 U15022 ( .INP(n14551), .ZN(n14550) );
  NOR2X0 U15023 ( .IN1(WX4748), .IN2(DFF_750_n1), .QN(n14551) );
  NAND2X0 U15024 ( .IN1(DFF_750_n1), .IN2(WX4748), .QN(n14549) );
  NOR2X0 U15025 ( .IN1(n10330), .IN2(n14552), .QN(WX5171) );
  NAND2X0 U15026 ( .IN1(n14553), .IN2(n14554), .QN(n14552) );
  INVX0 U15027 ( .INP(n14555), .ZN(n14554) );
  NOR2X0 U15028 ( .IN1(WX4750), .IN2(DFF_749_n1), .QN(n14555) );
  NAND2X0 U15029 ( .IN1(DFF_749_n1), .IN2(WX4750), .QN(n14553) );
  NOR2X0 U15030 ( .IN1(n10330), .IN2(n14556), .QN(WX5169) );
  NAND2X0 U15031 ( .IN1(n14557), .IN2(n14558), .QN(n14556) );
  INVX0 U15032 ( .INP(n14559), .ZN(n14558) );
  NOR2X0 U15033 ( .IN1(WX4752), .IN2(DFF_748_n1), .QN(n14559) );
  NAND2X0 U15034 ( .IN1(DFF_748_n1), .IN2(WX4752), .QN(n14557) );
  NOR2X0 U15035 ( .IN1(n10330), .IN2(n14560), .QN(WX5167) );
  NAND2X0 U15036 ( .IN1(n14561), .IN2(n14562), .QN(n14560) );
  INVX0 U15037 ( .INP(n14563), .ZN(n14562) );
  NOR2X0 U15038 ( .IN1(WX4754), .IN2(DFF_747_n1), .QN(n14563) );
  NAND2X0 U15039 ( .IN1(DFF_747_n1), .IN2(WX4754), .QN(n14561) );
  NOR2X0 U15040 ( .IN1(n10330), .IN2(n14564), .QN(WX5165) );
  NAND2X0 U15041 ( .IN1(n14565), .IN2(n14566), .QN(n14564) );
  INVX0 U15042 ( .INP(n14567), .ZN(n14566) );
  NOR2X0 U15043 ( .IN1(CRC_OUT_6_10), .IN2(n14568), .QN(n14567) );
  NAND2X0 U15044 ( .IN1(n14568), .IN2(CRC_OUT_6_10), .QN(n14565) );
  NAND2X0 U15045 ( .IN1(n14569), .IN2(n14570), .QN(n14568) );
  NAND2X0 U15046 ( .IN1(test_so41), .IN2(CRC_OUT_6_31), .QN(n14570) );
  NAND2X0 U15047 ( .IN1(DFF_767_n1), .IN2(n9850), .QN(n14569) );
  NOR2X0 U15048 ( .IN1(n10330), .IN2(n14571), .QN(WX5163) );
  NAND2X0 U15049 ( .IN1(n14572), .IN2(n14573), .QN(n14571) );
  INVX0 U15050 ( .INP(n14574), .ZN(n14573) );
  NOR2X0 U15051 ( .IN1(WX4758), .IN2(DFF_745_n1), .QN(n14574) );
  NAND2X0 U15052 ( .IN1(DFF_745_n1), .IN2(WX4758), .QN(n14572) );
  NOR2X0 U15053 ( .IN1(n10330), .IN2(n14575), .QN(WX5161) );
  NAND2X0 U15054 ( .IN1(n14576), .IN2(n14577), .QN(n14575) );
  INVX0 U15055 ( .INP(n14578), .ZN(n14577) );
  NOR2X0 U15056 ( .IN1(WX4760), .IN2(DFF_744_n1), .QN(n14578) );
  NAND2X0 U15057 ( .IN1(DFF_744_n1), .IN2(WX4760), .QN(n14576) );
  NOR2X0 U15058 ( .IN1(n10330), .IN2(n14579), .QN(WX5159) );
  NAND2X0 U15059 ( .IN1(n14580), .IN2(n14581), .QN(n14579) );
  INVX0 U15060 ( .INP(n14582), .ZN(n14581) );
  NOR2X0 U15061 ( .IN1(WX4762), .IN2(DFF_743_n1), .QN(n14582) );
  NAND2X0 U15062 ( .IN1(DFF_743_n1), .IN2(WX4762), .QN(n14580) );
  NOR2X0 U15063 ( .IN1(n10330), .IN2(n14583), .QN(WX5157) );
  NAND2X0 U15064 ( .IN1(n14584), .IN2(n14585), .QN(n14583) );
  INVX0 U15065 ( .INP(n14586), .ZN(n14585) );
  NOR2X0 U15066 ( .IN1(WX4764), .IN2(DFF_742_n1), .QN(n14586) );
  NAND2X0 U15067 ( .IN1(DFF_742_n1), .IN2(WX4764), .QN(n14584) );
  NOR2X0 U15068 ( .IN1(n10330), .IN2(n14587), .QN(WX5155) );
  NOR2X0 U15069 ( .IN1(n14588), .IN2(n14589), .QN(n14587) );
  NOR2X0 U15070 ( .IN1(test_so42), .IN2(WX4766), .QN(n14589) );
  NOR2X0 U15071 ( .IN1(n9680), .IN2(n9858), .QN(n14588) );
  NOR2X0 U15072 ( .IN1(n10330), .IN2(n14590), .QN(WX5153) );
  NAND2X0 U15073 ( .IN1(n14591), .IN2(n14592), .QN(n14590) );
  INVX0 U15074 ( .INP(n14593), .ZN(n14592) );
  NOR2X0 U15075 ( .IN1(WX4768), .IN2(DFF_740_n1), .QN(n14593) );
  NAND2X0 U15076 ( .IN1(DFF_740_n1), .IN2(WX4768), .QN(n14591) );
  NOR2X0 U15077 ( .IN1(n10331), .IN2(n14594), .QN(WX5151) );
  NOR2X0 U15078 ( .IN1(n14595), .IN2(n14596), .QN(n14594) );
  INVX0 U15079 ( .INP(n14597), .ZN(n14596) );
  NAND2X0 U15080 ( .IN1(CRC_OUT_6_3), .IN2(n14598), .QN(n14597) );
  NOR2X0 U15081 ( .IN1(n14598), .IN2(CRC_OUT_6_3), .QN(n14595) );
  NAND2X0 U15082 ( .IN1(n14599), .IN2(n14600), .QN(n14598) );
  NAND2X0 U15083 ( .IN1(n9510), .IN2(CRC_OUT_6_31), .QN(n14600) );
  NAND2X0 U15084 ( .IN1(DFF_767_n1), .IN2(WX4770), .QN(n14599) );
  NOR2X0 U15085 ( .IN1(n10331), .IN2(n14601), .QN(WX5149) );
  NAND2X0 U15086 ( .IN1(n14602), .IN2(n14603), .QN(n14601) );
  INVX0 U15087 ( .INP(n14604), .ZN(n14603) );
  NOR2X0 U15088 ( .IN1(WX4772), .IN2(DFF_738_n1), .QN(n14604) );
  NAND2X0 U15089 ( .IN1(DFF_738_n1), .IN2(WX4772), .QN(n14602) );
  NOR2X0 U15090 ( .IN1(n10331), .IN2(n14605), .QN(WX5147) );
  NAND2X0 U15091 ( .IN1(n14606), .IN2(n14607), .QN(n14605) );
  INVX0 U15092 ( .INP(n14608), .ZN(n14607) );
  NOR2X0 U15093 ( .IN1(WX4774), .IN2(DFF_737_n1), .QN(n14608) );
  NAND2X0 U15094 ( .IN1(DFF_737_n1), .IN2(WX4774), .QN(n14606) );
  NOR2X0 U15095 ( .IN1(n10331), .IN2(n14609), .QN(WX5145) );
  NAND2X0 U15096 ( .IN1(n14610), .IN2(n14611), .QN(n14609) );
  INVX0 U15097 ( .INP(n14612), .ZN(n14611) );
  NOR2X0 U15098 ( .IN1(WX4776), .IN2(DFF_736_n1), .QN(n14612) );
  NAND2X0 U15099 ( .IN1(DFF_736_n1), .IN2(WX4776), .QN(n14610) );
  NOR2X0 U15100 ( .IN1(n10331), .IN2(n14613), .QN(WX5143) );
  NAND2X0 U15101 ( .IN1(n14614), .IN2(n14615), .QN(n14613) );
  NAND2X0 U15102 ( .IN1(n9522), .IN2(CRC_OUT_6_31), .QN(n14615) );
  NAND2X0 U15103 ( .IN1(DFF_767_n1), .IN2(WX4778), .QN(n14614) );
  NOR2X0 U15104 ( .IN1(n18396), .IN2(n10292), .QN(WX4617) );
  NOR2X0 U15105 ( .IN1(n10331), .IN2(n9843), .QN(WX4615) );
  NOR2X0 U15106 ( .IN1(n18395), .IN2(n10291), .QN(WX4613) );
  NOR2X0 U15107 ( .IN1(n18394), .IN2(n10306), .QN(WX4611) );
  NOR2X0 U15108 ( .IN1(n18393), .IN2(n10243), .QN(WX4609) );
  NOR2X0 U15109 ( .IN1(n18392), .IN2(n10243), .QN(WX4607) );
  NOR2X0 U15110 ( .IN1(n18391), .IN2(n10243), .QN(WX4605) );
  NOR2X0 U15111 ( .IN1(n18390), .IN2(n10243), .QN(WX4603) );
  NOR2X0 U15112 ( .IN1(n18389), .IN2(n10243), .QN(WX4601) );
  NOR2X0 U15113 ( .IN1(n18388), .IN2(n10243), .QN(WX4599) );
  NOR2X0 U15114 ( .IN1(n18387), .IN2(n10243), .QN(WX4597) );
  NOR2X0 U15115 ( .IN1(n18386), .IN2(n10243), .QN(WX4595) );
  NOR2X0 U15116 ( .IN1(n18385), .IN2(n10243), .QN(WX4593) );
  NOR2X0 U15117 ( .IN1(n18384), .IN2(n10243), .QN(WX4591) );
  NOR2X0 U15118 ( .IN1(n18383), .IN2(n10243), .QN(WX4589) );
  NOR2X0 U15119 ( .IN1(n18382), .IN2(n10243), .QN(WX4587) );
  NAND2X0 U15120 ( .IN1(n14616), .IN2(n14617), .QN(WX4585) );
  NOR2X0 U15121 ( .IN1(n14618), .IN2(n14619), .QN(n14617) );
  NOR2X0 U15122 ( .IN1(n9943), .IN2(n14620), .QN(n14619) );
  NOR2X0 U15123 ( .IN1(n13795), .IN2(n9921), .QN(n14618) );
  INVX0 U15124 ( .INP(n14621), .ZN(n13795) );
  NAND2X0 U15125 ( .IN1(n14622), .IN2(n14623), .QN(n14621) );
  NAND2X0 U15126 ( .IN1(n14624), .IN2(n14625), .QN(n14623) );
  NAND2X0 U15127 ( .IN1(n14626), .IN2(n14627), .QN(n14625) );
  NAND2X0 U15128 ( .IN1(n9367), .IN2(WX5879), .QN(n14627) );
  NAND2X0 U15129 ( .IN1(n9366), .IN2(WX6007), .QN(n14626) );
  NOR2X0 U15130 ( .IN1(n14628), .IN2(n14629), .QN(n14624) );
  NOR2X0 U15131 ( .IN1(n9521), .IN2(WX5943), .QN(n14629) );
  NOR2X0 U15132 ( .IN1(n3659), .IN2(WX6071), .QN(n14628) );
  NAND2X0 U15133 ( .IN1(n14630), .IN2(n14631), .QN(n14622) );
  NAND2X0 U15134 ( .IN1(n14632), .IN2(n14633), .QN(n14631) );
  NAND2X0 U15135 ( .IN1(n9521), .IN2(WX5943), .QN(n14633) );
  NAND2X0 U15136 ( .IN1(n3659), .IN2(WX6071), .QN(n14632) );
  NOR2X0 U15137 ( .IN1(n14634), .IN2(n14635), .QN(n14630) );
  NOR2X0 U15138 ( .IN1(n9367), .IN2(WX5879), .QN(n14635) );
  NOR2X0 U15139 ( .IN1(n9366), .IN2(WX6007), .QN(n14634) );
  NOR2X0 U15140 ( .IN1(n14636), .IN2(n14637), .QN(n14616) );
  NOR2X0 U15141 ( .IN1(DFF_736_n1), .IN2(n9974), .QN(n14637) );
  NOR2X0 U15142 ( .IN1(n9988), .IN2(n10568), .QN(n14636) );
  NAND2X0 U15143 ( .IN1(n10207), .IN2(n8554), .QN(n10568) );
  NAND2X0 U15144 ( .IN1(n14638), .IN2(n14639), .QN(WX4583) );
  NOR2X0 U15145 ( .IN1(n14640), .IN2(n14641), .QN(n14639) );
  NOR2X0 U15146 ( .IN1(n14642), .IN2(n10563), .QN(n14641) );
  NOR2X0 U15147 ( .IN1(n9924), .IN2(n13817), .QN(n14640) );
  NAND2X0 U15148 ( .IN1(n14643), .IN2(n14644), .QN(n13817) );
  INVX0 U15149 ( .INP(n14645), .ZN(n14644) );
  NOR2X0 U15150 ( .IN1(n14646), .IN2(n14647), .QN(n14645) );
  NAND2X0 U15151 ( .IN1(n14647), .IN2(n14646), .QN(n14643) );
  NOR2X0 U15152 ( .IN1(n14648), .IN2(n14649), .QN(n14646) );
  INVX0 U15153 ( .INP(n14650), .ZN(n14649) );
  NAND2X0 U15154 ( .IN1(test_so51), .IN2(WX6069), .QN(n14650) );
  NOR2X0 U15155 ( .IN1(WX6069), .IN2(test_so51), .QN(n14648) );
  NAND2X0 U15156 ( .IN1(n14651), .IN2(n14652), .QN(n14647) );
  NAND2X0 U15157 ( .IN1(n9368), .IN2(WX5941), .QN(n14652) );
  INVX0 U15158 ( .INP(n14653), .ZN(n14651) );
  NOR2X0 U15159 ( .IN1(WX5941), .IN2(n9368), .QN(n14653) );
  NOR2X0 U15160 ( .IN1(n14654), .IN2(n14655), .QN(n14638) );
  NOR2X0 U15161 ( .IN1(DFF_737_n1), .IN2(n9974), .QN(n14655) );
  NOR2X0 U15162 ( .IN1(n9988), .IN2(n10569), .QN(n14654) );
  NAND2X0 U15163 ( .IN1(n10207), .IN2(n8555), .QN(n10569) );
  NAND2X0 U15164 ( .IN1(n14656), .IN2(n14657), .QN(WX4581) );
  NOR2X0 U15165 ( .IN1(n14658), .IN2(n14659), .QN(n14657) );
  NOR2X0 U15166 ( .IN1(n14660), .IN2(n9940), .QN(n14659) );
  NOR2X0 U15167 ( .IN1(n13839), .IN2(n9920), .QN(n14658) );
  INVX0 U15168 ( .INP(n14661), .ZN(n13839) );
  NAND2X0 U15169 ( .IN1(n14662), .IN2(n14663), .QN(n14661) );
  NAND2X0 U15170 ( .IN1(n14664), .IN2(n14665), .QN(n14663) );
  NAND2X0 U15171 ( .IN1(n14666), .IN2(n14667), .QN(n14665) );
  NAND2X0 U15172 ( .IN1(n9370), .IN2(WX5875), .QN(n14667) );
  NAND2X0 U15173 ( .IN1(n9369), .IN2(WX6003), .QN(n14666) );
  NOR2X0 U15174 ( .IN1(n14668), .IN2(n14669), .QN(n14664) );
  NOR2X0 U15175 ( .IN1(n9656), .IN2(WX5939), .QN(n14669) );
  NOR2X0 U15176 ( .IN1(n3663), .IN2(WX6067), .QN(n14668) );
  NAND2X0 U15177 ( .IN1(n14670), .IN2(n14671), .QN(n14662) );
  NAND2X0 U15178 ( .IN1(n14672), .IN2(n14673), .QN(n14671) );
  NAND2X0 U15179 ( .IN1(n9656), .IN2(WX5939), .QN(n14673) );
  NAND2X0 U15180 ( .IN1(n3663), .IN2(WX6067), .QN(n14672) );
  NOR2X0 U15181 ( .IN1(n14674), .IN2(n14675), .QN(n14670) );
  NOR2X0 U15182 ( .IN1(n9370), .IN2(WX5875), .QN(n14675) );
  NOR2X0 U15183 ( .IN1(n9369), .IN2(WX6003), .QN(n14674) );
  NOR2X0 U15184 ( .IN1(n14676), .IN2(n14677), .QN(n14656) );
  NOR2X0 U15185 ( .IN1(DFF_738_n1), .IN2(n9974), .QN(n14677) );
  NOR2X0 U15186 ( .IN1(n9988), .IN2(n10570), .QN(n14676) );
  NAND2X0 U15187 ( .IN1(test_so34), .IN2(n10214), .QN(n10570) );
  NAND2X0 U15188 ( .IN1(n14678), .IN2(n14679), .QN(WX4579) );
  NOR2X0 U15189 ( .IN1(n14680), .IN2(n14681), .QN(n14679) );
  NOR2X0 U15190 ( .IN1(n14682), .IN2(n9940), .QN(n14681) );
  NOR2X0 U15191 ( .IN1(n9924), .IN2(n13861), .QN(n14680) );
  NAND2X0 U15192 ( .IN1(n14683), .IN2(n14684), .QN(n13861) );
  INVX0 U15193 ( .INP(n14685), .ZN(n14684) );
  NOR2X0 U15194 ( .IN1(n14686), .IN2(n14687), .QN(n14685) );
  NAND2X0 U15195 ( .IN1(n14687), .IN2(n14686), .QN(n14683) );
  NOR2X0 U15196 ( .IN1(n14688), .IN2(n14689), .QN(n14686) );
  INVX0 U15197 ( .INP(n14690), .ZN(n14689) );
  NAND2X0 U15198 ( .IN1(test_so49), .IN2(WX6065), .QN(n14690) );
  NOR2X0 U15199 ( .IN1(WX6065), .IN2(test_so49), .QN(n14688) );
  NAND2X0 U15200 ( .IN1(n14691), .IN2(n14692), .QN(n14687) );
  NAND2X0 U15201 ( .IN1(n9372), .IN2(WX5873), .QN(n14692) );
  INVX0 U15202 ( .INP(n14693), .ZN(n14691) );
  NOR2X0 U15203 ( .IN1(WX5873), .IN2(n9372), .QN(n14693) );
  NOR2X0 U15204 ( .IN1(n14694), .IN2(n14695), .QN(n14678) );
  NOR2X0 U15205 ( .IN1(DFF_739_n1), .IN2(n9973), .QN(n14695) );
  NOR2X0 U15206 ( .IN1(n9988), .IN2(n10571), .QN(n14694) );
  NAND2X0 U15207 ( .IN1(n10207), .IN2(n8558), .QN(n10571) );
  NAND2X0 U15208 ( .IN1(n14696), .IN2(n14697), .QN(WX4577) );
  NOR2X0 U15209 ( .IN1(n14698), .IN2(n14699), .QN(n14697) );
  NOR2X0 U15210 ( .IN1(n14700), .IN2(n9940), .QN(n14699) );
  NOR2X0 U15211 ( .IN1(n13883), .IN2(n9920), .QN(n14698) );
  INVX0 U15212 ( .INP(n14701), .ZN(n13883) );
  NAND2X0 U15213 ( .IN1(n14702), .IN2(n14703), .QN(n14701) );
  NAND2X0 U15214 ( .IN1(n14704), .IN2(n14705), .QN(n14703) );
  NAND2X0 U15215 ( .IN1(n14706), .IN2(n14707), .QN(n14705) );
  NAND2X0 U15216 ( .IN1(n9374), .IN2(WX5871), .QN(n14707) );
  NAND2X0 U15217 ( .IN1(n9373), .IN2(WX5999), .QN(n14706) );
  NOR2X0 U15218 ( .IN1(n14708), .IN2(n14709), .QN(n14704) );
  NOR2X0 U15219 ( .IN1(n9508), .IN2(WX5935), .QN(n14709) );
  NOR2X0 U15220 ( .IN1(n3667), .IN2(WX6063), .QN(n14708) );
  NAND2X0 U15221 ( .IN1(n14710), .IN2(n14711), .QN(n14702) );
  NAND2X0 U15222 ( .IN1(n14712), .IN2(n14713), .QN(n14711) );
  NAND2X0 U15223 ( .IN1(n9508), .IN2(WX5935), .QN(n14713) );
  NAND2X0 U15224 ( .IN1(n3667), .IN2(WX6063), .QN(n14712) );
  NOR2X0 U15225 ( .IN1(n14714), .IN2(n14715), .QN(n14710) );
  NOR2X0 U15226 ( .IN1(n9374), .IN2(WX5871), .QN(n14715) );
  NOR2X0 U15227 ( .IN1(n9373), .IN2(WX5999), .QN(n14714) );
  NOR2X0 U15228 ( .IN1(n14716), .IN2(n14717), .QN(n14696) );
  NOR2X0 U15229 ( .IN1(DFF_740_n1), .IN2(n9974), .QN(n14717) );
  NOR2X0 U15230 ( .IN1(n9988), .IN2(n10572), .QN(n14716) );
  NAND2X0 U15231 ( .IN1(n10207), .IN2(n8559), .QN(n10572) );
  NAND2X0 U15232 ( .IN1(n14718), .IN2(n14719), .QN(WX4575) );
  NOR2X0 U15233 ( .IN1(n14720), .IN2(n14721), .QN(n14719) );
  NOR2X0 U15234 ( .IN1(n14722), .IN2(n9940), .QN(n14721) );
  NOR2X0 U15235 ( .IN1(n9923), .IN2(n13901), .QN(n14720) );
  NAND2X0 U15236 ( .IN1(n14723), .IN2(n14724), .QN(n13901) );
  INVX0 U15237 ( .INP(n14725), .ZN(n14724) );
  NOR2X0 U15238 ( .IN1(n14726), .IN2(n14727), .QN(n14725) );
  NAND2X0 U15239 ( .IN1(n14727), .IN2(n14726), .QN(n14723) );
  NOR2X0 U15240 ( .IN1(n14728), .IN2(n14729), .QN(n14726) );
  INVX0 U15241 ( .INP(n14730), .ZN(n14729) );
  NAND2X0 U15242 ( .IN1(test_so47), .IN2(WX6061), .QN(n14730) );
  NOR2X0 U15243 ( .IN1(WX6061), .IN2(test_so47), .QN(n14728) );
  NAND2X0 U15244 ( .IN1(n14731), .IN2(n14732), .QN(n14727) );
  NAND2X0 U15245 ( .IN1(n9375), .IN2(WX5933), .QN(n14732) );
  INVX0 U15246 ( .INP(n14733), .ZN(n14731) );
  NOR2X0 U15247 ( .IN1(WX5933), .IN2(n9375), .QN(n14733) );
  NOR2X0 U15248 ( .IN1(n14734), .IN2(n14735), .QN(n14718) );
  NOR2X0 U15249 ( .IN1(n9975), .IN2(n9858), .QN(n14735) );
  NOR2X0 U15250 ( .IN1(n9988), .IN2(n10573), .QN(n14734) );
  NAND2X0 U15251 ( .IN1(n10206), .IN2(n8560), .QN(n10573) );
  NAND2X0 U15252 ( .IN1(n14736), .IN2(n14737), .QN(WX4573) );
  NOR2X0 U15253 ( .IN1(n14738), .IN2(n14739), .QN(n14737) );
  NOR2X0 U15254 ( .IN1(n14740), .IN2(n10563), .QN(n14739) );
  NOR2X0 U15255 ( .IN1(n13923), .IN2(n9920), .QN(n14738) );
  INVX0 U15256 ( .INP(n14741), .ZN(n13923) );
  NAND2X0 U15257 ( .IN1(n14742), .IN2(n14743), .QN(n14741) );
  NAND2X0 U15258 ( .IN1(n14744), .IN2(n14745), .QN(n14743) );
  NAND2X0 U15259 ( .IN1(n14746), .IN2(n14747), .QN(n14745) );
  NAND2X0 U15260 ( .IN1(n9377), .IN2(WX5867), .QN(n14747) );
  NAND2X0 U15261 ( .IN1(n9376), .IN2(WX5995), .QN(n14746) );
  NOR2X0 U15262 ( .IN1(n14748), .IN2(n14749), .QN(n14744) );
  NOR2X0 U15263 ( .IN1(n9653), .IN2(WX5931), .QN(n14749) );
  NOR2X0 U15264 ( .IN1(n3671), .IN2(WX6059), .QN(n14748) );
  NAND2X0 U15265 ( .IN1(n14750), .IN2(n14751), .QN(n14742) );
  NAND2X0 U15266 ( .IN1(n14752), .IN2(n14753), .QN(n14751) );
  NAND2X0 U15267 ( .IN1(n9653), .IN2(WX5931), .QN(n14753) );
  NAND2X0 U15268 ( .IN1(n3671), .IN2(WX6059), .QN(n14752) );
  NOR2X0 U15269 ( .IN1(n14754), .IN2(n14755), .QN(n14750) );
  NOR2X0 U15270 ( .IN1(n9377), .IN2(WX5867), .QN(n14755) );
  NOR2X0 U15271 ( .IN1(n9376), .IN2(WX5995), .QN(n14754) );
  NOR2X0 U15272 ( .IN1(n14756), .IN2(n14757), .QN(n14736) );
  NOR2X0 U15273 ( .IN1(DFF_742_n1), .IN2(n9974), .QN(n14757) );
  NOR2X0 U15274 ( .IN1(n9988), .IN2(n10574), .QN(n14756) );
  NAND2X0 U15275 ( .IN1(n10206), .IN2(n8561), .QN(n10574) );
  NAND2X0 U15276 ( .IN1(n14758), .IN2(n14759), .QN(WX4571) );
  NOR2X0 U15277 ( .IN1(n14760), .IN2(n14761), .QN(n14759) );
  NOR2X0 U15278 ( .IN1(n14762), .IN2(n9940), .QN(n14761) );
  NOR2X0 U15279 ( .IN1(n13941), .IN2(n9920), .QN(n14760) );
  INVX0 U15280 ( .INP(n14763), .ZN(n13941) );
  NAND2X0 U15281 ( .IN1(n14764), .IN2(n14765), .QN(n14763) );
  NAND2X0 U15282 ( .IN1(n14766), .IN2(n14767), .QN(n14765) );
  NAND2X0 U15283 ( .IN1(n14768), .IN2(n14769), .QN(n14767) );
  NAND2X0 U15284 ( .IN1(n9379), .IN2(WX5865), .QN(n14769) );
  NAND2X0 U15285 ( .IN1(n9378), .IN2(WX5993), .QN(n14768) );
  NOR2X0 U15286 ( .IN1(n14770), .IN2(n14771), .QN(n14766) );
  NOR2X0 U15287 ( .IN1(n9652), .IN2(WX5929), .QN(n14771) );
  NOR2X0 U15288 ( .IN1(n3673), .IN2(WX6057), .QN(n14770) );
  NAND2X0 U15289 ( .IN1(n14772), .IN2(n14773), .QN(n14764) );
  NAND2X0 U15290 ( .IN1(n14774), .IN2(n14775), .QN(n14773) );
  NAND2X0 U15291 ( .IN1(n9652), .IN2(WX5929), .QN(n14775) );
  NAND2X0 U15292 ( .IN1(n3673), .IN2(WX6057), .QN(n14774) );
  NOR2X0 U15293 ( .IN1(n14776), .IN2(n14777), .QN(n14772) );
  NOR2X0 U15294 ( .IN1(n9379), .IN2(WX5865), .QN(n14777) );
  NOR2X0 U15295 ( .IN1(n9378), .IN2(WX5993), .QN(n14776) );
  NOR2X0 U15296 ( .IN1(n14778), .IN2(n14779), .QN(n14758) );
  NOR2X0 U15297 ( .IN1(DFF_743_n1), .IN2(n9974), .QN(n14779) );
  NOR2X0 U15298 ( .IN1(n9988), .IN2(n10575), .QN(n14778) );
  NAND2X0 U15299 ( .IN1(n10206), .IN2(n8562), .QN(n10575) );
  NAND2X0 U15300 ( .IN1(n14780), .IN2(n14781), .QN(WX4569) );
  NOR2X0 U15301 ( .IN1(n14782), .IN2(n14783), .QN(n14781) );
  NOR2X0 U15302 ( .IN1(n14784), .IN2(n9939), .QN(n14783) );
  NOR2X0 U15303 ( .IN1(n13963), .IN2(n9920), .QN(n14782) );
  INVX0 U15304 ( .INP(n14785), .ZN(n13963) );
  NAND2X0 U15305 ( .IN1(n14786), .IN2(n14787), .QN(n14785) );
  NAND2X0 U15306 ( .IN1(n14788), .IN2(n14789), .QN(n14787) );
  NAND2X0 U15307 ( .IN1(n14790), .IN2(n14791), .QN(n14789) );
  NAND2X0 U15308 ( .IN1(n9381), .IN2(WX5863), .QN(n14791) );
  NAND2X0 U15309 ( .IN1(n9380), .IN2(WX5991), .QN(n14790) );
  NOR2X0 U15310 ( .IN1(n14792), .IN2(n14793), .QN(n14788) );
  NOR2X0 U15311 ( .IN1(n9651), .IN2(WX5927), .QN(n14793) );
  NOR2X0 U15312 ( .IN1(n3675), .IN2(WX6055), .QN(n14792) );
  NAND2X0 U15313 ( .IN1(n14794), .IN2(n14795), .QN(n14786) );
  NAND2X0 U15314 ( .IN1(n14796), .IN2(n14797), .QN(n14795) );
  NAND2X0 U15315 ( .IN1(n9651), .IN2(WX5927), .QN(n14797) );
  NAND2X0 U15316 ( .IN1(n3675), .IN2(WX6055), .QN(n14796) );
  NOR2X0 U15317 ( .IN1(n14798), .IN2(n14799), .QN(n14794) );
  NOR2X0 U15318 ( .IN1(n9381), .IN2(WX5863), .QN(n14799) );
  NOR2X0 U15319 ( .IN1(n9380), .IN2(WX5991), .QN(n14798) );
  NOR2X0 U15320 ( .IN1(n14800), .IN2(n14801), .QN(n14780) );
  NOR2X0 U15321 ( .IN1(DFF_744_n1), .IN2(n9972), .QN(n14801) );
  NOR2X0 U15322 ( .IN1(n9988), .IN2(n10576), .QN(n14800) );
  NAND2X0 U15323 ( .IN1(n10206), .IN2(n8563), .QN(n10576) );
  NAND2X0 U15324 ( .IN1(n14802), .IN2(n14803), .QN(WX4567) );
  NOR2X0 U15325 ( .IN1(n14804), .IN2(n14805), .QN(n14803) );
  NOR2X0 U15326 ( .IN1(n14806), .IN2(n10563), .QN(n14805) );
  NOR2X0 U15327 ( .IN1(n13981), .IN2(n9921), .QN(n14804) );
  INVX0 U15328 ( .INP(n14807), .ZN(n13981) );
  NAND2X0 U15329 ( .IN1(n14808), .IN2(n14809), .QN(n14807) );
  NAND2X0 U15330 ( .IN1(n14810), .IN2(n14811), .QN(n14809) );
  NAND2X0 U15331 ( .IN1(n14812), .IN2(n14813), .QN(n14811) );
  NAND2X0 U15332 ( .IN1(n9383), .IN2(WX5861), .QN(n14813) );
  NAND2X0 U15333 ( .IN1(n9382), .IN2(WX5989), .QN(n14812) );
  NOR2X0 U15334 ( .IN1(n14814), .IN2(n14815), .QN(n14810) );
  NOR2X0 U15335 ( .IN1(n9650), .IN2(WX5925), .QN(n14815) );
  NOR2X0 U15336 ( .IN1(n3677), .IN2(WX6053), .QN(n14814) );
  NAND2X0 U15337 ( .IN1(n14816), .IN2(n14817), .QN(n14808) );
  NAND2X0 U15338 ( .IN1(n14818), .IN2(n14819), .QN(n14817) );
  NAND2X0 U15339 ( .IN1(n9650), .IN2(WX5925), .QN(n14819) );
  NAND2X0 U15340 ( .IN1(n3677), .IN2(WX6053), .QN(n14818) );
  NOR2X0 U15341 ( .IN1(n14820), .IN2(n14821), .QN(n14816) );
  NOR2X0 U15342 ( .IN1(n9383), .IN2(WX5861), .QN(n14821) );
  NOR2X0 U15343 ( .IN1(n9382), .IN2(WX5989), .QN(n14820) );
  NOR2X0 U15344 ( .IN1(n14822), .IN2(n14823), .QN(n14802) );
  NOR2X0 U15345 ( .IN1(DFF_745_n1), .IN2(n9974), .QN(n14823) );
  NOR2X0 U15346 ( .IN1(n9987), .IN2(n10577), .QN(n14822) );
  NAND2X0 U15347 ( .IN1(n10206), .IN2(n8564), .QN(n10577) );
  NAND2X0 U15348 ( .IN1(n14824), .IN2(n14825), .QN(WX4565) );
  NOR2X0 U15349 ( .IN1(n14826), .IN2(n14827), .QN(n14825) );
  NOR2X0 U15350 ( .IN1(n14828), .IN2(n9940), .QN(n14827) );
  NOR2X0 U15351 ( .IN1(n14003), .IN2(n9921), .QN(n14826) );
  INVX0 U15352 ( .INP(n14829), .ZN(n14003) );
  NAND2X0 U15353 ( .IN1(n14830), .IN2(n14831), .QN(n14829) );
  NAND2X0 U15354 ( .IN1(n14832), .IN2(n14833), .QN(n14831) );
  NAND2X0 U15355 ( .IN1(n14834), .IN2(n14835), .QN(n14833) );
  NAND2X0 U15356 ( .IN1(n9385), .IN2(WX5859), .QN(n14835) );
  NAND2X0 U15357 ( .IN1(n9384), .IN2(WX5987), .QN(n14834) );
  NOR2X0 U15358 ( .IN1(n14836), .IN2(n14837), .QN(n14832) );
  NOR2X0 U15359 ( .IN1(n9649), .IN2(WX5923), .QN(n14837) );
  NOR2X0 U15360 ( .IN1(n3679), .IN2(WX6051), .QN(n14836) );
  NAND2X0 U15361 ( .IN1(n14838), .IN2(n14839), .QN(n14830) );
  NAND2X0 U15362 ( .IN1(n14840), .IN2(n14841), .QN(n14839) );
  NAND2X0 U15363 ( .IN1(n9649), .IN2(WX5923), .QN(n14841) );
  NAND2X0 U15364 ( .IN1(n3679), .IN2(WX6051), .QN(n14840) );
  NOR2X0 U15365 ( .IN1(n14842), .IN2(n14843), .QN(n14838) );
  NOR2X0 U15366 ( .IN1(n9385), .IN2(WX5859), .QN(n14843) );
  NOR2X0 U15367 ( .IN1(n9384), .IN2(WX5987), .QN(n14842) );
  NOR2X0 U15368 ( .IN1(n14844), .IN2(n14845), .QN(n14824) );
  NOR2X0 U15369 ( .IN1(DFF_746_n1), .IN2(n9973), .QN(n14845) );
  NOR2X0 U15370 ( .IN1(n9987), .IN2(n10588), .QN(n14844) );
  NAND2X0 U15371 ( .IN1(n10206), .IN2(n8565), .QN(n10588) );
  NAND2X0 U15372 ( .IN1(n14846), .IN2(n14847), .QN(WX4563) );
  NOR2X0 U15373 ( .IN1(n14848), .IN2(n14849), .QN(n14847) );
  NOR2X0 U15374 ( .IN1(n9943), .IN2(n14850), .QN(n14849) );
  NOR2X0 U15375 ( .IN1(n14021), .IN2(n9921), .QN(n14848) );
  INVX0 U15376 ( .INP(n14851), .ZN(n14021) );
  NAND2X0 U15377 ( .IN1(n14852), .IN2(n14853), .QN(n14851) );
  NAND2X0 U15378 ( .IN1(n14854), .IN2(n14855), .QN(n14853) );
  NAND2X0 U15379 ( .IN1(n14856), .IN2(n14857), .QN(n14855) );
  NAND2X0 U15380 ( .IN1(n9387), .IN2(WX5857), .QN(n14857) );
  NAND2X0 U15381 ( .IN1(n9386), .IN2(WX5985), .QN(n14856) );
  NOR2X0 U15382 ( .IN1(n14858), .IN2(n14859), .QN(n14854) );
  NOR2X0 U15383 ( .IN1(n9507), .IN2(WX5921), .QN(n14859) );
  NOR2X0 U15384 ( .IN1(n3681), .IN2(WX6049), .QN(n14858) );
  NAND2X0 U15385 ( .IN1(n14860), .IN2(n14861), .QN(n14852) );
  NAND2X0 U15386 ( .IN1(n14862), .IN2(n14863), .QN(n14861) );
  NAND2X0 U15387 ( .IN1(n9507), .IN2(WX5921), .QN(n14863) );
  NAND2X0 U15388 ( .IN1(n3681), .IN2(WX6049), .QN(n14862) );
  NOR2X0 U15389 ( .IN1(n14864), .IN2(n14865), .QN(n14860) );
  NOR2X0 U15390 ( .IN1(n9387), .IN2(WX5857), .QN(n14865) );
  NOR2X0 U15391 ( .IN1(n9386), .IN2(WX5985), .QN(n14864) );
  NOR2X0 U15392 ( .IN1(n14866), .IN2(n14867), .QN(n14846) );
  NOR2X0 U15393 ( .IN1(DFF_747_n1), .IN2(n9973), .QN(n14867) );
  NOR2X0 U15394 ( .IN1(n9987), .IN2(n10589), .QN(n14866) );
  NAND2X0 U15395 ( .IN1(n10206), .IN2(n8566), .QN(n10589) );
  NAND2X0 U15396 ( .IN1(n14868), .IN2(n14869), .QN(WX4561) );
  NOR2X0 U15397 ( .IN1(n14870), .IN2(n14871), .QN(n14869) );
  NOR2X0 U15398 ( .IN1(n14872), .IN2(n9933), .QN(n14871) );
  NOR2X0 U15399 ( .IN1(n14043), .IN2(n9919), .QN(n14870) );
  INVX0 U15400 ( .INP(n14873), .ZN(n14043) );
  NAND2X0 U15401 ( .IN1(n14874), .IN2(n14875), .QN(n14873) );
  NAND2X0 U15402 ( .IN1(n14876), .IN2(n14877), .QN(n14875) );
  NAND2X0 U15403 ( .IN1(n14878), .IN2(n14879), .QN(n14877) );
  NAND2X0 U15404 ( .IN1(n9389), .IN2(WX5855), .QN(n14879) );
  NAND2X0 U15405 ( .IN1(n9388), .IN2(WX5983), .QN(n14878) );
  NOR2X0 U15406 ( .IN1(n14880), .IN2(n14881), .QN(n14876) );
  NOR2X0 U15407 ( .IN1(n9648), .IN2(WX5919), .QN(n14881) );
  NOR2X0 U15408 ( .IN1(n3683), .IN2(WX6047), .QN(n14880) );
  NAND2X0 U15409 ( .IN1(n14882), .IN2(n14883), .QN(n14874) );
  NAND2X0 U15410 ( .IN1(n14884), .IN2(n14885), .QN(n14883) );
  NAND2X0 U15411 ( .IN1(n9648), .IN2(WX5919), .QN(n14885) );
  NAND2X0 U15412 ( .IN1(n3683), .IN2(WX6047), .QN(n14884) );
  NOR2X0 U15413 ( .IN1(n14886), .IN2(n14887), .QN(n14882) );
  NOR2X0 U15414 ( .IN1(n9389), .IN2(WX5855), .QN(n14887) );
  NOR2X0 U15415 ( .IN1(n9388), .IN2(WX5983), .QN(n14886) );
  NOR2X0 U15416 ( .IN1(n14888), .IN2(n14889), .QN(n14868) );
  NOR2X0 U15417 ( .IN1(DFF_748_n1), .IN2(n9973), .QN(n14889) );
  NOR2X0 U15418 ( .IN1(n9987), .IN2(n10590), .QN(n14888) );
  NAND2X0 U15419 ( .IN1(n10206), .IN2(n8567), .QN(n10590) );
  NAND2X0 U15420 ( .IN1(n14890), .IN2(n14891), .QN(WX4559) );
  NOR2X0 U15421 ( .IN1(n14892), .IN2(n14893), .QN(n14891) );
  NOR2X0 U15422 ( .IN1(n9942), .IN2(n14894), .QN(n14893) );
  NOR2X0 U15423 ( .IN1(n14065), .IN2(n9921), .QN(n14892) );
  INVX0 U15424 ( .INP(n14895), .ZN(n14065) );
  NAND2X0 U15425 ( .IN1(n14896), .IN2(n14897), .QN(n14895) );
  NAND2X0 U15426 ( .IN1(n14898), .IN2(n14899), .QN(n14897) );
  NAND2X0 U15427 ( .IN1(n14900), .IN2(n14901), .QN(n14899) );
  NAND2X0 U15428 ( .IN1(n9391), .IN2(WX5853), .QN(n14901) );
  NAND2X0 U15429 ( .IN1(n9390), .IN2(WX5981), .QN(n14900) );
  NOR2X0 U15430 ( .IN1(n14902), .IN2(n14903), .QN(n14898) );
  NOR2X0 U15431 ( .IN1(n9647), .IN2(WX5917), .QN(n14903) );
  NOR2X0 U15432 ( .IN1(n3685), .IN2(WX6045), .QN(n14902) );
  NAND2X0 U15433 ( .IN1(n14904), .IN2(n14905), .QN(n14896) );
  NAND2X0 U15434 ( .IN1(n14906), .IN2(n14907), .QN(n14905) );
  NAND2X0 U15435 ( .IN1(n9647), .IN2(WX5917), .QN(n14907) );
  NAND2X0 U15436 ( .IN1(n3685), .IN2(WX6045), .QN(n14906) );
  NOR2X0 U15437 ( .IN1(n14908), .IN2(n14909), .QN(n14904) );
  NOR2X0 U15438 ( .IN1(n9391), .IN2(WX5853), .QN(n14909) );
  NOR2X0 U15439 ( .IN1(n9390), .IN2(WX5981), .QN(n14908) );
  NOR2X0 U15440 ( .IN1(n14910), .IN2(n14911), .QN(n14890) );
  NOR2X0 U15441 ( .IN1(DFF_749_n1), .IN2(n9973), .QN(n14911) );
  NOR2X0 U15442 ( .IN1(n9987), .IN2(n10591), .QN(n14910) );
  NAND2X0 U15443 ( .IN1(n10205), .IN2(n8568), .QN(n10591) );
  NAND2X0 U15444 ( .IN1(n14912), .IN2(n14913), .QN(WX4557) );
  NOR2X0 U15445 ( .IN1(n14914), .IN2(n14915), .QN(n14913) );
  NOR2X0 U15446 ( .IN1(n14916), .IN2(n9939), .QN(n14915) );
  NOR2X0 U15447 ( .IN1(n14087), .IN2(n9920), .QN(n14914) );
  INVX0 U15448 ( .INP(n14917), .ZN(n14087) );
  NAND2X0 U15449 ( .IN1(n14918), .IN2(n14919), .QN(n14917) );
  NAND2X0 U15450 ( .IN1(n14920), .IN2(n14921), .QN(n14919) );
  NAND2X0 U15451 ( .IN1(n14922), .IN2(n14923), .QN(n14921) );
  NAND2X0 U15452 ( .IN1(n9393), .IN2(WX5851), .QN(n14923) );
  NAND2X0 U15453 ( .IN1(n9392), .IN2(WX5979), .QN(n14922) );
  NOR2X0 U15454 ( .IN1(n14924), .IN2(n14925), .QN(n14920) );
  NOR2X0 U15455 ( .IN1(n9646), .IN2(WX5915), .QN(n14925) );
  NOR2X0 U15456 ( .IN1(n3687), .IN2(WX6043), .QN(n14924) );
  NAND2X0 U15457 ( .IN1(n14926), .IN2(n14927), .QN(n14918) );
  NAND2X0 U15458 ( .IN1(n14928), .IN2(n14929), .QN(n14927) );
  NAND2X0 U15459 ( .IN1(n9646), .IN2(WX5915), .QN(n14929) );
  NAND2X0 U15460 ( .IN1(n3687), .IN2(WX6043), .QN(n14928) );
  NOR2X0 U15461 ( .IN1(n14930), .IN2(n14931), .QN(n14926) );
  NOR2X0 U15462 ( .IN1(n9393), .IN2(WX5851), .QN(n14931) );
  NOR2X0 U15463 ( .IN1(n9392), .IN2(WX5979), .QN(n14930) );
  NOR2X0 U15464 ( .IN1(n14932), .IN2(n14933), .QN(n14912) );
  NOR2X0 U15465 ( .IN1(DFF_750_n1), .IN2(n9973), .QN(n14933) );
  NOR2X0 U15466 ( .IN1(n9987), .IN2(n10592), .QN(n14932) );
  NAND2X0 U15467 ( .IN1(n10205), .IN2(n8569), .QN(n10592) );
  NAND2X0 U15468 ( .IN1(n14934), .IN2(n14935), .QN(WX4555) );
  NOR2X0 U15469 ( .IN1(n14936), .IN2(n14937), .QN(n14935) );
  NOR2X0 U15470 ( .IN1(n9942), .IN2(n14938), .QN(n14937) );
  NOR2X0 U15471 ( .IN1(n14109), .IN2(n9920), .QN(n14936) );
  INVX0 U15472 ( .INP(n14939), .ZN(n14109) );
  NAND2X0 U15473 ( .IN1(n14940), .IN2(n14941), .QN(n14939) );
  NAND2X0 U15474 ( .IN1(n14942), .IN2(n14943), .QN(n14941) );
  NAND2X0 U15475 ( .IN1(n14944), .IN2(n14945), .QN(n14943) );
  NAND2X0 U15476 ( .IN1(n9395), .IN2(WX5849), .QN(n14945) );
  NAND2X0 U15477 ( .IN1(n9394), .IN2(WX5977), .QN(n14944) );
  NOR2X0 U15478 ( .IN1(n14946), .IN2(n14947), .QN(n14942) );
  NOR2X0 U15479 ( .IN1(n9645), .IN2(WX5913), .QN(n14947) );
  NOR2X0 U15480 ( .IN1(n3689), .IN2(WX6041), .QN(n14946) );
  NAND2X0 U15481 ( .IN1(n14948), .IN2(n14949), .QN(n14940) );
  NAND2X0 U15482 ( .IN1(n14950), .IN2(n14951), .QN(n14949) );
  NAND2X0 U15483 ( .IN1(n9645), .IN2(WX5913), .QN(n14951) );
  NAND2X0 U15484 ( .IN1(n3689), .IN2(WX6041), .QN(n14950) );
  NOR2X0 U15485 ( .IN1(n14952), .IN2(n14953), .QN(n14948) );
  NOR2X0 U15486 ( .IN1(n9395), .IN2(WX5849), .QN(n14953) );
  NOR2X0 U15487 ( .IN1(n9394), .IN2(WX5977), .QN(n14952) );
  NOR2X0 U15488 ( .IN1(n14954), .IN2(n14955), .QN(n14934) );
  NOR2X0 U15489 ( .IN1(DFF_751_n1), .IN2(n9972), .QN(n14955) );
  NOR2X0 U15490 ( .IN1(n9987), .IN2(n10593), .QN(n14954) );
  NAND2X0 U15491 ( .IN1(n10205), .IN2(n8570), .QN(n10593) );
  NAND2X0 U15492 ( .IN1(n14956), .IN2(n14957), .QN(WX4553) );
  NOR2X0 U15493 ( .IN1(n14958), .IN2(n14959), .QN(n14957) );
  NOR2X0 U15494 ( .IN1(n14960), .IN2(n10563), .QN(n14959) );
  NOR2X0 U15495 ( .IN1(n9922), .IN2(n14131), .QN(n14958) );
  NAND2X0 U15496 ( .IN1(n14961), .IN2(n14962), .QN(n14131) );
  NAND2X0 U15497 ( .IN1(n14963), .IN2(n14964), .QN(n14962) );
  INVX0 U15498 ( .INP(n14965), .ZN(n14961) );
  NOR2X0 U15499 ( .IN1(n14964), .IN2(n14963), .QN(n14965) );
  NAND2X0 U15500 ( .IN1(n14966), .IN2(n14967), .QN(n14963) );
  NAND2X0 U15501 ( .IN1(n14968), .IN2(WX5975), .QN(n14967) );
  NAND2X0 U15502 ( .IN1(n14969), .IN2(n14970), .QN(n14968) );
  NAND2X0 U15503 ( .IN1(test_so52), .IN2(WX5911), .QN(n14970) );
  NAND2X0 U15504 ( .IN1(n9131), .IN2(n9848), .QN(n14969) );
  NAND2X0 U15505 ( .IN1(n9132), .IN2(n14971), .QN(n14966) );
  NOR2X0 U15506 ( .IN1(n14972), .IN2(n14973), .QN(n14971) );
  NOR2X0 U15507 ( .IN1(test_so52), .IN2(WX5911), .QN(n14973) );
  NOR2X0 U15508 ( .IN1(n9131), .IN2(n9848), .QN(n14972) );
  NOR2X0 U15509 ( .IN1(n14974), .IN2(n14975), .QN(n14964) );
  INVX0 U15510 ( .INP(n14976), .ZN(n14975) );
  NAND2X0 U15511 ( .IN1(n18411), .IN2(n10018), .QN(n14976) );
  NOR2X0 U15512 ( .IN1(n10008), .IN2(n18411), .QN(n14974) );
  NOR2X0 U15513 ( .IN1(n14977), .IN2(n14978), .QN(n14956) );
  NOR2X0 U15514 ( .IN1(DFF_752_n1), .IN2(n9973), .QN(n14978) );
  NOR2X0 U15515 ( .IN1(n9987), .IN2(n10594), .QN(n14977) );
  NAND2X0 U15516 ( .IN1(n10205), .IN2(n8571), .QN(n10594) );
  NAND2X0 U15517 ( .IN1(n14979), .IN2(n14980), .QN(WX4551) );
  NOR2X0 U15518 ( .IN1(n14981), .IN2(n14982), .QN(n14980) );
  NOR2X0 U15519 ( .IN1(n9941), .IN2(n14983), .QN(n14982) );
  NOR2X0 U15520 ( .IN1(n14153), .IN2(n9920), .QN(n14981) );
  NOR2X0 U15521 ( .IN1(n14984), .IN2(n14985), .QN(n14153) );
  INVX0 U15522 ( .INP(n14986), .ZN(n14985) );
  NAND2X0 U15523 ( .IN1(n14987), .IN2(n14988), .QN(n14986) );
  NOR2X0 U15524 ( .IN1(n14988), .IN2(n14987), .QN(n14984) );
  NAND2X0 U15525 ( .IN1(n14989), .IN2(n14990), .QN(n14987) );
  NAND2X0 U15526 ( .IN1(n9134), .IN2(n14991), .QN(n14990) );
  INVX0 U15527 ( .INP(n14992), .ZN(n14989) );
  NOR2X0 U15528 ( .IN1(n14991), .IN2(n9134), .QN(n14992) );
  NOR2X0 U15529 ( .IN1(n14993), .IN2(n14994), .QN(n14991) );
  INVX0 U15530 ( .INP(n14995), .ZN(n14994) );
  NAND2X0 U15531 ( .IN1(n18410), .IN2(WX6037), .QN(n14995) );
  NOR2X0 U15532 ( .IN1(WX6037), .IN2(n18410), .QN(n14993) );
  NOR2X0 U15533 ( .IN1(n14996), .IN2(n14997), .QN(n14988) );
  INVX0 U15534 ( .INP(n14998), .ZN(n14997) );
  NAND2X0 U15535 ( .IN1(n9133), .IN2(n10018), .QN(n14998) );
  NOR2X0 U15536 ( .IN1(n10008), .IN2(n9133), .QN(n14996) );
  NOR2X0 U15537 ( .IN1(n14999), .IN2(n15000), .QN(n14979) );
  NOR2X0 U15538 ( .IN1(DFF_753_n1), .IN2(n9973), .QN(n15000) );
  NOR2X0 U15539 ( .IN1(n9987), .IN2(n10595), .QN(n14999) );
  NAND2X0 U15540 ( .IN1(n10205), .IN2(n8572), .QN(n10595) );
  NAND2X0 U15541 ( .IN1(n15001), .IN2(n15002), .QN(WX4549) );
  NOR2X0 U15542 ( .IN1(n15003), .IN2(n15004), .QN(n15002) );
  NOR2X0 U15543 ( .IN1(n15005), .IN2(n10563), .QN(n15004) );
  NOR2X0 U15544 ( .IN1(n9922), .IN2(n14175), .QN(n15003) );
  NAND2X0 U15545 ( .IN1(n15006), .IN2(n15007), .QN(n14175) );
  NAND2X0 U15546 ( .IN1(n15008), .IN2(n15009), .QN(n15007) );
  INVX0 U15547 ( .INP(n15010), .ZN(n15006) );
  NOR2X0 U15548 ( .IN1(n15009), .IN2(n15008), .QN(n15010) );
  NAND2X0 U15549 ( .IN1(n15011), .IN2(n15012), .QN(n15008) );
  NAND2X0 U15550 ( .IN1(n9643), .IN2(n15013), .QN(n15012) );
  INVX0 U15551 ( .INP(n15014), .ZN(n15013) );
  NAND2X0 U15552 ( .IN1(n15014), .IN2(WX6035), .QN(n15011) );
  NAND2X0 U15553 ( .IN1(n15015), .IN2(n15016), .QN(n15014) );
  INVX0 U15554 ( .INP(n15017), .ZN(n15016) );
  NOR2X0 U15555 ( .IN1(n9869), .IN2(n18409), .QN(n15017) );
  NAND2X0 U15556 ( .IN1(n18409), .IN2(n9869), .QN(n15015) );
  NOR2X0 U15557 ( .IN1(n15018), .IN2(n15019), .QN(n15009) );
  INVX0 U15558 ( .INP(n15020), .ZN(n15019) );
  NAND2X0 U15559 ( .IN1(n9135), .IN2(n10018), .QN(n15020) );
  NOR2X0 U15560 ( .IN1(n10008), .IN2(n9135), .QN(n15018) );
  NOR2X0 U15561 ( .IN1(n15021), .IN2(n15022), .QN(n15001) );
  NOR2X0 U15562 ( .IN1(DFF_754_n1), .IN2(n9972), .QN(n15022) );
  NOR2X0 U15563 ( .IN1(n9987), .IN2(n10596), .QN(n15021) );
  NAND2X0 U15564 ( .IN1(n10205), .IN2(n8573), .QN(n10596) );
  NAND2X0 U15565 ( .IN1(n15023), .IN2(n15024), .QN(WX4547) );
  NOR2X0 U15566 ( .IN1(n15025), .IN2(n15026), .QN(n15024) );
  NOR2X0 U15567 ( .IN1(n15027), .IN2(n10563), .QN(n15026) );
  NOR2X0 U15568 ( .IN1(n14197), .IN2(n9920), .QN(n15025) );
  NOR2X0 U15569 ( .IN1(n15028), .IN2(n15029), .QN(n14197) );
  INVX0 U15570 ( .INP(n15030), .ZN(n15029) );
  NAND2X0 U15571 ( .IN1(n15031), .IN2(n15032), .QN(n15030) );
  NOR2X0 U15572 ( .IN1(n15032), .IN2(n15031), .QN(n15028) );
  NAND2X0 U15573 ( .IN1(n15033), .IN2(n15034), .QN(n15031) );
  NAND2X0 U15574 ( .IN1(n9137), .IN2(n15035), .QN(n15034) );
  INVX0 U15575 ( .INP(n15036), .ZN(n15033) );
  NOR2X0 U15576 ( .IN1(n15035), .IN2(n9137), .QN(n15036) );
  NOR2X0 U15577 ( .IN1(n15037), .IN2(n15038), .QN(n15035) );
  INVX0 U15578 ( .INP(n15039), .ZN(n15038) );
  NAND2X0 U15579 ( .IN1(n18408), .IN2(WX6033), .QN(n15039) );
  NOR2X0 U15580 ( .IN1(WX6033), .IN2(n18408), .QN(n15037) );
  NOR2X0 U15581 ( .IN1(n15040), .IN2(n15041), .QN(n15032) );
  INVX0 U15582 ( .INP(n15042), .ZN(n15041) );
  NAND2X0 U15583 ( .IN1(n9136), .IN2(n10019), .QN(n15042) );
  NOR2X0 U15584 ( .IN1(n10008), .IN2(n9136), .QN(n15040) );
  NOR2X0 U15585 ( .IN1(n15043), .IN2(n15044), .QN(n15023) );
  NOR2X0 U15586 ( .IN1(DFF_755_n1), .IN2(n9973), .QN(n15044) );
  NOR2X0 U15587 ( .IN1(n9987), .IN2(n10597), .QN(n15043) );
  NAND2X0 U15588 ( .IN1(test_so33), .IN2(n10214), .QN(n10597) );
  NAND2X0 U15589 ( .IN1(n15045), .IN2(n15046), .QN(WX4545) );
  NOR2X0 U15590 ( .IN1(n15047), .IN2(n15048), .QN(n15046) );
  NOR2X0 U15591 ( .IN1(n15049), .IN2(n9939), .QN(n15048) );
  NOR2X0 U15592 ( .IN1(n9923), .IN2(n14219), .QN(n15047) );
  NAND2X0 U15593 ( .IN1(n15050), .IN2(n15051), .QN(n14219) );
  INVX0 U15594 ( .INP(n15052), .ZN(n15051) );
  NOR2X0 U15595 ( .IN1(n15053), .IN2(n15054), .QN(n15052) );
  NAND2X0 U15596 ( .IN1(n15054), .IN2(n15053), .QN(n15050) );
  NOR2X0 U15597 ( .IN1(n15055), .IN2(n15056), .QN(n15053) );
  INVX0 U15598 ( .INP(n15057), .ZN(n15056) );
  NAND2X0 U15599 ( .IN1(n9641), .IN2(n15058), .QN(n15057) );
  NOR2X0 U15600 ( .IN1(n15058), .IN2(n9641), .QN(n15055) );
  NOR2X0 U15601 ( .IN1(n15059), .IN2(n15060), .QN(n15058) );
  INVX0 U15602 ( .INP(n15061), .ZN(n15060) );
  NAND2X0 U15603 ( .IN1(test_so48), .IN2(n8483), .QN(n15061) );
  NOR2X0 U15604 ( .IN1(n8483), .IN2(test_so48), .QN(n15059) );
  NAND2X0 U15605 ( .IN1(n15062), .IN2(n15063), .QN(n15054) );
  NAND2X0 U15606 ( .IN1(n9138), .IN2(n10019), .QN(n15063) );
  INVX0 U15607 ( .INP(n15064), .ZN(n15062) );
  NOR2X0 U15608 ( .IN1(n10008), .IN2(n9138), .QN(n15064) );
  NOR2X0 U15609 ( .IN1(n15065), .IN2(n15066), .QN(n15045) );
  NOR2X0 U15610 ( .IN1(DFF_756_n1), .IN2(n9973), .QN(n15066) );
  NOR2X0 U15611 ( .IN1(n9987), .IN2(n10598), .QN(n15065) );
  NAND2X0 U15612 ( .IN1(n10205), .IN2(n8576), .QN(n10598) );
  NAND2X0 U15613 ( .IN1(n15067), .IN2(n15068), .QN(WX4543) );
  NOR2X0 U15614 ( .IN1(n15069), .IN2(n15070), .QN(n15068) );
  NOR2X0 U15615 ( .IN1(n15071), .IN2(n10563), .QN(n15070) );
  NOR2X0 U15616 ( .IN1(n14241), .IN2(n9920), .QN(n15069) );
  NOR2X0 U15617 ( .IN1(n15072), .IN2(n15073), .QN(n14241) );
  INVX0 U15618 ( .INP(n15074), .ZN(n15073) );
  NAND2X0 U15619 ( .IN1(n15075), .IN2(n15076), .QN(n15074) );
  NOR2X0 U15620 ( .IN1(n15076), .IN2(n15075), .QN(n15072) );
  NAND2X0 U15621 ( .IN1(n15077), .IN2(n15078), .QN(n15075) );
  NAND2X0 U15622 ( .IN1(n9140), .IN2(n15079), .QN(n15078) );
  INVX0 U15623 ( .INP(n15080), .ZN(n15077) );
  NOR2X0 U15624 ( .IN1(n15079), .IN2(n9140), .QN(n15080) );
  NOR2X0 U15625 ( .IN1(n15081), .IN2(n15082), .QN(n15079) );
  INVX0 U15626 ( .INP(n15083), .ZN(n15082) );
  NAND2X0 U15627 ( .IN1(n18406), .IN2(WX6029), .QN(n15083) );
  NOR2X0 U15628 ( .IN1(WX6029), .IN2(n18406), .QN(n15081) );
  NOR2X0 U15629 ( .IN1(n15084), .IN2(n15085), .QN(n15076) );
  INVX0 U15630 ( .INP(n15086), .ZN(n15085) );
  NAND2X0 U15631 ( .IN1(n9139), .IN2(n10019), .QN(n15086) );
  NOR2X0 U15632 ( .IN1(n10008), .IN2(n9139), .QN(n15084) );
  NOR2X0 U15633 ( .IN1(n15087), .IN2(n15088), .QN(n15067) );
  NOR2X0 U15634 ( .IN1(DFF_757_n1), .IN2(n9973), .QN(n15088) );
  NOR2X0 U15635 ( .IN1(n9986), .IN2(n10599), .QN(n15087) );
  NAND2X0 U15636 ( .IN1(n10205), .IN2(n8577), .QN(n10599) );
  NAND2X0 U15637 ( .IN1(n15089), .IN2(n15090), .QN(WX4541) );
  NOR2X0 U15638 ( .IN1(n15091), .IN2(n15092), .QN(n15090) );
  NOR2X0 U15639 ( .IN1(n15093), .IN2(n9932), .QN(n15092) );
  NOR2X0 U15640 ( .IN1(n9923), .IN2(n14264), .QN(n15091) );
  NAND2X0 U15641 ( .IN1(n15094), .IN2(n15095), .QN(n14264) );
  INVX0 U15642 ( .INP(n15096), .ZN(n15095) );
  NOR2X0 U15643 ( .IN1(n15097), .IN2(n15098), .QN(n15096) );
  NAND2X0 U15644 ( .IN1(n15098), .IN2(n15097), .QN(n15094) );
  INVX0 U15645 ( .INP(n15099), .ZN(n15097) );
  NAND2X0 U15646 ( .IN1(n15100), .IN2(n15101), .QN(n15099) );
  NAND2X0 U15647 ( .IN1(n15102), .IN2(WX5963), .QN(n15101) );
  NAND2X0 U15648 ( .IN1(n15103), .IN2(n15104), .QN(n15102) );
  NAND2X0 U15649 ( .IN1(test_so46), .IN2(WX5899), .QN(n15104) );
  NAND2X0 U15650 ( .IN1(n9141), .IN2(n9842), .QN(n15103) );
  NAND2X0 U15651 ( .IN1(n9142), .IN2(n15105), .QN(n15100) );
  NOR2X0 U15652 ( .IN1(n15106), .IN2(n15107), .QN(n15105) );
  NOR2X0 U15653 ( .IN1(test_so46), .IN2(WX5899), .QN(n15107) );
  NOR2X0 U15654 ( .IN1(n9141), .IN2(n9842), .QN(n15106) );
  NAND2X0 U15655 ( .IN1(n15108), .IN2(n15109), .QN(n15098) );
  NAND2X0 U15656 ( .IN1(n9639), .IN2(n10019), .QN(n15109) );
  NAND2X0 U15657 ( .IN1(TM1), .IN2(WX6027), .QN(n15108) );
  NOR2X0 U15658 ( .IN1(n15110), .IN2(n15111), .QN(n15089) );
  NOR2X0 U15659 ( .IN1(n9976), .IN2(n9859), .QN(n15111) );
  NOR2X0 U15660 ( .IN1(n9986), .IN2(n10600), .QN(n15110) );
  NAND2X0 U15661 ( .IN1(n10205), .IN2(n8578), .QN(n10600) );
  NAND2X0 U15662 ( .IN1(n15112), .IN2(n15113), .QN(WX4539) );
  NOR2X0 U15663 ( .IN1(n15114), .IN2(n15115), .QN(n15113) );
  NOR2X0 U15664 ( .IN1(n15116), .IN2(n9934), .QN(n15115) );
  NOR2X0 U15665 ( .IN1(n14286), .IN2(n9920), .QN(n15114) );
  NOR2X0 U15666 ( .IN1(n15117), .IN2(n15118), .QN(n14286) );
  INVX0 U15667 ( .INP(n15119), .ZN(n15118) );
  NAND2X0 U15668 ( .IN1(n15120), .IN2(n15121), .QN(n15119) );
  NOR2X0 U15669 ( .IN1(n15121), .IN2(n15120), .QN(n15117) );
  NAND2X0 U15670 ( .IN1(n15122), .IN2(n15123), .QN(n15120) );
  NAND2X0 U15671 ( .IN1(n9144), .IN2(n15124), .QN(n15123) );
  INVX0 U15672 ( .INP(n15125), .ZN(n15122) );
  NOR2X0 U15673 ( .IN1(n15124), .IN2(n9144), .QN(n15125) );
  NOR2X0 U15674 ( .IN1(n15126), .IN2(n15127), .QN(n15124) );
  INVX0 U15675 ( .INP(n15128), .ZN(n15127) );
  NAND2X0 U15676 ( .IN1(n18405), .IN2(WX6025), .QN(n15128) );
  NOR2X0 U15677 ( .IN1(WX6025), .IN2(n18405), .QN(n15126) );
  NOR2X0 U15678 ( .IN1(n15129), .IN2(n15130), .QN(n15121) );
  INVX0 U15679 ( .INP(n15131), .ZN(n15130) );
  NAND2X0 U15680 ( .IN1(n9143), .IN2(n10019), .QN(n15131) );
  NOR2X0 U15681 ( .IN1(n10008), .IN2(n9143), .QN(n15129) );
  NOR2X0 U15682 ( .IN1(n15132), .IN2(n15133), .QN(n15112) );
  NOR2X0 U15683 ( .IN1(DFF_759_n1), .IN2(n9972), .QN(n15133) );
  NOR2X0 U15684 ( .IN1(n9986), .IN2(n10601), .QN(n15132) );
  NAND2X0 U15685 ( .IN1(n10204), .IN2(n8579), .QN(n10601) );
  NAND2X0 U15686 ( .IN1(n15134), .IN2(n15135), .QN(WX4537) );
  NOR2X0 U15687 ( .IN1(n15136), .IN2(n15137), .QN(n15135) );
  NOR2X0 U15688 ( .IN1(n15138), .IN2(n9935), .QN(n15137) );
  NOR2X0 U15689 ( .IN1(n14308), .IN2(n9919), .QN(n15136) );
  NOR2X0 U15690 ( .IN1(n15139), .IN2(n15140), .QN(n14308) );
  INVX0 U15691 ( .INP(n15141), .ZN(n15140) );
  NAND2X0 U15692 ( .IN1(n15142), .IN2(n15143), .QN(n15141) );
  NOR2X0 U15693 ( .IN1(n15143), .IN2(n15142), .QN(n15139) );
  NAND2X0 U15694 ( .IN1(n15144), .IN2(n15145), .QN(n15142) );
  NAND2X0 U15695 ( .IN1(n9146), .IN2(n15146), .QN(n15145) );
  INVX0 U15696 ( .INP(n15147), .ZN(n15144) );
  NOR2X0 U15697 ( .IN1(n15146), .IN2(n9146), .QN(n15147) );
  NOR2X0 U15698 ( .IN1(n15148), .IN2(n15149), .QN(n15146) );
  INVX0 U15699 ( .INP(n15150), .ZN(n15149) );
  NAND2X0 U15700 ( .IN1(n18404), .IN2(WX6023), .QN(n15150) );
  NOR2X0 U15701 ( .IN1(WX6023), .IN2(n18404), .QN(n15148) );
  NOR2X0 U15702 ( .IN1(n15151), .IN2(n15152), .QN(n15143) );
  INVX0 U15703 ( .INP(n15153), .ZN(n15152) );
  NAND2X0 U15704 ( .IN1(n9145), .IN2(n10019), .QN(n15153) );
  NOR2X0 U15705 ( .IN1(n10008), .IN2(n9145), .QN(n15151) );
  NOR2X0 U15706 ( .IN1(n15154), .IN2(n15155), .QN(n15134) );
  NOR2X0 U15707 ( .IN1(DFF_760_n1), .IN2(n9972), .QN(n15155) );
  NOR2X0 U15708 ( .IN1(n9986), .IN2(n10602), .QN(n15154) );
  NAND2X0 U15709 ( .IN1(n10204), .IN2(n8580), .QN(n10602) );
  NAND2X0 U15710 ( .IN1(n15156), .IN2(n15157), .QN(WX4535) );
  NOR2X0 U15711 ( .IN1(n15158), .IN2(n15159), .QN(n15157) );
  NOR2X0 U15712 ( .IN1(n15160), .IN2(n9939), .QN(n15159) );
  NOR2X0 U15713 ( .IN1(n14330), .IN2(n9919), .QN(n15158) );
  NOR2X0 U15714 ( .IN1(n15161), .IN2(n15162), .QN(n14330) );
  INVX0 U15715 ( .INP(n15163), .ZN(n15162) );
  NAND2X0 U15716 ( .IN1(n15164), .IN2(n15165), .QN(n15163) );
  NOR2X0 U15717 ( .IN1(n15165), .IN2(n15164), .QN(n15161) );
  NAND2X0 U15718 ( .IN1(n15166), .IN2(n15167), .QN(n15164) );
  NAND2X0 U15719 ( .IN1(n9148), .IN2(n15168), .QN(n15167) );
  INVX0 U15720 ( .INP(n15169), .ZN(n15166) );
  NOR2X0 U15721 ( .IN1(n15168), .IN2(n9148), .QN(n15169) );
  NOR2X0 U15722 ( .IN1(n15170), .IN2(n15171), .QN(n15168) );
  INVX0 U15723 ( .INP(n15172), .ZN(n15171) );
  NAND2X0 U15724 ( .IN1(n18403), .IN2(WX6021), .QN(n15172) );
  NOR2X0 U15725 ( .IN1(WX6021), .IN2(n18403), .QN(n15170) );
  NOR2X0 U15726 ( .IN1(n15173), .IN2(n15174), .QN(n15165) );
  INVX0 U15727 ( .INP(n15175), .ZN(n15174) );
  NAND2X0 U15728 ( .IN1(n9147), .IN2(n10019), .QN(n15175) );
  NOR2X0 U15729 ( .IN1(n10008), .IN2(n9147), .QN(n15173) );
  NOR2X0 U15730 ( .IN1(n15176), .IN2(n15177), .QN(n15156) );
  NOR2X0 U15731 ( .IN1(DFF_761_n1), .IN2(n9972), .QN(n15177) );
  NOR2X0 U15732 ( .IN1(n9986), .IN2(n10603), .QN(n15176) );
  NAND2X0 U15733 ( .IN1(n10204), .IN2(n8581), .QN(n10603) );
  NAND2X0 U15734 ( .IN1(n15178), .IN2(n15179), .QN(WX4533) );
  NOR2X0 U15735 ( .IN1(n15180), .IN2(n15181), .QN(n15179) );
  NOR2X0 U15736 ( .IN1(n15182), .IN2(n9939), .QN(n15181) );
  NOR2X0 U15737 ( .IN1(n14352), .IN2(n9919), .QN(n15180) );
  NOR2X0 U15738 ( .IN1(n15183), .IN2(n15184), .QN(n14352) );
  INVX0 U15739 ( .INP(n15185), .ZN(n15184) );
  NAND2X0 U15740 ( .IN1(n15186), .IN2(n15187), .QN(n15185) );
  NOR2X0 U15741 ( .IN1(n15187), .IN2(n15186), .QN(n15183) );
  NAND2X0 U15742 ( .IN1(n15188), .IN2(n15189), .QN(n15186) );
  NAND2X0 U15743 ( .IN1(n9150), .IN2(n15190), .QN(n15189) );
  INVX0 U15744 ( .INP(n15191), .ZN(n15188) );
  NOR2X0 U15745 ( .IN1(n15190), .IN2(n9150), .QN(n15191) );
  NOR2X0 U15746 ( .IN1(n15192), .IN2(n15193), .QN(n15190) );
  INVX0 U15747 ( .INP(n15194), .ZN(n15193) );
  NAND2X0 U15748 ( .IN1(n18402), .IN2(WX6019), .QN(n15194) );
  NOR2X0 U15749 ( .IN1(WX6019), .IN2(n18402), .QN(n15192) );
  NOR2X0 U15750 ( .IN1(n15195), .IN2(n15196), .QN(n15187) );
  INVX0 U15751 ( .INP(n15197), .ZN(n15196) );
  NAND2X0 U15752 ( .IN1(n9149), .IN2(n10019), .QN(n15197) );
  NOR2X0 U15753 ( .IN1(n10008), .IN2(n9149), .QN(n15195) );
  NOR2X0 U15754 ( .IN1(n15198), .IN2(n15199), .QN(n15178) );
  NOR2X0 U15755 ( .IN1(DFF_762_n1), .IN2(n9972), .QN(n15199) );
  NOR2X0 U15756 ( .IN1(n9986), .IN2(n10604), .QN(n15198) );
  NAND2X0 U15757 ( .IN1(n10204), .IN2(n8582), .QN(n10604) );
  NAND2X0 U15758 ( .IN1(n15200), .IN2(n15201), .QN(WX4531) );
  NOR2X0 U15759 ( .IN1(n15202), .IN2(n15203), .QN(n15201) );
  NOR2X0 U15760 ( .IN1(n15204), .IN2(n9939), .QN(n15203) );
  NOR2X0 U15761 ( .IN1(n14374), .IN2(n9919), .QN(n15202) );
  NOR2X0 U15762 ( .IN1(n15205), .IN2(n15206), .QN(n14374) );
  INVX0 U15763 ( .INP(n15207), .ZN(n15206) );
  NAND2X0 U15764 ( .IN1(n15208), .IN2(n15209), .QN(n15207) );
  NOR2X0 U15765 ( .IN1(n15209), .IN2(n15208), .QN(n15205) );
  NAND2X0 U15766 ( .IN1(n15210), .IN2(n15211), .QN(n15208) );
  NAND2X0 U15767 ( .IN1(n9152), .IN2(n15212), .QN(n15211) );
  INVX0 U15768 ( .INP(n15213), .ZN(n15210) );
  NOR2X0 U15769 ( .IN1(n15212), .IN2(n9152), .QN(n15213) );
  NOR2X0 U15770 ( .IN1(n15214), .IN2(n15215), .QN(n15212) );
  INVX0 U15771 ( .INP(n15216), .ZN(n15215) );
  NAND2X0 U15772 ( .IN1(n18401), .IN2(WX6017), .QN(n15216) );
  NOR2X0 U15773 ( .IN1(WX6017), .IN2(n18401), .QN(n15214) );
  NOR2X0 U15774 ( .IN1(n15217), .IN2(n15218), .QN(n15209) );
  INVX0 U15775 ( .INP(n15219), .ZN(n15218) );
  NAND2X0 U15776 ( .IN1(n9151), .IN2(n10019), .QN(n15219) );
  NOR2X0 U15777 ( .IN1(n10008), .IN2(n9151), .QN(n15217) );
  NOR2X0 U15778 ( .IN1(n15220), .IN2(n15221), .QN(n15200) );
  NOR2X0 U15779 ( .IN1(DFF_763_n1), .IN2(n9972), .QN(n15221) );
  NOR2X0 U15780 ( .IN1(n9986), .IN2(n10605), .QN(n15220) );
  NAND2X0 U15781 ( .IN1(n10204), .IN2(n8583), .QN(n10605) );
  NAND2X0 U15782 ( .IN1(n15222), .IN2(n15223), .QN(WX4529) );
  NOR2X0 U15783 ( .IN1(n15224), .IN2(n15225), .QN(n15223) );
  NOR2X0 U15784 ( .IN1(n9941), .IN2(n15226), .QN(n15225) );
  NOR2X0 U15785 ( .IN1(n14397), .IN2(n9919), .QN(n15224) );
  NOR2X0 U15786 ( .IN1(n15227), .IN2(n15228), .QN(n14397) );
  INVX0 U15787 ( .INP(n15229), .ZN(n15228) );
  NAND2X0 U15788 ( .IN1(n15230), .IN2(n15231), .QN(n15229) );
  NOR2X0 U15789 ( .IN1(n15231), .IN2(n15230), .QN(n15227) );
  NAND2X0 U15790 ( .IN1(n15232), .IN2(n15233), .QN(n15230) );
  NAND2X0 U15791 ( .IN1(n9154), .IN2(n15234), .QN(n15233) );
  INVX0 U15792 ( .INP(n15235), .ZN(n15232) );
  NOR2X0 U15793 ( .IN1(n15234), .IN2(n9154), .QN(n15235) );
  NOR2X0 U15794 ( .IN1(n15236), .IN2(n15237), .QN(n15234) );
  INVX0 U15795 ( .INP(n15238), .ZN(n15237) );
  NAND2X0 U15796 ( .IN1(n18400), .IN2(WX6015), .QN(n15238) );
  NOR2X0 U15797 ( .IN1(WX6015), .IN2(n18400), .QN(n15236) );
  NOR2X0 U15798 ( .IN1(n15239), .IN2(n15240), .QN(n15231) );
  INVX0 U15799 ( .INP(n15241), .ZN(n15240) );
  NAND2X0 U15800 ( .IN1(n9153), .IN2(n10019), .QN(n15241) );
  NOR2X0 U15801 ( .IN1(n10008), .IN2(n9153), .QN(n15239) );
  NOR2X0 U15802 ( .IN1(n15242), .IN2(n15243), .QN(n15222) );
  NOR2X0 U15803 ( .IN1(DFF_764_n1), .IN2(n9972), .QN(n15243) );
  NOR2X0 U15804 ( .IN1(n9986), .IN2(n10606), .QN(n15242) );
  NAND2X0 U15805 ( .IN1(n10204), .IN2(n8584), .QN(n10606) );
  NAND2X0 U15806 ( .IN1(n15244), .IN2(n15245), .QN(WX4527) );
  NOR2X0 U15807 ( .IN1(n15246), .IN2(n15247), .QN(n15245) );
  NOR2X0 U15808 ( .IN1(n15248), .IN2(n9939), .QN(n15247) );
  NOR2X0 U15809 ( .IN1(n14419), .IN2(n9919), .QN(n15246) );
  NOR2X0 U15810 ( .IN1(n15249), .IN2(n15250), .QN(n14419) );
  INVX0 U15811 ( .INP(n15251), .ZN(n15250) );
  NAND2X0 U15812 ( .IN1(n15252), .IN2(n15253), .QN(n15251) );
  NOR2X0 U15813 ( .IN1(n15253), .IN2(n15252), .QN(n15249) );
  NAND2X0 U15814 ( .IN1(n15254), .IN2(n15255), .QN(n15252) );
  NAND2X0 U15815 ( .IN1(n9156), .IN2(n15256), .QN(n15255) );
  INVX0 U15816 ( .INP(n15257), .ZN(n15254) );
  NOR2X0 U15817 ( .IN1(n15256), .IN2(n9156), .QN(n15257) );
  NOR2X0 U15818 ( .IN1(n15258), .IN2(n15259), .QN(n15256) );
  INVX0 U15819 ( .INP(n15260), .ZN(n15259) );
  NAND2X0 U15820 ( .IN1(n18399), .IN2(WX6013), .QN(n15260) );
  NOR2X0 U15821 ( .IN1(WX6013), .IN2(n18399), .QN(n15258) );
  NOR2X0 U15822 ( .IN1(n15261), .IN2(n15262), .QN(n15253) );
  INVX0 U15823 ( .INP(n15263), .ZN(n15262) );
  NAND2X0 U15824 ( .IN1(n9155), .IN2(n10019), .QN(n15263) );
  NOR2X0 U15825 ( .IN1(n10009), .IN2(n9155), .QN(n15261) );
  NOR2X0 U15826 ( .IN1(n15264), .IN2(n15265), .QN(n15244) );
  NOR2X0 U15827 ( .IN1(DFF_765_n1), .IN2(n9972), .QN(n15265) );
  NOR2X0 U15828 ( .IN1(n9986), .IN2(n10607), .QN(n15264) );
  NAND2X0 U15829 ( .IN1(n10204), .IN2(n8585), .QN(n10607) );
  NAND2X0 U15830 ( .IN1(n15266), .IN2(n15267), .QN(WX4525) );
  NOR2X0 U15831 ( .IN1(n15268), .IN2(n15269), .QN(n15267) );
  NOR2X0 U15832 ( .IN1(n9941), .IN2(n15270), .QN(n15269) );
  NOR2X0 U15833 ( .IN1(n14441), .IN2(n9919), .QN(n15268) );
  NOR2X0 U15834 ( .IN1(n15271), .IN2(n15272), .QN(n14441) );
  INVX0 U15835 ( .INP(n15273), .ZN(n15272) );
  NAND2X0 U15836 ( .IN1(n15274), .IN2(n15275), .QN(n15273) );
  NOR2X0 U15837 ( .IN1(n15275), .IN2(n15274), .QN(n15271) );
  NAND2X0 U15838 ( .IN1(n15276), .IN2(n15277), .QN(n15274) );
  NAND2X0 U15839 ( .IN1(n9158), .IN2(n15278), .QN(n15277) );
  INVX0 U15840 ( .INP(n15279), .ZN(n15276) );
  NOR2X0 U15841 ( .IN1(n15278), .IN2(n9158), .QN(n15279) );
  NOR2X0 U15842 ( .IN1(n15280), .IN2(n15281), .QN(n15278) );
  INVX0 U15843 ( .INP(n15282), .ZN(n15281) );
  NAND2X0 U15844 ( .IN1(n18398), .IN2(WX6011), .QN(n15282) );
  NOR2X0 U15845 ( .IN1(WX6011), .IN2(n18398), .QN(n15280) );
  NOR2X0 U15846 ( .IN1(n15283), .IN2(n15284), .QN(n15275) );
  INVX0 U15847 ( .INP(n15285), .ZN(n15284) );
  NAND2X0 U15848 ( .IN1(n9157), .IN2(n10019), .QN(n15285) );
  NOR2X0 U15849 ( .IN1(n10009), .IN2(n9157), .QN(n15283) );
  NOR2X0 U15850 ( .IN1(n15286), .IN2(n15287), .QN(n15266) );
  NOR2X0 U15851 ( .IN1(DFF_766_n1), .IN2(n9972), .QN(n15287) );
  NOR2X0 U15852 ( .IN1(n9986), .IN2(n10608), .QN(n15286) );
  NAND2X0 U15853 ( .IN1(n10204), .IN2(n8586), .QN(n10608) );
  NAND2X0 U15854 ( .IN1(n15288), .IN2(n15289), .QN(WX4523) );
  NOR2X0 U15855 ( .IN1(n15290), .IN2(n15291), .QN(n15289) );
  NOR2X0 U15856 ( .IN1(n15292), .IN2(n9939), .QN(n15291) );
  NOR2X0 U15857 ( .IN1(n14463), .IN2(n9919), .QN(n15290) );
  NOR2X0 U15858 ( .IN1(n15293), .IN2(n15294), .QN(n14463) );
  INVX0 U15859 ( .INP(n15295), .ZN(n15294) );
  NAND2X0 U15860 ( .IN1(n15296), .IN2(n15297), .QN(n15295) );
  NOR2X0 U15861 ( .IN1(n15297), .IN2(n15296), .QN(n15293) );
  NAND2X0 U15862 ( .IN1(n15298), .IN2(n15299), .QN(n15296) );
  NAND2X0 U15863 ( .IN1(n9012), .IN2(n15300), .QN(n15299) );
  INVX0 U15864 ( .INP(n15301), .ZN(n15298) );
  NOR2X0 U15865 ( .IN1(n15300), .IN2(n9012), .QN(n15301) );
  NOR2X0 U15866 ( .IN1(n15302), .IN2(n15303), .QN(n15300) );
  INVX0 U15867 ( .INP(n15304), .ZN(n15303) );
  NAND2X0 U15868 ( .IN1(n18397), .IN2(WX6009), .QN(n15304) );
  NOR2X0 U15869 ( .IN1(WX6009), .IN2(n18397), .QN(n15302) );
  NOR2X0 U15870 ( .IN1(n15305), .IN2(n15306), .QN(n15297) );
  INVX0 U15871 ( .INP(n15307), .ZN(n15306) );
  NAND2X0 U15872 ( .IN1(n9011), .IN2(n10019), .QN(n15307) );
  NOR2X0 U15873 ( .IN1(n10009), .IN2(n9011), .QN(n15305) );
  NOR2X0 U15874 ( .IN1(n15308), .IN2(n15309), .QN(n15288) );
  NOR2X0 U15875 ( .IN1(n9493), .IN2(n11994), .QN(n15309) );
  NOR2X0 U15876 ( .IN1(DFF_767_n1), .IN2(n9972), .QN(n15308) );
  INVX0 U15877 ( .INP(n15310), .ZN(WX4425) );
  NAND2X0 U15878 ( .IN1(n10204), .IN2(n9493), .QN(n15310) );
  NOR2X0 U15879 ( .IN1(n10331), .IN2(n15311), .QN(WX3912) );
  NAND2X0 U15880 ( .IN1(n15312), .IN2(n15313), .QN(n15311) );
  INVX0 U15881 ( .INP(n15314), .ZN(n15313) );
  NOR2X0 U15882 ( .IN1(WX3423), .IN2(DFF_574_n1), .QN(n15314) );
  NAND2X0 U15883 ( .IN1(DFF_574_n1), .IN2(WX3423), .QN(n15312) );
  NOR2X0 U15884 ( .IN1(n10331), .IN2(n15315), .QN(WX3910) );
  NAND2X0 U15885 ( .IN1(n15316), .IN2(n15317), .QN(n15315) );
  INVX0 U15886 ( .INP(n15318), .ZN(n15317) );
  NOR2X0 U15887 ( .IN1(WX3425), .IN2(DFF_573_n1), .QN(n15318) );
  NAND2X0 U15888 ( .IN1(DFF_573_n1), .IN2(WX3425), .QN(n15316) );
  NOR2X0 U15889 ( .IN1(n10331), .IN2(n15319), .QN(WX3908) );
  NAND2X0 U15890 ( .IN1(n15320), .IN2(n15321), .QN(n15319) );
  INVX0 U15891 ( .INP(n15322), .ZN(n15321) );
  NOR2X0 U15892 ( .IN1(WX3427), .IN2(DFF_572_n1), .QN(n15322) );
  NAND2X0 U15893 ( .IN1(DFF_572_n1), .IN2(WX3427), .QN(n15320) );
  NOR2X0 U15894 ( .IN1(n10331), .IN2(n15323), .QN(WX3906) );
  NOR2X0 U15895 ( .IN1(n15324), .IN2(n15325), .QN(n15323) );
  NOR2X0 U15896 ( .IN1(test_so32), .IN2(WX3429), .QN(n15325) );
  NOR2X0 U15897 ( .IN1(n9688), .IN2(n9860), .QN(n15324) );
  NOR2X0 U15898 ( .IN1(n10331), .IN2(n15326), .QN(WX3904) );
  NAND2X0 U15899 ( .IN1(n15327), .IN2(n15328), .QN(n15326) );
  INVX0 U15900 ( .INP(n15329), .ZN(n15328) );
  NOR2X0 U15901 ( .IN1(WX3431), .IN2(DFF_570_n1), .QN(n15329) );
  NAND2X0 U15902 ( .IN1(DFF_570_n1), .IN2(WX3431), .QN(n15327) );
  NOR2X0 U15903 ( .IN1(n10331), .IN2(n15330), .QN(WX3902) );
  NAND2X0 U15904 ( .IN1(n15331), .IN2(n15332), .QN(n15330) );
  INVX0 U15905 ( .INP(n15333), .ZN(n15332) );
  NOR2X0 U15906 ( .IN1(WX3433), .IN2(DFF_569_n1), .QN(n15333) );
  NAND2X0 U15907 ( .IN1(DFF_569_n1), .IN2(WX3433), .QN(n15331) );
  NOR2X0 U15908 ( .IN1(n10331), .IN2(n15334), .QN(WX3900) );
  NAND2X0 U15909 ( .IN1(n15335), .IN2(n15336), .QN(n15334) );
  INVX0 U15910 ( .INP(n15337), .ZN(n15336) );
  NOR2X0 U15911 ( .IN1(WX3435), .IN2(DFF_568_n1), .QN(n15337) );
  NAND2X0 U15912 ( .IN1(DFF_568_n1), .IN2(WX3435), .QN(n15335) );
  NOR2X0 U15913 ( .IN1(n10332), .IN2(n15338), .QN(WX3898) );
  NAND2X0 U15914 ( .IN1(n15339), .IN2(n15340), .QN(n15338) );
  INVX0 U15915 ( .INP(n15341), .ZN(n15340) );
  NOR2X0 U15916 ( .IN1(WX3437), .IN2(DFF_567_n1), .QN(n15341) );
  NAND2X0 U15917 ( .IN1(DFF_567_n1), .IN2(WX3437), .QN(n15339) );
  NOR2X0 U15918 ( .IN1(n10332), .IN2(n15342), .QN(WX3896) );
  NOR2X0 U15919 ( .IN1(n15343), .IN2(n15344), .QN(n15342) );
  INVX0 U15920 ( .INP(n15345), .ZN(n15344) );
  NAND2X0 U15921 ( .IN1(n9831), .IN2(DFF_566_n1), .QN(n15345) );
  NOR2X0 U15922 ( .IN1(DFF_566_n1), .IN2(n9831), .QN(n15343) );
  NOR2X0 U15923 ( .IN1(n10332), .IN2(n15346), .QN(WX3894) );
  NAND2X0 U15924 ( .IN1(n15347), .IN2(n15348), .QN(n15346) );
  INVX0 U15925 ( .INP(n15349), .ZN(n15348) );
  NOR2X0 U15926 ( .IN1(WX3441), .IN2(DFF_565_n1), .QN(n15349) );
  NAND2X0 U15927 ( .IN1(DFF_565_n1), .IN2(WX3441), .QN(n15347) );
  NOR2X0 U15928 ( .IN1(n10332), .IN2(n15350), .QN(WX3892) );
  NAND2X0 U15929 ( .IN1(n15351), .IN2(n15352), .QN(n15350) );
  INVX0 U15930 ( .INP(n15353), .ZN(n15352) );
  NOR2X0 U15931 ( .IN1(WX3443), .IN2(DFF_564_n1), .QN(n15353) );
  NAND2X0 U15932 ( .IN1(DFF_564_n1), .IN2(WX3443), .QN(n15351) );
  NOR2X0 U15933 ( .IN1(n10332), .IN2(n15354), .QN(WX3890) );
  NAND2X0 U15934 ( .IN1(n15355), .IN2(n15356), .QN(n15354) );
  INVX0 U15935 ( .INP(n15357), .ZN(n15356) );
  NOR2X0 U15936 ( .IN1(WX3445), .IN2(DFF_563_n1), .QN(n15357) );
  NAND2X0 U15937 ( .IN1(DFF_563_n1), .IN2(WX3445), .QN(n15355) );
  NOR2X0 U15938 ( .IN1(n10332), .IN2(n15358), .QN(WX3888) );
  NAND2X0 U15939 ( .IN1(n15359), .IN2(n15360), .QN(n15358) );
  INVX0 U15940 ( .INP(n15361), .ZN(n15360) );
  NOR2X0 U15941 ( .IN1(WX3447), .IN2(DFF_562_n1), .QN(n15361) );
  NAND2X0 U15942 ( .IN1(DFF_562_n1), .IN2(WX3447), .QN(n15359) );
  NOR2X0 U15943 ( .IN1(n10332), .IN2(n15362), .QN(WX3886) );
  NAND2X0 U15944 ( .IN1(n15363), .IN2(n15364), .QN(n15362) );
  INVX0 U15945 ( .INP(n15365), .ZN(n15364) );
  NOR2X0 U15946 ( .IN1(WX3449), .IN2(DFF_561_n1), .QN(n15365) );
  NAND2X0 U15947 ( .IN1(DFF_561_n1), .IN2(WX3449), .QN(n15363) );
  NOR2X0 U15948 ( .IN1(n10332), .IN2(n15366), .QN(WX3884) );
  NAND2X0 U15949 ( .IN1(n15367), .IN2(n15368), .QN(n15366) );
  INVX0 U15950 ( .INP(n15369), .ZN(n15368) );
  NOR2X0 U15951 ( .IN1(WX3451), .IN2(DFF_560_n1), .QN(n15369) );
  NAND2X0 U15952 ( .IN1(DFF_560_n1), .IN2(WX3451), .QN(n15367) );
  NOR2X0 U15953 ( .IN1(n10332), .IN2(n15370), .QN(WX3882) );
  NOR2X0 U15954 ( .IN1(n15371), .IN2(n15372), .QN(n15370) );
  INVX0 U15955 ( .INP(n15373), .ZN(n15372) );
  NAND2X0 U15956 ( .IN1(CRC_OUT_7_15), .IN2(n15374), .QN(n15373) );
  NOR2X0 U15957 ( .IN1(n15374), .IN2(CRC_OUT_7_15), .QN(n15371) );
  NAND2X0 U15958 ( .IN1(n15375), .IN2(n15376), .QN(n15374) );
  NAND2X0 U15959 ( .IN1(n9511), .IN2(CRC_OUT_7_31), .QN(n15376) );
  NAND2X0 U15960 ( .IN1(DFF_575_n1), .IN2(WX3453), .QN(n15375) );
  NOR2X0 U15961 ( .IN1(n10332), .IN2(n15377), .QN(WX3880) );
  NAND2X0 U15962 ( .IN1(n15378), .IN2(n15379), .QN(n15377) );
  INVX0 U15963 ( .INP(n15380), .ZN(n15379) );
  NOR2X0 U15964 ( .IN1(WX3455), .IN2(DFF_558_n1), .QN(n15380) );
  NAND2X0 U15965 ( .IN1(DFF_558_n1), .IN2(WX3455), .QN(n15378) );
  NOR2X0 U15966 ( .IN1(n10332), .IN2(n15381), .QN(WX3878) );
  NAND2X0 U15967 ( .IN1(n15382), .IN2(n15383), .QN(n15381) );
  INVX0 U15968 ( .INP(n15384), .ZN(n15383) );
  NOR2X0 U15969 ( .IN1(WX3457), .IN2(DFF_557_n1), .QN(n15384) );
  NAND2X0 U15970 ( .IN1(DFF_557_n1), .IN2(WX3457), .QN(n15382) );
  NOR2X0 U15971 ( .IN1(n10332), .IN2(n15385), .QN(WX3876) );
  NAND2X0 U15972 ( .IN1(n15386), .IN2(n15387), .QN(n15385) );
  INVX0 U15973 ( .INP(n15388), .ZN(n15387) );
  NOR2X0 U15974 ( .IN1(WX3459), .IN2(DFF_556_n1), .QN(n15388) );
  NAND2X0 U15975 ( .IN1(DFF_556_n1), .IN2(WX3459), .QN(n15386) );
  NOR2X0 U15976 ( .IN1(n10332), .IN2(n15389), .QN(WX3874) );
  NAND2X0 U15977 ( .IN1(n15390), .IN2(n15391), .QN(n15389) );
  INVX0 U15978 ( .INP(n15392), .ZN(n15391) );
  NOR2X0 U15979 ( .IN1(WX3461), .IN2(DFF_555_n1), .QN(n15392) );
  NAND2X0 U15980 ( .IN1(DFF_555_n1), .IN2(WX3461), .QN(n15390) );
  NOR2X0 U15981 ( .IN1(n10295), .IN2(n15393), .QN(WX3872) );
  NAND2X0 U15982 ( .IN1(n15394), .IN2(n15395), .QN(n15393) );
  INVX0 U15983 ( .INP(n15396), .ZN(n15395) );
  NOR2X0 U15984 ( .IN1(CRC_OUT_7_31), .IN2(n15397), .QN(n15396) );
  NAND2X0 U15985 ( .IN1(n15397), .IN2(CRC_OUT_7_31), .QN(n15394) );
  NAND2X0 U15986 ( .IN1(n15398), .IN2(n15399), .QN(n15397) );
  NAND2X0 U15987 ( .IN1(test_so31), .IN2(WX3463), .QN(n15399) );
  NAND2X0 U15988 ( .IN1(n9512), .IN2(n9871), .QN(n15398) );
  NOR2X0 U15989 ( .IN1(n10296), .IN2(n15400), .QN(WX3870) );
  NAND2X0 U15990 ( .IN1(n15401), .IN2(n15402), .QN(n15400) );
  INVX0 U15991 ( .INP(n15403), .ZN(n15402) );
  NOR2X0 U15992 ( .IN1(WX3465), .IN2(DFF_553_n1), .QN(n15403) );
  NAND2X0 U15993 ( .IN1(DFF_553_n1), .IN2(WX3465), .QN(n15401) );
  NOR2X0 U15994 ( .IN1(n10297), .IN2(n15404), .QN(WX3868) );
  NAND2X0 U15995 ( .IN1(n15405), .IN2(n15406), .QN(n15404) );
  INVX0 U15996 ( .INP(n15407), .ZN(n15406) );
  NOR2X0 U15997 ( .IN1(WX3467), .IN2(DFF_552_n1), .QN(n15407) );
  NAND2X0 U15998 ( .IN1(DFF_552_n1), .IN2(WX3467), .QN(n15405) );
  NOR2X0 U15999 ( .IN1(n10298), .IN2(n15408), .QN(WX3866) );
  NAND2X0 U16000 ( .IN1(n15409), .IN2(n15410), .QN(n15408) );
  INVX0 U16001 ( .INP(n15411), .ZN(n15410) );
  NOR2X0 U16002 ( .IN1(WX3469), .IN2(DFF_551_n1), .QN(n15411) );
  NAND2X0 U16003 ( .IN1(DFF_551_n1), .IN2(WX3469), .QN(n15409) );
  NOR2X0 U16004 ( .IN1(n10311), .IN2(n15412), .QN(WX3864) );
  NAND2X0 U16005 ( .IN1(n15413), .IN2(n15414), .QN(n15412) );
  INVX0 U16006 ( .INP(n15415), .ZN(n15414) );
  NOR2X0 U16007 ( .IN1(WX3471), .IN2(DFF_550_n1), .QN(n15415) );
  NAND2X0 U16008 ( .IN1(DFF_550_n1), .IN2(WX3471), .QN(n15413) );
  NOR2X0 U16009 ( .IN1(n10310), .IN2(n15416), .QN(WX3862) );
  NOR2X0 U16010 ( .IN1(n15417), .IN2(n15418), .QN(n15416) );
  INVX0 U16011 ( .INP(n15419), .ZN(n15418) );
  NAND2X0 U16012 ( .IN1(n9835), .IN2(DFF_549_n1), .QN(n15419) );
  NOR2X0 U16013 ( .IN1(DFF_549_n1), .IN2(n9835), .QN(n15417) );
  NOR2X0 U16014 ( .IN1(n10311), .IN2(n15420), .QN(WX3860) );
  NAND2X0 U16015 ( .IN1(n15421), .IN2(n15422), .QN(n15420) );
  INVX0 U16016 ( .INP(n15423), .ZN(n15422) );
  NOR2X0 U16017 ( .IN1(WX3475), .IN2(DFF_548_n1), .QN(n15423) );
  NAND2X0 U16018 ( .IN1(DFF_548_n1), .IN2(WX3475), .QN(n15421) );
  NOR2X0 U16019 ( .IN1(n10311), .IN2(n15424), .QN(WX3858) );
  NOR2X0 U16020 ( .IN1(n15425), .IN2(n15426), .QN(n15424) );
  INVX0 U16021 ( .INP(n15427), .ZN(n15426) );
  NAND2X0 U16022 ( .IN1(CRC_OUT_7_3), .IN2(n15428), .QN(n15427) );
  NOR2X0 U16023 ( .IN1(n15428), .IN2(CRC_OUT_7_3), .QN(n15425) );
  NAND2X0 U16024 ( .IN1(n15429), .IN2(n15430), .QN(n15428) );
  NAND2X0 U16025 ( .IN1(n9513), .IN2(CRC_OUT_7_31), .QN(n15430) );
  NAND2X0 U16026 ( .IN1(DFF_575_n1), .IN2(WX3477), .QN(n15429) );
  NOR2X0 U16027 ( .IN1(n10310), .IN2(n15431), .QN(WX3856) );
  NAND2X0 U16028 ( .IN1(n15432), .IN2(n15433), .QN(n15431) );
  INVX0 U16029 ( .INP(n15434), .ZN(n15433) );
  NOR2X0 U16030 ( .IN1(WX3479), .IN2(DFF_546_n1), .QN(n15434) );
  NAND2X0 U16031 ( .IN1(DFF_546_n1), .IN2(WX3479), .QN(n15432) );
  NOR2X0 U16032 ( .IN1(n10311), .IN2(n15435), .QN(WX3854) );
  NAND2X0 U16033 ( .IN1(n15436), .IN2(n15437), .QN(n15435) );
  INVX0 U16034 ( .INP(n15438), .ZN(n15437) );
  NOR2X0 U16035 ( .IN1(WX3481), .IN2(DFF_545_n1), .QN(n15438) );
  NAND2X0 U16036 ( .IN1(DFF_545_n1), .IN2(WX3481), .QN(n15436) );
  NOR2X0 U16037 ( .IN1(n10310), .IN2(n15439), .QN(WX3852) );
  NAND2X0 U16038 ( .IN1(n15440), .IN2(n15441), .QN(n15439) );
  INVX0 U16039 ( .INP(n15442), .ZN(n15441) );
  NOR2X0 U16040 ( .IN1(WX3483), .IN2(DFF_544_n1), .QN(n15442) );
  NAND2X0 U16041 ( .IN1(DFF_544_n1), .IN2(WX3483), .QN(n15440) );
  NOR2X0 U16042 ( .IN1(n10311), .IN2(n15443), .QN(WX3850) );
  NAND2X0 U16043 ( .IN1(n15444), .IN2(n15445), .QN(n15443) );
  NAND2X0 U16044 ( .IN1(n9523), .IN2(CRC_OUT_7_31), .QN(n15445) );
  NAND2X0 U16045 ( .IN1(DFF_575_n1), .IN2(WX3485), .QN(n15444) );
  NOR2X0 U16046 ( .IN1(n10311), .IN2(n9844), .QN(WX3324) );
  NOR2X0 U16047 ( .IN1(n18381), .IN2(n10242), .QN(WX3322) );
  NOR2X0 U16048 ( .IN1(n18380), .IN2(n10242), .QN(WX3320) );
  NOR2X0 U16049 ( .IN1(n18379), .IN2(n10242), .QN(WX3318) );
  NOR2X0 U16050 ( .IN1(n18378), .IN2(n10242), .QN(WX3316) );
  NOR2X0 U16051 ( .IN1(n18377), .IN2(n10242), .QN(WX3314) );
  NOR2X0 U16052 ( .IN1(n18376), .IN2(n10242), .QN(WX3312) );
  NOR2X0 U16053 ( .IN1(n18375), .IN2(n10242), .QN(WX3310) );
  NOR2X0 U16054 ( .IN1(n18374), .IN2(n10242), .QN(WX3308) );
  NOR2X0 U16055 ( .IN1(n18373), .IN2(n10242), .QN(WX3306) );
  NOR2X0 U16056 ( .IN1(n18372), .IN2(n10242), .QN(WX3304) );
  NOR2X0 U16057 ( .IN1(n18371), .IN2(n10242), .QN(WX3302) );
  NOR2X0 U16058 ( .IN1(n18370), .IN2(n10242), .QN(WX3300) );
  NOR2X0 U16059 ( .IN1(n18369), .IN2(n10241), .QN(WX3298) );
  NOR2X0 U16060 ( .IN1(n18368), .IN2(n10241), .QN(WX3296) );
  NOR2X0 U16061 ( .IN1(n18367), .IN2(n10241), .QN(WX3294) );
  NAND2X0 U16062 ( .IN1(n15446), .IN2(n15447), .QN(WX3292) );
  NOR2X0 U16063 ( .IN1(n15448), .IN2(n15449), .QN(n15447) );
  NOR2X0 U16064 ( .IN1(n15450), .IN2(n9939), .QN(n15449) );
  NOR2X0 U16065 ( .IN1(n9922), .IN2(n14620), .QN(n15448) );
  NAND2X0 U16066 ( .IN1(n15451), .IN2(n15452), .QN(n14620) );
  INVX0 U16067 ( .INP(n15453), .ZN(n15452) );
  NOR2X0 U16068 ( .IN1(n15454), .IN2(n15455), .QN(n15453) );
  NAND2X0 U16069 ( .IN1(n15455), .IN2(n15454), .QN(n15451) );
  NOR2X0 U16070 ( .IN1(n15456), .IN2(n15457), .QN(n15454) );
  INVX0 U16071 ( .INP(n15458), .ZN(n15457) );
  NAND2X0 U16072 ( .IN1(test_so36), .IN2(WX4778), .QN(n15458) );
  NOR2X0 U16073 ( .IN1(WX4778), .IN2(test_so36), .QN(n15456) );
  NAND2X0 U16074 ( .IN1(n15459), .IN2(n15460), .QN(n15455) );
  NAND2X0 U16075 ( .IN1(n9396), .IN2(WX4650), .QN(n15460) );
  INVX0 U16076 ( .INP(n15461), .ZN(n15459) );
  NOR2X0 U16077 ( .IN1(WX4650), .IN2(n9396), .QN(n15461) );
  NOR2X0 U16078 ( .IN1(n15462), .IN2(n15463), .QN(n15446) );
  NOR2X0 U16079 ( .IN1(DFF_544_n1), .IN2(n9971), .QN(n15463) );
  NOR2X0 U16080 ( .IN1(n9986), .IN2(n10679), .QN(n15462) );
  NAND2X0 U16081 ( .IN1(n10203), .IN2(n8612), .QN(n10679) );
  NAND2X0 U16082 ( .IN1(n15464), .IN2(n15465), .QN(WX3290) );
  NOR2X0 U16083 ( .IN1(n15466), .IN2(n15467), .QN(n15465) );
  NOR2X0 U16084 ( .IN1(n15468), .IN2(n9939), .QN(n15467) );
  NOR2X0 U16085 ( .IN1(n14642), .IN2(n9919), .QN(n15466) );
  INVX0 U16086 ( .INP(n15469), .ZN(n14642) );
  NAND2X0 U16087 ( .IN1(n15470), .IN2(n15471), .QN(n15469) );
  NAND2X0 U16088 ( .IN1(n15472), .IN2(n15473), .QN(n15471) );
  NAND2X0 U16089 ( .IN1(n15474), .IN2(n15475), .QN(n15473) );
  NAND2X0 U16090 ( .IN1(n9398), .IN2(WX4584), .QN(n15475) );
  NAND2X0 U16091 ( .IN1(n9397), .IN2(WX4712), .QN(n15474) );
  NOR2X0 U16092 ( .IN1(n15476), .IN2(n15477), .QN(n15472) );
  NOR2X0 U16093 ( .IN1(n9684), .IN2(WX4648), .QN(n15477) );
  NOR2X0 U16094 ( .IN1(n3693), .IN2(WX4776), .QN(n15476) );
  NAND2X0 U16095 ( .IN1(n15478), .IN2(n15479), .QN(n15470) );
  NAND2X0 U16096 ( .IN1(n15480), .IN2(n15481), .QN(n15479) );
  NAND2X0 U16097 ( .IN1(n9684), .IN2(WX4648), .QN(n15481) );
  NAND2X0 U16098 ( .IN1(n3693), .IN2(WX4776), .QN(n15480) );
  NOR2X0 U16099 ( .IN1(n15482), .IN2(n15483), .QN(n15478) );
  NOR2X0 U16100 ( .IN1(n9398), .IN2(WX4584), .QN(n15483) );
  NOR2X0 U16101 ( .IN1(n9397), .IN2(WX4712), .QN(n15482) );
  NOR2X0 U16102 ( .IN1(n15484), .IN2(n15485), .QN(n15464) );
  NOR2X0 U16103 ( .IN1(DFF_545_n1), .IN2(n9971), .QN(n15485) );
  NOR2X0 U16104 ( .IN1(n9986), .IN2(n10680), .QN(n15484) );
  NAND2X0 U16105 ( .IN1(n10203), .IN2(n8613), .QN(n10680) );
  NAND2X0 U16106 ( .IN1(n15486), .IN2(n15487), .QN(WX3288) );
  NOR2X0 U16107 ( .IN1(n15488), .IN2(n15489), .QN(n15487) );
  NOR2X0 U16108 ( .IN1(n15490), .IN2(n9939), .QN(n15489) );
  NOR2X0 U16109 ( .IN1(n14660), .IN2(n9919), .QN(n15488) );
  INVX0 U16110 ( .INP(n15491), .ZN(n14660) );
  NAND2X0 U16111 ( .IN1(n15492), .IN2(n15493), .QN(n15491) );
  NAND2X0 U16112 ( .IN1(n15494), .IN2(n15495), .QN(n15493) );
  NAND2X0 U16113 ( .IN1(n15496), .IN2(n15497), .QN(n15495) );
  NAND2X0 U16114 ( .IN1(n9400), .IN2(WX4582), .QN(n15497) );
  NAND2X0 U16115 ( .IN1(n9399), .IN2(WX4710), .QN(n15496) );
  NOR2X0 U16116 ( .IN1(n15498), .IN2(n15499), .QN(n15494) );
  NOR2X0 U16117 ( .IN1(n9683), .IN2(WX4646), .QN(n15499) );
  NOR2X0 U16118 ( .IN1(n3695), .IN2(WX4774), .QN(n15498) );
  NAND2X0 U16119 ( .IN1(n15500), .IN2(n15501), .QN(n15492) );
  NAND2X0 U16120 ( .IN1(n15502), .IN2(n15503), .QN(n15501) );
  NAND2X0 U16121 ( .IN1(n9683), .IN2(WX4646), .QN(n15503) );
  NAND2X0 U16122 ( .IN1(n3695), .IN2(WX4774), .QN(n15502) );
  NOR2X0 U16123 ( .IN1(n15504), .IN2(n15505), .QN(n15500) );
  NOR2X0 U16124 ( .IN1(n9400), .IN2(WX4582), .QN(n15505) );
  NOR2X0 U16125 ( .IN1(n9399), .IN2(WX4710), .QN(n15504) );
  NOR2X0 U16126 ( .IN1(n15506), .IN2(n15507), .QN(n15486) );
  NOR2X0 U16127 ( .IN1(DFF_546_n1), .IN2(n9971), .QN(n15507) );
  NOR2X0 U16128 ( .IN1(n9985), .IN2(n10681), .QN(n15506) );
  NAND2X0 U16129 ( .IN1(test_so23), .IN2(n10214), .QN(n10681) );
  NAND2X0 U16130 ( .IN1(n15508), .IN2(n15509), .QN(WX3286) );
  NOR2X0 U16131 ( .IN1(n15510), .IN2(n15511), .QN(n15509) );
  NOR2X0 U16132 ( .IN1(n15512), .IN2(n9938), .QN(n15511) );
  NOR2X0 U16133 ( .IN1(n14682), .IN2(n9918), .QN(n15510) );
  INVX0 U16134 ( .INP(n15513), .ZN(n14682) );
  NAND2X0 U16135 ( .IN1(n15514), .IN2(n15515), .QN(n15513) );
  NAND2X0 U16136 ( .IN1(n15516), .IN2(n15517), .QN(n15515) );
  NAND2X0 U16137 ( .IN1(n15518), .IN2(n15519), .QN(n15517) );
  NAND2X0 U16138 ( .IN1(n9402), .IN2(WX4580), .QN(n15519) );
  NAND2X0 U16139 ( .IN1(n9401), .IN2(WX4708), .QN(n15518) );
  NOR2X0 U16140 ( .IN1(n15520), .IN2(n15521), .QN(n15516) );
  NOR2X0 U16141 ( .IN1(n9682), .IN2(WX4644), .QN(n15521) );
  NOR2X0 U16142 ( .IN1(n3697), .IN2(WX4772), .QN(n15520) );
  NAND2X0 U16143 ( .IN1(n15522), .IN2(n15523), .QN(n15514) );
  NAND2X0 U16144 ( .IN1(n15524), .IN2(n15525), .QN(n15523) );
  NAND2X0 U16145 ( .IN1(n9682), .IN2(WX4644), .QN(n15525) );
  NAND2X0 U16146 ( .IN1(n3697), .IN2(WX4772), .QN(n15524) );
  NOR2X0 U16147 ( .IN1(n15526), .IN2(n15527), .QN(n15522) );
  NOR2X0 U16148 ( .IN1(n9402), .IN2(WX4580), .QN(n15527) );
  NOR2X0 U16149 ( .IN1(n9401), .IN2(WX4708), .QN(n15526) );
  NOR2X0 U16150 ( .IN1(n15528), .IN2(n15529), .QN(n15508) );
  NOR2X0 U16151 ( .IN1(DFF_547_n1), .IN2(n9971), .QN(n15529) );
  NOR2X0 U16152 ( .IN1(n9985), .IN2(n10682), .QN(n15528) );
  NAND2X0 U16153 ( .IN1(n10203), .IN2(n8616), .QN(n10682) );
  NAND2X0 U16154 ( .IN1(n15530), .IN2(n15531), .QN(WX3284) );
  NOR2X0 U16155 ( .IN1(n15532), .IN2(n15533), .QN(n15531) );
  NOR2X0 U16156 ( .IN1(n15534), .IN2(n9938), .QN(n15533) );
  NOR2X0 U16157 ( .IN1(n14700), .IN2(n9918), .QN(n15532) );
  INVX0 U16158 ( .INP(n15535), .ZN(n14700) );
  NAND2X0 U16159 ( .IN1(n15536), .IN2(n15537), .QN(n15535) );
  NAND2X0 U16160 ( .IN1(n15538), .IN2(n15539), .QN(n15537) );
  NAND2X0 U16161 ( .IN1(n15540), .IN2(n15541), .QN(n15539) );
  NAND2X0 U16162 ( .IN1(n9404), .IN2(WX4578), .QN(n15541) );
  NAND2X0 U16163 ( .IN1(n9403), .IN2(WX4706), .QN(n15540) );
  NOR2X0 U16164 ( .IN1(n15542), .IN2(n15543), .QN(n15538) );
  NOR2X0 U16165 ( .IN1(n9510), .IN2(WX4642), .QN(n15543) );
  NOR2X0 U16166 ( .IN1(n3699), .IN2(WX4770), .QN(n15542) );
  NAND2X0 U16167 ( .IN1(n15544), .IN2(n15545), .QN(n15536) );
  NAND2X0 U16168 ( .IN1(n15546), .IN2(n15547), .QN(n15545) );
  NAND2X0 U16169 ( .IN1(n9510), .IN2(WX4642), .QN(n15547) );
  NAND2X0 U16170 ( .IN1(n3699), .IN2(WX4770), .QN(n15546) );
  NOR2X0 U16171 ( .IN1(n15548), .IN2(n15549), .QN(n15544) );
  NOR2X0 U16172 ( .IN1(n9404), .IN2(WX4578), .QN(n15549) );
  NOR2X0 U16173 ( .IN1(n9403), .IN2(WX4706), .QN(n15548) );
  NOR2X0 U16174 ( .IN1(n15550), .IN2(n15551), .QN(n15530) );
  NOR2X0 U16175 ( .IN1(DFF_548_n1), .IN2(n9971), .QN(n15551) );
  NOR2X0 U16176 ( .IN1(n9985), .IN2(n10683), .QN(n15550) );
  NAND2X0 U16177 ( .IN1(n10203), .IN2(n8617), .QN(n10683) );
  NAND2X0 U16178 ( .IN1(n15552), .IN2(n15553), .QN(WX3282) );
  NOR2X0 U16179 ( .IN1(n15554), .IN2(n15555), .QN(n15553) );
  NOR2X0 U16180 ( .IN1(n15556), .IN2(n9938), .QN(n15555) );
  NOR2X0 U16181 ( .IN1(n14722), .IN2(n9918), .QN(n15554) );
  INVX0 U16182 ( .INP(n15557), .ZN(n14722) );
  NAND2X0 U16183 ( .IN1(n15558), .IN2(n15559), .QN(n15557) );
  NAND2X0 U16184 ( .IN1(n15560), .IN2(n15561), .QN(n15559) );
  NAND2X0 U16185 ( .IN1(n15562), .IN2(n15563), .QN(n15561) );
  NAND2X0 U16186 ( .IN1(n9406), .IN2(WX4576), .QN(n15563) );
  NAND2X0 U16187 ( .IN1(n9405), .IN2(WX4704), .QN(n15562) );
  NOR2X0 U16188 ( .IN1(n15564), .IN2(n15565), .QN(n15560) );
  NOR2X0 U16189 ( .IN1(n9681), .IN2(WX4640), .QN(n15565) );
  NOR2X0 U16190 ( .IN1(n3701), .IN2(WX4768), .QN(n15564) );
  NAND2X0 U16191 ( .IN1(n15566), .IN2(n15567), .QN(n15558) );
  NAND2X0 U16192 ( .IN1(n15568), .IN2(n15569), .QN(n15567) );
  NAND2X0 U16193 ( .IN1(n9681), .IN2(WX4640), .QN(n15569) );
  NAND2X0 U16194 ( .IN1(n3701), .IN2(WX4768), .QN(n15568) );
  NOR2X0 U16195 ( .IN1(n15570), .IN2(n15571), .QN(n15566) );
  NOR2X0 U16196 ( .IN1(n9406), .IN2(WX4576), .QN(n15571) );
  NOR2X0 U16197 ( .IN1(n9405), .IN2(WX4704), .QN(n15570) );
  NOR2X0 U16198 ( .IN1(n15572), .IN2(n15573), .QN(n15552) );
  NOR2X0 U16199 ( .IN1(DFF_549_n1), .IN2(n9971), .QN(n15573) );
  NOR2X0 U16200 ( .IN1(n9985), .IN2(n10684), .QN(n15572) );
  NAND2X0 U16201 ( .IN1(n10203), .IN2(n8618), .QN(n10684) );
  NAND2X0 U16202 ( .IN1(n15574), .IN2(n15575), .QN(WX3280) );
  NOR2X0 U16203 ( .IN1(n15576), .IN2(n15577), .QN(n15575) );
  NOR2X0 U16204 ( .IN1(n9943), .IN2(n15578), .QN(n15577) );
  NOR2X0 U16205 ( .IN1(n14740), .IN2(n9918), .QN(n15576) );
  INVX0 U16206 ( .INP(n15579), .ZN(n14740) );
  NAND2X0 U16207 ( .IN1(n15580), .IN2(n15581), .QN(n15579) );
  NAND2X0 U16208 ( .IN1(n15582), .IN2(n15583), .QN(n15581) );
  NAND2X0 U16209 ( .IN1(n15584), .IN2(n15585), .QN(n15583) );
  NAND2X0 U16210 ( .IN1(n9408), .IN2(WX4574), .QN(n15585) );
  NAND2X0 U16211 ( .IN1(n9407), .IN2(WX4702), .QN(n15584) );
  NOR2X0 U16212 ( .IN1(n15586), .IN2(n15587), .QN(n15582) );
  NOR2X0 U16213 ( .IN1(n9680), .IN2(WX4638), .QN(n15587) );
  NOR2X0 U16214 ( .IN1(n3703), .IN2(WX4766), .QN(n15586) );
  NAND2X0 U16215 ( .IN1(n15588), .IN2(n15589), .QN(n15580) );
  NAND2X0 U16216 ( .IN1(n15590), .IN2(n15591), .QN(n15589) );
  NAND2X0 U16217 ( .IN1(n9680), .IN2(WX4638), .QN(n15591) );
  NAND2X0 U16218 ( .IN1(n3703), .IN2(WX4766), .QN(n15590) );
  NOR2X0 U16219 ( .IN1(n15592), .IN2(n15593), .QN(n15588) );
  NOR2X0 U16220 ( .IN1(n9408), .IN2(WX4574), .QN(n15593) );
  NOR2X0 U16221 ( .IN1(n9407), .IN2(WX4702), .QN(n15592) );
  NOR2X0 U16222 ( .IN1(n15594), .IN2(n15595), .QN(n15574) );
  NOR2X0 U16223 ( .IN1(DFF_550_n1), .IN2(n9971), .QN(n15595) );
  NOR2X0 U16224 ( .IN1(n9985), .IN2(n10685), .QN(n15594) );
  NAND2X0 U16225 ( .IN1(n10203), .IN2(n8619), .QN(n10685) );
  NAND2X0 U16226 ( .IN1(n15596), .IN2(n15597), .QN(WX3278) );
  NOR2X0 U16227 ( .IN1(n15598), .IN2(n15599), .QN(n15597) );
  NOR2X0 U16228 ( .IN1(n15600), .IN2(n9938), .QN(n15599) );
  NOR2X0 U16229 ( .IN1(n14762), .IN2(n9918), .QN(n15598) );
  INVX0 U16230 ( .INP(n15601), .ZN(n14762) );
  NAND2X0 U16231 ( .IN1(n15602), .IN2(n15603), .QN(n15601) );
  NAND2X0 U16232 ( .IN1(n15604), .IN2(n15605), .QN(n15603) );
  NAND2X0 U16233 ( .IN1(n15606), .IN2(n15607), .QN(n15605) );
  NAND2X0 U16234 ( .IN1(n9410), .IN2(WX4572), .QN(n15607) );
  NAND2X0 U16235 ( .IN1(n9409), .IN2(WX4700), .QN(n15606) );
  NOR2X0 U16236 ( .IN1(n15608), .IN2(n15609), .QN(n15604) );
  NOR2X0 U16237 ( .IN1(n9679), .IN2(WX4636), .QN(n15609) );
  NOR2X0 U16238 ( .IN1(n3705), .IN2(WX4764), .QN(n15608) );
  NAND2X0 U16239 ( .IN1(n15610), .IN2(n15611), .QN(n15602) );
  NAND2X0 U16240 ( .IN1(n15612), .IN2(n15613), .QN(n15611) );
  NAND2X0 U16241 ( .IN1(n9679), .IN2(WX4636), .QN(n15613) );
  NAND2X0 U16242 ( .IN1(n3705), .IN2(WX4764), .QN(n15612) );
  NOR2X0 U16243 ( .IN1(n15614), .IN2(n15615), .QN(n15610) );
  NOR2X0 U16244 ( .IN1(n9410), .IN2(WX4572), .QN(n15615) );
  NOR2X0 U16245 ( .IN1(n9409), .IN2(WX4700), .QN(n15614) );
  NOR2X0 U16246 ( .IN1(n15616), .IN2(n15617), .QN(n15596) );
  NOR2X0 U16247 ( .IN1(DFF_551_n1), .IN2(n9971), .QN(n15617) );
  NOR2X0 U16248 ( .IN1(n9985), .IN2(n10686), .QN(n15616) );
  NAND2X0 U16249 ( .IN1(n10203), .IN2(n8620), .QN(n10686) );
  NAND2X0 U16250 ( .IN1(n15618), .IN2(n15619), .QN(WX3276) );
  NOR2X0 U16251 ( .IN1(n15620), .IN2(n15621), .QN(n15619) );
  NOR2X0 U16252 ( .IN1(n9941), .IN2(n15622), .QN(n15621) );
  NOR2X0 U16253 ( .IN1(n14784), .IN2(n9918), .QN(n15620) );
  INVX0 U16254 ( .INP(n15623), .ZN(n14784) );
  NAND2X0 U16255 ( .IN1(n15624), .IN2(n15625), .QN(n15623) );
  NAND2X0 U16256 ( .IN1(n15626), .IN2(n15627), .QN(n15625) );
  NAND2X0 U16257 ( .IN1(n15628), .IN2(n15629), .QN(n15627) );
  NAND2X0 U16258 ( .IN1(n9412), .IN2(WX4570), .QN(n15629) );
  NAND2X0 U16259 ( .IN1(n9411), .IN2(WX4698), .QN(n15628) );
  NOR2X0 U16260 ( .IN1(n15630), .IN2(n15631), .QN(n15626) );
  NOR2X0 U16261 ( .IN1(n9678), .IN2(WX4634), .QN(n15631) );
  NOR2X0 U16262 ( .IN1(n3707), .IN2(WX4762), .QN(n15630) );
  NAND2X0 U16263 ( .IN1(n15632), .IN2(n15633), .QN(n15624) );
  NAND2X0 U16264 ( .IN1(n15634), .IN2(n15635), .QN(n15633) );
  NAND2X0 U16265 ( .IN1(n9678), .IN2(WX4634), .QN(n15635) );
  NAND2X0 U16266 ( .IN1(n3707), .IN2(WX4762), .QN(n15634) );
  NOR2X0 U16267 ( .IN1(n15636), .IN2(n15637), .QN(n15632) );
  NOR2X0 U16268 ( .IN1(n9412), .IN2(WX4570), .QN(n15637) );
  NOR2X0 U16269 ( .IN1(n9411), .IN2(WX4698), .QN(n15636) );
  NOR2X0 U16270 ( .IN1(n15638), .IN2(n15639), .QN(n15618) );
  NOR2X0 U16271 ( .IN1(DFF_552_n1), .IN2(n9971), .QN(n15639) );
  NOR2X0 U16272 ( .IN1(n9985), .IN2(n10687), .QN(n15638) );
  NAND2X0 U16273 ( .IN1(n10203), .IN2(n8621), .QN(n10687) );
  NAND2X0 U16274 ( .IN1(n15640), .IN2(n15641), .QN(WX3274) );
  NOR2X0 U16275 ( .IN1(n15642), .IN2(n15643), .QN(n15641) );
  NOR2X0 U16276 ( .IN1(n15644), .IN2(n9938), .QN(n15643) );
  NOR2X0 U16277 ( .IN1(n14806), .IN2(n9918), .QN(n15642) );
  INVX0 U16278 ( .INP(n15645), .ZN(n14806) );
  NAND2X0 U16279 ( .IN1(n15646), .IN2(n15647), .QN(n15645) );
  NAND2X0 U16280 ( .IN1(n15648), .IN2(n15649), .QN(n15647) );
  NAND2X0 U16281 ( .IN1(n15650), .IN2(n15651), .QN(n15649) );
  NAND2X0 U16282 ( .IN1(n9414), .IN2(WX4568), .QN(n15651) );
  NAND2X0 U16283 ( .IN1(n9413), .IN2(WX4696), .QN(n15650) );
  NOR2X0 U16284 ( .IN1(n15652), .IN2(n15653), .QN(n15648) );
  NOR2X0 U16285 ( .IN1(n9677), .IN2(WX4632), .QN(n15653) );
  NOR2X0 U16286 ( .IN1(n3709), .IN2(WX4760), .QN(n15652) );
  NAND2X0 U16287 ( .IN1(n15654), .IN2(n15655), .QN(n15646) );
  NAND2X0 U16288 ( .IN1(n15656), .IN2(n15657), .QN(n15655) );
  NAND2X0 U16289 ( .IN1(n9677), .IN2(WX4632), .QN(n15657) );
  NAND2X0 U16290 ( .IN1(n3709), .IN2(WX4760), .QN(n15656) );
  NOR2X0 U16291 ( .IN1(n15658), .IN2(n15659), .QN(n15654) );
  NOR2X0 U16292 ( .IN1(n9414), .IN2(WX4568), .QN(n15659) );
  NOR2X0 U16293 ( .IN1(n9413), .IN2(WX4696), .QN(n15658) );
  NOR2X0 U16294 ( .IN1(n15660), .IN2(n15661), .QN(n15640) );
  NOR2X0 U16295 ( .IN1(DFF_553_n1), .IN2(n9971), .QN(n15661) );
  NOR2X0 U16296 ( .IN1(n9985), .IN2(n10698), .QN(n15660) );
  NAND2X0 U16297 ( .IN1(n10203), .IN2(n8622), .QN(n10698) );
  NAND2X0 U16298 ( .IN1(n15662), .IN2(n15663), .QN(WX3272) );
  NOR2X0 U16299 ( .IN1(n15664), .IN2(n15665), .QN(n15663) );
  NOR2X0 U16300 ( .IN1(n15666), .IN2(n9938), .QN(n15665) );
  NOR2X0 U16301 ( .IN1(n14828), .IN2(n9918), .QN(n15664) );
  INVX0 U16302 ( .INP(n15667), .ZN(n14828) );
  NAND2X0 U16303 ( .IN1(n15668), .IN2(n15669), .QN(n15667) );
  NAND2X0 U16304 ( .IN1(n15670), .IN2(n15671), .QN(n15669) );
  NAND2X0 U16305 ( .IN1(n15672), .IN2(n15673), .QN(n15671) );
  NAND2X0 U16306 ( .IN1(n9416), .IN2(WX4566), .QN(n15673) );
  NAND2X0 U16307 ( .IN1(n9415), .IN2(WX4694), .QN(n15672) );
  NOR2X0 U16308 ( .IN1(n15674), .IN2(n15675), .QN(n15670) );
  NOR2X0 U16309 ( .IN1(n9676), .IN2(WX4630), .QN(n15675) );
  NOR2X0 U16310 ( .IN1(n3711), .IN2(WX4758), .QN(n15674) );
  NAND2X0 U16311 ( .IN1(n15676), .IN2(n15677), .QN(n15668) );
  NAND2X0 U16312 ( .IN1(n15678), .IN2(n15679), .QN(n15677) );
  NAND2X0 U16313 ( .IN1(n9676), .IN2(WX4630), .QN(n15679) );
  NAND2X0 U16314 ( .IN1(n3711), .IN2(WX4758), .QN(n15678) );
  NOR2X0 U16315 ( .IN1(n15680), .IN2(n15681), .QN(n15676) );
  NOR2X0 U16316 ( .IN1(n9416), .IN2(WX4566), .QN(n15681) );
  NOR2X0 U16317 ( .IN1(n9415), .IN2(WX4694), .QN(n15680) );
  NOR2X0 U16318 ( .IN1(n15682), .IN2(n15683), .QN(n15662) );
  NOR2X0 U16319 ( .IN1(n9975), .IN2(n9871), .QN(n15683) );
  NOR2X0 U16320 ( .IN1(n9985), .IN2(n10699), .QN(n15682) );
  NAND2X0 U16321 ( .IN1(n10202), .IN2(n8623), .QN(n10699) );
  NAND2X0 U16322 ( .IN1(n15684), .IN2(n15685), .QN(WX3270) );
  NOR2X0 U16323 ( .IN1(n15686), .IN2(n15687), .QN(n15685) );
  NOR2X0 U16324 ( .IN1(n15688), .IN2(n9938), .QN(n15687) );
  NOR2X0 U16325 ( .IN1(n9921), .IN2(n14850), .QN(n15686) );
  NAND2X0 U16326 ( .IN1(n15689), .IN2(n15690), .QN(n14850) );
  INVX0 U16327 ( .INP(n15691), .ZN(n15690) );
  NOR2X0 U16328 ( .IN1(n15692), .IN2(n15693), .QN(n15691) );
  NAND2X0 U16329 ( .IN1(n15693), .IN2(n15692), .QN(n15689) );
  NOR2X0 U16330 ( .IN1(n15694), .IN2(n15695), .QN(n15692) );
  NOR2X0 U16331 ( .IN1(n9850), .IN2(n9418), .QN(n15695) );
  INVX0 U16332 ( .INP(n15696), .ZN(n15694) );
  NAND2X0 U16333 ( .IN1(n9418), .IN2(n9850), .QN(n15696) );
  NAND2X0 U16334 ( .IN1(n15697), .IN2(n15698), .QN(n15693) );
  NAND2X0 U16335 ( .IN1(n9417), .IN2(WX4628), .QN(n15698) );
  INVX0 U16336 ( .INP(n15699), .ZN(n15697) );
  NOR2X0 U16337 ( .IN1(WX4628), .IN2(n9417), .QN(n15699) );
  NOR2X0 U16338 ( .IN1(n15700), .IN2(n15701), .QN(n15684) );
  NOR2X0 U16339 ( .IN1(DFF_555_n1), .IN2(n9971), .QN(n15701) );
  NOR2X0 U16340 ( .IN1(n9985), .IN2(n10700), .QN(n15700) );
  NAND2X0 U16341 ( .IN1(n10202), .IN2(n8624), .QN(n10700) );
  NAND2X0 U16342 ( .IN1(n15702), .IN2(n15703), .QN(WX3268) );
  NOR2X0 U16343 ( .IN1(n15704), .IN2(n15705), .QN(n15703) );
  NOR2X0 U16344 ( .IN1(n9941), .IN2(n15706), .QN(n15705) );
  NOR2X0 U16345 ( .IN1(n14872), .IN2(n9918), .QN(n15704) );
  INVX0 U16346 ( .INP(n15707), .ZN(n14872) );
  NAND2X0 U16347 ( .IN1(n15708), .IN2(n15709), .QN(n15707) );
  NAND2X0 U16348 ( .IN1(n15710), .IN2(n15711), .QN(n15709) );
  NAND2X0 U16349 ( .IN1(n15712), .IN2(n15713), .QN(n15711) );
  NAND2X0 U16350 ( .IN1(n9420), .IN2(WX4562), .QN(n15713) );
  NAND2X0 U16351 ( .IN1(n9419), .IN2(WX4690), .QN(n15712) );
  NOR2X0 U16352 ( .IN1(n15714), .IN2(n15715), .QN(n15710) );
  NOR2X0 U16353 ( .IN1(n9675), .IN2(WX4626), .QN(n15715) );
  NOR2X0 U16354 ( .IN1(n3715), .IN2(WX4754), .QN(n15714) );
  NAND2X0 U16355 ( .IN1(n15716), .IN2(n15717), .QN(n15708) );
  NAND2X0 U16356 ( .IN1(n15718), .IN2(n15719), .QN(n15717) );
  NAND2X0 U16357 ( .IN1(n9675), .IN2(WX4626), .QN(n15719) );
  NAND2X0 U16358 ( .IN1(n3715), .IN2(WX4754), .QN(n15718) );
  NOR2X0 U16359 ( .IN1(n15720), .IN2(n15721), .QN(n15716) );
  NOR2X0 U16360 ( .IN1(n9420), .IN2(WX4562), .QN(n15721) );
  NOR2X0 U16361 ( .IN1(n9419), .IN2(WX4690), .QN(n15720) );
  NOR2X0 U16362 ( .IN1(n15722), .IN2(n15723), .QN(n15702) );
  NOR2X0 U16363 ( .IN1(DFF_556_n1), .IN2(n9970), .QN(n15723) );
  NOR2X0 U16364 ( .IN1(n9985), .IN2(n10701), .QN(n15722) );
  NAND2X0 U16365 ( .IN1(n10202), .IN2(n8625), .QN(n10701) );
  NAND2X0 U16366 ( .IN1(n15724), .IN2(n15725), .QN(WX3266) );
  NOR2X0 U16367 ( .IN1(n15726), .IN2(n15727), .QN(n15725) );
  NOR2X0 U16368 ( .IN1(n15728), .IN2(n9938), .QN(n15727) );
  NOR2X0 U16369 ( .IN1(n9923), .IN2(n14894), .QN(n15726) );
  NAND2X0 U16370 ( .IN1(n15729), .IN2(n15730), .QN(n14894) );
  INVX0 U16371 ( .INP(n15731), .ZN(n15730) );
  NOR2X0 U16372 ( .IN1(n15732), .IN2(n15733), .QN(n15731) );
  NAND2X0 U16373 ( .IN1(n15733), .IN2(n15732), .QN(n15729) );
  NOR2X0 U16374 ( .IN1(n15734), .IN2(n15735), .QN(n15732) );
  INVX0 U16375 ( .INP(n15736), .ZN(n15735) );
  NAND2X0 U16376 ( .IN1(test_so39), .IN2(WX4752), .QN(n15736) );
  NOR2X0 U16377 ( .IN1(WX4752), .IN2(test_so39), .QN(n15734) );
  NAND2X0 U16378 ( .IN1(n15737), .IN2(n15738), .QN(n15733) );
  NAND2X0 U16379 ( .IN1(n9421), .IN2(WX4624), .QN(n15738) );
  INVX0 U16380 ( .INP(n15739), .ZN(n15737) );
  NOR2X0 U16381 ( .IN1(WX4624), .IN2(n9421), .QN(n15739) );
  NOR2X0 U16382 ( .IN1(n15740), .IN2(n15741), .QN(n15724) );
  NOR2X0 U16383 ( .IN1(DFF_557_n1), .IN2(n9970), .QN(n15741) );
  NOR2X0 U16384 ( .IN1(n9985), .IN2(n10702), .QN(n15740) );
  NAND2X0 U16385 ( .IN1(n10202), .IN2(n8626), .QN(n10702) );
  NAND2X0 U16386 ( .IN1(n15742), .IN2(n15743), .QN(WX3264) );
  NOR2X0 U16387 ( .IN1(n15744), .IN2(n15745), .QN(n15743) );
  NOR2X0 U16388 ( .IN1(n15746), .IN2(n9938), .QN(n15745) );
  NOR2X0 U16389 ( .IN1(n14916), .IN2(n9918), .QN(n15744) );
  INVX0 U16390 ( .INP(n15747), .ZN(n14916) );
  NAND2X0 U16391 ( .IN1(n15748), .IN2(n15749), .QN(n15747) );
  NAND2X0 U16392 ( .IN1(n15750), .IN2(n15751), .QN(n15749) );
  NAND2X0 U16393 ( .IN1(n15752), .IN2(n15753), .QN(n15751) );
  NAND2X0 U16394 ( .IN1(n9423), .IN2(WX4558), .QN(n15753) );
  NAND2X0 U16395 ( .IN1(n9422), .IN2(WX4686), .QN(n15752) );
  NOR2X0 U16396 ( .IN1(n15754), .IN2(n15755), .QN(n15750) );
  NOR2X0 U16397 ( .IN1(n9673), .IN2(WX4622), .QN(n15755) );
  NOR2X0 U16398 ( .IN1(n3719), .IN2(WX4750), .QN(n15754) );
  NAND2X0 U16399 ( .IN1(n15756), .IN2(n15757), .QN(n15748) );
  NAND2X0 U16400 ( .IN1(n15758), .IN2(n15759), .QN(n15757) );
  NAND2X0 U16401 ( .IN1(n9673), .IN2(WX4622), .QN(n15759) );
  NAND2X0 U16402 ( .IN1(n3719), .IN2(WX4750), .QN(n15758) );
  NOR2X0 U16403 ( .IN1(n15760), .IN2(n15761), .QN(n15756) );
  NOR2X0 U16404 ( .IN1(n9423), .IN2(WX4558), .QN(n15761) );
  NOR2X0 U16405 ( .IN1(n9422), .IN2(WX4686), .QN(n15760) );
  NOR2X0 U16406 ( .IN1(n15762), .IN2(n15763), .QN(n15742) );
  NOR2X0 U16407 ( .IN1(DFF_558_n1), .IN2(n9970), .QN(n15763) );
  NOR2X0 U16408 ( .IN1(n9984), .IN2(n10703), .QN(n15762) );
  NAND2X0 U16409 ( .IN1(n10202), .IN2(n8627), .QN(n10703) );
  NAND2X0 U16410 ( .IN1(n15764), .IN2(n15765), .QN(WX3262) );
  NOR2X0 U16411 ( .IN1(n15766), .IN2(n15767), .QN(n15765) );
  NOR2X0 U16412 ( .IN1(n15768), .IN2(n9938), .QN(n15767) );
  NOR2X0 U16413 ( .IN1(n9921), .IN2(n14938), .QN(n15766) );
  NAND2X0 U16414 ( .IN1(n15769), .IN2(n15770), .QN(n14938) );
  INVX0 U16415 ( .INP(n15771), .ZN(n15770) );
  NOR2X0 U16416 ( .IN1(n15772), .IN2(n15773), .QN(n15771) );
  NAND2X0 U16417 ( .IN1(n15773), .IN2(n15772), .QN(n15769) );
  NOR2X0 U16418 ( .IN1(n15774), .IN2(n15775), .QN(n15772) );
  INVX0 U16419 ( .INP(n15776), .ZN(n15775) );
  NAND2X0 U16420 ( .IN1(test_so37), .IN2(WX4748), .QN(n15776) );
  NOR2X0 U16421 ( .IN1(WX4748), .IN2(test_so37), .QN(n15774) );
  NAND2X0 U16422 ( .IN1(n15777), .IN2(n15778), .QN(n15773) );
  NAND2X0 U16423 ( .IN1(n9425), .IN2(WX4556), .QN(n15778) );
  INVX0 U16424 ( .INP(n15779), .ZN(n15777) );
  NOR2X0 U16425 ( .IN1(WX4556), .IN2(n9425), .QN(n15779) );
  NOR2X0 U16426 ( .IN1(n15780), .IN2(n15781), .QN(n15764) );
  NOR2X0 U16427 ( .IN1(DFF_559_n1), .IN2(n9970), .QN(n15781) );
  NOR2X0 U16428 ( .IN1(n9984), .IN2(n10704), .QN(n15780) );
  NAND2X0 U16429 ( .IN1(n10202), .IN2(n8628), .QN(n10704) );
  NAND2X0 U16430 ( .IN1(n15782), .IN2(n15783), .QN(WX3260) );
  NOR2X0 U16431 ( .IN1(n15784), .IN2(n15785), .QN(n15783) );
  NOR2X0 U16432 ( .IN1(n9942), .IN2(n15786), .QN(n15785) );
  NOR2X0 U16433 ( .IN1(n14960), .IN2(n9918), .QN(n15784) );
  NOR2X0 U16434 ( .IN1(n15787), .IN2(n15788), .QN(n14960) );
  INVX0 U16435 ( .INP(n15789), .ZN(n15788) );
  NAND2X0 U16436 ( .IN1(n15790), .IN2(n15791), .QN(n15789) );
  NOR2X0 U16437 ( .IN1(n15791), .IN2(n15790), .QN(n15787) );
  NAND2X0 U16438 ( .IN1(n15792), .IN2(n15793), .QN(n15790) );
  NAND2X0 U16439 ( .IN1(n9160), .IN2(n15794), .QN(n15793) );
  INVX0 U16440 ( .INP(n15795), .ZN(n15792) );
  NOR2X0 U16441 ( .IN1(n15794), .IN2(n9160), .QN(n15795) );
  NOR2X0 U16442 ( .IN1(n15796), .IN2(n15797), .QN(n15794) );
  INVX0 U16443 ( .INP(n15798), .ZN(n15797) );
  NAND2X0 U16444 ( .IN1(n18396), .IN2(WX4746), .QN(n15798) );
  NOR2X0 U16445 ( .IN1(WX4746), .IN2(n18396), .QN(n15796) );
  NOR2X0 U16446 ( .IN1(n15799), .IN2(n15800), .QN(n15791) );
  INVX0 U16447 ( .INP(n15801), .ZN(n15800) );
  NAND2X0 U16448 ( .IN1(n9159), .IN2(n10020), .QN(n15801) );
  NOR2X0 U16449 ( .IN1(n10009), .IN2(n9159), .QN(n15799) );
  NOR2X0 U16450 ( .IN1(n15802), .IN2(n15803), .QN(n15782) );
  NOR2X0 U16451 ( .IN1(DFF_560_n1), .IN2(n9970), .QN(n15803) );
  NOR2X0 U16452 ( .IN1(n9984), .IN2(n10705), .QN(n15802) );
  NAND2X0 U16453 ( .IN1(n10202), .IN2(n8629), .QN(n10705) );
  NAND2X0 U16454 ( .IN1(n15804), .IN2(n15805), .QN(WX3258) );
  NOR2X0 U16455 ( .IN1(n15806), .IN2(n15807), .QN(n15805) );
  NOR2X0 U16456 ( .IN1(n15808), .IN2(n9938), .QN(n15807) );
  NOR2X0 U16457 ( .IN1(n9922), .IN2(n14983), .QN(n15806) );
  NAND2X0 U16458 ( .IN1(n15809), .IN2(n15810), .QN(n14983) );
  INVX0 U16459 ( .INP(n15811), .ZN(n15810) );
  NOR2X0 U16460 ( .IN1(n15812), .IN2(n15813), .QN(n15811) );
  NAND2X0 U16461 ( .IN1(n15813), .IN2(n15812), .QN(n15809) );
  INVX0 U16462 ( .INP(n15814), .ZN(n15812) );
  NAND2X0 U16463 ( .IN1(n15815), .IN2(n15816), .QN(n15814) );
  NAND2X0 U16464 ( .IN1(n15817), .IN2(WX4680), .QN(n15816) );
  NAND2X0 U16465 ( .IN1(n15818), .IN2(n15819), .QN(n15817) );
  NAND2X0 U16466 ( .IN1(test_so35), .IN2(WX4616), .QN(n15819) );
  NAND2X0 U16467 ( .IN1(n9161), .IN2(n9843), .QN(n15818) );
  NAND2X0 U16468 ( .IN1(n9162), .IN2(n15820), .QN(n15815) );
  NOR2X0 U16469 ( .IN1(n15821), .IN2(n15822), .QN(n15820) );
  NOR2X0 U16470 ( .IN1(test_so35), .IN2(WX4616), .QN(n15822) );
  NOR2X0 U16471 ( .IN1(n9161), .IN2(n9843), .QN(n15821) );
  NAND2X0 U16472 ( .IN1(n15823), .IN2(n15824), .QN(n15813) );
  NAND2X0 U16473 ( .IN1(n9671), .IN2(n10020), .QN(n15824) );
  NAND2X0 U16474 ( .IN1(TM1), .IN2(WX4744), .QN(n15823) );
  NOR2X0 U16475 ( .IN1(n15825), .IN2(n15826), .QN(n15804) );
  NOR2X0 U16476 ( .IN1(DFF_561_n1), .IN2(n9970), .QN(n15826) );
  NOR2X0 U16477 ( .IN1(n9984), .IN2(n10706), .QN(n15825) );
  NAND2X0 U16478 ( .IN1(n10202), .IN2(n8630), .QN(n10706) );
  NAND2X0 U16479 ( .IN1(n15827), .IN2(n15828), .QN(WX3256) );
  NOR2X0 U16480 ( .IN1(n15829), .IN2(n15830), .QN(n15828) );
  NOR2X0 U16481 ( .IN1(n15831), .IN2(n9938), .QN(n15830) );
  NOR2X0 U16482 ( .IN1(n15005), .IN2(n9918), .QN(n15829) );
  NOR2X0 U16483 ( .IN1(n15832), .IN2(n15833), .QN(n15005) );
  INVX0 U16484 ( .INP(n15834), .ZN(n15833) );
  NAND2X0 U16485 ( .IN1(n15835), .IN2(n15836), .QN(n15834) );
  NOR2X0 U16486 ( .IN1(n15836), .IN2(n15835), .QN(n15832) );
  NAND2X0 U16487 ( .IN1(n15837), .IN2(n15838), .QN(n15835) );
  NAND2X0 U16488 ( .IN1(n9164), .IN2(n15839), .QN(n15838) );
  INVX0 U16489 ( .INP(n15840), .ZN(n15837) );
  NOR2X0 U16490 ( .IN1(n15839), .IN2(n9164), .QN(n15840) );
  NOR2X0 U16491 ( .IN1(n15841), .IN2(n15842), .QN(n15839) );
  INVX0 U16492 ( .INP(n15843), .ZN(n15842) );
  NAND2X0 U16493 ( .IN1(n18395), .IN2(WX4742), .QN(n15843) );
  NOR2X0 U16494 ( .IN1(WX4742), .IN2(n18395), .QN(n15841) );
  NOR2X0 U16495 ( .IN1(n15844), .IN2(n15845), .QN(n15836) );
  INVX0 U16496 ( .INP(n15846), .ZN(n15845) );
  NAND2X0 U16497 ( .IN1(n9163), .IN2(n10020), .QN(n15846) );
  NOR2X0 U16498 ( .IN1(n10009), .IN2(n9163), .QN(n15844) );
  NOR2X0 U16499 ( .IN1(n15847), .IN2(n15848), .QN(n15827) );
  NOR2X0 U16500 ( .IN1(DFF_562_n1), .IN2(n9970), .QN(n15848) );
  NOR2X0 U16501 ( .IN1(n9984), .IN2(n10707), .QN(n15847) );
  NAND2X0 U16502 ( .IN1(n10202), .IN2(n8631), .QN(n10707) );
  NAND2X0 U16503 ( .IN1(n15849), .IN2(n15850), .QN(WX3254) );
  NOR2X0 U16504 ( .IN1(n15851), .IN2(n15852), .QN(n15850) );
  NOR2X0 U16505 ( .IN1(n15853), .IN2(n9937), .QN(n15852) );
  NOR2X0 U16506 ( .IN1(n15027), .IN2(n9917), .QN(n15851) );
  NOR2X0 U16507 ( .IN1(n15854), .IN2(n15855), .QN(n15027) );
  INVX0 U16508 ( .INP(n15856), .ZN(n15855) );
  NAND2X0 U16509 ( .IN1(n15857), .IN2(n15858), .QN(n15856) );
  NOR2X0 U16510 ( .IN1(n15858), .IN2(n15857), .QN(n15854) );
  NAND2X0 U16511 ( .IN1(n15859), .IN2(n15860), .QN(n15857) );
  NAND2X0 U16512 ( .IN1(n9166), .IN2(n15861), .QN(n15860) );
  INVX0 U16513 ( .INP(n15862), .ZN(n15859) );
  NOR2X0 U16514 ( .IN1(n15861), .IN2(n9166), .QN(n15862) );
  NOR2X0 U16515 ( .IN1(n15863), .IN2(n15864), .QN(n15861) );
  INVX0 U16516 ( .INP(n15865), .ZN(n15864) );
  NAND2X0 U16517 ( .IN1(n18394), .IN2(WX4740), .QN(n15865) );
  NOR2X0 U16518 ( .IN1(WX4740), .IN2(n18394), .QN(n15863) );
  NOR2X0 U16519 ( .IN1(n15866), .IN2(n15867), .QN(n15858) );
  INVX0 U16520 ( .INP(n15868), .ZN(n15867) );
  NAND2X0 U16521 ( .IN1(n9165), .IN2(n10020), .QN(n15868) );
  NOR2X0 U16522 ( .IN1(n10009), .IN2(n9165), .QN(n15866) );
  NOR2X0 U16523 ( .IN1(n15869), .IN2(n15870), .QN(n15849) );
  NOR2X0 U16524 ( .IN1(DFF_563_n1), .IN2(n9970), .QN(n15870) );
  NOR2X0 U16525 ( .IN1(n9984), .IN2(n10708), .QN(n15869) );
  NAND2X0 U16526 ( .IN1(n10201), .IN2(n8632), .QN(n10708) );
  NAND2X0 U16527 ( .IN1(n15871), .IN2(n15872), .QN(WX3252) );
  NOR2X0 U16528 ( .IN1(n15873), .IN2(n15874), .QN(n15872) );
  NOR2X0 U16529 ( .IN1(n15875), .IN2(n9937), .QN(n15874) );
  NOR2X0 U16530 ( .IN1(n15049), .IN2(n9917), .QN(n15873) );
  NOR2X0 U16531 ( .IN1(n15876), .IN2(n15877), .QN(n15049) );
  INVX0 U16532 ( .INP(n15878), .ZN(n15877) );
  NAND2X0 U16533 ( .IN1(n15879), .IN2(n15880), .QN(n15878) );
  NOR2X0 U16534 ( .IN1(n15880), .IN2(n15879), .QN(n15876) );
  NAND2X0 U16535 ( .IN1(n15881), .IN2(n15882), .QN(n15879) );
  NAND2X0 U16536 ( .IN1(n9168), .IN2(n15883), .QN(n15882) );
  INVX0 U16537 ( .INP(n15884), .ZN(n15881) );
  NOR2X0 U16538 ( .IN1(n15883), .IN2(n9168), .QN(n15884) );
  NOR2X0 U16539 ( .IN1(n15885), .IN2(n15886), .QN(n15883) );
  INVX0 U16540 ( .INP(n15887), .ZN(n15886) );
  NAND2X0 U16541 ( .IN1(n18393), .IN2(WX4738), .QN(n15887) );
  NOR2X0 U16542 ( .IN1(WX4738), .IN2(n18393), .QN(n15885) );
  NOR2X0 U16543 ( .IN1(n15888), .IN2(n15889), .QN(n15880) );
  INVX0 U16544 ( .INP(n15890), .ZN(n15889) );
  NAND2X0 U16545 ( .IN1(n9167), .IN2(n10020), .QN(n15890) );
  NOR2X0 U16546 ( .IN1(n10009), .IN2(n9167), .QN(n15888) );
  NOR2X0 U16547 ( .IN1(n15891), .IN2(n15892), .QN(n15871) );
  NOR2X0 U16548 ( .IN1(DFF_564_n1), .IN2(n9970), .QN(n15892) );
  NOR2X0 U16549 ( .IN1(n9984), .IN2(n10709), .QN(n15891) );
  NAND2X0 U16550 ( .IN1(test_so22), .IN2(n10214), .QN(n10709) );
  NAND2X0 U16551 ( .IN1(n15893), .IN2(n15894), .QN(WX3250) );
  NOR2X0 U16552 ( .IN1(n15895), .IN2(n15896), .QN(n15894) );
  NOR2X0 U16553 ( .IN1(n15897), .IN2(n9937), .QN(n15896) );
  NOR2X0 U16554 ( .IN1(n15071), .IN2(n9917), .QN(n15895) );
  NOR2X0 U16555 ( .IN1(n15898), .IN2(n15899), .QN(n15071) );
  INVX0 U16556 ( .INP(n15900), .ZN(n15899) );
  NAND2X0 U16557 ( .IN1(n15901), .IN2(n15902), .QN(n15900) );
  NOR2X0 U16558 ( .IN1(n15902), .IN2(n15901), .QN(n15898) );
  NAND2X0 U16559 ( .IN1(n15903), .IN2(n15904), .QN(n15901) );
  NAND2X0 U16560 ( .IN1(n9170), .IN2(n15905), .QN(n15904) );
  INVX0 U16561 ( .INP(n15906), .ZN(n15903) );
  NOR2X0 U16562 ( .IN1(n15905), .IN2(n9170), .QN(n15906) );
  NOR2X0 U16563 ( .IN1(n15907), .IN2(n15908), .QN(n15905) );
  INVX0 U16564 ( .INP(n15909), .ZN(n15908) );
  NAND2X0 U16565 ( .IN1(n18392), .IN2(WX4736), .QN(n15909) );
  NOR2X0 U16566 ( .IN1(WX4736), .IN2(n18392), .QN(n15907) );
  NOR2X0 U16567 ( .IN1(n15910), .IN2(n15911), .QN(n15902) );
  INVX0 U16568 ( .INP(n15912), .ZN(n15911) );
  NAND2X0 U16569 ( .IN1(n9169), .IN2(n10020), .QN(n15912) );
  NOR2X0 U16570 ( .IN1(n10009), .IN2(n9169), .QN(n15910) );
  NOR2X0 U16571 ( .IN1(n15913), .IN2(n15914), .QN(n15893) );
  NOR2X0 U16572 ( .IN1(DFF_565_n1), .IN2(n9970), .QN(n15914) );
  NOR2X0 U16573 ( .IN1(n9984), .IN2(n10710), .QN(n15913) );
  NAND2X0 U16574 ( .IN1(n10201), .IN2(n8635), .QN(n10710) );
  NAND2X0 U16575 ( .IN1(n15915), .IN2(n15916), .QN(WX3248) );
  NOR2X0 U16576 ( .IN1(n15917), .IN2(n15918), .QN(n15916) );
  NOR2X0 U16577 ( .IN1(n15919), .IN2(n9937), .QN(n15918) );
  NOR2X0 U16578 ( .IN1(n15093), .IN2(n9917), .QN(n15917) );
  NOR2X0 U16579 ( .IN1(n15920), .IN2(n15921), .QN(n15093) );
  INVX0 U16580 ( .INP(n15922), .ZN(n15921) );
  NAND2X0 U16581 ( .IN1(n15923), .IN2(n15924), .QN(n15922) );
  NOR2X0 U16582 ( .IN1(n15924), .IN2(n15923), .QN(n15920) );
  NAND2X0 U16583 ( .IN1(n15925), .IN2(n15926), .QN(n15923) );
  NAND2X0 U16584 ( .IN1(n9172), .IN2(n15927), .QN(n15926) );
  INVX0 U16585 ( .INP(n15928), .ZN(n15925) );
  NOR2X0 U16586 ( .IN1(n15927), .IN2(n9172), .QN(n15928) );
  NOR2X0 U16587 ( .IN1(n15929), .IN2(n15930), .QN(n15927) );
  INVX0 U16588 ( .INP(n15931), .ZN(n15930) );
  NAND2X0 U16589 ( .IN1(n18391), .IN2(WX4734), .QN(n15931) );
  NOR2X0 U16590 ( .IN1(WX4734), .IN2(n18391), .QN(n15929) );
  NOR2X0 U16591 ( .IN1(n15932), .IN2(n15933), .QN(n15924) );
  INVX0 U16592 ( .INP(n15934), .ZN(n15933) );
  NAND2X0 U16593 ( .IN1(n9171), .IN2(n10020), .QN(n15934) );
  NOR2X0 U16594 ( .IN1(n10009), .IN2(n9171), .QN(n15932) );
  NOR2X0 U16595 ( .IN1(n15935), .IN2(n15936), .QN(n15915) );
  NOR2X0 U16596 ( .IN1(DFF_566_n1), .IN2(n9970), .QN(n15936) );
  NOR2X0 U16597 ( .IN1(n9984), .IN2(n10711), .QN(n15935) );
  NAND2X0 U16598 ( .IN1(n10201), .IN2(n8636), .QN(n10711) );
  NAND2X0 U16599 ( .IN1(n15937), .IN2(n15938), .QN(WX3246) );
  NOR2X0 U16600 ( .IN1(n15939), .IN2(n15940), .QN(n15938) );
  NOR2X0 U16601 ( .IN1(n9943), .IN2(n15941), .QN(n15940) );
  NOR2X0 U16602 ( .IN1(n15116), .IN2(n9917), .QN(n15939) );
  NOR2X0 U16603 ( .IN1(n15942), .IN2(n15943), .QN(n15116) );
  INVX0 U16604 ( .INP(n15944), .ZN(n15943) );
  NAND2X0 U16605 ( .IN1(n15945), .IN2(n15946), .QN(n15944) );
  NOR2X0 U16606 ( .IN1(n15946), .IN2(n15945), .QN(n15942) );
  NAND2X0 U16607 ( .IN1(n15947), .IN2(n15948), .QN(n15945) );
  NAND2X0 U16608 ( .IN1(n9174), .IN2(n15949), .QN(n15948) );
  INVX0 U16609 ( .INP(n15950), .ZN(n15947) );
  NOR2X0 U16610 ( .IN1(n15949), .IN2(n9174), .QN(n15950) );
  NOR2X0 U16611 ( .IN1(n15951), .IN2(n15952), .QN(n15949) );
  INVX0 U16612 ( .INP(n15953), .ZN(n15952) );
  NAND2X0 U16613 ( .IN1(n18390), .IN2(WX4732), .QN(n15953) );
  NOR2X0 U16614 ( .IN1(WX4732), .IN2(n18390), .QN(n15951) );
  NOR2X0 U16615 ( .IN1(n15954), .IN2(n15955), .QN(n15946) );
  INVX0 U16616 ( .INP(n15956), .ZN(n15955) );
  NAND2X0 U16617 ( .IN1(n9173), .IN2(n10020), .QN(n15956) );
  NOR2X0 U16618 ( .IN1(n10009), .IN2(n9173), .QN(n15954) );
  NOR2X0 U16619 ( .IN1(n15957), .IN2(n15958), .QN(n15937) );
  NOR2X0 U16620 ( .IN1(DFF_567_n1), .IN2(n9970), .QN(n15958) );
  NOR2X0 U16621 ( .IN1(n9984), .IN2(n10712), .QN(n15957) );
  NAND2X0 U16622 ( .IN1(n10201), .IN2(n8637), .QN(n10712) );
  NAND2X0 U16623 ( .IN1(n15959), .IN2(n15960), .QN(WX3244) );
  NOR2X0 U16624 ( .IN1(n15961), .IN2(n15962), .QN(n15960) );
  NOR2X0 U16625 ( .IN1(n15963), .IN2(n9937), .QN(n15962) );
  NOR2X0 U16626 ( .IN1(n15138), .IN2(n9917), .QN(n15961) );
  NOR2X0 U16627 ( .IN1(n15964), .IN2(n15965), .QN(n15138) );
  INVX0 U16628 ( .INP(n15966), .ZN(n15965) );
  NAND2X0 U16629 ( .IN1(n15967), .IN2(n15968), .QN(n15966) );
  NOR2X0 U16630 ( .IN1(n15968), .IN2(n15967), .QN(n15964) );
  NAND2X0 U16631 ( .IN1(n15969), .IN2(n15970), .QN(n15967) );
  NAND2X0 U16632 ( .IN1(n9176), .IN2(n15971), .QN(n15970) );
  INVX0 U16633 ( .INP(n15972), .ZN(n15969) );
  NOR2X0 U16634 ( .IN1(n15971), .IN2(n9176), .QN(n15972) );
  NOR2X0 U16635 ( .IN1(n15973), .IN2(n15974), .QN(n15971) );
  INVX0 U16636 ( .INP(n15975), .ZN(n15974) );
  NAND2X0 U16637 ( .IN1(n18389), .IN2(WX4730), .QN(n15975) );
  NOR2X0 U16638 ( .IN1(WX4730), .IN2(n18389), .QN(n15973) );
  NOR2X0 U16639 ( .IN1(n15976), .IN2(n15977), .QN(n15968) );
  INVX0 U16640 ( .INP(n15978), .ZN(n15977) );
  NAND2X0 U16641 ( .IN1(n9175), .IN2(n10020), .QN(n15978) );
  NOR2X0 U16642 ( .IN1(n10009), .IN2(n9175), .QN(n15976) );
  NOR2X0 U16643 ( .IN1(n15979), .IN2(n15980), .QN(n15959) );
  NOR2X0 U16644 ( .IN1(DFF_568_n1), .IN2(n9969), .QN(n15980) );
  NOR2X0 U16645 ( .IN1(n9984), .IN2(n10713), .QN(n15979) );
  NAND2X0 U16646 ( .IN1(n10201), .IN2(n8638), .QN(n10713) );
  NAND2X0 U16647 ( .IN1(n15981), .IN2(n15982), .QN(WX3242) );
  NOR2X0 U16648 ( .IN1(n15983), .IN2(n15984), .QN(n15982) );
  NOR2X0 U16649 ( .IN1(n15985), .IN2(n9937), .QN(n15984) );
  NOR2X0 U16650 ( .IN1(n15160), .IN2(n9917), .QN(n15983) );
  NOR2X0 U16651 ( .IN1(n15986), .IN2(n15987), .QN(n15160) );
  INVX0 U16652 ( .INP(n15988), .ZN(n15987) );
  NAND2X0 U16653 ( .IN1(n15989), .IN2(n15990), .QN(n15988) );
  NOR2X0 U16654 ( .IN1(n15990), .IN2(n15989), .QN(n15986) );
  NAND2X0 U16655 ( .IN1(n15991), .IN2(n15992), .QN(n15989) );
  NAND2X0 U16656 ( .IN1(n9178), .IN2(n15993), .QN(n15992) );
  INVX0 U16657 ( .INP(n15994), .ZN(n15991) );
  NOR2X0 U16658 ( .IN1(n15993), .IN2(n9178), .QN(n15994) );
  NOR2X0 U16659 ( .IN1(n15995), .IN2(n15996), .QN(n15993) );
  INVX0 U16660 ( .INP(n15997), .ZN(n15996) );
  NAND2X0 U16661 ( .IN1(n18388), .IN2(WX4728), .QN(n15997) );
  NOR2X0 U16662 ( .IN1(WX4728), .IN2(n18388), .QN(n15995) );
  NOR2X0 U16663 ( .IN1(n15998), .IN2(n15999), .QN(n15990) );
  INVX0 U16664 ( .INP(n16000), .ZN(n15999) );
  NAND2X0 U16665 ( .IN1(n9177), .IN2(n10020), .QN(n16000) );
  NOR2X0 U16666 ( .IN1(n10009), .IN2(n9177), .QN(n15998) );
  NOR2X0 U16667 ( .IN1(n16001), .IN2(n16002), .QN(n15981) );
  NOR2X0 U16668 ( .IN1(DFF_569_n1), .IN2(n9969), .QN(n16002) );
  NOR2X0 U16669 ( .IN1(n9984), .IN2(n10714), .QN(n16001) );
  NAND2X0 U16670 ( .IN1(n10201), .IN2(n8639), .QN(n10714) );
  NAND2X0 U16671 ( .IN1(n16003), .IN2(n16004), .QN(WX3240) );
  NOR2X0 U16672 ( .IN1(n16005), .IN2(n16006), .QN(n16004) );
  NOR2X0 U16673 ( .IN1(n9942), .IN2(n16007), .QN(n16006) );
  NOR2X0 U16674 ( .IN1(n15182), .IN2(n9917), .QN(n16005) );
  NOR2X0 U16675 ( .IN1(n16008), .IN2(n16009), .QN(n15182) );
  INVX0 U16676 ( .INP(n16010), .ZN(n16009) );
  NAND2X0 U16677 ( .IN1(n16011), .IN2(n16012), .QN(n16010) );
  NOR2X0 U16678 ( .IN1(n16012), .IN2(n16011), .QN(n16008) );
  NAND2X0 U16679 ( .IN1(n16013), .IN2(n16014), .QN(n16011) );
  NAND2X0 U16680 ( .IN1(n9180), .IN2(n16015), .QN(n16014) );
  INVX0 U16681 ( .INP(n16016), .ZN(n16013) );
  NOR2X0 U16682 ( .IN1(n16015), .IN2(n9180), .QN(n16016) );
  NOR2X0 U16683 ( .IN1(n16017), .IN2(n16018), .QN(n16015) );
  INVX0 U16684 ( .INP(n16019), .ZN(n16018) );
  NAND2X0 U16685 ( .IN1(n18387), .IN2(WX4726), .QN(n16019) );
  NOR2X0 U16686 ( .IN1(WX4726), .IN2(n18387), .QN(n16017) );
  NOR2X0 U16687 ( .IN1(n16020), .IN2(n16021), .QN(n16012) );
  INVX0 U16688 ( .INP(n16022), .ZN(n16021) );
  NAND2X0 U16689 ( .IN1(n9179), .IN2(n10020), .QN(n16022) );
  NOR2X0 U16690 ( .IN1(n10009), .IN2(n9179), .QN(n16020) );
  NOR2X0 U16691 ( .IN1(n16023), .IN2(n16024), .QN(n16003) );
  NOR2X0 U16692 ( .IN1(DFF_570_n1), .IN2(n9969), .QN(n16024) );
  NOR2X0 U16693 ( .IN1(n9983), .IN2(n10715), .QN(n16023) );
  NAND2X0 U16694 ( .IN1(n10201), .IN2(n8640), .QN(n10715) );
  NAND2X0 U16695 ( .IN1(n16025), .IN2(n16026), .QN(WX3238) );
  NOR2X0 U16696 ( .IN1(n16027), .IN2(n16028), .QN(n16026) );
  NOR2X0 U16697 ( .IN1(n16029), .IN2(n9937), .QN(n16028) );
  NOR2X0 U16698 ( .IN1(n15204), .IN2(n9917), .QN(n16027) );
  NOR2X0 U16699 ( .IN1(n16030), .IN2(n16031), .QN(n15204) );
  INVX0 U16700 ( .INP(n16032), .ZN(n16031) );
  NAND2X0 U16701 ( .IN1(n16033), .IN2(n16034), .QN(n16032) );
  NOR2X0 U16702 ( .IN1(n16034), .IN2(n16033), .QN(n16030) );
  NAND2X0 U16703 ( .IN1(n16035), .IN2(n16036), .QN(n16033) );
  NAND2X0 U16704 ( .IN1(n9182), .IN2(n16037), .QN(n16036) );
  INVX0 U16705 ( .INP(n16038), .ZN(n16035) );
  NOR2X0 U16706 ( .IN1(n16037), .IN2(n9182), .QN(n16038) );
  NOR2X0 U16707 ( .IN1(n16039), .IN2(n16040), .QN(n16037) );
  INVX0 U16708 ( .INP(n16041), .ZN(n16040) );
  NAND2X0 U16709 ( .IN1(n18386), .IN2(WX4724), .QN(n16041) );
  NOR2X0 U16710 ( .IN1(WX4724), .IN2(n18386), .QN(n16039) );
  NOR2X0 U16711 ( .IN1(n16042), .IN2(n16043), .QN(n16034) );
  INVX0 U16712 ( .INP(n16044), .ZN(n16043) );
  NAND2X0 U16713 ( .IN1(n9181), .IN2(n10020), .QN(n16044) );
  NOR2X0 U16714 ( .IN1(n10010), .IN2(n9181), .QN(n16042) );
  NOR2X0 U16715 ( .IN1(n16045), .IN2(n16046), .QN(n16025) );
  NOR2X0 U16716 ( .IN1(n9975), .IN2(n9860), .QN(n16046) );
  NOR2X0 U16717 ( .IN1(n9983), .IN2(n10716), .QN(n16045) );
  NAND2X0 U16718 ( .IN1(n10201), .IN2(n8641), .QN(n10716) );
  NAND2X0 U16719 ( .IN1(n16047), .IN2(n16048), .QN(WX3236) );
  NOR2X0 U16720 ( .IN1(n16049), .IN2(n16050), .QN(n16048) );
  NOR2X0 U16721 ( .IN1(n16051), .IN2(n9937), .QN(n16050) );
  NOR2X0 U16722 ( .IN1(n9922), .IN2(n15226), .QN(n16049) );
  NAND2X0 U16723 ( .IN1(n16052), .IN2(n16053), .QN(n15226) );
  NAND2X0 U16724 ( .IN1(n16054), .IN2(n16055), .QN(n16053) );
  INVX0 U16725 ( .INP(n16056), .ZN(n16052) );
  NOR2X0 U16726 ( .IN1(n16055), .IN2(n16054), .QN(n16056) );
  NAND2X0 U16727 ( .IN1(n16057), .IN2(n16058), .QN(n16054) );
  NAND2X0 U16728 ( .IN1(n16059), .IN2(WX4658), .QN(n16058) );
  NAND2X0 U16729 ( .IN1(n16060), .IN2(n16061), .QN(n16059) );
  NAND2X0 U16730 ( .IN1(test_so40), .IN2(WX4594), .QN(n16061) );
  NAND2X0 U16731 ( .IN1(n9183), .IN2(n9830), .QN(n16060) );
  NAND2X0 U16732 ( .IN1(n9184), .IN2(n16062), .QN(n16057) );
  NOR2X0 U16733 ( .IN1(n16063), .IN2(n16064), .QN(n16062) );
  NOR2X0 U16734 ( .IN1(test_so40), .IN2(WX4594), .QN(n16064) );
  NOR2X0 U16735 ( .IN1(n9183), .IN2(n9830), .QN(n16063) );
  NOR2X0 U16736 ( .IN1(n16065), .IN2(n16066), .QN(n16055) );
  INVX0 U16737 ( .INP(n16067), .ZN(n16066) );
  NAND2X0 U16738 ( .IN1(n18385), .IN2(n10020), .QN(n16067) );
  NOR2X0 U16739 ( .IN1(n10010), .IN2(n18385), .QN(n16065) );
  NOR2X0 U16740 ( .IN1(n16068), .IN2(n16069), .QN(n16047) );
  NOR2X0 U16741 ( .IN1(DFF_572_n1), .IN2(n9969), .QN(n16069) );
  NOR2X0 U16742 ( .IN1(n9983), .IN2(n10717), .QN(n16068) );
  NAND2X0 U16743 ( .IN1(n10201), .IN2(n8642), .QN(n10717) );
  NAND2X0 U16744 ( .IN1(n16070), .IN2(n16071), .QN(WX3234) );
  NOR2X0 U16745 ( .IN1(n16072), .IN2(n16073), .QN(n16071) );
  NOR2X0 U16746 ( .IN1(n16074), .IN2(n9937), .QN(n16073) );
  NOR2X0 U16747 ( .IN1(n15248), .IN2(n9917), .QN(n16072) );
  NOR2X0 U16748 ( .IN1(n16075), .IN2(n16076), .QN(n15248) );
  INVX0 U16749 ( .INP(n16077), .ZN(n16076) );
  NAND2X0 U16750 ( .IN1(n16078), .IN2(n16079), .QN(n16077) );
  NOR2X0 U16751 ( .IN1(n16079), .IN2(n16078), .QN(n16075) );
  NAND2X0 U16752 ( .IN1(n16080), .IN2(n16081), .QN(n16078) );
  NAND2X0 U16753 ( .IN1(n9186), .IN2(n16082), .QN(n16081) );
  INVX0 U16754 ( .INP(n16083), .ZN(n16080) );
  NOR2X0 U16755 ( .IN1(n16082), .IN2(n9186), .QN(n16083) );
  NOR2X0 U16756 ( .IN1(n16084), .IN2(n16085), .QN(n16082) );
  INVX0 U16757 ( .INP(n16086), .ZN(n16085) );
  NAND2X0 U16758 ( .IN1(n18384), .IN2(WX4720), .QN(n16086) );
  NOR2X0 U16759 ( .IN1(WX4720), .IN2(n18384), .QN(n16084) );
  NOR2X0 U16760 ( .IN1(n16087), .IN2(n16088), .QN(n16079) );
  INVX0 U16761 ( .INP(n16089), .ZN(n16088) );
  NAND2X0 U16762 ( .IN1(n9185), .IN2(n10021), .QN(n16089) );
  NOR2X0 U16763 ( .IN1(n10010), .IN2(n9185), .QN(n16087) );
  NOR2X0 U16764 ( .IN1(n16090), .IN2(n16091), .QN(n16070) );
  NOR2X0 U16765 ( .IN1(DFF_573_n1), .IN2(n9969), .QN(n16091) );
  NOR2X0 U16766 ( .IN1(n9983), .IN2(n10718), .QN(n16090) );
  NAND2X0 U16767 ( .IN1(n10200), .IN2(n8643), .QN(n10718) );
  NAND2X0 U16768 ( .IN1(n16092), .IN2(n16093), .QN(WX3232) );
  NOR2X0 U16769 ( .IN1(n16094), .IN2(n16095), .QN(n16093) );
  NOR2X0 U16770 ( .IN1(n9942), .IN2(n16096), .QN(n16095) );
  NOR2X0 U16771 ( .IN1(n9923), .IN2(n15270), .QN(n16094) );
  NAND2X0 U16772 ( .IN1(n16097), .IN2(n16098), .QN(n15270) );
  INVX0 U16773 ( .INP(n16099), .ZN(n16098) );
  NOR2X0 U16774 ( .IN1(n16100), .IN2(n16101), .QN(n16099) );
  NAND2X0 U16775 ( .IN1(n16101), .IN2(n16100), .QN(n16097) );
  NOR2X0 U16776 ( .IN1(n16102), .IN2(n16103), .QN(n16100) );
  INVX0 U16777 ( .INP(n16104), .ZN(n16103) );
  NAND2X0 U16778 ( .IN1(n9659), .IN2(n16105), .QN(n16104) );
  NOR2X0 U16779 ( .IN1(n16105), .IN2(n9659), .QN(n16102) );
  NOR2X0 U16780 ( .IN1(n16106), .IN2(n16107), .QN(n16105) );
  INVX0 U16781 ( .INP(n16108), .ZN(n16107) );
  NAND2X0 U16782 ( .IN1(test_so38), .IN2(n8552), .QN(n16108) );
  NOR2X0 U16783 ( .IN1(n8552), .IN2(test_so38), .QN(n16106) );
  NAND2X0 U16784 ( .IN1(n16109), .IN2(n16110), .QN(n16101) );
  NAND2X0 U16785 ( .IN1(n9187), .IN2(n10021), .QN(n16110) );
  INVX0 U16786 ( .INP(n16111), .ZN(n16109) );
  NOR2X0 U16787 ( .IN1(n10010), .IN2(n9187), .QN(n16111) );
  NOR2X0 U16788 ( .IN1(n16112), .IN2(n16113), .QN(n16092) );
  NOR2X0 U16789 ( .IN1(DFF_574_n1), .IN2(n9969), .QN(n16113) );
  NOR2X0 U16790 ( .IN1(n9983), .IN2(n10719), .QN(n16112) );
  NAND2X0 U16791 ( .IN1(n10200), .IN2(n8644), .QN(n10719) );
  NAND2X0 U16792 ( .IN1(n16114), .IN2(n16115), .QN(WX3230) );
  NOR2X0 U16793 ( .IN1(n16116), .IN2(n16117), .QN(n16115) );
  NOR2X0 U16794 ( .IN1(n16118), .IN2(n9937), .QN(n16117) );
  NOR2X0 U16795 ( .IN1(n15292), .IN2(n9917), .QN(n16116) );
  NOR2X0 U16796 ( .IN1(n16119), .IN2(n16120), .QN(n15292) );
  INVX0 U16797 ( .INP(n16121), .ZN(n16120) );
  NAND2X0 U16798 ( .IN1(n16122), .IN2(n16123), .QN(n16121) );
  NOR2X0 U16799 ( .IN1(n16123), .IN2(n16122), .QN(n16119) );
  NAND2X0 U16800 ( .IN1(n16124), .IN2(n16125), .QN(n16122) );
  NAND2X0 U16801 ( .IN1(n9014), .IN2(n16126), .QN(n16125) );
  INVX0 U16802 ( .INP(n16127), .ZN(n16124) );
  NOR2X0 U16803 ( .IN1(n16126), .IN2(n9014), .QN(n16127) );
  NOR2X0 U16804 ( .IN1(n16128), .IN2(n16129), .QN(n16126) );
  INVX0 U16805 ( .INP(n16130), .ZN(n16129) );
  NAND2X0 U16806 ( .IN1(n18382), .IN2(WX4716), .QN(n16130) );
  NOR2X0 U16807 ( .IN1(WX4716), .IN2(n18382), .QN(n16128) );
  NOR2X0 U16808 ( .IN1(n16131), .IN2(n16132), .QN(n16123) );
  INVX0 U16809 ( .INP(n16133), .ZN(n16132) );
  NAND2X0 U16810 ( .IN1(n9013), .IN2(n10013), .QN(n16133) );
  NOR2X0 U16811 ( .IN1(n10010), .IN2(n9013), .QN(n16131) );
  NOR2X0 U16812 ( .IN1(n16134), .IN2(n16135), .QN(n16114) );
  NOR2X0 U16813 ( .IN1(n9494), .IN2(n11994), .QN(n16135) );
  NOR2X0 U16814 ( .IN1(DFF_575_n1), .IN2(n9969), .QN(n16134) );
  INVX0 U16815 ( .INP(n16136), .ZN(WX3132) );
  NAND2X0 U16816 ( .IN1(n10200), .IN2(n9494), .QN(n16136) );
  NOR2X0 U16817 ( .IN1(n10309), .IN2(n16137), .QN(WX2619) );
  NAND2X0 U16818 ( .IN1(n16138), .IN2(n16139), .QN(n16137) );
  INVX0 U16819 ( .INP(n16140), .ZN(n16139) );
  NOR2X0 U16820 ( .IN1(WX2130), .IN2(DFF_382_n1), .QN(n16140) );
  NAND2X0 U16821 ( .IN1(DFF_382_n1), .IN2(WX2130), .QN(n16138) );
  NOR2X0 U16822 ( .IN1(n10308), .IN2(n16141), .QN(WX2617) );
  NAND2X0 U16823 ( .IN1(n16142), .IN2(n16143), .QN(n16141) );
  INVX0 U16824 ( .INP(n16144), .ZN(n16143) );
  NOR2X0 U16825 ( .IN1(WX2132), .IN2(DFF_381_n1), .QN(n16144) );
  NAND2X0 U16826 ( .IN1(DFF_381_n1), .IN2(WX2132), .QN(n16142) );
  NOR2X0 U16827 ( .IN1(n10308), .IN2(n16145), .QN(WX2615) );
  NAND2X0 U16828 ( .IN1(n16146), .IN2(n16147), .QN(n16145) );
  INVX0 U16829 ( .INP(n16148), .ZN(n16147) );
  NOR2X0 U16830 ( .IN1(WX2134), .IN2(DFF_380_n1), .QN(n16148) );
  NAND2X0 U16831 ( .IN1(DFF_380_n1), .IN2(WX2134), .QN(n16146) );
  NOR2X0 U16832 ( .IN1(n10309), .IN2(n16149), .QN(WX2613) );
  NOR2X0 U16833 ( .IN1(n16150), .IN2(n16151), .QN(n16149) );
  INVX0 U16834 ( .INP(n16152), .ZN(n16151) );
  NAND2X0 U16835 ( .IN1(n9832), .IN2(DFF_379_n1), .QN(n16152) );
  NOR2X0 U16836 ( .IN1(DFF_379_n1), .IN2(n9832), .QN(n16150) );
  NOR2X0 U16837 ( .IN1(n10308), .IN2(n16153), .QN(WX2611) );
  NAND2X0 U16838 ( .IN1(n16154), .IN2(n16155), .QN(n16153) );
  INVX0 U16839 ( .INP(n16156), .ZN(n16155) );
  NOR2X0 U16840 ( .IN1(WX2138), .IN2(DFF_378_n1), .QN(n16156) );
  NAND2X0 U16841 ( .IN1(DFF_378_n1), .IN2(WX2138), .QN(n16154) );
  NOR2X0 U16842 ( .IN1(n10308), .IN2(n16157), .QN(WX2609) );
  NOR2X0 U16843 ( .IN1(n16158), .IN2(n16159), .QN(n16157) );
  NOR2X0 U16844 ( .IN1(test_so21), .IN2(WX2140), .QN(n16159) );
  NOR2X0 U16845 ( .IN1(n9715), .IN2(n9862), .QN(n16158) );
  NOR2X0 U16846 ( .IN1(n10310), .IN2(n16160), .QN(WX2607) );
  NAND2X0 U16847 ( .IN1(n16161), .IN2(n16162), .QN(n16160) );
  INVX0 U16848 ( .INP(n16163), .ZN(n16162) );
  NOR2X0 U16849 ( .IN1(WX2142), .IN2(DFF_376_n1), .QN(n16163) );
  NAND2X0 U16850 ( .IN1(DFF_376_n1), .IN2(WX2142), .QN(n16161) );
  NOR2X0 U16851 ( .IN1(n10310), .IN2(n16164), .QN(WX2605) );
  NAND2X0 U16852 ( .IN1(n16165), .IN2(n16166), .QN(n16164) );
  INVX0 U16853 ( .INP(n16167), .ZN(n16166) );
  NOR2X0 U16854 ( .IN1(WX2144), .IN2(DFF_375_n1), .QN(n16167) );
  NAND2X0 U16855 ( .IN1(DFF_375_n1), .IN2(WX2144), .QN(n16165) );
  NOR2X0 U16856 ( .IN1(n10308), .IN2(n16168), .QN(WX2603) );
  NAND2X0 U16857 ( .IN1(n16169), .IN2(n16170), .QN(n16168) );
  INVX0 U16858 ( .INP(n16171), .ZN(n16170) );
  NOR2X0 U16859 ( .IN1(WX2146), .IN2(DFF_374_n1), .QN(n16171) );
  NAND2X0 U16860 ( .IN1(DFF_374_n1), .IN2(WX2146), .QN(n16169) );
  NOR2X0 U16861 ( .IN1(n10309), .IN2(n16172), .QN(WX2601) );
  NAND2X0 U16862 ( .IN1(n16173), .IN2(n16174), .QN(n16172) );
  INVX0 U16863 ( .INP(n16175), .ZN(n16174) );
  NOR2X0 U16864 ( .IN1(WX2148), .IN2(DFF_373_n1), .QN(n16175) );
  NAND2X0 U16865 ( .IN1(DFF_373_n1), .IN2(WX2148), .QN(n16173) );
  NOR2X0 U16866 ( .IN1(n10309), .IN2(n16176), .QN(WX2599) );
  NAND2X0 U16867 ( .IN1(n16177), .IN2(n16178), .QN(n16176) );
  INVX0 U16868 ( .INP(n16179), .ZN(n16178) );
  NOR2X0 U16869 ( .IN1(WX2150), .IN2(DFF_372_n1), .QN(n16179) );
  NAND2X0 U16870 ( .IN1(DFF_372_n1), .IN2(WX2150), .QN(n16177) );
  NOR2X0 U16871 ( .IN1(n10308), .IN2(n16180), .QN(WX2597) );
  NAND2X0 U16872 ( .IN1(n16181), .IN2(n16182), .QN(n16180) );
  INVX0 U16873 ( .INP(n16183), .ZN(n16182) );
  NOR2X0 U16874 ( .IN1(WX2152), .IN2(DFF_371_n1), .QN(n16183) );
  NAND2X0 U16875 ( .IN1(DFF_371_n1), .IN2(WX2152), .QN(n16181) );
  NOR2X0 U16876 ( .IN1(n10309), .IN2(n16184), .QN(WX2595) );
  NAND2X0 U16877 ( .IN1(n16185), .IN2(n16186), .QN(n16184) );
  INVX0 U16878 ( .INP(n16187), .ZN(n16186) );
  NOR2X0 U16879 ( .IN1(WX2154), .IN2(DFF_370_n1), .QN(n16187) );
  NAND2X0 U16880 ( .IN1(DFF_370_n1), .IN2(WX2154), .QN(n16185) );
  NOR2X0 U16881 ( .IN1(n10308), .IN2(n16188), .QN(WX2593) );
  NAND2X0 U16882 ( .IN1(n16189), .IN2(n16190), .QN(n16188) );
  NAND2X0 U16883 ( .IN1(n9723), .IN2(CRC_OUT_8_17), .QN(n16190) );
  NAND2X0 U16884 ( .IN1(DFF_369_n1), .IN2(WX2156), .QN(n16189) );
  NOR2X0 U16885 ( .IN1(n10308), .IN2(n16191), .QN(WX2591) );
  NAND2X0 U16886 ( .IN1(n16192), .IN2(n16193), .QN(n16191) );
  INVX0 U16887 ( .INP(n16194), .ZN(n16193) );
  NOR2X0 U16888 ( .IN1(WX2158), .IN2(DFF_368_n1), .QN(n16194) );
  NAND2X0 U16889 ( .IN1(DFF_368_n1), .IN2(WX2158), .QN(n16192) );
  NOR2X0 U16890 ( .IN1(n10310), .IN2(n16195), .QN(WX2589) );
  NOR2X0 U16891 ( .IN1(n16196), .IN2(n16197), .QN(n16195) );
  INVX0 U16892 ( .INP(n16198), .ZN(n16197) );
  NAND2X0 U16893 ( .IN1(CRC_OUT_8_15), .IN2(n16199), .QN(n16198) );
  NOR2X0 U16894 ( .IN1(n16199), .IN2(CRC_OUT_8_15), .QN(n16196) );
  NAND2X0 U16895 ( .IN1(n16200), .IN2(n16201), .QN(n16199) );
  NAND2X0 U16896 ( .IN1(n9514), .IN2(CRC_OUT_8_31), .QN(n16201) );
  NAND2X0 U16897 ( .IN1(DFF_383_n1), .IN2(WX2160), .QN(n16200) );
  NOR2X0 U16898 ( .IN1(n10308), .IN2(n16202), .QN(WX2587) );
  NAND2X0 U16899 ( .IN1(n16203), .IN2(n16204), .QN(n16202) );
  INVX0 U16900 ( .INP(n16205), .ZN(n16204) );
  NOR2X0 U16901 ( .IN1(WX2162), .IN2(DFF_366_n1), .QN(n16205) );
  NAND2X0 U16902 ( .IN1(DFF_366_n1), .IN2(WX2162), .QN(n16203) );
  NOR2X0 U16903 ( .IN1(n10308), .IN2(n16206), .QN(WX2585) );
  NAND2X0 U16904 ( .IN1(n16207), .IN2(n16208), .QN(n16206) );
  INVX0 U16905 ( .INP(n16209), .ZN(n16208) );
  NOR2X0 U16906 ( .IN1(WX2164), .IN2(DFF_365_n1), .QN(n16209) );
  NAND2X0 U16907 ( .IN1(DFF_365_n1), .IN2(WX2164), .QN(n16207) );
  NOR2X0 U16908 ( .IN1(n10309), .IN2(n16210), .QN(WX2583) );
  NAND2X0 U16909 ( .IN1(n16211), .IN2(n16212), .QN(n16210) );
  INVX0 U16910 ( .INP(n16213), .ZN(n16212) );
  NOR2X0 U16911 ( .IN1(WX2166), .IN2(DFF_364_n1), .QN(n16213) );
  NAND2X0 U16912 ( .IN1(DFF_364_n1), .IN2(WX2166), .QN(n16211) );
  NOR2X0 U16913 ( .IN1(n10309), .IN2(n16214), .QN(WX2581) );
  NAND2X0 U16914 ( .IN1(n16215), .IN2(n16216), .QN(n16214) );
  INVX0 U16915 ( .INP(n16217), .ZN(n16216) );
  NOR2X0 U16916 ( .IN1(WX2168), .IN2(DFF_363_n1), .QN(n16217) );
  NAND2X0 U16917 ( .IN1(DFF_363_n1), .IN2(WX2168), .QN(n16215) );
  NOR2X0 U16918 ( .IN1(n10309), .IN2(n16218), .QN(WX2579) );
  NOR2X0 U16919 ( .IN1(n16219), .IN2(n16220), .QN(n16218) );
  INVX0 U16920 ( .INP(n16221), .ZN(n16220) );
  NAND2X0 U16921 ( .IN1(CRC_OUT_8_10), .IN2(n16222), .QN(n16221) );
  NOR2X0 U16922 ( .IN1(n16222), .IN2(CRC_OUT_8_10), .QN(n16219) );
  NAND2X0 U16923 ( .IN1(n16223), .IN2(n16224), .QN(n16222) );
  NAND2X0 U16924 ( .IN1(n9515), .IN2(CRC_OUT_8_31), .QN(n16224) );
  NAND2X0 U16925 ( .IN1(DFF_383_n1), .IN2(WX2170), .QN(n16223) );
  NOR2X0 U16926 ( .IN1(n10310), .IN2(n16225), .QN(WX2577) );
  NOR2X0 U16927 ( .IN1(n16226), .IN2(n16227), .QN(n16225) );
  INVX0 U16928 ( .INP(n16228), .ZN(n16227) );
  NAND2X0 U16929 ( .IN1(n9836), .IN2(DFF_361_n1), .QN(n16228) );
  NOR2X0 U16930 ( .IN1(DFF_361_n1), .IN2(n9836), .QN(n16226) );
  NOR2X0 U16931 ( .IN1(n10310), .IN2(n16229), .QN(WX2575) );
  NAND2X0 U16932 ( .IN1(n16230), .IN2(n16231), .QN(n16229) );
  INVX0 U16933 ( .INP(n16232), .ZN(n16231) );
  NOR2X0 U16934 ( .IN1(WX2174), .IN2(DFF_360_n1), .QN(n16232) );
  NAND2X0 U16935 ( .IN1(DFF_360_n1), .IN2(WX2174), .QN(n16230) );
  NOR2X0 U16936 ( .IN1(n10309), .IN2(n16233), .QN(WX2573) );
  NOR2X0 U16937 ( .IN1(n16234), .IN2(n16235), .QN(n16233) );
  NOR2X0 U16938 ( .IN1(test_so20), .IN2(WX2176), .QN(n16235) );
  NOR2X0 U16939 ( .IN1(n9730), .IN2(n9861), .QN(n16234) );
  NOR2X0 U16940 ( .IN1(n10310), .IN2(n16236), .QN(WX2571) );
  NAND2X0 U16941 ( .IN1(n16237), .IN2(n16238), .QN(n16236) );
  INVX0 U16942 ( .INP(n16239), .ZN(n16238) );
  NOR2X0 U16943 ( .IN1(WX2178), .IN2(DFF_358_n1), .QN(n16239) );
  NAND2X0 U16944 ( .IN1(DFF_358_n1), .IN2(WX2178), .QN(n16237) );
  NOR2X0 U16945 ( .IN1(n10309), .IN2(n16240), .QN(WX2569) );
  NAND2X0 U16946 ( .IN1(n16241), .IN2(n16242), .QN(n16240) );
  INVX0 U16947 ( .INP(n16243), .ZN(n16242) );
  NOR2X0 U16948 ( .IN1(WX2180), .IN2(DFF_357_n1), .QN(n16243) );
  NAND2X0 U16949 ( .IN1(DFF_357_n1), .IN2(WX2180), .QN(n16241) );
  NOR2X0 U16950 ( .IN1(n10309), .IN2(n16244), .QN(WX2567) );
  NAND2X0 U16951 ( .IN1(n16245), .IN2(n16246), .QN(n16244) );
  INVX0 U16952 ( .INP(n16247), .ZN(n16246) );
  NOR2X0 U16953 ( .IN1(WX2182), .IN2(DFF_356_n1), .QN(n16247) );
  NAND2X0 U16954 ( .IN1(DFF_356_n1), .IN2(WX2182), .QN(n16245) );
  NOR2X0 U16955 ( .IN1(n10310), .IN2(n16248), .QN(WX2565) );
  NOR2X0 U16956 ( .IN1(n16249), .IN2(n16250), .QN(n16248) );
  INVX0 U16957 ( .INP(n16251), .ZN(n16250) );
  NAND2X0 U16958 ( .IN1(CRC_OUT_8_3), .IN2(n16252), .QN(n16251) );
  NOR2X0 U16959 ( .IN1(n16252), .IN2(CRC_OUT_8_3), .QN(n16249) );
  NAND2X0 U16960 ( .IN1(n16253), .IN2(n16254), .QN(n16252) );
  NAND2X0 U16961 ( .IN1(n9516), .IN2(CRC_OUT_8_31), .QN(n16254) );
  NAND2X0 U16962 ( .IN1(DFF_383_n1), .IN2(WX2184), .QN(n16253) );
  NOR2X0 U16963 ( .IN1(n10309), .IN2(n16255), .QN(WX2563) );
  NAND2X0 U16964 ( .IN1(n16256), .IN2(n16257), .QN(n16255) );
  INVX0 U16965 ( .INP(n16258), .ZN(n16257) );
  NOR2X0 U16966 ( .IN1(WX2186), .IN2(DFF_354_n1), .QN(n16258) );
  NAND2X0 U16967 ( .IN1(DFF_354_n1), .IN2(WX2186), .QN(n16256) );
  NOR2X0 U16968 ( .IN1(n10310), .IN2(n16259), .QN(WX2561) );
  NAND2X0 U16969 ( .IN1(n16260), .IN2(n16261), .QN(n16259) );
  INVX0 U16970 ( .INP(n16262), .ZN(n16261) );
  NOR2X0 U16971 ( .IN1(WX2188), .IN2(DFF_353_n1), .QN(n16262) );
  NAND2X0 U16972 ( .IN1(DFF_353_n1), .IN2(WX2188), .QN(n16260) );
  NOR2X0 U16973 ( .IN1(n10310), .IN2(n16263), .QN(WX2559) );
  NAND2X0 U16974 ( .IN1(n16264), .IN2(n16265), .QN(n16263) );
  INVX0 U16975 ( .INP(n16266), .ZN(n16265) );
  NOR2X0 U16976 ( .IN1(WX2190), .IN2(DFF_352_n1), .QN(n16266) );
  NAND2X0 U16977 ( .IN1(DFF_352_n1), .IN2(WX2190), .QN(n16264) );
  NOR2X0 U16978 ( .IN1(n10309), .IN2(n16267), .QN(WX2557) );
  NAND2X0 U16979 ( .IN1(n16268), .IN2(n16269), .QN(n16267) );
  NAND2X0 U16980 ( .IN1(n9524), .IN2(CRC_OUT_8_31), .QN(n16269) );
  NAND2X0 U16981 ( .IN1(DFF_383_n1), .IN2(WX2192), .QN(n16268) );
  NOR2X0 U16982 ( .IN1(n18366), .IN2(n10241), .QN(WX2031) );
  NOR2X0 U16983 ( .IN1(n18365), .IN2(n10241), .QN(WX2029) );
  NOR2X0 U16984 ( .IN1(n18364), .IN2(n10241), .QN(WX2027) );
  NOR2X0 U16985 ( .IN1(n18363), .IN2(n10241), .QN(WX2025) );
  NOR2X0 U16986 ( .IN1(n18362), .IN2(n10241), .QN(WX2023) );
  NOR2X0 U16987 ( .IN1(n18361), .IN2(n10241), .QN(WX2021) );
  NOR2X0 U16988 ( .IN1(n10310), .IN2(n9845), .QN(WX2019) );
  NOR2X0 U16989 ( .IN1(n18360), .IN2(n10241), .QN(WX2017) );
  NOR2X0 U16990 ( .IN1(n18359), .IN2(n10241), .QN(WX2015) );
  NOR2X0 U16991 ( .IN1(n18358), .IN2(n10240), .QN(WX2013) );
  NOR2X0 U16992 ( .IN1(n18357), .IN2(n10240), .QN(WX2011) );
  NOR2X0 U16993 ( .IN1(n18356), .IN2(n10240), .QN(WX2009) );
  NOR2X0 U16994 ( .IN1(n18355), .IN2(n10240), .QN(WX2007) );
  NOR2X0 U16995 ( .IN1(n18354), .IN2(n10240), .QN(WX2005) );
  NOR2X0 U16996 ( .IN1(n18353), .IN2(n10240), .QN(WX2003) );
  NOR2X0 U16997 ( .IN1(n18352), .IN2(n10240), .QN(WX2001) );
  NAND2X0 U16998 ( .IN1(n16270), .IN2(n16271), .QN(WX1999) );
  NOR2X0 U16999 ( .IN1(n16272), .IN2(n16273), .QN(n16271) );
  NOR2X0 U17000 ( .IN1(n15450), .IN2(n9917), .QN(n16273) );
  INVX0 U17001 ( .INP(n16274), .ZN(n15450) );
  NAND2X0 U17002 ( .IN1(n16275), .IN2(n16276), .QN(n16274) );
  NAND2X0 U17003 ( .IN1(n16277), .IN2(n16278), .QN(n16276) );
  NAND2X0 U17004 ( .IN1(n16279), .IN2(n16280), .QN(n16278) );
  NAND2X0 U17005 ( .IN1(n9427), .IN2(WX3293), .QN(n16280) );
  NAND2X0 U17006 ( .IN1(n9426), .IN2(WX3421), .QN(n16279) );
  NOR2X0 U17007 ( .IN1(n16281), .IN2(n16282), .QN(n16277) );
  NOR2X0 U17008 ( .IN1(n9523), .IN2(WX3357), .QN(n16282) );
  NOR2X0 U17009 ( .IN1(n3723), .IN2(WX3485), .QN(n16281) );
  NAND2X0 U17010 ( .IN1(n16283), .IN2(n16284), .QN(n16275) );
  NAND2X0 U17011 ( .IN1(n16285), .IN2(n16286), .QN(n16284) );
  NAND2X0 U17012 ( .IN1(n9523), .IN2(WX3357), .QN(n16286) );
  NAND2X0 U17013 ( .IN1(n3723), .IN2(WX3485), .QN(n16285) );
  NOR2X0 U17014 ( .IN1(n16287), .IN2(n16288), .QN(n16283) );
  NOR2X0 U17015 ( .IN1(n9427), .IN2(WX3293), .QN(n16288) );
  NOR2X0 U17016 ( .IN1(n9426), .IN2(WX3421), .QN(n16287) );
  INVX0 U17017 ( .INP(n16289), .ZN(n16272) );
  NAND2X0 U17018 ( .IN1(n9951), .IN2(n11151), .QN(n16289) );
  NOR2X0 U17019 ( .IN1(n16290), .IN2(n16291), .QN(n11151) );
  INVX0 U17020 ( .INP(n16292), .ZN(n16291) );
  NAND2X0 U17021 ( .IN1(n16293), .IN2(n16294), .QN(n16292) );
  NOR2X0 U17022 ( .IN1(n16294), .IN2(n16293), .QN(n16290) );
  INVX0 U17023 ( .INP(n16295), .ZN(n16293) );
  NOR2X0 U17024 ( .IN1(n16296), .IN2(n16297), .QN(n16295) );
  INVX0 U17025 ( .INP(n16298), .ZN(n16297) );
  NAND2X0 U17026 ( .IN1(test_so16), .IN2(WX2192), .QN(n16298) );
  NOR2X0 U17027 ( .IN1(WX2192), .IN2(test_so16), .QN(n16296) );
  NOR2X0 U17028 ( .IN1(n16299), .IN2(n16300), .QN(n16294) );
  INVX0 U17029 ( .INP(n16301), .ZN(n16300) );
  NAND2X0 U17030 ( .IN1(n9458), .IN2(WX2000), .QN(n16301) );
  NOR2X0 U17031 ( .IN1(WX2000), .IN2(n9458), .QN(n16299) );
  NOR2X0 U17032 ( .IN1(n16302), .IN2(n16303), .QN(n16270) );
  NOR2X0 U17033 ( .IN1(DFF_352_n1), .IN2(n9969), .QN(n16303) );
  NOR2X0 U17034 ( .IN1(n9983), .IN2(n10770), .QN(n16302) );
  NAND2X0 U17035 ( .IN1(n10200), .IN2(n8670), .QN(n10770) );
  NAND2X0 U17036 ( .IN1(n16304), .IN2(n16305), .QN(WX1997) );
  NOR2X0 U17037 ( .IN1(n16306), .IN2(n16307), .QN(n16305) );
  NOR2X0 U17038 ( .IN1(n15468), .IN2(n9916), .QN(n16307) );
  INVX0 U17039 ( .INP(n16308), .ZN(n15468) );
  NAND2X0 U17040 ( .IN1(n16309), .IN2(n16310), .QN(n16308) );
  NAND2X0 U17041 ( .IN1(n16311), .IN2(n16312), .QN(n16310) );
  NAND2X0 U17042 ( .IN1(n16313), .IN2(n16314), .QN(n16312) );
  NAND2X0 U17043 ( .IN1(n9429), .IN2(WX3291), .QN(n16314) );
  NAND2X0 U17044 ( .IN1(n9428), .IN2(WX3419), .QN(n16313) );
  NOR2X0 U17045 ( .IN1(n16315), .IN2(n16316), .QN(n16311) );
  NOR2X0 U17046 ( .IN1(n9710), .IN2(WX3355), .QN(n16316) );
  NOR2X0 U17047 ( .IN1(n3725), .IN2(WX3483), .QN(n16315) );
  NAND2X0 U17048 ( .IN1(n16317), .IN2(n16318), .QN(n16309) );
  NAND2X0 U17049 ( .IN1(n16319), .IN2(n16320), .QN(n16318) );
  NAND2X0 U17050 ( .IN1(n9710), .IN2(WX3355), .QN(n16320) );
  NAND2X0 U17051 ( .IN1(n3725), .IN2(WX3483), .QN(n16319) );
  NOR2X0 U17052 ( .IN1(n16321), .IN2(n16322), .QN(n16317) );
  NOR2X0 U17053 ( .IN1(n9429), .IN2(WX3291), .QN(n16322) );
  NOR2X0 U17054 ( .IN1(n9428), .IN2(WX3419), .QN(n16321) );
  NOR2X0 U17055 ( .IN1(n11162), .IN2(n9937), .QN(n16306) );
  NOR2X0 U17056 ( .IN1(n16323), .IN2(n16324), .QN(n11162) );
  INVX0 U17057 ( .INP(n16325), .ZN(n16324) );
  NAND2X0 U17058 ( .IN1(n16326), .IN2(n16327), .QN(n16325) );
  NOR2X0 U17059 ( .IN1(n16327), .IN2(n16326), .QN(n16323) );
  INVX0 U17060 ( .INP(n16328), .ZN(n16326) );
  NOR2X0 U17061 ( .IN1(n16329), .IN2(n16330), .QN(n16328) );
  NOR2X0 U17062 ( .IN1(WX2190), .IN2(n9460), .QN(n16330) );
  INVX0 U17063 ( .INP(n16331), .ZN(n16329) );
  NAND2X0 U17064 ( .IN1(n9460), .IN2(WX2190), .QN(n16331) );
  NOR2X0 U17065 ( .IN1(n16332), .IN2(n16333), .QN(n16327) );
  INVX0 U17066 ( .INP(n16334), .ZN(n16333) );
  NAND2X0 U17067 ( .IN1(n9459), .IN2(WX2062), .QN(n16334) );
  NOR2X0 U17068 ( .IN1(WX2062), .IN2(n9459), .QN(n16332) );
  NOR2X0 U17069 ( .IN1(n16335), .IN2(n16336), .QN(n16304) );
  NOR2X0 U17070 ( .IN1(DFF_353_n1), .IN2(n9969), .QN(n16336) );
  NOR2X0 U17071 ( .IN1(n9983), .IN2(n10771), .QN(n16335) );
  NAND2X0 U17072 ( .IN1(n10200), .IN2(n8671), .QN(n10771) );
  NAND2X0 U17073 ( .IN1(n16337), .IN2(n16338), .QN(WX1995) );
  NOR2X0 U17074 ( .IN1(n16339), .IN2(n16340), .QN(n16338) );
  NOR2X0 U17075 ( .IN1(n15490), .IN2(n9916), .QN(n16340) );
  INVX0 U17076 ( .INP(n16341), .ZN(n15490) );
  NAND2X0 U17077 ( .IN1(n16342), .IN2(n16343), .QN(n16341) );
  NAND2X0 U17078 ( .IN1(n16344), .IN2(n16345), .QN(n16343) );
  NAND2X0 U17079 ( .IN1(n16346), .IN2(n16347), .QN(n16345) );
  NAND2X0 U17080 ( .IN1(n9431), .IN2(WX3289), .QN(n16347) );
  NAND2X0 U17081 ( .IN1(n9430), .IN2(WX3417), .QN(n16346) );
  NOR2X0 U17082 ( .IN1(n16348), .IN2(n16349), .QN(n16344) );
  NOR2X0 U17083 ( .IN1(n9709), .IN2(WX3353), .QN(n16349) );
  NOR2X0 U17084 ( .IN1(n3727), .IN2(WX3481), .QN(n16348) );
  NAND2X0 U17085 ( .IN1(n16350), .IN2(n16351), .QN(n16342) );
  NAND2X0 U17086 ( .IN1(n16352), .IN2(n16353), .QN(n16351) );
  NAND2X0 U17087 ( .IN1(n9709), .IN2(WX3353), .QN(n16353) );
  NAND2X0 U17088 ( .IN1(n3727), .IN2(WX3481), .QN(n16352) );
  NOR2X0 U17089 ( .IN1(n16354), .IN2(n16355), .QN(n16350) );
  NOR2X0 U17090 ( .IN1(n9431), .IN2(WX3289), .QN(n16355) );
  NOR2X0 U17091 ( .IN1(n9430), .IN2(WX3417), .QN(n16354) );
  NOR2X0 U17092 ( .IN1(n11203), .IN2(n9937), .QN(n16339) );
  NOR2X0 U17093 ( .IN1(n16356), .IN2(n16357), .QN(n11203) );
  INVX0 U17094 ( .INP(n16358), .ZN(n16357) );
  NAND2X0 U17095 ( .IN1(n16359), .IN2(n16360), .QN(n16358) );
  NOR2X0 U17096 ( .IN1(n16360), .IN2(n16359), .QN(n16356) );
  INVX0 U17097 ( .INP(n16361), .ZN(n16359) );
  NOR2X0 U17098 ( .IN1(n16362), .IN2(n16363), .QN(n16361) );
  NOR2X0 U17099 ( .IN1(WX2188), .IN2(n9462), .QN(n16363) );
  INVX0 U17100 ( .INP(n16364), .ZN(n16362) );
  NAND2X0 U17101 ( .IN1(n9462), .IN2(WX2188), .QN(n16364) );
  NOR2X0 U17102 ( .IN1(n16365), .IN2(n16366), .QN(n16360) );
  INVX0 U17103 ( .INP(n16367), .ZN(n16366) );
  NAND2X0 U17104 ( .IN1(n9461), .IN2(WX2060), .QN(n16367) );
  NOR2X0 U17105 ( .IN1(WX2060), .IN2(n9461), .QN(n16365) );
  NOR2X0 U17106 ( .IN1(n16368), .IN2(n16369), .QN(n16337) );
  NOR2X0 U17107 ( .IN1(DFF_354_n1), .IN2(n9969), .QN(n16369) );
  NOR2X0 U17108 ( .IN1(n9983), .IN2(n10772), .QN(n16368) );
  NAND2X0 U17109 ( .IN1(n10200), .IN2(n8672), .QN(n10772) );
  NAND2X0 U17110 ( .IN1(n16370), .IN2(n16371), .QN(WX1993) );
  NOR2X0 U17111 ( .IN1(n16372), .IN2(n16373), .QN(n16371) );
  NOR2X0 U17112 ( .IN1(n15512), .IN2(n9916), .QN(n16373) );
  INVX0 U17113 ( .INP(n16374), .ZN(n15512) );
  NAND2X0 U17114 ( .IN1(n16375), .IN2(n16376), .QN(n16374) );
  NAND2X0 U17115 ( .IN1(n16377), .IN2(n16378), .QN(n16376) );
  NAND2X0 U17116 ( .IN1(n16379), .IN2(n16380), .QN(n16378) );
  NAND2X0 U17117 ( .IN1(n9433), .IN2(WX3287), .QN(n16380) );
  NAND2X0 U17118 ( .IN1(n9432), .IN2(WX3415), .QN(n16379) );
  NOR2X0 U17119 ( .IN1(n16381), .IN2(n16382), .QN(n16377) );
  NOR2X0 U17120 ( .IN1(n9708), .IN2(WX3351), .QN(n16382) );
  NOR2X0 U17121 ( .IN1(n3729), .IN2(WX3479), .QN(n16381) );
  NAND2X0 U17122 ( .IN1(n16383), .IN2(n16384), .QN(n16375) );
  NAND2X0 U17123 ( .IN1(n16385), .IN2(n16386), .QN(n16384) );
  NAND2X0 U17124 ( .IN1(n9708), .IN2(WX3351), .QN(n16386) );
  NAND2X0 U17125 ( .IN1(n3729), .IN2(WX3479), .QN(n16385) );
  NOR2X0 U17126 ( .IN1(n16387), .IN2(n16388), .QN(n16383) );
  NOR2X0 U17127 ( .IN1(n9433), .IN2(WX3287), .QN(n16388) );
  NOR2X0 U17128 ( .IN1(n9432), .IN2(WX3415), .QN(n16387) );
  NOR2X0 U17129 ( .IN1(n11213), .IN2(n9936), .QN(n16372) );
  NOR2X0 U17130 ( .IN1(n16389), .IN2(n16390), .QN(n11213) );
  INVX0 U17131 ( .INP(n16391), .ZN(n16390) );
  NAND2X0 U17132 ( .IN1(n16392), .IN2(n16393), .QN(n16391) );
  NOR2X0 U17133 ( .IN1(n16393), .IN2(n16392), .QN(n16389) );
  INVX0 U17134 ( .INP(n16394), .ZN(n16392) );
  NOR2X0 U17135 ( .IN1(n16395), .IN2(n16396), .QN(n16394) );
  NOR2X0 U17136 ( .IN1(WX2186), .IN2(n9464), .QN(n16396) );
  INVX0 U17137 ( .INP(n16397), .ZN(n16395) );
  NAND2X0 U17138 ( .IN1(n9464), .IN2(WX2186), .QN(n16397) );
  NOR2X0 U17139 ( .IN1(n16398), .IN2(n16399), .QN(n16393) );
  INVX0 U17140 ( .INP(n16400), .ZN(n16399) );
  NAND2X0 U17141 ( .IN1(n9463), .IN2(WX2058), .QN(n16400) );
  NOR2X0 U17142 ( .IN1(WX2058), .IN2(n9463), .QN(n16398) );
  NOR2X0 U17143 ( .IN1(n16401), .IN2(n16402), .QN(n16370) );
  NOR2X0 U17144 ( .IN1(DFF_355_n1), .IN2(n9969), .QN(n16402) );
  NOR2X0 U17145 ( .IN1(n9983), .IN2(n10773), .QN(n16401) );
  NAND2X0 U17146 ( .IN1(n10200), .IN2(n8673), .QN(n10773) );
  NAND2X0 U17147 ( .IN1(n16403), .IN2(n16404), .QN(WX1991) );
  NOR2X0 U17148 ( .IN1(n16405), .IN2(n16406), .QN(n16404) );
  NOR2X0 U17149 ( .IN1(n15534), .IN2(n9916), .QN(n16406) );
  INVX0 U17150 ( .INP(n16407), .ZN(n15534) );
  NAND2X0 U17151 ( .IN1(n16408), .IN2(n16409), .QN(n16407) );
  NAND2X0 U17152 ( .IN1(n16410), .IN2(n16411), .QN(n16409) );
  NAND2X0 U17153 ( .IN1(n16412), .IN2(n16413), .QN(n16411) );
  NAND2X0 U17154 ( .IN1(n9435), .IN2(WX3285), .QN(n16413) );
  NAND2X0 U17155 ( .IN1(n9434), .IN2(WX3413), .QN(n16412) );
  NOR2X0 U17156 ( .IN1(n16414), .IN2(n16415), .QN(n16410) );
  NOR2X0 U17157 ( .IN1(n9513), .IN2(WX3349), .QN(n16415) );
  NOR2X0 U17158 ( .IN1(n3731), .IN2(WX3477), .QN(n16414) );
  NAND2X0 U17159 ( .IN1(n16416), .IN2(n16417), .QN(n16408) );
  NAND2X0 U17160 ( .IN1(n16418), .IN2(n16419), .QN(n16417) );
  NAND2X0 U17161 ( .IN1(n9513), .IN2(WX3349), .QN(n16419) );
  NAND2X0 U17162 ( .IN1(n3731), .IN2(WX3477), .QN(n16418) );
  NOR2X0 U17163 ( .IN1(n16420), .IN2(n16421), .QN(n16416) );
  NOR2X0 U17164 ( .IN1(n9435), .IN2(WX3285), .QN(n16421) );
  NOR2X0 U17165 ( .IN1(n9434), .IN2(WX3413), .QN(n16420) );
  INVX0 U17166 ( .INP(n16422), .ZN(n16405) );
  NAND2X0 U17167 ( .IN1(n9951), .IN2(n11222), .QN(n16422) );
  NOR2X0 U17168 ( .IN1(n16423), .IN2(n16424), .QN(n11222) );
  INVX0 U17169 ( .INP(n16425), .ZN(n16424) );
  NAND2X0 U17170 ( .IN1(n16426), .IN2(n16427), .QN(n16425) );
  NOR2X0 U17171 ( .IN1(n16427), .IN2(n16426), .QN(n16423) );
  INVX0 U17172 ( .INP(n16428), .ZN(n16426) );
  NOR2X0 U17173 ( .IN1(n16429), .IN2(n16430), .QN(n16428) );
  INVX0 U17174 ( .INP(n16431), .ZN(n16430) );
  NAND2X0 U17175 ( .IN1(test_so14), .IN2(WX2184), .QN(n16431) );
  NOR2X0 U17176 ( .IN1(WX2184), .IN2(test_so14), .QN(n16429) );
  NOR2X0 U17177 ( .IN1(n16432), .IN2(n16433), .QN(n16427) );
  INVX0 U17178 ( .INP(n16434), .ZN(n16433) );
  NAND2X0 U17179 ( .IN1(n9465), .IN2(WX2056), .QN(n16434) );
  NOR2X0 U17180 ( .IN1(WX2056), .IN2(n9465), .QN(n16432) );
  NOR2X0 U17181 ( .IN1(n16435), .IN2(n16436), .QN(n16403) );
  NOR2X0 U17182 ( .IN1(DFF_356_n1), .IN2(n9969), .QN(n16436) );
  NOR2X0 U17183 ( .IN1(n9983), .IN2(n10774), .QN(n16435) );
  NAND2X0 U17184 ( .IN1(n10200), .IN2(n8674), .QN(n10774) );
  NAND2X0 U17185 ( .IN1(n16437), .IN2(n16438), .QN(WX1989) );
  NOR2X0 U17186 ( .IN1(n16439), .IN2(n16440), .QN(n16438) );
  NOR2X0 U17187 ( .IN1(n15556), .IN2(n9916), .QN(n16440) );
  INVX0 U17188 ( .INP(n16441), .ZN(n15556) );
  NAND2X0 U17189 ( .IN1(n16442), .IN2(n16443), .QN(n16441) );
  NAND2X0 U17190 ( .IN1(n16444), .IN2(n16445), .QN(n16443) );
  NAND2X0 U17191 ( .IN1(n16446), .IN2(n16447), .QN(n16445) );
  NAND2X0 U17192 ( .IN1(n9437), .IN2(WX3283), .QN(n16447) );
  NAND2X0 U17193 ( .IN1(n9436), .IN2(WX3411), .QN(n16446) );
  NOR2X0 U17194 ( .IN1(n16448), .IN2(n16449), .QN(n16444) );
  NOR2X0 U17195 ( .IN1(n9707), .IN2(WX3347), .QN(n16449) );
  NOR2X0 U17196 ( .IN1(n3733), .IN2(WX3475), .QN(n16448) );
  NAND2X0 U17197 ( .IN1(n16450), .IN2(n16451), .QN(n16442) );
  NAND2X0 U17198 ( .IN1(n16452), .IN2(n16453), .QN(n16451) );
  NAND2X0 U17199 ( .IN1(n9707), .IN2(WX3347), .QN(n16453) );
  NAND2X0 U17200 ( .IN1(n3733), .IN2(WX3475), .QN(n16452) );
  NOR2X0 U17201 ( .IN1(n16454), .IN2(n16455), .QN(n16450) );
  NOR2X0 U17202 ( .IN1(n9437), .IN2(WX3283), .QN(n16455) );
  NOR2X0 U17203 ( .IN1(n9436), .IN2(WX3411), .QN(n16454) );
  NOR2X0 U17204 ( .IN1(n11232), .IN2(n9936), .QN(n16439) );
  NOR2X0 U17205 ( .IN1(n16456), .IN2(n16457), .QN(n11232) );
  INVX0 U17206 ( .INP(n16458), .ZN(n16457) );
  NAND2X0 U17207 ( .IN1(n16459), .IN2(n16460), .QN(n16458) );
  NOR2X0 U17208 ( .IN1(n16460), .IN2(n16459), .QN(n16456) );
  INVX0 U17209 ( .INP(n16461), .ZN(n16459) );
  NOR2X0 U17210 ( .IN1(n16462), .IN2(n16463), .QN(n16461) );
  NOR2X0 U17211 ( .IN1(WX2182), .IN2(n9467), .QN(n16463) );
  INVX0 U17212 ( .INP(n16464), .ZN(n16462) );
  NAND2X0 U17213 ( .IN1(n9467), .IN2(WX2182), .QN(n16464) );
  NOR2X0 U17214 ( .IN1(n16465), .IN2(n16466), .QN(n16460) );
  INVX0 U17215 ( .INP(n16467), .ZN(n16466) );
  NAND2X0 U17216 ( .IN1(n9466), .IN2(WX2054), .QN(n16467) );
  NOR2X0 U17217 ( .IN1(WX2054), .IN2(n9466), .QN(n16465) );
  NOR2X0 U17218 ( .IN1(n16468), .IN2(n16469), .QN(n16437) );
  NOR2X0 U17219 ( .IN1(DFF_357_n1), .IN2(n9968), .QN(n16469) );
  NOR2X0 U17220 ( .IN1(n9983), .IN2(n10775), .QN(n16468) );
  NAND2X0 U17221 ( .IN1(n10200), .IN2(n8675), .QN(n10775) );
  NAND2X0 U17222 ( .IN1(n16470), .IN2(n16471), .QN(WX1987) );
  NOR2X0 U17223 ( .IN1(n16472), .IN2(n16473), .QN(n16471) );
  NOR2X0 U17224 ( .IN1(n9923), .IN2(n15578), .QN(n16473) );
  NAND2X0 U17225 ( .IN1(n16474), .IN2(n16475), .QN(n15578) );
  INVX0 U17226 ( .INP(n16476), .ZN(n16475) );
  NOR2X0 U17227 ( .IN1(n16477), .IN2(n16478), .QN(n16476) );
  NAND2X0 U17228 ( .IN1(n16478), .IN2(n16477), .QN(n16474) );
  NOR2X0 U17229 ( .IN1(n16479), .IN2(n16480), .QN(n16477) );
  NOR2X0 U17230 ( .IN1(n9835), .IN2(n9439), .QN(n16480) );
  INVX0 U17231 ( .INP(n16481), .ZN(n16479) );
  NAND2X0 U17232 ( .IN1(n9439), .IN2(n9835), .QN(n16481) );
  NAND2X0 U17233 ( .IN1(n16482), .IN2(n16483), .QN(n16478) );
  NAND2X0 U17234 ( .IN1(n9438), .IN2(WX3345), .QN(n16483) );
  INVX0 U17235 ( .INP(n16484), .ZN(n16482) );
  NOR2X0 U17236 ( .IN1(WX3345), .IN2(n9438), .QN(n16484) );
  NOR2X0 U17237 ( .IN1(n11243), .IN2(n9936), .QN(n16472) );
  NOR2X0 U17238 ( .IN1(n16485), .IN2(n16486), .QN(n11243) );
  INVX0 U17239 ( .INP(n16487), .ZN(n16486) );
  NAND2X0 U17240 ( .IN1(n16488), .IN2(n16489), .QN(n16487) );
  NOR2X0 U17241 ( .IN1(n16489), .IN2(n16488), .QN(n16485) );
  INVX0 U17242 ( .INP(n16490), .ZN(n16488) );
  NOR2X0 U17243 ( .IN1(n16491), .IN2(n16492), .QN(n16490) );
  NOR2X0 U17244 ( .IN1(WX2180), .IN2(n9469), .QN(n16492) );
  INVX0 U17245 ( .INP(n16493), .ZN(n16491) );
  NAND2X0 U17246 ( .IN1(n9469), .IN2(WX2180), .QN(n16493) );
  NOR2X0 U17247 ( .IN1(n16494), .IN2(n16495), .QN(n16489) );
  INVX0 U17248 ( .INP(n16496), .ZN(n16495) );
  NAND2X0 U17249 ( .IN1(n9468), .IN2(WX2052), .QN(n16496) );
  NOR2X0 U17250 ( .IN1(WX2052), .IN2(n9468), .QN(n16494) );
  NOR2X0 U17251 ( .IN1(n16497), .IN2(n16498), .QN(n16470) );
  NOR2X0 U17252 ( .IN1(DFF_358_n1), .IN2(n9968), .QN(n16498) );
  NOR2X0 U17253 ( .IN1(n9983), .IN2(n10776), .QN(n16497) );
  NAND2X0 U17254 ( .IN1(n10199), .IN2(n8676), .QN(n10776) );
  NAND2X0 U17255 ( .IN1(n16499), .IN2(n16500), .QN(WX1985) );
  NOR2X0 U17256 ( .IN1(n16501), .IN2(n16502), .QN(n16500) );
  NOR2X0 U17257 ( .IN1(n15600), .IN2(n9916), .QN(n16502) );
  INVX0 U17258 ( .INP(n16503), .ZN(n15600) );
  NAND2X0 U17259 ( .IN1(n16504), .IN2(n16505), .QN(n16503) );
  NAND2X0 U17260 ( .IN1(n16506), .IN2(n16507), .QN(n16505) );
  NAND2X0 U17261 ( .IN1(n16508), .IN2(n16509), .QN(n16507) );
  NAND2X0 U17262 ( .IN1(n9441), .IN2(WX3279), .QN(n16509) );
  NAND2X0 U17263 ( .IN1(n9440), .IN2(WX3407), .QN(n16508) );
  NOR2X0 U17264 ( .IN1(n16510), .IN2(n16511), .QN(n16506) );
  NOR2X0 U17265 ( .IN1(n9706), .IN2(WX3343), .QN(n16511) );
  NOR2X0 U17266 ( .IN1(n3737), .IN2(WX3471), .QN(n16510) );
  NAND2X0 U17267 ( .IN1(n16512), .IN2(n16513), .QN(n16504) );
  NAND2X0 U17268 ( .IN1(n16514), .IN2(n16515), .QN(n16513) );
  NAND2X0 U17269 ( .IN1(n9706), .IN2(WX3343), .QN(n16515) );
  NAND2X0 U17270 ( .IN1(n3737), .IN2(WX3471), .QN(n16514) );
  NOR2X0 U17271 ( .IN1(n16516), .IN2(n16517), .QN(n16512) );
  NOR2X0 U17272 ( .IN1(n9441), .IN2(WX3279), .QN(n16517) );
  NOR2X0 U17273 ( .IN1(n9440), .IN2(WX3407), .QN(n16516) );
  NOR2X0 U17274 ( .IN1(n11253), .IN2(n9936), .QN(n16501) );
  NOR2X0 U17275 ( .IN1(n16518), .IN2(n16519), .QN(n11253) );
  INVX0 U17276 ( .INP(n16520), .ZN(n16519) );
  NAND2X0 U17277 ( .IN1(n16521), .IN2(n16522), .QN(n16520) );
  NOR2X0 U17278 ( .IN1(n16522), .IN2(n16521), .QN(n16518) );
  INVX0 U17279 ( .INP(n16523), .ZN(n16521) );
  NOR2X0 U17280 ( .IN1(n16524), .IN2(n16525), .QN(n16523) );
  NOR2X0 U17281 ( .IN1(WX2178), .IN2(n9471), .QN(n16525) );
  INVX0 U17282 ( .INP(n16526), .ZN(n16524) );
  NAND2X0 U17283 ( .IN1(n9471), .IN2(WX2178), .QN(n16526) );
  NOR2X0 U17284 ( .IN1(n16527), .IN2(n16528), .QN(n16522) );
  INVX0 U17285 ( .INP(n16529), .ZN(n16528) );
  NAND2X0 U17286 ( .IN1(n9470), .IN2(WX2050), .QN(n16529) );
  NOR2X0 U17287 ( .IN1(WX2050), .IN2(n9470), .QN(n16527) );
  NOR2X0 U17288 ( .IN1(n16530), .IN2(n16531), .QN(n16499) );
  NOR2X0 U17289 ( .IN1(n9976), .IN2(n9861), .QN(n16531) );
  NOR2X0 U17290 ( .IN1(n9982), .IN2(n10777), .QN(n16530) );
  NAND2X0 U17291 ( .IN1(n10199), .IN2(n8677), .QN(n10777) );
  NAND2X0 U17292 ( .IN1(n16532), .IN2(n16533), .QN(WX1983) );
  NOR2X0 U17293 ( .IN1(n16534), .IN2(n16535), .QN(n16533) );
  NOR2X0 U17294 ( .IN1(n9924), .IN2(n15622), .QN(n16535) );
  NAND2X0 U17295 ( .IN1(n16536), .IN2(n16537), .QN(n15622) );
  INVX0 U17296 ( .INP(n16538), .ZN(n16537) );
  NOR2X0 U17297 ( .IN1(n16539), .IN2(n16540), .QN(n16538) );
  NAND2X0 U17298 ( .IN1(n16540), .IN2(n16539), .QN(n16536) );
  NOR2X0 U17299 ( .IN1(n16541), .IN2(n16542), .QN(n16539) );
  INVX0 U17300 ( .INP(n16543), .ZN(n16542) );
  NAND2X0 U17301 ( .IN1(test_so28), .IN2(WX3469), .QN(n16543) );
  NOR2X0 U17302 ( .IN1(WX3469), .IN2(test_so28), .QN(n16541) );
  NAND2X0 U17303 ( .IN1(n16544), .IN2(n16545), .QN(n16540) );
  NAND2X0 U17304 ( .IN1(n9442), .IN2(WX3341), .QN(n16545) );
  INVX0 U17305 ( .INP(n16546), .ZN(n16544) );
  NOR2X0 U17306 ( .IN1(WX3341), .IN2(n9442), .QN(n16546) );
  NOR2X0 U17307 ( .IN1(n11263), .IN2(n9936), .QN(n16534) );
  NOR2X0 U17308 ( .IN1(n16547), .IN2(n16548), .QN(n11263) );
  INVX0 U17309 ( .INP(n16549), .ZN(n16548) );
  NAND2X0 U17310 ( .IN1(n16550), .IN2(n16551), .QN(n16549) );
  NOR2X0 U17311 ( .IN1(n16551), .IN2(n16550), .QN(n16547) );
  INVX0 U17312 ( .INP(n16552), .ZN(n16550) );
  NOR2X0 U17313 ( .IN1(n16553), .IN2(n16554), .QN(n16552) );
  NOR2X0 U17314 ( .IN1(WX2176), .IN2(n9473), .QN(n16554) );
  INVX0 U17315 ( .INP(n16555), .ZN(n16553) );
  NAND2X0 U17316 ( .IN1(n9473), .IN2(WX2176), .QN(n16555) );
  NOR2X0 U17317 ( .IN1(n16556), .IN2(n16557), .QN(n16551) );
  INVX0 U17318 ( .INP(n16558), .ZN(n16557) );
  NAND2X0 U17319 ( .IN1(n9472), .IN2(WX2048), .QN(n16558) );
  NOR2X0 U17320 ( .IN1(WX2048), .IN2(n9472), .QN(n16556) );
  NOR2X0 U17321 ( .IN1(n16559), .IN2(n16560), .QN(n16532) );
  NOR2X0 U17322 ( .IN1(DFF_360_n1), .IN2(n9968), .QN(n16560) );
  NOR2X0 U17323 ( .IN1(n9982), .IN2(n10778), .QN(n16559) );
  NAND2X0 U17324 ( .IN1(test_so12), .IN2(n10215), .QN(n10778) );
  NAND2X0 U17325 ( .IN1(n16561), .IN2(n16562), .QN(WX1981) );
  NOR2X0 U17326 ( .IN1(n16563), .IN2(n16564), .QN(n16562) );
  NOR2X0 U17327 ( .IN1(n15644), .IN2(n9916), .QN(n16564) );
  INVX0 U17328 ( .INP(n16565), .ZN(n15644) );
  NAND2X0 U17329 ( .IN1(n16566), .IN2(n16567), .QN(n16565) );
  NAND2X0 U17330 ( .IN1(n16568), .IN2(n16569), .QN(n16567) );
  NAND2X0 U17331 ( .IN1(n16570), .IN2(n16571), .QN(n16569) );
  NAND2X0 U17332 ( .IN1(n9444), .IN2(WX3275), .QN(n16571) );
  NAND2X0 U17333 ( .IN1(n9443), .IN2(WX3403), .QN(n16570) );
  NOR2X0 U17334 ( .IN1(n16572), .IN2(n16573), .QN(n16568) );
  NOR2X0 U17335 ( .IN1(n9704), .IN2(WX3339), .QN(n16573) );
  NOR2X0 U17336 ( .IN1(n3741), .IN2(WX3467), .QN(n16572) );
  NAND2X0 U17337 ( .IN1(n16574), .IN2(n16575), .QN(n16566) );
  NAND2X0 U17338 ( .IN1(n16576), .IN2(n16577), .QN(n16575) );
  NAND2X0 U17339 ( .IN1(n9704), .IN2(WX3339), .QN(n16577) );
  NAND2X0 U17340 ( .IN1(n3741), .IN2(WX3467), .QN(n16576) );
  NOR2X0 U17341 ( .IN1(n16578), .IN2(n16579), .QN(n16574) );
  NOR2X0 U17342 ( .IN1(n9444), .IN2(WX3275), .QN(n16579) );
  NOR2X0 U17343 ( .IN1(n9443), .IN2(WX3403), .QN(n16578) );
  NOR2X0 U17344 ( .IN1(n11273), .IN2(n9936), .QN(n16563) );
  NOR2X0 U17345 ( .IN1(n16580), .IN2(n16581), .QN(n11273) );
  INVX0 U17346 ( .INP(n16582), .ZN(n16581) );
  NAND2X0 U17347 ( .IN1(n16583), .IN2(n16584), .QN(n16582) );
  NOR2X0 U17348 ( .IN1(n16584), .IN2(n16583), .QN(n16580) );
  INVX0 U17349 ( .INP(n16585), .ZN(n16583) );
  NOR2X0 U17350 ( .IN1(n16586), .IN2(n16587), .QN(n16585) );
  NOR2X0 U17351 ( .IN1(WX2174), .IN2(n9475), .QN(n16587) );
  INVX0 U17352 ( .INP(n16588), .ZN(n16586) );
  NAND2X0 U17353 ( .IN1(n9475), .IN2(WX2174), .QN(n16588) );
  NOR2X0 U17354 ( .IN1(n16589), .IN2(n16590), .QN(n16584) );
  INVX0 U17355 ( .INP(n16591), .ZN(n16590) );
  NAND2X0 U17356 ( .IN1(n9474), .IN2(WX2046), .QN(n16591) );
  NOR2X0 U17357 ( .IN1(WX2046), .IN2(n9474), .QN(n16589) );
  NOR2X0 U17358 ( .IN1(n16592), .IN2(n16593), .QN(n16561) );
  NOR2X0 U17359 ( .IN1(DFF_361_n1), .IN2(n9968), .QN(n16593) );
  NOR2X0 U17360 ( .IN1(n9982), .IN2(n10779), .QN(n16592) );
  NAND2X0 U17361 ( .IN1(n10199), .IN2(n8680), .QN(n10779) );
  NAND2X0 U17362 ( .IN1(n16594), .IN2(n16595), .QN(WX1979) );
  NOR2X0 U17363 ( .IN1(n16596), .IN2(n16597), .QN(n16595) );
  NOR2X0 U17364 ( .IN1(n15666), .IN2(n9916), .QN(n16597) );
  INVX0 U17365 ( .INP(n16598), .ZN(n15666) );
  NAND2X0 U17366 ( .IN1(n16599), .IN2(n16600), .QN(n16598) );
  NAND2X0 U17367 ( .IN1(n16601), .IN2(n16602), .QN(n16600) );
  NAND2X0 U17368 ( .IN1(n16603), .IN2(n16604), .QN(n16602) );
  NAND2X0 U17369 ( .IN1(n9446), .IN2(WX3273), .QN(n16604) );
  NAND2X0 U17370 ( .IN1(n9445), .IN2(WX3401), .QN(n16603) );
  NOR2X0 U17371 ( .IN1(n16605), .IN2(n16606), .QN(n16601) );
  NOR2X0 U17372 ( .IN1(n9703), .IN2(WX3337), .QN(n16606) );
  NOR2X0 U17373 ( .IN1(n3743), .IN2(WX3465), .QN(n16605) );
  NAND2X0 U17374 ( .IN1(n16607), .IN2(n16608), .QN(n16599) );
  NAND2X0 U17375 ( .IN1(n16609), .IN2(n16610), .QN(n16608) );
  NAND2X0 U17376 ( .IN1(n9703), .IN2(WX3337), .QN(n16610) );
  NAND2X0 U17377 ( .IN1(n3743), .IN2(WX3465), .QN(n16609) );
  NOR2X0 U17378 ( .IN1(n16611), .IN2(n16612), .QN(n16607) );
  NOR2X0 U17379 ( .IN1(n9446), .IN2(WX3273), .QN(n16612) );
  NOR2X0 U17380 ( .IN1(n9445), .IN2(WX3401), .QN(n16611) );
  INVX0 U17381 ( .INP(n16613), .ZN(n16596) );
  NAND2X0 U17382 ( .IN1(n9951), .IN2(n11314), .QN(n16613) );
  NOR2X0 U17383 ( .IN1(n16614), .IN2(n16615), .QN(n11314) );
  INVX0 U17384 ( .INP(n16616), .ZN(n16615) );
  NAND2X0 U17385 ( .IN1(n16617), .IN2(n16618), .QN(n16616) );
  NOR2X0 U17386 ( .IN1(n16618), .IN2(n16617), .QN(n16614) );
  INVX0 U17387 ( .INP(n16619), .ZN(n16617) );
  NOR2X0 U17388 ( .IN1(n16620), .IN2(n16621), .QN(n16619) );
  NOR2X0 U17389 ( .IN1(n9836), .IN2(n9477), .QN(n16621) );
  INVX0 U17390 ( .INP(n16622), .ZN(n16620) );
  NAND2X0 U17391 ( .IN1(n9477), .IN2(n9836), .QN(n16622) );
  NOR2X0 U17392 ( .IN1(n16623), .IN2(n16624), .QN(n16618) );
  INVX0 U17393 ( .INP(n16625), .ZN(n16624) );
  NAND2X0 U17394 ( .IN1(n9476), .IN2(WX2044), .QN(n16625) );
  NOR2X0 U17395 ( .IN1(WX2044), .IN2(n9476), .QN(n16623) );
  NOR2X0 U17396 ( .IN1(n16626), .IN2(n16627), .QN(n16594) );
  NOR2X0 U17397 ( .IN1(DFF_362_n1), .IN2(n9968), .QN(n16627) );
  NOR2X0 U17398 ( .IN1(n9982), .IN2(n10780), .QN(n16626) );
  NAND2X0 U17399 ( .IN1(n10199), .IN2(n8681), .QN(n10780) );
  NAND2X0 U17400 ( .IN1(n16628), .IN2(n16629), .QN(WX1977) );
  NOR2X0 U17401 ( .IN1(n16630), .IN2(n16631), .QN(n16629) );
  NOR2X0 U17402 ( .IN1(n15688), .IN2(n9916), .QN(n16631) );
  INVX0 U17403 ( .INP(n16632), .ZN(n15688) );
  NAND2X0 U17404 ( .IN1(n16633), .IN2(n16634), .QN(n16632) );
  NAND2X0 U17405 ( .IN1(n16635), .IN2(n16636), .QN(n16634) );
  NAND2X0 U17406 ( .IN1(n16637), .IN2(n16638), .QN(n16636) );
  NAND2X0 U17407 ( .IN1(n9448), .IN2(WX3271), .QN(n16638) );
  NAND2X0 U17408 ( .IN1(n9447), .IN2(WX3399), .QN(n16637) );
  NOR2X0 U17409 ( .IN1(n16639), .IN2(n16640), .QN(n16635) );
  NOR2X0 U17410 ( .IN1(n9512), .IN2(WX3335), .QN(n16640) );
  NOR2X0 U17411 ( .IN1(n3745), .IN2(WX3463), .QN(n16639) );
  NAND2X0 U17412 ( .IN1(n16641), .IN2(n16642), .QN(n16633) );
  NAND2X0 U17413 ( .IN1(n16643), .IN2(n16644), .QN(n16642) );
  NAND2X0 U17414 ( .IN1(n9512), .IN2(WX3335), .QN(n16644) );
  NAND2X0 U17415 ( .IN1(n3745), .IN2(WX3463), .QN(n16643) );
  NOR2X0 U17416 ( .IN1(n16645), .IN2(n16646), .QN(n16641) );
  NOR2X0 U17417 ( .IN1(n9448), .IN2(WX3271), .QN(n16646) );
  NOR2X0 U17418 ( .IN1(n9447), .IN2(WX3399), .QN(n16645) );
  NOR2X0 U17419 ( .IN1(n11324), .IN2(n9936), .QN(n16630) );
  NOR2X0 U17420 ( .IN1(n16647), .IN2(n16648), .QN(n11324) );
  INVX0 U17421 ( .INP(n16649), .ZN(n16648) );
  NAND2X0 U17422 ( .IN1(n16650), .IN2(n16651), .QN(n16649) );
  NOR2X0 U17423 ( .IN1(n16651), .IN2(n16650), .QN(n16647) );
  INVX0 U17424 ( .INP(n16652), .ZN(n16650) );
  NOR2X0 U17425 ( .IN1(n16653), .IN2(n16654), .QN(n16652) );
  NOR2X0 U17426 ( .IN1(WX2170), .IN2(n9479), .QN(n16654) );
  INVX0 U17427 ( .INP(n16655), .ZN(n16653) );
  NAND2X0 U17428 ( .IN1(n9479), .IN2(WX2170), .QN(n16655) );
  NOR2X0 U17429 ( .IN1(n16656), .IN2(n16657), .QN(n16651) );
  INVX0 U17430 ( .INP(n16658), .ZN(n16657) );
  NAND2X0 U17431 ( .IN1(n9478), .IN2(WX2042), .QN(n16658) );
  NOR2X0 U17432 ( .IN1(WX2042), .IN2(n9478), .QN(n16656) );
  NOR2X0 U17433 ( .IN1(n16659), .IN2(n16660), .QN(n16628) );
  NOR2X0 U17434 ( .IN1(DFF_363_n1), .IN2(n9968), .QN(n16660) );
  NOR2X0 U17435 ( .IN1(n9982), .IN2(n10781), .QN(n16659) );
  NAND2X0 U17436 ( .IN1(n10199), .IN2(n8682), .QN(n10781) );
  NAND2X0 U17437 ( .IN1(n16661), .IN2(n16662), .QN(WX1975) );
  NOR2X0 U17438 ( .IN1(n16663), .IN2(n16664), .QN(n16662) );
  NOR2X0 U17439 ( .IN1(n9923), .IN2(n15706), .QN(n16664) );
  NAND2X0 U17440 ( .IN1(n16665), .IN2(n16666), .QN(n15706) );
  INVX0 U17441 ( .INP(n16667), .ZN(n16666) );
  NOR2X0 U17442 ( .IN1(n16668), .IN2(n16669), .QN(n16667) );
  NAND2X0 U17443 ( .IN1(n16669), .IN2(n16668), .QN(n16665) );
  NOR2X0 U17444 ( .IN1(n16670), .IN2(n16671), .QN(n16668) );
  INVX0 U17445 ( .INP(n16672), .ZN(n16671) );
  NAND2X0 U17446 ( .IN1(test_so26), .IN2(WX3461), .QN(n16672) );
  NOR2X0 U17447 ( .IN1(WX3461), .IN2(test_so26), .QN(n16670) );
  NAND2X0 U17448 ( .IN1(n16673), .IN2(n16674), .QN(n16669) );
  NAND2X0 U17449 ( .IN1(n9450), .IN2(WX3269), .QN(n16674) );
  INVX0 U17450 ( .INP(n16675), .ZN(n16673) );
  NOR2X0 U17451 ( .IN1(WX3269), .IN2(n9450), .QN(n16675) );
  NOR2X0 U17452 ( .IN1(n10526), .IN2(n9936), .QN(n16663) );
  NOR2X0 U17453 ( .IN1(n16676), .IN2(n16677), .QN(n10526) );
  INVX0 U17454 ( .INP(n16678), .ZN(n16677) );
  NAND2X0 U17455 ( .IN1(n16679), .IN2(n16680), .QN(n16678) );
  NOR2X0 U17456 ( .IN1(n16680), .IN2(n16679), .QN(n16676) );
  INVX0 U17457 ( .INP(n16681), .ZN(n16679) );
  NOR2X0 U17458 ( .IN1(n16682), .IN2(n16683), .QN(n16681) );
  NOR2X0 U17459 ( .IN1(WX2168), .IN2(n9481), .QN(n16683) );
  INVX0 U17460 ( .INP(n16684), .ZN(n16682) );
  NAND2X0 U17461 ( .IN1(n9481), .IN2(WX2168), .QN(n16684) );
  NOR2X0 U17462 ( .IN1(n16685), .IN2(n16686), .QN(n16680) );
  INVX0 U17463 ( .INP(n16687), .ZN(n16686) );
  NAND2X0 U17464 ( .IN1(n9480), .IN2(WX2040), .QN(n16687) );
  NOR2X0 U17465 ( .IN1(WX2040), .IN2(n9480), .QN(n16685) );
  NOR2X0 U17466 ( .IN1(n16688), .IN2(n16689), .QN(n16661) );
  NOR2X0 U17467 ( .IN1(DFF_364_n1), .IN2(n9968), .QN(n16689) );
  NOR2X0 U17468 ( .IN1(n9982), .IN2(n10782), .QN(n16688) );
  NAND2X0 U17469 ( .IN1(n10199), .IN2(n8683), .QN(n10782) );
  NAND2X0 U17470 ( .IN1(n16690), .IN2(n16691), .QN(WX1973) );
  NOR2X0 U17471 ( .IN1(n16692), .IN2(n16693), .QN(n16691) );
  NOR2X0 U17472 ( .IN1(n15728), .IN2(n9916), .QN(n16693) );
  INVX0 U17473 ( .INP(n16694), .ZN(n15728) );
  NAND2X0 U17474 ( .IN1(n16695), .IN2(n16696), .QN(n16694) );
  NAND2X0 U17475 ( .IN1(n16697), .IN2(n16698), .QN(n16696) );
  NAND2X0 U17476 ( .IN1(n16699), .IN2(n16700), .QN(n16698) );
  NAND2X0 U17477 ( .IN1(n9452), .IN2(WX3267), .QN(n16700) );
  NAND2X0 U17478 ( .IN1(n9451), .IN2(WX3395), .QN(n16699) );
  NOR2X0 U17479 ( .IN1(n16701), .IN2(n16702), .QN(n16697) );
  NOR2X0 U17480 ( .IN1(n9701), .IN2(WX3331), .QN(n16702) );
  NOR2X0 U17481 ( .IN1(n3749), .IN2(WX3459), .QN(n16701) );
  NAND2X0 U17482 ( .IN1(n16703), .IN2(n16704), .QN(n16695) );
  NAND2X0 U17483 ( .IN1(n16705), .IN2(n16706), .QN(n16704) );
  NAND2X0 U17484 ( .IN1(n9701), .IN2(WX3331), .QN(n16706) );
  NAND2X0 U17485 ( .IN1(n3749), .IN2(WX3459), .QN(n16705) );
  NOR2X0 U17486 ( .IN1(n16707), .IN2(n16708), .QN(n16703) );
  NOR2X0 U17487 ( .IN1(n9452), .IN2(WX3267), .QN(n16708) );
  NOR2X0 U17488 ( .IN1(n9451), .IN2(WX3395), .QN(n16707) );
  NOR2X0 U17489 ( .IN1(n10536), .IN2(n9936), .QN(n16692) );
  NOR2X0 U17490 ( .IN1(n16709), .IN2(n16710), .QN(n10536) );
  INVX0 U17491 ( .INP(n16711), .ZN(n16710) );
  NAND2X0 U17492 ( .IN1(n16712), .IN2(n16713), .QN(n16711) );
  NOR2X0 U17493 ( .IN1(n16713), .IN2(n16712), .QN(n16709) );
  INVX0 U17494 ( .INP(n16714), .ZN(n16712) );
  NOR2X0 U17495 ( .IN1(n16715), .IN2(n16716), .QN(n16714) );
  NOR2X0 U17496 ( .IN1(WX2166), .IN2(n9483), .QN(n16716) );
  INVX0 U17497 ( .INP(n16717), .ZN(n16715) );
  NAND2X0 U17498 ( .IN1(n9483), .IN2(WX2166), .QN(n16717) );
  NOR2X0 U17499 ( .IN1(n16718), .IN2(n16719), .QN(n16713) );
  INVX0 U17500 ( .INP(n16720), .ZN(n16719) );
  NAND2X0 U17501 ( .IN1(n9482), .IN2(WX2038), .QN(n16720) );
  NOR2X0 U17502 ( .IN1(WX2038), .IN2(n9482), .QN(n16718) );
  NOR2X0 U17503 ( .IN1(n16721), .IN2(n16722), .QN(n16690) );
  NOR2X0 U17504 ( .IN1(DFF_365_n1), .IN2(n9968), .QN(n16722) );
  NOR2X0 U17505 ( .IN1(n9982), .IN2(n10783), .QN(n16721) );
  NAND2X0 U17506 ( .IN1(n10199), .IN2(n8684), .QN(n10783) );
  NAND2X0 U17507 ( .IN1(n16723), .IN2(n16724), .QN(WX1971) );
  NOR2X0 U17508 ( .IN1(n16725), .IN2(n16726), .QN(n16724) );
  NOR2X0 U17509 ( .IN1(n15746), .IN2(n9916), .QN(n16726) );
  INVX0 U17510 ( .INP(n16727), .ZN(n15746) );
  NAND2X0 U17511 ( .IN1(n16728), .IN2(n16729), .QN(n16727) );
  NAND2X0 U17512 ( .IN1(n16730), .IN2(n16731), .QN(n16729) );
  NAND2X0 U17513 ( .IN1(n16732), .IN2(n16733), .QN(n16731) );
  NAND2X0 U17514 ( .IN1(n9454), .IN2(WX3265), .QN(n16733) );
  NAND2X0 U17515 ( .IN1(n9453), .IN2(WX3393), .QN(n16732) );
  NOR2X0 U17516 ( .IN1(n16734), .IN2(n16735), .QN(n16730) );
  NOR2X0 U17517 ( .IN1(n9700), .IN2(WX3329), .QN(n16735) );
  NOR2X0 U17518 ( .IN1(n3751), .IN2(WX3457), .QN(n16734) );
  NAND2X0 U17519 ( .IN1(n16736), .IN2(n16737), .QN(n16728) );
  NAND2X0 U17520 ( .IN1(n16738), .IN2(n16739), .QN(n16737) );
  NAND2X0 U17521 ( .IN1(n9700), .IN2(WX3329), .QN(n16739) );
  NAND2X0 U17522 ( .IN1(n3751), .IN2(WX3457), .QN(n16738) );
  NOR2X0 U17523 ( .IN1(n16740), .IN2(n16741), .QN(n16736) );
  NOR2X0 U17524 ( .IN1(n9454), .IN2(WX3265), .QN(n16741) );
  NOR2X0 U17525 ( .IN1(n9453), .IN2(WX3393), .QN(n16740) );
  INVX0 U17526 ( .INP(n16742), .ZN(n16725) );
  NAND2X0 U17527 ( .IN1(n9951), .IN2(n10545), .QN(n16742) );
  NOR2X0 U17528 ( .IN1(n16743), .IN2(n16744), .QN(n10545) );
  INVX0 U17529 ( .INP(n16745), .ZN(n16744) );
  NAND2X0 U17530 ( .IN1(n16746), .IN2(n16747), .QN(n16745) );
  NOR2X0 U17531 ( .IN1(n16747), .IN2(n16746), .QN(n16743) );
  INVX0 U17532 ( .INP(n16748), .ZN(n16746) );
  NOR2X0 U17533 ( .IN1(n16749), .IN2(n16750), .QN(n16748) );
  INVX0 U17534 ( .INP(n16751), .ZN(n16750) );
  NAND2X0 U17535 ( .IN1(test_so17), .IN2(WX2164), .QN(n16751) );
  NOR2X0 U17536 ( .IN1(WX2164), .IN2(test_so17), .QN(n16749) );
  NOR2X0 U17537 ( .IN1(n16752), .IN2(n16753), .QN(n16747) );
  INVX0 U17538 ( .INP(n16754), .ZN(n16753) );
  NAND2X0 U17539 ( .IN1(n9484), .IN2(WX2036), .QN(n16754) );
  NOR2X0 U17540 ( .IN1(WX2036), .IN2(n9484), .QN(n16752) );
  NOR2X0 U17541 ( .IN1(n16755), .IN2(n16756), .QN(n16723) );
  NOR2X0 U17542 ( .IN1(DFF_366_n1), .IN2(n9968), .QN(n16756) );
  NOR2X0 U17543 ( .IN1(n9982), .IN2(n10784), .QN(n16755) );
  NAND2X0 U17544 ( .IN1(n10199), .IN2(n8685), .QN(n10784) );
  NAND2X0 U17545 ( .IN1(n16757), .IN2(n16758), .QN(WX1969) );
  NOR2X0 U17546 ( .IN1(n16759), .IN2(n16760), .QN(n16758) );
  NOR2X0 U17547 ( .IN1(n15768), .IN2(n9916), .QN(n16760) );
  INVX0 U17548 ( .INP(n16761), .ZN(n15768) );
  NAND2X0 U17549 ( .IN1(n16762), .IN2(n16763), .QN(n16761) );
  NAND2X0 U17550 ( .IN1(n16764), .IN2(n16765), .QN(n16763) );
  NAND2X0 U17551 ( .IN1(n16766), .IN2(n16767), .QN(n16765) );
  NAND2X0 U17552 ( .IN1(n9456), .IN2(WX3263), .QN(n16767) );
  NAND2X0 U17553 ( .IN1(n9455), .IN2(WX3391), .QN(n16766) );
  NOR2X0 U17554 ( .IN1(n16768), .IN2(n16769), .QN(n16764) );
  NOR2X0 U17555 ( .IN1(n9699), .IN2(WX3327), .QN(n16769) );
  NOR2X0 U17556 ( .IN1(n3753), .IN2(WX3455), .QN(n16768) );
  NAND2X0 U17557 ( .IN1(n16770), .IN2(n16771), .QN(n16762) );
  NAND2X0 U17558 ( .IN1(n16772), .IN2(n16773), .QN(n16771) );
  NAND2X0 U17559 ( .IN1(n9699), .IN2(WX3327), .QN(n16773) );
  NAND2X0 U17560 ( .IN1(n3753), .IN2(WX3455), .QN(n16772) );
  NOR2X0 U17561 ( .IN1(n16774), .IN2(n16775), .QN(n16770) );
  NOR2X0 U17562 ( .IN1(n9456), .IN2(WX3263), .QN(n16775) );
  NOR2X0 U17563 ( .IN1(n9455), .IN2(WX3391), .QN(n16774) );
  NOR2X0 U17564 ( .IN1(n10555), .IN2(n9936), .QN(n16759) );
  NOR2X0 U17565 ( .IN1(n16776), .IN2(n16777), .QN(n10555) );
  INVX0 U17566 ( .INP(n16778), .ZN(n16777) );
  NAND2X0 U17567 ( .IN1(n16779), .IN2(n16780), .QN(n16778) );
  NOR2X0 U17568 ( .IN1(n16780), .IN2(n16779), .QN(n16776) );
  INVX0 U17569 ( .INP(n16781), .ZN(n16779) );
  NOR2X0 U17570 ( .IN1(n16782), .IN2(n16783), .QN(n16781) );
  NOR2X0 U17571 ( .IN1(WX2162), .IN2(n9486), .QN(n16783) );
  INVX0 U17572 ( .INP(n16784), .ZN(n16782) );
  NAND2X0 U17573 ( .IN1(n9486), .IN2(WX2162), .QN(n16784) );
  NOR2X0 U17574 ( .IN1(n16785), .IN2(n16786), .QN(n16780) );
  INVX0 U17575 ( .INP(n16787), .ZN(n16786) );
  NAND2X0 U17576 ( .IN1(n9485), .IN2(WX2034), .QN(n16787) );
  NOR2X0 U17577 ( .IN1(WX2034), .IN2(n9485), .QN(n16785) );
  NOR2X0 U17578 ( .IN1(n16788), .IN2(n16789), .QN(n16757) );
  NOR2X0 U17579 ( .IN1(DFF_367_n1), .IN2(n9968), .QN(n16789) );
  NOR2X0 U17580 ( .IN1(n9982), .IN2(n10785), .QN(n16788) );
  NAND2X0 U17581 ( .IN1(n10199), .IN2(n8686), .QN(n10785) );
  NAND2X0 U17582 ( .IN1(n16790), .IN2(n16791), .QN(WX1967) );
  NOR2X0 U17583 ( .IN1(n16792), .IN2(n16793), .QN(n16791) );
  NOR2X0 U17584 ( .IN1(n9923), .IN2(n15786), .QN(n16793) );
  NAND2X0 U17585 ( .IN1(n16794), .IN2(n16795), .QN(n15786) );
  INVX0 U17586 ( .INP(n16796), .ZN(n16795) );
  NOR2X0 U17587 ( .IN1(n16797), .IN2(n16798), .QN(n16796) );
  NAND2X0 U17588 ( .IN1(n16798), .IN2(n16797), .QN(n16794) );
  INVX0 U17589 ( .INP(n16799), .ZN(n16797) );
  NAND2X0 U17590 ( .IN1(n16800), .IN2(n16801), .QN(n16799) );
  NAND2X0 U17591 ( .IN1(n16802), .IN2(WX3389), .QN(n16801) );
  NAND2X0 U17592 ( .IN1(n16803), .IN2(n16804), .QN(n16802) );
  NAND2X0 U17593 ( .IN1(test_so24), .IN2(WX3325), .QN(n16804) );
  NAND2X0 U17594 ( .IN1(n9188), .IN2(n9844), .QN(n16803) );
  NAND2X0 U17595 ( .IN1(n9189), .IN2(n16805), .QN(n16800) );
  NOR2X0 U17596 ( .IN1(n16806), .IN2(n16807), .QN(n16805) );
  NOR2X0 U17597 ( .IN1(test_so24), .IN2(WX3325), .QN(n16807) );
  NOR2X0 U17598 ( .IN1(n9188), .IN2(n9844), .QN(n16806) );
  NAND2X0 U17599 ( .IN1(n16808), .IN2(n16809), .QN(n16798) );
  NAND2X0 U17600 ( .IN1(n9511), .IN2(n10021), .QN(n16809) );
  NAND2X0 U17601 ( .IN1(TM1), .IN2(WX3453), .QN(n16808) );
  NOR2X0 U17602 ( .IN1(n10567), .IN2(n9936), .QN(n16792) );
  NOR2X0 U17603 ( .IN1(n16810), .IN2(n16811), .QN(n10567) );
  INVX0 U17604 ( .INP(n16812), .ZN(n16811) );
  NAND2X0 U17605 ( .IN1(n16813), .IN2(n16814), .QN(n16812) );
  NOR2X0 U17606 ( .IN1(n16814), .IN2(n16813), .QN(n16810) );
  NAND2X0 U17607 ( .IN1(n16815), .IN2(n16816), .QN(n16813) );
  NAND2X0 U17608 ( .IN1(n9217), .IN2(n16817), .QN(n16816) );
  INVX0 U17609 ( .INP(n16818), .ZN(n16815) );
  NOR2X0 U17610 ( .IN1(n16817), .IN2(n9217), .QN(n16818) );
  NOR2X0 U17611 ( .IN1(n16819), .IN2(n16820), .QN(n16817) );
  INVX0 U17612 ( .INP(n16821), .ZN(n16820) );
  NAND2X0 U17613 ( .IN1(n18366), .IN2(WX2160), .QN(n16821) );
  NOR2X0 U17614 ( .IN1(WX2160), .IN2(n18366), .QN(n16819) );
  NOR2X0 U17615 ( .IN1(n16822), .IN2(n16823), .QN(n16814) );
  INVX0 U17616 ( .INP(n16824), .ZN(n16823) );
  NAND2X0 U17617 ( .IN1(n9216), .IN2(n10021), .QN(n16824) );
  NOR2X0 U17618 ( .IN1(n10010), .IN2(n9216), .QN(n16822) );
  NOR2X0 U17619 ( .IN1(n16825), .IN2(n16826), .QN(n16790) );
  NOR2X0 U17620 ( .IN1(DFF_368_n1), .IN2(n9968), .QN(n16826) );
  NOR2X0 U17621 ( .IN1(n9982), .IN2(n10786), .QN(n16825) );
  NAND2X0 U17622 ( .IN1(n10198), .IN2(n8687), .QN(n10786) );
  NAND2X0 U17623 ( .IN1(n16827), .IN2(n16828), .QN(WX1965) );
  NOR2X0 U17624 ( .IN1(n16829), .IN2(n16830), .QN(n16828) );
  NOR2X0 U17625 ( .IN1(n15808), .IN2(n9915), .QN(n16830) );
  NOR2X0 U17626 ( .IN1(n16831), .IN2(n16832), .QN(n15808) );
  INVX0 U17627 ( .INP(n16833), .ZN(n16832) );
  NAND2X0 U17628 ( .IN1(n16834), .IN2(n16835), .QN(n16833) );
  NOR2X0 U17629 ( .IN1(n16835), .IN2(n16834), .QN(n16831) );
  NAND2X0 U17630 ( .IN1(n16836), .IN2(n16837), .QN(n16834) );
  NAND2X0 U17631 ( .IN1(n9191), .IN2(n16838), .QN(n16837) );
  INVX0 U17632 ( .INP(n16839), .ZN(n16836) );
  NOR2X0 U17633 ( .IN1(n16838), .IN2(n9191), .QN(n16839) );
  NOR2X0 U17634 ( .IN1(n16840), .IN2(n16841), .QN(n16838) );
  INVX0 U17635 ( .INP(n16842), .ZN(n16841) );
  NAND2X0 U17636 ( .IN1(n18381), .IN2(WX3451), .QN(n16842) );
  NOR2X0 U17637 ( .IN1(WX3451), .IN2(n18381), .QN(n16840) );
  NOR2X0 U17638 ( .IN1(n16843), .IN2(n16844), .QN(n16835) );
  INVX0 U17639 ( .INP(n16845), .ZN(n16844) );
  NAND2X0 U17640 ( .IN1(n9190), .IN2(n10020), .QN(n16845) );
  NOR2X0 U17641 ( .IN1(n10011), .IN2(n9190), .QN(n16843) );
  NOR2X0 U17642 ( .IN1(n10587), .IN2(n9936), .QN(n16829) );
  NOR2X0 U17643 ( .IN1(n16846), .IN2(n16847), .QN(n10587) );
  INVX0 U17644 ( .INP(n16848), .ZN(n16847) );
  NAND2X0 U17645 ( .IN1(n16849), .IN2(n16850), .QN(n16848) );
  NOR2X0 U17646 ( .IN1(n16850), .IN2(n16849), .QN(n16846) );
  NAND2X0 U17647 ( .IN1(n16851), .IN2(n16852), .QN(n16849) );
  NAND2X0 U17648 ( .IN1(n9219), .IN2(n16853), .QN(n16852) );
  INVX0 U17649 ( .INP(n16854), .ZN(n16851) );
  NOR2X0 U17650 ( .IN1(n16853), .IN2(n9219), .QN(n16854) );
  NOR2X0 U17651 ( .IN1(n16855), .IN2(n16856), .QN(n16853) );
  INVX0 U17652 ( .INP(n16857), .ZN(n16856) );
  NAND2X0 U17653 ( .IN1(n18365), .IN2(WX2158), .QN(n16857) );
  NOR2X0 U17654 ( .IN1(WX2158), .IN2(n18365), .QN(n16855) );
  NOR2X0 U17655 ( .IN1(n16858), .IN2(n16859), .QN(n16850) );
  INVX0 U17656 ( .INP(n16860), .ZN(n16859) );
  NAND2X0 U17657 ( .IN1(n9218), .IN2(n10020), .QN(n16860) );
  NOR2X0 U17658 ( .IN1(n10011), .IN2(n9218), .QN(n16858) );
  NOR2X0 U17659 ( .IN1(n16861), .IN2(n16862), .QN(n16827) );
  NOR2X0 U17660 ( .IN1(DFF_369_n1), .IN2(n9968), .QN(n16862) );
  NOR2X0 U17661 ( .IN1(n9982), .IN2(n10787), .QN(n16861) );
  NAND2X0 U17662 ( .IN1(n10198), .IN2(n8688), .QN(n10787) );
  NAND2X0 U17663 ( .IN1(n16863), .IN2(n16864), .QN(WX1963) );
  NOR2X0 U17664 ( .IN1(n16865), .IN2(n16866), .QN(n16864) );
  NOR2X0 U17665 ( .IN1(n15831), .IN2(n9915), .QN(n16866) );
  NOR2X0 U17666 ( .IN1(n16867), .IN2(n16868), .QN(n15831) );
  INVX0 U17667 ( .INP(n16869), .ZN(n16868) );
  NAND2X0 U17668 ( .IN1(n16870), .IN2(n16871), .QN(n16869) );
  NOR2X0 U17669 ( .IN1(n16871), .IN2(n16870), .QN(n16867) );
  NAND2X0 U17670 ( .IN1(n16872), .IN2(n16873), .QN(n16870) );
  NAND2X0 U17671 ( .IN1(n9193), .IN2(n16874), .QN(n16873) );
  INVX0 U17672 ( .INP(n16875), .ZN(n16872) );
  NOR2X0 U17673 ( .IN1(n16874), .IN2(n9193), .QN(n16875) );
  NOR2X0 U17674 ( .IN1(n16876), .IN2(n16877), .QN(n16874) );
  INVX0 U17675 ( .INP(n16878), .ZN(n16877) );
  NAND2X0 U17676 ( .IN1(n18380), .IN2(WX3449), .QN(n16878) );
  NOR2X0 U17677 ( .IN1(WX3449), .IN2(n18380), .QN(n16876) );
  NOR2X0 U17678 ( .IN1(n16879), .IN2(n16880), .QN(n16871) );
  INVX0 U17679 ( .INP(n16881), .ZN(n16880) );
  NAND2X0 U17680 ( .IN1(n9192), .IN2(n10020), .QN(n16881) );
  NOR2X0 U17681 ( .IN1(n10011), .IN2(n9192), .QN(n16879) );
  INVX0 U17682 ( .INP(n16882), .ZN(n16865) );
  NAND2X0 U17683 ( .IN1(n9951), .IN2(n10617), .QN(n16882) );
  NOR2X0 U17684 ( .IN1(n16883), .IN2(n16884), .QN(n10617) );
  INVX0 U17685 ( .INP(n16885), .ZN(n16884) );
  NAND2X0 U17686 ( .IN1(n16886), .IN2(n16887), .QN(n16885) );
  NOR2X0 U17687 ( .IN1(n16887), .IN2(n16886), .QN(n16883) );
  NAND2X0 U17688 ( .IN1(n16888), .IN2(n16889), .QN(n16886) );
  NAND2X0 U17689 ( .IN1(n9723), .IN2(n16890), .QN(n16889) );
  INVX0 U17690 ( .INP(n16891), .ZN(n16890) );
  NAND2X0 U17691 ( .IN1(n16891), .IN2(WX2156), .QN(n16888) );
  NAND2X0 U17692 ( .IN1(n16892), .IN2(n16893), .QN(n16891) );
  INVX0 U17693 ( .INP(n16894), .ZN(n16893) );
  NOR2X0 U17694 ( .IN1(n9870), .IN2(n18364), .QN(n16894) );
  NAND2X0 U17695 ( .IN1(n18364), .IN2(n9870), .QN(n16892) );
  NOR2X0 U17696 ( .IN1(n16895), .IN2(n16896), .QN(n16887) );
  INVX0 U17697 ( .INP(n16897), .ZN(n16896) );
  NAND2X0 U17698 ( .IN1(n9220), .IN2(n10020), .QN(n16897) );
  NOR2X0 U17699 ( .IN1(n10011), .IN2(n9220), .QN(n16895) );
  NOR2X0 U17700 ( .IN1(n16898), .IN2(n16899), .QN(n16863) );
  NOR2X0 U17701 ( .IN1(DFF_370_n1), .IN2(n9967), .QN(n16899) );
  NOR2X0 U17702 ( .IN1(n9982), .IN2(n10788), .QN(n16898) );
  NAND2X0 U17703 ( .IN1(n10198), .IN2(n8689), .QN(n10788) );
  NAND2X0 U17704 ( .IN1(n16900), .IN2(n16901), .QN(WX1961) );
  NOR2X0 U17705 ( .IN1(n16902), .IN2(n16903), .QN(n16901) );
  NOR2X0 U17706 ( .IN1(n15853), .IN2(n9915), .QN(n16903) );
  NOR2X0 U17707 ( .IN1(n16904), .IN2(n16905), .QN(n15853) );
  INVX0 U17708 ( .INP(n16906), .ZN(n16905) );
  NAND2X0 U17709 ( .IN1(n16907), .IN2(n16908), .QN(n16906) );
  NOR2X0 U17710 ( .IN1(n16908), .IN2(n16907), .QN(n16904) );
  NAND2X0 U17711 ( .IN1(n16909), .IN2(n16910), .QN(n16907) );
  NAND2X0 U17712 ( .IN1(n9195), .IN2(n16911), .QN(n16910) );
  INVX0 U17713 ( .INP(n16912), .ZN(n16909) );
  NOR2X0 U17714 ( .IN1(n16911), .IN2(n9195), .QN(n16912) );
  NOR2X0 U17715 ( .IN1(n16913), .IN2(n16914), .QN(n16911) );
  INVX0 U17716 ( .INP(n16915), .ZN(n16914) );
  NAND2X0 U17717 ( .IN1(n18379), .IN2(WX3447), .QN(n16915) );
  NOR2X0 U17718 ( .IN1(WX3447), .IN2(n18379), .QN(n16913) );
  NOR2X0 U17719 ( .IN1(n16916), .IN2(n16917), .QN(n16908) );
  INVX0 U17720 ( .INP(n16918), .ZN(n16917) );
  NAND2X0 U17721 ( .IN1(n9194), .IN2(n10020), .QN(n16918) );
  NOR2X0 U17722 ( .IN1(n10011), .IN2(n9194), .QN(n16916) );
  NOR2X0 U17723 ( .IN1(n10627), .IN2(n9935), .QN(n16902) );
  NOR2X0 U17724 ( .IN1(n16919), .IN2(n16920), .QN(n10627) );
  INVX0 U17725 ( .INP(n16921), .ZN(n16920) );
  NAND2X0 U17726 ( .IN1(n16922), .IN2(n16923), .QN(n16921) );
  NOR2X0 U17727 ( .IN1(n16923), .IN2(n16922), .QN(n16919) );
  NAND2X0 U17728 ( .IN1(n16924), .IN2(n16925), .QN(n16922) );
  NAND2X0 U17729 ( .IN1(n9222), .IN2(n16926), .QN(n16925) );
  INVX0 U17730 ( .INP(n16927), .ZN(n16924) );
  NOR2X0 U17731 ( .IN1(n16926), .IN2(n9222), .QN(n16927) );
  NOR2X0 U17732 ( .IN1(n16928), .IN2(n16929), .QN(n16926) );
  INVX0 U17733 ( .INP(n16930), .ZN(n16929) );
  NAND2X0 U17734 ( .IN1(n18363), .IN2(WX2154), .QN(n16930) );
  NOR2X0 U17735 ( .IN1(WX2154), .IN2(n18363), .QN(n16928) );
  NOR2X0 U17736 ( .IN1(n16931), .IN2(n16932), .QN(n16923) );
  INVX0 U17737 ( .INP(n16933), .ZN(n16932) );
  NAND2X0 U17738 ( .IN1(n9221), .IN2(n10020), .QN(n16933) );
  NOR2X0 U17739 ( .IN1(n10011), .IN2(n9221), .QN(n16931) );
  NOR2X0 U17740 ( .IN1(n16934), .IN2(n16935), .QN(n16900) );
  NOR2X0 U17741 ( .IN1(DFF_371_n1), .IN2(n9967), .QN(n16935) );
  NOR2X0 U17742 ( .IN1(n9981), .IN2(n10789), .QN(n16934) );
  NAND2X0 U17743 ( .IN1(n10198), .IN2(n8690), .QN(n10789) );
  NAND2X0 U17744 ( .IN1(n16936), .IN2(n16937), .QN(WX1959) );
  NOR2X0 U17745 ( .IN1(n16938), .IN2(n16939), .QN(n16937) );
  NOR2X0 U17746 ( .IN1(n15875), .IN2(n9915), .QN(n16939) );
  NOR2X0 U17747 ( .IN1(n16940), .IN2(n16941), .QN(n15875) );
  INVX0 U17748 ( .INP(n16942), .ZN(n16941) );
  NAND2X0 U17749 ( .IN1(n16943), .IN2(n16944), .QN(n16942) );
  NOR2X0 U17750 ( .IN1(n16944), .IN2(n16943), .QN(n16940) );
  NAND2X0 U17751 ( .IN1(n16945), .IN2(n16946), .QN(n16943) );
  NAND2X0 U17752 ( .IN1(n9197), .IN2(n16947), .QN(n16946) );
  INVX0 U17753 ( .INP(n16948), .ZN(n16945) );
  NOR2X0 U17754 ( .IN1(n16947), .IN2(n9197), .QN(n16948) );
  NOR2X0 U17755 ( .IN1(n16949), .IN2(n16950), .QN(n16947) );
  INVX0 U17756 ( .INP(n16951), .ZN(n16950) );
  NAND2X0 U17757 ( .IN1(n18378), .IN2(WX3445), .QN(n16951) );
  NOR2X0 U17758 ( .IN1(WX3445), .IN2(n18378), .QN(n16949) );
  NOR2X0 U17759 ( .IN1(n16952), .IN2(n16953), .QN(n16944) );
  INVX0 U17760 ( .INP(n16954), .ZN(n16953) );
  NAND2X0 U17761 ( .IN1(n9196), .IN2(n10019), .QN(n16954) );
  NOR2X0 U17762 ( .IN1(n10012), .IN2(n9196), .QN(n16952) );
  NOR2X0 U17763 ( .IN1(n10638), .IN2(n9935), .QN(n16938) );
  NOR2X0 U17764 ( .IN1(n16955), .IN2(n16956), .QN(n10638) );
  INVX0 U17765 ( .INP(n16957), .ZN(n16956) );
  NAND2X0 U17766 ( .IN1(n16958), .IN2(n16959), .QN(n16957) );
  NOR2X0 U17767 ( .IN1(n16959), .IN2(n16958), .QN(n16955) );
  NAND2X0 U17768 ( .IN1(n16960), .IN2(n16961), .QN(n16958) );
  NAND2X0 U17769 ( .IN1(n9224), .IN2(n16962), .QN(n16961) );
  INVX0 U17770 ( .INP(n16963), .ZN(n16960) );
  NOR2X0 U17771 ( .IN1(n16962), .IN2(n9224), .QN(n16963) );
  NOR2X0 U17772 ( .IN1(n16964), .IN2(n16965), .QN(n16962) );
  INVX0 U17773 ( .INP(n16966), .ZN(n16965) );
  NAND2X0 U17774 ( .IN1(n18362), .IN2(WX2152), .QN(n16966) );
  NOR2X0 U17775 ( .IN1(WX2152), .IN2(n18362), .QN(n16964) );
  NOR2X0 U17776 ( .IN1(n16967), .IN2(n16968), .QN(n16959) );
  INVX0 U17777 ( .INP(n16969), .ZN(n16968) );
  NAND2X0 U17778 ( .IN1(n9223), .IN2(n10019), .QN(n16969) );
  NOR2X0 U17779 ( .IN1(n10012), .IN2(n9223), .QN(n16967) );
  NOR2X0 U17780 ( .IN1(n16970), .IN2(n16971), .QN(n16936) );
  NOR2X0 U17781 ( .IN1(DFF_372_n1), .IN2(n9967), .QN(n16971) );
  NOR2X0 U17782 ( .IN1(n9981), .IN2(n10790), .QN(n16970) );
  NAND2X0 U17783 ( .IN1(n10198), .IN2(n8691), .QN(n10790) );
  NAND2X0 U17784 ( .IN1(n16972), .IN2(n16973), .QN(WX1957) );
  NOR2X0 U17785 ( .IN1(n16974), .IN2(n16975), .QN(n16973) );
  NOR2X0 U17786 ( .IN1(n15897), .IN2(n9915), .QN(n16975) );
  NOR2X0 U17787 ( .IN1(n16976), .IN2(n16977), .QN(n15897) );
  INVX0 U17788 ( .INP(n16978), .ZN(n16977) );
  NAND2X0 U17789 ( .IN1(n16979), .IN2(n16980), .QN(n16978) );
  NOR2X0 U17790 ( .IN1(n16980), .IN2(n16979), .QN(n16976) );
  NAND2X0 U17791 ( .IN1(n16981), .IN2(n16982), .QN(n16979) );
  NAND2X0 U17792 ( .IN1(n9199), .IN2(n16983), .QN(n16982) );
  INVX0 U17793 ( .INP(n16984), .ZN(n16981) );
  NOR2X0 U17794 ( .IN1(n16983), .IN2(n9199), .QN(n16984) );
  NOR2X0 U17795 ( .IN1(n16985), .IN2(n16986), .QN(n16983) );
  INVX0 U17796 ( .INP(n16987), .ZN(n16986) );
  NAND2X0 U17797 ( .IN1(n18377), .IN2(WX3443), .QN(n16987) );
  NOR2X0 U17798 ( .IN1(WX3443), .IN2(n18377), .QN(n16985) );
  NOR2X0 U17799 ( .IN1(n16988), .IN2(n16989), .QN(n16980) );
  INVX0 U17800 ( .INP(n16990), .ZN(n16989) );
  NAND2X0 U17801 ( .IN1(n9198), .IN2(n10019), .QN(n16990) );
  NOR2X0 U17802 ( .IN1(n10012), .IN2(n9198), .QN(n16988) );
  NOR2X0 U17803 ( .IN1(n10648), .IN2(n9935), .QN(n16974) );
  NOR2X0 U17804 ( .IN1(n16991), .IN2(n16992), .QN(n10648) );
  INVX0 U17805 ( .INP(n16993), .ZN(n16992) );
  NAND2X0 U17806 ( .IN1(n16994), .IN2(n16995), .QN(n16993) );
  NOR2X0 U17807 ( .IN1(n16995), .IN2(n16994), .QN(n16991) );
  NAND2X0 U17808 ( .IN1(n16996), .IN2(n16997), .QN(n16994) );
  NAND2X0 U17809 ( .IN1(n9226), .IN2(n16998), .QN(n16997) );
  INVX0 U17810 ( .INP(n16999), .ZN(n16996) );
  NOR2X0 U17811 ( .IN1(n16998), .IN2(n9226), .QN(n16999) );
  NOR2X0 U17812 ( .IN1(n17000), .IN2(n17001), .QN(n16998) );
  INVX0 U17813 ( .INP(n17002), .ZN(n17001) );
  NAND2X0 U17814 ( .IN1(n18361), .IN2(WX2150), .QN(n17002) );
  NOR2X0 U17815 ( .IN1(WX2150), .IN2(n18361), .QN(n17000) );
  NOR2X0 U17816 ( .IN1(n17003), .IN2(n17004), .QN(n16995) );
  INVX0 U17817 ( .INP(n17005), .ZN(n17004) );
  NAND2X0 U17818 ( .IN1(n9225), .IN2(n10019), .QN(n17005) );
  NOR2X0 U17819 ( .IN1(n10011), .IN2(n9225), .QN(n17003) );
  NOR2X0 U17820 ( .IN1(n17006), .IN2(n17007), .QN(n16972) );
  NOR2X0 U17821 ( .IN1(DFF_373_n1), .IN2(n9967), .QN(n17007) );
  NOR2X0 U17822 ( .IN1(n9981), .IN2(n10791), .QN(n17006) );
  NAND2X0 U17823 ( .IN1(n10198), .IN2(n8692), .QN(n10791) );
  NAND2X0 U17824 ( .IN1(n17008), .IN2(n17009), .QN(WX1955) );
  NOR2X0 U17825 ( .IN1(n17010), .IN2(n17011), .QN(n17009) );
  NOR2X0 U17826 ( .IN1(n15919), .IN2(n9915), .QN(n17011) );
  NOR2X0 U17827 ( .IN1(n17012), .IN2(n17013), .QN(n15919) );
  INVX0 U17828 ( .INP(n17014), .ZN(n17013) );
  NAND2X0 U17829 ( .IN1(n17015), .IN2(n17016), .QN(n17014) );
  NOR2X0 U17830 ( .IN1(n17016), .IN2(n17015), .QN(n17012) );
  NAND2X0 U17831 ( .IN1(n17017), .IN2(n17018), .QN(n17015) );
  NAND2X0 U17832 ( .IN1(n9201), .IN2(n17019), .QN(n17018) );
  INVX0 U17833 ( .INP(n17020), .ZN(n17017) );
  NOR2X0 U17834 ( .IN1(n17019), .IN2(n9201), .QN(n17020) );
  NOR2X0 U17835 ( .IN1(n17021), .IN2(n17022), .QN(n17019) );
  INVX0 U17836 ( .INP(n17023), .ZN(n17022) );
  NAND2X0 U17837 ( .IN1(n18376), .IN2(WX3441), .QN(n17023) );
  NOR2X0 U17838 ( .IN1(WX3441), .IN2(n18376), .QN(n17021) );
  NOR2X0 U17839 ( .IN1(n17024), .IN2(n17025), .QN(n17016) );
  INVX0 U17840 ( .INP(n17026), .ZN(n17025) );
  NAND2X0 U17841 ( .IN1(n9200), .IN2(n10019), .QN(n17026) );
  NOR2X0 U17842 ( .IN1(n10010), .IN2(n9200), .QN(n17024) );
  INVX0 U17843 ( .INP(n17027), .ZN(n17010) );
  NAND2X0 U17844 ( .IN1(n9951), .IN2(n10657), .QN(n17027) );
  NOR2X0 U17845 ( .IN1(n17028), .IN2(n17029), .QN(n10657) );
  INVX0 U17846 ( .INP(n17030), .ZN(n17029) );
  NAND2X0 U17847 ( .IN1(n17031), .IN2(n17032), .QN(n17030) );
  NOR2X0 U17848 ( .IN1(n17032), .IN2(n17031), .QN(n17028) );
  NAND2X0 U17849 ( .IN1(n17033), .IN2(n17034), .QN(n17031) );
  NAND2X0 U17850 ( .IN1(n17035), .IN2(WX2084), .QN(n17034) );
  NAND2X0 U17851 ( .IN1(n17036), .IN2(n17037), .QN(n17035) );
  NAND2X0 U17852 ( .IN1(test_so13), .IN2(WX2020), .QN(n17037) );
  NAND2X0 U17853 ( .IN1(n9227), .IN2(n9845), .QN(n17036) );
  NAND2X0 U17854 ( .IN1(n9228), .IN2(n17038), .QN(n17033) );
  NOR2X0 U17855 ( .IN1(n17039), .IN2(n17040), .QN(n17038) );
  NOR2X0 U17856 ( .IN1(test_so13), .IN2(WX2020), .QN(n17040) );
  NOR2X0 U17857 ( .IN1(n9227), .IN2(n9845), .QN(n17039) );
  INVX0 U17858 ( .INP(n17041), .ZN(n17032) );
  NAND2X0 U17859 ( .IN1(n17042), .IN2(n17043), .QN(n17041) );
  NAND2X0 U17860 ( .IN1(n9719), .IN2(n10018), .QN(n17043) );
  NAND2X0 U17861 ( .IN1(TM1), .IN2(WX2148), .QN(n17042) );
  NOR2X0 U17862 ( .IN1(n17044), .IN2(n17045), .QN(n17008) );
  NOR2X0 U17863 ( .IN1(DFF_374_n1), .IN2(n9967), .QN(n17045) );
  NOR2X0 U17864 ( .IN1(n9981), .IN2(n10792), .QN(n17044) );
  NAND2X0 U17865 ( .IN1(n10198), .IN2(n8693), .QN(n10792) );
  NAND2X0 U17866 ( .IN1(n17046), .IN2(n17047), .QN(WX1953) );
  NOR2X0 U17867 ( .IN1(n17048), .IN2(n17049), .QN(n17047) );
  NOR2X0 U17868 ( .IN1(n9924), .IN2(n15941), .QN(n17049) );
  NAND2X0 U17869 ( .IN1(n17050), .IN2(n17051), .QN(n15941) );
  NAND2X0 U17870 ( .IN1(n17052), .IN2(n17053), .QN(n17051) );
  INVX0 U17871 ( .INP(n17054), .ZN(n17050) );
  NOR2X0 U17872 ( .IN1(n17053), .IN2(n17052), .QN(n17054) );
  NAND2X0 U17873 ( .IN1(n17055), .IN2(n17056), .QN(n17052) );
  NAND2X0 U17874 ( .IN1(n17057), .IN2(WX3375), .QN(n17056) );
  NAND2X0 U17875 ( .IN1(n17058), .IN2(n17059), .QN(n17057) );
  NAND2X0 U17876 ( .IN1(test_so29), .IN2(WX3311), .QN(n17059) );
  NAND2X0 U17877 ( .IN1(n9202), .IN2(n9831), .QN(n17058) );
  NAND2X0 U17878 ( .IN1(n9203), .IN2(n17060), .QN(n17055) );
  NOR2X0 U17879 ( .IN1(n17061), .IN2(n17062), .QN(n17060) );
  NOR2X0 U17880 ( .IN1(test_so29), .IN2(WX3311), .QN(n17062) );
  NOR2X0 U17881 ( .IN1(n9202), .IN2(n9831), .QN(n17061) );
  NOR2X0 U17882 ( .IN1(n17063), .IN2(n17064), .QN(n17053) );
  INVX0 U17883 ( .INP(n17065), .ZN(n17064) );
  NAND2X0 U17884 ( .IN1(n18375), .IN2(n10018), .QN(n17065) );
  NOR2X0 U17885 ( .IN1(n10012), .IN2(n18375), .QN(n17063) );
  NOR2X0 U17886 ( .IN1(n10667), .IN2(n9935), .QN(n17048) );
  NOR2X0 U17887 ( .IN1(n17066), .IN2(n17067), .QN(n10667) );
  INVX0 U17888 ( .INP(n17068), .ZN(n17067) );
  NAND2X0 U17889 ( .IN1(n17069), .IN2(n17070), .QN(n17068) );
  NOR2X0 U17890 ( .IN1(n17070), .IN2(n17069), .QN(n17066) );
  NAND2X0 U17891 ( .IN1(n17071), .IN2(n17072), .QN(n17069) );
  NAND2X0 U17892 ( .IN1(n9230), .IN2(n17073), .QN(n17072) );
  INVX0 U17893 ( .INP(n17074), .ZN(n17071) );
  NOR2X0 U17894 ( .IN1(n17073), .IN2(n9230), .QN(n17074) );
  NOR2X0 U17895 ( .IN1(n17075), .IN2(n17076), .QN(n17073) );
  INVX0 U17896 ( .INP(n17077), .ZN(n17076) );
  NAND2X0 U17897 ( .IN1(n18360), .IN2(WX2146), .QN(n17077) );
  NOR2X0 U17898 ( .IN1(WX2146), .IN2(n18360), .QN(n17075) );
  NOR2X0 U17899 ( .IN1(n17078), .IN2(n17079), .QN(n17070) );
  INVX0 U17900 ( .INP(n17080), .ZN(n17079) );
  NAND2X0 U17901 ( .IN1(n9229), .IN2(n10018), .QN(n17080) );
  NOR2X0 U17902 ( .IN1(n10013), .IN2(n9229), .QN(n17078) );
  NOR2X0 U17903 ( .IN1(n17081), .IN2(n17082), .QN(n17046) );
  NOR2X0 U17904 ( .IN1(DFF_375_n1), .IN2(n9967), .QN(n17082) );
  NOR2X0 U17905 ( .IN1(n9981), .IN2(n10793), .QN(n17081) );
  NAND2X0 U17906 ( .IN1(n10198), .IN2(n8694), .QN(n10793) );
  NAND2X0 U17907 ( .IN1(n17083), .IN2(n17084), .QN(WX1951) );
  NOR2X0 U17908 ( .IN1(n17085), .IN2(n17086), .QN(n17084) );
  NOR2X0 U17909 ( .IN1(n15963), .IN2(n9915), .QN(n17086) );
  NOR2X0 U17910 ( .IN1(n17087), .IN2(n17088), .QN(n15963) );
  INVX0 U17911 ( .INP(n17089), .ZN(n17088) );
  NAND2X0 U17912 ( .IN1(n17090), .IN2(n17091), .QN(n17089) );
  NOR2X0 U17913 ( .IN1(n17091), .IN2(n17090), .QN(n17087) );
  NAND2X0 U17914 ( .IN1(n17092), .IN2(n17093), .QN(n17090) );
  NAND2X0 U17915 ( .IN1(n9205), .IN2(n17094), .QN(n17093) );
  INVX0 U17916 ( .INP(n17095), .ZN(n17092) );
  NOR2X0 U17917 ( .IN1(n17094), .IN2(n9205), .QN(n17095) );
  NOR2X0 U17918 ( .IN1(n17096), .IN2(n17097), .QN(n17094) );
  INVX0 U17919 ( .INP(n17098), .ZN(n17097) );
  NAND2X0 U17920 ( .IN1(n18374), .IN2(WX3437), .QN(n17098) );
  NOR2X0 U17921 ( .IN1(WX3437), .IN2(n18374), .QN(n17096) );
  NOR2X0 U17922 ( .IN1(n17099), .IN2(n17100), .QN(n17091) );
  INVX0 U17923 ( .INP(n17101), .ZN(n17100) );
  NAND2X0 U17924 ( .IN1(n9204), .IN2(n10018), .QN(n17101) );
  NOR2X0 U17925 ( .IN1(n10012), .IN2(n9204), .QN(n17099) );
  NOR2X0 U17926 ( .IN1(n10678), .IN2(n9935), .QN(n17085) );
  NOR2X0 U17927 ( .IN1(n17102), .IN2(n17103), .QN(n10678) );
  INVX0 U17928 ( .INP(n17104), .ZN(n17103) );
  NAND2X0 U17929 ( .IN1(n17105), .IN2(n17106), .QN(n17104) );
  NOR2X0 U17930 ( .IN1(n17106), .IN2(n17105), .QN(n17102) );
  NAND2X0 U17931 ( .IN1(n17107), .IN2(n17108), .QN(n17105) );
  NAND2X0 U17932 ( .IN1(n9232), .IN2(n17109), .QN(n17108) );
  INVX0 U17933 ( .INP(n17110), .ZN(n17107) );
  NOR2X0 U17934 ( .IN1(n17109), .IN2(n9232), .QN(n17110) );
  NOR2X0 U17935 ( .IN1(n17111), .IN2(n17112), .QN(n17109) );
  INVX0 U17936 ( .INP(n17113), .ZN(n17112) );
  NAND2X0 U17937 ( .IN1(n18359), .IN2(WX2144), .QN(n17113) );
  NOR2X0 U17938 ( .IN1(WX2144), .IN2(n18359), .QN(n17111) );
  NOR2X0 U17939 ( .IN1(n17114), .IN2(n17115), .QN(n17106) );
  INVX0 U17940 ( .INP(n17116), .ZN(n17115) );
  NAND2X0 U17941 ( .IN1(n9231), .IN2(n10018), .QN(n17116) );
  NOR2X0 U17942 ( .IN1(n10013), .IN2(n9231), .QN(n17114) );
  NOR2X0 U17943 ( .IN1(n17117), .IN2(n17118), .QN(n17083) );
  NOR2X0 U17944 ( .IN1(DFF_376_n1), .IN2(n9967), .QN(n17118) );
  NOR2X0 U17945 ( .IN1(n9981), .IN2(n10794), .QN(n17117) );
  NAND2X0 U17946 ( .IN1(n10198), .IN2(n8695), .QN(n10794) );
  NAND2X0 U17947 ( .IN1(n17119), .IN2(n17120), .QN(WX1949) );
  NOR2X0 U17948 ( .IN1(n17121), .IN2(n17122), .QN(n17120) );
  NOR2X0 U17949 ( .IN1(n15985), .IN2(n9915), .QN(n17122) );
  NOR2X0 U17950 ( .IN1(n17123), .IN2(n17124), .QN(n15985) );
  INVX0 U17951 ( .INP(n17125), .ZN(n17124) );
  NAND2X0 U17952 ( .IN1(n17126), .IN2(n17127), .QN(n17125) );
  NOR2X0 U17953 ( .IN1(n17127), .IN2(n17126), .QN(n17123) );
  NAND2X0 U17954 ( .IN1(n17128), .IN2(n17129), .QN(n17126) );
  NAND2X0 U17955 ( .IN1(n9207), .IN2(n17130), .QN(n17129) );
  INVX0 U17956 ( .INP(n17131), .ZN(n17128) );
  NOR2X0 U17957 ( .IN1(n17130), .IN2(n9207), .QN(n17131) );
  NOR2X0 U17958 ( .IN1(n17132), .IN2(n17133), .QN(n17130) );
  INVX0 U17959 ( .INP(n17134), .ZN(n17133) );
  NAND2X0 U17960 ( .IN1(n18373), .IN2(WX3435), .QN(n17134) );
  NOR2X0 U17961 ( .IN1(WX3435), .IN2(n18373), .QN(n17132) );
  NOR2X0 U17962 ( .IN1(n17135), .IN2(n17136), .QN(n17127) );
  INVX0 U17963 ( .INP(n17137), .ZN(n17136) );
  NAND2X0 U17964 ( .IN1(n9206), .IN2(n10018), .QN(n17137) );
  NOR2X0 U17965 ( .IN1(n10013), .IN2(n9206), .QN(n17135) );
  NOR2X0 U17966 ( .IN1(n10697), .IN2(n9935), .QN(n17121) );
  NOR2X0 U17967 ( .IN1(n17138), .IN2(n17139), .QN(n10697) );
  INVX0 U17968 ( .INP(n17140), .ZN(n17139) );
  NAND2X0 U17969 ( .IN1(n17141), .IN2(n17142), .QN(n17140) );
  NOR2X0 U17970 ( .IN1(n17142), .IN2(n17141), .QN(n17138) );
  NAND2X0 U17971 ( .IN1(n17143), .IN2(n17144), .QN(n17141) );
  NAND2X0 U17972 ( .IN1(n9234), .IN2(n17145), .QN(n17144) );
  INVX0 U17973 ( .INP(n17146), .ZN(n17143) );
  NOR2X0 U17974 ( .IN1(n17145), .IN2(n9234), .QN(n17146) );
  NOR2X0 U17975 ( .IN1(n17147), .IN2(n17148), .QN(n17145) );
  INVX0 U17976 ( .INP(n17149), .ZN(n17148) );
  NAND2X0 U17977 ( .IN1(n18358), .IN2(WX2142), .QN(n17149) );
  NOR2X0 U17978 ( .IN1(WX2142), .IN2(n18358), .QN(n17147) );
  NOR2X0 U17979 ( .IN1(n17150), .IN2(n17151), .QN(n17142) );
  INVX0 U17980 ( .INP(n17152), .ZN(n17151) );
  NAND2X0 U17981 ( .IN1(n9233), .IN2(n10018), .QN(n17152) );
  NOR2X0 U17982 ( .IN1(n10013), .IN2(n9233), .QN(n17150) );
  NOR2X0 U17983 ( .IN1(n17153), .IN2(n17154), .QN(n17119) );
  NOR2X0 U17984 ( .IN1(n9976), .IN2(n9862), .QN(n17154) );
  NOR2X0 U17985 ( .IN1(n9981), .IN2(n10795), .QN(n17153) );
  NAND2X0 U17986 ( .IN1(n10197), .IN2(n8696), .QN(n10795) );
  NAND2X0 U17987 ( .IN1(n17155), .IN2(n17156), .QN(WX1947) );
  NOR2X0 U17988 ( .IN1(n17157), .IN2(n17158), .QN(n17156) );
  NOR2X0 U17989 ( .IN1(n9924), .IN2(n16007), .QN(n17158) );
  NAND2X0 U17990 ( .IN1(n17159), .IN2(n17160), .QN(n16007) );
  INVX0 U17991 ( .INP(n17161), .ZN(n17160) );
  NOR2X0 U17992 ( .IN1(n17162), .IN2(n17163), .QN(n17161) );
  NAND2X0 U17993 ( .IN1(n17163), .IN2(n17162), .QN(n17159) );
  NOR2X0 U17994 ( .IN1(n17164), .IN2(n17165), .QN(n17162) );
  INVX0 U17995 ( .INP(n17166), .ZN(n17165) );
  NAND2X0 U17996 ( .IN1(n9690), .IN2(n17167), .QN(n17166) );
  NOR2X0 U17997 ( .IN1(n17167), .IN2(n9690), .QN(n17164) );
  NOR2X0 U17998 ( .IN1(n17168), .IN2(n17169), .QN(n17167) );
  INVX0 U17999 ( .INP(n17170), .ZN(n17169) );
  NAND2X0 U18000 ( .IN1(test_so27), .IN2(n8606), .QN(n17170) );
  NOR2X0 U18001 ( .IN1(n8606), .IN2(test_so27), .QN(n17168) );
  NAND2X0 U18002 ( .IN1(n17171), .IN2(n17172), .QN(n17163) );
  NAND2X0 U18003 ( .IN1(n9208), .IN2(n10017), .QN(n17172) );
  INVX0 U18004 ( .INP(n17173), .ZN(n17171) );
  NOR2X0 U18005 ( .IN1(n10011), .IN2(n9208), .QN(n17173) );
  NOR2X0 U18006 ( .IN1(n10729), .IN2(n9935), .QN(n17157) );
  NOR2X0 U18007 ( .IN1(n17174), .IN2(n17175), .QN(n10729) );
  INVX0 U18008 ( .INP(n17176), .ZN(n17175) );
  NAND2X0 U18009 ( .IN1(n17177), .IN2(n17178), .QN(n17176) );
  NOR2X0 U18010 ( .IN1(n17178), .IN2(n17177), .QN(n17174) );
  NAND2X0 U18011 ( .IN1(n17179), .IN2(n17180), .QN(n17177) );
  NAND2X0 U18012 ( .IN1(n9236), .IN2(n17181), .QN(n17180) );
  INVX0 U18013 ( .INP(n17182), .ZN(n17179) );
  NOR2X0 U18014 ( .IN1(n17181), .IN2(n9236), .QN(n17182) );
  NOR2X0 U18015 ( .IN1(n17183), .IN2(n17184), .QN(n17181) );
  INVX0 U18016 ( .INP(n17185), .ZN(n17184) );
  NAND2X0 U18017 ( .IN1(n18357), .IN2(WX2140), .QN(n17185) );
  NOR2X0 U18018 ( .IN1(WX2140), .IN2(n18357), .QN(n17183) );
  NOR2X0 U18019 ( .IN1(n17186), .IN2(n17187), .QN(n17178) );
  INVX0 U18020 ( .INP(n17188), .ZN(n17187) );
  NAND2X0 U18021 ( .IN1(n9235), .IN2(n10017), .QN(n17188) );
  NOR2X0 U18022 ( .IN1(n10012), .IN2(n9235), .QN(n17186) );
  NOR2X0 U18023 ( .IN1(n17189), .IN2(n17190), .QN(n17155) );
  NOR2X0 U18024 ( .IN1(DFF_378_n1), .IN2(n9967), .QN(n17190) );
  NOR2X0 U18025 ( .IN1(n9981), .IN2(n10796), .QN(n17189) );
  NAND2X0 U18026 ( .IN1(test_so11), .IN2(n10215), .QN(n10796) );
  NAND2X0 U18027 ( .IN1(n17191), .IN2(n17192), .QN(WX1945) );
  NOR2X0 U18028 ( .IN1(n17193), .IN2(n17194), .QN(n17192) );
  NOR2X0 U18029 ( .IN1(n16029), .IN2(n9915), .QN(n17194) );
  NOR2X0 U18030 ( .IN1(n17195), .IN2(n17196), .QN(n16029) );
  INVX0 U18031 ( .INP(n17197), .ZN(n17196) );
  NAND2X0 U18032 ( .IN1(n17198), .IN2(n17199), .QN(n17197) );
  NOR2X0 U18033 ( .IN1(n17199), .IN2(n17198), .QN(n17195) );
  NAND2X0 U18034 ( .IN1(n17200), .IN2(n17201), .QN(n17198) );
  NAND2X0 U18035 ( .IN1(n9210), .IN2(n17202), .QN(n17201) );
  INVX0 U18036 ( .INP(n17203), .ZN(n17200) );
  NOR2X0 U18037 ( .IN1(n17202), .IN2(n9210), .QN(n17203) );
  NOR2X0 U18038 ( .IN1(n17204), .IN2(n17205), .QN(n17202) );
  INVX0 U18039 ( .INP(n17206), .ZN(n17205) );
  NAND2X0 U18040 ( .IN1(n18371), .IN2(WX3431), .QN(n17206) );
  NOR2X0 U18041 ( .IN1(WX3431), .IN2(n18371), .QN(n17204) );
  NOR2X0 U18042 ( .IN1(n17207), .IN2(n17208), .QN(n17199) );
  INVX0 U18043 ( .INP(n17209), .ZN(n17208) );
  NAND2X0 U18044 ( .IN1(n9209), .IN2(n10017), .QN(n17209) );
  NOR2X0 U18045 ( .IN1(n10011), .IN2(n9209), .QN(n17207) );
  NOR2X0 U18046 ( .IN1(n10739), .IN2(n9935), .QN(n17193) );
  NOR2X0 U18047 ( .IN1(n17210), .IN2(n17211), .QN(n10739) );
  INVX0 U18048 ( .INP(n17212), .ZN(n17211) );
  NAND2X0 U18049 ( .IN1(n17213), .IN2(n17214), .QN(n17212) );
  NOR2X0 U18050 ( .IN1(n17214), .IN2(n17213), .QN(n17210) );
  NAND2X0 U18051 ( .IN1(n17215), .IN2(n17216), .QN(n17213) );
  NAND2X0 U18052 ( .IN1(n9238), .IN2(n17217), .QN(n17216) );
  INVX0 U18053 ( .INP(n17218), .ZN(n17215) );
  NOR2X0 U18054 ( .IN1(n17217), .IN2(n9238), .QN(n17218) );
  NOR2X0 U18055 ( .IN1(n17219), .IN2(n17220), .QN(n17217) );
  INVX0 U18056 ( .INP(n17221), .ZN(n17220) );
  NAND2X0 U18057 ( .IN1(n18356), .IN2(WX2138), .QN(n17221) );
  NOR2X0 U18058 ( .IN1(WX2138), .IN2(n18356), .QN(n17219) );
  NOR2X0 U18059 ( .IN1(n17222), .IN2(n17223), .QN(n17214) );
  INVX0 U18060 ( .INP(n17224), .ZN(n17223) );
  NAND2X0 U18061 ( .IN1(n9237), .IN2(n10017), .QN(n17224) );
  NOR2X0 U18062 ( .IN1(n10010), .IN2(n9237), .QN(n17222) );
  NOR2X0 U18063 ( .IN1(n17225), .IN2(n17226), .QN(n17191) );
  NOR2X0 U18064 ( .IN1(DFF_379_n1), .IN2(n9967), .QN(n17226) );
  NOR2X0 U18065 ( .IN1(n9981), .IN2(n10797), .QN(n17225) );
  NAND2X0 U18066 ( .IN1(n10197), .IN2(n8699), .QN(n10797) );
  NAND2X0 U18067 ( .IN1(n17227), .IN2(n17228), .QN(WX1943) );
  NOR2X0 U18068 ( .IN1(n17229), .IN2(n17230), .QN(n17228) );
  NOR2X0 U18069 ( .IN1(n16051), .IN2(n9915), .QN(n17230) );
  NOR2X0 U18070 ( .IN1(n17231), .IN2(n17232), .QN(n16051) );
  INVX0 U18071 ( .INP(n17233), .ZN(n17232) );
  NAND2X0 U18072 ( .IN1(n17234), .IN2(n17235), .QN(n17233) );
  NOR2X0 U18073 ( .IN1(n17235), .IN2(n17234), .QN(n17231) );
  NAND2X0 U18074 ( .IN1(n17236), .IN2(n17237), .QN(n17234) );
  NAND2X0 U18075 ( .IN1(n9212), .IN2(n17238), .QN(n17237) );
  INVX0 U18076 ( .INP(n17239), .ZN(n17236) );
  NOR2X0 U18077 ( .IN1(n17238), .IN2(n9212), .QN(n17239) );
  NOR2X0 U18078 ( .IN1(n17240), .IN2(n17241), .QN(n17238) );
  INVX0 U18079 ( .INP(n17242), .ZN(n17241) );
  NAND2X0 U18080 ( .IN1(n18370), .IN2(WX3429), .QN(n17242) );
  NOR2X0 U18081 ( .IN1(WX3429), .IN2(n18370), .QN(n17240) );
  NOR2X0 U18082 ( .IN1(n17243), .IN2(n17244), .QN(n17235) );
  INVX0 U18083 ( .INP(n17245), .ZN(n17244) );
  NAND2X0 U18084 ( .IN1(n9211), .IN2(n10017), .QN(n17245) );
  NOR2X0 U18085 ( .IN1(n10010), .IN2(n9211), .QN(n17243) );
  INVX0 U18086 ( .INP(n17246), .ZN(n17229) );
  NAND2X0 U18087 ( .IN1(n9948), .IN2(n10749), .QN(n17246) );
  NOR2X0 U18088 ( .IN1(n17247), .IN2(n17248), .QN(n10749) );
  INVX0 U18089 ( .INP(n17249), .ZN(n17248) );
  NAND2X0 U18090 ( .IN1(n17250), .IN2(n17251), .QN(n17249) );
  NOR2X0 U18091 ( .IN1(n17251), .IN2(n17250), .QN(n17247) );
  NAND2X0 U18092 ( .IN1(n17252), .IN2(n17253), .QN(n17250) );
  NAND2X0 U18093 ( .IN1(n17254), .IN2(WX2072), .QN(n17253) );
  NAND2X0 U18094 ( .IN1(n17255), .IN2(n17256), .QN(n17254) );
  NAND2X0 U18095 ( .IN1(test_so18), .IN2(WX2008), .QN(n17256) );
  NAND2X0 U18096 ( .IN1(n9239), .IN2(n9832), .QN(n17255) );
  NAND2X0 U18097 ( .IN1(n9240), .IN2(n17257), .QN(n17252) );
  NOR2X0 U18098 ( .IN1(n17258), .IN2(n17259), .QN(n17257) );
  NOR2X0 U18099 ( .IN1(test_so18), .IN2(WX2008), .QN(n17259) );
  NOR2X0 U18100 ( .IN1(n9239), .IN2(n9832), .QN(n17258) );
  NOR2X0 U18101 ( .IN1(n17260), .IN2(n17261), .QN(n17251) );
  INVX0 U18102 ( .INP(n17262), .ZN(n17261) );
  NAND2X0 U18103 ( .IN1(n18355), .IN2(n10017), .QN(n17262) );
  NOR2X0 U18104 ( .IN1(n10013), .IN2(n18355), .QN(n17260) );
  NOR2X0 U18105 ( .IN1(n17263), .IN2(n17264), .QN(n17227) );
  NOR2X0 U18106 ( .IN1(DFF_380_n1), .IN2(n9967), .QN(n17264) );
  NOR2X0 U18107 ( .IN1(n9981), .IN2(n10798), .QN(n17263) );
  NAND2X0 U18108 ( .IN1(n10197), .IN2(n8700), .QN(n10798) );
  NAND2X0 U18109 ( .IN1(n17265), .IN2(n17266), .QN(WX1941) );
  NOR2X0 U18110 ( .IN1(n17267), .IN2(n17268), .QN(n17266) );
  NOR2X0 U18111 ( .IN1(n16074), .IN2(n9915), .QN(n17268) );
  NOR2X0 U18112 ( .IN1(n17269), .IN2(n17270), .QN(n16074) );
  INVX0 U18113 ( .INP(n17271), .ZN(n17270) );
  NAND2X0 U18114 ( .IN1(n17272), .IN2(n17273), .QN(n17271) );
  NOR2X0 U18115 ( .IN1(n17273), .IN2(n17272), .QN(n17269) );
  NAND2X0 U18116 ( .IN1(n17274), .IN2(n17275), .QN(n17272) );
  NAND2X0 U18117 ( .IN1(n9214), .IN2(n17276), .QN(n17275) );
  INVX0 U18118 ( .INP(n17277), .ZN(n17274) );
  NOR2X0 U18119 ( .IN1(n17276), .IN2(n9214), .QN(n17277) );
  NOR2X0 U18120 ( .IN1(n17278), .IN2(n17279), .QN(n17276) );
  INVX0 U18121 ( .INP(n17280), .ZN(n17279) );
  NAND2X0 U18122 ( .IN1(n18369), .IN2(WX3427), .QN(n17280) );
  NOR2X0 U18123 ( .IN1(WX3427), .IN2(n18369), .QN(n17278) );
  NOR2X0 U18124 ( .IN1(n17281), .IN2(n17282), .QN(n17273) );
  INVX0 U18125 ( .INP(n17283), .ZN(n17282) );
  NAND2X0 U18126 ( .IN1(n9213), .IN2(n10014), .QN(n17283) );
  NOR2X0 U18127 ( .IN1(n10010), .IN2(n9213), .QN(n17281) );
  NOR2X0 U18128 ( .IN1(n10759), .IN2(n9935), .QN(n17267) );
  NOR2X0 U18129 ( .IN1(n17284), .IN2(n17285), .QN(n10759) );
  INVX0 U18130 ( .INP(n17286), .ZN(n17285) );
  NAND2X0 U18131 ( .IN1(n17287), .IN2(n17288), .QN(n17286) );
  NOR2X0 U18132 ( .IN1(n17288), .IN2(n17287), .QN(n17284) );
  NAND2X0 U18133 ( .IN1(n17289), .IN2(n17290), .QN(n17287) );
  NAND2X0 U18134 ( .IN1(n9242), .IN2(n17291), .QN(n17290) );
  INVX0 U18135 ( .INP(n17292), .ZN(n17289) );
  NOR2X0 U18136 ( .IN1(n17291), .IN2(n9242), .QN(n17292) );
  NOR2X0 U18137 ( .IN1(n17293), .IN2(n17294), .QN(n17291) );
  INVX0 U18138 ( .INP(n17295), .ZN(n17294) );
  NAND2X0 U18139 ( .IN1(n18354), .IN2(WX2134), .QN(n17295) );
  NOR2X0 U18140 ( .IN1(WX2134), .IN2(n18354), .QN(n17293) );
  NOR2X0 U18141 ( .IN1(n17296), .IN2(n17297), .QN(n17288) );
  INVX0 U18142 ( .INP(n17298), .ZN(n17297) );
  NAND2X0 U18143 ( .IN1(n9241), .IN2(n10013), .QN(n17298) );
  NOR2X0 U18144 ( .IN1(n10011), .IN2(n9241), .QN(n17296) );
  NOR2X0 U18145 ( .IN1(n17299), .IN2(n17300), .QN(n17265) );
  NOR2X0 U18146 ( .IN1(DFF_381_n1), .IN2(n9967), .QN(n17300) );
  NOR2X0 U18147 ( .IN1(n9981), .IN2(n10799), .QN(n17299) );
  NAND2X0 U18148 ( .IN1(n10206), .IN2(n8701), .QN(n10799) );
  NAND2X0 U18149 ( .IN1(n17301), .IN2(n17302), .QN(WX1939) );
  NOR2X0 U18150 ( .IN1(n17303), .IN2(n17304), .QN(n17302) );
  NOR2X0 U18151 ( .IN1(n9926), .IN2(n16096), .QN(n17304) );
  NAND2X0 U18152 ( .IN1(n17305), .IN2(n17306), .QN(n16096) );
  INVX0 U18153 ( .INP(n17307), .ZN(n17306) );
  NOR2X0 U18154 ( .IN1(n17308), .IN2(n17309), .QN(n17307) );
  NAND2X0 U18155 ( .IN1(n17309), .IN2(n17308), .QN(n17305) );
  NOR2X0 U18156 ( .IN1(n17310), .IN2(n17311), .QN(n17308) );
  INVX0 U18157 ( .INP(n17312), .ZN(n17311) );
  NAND2X0 U18158 ( .IN1(n9686), .IN2(n17313), .QN(n17312) );
  NOR2X0 U18159 ( .IN1(n17313), .IN2(n9686), .QN(n17310) );
  NOR2X0 U18160 ( .IN1(n17314), .IN2(n17315), .QN(n17313) );
  INVX0 U18161 ( .INP(n17316), .ZN(n17315) );
  NAND2X0 U18162 ( .IN1(test_so25), .IN2(n8610), .QN(n17316) );
  NOR2X0 U18163 ( .IN1(n8610), .IN2(test_so25), .QN(n17314) );
  NAND2X0 U18164 ( .IN1(n17317), .IN2(n17318), .QN(n17309) );
  NAND2X0 U18165 ( .IN1(n9215), .IN2(n10014), .QN(n17318) );
  INVX0 U18166 ( .INP(n17319), .ZN(n17317) );
  NOR2X0 U18167 ( .IN1(n10012), .IN2(n9215), .QN(n17319) );
  NOR2X0 U18168 ( .IN1(n10769), .IN2(n9939), .QN(n17303) );
  NOR2X0 U18169 ( .IN1(n17320), .IN2(n17321), .QN(n10769) );
  INVX0 U18170 ( .INP(n17322), .ZN(n17321) );
  NAND2X0 U18171 ( .IN1(n17323), .IN2(n17324), .QN(n17322) );
  NOR2X0 U18172 ( .IN1(n17324), .IN2(n17323), .QN(n17320) );
  NAND2X0 U18173 ( .IN1(n17325), .IN2(n17326), .QN(n17323) );
  NAND2X0 U18174 ( .IN1(n9244), .IN2(n17327), .QN(n17326) );
  INVX0 U18175 ( .INP(n17328), .ZN(n17325) );
  NOR2X0 U18176 ( .IN1(n17327), .IN2(n9244), .QN(n17328) );
  NOR2X0 U18177 ( .IN1(n17329), .IN2(n17330), .QN(n17327) );
  INVX0 U18178 ( .INP(n17331), .ZN(n17330) );
  NAND2X0 U18179 ( .IN1(n18353), .IN2(WX2132), .QN(n17331) );
  NOR2X0 U18180 ( .IN1(WX2132), .IN2(n18353), .QN(n17329) );
  NOR2X0 U18181 ( .IN1(n17332), .IN2(n17333), .QN(n17324) );
  INVX0 U18182 ( .INP(n17334), .ZN(n17333) );
  NAND2X0 U18183 ( .IN1(n9243), .IN2(n10014), .QN(n17334) );
  NOR2X0 U18184 ( .IN1(n10012), .IN2(n9243), .QN(n17332) );
  NOR2X0 U18185 ( .IN1(n17335), .IN2(n17336), .QN(n17301) );
  NOR2X0 U18186 ( .IN1(DFF_382_n1), .IN2(n9971), .QN(n17336) );
  NOR2X0 U18187 ( .IN1(n9981), .IN2(n10800), .QN(n17335) );
  NAND2X0 U18188 ( .IN1(n10191), .IN2(n8702), .QN(n10800) );
  INVX0 U18189 ( .INP(n2339), .ZN(n11345) );
  NOR2X0 U18190 ( .IN1(n10012), .IN2(n2340), .QN(n2339) );
  NAND2X0 U18191 ( .IN1(n17337), .IN2(n17338), .QN(WX1937) );
  NOR2X0 U18192 ( .IN1(n17339), .IN2(n17340), .QN(n17338) );
  NOR2X0 U18193 ( .IN1(n13782), .IN2(n9927), .QN(n17340) );
  NAND2X0 U18194 ( .IN1(n17341), .IN2(TM1), .QN(n10563) );
  NOR2X0 U18195 ( .IN1(TM0), .IN2(n10240), .QN(n17341) );
  NOR2X0 U18196 ( .IN1(n17342), .IN2(n17343), .QN(n13782) );
  INVX0 U18197 ( .INP(n17344), .ZN(n17343) );
  NAND2X0 U18198 ( .IN1(n17345), .IN2(n17346), .QN(n17344) );
  NOR2X0 U18199 ( .IN1(n17346), .IN2(n17345), .QN(n17342) );
  NAND2X0 U18200 ( .IN1(n17347), .IN2(n17348), .QN(n17345) );
  NAND2X0 U18201 ( .IN1(n9018), .IN2(n17349), .QN(n17348) );
  INVX0 U18202 ( .INP(n17350), .ZN(n17347) );
  NOR2X0 U18203 ( .IN1(n17349), .IN2(n9018), .QN(n17350) );
  NOR2X0 U18204 ( .IN1(n17351), .IN2(n17352), .QN(n17349) );
  INVX0 U18205 ( .INP(n17353), .ZN(n17352) );
  NAND2X0 U18206 ( .IN1(n18352), .IN2(WX2130), .QN(n17353) );
  NOR2X0 U18207 ( .IN1(WX2130), .IN2(n18352), .QN(n17351) );
  NOR2X0 U18208 ( .IN1(n17354), .IN2(n17355), .QN(n17346) );
  INVX0 U18209 ( .INP(n17356), .ZN(n17355) );
  NAND2X0 U18210 ( .IN1(n9017), .IN2(n10014), .QN(n17356) );
  NOR2X0 U18211 ( .IN1(n10012), .IN2(n9017), .QN(n17354) );
  NOR2X0 U18212 ( .IN1(n16118), .IN2(n9907), .QN(n17339) );
  INVX0 U18213 ( .INP(n2153), .ZN(n10525) );
  NOR2X0 U18214 ( .IN1(n17357), .IN2(n17358), .QN(n16118) );
  INVX0 U18215 ( .INP(n17359), .ZN(n17358) );
  NAND2X0 U18216 ( .IN1(n17360), .IN2(n17361), .QN(n17359) );
  NOR2X0 U18217 ( .IN1(n17361), .IN2(n17360), .QN(n17357) );
  NAND2X0 U18218 ( .IN1(n17362), .IN2(n17363), .QN(n17360) );
  NAND2X0 U18219 ( .IN1(n9016), .IN2(n17364), .QN(n17363) );
  INVX0 U18220 ( .INP(n17365), .ZN(n17362) );
  NOR2X0 U18221 ( .IN1(n17364), .IN2(n9016), .QN(n17365) );
  NOR2X0 U18222 ( .IN1(n17366), .IN2(n17367), .QN(n17364) );
  INVX0 U18223 ( .INP(n17368), .ZN(n17367) );
  NAND2X0 U18224 ( .IN1(n18367), .IN2(WX3423), .QN(n17368) );
  NOR2X0 U18225 ( .IN1(WX3423), .IN2(n18367), .QN(n17366) );
  NOR2X0 U18226 ( .IN1(n17369), .IN2(n17370), .QN(n17361) );
  INVX0 U18227 ( .INP(n17371), .ZN(n17370) );
  NAND2X0 U18228 ( .IN1(n9015), .IN2(n10014), .QN(n17371) );
  NOR2X0 U18229 ( .IN1(n10013), .IN2(n9015), .QN(n17369) );
  NOR2X0 U18230 ( .IN1(n17372), .IN2(n17373), .QN(n17337) );
  NOR2X0 U18231 ( .IN1(n9495), .IN2(n11994), .QN(n17373) );
  INVX0 U18232 ( .INP(n2245), .ZN(n11994) );
  NOR2X0 U18233 ( .IN1(DFF_383_n1), .IN2(n9958), .QN(n17372) );
  INVX0 U18234 ( .INP(n2152), .ZN(n11344) );
  INVX0 U18235 ( .INP(n17374), .ZN(WX1839) );
  NAND2X0 U18236 ( .IN1(n10197), .IN2(n9495), .QN(n17374) );
  NOR2X0 U18237 ( .IN1(n10311), .IN2(n17375), .QN(WX1326) );
  NAND2X0 U18238 ( .IN1(n17376), .IN2(n17377), .QN(n17375) );
  NAND2X0 U18239 ( .IN1(n9813), .IN2(CRC_OUT_9_30), .QN(n17377) );
  NAND2X0 U18240 ( .IN1(DFF_190_n1), .IN2(WX837), .QN(n17376) );
  NOR2X0 U18241 ( .IN1(n10311), .IN2(n17378), .QN(WX1324) );
  NAND2X0 U18242 ( .IN1(n17379), .IN2(n17380), .QN(n17378) );
  NAND2X0 U18243 ( .IN1(n9739), .IN2(CRC_OUT_9_29), .QN(n17380) );
  NAND2X0 U18244 ( .IN1(DFF_189_n1), .IN2(WX839), .QN(n17379) );
  NOR2X0 U18245 ( .IN1(n10311), .IN2(n17381), .QN(WX1322) );
  NAND2X0 U18246 ( .IN1(n17382), .IN2(n17383), .QN(n17381) );
  NAND2X0 U18247 ( .IN1(n9747), .IN2(CRC_OUT_9_28), .QN(n17383) );
  NAND2X0 U18248 ( .IN1(DFF_188_n1), .IN2(WX841), .QN(n17382) );
  NOR2X0 U18249 ( .IN1(n10311), .IN2(n17384), .QN(WX1320) );
  NAND2X0 U18250 ( .IN1(n17385), .IN2(n17386), .QN(n17384) );
  NAND2X0 U18251 ( .IN1(n9756), .IN2(CRC_OUT_9_27), .QN(n17386) );
  NAND2X0 U18252 ( .IN1(DFF_187_n1), .IN2(WX843), .QN(n17385) );
  NOR2X0 U18253 ( .IN1(n10311), .IN2(n17387), .QN(WX1318) );
  NAND2X0 U18254 ( .IN1(n17388), .IN2(n17389), .QN(n17387) );
  NAND2X0 U18255 ( .IN1(n9762), .IN2(CRC_OUT_9_26), .QN(n17389) );
  NAND2X0 U18256 ( .IN1(DFF_186_n1), .IN2(WX845), .QN(n17388) );
  NOR2X0 U18257 ( .IN1(n10311), .IN2(n17390), .QN(WX1316) );
  NAND2X0 U18258 ( .IN1(n17391), .IN2(n17392), .QN(n17390) );
  NAND2X0 U18259 ( .IN1(n9765), .IN2(CRC_OUT_9_25), .QN(n17392) );
  NAND2X0 U18260 ( .IN1(DFF_185_n1), .IN2(WX847), .QN(n17391) );
  NOR2X0 U18261 ( .IN1(n10312), .IN2(n17393), .QN(WX1314) );
  NAND2X0 U18262 ( .IN1(n17394), .IN2(n17395), .QN(n17393) );
  NAND2X0 U18263 ( .IN1(n9774), .IN2(CRC_OUT_9_24), .QN(n17395) );
  NAND2X0 U18264 ( .IN1(DFF_184_n1), .IN2(WX849), .QN(n17394) );
  NOR2X0 U18265 ( .IN1(n10312), .IN2(n17396), .QN(WX1312) );
  NAND2X0 U18266 ( .IN1(n17397), .IN2(n17398), .QN(n17396) );
  NAND2X0 U18267 ( .IN1(n9783), .IN2(CRC_OUT_9_23), .QN(n17398) );
  NAND2X0 U18268 ( .IN1(DFF_183_n1), .IN2(WX851), .QN(n17397) );
  NOR2X0 U18269 ( .IN1(n10312), .IN2(n17399), .QN(WX1310) );
  NAND2X0 U18270 ( .IN1(n17400), .IN2(n17401), .QN(n17399) );
  NAND2X0 U18271 ( .IN1(n9785), .IN2(CRC_OUT_9_22), .QN(n17401) );
  NAND2X0 U18272 ( .IN1(DFF_182_n1), .IN2(WX853), .QN(n17400) );
  NOR2X0 U18273 ( .IN1(n10312), .IN2(n17402), .QN(WX1308) );
  NAND2X0 U18274 ( .IN1(n17403), .IN2(n17404), .QN(n17402) );
  NAND2X0 U18275 ( .IN1(n9800), .IN2(CRC_OUT_9_21), .QN(n17404) );
  NAND2X0 U18276 ( .IN1(DFF_181_n1), .IN2(WX855), .QN(n17403) );
  NOR2X0 U18277 ( .IN1(n10312), .IN2(n17405), .QN(WX1306) );
  NAND2X0 U18278 ( .IN1(n17406), .IN2(n17407), .QN(n17405) );
  NAND2X0 U18279 ( .IN1(n9806), .IN2(CRC_OUT_9_20), .QN(n17407) );
  NAND2X0 U18280 ( .IN1(DFF_180_n1), .IN2(WX857), .QN(n17406) );
  NOR2X0 U18281 ( .IN1(n10312), .IN2(n17408), .QN(WX1304) );
  NOR2X0 U18282 ( .IN1(n17409), .IN2(n17410), .QN(n17408) );
  NOR2X0 U18283 ( .IN1(test_so10), .IN2(WX859), .QN(n17410) );
  INVX0 U18284 ( .INP(n17411), .ZN(n17409) );
  NAND2X0 U18285 ( .IN1(WX859), .IN2(test_so10), .QN(n17411) );
  NOR2X0 U18286 ( .IN1(n10312), .IN2(n17412), .QN(WX1302) );
  NAND2X0 U18287 ( .IN1(n17413), .IN2(n17414), .QN(n17412) );
  NAND2X0 U18288 ( .IN1(n9744), .IN2(CRC_OUT_9_18), .QN(n17414) );
  NAND2X0 U18289 ( .IN1(DFF_178_n1), .IN2(WX861), .QN(n17413) );
  NOR2X0 U18290 ( .IN1(n10312), .IN2(n17415), .QN(WX1300) );
  NAND2X0 U18291 ( .IN1(n17416), .IN2(n17417), .QN(n17415) );
  NAND2X0 U18292 ( .IN1(n9759), .IN2(CRC_OUT_9_17), .QN(n17417) );
  NAND2X0 U18293 ( .IN1(DFF_177_n1), .IN2(WX863), .QN(n17416) );
  NOR2X0 U18294 ( .IN1(n10312), .IN2(n17418), .QN(WX1298) );
  NAND2X0 U18295 ( .IN1(n17419), .IN2(n17420), .QN(n17418) );
  NAND2X0 U18296 ( .IN1(n9771), .IN2(CRC_OUT_9_16), .QN(n17420) );
  NAND2X0 U18297 ( .IN1(DFF_176_n1), .IN2(WX865), .QN(n17419) );
  NOR2X0 U18298 ( .IN1(n10312), .IN2(n17421), .QN(WX1296) );
  NAND2X0 U18299 ( .IN1(n17422), .IN2(n17423), .QN(n17421) );
  INVX0 U18300 ( .INP(n17424), .ZN(n17423) );
  NOR2X0 U18301 ( .IN1(CRC_OUT_9_15), .IN2(n17425), .QN(n17424) );
  NAND2X0 U18302 ( .IN1(n17425), .IN2(CRC_OUT_9_15), .QN(n17422) );
  NAND2X0 U18303 ( .IN1(n17426), .IN2(n17427), .QN(n17425) );
  NAND2X0 U18304 ( .IN1(test_so8), .IN2(CRC_OUT_9_31), .QN(n17427) );
  NAND2X0 U18305 ( .IN1(DFF_191_n1), .IN2(n9851), .QN(n17426) );
  NOR2X0 U18306 ( .IN1(n10312), .IN2(n17428), .QN(WX1294) );
  NAND2X0 U18307 ( .IN1(n17429), .IN2(n17430), .QN(n17428) );
  NAND2X0 U18308 ( .IN1(n9803), .IN2(CRC_OUT_9_14), .QN(n17430) );
  NAND2X0 U18309 ( .IN1(DFF_174_n1), .IN2(WX869), .QN(n17429) );
  NOR2X0 U18310 ( .IN1(n10312), .IN2(n17431), .QN(WX1292) );
  NAND2X0 U18311 ( .IN1(n17432), .IN2(n17433), .QN(n17431) );
  NAND2X0 U18312 ( .IN1(n9815), .IN2(CRC_OUT_9_13), .QN(n17433) );
  NAND2X0 U18313 ( .IN1(DFF_173_n1), .IN2(WX871), .QN(n17432) );
  NOR2X0 U18314 ( .IN1(n10312), .IN2(n17434), .QN(WX1290) );
  NAND2X0 U18315 ( .IN1(n17435), .IN2(n17436), .QN(n17434) );
  NAND2X0 U18316 ( .IN1(n9750), .IN2(CRC_OUT_9_12), .QN(n17436) );
  NAND2X0 U18317 ( .IN1(DFF_172_n1), .IN2(WX873), .QN(n17435) );
  NOR2X0 U18318 ( .IN1(n10313), .IN2(n17437), .QN(WX1288) );
  NAND2X0 U18319 ( .IN1(n17438), .IN2(n17439), .QN(n17437) );
  NAND2X0 U18320 ( .IN1(n9777), .IN2(CRC_OUT_9_11), .QN(n17439) );
  NAND2X0 U18321 ( .IN1(DFF_171_n1), .IN2(WX875), .QN(n17438) );
  NOR2X0 U18322 ( .IN1(n10313), .IN2(n17440), .QN(WX1286) );
  NOR2X0 U18323 ( .IN1(n17441), .IN2(n17442), .QN(n17440) );
  INVX0 U18324 ( .INP(n17443), .ZN(n17442) );
  NAND2X0 U18325 ( .IN1(CRC_OUT_9_10), .IN2(n17444), .QN(n17443) );
  NOR2X0 U18326 ( .IN1(n17444), .IN2(CRC_OUT_9_10), .QN(n17441) );
  NAND2X0 U18327 ( .IN1(n17445), .IN2(n17446), .QN(n17444) );
  NAND2X0 U18328 ( .IN1(n9823), .IN2(CRC_OUT_9_31), .QN(n17446) );
  NAND2X0 U18329 ( .IN1(DFF_191_n1), .IN2(WX877), .QN(n17445) );
  NOR2X0 U18330 ( .IN1(n10313), .IN2(n17447), .QN(WX1284) );
  NAND2X0 U18331 ( .IN1(n17448), .IN2(n17449), .QN(n17447) );
  NAND2X0 U18332 ( .IN1(n9768), .IN2(CRC_OUT_9_9), .QN(n17449) );
  NAND2X0 U18333 ( .IN1(DFF_169_n1), .IN2(WX879), .QN(n17448) );
  NOR2X0 U18334 ( .IN1(n10313), .IN2(n17450), .QN(WX1282) );
  NAND2X0 U18335 ( .IN1(n17451), .IN2(n17452), .QN(n17450) );
  NAND2X0 U18336 ( .IN1(n9781), .IN2(CRC_OUT_9_8), .QN(n17452) );
  NAND2X0 U18337 ( .IN1(DFF_168_n1), .IN2(WX881), .QN(n17451) );
  NOR2X0 U18338 ( .IN1(n10313), .IN2(n17453), .QN(WX1280) );
  NAND2X0 U18339 ( .IN1(n17454), .IN2(n17455), .QN(n17453) );
  NAND2X0 U18340 ( .IN1(n9790), .IN2(CRC_OUT_9_7), .QN(n17455) );
  NAND2X0 U18341 ( .IN1(DFF_167_n1), .IN2(WX883), .QN(n17454) );
  NOR2X0 U18342 ( .IN1(n10313), .IN2(n17456), .QN(WX1278) );
  NAND2X0 U18343 ( .IN1(n17457), .IN2(n17458), .QN(n17456) );
  NAND2X0 U18344 ( .IN1(n9821), .IN2(CRC_OUT_9_6), .QN(n17458) );
  NAND2X0 U18345 ( .IN1(DFF_166_n1), .IN2(WX885), .QN(n17457) );
  NOR2X0 U18346 ( .IN1(n10313), .IN2(n17459), .QN(WX1276) );
  NAND2X0 U18347 ( .IN1(n17460), .IN2(n17461), .QN(n17459) );
  NAND2X0 U18348 ( .IN1(n9808), .IN2(CRC_OUT_9_5), .QN(n17461) );
  NAND2X0 U18349 ( .IN1(DFF_165_n1), .IN2(WX887), .QN(n17460) );
  NOR2X0 U18350 ( .IN1(n10313), .IN2(n17462), .QN(WX1274) );
  NAND2X0 U18351 ( .IN1(n17463), .IN2(n17464), .QN(n17462) );
  NAND2X0 U18352 ( .IN1(n9793), .IN2(CRC_OUT_9_4), .QN(n17464) );
  NAND2X0 U18353 ( .IN1(DFF_164_n1), .IN2(WX889), .QN(n17463) );
  NOR2X0 U18354 ( .IN1(n10313), .IN2(n17465), .QN(WX1272) );
  NOR2X0 U18355 ( .IN1(n17466), .IN2(n17467), .QN(n17465) );
  INVX0 U18356 ( .INP(n17468), .ZN(n17467) );
  NAND2X0 U18357 ( .IN1(CRC_OUT_9_3), .IN2(n17469), .QN(n17468) );
  NOR2X0 U18358 ( .IN1(n17469), .IN2(CRC_OUT_9_3), .QN(n17466) );
  NAND2X0 U18359 ( .IN1(n17470), .IN2(n17471), .QN(n17469) );
  NAND2X0 U18360 ( .IN1(n9796), .IN2(CRC_OUT_9_31), .QN(n17471) );
  NAND2X0 U18361 ( .IN1(DFF_191_n1), .IN2(WX891), .QN(n17470) );
  NOR2X0 U18362 ( .IN1(n10313), .IN2(n17472), .QN(WX1270) );
  NAND2X0 U18363 ( .IN1(n17473), .IN2(n17474), .QN(n17472) );
  NAND2X0 U18364 ( .IN1(n9741), .IN2(CRC_OUT_9_2), .QN(n17474) );
  NAND2X0 U18365 ( .IN1(DFF_162_n1), .IN2(WX893), .QN(n17473) );
  NOR2X0 U18366 ( .IN1(n10313), .IN2(n17475), .QN(WX1268) );
  NOR2X0 U18367 ( .IN1(n17476), .IN2(n17477), .QN(n17475) );
  NOR2X0 U18368 ( .IN1(test_so9), .IN2(WX895), .QN(n17477) );
  INVX0 U18369 ( .INP(n17478), .ZN(n17476) );
  NAND2X0 U18370 ( .IN1(WX895), .IN2(test_so9), .QN(n17478) );
  NOR2X0 U18371 ( .IN1(n10313), .IN2(n17479), .QN(WX1266) );
  NAND2X0 U18372 ( .IN1(n17480), .IN2(n17481), .QN(n17479) );
  NAND2X0 U18373 ( .IN1(n9752), .IN2(CRC_OUT_9_0), .QN(n17481) );
  NAND2X0 U18374 ( .IN1(DFF_160_n1), .IN2(WX897), .QN(n17480) );
  NOR2X0 U18375 ( .IN1(n10313), .IN2(n17482), .QN(WX1264) );
  NAND2X0 U18376 ( .IN1(n17483), .IN2(n17484), .QN(n17482) );
  NAND2X0 U18377 ( .IN1(n9827), .IN2(CRC_OUT_9_31), .QN(n17484) );
  NAND2X0 U18378 ( .IN1(DFF_191_n1), .IN2(WX899), .QN(n17483) );
  NOR2X0 U18379 ( .IN1(n10314), .IN2(n17485), .QN(WX11670) );
  NAND2X0 U18380 ( .IN1(n17486), .IN2(n17487), .QN(n17485) );
  NAND2X0 U18381 ( .IN1(n9525), .IN2(CRC_OUT_1_30), .QN(n17487) );
  NAND2X0 U18382 ( .IN1(DFF_1726_n1), .IN2(WX11181), .QN(n17486) );
  NOR2X0 U18383 ( .IN1(n10314), .IN2(n17488), .QN(WX11668) );
  NAND2X0 U18384 ( .IN1(n17489), .IN2(n17490), .QN(n17488) );
  NAND2X0 U18385 ( .IN1(n9526), .IN2(CRC_OUT_1_29), .QN(n17490) );
  NAND2X0 U18386 ( .IN1(DFF_1725_n1), .IN2(WX11183), .QN(n17489) );
  NOR2X0 U18387 ( .IN1(n10314), .IN2(n17491), .QN(WX11666) );
  NAND2X0 U18388 ( .IN1(n17492), .IN2(n17493), .QN(n17491) );
  NAND2X0 U18389 ( .IN1(n9527), .IN2(CRC_OUT_1_28), .QN(n17493) );
  NAND2X0 U18390 ( .IN1(DFF_1724_n1), .IN2(WX11185), .QN(n17492) );
  NOR2X0 U18391 ( .IN1(n10314), .IN2(n17494), .QN(WX11664) );
  NAND2X0 U18392 ( .IN1(n17495), .IN2(n17496), .QN(n17494) );
  NAND2X0 U18393 ( .IN1(n9528), .IN2(CRC_OUT_1_27), .QN(n17496) );
  NAND2X0 U18394 ( .IN1(DFF_1723_n1), .IN2(WX11187), .QN(n17495) );
  NOR2X0 U18395 ( .IN1(n10314), .IN2(n17497), .QN(WX11662) );
  NAND2X0 U18396 ( .IN1(n17498), .IN2(n17499), .QN(n17497) );
  NAND2X0 U18397 ( .IN1(n9529), .IN2(CRC_OUT_1_26), .QN(n17499) );
  NAND2X0 U18398 ( .IN1(DFF_1722_n1), .IN2(WX11189), .QN(n17498) );
  NOR2X0 U18399 ( .IN1(n10314), .IN2(n17500), .QN(WX11660) );
  NAND2X0 U18400 ( .IN1(n17501), .IN2(n17502), .QN(n17500) );
  NAND2X0 U18401 ( .IN1(n9530), .IN2(CRC_OUT_1_25), .QN(n17502) );
  NAND2X0 U18402 ( .IN1(DFF_1721_n1), .IN2(WX11191), .QN(n17501) );
  NOR2X0 U18403 ( .IN1(n10314), .IN2(n17503), .QN(WX11658) );
  NAND2X0 U18404 ( .IN1(n17504), .IN2(n17505), .QN(n17503) );
  NAND2X0 U18405 ( .IN1(n9531), .IN2(CRC_OUT_1_24), .QN(n17505) );
  NAND2X0 U18406 ( .IN1(DFF_1720_n1), .IN2(WX11193), .QN(n17504) );
  NOR2X0 U18407 ( .IN1(n10314), .IN2(n17506), .QN(WX11656) );
  NAND2X0 U18408 ( .IN1(n17507), .IN2(n17508), .QN(n17506) );
  NAND2X0 U18409 ( .IN1(n9532), .IN2(CRC_OUT_1_23), .QN(n17508) );
  NAND2X0 U18410 ( .IN1(DFF_1719_n1), .IN2(WX11195), .QN(n17507) );
  NOR2X0 U18411 ( .IN1(n10314), .IN2(n17509), .QN(WX11654) );
  NAND2X0 U18412 ( .IN1(n17510), .IN2(n17511), .QN(n17509) );
  NAND2X0 U18413 ( .IN1(n9533), .IN2(CRC_OUT_1_22), .QN(n17511) );
  NAND2X0 U18414 ( .IN1(DFF_1718_n1), .IN2(WX11197), .QN(n17510) );
  NOR2X0 U18415 ( .IN1(n10314), .IN2(n17512), .QN(WX11652) );
  NAND2X0 U18416 ( .IN1(n17513), .IN2(n17514), .QN(n17512) );
  NAND2X0 U18417 ( .IN1(n9534), .IN2(CRC_OUT_1_21), .QN(n17514) );
  NAND2X0 U18418 ( .IN1(DFF_1717_n1), .IN2(WX11199), .QN(n17513) );
  NOR2X0 U18419 ( .IN1(n10314), .IN2(n17515), .QN(WX11650) );
  NAND2X0 U18420 ( .IN1(n17516), .IN2(n17517), .QN(n17515) );
  NAND2X0 U18421 ( .IN1(n9535), .IN2(CRC_OUT_1_20), .QN(n17517) );
  NAND2X0 U18422 ( .IN1(DFF_1716_n1), .IN2(WX11201), .QN(n17516) );
  NOR2X0 U18423 ( .IN1(n10314), .IN2(n17518), .QN(WX11648) );
  NAND2X0 U18424 ( .IN1(n17519), .IN2(n17520), .QN(n17518) );
  NAND2X0 U18425 ( .IN1(n9536), .IN2(CRC_OUT_1_19), .QN(n17520) );
  NAND2X0 U18426 ( .IN1(DFF_1715_n1), .IN2(WX11203), .QN(n17519) );
  NOR2X0 U18427 ( .IN1(n10314), .IN2(n17521), .QN(WX11646) );
  NOR2X0 U18428 ( .IN1(n17522), .IN2(n17523), .QN(n17521) );
  NOR2X0 U18429 ( .IN1(test_so97), .IN2(CRC_OUT_1_18), .QN(n17523) );
  NOR2X0 U18430 ( .IN1(DFF_1714_n1), .IN2(n9839), .QN(n17522) );
  NOR2X0 U18431 ( .IN1(n10315), .IN2(n17524), .QN(WX11644) );
  NAND2X0 U18432 ( .IN1(n17525), .IN2(n17526), .QN(n17524) );
  NAND2X0 U18433 ( .IN1(n9537), .IN2(CRC_OUT_1_17), .QN(n17526) );
  NAND2X0 U18434 ( .IN1(DFF_1713_n1), .IN2(WX11207), .QN(n17525) );
  NOR2X0 U18435 ( .IN1(n10315), .IN2(n17527), .QN(WX11642) );
  NAND2X0 U18436 ( .IN1(n17528), .IN2(n17529), .QN(n17527) );
  NAND2X0 U18437 ( .IN1(n9538), .IN2(CRC_OUT_1_16), .QN(n17529) );
  NAND2X0 U18438 ( .IN1(DFF_1712_n1), .IN2(WX11209), .QN(n17528) );
  NOR2X0 U18439 ( .IN1(n10315), .IN2(n17530), .QN(WX11640) );
  NAND2X0 U18440 ( .IN1(n17531), .IN2(n17532), .QN(n17530) );
  INVX0 U18441 ( .INP(n17533), .ZN(n17532) );
  NOR2X0 U18442 ( .IN1(CRC_OUT_1_15), .IN2(n17534), .QN(n17533) );
  NAND2X0 U18443 ( .IN1(n17534), .IN2(CRC_OUT_1_15), .QN(n17531) );
  NAND2X0 U18444 ( .IN1(n17535), .IN2(n17536), .QN(n17534) );
  NAND2X0 U18445 ( .IN1(test_so100), .IN2(WX11211), .QN(n17536) );
  NAND2X0 U18446 ( .IN1(n9496), .IN2(n9838), .QN(n17535) );
  NOR2X0 U18447 ( .IN1(n10315), .IN2(n17537), .QN(WX11638) );
  NOR2X0 U18448 ( .IN1(n17538), .IN2(n17539), .QN(n17537) );
  NOR2X0 U18449 ( .IN1(test_so99), .IN2(WX11213), .QN(n17539) );
  INVX0 U18450 ( .INP(n17540), .ZN(n17538) );
  NAND2X0 U18451 ( .IN1(WX11213), .IN2(test_so99), .QN(n17540) );
  NOR2X0 U18452 ( .IN1(n10315), .IN2(n17541), .QN(WX11636) );
  NAND2X0 U18453 ( .IN1(n17542), .IN2(n17543), .QN(n17541) );
  NAND2X0 U18454 ( .IN1(n9540), .IN2(CRC_OUT_1_13), .QN(n17543) );
  NAND2X0 U18455 ( .IN1(DFF_1709_n1), .IN2(WX11215), .QN(n17542) );
  NOR2X0 U18456 ( .IN1(n10315), .IN2(n17544), .QN(WX11634) );
  NAND2X0 U18457 ( .IN1(n17545), .IN2(n17546), .QN(n17544) );
  NAND2X0 U18458 ( .IN1(n9541), .IN2(CRC_OUT_1_12), .QN(n17546) );
  NAND2X0 U18459 ( .IN1(DFF_1708_n1), .IN2(WX11217), .QN(n17545) );
  NOR2X0 U18460 ( .IN1(n10315), .IN2(n17547), .QN(WX11632) );
  NAND2X0 U18461 ( .IN1(n17548), .IN2(n17549), .QN(n17547) );
  NAND2X0 U18462 ( .IN1(n9542), .IN2(CRC_OUT_1_11), .QN(n17549) );
  NAND2X0 U18463 ( .IN1(DFF_1707_n1), .IN2(WX11219), .QN(n17548) );
  NOR2X0 U18464 ( .IN1(n10315), .IN2(n17550), .QN(WX11630) );
  NAND2X0 U18465 ( .IN1(n17551), .IN2(n17552), .QN(n17550) );
  INVX0 U18466 ( .INP(n17553), .ZN(n17552) );
  NOR2X0 U18467 ( .IN1(CRC_OUT_1_10), .IN2(n17554), .QN(n17553) );
  NAND2X0 U18468 ( .IN1(n17554), .IN2(CRC_OUT_1_10), .QN(n17551) );
  NAND2X0 U18469 ( .IN1(n17555), .IN2(n17556), .QN(n17554) );
  NAND2X0 U18470 ( .IN1(test_so100), .IN2(WX11221), .QN(n17556) );
  NAND2X0 U18471 ( .IN1(n9497), .IN2(n9838), .QN(n17555) );
  NOR2X0 U18472 ( .IN1(n10315), .IN2(n17557), .QN(WX11628) );
  NAND2X0 U18473 ( .IN1(n17558), .IN2(n17559), .QN(n17557) );
  NAND2X0 U18474 ( .IN1(n9543), .IN2(CRC_OUT_1_9), .QN(n17559) );
  NAND2X0 U18475 ( .IN1(DFF_1705_n1), .IN2(WX11223), .QN(n17558) );
  NOR2X0 U18476 ( .IN1(n10315), .IN2(n17560), .QN(WX11626) );
  NAND2X0 U18477 ( .IN1(n17561), .IN2(n17562), .QN(n17560) );
  NAND2X0 U18478 ( .IN1(n9544), .IN2(CRC_OUT_1_8), .QN(n17562) );
  NAND2X0 U18479 ( .IN1(DFF_1704_n1), .IN2(WX11225), .QN(n17561) );
  NOR2X0 U18480 ( .IN1(n10315), .IN2(n17563), .QN(WX11624) );
  NAND2X0 U18481 ( .IN1(n17564), .IN2(n17565), .QN(n17563) );
  NAND2X0 U18482 ( .IN1(n9545), .IN2(CRC_OUT_1_7), .QN(n17565) );
  NAND2X0 U18483 ( .IN1(DFF_1703_n1), .IN2(WX11227), .QN(n17564) );
  NOR2X0 U18484 ( .IN1(n10315), .IN2(n17566), .QN(WX11622) );
  NAND2X0 U18485 ( .IN1(n17567), .IN2(n17568), .QN(n17566) );
  NAND2X0 U18486 ( .IN1(n9546), .IN2(CRC_OUT_1_6), .QN(n17568) );
  NAND2X0 U18487 ( .IN1(DFF_1702_n1), .IN2(WX11229), .QN(n17567) );
  NOR2X0 U18488 ( .IN1(n10315), .IN2(n17569), .QN(WX11620) );
  NAND2X0 U18489 ( .IN1(n17570), .IN2(n17571), .QN(n17569) );
  NAND2X0 U18490 ( .IN1(n9547), .IN2(CRC_OUT_1_5), .QN(n17571) );
  NAND2X0 U18491 ( .IN1(DFF_1701_n1), .IN2(WX11231), .QN(n17570) );
  NOR2X0 U18492 ( .IN1(n10316), .IN2(n17572), .QN(WX11618) );
  NAND2X0 U18493 ( .IN1(n17573), .IN2(n17574), .QN(n17572) );
  NAND2X0 U18494 ( .IN1(n9548), .IN2(CRC_OUT_1_4), .QN(n17574) );
  NAND2X0 U18495 ( .IN1(DFF_1700_n1), .IN2(WX11233), .QN(n17573) );
  NOR2X0 U18496 ( .IN1(n10316), .IN2(n17575), .QN(WX11616) );
  NAND2X0 U18497 ( .IN1(n17576), .IN2(n17577), .QN(n17575) );
  INVX0 U18498 ( .INP(n17578), .ZN(n17577) );
  NOR2X0 U18499 ( .IN1(CRC_OUT_1_3), .IN2(n17579), .QN(n17578) );
  NAND2X0 U18500 ( .IN1(n17579), .IN2(CRC_OUT_1_3), .QN(n17576) );
  NAND2X0 U18501 ( .IN1(n17580), .IN2(n17581), .QN(n17579) );
  NAND2X0 U18502 ( .IN1(test_so100), .IN2(WX11235), .QN(n17581) );
  NAND2X0 U18503 ( .IN1(n9498), .IN2(n9838), .QN(n17580) );
  NOR2X0 U18504 ( .IN1(n10316), .IN2(n17582), .QN(WX11614) );
  NAND2X0 U18505 ( .IN1(n17583), .IN2(n17584), .QN(n17582) );
  NAND2X0 U18506 ( .IN1(n9549), .IN2(CRC_OUT_1_2), .QN(n17584) );
  NAND2X0 U18507 ( .IN1(DFF_1698_n1), .IN2(WX11237), .QN(n17583) );
  NOR2X0 U18508 ( .IN1(n10316), .IN2(n17585), .QN(WX11612) );
  NOR2X0 U18509 ( .IN1(n17586), .IN2(n17587), .QN(n17585) );
  NOR2X0 U18510 ( .IN1(test_so98), .IN2(CRC_OUT_1_1), .QN(n17587) );
  NOR2X0 U18511 ( .IN1(DFF_1697_n1), .IN2(n9847), .QN(n17586) );
  NOR2X0 U18512 ( .IN1(n10316), .IN2(n17588), .QN(WX11610) );
  NAND2X0 U18513 ( .IN1(n17589), .IN2(n17590), .QN(n17588) );
  NAND2X0 U18514 ( .IN1(n9550), .IN2(CRC_OUT_1_0), .QN(n17590) );
  NAND2X0 U18515 ( .IN1(DFF_1696_n1), .IN2(WX11241), .QN(n17589) );
  NOR2X0 U18516 ( .IN1(n10316), .IN2(n17591), .QN(WX11608) );
  NOR2X0 U18517 ( .IN1(n17592), .IN2(n17593), .QN(n17591) );
  NOR2X0 U18518 ( .IN1(test_so100), .IN2(WX11243), .QN(n17593) );
  NOR2X0 U18519 ( .IN1(n9517), .IN2(n9838), .QN(n17592) );
  NOR2X0 U18520 ( .IN1(n18472), .IN2(n10240), .QN(WX11082) );
  NOR2X0 U18521 ( .IN1(n18471), .IN2(n10240), .QN(WX11080) );
  NOR2X0 U18522 ( .IN1(n18470), .IN2(n10240), .QN(WX11078) );
  NOR2X0 U18523 ( .IN1(n18469), .IN2(n10240), .QN(WX11076) );
  NOR2X0 U18524 ( .IN1(n18468), .IN2(n10239), .QN(WX11074) );
  NOR2X0 U18525 ( .IN1(n18467), .IN2(n10239), .QN(WX11072) );
  NOR2X0 U18526 ( .IN1(n18466), .IN2(n10239), .QN(WX11070) );
  NOR2X0 U18527 ( .IN1(n18465), .IN2(n10239), .QN(WX11068) );
  NOR2X0 U18528 ( .IN1(n18464), .IN2(n10239), .QN(WX11066) );
  NOR2X0 U18529 ( .IN1(n10316), .IN2(n9846), .QN(WX11064) );
  NOR2X0 U18530 ( .IN1(n18463), .IN2(n10239), .QN(WX11062) );
  NOR2X0 U18531 ( .IN1(n18462), .IN2(n10239), .QN(WX11060) );
  NOR2X0 U18532 ( .IN1(n18461), .IN2(n10239), .QN(WX11058) );
  NOR2X0 U18533 ( .IN1(n18460), .IN2(n10239), .QN(WX11056) );
  NOR2X0 U18534 ( .IN1(n18459), .IN2(n10239), .QN(WX11054) );
  NOR2X0 U18535 ( .IN1(n18458), .IN2(n10241), .QN(WX11052) );
  NOR2X0 U18536 ( .IN1(n10316), .IN2(WX10829), .QN(WX10890) );
  NOR2X0 U18537 ( .IN1(n10316), .IN2(n17594), .QN(WX10377) );
  NOR2X0 U18538 ( .IN1(n17595), .IN2(n17596), .QN(n17594) );
  INVX0 U18539 ( .INP(n17597), .ZN(n17596) );
  NAND2X0 U18540 ( .IN1(n9833), .IN2(DFF_1534_n1), .QN(n17597) );
  NOR2X0 U18541 ( .IN1(DFF_1534_n1), .IN2(n9833), .QN(n17595) );
  NOR2X0 U18542 ( .IN1(n10316), .IN2(n17598), .QN(WX10375) );
  NAND2X0 U18543 ( .IN1(n17599), .IN2(n17600), .QN(n17598) );
  INVX0 U18544 ( .INP(n17601), .ZN(n17600) );
  NOR2X0 U18545 ( .IN1(WX9890), .IN2(DFF_1533_n1), .QN(n17601) );
  NAND2X0 U18546 ( .IN1(DFF_1533_n1), .IN2(WX9890), .QN(n17599) );
  NOR2X0 U18547 ( .IN1(n10316), .IN2(n17602), .QN(WX10373) );
  NAND2X0 U18548 ( .IN1(n17603), .IN2(n17604), .QN(n17602) );
  INVX0 U18549 ( .INP(n17605), .ZN(n17604) );
  NOR2X0 U18550 ( .IN1(WX9892), .IN2(DFF_1532_n1), .QN(n17605) );
  NAND2X0 U18551 ( .IN1(DFF_1532_n1), .IN2(WX9892), .QN(n17603) );
  NOR2X0 U18552 ( .IN1(n10316), .IN2(n17606), .QN(WX10371) );
  NAND2X0 U18553 ( .IN1(n17607), .IN2(n17608), .QN(n17606) );
  INVX0 U18554 ( .INP(n17609), .ZN(n17608) );
  NOR2X0 U18555 ( .IN1(WX9894), .IN2(DFF_1531_n1), .QN(n17609) );
  NAND2X0 U18556 ( .IN1(DFF_1531_n1), .IN2(WX9894), .QN(n17607) );
  NOR2X0 U18557 ( .IN1(n10316), .IN2(n17610), .QN(WX10369) );
  NAND2X0 U18558 ( .IN1(n17611), .IN2(n17612), .QN(n17610) );
  INVX0 U18559 ( .INP(n17613), .ZN(n17612) );
  NOR2X0 U18560 ( .IN1(WX9896), .IN2(DFF_1530_n1), .QN(n17613) );
  NAND2X0 U18561 ( .IN1(DFF_1530_n1), .IN2(WX9896), .QN(n17611) );
  NOR2X0 U18562 ( .IN1(n10317), .IN2(n17614), .QN(WX10367) );
  NAND2X0 U18563 ( .IN1(n17615), .IN2(n17616), .QN(n17614) );
  INVX0 U18564 ( .INP(n17617), .ZN(n17616) );
  NOR2X0 U18565 ( .IN1(WX9898), .IN2(DFF_1529_n1), .QN(n17617) );
  NAND2X0 U18566 ( .IN1(DFF_1529_n1), .IN2(WX9898), .QN(n17615) );
  NOR2X0 U18567 ( .IN1(n10317), .IN2(n17618), .QN(WX10365) );
  NAND2X0 U18568 ( .IN1(n17619), .IN2(n17620), .QN(n17618) );
  INVX0 U18569 ( .INP(n17621), .ZN(n17620) );
  NOR2X0 U18570 ( .IN1(WX9900), .IN2(DFF_1528_n1), .QN(n17621) );
  NAND2X0 U18571 ( .IN1(DFF_1528_n1), .IN2(WX9900), .QN(n17619) );
  NOR2X0 U18572 ( .IN1(n10317), .IN2(n17622), .QN(WX10363) );
  NAND2X0 U18573 ( .IN1(n17623), .IN2(n17624), .QN(n17622) );
  INVX0 U18574 ( .INP(n17625), .ZN(n17624) );
  NOR2X0 U18575 ( .IN1(WX9902), .IN2(DFF_1527_n1), .QN(n17625) );
  NAND2X0 U18576 ( .IN1(DFF_1527_n1), .IN2(WX9902), .QN(n17623) );
  NOR2X0 U18577 ( .IN1(n10317), .IN2(n17626), .QN(WX10361) );
  NAND2X0 U18578 ( .IN1(n17627), .IN2(n17628), .QN(n17626) );
  INVX0 U18579 ( .INP(n17629), .ZN(n17628) );
  NOR2X0 U18580 ( .IN1(WX9904), .IN2(DFF_1526_n1), .QN(n17629) );
  NAND2X0 U18581 ( .IN1(DFF_1526_n1), .IN2(WX9904), .QN(n17627) );
  NOR2X0 U18582 ( .IN1(n10317), .IN2(n17630), .QN(WX10359) );
  NAND2X0 U18583 ( .IN1(n17631), .IN2(n17632), .QN(n17630) );
  INVX0 U18584 ( .INP(n17633), .ZN(n17632) );
  NOR2X0 U18585 ( .IN1(WX9906), .IN2(DFF_1525_n1), .QN(n17633) );
  NAND2X0 U18586 ( .IN1(DFF_1525_n1), .IN2(WX9906), .QN(n17631) );
  NOR2X0 U18587 ( .IN1(n10317), .IN2(n17634), .QN(WX10357) );
  NAND2X0 U18588 ( .IN1(n17635), .IN2(n17636), .QN(n17634) );
  INVX0 U18589 ( .INP(n17637), .ZN(n17636) );
  NOR2X0 U18590 ( .IN1(WX9908), .IN2(DFF_1524_n1), .QN(n17637) );
  NAND2X0 U18591 ( .IN1(DFF_1524_n1), .IN2(WX9908), .QN(n17635) );
  NOR2X0 U18592 ( .IN1(n10317), .IN2(n17638), .QN(WX10355) );
  NOR2X0 U18593 ( .IN1(n17639), .IN2(n17640), .QN(n17638) );
  NOR2X0 U18594 ( .IN1(test_so88), .IN2(WX9910), .QN(n17640) );
  NOR2X0 U18595 ( .IN1(n9561), .IN2(n9863), .QN(n17639) );
  NOR2X0 U18596 ( .IN1(n10317), .IN2(n17641), .QN(WX10353) );
  NAND2X0 U18597 ( .IN1(n17642), .IN2(n17643), .QN(n17641) );
  INVX0 U18598 ( .INP(n17644), .ZN(n17643) );
  NOR2X0 U18599 ( .IN1(WX9912), .IN2(DFF_1522_n1), .QN(n17644) );
  NAND2X0 U18600 ( .IN1(DFF_1522_n1), .IN2(WX9912), .QN(n17642) );
  NOR2X0 U18601 ( .IN1(n10317), .IN2(n17645), .QN(WX10351) );
  NAND2X0 U18602 ( .IN1(n17646), .IN2(n17647), .QN(n17645) );
  NAND2X0 U18603 ( .IN1(n9563), .IN2(CRC_OUT_2_17), .QN(n17647) );
  NAND2X0 U18604 ( .IN1(DFF_1521_n1), .IN2(WX9914), .QN(n17646) );
  NOR2X0 U18605 ( .IN1(n10317), .IN2(n17648), .QN(WX10349) );
  NAND2X0 U18606 ( .IN1(n17649), .IN2(n17650), .QN(n17648) );
  INVX0 U18607 ( .INP(n17651), .ZN(n17650) );
  NOR2X0 U18608 ( .IN1(WX9916), .IN2(DFF_1520_n1), .QN(n17651) );
  NAND2X0 U18609 ( .IN1(DFF_1520_n1), .IN2(WX9916), .QN(n17649) );
  NOR2X0 U18610 ( .IN1(n10317), .IN2(n17652), .QN(WX10347) );
  NOR2X0 U18611 ( .IN1(n17653), .IN2(n17654), .QN(n17652) );
  NOR2X0 U18612 ( .IN1(DFF_1519_n1), .IN2(n17655), .QN(n17654) );
  INVX0 U18613 ( .INP(n17656), .ZN(n17653) );
  NAND2X0 U18614 ( .IN1(n17655), .IN2(DFF_1519_n1), .QN(n17656) );
  NOR2X0 U18615 ( .IN1(n17657), .IN2(n17658), .QN(n17655) );
  NOR2X0 U18616 ( .IN1(WX9918), .IN2(DFF_1535_n1), .QN(n17658) );
  NOR2X0 U18617 ( .IN1(CRC_OUT_2_31), .IN2(n9499), .QN(n17657) );
  NOR2X0 U18618 ( .IN1(n10317), .IN2(n17659), .QN(WX10345) );
  NAND2X0 U18619 ( .IN1(n17660), .IN2(n17661), .QN(n17659) );
  INVX0 U18620 ( .INP(n17662), .ZN(n17661) );
  NOR2X0 U18621 ( .IN1(WX9920), .IN2(DFF_1518_n1), .QN(n17662) );
  NAND2X0 U18622 ( .IN1(DFF_1518_n1), .IN2(WX9920), .QN(n17660) );
  NOR2X0 U18623 ( .IN1(n10317), .IN2(n17663), .QN(WX10343) );
  NOR2X0 U18624 ( .IN1(n17664), .IN2(n17665), .QN(n17663) );
  INVX0 U18625 ( .INP(n17666), .ZN(n17665) );
  NAND2X0 U18626 ( .IN1(n9837), .IN2(DFF_1517_n1), .QN(n17666) );
  NOR2X0 U18627 ( .IN1(DFF_1517_n1), .IN2(n9837), .QN(n17664) );
  NOR2X0 U18628 ( .IN1(n10318), .IN2(n17667), .QN(WX10341) );
  NAND2X0 U18629 ( .IN1(n17668), .IN2(n17669), .QN(n17667) );
  INVX0 U18630 ( .INP(n17670), .ZN(n17669) );
  NOR2X0 U18631 ( .IN1(WX9924), .IN2(DFF_1516_n1), .QN(n17670) );
  NAND2X0 U18632 ( .IN1(DFF_1516_n1), .IN2(WX9924), .QN(n17668) );
  NOR2X0 U18633 ( .IN1(n10318), .IN2(n17671), .QN(WX10339) );
  NAND2X0 U18634 ( .IN1(n17672), .IN2(n17673), .QN(n17671) );
  INVX0 U18635 ( .INP(n17674), .ZN(n17673) );
  NOR2X0 U18636 ( .IN1(WX9926), .IN2(DFF_1515_n1), .QN(n17674) );
  NAND2X0 U18637 ( .IN1(DFF_1515_n1), .IN2(WX9926), .QN(n17672) );
  NOR2X0 U18638 ( .IN1(n10318), .IN2(n17675), .QN(WX10337) );
  NOR2X0 U18639 ( .IN1(n17676), .IN2(n17677), .QN(n17675) );
  INVX0 U18640 ( .INP(n17678), .ZN(n17677) );
  NAND2X0 U18641 ( .IN1(CRC_OUT_2_10), .IN2(n17679), .QN(n17678) );
  NOR2X0 U18642 ( .IN1(n17679), .IN2(CRC_OUT_2_10), .QN(n17676) );
  NAND2X0 U18643 ( .IN1(n17680), .IN2(n17681), .QN(n17679) );
  NAND2X0 U18644 ( .IN1(n9500), .IN2(CRC_OUT_2_31), .QN(n17681) );
  NAND2X0 U18645 ( .IN1(DFF_1535_n1), .IN2(WX9928), .QN(n17680) );
  NOR2X0 U18646 ( .IN1(n10318), .IN2(n17682), .QN(WX10335) );
  NAND2X0 U18647 ( .IN1(n17683), .IN2(n17684), .QN(n17682) );
  INVX0 U18648 ( .INP(n17685), .ZN(n17684) );
  NOR2X0 U18649 ( .IN1(WX9930), .IN2(DFF_1513_n1), .QN(n17685) );
  NAND2X0 U18650 ( .IN1(DFF_1513_n1), .IN2(WX9930), .QN(n17683) );
  NOR2X0 U18651 ( .IN1(n10318), .IN2(n17686), .QN(WX10333) );
  NAND2X0 U18652 ( .IN1(n17687), .IN2(n17688), .QN(n17686) );
  INVX0 U18653 ( .INP(n17689), .ZN(n17688) );
  NOR2X0 U18654 ( .IN1(WX9932), .IN2(DFF_1512_n1), .QN(n17689) );
  NAND2X0 U18655 ( .IN1(DFF_1512_n1), .IN2(WX9932), .QN(n17687) );
  NOR2X0 U18656 ( .IN1(n10318), .IN2(n17690), .QN(WX10331) );
  NAND2X0 U18657 ( .IN1(n17691), .IN2(n17692), .QN(n17690) );
  INVX0 U18658 ( .INP(n17693), .ZN(n17692) );
  NOR2X0 U18659 ( .IN1(WX9934), .IN2(DFF_1511_n1), .QN(n17693) );
  NAND2X0 U18660 ( .IN1(DFF_1511_n1), .IN2(WX9934), .QN(n17691) );
  NOR2X0 U18661 ( .IN1(n10318), .IN2(n17694), .QN(WX10329) );
  NAND2X0 U18662 ( .IN1(n17695), .IN2(n17696), .QN(n17694) );
  INVX0 U18663 ( .INP(n17697), .ZN(n17696) );
  NOR2X0 U18664 ( .IN1(WX9936), .IN2(DFF_1510_n1), .QN(n17697) );
  NAND2X0 U18665 ( .IN1(DFF_1510_n1), .IN2(WX9936), .QN(n17695) );
  NOR2X0 U18666 ( .IN1(n10318), .IN2(n17698), .QN(WX10327) );
  NAND2X0 U18667 ( .IN1(n17699), .IN2(n17700), .QN(n17698) );
  INVX0 U18668 ( .INP(n17701), .ZN(n17700) );
  NOR2X0 U18669 ( .IN1(WX9938), .IN2(DFF_1509_n1), .QN(n17701) );
  NAND2X0 U18670 ( .IN1(DFF_1509_n1), .IN2(WX9938), .QN(n17699) );
  NOR2X0 U18671 ( .IN1(n10318), .IN2(n17702), .QN(WX10325) );
  NAND2X0 U18672 ( .IN1(n17703), .IN2(n17704), .QN(n17702) );
  INVX0 U18673 ( .INP(n17705), .ZN(n17704) );
  NOR2X0 U18674 ( .IN1(WX9940), .IN2(DFF_1508_n1), .QN(n17705) );
  NAND2X0 U18675 ( .IN1(DFF_1508_n1), .IN2(WX9940), .QN(n17703) );
  NOR2X0 U18676 ( .IN1(n10318), .IN2(n17706), .QN(WX10323) );
  NOR2X0 U18677 ( .IN1(n17707), .IN2(n17708), .QN(n17706) );
  INVX0 U18678 ( .INP(n17709), .ZN(n17708) );
  NAND2X0 U18679 ( .IN1(CRC_OUT_2_3), .IN2(n17710), .QN(n17709) );
  NOR2X0 U18680 ( .IN1(n17710), .IN2(CRC_OUT_2_3), .QN(n17707) );
  NAND2X0 U18681 ( .IN1(n17711), .IN2(n17712), .QN(n17710) );
  NAND2X0 U18682 ( .IN1(n9501), .IN2(CRC_OUT_2_31), .QN(n17712) );
  NAND2X0 U18683 ( .IN1(DFF_1535_n1), .IN2(WX9942), .QN(n17711) );
  NOR2X0 U18684 ( .IN1(n10318), .IN2(n17713), .QN(WX10321) );
  NOR2X0 U18685 ( .IN1(n17714), .IN2(n17715), .QN(n17713) );
  NOR2X0 U18686 ( .IN1(test_so87), .IN2(WX9944), .QN(n17715) );
  NOR2X0 U18687 ( .IN1(n9574), .IN2(n9864), .QN(n17714) );
  NOR2X0 U18688 ( .IN1(n10318), .IN2(n17716), .QN(WX10319) );
  NAND2X0 U18689 ( .IN1(n17717), .IN2(n17718), .QN(n17716) );
  INVX0 U18690 ( .INP(n17719), .ZN(n17718) );
  NOR2X0 U18691 ( .IN1(WX9946), .IN2(DFF_1505_n1), .QN(n17719) );
  NAND2X0 U18692 ( .IN1(DFF_1505_n1), .IN2(WX9946), .QN(n17717) );
  NOR2X0 U18693 ( .IN1(n10318), .IN2(n17720), .QN(WX10317) );
  NAND2X0 U18694 ( .IN1(n17721), .IN2(n17722), .QN(n17720) );
  INVX0 U18695 ( .INP(n17723), .ZN(n17722) );
  NOR2X0 U18696 ( .IN1(WX9948), .IN2(DFF_1504_n1), .QN(n17723) );
  NAND2X0 U18697 ( .IN1(DFF_1504_n1), .IN2(WX9948), .QN(n17721) );
  NOR2X0 U18698 ( .IN1(n10319), .IN2(n17724), .QN(WX10315) );
  NAND2X0 U18699 ( .IN1(n17725), .IN2(n17726), .QN(n17724) );
  NAND2X0 U18700 ( .IN1(n9518), .IN2(CRC_OUT_2_31), .QN(n17726) );
  NAND2X0 U18701 ( .IN1(DFF_1535_n1), .IN2(WX9950), .QN(n17725) );
  NAND2X0 U18702 ( .IN1(n17727), .IN2(n17728), .QN(DATA_9_9) );
  INVX0 U18703 ( .INP(n17729), .ZN(n17728) );
  NOR2X0 U18704 ( .IN1(n17730), .IN2(n11269), .QN(n17729) );
  NAND2X0 U18705 ( .IN1(n11269), .IN2(n17730), .QN(n17727) );
  NAND2X0 U18706 ( .IN1(TM0), .IN2(WX529), .QN(n17730) );
  NAND2X0 U18707 ( .IN1(n17731), .IN2(n17732), .QN(n11269) );
  NAND2X0 U18708 ( .IN1(n17733), .IN2(n17734), .QN(n17732) );
  INVX0 U18709 ( .INP(n17735), .ZN(n17731) );
  NOR2X0 U18710 ( .IN1(n17734), .IN2(n17733), .QN(n17735) );
  NAND2X0 U18711 ( .IN1(n17736), .IN2(n17737), .QN(n17733) );
  NAND2X0 U18712 ( .IN1(n9779), .IN2(n17738), .QN(n17737) );
  INVX0 U18713 ( .INP(n17739), .ZN(n17736) );
  NOR2X0 U18714 ( .IN1(n17738), .IN2(n9779), .QN(n17739) );
  NOR2X0 U18715 ( .IN1(n17740), .IN2(n17741), .QN(n17738) );
  NOR2X0 U18716 ( .IN1(WX881), .IN2(n9780), .QN(n17741) );
  INVX0 U18717 ( .INP(n17742), .ZN(n17740) );
  NAND2X0 U18718 ( .IN1(n9780), .IN2(WX881), .QN(n17742) );
  NOR2X0 U18719 ( .IN1(n17743), .IN2(n17744), .QN(n17734) );
  INVX0 U18720 ( .INP(n17745), .ZN(n17744) );
  NAND2X0 U18721 ( .IN1(n3485), .IN2(n2340), .QN(n17745) );
  NOR2X0 U18722 ( .IN1(n2340), .IN2(n3485), .QN(n17743) );
  NAND2X0 U18723 ( .IN1(n17746), .IN2(n17747), .QN(DATA_9_8) );
  INVX0 U18724 ( .INP(n17748), .ZN(n17747) );
  NOR2X0 U18725 ( .IN1(n17749), .IN2(n11259), .QN(n17748) );
  NAND2X0 U18726 ( .IN1(n11259), .IN2(n17749), .QN(n17746) );
  NAND2X0 U18727 ( .IN1(TM0), .IN2(WX531), .QN(n17749) );
  NAND2X0 U18728 ( .IN1(n17750), .IN2(n17751), .QN(n11259) );
  NAND2X0 U18729 ( .IN1(n17752), .IN2(n17753), .QN(n17751) );
  INVX0 U18730 ( .INP(n17754), .ZN(n17750) );
  NOR2X0 U18731 ( .IN1(n17753), .IN2(n17752), .QN(n17754) );
  NAND2X0 U18732 ( .IN1(n17755), .IN2(n17756), .QN(n17752) );
  NAND2X0 U18733 ( .IN1(n9789), .IN2(n17757), .QN(n17756) );
  INVX0 U18734 ( .INP(n17758), .ZN(n17755) );
  NOR2X0 U18735 ( .IN1(n17757), .IN2(n9789), .QN(n17758) );
  NOR2X0 U18736 ( .IN1(n17759), .IN2(n17760), .QN(n17757) );
  INVX0 U18737 ( .INP(n17761), .ZN(n17760) );
  NAND2X0 U18738 ( .IN1(n9791), .IN2(WX883), .QN(n17761) );
  NOR2X0 U18739 ( .IN1(WX883), .IN2(n9791), .QN(n17759) );
  NOR2X0 U18740 ( .IN1(n17762), .IN2(n17763), .QN(n17753) );
  INVX0 U18741 ( .INP(n17764), .ZN(n17763) );
  NAND2X0 U18742 ( .IN1(n3483), .IN2(n2340), .QN(n17764) );
  NOR2X0 U18743 ( .IN1(n2340), .IN2(n3483), .QN(n17762) );
  NAND2X0 U18744 ( .IN1(n17765), .IN2(n17766), .QN(DATA_9_7) );
  INVX0 U18745 ( .INP(n17767), .ZN(n17766) );
  NOR2X0 U18746 ( .IN1(n17768), .IN2(n11249), .QN(n17767) );
  NAND2X0 U18747 ( .IN1(n11249), .IN2(n17768), .QN(n17765) );
  NAND2X0 U18748 ( .IN1(TM0), .IN2(WX533), .QN(n17768) );
  NAND2X0 U18749 ( .IN1(n17769), .IN2(n17770), .QN(n11249) );
  NAND2X0 U18750 ( .IN1(n17771), .IN2(n17772), .QN(n17770) );
  INVX0 U18751 ( .INP(n17773), .ZN(n17769) );
  NOR2X0 U18752 ( .IN1(n17772), .IN2(n17771), .QN(n17773) );
  NAND2X0 U18753 ( .IN1(n17774), .IN2(n17775), .QN(n17771) );
  NAND2X0 U18754 ( .IN1(n9819), .IN2(n17776), .QN(n17775) );
  INVX0 U18755 ( .INP(n17777), .ZN(n17774) );
  NOR2X0 U18756 ( .IN1(n17776), .IN2(n9819), .QN(n17777) );
  NOR2X0 U18757 ( .IN1(n17778), .IN2(n17779), .QN(n17776) );
  NOR2X0 U18758 ( .IN1(WX885), .IN2(n9820), .QN(n17779) );
  INVX0 U18759 ( .INP(n17780), .ZN(n17778) );
  NAND2X0 U18760 ( .IN1(n9820), .IN2(WX885), .QN(n17780) );
  NOR2X0 U18761 ( .IN1(n17781), .IN2(n17782), .QN(n17772) );
  INVX0 U18762 ( .INP(n17783), .ZN(n17782) );
  NAND2X0 U18763 ( .IN1(n3481), .IN2(n2340), .QN(n17783) );
  NOR2X0 U18764 ( .IN1(n2340), .IN2(n3481), .QN(n17781) );
  NOR2X0 U18765 ( .IN1(n17784), .IN2(n17785), .QN(DATA_9_6) );
  INVX0 U18766 ( .INP(n17786), .ZN(n17785) );
  NAND2X0 U18767 ( .IN1(n17787), .IN2(n11239), .QN(n17786) );
  NOR2X0 U18768 ( .IN1(n11239), .IN2(n17787), .QN(n17784) );
  NAND2X0 U18769 ( .IN1(TM0), .IN2(WX535), .QN(n17787) );
  NAND2X0 U18770 ( .IN1(n17788), .IN2(n17789), .QN(n11239) );
  NAND2X0 U18771 ( .IN1(n17790), .IN2(n17791), .QN(n17789) );
  NAND2X0 U18772 ( .IN1(n17792), .IN2(n17793), .QN(n17790) );
  NAND2X0 U18773 ( .IN1(n3479), .IN2(n2340), .QN(n17793) );
  NAND2X0 U18774 ( .IN1(TM0), .IN2(WX695), .QN(n17792) );
  NAND2X0 U18775 ( .IN1(n17794), .IN2(n17795), .QN(n17788) );
  NOR2X0 U18776 ( .IN1(n17796), .IN2(n17797), .QN(n17795) );
  NOR2X0 U18777 ( .IN1(n3479), .IN2(n2340), .QN(n17797) );
  NOR2X0 U18778 ( .IN1(TM0), .IN2(WX695), .QN(n17796) );
  INVX0 U18779 ( .INP(n17791), .ZN(n17794) );
  NOR2X0 U18780 ( .IN1(n17798), .IN2(n17799), .QN(n17791) );
  INVX0 U18781 ( .INP(n17800), .ZN(n17799) );
  NAND2X0 U18782 ( .IN1(n9807), .IN2(n17801), .QN(n17800) );
  NOR2X0 U18783 ( .IN1(n17801), .IN2(n9807), .QN(n17798) );
  NOR2X0 U18784 ( .IN1(n17802), .IN2(n17803), .QN(n17801) );
  INVX0 U18785 ( .INP(n17804), .ZN(n17803) );
  NAND2X0 U18786 ( .IN1(test_so5), .IN2(WX887), .QN(n17804) );
  NOR2X0 U18787 ( .IN1(WX887), .IN2(test_so5), .QN(n17802) );
  NAND2X0 U18788 ( .IN1(n17805), .IN2(n17806), .QN(DATA_9_5) );
  INVX0 U18789 ( .INP(n17807), .ZN(n17806) );
  NOR2X0 U18790 ( .IN1(n17808), .IN2(n11228), .QN(n17807) );
  NAND2X0 U18791 ( .IN1(n11228), .IN2(n17808), .QN(n17805) );
  NAND2X0 U18792 ( .IN1(TM0), .IN2(WX537), .QN(n17808) );
  NAND2X0 U18793 ( .IN1(n17809), .IN2(n17810), .QN(n11228) );
  NAND2X0 U18794 ( .IN1(n17811), .IN2(n17812), .QN(n17810) );
  INVX0 U18795 ( .INP(n17813), .ZN(n17809) );
  NOR2X0 U18796 ( .IN1(n17812), .IN2(n17811), .QN(n17813) );
  NAND2X0 U18797 ( .IN1(n17814), .IN2(n17815), .QN(n17811) );
  NAND2X0 U18798 ( .IN1(n9792), .IN2(n17816), .QN(n17815) );
  INVX0 U18799 ( .INP(n17817), .ZN(n17814) );
  NOR2X0 U18800 ( .IN1(n17816), .IN2(n9792), .QN(n17817) );
  NOR2X0 U18801 ( .IN1(n17818), .IN2(n17819), .QN(n17816) );
  INVX0 U18802 ( .INP(n17820), .ZN(n17819) );
  NAND2X0 U18803 ( .IN1(n9794), .IN2(WX889), .QN(n17820) );
  NOR2X0 U18804 ( .IN1(WX889), .IN2(n9794), .QN(n17818) );
  NOR2X0 U18805 ( .IN1(n17821), .IN2(n17822), .QN(n17812) );
  INVX0 U18806 ( .INP(n17823), .ZN(n17822) );
  NAND2X0 U18807 ( .IN1(n3477), .IN2(n2340), .QN(n17823) );
  NOR2X0 U18808 ( .IN1(n2340), .IN2(n3477), .QN(n17821) );
  NAND2X0 U18809 ( .IN1(n17824), .IN2(n17825), .QN(DATA_9_4) );
  INVX0 U18810 ( .INP(n17826), .ZN(n17825) );
  NOR2X0 U18811 ( .IN1(n17827), .IN2(n11219), .QN(n17826) );
  NAND2X0 U18812 ( .IN1(n11219), .IN2(n17827), .QN(n17824) );
  NAND2X0 U18813 ( .IN1(TM0), .IN2(WX539), .QN(n17827) );
  NAND2X0 U18814 ( .IN1(n17828), .IN2(n17829), .QN(n11219) );
  NAND2X0 U18815 ( .IN1(n17830), .IN2(n17831), .QN(n17829) );
  INVX0 U18816 ( .INP(n17832), .ZN(n17828) );
  NOR2X0 U18817 ( .IN1(n17831), .IN2(n17830), .QN(n17832) );
  NAND2X0 U18818 ( .IN1(n17833), .IN2(n17834), .QN(n17830) );
  NAND2X0 U18819 ( .IN1(n9795), .IN2(n17835), .QN(n17834) );
  INVX0 U18820 ( .INP(n17836), .ZN(n17833) );
  NOR2X0 U18821 ( .IN1(n17835), .IN2(n9795), .QN(n17836) );
  NOR2X0 U18822 ( .IN1(n17837), .IN2(n17838), .QN(n17835) );
  INVX0 U18823 ( .INP(n17839), .ZN(n17838) );
  NAND2X0 U18824 ( .IN1(n9797), .IN2(WX891), .QN(n17839) );
  NOR2X0 U18825 ( .IN1(WX891), .IN2(n9797), .QN(n17837) );
  NOR2X0 U18826 ( .IN1(n17840), .IN2(n17841), .QN(n17831) );
  INVX0 U18827 ( .INP(n17842), .ZN(n17841) );
  NAND2X0 U18828 ( .IN1(n3475), .IN2(n2340), .QN(n17842) );
  NOR2X0 U18829 ( .IN1(n2340), .IN2(n3475), .QN(n17840) );
  NAND2X0 U18830 ( .IN1(n17843), .IN2(n17844), .QN(DATA_9_31) );
  NAND2X0 U18831 ( .IN1(n17845), .IN2(n13781), .QN(n17844) );
  INVX0 U18832 ( .INP(n17846), .ZN(n13781) );
  INVX0 U18833 ( .INP(n17847), .ZN(n17845) );
  NAND2X0 U18834 ( .IN1(n17846), .IN2(n17847), .QN(n17843) );
  NAND2X0 U18835 ( .IN1(TM0), .IN2(WX485), .QN(n17847) );
  NAND2X0 U18836 ( .IN1(n17848), .IN2(n17849), .QN(n17846) );
  NAND2X0 U18837 ( .IN1(n17850), .IN2(n17851), .QN(n17849) );
  NAND2X0 U18838 ( .IN1(n17852), .IN2(n17853), .QN(n17850) );
  NAND2X0 U18839 ( .IN1(n3529), .IN2(n10014), .QN(n17853) );
  NAND2X0 U18840 ( .IN1(TM1), .IN2(WX645), .QN(n17852) );
  NAND2X0 U18841 ( .IN1(n17854), .IN2(n17855), .QN(n17848) );
  NOR2X0 U18842 ( .IN1(n17856), .IN2(n17857), .QN(n17855) );
  NOR2X0 U18843 ( .IN1(n3529), .IN2(n10003), .QN(n17857) );
  NOR2X0 U18844 ( .IN1(TM1), .IN2(WX645), .QN(n17856) );
  INVX0 U18845 ( .INP(n17851), .ZN(n17854) );
  NOR2X0 U18846 ( .IN1(n17858), .IN2(n17859), .QN(n17851) );
  INVX0 U18847 ( .INP(n17860), .ZN(n17859) );
  NAND2X0 U18848 ( .IN1(n9811), .IN2(n17861), .QN(n17860) );
  NOR2X0 U18849 ( .IN1(n17861), .IN2(n9811), .QN(n17858) );
  NOR2X0 U18850 ( .IN1(n17862), .IN2(n17863), .QN(n17861) );
  NOR2X0 U18851 ( .IN1(WX837), .IN2(n9812), .QN(n17863) );
  INVX0 U18852 ( .INP(n17864), .ZN(n17862) );
  NAND2X0 U18853 ( .IN1(n9812), .IN2(WX837), .QN(n17864) );
  NAND2X0 U18854 ( .IN1(n17865), .IN2(n17866), .QN(DATA_9_30) );
  INVX0 U18855 ( .INP(n17867), .ZN(n17866) );
  NOR2X0 U18856 ( .IN1(n17868), .IN2(n10765), .QN(n17867) );
  NAND2X0 U18857 ( .IN1(n10765), .IN2(n17868), .QN(n17865) );
  NAND2X0 U18858 ( .IN1(TM0), .IN2(WX487), .QN(n17868) );
  NAND2X0 U18859 ( .IN1(n17869), .IN2(n17870), .QN(n10765) );
  NAND2X0 U18860 ( .IN1(n17871), .IN2(n17872), .QN(n17870) );
  INVX0 U18861 ( .INP(n17873), .ZN(n17869) );
  NOR2X0 U18862 ( .IN1(n17872), .IN2(n17871), .QN(n17873) );
  NAND2X0 U18863 ( .IN1(n17874), .IN2(n17875), .QN(n17871) );
  NAND2X0 U18864 ( .IN1(n9737), .IN2(n17876), .QN(n17875) );
  INVX0 U18865 ( .INP(n17877), .ZN(n17874) );
  NOR2X0 U18866 ( .IN1(n17876), .IN2(n9737), .QN(n17877) );
  NOR2X0 U18867 ( .IN1(n17878), .IN2(n17879), .QN(n17876) );
  NOR2X0 U18868 ( .IN1(WX839), .IN2(n9738), .QN(n17879) );
  INVX0 U18869 ( .INP(n17880), .ZN(n17878) );
  NAND2X0 U18870 ( .IN1(n9738), .IN2(WX839), .QN(n17880) );
  NOR2X0 U18871 ( .IN1(n17881), .IN2(n17882), .QN(n17872) );
  INVX0 U18872 ( .INP(n17883), .ZN(n17882) );
  NAND2X0 U18873 ( .IN1(n3527), .IN2(n10014), .QN(n17883) );
  NOR2X0 U18874 ( .IN1(n10012), .IN2(n3527), .QN(n17881) );
  NAND2X0 U18875 ( .IN1(n17884), .IN2(n17885), .QN(DATA_9_3) );
  INVX0 U18876 ( .INP(n17886), .ZN(n17885) );
  NOR2X0 U18877 ( .IN1(n17887), .IN2(n11209), .QN(n17886) );
  NAND2X0 U18878 ( .IN1(n11209), .IN2(n17887), .QN(n17884) );
  NAND2X0 U18879 ( .IN1(TM0), .IN2(WX541), .QN(n17887) );
  NAND2X0 U18880 ( .IN1(n17888), .IN2(n17889), .QN(n11209) );
  NAND2X0 U18881 ( .IN1(n17890), .IN2(n17891), .QN(n17889) );
  INVX0 U18882 ( .INP(n17892), .ZN(n17888) );
  NOR2X0 U18883 ( .IN1(n17891), .IN2(n17890), .QN(n17892) );
  NAND2X0 U18884 ( .IN1(n17893), .IN2(n17894), .QN(n17890) );
  NAND2X0 U18885 ( .IN1(n9740), .IN2(n17895), .QN(n17894) );
  INVX0 U18886 ( .INP(n17896), .ZN(n17893) );
  NOR2X0 U18887 ( .IN1(n17895), .IN2(n9740), .QN(n17896) );
  NOR2X0 U18888 ( .IN1(n17897), .IN2(n17898), .QN(n17895) );
  INVX0 U18889 ( .INP(n17899), .ZN(n17898) );
  NAND2X0 U18890 ( .IN1(n9742), .IN2(WX893), .QN(n17899) );
  NOR2X0 U18891 ( .IN1(WX893), .IN2(n9742), .QN(n17897) );
  NOR2X0 U18892 ( .IN1(n17900), .IN2(n17901), .QN(n17891) );
  INVX0 U18893 ( .INP(n17902), .ZN(n17901) );
  NAND2X0 U18894 ( .IN1(n3473), .IN2(n2340), .QN(n17902) );
  NOR2X0 U18895 ( .IN1(n2340), .IN2(n3473), .QN(n17900) );
  NAND2X0 U18896 ( .IN1(n17903), .IN2(n17904), .QN(DATA_9_29) );
  INVX0 U18897 ( .INP(n17905), .ZN(n17904) );
  NOR2X0 U18898 ( .IN1(n17906), .IN2(n10755), .QN(n17905) );
  NAND2X0 U18899 ( .IN1(n10755), .IN2(n17906), .QN(n17903) );
  NAND2X0 U18900 ( .IN1(TM0), .IN2(WX489), .QN(n17906) );
  NAND2X0 U18901 ( .IN1(n17907), .IN2(n17908), .QN(n10755) );
  NAND2X0 U18902 ( .IN1(n17909), .IN2(n17910), .QN(n17908) );
  INVX0 U18903 ( .INP(n17911), .ZN(n17907) );
  NOR2X0 U18904 ( .IN1(n17910), .IN2(n17909), .QN(n17911) );
  NAND2X0 U18905 ( .IN1(n17912), .IN2(n17913), .QN(n17909) );
  NAND2X0 U18906 ( .IN1(n9746), .IN2(n17914), .QN(n17913) );
  INVX0 U18907 ( .INP(n17915), .ZN(n17912) );
  NOR2X0 U18908 ( .IN1(n17914), .IN2(n9746), .QN(n17915) );
  NOR2X0 U18909 ( .IN1(n17916), .IN2(n17917), .QN(n17914) );
  INVX0 U18910 ( .INP(n17918), .ZN(n17917) );
  NAND2X0 U18911 ( .IN1(n9748), .IN2(WX841), .QN(n17918) );
  NOR2X0 U18912 ( .IN1(WX841), .IN2(n9748), .QN(n17916) );
  NOR2X0 U18913 ( .IN1(n17919), .IN2(n17920), .QN(n17910) );
  INVX0 U18914 ( .INP(n17921), .ZN(n17920) );
  NAND2X0 U18915 ( .IN1(n3525), .IN2(n10015), .QN(n17921) );
  NOR2X0 U18916 ( .IN1(n10013), .IN2(n3525), .QN(n17919) );
  NOR2X0 U18917 ( .IN1(n17922), .IN2(n17923), .QN(DATA_9_28) );
  INVX0 U18918 ( .INP(n17924), .ZN(n17923) );
  NAND2X0 U18919 ( .IN1(n17925), .IN2(n10746), .QN(n17924) );
  NOR2X0 U18920 ( .IN1(n10746), .IN2(n17925), .QN(n17922) );
  NAND2X0 U18921 ( .IN1(TM0), .IN2(WX491), .QN(n17925) );
  NAND2X0 U18922 ( .IN1(n17926), .IN2(n17927), .QN(n10746) );
  NAND2X0 U18923 ( .IN1(n17928), .IN2(n17929), .QN(n17927) );
  NAND2X0 U18924 ( .IN1(n17930), .IN2(n17931), .QN(n17928) );
  NAND2X0 U18925 ( .IN1(n9757), .IN2(n10015), .QN(n17931) );
  NAND2X0 U18926 ( .IN1(TM1), .IN2(WX715), .QN(n17930) );
  NAND2X0 U18927 ( .IN1(n17932), .IN2(n17933), .QN(n17926) );
  NOR2X0 U18928 ( .IN1(n17934), .IN2(n17935), .QN(n17933) );
  NOR2X0 U18929 ( .IN1(n9757), .IN2(n10003), .QN(n17935) );
  NOR2X0 U18930 ( .IN1(TM1), .IN2(WX715), .QN(n17934) );
  INVX0 U18931 ( .INP(n17929), .ZN(n17932) );
  NOR2X0 U18932 ( .IN1(n17936), .IN2(n17937), .QN(n17929) );
  INVX0 U18933 ( .INP(n17938), .ZN(n17937) );
  NAND2X0 U18934 ( .IN1(n9755), .IN2(n17939), .QN(n17938) );
  NOR2X0 U18935 ( .IN1(n17939), .IN2(n9755), .QN(n17936) );
  NOR2X0 U18936 ( .IN1(n17940), .IN2(n17941), .QN(n17939) );
  INVX0 U18937 ( .INP(n17942), .ZN(n17941) );
  NAND2X0 U18938 ( .IN1(test_so2), .IN2(WX843), .QN(n17942) );
  NOR2X0 U18939 ( .IN1(WX843), .IN2(test_so2), .QN(n17940) );
  NAND2X0 U18940 ( .IN1(n17943), .IN2(n17944), .QN(DATA_9_27) );
  INVX0 U18941 ( .INP(n17945), .ZN(n17944) );
  NOR2X0 U18942 ( .IN1(n17946), .IN2(n10735), .QN(n17945) );
  NAND2X0 U18943 ( .IN1(n10735), .IN2(n17946), .QN(n17943) );
  NAND2X0 U18944 ( .IN1(TM0), .IN2(WX493), .QN(n17946) );
  NAND2X0 U18945 ( .IN1(n17947), .IN2(n17948), .QN(n10735) );
  NAND2X0 U18946 ( .IN1(n17949), .IN2(n17950), .QN(n17948) );
  INVX0 U18947 ( .INP(n17951), .ZN(n17947) );
  NOR2X0 U18948 ( .IN1(n17950), .IN2(n17949), .QN(n17951) );
  NAND2X0 U18949 ( .IN1(n17952), .IN2(n17953), .QN(n17949) );
  NAND2X0 U18950 ( .IN1(n9761), .IN2(n17954), .QN(n17953) );
  INVX0 U18951 ( .INP(n17955), .ZN(n17952) );
  NOR2X0 U18952 ( .IN1(n17954), .IN2(n9761), .QN(n17955) );
  NOR2X0 U18953 ( .IN1(n17956), .IN2(n17957), .QN(n17954) );
  INVX0 U18954 ( .INP(n17958), .ZN(n17957) );
  NAND2X0 U18955 ( .IN1(n9763), .IN2(WX845), .QN(n17958) );
  NOR2X0 U18956 ( .IN1(WX845), .IN2(n9763), .QN(n17956) );
  NOR2X0 U18957 ( .IN1(n17959), .IN2(n17960), .QN(n17950) );
  INVX0 U18958 ( .INP(n17961), .ZN(n17960) );
  NAND2X0 U18959 ( .IN1(n3521), .IN2(n10015), .QN(n17961) );
  NOR2X0 U18960 ( .IN1(n10012), .IN2(n3521), .QN(n17959) );
  NAND2X0 U18961 ( .IN1(n17962), .IN2(n17963), .QN(DATA_9_26) );
  INVX0 U18962 ( .INP(n17964), .ZN(n17963) );
  NOR2X0 U18963 ( .IN1(n17965), .IN2(n10725), .QN(n17964) );
  NAND2X0 U18964 ( .IN1(n10725), .IN2(n17965), .QN(n17962) );
  NAND2X0 U18965 ( .IN1(TM0), .IN2(WX495), .QN(n17965) );
  NAND2X0 U18966 ( .IN1(n17966), .IN2(n17967), .QN(n10725) );
  NAND2X0 U18967 ( .IN1(n17968), .IN2(n17969), .QN(n17967) );
  INVX0 U18968 ( .INP(n17970), .ZN(n17966) );
  NOR2X0 U18969 ( .IN1(n17969), .IN2(n17968), .QN(n17970) );
  NAND2X0 U18970 ( .IN1(n17971), .IN2(n17972), .QN(n17968) );
  NAND2X0 U18971 ( .IN1(n9764), .IN2(n17973), .QN(n17972) );
  INVX0 U18972 ( .INP(n17974), .ZN(n17971) );
  NOR2X0 U18973 ( .IN1(n17973), .IN2(n9764), .QN(n17974) );
  NOR2X0 U18974 ( .IN1(n17975), .IN2(n17976), .QN(n17973) );
  INVX0 U18975 ( .INP(n17977), .ZN(n17976) );
  NAND2X0 U18976 ( .IN1(n9766), .IN2(WX847), .QN(n17977) );
  NOR2X0 U18977 ( .IN1(WX847), .IN2(n9766), .QN(n17975) );
  NOR2X0 U18978 ( .IN1(n17978), .IN2(n17979), .QN(n17969) );
  INVX0 U18979 ( .INP(n17980), .ZN(n17979) );
  NAND2X0 U18980 ( .IN1(n3519), .IN2(n10015), .QN(n17980) );
  NOR2X0 U18981 ( .IN1(n10013), .IN2(n3519), .QN(n17978) );
  NAND2X0 U18982 ( .IN1(n17981), .IN2(n17982), .QN(DATA_9_25) );
  INVX0 U18983 ( .INP(n17983), .ZN(n17982) );
  NOR2X0 U18984 ( .IN1(n17984), .IN2(n10693), .QN(n17983) );
  NAND2X0 U18985 ( .IN1(n10693), .IN2(n17984), .QN(n17981) );
  NAND2X0 U18986 ( .IN1(TM0), .IN2(WX497), .QN(n17984) );
  NAND2X0 U18987 ( .IN1(n17985), .IN2(n17986), .QN(n10693) );
  NAND2X0 U18988 ( .IN1(n17987), .IN2(n17988), .QN(n17986) );
  INVX0 U18989 ( .INP(n17989), .ZN(n17985) );
  NOR2X0 U18990 ( .IN1(n17988), .IN2(n17987), .QN(n17989) );
  NAND2X0 U18991 ( .IN1(n17990), .IN2(n17991), .QN(n17987) );
  NAND2X0 U18992 ( .IN1(n9773), .IN2(n17992), .QN(n17991) );
  INVX0 U18993 ( .INP(n17993), .ZN(n17990) );
  NOR2X0 U18994 ( .IN1(n17992), .IN2(n9773), .QN(n17993) );
  NOR2X0 U18995 ( .IN1(n17994), .IN2(n17995), .QN(n17992) );
  INVX0 U18996 ( .INP(n17996), .ZN(n17995) );
  NAND2X0 U18997 ( .IN1(n9775), .IN2(WX849), .QN(n17996) );
  NOR2X0 U18998 ( .IN1(WX849), .IN2(n9775), .QN(n17994) );
  NOR2X0 U18999 ( .IN1(n17997), .IN2(n17998), .QN(n17988) );
  INVX0 U19000 ( .INP(n17999), .ZN(n17998) );
  NAND2X0 U19001 ( .IN1(n3517), .IN2(n10015), .QN(n17999) );
  NOR2X0 U19002 ( .IN1(n10011), .IN2(n3517), .QN(n17997) );
  NOR2X0 U19003 ( .IN1(n18000), .IN2(n18001), .QN(DATA_9_24) );
  INVX0 U19004 ( .INP(n18002), .ZN(n18001) );
  NAND2X0 U19005 ( .IN1(n18003), .IN2(n10674), .QN(n18002) );
  NOR2X0 U19006 ( .IN1(n10674), .IN2(n18003), .QN(n18000) );
  NAND2X0 U19007 ( .IN1(TM0), .IN2(WX499), .QN(n18003) );
  NAND2X0 U19008 ( .IN1(n18004), .IN2(n18005), .QN(n10674) );
  NAND2X0 U19009 ( .IN1(n18006), .IN2(n18007), .QN(n18005) );
  NAND2X0 U19010 ( .IN1(n18008), .IN2(n18009), .QN(n18006) );
  NAND2X0 U19011 ( .IN1(n3515), .IN2(n10015), .QN(n18009) );
  NAND2X0 U19012 ( .IN1(TM1), .IN2(WX659), .QN(n18008) );
  NAND2X0 U19013 ( .IN1(n18010), .IN2(n18011), .QN(n18004) );
  NOR2X0 U19014 ( .IN1(n18012), .IN2(n18013), .QN(n18011) );
  NOR2X0 U19015 ( .IN1(n3515), .IN2(n10003), .QN(n18013) );
  NOR2X0 U19016 ( .IN1(TM1), .IN2(WX659), .QN(n18012) );
  INVX0 U19017 ( .INP(n18007), .ZN(n18010) );
  NOR2X0 U19018 ( .IN1(n18014), .IN2(n18015), .QN(n18007) );
  INVX0 U19019 ( .INP(n18016), .ZN(n18015) );
  NAND2X0 U19020 ( .IN1(n9782), .IN2(n18017), .QN(n18016) );
  NOR2X0 U19021 ( .IN1(n18017), .IN2(n9782), .QN(n18014) );
  NOR2X0 U19022 ( .IN1(n18018), .IN2(n18019), .QN(n18017) );
  INVX0 U19023 ( .INP(n18020), .ZN(n18019) );
  NAND2X0 U19024 ( .IN1(test_so4), .IN2(WX851), .QN(n18020) );
  NOR2X0 U19025 ( .IN1(WX851), .IN2(test_so4), .QN(n18018) );
  NAND2X0 U19026 ( .IN1(n18021), .IN2(n18022), .QN(DATA_9_23) );
  INVX0 U19027 ( .INP(n18023), .ZN(n18022) );
  NOR2X0 U19028 ( .IN1(n18024), .IN2(n10663), .QN(n18023) );
  NAND2X0 U19029 ( .IN1(n10663), .IN2(n18024), .QN(n18021) );
  NAND2X0 U19030 ( .IN1(TM0), .IN2(WX501), .QN(n18024) );
  NAND2X0 U19031 ( .IN1(n18025), .IN2(n18026), .QN(n10663) );
  NAND2X0 U19032 ( .IN1(n18027), .IN2(n18028), .QN(n18026) );
  INVX0 U19033 ( .INP(n18029), .ZN(n18025) );
  NOR2X0 U19034 ( .IN1(n18028), .IN2(n18027), .QN(n18029) );
  NAND2X0 U19035 ( .IN1(n18030), .IN2(n18031), .QN(n18027) );
  NAND2X0 U19036 ( .IN1(n9784), .IN2(n18032), .QN(n18031) );
  INVX0 U19037 ( .INP(n18033), .ZN(n18030) );
  NOR2X0 U19038 ( .IN1(n18032), .IN2(n9784), .QN(n18033) );
  NOR2X0 U19039 ( .IN1(n18034), .IN2(n18035), .QN(n18032) );
  INVX0 U19040 ( .INP(n18036), .ZN(n18035) );
  NAND2X0 U19041 ( .IN1(n9786), .IN2(WX853), .QN(n18036) );
  NOR2X0 U19042 ( .IN1(WX853), .IN2(n9786), .QN(n18034) );
  NOR2X0 U19043 ( .IN1(n18037), .IN2(n18038), .QN(n18028) );
  INVX0 U19044 ( .INP(n18039), .ZN(n18038) );
  NAND2X0 U19045 ( .IN1(n3513), .IN2(n10015), .QN(n18039) );
  NOR2X0 U19046 ( .IN1(n10012), .IN2(n3513), .QN(n18037) );
  NAND2X0 U19047 ( .IN1(n18040), .IN2(n18041), .QN(DATA_9_22) );
  INVX0 U19048 ( .INP(n18042), .ZN(n18041) );
  NOR2X0 U19049 ( .IN1(n18043), .IN2(n10654), .QN(n18042) );
  NAND2X0 U19050 ( .IN1(n10654), .IN2(n18043), .QN(n18040) );
  NAND2X0 U19051 ( .IN1(TM0), .IN2(WX503), .QN(n18043) );
  NAND2X0 U19052 ( .IN1(n18044), .IN2(n18045), .QN(n10654) );
  NAND2X0 U19053 ( .IN1(n18046), .IN2(n18047), .QN(n18045) );
  INVX0 U19054 ( .INP(n18048), .ZN(n18044) );
  NOR2X0 U19055 ( .IN1(n18047), .IN2(n18046), .QN(n18048) );
  NAND2X0 U19056 ( .IN1(n18049), .IN2(n18050), .QN(n18046) );
  NAND2X0 U19057 ( .IN1(n9798), .IN2(n18051), .QN(n18050) );
  INVX0 U19058 ( .INP(n18052), .ZN(n18049) );
  NOR2X0 U19059 ( .IN1(n18051), .IN2(n9798), .QN(n18052) );
  NOR2X0 U19060 ( .IN1(n18053), .IN2(n18054), .QN(n18051) );
  NOR2X0 U19061 ( .IN1(WX855), .IN2(n9799), .QN(n18054) );
  INVX0 U19062 ( .INP(n18055), .ZN(n18053) );
  NAND2X0 U19063 ( .IN1(n9799), .IN2(WX855), .QN(n18055) );
  NOR2X0 U19064 ( .IN1(n18056), .IN2(n18057), .QN(n18047) );
  INVX0 U19065 ( .INP(n18058), .ZN(n18057) );
  NAND2X0 U19066 ( .IN1(n3511), .IN2(n10016), .QN(n18058) );
  NOR2X0 U19067 ( .IN1(n10011), .IN2(n3511), .QN(n18056) );
  NAND2X0 U19068 ( .IN1(n18059), .IN2(n18060), .QN(DATA_9_21) );
  INVX0 U19069 ( .INP(n18061), .ZN(n18060) );
  NOR2X0 U19070 ( .IN1(n18062), .IN2(n10644), .QN(n18061) );
  NAND2X0 U19071 ( .IN1(n10644), .IN2(n18062), .QN(n18059) );
  NAND2X0 U19072 ( .IN1(TM0), .IN2(WX505), .QN(n18062) );
  NAND2X0 U19073 ( .IN1(n18063), .IN2(n18064), .QN(n10644) );
  NAND2X0 U19074 ( .IN1(n18065), .IN2(n18066), .QN(n18064) );
  INVX0 U19075 ( .INP(n18067), .ZN(n18063) );
  NOR2X0 U19076 ( .IN1(n18066), .IN2(n18065), .QN(n18067) );
  NAND2X0 U19077 ( .IN1(n18068), .IN2(n18069), .QN(n18065) );
  NAND2X0 U19078 ( .IN1(n9804), .IN2(n18070), .QN(n18069) );
  INVX0 U19079 ( .INP(n18071), .ZN(n18068) );
  NOR2X0 U19080 ( .IN1(n18070), .IN2(n9804), .QN(n18071) );
  NOR2X0 U19081 ( .IN1(n18072), .IN2(n18073), .QN(n18070) );
  NOR2X0 U19082 ( .IN1(WX857), .IN2(n9805), .QN(n18073) );
  INVX0 U19083 ( .INP(n18074), .ZN(n18072) );
  NAND2X0 U19084 ( .IN1(n9805), .IN2(WX857), .QN(n18074) );
  NOR2X0 U19085 ( .IN1(n18075), .IN2(n18076), .QN(n18066) );
  INVX0 U19086 ( .INP(n18077), .ZN(n18076) );
  NAND2X0 U19087 ( .IN1(n3509), .IN2(n10016), .QN(n18077) );
  NOR2X0 U19088 ( .IN1(n10011), .IN2(n3509), .QN(n18075) );
  NOR2X0 U19089 ( .IN1(n18078), .IN2(n18079), .QN(DATA_9_20) );
  INVX0 U19090 ( .INP(n18080), .ZN(n18079) );
  NAND2X0 U19091 ( .IN1(n18081), .IN2(n10634), .QN(n18080) );
  NOR2X0 U19092 ( .IN1(n10634), .IN2(n18081), .QN(n18078) );
  NAND2X0 U19093 ( .IN1(TM0), .IN2(WX507), .QN(n18081) );
  NAND2X0 U19094 ( .IN1(n18082), .IN2(n18083), .QN(n10634) );
  NAND2X0 U19095 ( .IN1(n18084), .IN2(n18085), .QN(n18083) );
  NAND2X0 U19096 ( .IN1(n18086), .IN2(n18087), .QN(n18084) );
  NAND2X0 U19097 ( .IN1(n3507), .IN2(n10016), .QN(n18087) );
  NAND2X0 U19098 ( .IN1(TM1), .IN2(WX667), .QN(n18086) );
  NAND2X0 U19099 ( .IN1(n18088), .IN2(n18089), .QN(n18082) );
  NOR2X0 U19100 ( .IN1(n18090), .IN2(n18091), .QN(n18089) );
  NOR2X0 U19101 ( .IN1(n3507), .IN2(n10003), .QN(n18091) );
  NOR2X0 U19102 ( .IN1(TM1), .IN2(WX667), .QN(n18090) );
  INVX0 U19103 ( .INP(n18085), .ZN(n18088) );
  NOR2X0 U19104 ( .IN1(n18092), .IN2(n18093), .QN(n18085) );
  INVX0 U19105 ( .INP(n18094), .ZN(n18093) );
  NAND2X0 U19106 ( .IN1(n9809), .IN2(n18095), .QN(n18094) );
  NOR2X0 U19107 ( .IN1(n18095), .IN2(n9809), .QN(n18092) );
  NOR2X0 U19108 ( .IN1(n18096), .IN2(n18097), .QN(n18095) );
  INVX0 U19109 ( .INP(n18098), .ZN(n18097) );
  NAND2X0 U19110 ( .IN1(test_so6), .IN2(WX731), .QN(n18098) );
  NOR2X0 U19111 ( .IN1(WX731), .IN2(test_so6), .QN(n18096) );
  NOR2X0 U19112 ( .IN1(n18099), .IN2(n18100), .QN(DATA_9_2) );
  INVX0 U19113 ( .INP(n18101), .ZN(n18100) );
  NAND2X0 U19114 ( .IN1(n18102), .IN2(n11199), .QN(n18101) );
  NOR2X0 U19115 ( .IN1(n11199), .IN2(n18102), .QN(n18099) );
  NAND2X0 U19116 ( .IN1(TM0), .IN2(WX543), .QN(n18102) );
  NAND2X0 U19117 ( .IN1(n18103), .IN2(n18104), .QN(n11199) );
  NAND2X0 U19118 ( .IN1(n18105), .IN2(n18106), .QN(n18104) );
  NAND2X0 U19119 ( .IN1(n18107), .IN2(n18108), .QN(n18105) );
  NAND2X0 U19120 ( .IN1(n3471), .IN2(n2340), .QN(n18108) );
  NAND2X0 U19121 ( .IN1(TM0), .IN2(WX703), .QN(n18107) );
  NAND2X0 U19122 ( .IN1(n18109), .IN2(n18110), .QN(n18103) );
  NOR2X0 U19123 ( .IN1(n18111), .IN2(n18112), .QN(n18110) );
  NOR2X0 U19124 ( .IN1(n3471), .IN2(n2340), .QN(n18112) );
  NOR2X0 U19125 ( .IN1(TM0), .IN2(WX703), .QN(n18111) );
  INVX0 U19126 ( .INP(n18106), .ZN(n18109) );
  NOR2X0 U19127 ( .IN1(n18113), .IN2(n18114), .QN(n18106) );
  INVX0 U19128 ( .INP(n18115), .ZN(n18114) );
  NAND2X0 U19129 ( .IN1(n9817), .IN2(n18116), .QN(n18115) );
  NOR2X0 U19130 ( .IN1(n18116), .IN2(n9817), .QN(n18113) );
  NOR2X0 U19131 ( .IN1(n18117), .IN2(n18118), .QN(n18116) );
  INVX0 U19132 ( .INP(n18119), .ZN(n18118) );
  NAND2X0 U19133 ( .IN1(test_so7), .IN2(WX895), .QN(n18119) );
  NOR2X0 U19134 ( .IN1(WX895), .IN2(test_so7), .QN(n18117) );
  NAND2X0 U19135 ( .IN1(n18120), .IN2(n18121), .QN(DATA_9_19) );
  INVX0 U19136 ( .INP(n18122), .ZN(n18121) );
  NOR2X0 U19137 ( .IN1(n18123), .IN2(n10623), .QN(n18122) );
  NAND2X0 U19138 ( .IN1(n10623), .IN2(n18123), .QN(n18120) );
  NAND2X0 U19139 ( .IN1(TM0), .IN2(WX509), .QN(n18123) );
  NAND2X0 U19140 ( .IN1(n18124), .IN2(n18125), .QN(n10623) );
  NAND2X0 U19141 ( .IN1(n18126), .IN2(n18127), .QN(n18125) );
  INVX0 U19142 ( .INP(n18128), .ZN(n18124) );
  NOR2X0 U19143 ( .IN1(n18127), .IN2(n18126), .QN(n18128) );
  NAND2X0 U19144 ( .IN1(n18129), .IN2(n18130), .QN(n18126) );
  NAND2X0 U19145 ( .IN1(n9743), .IN2(n18131), .QN(n18130) );
  INVX0 U19146 ( .INP(n18132), .ZN(n18129) );
  NOR2X0 U19147 ( .IN1(n18131), .IN2(n9743), .QN(n18132) );
  NOR2X0 U19148 ( .IN1(n18133), .IN2(n18134), .QN(n18131) );
  INVX0 U19149 ( .INP(n18135), .ZN(n18134) );
  NAND2X0 U19150 ( .IN1(n9745), .IN2(WX861), .QN(n18135) );
  NOR2X0 U19151 ( .IN1(WX861), .IN2(n9745), .QN(n18133) );
  NOR2X0 U19152 ( .IN1(n18136), .IN2(n18137), .QN(n18127) );
  INVX0 U19153 ( .INP(n18138), .ZN(n18137) );
  NAND2X0 U19154 ( .IN1(n3505), .IN2(n10016), .QN(n18138) );
  NOR2X0 U19155 ( .IN1(n10010), .IN2(n3505), .QN(n18136) );
  NAND2X0 U19156 ( .IN1(n18139), .IN2(n18140), .QN(DATA_9_18) );
  INVX0 U19157 ( .INP(n18141), .ZN(n18140) );
  NOR2X0 U19158 ( .IN1(n18142), .IN2(n10614), .QN(n18141) );
  NAND2X0 U19159 ( .IN1(n10614), .IN2(n18142), .QN(n18139) );
  NAND2X0 U19160 ( .IN1(TM0), .IN2(WX511), .QN(n18142) );
  NAND2X0 U19161 ( .IN1(n18143), .IN2(n18144), .QN(n10614) );
  NAND2X0 U19162 ( .IN1(n18145), .IN2(n18146), .QN(n18144) );
  INVX0 U19163 ( .INP(n18147), .ZN(n18143) );
  NOR2X0 U19164 ( .IN1(n18146), .IN2(n18145), .QN(n18147) );
  NAND2X0 U19165 ( .IN1(n18148), .IN2(n18149), .QN(n18145) );
  NAND2X0 U19166 ( .IN1(n9758), .IN2(n18150), .QN(n18149) );
  INVX0 U19167 ( .INP(n18151), .ZN(n18148) );
  NOR2X0 U19168 ( .IN1(n18150), .IN2(n9758), .QN(n18151) );
  NOR2X0 U19169 ( .IN1(n18152), .IN2(n18153), .QN(n18150) );
  INVX0 U19170 ( .INP(n18154), .ZN(n18153) );
  NAND2X0 U19171 ( .IN1(n9760), .IN2(WX863), .QN(n18154) );
  NOR2X0 U19172 ( .IN1(WX863), .IN2(n9760), .QN(n18152) );
  NOR2X0 U19173 ( .IN1(n18155), .IN2(n18156), .QN(n18146) );
  INVX0 U19174 ( .INP(n18157), .ZN(n18156) );
  NAND2X0 U19175 ( .IN1(n3503), .IN2(n10016), .QN(n18157) );
  NOR2X0 U19176 ( .IN1(n10010), .IN2(n3503), .QN(n18155) );
  NAND2X0 U19177 ( .IN1(n18158), .IN2(n18159), .QN(DATA_9_17) );
  INVX0 U19178 ( .INP(n18160), .ZN(n18159) );
  NOR2X0 U19179 ( .IN1(n18161), .IN2(n10583), .QN(n18160) );
  NAND2X0 U19180 ( .IN1(n10583), .IN2(n18161), .QN(n18158) );
  NAND2X0 U19181 ( .IN1(TM0), .IN2(WX513), .QN(n18161) );
  NAND2X0 U19182 ( .IN1(n18162), .IN2(n18163), .QN(n10583) );
  NAND2X0 U19183 ( .IN1(n18164), .IN2(n18165), .QN(n18163) );
  INVX0 U19184 ( .INP(n18166), .ZN(n18162) );
  NOR2X0 U19185 ( .IN1(n18165), .IN2(n18164), .QN(n18166) );
  NAND2X0 U19186 ( .IN1(n18167), .IN2(n18168), .QN(n18164) );
  NAND2X0 U19187 ( .IN1(n9770), .IN2(n18169), .QN(n18168) );
  INVX0 U19188 ( .INP(n18170), .ZN(n18167) );
  NOR2X0 U19189 ( .IN1(n18169), .IN2(n9770), .QN(n18170) );
  NOR2X0 U19190 ( .IN1(n18171), .IN2(n18172), .QN(n18169) );
  INVX0 U19191 ( .INP(n18173), .ZN(n18172) );
  NAND2X0 U19192 ( .IN1(n9772), .IN2(WX865), .QN(n18173) );
  NOR2X0 U19193 ( .IN1(WX865), .IN2(n9772), .QN(n18171) );
  NOR2X0 U19194 ( .IN1(n18174), .IN2(n18175), .QN(n18165) );
  INVX0 U19195 ( .INP(n18176), .ZN(n18175) );
  NAND2X0 U19196 ( .IN1(n3501), .IN2(n10016), .QN(n18176) );
  NOR2X0 U19197 ( .IN1(n10010), .IN2(n3501), .QN(n18174) );
  NOR2X0 U19198 ( .IN1(n18177), .IN2(n18178), .QN(DATA_9_16) );
  INVX0 U19199 ( .INP(n18179), .ZN(n18178) );
  NAND2X0 U19200 ( .IN1(n18180), .IN2(n10562), .QN(n18179) );
  NOR2X0 U19201 ( .IN1(n10562), .IN2(n18180), .QN(n18177) );
  NAND2X0 U19202 ( .IN1(TM0), .IN2(WX515), .QN(n18180) );
  NAND2X0 U19203 ( .IN1(n18181), .IN2(n18182), .QN(n10562) );
  NAND2X0 U19204 ( .IN1(n18183), .IN2(n18184), .QN(n18182) );
  NAND2X0 U19205 ( .IN1(n18185), .IN2(n18186), .QN(n18183) );
  NAND2X0 U19206 ( .IN1(n3499), .IN2(n10016), .QN(n18186) );
  NAND2X0 U19207 ( .IN1(TM1), .IN2(WX675), .QN(n18185) );
  NAND2X0 U19208 ( .IN1(n18187), .IN2(n18188), .QN(n18181) );
  NOR2X0 U19209 ( .IN1(n18189), .IN2(n18190), .QN(n18188) );
  NOR2X0 U19210 ( .IN1(n3499), .IN2(n10003), .QN(n18190) );
  INVX0 U19211 ( .INP(TM1), .ZN(n11655) );
  NOR2X0 U19212 ( .IN1(TM1), .IN2(WX675), .QN(n18189) );
  INVX0 U19213 ( .INP(n18184), .ZN(n18187) );
  NOR2X0 U19214 ( .IN1(n18191), .IN2(n18192), .QN(n18184) );
  INVX0 U19215 ( .INP(n18193), .ZN(n18192) );
  NAND2X0 U19216 ( .IN1(n9787), .IN2(n18194), .QN(n18193) );
  NOR2X0 U19217 ( .IN1(n18194), .IN2(n9787), .QN(n18191) );
  NOR2X0 U19218 ( .IN1(n18195), .IN2(n18196), .QN(n18194) );
  NOR2X0 U19219 ( .IN1(n9851), .IN2(n9788), .QN(n18196) );
  INVX0 U19220 ( .INP(n18197), .ZN(n18195) );
  NAND2X0 U19221 ( .IN1(n9788), .IN2(n9851), .QN(n18197) );
  NAND2X0 U19222 ( .IN1(n18198), .IN2(n18199), .QN(DATA_9_15) );
  INVX0 U19223 ( .INP(n18200), .ZN(n18199) );
  NOR2X0 U19224 ( .IN1(n18201), .IN2(n10551), .QN(n18200) );
  NAND2X0 U19225 ( .IN1(n10551), .IN2(n18201), .QN(n18198) );
  NAND2X0 U19226 ( .IN1(TM0), .IN2(WX517), .QN(n18201) );
  NAND2X0 U19227 ( .IN1(n18202), .IN2(n18203), .QN(n10551) );
  NAND2X0 U19228 ( .IN1(n18204), .IN2(n18205), .QN(n18203) );
  INVX0 U19229 ( .INP(n18206), .ZN(n18202) );
  NOR2X0 U19230 ( .IN1(n18205), .IN2(n18204), .QN(n18206) );
  NAND2X0 U19231 ( .IN1(n18207), .IN2(n18208), .QN(n18204) );
  NAND2X0 U19232 ( .IN1(n9801), .IN2(n18209), .QN(n18208) );
  INVX0 U19233 ( .INP(n18210), .ZN(n18207) );
  NOR2X0 U19234 ( .IN1(n18209), .IN2(n9801), .QN(n18210) );
  NOR2X0 U19235 ( .IN1(n18211), .IN2(n18212), .QN(n18209) );
  NOR2X0 U19236 ( .IN1(WX869), .IN2(n9802), .QN(n18212) );
  INVX0 U19237 ( .INP(n18213), .ZN(n18211) );
  NAND2X0 U19238 ( .IN1(n9802), .IN2(WX869), .QN(n18213) );
  NOR2X0 U19239 ( .IN1(n18214), .IN2(n18215), .QN(n18205) );
  INVX0 U19240 ( .INP(n18216), .ZN(n18215) );
  NAND2X0 U19241 ( .IN1(n3497), .IN2(n2340), .QN(n18216) );
  NOR2X0 U19242 ( .IN1(n2340), .IN2(n3497), .QN(n18214) );
  NAND2X0 U19243 ( .IN1(n18217), .IN2(n18218), .QN(DATA_9_14) );
  INVX0 U19244 ( .INP(n18219), .ZN(n18218) );
  NOR2X0 U19245 ( .IN1(n18220), .IN2(n10542), .QN(n18219) );
  NAND2X0 U19246 ( .IN1(n10542), .IN2(n18220), .QN(n18217) );
  NAND2X0 U19247 ( .IN1(test_so1), .IN2(TM0), .QN(n18220) );
  NAND2X0 U19248 ( .IN1(n18221), .IN2(n18222), .QN(n10542) );
  NAND2X0 U19249 ( .IN1(n18223), .IN2(n18224), .QN(n18222) );
  INVX0 U19250 ( .INP(n18225), .ZN(n18221) );
  NOR2X0 U19251 ( .IN1(n18224), .IN2(n18223), .QN(n18225) );
  NAND2X0 U19252 ( .IN1(n18226), .IN2(n18227), .QN(n18223) );
  NAND2X0 U19253 ( .IN1(n9814), .IN2(n18228), .QN(n18227) );
  INVX0 U19254 ( .INP(n18229), .ZN(n18226) );
  NOR2X0 U19255 ( .IN1(n18228), .IN2(n9814), .QN(n18229) );
  NOR2X0 U19256 ( .IN1(n18230), .IN2(n18231), .QN(n18228) );
  INVX0 U19257 ( .INP(n18232), .ZN(n18231) );
  NAND2X0 U19258 ( .IN1(n9816), .IN2(WX871), .QN(n18232) );
  NOR2X0 U19259 ( .IN1(WX871), .IN2(n9816), .QN(n18230) );
  NOR2X0 U19260 ( .IN1(n18233), .IN2(n18234), .QN(n18224) );
  INVX0 U19261 ( .INP(n18235), .ZN(n18234) );
  NAND2X0 U19262 ( .IN1(n3495), .IN2(n2340), .QN(n18235) );
  NOR2X0 U19263 ( .IN1(n2340), .IN2(n3495), .QN(n18233) );
  NAND2X0 U19264 ( .IN1(n18236), .IN2(n18237), .QN(DATA_9_13) );
  INVX0 U19265 ( .INP(n18238), .ZN(n18237) );
  NOR2X0 U19266 ( .IN1(n18239), .IN2(n10532), .QN(n18238) );
  NAND2X0 U19267 ( .IN1(n10532), .IN2(n18239), .QN(n18236) );
  NAND2X0 U19268 ( .IN1(TM0), .IN2(WX521), .QN(n18239) );
  NAND2X0 U19269 ( .IN1(n18240), .IN2(n18241), .QN(n10532) );
  NAND2X0 U19270 ( .IN1(n18242), .IN2(n18243), .QN(n18241) );
  INVX0 U19271 ( .INP(n18244), .ZN(n18240) );
  NOR2X0 U19272 ( .IN1(n18243), .IN2(n18242), .QN(n18244) );
  NAND2X0 U19273 ( .IN1(n18245), .IN2(n18246), .QN(n18242) );
  NAND2X0 U19274 ( .IN1(n9749), .IN2(n18247), .QN(n18246) );
  INVX0 U19275 ( .INP(n18248), .ZN(n18245) );
  NOR2X0 U19276 ( .IN1(n18247), .IN2(n9749), .QN(n18248) );
  NOR2X0 U19277 ( .IN1(n18249), .IN2(n18250), .QN(n18247) );
  INVX0 U19278 ( .INP(n18251), .ZN(n18250) );
  NAND2X0 U19279 ( .IN1(n9751), .IN2(WX873), .QN(n18251) );
  NOR2X0 U19280 ( .IN1(WX873), .IN2(n9751), .QN(n18249) );
  NOR2X0 U19281 ( .IN1(n18252), .IN2(n18253), .QN(n18243) );
  INVX0 U19282 ( .INP(n18254), .ZN(n18253) );
  NAND2X0 U19283 ( .IN1(n3493), .IN2(n2340), .QN(n18254) );
  NOR2X0 U19284 ( .IN1(n2340), .IN2(n3493), .QN(n18252) );
  NAND2X0 U19285 ( .IN1(n18255), .IN2(n18256), .QN(DATA_9_12) );
  INVX0 U19286 ( .INP(n18257), .ZN(n18256) );
  NOR2X0 U19287 ( .IN1(n18258), .IN2(n10521), .QN(n18257) );
  NAND2X0 U19288 ( .IN1(n10521), .IN2(n18258), .QN(n18255) );
  NAND2X0 U19289 ( .IN1(TM0), .IN2(WX523), .QN(n18258) );
  NAND2X0 U19290 ( .IN1(n18259), .IN2(n18260), .QN(n10521) );
  NAND2X0 U19291 ( .IN1(n18261), .IN2(n18262), .QN(n18260) );
  INVX0 U19292 ( .INP(n18263), .ZN(n18259) );
  NOR2X0 U19293 ( .IN1(n18262), .IN2(n18261), .QN(n18263) );
  NAND2X0 U19294 ( .IN1(n18264), .IN2(n18265), .QN(n18261) );
  NAND2X0 U19295 ( .IN1(n9776), .IN2(n18266), .QN(n18265) );
  INVX0 U19296 ( .INP(n18267), .ZN(n18264) );
  NOR2X0 U19297 ( .IN1(n18266), .IN2(n9776), .QN(n18267) );
  NOR2X0 U19298 ( .IN1(n18268), .IN2(n18269), .QN(n18266) );
  INVX0 U19299 ( .INP(n18270), .ZN(n18269) );
  NAND2X0 U19300 ( .IN1(n9778), .IN2(WX875), .QN(n18270) );
  NOR2X0 U19301 ( .IN1(WX875), .IN2(n9778), .QN(n18268) );
  NOR2X0 U19302 ( .IN1(n18271), .IN2(n18272), .QN(n18262) );
  INVX0 U19303 ( .INP(n18273), .ZN(n18272) );
  NAND2X0 U19304 ( .IN1(n3491), .IN2(n2340), .QN(n18273) );
  NOR2X0 U19305 ( .IN1(n2340), .IN2(n3491), .QN(n18271) );
  NAND2X0 U19306 ( .IN1(n18274), .IN2(n18275), .QN(DATA_9_11) );
  INVX0 U19307 ( .INP(n18276), .ZN(n18275) );
  NOR2X0 U19308 ( .IN1(n18277), .IN2(n11320), .QN(n18276) );
  NAND2X0 U19309 ( .IN1(n11320), .IN2(n18277), .QN(n18274) );
  NAND2X0 U19310 ( .IN1(TM0), .IN2(WX525), .QN(n18277) );
  NAND2X0 U19311 ( .IN1(n18278), .IN2(n18279), .QN(n11320) );
  NAND2X0 U19312 ( .IN1(n18280), .IN2(n18281), .QN(n18279) );
  INVX0 U19313 ( .INP(n18282), .ZN(n18278) );
  NOR2X0 U19314 ( .IN1(n18281), .IN2(n18280), .QN(n18282) );
  NAND2X0 U19315 ( .IN1(n18283), .IN2(n18284), .QN(n18280) );
  NAND2X0 U19316 ( .IN1(n9822), .IN2(n18285), .QN(n18284) );
  INVX0 U19317 ( .INP(n18286), .ZN(n18283) );
  NOR2X0 U19318 ( .IN1(n18285), .IN2(n9822), .QN(n18286) );
  NOR2X0 U19319 ( .IN1(n18287), .IN2(n18288), .QN(n18285) );
  INVX0 U19320 ( .INP(n18289), .ZN(n18288) );
  NAND2X0 U19321 ( .IN1(n9824), .IN2(WX877), .QN(n18289) );
  NOR2X0 U19322 ( .IN1(WX877), .IN2(n9824), .QN(n18287) );
  NOR2X0 U19323 ( .IN1(n18290), .IN2(n18291), .QN(n18281) );
  INVX0 U19324 ( .INP(n18292), .ZN(n18291) );
  NAND2X0 U19325 ( .IN1(n3489), .IN2(n2340), .QN(n18292) );
  NOR2X0 U19326 ( .IN1(n2340), .IN2(n3489), .QN(n18290) );
  NOR2X0 U19327 ( .IN1(n18293), .IN2(n18294), .QN(DATA_9_10) );
  INVX0 U19328 ( .INP(n18295), .ZN(n18294) );
  NAND2X0 U19329 ( .IN1(n18296), .IN2(n11311), .QN(n18295) );
  NOR2X0 U19330 ( .IN1(n11311), .IN2(n18296), .QN(n18293) );
  NAND2X0 U19331 ( .IN1(TM0), .IN2(WX527), .QN(n18296) );
  NAND2X0 U19332 ( .IN1(n18297), .IN2(n18298), .QN(n11311) );
  NAND2X0 U19333 ( .IN1(n18299), .IN2(n18300), .QN(n18298) );
  NAND2X0 U19334 ( .IN1(n18301), .IN2(n18302), .QN(n18299) );
  NAND2X0 U19335 ( .IN1(n9769), .IN2(n2340), .QN(n18302) );
  NAND2X0 U19336 ( .IN1(TM0), .IN2(WX751), .QN(n18301) );
  NAND2X0 U19337 ( .IN1(n18303), .IN2(n18304), .QN(n18297) );
  NOR2X0 U19338 ( .IN1(n18305), .IN2(n18306), .QN(n18304) );
  NOR2X0 U19339 ( .IN1(n9769), .IN2(n2340), .QN(n18306) );
  NOR2X0 U19340 ( .IN1(TM0), .IN2(WX751), .QN(n18305) );
  INVX0 U19341 ( .INP(n18300), .ZN(n18303) );
  NOR2X0 U19342 ( .IN1(n18307), .IN2(n18308), .QN(n18300) );
  INVX0 U19343 ( .INP(n18309), .ZN(n18308) );
  NAND2X0 U19344 ( .IN1(n9767), .IN2(n18310), .QN(n18309) );
  NOR2X0 U19345 ( .IN1(n18310), .IN2(n9767), .QN(n18307) );
  NOR2X0 U19346 ( .IN1(n18311), .IN2(n18312), .QN(n18310) );
  INVX0 U19347 ( .INP(n18313), .ZN(n18312) );
  NAND2X0 U19348 ( .IN1(test_so3), .IN2(WX879), .QN(n18313) );
  NOR2X0 U19349 ( .IN1(WX879), .IN2(test_so3), .QN(n18311) );
  NAND2X0 U19350 ( .IN1(n18314), .IN2(n18315), .QN(DATA_9_1) );
  INVX0 U19351 ( .INP(n18316), .ZN(n18315) );
  NOR2X0 U19352 ( .IN1(n18317), .IN2(n11158), .QN(n18316) );
  NAND2X0 U19353 ( .IN1(n11158), .IN2(n18317), .QN(n18314) );
  NAND2X0 U19354 ( .IN1(TM0), .IN2(WX545), .QN(n18317) );
  NAND2X0 U19355 ( .IN1(n18318), .IN2(n18319), .QN(n11158) );
  NAND2X0 U19356 ( .IN1(n18320), .IN2(n18321), .QN(n18319) );
  INVX0 U19357 ( .INP(n18322), .ZN(n18318) );
  NOR2X0 U19358 ( .IN1(n18321), .IN2(n18320), .QN(n18322) );
  NAND2X0 U19359 ( .IN1(n18323), .IN2(n18324), .QN(n18320) );
  NAND2X0 U19360 ( .IN1(n9752), .IN2(n18325), .QN(n18324) );
  INVX0 U19361 ( .INP(n18326), .ZN(n18325) );
  NAND2X0 U19362 ( .IN1(n18326), .IN2(WX897), .QN(n18323) );
  NAND2X0 U19363 ( .IN1(n18327), .IN2(n18328), .QN(n18326) );
  INVX0 U19364 ( .INP(n18329), .ZN(n18328) );
  NOR2X0 U19365 ( .IN1(WX833), .IN2(n9753), .QN(n18329) );
  NAND2X0 U19366 ( .IN1(n9753), .IN2(WX833), .QN(n18327) );
  NOR2X0 U19367 ( .IN1(n18330), .IN2(n18331), .QN(n18321) );
  INVX0 U19368 ( .INP(n18332), .ZN(n18331) );
  NAND2X0 U19369 ( .IN1(n3469), .IN2(n2340), .QN(n18332) );
  NOR2X0 U19370 ( .IN1(n2340), .IN2(n3469), .QN(n18330) );
  NAND2X0 U19371 ( .IN1(n18333), .IN2(n18334), .QN(DATA_9_0) );
  INVX0 U19372 ( .INP(n18335), .ZN(n18334) );
  NOR2X0 U19373 ( .IN1(n18336), .IN2(n11148), .QN(n18335) );
  NAND2X0 U19374 ( .IN1(n11148), .IN2(n18336), .QN(n18333) );
  NAND2X0 U19375 ( .IN1(TM0), .IN2(WX547), .QN(n18336) );
  NAND2X0 U19376 ( .IN1(n18337), .IN2(n18338), .QN(n11148) );
  NAND2X0 U19377 ( .IN1(n18339), .IN2(n18340), .QN(n18338) );
  INVX0 U19378 ( .INP(n18341), .ZN(n18337) );
  NOR2X0 U19379 ( .IN1(n18340), .IN2(n18339), .QN(n18341) );
  NAND2X0 U19380 ( .IN1(n18342), .IN2(n18343), .QN(n18339) );
  NAND2X0 U19381 ( .IN1(n9825), .IN2(n18344), .QN(n18343) );
  INVX0 U19382 ( .INP(n18345), .ZN(n18342) );
  NOR2X0 U19383 ( .IN1(n18344), .IN2(n9825), .QN(n18345) );
  NOR2X0 U19384 ( .IN1(n18346), .IN2(n18347), .QN(n18344) );
  NOR2X0 U19385 ( .IN1(WX899), .IN2(n9826), .QN(n18347) );
  INVX0 U19386 ( .INP(n18348), .ZN(n18346) );
  NAND2X0 U19387 ( .IN1(n9826), .IN2(WX899), .QN(n18348) );
  NOR2X0 U19388 ( .IN1(n18349), .IN2(n18350), .QN(n18340) );
  INVX0 U19389 ( .INP(n18351), .ZN(n18350) );
  NAND2X0 U19390 ( .IN1(n3467), .IN2(n2340), .QN(n18351) );
  NOR2X0 U19391 ( .IN1(n2340), .IN2(n3467), .QN(n18349) );
  INVX0 U19392 ( .INP(TM0), .ZN(n2340) );
  INVX0 U3558_U2 ( .INP(n2339), .ZN(U3558_n1) );
  NOR2X0 U3558_U1 ( .IN1(n10300), .IN2(U3558_n1), .QN(n2245) );
  INVX0 U3871_U2 ( .INP(n3278), .ZN(U3871_n1) );
  NOR2X0 U3871_U1 ( .IN1(TM0), .IN2(U3871_n1), .QN(n2153) );
  INVX0 U3991_U2 ( .INP(n3278), .ZN(U3991_n1) );
  NOR2X1 U3991_U1 ( .IN1(n2340), .IN2(U3991_n1), .QN(n2152) );
  INVX0 U5716_U2 ( .INP(WX547), .ZN(U5716_n1) );
  NOR2X0 U5716_U1 ( .IN1(n10287), .IN2(U5716_n1), .QN(WX544) );
  INVX0 U5717_U2 ( .INP(WX545), .ZN(U5717_n1) );
  NOR2X0 U5717_U1 ( .IN1(n10287), .IN2(U5717_n1), .QN(WX542) );
  INVX0 U5718_U2 ( .INP(WX543), .ZN(U5718_n1) );
  NOR2X0 U5718_U1 ( .IN1(n10287), .IN2(U5718_n1), .QN(WX540) );
  INVX0 U5719_U2 ( .INP(WX541), .ZN(U5719_n1) );
  NOR2X0 U5719_U1 ( .IN1(n10287), .IN2(U5719_n1), .QN(WX538) );
  INVX0 U5720_U2 ( .INP(WX539), .ZN(U5720_n1) );
  NOR2X0 U5720_U1 ( .IN1(n10287), .IN2(U5720_n1), .QN(WX536) );
  INVX0 U5721_U2 ( .INP(WX537), .ZN(U5721_n1) );
  NOR2X0 U5721_U1 ( .IN1(n10287), .IN2(U5721_n1), .QN(WX534) );
  INVX0 U5722_U2 ( .INP(WX535), .ZN(U5722_n1) );
  NOR2X0 U5722_U1 ( .IN1(n10286), .IN2(U5722_n1), .QN(WX532) );
  INVX0 U5723_U2 ( .INP(WX533), .ZN(U5723_n1) );
  NOR2X0 U5723_U1 ( .IN1(n10286), .IN2(U5723_n1), .QN(WX530) );
  INVX0 U5724_U2 ( .INP(WX531), .ZN(U5724_n1) );
  NOR2X0 U5724_U1 ( .IN1(n10286), .IN2(U5724_n1), .QN(WX528) );
  INVX0 U5725_U2 ( .INP(WX529), .ZN(U5725_n1) );
  NOR2X0 U5725_U1 ( .IN1(n10286), .IN2(U5725_n1), .QN(WX526) );
  INVX0 U5726_U2 ( .INP(WX527), .ZN(U5726_n1) );
  NOR2X0 U5726_U1 ( .IN1(n10286), .IN2(U5726_n1), .QN(WX524) );
  INVX0 U5727_U2 ( .INP(WX525), .ZN(U5727_n1) );
  NOR2X0 U5727_U1 ( .IN1(n10286), .IN2(U5727_n1), .QN(WX522) );
  INVX0 U5728_U2 ( .INP(WX523), .ZN(U5728_n1) );
  NOR2X0 U5728_U1 ( .IN1(n10286), .IN2(U5728_n1), .QN(WX520) );
  INVX0 U5729_U2 ( .INP(WX521), .ZN(U5729_n1) );
  NOR2X0 U5729_U1 ( .IN1(n10286), .IN2(U5729_n1), .QN(WX518) );
  INVX0 U5730_U2 ( .INP(test_so1), .ZN(U5730_n1) );
  NOR2X0 U5730_U1 ( .IN1(n10286), .IN2(U5730_n1), .QN(WX516) );
  INVX0 U5731_U2 ( .INP(WX517), .ZN(U5731_n1) );
  NOR2X0 U5731_U1 ( .IN1(n10286), .IN2(U5731_n1), .QN(WX514) );
  INVX0 U5732_U2 ( .INP(WX515), .ZN(U5732_n1) );
  NOR2X0 U5732_U1 ( .IN1(n10283), .IN2(U5732_n1), .QN(WX512) );
  INVX0 U5733_U2 ( .INP(WX513), .ZN(U5733_n1) );
  NOR2X0 U5733_U1 ( .IN1(n10283), .IN2(U5733_n1), .QN(WX510) );
  INVX0 U5734_U2 ( .INP(WX511), .ZN(U5734_n1) );
  NOR2X0 U5734_U1 ( .IN1(n10283), .IN2(U5734_n1), .QN(WX508) );
  INVX0 U5735_U2 ( .INP(WX509), .ZN(U5735_n1) );
  NOR2X0 U5735_U1 ( .IN1(n10282), .IN2(U5735_n1), .QN(WX506) );
  INVX0 U5736_U2 ( .INP(WX507), .ZN(U5736_n1) );
  NOR2X0 U5736_U1 ( .IN1(n10282), .IN2(U5736_n1), .QN(WX504) );
  INVX0 U5737_U2 ( .INP(WX505), .ZN(U5737_n1) );
  NOR2X0 U5737_U1 ( .IN1(n10282), .IN2(U5737_n1), .QN(WX502) );
  INVX0 U5738_U2 ( .INP(WX503), .ZN(U5738_n1) );
  NOR2X0 U5738_U1 ( .IN1(n10282), .IN2(U5738_n1), .QN(WX500) );
  INVX0 U5739_U2 ( .INP(WX501), .ZN(U5739_n1) );
  NOR2X0 U5739_U1 ( .IN1(n10282), .IN2(U5739_n1), .QN(WX498) );
  INVX0 U5740_U2 ( .INP(WX499), .ZN(U5740_n1) );
  NOR2X0 U5740_U1 ( .IN1(n10282), .IN2(U5740_n1), .QN(WX496) );
  INVX0 U5741_U2 ( .INP(WX497), .ZN(U5741_n1) );
  NOR2X0 U5741_U1 ( .IN1(n10282), .IN2(U5741_n1), .QN(WX494) );
  INVX0 U5742_U2 ( .INP(WX495), .ZN(U5742_n1) );
  NOR2X0 U5742_U1 ( .IN1(n10282), .IN2(U5742_n1), .QN(WX492) );
  INVX0 U5743_U2 ( .INP(WX493), .ZN(U5743_n1) );
  NOR2X0 U5743_U1 ( .IN1(n10282), .IN2(U5743_n1), .QN(WX490) );
  INVX0 U5744_U2 ( .INP(WX491), .ZN(U5744_n1) );
  NOR2X0 U5744_U1 ( .IN1(n10282), .IN2(U5744_n1), .QN(WX488) );
  INVX0 U5745_U2 ( .INP(WX489), .ZN(U5745_n1) );
  NOR2X0 U5745_U1 ( .IN1(n10281), .IN2(U5745_n1), .QN(WX486) );
  INVX0 U5746_U2 ( .INP(WX487), .ZN(U5746_n1) );
  NOR2X0 U5746_U1 ( .IN1(n10281), .IN2(U5746_n1), .QN(WX484) );
  INVX0 U5747_U2 ( .INP(WX5939), .ZN(U5747_n1) );
  NOR2X0 U5747_U1 ( .IN1(n10280), .IN2(U5747_n1), .QN(WX6002) );
  INVX0 U5748_U2 ( .INP(test_so49), .ZN(U5748_n1) );
  NOR2X0 U5748_U1 ( .IN1(n10278), .IN2(U5748_n1), .QN(WX6000) );
  INVX0 U5749_U2 ( .INP(WX5935), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n10278), .IN2(U5749_n1), .QN(WX5998) );
  INVX0 U5750_U2 ( .INP(WX5933), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n10278), .IN2(U5750_n1), .QN(WX5996) );
  INVX0 U5751_U2 ( .INP(WX5931), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n10278), .IN2(U5751_n1), .QN(WX5994) );
  INVX0 U5752_U2 ( .INP(WX3269), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n10278), .IN2(U5752_n1), .QN(WX3332) );
  INVX0 U5753_U2 ( .INP(WX3265), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n10278), .IN2(U5753_n1), .QN(WX3328) );
  INVX0 U5754_U2 ( .INP(WX3263), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n10278), .IN2(U5754_n1), .QN(WX3326) );
  INVX0 U5755_U2 ( .INP(WX11179), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n10278), .IN2(U5755_n1), .QN(WX11242) );
  INVX0 U5756_U2 ( .INP(WX11177), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n10278), .IN2(U5756_n1), .QN(WX11240) );
  INVX0 U5757_U2 ( .INP(WX11175), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n10278), .IN2(U5757_n1), .QN(WX11238) );
  INVX0 U5758_U2 ( .INP(WX11173), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n10278), .IN2(U5758_n1), .QN(WX11236) );
  INVX0 U5759_U2 ( .INP(test_so96), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n10277), .IN2(U5759_n1), .QN(WX11234) );
  INVX0 U5760_U2 ( .INP(WX11169), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n10277), .IN2(U5760_n1), .QN(WX11232) );
  INVX0 U5761_U2 ( .INP(WX11167), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n10282), .IN2(U5761_n1), .QN(WX11230) );
  INVX0 U5762_U2 ( .INP(WX11165), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n10267), .IN2(U5762_n1), .QN(WX11228) );
  INVX0 U5763_U2 ( .INP(WX11163), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n10279), .IN2(U5763_n1), .QN(WX11226) );
  INVX0 U5764_U2 ( .INP(WX11161), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n10279), .IN2(U5764_n1), .QN(WX11224) );
  INVX0 U5765_U2 ( .INP(WX11159), .ZN(U5765_n1) );
  NOR2X0 U5765_U1 ( .IN1(n10279), .IN2(U5765_n1), .QN(WX11222) );
  INVX0 U5766_U2 ( .INP(WX11157), .ZN(U5766_n1) );
  NOR2X0 U5766_U1 ( .IN1(n10279), .IN2(U5766_n1), .QN(WX11220) );
  INVX0 U5767_U2 ( .INP(WX11155), .ZN(U5767_n1) );
  NOR2X0 U5767_U1 ( .IN1(n10279), .IN2(U5767_n1), .QN(WX11218) );
  INVX0 U5768_U2 ( .INP(WX11153), .ZN(U5768_n1) );
  NOR2X0 U5768_U1 ( .IN1(n10279), .IN2(U5768_n1), .QN(WX11216) );
  INVX0 U5769_U2 ( .INP(WX11151), .ZN(U5769_n1) );
  NOR2X0 U5769_U1 ( .IN1(n10279), .IN2(U5769_n1), .QN(WX11214) );
  INVX0 U5770_U2 ( .INP(WX11149), .ZN(U5770_n1) );
  NOR2X0 U5770_U1 ( .IN1(n10279), .IN2(U5770_n1), .QN(WX11212) );
  INVX0 U5771_U2 ( .INP(WX11147), .ZN(U5771_n1) );
  NOR2X0 U5771_U1 ( .IN1(n10279), .IN2(U5771_n1), .QN(WX11210) );
  INVX0 U5772_U2 ( .INP(WX11145), .ZN(U5772_n1) );
  NOR2X0 U5772_U1 ( .IN1(n10279), .IN2(U5772_n1), .QN(WX11208) );
  INVX0 U5773_U2 ( .INP(WX11143), .ZN(U5773_n1) );
  NOR2X0 U5773_U1 ( .IN1(n10279), .IN2(U5773_n1), .QN(WX11206) );
  INVX0 U5774_U2 ( .INP(WX11141), .ZN(U5774_n1) );
  NOR2X0 U5774_U1 ( .IN1(n10280), .IN2(U5774_n1), .QN(WX11204) );
  INVX0 U5775_U2 ( .INP(WX11139), .ZN(U5775_n1) );
  NOR2X0 U5775_U1 ( .IN1(n10280), .IN2(U5775_n1), .QN(WX11202) );
  INVX0 U5776_U2 ( .INP(test_so95), .ZN(U5776_n1) );
  NOR2X0 U5776_U1 ( .IN1(n10280), .IN2(U5776_n1), .QN(WX11200) );
  INVX0 U5777_U2 ( .INP(WX11135), .ZN(U5777_n1) );
  NOR2X0 U5777_U1 ( .IN1(n10280), .IN2(U5777_n1), .QN(WX11198) );
  INVX0 U5778_U2 ( .INP(WX11133), .ZN(U5778_n1) );
  NOR2X0 U5778_U1 ( .IN1(n10280), .IN2(U5778_n1), .QN(WX11196) );
  INVX0 U5779_U2 ( .INP(WX11131), .ZN(U5779_n1) );
  NOR2X0 U5779_U1 ( .IN1(n10280), .IN2(U5779_n1), .QN(WX11194) );
  INVX0 U5780_U2 ( .INP(WX11129), .ZN(U5780_n1) );
  NOR2X0 U5780_U1 ( .IN1(n10280), .IN2(U5780_n1), .QN(WX11192) );
  INVX0 U5781_U2 ( .INP(WX11127), .ZN(U5781_n1) );
  NOR2X0 U5781_U1 ( .IN1(n10280), .IN2(U5781_n1), .QN(WX11190) );
  INVX0 U5782_U2 ( .INP(WX11125), .ZN(U5782_n1) );
  NOR2X0 U5782_U1 ( .IN1(n10280), .IN2(U5782_n1), .QN(WX11188) );
  INVX0 U5783_U2 ( .INP(WX11123), .ZN(U5783_n1) );
  NOR2X0 U5783_U1 ( .IN1(n10280), .IN2(U5783_n1), .QN(WX11186) );
  INVX0 U5784_U2 ( .INP(WX11121), .ZN(U5784_n1) );
  NOR2X0 U5784_U1 ( .IN1(n10281), .IN2(U5784_n1), .QN(WX11184) );
  INVX0 U5785_U2 ( .INP(WX11119), .ZN(U5785_n1) );
  NOR2X0 U5785_U1 ( .IN1(n10281), .IN2(U5785_n1), .QN(WX11182) );
  INVX0 U5786_U2 ( .INP(WX11117), .ZN(U5786_n1) );
  NOR2X0 U5786_U1 ( .IN1(n10281), .IN2(U5786_n1), .QN(WX11180) );
  INVX0 U5787_U2 ( .INP(WX11115), .ZN(U5787_n1) );
  NOR2X0 U5787_U1 ( .IN1(n10281), .IN2(U5787_n1), .QN(WX11178) );
  INVX0 U5788_U2 ( .INP(WX11113), .ZN(U5788_n1) );
  NOR2X0 U5788_U1 ( .IN1(n10281), .IN2(U5788_n1), .QN(WX11176) );
  INVX0 U5789_U2 ( .INP(WX11111), .ZN(U5789_n1) );
  NOR2X0 U5789_U1 ( .IN1(n10281), .IN2(U5789_n1), .QN(WX11174) );
  INVX0 U5790_U2 ( .INP(WX11109), .ZN(U5790_n1) );
  NOR2X0 U5790_U1 ( .IN1(n10281), .IN2(U5790_n1), .QN(WX11172) );
  INVX0 U5791_U2 ( .INP(WX11107), .ZN(U5791_n1) );
  NOR2X0 U5791_U1 ( .IN1(n10281), .IN2(U5791_n1), .QN(WX11170) );
  INVX0 U5792_U2 ( .INP(WX11105), .ZN(U5792_n1) );
  NOR2X0 U5792_U1 ( .IN1(n10281), .IN2(U5792_n1), .QN(WX11168) );
  INVX0 U5793_U2 ( .INP(test_so94), .ZN(U5793_n1) );
  NOR2X0 U5793_U1 ( .IN1(n10283), .IN2(U5793_n1), .QN(WX11166) );
  INVX0 U5794_U2 ( .INP(WX11101), .ZN(U5794_n1) );
  NOR2X0 U5794_U1 ( .IN1(n10283), .IN2(U5794_n1), .QN(WX11164) );
  INVX0 U5795_U2 ( .INP(WX11099), .ZN(U5795_n1) );
  NOR2X0 U5795_U1 ( .IN1(n10283), .IN2(U5795_n1), .QN(WX11162) );
  INVX0 U5796_U2 ( .INP(WX11097), .ZN(U5796_n1) );
  NOR2X0 U5796_U1 ( .IN1(n10283), .IN2(U5796_n1), .QN(WX11160) );
  INVX0 U5797_U2 ( .INP(WX11095), .ZN(U5797_n1) );
  NOR2X0 U5797_U1 ( .IN1(n10283), .IN2(U5797_n1), .QN(WX11158) );
  INVX0 U5798_U2 ( .INP(WX11093), .ZN(U5798_n1) );
  NOR2X0 U5798_U1 ( .IN1(n10283), .IN2(U5798_n1), .QN(WX11156) );
  INVX0 U5799_U2 ( .INP(WX11091), .ZN(U5799_n1) );
  NOR2X0 U5799_U1 ( .IN1(n10283), .IN2(U5799_n1), .QN(WX11154) );
  INVX0 U5800_U2 ( .INP(WX11089), .ZN(U5800_n1) );
  NOR2X0 U5800_U1 ( .IN1(n10283), .IN2(U5800_n1), .QN(WX11152) );
  INVX0 U5801_U2 ( .INP(WX11087), .ZN(U5801_n1) );
  NOR2X0 U5801_U1 ( .IN1(n10284), .IN2(U5801_n1), .QN(WX11150) );
  INVX0 U5802_U2 ( .INP(WX11085), .ZN(U5802_n1) );
  NOR2X0 U5802_U1 ( .IN1(n10284), .IN2(U5802_n1), .QN(WX11148) );
  INVX0 U5803_U2 ( .INP(WX11083), .ZN(U5803_n1) );
  NOR2X0 U5803_U1 ( .IN1(n10284), .IN2(U5803_n1), .QN(WX11146) );
  INVX0 U5804_U2 ( .INP(WX11081), .ZN(U5804_n1) );
  NOR2X0 U5804_U1 ( .IN1(n10284), .IN2(U5804_n1), .QN(WX11144) );
  INVX0 U5805_U2 ( .INP(WX11079), .ZN(U5805_n1) );
  NOR2X0 U5805_U1 ( .IN1(n10284), .IN2(U5805_n1), .QN(WX11142) );
  INVX0 U5806_U2 ( .INP(WX11077), .ZN(U5806_n1) );
  NOR2X0 U5806_U1 ( .IN1(n10284), .IN2(U5806_n1), .QN(WX11140) );
  INVX0 U5807_U2 ( .INP(WX11075), .ZN(U5807_n1) );
  NOR2X0 U5807_U1 ( .IN1(n10284), .IN2(U5807_n1), .QN(WX11138) );
  INVX0 U5808_U2 ( .INP(WX11073), .ZN(U5808_n1) );
  NOR2X0 U5808_U1 ( .IN1(n10284), .IN2(U5808_n1), .QN(WX11136) );
  INVX0 U5809_U2 ( .INP(WX11071), .ZN(U5809_n1) );
  NOR2X0 U5809_U1 ( .IN1(n10284), .IN2(U5809_n1), .QN(WX11134) );
  INVX0 U5810_U2 ( .INP(test_so93), .ZN(U5810_n1) );
  NOR2X0 U5810_U1 ( .IN1(n10284), .IN2(U5810_n1), .QN(WX11132) );
  INVX0 U5811_U2 ( .INP(WX11067), .ZN(U5811_n1) );
  NOR2X0 U5811_U1 ( .IN1(n10284), .IN2(U5811_n1), .QN(WX11130) );
  INVX0 U5812_U2 ( .INP(WX11065), .ZN(U5812_n1) );
  NOR2X0 U5812_U1 ( .IN1(n10285), .IN2(U5812_n1), .QN(WX11128) );
  INVX0 U5813_U2 ( .INP(WX11063), .ZN(U5813_n1) );
  NOR2X0 U5813_U1 ( .IN1(n10285), .IN2(U5813_n1), .QN(WX11126) );
  INVX0 U5814_U2 ( .INP(WX11061), .ZN(U5814_n1) );
  NOR2X0 U5814_U1 ( .IN1(n10285), .IN2(U5814_n1), .QN(WX11124) );
  INVX0 U5815_U2 ( .INP(WX11059), .ZN(U5815_n1) );
  NOR2X0 U5815_U1 ( .IN1(n10285), .IN2(U5815_n1), .QN(WX11122) );
  INVX0 U5816_U2 ( .INP(WX11057), .ZN(U5816_n1) );
  NOR2X0 U5816_U1 ( .IN1(n10285), .IN2(U5816_n1), .QN(WX11120) );
  INVX0 U5817_U2 ( .INP(WX11055), .ZN(U5817_n1) );
  NOR2X0 U5817_U1 ( .IN1(n10285), .IN2(U5817_n1), .QN(WX11118) );
  INVX0 U5818_U2 ( .INP(WX11053), .ZN(U5818_n1) );
  NOR2X0 U5818_U1 ( .IN1(n10285), .IN2(U5818_n1), .QN(WX11116) );
  INVX0 U5819_U2 ( .INP(WX11051), .ZN(U5819_n1) );
  NOR2X0 U5819_U1 ( .IN1(n10285), .IN2(U5819_n1), .QN(WX11114) );
  INVX0 U5820_U2 ( .INP(WX11049), .ZN(U5820_n1) );
  NOR2X0 U5820_U1 ( .IN1(n10285), .IN2(U5820_n1), .QN(WX11112) );
  INVX0 U5821_U2 ( .INP(WX11047), .ZN(U5821_n1) );
  NOR2X0 U5821_U1 ( .IN1(n10285), .IN2(U5821_n1), .QN(WX11110) );
  INVX0 U5822_U2 ( .INP(WX11045), .ZN(U5822_n1) );
  NOR2X0 U5822_U1 ( .IN1(n10285), .IN2(U5822_n1), .QN(WX11108) );
  INVX0 U5823_U2 ( .INP(WX11043), .ZN(U5823_n1) );
  NOR2X0 U5823_U1 ( .IN1(n10286), .IN2(U5823_n1), .QN(WX11106) );
  INVX0 U5824_U2 ( .INP(WX11041), .ZN(U5824_n1) );
  NOR2X0 U5824_U1 ( .IN1(n10287), .IN2(U5824_n1), .QN(WX11104) );
  INVX0 U5825_U2 ( .INP(WX11039), .ZN(U5825_n1) );
  NOR2X0 U5825_U1 ( .IN1(n10287), .IN2(U5825_n1), .QN(WX11102) );
  INVX0 U5826_U2 ( .INP(WX11037), .ZN(U5826_n1) );
  NOR2X0 U5826_U1 ( .IN1(n10287), .IN2(U5826_n1), .QN(WX11100) );
  INVX0 U5827_U2 ( .INP(test_so92), .ZN(U5827_n1) );
  NOR2X0 U5827_U1 ( .IN1(n10287), .IN2(U5827_n1), .QN(WX11098) );
  INVX0 U5828_U2 ( .INP(WX11033), .ZN(U5828_n1) );
  NOR2X0 U5828_U1 ( .IN1(n10287), .IN2(U5828_n1), .QN(WX11096) );
  INVX0 U5829_U2 ( .INP(WX11031), .ZN(U5829_n1) );
  NOR2X0 U5829_U1 ( .IN1(n10272), .IN2(U5829_n1), .QN(WX11094) );
  INVX0 U5830_U2 ( .INP(WX11029), .ZN(U5830_n1) );
  NOR2X0 U5830_U1 ( .IN1(n10267), .IN2(U5830_n1), .QN(WX11092) );
  INVX0 U5831_U2 ( .INP(WX11027), .ZN(U5831_n1) );
  NOR2X0 U5831_U1 ( .IN1(n10267), .IN2(U5831_n1), .QN(WX11090) );
  INVX0 U5832_U2 ( .INP(WX11025), .ZN(U5832_n1) );
  NOR2X0 U5832_U1 ( .IN1(n10267), .IN2(U5832_n1), .QN(WX11088) );
  INVX0 U5833_U2 ( .INP(WX11023), .ZN(U5833_n1) );
  NOR2X0 U5833_U1 ( .IN1(n10268), .IN2(U5833_n1), .QN(WX11086) );
  INVX0 U5834_U2 ( .INP(WX11021), .ZN(U5834_n1) );
  NOR2X0 U5834_U1 ( .IN1(n10268), .IN2(U5834_n1), .QN(WX11084) );
  INVX0 U5835_U2 ( .INP(WX9886), .ZN(U5835_n1) );
  NOR2X0 U5835_U1 ( .IN1(n10268), .IN2(U5835_n1), .QN(WX9949) );
  INVX0 U5836_U2 ( .INP(WX9884), .ZN(U5836_n1) );
  NOR2X0 U5836_U1 ( .IN1(n10268), .IN2(U5836_n1), .QN(WX9947) );
  INVX0 U5837_U2 ( .INP(WX9882), .ZN(U5837_n1) );
  NOR2X0 U5837_U1 ( .IN1(n10268), .IN2(U5837_n1), .QN(WX9945) );
  INVX0 U5838_U2 ( .INP(WX9880), .ZN(U5838_n1) );
  NOR2X0 U5838_U1 ( .IN1(n10268), .IN2(U5838_n1), .QN(WX9943) );
  INVX0 U5839_U2 ( .INP(WX9878), .ZN(U5839_n1) );
  NOR2X0 U5839_U1 ( .IN1(n10268), .IN2(U5839_n1), .QN(WX9941) );
  INVX0 U5840_U2 ( .INP(WX9876), .ZN(U5840_n1) );
  NOR2X0 U5840_U1 ( .IN1(n10268), .IN2(U5840_n1), .QN(WX9939) );
  INVX0 U5841_U2 ( .INP(WX9874), .ZN(U5841_n1) );
  NOR2X0 U5841_U1 ( .IN1(n10268), .IN2(U5841_n1), .QN(WX9937) );
  INVX0 U5842_U2 ( .INP(WX9872), .ZN(U5842_n1) );
  NOR2X0 U5842_U1 ( .IN1(n10268), .IN2(U5842_n1), .QN(WX9935) );
  INVX0 U5843_U2 ( .INP(WX9870), .ZN(U5843_n1) );
  NOR2X0 U5843_U1 ( .IN1(n10268), .IN2(U5843_n1), .QN(WX9933) );
  INVX0 U5844_U2 ( .INP(WX9868), .ZN(U5844_n1) );
  NOR2X0 U5844_U1 ( .IN1(n10269), .IN2(U5844_n1), .QN(WX9931) );
  INVX0 U5845_U2 ( .INP(WX9866), .ZN(U5845_n1) );
  NOR2X0 U5845_U1 ( .IN1(n10269), .IN2(U5845_n1), .QN(WX9929) );
  INVX0 U5846_U2 ( .INP(WX9864), .ZN(U5846_n1) );
  NOR2X0 U5846_U1 ( .IN1(n10269), .IN2(U5846_n1), .QN(WX9927) );
  INVX0 U5847_U2 ( .INP(WX9862), .ZN(U5847_n1) );
  NOR2X0 U5847_U1 ( .IN1(n10269), .IN2(U5847_n1), .QN(WX9925) );
  INVX0 U5848_U2 ( .INP(WX9860), .ZN(U5848_n1) );
  NOR2X0 U5848_U1 ( .IN1(n10269), .IN2(U5848_n1), .QN(WX9923) );
  INVX0 U5849_U2 ( .INP(WX9858), .ZN(U5849_n1) );
  NOR2X0 U5849_U1 ( .IN1(n10269), .IN2(U5849_n1), .QN(WX9921) );
  INVX0 U5850_U2 ( .INP(WX9856), .ZN(U5850_n1) );
  NOR2X0 U5850_U1 ( .IN1(n10269), .IN2(U5850_n1), .QN(WX9919) );
  INVX0 U5851_U2 ( .INP(test_so84), .ZN(U5851_n1) );
  NOR2X0 U5851_U1 ( .IN1(n10269), .IN2(U5851_n1), .QN(WX9917) );
  INVX0 U5852_U2 ( .INP(WX9852), .ZN(U5852_n1) );
  NOR2X0 U5852_U1 ( .IN1(n10269), .IN2(U5852_n1), .QN(WX9915) );
  INVX0 U5853_U2 ( .INP(WX9850), .ZN(U5853_n1) );
  NOR2X0 U5853_U1 ( .IN1(n10269), .IN2(U5853_n1), .QN(WX9913) );
  INVX0 U5854_U2 ( .INP(WX9848), .ZN(U5854_n1) );
  NOR2X0 U5854_U1 ( .IN1(n10269), .IN2(U5854_n1), .QN(WX9911) );
  INVX0 U5855_U2 ( .INP(WX9846), .ZN(U5855_n1) );
  NOR2X0 U5855_U1 ( .IN1(n10270), .IN2(U5855_n1), .QN(WX9909) );
  INVX0 U5856_U2 ( .INP(WX9844), .ZN(U5856_n1) );
  NOR2X0 U5856_U1 ( .IN1(n10270), .IN2(U5856_n1), .QN(WX9907) );
  INVX0 U5857_U2 ( .INP(WX9842), .ZN(U5857_n1) );
  NOR2X0 U5857_U1 ( .IN1(n10270), .IN2(U5857_n1), .QN(WX9905) );
  INVX0 U5858_U2 ( .INP(WX9840), .ZN(U5858_n1) );
  NOR2X0 U5858_U1 ( .IN1(n10270), .IN2(U5858_n1), .QN(WX9903) );
  INVX0 U5859_U2 ( .INP(WX9838), .ZN(U5859_n1) );
  NOR2X0 U5859_U1 ( .IN1(n10270), .IN2(U5859_n1), .QN(WX9901) );
  INVX0 U5860_U2 ( .INP(WX9836), .ZN(U5860_n1) );
  NOR2X0 U5860_U1 ( .IN1(n10270), .IN2(U5860_n1), .QN(WX9899) );
  INVX0 U5861_U2 ( .INP(WX9834), .ZN(U5861_n1) );
  NOR2X0 U5861_U1 ( .IN1(n10270), .IN2(U5861_n1), .QN(WX9897) );
  INVX0 U5862_U2 ( .INP(WX9832), .ZN(U5862_n1) );
  NOR2X0 U5862_U1 ( .IN1(n10270), .IN2(U5862_n1), .QN(WX9895) );
  INVX0 U5863_U2 ( .INP(WX9830), .ZN(U5863_n1) );
  NOR2X0 U5863_U1 ( .IN1(n10270), .IN2(U5863_n1), .QN(WX9893) );
  INVX0 U5864_U2 ( .INP(WX9828), .ZN(U5864_n1) );
  NOR2X0 U5864_U1 ( .IN1(n10270), .IN2(U5864_n1), .QN(WX9891) );
  INVX0 U5865_U2 ( .INP(WX9826), .ZN(U5865_n1) );
  NOR2X0 U5865_U1 ( .IN1(n10270), .IN2(U5865_n1), .QN(WX9889) );
  INVX0 U5866_U2 ( .INP(WX9824), .ZN(U5866_n1) );
  NOR2X0 U5866_U1 ( .IN1(n10271), .IN2(U5866_n1), .QN(WX9887) );
  INVX0 U5867_U2 ( .INP(WX9822), .ZN(U5867_n1) );
  NOR2X0 U5867_U1 ( .IN1(n10271), .IN2(U5867_n1), .QN(WX9885) );
  INVX0 U5868_U2 ( .INP(test_so83), .ZN(U5868_n1) );
  NOR2X0 U5868_U1 ( .IN1(n10271), .IN2(U5868_n1), .QN(WX9883) );
  INVX0 U5869_U2 ( .INP(WX9818), .ZN(U5869_n1) );
  NOR2X0 U5869_U1 ( .IN1(n10271), .IN2(U5869_n1), .QN(WX9881) );
  INVX0 U5870_U2 ( .INP(WX9816), .ZN(U5870_n1) );
  NOR2X0 U5870_U1 ( .IN1(n10271), .IN2(U5870_n1), .QN(WX9879) );
  INVX0 U5871_U2 ( .INP(WX9814), .ZN(U5871_n1) );
  NOR2X0 U5871_U1 ( .IN1(n10271), .IN2(U5871_n1), .QN(WX9877) );
  INVX0 U5872_U2 ( .INP(WX9812), .ZN(U5872_n1) );
  NOR2X0 U5872_U1 ( .IN1(n10271), .IN2(U5872_n1), .QN(WX9875) );
  INVX0 U5873_U2 ( .INP(WX9810), .ZN(U5873_n1) );
  NOR2X0 U5873_U1 ( .IN1(n10271), .IN2(U5873_n1), .QN(WX9873) );
  INVX0 U5874_U2 ( .INP(WX9808), .ZN(U5874_n1) );
  NOR2X0 U5874_U1 ( .IN1(n10271), .IN2(U5874_n1), .QN(WX9871) );
  INVX0 U5875_U2 ( .INP(WX9806), .ZN(U5875_n1) );
  NOR2X0 U5875_U1 ( .IN1(n10271), .IN2(U5875_n1), .QN(WX9869) );
  INVX0 U5876_U2 ( .INP(WX9804), .ZN(U5876_n1) );
  NOR2X0 U5876_U1 ( .IN1(n10271), .IN2(U5876_n1), .QN(WX9867) );
  INVX0 U5877_U2 ( .INP(WX9802), .ZN(U5877_n1) );
  NOR2X0 U5877_U1 ( .IN1(n10272), .IN2(U5877_n1), .QN(WX9865) );
  INVX0 U5878_U2 ( .INP(WX9800), .ZN(U5878_n1) );
  NOR2X0 U5878_U1 ( .IN1(n10272), .IN2(U5878_n1), .QN(WX9863) );
  INVX0 U5879_U2 ( .INP(WX9798), .ZN(U5879_n1) );
  NOR2X0 U5879_U1 ( .IN1(n10272), .IN2(U5879_n1), .QN(WX9861) );
  INVX0 U5880_U2 ( .INP(WX9796), .ZN(U5880_n1) );
  NOR2X0 U5880_U1 ( .IN1(n10272), .IN2(U5880_n1), .QN(WX9859) );
  INVX0 U5881_U2 ( .INP(WX9794), .ZN(U5881_n1) );
  NOR2X0 U5881_U1 ( .IN1(n10272), .IN2(U5881_n1), .QN(WX9857) );
  INVX0 U5882_U2 ( .INP(WX9792), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(n10272), .IN2(U5882_n1), .QN(WX9855) );
  INVX0 U5883_U2 ( .INP(WX9790), .ZN(U5883_n1) );
  NOR2X0 U5883_U1 ( .IN1(n10272), .IN2(U5883_n1), .QN(WX9853) );
  INVX0 U5884_U2 ( .INP(WX9788), .ZN(U5884_n1) );
  NOR2X0 U5884_U1 ( .IN1(n10272), .IN2(U5884_n1), .QN(WX9851) );
  INVX0 U5885_U2 ( .INP(test_so82), .ZN(U5885_n1) );
  NOR2X0 U5885_U1 ( .IN1(n10272), .IN2(U5885_n1), .QN(WX9849) );
  INVX0 U5886_U2 ( .INP(WX9784), .ZN(U5886_n1) );
  NOR2X0 U5886_U1 ( .IN1(n10272), .IN2(U5886_n1), .QN(WX9847) );
  INVX0 U5887_U2 ( .INP(WX9782), .ZN(U5887_n1) );
  NOR2X0 U5887_U1 ( .IN1(n10273), .IN2(U5887_n1), .QN(WX9845) );
  INVX0 U5888_U2 ( .INP(WX9780), .ZN(U5888_n1) );
  NOR2X0 U5888_U1 ( .IN1(n10273), .IN2(U5888_n1), .QN(WX9843) );
  INVX0 U5889_U2 ( .INP(WX9778), .ZN(U5889_n1) );
  NOR2X0 U5889_U1 ( .IN1(n10273), .IN2(U5889_n1), .QN(WX9841) );
  INVX0 U5890_U2 ( .INP(WX9776), .ZN(U5890_n1) );
  NOR2X0 U5890_U1 ( .IN1(n10273), .IN2(U5890_n1), .QN(WX9839) );
  INVX0 U5891_U2 ( .INP(WX9774), .ZN(U5891_n1) );
  NOR2X0 U5891_U1 ( .IN1(n10273), .IN2(U5891_n1), .QN(WX9837) );
  INVX0 U5892_U2 ( .INP(WX9772), .ZN(U5892_n1) );
  NOR2X0 U5892_U1 ( .IN1(n10273), .IN2(U5892_n1), .QN(WX9835) );
  INVX0 U5893_U2 ( .INP(WX9770), .ZN(U5893_n1) );
  NOR2X0 U5893_U1 ( .IN1(n10273), .IN2(U5893_n1), .QN(WX9833) );
  INVX0 U5894_U2 ( .INP(WX9768), .ZN(U5894_n1) );
  NOR2X0 U5894_U1 ( .IN1(n10273), .IN2(U5894_n1), .QN(WX9831) );
  INVX0 U5895_U2 ( .INP(WX9766), .ZN(U5895_n1) );
  NOR2X0 U5895_U1 ( .IN1(n10273), .IN2(U5895_n1), .QN(WX9829) );
  INVX0 U5896_U2 ( .INP(WX9764), .ZN(U5896_n1) );
  NOR2X0 U5896_U1 ( .IN1(n10273), .IN2(U5896_n1), .QN(WX9827) );
  INVX0 U5897_U2 ( .INP(WX9762), .ZN(U5897_n1) );
  NOR2X0 U5897_U1 ( .IN1(n10273), .IN2(U5897_n1), .QN(WX9825) );
  INVX0 U5898_U2 ( .INP(WX9760), .ZN(U5898_n1) );
  NOR2X0 U5898_U1 ( .IN1(n10274), .IN2(U5898_n1), .QN(WX9823) );
  INVX0 U5899_U2 ( .INP(WX9758), .ZN(U5899_n1) );
  NOR2X0 U5899_U1 ( .IN1(n10274), .IN2(U5899_n1), .QN(WX9821) );
  INVX0 U5900_U2 ( .INP(WX9756), .ZN(U5900_n1) );
  NOR2X0 U5900_U1 ( .IN1(n10274), .IN2(U5900_n1), .QN(WX9819) );
  INVX0 U5901_U2 ( .INP(WX9754), .ZN(U5901_n1) );
  NOR2X0 U5901_U1 ( .IN1(n10274), .IN2(U5901_n1), .QN(WX9817) );
  INVX0 U5902_U2 ( .INP(test_so81), .ZN(U5902_n1) );
  NOR2X0 U5902_U1 ( .IN1(n10274), .IN2(U5902_n1), .QN(WX9815) );
  INVX0 U5903_U2 ( .INP(WX9750), .ZN(U5903_n1) );
  NOR2X0 U5903_U1 ( .IN1(n10274), .IN2(U5903_n1), .QN(WX9813) );
  INVX0 U5904_U2 ( .INP(WX9748), .ZN(U5904_n1) );
  NOR2X0 U5904_U1 ( .IN1(n10274), .IN2(U5904_n1), .QN(WX9811) );
  INVX0 U5905_U2 ( .INP(WX9746), .ZN(U5905_n1) );
  NOR2X0 U5905_U1 ( .IN1(n10274), .IN2(U5905_n1), .QN(WX9809) );
  INVX0 U5906_U2 ( .INP(WX9744), .ZN(U5906_n1) );
  NOR2X0 U5906_U1 ( .IN1(n10274), .IN2(U5906_n1), .QN(WX9807) );
  INVX0 U5907_U2 ( .INP(WX9742), .ZN(U5907_n1) );
  NOR2X0 U5907_U1 ( .IN1(n10274), .IN2(U5907_n1), .QN(WX9805) );
  INVX0 U5908_U2 ( .INP(WX9740), .ZN(U5908_n1) );
  NOR2X0 U5908_U1 ( .IN1(n10274), .IN2(U5908_n1), .QN(WX9803) );
  INVX0 U5909_U2 ( .INP(WX9738), .ZN(U5909_n1) );
  NOR2X0 U5909_U1 ( .IN1(n10275), .IN2(U5909_n1), .QN(WX9801) );
  INVX0 U5910_U2 ( .INP(WX9736), .ZN(U5910_n1) );
  NOR2X0 U5910_U1 ( .IN1(n10275), .IN2(U5910_n1), .QN(WX9799) );
  INVX0 U5911_U2 ( .INP(WX9734), .ZN(U5911_n1) );
  NOR2X0 U5911_U1 ( .IN1(n10275), .IN2(U5911_n1), .QN(WX9797) );
  INVX0 U5912_U2 ( .INP(WX9732), .ZN(U5912_n1) );
  NOR2X0 U5912_U1 ( .IN1(n10275), .IN2(U5912_n1), .QN(WX9795) );
  INVX0 U5913_U2 ( .INP(WX9730), .ZN(U5913_n1) );
  NOR2X0 U5913_U1 ( .IN1(n10275), .IN2(U5913_n1), .QN(WX9793) );
  INVX0 U5914_U2 ( .INP(WX9728), .ZN(U5914_n1) );
  NOR2X0 U5914_U1 ( .IN1(n10275), .IN2(U5914_n1), .QN(WX9791) );
  INVX0 U5915_U2 ( .INP(WX8593), .ZN(U5915_n1) );
  NOR2X0 U5915_U1 ( .IN1(n10275), .IN2(U5915_n1), .QN(WX8656) );
  INVX0 U5916_U2 ( .INP(WX8591), .ZN(U5916_n1) );
  NOR2X0 U5916_U1 ( .IN1(n10275), .IN2(U5916_n1), .QN(WX8654) );
  INVX0 U5917_U2 ( .INP(WX8589), .ZN(U5917_n1) );
  NOR2X0 U5917_U1 ( .IN1(n10275), .IN2(U5917_n1), .QN(WX8652) );
  INVX0 U5918_U2 ( .INP(WX8587), .ZN(U5918_n1) );
  NOR2X0 U5918_U1 ( .IN1(n10275), .IN2(U5918_n1), .QN(WX8650) );
  INVX0 U5919_U2 ( .INP(WX8585), .ZN(U5919_n1) );
  NOR2X0 U5919_U1 ( .IN1(n10275), .IN2(U5919_n1), .QN(WX8648) );
  INVX0 U5920_U2 ( .INP(WX8583), .ZN(U5920_n1) );
  NOR2X0 U5920_U1 ( .IN1(n10276), .IN2(U5920_n1), .QN(WX8646) );
  INVX0 U5921_U2 ( .INP(WX8581), .ZN(U5921_n1) );
  NOR2X0 U5921_U1 ( .IN1(n10276), .IN2(U5921_n1), .QN(WX8644) );
  INVX0 U5922_U2 ( .INP(WX8579), .ZN(U5922_n1) );
  NOR2X0 U5922_U1 ( .IN1(n10276), .IN2(U5922_n1), .QN(WX8642) );
  INVX0 U5923_U2 ( .INP(WX8577), .ZN(U5923_n1) );
  NOR2X0 U5923_U1 ( .IN1(n10276), .IN2(U5923_n1), .QN(WX8640) );
  INVX0 U5924_U2 ( .INP(WX8575), .ZN(U5924_n1) );
  NOR2X0 U5924_U1 ( .IN1(n10276), .IN2(U5924_n1), .QN(WX8638) );
  INVX0 U5925_U2 ( .INP(WX8573), .ZN(U5925_n1) );
  NOR2X0 U5925_U1 ( .IN1(n10276), .IN2(U5925_n1), .QN(WX8636) );
  INVX0 U5926_U2 ( .INP(test_so73), .ZN(U5926_n1) );
  NOR2X0 U5926_U1 ( .IN1(n10276), .IN2(U5926_n1), .QN(WX8634) );
  INVX0 U5927_U2 ( .INP(WX8569), .ZN(U5927_n1) );
  NOR2X0 U5927_U1 ( .IN1(n10276), .IN2(U5927_n1), .QN(WX8632) );
  INVX0 U5928_U2 ( .INP(WX8567), .ZN(U5928_n1) );
  NOR2X0 U5928_U1 ( .IN1(n10276), .IN2(U5928_n1), .QN(WX8630) );
  INVX0 U5929_U2 ( .INP(WX8565), .ZN(U5929_n1) );
  NOR2X0 U5929_U1 ( .IN1(n10276), .IN2(U5929_n1), .QN(WX8628) );
  INVX0 U5930_U2 ( .INP(WX8563), .ZN(U5930_n1) );
  NOR2X0 U5930_U1 ( .IN1(n10276), .IN2(U5930_n1), .QN(WX8626) );
  INVX0 U5931_U2 ( .INP(WX8561), .ZN(U5931_n1) );
  NOR2X0 U5931_U1 ( .IN1(n10277), .IN2(U5931_n1), .QN(WX8624) );
  INVX0 U5932_U2 ( .INP(WX8559), .ZN(U5932_n1) );
  NOR2X0 U5932_U1 ( .IN1(n10277), .IN2(U5932_n1), .QN(WX8622) );
  INVX0 U5933_U2 ( .INP(WX8557), .ZN(U5933_n1) );
  NOR2X0 U5933_U1 ( .IN1(n10277), .IN2(U5933_n1), .QN(WX8620) );
  INVX0 U5934_U2 ( .INP(WX8555), .ZN(U5934_n1) );
  NOR2X0 U5934_U1 ( .IN1(n10277), .IN2(U5934_n1), .QN(WX8618) );
  INVX0 U5935_U2 ( .INP(WX8553), .ZN(U5935_n1) );
  NOR2X0 U5935_U1 ( .IN1(n10277), .IN2(U5935_n1), .QN(WX8616) );
  INVX0 U5936_U2 ( .INP(WX8551), .ZN(U5936_n1) );
  NOR2X0 U5936_U1 ( .IN1(n10277), .IN2(U5936_n1), .QN(WX8614) );
  INVX0 U5937_U2 ( .INP(WX8549), .ZN(U5937_n1) );
  NOR2X0 U5937_U1 ( .IN1(n10277), .IN2(U5937_n1), .QN(WX8612) );
  INVX0 U5938_U2 ( .INP(WX8547), .ZN(U5938_n1) );
  NOR2X0 U5938_U1 ( .IN1(n10277), .IN2(U5938_n1), .QN(WX8610) );
  INVX0 U5939_U2 ( .INP(WX8545), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n10277), .IN2(U5939_n1), .QN(WX8608) );
  INVX0 U5940_U2 ( .INP(WX8543), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n10304), .IN2(U5940_n1), .QN(WX8606) );
  INVX0 U5941_U2 ( .INP(WX8541), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n10298), .IN2(U5941_n1), .QN(WX8604) );
  INVX0 U5942_U2 ( .INP(WX8539), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n10298), .IN2(U5942_n1), .QN(WX8602) );
  INVX0 U5943_U2 ( .INP(test_so72), .ZN(U5943_n1) );
  NOR2X0 U5943_U1 ( .IN1(n10298), .IN2(U5943_n1), .QN(WX8600) );
  INVX0 U5944_U2 ( .INP(WX8535), .ZN(U5944_n1) );
  NOR2X0 U5944_U1 ( .IN1(n10298), .IN2(U5944_n1), .QN(WX8598) );
  INVX0 U5945_U2 ( .INP(WX8533), .ZN(U5945_n1) );
  NOR2X0 U5945_U1 ( .IN1(n10298), .IN2(U5945_n1), .QN(WX8596) );
  INVX0 U5946_U2 ( .INP(WX8531), .ZN(U5946_n1) );
  NOR2X0 U5946_U1 ( .IN1(n10299), .IN2(U5946_n1), .QN(WX8594) );
  INVX0 U5947_U2 ( .INP(WX8529), .ZN(U5947_n1) );
  NOR2X0 U5947_U1 ( .IN1(n10299), .IN2(U5947_n1), .QN(WX8592) );
  INVX0 U5948_U2 ( .INP(WX8527), .ZN(U5948_n1) );
  NOR2X0 U5948_U1 ( .IN1(n10299), .IN2(U5948_n1), .QN(WX8590) );
  INVX0 U5949_U2 ( .INP(WX8525), .ZN(U5949_n1) );
  NOR2X0 U5949_U1 ( .IN1(n10299), .IN2(U5949_n1), .QN(WX8588) );
  INVX0 U5950_U2 ( .INP(WX8523), .ZN(U5950_n1) );
  NOR2X0 U5950_U1 ( .IN1(n10299), .IN2(U5950_n1), .QN(WX8586) );
  INVX0 U5951_U2 ( .INP(WX8521), .ZN(U5951_n1) );
  NOR2X0 U5951_U1 ( .IN1(n10299), .IN2(U5951_n1), .QN(WX8584) );
  INVX0 U5952_U2 ( .INP(WX8519), .ZN(U5952_n1) );
  NOR2X0 U5952_U1 ( .IN1(n10299), .IN2(U5952_n1), .QN(WX8582) );
  INVX0 U5953_U2 ( .INP(WX8517), .ZN(U5953_n1) );
  NOR2X0 U5953_U1 ( .IN1(n10299), .IN2(U5953_n1), .QN(WX8580) );
  INVX0 U5954_U2 ( .INP(WX8515), .ZN(U5954_n1) );
  NOR2X0 U5954_U1 ( .IN1(n10299), .IN2(U5954_n1), .QN(WX8578) );
  INVX0 U5955_U2 ( .INP(WX8513), .ZN(U5955_n1) );
  NOR2X0 U5955_U1 ( .IN1(n10299), .IN2(U5955_n1), .QN(WX8576) );
  INVX0 U5956_U2 ( .INP(WX8511), .ZN(U5956_n1) );
  NOR2X0 U5956_U1 ( .IN1(n10299), .IN2(U5956_n1), .QN(WX8574) );
  INVX0 U5957_U2 ( .INP(WX8509), .ZN(U5957_n1) );
  NOR2X0 U5957_U1 ( .IN1(n10300), .IN2(U5957_n1), .QN(WX8572) );
  INVX0 U5958_U2 ( .INP(WX8507), .ZN(U5958_n1) );
  NOR2X0 U5958_U1 ( .IN1(n10300), .IN2(U5958_n1), .QN(WX8570) );
  INVX0 U5959_U2 ( .INP(WX8505), .ZN(U5959_n1) );
  NOR2X0 U5959_U1 ( .IN1(n10300), .IN2(U5959_n1), .QN(WX8568) );
  INVX0 U5960_U2 ( .INP(test_so71), .ZN(U5960_n1) );
  NOR2X0 U5960_U1 ( .IN1(n10300), .IN2(U5960_n1), .QN(WX8566) );
  INVX0 U5961_U2 ( .INP(WX8501), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n10300), .IN2(U5961_n1), .QN(WX8564) );
  INVX0 U5962_U2 ( .INP(WX8499), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n10300), .IN2(U5962_n1), .QN(WX8562) );
  INVX0 U5963_U2 ( .INP(WX8497), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n10300), .IN2(U5963_n1), .QN(WX8560) );
  INVX0 U5964_U2 ( .INP(WX8495), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n10300), .IN2(U5964_n1), .QN(WX8558) );
  INVX0 U5965_U2 ( .INP(WX8493), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n10300), .IN2(U5965_n1), .QN(WX8556) );
  INVX0 U5966_U2 ( .INP(WX8491), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n10300), .IN2(U5966_n1), .QN(WX8554) );
  INVX0 U5967_U2 ( .INP(WX8489), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n10300), .IN2(U5967_n1), .QN(WX8552) );
  INVX0 U5968_U2 ( .INP(WX8487), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n10301), .IN2(U5968_n1), .QN(WX8550) );
  INVX0 U5969_U2 ( .INP(WX8485), .ZN(U5969_n1) );
  NOR2X0 U5969_U1 ( .IN1(n10301), .IN2(U5969_n1), .QN(WX8548) );
  INVX0 U5970_U2 ( .INP(WX8483), .ZN(U5970_n1) );
  NOR2X0 U5970_U1 ( .IN1(n10301), .IN2(U5970_n1), .QN(WX8546) );
  INVX0 U5971_U2 ( .INP(WX8481), .ZN(U5971_n1) );
  NOR2X0 U5971_U1 ( .IN1(n10301), .IN2(U5971_n1), .QN(WX8544) );
  INVX0 U5972_U2 ( .INP(WX8479), .ZN(U5972_n1) );
  NOR2X0 U5972_U1 ( .IN1(n10301), .IN2(U5972_n1), .QN(WX8542) );
  INVX0 U5973_U2 ( .INP(WX8477), .ZN(U5973_n1) );
  NOR2X0 U5973_U1 ( .IN1(n10301), .IN2(U5973_n1), .QN(WX8540) );
  INVX0 U5974_U2 ( .INP(WX8475), .ZN(U5974_n1) );
  NOR2X0 U5974_U1 ( .IN1(n10301), .IN2(U5974_n1), .QN(WX8538) );
  INVX0 U5975_U2 ( .INP(WX8473), .ZN(U5975_n1) );
  NOR2X0 U5975_U1 ( .IN1(n10301), .IN2(U5975_n1), .QN(WX8536) );
  INVX0 U5976_U2 ( .INP(WX8471), .ZN(U5976_n1) );
  NOR2X0 U5976_U1 ( .IN1(n10301), .IN2(U5976_n1), .QN(WX8534) );
  INVX0 U5977_U2 ( .INP(test_so70), .ZN(U5977_n1) );
  NOR2X0 U5977_U1 ( .IN1(n10301), .IN2(U5977_n1), .QN(WX8532) );
  INVX0 U5978_U2 ( .INP(WX8467), .ZN(U5978_n1) );
  NOR2X0 U5978_U1 ( .IN1(n10301), .IN2(U5978_n1), .QN(WX8530) );
  INVX0 U5979_U2 ( .INP(WX8465), .ZN(U5979_n1) );
  NOR2X0 U5979_U1 ( .IN1(n10302), .IN2(U5979_n1), .QN(WX8528) );
  INVX0 U5980_U2 ( .INP(WX8463), .ZN(U5980_n1) );
  NOR2X0 U5980_U1 ( .IN1(n10302), .IN2(U5980_n1), .QN(WX8526) );
  INVX0 U5981_U2 ( .INP(WX8461), .ZN(U5981_n1) );
  NOR2X0 U5981_U1 ( .IN1(n10302), .IN2(U5981_n1), .QN(WX8524) );
  INVX0 U5982_U2 ( .INP(WX8459), .ZN(U5982_n1) );
  NOR2X0 U5982_U1 ( .IN1(n10302), .IN2(U5982_n1), .QN(WX8522) );
  INVX0 U5983_U2 ( .INP(WX8457), .ZN(U5983_n1) );
  NOR2X0 U5983_U1 ( .IN1(n10302), .IN2(U5983_n1), .QN(WX8520) );
  INVX0 U5984_U2 ( .INP(WX8455), .ZN(U5984_n1) );
  NOR2X0 U5984_U1 ( .IN1(n10302), .IN2(U5984_n1), .QN(WX8518) );
  INVX0 U5985_U2 ( .INP(WX8453), .ZN(U5985_n1) );
  NOR2X0 U5985_U1 ( .IN1(n10302), .IN2(U5985_n1), .QN(WX8516) );
  INVX0 U5986_U2 ( .INP(WX8451), .ZN(U5986_n1) );
  NOR2X0 U5986_U1 ( .IN1(n10302), .IN2(U5986_n1), .QN(WX8514) );
  INVX0 U5987_U2 ( .INP(WX8449), .ZN(U5987_n1) );
  NOR2X0 U5987_U1 ( .IN1(n10302), .IN2(U5987_n1), .QN(WX8512) );
  INVX0 U5988_U2 ( .INP(WX8447), .ZN(U5988_n1) );
  NOR2X0 U5988_U1 ( .IN1(n10302), .IN2(U5988_n1), .QN(WX8510) );
  INVX0 U5989_U2 ( .INP(WX8445), .ZN(U5989_n1) );
  NOR2X0 U5989_U1 ( .IN1(n10302), .IN2(U5989_n1), .QN(WX8508) );
  INVX0 U5990_U2 ( .INP(WX8443), .ZN(U5990_n1) );
  NOR2X0 U5990_U1 ( .IN1(n10303), .IN2(U5990_n1), .QN(WX8506) );
  INVX0 U5991_U2 ( .INP(WX8441), .ZN(U5991_n1) );
  NOR2X0 U5991_U1 ( .IN1(n10303), .IN2(U5991_n1), .QN(WX8504) );
  INVX0 U5992_U2 ( .INP(WX8439), .ZN(U5992_n1) );
  NOR2X0 U5992_U1 ( .IN1(n10303), .IN2(U5992_n1), .QN(WX8502) );
  INVX0 U5993_U2 ( .INP(WX8437), .ZN(U5993_n1) );
  NOR2X0 U5993_U1 ( .IN1(n10303), .IN2(U5993_n1), .QN(WX8500) );
  INVX0 U5994_U2 ( .INP(test_so69), .ZN(U5994_n1) );
  NOR2X0 U5994_U1 ( .IN1(n10303), .IN2(U5994_n1), .QN(WX8498) );
  INVX0 U5995_U2 ( .INP(WX7300), .ZN(U5995_n1) );
  NOR2X0 U5995_U1 ( .IN1(n10303), .IN2(U5995_n1), .QN(WX7363) );
  INVX0 U5996_U2 ( .INP(WX7298), .ZN(U5996_n1) );
  NOR2X0 U5996_U1 ( .IN1(n10303), .IN2(U5996_n1), .QN(WX7361) );
  INVX0 U5997_U2 ( .INP(WX7296), .ZN(U5997_n1) );
  NOR2X0 U5997_U1 ( .IN1(n10303), .IN2(U5997_n1), .QN(WX7359) );
  INVX0 U5998_U2 ( .INP(WX7294), .ZN(U5998_n1) );
  NOR2X0 U5998_U1 ( .IN1(n10303), .IN2(U5998_n1), .QN(WX7357) );
  INVX0 U5999_U2 ( .INP(WX7292), .ZN(U5999_n1) );
  NOR2X0 U5999_U1 ( .IN1(n10303), .IN2(U5999_n1), .QN(WX7355) );
  INVX0 U6000_U2 ( .INP(WX7290), .ZN(U6000_n1) );
  NOR2X0 U6000_U1 ( .IN1(n10303), .IN2(U6000_n1), .QN(WX7353) );
  INVX0 U6001_U2 ( .INP(test_so62), .ZN(U6001_n1) );
  NOR2X0 U6001_U1 ( .IN1(n10304), .IN2(U6001_n1), .QN(WX7351) );
  INVX0 U6002_U2 ( .INP(WX7286), .ZN(U6002_n1) );
  NOR2X0 U6002_U1 ( .IN1(n10304), .IN2(U6002_n1), .QN(WX7349) );
  INVX0 U6003_U2 ( .INP(WX7284), .ZN(U6003_n1) );
  NOR2X0 U6003_U1 ( .IN1(n10304), .IN2(U6003_n1), .QN(WX7347) );
  INVX0 U6004_U2 ( .INP(WX7282), .ZN(U6004_n1) );
  NOR2X0 U6004_U1 ( .IN1(n10304), .IN2(U6004_n1), .QN(WX7345) );
  INVX0 U6005_U2 ( .INP(WX7280), .ZN(U6005_n1) );
  NOR2X0 U6005_U1 ( .IN1(n10304), .IN2(U6005_n1), .QN(WX7343) );
  INVX0 U6006_U2 ( .INP(WX7278), .ZN(U6006_n1) );
  NOR2X0 U6006_U1 ( .IN1(n10304), .IN2(U6006_n1), .QN(WX7341) );
  INVX0 U6007_U2 ( .INP(WX7276), .ZN(U6007_n1) );
  NOR2X0 U6007_U1 ( .IN1(n10304), .IN2(U6007_n1), .QN(WX7339) );
  INVX0 U6008_U2 ( .INP(WX7274), .ZN(U6008_n1) );
  NOR2X0 U6008_U1 ( .IN1(n10305), .IN2(U6008_n1), .QN(WX7337) );
  INVX0 U6009_U2 ( .INP(WX7272), .ZN(U6009_n1) );
  NOR2X0 U6009_U1 ( .IN1(n10304), .IN2(U6009_n1), .QN(WX7335) );
  INVX0 U6010_U2 ( .INP(WX7270), .ZN(U6010_n1) );
  NOR2X0 U6010_U1 ( .IN1(n10306), .IN2(U6010_n1), .QN(WX7333) );
  INVX0 U6011_U2 ( .INP(WX7268), .ZN(U6011_n1) );
  NOR2X0 U6011_U1 ( .IN1(n10305), .IN2(U6011_n1), .QN(WX7331) );
  INVX0 U6012_U2 ( .INP(WX7266), .ZN(U6012_n1) );
  NOR2X0 U6012_U1 ( .IN1(n10306), .IN2(U6012_n1), .QN(WX7329) );
  INVX0 U6013_U2 ( .INP(WX7264), .ZN(U6013_n1) );
  NOR2X0 U6013_U1 ( .IN1(n10306), .IN2(U6013_n1), .QN(WX7327) );
  INVX0 U6014_U2 ( .INP(WX7262), .ZN(U6014_n1) );
  NOR2X0 U6014_U1 ( .IN1(n10304), .IN2(U6014_n1), .QN(WX7325) );
  INVX0 U6015_U2 ( .INP(WX7260), .ZN(U6015_n1) );
  NOR2X0 U6015_U1 ( .IN1(n10306), .IN2(U6015_n1), .QN(WX7323) );
  INVX0 U6016_U2 ( .INP(WX7258), .ZN(U6016_n1) );
  NOR2X0 U6016_U1 ( .IN1(n10306), .IN2(U6016_n1), .QN(WX7321) );
  INVX0 U6017_U2 ( .INP(WX7256), .ZN(U6017_n1) );
  NOR2X0 U6017_U1 ( .IN1(n10305), .IN2(U6017_n1), .QN(WX7319) );
  INVX0 U6018_U2 ( .INP(test_so61), .ZN(U6018_n1) );
  NOR2X0 U6018_U1 ( .IN1(n10306), .IN2(U6018_n1), .QN(WX7317) );
  INVX0 U6019_U2 ( .INP(WX7252), .ZN(U6019_n1) );
  NOR2X0 U6019_U1 ( .IN1(n10307), .IN2(U6019_n1), .QN(WX7315) );
  INVX0 U6020_U2 ( .INP(WX7250), .ZN(U6020_n1) );
  NOR2X0 U6020_U1 ( .IN1(n10305), .IN2(U6020_n1), .QN(WX7313) );
  INVX0 U6021_U2 ( .INP(WX7248), .ZN(U6021_n1) );
  NOR2X0 U6021_U1 ( .IN1(n10305), .IN2(U6021_n1), .QN(WX7311) );
  INVX0 U6022_U2 ( .INP(WX7246), .ZN(U6022_n1) );
  NOR2X0 U6022_U1 ( .IN1(n10304), .IN2(U6022_n1), .QN(WX7309) );
  INVX0 U6023_U2 ( .INP(WX7244), .ZN(U6023_n1) );
  NOR2X0 U6023_U1 ( .IN1(n10305), .IN2(U6023_n1), .QN(WX7307) );
  INVX0 U6024_U2 ( .INP(WX7242), .ZN(U6024_n1) );
  NOR2X0 U6024_U1 ( .IN1(n10307), .IN2(U6024_n1), .QN(WX7305) );
  INVX0 U6025_U2 ( .INP(WX7240), .ZN(U6025_n1) );
  NOR2X0 U6025_U1 ( .IN1(n10307), .IN2(U6025_n1), .QN(WX7303) );
  INVX0 U6026_U2 ( .INP(WX7238), .ZN(U6026_n1) );
  NOR2X0 U6026_U1 ( .IN1(n10305), .IN2(U6026_n1), .QN(WX7301) );
  INVX0 U6027_U2 ( .INP(WX7236), .ZN(U6027_n1) );
  NOR2X0 U6027_U1 ( .IN1(n10307), .IN2(U6027_n1), .QN(WX7299) );
  INVX0 U6028_U2 ( .INP(WX7234), .ZN(U6028_n1) );
  NOR2X0 U6028_U1 ( .IN1(n10305), .IN2(U6028_n1), .QN(WX7297) );
  INVX0 U6029_U2 ( .INP(WX7232), .ZN(U6029_n1) );
  NOR2X0 U6029_U1 ( .IN1(n10305), .IN2(U6029_n1), .QN(WX7295) );
  INVX0 U6030_U2 ( .INP(WX7230), .ZN(U6030_n1) );
  NOR2X0 U6030_U1 ( .IN1(n10307), .IN2(U6030_n1), .QN(WX7293) );
  INVX0 U6031_U2 ( .INP(WX7228), .ZN(U6031_n1) );
  NOR2X0 U6031_U1 ( .IN1(n10307), .IN2(U6031_n1), .QN(WX7291) );
  INVX0 U6032_U2 ( .INP(WX7226), .ZN(U6032_n1) );
  NOR2X0 U6032_U1 ( .IN1(n10306), .IN2(U6032_n1), .QN(WX7289) );
  INVX0 U6033_U2 ( .INP(WX7224), .ZN(U6033_n1) );
  NOR2X0 U6033_U1 ( .IN1(n10307), .IN2(U6033_n1), .QN(WX7287) );
  INVX0 U6034_U2 ( .INP(WX7222), .ZN(U6034_n1) );
  NOR2X0 U6034_U1 ( .IN1(n10307), .IN2(U6034_n1), .QN(WX7285) );
  INVX0 U6035_U2 ( .INP(test_so60), .ZN(U6035_n1) );
  NOR2X0 U6035_U1 ( .IN1(n10305), .IN2(U6035_n1), .QN(WX7283) );
  INVX0 U6036_U2 ( .INP(WX7218), .ZN(U6036_n1) );
  NOR2X0 U6036_U1 ( .IN1(n10307), .IN2(U6036_n1), .QN(WX7281) );
  INVX0 U6037_U2 ( .INP(WX7216), .ZN(U6037_n1) );
  NOR2X0 U6037_U1 ( .IN1(n10307), .IN2(U6037_n1), .QN(WX7279) );
  INVX0 U6038_U2 ( .INP(WX7214), .ZN(U6038_n1) );
  NOR2X0 U6038_U1 ( .IN1(n10306), .IN2(U6038_n1), .QN(WX7277) );
  INVX0 U6039_U2 ( .INP(WX7212), .ZN(U6039_n1) );
  NOR2X0 U6039_U1 ( .IN1(n10306), .IN2(U6039_n1), .QN(WX7275) );
  INVX0 U6040_U2 ( .INP(WX7210), .ZN(U6040_n1) );
  NOR2X0 U6040_U1 ( .IN1(n10288), .IN2(U6040_n1), .QN(WX7273) );
  INVX0 U6041_U2 ( .INP(WX7208), .ZN(U6041_n1) );
  NOR2X0 U6041_U1 ( .IN1(n10289), .IN2(U6041_n1), .QN(WX7271) );
  INVX0 U6042_U2 ( .INP(WX7206), .ZN(U6042_n1) );
  NOR2X0 U6042_U1 ( .IN1(n10289), .IN2(U6042_n1), .QN(WX7269) );
  INVX0 U6043_U2 ( .INP(WX7204), .ZN(U6043_n1) );
  NOR2X0 U6043_U1 ( .IN1(n10289), .IN2(U6043_n1), .QN(WX7267) );
  INVX0 U6044_U2 ( .INP(WX7202), .ZN(U6044_n1) );
  NOR2X0 U6044_U1 ( .IN1(n10289), .IN2(U6044_n1), .QN(WX7265) );
  INVX0 U6045_U2 ( .INP(WX7200), .ZN(U6045_n1) );
  NOR2X0 U6045_U1 ( .IN1(n10289), .IN2(U6045_n1), .QN(WX7263) );
  INVX0 U6046_U2 ( .INP(WX7198), .ZN(U6046_n1) );
  NOR2X0 U6046_U1 ( .IN1(n10289), .IN2(U6046_n1), .QN(WX7261) );
  INVX0 U6047_U2 ( .INP(WX7196), .ZN(U6047_n1) );
  NOR2X0 U6047_U1 ( .IN1(n10289), .IN2(U6047_n1), .QN(WX7259) );
  INVX0 U6048_U2 ( .INP(WX7194), .ZN(U6048_n1) );
  NOR2X0 U6048_U1 ( .IN1(n10290), .IN2(U6048_n1), .QN(WX7257) );
  INVX0 U6049_U2 ( .INP(WX7192), .ZN(U6049_n1) );
  NOR2X0 U6049_U1 ( .IN1(n10290), .IN2(U6049_n1), .QN(WX7255) );
  INVX0 U6050_U2 ( .INP(WX7190), .ZN(U6050_n1) );
  NOR2X0 U6050_U1 ( .IN1(n10290), .IN2(U6050_n1), .QN(WX7253) );
  INVX0 U6051_U2 ( .INP(WX7188), .ZN(U6051_n1) );
  NOR2X0 U6051_U1 ( .IN1(n10290), .IN2(U6051_n1), .QN(WX7251) );
  INVX0 U6052_U2 ( .INP(test_so59), .ZN(U6052_n1) );
  NOR2X0 U6052_U1 ( .IN1(n10290), .IN2(U6052_n1), .QN(WX7249) );
  INVX0 U6053_U2 ( .INP(WX7184), .ZN(U6053_n1) );
  NOR2X0 U6053_U1 ( .IN1(n10290), .IN2(U6053_n1), .QN(WX7247) );
  INVX0 U6054_U2 ( .INP(WX7182), .ZN(U6054_n1) );
  NOR2X0 U6054_U1 ( .IN1(n10290), .IN2(U6054_n1), .QN(WX7245) );
  INVX0 U6055_U2 ( .INP(WX7180), .ZN(U6055_n1) );
  NOR2X0 U6055_U1 ( .IN1(n10290), .IN2(U6055_n1), .QN(WX7243) );
  INVX0 U6056_U2 ( .INP(WX7178), .ZN(U6056_n1) );
  NOR2X0 U6056_U1 ( .IN1(n10290), .IN2(U6056_n1), .QN(WX7241) );
  INVX0 U6057_U2 ( .INP(WX7176), .ZN(U6057_n1) );
  NOR2X0 U6057_U1 ( .IN1(n10291), .IN2(U6057_n1), .QN(WX7239) );
  INVX0 U6058_U2 ( .INP(WX7174), .ZN(U6058_n1) );
  NOR2X0 U6058_U1 ( .IN1(n10291), .IN2(U6058_n1), .QN(WX7237) );
  INVX0 U6059_U2 ( .INP(WX7172), .ZN(U6059_n1) );
  NOR2X0 U6059_U1 ( .IN1(n10291), .IN2(U6059_n1), .QN(WX7235) );
  INVX0 U6060_U2 ( .INP(WX7170), .ZN(U6060_n1) );
  NOR2X0 U6060_U1 ( .IN1(n10291), .IN2(U6060_n1), .QN(WX7233) );
  INVX0 U6061_U2 ( .INP(WX7168), .ZN(U6061_n1) );
  NOR2X0 U6061_U1 ( .IN1(n10291), .IN2(U6061_n1), .QN(WX7231) );
  INVX0 U6062_U2 ( .INP(WX7166), .ZN(U6062_n1) );
  NOR2X0 U6062_U1 ( .IN1(n10291), .IN2(U6062_n1), .QN(WX7229) );
  INVX0 U6063_U2 ( .INP(WX7164), .ZN(U6063_n1) );
  NOR2X0 U6063_U1 ( .IN1(n10291), .IN2(U6063_n1), .QN(WX7227) );
  INVX0 U6064_U2 ( .INP(WX7162), .ZN(U6064_n1) );
  NOR2X0 U6064_U1 ( .IN1(n10291), .IN2(U6064_n1), .QN(WX7225) );
  INVX0 U6065_U2 ( .INP(WX7160), .ZN(U6065_n1) );
  NOR2X0 U6065_U1 ( .IN1(n10291), .IN2(U6065_n1), .QN(WX7223) );
  INVX0 U6066_U2 ( .INP(WX7158), .ZN(U6066_n1) );
  NOR2X0 U6066_U1 ( .IN1(n10291), .IN2(U6066_n1), .QN(WX7221) );
  INVX0 U6067_U2 ( .INP(WX7156), .ZN(U6067_n1) );
  NOR2X0 U6067_U1 ( .IN1(n10292), .IN2(U6067_n1), .QN(WX7219) );
  INVX0 U6068_U2 ( .INP(WX7154), .ZN(U6068_n1) );
  NOR2X0 U6068_U1 ( .IN1(n10292), .IN2(U6068_n1), .QN(WX7217) );
  INVX0 U6069_U2 ( .INP(test_so58), .ZN(U6069_n1) );
  NOR2X0 U6069_U1 ( .IN1(n10292), .IN2(U6069_n1), .QN(WX7215) );
  INVX0 U6070_U2 ( .INP(WX7150), .ZN(U6070_n1) );
  NOR2X0 U6070_U1 ( .IN1(n10292), .IN2(U6070_n1), .QN(WX7213) );
  INVX0 U6071_U2 ( .INP(WX7148), .ZN(U6071_n1) );
  NOR2X0 U6071_U1 ( .IN1(n10292), .IN2(U6071_n1), .QN(WX7211) );
  INVX0 U6072_U2 ( .INP(WX7146), .ZN(U6072_n1) );
  NOR2X0 U6072_U1 ( .IN1(n10292), .IN2(U6072_n1), .QN(WX7209) );
  INVX0 U6073_U2 ( .INP(WX7144), .ZN(U6073_n1) );
  NOR2X0 U6073_U1 ( .IN1(n10293), .IN2(U6073_n1), .QN(WX7207) );
  INVX0 U6074_U2 ( .INP(WX7142), .ZN(U6074_n1) );
  NOR2X0 U6074_U1 ( .IN1(n10293), .IN2(U6074_n1), .QN(WX7205) );
  INVX0 U6075_U2 ( .INP(WX6007), .ZN(U6075_n1) );
  NOR2X0 U6075_U1 ( .IN1(n10293), .IN2(U6075_n1), .QN(WX6070) );
  INVX0 U6076_U2 ( .INP(test_so51), .ZN(U6076_n1) );
  NOR2X0 U6076_U1 ( .IN1(n10293), .IN2(U6076_n1), .QN(WX6068) );
  INVX0 U6077_U2 ( .INP(WX6003), .ZN(U6077_n1) );
  NOR2X0 U6077_U1 ( .IN1(n10293), .IN2(U6077_n1), .QN(WX6066) );
  INVX0 U6078_U2 ( .INP(WX6001), .ZN(U6078_n1) );
  NOR2X0 U6078_U1 ( .IN1(n10293), .IN2(U6078_n1), .QN(WX6064) );
  INVX0 U6079_U2 ( .INP(WX5999), .ZN(U6079_n1) );
  NOR2X0 U6079_U1 ( .IN1(n10293), .IN2(U6079_n1), .QN(WX6062) );
  INVX0 U6080_U2 ( .INP(WX5997), .ZN(U6080_n1) );
  NOR2X0 U6080_U1 ( .IN1(n10293), .IN2(U6080_n1), .QN(WX6060) );
  INVX0 U6081_U2 ( .INP(WX5995), .ZN(U6081_n1) );
  NOR2X0 U6081_U1 ( .IN1(n10293), .IN2(U6081_n1), .QN(WX6058) );
  INVX0 U6082_U2 ( .INP(WX5993), .ZN(U6082_n1) );
  NOR2X0 U6082_U1 ( .IN1(n10293), .IN2(U6082_n1), .QN(WX6056) );
  INVX0 U6083_U2 ( .INP(WX5991), .ZN(U6083_n1) );
  NOR2X0 U6083_U1 ( .IN1(n10294), .IN2(U6083_n1), .QN(WX6054) );
  INVX0 U6084_U2 ( .INP(WX5989), .ZN(U6084_n1) );
  NOR2X0 U6084_U1 ( .IN1(n10294), .IN2(U6084_n1), .QN(WX6052) );
  INVX0 U6085_U2 ( .INP(WX5987), .ZN(U6085_n1) );
  NOR2X0 U6085_U1 ( .IN1(n10294), .IN2(U6085_n1), .QN(WX6050) );
  INVX0 U6086_U2 ( .INP(WX5985), .ZN(U6086_n1) );
  NOR2X0 U6086_U1 ( .IN1(n10294), .IN2(U6086_n1), .QN(WX6048) );
  INVX0 U6087_U2 ( .INP(WX5983), .ZN(U6087_n1) );
  NOR2X0 U6087_U1 ( .IN1(n10295), .IN2(U6087_n1), .QN(WX6046) );
  INVX0 U6088_U2 ( .INP(WX5981), .ZN(U6088_n1) );
  NOR2X0 U6088_U1 ( .IN1(n10295), .IN2(U6088_n1), .QN(WX6044) );
  INVX0 U6089_U2 ( .INP(WX5979), .ZN(U6089_n1) );
  NOR2X0 U6089_U1 ( .IN1(n10295), .IN2(U6089_n1), .QN(WX6042) );
  INVX0 U6090_U2 ( .INP(WX5977), .ZN(U6090_n1) );
  NOR2X0 U6090_U1 ( .IN1(n10295), .IN2(U6090_n1), .QN(WX6040) );
  INVX0 U6091_U2 ( .INP(WX5975), .ZN(U6091_n1) );
  NOR2X0 U6091_U1 ( .IN1(n10298), .IN2(U6091_n1), .QN(WX6038) );
  INVX0 U6092_U2 ( .INP(WX5973), .ZN(U6092_n1) );
  NOR2X0 U6092_U1 ( .IN1(n10295), .IN2(U6092_n1), .QN(WX6036) );
  INVX0 U6093_U2 ( .INP(test_so50), .ZN(U6093_n1) );
  NOR2X0 U6093_U1 ( .IN1(n10295), .IN2(U6093_n1), .QN(WX6034) );
  INVX0 U6094_U2 ( .INP(WX5969), .ZN(U6094_n1) );
  NOR2X0 U6094_U1 ( .IN1(n10295), .IN2(U6094_n1), .QN(WX6032) );
  INVX0 U6095_U2 ( .INP(WX5967), .ZN(U6095_n1) );
  NOR2X0 U6095_U1 ( .IN1(n10295), .IN2(U6095_n1), .QN(WX6030) );
  INVX0 U6096_U2 ( .INP(WX5965), .ZN(U6096_n1) );
  NOR2X0 U6096_U1 ( .IN1(n10296), .IN2(U6096_n1), .QN(WX6028) );
  INVX0 U6097_U2 ( .INP(WX5963), .ZN(U6097_n1) );
  NOR2X0 U6097_U1 ( .IN1(n10296), .IN2(U6097_n1), .QN(WX6026) );
  INVX0 U6098_U2 ( .INP(WX5961), .ZN(U6098_n1) );
  NOR2X0 U6098_U1 ( .IN1(n10296), .IN2(U6098_n1), .QN(WX6024) );
  INVX0 U6099_U2 ( .INP(WX5959), .ZN(U6099_n1) );
  NOR2X0 U6099_U1 ( .IN1(n10296), .IN2(U6099_n1), .QN(WX6022) );
  INVX0 U6100_U2 ( .INP(WX5957), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n10296), .IN2(U6100_n1), .QN(WX6020) );
  INVX0 U6101_U2 ( .INP(WX5955), .ZN(U6101_n1) );
  NOR2X0 U6101_U1 ( .IN1(n10296), .IN2(U6101_n1), .QN(WX6018) );
  INVX0 U6102_U2 ( .INP(WX5953), .ZN(U6102_n1) );
  NOR2X0 U6102_U1 ( .IN1(n10298), .IN2(U6102_n1), .QN(WX6016) );
  INVX0 U6103_U2 ( .INP(WX5951), .ZN(U6103_n1) );
  NOR2X0 U6103_U1 ( .IN1(n10298), .IN2(U6103_n1), .QN(WX6014) );
  INVX0 U6104_U2 ( .INP(WX5949), .ZN(U6104_n1) );
  NOR2X0 U6104_U1 ( .IN1(n10298), .IN2(U6104_n1), .QN(WX6012) );
  INVX0 U6105_U2 ( .INP(WX5947), .ZN(U6105_n1) );
  NOR2X0 U6105_U1 ( .IN1(n10298), .IN2(U6105_n1), .QN(WX6010) );
  INVX0 U6106_U2 ( .INP(WX5945), .ZN(U6106_n1) );
  NOR2X0 U6106_U1 ( .IN1(n10295), .IN2(U6106_n1), .QN(WX6008) );
  INVX0 U6107_U2 ( .INP(WX5943), .ZN(U6107_n1) );
  NOR2X0 U6107_U1 ( .IN1(n10298), .IN2(U6107_n1), .QN(WX6006) );
  INVX0 U6108_U2 ( .INP(WX5941), .ZN(U6108_n1) );
  NOR2X0 U6108_U1 ( .IN1(n10297), .IN2(U6108_n1), .QN(WX6004) );
  INVX0 U6109_U2 ( .INP(WX5929), .ZN(U6109_n1) );
  NOR2X0 U6109_U1 ( .IN1(n10297), .IN2(U6109_n1), .QN(WX5992) );
  INVX0 U6110_U2 ( .INP(WX5927), .ZN(U6110_n1) );
  NOR2X0 U6110_U1 ( .IN1(n10297), .IN2(U6110_n1), .QN(WX5990) );
  INVX0 U6111_U2 ( .INP(WX5925), .ZN(U6111_n1) );
  NOR2X0 U6111_U1 ( .IN1(n10297), .IN2(U6111_n1), .QN(WX5988) );
  INVX0 U6112_U2 ( .INP(WX5923), .ZN(U6112_n1) );
  NOR2X0 U6112_U1 ( .IN1(n10297), .IN2(U6112_n1), .QN(WX5986) );
  INVX0 U6113_U2 ( .INP(WX5921), .ZN(U6113_n1) );
  NOR2X0 U6113_U1 ( .IN1(n10297), .IN2(U6113_n1), .QN(WX5984) );
  INVX0 U6114_U2 ( .INP(WX5919), .ZN(U6114_n1) );
  NOR2X0 U6114_U1 ( .IN1(n10297), .IN2(U6114_n1), .QN(WX5982) );
  INVX0 U6115_U2 ( .INP(WX5917), .ZN(U6115_n1) );
  NOR2X0 U6115_U1 ( .IN1(n10297), .IN2(U6115_n1), .QN(WX5980) );
  INVX0 U6116_U2 ( .INP(WX5915), .ZN(U6116_n1) );
  NOR2X0 U6116_U1 ( .IN1(n10297), .IN2(U6116_n1), .QN(WX5978) );
  INVX0 U6117_U2 ( .INP(WX5913), .ZN(U6117_n1) );
  NOR2X0 U6117_U1 ( .IN1(n10297), .IN2(U6117_n1), .QN(WX5976) );
  INVX0 U6118_U2 ( .INP(WX5911), .ZN(U6118_n1) );
  NOR2X0 U6118_U1 ( .IN1(n10297), .IN2(U6118_n1), .QN(WX5974) );
  INVX0 U6119_U2 ( .INP(WX5909), .ZN(U6119_n1) );
  NOR2X0 U6119_U1 ( .IN1(n10296), .IN2(U6119_n1), .QN(WX5972) );
  INVX0 U6120_U2 ( .INP(WX5907), .ZN(U6120_n1) );
  NOR2X0 U6120_U1 ( .IN1(n10296), .IN2(U6120_n1), .QN(WX5970) );
  INVX0 U6121_U2 ( .INP(WX5905), .ZN(U6121_n1) );
  NOR2X0 U6121_U1 ( .IN1(n10296), .IN2(U6121_n1), .QN(WX5968) );
  INVX0 U6122_U2 ( .INP(test_so48), .ZN(U6122_n1) );
  NOR2X0 U6122_U1 ( .IN1(n10296), .IN2(U6122_n1), .QN(WX5966) );
  INVX0 U6123_U2 ( .INP(WX5901), .ZN(U6123_n1) );
  NOR2X0 U6123_U1 ( .IN1(n10296), .IN2(U6123_n1), .QN(WX5964) );
  INVX0 U6124_U2 ( .INP(WX5899), .ZN(U6124_n1) );
  NOR2X0 U6124_U1 ( .IN1(n10295), .IN2(U6124_n1), .QN(WX5962) );
  INVX0 U6125_U2 ( .INP(WX5897), .ZN(U6125_n1) );
  NOR2X0 U6125_U1 ( .IN1(n10295), .IN2(U6125_n1), .QN(WX5960) );
  INVX0 U6126_U2 ( .INP(WX5895), .ZN(U6126_n1) );
  NOR2X0 U6126_U1 ( .IN1(n10294), .IN2(U6126_n1), .QN(WX5958) );
  INVX0 U6127_U2 ( .INP(WX5893), .ZN(U6127_n1) );
  NOR2X0 U6127_U1 ( .IN1(n10294), .IN2(U6127_n1), .QN(WX5956) );
  INVX0 U6128_U2 ( .INP(WX5891), .ZN(U6128_n1) );
  NOR2X0 U6128_U1 ( .IN1(n10294), .IN2(U6128_n1), .QN(WX5954) );
  INVX0 U6129_U2 ( .INP(WX5889), .ZN(U6129_n1) );
  NOR2X0 U6129_U1 ( .IN1(n10294), .IN2(U6129_n1), .QN(WX5952) );
  INVX0 U6130_U2 ( .INP(WX5887), .ZN(U6130_n1) );
  NOR2X0 U6130_U1 ( .IN1(n10294), .IN2(U6130_n1), .QN(WX5950) );
  INVX0 U6131_U2 ( .INP(WX5885), .ZN(U6131_n1) );
  NOR2X0 U6131_U1 ( .IN1(n10294), .IN2(U6131_n1), .QN(WX5948) );
  INVX0 U6132_U2 ( .INP(WX5883), .ZN(U6132_n1) );
  NOR2X0 U6132_U1 ( .IN1(n10294), .IN2(U6132_n1), .QN(WX5946) );
  INVX0 U6133_U2 ( .INP(WX5881), .ZN(U6133_n1) );
  NOR2X0 U6133_U1 ( .IN1(n10292), .IN2(U6133_n1), .QN(WX5944) );
  INVX0 U6134_U2 ( .INP(WX5879), .ZN(U6134_n1) );
  NOR2X0 U6134_U1 ( .IN1(n10292), .IN2(U6134_n1), .QN(WX5942) );
  INVX0 U6135_U2 ( .INP(WX5877), .ZN(U6135_n1) );
  NOR2X0 U6135_U1 ( .IN1(n10292), .IN2(U6135_n1), .QN(WX5940) );
  INVX0 U6136_U2 ( .INP(WX5875), .ZN(U6136_n1) );
  NOR2X0 U6136_U1 ( .IN1(n10292), .IN2(U6136_n1), .QN(WX5938) );
  INVX0 U6137_U2 ( .INP(WX5873), .ZN(U6137_n1) );
  NOR2X0 U6137_U1 ( .IN1(n10292), .IN2(U6137_n1), .QN(WX5936) );
  INVX0 U6138_U2 ( .INP(WX5871), .ZN(U6138_n1) );
  NOR2X0 U6138_U1 ( .IN1(n10291), .IN2(U6138_n1), .QN(WX5934) );
  INVX0 U6139_U2 ( .INP(test_so47), .ZN(U6139_n1) );
  NOR2X0 U6139_U1 ( .IN1(n10290), .IN2(U6139_n1), .QN(WX5932) );
  INVX0 U6140_U2 ( .INP(WX5867), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n10290), .IN2(U6140_n1), .QN(WX5930) );
  INVX0 U6141_U2 ( .INP(WX5865), .ZN(U6141_n1) );
  NOR2X0 U6141_U1 ( .IN1(n10289), .IN2(U6141_n1), .QN(WX5928) );
  INVX0 U6142_U2 ( .INP(WX5863), .ZN(U6142_n1) );
  NOR2X0 U6142_U1 ( .IN1(n10289), .IN2(U6142_n1), .QN(WX5926) );
  INVX0 U6143_U2 ( .INP(WX5861), .ZN(U6143_n1) );
  NOR2X0 U6143_U1 ( .IN1(n10289), .IN2(U6143_n1), .QN(WX5924) );
  INVX0 U6144_U2 ( .INP(WX5859), .ZN(U6144_n1) );
  NOR2X0 U6144_U1 ( .IN1(n10289), .IN2(U6144_n1), .QN(WX5922) );
  INVX0 U6145_U2 ( .INP(WX5857), .ZN(U6145_n1) );
  NOR2X0 U6145_U1 ( .IN1(n10288), .IN2(U6145_n1), .QN(WX5920) );
  INVX0 U6146_U2 ( .INP(WX5855), .ZN(U6146_n1) );
  NOR2X0 U6146_U1 ( .IN1(n10288), .IN2(U6146_n1), .QN(WX5918) );
  INVX0 U6147_U2 ( .INP(WX5853), .ZN(U6147_n1) );
  NOR2X0 U6147_U1 ( .IN1(n10288), .IN2(U6147_n1), .QN(WX5916) );
  INVX0 U6148_U2 ( .INP(WX5851), .ZN(U6148_n1) );
  NOR2X0 U6148_U1 ( .IN1(n10288), .IN2(U6148_n1), .QN(WX5914) );
  INVX0 U6149_U2 ( .INP(WX5849), .ZN(U6149_n1) );
  NOR2X0 U6149_U1 ( .IN1(n10288), .IN2(U6149_n1), .QN(WX5912) );
  INVX0 U6150_U2 ( .INP(WX4714), .ZN(U6150_n1) );
  NOR2X0 U6150_U1 ( .IN1(n10288), .IN2(U6150_n1), .QN(WX4777) );
  INVX0 U6151_U2 ( .INP(WX4712), .ZN(U6151_n1) );
  NOR2X0 U6151_U1 ( .IN1(n10288), .IN2(U6151_n1), .QN(WX4775) );
  INVX0 U6152_U2 ( .INP(WX4710), .ZN(U6152_n1) );
  NOR2X0 U6152_U1 ( .IN1(n10288), .IN2(U6152_n1), .QN(WX4773) );
  INVX0 U6153_U2 ( .INP(WX4708), .ZN(U6153_n1) );
  NOR2X0 U6153_U1 ( .IN1(n10288), .IN2(U6153_n1), .QN(WX4771) );
  INVX0 U6154_U2 ( .INP(WX4706), .ZN(U6154_n1) );
  NOR2X0 U6154_U1 ( .IN1(n10288), .IN2(U6154_n1), .QN(WX4769) );
  INVX0 U6155_U2 ( .INP(WX4704), .ZN(U6155_n1) );
  NOR2X0 U6155_U1 ( .IN1(n10293), .IN2(U6155_n1), .QN(WX4767) );
  INVX0 U6156_U2 ( .INP(WX4702), .ZN(U6156_n1) );
  NOR2X0 U6156_U1 ( .IN1(n10305), .IN2(U6156_n1), .QN(WX4765) );
  INVX0 U6157_U2 ( .INP(WX4700), .ZN(U6157_n1) );
  NOR2X0 U6157_U1 ( .IN1(n10308), .IN2(U6157_n1), .QN(WX4763) );
  INVX0 U6158_U2 ( .INP(WX4698), .ZN(U6158_n1) );
  NOR2X0 U6158_U1 ( .IN1(n10308), .IN2(U6158_n1), .QN(WX4761) );
  INVX0 U6159_U2 ( .INP(WX4696), .ZN(U6159_n1) );
  NOR2X0 U6159_U1 ( .IN1(n10306), .IN2(U6159_n1), .QN(WX4759) );
  INVX0 U6160_U2 ( .INP(WX4694), .ZN(U6160_n1) );
  NOR2X0 U6160_U1 ( .IN1(n10308), .IN2(U6160_n1), .QN(WX4757) );
  INVX0 U6161_U2 ( .INP(WX4692), .ZN(U6161_n1) );
  NOR2X0 U6161_U1 ( .IN1(n10307), .IN2(U6161_n1), .QN(WX4755) );
  INVX0 U6162_U2 ( .INP(WX4690), .ZN(U6162_n1) );
  NOR2X0 U6162_U1 ( .IN1(n10306), .IN2(U6162_n1), .QN(WX4753) );
  INVX0 U6163_U2 ( .INP(test_so39), .ZN(U6163_n1) );
  NOR2X0 U6163_U1 ( .IN1(n10254), .IN2(U6163_n1), .QN(WX4751) );
  INVX0 U6164_U2 ( .INP(WX4686), .ZN(U6164_n1) );
  NOR2X0 U6164_U1 ( .IN1(n10253), .IN2(U6164_n1), .QN(WX4749) );
  INVX0 U6165_U2 ( .INP(WX4684), .ZN(U6165_n1) );
  NOR2X0 U6165_U1 ( .IN1(n10253), .IN2(U6165_n1), .QN(WX4747) );
  INVX0 U6166_U2 ( .INP(WX4682), .ZN(U6166_n1) );
  NOR2X0 U6166_U1 ( .IN1(n10253), .IN2(U6166_n1), .QN(WX4745) );
  INVX0 U6167_U2 ( .INP(WX4680), .ZN(U6167_n1) );
  NOR2X0 U6167_U1 ( .IN1(n10253), .IN2(U6167_n1), .QN(WX4743) );
  INVX0 U6168_U2 ( .INP(WX4678), .ZN(U6168_n1) );
  NOR2X0 U6168_U1 ( .IN1(n10253), .IN2(U6168_n1), .QN(WX4741) );
  INVX0 U6169_U2 ( .INP(WX4676), .ZN(U6169_n1) );
  NOR2X0 U6169_U1 ( .IN1(n10253), .IN2(U6169_n1), .QN(WX4739) );
  INVX0 U6170_U2 ( .INP(WX4674), .ZN(U6170_n1) );
  NOR2X0 U6170_U1 ( .IN1(n10253), .IN2(U6170_n1), .QN(WX4737) );
  INVX0 U6171_U2 ( .INP(WX4672), .ZN(U6171_n1) );
  NOR2X0 U6171_U1 ( .IN1(n10253), .IN2(U6171_n1), .QN(WX4735) );
  INVX0 U6172_U2 ( .INP(WX4670), .ZN(U6172_n1) );
  NOR2X0 U6172_U1 ( .IN1(n10253), .IN2(U6172_n1), .QN(WX4733) );
  INVX0 U6173_U2 ( .INP(WX4668), .ZN(U6173_n1) );
  NOR2X0 U6173_U1 ( .IN1(n10253), .IN2(U6173_n1), .QN(WX4731) );
  INVX0 U6174_U2 ( .INP(WX4666), .ZN(U6174_n1) );
  NOR2X0 U6174_U1 ( .IN1(n10253), .IN2(U6174_n1), .QN(WX4729) );
  INVX0 U6175_U2 ( .INP(WX4664), .ZN(U6175_n1) );
  NOR2X0 U6175_U1 ( .IN1(n10252), .IN2(U6175_n1), .QN(WX4727) );
  INVX0 U6176_U2 ( .INP(WX4662), .ZN(U6176_n1) );
  NOR2X0 U6176_U1 ( .IN1(n10252), .IN2(U6176_n1), .QN(WX4725) );
  INVX0 U6177_U2 ( .INP(WX4660), .ZN(U6177_n1) );
  NOR2X0 U6177_U1 ( .IN1(n10252), .IN2(U6177_n1), .QN(WX4723) );
  INVX0 U6178_U2 ( .INP(WX4658), .ZN(U6178_n1) );
  NOR2X0 U6178_U1 ( .IN1(n10252), .IN2(U6178_n1), .QN(WX4721) );
  INVX0 U6179_U2 ( .INP(WX4656), .ZN(U6179_n1) );
  NOR2X0 U6179_U1 ( .IN1(n10252), .IN2(U6179_n1), .QN(WX4719) );
  INVX0 U6180_U2 ( .INP(test_so38), .ZN(U6180_n1) );
  NOR2X0 U6180_U1 ( .IN1(n10252), .IN2(U6180_n1), .QN(WX4717) );
  INVX0 U6181_U2 ( .INP(WX4652), .ZN(U6181_n1) );
  NOR2X0 U6181_U1 ( .IN1(n10252), .IN2(U6181_n1), .QN(WX4715) );
  INVX0 U6182_U2 ( .INP(WX4650), .ZN(U6182_n1) );
  NOR2X0 U6182_U1 ( .IN1(n10252), .IN2(U6182_n1), .QN(WX4713) );
  INVX0 U6183_U2 ( .INP(WX4648), .ZN(U6183_n1) );
  NOR2X0 U6183_U1 ( .IN1(n10252), .IN2(U6183_n1), .QN(WX4711) );
  INVX0 U6184_U2 ( .INP(WX4646), .ZN(U6184_n1) );
  NOR2X0 U6184_U1 ( .IN1(n10252), .IN2(U6184_n1), .QN(WX4709) );
  INVX0 U6185_U2 ( .INP(WX4644), .ZN(U6185_n1) );
  NOR2X0 U6185_U1 ( .IN1(n10252), .IN2(U6185_n1), .QN(WX4707) );
  INVX0 U6186_U2 ( .INP(WX4642), .ZN(U6186_n1) );
  NOR2X0 U6186_U1 ( .IN1(n10251), .IN2(U6186_n1), .QN(WX4705) );
  INVX0 U6187_U2 ( .INP(WX4640), .ZN(U6187_n1) );
  NOR2X0 U6187_U1 ( .IN1(n10251), .IN2(U6187_n1), .QN(WX4703) );
  INVX0 U6188_U2 ( .INP(WX4638), .ZN(U6188_n1) );
  NOR2X0 U6188_U1 ( .IN1(n10251), .IN2(U6188_n1), .QN(WX4701) );
  INVX0 U6189_U2 ( .INP(WX4636), .ZN(U6189_n1) );
  NOR2X0 U6189_U1 ( .IN1(n10251), .IN2(U6189_n1), .QN(WX4699) );
  INVX0 U6190_U2 ( .INP(WX4634), .ZN(U6190_n1) );
  NOR2X0 U6190_U1 ( .IN1(n10251), .IN2(U6190_n1), .QN(WX4697) );
  INVX0 U6191_U2 ( .INP(WX4632), .ZN(U6191_n1) );
  NOR2X0 U6191_U1 ( .IN1(n10251), .IN2(U6191_n1), .QN(WX4695) );
  INVX0 U6192_U2 ( .INP(WX4630), .ZN(U6192_n1) );
  NOR2X0 U6192_U1 ( .IN1(n10251), .IN2(U6192_n1), .QN(WX4693) );
  INVX0 U6193_U2 ( .INP(WX4628), .ZN(U6193_n1) );
  NOR2X0 U6193_U1 ( .IN1(n10251), .IN2(U6193_n1), .QN(WX4691) );
  INVX0 U6194_U2 ( .INP(WX4626), .ZN(U6194_n1) );
  NOR2X0 U6194_U1 ( .IN1(n10251), .IN2(U6194_n1), .QN(WX4689) );
  INVX0 U6195_U2 ( .INP(WX4624), .ZN(U6195_n1) );
  NOR2X0 U6195_U1 ( .IN1(n10251), .IN2(U6195_n1), .QN(WX4687) );
  INVX0 U6196_U2 ( .INP(WX4622), .ZN(U6196_n1) );
  NOR2X0 U6196_U1 ( .IN1(n10251), .IN2(U6196_n1), .QN(WX4685) );
  INVX0 U6197_U2 ( .INP(test_so37), .ZN(U6197_n1) );
  NOR2X0 U6197_U1 ( .IN1(n10250), .IN2(U6197_n1), .QN(WX4683) );
  INVX0 U6198_U2 ( .INP(WX4618), .ZN(U6198_n1) );
  NOR2X0 U6198_U1 ( .IN1(n10250), .IN2(U6198_n1), .QN(WX4681) );
  INVX0 U6199_U2 ( .INP(WX4616), .ZN(U6199_n1) );
  NOR2X0 U6199_U1 ( .IN1(n10250), .IN2(U6199_n1), .QN(WX4679) );
  INVX0 U6200_U2 ( .INP(WX4614), .ZN(U6200_n1) );
  NOR2X0 U6200_U1 ( .IN1(n10250), .IN2(U6200_n1), .QN(WX4677) );
  INVX0 U6201_U2 ( .INP(WX4612), .ZN(U6201_n1) );
  NOR2X0 U6201_U1 ( .IN1(n10250), .IN2(U6201_n1), .QN(WX4675) );
  INVX0 U6202_U2 ( .INP(WX4610), .ZN(U6202_n1) );
  NOR2X0 U6202_U1 ( .IN1(n10250), .IN2(U6202_n1), .QN(WX4673) );
  INVX0 U6203_U2 ( .INP(WX4608), .ZN(U6203_n1) );
  NOR2X0 U6203_U1 ( .IN1(n10250), .IN2(U6203_n1), .QN(WX4671) );
  INVX0 U6204_U2 ( .INP(WX4606), .ZN(U6204_n1) );
  NOR2X0 U6204_U1 ( .IN1(n10250), .IN2(U6204_n1), .QN(WX4669) );
  INVX0 U6205_U2 ( .INP(WX4604), .ZN(U6205_n1) );
  NOR2X0 U6205_U1 ( .IN1(n10250), .IN2(U6205_n1), .QN(WX4667) );
  INVX0 U6206_U2 ( .INP(WX4602), .ZN(U6206_n1) );
  NOR2X0 U6206_U1 ( .IN1(n10250), .IN2(U6206_n1), .QN(WX4665) );
  INVX0 U6207_U2 ( .INP(WX4600), .ZN(U6207_n1) );
  NOR2X0 U6207_U1 ( .IN1(n10250), .IN2(U6207_n1), .QN(WX4663) );
  INVX0 U6208_U2 ( .INP(WX4598), .ZN(U6208_n1) );
  NOR2X0 U6208_U1 ( .IN1(n10249), .IN2(U6208_n1), .QN(WX4661) );
  INVX0 U6209_U2 ( .INP(WX4596), .ZN(U6209_n1) );
  NOR2X0 U6209_U1 ( .IN1(n10249), .IN2(U6209_n1), .QN(WX4659) );
  INVX0 U6210_U2 ( .INP(WX4594), .ZN(U6210_n1) );
  NOR2X0 U6210_U1 ( .IN1(n10249), .IN2(U6210_n1), .QN(WX4657) );
  INVX0 U6211_U2 ( .INP(WX4592), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n10249), .IN2(U6211_n1), .QN(WX4655) );
  INVX0 U6212_U2 ( .INP(WX4590), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n10249), .IN2(U6212_n1), .QN(WX4653) );
  INVX0 U6213_U2 ( .INP(WX4588), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n10249), .IN2(U6213_n1), .QN(WX4651) );
  INVX0 U6214_U2 ( .INP(test_so36), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n10249), .IN2(U6214_n1), .QN(WX4649) );
  INVX0 U6215_U2 ( .INP(WX4584), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n10249), .IN2(U6215_n1), .QN(WX4647) );
  INVX0 U6216_U2 ( .INP(WX4582), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n10249), .IN2(U6216_n1), .QN(WX4645) );
  INVX0 U6217_U2 ( .INP(WX4580), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n10249), .IN2(U6217_n1), .QN(WX4643) );
  INVX0 U6218_U2 ( .INP(WX4578), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n10249), .IN2(U6218_n1), .QN(WX4641) );
  INVX0 U6219_U2 ( .INP(WX4576), .ZN(U6219_n1) );
  NOR2X0 U6219_U1 ( .IN1(n10248), .IN2(U6219_n1), .QN(WX4639) );
  INVX0 U6220_U2 ( .INP(WX4574), .ZN(U6220_n1) );
  NOR2X0 U6220_U1 ( .IN1(n10248), .IN2(U6220_n1), .QN(WX4637) );
  INVX0 U6221_U2 ( .INP(WX4572), .ZN(U6221_n1) );
  NOR2X0 U6221_U1 ( .IN1(n10248), .IN2(U6221_n1), .QN(WX4635) );
  INVX0 U6222_U2 ( .INP(WX4570), .ZN(U6222_n1) );
  NOR2X0 U6222_U1 ( .IN1(n10248), .IN2(U6222_n1), .QN(WX4633) );
  INVX0 U6223_U2 ( .INP(WX4568), .ZN(U6223_n1) );
  NOR2X0 U6223_U1 ( .IN1(n10248), .IN2(U6223_n1), .QN(WX4631) );
  INVX0 U6224_U2 ( .INP(WX4566), .ZN(U6224_n1) );
  NOR2X0 U6224_U1 ( .IN1(n10248), .IN2(U6224_n1), .QN(WX4629) );
  INVX0 U6225_U2 ( .INP(WX4564), .ZN(U6225_n1) );
  NOR2X0 U6225_U1 ( .IN1(n10248), .IN2(U6225_n1), .QN(WX4627) );
  INVX0 U6226_U2 ( .INP(WX4562), .ZN(U6226_n1) );
  NOR2X0 U6226_U1 ( .IN1(n10248), .IN2(U6226_n1), .QN(WX4625) );
  INVX0 U6227_U2 ( .INP(WX4560), .ZN(U6227_n1) );
  NOR2X0 U6227_U1 ( .IN1(n10248), .IN2(U6227_n1), .QN(WX4623) );
  INVX0 U6228_U2 ( .INP(WX4558), .ZN(U6228_n1) );
  NOR2X0 U6228_U1 ( .IN1(n10248), .IN2(U6228_n1), .QN(WX4621) );
  INVX0 U6229_U2 ( .INP(WX4556), .ZN(U6229_n1) );
  NOR2X0 U6229_U1 ( .IN1(n10248), .IN2(U6229_n1), .QN(WX4619) );
  INVX0 U6230_U2 ( .INP(WX3421), .ZN(U6230_n1) );
  NOR2X0 U6230_U1 ( .IN1(n10247), .IN2(U6230_n1), .QN(WX3484) );
  INVX0 U6231_U2 ( .INP(WX3419), .ZN(U6231_n1) );
  NOR2X0 U6231_U1 ( .IN1(n10247), .IN2(U6231_n1), .QN(WX3482) );
  INVX0 U6232_U2 ( .INP(WX3417), .ZN(U6232_n1) );
  NOR2X0 U6232_U1 ( .IN1(n10247), .IN2(U6232_n1), .QN(WX3480) );
  INVX0 U6233_U2 ( .INP(WX3415), .ZN(U6233_n1) );
  NOR2X0 U6233_U1 ( .IN1(n10247), .IN2(U6233_n1), .QN(WX3478) );
  INVX0 U6234_U2 ( .INP(WX3413), .ZN(U6234_n1) );
  NOR2X0 U6234_U1 ( .IN1(n10247), .IN2(U6234_n1), .QN(WX3476) );
  INVX0 U6235_U2 ( .INP(WX3411), .ZN(U6235_n1) );
  NOR2X0 U6235_U1 ( .IN1(n10247), .IN2(U6235_n1), .QN(WX3474) );
  INVX0 U6236_U2 ( .INP(WX3409), .ZN(U6236_n1) );
  NOR2X0 U6236_U1 ( .IN1(n10247), .IN2(U6236_n1), .QN(WX3472) );
  INVX0 U6237_U2 ( .INP(WX3407), .ZN(U6237_n1) );
  NOR2X0 U6237_U1 ( .IN1(n10247), .IN2(U6237_n1), .QN(WX3470) );
  INVX0 U6238_U2 ( .INP(test_so28), .ZN(U6238_n1) );
  NOR2X0 U6238_U1 ( .IN1(n10247), .IN2(U6238_n1), .QN(WX3468) );
  INVX0 U6239_U2 ( .INP(WX3403), .ZN(U6239_n1) );
  NOR2X0 U6239_U1 ( .IN1(n10247), .IN2(U6239_n1), .QN(WX3466) );
  INVX0 U6240_U2 ( .INP(WX3401), .ZN(U6240_n1) );
  NOR2X0 U6240_U1 ( .IN1(n10247), .IN2(U6240_n1), .QN(WX3464) );
  INVX0 U6241_U2 ( .INP(WX3399), .ZN(U6241_n1) );
  NOR2X0 U6241_U1 ( .IN1(n10246), .IN2(U6241_n1), .QN(WX3462) );
  INVX0 U6242_U2 ( .INP(WX3397), .ZN(U6242_n1) );
  NOR2X0 U6242_U1 ( .IN1(n10246), .IN2(U6242_n1), .QN(WX3460) );
  INVX0 U6243_U2 ( .INP(WX3395), .ZN(U6243_n1) );
  NOR2X0 U6243_U1 ( .IN1(n10287), .IN2(U6243_n1), .QN(WX3458) );
  INVX0 U6244_U2 ( .INP(WX3393), .ZN(U6244_n1) );
  NOR2X0 U6244_U1 ( .IN1(n10301), .IN2(U6244_n1), .QN(WX3456) );
  INVX0 U6245_U2 ( .INP(WX3391), .ZN(U6245_n1) );
  NOR2X0 U6245_U1 ( .IN1(n10302), .IN2(U6245_n1), .QN(WX3454) );
  INVX0 U6246_U2 ( .INP(WX3389), .ZN(U6246_n1) );
  NOR2X0 U6246_U1 ( .IN1(n10303), .IN2(U6246_n1), .QN(WX3452) );
  INVX0 U6247_U2 ( .INP(WX3387), .ZN(U6247_n1) );
  NOR2X0 U6247_U1 ( .IN1(n10304), .IN2(U6247_n1), .QN(WX3450) );
  INVX0 U6248_U2 ( .INP(WX3385), .ZN(U6248_n1) );
  NOR2X0 U6248_U1 ( .IN1(n10305), .IN2(U6248_n1), .QN(WX3448) );
  INVX0 U6249_U2 ( .INP(WX3383), .ZN(U6249_n1) );
  NOR2X0 U6249_U1 ( .IN1(n10244), .IN2(U6249_n1), .QN(WX3446) );
  INVX0 U6250_U2 ( .INP(WX3381), .ZN(U6250_n1) );
  NOR2X0 U6250_U1 ( .IN1(n10244), .IN2(U6250_n1), .QN(WX3444) );
  INVX0 U6251_U2 ( .INP(WX3379), .ZN(U6251_n1) );
  NOR2X0 U6251_U1 ( .IN1(n10244), .IN2(U6251_n1), .QN(WX3442) );
  INVX0 U6252_U2 ( .INP(WX3377), .ZN(U6252_n1) );
  NOR2X0 U6252_U1 ( .IN1(n10244), .IN2(U6252_n1), .QN(WX3440) );
  INVX0 U6253_U2 ( .INP(WX3375), .ZN(U6253_n1) );
  NOR2X0 U6253_U1 ( .IN1(n10244), .IN2(U6253_n1), .QN(WX3438) );
  INVX0 U6254_U2 ( .INP(WX3373), .ZN(U6254_n1) );
  NOR2X0 U6254_U1 ( .IN1(n10244), .IN2(U6254_n1), .QN(WX3436) );
  INVX0 U6255_U2 ( .INP(WX3371), .ZN(U6255_n1) );
  NOR2X0 U6255_U1 ( .IN1(n10244), .IN2(U6255_n1), .QN(WX3434) );
  INVX0 U6256_U2 ( .INP(test_so27), .ZN(U6256_n1) );
  NOR2X0 U6256_U1 ( .IN1(n10244), .IN2(U6256_n1), .QN(WX3432) );
  INVX0 U6257_U2 ( .INP(WX3367), .ZN(U6257_n1) );
  NOR2X0 U6257_U1 ( .IN1(n10244), .IN2(U6257_n1), .QN(WX3430) );
  INVX0 U6258_U2 ( .INP(WX3365), .ZN(U6258_n1) );
  NOR2X0 U6258_U1 ( .IN1(n10244), .IN2(U6258_n1), .QN(WX3428) );
  INVX0 U6259_U2 ( .INP(WX3363), .ZN(U6259_n1) );
  NOR2X0 U6259_U1 ( .IN1(n10244), .IN2(U6259_n1), .QN(WX3426) );
  INVX0 U6260_U2 ( .INP(WX3361), .ZN(U6260_n1) );
  NOR2X0 U6260_U1 ( .IN1(n10265), .IN2(U6260_n1), .QN(WX3424) );
  INVX0 U6261_U2 ( .INP(WX3359), .ZN(U6261_n1) );
  NOR2X0 U6261_U1 ( .IN1(n10266), .IN2(U6261_n1), .QN(WX3422) );
  INVX0 U6262_U2 ( .INP(WX3357), .ZN(U6262_n1) );
  NOR2X0 U6262_U1 ( .IN1(n10267), .IN2(U6262_n1), .QN(WX3420) );
  INVX0 U6263_U2 ( .INP(WX3355), .ZN(U6263_n1) );
  NOR2X0 U6263_U1 ( .IN1(n10253), .IN2(U6263_n1), .QN(WX3418) );
  INVX0 U6264_U2 ( .INP(WX3353), .ZN(U6264_n1) );
  NOR2X0 U6264_U1 ( .IN1(n10254), .IN2(U6264_n1), .QN(WX3416) );
  INVX0 U6265_U2 ( .INP(WX3351), .ZN(U6265_n1) );
  NOR2X0 U6265_U1 ( .IN1(n10255), .IN2(U6265_n1), .QN(WX3414) );
  INVX0 U6266_U2 ( .INP(WX3349), .ZN(U6266_n1) );
  NOR2X0 U6266_U1 ( .IN1(n10256), .IN2(U6266_n1), .QN(WX3412) );
  INVX0 U6267_U2 ( .INP(WX3347), .ZN(U6267_n1) );
  NOR2X0 U6267_U1 ( .IN1(n10257), .IN2(U6267_n1), .QN(WX3410) );
  INVX0 U6268_U2 ( .INP(WX3345), .ZN(U6268_n1) );
  NOR2X0 U6268_U1 ( .IN1(n10258), .IN2(U6268_n1), .QN(WX3408) );
  INVX0 U6269_U2 ( .INP(WX3343), .ZN(U6269_n1) );
  NOR2X0 U6269_U1 ( .IN1(n10259), .IN2(U6269_n1), .QN(WX3406) );
  INVX0 U6270_U2 ( .INP(WX3341), .ZN(U6270_n1) );
  NOR2X0 U6270_U1 ( .IN1(n10260), .IN2(U6270_n1), .QN(WX3404) );
  INVX0 U6271_U2 ( .INP(WX3339), .ZN(U6271_n1) );
  NOR2X0 U6271_U1 ( .IN1(n10245), .IN2(U6271_n1), .QN(WX3402) );
  INVX0 U6272_U2 ( .INP(WX3337), .ZN(U6272_n1) );
  NOR2X0 U6272_U1 ( .IN1(n10246), .IN2(U6272_n1), .QN(WX3400) );
  INVX0 U6273_U2 ( .INP(WX3335), .ZN(U6273_n1) );
  NOR2X0 U6273_U1 ( .IN1(n10247), .IN2(U6273_n1), .QN(WX3398) );
  INVX0 U6274_U2 ( .INP(test_so26), .ZN(U6274_n1) );
  NOR2X0 U6274_U1 ( .IN1(n10248), .IN2(U6274_n1), .QN(WX3396) );
  INVX0 U6275_U2 ( .INP(WX3331), .ZN(U6275_n1) );
  NOR2X0 U6275_U1 ( .IN1(n10249), .IN2(U6275_n1), .QN(WX3394) );
  INVX0 U6276_U2 ( .INP(WX3329), .ZN(U6276_n1) );
  NOR2X0 U6276_U1 ( .IN1(n10250), .IN2(U6276_n1), .QN(WX3392) );
  INVX0 U6277_U2 ( .INP(WX3327), .ZN(U6277_n1) );
  NOR2X0 U6277_U1 ( .IN1(n10251), .IN2(U6277_n1), .QN(WX3390) );
  INVX0 U6278_U2 ( .INP(WX3325), .ZN(U6278_n1) );
  NOR2X0 U6278_U1 ( .IN1(n10252), .IN2(U6278_n1), .QN(WX3388) );
  INVX0 U6279_U2 ( .INP(WX3323), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n10283), .IN2(U6279_n1), .QN(WX3386) );
  INVX0 U6280_U2 ( .INP(WX3321), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n10284), .IN2(U6280_n1), .QN(WX3384) );
  INVX0 U6281_U2 ( .INP(WX3319), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n10285), .IN2(U6281_n1), .QN(WX3382) );
  INVX0 U6282_U2 ( .INP(WX3317), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n10286), .IN2(U6282_n1), .QN(WX3380) );
  INVX0 U6283_U2 ( .INP(WX3315), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n10288), .IN2(U6283_n1), .QN(WX3378) );
  INVX0 U6284_U2 ( .INP(WX3313), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n10289), .IN2(U6284_n1), .QN(WX3376) );
  INVX0 U6285_U2 ( .INP(WX3311), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n10290), .IN2(U6285_n1), .QN(WX3374) );
  INVX0 U6286_U2 ( .INP(WX3309), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n10276), .IN2(U6286_n1), .QN(WX3372) );
  INVX0 U6287_U2 ( .INP(WX3307), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n10277), .IN2(U6287_n1), .QN(WX3370) );
  INVX0 U6288_U2 ( .INP(WX3305), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n10278), .IN2(U6288_n1), .QN(WX3368) );
  INVX0 U6289_U2 ( .INP(WX3303), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n10279), .IN2(U6289_n1), .QN(WX3366) );
  INVX0 U6290_U2 ( .INP(WX3301), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n10280), .IN2(U6290_n1), .QN(WX3364) );
  INVX0 U6291_U2 ( .INP(WX3299), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n10281), .IN2(U6291_n1), .QN(WX3362) );
  INVX0 U6292_U2 ( .INP(test_so25), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n10282), .IN2(U6292_n1), .QN(WX3360) );
  INVX0 U6293_U2 ( .INP(WX3295), .ZN(U6293_n1) );
  NOR2X0 U6293_U1 ( .IN1(n10268), .IN2(U6293_n1), .QN(WX3358) );
  INVX0 U6294_U2 ( .INP(WX3293), .ZN(U6294_n1) );
  NOR2X0 U6294_U1 ( .IN1(n10269), .IN2(U6294_n1), .QN(WX3356) );
  INVX0 U6295_U2 ( .INP(WX3291), .ZN(U6295_n1) );
  NOR2X0 U6295_U1 ( .IN1(n10270), .IN2(U6295_n1), .QN(WX3354) );
  INVX0 U6296_U2 ( .INP(WX3289), .ZN(U6296_n1) );
  NOR2X0 U6296_U1 ( .IN1(n10271), .IN2(U6296_n1), .QN(WX3352) );
  INVX0 U6297_U2 ( .INP(WX3287), .ZN(U6297_n1) );
  NOR2X0 U6297_U1 ( .IN1(n10272), .IN2(U6297_n1), .QN(WX3350) );
  INVX0 U6298_U2 ( .INP(WX3285), .ZN(U6298_n1) );
  NOR2X0 U6298_U1 ( .IN1(n10273), .IN2(U6298_n1), .QN(WX3348) );
  INVX0 U6299_U2 ( .INP(WX3283), .ZN(U6299_n1) );
  NOR2X0 U6299_U1 ( .IN1(n10274), .IN2(U6299_n1), .QN(WX3346) );
  INVX0 U6300_U2 ( .INP(WX3281), .ZN(U6300_n1) );
  NOR2X0 U6300_U1 ( .IN1(n10275), .IN2(U6300_n1), .QN(WX3344) );
  INVX0 U6301_U2 ( .INP(WX3279), .ZN(U6301_n1) );
  NOR2X0 U6301_U1 ( .IN1(n10307), .IN2(U6301_n1), .QN(WX3342) );
  INVX0 U6302_U2 ( .INP(WX3277), .ZN(U6302_n1) );
  NOR2X0 U6302_U1 ( .IN1(n10299), .IN2(U6302_n1), .QN(WX3340) );
  INVX0 U6303_U2 ( .INP(WX3275), .ZN(U6303_n1) );
  NOR2X0 U6303_U1 ( .IN1(n10245), .IN2(U6303_n1), .QN(WX3338) );
  INVX0 U6304_U2 ( .INP(WX3273), .ZN(U6304_n1) );
  NOR2X0 U6304_U1 ( .IN1(n10245), .IN2(U6304_n1), .QN(WX3336) );
  INVX0 U6305_U2 ( .INP(WX3271), .ZN(U6305_n1) );
  NOR2X0 U6305_U1 ( .IN1(n10245), .IN2(U6305_n1), .QN(WX3334) );
  INVX0 U6306_U2 ( .INP(WX3267), .ZN(U6306_n1) );
  NOR2X0 U6306_U1 ( .IN1(n10245), .IN2(U6306_n1), .QN(WX3330) );
  INVX0 U6307_U2 ( .INP(WX2128), .ZN(U6307_n1) );
  NOR2X0 U6307_U1 ( .IN1(n10245), .IN2(U6307_n1), .QN(WX2191) );
  INVX0 U6308_U2 ( .INP(WX2126), .ZN(U6308_n1) );
  NOR2X0 U6308_U1 ( .IN1(n10245), .IN2(U6308_n1), .QN(WX2189) );
  INVX0 U6309_U2 ( .INP(WX2124), .ZN(U6309_n1) );
  NOR2X0 U6309_U1 ( .IN1(n10245), .IN2(U6309_n1), .QN(WX2187) );
  INVX0 U6310_U2 ( .INP(WX2122), .ZN(U6310_n1) );
  NOR2X0 U6310_U1 ( .IN1(n10245), .IN2(U6310_n1), .QN(WX2185) );
  INVX0 U6311_U2 ( .INP(WX2120), .ZN(U6311_n1) );
  NOR2X0 U6311_U1 ( .IN1(n10245), .IN2(U6311_n1), .QN(WX2183) );
  INVX0 U6312_U2 ( .INP(WX2118), .ZN(U6312_n1) );
  NOR2X0 U6312_U1 ( .IN1(n10245), .IN2(U6312_n1), .QN(WX2181) );
  INVX0 U6313_U2 ( .INP(WX2116), .ZN(U6313_n1) );
  NOR2X0 U6313_U1 ( .IN1(n10245), .IN2(U6313_n1), .QN(WX2179) );
  INVX0 U6314_U2 ( .INP(WX2114), .ZN(U6314_n1) );
  NOR2X0 U6314_U1 ( .IN1(n10246), .IN2(U6314_n1), .QN(WX2177) );
  INVX0 U6315_U2 ( .INP(WX2112), .ZN(U6315_n1) );
  NOR2X0 U6315_U1 ( .IN1(n10246), .IN2(U6315_n1), .QN(WX2175) );
  INVX0 U6316_U2 ( .INP(WX2110), .ZN(U6316_n1) );
  NOR2X0 U6316_U1 ( .IN1(n10246), .IN2(U6316_n1), .QN(WX2173) );
  INVX0 U6317_U2 ( .INP(WX2108), .ZN(U6317_n1) );
  NOR2X0 U6317_U1 ( .IN1(n10246), .IN2(U6317_n1), .QN(WX2171) );
  INVX0 U6318_U2 ( .INP(WX2106), .ZN(U6318_n1) );
  NOR2X0 U6318_U1 ( .IN1(n10246), .IN2(U6318_n1), .QN(WX2169) );
  INVX0 U6319_U2 ( .INP(WX2104), .ZN(U6319_n1) );
  NOR2X0 U6319_U1 ( .IN1(n10246), .IN2(U6319_n1), .QN(WX2167) );
  INVX0 U6320_U2 ( .INP(WX2102), .ZN(U6320_n1) );
  NOR2X0 U6320_U1 ( .IN1(n10246), .IN2(U6320_n1), .QN(WX2165) );
  INVX0 U6321_U2 ( .INP(test_so17), .ZN(U6321_n1) );
  NOR2X0 U6321_U1 ( .IN1(n10246), .IN2(U6321_n1), .QN(WX2163) );
  INVX0 U6322_U2 ( .INP(WX2098), .ZN(U6322_n1) );
  NOR2X0 U6322_U1 ( .IN1(n10246), .IN2(U6322_n1), .QN(WX2161) );
  INVX0 U6323_U2 ( .INP(WX2096), .ZN(U6323_n1) );
  NOR2X0 U6323_U1 ( .IN1(n10267), .IN2(U6323_n1), .QN(WX2159) );
  INVX0 U6324_U2 ( .INP(WX2094), .ZN(U6324_n1) );
  NOR2X0 U6324_U1 ( .IN1(n10267), .IN2(U6324_n1), .QN(WX2157) );
  INVX0 U6325_U2 ( .INP(WX2092), .ZN(U6325_n1) );
  NOR2X0 U6325_U1 ( .IN1(n10267), .IN2(U6325_n1), .QN(WX2155) );
  INVX0 U6326_U2 ( .INP(WX2090), .ZN(U6326_n1) );
  NOR2X0 U6326_U1 ( .IN1(n10267), .IN2(U6326_n1), .QN(WX2153) );
  INVX0 U6327_U2 ( .INP(WX2088), .ZN(U6327_n1) );
  NOR2X0 U6327_U1 ( .IN1(n10267), .IN2(U6327_n1), .QN(WX2151) );
  INVX0 U6328_U2 ( .INP(WX2086), .ZN(U6328_n1) );
  NOR2X0 U6328_U1 ( .IN1(n10267), .IN2(U6328_n1), .QN(WX2149) );
  INVX0 U6329_U2 ( .INP(WX2084), .ZN(U6329_n1) );
  NOR2X0 U6329_U1 ( .IN1(n10267), .IN2(U6329_n1), .QN(WX2147) );
  INVX0 U6330_U2 ( .INP(WX2082), .ZN(U6330_n1) );
  NOR2X0 U6330_U1 ( .IN1(n10266), .IN2(U6330_n1), .QN(WX2145) );
  INVX0 U6331_U2 ( .INP(WX2080), .ZN(U6331_n1) );
  NOR2X0 U6331_U1 ( .IN1(n10266), .IN2(U6331_n1), .QN(WX2143) );
  INVX0 U6332_U2 ( .INP(WX2078), .ZN(U6332_n1) );
  NOR2X0 U6332_U1 ( .IN1(n10266), .IN2(U6332_n1), .QN(WX2141) );
  INVX0 U6333_U2 ( .INP(WX2076), .ZN(U6333_n1) );
  NOR2X0 U6333_U1 ( .IN1(n10266), .IN2(U6333_n1), .QN(WX2139) );
  INVX0 U6334_U2 ( .INP(WX2074), .ZN(U6334_n1) );
  NOR2X0 U6334_U1 ( .IN1(n10266), .IN2(U6334_n1), .QN(WX2137) );
  INVX0 U6335_U2 ( .INP(WX2072), .ZN(U6335_n1) );
  NOR2X0 U6335_U1 ( .IN1(n10266), .IN2(U6335_n1), .QN(WX2135) );
  INVX0 U6336_U2 ( .INP(WX2070), .ZN(U6336_n1) );
  NOR2X0 U6336_U1 ( .IN1(n10266), .IN2(U6336_n1), .QN(WX2133) );
  INVX0 U6337_U2 ( .INP(WX2068), .ZN(U6337_n1) );
  NOR2X0 U6337_U1 ( .IN1(n10266), .IN2(U6337_n1), .QN(WX2131) );
  INVX0 U6338_U2 ( .INP(WX2066), .ZN(U6338_n1) );
  NOR2X0 U6338_U1 ( .IN1(n10266), .IN2(U6338_n1), .QN(WX2129) );
  INVX0 U6339_U2 ( .INP(test_so16), .ZN(U6339_n1) );
  NOR2X0 U6339_U1 ( .IN1(n10266), .IN2(U6339_n1), .QN(WX2127) );
  INVX0 U6340_U2 ( .INP(WX2062), .ZN(U6340_n1) );
  NOR2X0 U6340_U1 ( .IN1(n10266), .IN2(U6340_n1), .QN(WX2125) );
  INVX0 U6341_U2 ( .INP(WX2060), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n10265), .IN2(U6341_n1), .QN(WX2123) );
  INVX0 U6342_U2 ( .INP(WX2058), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n10265), .IN2(U6342_n1), .QN(WX2121) );
  INVX0 U6343_U2 ( .INP(WX2056), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n10265), .IN2(U6343_n1), .QN(WX2119) );
  INVX0 U6344_U2 ( .INP(WX2054), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n10265), .IN2(U6344_n1), .QN(WX2117) );
  INVX0 U6345_U2 ( .INP(WX2052), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n10265), .IN2(U6345_n1), .QN(WX2115) );
  INVX0 U6346_U2 ( .INP(WX2050), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n10265), .IN2(U6346_n1), .QN(WX2113) );
  INVX0 U6347_U2 ( .INP(WX2048), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n10265), .IN2(U6347_n1), .QN(WX2111) );
  INVX0 U6348_U2 ( .INP(WX2046), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n10265), .IN2(U6348_n1), .QN(WX2109) );
  INVX0 U6349_U2 ( .INP(WX2044), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n10265), .IN2(U6349_n1), .QN(WX2107) );
  INVX0 U6350_U2 ( .INP(WX2042), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n10265), .IN2(U6350_n1), .QN(WX2105) );
  INVX0 U6351_U2 ( .INP(WX2040), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n10265), .IN2(U6351_n1), .QN(WX2103) );
  INVX0 U6352_U2 ( .INP(WX2038), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n10264), .IN2(U6352_n1), .QN(WX2101) );
  INVX0 U6353_U2 ( .INP(WX2036), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n10264), .IN2(U6353_n1), .QN(WX2099) );
  INVX0 U6354_U2 ( .INP(WX2034), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n10264), .IN2(U6354_n1), .QN(WX2097) );
  INVX0 U6355_U2 ( .INP(WX2032), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n10264), .IN2(U6355_n1), .QN(WX2095) );
  INVX0 U6356_U2 ( .INP(WX2030), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n10264), .IN2(U6356_n1), .QN(WX2093) );
  INVX0 U6357_U2 ( .INP(test_so15), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n10264), .IN2(U6357_n1), .QN(WX2091) );
  INVX0 U6358_U2 ( .INP(WX2026), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n10264), .IN2(U6358_n1), .QN(WX2089) );
  INVX0 U6359_U2 ( .INP(WX2024), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n10264), .IN2(U6359_n1), .QN(WX2087) );
  INVX0 U6360_U2 ( .INP(WX2022), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n10264), .IN2(U6360_n1), .QN(WX2085) );
  INVX0 U6361_U2 ( .INP(WX2020), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n10264), .IN2(U6361_n1), .QN(WX2083) );
  INVX0 U6362_U2 ( .INP(WX2018), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n10264), .IN2(U6362_n1), .QN(WX2081) );
  INVX0 U6363_U2 ( .INP(WX2016), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n10263), .IN2(U6363_n1), .QN(WX2079) );
  INVX0 U6364_U2 ( .INP(WX2014), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n10263), .IN2(U6364_n1), .QN(WX2077) );
  INVX0 U6365_U2 ( .INP(WX2012), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n10263), .IN2(U6365_n1), .QN(WX2075) );
  INVX0 U6366_U2 ( .INP(WX2010), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n10263), .IN2(U6366_n1), .QN(WX2073) );
  INVX0 U6367_U2 ( .INP(WX2008), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n10263), .IN2(U6367_n1), .QN(WX2071) );
  INVX0 U6368_U2 ( .INP(WX2006), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n10263), .IN2(U6368_n1), .QN(WX2069) );
  INVX0 U6369_U2 ( .INP(WX2004), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n10263), .IN2(U6369_n1), .QN(WX2067) );
  INVX0 U6370_U2 ( .INP(WX2002), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n10263), .IN2(U6370_n1), .QN(WX2065) );
  INVX0 U6371_U2 ( .INP(WX2000), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n10263), .IN2(U6371_n1), .QN(WX2063) );
  INVX0 U6372_U2 ( .INP(WX1998), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n10263), .IN2(U6372_n1), .QN(WX2061) );
  INVX0 U6373_U2 ( .INP(WX1996), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n10263), .IN2(U6373_n1), .QN(WX2059) );
  INVX0 U6374_U2 ( .INP(WX1994), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n10262), .IN2(U6374_n1), .QN(WX2057) );
  INVX0 U6375_U2 ( .INP(test_so14), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n10262), .IN2(U6375_n1), .QN(WX2055) );
  INVX0 U6376_U2 ( .INP(WX1990), .ZN(U6376_n1) );
  NOR2X0 U6376_U1 ( .IN1(n10262), .IN2(U6376_n1), .QN(WX2053) );
  INVX0 U6377_U2 ( .INP(WX1988), .ZN(U6377_n1) );
  NOR2X0 U6377_U1 ( .IN1(n10262), .IN2(U6377_n1), .QN(WX2051) );
  INVX0 U6378_U2 ( .INP(WX1986), .ZN(U6378_n1) );
  NOR2X0 U6378_U1 ( .IN1(n10262), .IN2(U6378_n1), .QN(WX2049) );
  INVX0 U6379_U2 ( .INP(WX1984), .ZN(U6379_n1) );
  NOR2X0 U6379_U1 ( .IN1(n10262), .IN2(U6379_n1), .QN(WX2047) );
  INVX0 U6380_U2 ( .INP(WX1982), .ZN(U6380_n1) );
  NOR2X0 U6380_U1 ( .IN1(n10262), .IN2(U6380_n1), .QN(WX2045) );
  INVX0 U6381_U2 ( .INP(WX1980), .ZN(U6381_n1) );
  NOR2X0 U6381_U1 ( .IN1(n10262), .IN2(U6381_n1), .QN(WX2043) );
  INVX0 U6382_U2 ( .INP(WX1978), .ZN(U6382_n1) );
  NOR2X0 U6382_U1 ( .IN1(n10262), .IN2(U6382_n1), .QN(WX2041) );
  INVX0 U6383_U2 ( .INP(WX1976), .ZN(U6383_n1) );
  NOR2X0 U6383_U1 ( .IN1(n10262), .IN2(U6383_n1), .QN(WX2039) );
  INVX0 U6384_U2 ( .INP(WX1974), .ZN(U6384_n1) );
  NOR2X0 U6384_U1 ( .IN1(n10262), .IN2(U6384_n1), .QN(WX2037) );
  INVX0 U6385_U2 ( .INP(WX1972), .ZN(U6385_n1) );
  NOR2X0 U6385_U1 ( .IN1(n10261), .IN2(U6385_n1), .QN(WX2035) );
  INVX0 U6386_U2 ( .INP(WX1970), .ZN(U6386_n1) );
  NOR2X0 U6386_U1 ( .IN1(n10261), .IN2(U6386_n1), .QN(WX2033) );
  INVX0 U6387_U2 ( .INP(WX835), .ZN(U6387_n1) );
  NOR2X0 U6387_U1 ( .IN1(n10261), .IN2(U6387_n1), .QN(WX898) );
  INVX0 U6388_U2 ( .INP(WX833), .ZN(U6388_n1) );
  NOR2X0 U6388_U1 ( .IN1(n10261), .IN2(U6388_n1), .QN(WX896) );
  INVX0 U6389_U2 ( .INP(test_so7), .ZN(U6389_n1) );
  NOR2X0 U6389_U1 ( .IN1(n10261), .IN2(U6389_n1), .QN(WX894) );
  INVX0 U6390_U2 ( .INP(WX829), .ZN(U6390_n1) );
  NOR2X0 U6390_U1 ( .IN1(n10261), .IN2(U6390_n1), .QN(WX892) );
  INVX0 U6391_U2 ( .INP(WX827), .ZN(U6391_n1) );
  NOR2X0 U6391_U1 ( .IN1(n10261), .IN2(U6391_n1), .QN(WX890) );
  INVX0 U6392_U2 ( .INP(WX825), .ZN(U6392_n1) );
  NOR2X0 U6392_U1 ( .IN1(n10261), .IN2(U6392_n1), .QN(WX888) );
  INVX0 U6393_U2 ( .INP(WX823), .ZN(U6393_n1) );
  NOR2X0 U6393_U1 ( .IN1(n10261), .IN2(U6393_n1), .QN(WX886) );
  INVX0 U6394_U2 ( .INP(WX821), .ZN(U6394_n1) );
  NOR2X0 U6394_U1 ( .IN1(n10261), .IN2(U6394_n1), .QN(WX884) );
  INVX0 U6395_U2 ( .INP(WX819), .ZN(U6395_n1) );
  NOR2X0 U6395_U1 ( .IN1(n10261), .IN2(U6395_n1), .QN(WX882) );
  INVX0 U6396_U2 ( .INP(WX817), .ZN(U6396_n1) );
  NOR2X0 U6396_U1 ( .IN1(n10244), .IN2(U6396_n1), .QN(WX880) );
  INVX0 U6397_U2 ( .INP(WX815), .ZN(U6397_n1) );
  NOR2X0 U6397_U1 ( .IN1(n10264), .IN2(U6397_n1), .QN(WX878) );
  INVX0 U6398_U2 ( .INP(WX813), .ZN(U6398_n1) );
  NOR2X0 U6398_U1 ( .IN1(n10263), .IN2(U6398_n1), .QN(WX876) );
  INVX0 U6399_U2 ( .INP(WX811), .ZN(U6399_n1) );
  NOR2X0 U6399_U1 ( .IN1(n10262), .IN2(U6399_n1), .QN(WX874) );
  INVX0 U6400_U2 ( .INP(WX809), .ZN(U6400_n1) );
  NOR2X0 U6400_U1 ( .IN1(n10261), .IN2(U6400_n1), .QN(WX872) );
  INVX0 U6401_U2 ( .INP(WX807), .ZN(U6401_n1) );
  NOR2X0 U6401_U1 ( .IN1(n10298), .IN2(U6401_n1), .QN(WX870) );
  INVX0 U6402_U2 ( .INP(WX805), .ZN(U6402_n1) );
  NOR2X0 U6402_U1 ( .IN1(n10297), .IN2(U6402_n1), .QN(WX868) );
  INVX0 U6403_U2 ( .INP(WX803), .ZN(U6403_n1) );
  NOR2X0 U6403_U1 ( .IN1(n10295), .IN2(U6403_n1), .QN(WX866) );
  INVX0 U6404_U2 ( .INP(WX801), .ZN(U6404_n1) );
  NOR2X0 U6404_U1 ( .IN1(n10305), .IN2(U6404_n1), .QN(WX864) );
  INVX0 U6405_U2 ( .INP(WX799), .ZN(U6405_n1) );
  NOR2X0 U6405_U1 ( .IN1(n10304), .IN2(U6405_n1), .QN(WX862) );
  INVX0 U6406_U2 ( .INP(WX797), .ZN(U6406_n1) );
  NOR2X0 U6406_U1 ( .IN1(n10260), .IN2(U6406_n1), .QN(WX860) );
  INVX0 U6407_U2 ( .INP(test_so6), .ZN(U6407_n1) );
  NOR2X0 U6407_U1 ( .IN1(n10260), .IN2(U6407_n1), .QN(WX858) );
  INVX0 U6408_U2 ( .INP(WX793), .ZN(U6408_n1) );
  NOR2X0 U6408_U1 ( .IN1(n10260), .IN2(U6408_n1), .QN(WX856) );
  INVX0 U6409_U2 ( .INP(WX791), .ZN(U6409_n1) );
  NOR2X0 U6409_U1 ( .IN1(n10260), .IN2(U6409_n1), .QN(WX854) );
  INVX0 U6410_U2 ( .INP(WX789), .ZN(U6410_n1) );
  NOR2X0 U6410_U1 ( .IN1(n10260), .IN2(U6410_n1), .QN(WX852) );
  INVX0 U6411_U2 ( .INP(WX787), .ZN(U6411_n1) );
  NOR2X0 U6411_U1 ( .IN1(n10260), .IN2(U6411_n1), .QN(WX850) );
  INVX0 U6412_U2 ( .INP(WX785), .ZN(U6412_n1) );
  NOR2X0 U6412_U1 ( .IN1(n10260), .IN2(U6412_n1), .QN(WX848) );
  INVX0 U6413_U2 ( .INP(WX783), .ZN(U6413_n1) );
  NOR2X0 U6413_U1 ( .IN1(n10260), .IN2(U6413_n1), .QN(WX846) );
  INVX0 U6414_U2 ( .INP(WX781), .ZN(U6414_n1) );
  NOR2X0 U6414_U1 ( .IN1(n10260), .IN2(U6414_n1), .QN(WX844) );
  INVX0 U6415_U2 ( .INP(WX779), .ZN(U6415_n1) );
  NOR2X0 U6415_U1 ( .IN1(n10260), .IN2(U6415_n1), .QN(WX842) );
  INVX0 U6416_U2 ( .INP(WX777), .ZN(U6416_n1) );
  NOR2X0 U6416_U1 ( .IN1(n10260), .IN2(U6416_n1), .QN(WX840) );
  INVX0 U6417_U2 ( .INP(WX775), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n10259), .IN2(U6417_n1), .QN(WX838) );
  INVX0 U6418_U2 ( .INP(WX773), .ZN(U6418_n1) );
  NOR2X0 U6418_U1 ( .IN1(n10259), .IN2(U6418_n1), .QN(WX836) );
  INVX0 U6419_U2 ( .INP(WX771), .ZN(U6419_n1) );
  NOR2X0 U6419_U1 ( .IN1(n10259), .IN2(U6419_n1), .QN(WX834) );
  INVX0 U6420_U2 ( .INP(WX769), .ZN(U6420_n1) );
  NOR2X0 U6420_U1 ( .IN1(n10259), .IN2(U6420_n1), .QN(WX832) );
  INVX0 U6421_U2 ( .INP(WX767), .ZN(U6421_n1) );
  NOR2X0 U6421_U1 ( .IN1(n10259), .IN2(U6421_n1), .QN(WX830) );
  INVX0 U6422_U2 ( .INP(WX765), .ZN(U6422_n1) );
  NOR2X0 U6422_U1 ( .IN1(n10259), .IN2(U6422_n1), .QN(WX828) );
  INVX0 U6423_U2 ( .INP(WX763), .ZN(U6423_n1) );
  NOR2X0 U6423_U1 ( .IN1(n10259), .IN2(U6423_n1), .QN(WX826) );
  INVX0 U6424_U2 ( .INP(WX761), .ZN(U6424_n1) );
  NOR2X0 U6424_U1 ( .IN1(n10259), .IN2(U6424_n1), .QN(WX824) );
  INVX0 U6425_U2 ( .INP(test_so5), .ZN(U6425_n1) );
  NOR2X0 U6425_U1 ( .IN1(n10259), .IN2(U6425_n1), .QN(WX822) );
  INVX0 U6426_U2 ( .INP(WX757), .ZN(U6426_n1) );
  NOR2X0 U6426_U1 ( .IN1(n10259), .IN2(U6426_n1), .QN(WX820) );
  INVX0 U6427_U2 ( .INP(WX755), .ZN(U6427_n1) );
  NOR2X0 U6427_U1 ( .IN1(n10259), .IN2(U6427_n1), .QN(WX818) );
  INVX0 U6428_U2 ( .INP(WX753), .ZN(U6428_n1) );
  NOR2X0 U6428_U1 ( .IN1(n10258), .IN2(U6428_n1), .QN(WX816) );
  INVX0 U6429_U2 ( .INP(WX751), .ZN(U6429_n1) );
  NOR2X0 U6429_U1 ( .IN1(n10258), .IN2(U6429_n1), .QN(WX814) );
  INVX0 U6430_U2 ( .INP(WX749), .ZN(U6430_n1) );
  NOR2X0 U6430_U1 ( .IN1(n10258), .IN2(U6430_n1), .QN(WX812) );
  INVX0 U6431_U2 ( .INP(WX747), .ZN(U6431_n1) );
  NOR2X0 U6431_U1 ( .IN1(n10258), .IN2(U6431_n1), .QN(WX810) );
  INVX0 U6432_U2 ( .INP(WX745), .ZN(U6432_n1) );
  NOR2X0 U6432_U1 ( .IN1(n10258), .IN2(U6432_n1), .QN(WX808) );
  INVX0 U6433_U2 ( .INP(WX743), .ZN(U6433_n1) );
  NOR2X0 U6433_U1 ( .IN1(n10258), .IN2(U6433_n1), .QN(WX806) );
  INVX0 U6434_U2 ( .INP(WX741), .ZN(U6434_n1) );
  NOR2X0 U6434_U1 ( .IN1(n10258), .IN2(U6434_n1), .QN(WX804) );
  INVX0 U6435_U2 ( .INP(WX739), .ZN(U6435_n1) );
  NOR2X0 U6435_U1 ( .IN1(n10258), .IN2(U6435_n1), .QN(WX802) );
  INVX0 U6436_U2 ( .INP(WX737), .ZN(U6436_n1) );
  NOR2X0 U6436_U1 ( .IN1(n10258), .IN2(U6436_n1), .QN(WX800) );
  INVX0 U6437_U2 ( .INP(WX735), .ZN(U6437_n1) );
  NOR2X0 U6437_U1 ( .IN1(n10258), .IN2(U6437_n1), .QN(WX798) );
  INVX0 U6438_U2 ( .INP(WX733), .ZN(U6438_n1) );
  NOR2X0 U6438_U1 ( .IN1(n10258), .IN2(U6438_n1), .QN(WX796) );
  INVX0 U6439_U2 ( .INP(WX731), .ZN(U6439_n1) );
  NOR2X0 U6439_U1 ( .IN1(n10257), .IN2(U6439_n1), .QN(WX794) );
  INVX0 U6440_U2 ( .INP(WX729), .ZN(U6440_n1) );
  NOR2X0 U6440_U1 ( .IN1(n10257), .IN2(U6440_n1), .QN(WX792) );
  INVX0 U6441_U2 ( .INP(WX727), .ZN(U6441_n1) );
  NOR2X0 U6441_U1 ( .IN1(n10257), .IN2(U6441_n1), .QN(WX790) );
  INVX0 U6442_U2 ( .INP(WX725), .ZN(U6442_n1) );
  NOR2X0 U6442_U1 ( .IN1(n10257), .IN2(U6442_n1), .QN(WX788) );
  INVX0 U6443_U2 ( .INP(test_so4), .ZN(U6443_n1) );
  NOR2X0 U6443_U1 ( .IN1(n10257), .IN2(U6443_n1), .QN(WX786) );
  INVX0 U6444_U2 ( .INP(WX721), .ZN(U6444_n1) );
  NOR2X0 U6444_U1 ( .IN1(n10257), .IN2(U6444_n1), .QN(WX784) );
  INVX0 U6445_U2 ( .INP(WX719), .ZN(U6445_n1) );
  NOR2X0 U6445_U1 ( .IN1(n10257), .IN2(U6445_n1), .QN(WX782) );
  INVX0 U6446_U2 ( .INP(WX717), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n10257), .IN2(U6446_n1), .QN(WX780) );
  INVX0 U6447_U2 ( .INP(WX715), .ZN(U6447_n1) );
  NOR2X0 U6447_U1 ( .IN1(n10257), .IN2(U6447_n1), .QN(WX778) );
  INVX0 U6448_U2 ( .INP(WX713), .ZN(U6448_n1) );
  NOR2X0 U6448_U1 ( .IN1(n10257), .IN2(U6448_n1), .QN(WX776) );
  INVX0 U6449_U2 ( .INP(WX711), .ZN(U6449_n1) );
  NOR2X0 U6449_U1 ( .IN1(n10257), .IN2(U6449_n1), .QN(WX774) );
  INVX0 U6450_U2 ( .INP(WX709), .ZN(U6450_n1) );
  NOR2X0 U6450_U1 ( .IN1(n10256), .IN2(U6450_n1), .QN(WX772) );
  INVX0 U6451_U2 ( .INP(WX707), .ZN(U6451_n1) );
  NOR2X0 U6451_U1 ( .IN1(n10256), .IN2(U6451_n1), .QN(WX770) );
  INVX0 U6452_U2 ( .INP(WX705), .ZN(U6452_n1) );
  NOR2X0 U6452_U1 ( .IN1(n10256), .IN2(U6452_n1), .QN(WX768) );
  INVX0 U6453_U2 ( .INP(WX703), .ZN(U6453_n1) );
  NOR2X0 U6453_U1 ( .IN1(n10256), .IN2(U6453_n1), .QN(WX766) );
  INVX0 U6454_U2 ( .INP(WX701), .ZN(U6454_n1) );
  NOR2X0 U6454_U1 ( .IN1(n10256), .IN2(U6454_n1), .QN(WX764) );
  INVX0 U6455_U2 ( .INP(WX699), .ZN(U6455_n1) );
  NOR2X0 U6455_U1 ( .IN1(n10256), .IN2(U6455_n1), .QN(WX762) );
  INVX0 U6456_U2 ( .INP(WX697), .ZN(U6456_n1) );
  NOR2X0 U6456_U1 ( .IN1(n10256), .IN2(U6456_n1), .QN(WX760) );
  INVX0 U6457_U2 ( .INP(WX695), .ZN(U6457_n1) );
  NOR2X0 U6457_U1 ( .IN1(n10256), .IN2(U6457_n1), .QN(WX758) );
  INVX0 U6458_U2 ( .INP(WX693), .ZN(U6458_n1) );
  NOR2X0 U6458_U1 ( .IN1(n10256), .IN2(U6458_n1), .QN(WX756) );
  INVX0 U6459_U2 ( .INP(WX691), .ZN(U6459_n1) );
  NOR2X0 U6459_U1 ( .IN1(n10256), .IN2(U6459_n1), .QN(WX754) );
  INVX0 U6460_U2 ( .INP(WX689), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(n10256), .IN2(U6460_n1), .QN(WX752) );
  INVX0 U6461_U2 ( .INP(test_so3), .ZN(U6461_n1) );
  NOR2X0 U6461_U1 ( .IN1(n10255), .IN2(U6461_n1), .QN(WX750) );
  INVX0 U6462_U2 ( .INP(WX685), .ZN(U6462_n1) );
  NOR2X0 U6462_U1 ( .IN1(n10255), .IN2(U6462_n1), .QN(WX748) );
  INVX0 U6463_U2 ( .INP(WX683), .ZN(U6463_n1) );
  NOR2X0 U6463_U1 ( .IN1(n10255), .IN2(U6463_n1), .QN(WX746) );
  INVX0 U6464_U2 ( .INP(WX681), .ZN(U6464_n1) );
  NOR2X0 U6464_U1 ( .IN1(n10255), .IN2(U6464_n1), .QN(WX744) );
  INVX0 U6465_U2 ( .INP(WX679), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n10255), .IN2(U6465_n1), .QN(WX742) );
  INVX0 U6466_U2 ( .INP(WX677), .ZN(U6466_n1) );
  NOR2X0 U6466_U1 ( .IN1(n10255), .IN2(U6466_n1), .QN(WX740) );
  INVX0 U6467_U2 ( .INP(WX675), .ZN(U6467_n1) );
  NOR2X0 U6467_U1 ( .IN1(n10255), .IN2(U6467_n1), .QN(WX738) );
  INVX0 U6468_U2 ( .INP(WX673), .ZN(U6468_n1) );
  NOR2X0 U6468_U1 ( .IN1(n10255), .IN2(U6468_n1), .QN(WX736) );
  INVX0 U6469_U2 ( .INP(WX671), .ZN(U6469_n1) );
  NOR2X0 U6469_U1 ( .IN1(n10255), .IN2(U6469_n1), .QN(WX734) );
  INVX0 U6470_U2 ( .INP(WX669), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n10255), .IN2(U6470_n1), .QN(WX732) );
  INVX0 U6471_U2 ( .INP(WX667), .ZN(U6471_n1) );
  NOR2X0 U6471_U1 ( .IN1(n10255), .IN2(U6471_n1), .QN(WX730) );
  INVX0 U6472_U2 ( .INP(WX665), .ZN(U6472_n1) );
  NOR2X0 U6472_U1 ( .IN1(n10254), .IN2(U6472_n1), .QN(WX728) );
  INVX0 U6473_U2 ( .INP(WX663), .ZN(U6473_n1) );
  NOR2X0 U6473_U1 ( .IN1(n10254), .IN2(U6473_n1), .QN(WX726) );
  INVX0 U6474_U2 ( .INP(WX661), .ZN(U6474_n1) );
  NOR2X0 U6474_U1 ( .IN1(n10254), .IN2(U6474_n1), .QN(WX724) );
  INVX0 U6475_U2 ( .INP(WX659), .ZN(U6475_n1) );
  NOR2X0 U6475_U1 ( .IN1(n10254), .IN2(U6475_n1), .QN(WX722) );
  INVX0 U6476_U2 ( .INP(WX657), .ZN(U6476_n1) );
  NOR2X0 U6476_U1 ( .IN1(n10254), .IN2(U6476_n1), .QN(WX720) );
  INVX0 U6477_U2 ( .INP(WX655), .ZN(U6477_n1) );
  NOR2X0 U6477_U1 ( .IN1(n10254), .IN2(U6477_n1), .QN(WX718) );
  INVX0 U6478_U2 ( .INP(WX653), .ZN(U6478_n1) );
  NOR2X0 U6478_U1 ( .IN1(n10254), .IN2(U6478_n1), .QN(WX716) );
  INVX0 U6479_U2 ( .INP(test_so2), .ZN(U6479_n1) );
  NOR2X0 U6479_U1 ( .IN1(n10254), .IN2(U6479_n1), .QN(WX714) );
  INVX0 U6480_U2 ( .INP(WX649), .ZN(U6480_n1) );
  NOR2X0 U6480_U1 ( .IN1(n10254), .IN2(U6480_n1), .QN(WX712) );
  INVX0 U6481_U2 ( .INP(WX647), .ZN(U6481_n1) );
  NOR2X0 U6481_U1 ( .IN1(n10254), .IN2(U6481_n1), .QN(WX710) );
  INVX0 U6482_U2 ( .INP(WX645), .ZN(U6482_n1) );
  NOR2X0 U6482_U1 ( .IN1(n10296), .IN2(U6482_n1), .QN(WX708) );
endmodule

