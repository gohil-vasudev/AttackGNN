module add_mul_combine_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, Result_mul_0_, Result_mul_1_, 
        Result_mul_2_, Result_mul_3_, Result_mul_4_, Result_mul_5_, 
        Result_mul_6_, Result_mul_7_, Result_mul_8_, Result_mul_9_, 
        Result_mul_10_, Result_mul_11_, Result_mul_12_, Result_mul_13_, 
        Result_mul_14_, Result_mul_15_, Result_mul_16_, Result_mul_17_, 
        Result_mul_18_, Result_mul_19_, Result_mul_20_, Result_mul_21_, 
        Result_mul_22_, Result_mul_23_, Result_mul_24_, Result_mul_25_, 
        Result_mul_26_, Result_mul_27_, Result_mul_28_, Result_mul_29_, 
        Result_mul_30_, Result_mul_31_, Result_mul_32_, Result_mul_33_, 
        Result_mul_34_, Result_mul_35_, Result_mul_36_, Result_mul_37_, 
        Result_mul_38_, Result_mul_39_, Result_mul_40_, Result_mul_41_, 
        Result_mul_42_, Result_mul_43_, Result_mul_44_, Result_mul_45_, 
        Result_mul_46_, Result_mul_47_, Result_mul_48_, Result_mul_49_, 
        Result_mul_50_, Result_mul_51_, Result_mul_52_, Result_mul_53_, 
        Result_mul_54_, Result_mul_55_, Result_mul_56_, Result_mul_57_, 
        Result_mul_58_, Result_mul_59_, Result_mul_60_, Result_mul_61_, 
        Result_mul_62_, Result_mul_63_, Result_add_0_, Result_add_1_, 
        Result_add_2_, Result_add_3_, Result_add_4_, Result_add_5_, 
        Result_add_6_, Result_add_7_, Result_add_8_, Result_add_9_, 
        Result_add_10_, Result_add_11_, Result_add_12_, Result_add_13_, 
        Result_add_14_, Result_add_15_, Result_add_16_, Result_add_17_, 
        Result_add_18_, Result_add_19_, Result_add_20_, Result_add_21_, 
        Result_add_22_, Result_add_23_, Result_add_24_, Result_add_25_, 
        Result_add_26_, Result_add_27_, Result_add_28_, Result_add_29_, 
        Result_add_30_, Result_add_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_mul_32_, Result_mul_33_, Result_mul_34_, Result_mul_35_,
         Result_mul_36_, Result_mul_37_, Result_mul_38_, Result_mul_39_,
         Result_mul_40_, Result_mul_41_, Result_mul_42_, Result_mul_43_,
         Result_mul_44_, Result_mul_45_, Result_mul_46_, Result_mul_47_,
         Result_mul_48_, Result_mul_49_, Result_mul_50_, Result_mul_51_,
         Result_mul_52_, Result_mul_53_, Result_mul_54_, Result_mul_55_,
         Result_mul_56_, Result_mul_57_, Result_mul_58_, Result_mul_59_,
         Result_mul_60_, Result_mul_61_, Result_mul_62_, Result_mul_63_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_,
         Result_add_16_, Result_add_17_, Result_add_18_, Result_add_19_,
         Result_add_20_, Result_add_21_, Result_add_22_, Result_add_23_,
         Result_add_24_, Result_add_25_, Result_add_26_, Result_add_27_,
         Result_add_28_, Result_add_29_, Result_add_30_, Result_add_31_;
  wire   n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610;

  INV_X2 U7384 ( .A(b_21_), .ZN(n9875) );
  INV_X2 U7385 ( .A(b_29_), .ZN(n8110) );
  INV_X2 U7386 ( .A(b_19_), .ZN(n7909) );
  INV_X2 U7387 ( .A(b_3_), .ZN(n7620) );
  INV_X2 U7388 ( .A(b_5_), .ZN(n7674) );
  INV_X2 U7389 ( .A(b_7_), .ZN(n7755) );
  INV_X2 U7390 ( .A(b_9_), .ZN(n12396) );
  INV_X2 U7391 ( .A(b_11_), .ZN(n11958) );
  INV_X2 U7392 ( .A(b_13_), .ZN(n11530) );
  INV_X2 U7393 ( .A(b_17_), .ZN(n7852) );
  INV_X2 U7394 ( .A(b_15_), .ZN(n11108) );
  XOR2_X1 U7395 ( .A(n7288), .B(n7289), .Z(Result_mul_9_) );
  AND2_X1 U7396 ( .A1(n7290), .A2(n7291), .ZN(n7289) );
  OR2_X1 U7397 ( .A1(n7292), .A2(n7293), .ZN(n7291) );
  AND2_X1 U7398 ( .A1(n7294), .A2(n7295), .ZN(n7293) );
  INV_X1 U7399 ( .A(n7296), .ZN(n7290) );
  XOR2_X1 U7400 ( .A(n7297), .B(n7298), .Z(Result_mul_8_) );
  XOR2_X1 U7401 ( .A(n7299), .B(n7300), .Z(Result_mul_7_) );
  AND2_X1 U7402 ( .A1(n7301), .A2(n7302), .ZN(n7300) );
  OR2_X1 U7403 ( .A1(n7303), .A2(n7304), .ZN(n7302) );
  AND2_X1 U7404 ( .A1(n7305), .A2(n7306), .ZN(n7304) );
  INV_X1 U7405 ( .A(n7307), .ZN(n7301) );
  XOR2_X1 U7406 ( .A(n7308), .B(n7309), .Z(Result_mul_6_) );
  OR2_X1 U7407 ( .A1(n7310), .A2(n7311), .ZN(Result_mul_62_) );
  AND2_X1 U7408 ( .A1(b_31_), .A2(n7312), .ZN(n7311) );
  OR2_X1 U7409 ( .A1(n7313), .A2(n7314), .ZN(n7312) );
  AND2_X1 U7410 ( .A1(a_30_), .A2(n7315), .ZN(n7313) );
  AND2_X1 U7411 ( .A1(b_30_), .A2(n7316), .ZN(n7310) );
  OR2_X1 U7412 ( .A1(n7317), .A2(n7318), .ZN(n7316) );
  AND2_X1 U7413 ( .A1(a_31_), .A2(n7319), .ZN(n7317) );
  XNOR2_X1 U7414 ( .A(n7320), .B(n7321), .ZN(Result_mul_61_) );
  XNOR2_X1 U7415 ( .A(n7322), .B(n7323), .ZN(n7320) );
  XOR2_X1 U7416 ( .A(n7324), .B(n7325), .Z(Result_mul_60_) );
  XNOR2_X1 U7417 ( .A(n7326), .B(n7327), .ZN(n7324) );
  XOR2_X1 U7418 ( .A(n7328), .B(n7329), .Z(Result_mul_5_) );
  AND2_X1 U7419 ( .A1(n7330), .A2(n7331), .ZN(n7329) );
  OR2_X1 U7420 ( .A1(n7332), .A2(n7333), .ZN(n7331) );
  AND2_X1 U7421 ( .A1(n7334), .A2(n7335), .ZN(n7333) );
  INV_X1 U7422 ( .A(n7336), .ZN(n7330) );
  XOR2_X1 U7423 ( .A(n7337), .B(n7338), .Z(Result_mul_59_) );
  XNOR2_X1 U7424 ( .A(n7339), .B(n7340), .ZN(n7337) );
  XOR2_X1 U7425 ( .A(n7341), .B(n7342), .Z(Result_mul_58_) );
  XNOR2_X1 U7426 ( .A(n7343), .B(n7344), .ZN(n7341) );
  XNOR2_X1 U7427 ( .A(n7345), .B(n7346), .ZN(Result_mul_57_) );
  XOR2_X1 U7428 ( .A(n7347), .B(n7348), .Z(n7346) );
  XNOR2_X1 U7429 ( .A(n7349), .B(n7350), .ZN(Result_mul_56_) );
  XOR2_X1 U7430 ( .A(n7351), .B(n7352), .Z(n7350) );
  XNOR2_X1 U7431 ( .A(n7353), .B(n7354), .ZN(Result_mul_55_) );
  XOR2_X1 U7432 ( .A(n7355), .B(n7356), .Z(n7354) );
  XNOR2_X1 U7433 ( .A(n7357), .B(n7358), .ZN(Result_mul_54_) );
  XOR2_X1 U7434 ( .A(n7359), .B(n7360), .Z(n7358) );
  XNOR2_X1 U7435 ( .A(n7361), .B(n7362), .ZN(Result_mul_53_) );
  XOR2_X1 U7436 ( .A(n7363), .B(n7364), .Z(n7362) );
  XNOR2_X1 U7437 ( .A(n7365), .B(n7366), .ZN(Result_mul_52_) );
  XOR2_X1 U7438 ( .A(n7367), .B(n7368), .Z(n7366) );
  XNOR2_X1 U7439 ( .A(n7369), .B(n7370), .ZN(Result_mul_51_) );
  XOR2_X1 U7440 ( .A(n7371), .B(n7372), .Z(n7370) );
  XNOR2_X1 U7441 ( .A(n7373), .B(n7374), .ZN(Result_mul_50_) );
  XOR2_X1 U7442 ( .A(n7375), .B(n7376), .Z(n7374) );
  XOR2_X1 U7443 ( .A(n7377), .B(n7378), .Z(Result_mul_4_) );
  XNOR2_X1 U7444 ( .A(n7379), .B(n7380), .ZN(Result_mul_49_) );
  XOR2_X1 U7445 ( .A(n7381), .B(n7382), .Z(n7380) );
  XNOR2_X1 U7446 ( .A(n7383), .B(n7384), .ZN(Result_mul_48_) );
  XOR2_X1 U7447 ( .A(n7385), .B(n7386), .Z(n7384) );
  XNOR2_X1 U7448 ( .A(n7387), .B(n7388), .ZN(Result_mul_47_) );
  XOR2_X1 U7449 ( .A(n7389), .B(n7390), .Z(n7388) );
  XNOR2_X1 U7450 ( .A(n7391), .B(n7392), .ZN(Result_mul_46_) );
  XOR2_X1 U7451 ( .A(n7393), .B(n7394), .Z(n7392) );
  XNOR2_X1 U7452 ( .A(n7395), .B(n7396), .ZN(Result_mul_45_) );
  XOR2_X1 U7453 ( .A(n7397), .B(n7398), .Z(n7396) );
  XNOR2_X1 U7454 ( .A(n7399), .B(n7400), .ZN(Result_mul_44_) );
  XOR2_X1 U7455 ( .A(n7401), .B(n7402), .Z(n7400) );
  XNOR2_X1 U7456 ( .A(n7403), .B(n7404), .ZN(Result_mul_43_) );
  XOR2_X1 U7457 ( .A(n7405), .B(n7406), .Z(n7404) );
  XNOR2_X1 U7458 ( .A(n7407), .B(n7408), .ZN(Result_mul_42_) );
  XOR2_X1 U7459 ( .A(n7409), .B(n7410), .Z(n7408) );
  XNOR2_X1 U7460 ( .A(n7411), .B(n7412), .ZN(Result_mul_41_) );
  XOR2_X1 U7461 ( .A(n7413), .B(n7414), .Z(n7412) );
  XNOR2_X1 U7462 ( .A(n7415), .B(n7416), .ZN(Result_mul_40_) );
  XOR2_X1 U7463 ( .A(n7417), .B(n7418), .Z(n7416) );
  XOR2_X1 U7464 ( .A(n7419), .B(n7420), .Z(Result_mul_3_) );
  AND2_X1 U7465 ( .A1(n7421), .A2(n7422), .ZN(n7420) );
  OR2_X1 U7466 ( .A1(n7423), .A2(n7424), .ZN(n7422) );
  AND2_X1 U7467 ( .A1(n7425), .A2(n7426), .ZN(n7424) );
  INV_X1 U7468 ( .A(n7427), .ZN(n7421) );
  XNOR2_X1 U7469 ( .A(n7428), .B(n7429), .ZN(Result_mul_39_) );
  XOR2_X1 U7470 ( .A(n7430), .B(n7431), .Z(n7429) );
  XNOR2_X1 U7471 ( .A(n7432), .B(n7433), .ZN(Result_mul_38_) );
  XOR2_X1 U7472 ( .A(n7434), .B(n7435), .Z(n7433) );
  XNOR2_X1 U7473 ( .A(n7436), .B(n7437), .ZN(Result_mul_37_) );
  XOR2_X1 U7474 ( .A(n7438), .B(n7439), .Z(n7437) );
  XNOR2_X1 U7475 ( .A(n7440), .B(n7441), .ZN(Result_mul_36_) );
  XOR2_X1 U7476 ( .A(n7442), .B(n7443), .Z(n7441) );
  XNOR2_X1 U7477 ( .A(n7444), .B(n7445), .ZN(Result_mul_35_) );
  XOR2_X1 U7478 ( .A(n7446), .B(n7447), .Z(n7445) );
  XNOR2_X1 U7479 ( .A(n7448), .B(n7449), .ZN(Result_mul_34_) );
  XOR2_X1 U7480 ( .A(n7450), .B(n7451), .Z(n7449) );
  XNOR2_X1 U7481 ( .A(n7452), .B(n7453), .ZN(Result_mul_33_) );
  XOR2_X1 U7482 ( .A(n7454), .B(n7455), .Z(n7453) );
  XNOR2_X1 U7483 ( .A(n7456), .B(n7457), .ZN(Result_mul_32_) );
  XOR2_X1 U7484 ( .A(n7458), .B(n7459), .Z(n7457) );
  XNOR2_X1 U7485 ( .A(n7460), .B(n7461), .ZN(Result_mul_31_) );
  AND2_X1 U7486 ( .A1(n7462), .A2(n7463), .ZN(Result_mul_30_) );
  OR2_X1 U7487 ( .A1(n7464), .A2(n7465), .ZN(n7462) );
  AND2_X1 U7488 ( .A1(n7466), .A2(n7461), .ZN(n7464) );
  XOR2_X1 U7489 ( .A(n7467), .B(n7468), .Z(Result_mul_2_) );
  XNOR2_X1 U7490 ( .A(n7463), .B(n7469), .ZN(Result_mul_29_) );
  AND2_X1 U7491 ( .A1(n7470), .A2(n7471), .ZN(n7469) );
  INV_X1 U7492 ( .A(n7472), .ZN(n7463) );
  XOR2_X1 U7493 ( .A(n7473), .B(n7474), .Z(Result_mul_28_) );
  AND2_X1 U7494 ( .A1(n7475), .A2(n7476), .ZN(n7474) );
  INV_X1 U7495 ( .A(n7477), .ZN(n7476) );
  XOR2_X1 U7496 ( .A(n7478), .B(n7479), .Z(Result_mul_27_) );
  AND2_X1 U7497 ( .A1(n7480), .A2(n7481), .ZN(n7479) );
  INV_X1 U7498 ( .A(n7482), .ZN(n7481) );
  XOR2_X1 U7499 ( .A(n7483), .B(n7484), .Z(Result_mul_26_) );
  AND2_X1 U7500 ( .A1(n7485), .A2(n7486), .ZN(n7484) );
  INV_X1 U7501 ( .A(n7487), .ZN(n7486) );
  XOR2_X1 U7502 ( .A(n7488), .B(n7489), .Z(Result_mul_25_) );
  AND2_X1 U7503 ( .A1(n7490), .A2(n7491), .ZN(n7489) );
  INV_X1 U7504 ( .A(n7492), .ZN(n7490) );
  XOR2_X1 U7505 ( .A(n7493), .B(n7494), .Z(Result_mul_24_) );
  AND2_X1 U7506 ( .A1(n7495), .A2(n7496), .ZN(n7494) );
  XOR2_X1 U7507 ( .A(n7497), .B(n7498), .Z(Result_mul_23_) );
  AND2_X1 U7508 ( .A1(n7499), .A2(n7500), .ZN(n7498) );
  XOR2_X1 U7509 ( .A(n7501), .B(n7502), .Z(Result_mul_22_) );
  AND2_X1 U7510 ( .A1(n7503), .A2(n7504), .ZN(n7502) );
  XOR2_X1 U7511 ( .A(n7505), .B(n7506), .Z(Result_mul_21_) );
  AND2_X1 U7512 ( .A1(n7507), .A2(n7508), .ZN(n7506) );
  INV_X1 U7513 ( .A(n7509), .ZN(n7507) );
  XOR2_X1 U7514 ( .A(n7510), .B(n7511), .Z(Result_mul_20_) );
  AND2_X1 U7515 ( .A1(n7512), .A2(n7513), .ZN(n7511) );
  XOR2_X1 U7516 ( .A(n7514), .B(n7515), .Z(Result_mul_1_) );
  AND2_X1 U7517 ( .A1(n7516), .A2(n7517), .ZN(n7515) );
  OR2_X1 U7518 ( .A1(n7518), .A2(n7519), .ZN(n7517) );
  AND2_X1 U7519 ( .A1(n7520), .A2(n7521), .ZN(n7518) );
  INV_X1 U7520 ( .A(n7522), .ZN(n7516) );
  XOR2_X1 U7521 ( .A(n7523), .B(n7524), .Z(Result_mul_19_) );
  AND2_X1 U7522 ( .A1(n7525), .A2(n7526), .ZN(n7524) );
  XOR2_X1 U7523 ( .A(n7527), .B(n7528), .Z(Result_mul_18_) );
  AND2_X1 U7524 ( .A1(n7529), .A2(n7530), .ZN(n7528) );
  XOR2_X1 U7525 ( .A(n7531), .B(n7532), .Z(Result_mul_17_) );
  AND2_X1 U7526 ( .A1(n7533), .A2(n7534), .ZN(n7532) );
  XOR2_X1 U7527 ( .A(n7535), .B(n7536), .Z(Result_mul_16_) );
  AND2_X1 U7528 ( .A1(n7537), .A2(n7538), .ZN(n7536) );
  XOR2_X1 U7529 ( .A(n7539), .B(n7540), .Z(Result_mul_15_) );
  AND2_X1 U7530 ( .A1(n7541), .A2(n7542), .ZN(n7540) );
  INV_X1 U7531 ( .A(n7543), .ZN(n7542) );
  XOR2_X1 U7532 ( .A(n7544), .B(n7545), .Z(Result_mul_14_) );
  AND2_X1 U7533 ( .A1(n7546), .A2(n7547), .ZN(n7545) );
  INV_X1 U7534 ( .A(n7548), .ZN(n7547) );
  OR2_X1 U7535 ( .A1(n7549), .A2(n7550), .ZN(n7546) );
  AND2_X1 U7536 ( .A1(n7551), .A2(n7552), .ZN(n7549) );
  XOR2_X1 U7537 ( .A(n7553), .B(n7554), .Z(Result_mul_13_) );
  AND2_X1 U7538 ( .A1(n7555), .A2(n7556), .ZN(n7554) );
  INV_X1 U7539 ( .A(n7557), .ZN(n7556) );
  OR2_X1 U7540 ( .A1(n7558), .A2(n7559), .ZN(n7555) );
  AND2_X1 U7541 ( .A1(n7560), .A2(n7561), .ZN(n7558) );
  XOR2_X1 U7542 ( .A(n7562), .B(n7563), .Z(Result_mul_12_) );
  AND2_X1 U7543 ( .A1(n7564), .A2(n7565), .ZN(n7563) );
  INV_X1 U7544 ( .A(n7566), .ZN(n7565) );
  OR2_X1 U7545 ( .A1(n7567), .A2(n7568), .ZN(n7564) );
  AND2_X1 U7546 ( .A1(n7569), .A2(n7570), .ZN(n7567) );
  XOR2_X1 U7547 ( .A(n7571), .B(n7572), .Z(Result_mul_11_) );
  AND2_X1 U7548 ( .A1(n7573), .A2(n7574), .ZN(n7572) );
  INV_X1 U7549 ( .A(n7575), .ZN(n7574) );
  OR2_X1 U7550 ( .A1(n7576), .A2(n7577), .ZN(n7573) );
  AND2_X1 U7551 ( .A1(n7578), .A2(n7579), .ZN(n7576) );
  XOR2_X1 U7552 ( .A(n7580), .B(n7581), .Z(Result_mul_10_) );
  AND2_X1 U7553 ( .A1(n7582), .A2(n7583), .ZN(n7581) );
  INV_X1 U7554 ( .A(n7584), .ZN(n7583) );
  OR2_X1 U7555 ( .A1(n7585), .A2(n7586), .ZN(n7582) );
  AND2_X1 U7556 ( .A1(n7587), .A2(n7588), .ZN(n7585) );
  OR3_X1 U7557 ( .A1(n7522), .A2(n7589), .A3(n7590), .ZN(Result_mul_0_) );
  AND2_X1 U7558 ( .A1(n7591), .A2(a_0_), .ZN(n7590) );
  INV_X1 U7559 ( .A(n7592), .ZN(n7591) );
  AND2_X1 U7560 ( .A1(n7514), .A2(n7519), .ZN(n7589) );
  AND2_X1 U7561 ( .A1(n7467), .A2(n7468), .ZN(n7514) );
  XNOR2_X1 U7562 ( .A(n7521), .B(n7593), .ZN(n7468) );
  OR2_X1 U7563 ( .A1(n7594), .A2(n7595), .ZN(n7467) );
  OR2_X1 U7564 ( .A1(n7596), .A2(n7427), .ZN(n7594) );
  AND3_X1 U7565 ( .A1(n7426), .A2(n7425), .A3(n7423), .ZN(n7427) );
  INV_X1 U7566 ( .A(n7597), .ZN(n7425) );
  AND2_X1 U7567 ( .A1(n7419), .A2(n7423), .ZN(n7596) );
  INV_X1 U7568 ( .A(n7598), .ZN(n7423) );
  OR2_X1 U7569 ( .A1(n7599), .A2(n7595), .ZN(n7598) );
  INV_X1 U7570 ( .A(n7600), .ZN(n7595) );
  OR2_X1 U7571 ( .A1(n7601), .A2(n7602), .ZN(n7600) );
  AND2_X1 U7572 ( .A1(n7601), .A2(n7602), .ZN(n7599) );
  OR2_X1 U7573 ( .A1(n7603), .A2(n7604), .ZN(n7602) );
  AND2_X1 U7574 ( .A1(n7605), .A2(n7606), .ZN(n7604) );
  AND2_X1 U7575 ( .A1(n7607), .A2(n7608), .ZN(n7603) );
  OR2_X1 U7576 ( .A1(n7606), .A2(n7605), .ZN(n7608) );
  XOR2_X1 U7577 ( .A(n7609), .B(n7610), .Z(n7601) );
  XOR2_X1 U7578 ( .A(n7611), .B(n7612), .Z(n7610) );
  AND2_X1 U7579 ( .A1(n7377), .A2(n7378), .ZN(n7419) );
  XNOR2_X1 U7580 ( .A(n7426), .B(n7597), .ZN(n7378) );
  OR2_X1 U7581 ( .A1(n7613), .A2(n7614), .ZN(n7597) );
  AND2_X1 U7582 ( .A1(n7615), .A2(n7616), .ZN(n7614) );
  AND2_X1 U7583 ( .A1(n7617), .A2(n7618), .ZN(n7613) );
  OR2_X1 U7584 ( .A1(n7616), .A2(n7615), .ZN(n7618) );
  XNOR2_X1 U7585 ( .A(n7607), .B(n7619), .ZN(n7426) );
  XOR2_X1 U7586 ( .A(n7606), .B(n7605), .Z(n7619) );
  OR2_X1 U7587 ( .A1(n7620), .A2(n7621), .ZN(n7605) );
  OR2_X1 U7588 ( .A1(n7622), .A2(n7623), .ZN(n7606) );
  AND2_X1 U7589 ( .A1(n7624), .A2(n7625), .ZN(n7623) );
  AND2_X1 U7590 ( .A1(n7626), .A2(n7627), .ZN(n7622) );
  OR2_X1 U7591 ( .A1(n7625), .A2(n7624), .ZN(n7627) );
  XOR2_X1 U7592 ( .A(n7628), .B(n7629), .Z(n7607) );
  XOR2_X1 U7593 ( .A(n7630), .B(n7631), .Z(n7629) );
  OR2_X1 U7594 ( .A1(n7632), .A2(n7633), .ZN(n7377) );
  OR2_X1 U7595 ( .A1(n7634), .A2(n7336), .ZN(n7632) );
  AND3_X1 U7596 ( .A1(n7335), .A2(n7334), .A3(n7332), .ZN(n7336) );
  INV_X1 U7597 ( .A(n7635), .ZN(n7334) );
  AND2_X1 U7598 ( .A1(n7328), .A2(n7332), .ZN(n7634) );
  INV_X1 U7599 ( .A(n7636), .ZN(n7332) );
  OR2_X1 U7600 ( .A1(n7637), .A2(n7633), .ZN(n7636) );
  INV_X1 U7601 ( .A(n7638), .ZN(n7633) );
  OR2_X1 U7602 ( .A1(n7639), .A2(n7640), .ZN(n7638) );
  AND2_X1 U7603 ( .A1(n7639), .A2(n7640), .ZN(n7637) );
  OR2_X1 U7604 ( .A1(n7641), .A2(n7642), .ZN(n7640) );
  AND2_X1 U7605 ( .A1(n7643), .A2(n7644), .ZN(n7642) );
  AND2_X1 U7606 ( .A1(n7645), .A2(n7646), .ZN(n7641) );
  OR2_X1 U7607 ( .A1(n7644), .A2(n7643), .ZN(n7646) );
  XOR2_X1 U7608 ( .A(n7617), .B(n7647), .Z(n7639) );
  XOR2_X1 U7609 ( .A(n7616), .B(n7615), .Z(n7647) );
  OR2_X1 U7610 ( .A1(n7648), .A2(n7621), .ZN(n7615) );
  OR2_X1 U7611 ( .A1(n7649), .A2(n7650), .ZN(n7616) );
  AND2_X1 U7612 ( .A1(n7651), .A2(n7652), .ZN(n7650) );
  AND2_X1 U7613 ( .A1(n7653), .A2(n7654), .ZN(n7649) );
  OR2_X1 U7614 ( .A1(n7652), .A2(n7651), .ZN(n7654) );
  XOR2_X1 U7615 ( .A(n7626), .B(n7655), .Z(n7617) );
  XOR2_X1 U7616 ( .A(n7625), .B(n7624), .Z(n7655) );
  OR2_X1 U7617 ( .A1(n7620), .A2(n7656), .ZN(n7624) );
  OR2_X1 U7618 ( .A1(n7657), .A2(n7658), .ZN(n7625) );
  AND2_X1 U7619 ( .A1(n7659), .A2(n7660), .ZN(n7658) );
  AND2_X1 U7620 ( .A1(n7661), .A2(n7662), .ZN(n7657) );
  OR2_X1 U7621 ( .A1(n7660), .A2(n7659), .ZN(n7662) );
  XNOR2_X1 U7622 ( .A(n7663), .B(n7664), .ZN(n7626) );
  XNOR2_X1 U7623 ( .A(n7665), .B(n7666), .ZN(n7663) );
  AND2_X1 U7624 ( .A1(n7308), .A2(n7309), .ZN(n7328) );
  XNOR2_X1 U7625 ( .A(n7335), .B(n7635), .ZN(n7309) );
  OR2_X1 U7626 ( .A1(n7667), .A2(n7668), .ZN(n7635) );
  AND2_X1 U7627 ( .A1(n7669), .A2(n7670), .ZN(n7668) );
  AND2_X1 U7628 ( .A1(n7671), .A2(n7672), .ZN(n7667) );
  OR2_X1 U7629 ( .A1(n7670), .A2(n7669), .ZN(n7672) );
  XNOR2_X1 U7630 ( .A(n7645), .B(n7673), .ZN(n7335) );
  XOR2_X1 U7631 ( .A(n7644), .B(n7643), .Z(n7673) );
  OR2_X1 U7632 ( .A1(n7674), .A2(n7621), .ZN(n7643) );
  OR2_X1 U7633 ( .A1(n7675), .A2(n7676), .ZN(n7644) );
  AND2_X1 U7634 ( .A1(n7677), .A2(n7678), .ZN(n7676) );
  AND2_X1 U7635 ( .A1(n7679), .A2(n7680), .ZN(n7675) );
  OR2_X1 U7636 ( .A1(n7678), .A2(n7677), .ZN(n7680) );
  XOR2_X1 U7637 ( .A(n7653), .B(n7681), .Z(n7645) );
  XOR2_X1 U7638 ( .A(n7652), .B(n7651), .Z(n7681) );
  OR2_X1 U7639 ( .A1(n7648), .A2(n7656), .ZN(n7651) );
  OR2_X1 U7640 ( .A1(n7682), .A2(n7683), .ZN(n7652) );
  AND2_X1 U7641 ( .A1(n7684), .A2(n7685), .ZN(n7683) );
  AND2_X1 U7642 ( .A1(n7686), .A2(n7687), .ZN(n7682) );
  OR2_X1 U7643 ( .A1(n7685), .A2(n7684), .ZN(n7687) );
  XOR2_X1 U7644 ( .A(n7661), .B(n7688), .Z(n7653) );
  XOR2_X1 U7645 ( .A(n7660), .B(n7659), .Z(n7688) );
  OR2_X1 U7646 ( .A1(n7620), .A2(n7689), .ZN(n7659) );
  OR2_X1 U7647 ( .A1(n7690), .A2(n7691), .ZN(n7660) );
  AND2_X1 U7648 ( .A1(n7692), .A2(n7693), .ZN(n7691) );
  AND2_X1 U7649 ( .A1(n7694), .A2(n7695), .ZN(n7690) );
  OR2_X1 U7650 ( .A1(n7692), .A2(n7693), .ZN(n7694) );
  XOR2_X1 U7651 ( .A(n7696), .B(n7697), .Z(n7661) );
  XOR2_X1 U7652 ( .A(n7698), .B(n7699), .Z(n7697) );
  OR2_X1 U7653 ( .A1(n7700), .A2(n7701), .ZN(n7308) );
  OR2_X1 U7654 ( .A1(n7702), .A2(n7307), .ZN(n7700) );
  AND3_X1 U7655 ( .A1(n7306), .A2(n7305), .A3(n7303), .ZN(n7307) );
  INV_X1 U7656 ( .A(n7703), .ZN(n7305) );
  AND2_X1 U7657 ( .A1(n7299), .A2(n7303), .ZN(n7702) );
  INV_X1 U7658 ( .A(n7704), .ZN(n7303) );
  OR2_X1 U7659 ( .A1(n7705), .A2(n7701), .ZN(n7704) );
  INV_X1 U7660 ( .A(n7706), .ZN(n7701) );
  OR2_X1 U7661 ( .A1(n7707), .A2(n7708), .ZN(n7706) );
  AND2_X1 U7662 ( .A1(n7707), .A2(n7708), .ZN(n7705) );
  OR2_X1 U7663 ( .A1(n7709), .A2(n7710), .ZN(n7708) );
  AND2_X1 U7664 ( .A1(n7711), .A2(n7712), .ZN(n7710) );
  AND2_X1 U7665 ( .A1(n7713), .A2(n7714), .ZN(n7709) );
  OR2_X1 U7666 ( .A1(n7712), .A2(n7711), .ZN(n7714) );
  XOR2_X1 U7667 ( .A(n7671), .B(n7715), .Z(n7707) );
  XOR2_X1 U7668 ( .A(n7670), .B(n7669), .Z(n7715) );
  OR2_X1 U7669 ( .A1(n7716), .A2(n7621), .ZN(n7669) );
  OR2_X1 U7670 ( .A1(n7717), .A2(n7718), .ZN(n7670) );
  AND2_X1 U7671 ( .A1(n7719), .A2(n7720), .ZN(n7718) );
  AND2_X1 U7672 ( .A1(n7721), .A2(n7722), .ZN(n7717) );
  OR2_X1 U7673 ( .A1(n7720), .A2(n7719), .ZN(n7722) );
  XOR2_X1 U7674 ( .A(n7679), .B(n7723), .Z(n7671) );
  XOR2_X1 U7675 ( .A(n7678), .B(n7677), .Z(n7723) );
  OR2_X1 U7676 ( .A1(n7674), .A2(n7656), .ZN(n7677) );
  OR2_X1 U7677 ( .A1(n7724), .A2(n7725), .ZN(n7678) );
  AND2_X1 U7678 ( .A1(n7726), .A2(n7727), .ZN(n7725) );
  AND2_X1 U7679 ( .A1(n7728), .A2(n7729), .ZN(n7724) );
  OR2_X1 U7680 ( .A1(n7727), .A2(n7726), .ZN(n7729) );
  XOR2_X1 U7681 ( .A(n7686), .B(n7730), .Z(n7679) );
  XOR2_X1 U7682 ( .A(n7685), .B(n7684), .Z(n7730) );
  OR2_X1 U7683 ( .A1(n7648), .A2(n7689), .ZN(n7684) );
  OR2_X1 U7684 ( .A1(n7731), .A2(n7732), .ZN(n7685) );
  AND2_X1 U7685 ( .A1(n7733), .A2(n7734), .ZN(n7732) );
  AND2_X1 U7686 ( .A1(n7735), .A2(n7736), .ZN(n7731) );
  OR2_X1 U7687 ( .A1(n7734), .A2(n7733), .ZN(n7736) );
  XNOR2_X1 U7688 ( .A(n7737), .B(n7692), .ZN(n7686) );
  XOR2_X1 U7689 ( .A(n7738), .B(n7739), .Z(n7692) );
  XOR2_X1 U7690 ( .A(n7740), .B(n7741), .Z(n7739) );
  XNOR2_X1 U7691 ( .A(n7695), .B(n7693), .ZN(n7737) );
  OR2_X1 U7692 ( .A1(n7742), .A2(n7743), .ZN(n7693) );
  AND2_X1 U7693 ( .A1(n7744), .A2(n7745), .ZN(n7743) );
  AND2_X1 U7694 ( .A1(n7746), .A2(n7747), .ZN(n7742) );
  OR2_X1 U7695 ( .A1(n7745), .A2(n7744), .ZN(n7747) );
  AND2_X1 U7696 ( .A1(n7297), .A2(n7298), .ZN(n7299) );
  XNOR2_X1 U7697 ( .A(n7306), .B(n7703), .ZN(n7298) );
  OR2_X1 U7698 ( .A1(n7748), .A2(n7749), .ZN(n7703) );
  AND2_X1 U7699 ( .A1(n7750), .A2(n7751), .ZN(n7749) );
  AND2_X1 U7700 ( .A1(n7752), .A2(n7753), .ZN(n7748) );
  OR2_X1 U7701 ( .A1(n7751), .A2(n7750), .ZN(n7753) );
  XNOR2_X1 U7702 ( .A(n7713), .B(n7754), .ZN(n7306) );
  XOR2_X1 U7703 ( .A(n7712), .B(n7711), .Z(n7754) );
  OR2_X1 U7704 ( .A1(n7755), .A2(n7621), .ZN(n7711) );
  OR2_X1 U7705 ( .A1(n7756), .A2(n7757), .ZN(n7712) );
  AND2_X1 U7706 ( .A1(n7758), .A2(n7759), .ZN(n7757) );
  AND2_X1 U7707 ( .A1(n7760), .A2(n7761), .ZN(n7756) );
  OR2_X1 U7708 ( .A1(n7759), .A2(n7758), .ZN(n7761) );
  XOR2_X1 U7709 ( .A(n7721), .B(n7762), .Z(n7713) );
  XOR2_X1 U7710 ( .A(n7720), .B(n7719), .Z(n7762) );
  OR2_X1 U7711 ( .A1(n7716), .A2(n7656), .ZN(n7719) );
  OR2_X1 U7712 ( .A1(n7763), .A2(n7764), .ZN(n7720) );
  AND2_X1 U7713 ( .A1(n7765), .A2(n7766), .ZN(n7764) );
  AND2_X1 U7714 ( .A1(n7767), .A2(n7768), .ZN(n7763) );
  OR2_X1 U7715 ( .A1(n7766), .A2(n7765), .ZN(n7768) );
  XOR2_X1 U7716 ( .A(n7728), .B(n7769), .Z(n7721) );
  XOR2_X1 U7717 ( .A(n7727), .B(n7726), .Z(n7769) );
  OR2_X1 U7718 ( .A1(n7674), .A2(n7689), .ZN(n7726) );
  OR2_X1 U7719 ( .A1(n7770), .A2(n7771), .ZN(n7727) );
  AND2_X1 U7720 ( .A1(n7772), .A2(n7773), .ZN(n7771) );
  AND2_X1 U7721 ( .A1(n7774), .A2(n7775), .ZN(n7770) );
  OR2_X1 U7722 ( .A1(n7773), .A2(n7772), .ZN(n7775) );
  XOR2_X1 U7723 ( .A(n7735), .B(n7776), .Z(n7728) );
  XOR2_X1 U7724 ( .A(n7734), .B(n7733), .Z(n7776) );
  OR2_X1 U7725 ( .A1(n7648), .A2(n7777), .ZN(n7733) );
  OR2_X1 U7726 ( .A1(n7778), .A2(n7779), .ZN(n7734) );
  AND2_X1 U7727 ( .A1(n7780), .A2(n7781), .ZN(n7779) );
  AND2_X1 U7728 ( .A1(n7782), .A2(n7783), .ZN(n7778) );
  OR2_X1 U7729 ( .A1(n7780), .A2(n7781), .ZN(n7782) );
  XOR2_X1 U7730 ( .A(n7746), .B(n7784), .Z(n7735) );
  XOR2_X1 U7731 ( .A(n7745), .B(n7744), .Z(n7784) );
  OR2_X1 U7732 ( .A1(n7620), .A2(n7785), .ZN(n7744) );
  OR2_X1 U7733 ( .A1(n7786), .A2(n7787), .ZN(n7745) );
  AND2_X1 U7734 ( .A1(n7788), .A2(n7789), .ZN(n7787) );
  AND2_X1 U7735 ( .A1(n7790), .A2(n7791), .ZN(n7786) );
  OR2_X1 U7736 ( .A1(n7789), .A2(n7788), .ZN(n7791) );
  XOR2_X1 U7737 ( .A(n7792), .B(n7793), .Z(n7746) );
  XOR2_X1 U7738 ( .A(n7794), .B(n7795), .Z(n7793) );
  OR2_X1 U7739 ( .A1(n7796), .A2(n7797), .ZN(n7297) );
  OR2_X1 U7740 ( .A1(n7798), .A2(n7296), .ZN(n7796) );
  AND3_X1 U7741 ( .A1(n7295), .A2(n7294), .A3(n7292), .ZN(n7296) );
  INV_X1 U7742 ( .A(n7799), .ZN(n7294) );
  AND2_X1 U7743 ( .A1(n7292), .A2(n7288), .ZN(n7798) );
  OR2_X1 U7744 ( .A1(n7800), .A2(n7584), .ZN(n7288) );
  AND3_X1 U7745 ( .A1(n7588), .A2(n7586), .A3(n7587), .ZN(n7584) );
  INV_X1 U7746 ( .A(n7801), .ZN(n7587) );
  AND2_X1 U7747 ( .A1(n7586), .A2(n7580), .ZN(n7800) );
  OR2_X1 U7748 ( .A1(n7802), .A2(n7575), .ZN(n7580) );
  AND3_X1 U7749 ( .A1(n7579), .A2(n7577), .A3(n7578), .ZN(n7575) );
  INV_X1 U7750 ( .A(n7803), .ZN(n7578) );
  AND2_X1 U7751 ( .A1(n7577), .A2(n7571), .ZN(n7802) );
  OR2_X1 U7752 ( .A1(n7804), .A2(n7566), .ZN(n7571) );
  AND3_X1 U7753 ( .A1(n7570), .A2(n7568), .A3(n7569), .ZN(n7566) );
  INV_X1 U7754 ( .A(n7805), .ZN(n7569) );
  AND2_X1 U7755 ( .A1(n7568), .A2(n7562), .ZN(n7804) );
  OR2_X1 U7756 ( .A1(n7806), .A2(n7557), .ZN(n7562) );
  AND3_X1 U7757 ( .A1(n7561), .A2(n7559), .A3(n7560), .ZN(n7557) );
  INV_X1 U7758 ( .A(n7807), .ZN(n7560) );
  AND2_X1 U7759 ( .A1(n7559), .A2(n7553), .ZN(n7806) );
  OR2_X1 U7760 ( .A1(n7808), .A2(n7548), .ZN(n7553) );
  AND3_X1 U7761 ( .A1(n7552), .A2(n7550), .A3(n7551), .ZN(n7548) );
  INV_X1 U7762 ( .A(n7809), .ZN(n7551) );
  AND2_X1 U7763 ( .A1(n7550), .A2(n7544), .ZN(n7808) );
  OR2_X1 U7764 ( .A1(n7810), .A2(n7543), .ZN(n7544) );
  AND3_X1 U7765 ( .A1(n7811), .A2(n7812), .A3(n7813), .ZN(n7543) );
  AND2_X1 U7766 ( .A1(n7541), .A2(n7539), .ZN(n7810) );
  OR2_X1 U7767 ( .A1(n7814), .A2(n7815), .ZN(n7539) );
  INV_X1 U7768 ( .A(n7537), .ZN(n7815) );
  OR3_X1 U7769 ( .A1(n7816), .A2(n7817), .A3(n7818), .ZN(n7537) );
  AND2_X1 U7770 ( .A1(n7535), .A2(n7538), .ZN(n7814) );
  INV_X1 U7771 ( .A(n7819), .ZN(n7538) );
  AND2_X1 U7772 ( .A1(n7820), .A2(n7817), .ZN(n7819) );
  XNOR2_X1 U7773 ( .A(n7811), .B(n7813), .ZN(n7817) );
  OR2_X1 U7774 ( .A1(n7818), .A2(n7816), .ZN(n7820) );
  OR2_X1 U7775 ( .A1(n7821), .A2(n7822), .ZN(n7535) );
  INV_X1 U7776 ( .A(n7533), .ZN(n7822) );
  OR3_X1 U7777 ( .A1(n7823), .A2(n7824), .A3(n7825), .ZN(n7533) );
  AND2_X1 U7778 ( .A1(n7531), .A2(n7534), .ZN(n7821) );
  INV_X1 U7779 ( .A(n7826), .ZN(n7534) );
  AND2_X1 U7780 ( .A1(n7827), .A2(n7824), .ZN(n7826) );
  XNOR2_X1 U7781 ( .A(n7816), .B(n7818), .ZN(n7824) );
  OR2_X1 U7782 ( .A1(n7828), .A2(n7829), .ZN(n7818) );
  AND2_X1 U7783 ( .A1(n7830), .A2(n7831), .ZN(n7829) );
  AND2_X1 U7784 ( .A1(n7832), .A2(n7833), .ZN(n7828) );
  OR2_X1 U7785 ( .A1(n7830), .A2(n7831), .ZN(n7833) );
  XOR2_X1 U7786 ( .A(n7834), .B(n7835), .Z(n7816) );
  XOR2_X1 U7787 ( .A(n7836), .B(n7837), .Z(n7835) );
  OR2_X1 U7788 ( .A1(n7825), .A2(n7823), .ZN(n7827) );
  OR2_X1 U7789 ( .A1(n7838), .A2(n7839), .ZN(n7531) );
  INV_X1 U7790 ( .A(n7530), .ZN(n7839) );
  OR3_X1 U7791 ( .A1(n7840), .A2(n7841), .A3(n7842), .ZN(n7530) );
  AND2_X1 U7792 ( .A1(n7527), .A2(n7529), .ZN(n7838) );
  INV_X1 U7793 ( .A(n7843), .ZN(n7529) );
  AND2_X1 U7794 ( .A1(n7844), .A2(n7841), .ZN(n7843) );
  XNOR2_X1 U7795 ( .A(n7823), .B(n7825), .ZN(n7841) );
  OR2_X1 U7796 ( .A1(n7845), .A2(n7846), .ZN(n7825) );
  AND2_X1 U7797 ( .A1(n7847), .A2(n7848), .ZN(n7846) );
  AND2_X1 U7798 ( .A1(n7849), .A2(n7850), .ZN(n7845) );
  OR2_X1 U7799 ( .A1(n7847), .A2(n7848), .ZN(n7850) );
  XOR2_X1 U7800 ( .A(n7832), .B(n7851), .Z(n7823) );
  XOR2_X1 U7801 ( .A(n7831), .B(n7830), .Z(n7851) );
  OR2_X1 U7802 ( .A1(n7852), .A2(n7621), .ZN(n7830) );
  OR2_X1 U7803 ( .A1(n7853), .A2(n7854), .ZN(n7831) );
  AND2_X1 U7804 ( .A1(n7855), .A2(n7856), .ZN(n7854) );
  AND2_X1 U7805 ( .A1(n7857), .A2(n7858), .ZN(n7853) );
  OR2_X1 U7806 ( .A1(n7855), .A2(n7856), .ZN(n7858) );
  XOR2_X1 U7807 ( .A(n7859), .B(n7860), .Z(n7832) );
  XOR2_X1 U7808 ( .A(n7861), .B(n7862), .Z(n7860) );
  OR2_X1 U7809 ( .A1(n7842), .A2(n7840), .ZN(n7844) );
  OR2_X1 U7810 ( .A1(n7863), .A2(n7864), .ZN(n7527) );
  INV_X1 U7811 ( .A(n7525), .ZN(n7864) );
  OR3_X1 U7812 ( .A1(n7865), .A2(n7866), .A3(n7867), .ZN(n7525) );
  AND2_X1 U7813 ( .A1(n7523), .A2(n7526), .ZN(n7863) );
  INV_X1 U7814 ( .A(n7868), .ZN(n7526) );
  AND2_X1 U7815 ( .A1(n7869), .A2(n7866), .ZN(n7868) );
  XNOR2_X1 U7816 ( .A(n7840), .B(n7842), .ZN(n7866) );
  OR2_X1 U7817 ( .A1(n7870), .A2(n7871), .ZN(n7842) );
  AND2_X1 U7818 ( .A1(n7872), .A2(n7873), .ZN(n7871) );
  AND2_X1 U7819 ( .A1(n7874), .A2(n7875), .ZN(n7870) );
  OR2_X1 U7820 ( .A1(n7872), .A2(n7873), .ZN(n7875) );
  XOR2_X1 U7821 ( .A(n7849), .B(n7876), .Z(n7840) );
  XOR2_X1 U7822 ( .A(n7848), .B(n7847), .Z(n7876) );
  OR2_X1 U7823 ( .A1(n7621), .A2(n7877), .ZN(n7847) );
  OR2_X1 U7824 ( .A1(n7878), .A2(n7879), .ZN(n7848) );
  AND2_X1 U7825 ( .A1(n7880), .A2(n7881), .ZN(n7879) );
  AND2_X1 U7826 ( .A1(n7882), .A2(n7883), .ZN(n7878) );
  OR2_X1 U7827 ( .A1(n7880), .A2(n7881), .ZN(n7883) );
  XOR2_X1 U7828 ( .A(n7857), .B(n7884), .Z(n7849) );
  XOR2_X1 U7829 ( .A(n7856), .B(n7855), .Z(n7884) );
  OR2_X1 U7830 ( .A1(n7852), .A2(n7656), .ZN(n7855) );
  OR2_X1 U7831 ( .A1(n7885), .A2(n7886), .ZN(n7856) );
  AND2_X1 U7832 ( .A1(n7887), .A2(n7888), .ZN(n7886) );
  AND2_X1 U7833 ( .A1(n7889), .A2(n7890), .ZN(n7885) );
  OR2_X1 U7834 ( .A1(n7887), .A2(n7888), .ZN(n7890) );
  XOR2_X1 U7835 ( .A(n7891), .B(n7892), .Z(n7857) );
  XOR2_X1 U7836 ( .A(n7893), .B(n7894), .Z(n7892) );
  OR2_X1 U7837 ( .A1(n7867), .A2(n7865), .ZN(n7869) );
  OR2_X1 U7838 ( .A1(n7895), .A2(n7896), .ZN(n7523) );
  INV_X1 U7839 ( .A(n7512), .ZN(n7896) );
  OR3_X1 U7840 ( .A1(n7897), .A2(n7898), .A3(n7899), .ZN(n7512) );
  AND2_X1 U7841 ( .A1(n7510), .A2(n7513), .ZN(n7895) );
  INV_X1 U7842 ( .A(n7900), .ZN(n7513) );
  AND2_X1 U7843 ( .A1(n7901), .A2(n7898), .ZN(n7900) );
  XNOR2_X1 U7844 ( .A(n7865), .B(n7867), .ZN(n7898) );
  OR2_X1 U7845 ( .A1(n7902), .A2(n7903), .ZN(n7867) );
  AND2_X1 U7846 ( .A1(n7904), .A2(n7905), .ZN(n7903) );
  AND2_X1 U7847 ( .A1(n7906), .A2(n7907), .ZN(n7902) );
  OR2_X1 U7848 ( .A1(n7904), .A2(n7905), .ZN(n7907) );
  XOR2_X1 U7849 ( .A(n7874), .B(n7908), .Z(n7865) );
  XOR2_X1 U7850 ( .A(n7873), .B(n7872), .Z(n7908) );
  OR2_X1 U7851 ( .A1(n7621), .A2(n7909), .ZN(n7872) );
  OR2_X1 U7852 ( .A1(n7910), .A2(n7911), .ZN(n7873) );
  AND2_X1 U7853 ( .A1(n7912), .A2(n7913), .ZN(n7911) );
  AND2_X1 U7854 ( .A1(n7914), .A2(n7915), .ZN(n7910) );
  OR2_X1 U7855 ( .A1(n7912), .A2(n7913), .ZN(n7915) );
  XOR2_X1 U7856 ( .A(n7882), .B(n7916), .Z(n7874) );
  XOR2_X1 U7857 ( .A(n7881), .B(n7880), .Z(n7916) );
  OR2_X1 U7858 ( .A1(n7656), .A2(n7877), .ZN(n7880) );
  OR2_X1 U7859 ( .A1(n7917), .A2(n7918), .ZN(n7881) );
  AND2_X1 U7860 ( .A1(n7919), .A2(n7920), .ZN(n7918) );
  AND2_X1 U7861 ( .A1(n7921), .A2(n7922), .ZN(n7917) );
  OR2_X1 U7862 ( .A1(n7919), .A2(n7920), .ZN(n7922) );
  XOR2_X1 U7863 ( .A(n7889), .B(n7923), .Z(n7882) );
  XOR2_X1 U7864 ( .A(n7888), .B(n7887), .Z(n7923) );
  OR2_X1 U7865 ( .A1(n7852), .A2(n7689), .ZN(n7887) );
  OR2_X1 U7866 ( .A1(n7924), .A2(n7925), .ZN(n7888) );
  AND2_X1 U7867 ( .A1(n7926), .A2(n7927), .ZN(n7925) );
  AND2_X1 U7868 ( .A1(n7928), .A2(n7929), .ZN(n7924) );
  OR2_X1 U7869 ( .A1(n7926), .A2(n7927), .ZN(n7929) );
  XOR2_X1 U7870 ( .A(n7930), .B(n7931), .Z(n7889) );
  XOR2_X1 U7871 ( .A(n7932), .B(n7933), .Z(n7931) );
  OR2_X1 U7872 ( .A1(n7899), .A2(n7897), .ZN(n7901) );
  OR2_X1 U7873 ( .A1(n7934), .A2(n7509), .ZN(n7510) );
  AND3_X1 U7874 ( .A1(n7935), .A2(n7936), .A3(n7937), .ZN(n7509) );
  AND2_X1 U7875 ( .A1(n7508), .A2(n7505), .ZN(n7934) );
  OR2_X1 U7876 ( .A1(n7938), .A2(n7939), .ZN(n7505) );
  INV_X1 U7877 ( .A(n7504), .ZN(n7939) );
  OR3_X1 U7878 ( .A1(n7940), .A2(n7941), .A3(n7942), .ZN(n7504) );
  AND2_X1 U7879 ( .A1(n7501), .A2(n7503), .ZN(n7938) );
  INV_X1 U7880 ( .A(n7943), .ZN(n7503) );
  AND2_X1 U7881 ( .A1(n7944), .A2(n7941), .ZN(n7943) );
  XNOR2_X1 U7882 ( .A(n7935), .B(n7937), .ZN(n7941) );
  OR2_X1 U7883 ( .A1(n7942), .A2(n7940), .ZN(n7944) );
  OR2_X1 U7884 ( .A1(n7945), .A2(n7946), .ZN(n7501) );
  INV_X1 U7885 ( .A(n7499), .ZN(n7946) );
  OR3_X1 U7886 ( .A1(n7947), .A2(n7948), .A3(n7949), .ZN(n7499) );
  AND2_X1 U7887 ( .A1(n7497), .A2(n7500), .ZN(n7945) );
  INV_X1 U7888 ( .A(n7950), .ZN(n7500) );
  AND2_X1 U7889 ( .A1(n7951), .A2(n7948), .ZN(n7950) );
  XNOR2_X1 U7890 ( .A(n7940), .B(n7942), .ZN(n7948) );
  OR2_X1 U7891 ( .A1(n7952), .A2(n7953), .ZN(n7942) );
  AND2_X1 U7892 ( .A1(n7954), .A2(n7955), .ZN(n7953) );
  AND2_X1 U7893 ( .A1(n7956), .A2(n7957), .ZN(n7952) );
  OR2_X1 U7894 ( .A1(n7954), .A2(n7955), .ZN(n7957) );
  XOR2_X1 U7895 ( .A(n7958), .B(n7959), .Z(n7940) );
  XOR2_X1 U7896 ( .A(n7960), .B(n7961), .Z(n7959) );
  OR2_X1 U7897 ( .A1(n7949), .A2(n7947), .ZN(n7951) );
  OR2_X1 U7898 ( .A1(n7962), .A2(n7963), .ZN(n7497) );
  INV_X1 U7899 ( .A(n7495), .ZN(n7963) );
  OR3_X1 U7900 ( .A1(n7964), .A2(n7965), .A3(n7966), .ZN(n7495) );
  AND2_X1 U7901 ( .A1(n7493), .A2(n7496), .ZN(n7962) );
  INV_X1 U7902 ( .A(n7967), .ZN(n7496) );
  AND2_X1 U7903 ( .A1(n7968), .A2(n7965), .ZN(n7967) );
  XNOR2_X1 U7904 ( .A(n7947), .B(n7949), .ZN(n7965) );
  OR2_X1 U7905 ( .A1(n7969), .A2(n7970), .ZN(n7949) );
  AND2_X1 U7906 ( .A1(n7971), .A2(n7972), .ZN(n7970) );
  AND2_X1 U7907 ( .A1(n7973), .A2(n7974), .ZN(n7969) );
  OR2_X1 U7908 ( .A1(n7971), .A2(n7972), .ZN(n7974) );
  XOR2_X1 U7909 ( .A(n7956), .B(n7975), .Z(n7947) );
  XOR2_X1 U7910 ( .A(n7955), .B(n7954), .Z(n7975) );
  OR2_X1 U7911 ( .A1(n7621), .A2(n7976), .ZN(n7954) );
  OR2_X1 U7912 ( .A1(n7977), .A2(n7978), .ZN(n7955) );
  AND2_X1 U7913 ( .A1(n7979), .A2(n7980), .ZN(n7978) );
  AND2_X1 U7914 ( .A1(n7981), .A2(n7982), .ZN(n7977) );
  OR2_X1 U7915 ( .A1(n7979), .A2(n7980), .ZN(n7982) );
  XOR2_X1 U7916 ( .A(n7983), .B(n7984), .Z(n7956) );
  XOR2_X1 U7917 ( .A(n7985), .B(n7986), .Z(n7984) );
  OR2_X1 U7918 ( .A1(n7966), .A2(n7964), .ZN(n7968) );
  OR2_X1 U7919 ( .A1(n7987), .A2(n7492), .ZN(n7493) );
  AND3_X1 U7920 ( .A1(n7988), .A2(n7989), .A3(n7990), .ZN(n7492) );
  AND2_X1 U7921 ( .A1(n7491), .A2(n7488), .ZN(n7987) );
  OR2_X1 U7922 ( .A1(n7991), .A2(n7487), .ZN(n7488) );
  AND2_X1 U7923 ( .A1(n7992), .A2(n7993), .ZN(n7487) );
  AND2_X1 U7924 ( .A1(n7485), .A2(n7483), .ZN(n7991) );
  OR2_X1 U7925 ( .A1(n7994), .A2(n7482), .ZN(n7483) );
  AND3_X1 U7926 ( .A1(n7995), .A2(n7996), .A3(n7997), .ZN(n7482) );
  AND2_X1 U7927 ( .A1(n7480), .A2(n7478), .ZN(n7994) );
  OR2_X1 U7928 ( .A1(n7998), .A2(n7477), .ZN(n7478) );
  AND3_X1 U7929 ( .A1(n7999), .A2(n8000), .A3(n8001), .ZN(n7477) );
  AND2_X1 U7930 ( .A1(n7475), .A2(n7473), .ZN(n7998) );
  OR2_X1 U7931 ( .A1(n8002), .A2(n8003), .ZN(n7473) );
  INV_X1 U7932 ( .A(n7471), .ZN(n8003) );
  OR3_X1 U7933 ( .A1(n8004), .A2(n8005), .A3(n8006), .ZN(n7471) );
  XNOR2_X1 U7934 ( .A(n7999), .B(n8001), .ZN(n8004) );
  AND2_X1 U7935 ( .A1(n7472), .A2(n7470), .ZN(n8002) );
  OR2_X1 U7936 ( .A1(n8007), .A2(n8008), .ZN(n7470) );
  XNOR2_X1 U7937 ( .A(n8009), .B(n7999), .ZN(n8008) );
  INV_X1 U7938 ( .A(n8010), .ZN(n8007) );
  OR2_X1 U7939 ( .A1(n8006), .A2(n8005), .ZN(n8010) );
  AND3_X1 U7940 ( .A1(n7461), .A2(n7465), .A3(n7466), .ZN(n7472) );
  INV_X1 U7941 ( .A(n7460), .ZN(n7466) );
  OR2_X1 U7942 ( .A1(n8011), .A2(n8012), .ZN(n7460) );
  AND2_X1 U7943 ( .A1(n7459), .A2(n7458), .ZN(n8012) );
  AND2_X1 U7944 ( .A1(n7456), .A2(n8013), .ZN(n8011) );
  OR2_X1 U7945 ( .A1(n7459), .A2(n7458), .ZN(n8013) );
  OR2_X1 U7946 ( .A1(n8014), .A2(n8015), .ZN(n7458) );
  AND2_X1 U7947 ( .A1(n7455), .A2(n7454), .ZN(n8015) );
  AND2_X1 U7948 ( .A1(n7452), .A2(n8016), .ZN(n8014) );
  OR2_X1 U7949 ( .A1(n7455), .A2(n7454), .ZN(n8016) );
  OR2_X1 U7950 ( .A1(n8017), .A2(n8018), .ZN(n7454) );
  AND2_X1 U7951 ( .A1(n7451), .A2(n7450), .ZN(n8018) );
  AND2_X1 U7952 ( .A1(n7448), .A2(n8019), .ZN(n8017) );
  OR2_X1 U7953 ( .A1(n7451), .A2(n7450), .ZN(n8019) );
  OR2_X1 U7954 ( .A1(n8020), .A2(n8021), .ZN(n7450) );
  AND2_X1 U7955 ( .A1(n7447), .A2(n7446), .ZN(n8021) );
  AND2_X1 U7956 ( .A1(n7444), .A2(n8022), .ZN(n8020) );
  OR2_X1 U7957 ( .A1(n7447), .A2(n7446), .ZN(n8022) );
  OR2_X1 U7958 ( .A1(n8023), .A2(n8024), .ZN(n7446) );
  AND2_X1 U7959 ( .A1(n7443), .A2(n7442), .ZN(n8024) );
  AND2_X1 U7960 ( .A1(n7440), .A2(n8025), .ZN(n8023) );
  OR2_X1 U7961 ( .A1(n7443), .A2(n7442), .ZN(n8025) );
  OR2_X1 U7962 ( .A1(n8026), .A2(n8027), .ZN(n7442) );
  AND2_X1 U7963 ( .A1(n7439), .A2(n7438), .ZN(n8027) );
  AND2_X1 U7964 ( .A1(n7436), .A2(n8028), .ZN(n8026) );
  OR2_X1 U7965 ( .A1(n7439), .A2(n7438), .ZN(n8028) );
  OR2_X1 U7966 ( .A1(n8029), .A2(n8030), .ZN(n7438) );
  AND2_X1 U7967 ( .A1(n7435), .A2(n7434), .ZN(n8030) );
  AND2_X1 U7968 ( .A1(n7432), .A2(n8031), .ZN(n8029) );
  OR2_X1 U7969 ( .A1(n7435), .A2(n7434), .ZN(n8031) );
  OR2_X1 U7970 ( .A1(n8032), .A2(n8033), .ZN(n7434) );
  AND2_X1 U7971 ( .A1(n7431), .A2(n7430), .ZN(n8033) );
  AND2_X1 U7972 ( .A1(n7428), .A2(n8034), .ZN(n8032) );
  OR2_X1 U7973 ( .A1(n7431), .A2(n7430), .ZN(n8034) );
  OR2_X1 U7974 ( .A1(n8035), .A2(n8036), .ZN(n7430) );
  AND2_X1 U7975 ( .A1(n7418), .A2(n7417), .ZN(n8036) );
  AND2_X1 U7976 ( .A1(n7415), .A2(n8037), .ZN(n8035) );
  OR2_X1 U7977 ( .A1(n7418), .A2(n7417), .ZN(n8037) );
  OR2_X1 U7978 ( .A1(n8038), .A2(n8039), .ZN(n7417) );
  AND2_X1 U7979 ( .A1(n7414), .A2(n7413), .ZN(n8039) );
  AND2_X1 U7980 ( .A1(n7411), .A2(n8040), .ZN(n8038) );
  OR2_X1 U7981 ( .A1(n7414), .A2(n7413), .ZN(n8040) );
  OR2_X1 U7982 ( .A1(n8041), .A2(n8042), .ZN(n7413) );
  AND2_X1 U7983 ( .A1(n7410), .A2(n7409), .ZN(n8042) );
  AND2_X1 U7984 ( .A1(n7407), .A2(n8043), .ZN(n8041) );
  OR2_X1 U7985 ( .A1(n7410), .A2(n7409), .ZN(n8043) );
  OR2_X1 U7986 ( .A1(n8044), .A2(n8045), .ZN(n7409) );
  AND2_X1 U7987 ( .A1(n7406), .A2(n7405), .ZN(n8045) );
  AND2_X1 U7988 ( .A1(n7403), .A2(n8046), .ZN(n8044) );
  OR2_X1 U7989 ( .A1(n7406), .A2(n7405), .ZN(n8046) );
  OR2_X1 U7990 ( .A1(n8047), .A2(n8048), .ZN(n7405) );
  AND2_X1 U7991 ( .A1(n7402), .A2(n7401), .ZN(n8048) );
  AND2_X1 U7992 ( .A1(n7399), .A2(n8049), .ZN(n8047) );
  OR2_X1 U7993 ( .A1(n7402), .A2(n7401), .ZN(n8049) );
  OR2_X1 U7994 ( .A1(n8050), .A2(n8051), .ZN(n7401) );
  AND2_X1 U7995 ( .A1(n7398), .A2(n7397), .ZN(n8051) );
  AND2_X1 U7996 ( .A1(n7395), .A2(n8052), .ZN(n8050) );
  OR2_X1 U7997 ( .A1(n7398), .A2(n7397), .ZN(n8052) );
  OR2_X1 U7998 ( .A1(n8053), .A2(n8054), .ZN(n7397) );
  AND2_X1 U7999 ( .A1(n7394), .A2(n7393), .ZN(n8054) );
  AND2_X1 U8000 ( .A1(n7391), .A2(n8055), .ZN(n8053) );
  OR2_X1 U8001 ( .A1(n7394), .A2(n7393), .ZN(n8055) );
  OR2_X1 U8002 ( .A1(n8056), .A2(n8057), .ZN(n7393) );
  AND2_X1 U8003 ( .A1(n7390), .A2(n7389), .ZN(n8057) );
  AND2_X1 U8004 ( .A1(n7387), .A2(n8058), .ZN(n8056) );
  OR2_X1 U8005 ( .A1(n7390), .A2(n7389), .ZN(n8058) );
  OR2_X1 U8006 ( .A1(n8059), .A2(n8060), .ZN(n7389) );
  AND2_X1 U8007 ( .A1(n7386), .A2(n7385), .ZN(n8060) );
  AND2_X1 U8008 ( .A1(n7383), .A2(n8061), .ZN(n8059) );
  OR2_X1 U8009 ( .A1(n7386), .A2(n7385), .ZN(n8061) );
  OR2_X1 U8010 ( .A1(n8062), .A2(n8063), .ZN(n7385) );
  AND2_X1 U8011 ( .A1(n7382), .A2(n7381), .ZN(n8063) );
  AND2_X1 U8012 ( .A1(n7379), .A2(n8064), .ZN(n8062) );
  OR2_X1 U8013 ( .A1(n7382), .A2(n7381), .ZN(n8064) );
  OR2_X1 U8014 ( .A1(n8065), .A2(n8066), .ZN(n7381) );
  AND2_X1 U8015 ( .A1(n7376), .A2(n7375), .ZN(n8066) );
  AND2_X1 U8016 ( .A1(n7373), .A2(n8067), .ZN(n8065) );
  OR2_X1 U8017 ( .A1(n7376), .A2(n7375), .ZN(n8067) );
  OR2_X1 U8018 ( .A1(n8068), .A2(n8069), .ZN(n7375) );
  AND2_X1 U8019 ( .A1(n7372), .A2(n7371), .ZN(n8069) );
  AND2_X1 U8020 ( .A1(n7369), .A2(n8070), .ZN(n8068) );
  OR2_X1 U8021 ( .A1(n7372), .A2(n7371), .ZN(n8070) );
  OR2_X1 U8022 ( .A1(n8071), .A2(n8072), .ZN(n7371) );
  AND2_X1 U8023 ( .A1(n7368), .A2(n7367), .ZN(n8072) );
  AND2_X1 U8024 ( .A1(n7365), .A2(n8073), .ZN(n8071) );
  OR2_X1 U8025 ( .A1(n7368), .A2(n7367), .ZN(n8073) );
  OR2_X1 U8026 ( .A1(n8074), .A2(n8075), .ZN(n7367) );
  AND2_X1 U8027 ( .A1(n7364), .A2(n7363), .ZN(n8075) );
  AND2_X1 U8028 ( .A1(n7361), .A2(n8076), .ZN(n8074) );
  OR2_X1 U8029 ( .A1(n7364), .A2(n7363), .ZN(n8076) );
  OR2_X1 U8030 ( .A1(n8077), .A2(n8078), .ZN(n7363) );
  AND2_X1 U8031 ( .A1(n7360), .A2(n7359), .ZN(n8078) );
  AND2_X1 U8032 ( .A1(n7357), .A2(n8079), .ZN(n8077) );
  OR2_X1 U8033 ( .A1(n7360), .A2(n7359), .ZN(n8079) );
  OR2_X1 U8034 ( .A1(n8080), .A2(n8081), .ZN(n7359) );
  AND2_X1 U8035 ( .A1(n7356), .A2(n7355), .ZN(n8081) );
  AND2_X1 U8036 ( .A1(n7353), .A2(n8082), .ZN(n8080) );
  OR2_X1 U8037 ( .A1(n7356), .A2(n7355), .ZN(n8082) );
  OR2_X1 U8038 ( .A1(n8083), .A2(n8084), .ZN(n7355) );
  AND2_X1 U8039 ( .A1(n7352), .A2(n7351), .ZN(n8084) );
  AND2_X1 U8040 ( .A1(n7349), .A2(n8085), .ZN(n8083) );
  OR2_X1 U8041 ( .A1(n7352), .A2(n7351), .ZN(n8085) );
  OR2_X1 U8042 ( .A1(n8086), .A2(n8087), .ZN(n7351) );
  AND2_X1 U8043 ( .A1(n7348), .A2(n7347), .ZN(n8087) );
  AND2_X1 U8044 ( .A1(n7345), .A2(n8088), .ZN(n8086) );
  OR2_X1 U8045 ( .A1(n7348), .A2(n7347), .ZN(n8088) );
  OR2_X1 U8046 ( .A1(n8089), .A2(n8090), .ZN(n7347) );
  AND2_X1 U8047 ( .A1(n7344), .A2(n7343), .ZN(n8090) );
  AND2_X1 U8048 ( .A1(n7342), .A2(n8091), .ZN(n8089) );
  OR2_X1 U8049 ( .A1(n7344), .A2(n7343), .ZN(n8091) );
  OR2_X1 U8050 ( .A1(n8092), .A2(n8093), .ZN(n7343) );
  AND2_X1 U8051 ( .A1(n7340), .A2(n7339), .ZN(n8093) );
  AND2_X1 U8052 ( .A1(n7338), .A2(n8094), .ZN(n8092) );
  OR2_X1 U8053 ( .A1(n7340), .A2(n7339), .ZN(n8094) );
  OR2_X1 U8054 ( .A1(n8095), .A2(n8096), .ZN(n7339) );
  AND2_X1 U8055 ( .A1(n7327), .A2(n7326), .ZN(n8096) );
  AND2_X1 U8056 ( .A1(n7325), .A2(n8097), .ZN(n8095) );
  OR2_X1 U8057 ( .A1(n7327), .A2(n7326), .ZN(n8097) );
  OR2_X1 U8058 ( .A1(n8098), .A2(n8099), .ZN(n7326) );
  AND2_X1 U8059 ( .A1(n7321), .A2(n8100), .ZN(n8099) );
  AND2_X1 U8060 ( .A1(n7323), .A2(n8101), .ZN(n8098) );
  OR2_X1 U8061 ( .A1(n7321), .A2(n8100), .ZN(n8101) );
  INV_X1 U8062 ( .A(n7322), .ZN(n8100) );
  OR2_X1 U8063 ( .A1(n8102), .A2(n7319), .ZN(n7321) );
  INV_X1 U8064 ( .A(n8103), .ZN(n7323) );
  OR3_X1 U8065 ( .A1(n8104), .A2(n8105), .A3(n8106), .ZN(n8103) );
  AND2_X1 U8066 ( .A1(b_30_), .A2(n7314), .ZN(n8106) );
  AND2_X1 U8067 ( .A1(b_29_), .A2(n8107), .ZN(n8105) );
  OR2_X1 U8068 ( .A1(n8108), .A2(n7318), .ZN(n8107) );
  AND2_X1 U8069 ( .A1(a_31_), .A2(n7315), .ZN(n8108) );
  AND2_X1 U8070 ( .A1(n8109), .A2(n8110), .ZN(n8104) );
  OR2_X1 U8071 ( .A1(n8111), .A2(n7319), .ZN(n7327) );
  XNOR2_X1 U8072 ( .A(n8112), .B(n8113), .ZN(n7325) );
  XNOR2_X1 U8073 ( .A(n8114), .B(n8115), .ZN(n8113) );
  OR2_X1 U8074 ( .A1(n8116), .A2(n7319), .ZN(n7340) );
  XOR2_X1 U8075 ( .A(n8117), .B(n8118), .Z(n7338) );
  XOR2_X1 U8076 ( .A(n8119), .B(n8120), .Z(n8118) );
  OR2_X1 U8077 ( .A1(n8121), .A2(n7319), .ZN(n7344) );
  XOR2_X1 U8078 ( .A(n8122), .B(n8123), .Z(n7342) );
  XOR2_X1 U8079 ( .A(n8124), .B(n8125), .Z(n8123) );
  OR2_X1 U8080 ( .A1(n8126), .A2(n7319), .ZN(n7348) );
  XOR2_X1 U8081 ( .A(n8127), .B(n8128), .Z(n7345) );
  XOR2_X1 U8082 ( .A(n8129), .B(n8130), .Z(n8128) );
  OR2_X1 U8083 ( .A1(n8131), .A2(n7319), .ZN(n7352) );
  XOR2_X1 U8084 ( .A(n8132), .B(n8133), .Z(n7349) );
  XOR2_X1 U8085 ( .A(n8134), .B(n8135), .Z(n8133) );
  OR2_X1 U8086 ( .A1(n8136), .A2(n7319), .ZN(n7356) );
  XOR2_X1 U8087 ( .A(n8137), .B(n8138), .Z(n7353) );
  XOR2_X1 U8088 ( .A(n8139), .B(n8140), .Z(n8138) );
  OR2_X1 U8089 ( .A1(n8141), .A2(n7319), .ZN(n7360) );
  XOR2_X1 U8090 ( .A(n8142), .B(n8143), .Z(n7357) );
  XOR2_X1 U8091 ( .A(n8144), .B(n8145), .Z(n8143) );
  OR2_X1 U8092 ( .A1(n8146), .A2(n7319), .ZN(n7364) );
  XOR2_X1 U8093 ( .A(n8147), .B(n8148), .Z(n7361) );
  XOR2_X1 U8094 ( .A(n8149), .B(n8150), .Z(n8148) );
  OR2_X1 U8095 ( .A1(n8151), .A2(n7319), .ZN(n7368) );
  XOR2_X1 U8096 ( .A(n8152), .B(n8153), .Z(n7365) );
  XOR2_X1 U8097 ( .A(n8154), .B(n8155), .Z(n8153) );
  OR2_X1 U8098 ( .A1(n8156), .A2(n7319), .ZN(n7372) );
  XOR2_X1 U8099 ( .A(n8157), .B(n8158), .Z(n7369) );
  XOR2_X1 U8100 ( .A(n8159), .B(n8160), .Z(n8158) );
  OR2_X1 U8101 ( .A1(n8161), .A2(n7319), .ZN(n7376) );
  XOR2_X1 U8102 ( .A(n8162), .B(n8163), .Z(n7373) );
  XOR2_X1 U8103 ( .A(n8164), .B(n8165), .Z(n8163) );
  OR2_X1 U8104 ( .A1(n8166), .A2(n7319), .ZN(n7382) );
  XOR2_X1 U8105 ( .A(n8167), .B(n8168), .Z(n7379) );
  XOR2_X1 U8106 ( .A(n8169), .B(n8170), .Z(n8168) );
  OR2_X1 U8107 ( .A1(n8171), .A2(n7319), .ZN(n7386) );
  XOR2_X1 U8108 ( .A(n8172), .B(n8173), .Z(n7383) );
  XOR2_X1 U8109 ( .A(n8174), .B(n8175), .Z(n8173) );
  OR2_X1 U8110 ( .A1(n8176), .A2(n7319), .ZN(n7390) );
  XOR2_X1 U8111 ( .A(n8177), .B(n8178), .Z(n7387) );
  XOR2_X1 U8112 ( .A(n8179), .B(n8180), .Z(n8178) );
  OR2_X1 U8113 ( .A1(n8181), .A2(n7319), .ZN(n7394) );
  XOR2_X1 U8114 ( .A(n8182), .B(n8183), .Z(n7391) );
  XOR2_X1 U8115 ( .A(n8184), .B(n8185), .Z(n8183) );
  OR2_X1 U8116 ( .A1(n8186), .A2(n7319), .ZN(n7398) );
  XOR2_X1 U8117 ( .A(n8187), .B(n8188), .Z(n7395) );
  XOR2_X1 U8118 ( .A(n8189), .B(n8190), .Z(n8188) );
  OR2_X1 U8119 ( .A1(n8191), .A2(n7319), .ZN(n7402) );
  XOR2_X1 U8120 ( .A(n8192), .B(n8193), .Z(n7399) );
  XOR2_X1 U8121 ( .A(n8194), .B(n8195), .Z(n8193) );
  OR2_X1 U8122 ( .A1(n8196), .A2(n7319), .ZN(n7406) );
  XOR2_X1 U8123 ( .A(n8197), .B(n8198), .Z(n7403) );
  XOR2_X1 U8124 ( .A(n8199), .B(n8200), .Z(n8198) );
  OR2_X1 U8125 ( .A1(n8201), .A2(n7319), .ZN(n7410) );
  XOR2_X1 U8126 ( .A(n8202), .B(n8203), .Z(n7407) );
  XOR2_X1 U8127 ( .A(n8204), .B(n8205), .Z(n8203) );
  OR2_X1 U8128 ( .A1(n8206), .A2(n7319), .ZN(n7414) );
  XOR2_X1 U8129 ( .A(n8207), .B(n8208), .Z(n7411) );
  XOR2_X1 U8130 ( .A(n8209), .B(n8210), .Z(n8208) );
  OR2_X1 U8131 ( .A1(n8211), .A2(n7319), .ZN(n7418) );
  XOR2_X1 U8132 ( .A(n8212), .B(n8213), .Z(n7415) );
  XOR2_X1 U8133 ( .A(n8214), .B(n8215), .Z(n8213) );
  OR2_X1 U8134 ( .A1(n8216), .A2(n7319), .ZN(n7431) );
  XOR2_X1 U8135 ( .A(n8217), .B(n8218), .Z(n7428) );
  XOR2_X1 U8136 ( .A(n8219), .B(n8220), .Z(n8218) );
  OR2_X1 U8137 ( .A1(n8221), .A2(n7319), .ZN(n7435) );
  XOR2_X1 U8138 ( .A(n8222), .B(n8223), .Z(n7432) );
  XOR2_X1 U8139 ( .A(n8224), .B(n8225), .Z(n8223) );
  OR2_X1 U8140 ( .A1(n8226), .A2(n7319), .ZN(n7439) );
  XOR2_X1 U8141 ( .A(n8227), .B(n8228), .Z(n7436) );
  XOR2_X1 U8142 ( .A(n8229), .B(n8230), .Z(n8228) );
  OR2_X1 U8143 ( .A1(n7785), .A2(n7319), .ZN(n7443) );
  XOR2_X1 U8144 ( .A(n8231), .B(n8232), .Z(n7440) );
  XOR2_X1 U8145 ( .A(n8233), .B(n8234), .Z(n8232) );
  OR2_X1 U8146 ( .A1(n7777), .A2(n7319), .ZN(n7447) );
  XOR2_X1 U8147 ( .A(n8235), .B(n8236), .Z(n7444) );
  XOR2_X1 U8148 ( .A(n8237), .B(n8238), .Z(n8236) );
  OR2_X1 U8149 ( .A1(n7689), .A2(n7319), .ZN(n7451) );
  XOR2_X1 U8150 ( .A(n8239), .B(n8240), .Z(n7448) );
  XOR2_X1 U8151 ( .A(n8241), .B(n8242), .Z(n8240) );
  OR2_X1 U8152 ( .A1(n7656), .A2(n7319), .ZN(n7455) );
  XOR2_X1 U8153 ( .A(n8243), .B(n8244), .Z(n7452) );
  XOR2_X1 U8154 ( .A(n8245), .B(n8246), .Z(n8244) );
  OR2_X1 U8155 ( .A1(n7621), .A2(n7319), .ZN(n7459) );
  INV_X1 U8156 ( .A(b_31_), .ZN(n7319) );
  XOR2_X1 U8157 ( .A(n8247), .B(n8248), .Z(n7456) );
  XOR2_X1 U8158 ( .A(n8249), .B(n8250), .Z(n8248) );
  XOR2_X1 U8159 ( .A(n8005), .B(n8006), .Z(n7465) );
  OR2_X1 U8160 ( .A1(n8251), .A2(n8252), .ZN(n8006) );
  AND2_X1 U8161 ( .A1(n8253), .A2(n8254), .ZN(n8252) );
  AND2_X1 U8162 ( .A1(n8255), .A2(n8256), .ZN(n8251) );
  OR2_X1 U8163 ( .A1(n8253), .A2(n8254), .ZN(n8256) );
  XOR2_X1 U8164 ( .A(n8257), .B(n8258), .Z(n8005) );
  XOR2_X1 U8165 ( .A(n8259), .B(n8260), .Z(n8258) );
  XNOR2_X1 U8166 ( .A(n8255), .B(n8261), .ZN(n7461) );
  XOR2_X1 U8167 ( .A(n8254), .B(n8253), .Z(n8261) );
  OR2_X1 U8168 ( .A1(n7621), .A2(n7315), .ZN(n8253) );
  OR2_X1 U8169 ( .A1(n8262), .A2(n8263), .ZN(n8254) );
  AND2_X1 U8170 ( .A1(n8247), .A2(n8250), .ZN(n8263) );
  AND2_X1 U8171 ( .A1(n8264), .A2(n8249), .ZN(n8262) );
  OR2_X1 U8172 ( .A1(n8265), .A2(n8266), .ZN(n8249) );
  AND2_X1 U8173 ( .A1(n8243), .A2(n8246), .ZN(n8266) );
  AND2_X1 U8174 ( .A1(n8267), .A2(n8245), .ZN(n8265) );
  OR2_X1 U8175 ( .A1(n8268), .A2(n8269), .ZN(n8245) );
  AND2_X1 U8176 ( .A1(n8239), .A2(n8242), .ZN(n8269) );
  AND2_X1 U8177 ( .A1(n8270), .A2(n8241), .ZN(n8268) );
  OR2_X1 U8178 ( .A1(n8271), .A2(n8272), .ZN(n8241) );
  AND2_X1 U8179 ( .A1(n8235), .A2(n8238), .ZN(n8272) );
  AND2_X1 U8180 ( .A1(n8273), .A2(n8237), .ZN(n8271) );
  OR2_X1 U8181 ( .A1(n8274), .A2(n8275), .ZN(n8237) );
  AND2_X1 U8182 ( .A1(n8231), .A2(n8234), .ZN(n8275) );
  AND2_X1 U8183 ( .A1(n8276), .A2(n8233), .ZN(n8274) );
  OR2_X1 U8184 ( .A1(n8277), .A2(n8278), .ZN(n8233) );
  AND2_X1 U8185 ( .A1(n8227), .A2(n8230), .ZN(n8278) );
  AND2_X1 U8186 ( .A1(n8279), .A2(n8229), .ZN(n8277) );
  OR2_X1 U8187 ( .A1(n8280), .A2(n8281), .ZN(n8229) );
  AND2_X1 U8188 ( .A1(n8222), .A2(n8225), .ZN(n8281) );
  AND2_X1 U8189 ( .A1(n8282), .A2(n8224), .ZN(n8280) );
  OR2_X1 U8190 ( .A1(n8283), .A2(n8284), .ZN(n8224) );
  AND2_X1 U8191 ( .A1(n8217), .A2(n8220), .ZN(n8284) );
  AND2_X1 U8192 ( .A1(n8285), .A2(n8219), .ZN(n8283) );
  OR2_X1 U8193 ( .A1(n8286), .A2(n8287), .ZN(n8219) );
  AND2_X1 U8194 ( .A1(n8212), .A2(n8215), .ZN(n8287) );
  AND2_X1 U8195 ( .A1(n8288), .A2(n8214), .ZN(n8286) );
  OR2_X1 U8196 ( .A1(n8289), .A2(n8290), .ZN(n8214) );
  AND2_X1 U8197 ( .A1(n8207), .A2(n8210), .ZN(n8290) );
  AND2_X1 U8198 ( .A1(n8291), .A2(n8209), .ZN(n8289) );
  OR2_X1 U8199 ( .A1(n8292), .A2(n8293), .ZN(n8209) );
  AND2_X1 U8200 ( .A1(n8202), .A2(n8205), .ZN(n8293) );
  AND2_X1 U8201 ( .A1(n8294), .A2(n8204), .ZN(n8292) );
  OR2_X1 U8202 ( .A1(n8295), .A2(n8296), .ZN(n8204) );
  AND2_X1 U8203 ( .A1(n8197), .A2(n8200), .ZN(n8296) );
  AND2_X1 U8204 ( .A1(n8297), .A2(n8199), .ZN(n8295) );
  OR2_X1 U8205 ( .A1(n8298), .A2(n8299), .ZN(n8199) );
  AND2_X1 U8206 ( .A1(n8192), .A2(n8195), .ZN(n8299) );
  AND2_X1 U8207 ( .A1(n8300), .A2(n8194), .ZN(n8298) );
  OR2_X1 U8208 ( .A1(n8301), .A2(n8302), .ZN(n8194) );
  AND2_X1 U8209 ( .A1(n8187), .A2(n8190), .ZN(n8302) );
  AND2_X1 U8210 ( .A1(n8303), .A2(n8189), .ZN(n8301) );
  OR2_X1 U8211 ( .A1(n8304), .A2(n8305), .ZN(n8189) );
  AND2_X1 U8212 ( .A1(n8182), .A2(n8185), .ZN(n8305) );
  AND2_X1 U8213 ( .A1(n8306), .A2(n8184), .ZN(n8304) );
  OR2_X1 U8214 ( .A1(n8307), .A2(n8308), .ZN(n8184) );
  AND2_X1 U8215 ( .A1(n8177), .A2(n8180), .ZN(n8308) );
  AND2_X1 U8216 ( .A1(n8309), .A2(n8179), .ZN(n8307) );
  OR2_X1 U8217 ( .A1(n8310), .A2(n8311), .ZN(n8179) );
  AND2_X1 U8218 ( .A1(n8172), .A2(n8175), .ZN(n8311) );
  AND2_X1 U8219 ( .A1(n8312), .A2(n8174), .ZN(n8310) );
  OR2_X1 U8220 ( .A1(n8313), .A2(n8314), .ZN(n8174) );
  AND2_X1 U8221 ( .A1(n8167), .A2(n8170), .ZN(n8314) );
  AND2_X1 U8222 ( .A1(n8315), .A2(n8169), .ZN(n8313) );
  OR2_X1 U8223 ( .A1(n8316), .A2(n8317), .ZN(n8169) );
  AND2_X1 U8224 ( .A1(n8162), .A2(n8165), .ZN(n8317) );
  AND2_X1 U8225 ( .A1(n8318), .A2(n8164), .ZN(n8316) );
  OR2_X1 U8226 ( .A1(n8319), .A2(n8320), .ZN(n8164) );
  AND2_X1 U8227 ( .A1(n8157), .A2(n8160), .ZN(n8320) );
  AND2_X1 U8228 ( .A1(n8321), .A2(n8159), .ZN(n8319) );
  OR2_X1 U8229 ( .A1(n8322), .A2(n8323), .ZN(n8159) );
  AND2_X1 U8230 ( .A1(n8152), .A2(n8155), .ZN(n8323) );
  AND2_X1 U8231 ( .A1(n8324), .A2(n8154), .ZN(n8322) );
  OR2_X1 U8232 ( .A1(n8325), .A2(n8326), .ZN(n8154) );
  AND2_X1 U8233 ( .A1(n8147), .A2(n8150), .ZN(n8326) );
  AND2_X1 U8234 ( .A1(n8327), .A2(n8149), .ZN(n8325) );
  OR2_X1 U8235 ( .A1(n8328), .A2(n8329), .ZN(n8149) );
  AND2_X1 U8236 ( .A1(n8142), .A2(n8145), .ZN(n8329) );
  AND2_X1 U8237 ( .A1(n8330), .A2(n8144), .ZN(n8328) );
  OR2_X1 U8238 ( .A1(n8331), .A2(n8332), .ZN(n8144) );
  AND2_X1 U8239 ( .A1(n8137), .A2(n8140), .ZN(n8332) );
  AND2_X1 U8240 ( .A1(n8333), .A2(n8139), .ZN(n8331) );
  OR2_X1 U8241 ( .A1(n8334), .A2(n8335), .ZN(n8139) );
  AND2_X1 U8242 ( .A1(n8132), .A2(n8135), .ZN(n8335) );
  AND2_X1 U8243 ( .A1(n8336), .A2(n8134), .ZN(n8334) );
  OR2_X1 U8244 ( .A1(n8337), .A2(n8338), .ZN(n8134) );
  AND2_X1 U8245 ( .A1(n8127), .A2(n8130), .ZN(n8338) );
  AND2_X1 U8246 ( .A1(n8339), .A2(n8129), .ZN(n8337) );
  OR2_X1 U8247 ( .A1(n8340), .A2(n8341), .ZN(n8129) );
  AND2_X1 U8248 ( .A1(n8122), .A2(n8125), .ZN(n8341) );
  AND2_X1 U8249 ( .A1(n8342), .A2(n8124), .ZN(n8340) );
  OR2_X1 U8250 ( .A1(n8343), .A2(n8344), .ZN(n8124) );
  AND2_X1 U8251 ( .A1(n8117), .A2(n8120), .ZN(n8344) );
  AND2_X1 U8252 ( .A1(n8345), .A2(n8119), .ZN(n8343) );
  OR2_X1 U8253 ( .A1(n8346), .A2(n8347), .ZN(n8119) );
  AND2_X1 U8254 ( .A1(n8112), .A2(n8115), .ZN(n8347) );
  AND2_X1 U8255 ( .A1(n8114), .A2(n8348), .ZN(n8346) );
  OR2_X1 U8256 ( .A1(n8115), .A2(n8112), .ZN(n8348) );
  OR2_X1 U8257 ( .A1(n8102), .A2(n7315), .ZN(n8112) );
  OR3_X1 U8258 ( .A1(n8349), .A2(n7315), .A3(n8110), .ZN(n8115) );
  INV_X1 U8259 ( .A(n8350), .ZN(n8114) );
  OR2_X1 U8260 ( .A1(n8351), .A2(n8352), .ZN(n8350) );
  AND2_X1 U8261 ( .A1(b_29_), .A2(n8353), .ZN(n8352) );
  OR2_X1 U8262 ( .A1(n8354), .A2(n7314), .ZN(n8353) );
  AND2_X1 U8263 ( .A1(a_30_), .A2(n8355), .ZN(n8354) );
  AND2_X1 U8264 ( .A1(b_28_), .A2(n8356), .ZN(n8351) );
  OR2_X1 U8265 ( .A1(n8357), .A2(n7318), .ZN(n8356) );
  AND2_X1 U8266 ( .A1(a_31_), .A2(n8110), .ZN(n8357) );
  OR2_X1 U8267 ( .A1(n8120), .A2(n8117), .ZN(n8345) );
  XOR2_X1 U8268 ( .A(n8358), .B(n8359), .Z(n8117) );
  XNOR2_X1 U8269 ( .A(n8360), .B(n8361), .ZN(n8358) );
  OR2_X1 U8270 ( .A1(n8111), .A2(n7315), .ZN(n8120) );
  OR2_X1 U8271 ( .A1(n8125), .A2(n8122), .ZN(n8342) );
  XOR2_X1 U8272 ( .A(n8362), .B(n8363), .Z(n8122) );
  XOR2_X1 U8273 ( .A(n8364), .B(n8365), .Z(n8363) );
  OR2_X1 U8274 ( .A1(n8116), .A2(n7315), .ZN(n8125) );
  OR2_X1 U8275 ( .A1(n8130), .A2(n8127), .ZN(n8339) );
  XOR2_X1 U8276 ( .A(n8366), .B(n8367), .Z(n8127) );
  XOR2_X1 U8277 ( .A(n8368), .B(n8369), .Z(n8367) );
  OR2_X1 U8278 ( .A1(n8121), .A2(n7315), .ZN(n8130) );
  OR2_X1 U8279 ( .A1(n8135), .A2(n8132), .ZN(n8336) );
  XOR2_X1 U8280 ( .A(n8370), .B(n8371), .Z(n8132) );
  XOR2_X1 U8281 ( .A(n8372), .B(n8373), .Z(n8371) );
  OR2_X1 U8282 ( .A1(n8126), .A2(n7315), .ZN(n8135) );
  OR2_X1 U8283 ( .A1(n8140), .A2(n8137), .ZN(n8333) );
  XOR2_X1 U8284 ( .A(n8374), .B(n8375), .Z(n8137) );
  XOR2_X1 U8285 ( .A(n8376), .B(n8377), .Z(n8375) );
  OR2_X1 U8286 ( .A1(n8131), .A2(n7315), .ZN(n8140) );
  OR2_X1 U8287 ( .A1(n8145), .A2(n8142), .ZN(n8330) );
  XOR2_X1 U8288 ( .A(n8378), .B(n8379), .Z(n8142) );
  XOR2_X1 U8289 ( .A(n8380), .B(n8381), .Z(n8379) );
  OR2_X1 U8290 ( .A1(n8136), .A2(n7315), .ZN(n8145) );
  OR2_X1 U8291 ( .A1(n8150), .A2(n8147), .ZN(n8327) );
  XOR2_X1 U8292 ( .A(n8382), .B(n8383), .Z(n8147) );
  XOR2_X1 U8293 ( .A(n8384), .B(n8385), .Z(n8383) );
  OR2_X1 U8294 ( .A1(n8141), .A2(n7315), .ZN(n8150) );
  OR2_X1 U8295 ( .A1(n8155), .A2(n8152), .ZN(n8324) );
  XOR2_X1 U8296 ( .A(n8386), .B(n8387), .Z(n8152) );
  XOR2_X1 U8297 ( .A(n8388), .B(n8389), .Z(n8387) );
  OR2_X1 U8298 ( .A1(n8146), .A2(n7315), .ZN(n8155) );
  OR2_X1 U8299 ( .A1(n8160), .A2(n8157), .ZN(n8321) );
  XOR2_X1 U8300 ( .A(n8390), .B(n8391), .Z(n8157) );
  XOR2_X1 U8301 ( .A(n8392), .B(n8393), .Z(n8391) );
  OR2_X1 U8302 ( .A1(n8151), .A2(n7315), .ZN(n8160) );
  OR2_X1 U8303 ( .A1(n8165), .A2(n8162), .ZN(n8318) );
  XOR2_X1 U8304 ( .A(n8394), .B(n8395), .Z(n8162) );
  XOR2_X1 U8305 ( .A(n8396), .B(n8397), .Z(n8395) );
  OR2_X1 U8306 ( .A1(n8156), .A2(n7315), .ZN(n8165) );
  OR2_X1 U8307 ( .A1(n8170), .A2(n8167), .ZN(n8315) );
  XOR2_X1 U8308 ( .A(n8398), .B(n8399), .Z(n8167) );
  XOR2_X1 U8309 ( .A(n8400), .B(n8401), .Z(n8399) );
  OR2_X1 U8310 ( .A1(n8161), .A2(n7315), .ZN(n8170) );
  OR2_X1 U8311 ( .A1(n8175), .A2(n8172), .ZN(n8312) );
  XOR2_X1 U8312 ( .A(n8402), .B(n8403), .Z(n8172) );
  XOR2_X1 U8313 ( .A(n8404), .B(n8405), .Z(n8403) );
  OR2_X1 U8314 ( .A1(n8166), .A2(n7315), .ZN(n8175) );
  OR2_X1 U8315 ( .A1(n8180), .A2(n8177), .ZN(n8309) );
  XOR2_X1 U8316 ( .A(n8406), .B(n8407), .Z(n8177) );
  XOR2_X1 U8317 ( .A(n8408), .B(n8409), .Z(n8407) );
  OR2_X1 U8318 ( .A1(n8171), .A2(n7315), .ZN(n8180) );
  OR2_X1 U8319 ( .A1(n8185), .A2(n8182), .ZN(n8306) );
  XOR2_X1 U8320 ( .A(n8410), .B(n8411), .Z(n8182) );
  XOR2_X1 U8321 ( .A(n8412), .B(n8413), .Z(n8411) );
  OR2_X1 U8322 ( .A1(n8176), .A2(n7315), .ZN(n8185) );
  OR2_X1 U8323 ( .A1(n8190), .A2(n8187), .ZN(n8303) );
  XOR2_X1 U8324 ( .A(n8414), .B(n8415), .Z(n8187) );
  XOR2_X1 U8325 ( .A(n8416), .B(n8417), .Z(n8415) );
  OR2_X1 U8326 ( .A1(n8181), .A2(n7315), .ZN(n8190) );
  OR2_X1 U8327 ( .A1(n8195), .A2(n8192), .ZN(n8300) );
  XOR2_X1 U8328 ( .A(n8418), .B(n8419), .Z(n8192) );
  XOR2_X1 U8329 ( .A(n8420), .B(n8421), .Z(n8419) );
  OR2_X1 U8330 ( .A1(n8186), .A2(n7315), .ZN(n8195) );
  OR2_X1 U8331 ( .A1(n8200), .A2(n8197), .ZN(n8297) );
  XOR2_X1 U8332 ( .A(n8422), .B(n8423), .Z(n8197) );
  XOR2_X1 U8333 ( .A(n8424), .B(n8425), .Z(n8423) );
  OR2_X1 U8334 ( .A1(n8191), .A2(n7315), .ZN(n8200) );
  OR2_X1 U8335 ( .A1(n8205), .A2(n8202), .ZN(n8294) );
  XOR2_X1 U8336 ( .A(n8426), .B(n8427), .Z(n8202) );
  XOR2_X1 U8337 ( .A(n8428), .B(n8429), .Z(n8427) );
  OR2_X1 U8338 ( .A1(n8196), .A2(n7315), .ZN(n8205) );
  OR2_X1 U8339 ( .A1(n8210), .A2(n8207), .ZN(n8291) );
  XOR2_X1 U8340 ( .A(n8430), .B(n8431), .Z(n8207) );
  XOR2_X1 U8341 ( .A(n8432), .B(n8433), .Z(n8431) );
  OR2_X1 U8342 ( .A1(n8201), .A2(n7315), .ZN(n8210) );
  OR2_X1 U8343 ( .A1(n8215), .A2(n8212), .ZN(n8288) );
  XOR2_X1 U8344 ( .A(n8434), .B(n8435), .Z(n8212) );
  XOR2_X1 U8345 ( .A(n8436), .B(n8437), .Z(n8435) );
  OR2_X1 U8346 ( .A1(n8206), .A2(n7315), .ZN(n8215) );
  OR2_X1 U8347 ( .A1(n8220), .A2(n8217), .ZN(n8285) );
  XOR2_X1 U8348 ( .A(n8438), .B(n8439), .Z(n8217) );
  XOR2_X1 U8349 ( .A(n8440), .B(n8441), .Z(n8439) );
  OR2_X1 U8350 ( .A1(n8211), .A2(n7315), .ZN(n8220) );
  OR2_X1 U8351 ( .A1(n8225), .A2(n8222), .ZN(n8282) );
  XOR2_X1 U8352 ( .A(n8442), .B(n8443), .Z(n8222) );
  XOR2_X1 U8353 ( .A(n8444), .B(n8445), .Z(n8443) );
  OR2_X1 U8354 ( .A1(n8216), .A2(n7315), .ZN(n8225) );
  OR2_X1 U8355 ( .A1(n8230), .A2(n8227), .ZN(n8279) );
  XOR2_X1 U8356 ( .A(n8446), .B(n8447), .Z(n8227) );
  XOR2_X1 U8357 ( .A(n8448), .B(n8449), .Z(n8447) );
  OR2_X1 U8358 ( .A1(n8221), .A2(n7315), .ZN(n8230) );
  OR2_X1 U8359 ( .A1(n8234), .A2(n8231), .ZN(n8276) );
  XOR2_X1 U8360 ( .A(n8450), .B(n8451), .Z(n8231) );
  XOR2_X1 U8361 ( .A(n8452), .B(n8453), .Z(n8451) );
  OR2_X1 U8362 ( .A1(n8226), .A2(n7315), .ZN(n8234) );
  OR2_X1 U8363 ( .A1(n8238), .A2(n8235), .ZN(n8273) );
  XOR2_X1 U8364 ( .A(n8454), .B(n8455), .Z(n8235) );
  XOR2_X1 U8365 ( .A(n8456), .B(n8457), .Z(n8455) );
  OR2_X1 U8366 ( .A1(n7785), .A2(n7315), .ZN(n8238) );
  OR2_X1 U8367 ( .A1(n8242), .A2(n8239), .ZN(n8270) );
  XOR2_X1 U8368 ( .A(n8458), .B(n8459), .Z(n8239) );
  XOR2_X1 U8369 ( .A(n8460), .B(n8461), .Z(n8459) );
  OR2_X1 U8370 ( .A1(n7777), .A2(n7315), .ZN(n8242) );
  OR2_X1 U8371 ( .A1(n8246), .A2(n8243), .ZN(n8267) );
  XOR2_X1 U8372 ( .A(n8462), .B(n8463), .Z(n8243) );
  XOR2_X1 U8373 ( .A(n8464), .B(n8465), .Z(n8463) );
  OR2_X1 U8374 ( .A1(n7689), .A2(n7315), .ZN(n8246) );
  OR2_X1 U8375 ( .A1(n8250), .A2(n8247), .ZN(n8264) );
  XNOR2_X1 U8376 ( .A(n8466), .B(n8467), .ZN(n8247) );
  XNOR2_X1 U8377 ( .A(n8468), .B(n8469), .ZN(n8466) );
  OR2_X1 U8378 ( .A1(n7656), .A2(n7315), .ZN(n8250) );
  XOR2_X1 U8379 ( .A(n8470), .B(n8471), .Z(n8255) );
  XOR2_X1 U8380 ( .A(n8472), .B(n8473), .Z(n8471) );
  OR2_X1 U8381 ( .A1(n8474), .A2(n8000), .ZN(n7475) );
  XNOR2_X1 U8382 ( .A(n7995), .B(n8475), .ZN(n8000) );
  AND2_X1 U8383 ( .A1(n8001), .A2(n7999), .ZN(n8474) );
  XNOR2_X1 U8384 ( .A(n8476), .B(n8477), .ZN(n7999) );
  XOR2_X1 U8385 ( .A(n8478), .B(n8479), .Z(n8477) );
  INV_X1 U8386 ( .A(n8009), .ZN(n8001) );
  OR2_X1 U8387 ( .A1(n8480), .A2(n8481), .ZN(n8009) );
  AND2_X1 U8388 ( .A1(n8260), .A2(n8259), .ZN(n8481) );
  AND2_X1 U8389 ( .A1(n8257), .A2(n8482), .ZN(n8480) );
  OR2_X1 U8390 ( .A1(n8259), .A2(n8260), .ZN(n8482) );
  OR2_X1 U8391 ( .A1(n7621), .A2(n8110), .ZN(n8260) );
  OR2_X1 U8392 ( .A1(n8483), .A2(n8484), .ZN(n8259) );
  AND2_X1 U8393 ( .A1(n8473), .A2(n8472), .ZN(n8484) );
  AND2_X1 U8394 ( .A1(n8470), .A2(n8485), .ZN(n8483) );
  OR2_X1 U8395 ( .A1(n8472), .A2(n8473), .ZN(n8485) );
  OR2_X1 U8396 ( .A1(n7656), .A2(n8110), .ZN(n8473) );
  OR2_X1 U8397 ( .A1(n8486), .A2(n8487), .ZN(n8472) );
  AND2_X1 U8398 ( .A1(n8469), .A2(n8468), .ZN(n8487) );
  AND2_X1 U8399 ( .A1(n8467), .A2(n8488), .ZN(n8486) );
  OR2_X1 U8400 ( .A1(n8468), .A2(n8469), .ZN(n8488) );
  OR2_X1 U8401 ( .A1(n8489), .A2(n8490), .ZN(n8469) );
  AND2_X1 U8402 ( .A1(n8465), .A2(n8464), .ZN(n8490) );
  AND2_X1 U8403 ( .A1(n8462), .A2(n8491), .ZN(n8489) );
  OR2_X1 U8404 ( .A1(n8464), .A2(n8465), .ZN(n8491) );
  OR2_X1 U8405 ( .A1(n7777), .A2(n8110), .ZN(n8465) );
  OR2_X1 U8406 ( .A1(n8492), .A2(n8493), .ZN(n8464) );
  AND2_X1 U8407 ( .A1(n8461), .A2(n8460), .ZN(n8493) );
  AND2_X1 U8408 ( .A1(n8458), .A2(n8494), .ZN(n8492) );
  OR2_X1 U8409 ( .A1(n8460), .A2(n8461), .ZN(n8494) );
  OR2_X1 U8410 ( .A1(n7785), .A2(n8110), .ZN(n8461) );
  OR2_X1 U8411 ( .A1(n8495), .A2(n8496), .ZN(n8460) );
  AND2_X1 U8412 ( .A1(n8457), .A2(n8456), .ZN(n8496) );
  AND2_X1 U8413 ( .A1(n8454), .A2(n8497), .ZN(n8495) );
  OR2_X1 U8414 ( .A1(n8456), .A2(n8457), .ZN(n8497) );
  OR2_X1 U8415 ( .A1(n8226), .A2(n8110), .ZN(n8457) );
  OR2_X1 U8416 ( .A1(n8498), .A2(n8499), .ZN(n8456) );
  AND2_X1 U8417 ( .A1(n8453), .A2(n8452), .ZN(n8499) );
  AND2_X1 U8418 ( .A1(n8450), .A2(n8500), .ZN(n8498) );
  OR2_X1 U8419 ( .A1(n8452), .A2(n8453), .ZN(n8500) );
  OR2_X1 U8420 ( .A1(n8221), .A2(n8110), .ZN(n8453) );
  OR2_X1 U8421 ( .A1(n8501), .A2(n8502), .ZN(n8452) );
  AND2_X1 U8422 ( .A1(n8449), .A2(n8448), .ZN(n8502) );
  AND2_X1 U8423 ( .A1(n8446), .A2(n8503), .ZN(n8501) );
  OR2_X1 U8424 ( .A1(n8448), .A2(n8449), .ZN(n8503) );
  OR2_X1 U8425 ( .A1(n8216), .A2(n8110), .ZN(n8449) );
  OR2_X1 U8426 ( .A1(n8504), .A2(n8505), .ZN(n8448) );
  AND2_X1 U8427 ( .A1(n8445), .A2(n8444), .ZN(n8505) );
  AND2_X1 U8428 ( .A1(n8442), .A2(n8506), .ZN(n8504) );
  OR2_X1 U8429 ( .A1(n8444), .A2(n8445), .ZN(n8506) );
  OR2_X1 U8430 ( .A1(n8211), .A2(n8110), .ZN(n8445) );
  OR2_X1 U8431 ( .A1(n8507), .A2(n8508), .ZN(n8444) );
  AND2_X1 U8432 ( .A1(n8441), .A2(n8440), .ZN(n8508) );
  AND2_X1 U8433 ( .A1(n8438), .A2(n8509), .ZN(n8507) );
  OR2_X1 U8434 ( .A1(n8440), .A2(n8441), .ZN(n8509) );
  OR2_X1 U8435 ( .A1(n8206), .A2(n8110), .ZN(n8441) );
  OR2_X1 U8436 ( .A1(n8510), .A2(n8511), .ZN(n8440) );
  AND2_X1 U8437 ( .A1(n8437), .A2(n8436), .ZN(n8511) );
  AND2_X1 U8438 ( .A1(n8434), .A2(n8512), .ZN(n8510) );
  OR2_X1 U8439 ( .A1(n8436), .A2(n8437), .ZN(n8512) );
  OR2_X1 U8440 ( .A1(n8201), .A2(n8110), .ZN(n8437) );
  OR2_X1 U8441 ( .A1(n8513), .A2(n8514), .ZN(n8436) );
  AND2_X1 U8442 ( .A1(n8433), .A2(n8432), .ZN(n8514) );
  AND2_X1 U8443 ( .A1(n8430), .A2(n8515), .ZN(n8513) );
  OR2_X1 U8444 ( .A1(n8432), .A2(n8433), .ZN(n8515) );
  OR2_X1 U8445 ( .A1(n8196), .A2(n8110), .ZN(n8433) );
  OR2_X1 U8446 ( .A1(n8516), .A2(n8517), .ZN(n8432) );
  AND2_X1 U8447 ( .A1(n8429), .A2(n8428), .ZN(n8517) );
  AND2_X1 U8448 ( .A1(n8426), .A2(n8518), .ZN(n8516) );
  OR2_X1 U8449 ( .A1(n8428), .A2(n8429), .ZN(n8518) );
  OR2_X1 U8450 ( .A1(n8191), .A2(n8110), .ZN(n8429) );
  OR2_X1 U8451 ( .A1(n8519), .A2(n8520), .ZN(n8428) );
  AND2_X1 U8452 ( .A1(n8425), .A2(n8424), .ZN(n8520) );
  AND2_X1 U8453 ( .A1(n8422), .A2(n8521), .ZN(n8519) );
  OR2_X1 U8454 ( .A1(n8424), .A2(n8425), .ZN(n8521) );
  OR2_X1 U8455 ( .A1(n8186), .A2(n8110), .ZN(n8425) );
  OR2_X1 U8456 ( .A1(n8522), .A2(n8523), .ZN(n8424) );
  AND2_X1 U8457 ( .A1(n8421), .A2(n8420), .ZN(n8523) );
  AND2_X1 U8458 ( .A1(n8418), .A2(n8524), .ZN(n8522) );
  OR2_X1 U8459 ( .A1(n8420), .A2(n8421), .ZN(n8524) );
  OR2_X1 U8460 ( .A1(n8181), .A2(n8110), .ZN(n8421) );
  OR2_X1 U8461 ( .A1(n8525), .A2(n8526), .ZN(n8420) );
  AND2_X1 U8462 ( .A1(n8417), .A2(n8416), .ZN(n8526) );
  AND2_X1 U8463 ( .A1(n8414), .A2(n8527), .ZN(n8525) );
  OR2_X1 U8464 ( .A1(n8416), .A2(n8417), .ZN(n8527) );
  OR2_X1 U8465 ( .A1(n8176), .A2(n8110), .ZN(n8417) );
  OR2_X1 U8466 ( .A1(n8528), .A2(n8529), .ZN(n8416) );
  AND2_X1 U8467 ( .A1(n8413), .A2(n8412), .ZN(n8529) );
  AND2_X1 U8468 ( .A1(n8410), .A2(n8530), .ZN(n8528) );
  OR2_X1 U8469 ( .A1(n8412), .A2(n8413), .ZN(n8530) );
  OR2_X1 U8470 ( .A1(n8171), .A2(n8110), .ZN(n8413) );
  OR2_X1 U8471 ( .A1(n8531), .A2(n8532), .ZN(n8412) );
  AND2_X1 U8472 ( .A1(n8409), .A2(n8408), .ZN(n8532) );
  AND2_X1 U8473 ( .A1(n8406), .A2(n8533), .ZN(n8531) );
  OR2_X1 U8474 ( .A1(n8408), .A2(n8409), .ZN(n8533) );
  OR2_X1 U8475 ( .A1(n8166), .A2(n8110), .ZN(n8409) );
  OR2_X1 U8476 ( .A1(n8534), .A2(n8535), .ZN(n8408) );
  AND2_X1 U8477 ( .A1(n8405), .A2(n8404), .ZN(n8535) );
  AND2_X1 U8478 ( .A1(n8402), .A2(n8536), .ZN(n8534) );
  OR2_X1 U8479 ( .A1(n8404), .A2(n8405), .ZN(n8536) );
  OR2_X1 U8480 ( .A1(n8161), .A2(n8110), .ZN(n8405) );
  OR2_X1 U8481 ( .A1(n8537), .A2(n8538), .ZN(n8404) );
  AND2_X1 U8482 ( .A1(n8401), .A2(n8400), .ZN(n8538) );
  AND2_X1 U8483 ( .A1(n8398), .A2(n8539), .ZN(n8537) );
  OR2_X1 U8484 ( .A1(n8400), .A2(n8401), .ZN(n8539) );
  OR2_X1 U8485 ( .A1(n8156), .A2(n8110), .ZN(n8401) );
  OR2_X1 U8486 ( .A1(n8540), .A2(n8541), .ZN(n8400) );
  AND2_X1 U8487 ( .A1(n8397), .A2(n8396), .ZN(n8541) );
  AND2_X1 U8488 ( .A1(n8394), .A2(n8542), .ZN(n8540) );
  OR2_X1 U8489 ( .A1(n8396), .A2(n8397), .ZN(n8542) );
  OR2_X1 U8490 ( .A1(n8151), .A2(n8110), .ZN(n8397) );
  OR2_X1 U8491 ( .A1(n8543), .A2(n8544), .ZN(n8396) );
  AND2_X1 U8492 ( .A1(n8393), .A2(n8392), .ZN(n8544) );
  AND2_X1 U8493 ( .A1(n8390), .A2(n8545), .ZN(n8543) );
  OR2_X1 U8494 ( .A1(n8392), .A2(n8393), .ZN(n8545) );
  OR2_X1 U8495 ( .A1(n8146), .A2(n8110), .ZN(n8393) );
  OR2_X1 U8496 ( .A1(n8546), .A2(n8547), .ZN(n8392) );
  AND2_X1 U8497 ( .A1(n8389), .A2(n8388), .ZN(n8547) );
  AND2_X1 U8498 ( .A1(n8386), .A2(n8548), .ZN(n8546) );
  OR2_X1 U8499 ( .A1(n8388), .A2(n8389), .ZN(n8548) );
  OR2_X1 U8500 ( .A1(n8141), .A2(n8110), .ZN(n8389) );
  OR2_X1 U8501 ( .A1(n8549), .A2(n8550), .ZN(n8388) );
  AND2_X1 U8502 ( .A1(n8385), .A2(n8384), .ZN(n8550) );
  AND2_X1 U8503 ( .A1(n8382), .A2(n8551), .ZN(n8549) );
  OR2_X1 U8504 ( .A1(n8384), .A2(n8385), .ZN(n8551) );
  OR2_X1 U8505 ( .A1(n8136), .A2(n8110), .ZN(n8385) );
  OR2_X1 U8506 ( .A1(n8552), .A2(n8553), .ZN(n8384) );
  AND2_X1 U8507 ( .A1(n8381), .A2(n8380), .ZN(n8553) );
  AND2_X1 U8508 ( .A1(n8378), .A2(n8554), .ZN(n8552) );
  OR2_X1 U8509 ( .A1(n8380), .A2(n8381), .ZN(n8554) );
  OR2_X1 U8510 ( .A1(n8131), .A2(n8110), .ZN(n8381) );
  OR2_X1 U8511 ( .A1(n8555), .A2(n8556), .ZN(n8380) );
  AND2_X1 U8512 ( .A1(n8377), .A2(n8376), .ZN(n8556) );
  AND2_X1 U8513 ( .A1(n8374), .A2(n8557), .ZN(n8555) );
  OR2_X1 U8514 ( .A1(n8376), .A2(n8377), .ZN(n8557) );
  OR2_X1 U8515 ( .A1(n8126), .A2(n8110), .ZN(n8377) );
  OR2_X1 U8516 ( .A1(n8558), .A2(n8559), .ZN(n8376) );
  AND2_X1 U8517 ( .A1(n8373), .A2(n8372), .ZN(n8559) );
  AND2_X1 U8518 ( .A1(n8370), .A2(n8560), .ZN(n8558) );
  OR2_X1 U8519 ( .A1(n8372), .A2(n8373), .ZN(n8560) );
  OR2_X1 U8520 ( .A1(n8121), .A2(n8110), .ZN(n8373) );
  OR2_X1 U8521 ( .A1(n8561), .A2(n8562), .ZN(n8372) );
  AND2_X1 U8522 ( .A1(n8369), .A2(n8368), .ZN(n8562) );
  AND2_X1 U8523 ( .A1(n8366), .A2(n8563), .ZN(n8561) );
  OR2_X1 U8524 ( .A1(n8368), .A2(n8369), .ZN(n8563) );
  OR2_X1 U8525 ( .A1(n8116), .A2(n8110), .ZN(n8369) );
  OR2_X1 U8526 ( .A1(n8564), .A2(n8565), .ZN(n8368) );
  AND2_X1 U8527 ( .A1(n8365), .A2(n8364), .ZN(n8565) );
  AND2_X1 U8528 ( .A1(n8362), .A2(n8566), .ZN(n8564) );
  OR2_X1 U8529 ( .A1(n8364), .A2(n8365), .ZN(n8566) );
  OR2_X1 U8530 ( .A1(n8111), .A2(n8110), .ZN(n8365) );
  OR2_X1 U8531 ( .A1(n8567), .A2(n8568), .ZN(n8364) );
  AND2_X1 U8532 ( .A1(n8569), .A2(n8359), .ZN(n8568) );
  AND2_X1 U8533 ( .A1(n8570), .A2(n8360), .ZN(n8567) );
  OR2_X1 U8534 ( .A1(n8569), .A2(n8359), .ZN(n8570) );
  OR3_X1 U8535 ( .A1(n8349), .A2(n8110), .A3(n8355), .ZN(n8359) );
  INV_X1 U8536 ( .A(n8361), .ZN(n8569) );
  OR2_X1 U8537 ( .A1(n8571), .A2(n8572), .ZN(n8361) );
  AND2_X1 U8538 ( .A1(b_28_), .A2(n8573), .ZN(n8572) );
  OR2_X1 U8539 ( .A1(n8574), .A2(n7314), .ZN(n8573) );
  AND2_X1 U8540 ( .A1(a_30_), .A2(n8575), .ZN(n8574) );
  AND2_X1 U8541 ( .A1(b_27_), .A2(n8576), .ZN(n8571) );
  OR2_X1 U8542 ( .A1(n8577), .A2(n7318), .ZN(n8576) );
  AND2_X1 U8543 ( .A1(a_31_), .A2(n8355), .ZN(n8577) );
  XNOR2_X1 U8544 ( .A(n8578), .B(n8579), .ZN(n8362) );
  XNOR2_X1 U8545 ( .A(n8580), .B(n8581), .ZN(n8579) );
  XNOR2_X1 U8546 ( .A(n8582), .B(n8583), .ZN(n8366) );
  XNOR2_X1 U8547 ( .A(n8584), .B(n8585), .ZN(n8582) );
  XOR2_X1 U8548 ( .A(n8586), .B(n8587), .Z(n8370) );
  XOR2_X1 U8549 ( .A(n8588), .B(n8589), .Z(n8587) );
  XOR2_X1 U8550 ( .A(n8590), .B(n8591), .Z(n8374) );
  XOR2_X1 U8551 ( .A(n8592), .B(n8593), .Z(n8591) );
  XOR2_X1 U8552 ( .A(n8594), .B(n8595), .Z(n8378) );
  XOR2_X1 U8553 ( .A(n8596), .B(n8597), .Z(n8595) );
  XOR2_X1 U8554 ( .A(n8598), .B(n8599), .Z(n8382) );
  XOR2_X1 U8555 ( .A(n8600), .B(n8601), .Z(n8599) );
  XOR2_X1 U8556 ( .A(n8602), .B(n8603), .Z(n8386) );
  XOR2_X1 U8557 ( .A(n8604), .B(n8605), .Z(n8603) );
  XOR2_X1 U8558 ( .A(n8606), .B(n8607), .Z(n8390) );
  XOR2_X1 U8559 ( .A(n8608), .B(n8609), .Z(n8607) );
  XOR2_X1 U8560 ( .A(n8610), .B(n8611), .Z(n8394) );
  XOR2_X1 U8561 ( .A(n8612), .B(n8613), .Z(n8611) );
  XOR2_X1 U8562 ( .A(n8614), .B(n8615), .Z(n8398) );
  XOR2_X1 U8563 ( .A(n8616), .B(n8617), .Z(n8615) );
  XOR2_X1 U8564 ( .A(n8618), .B(n8619), .Z(n8402) );
  XOR2_X1 U8565 ( .A(n8620), .B(n8621), .Z(n8619) );
  XOR2_X1 U8566 ( .A(n8622), .B(n8623), .Z(n8406) );
  XOR2_X1 U8567 ( .A(n8624), .B(n8625), .Z(n8623) );
  XOR2_X1 U8568 ( .A(n8626), .B(n8627), .Z(n8410) );
  XOR2_X1 U8569 ( .A(n8628), .B(n8629), .Z(n8627) );
  XOR2_X1 U8570 ( .A(n8630), .B(n8631), .Z(n8414) );
  XOR2_X1 U8571 ( .A(n8632), .B(n8633), .Z(n8631) );
  XOR2_X1 U8572 ( .A(n8634), .B(n8635), .Z(n8418) );
  XOR2_X1 U8573 ( .A(n8636), .B(n8637), .Z(n8635) );
  XOR2_X1 U8574 ( .A(n8638), .B(n8639), .Z(n8422) );
  XOR2_X1 U8575 ( .A(n8640), .B(n8641), .Z(n8639) );
  XOR2_X1 U8576 ( .A(n8642), .B(n8643), .Z(n8426) );
  XOR2_X1 U8577 ( .A(n8644), .B(n8645), .Z(n8643) );
  XOR2_X1 U8578 ( .A(n8646), .B(n8647), .Z(n8430) );
  XOR2_X1 U8579 ( .A(n8648), .B(n8649), .Z(n8647) );
  XOR2_X1 U8580 ( .A(n8650), .B(n8651), .Z(n8434) );
  XOR2_X1 U8581 ( .A(n8652), .B(n8653), .Z(n8651) );
  XOR2_X1 U8582 ( .A(n8654), .B(n8655), .Z(n8438) );
  XOR2_X1 U8583 ( .A(n8656), .B(n8657), .Z(n8655) );
  XOR2_X1 U8584 ( .A(n8658), .B(n8659), .Z(n8442) );
  XOR2_X1 U8585 ( .A(n8660), .B(n8661), .Z(n8659) );
  XOR2_X1 U8586 ( .A(n8662), .B(n8663), .Z(n8446) );
  XOR2_X1 U8587 ( .A(n8664), .B(n8665), .Z(n8663) );
  XOR2_X1 U8588 ( .A(n8666), .B(n8667), .Z(n8450) );
  XOR2_X1 U8589 ( .A(n8668), .B(n8669), .Z(n8667) );
  XOR2_X1 U8590 ( .A(n8670), .B(n8671), .Z(n8454) );
  XOR2_X1 U8591 ( .A(n8672), .B(n8673), .Z(n8671) );
  XOR2_X1 U8592 ( .A(n8674), .B(n8675), .Z(n8458) );
  XOR2_X1 U8593 ( .A(n8676), .B(n8677), .Z(n8675) );
  XOR2_X1 U8594 ( .A(n8678), .B(n8679), .Z(n8462) );
  XOR2_X1 U8595 ( .A(n8680), .B(n8681), .Z(n8679) );
  OR2_X1 U8596 ( .A1(n7689), .A2(n8110), .ZN(n8468) );
  XOR2_X1 U8597 ( .A(n8682), .B(n8683), .Z(n8467) );
  XOR2_X1 U8598 ( .A(n8684), .B(n8685), .Z(n8683) );
  XNOR2_X1 U8599 ( .A(n8686), .B(n8687), .ZN(n8470) );
  XNOR2_X1 U8600 ( .A(n8688), .B(n8689), .ZN(n8686) );
  XOR2_X1 U8601 ( .A(n8690), .B(n8691), .Z(n8257) );
  XOR2_X1 U8602 ( .A(n8692), .B(n8693), .Z(n8691) );
  OR2_X1 U8603 ( .A1(n8694), .A2(n7997), .ZN(n7480) );
  INV_X1 U8604 ( .A(n8695), .ZN(n7997) );
  OR2_X1 U8605 ( .A1(n8696), .A2(n7993), .ZN(n8695) );
  AND2_X1 U8606 ( .A1(n8697), .A2(n8698), .ZN(n8696) );
  AND2_X1 U8607 ( .A1(n7996), .A2(n7995), .ZN(n8694) );
  XNOR2_X1 U8608 ( .A(n8699), .B(n8700), .ZN(n7995) );
  XOR2_X1 U8609 ( .A(n8701), .B(n8702), .Z(n8700) );
  INV_X1 U8610 ( .A(n8475), .ZN(n7996) );
  OR2_X1 U8611 ( .A1(n8703), .A2(n8704), .ZN(n8475) );
  AND2_X1 U8612 ( .A1(n8479), .A2(n8478), .ZN(n8704) );
  AND2_X1 U8613 ( .A1(n8476), .A2(n8705), .ZN(n8703) );
  OR2_X1 U8614 ( .A1(n8478), .A2(n8479), .ZN(n8705) );
  OR2_X1 U8615 ( .A1(n7621), .A2(n8355), .ZN(n8479) );
  OR2_X1 U8616 ( .A1(n8706), .A2(n8707), .ZN(n8478) );
  AND2_X1 U8617 ( .A1(n8693), .A2(n8692), .ZN(n8707) );
  AND2_X1 U8618 ( .A1(n8690), .A2(n8708), .ZN(n8706) );
  OR2_X1 U8619 ( .A1(n8692), .A2(n8693), .ZN(n8708) );
  OR2_X1 U8620 ( .A1(n7656), .A2(n8355), .ZN(n8693) );
  OR2_X1 U8621 ( .A1(n8709), .A2(n8710), .ZN(n8692) );
  AND2_X1 U8622 ( .A1(n8689), .A2(n8688), .ZN(n8710) );
  AND2_X1 U8623 ( .A1(n8687), .A2(n8711), .ZN(n8709) );
  OR2_X1 U8624 ( .A1(n8688), .A2(n8689), .ZN(n8711) );
  OR2_X1 U8625 ( .A1(n8712), .A2(n8713), .ZN(n8689) );
  AND2_X1 U8626 ( .A1(n8685), .A2(n8684), .ZN(n8713) );
  AND2_X1 U8627 ( .A1(n8682), .A2(n8714), .ZN(n8712) );
  OR2_X1 U8628 ( .A1(n8684), .A2(n8685), .ZN(n8714) );
  OR2_X1 U8629 ( .A1(n7777), .A2(n8355), .ZN(n8685) );
  OR2_X1 U8630 ( .A1(n8715), .A2(n8716), .ZN(n8684) );
  AND2_X1 U8631 ( .A1(n8681), .A2(n8680), .ZN(n8716) );
  AND2_X1 U8632 ( .A1(n8678), .A2(n8717), .ZN(n8715) );
  OR2_X1 U8633 ( .A1(n8680), .A2(n8681), .ZN(n8717) );
  OR2_X1 U8634 ( .A1(n7785), .A2(n8355), .ZN(n8681) );
  OR2_X1 U8635 ( .A1(n8718), .A2(n8719), .ZN(n8680) );
  AND2_X1 U8636 ( .A1(n8677), .A2(n8676), .ZN(n8719) );
  AND2_X1 U8637 ( .A1(n8674), .A2(n8720), .ZN(n8718) );
  OR2_X1 U8638 ( .A1(n8676), .A2(n8677), .ZN(n8720) );
  OR2_X1 U8639 ( .A1(n8226), .A2(n8355), .ZN(n8677) );
  OR2_X1 U8640 ( .A1(n8721), .A2(n8722), .ZN(n8676) );
  AND2_X1 U8641 ( .A1(n8673), .A2(n8672), .ZN(n8722) );
  AND2_X1 U8642 ( .A1(n8670), .A2(n8723), .ZN(n8721) );
  OR2_X1 U8643 ( .A1(n8672), .A2(n8673), .ZN(n8723) );
  OR2_X1 U8644 ( .A1(n8221), .A2(n8355), .ZN(n8673) );
  OR2_X1 U8645 ( .A1(n8724), .A2(n8725), .ZN(n8672) );
  AND2_X1 U8646 ( .A1(n8669), .A2(n8668), .ZN(n8725) );
  AND2_X1 U8647 ( .A1(n8666), .A2(n8726), .ZN(n8724) );
  OR2_X1 U8648 ( .A1(n8668), .A2(n8669), .ZN(n8726) );
  OR2_X1 U8649 ( .A1(n8216), .A2(n8355), .ZN(n8669) );
  OR2_X1 U8650 ( .A1(n8727), .A2(n8728), .ZN(n8668) );
  AND2_X1 U8651 ( .A1(n8665), .A2(n8664), .ZN(n8728) );
  AND2_X1 U8652 ( .A1(n8662), .A2(n8729), .ZN(n8727) );
  OR2_X1 U8653 ( .A1(n8664), .A2(n8665), .ZN(n8729) );
  OR2_X1 U8654 ( .A1(n8211), .A2(n8355), .ZN(n8665) );
  OR2_X1 U8655 ( .A1(n8730), .A2(n8731), .ZN(n8664) );
  AND2_X1 U8656 ( .A1(n8661), .A2(n8660), .ZN(n8731) );
  AND2_X1 U8657 ( .A1(n8658), .A2(n8732), .ZN(n8730) );
  OR2_X1 U8658 ( .A1(n8660), .A2(n8661), .ZN(n8732) );
  OR2_X1 U8659 ( .A1(n8206), .A2(n8355), .ZN(n8661) );
  OR2_X1 U8660 ( .A1(n8733), .A2(n8734), .ZN(n8660) );
  AND2_X1 U8661 ( .A1(n8657), .A2(n8656), .ZN(n8734) );
  AND2_X1 U8662 ( .A1(n8654), .A2(n8735), .ZN(n8733) );
  OR2_X1 U8663 ( .A1(n8656), .A2(n8657), .ZN(n8735) );
  OR2_X1 U8664 ( .A1(n8201), .A2(n8355), .ZN(n8657) );
  OR2_X1 U8665 ( .A1(n8736), .A2(n8737), .ZN(n8656) );
  AND2_X1 U8666 ( .A1(n8653), .A2(n8652), .ZN(n8737) );
  AND2_X1 U8667 ( .A1(n8650), .A2(n8738), .ZN(n8736) );
  OR2_X1 U8668 ( .A1(n8652), .A2(n8653), .ZN(n8738) );
  OR2_X1 U8669 ( .A1(n8196), .A2(n8355), .ZN(n8653) );
  OR2_X1 U8670 ( .A1(n8739), .A2(n8740), .ZN(n8652) );
  AND2_X1 U8671 ( .A1(n8649), .A2(n8648), .ZN(n8740) );
  AND2_X1 U8672 ( .A1(n8646), .A2(n8741), .ZN(n8739) );
  OR2_X1 U8673 ( .A1(n8648), .A2(n8649), .ZN(n8741) );
  OR2_X1 U8674 ( .A1(n8191), .A2(n8355), .ZN(n8649) );
  OR2_X1 U8675 ( .A1(n8742), .A2(n8743), .ZN(n8648) );
  AND2_X1 U8676 ( .A1(n8645), .A2(n8644), .ZN(n8743) );
  AND2_X1 U8677 ( .A1(n8642), .A2(n8744), .ZN(n8742) );
  OR2_X1 U8678 ( .A1(n8644), .A2(n8645), .ZN(n8744) );
  OR2_X1 U8679 ( .A1(n8186), .A2(n8355), .ZN(n8645) );
  OR2_X1 U8680 ( .A1(n8745), .A2(n8746), .ZN(n8644) );
  AND2_X1 U8681 ( .A1(n8641), .A2(n8640), .ZN(n8746) );
  AND2_X1 U8682 ( .A1(n8638), .A2(n8747), .ZN(n8745) );
  OR2_X1 U8683 ( .A1(n8640), .A2(n8641), .ZN(n8747) );
  OR2_X1 U8684 ( .A1(n8181), .A2(n8355), .ZN(n8641) );
  OR2_X1 U8685 ( .A1(n8748), .A2(n8749), .ZN(n8640) );
  AND2_X1 U8686 ( .A1(n8637), .A2(n8636), .ZN(n8749) );
  AND2_X1 U8687 ( .A1(n8634), .A2(n8750), .ZN(n8748) );
  OR2_X1 U8688 ( .A1(n8636), .A2(n8637), .ZN(n8750) );
  OR2_X1 U8689 ( .A1(n8176), .A2(n8355), .ZN(n8637) );
  OR2_X1 U8690 ( .A1(n8751), .A2(n8752), .ZN(n8636) );
  AND2_X1 U8691 ( .A1(n8633), .A2(n8632), .ZN(n8752) );
  AND2_X1 U8692 ( .A1(n8630), .A2(n8753), .ZN(n8751) );
  OR2_X1 U8693 ( .A1(n8632), .A2(n8633), .ZN(n8753) );
  OR2_X1 U8694 ( .A1(n8171), .A2(n8355), .ZN(n8633) );
  OR2_X1 U8695 ( .A1(n8754), .A2(n8755), .ZN(n8632) );
  AND2_X1 U8696 ( .A1(n8629), .A2(n8628), .ZN(n8755) );
  AND2_X1 U8697 ( .A1(n8626), .A2(n8756), .ZN(n8754) );
  OR2_X1 U8698 ( .A1(n8628), .A2(n8629), .ZN(n8756) );
  OR2_X1 U8699 ( .A1(n8166), .A2(n8355), .ZN(n8629) );
  OR2_X1 U8700 ( .A1(n8757), .A2(n8758), .ZN(n8628) );
  AND2_X1 U8701 ( .A1(n8625), .A2(n8624), .ZN(n8758) );
  AND2_X1 U8702 ( .A1(n8622), .A2(n8759), .ZN(n8757) );
  OR2_X1 U8703 ( .A1(n8624), .A2(n8625), .ZN(n8759) );
  OR2_X1 U8704 ( .A1(n8161), .A2(n8355), .ZN(n8625) );
  OR2_X1 U8705 ( .A1(n8760), .A2(n8761), .ZN(n8624) );
  AND2_X1 U8706 ( .A1(n8621), .A2(n8620), .ZN(n8761) );
  AND2_X1 U8707 ( .A1(n8618), .A2(n8762), .ZN(n8760) );
  OR2_X1 U8708 ( .A1(n8620), .A2(n8621), .ZN(n8762) );
  OR2_X1 U8709 ( .A1(n8156), .A2(n8355), .ZN(n8621) );
  OR2_X1 U8710 ( .A1(n8763), .A2(n8764), .ZN(n8620) );
  AND2_X1 U8711 ( .A1(n8617), .A2(n8616), .ZN(n8764) );
  AND2_X1 U8712 ( .A1(n8614), .A2(n8765), .ZN(n8763) );
  OR2_X1 U8713 ( .A1(n8616), .A2(n8617), .ZN(n8765) );
  OR2_X1 U8714 ( .A1(n8151), .A2(n8355), .ZN(n8617) );
  OR2_X1 U8715 ( .A1(n8766), .A2(n8767), .ZN(n8616) );
  AND2_X1 U8716 ( .A1(n8613), .A2(n8612), .ZN(n8767) );
  AND2_X1 U8717 ( .A1(n8610), .A2(n8768), .ZN(n8766) );
  OR2_X1 U8718 ( .A1(n8612), .A2(n8613), .ZN(n8768) );
  OR2_X1 U8719 ( .A1(n8146), .A2(n8355), .ZN(n8613) );
  OR2_X1 U8720 ( .A1(n8769), .A2(n8770), .ZN(n8612) );
  AND2_X1 U8721 ( .A1(n8609), .A2(n8608), .ZN(n8770) );
  AND2_X1 U8722 ( .A1(n8606), .A2(n8771), .ZN(n8769) );
  OR2_X1 U8723 ( .A1(n8608), .A2(n8609), .ZN(n8771) );
  OR2_X1 U8724 ( .A1(n8141), .A2(n8355), .ZN(n8609) );
  OR2_X1 U8725 ( .A1(n8772), .A2(n8773), .ZN(n8608) );
  AND2_X1 U8726 ( .A1(n8605), .A2(n8604), .ZN(n8773) );
  AND2_X1 U8727 ( .A1(n8602), .A2(n8774), .ZN(n8772) );
  OR2_X1 U8728 ( .A1(n8604), .A2(n8605), .ZN(n8774) );
  OR2_X1 U8729 ( .A1(n8136), .A2(n8355), .ZN(n8605) );
  OR2_X1 U8730 ( .A1(n8775), .A2(n8776), .ZN(n8604) );
  AND2_X1 U8731 ( .A1(n8601), .A2(n8600), .ZN(n8776) );
  AND2_X1 U8732 ( .A1(n8598), .A2(n8777), .ZN(n8775) );
  OR2_X1 U8733 ( .A1(n8600), .A2(n8601), .ZN(n8777) );
  OR2_X1 U8734 ( .A1(n8131), .A2(n8355), .ZN(n8601) );
  OR2_X1 U8735 ( .A1(n8778), .A2(n8779), .ZN(n8600) );
  AND2_X1 U8736 ( .A1(n8597), .A2(n8596), .ZN(n8779) );
  AND2_X1 U8737 ( .A1(n8594), .A2(n8780), .ZN(n8778) );
  OR2_X1 U8738 ( .A1(n8596), .A2(n8597), .ZN(n8780) );
  OR2_X1 U8739 ( .A1(n8126), .A2(n8355), .ZN(n8597) );
  OR2_X1 U8740 ( .A1(n8781), .A2(n8782), .ZN(n8596) );
  AND2_X1 U8741 ( .A1(n8593), .A2(n8592), .ZN(n8782) );
  AND2_X1 U8742 ( .A1(n8590), .A2(n8783), .ZN(n8781) );
  OR2_X1 U8743 ( .A1(n8592), .A2(n8593), .ZN(n8783) );
  OR2_X1 U8744 ( .A1(n8121), .A2(n8355), .ZN(n8593) );
  OR2_X1 U8745 ( .A1(n8784), .A2(n8785), .ZN(n8592) );
  AND2_X1 U8746 ( .A1(n8589), .A2(n8588), .ZN(n8785) );
  AND2_X1 U8747 ( .A1(n8586), .A2(n8786), .ZN(n8784) );
  OR2_X1 U8748 ( .A1(n8588), .A2(n8589), .ZN(n8786) );
  OR2_X1 U8749 ( .A1(n8116), .A2(n8355), .ZN(n8589) );
  OR2_X1 U8750 ( .A1(n8787), .A2(n8788), .ZN(n8588) );
  AND2_X1 U8751 ( .A1(n8583), .A2(n8585), .ZN(n8788) );
  AND2_X1 U8752 ( .A1(n8789), .A2(n8584), .ZN(n8787) );
  OR2_X1 U8753 ( .A1(n8585), .A2(n8583), .ZN(n8789) );
  XNOR2_X1 U8754 ( .A(n8790), .B(n8791), .ZN(n8583) );
  XNOR2_X1 U8755 ( .A(n8792), .B(n8793), .ZN(n8791) );
  OR2_X1 U8756 ( .A1(n8794), .A2(n8795), .ZN(n8585) );
  AND2_X1 U8757 ( .A1(n8578), .A2(n8581), .ZN(n8795) );
  AND2_X1 U8758 ( .A1(n8580), .A2(n8796), .ZN(n8794) );
  OR2_X1 U8759 ( .A1(n8581), .A2(n8578), .ZN(n8796) );
  OR2_X1 U8760 ( .A1(n8102), .A2(n8355), .ZN(n8578) );
  OR3_X1 U8761 ( .A1(n8349), .A2(n8355), .A3(n8575), .ZN(n8581) );
  INV_X1 U8762 ( .A(n8797), .ZN(n8580) );
  OR2_X1 U8763 ( .A1(n8798), .A2(n8799), .ZN(n8797) );
  AND2_X1 U8764 ( .A1(b_27_), .A2(n8800), .ZN(n8799) );
  OR2_X1 U8765 ( .A1(n8801), .A2(n7314), .ZN(n8800) );
  AND2_X1 U8766 ( .A1(a_30_), .A2(n8802), .ZN(n8801) );
  AND2_X1 U8767 ( .A1(b_26_), .A2(n8803), .ZN(n8798) );
  OR2_X1 U8768 ( .A1(n8804), .A2(n7318), .ZN(n8803) );
  AND2_X1 U8769 ( .A1(a_31_), .A2(n8575), .ZN(n8804) );
  XOR2_X1 U8770 ( .A(n8805), .B(n8806), .Z(n8586) );
  XOR2_X1 U8771 ( .A(n8807), .B(n8808), .Z(n8806) );
  XNOR2_X1 U8772 ( .A(n8809), .B(n8810), .ZN(n8590) );
  XNOR2_X1 U8773 ( .A(n8811), .B(n8812), .ZN(n8809) );
  XOR2_X1 U8774 ( .A(n8813), .B(n8814), .Z(n8594) );
  XOR2_X1 U8775 ( .A(n8815), .B(n8816), .Z(n8814) );
  XOR2_X1 U8776 ( .A(n8817), .B(n8818), .Z(n8598) );
  XOR2_X1 U8777 ( .A(n8819), .B(n8820), .Z(n8818) );
  XOR2_X1 U8778 ( .A(n8821), .B(n8822), .Z(n8602) );
  XOR2_X1 U8779 ( .A(n8823), .B(n8824), .Z(n8822) );
  XOR2_X1 U8780 ( .A(n8825), .B(n8826), .Z(n8606) );
  XOR2_X1 U8781 ( .A(n8827), .B(n8828), .Z(n8826) );
  XOR2_X1 U8782 ( .A(n8829), .B(n8830), .Z(n8610) );
  XOR2_X1 U8783 ( .A(n8831), .B(n8832), .Z(n8830) );
  XOR2_X1 U8784 ( .A(n8833), .B(n8834), .Z(n8614) );
  XOR2_X1 U8785 ( .A(n8835), .B(n8836), .Z(n8834) );
  XOR2_X1 U8786 ( .A(n8837), .B(n8838), .Z(n8618) );
  XOR2_X1 U8787 ( .A(n8839), .B(n8840), .Z(n8838) );
  XOR2_X1 U8788 ( .A(n8841), .B(n8842), .Z(n8622) );
  XOR2_X1 U8789 ( .A(n8843), .B(n8844), .Z(n8842) );
  XOR2_X1 U8790 ( .A(n8845), .B(n8846), .Z(n8626) );
  XOR2_X1 U8791 ( .A(n8847), .B(n8848), .Z(n8846) );
  XOR2_X1 U8792 ( .A(n8849), .B(n8850), .Z(n8630) );
  XOR2_X1 U8793 ( .A(n8851), .B(n8852), .Z(n8850) );
  XOR2_X1 U8794 ( .A(n8853), .B(n8854), .Z(n8634) );
  XOR2_X1 U8795 ( .A(n8855), .B(n8856), .Z(n8854) );
  XOR2_X1 U8796 ( .A(n8857), .B(n8858), .Z(n8638) );
  XOR2_X1 U8797 ( .A(n8859), .B(n8860), .Z(n8858) );
  XOR2_X1 U8798 ( .A(n8861), .B(n8862), .Z(n8642) );
  XOR2_X1 U8799 ( .A(n8863), .B(n8864), .Z(n8862) );
  XOR2_X1 U8800 ( .A(n8865), .B(n8866), .Z(n8646) );
  XOR2_X1 U8801 ( .A(n8867), .B(n8868), .Z(n8866) );
  XOR2_X1 U8802 ( .A(n8869), .B(n8870), .Z(n8650) );
  XOR2_X1 U8803 ( .A(n8871), .B(n8872), .Z(n8870) );
  XOR2_X1 U8804 ( .A(n8873), .B(n8874), .Z(n8654) );
  XOR2_X1 U8805 ( .A(n8875), .B(n8876), .Z(n8874) );
  XOR2_X1 U8806 ( .A(n8877), .B(n8878), .Z(n8658) );
  XOR2_X1 U8807 ( .A(n8879), .B(n8880), .Z(n8878) );
  XOR2_X1 U8808 ( .A(n8881), .B(n8882), .Z(n8662) );
  XOR2_X1 U8809 ( .A(n8883), .B(n8884), .Z(n8882) );
  XOR2_X1 U8810 ( .A(n8885), .B(n8886), .Z(n8666) );
  XOR2_X1 U8811 ( .A(n8887), .B(n8888), .Z(n8886) );
  XOR2_X1 U8812 ( .A(n8889), .B(n8890), .Z(n8670) );
  XOR2_X1 U8813 ( .A(n8891), .B(n8892), .Z(n8890) );
  XNOR2_X1 U8814 ( .A(n8893), .B(n8894), .ZN(n8674) );
  XNOR2_X1 U8815 ( .A(n8895), .B(n8896), .ZN(n8893) );
  XOR2_X1 U8816 ( .A(n8897), .B(n8898), .Z(n8678) );
  XOR2_X1 U8817 ( .A(n8899), .B(n8900), .Z(n8898) );
  XOR2_X1 U8818 ( .A(n8901), .B(n8902), .Z(n8682) );
  XOR2_X1 U8819 ( .A(n8903), .B(n8904), .Z(n8902) );
  OR2_X1 U8820 ( .A1(n7689), .A2(n8355), .ZN(n8688) );
  XOR2_X1 U8821 ( .A(n8905), .B(n8906), .Z(n8687) );
  XOR2_X1 U8822 ( .A(n8907), .B(n8908), .Z(n8906) );
  XNOR2_X1 U8823 ( .A(n8909), .B(n8910), .ZN(n8690) );
  XNOR2_X1 U8824 ( .A(n8911), .B(n8912), .ZN(n8909) );
  XOR2_X1 U8825 ( .A(n8913), .B(n8914), .Z(n8476) );
  XOR2_X1 U8826 ( .A(n8915), .B(n8916), .Z(n8914) );
  OR2_X1 U8827 ( .A1(n7993), .A2(n7992), .ZN(n7485) );
  XNOR2_X1 U8828 ( .A(n7988), .B(n8917), .ZN(n7992) );
  INV_X1 U8829 ( .A(n8918), .ZN(n7993) );
  OR2_X1 U8830 ( .A1(n8697), .A2(n8698), .ZN(n8918) );
  OR2_X1 U8831 ( .A1(n8919), .A2(n8920), .ZN(n8698) );
  AND2_X1 U8832 ( .A1(n8699), .A2(n8702), .ZN(n8920) );
  AND2_X1 U8833 ( .A1(n8921), .A2(n8701), .ZN(n8919) );
  OR2_X1 U8834 ( .A1(n8922), .A2(n8923), .ZN(n8701) );
  AND2_X1 U8835 ( .A1(n8913), .A2(n8916), .ZN(n8923) );
  AND2_X1 U8836 ( .A1(n8924), .A2(n8915), .ZN(n8922) );
  OR2_X1 U8837 ( .A1(n8925), .A2(n8926), .ZN(n8915) );
  AND2_X1 U8838 ( .A1(n8912), .A2(n8911), .ZN(n8926) );
  AND2_X1 U8839 ( .A1(n8910), .A2(n8927), .ZN(n8925) );
  OR2_X1 U8840 ( .A1(n8911), .A2(n8912), .ZN(n8927) );
  OR2_X1 U8841 ( .A1(n8928), .A2(n8929), .ZN(n8912) );
  AND2_X1 U8842 ( .A1(n8908), .A2(n8907), .ZN(n8929) );
  AND2_X1 U8843 ( .A1(n8905), .A2(n8930), .ZN(n8928) );
  OR2_X1 U8844 ( .A1(n8907), .A2(n8908), .ZN(n8930) );
  OR2_X1 U8845 ( .A1(n7777), .A2(n8575), .ZN(n8908) );
  OR2_X1 U8846 ( .A1(n8931), .A2(n8932), .ZN(n8907) );
  AND2_X1 U8847 ( .A1(n8904), .A2(n8903), .ZN(n8932) );
  AND2_X1 U8848 ( .A1(n8901), .A2(n8933), .ZN(n8931) );
  OR2_X1 U8849 ( .A1(n8903), .A2(n8904), .ZN(n8933) );
  OR2_X1 U8850 ( .A1(n7785), .A2(n8575), .ZN(n8904) );
  OR2_X1 U8851 ( .A1(n8934), .A2(n8935), .ZN(n8903) );
  AND2_X1 U8852 ( .A1(n8900), .A2(n8899), .ZN(n8935) );
  AND2_X1 U8853 ( .A1(n8897), .A2(n8936), .ZN(n8934) );
  OR2_X1 U8854 ( .A1(n8899), .A2(n8900), .ZN(n8936) );
  OR2_X1 U8855 ( .A1(n8226), .A2(n8575), .ZN(n8900) );
  OR2_X1 U8856 ( .A1(n8937), .A2(n8938), .ZN(n8899) );
  AND2_X1 U8857 ( .A1(n8896), .A2(n8895), .ZN(n8938) );
  AND2_X1 U8858 ( .A1(n8894), .A2(n8939), .ZN(n8937) );
  OR2_X1 U8859 ( .A1(n8895), .A2(n8896), .ZN(n8939) );
  OR2_X1 U8860 ( .A1(n8940), .A2(n8941), .ZN(n8896) );
  AND2_X1 U8861 ( .A1(n8892), .A2(n8891), .ZN(n8941) );
  AND2_X1 U8862 ( .A1(n8889), .A2(n8942), .ZN(n8940) );
  OR2_X1 U8863 ( .A1(n8891), .A2(n8892), .ZN(n8942) );
  OR2_X1 U8864 ( .A1(n8216), .A2(n8575), .ZN(n8892) );
  OR2_X1 U8865 ( .A1(n8943), .A2(n8944), .ZN(n8891) );
  AND2_X1 U8866 ( .A1(n8888), .A2(n8887), .ZN(n8944) );
  AND2_X1 U8867 ( .A1(n8885), .A2(n8945), .ZN(n8943) );
  OR2_X1 U8868 ( .A1(n8887), .A2(n8888), .ZN(n8945) );
  OR2_X1 U8869 ( .A1(n8211), .A2(n8575), .ZN(n8888) );
  OR2_X1 U8870 ( .A1(n8946), .A2(n8947), .ZN(n8887) );
  AND2_X1 U8871 ( .A1(n8884), .A2(n8883), .ZN(n8947) );
  AND2_X1 U8872 ( .A1(n8881), .A2(n8948), .ZN(n8946) );
  OR2_X1 U8873 ( .A1(n8883), .A2(n8884), .ZN(n8948) );
  OR2_X1 U8874 ( .A1(n8206), .A2(n8575), .ZN(n8884) );
  OR2_X1 U8875 ( .A1(n8949), .A2(n8950), .ZN(n8883) );
  AND2_X1 U8876 ( .A1(n8880), .A2(n8879), .ZN(n8950) );
  AND2_X1 U8877 ( .A1(n8877), .A2(n8951), .ZN(n8949) );
  OR2_X1 U8878 ( .A1(n8879), .A2(n8880), .ZN(n8951) );
  OR2_X1 U8879 ( .A1(n8201), .A2(n8575), .ZN(n8880) );
  OR2_X1 U8880 ( .A1(n8952), .A2(n8953), .ZN(n8879) );
  AND2_X1 U8881 ( .A1(n8876), .A2(n8875), .ZN(n8953) );
  AND2_X1 U8882 ( .A1(n8873), .A2(n8954), .ZN(n8952) );
  OR2_X1 U8883 ( .A1(n8875), .A2(n8876), .ZN(n8954) );
  OR2_X1 U8884 ( .A1(n8196), .A2(n8575), .ZN(n8876) );
  OR2_X1 U8885 ( .A1(n8955), .A2(n8956), .ZN(n8875) );
  AND2_X1 U8886 ( .A1(n8872), .A2(n8871), .ZN(n8956) );
  AND2_X1 U8887 ( .A1(n8869), .A2(n8957), .ZN(n8955) );
  OR2_X1 U8888 ( .A1(n8871), .A2(n8872), .ZN(n8957) );
  OR2_X1 U8889 ( .A1(n8191), .A2(n8575), .ZN(n8872) );
  OR2_X1 U8890 ( .A1(n8958), .A2(n8959), .ZN(n8871) );
  AND2_X1 U8891 ( .A1(n8868), .A2(n8867), .ZN(n8959) );
  AND2_X1 U8892 ( .A1(n8865), .A2(n8960), .ZN(n8958) );
  OR2_X1 U8893 ( .A1(n8867), .A2(n8868), .ZN(n8960) );
  OR2_X1 U8894 ( .A1(n8186), .A2(n8575), .ZN(n8868) );
  OR2_X1 U8895 ( .A1(n8961), .A2(n8962), .ZN(n8867) );
  AND2_X1 U8896 ( .A1(n8864), .A2(n8863), .ZN(n8962) );
  AND2_X1 U8897 ( .A1(n8861), .A2(n8963), .ZN(n8961) );
  OR2_X1 U8898 ( .A1(n8863), .A2(n8864), .ZN(n8963) );
  OR2_X1 U8899 ( .A1(n8181), .A2(n8575), .ZN(n8864) );
  OR2_X1 U8900 ( .A1(n8964), .A2(n8965), .ZN(n8863) );
  AND2_X1 U8901 ( .A1(n8860), .A2(n8859), .ZN(n8965) );
  AND2_X1 U8902 ( .A1(n8857), .A2(n8966), .ZN(n8964) );
  OR2_X1 U8903 ( .A1(n8859), .A2(n8860), .ZN(n8966) );
  OR2_X1 U8904 ( .A1(n8176), .A2(n8575), .ZN(n8860) );
  OR2_X1 U8905 ( .A1(n8967), .A2(n8968), .ZN(n8859) );
  AND2_X1 U8906 ( .A1(n8856), .A2(n8855), .ZN(n8968) );
  AND2_X1 U8907 ( .A1(n8853), .A2(n8969), .ZN(n8967) );
  OR2_X1 U8908 ( .A1(n8855), .A2(n8856), .ZN(n8969) );
  OR2_X1 U8909 ( .A1(n8171), .A2(n8575), .ZN(n8856) );
  OR2_X1 U8910 ( .A1(n8970), .A2(n8971), .ZN(n8855) );
  AND2_X1 U8911 ( .A1(n8852), .A2(n8851), .ZN(n8971) );
  AND2_X1 U8912 ( .A1(n8849), .A2(n8972), .ZN(n8970) );
  OR2_X1 U8913 ( .A1(n8851), .A2(n8852), .ZN(n8972) );
  OR2_X1 U8914 ( .A1(n8166), .A2(n8575), .ZN(n8852) );
  OR2_X1 U8915 ( .A1(n8973), .A2(n8974), .ZN(n8851) );
  AND2_X1 U8916 ( .A1(n8848), .A2(n8847), .ZN(n8974) );
  AND2_X1 U8917 ( .A1(n8845), .A2(n8975), .ZN(n8973) );
  OR2_X1 U8918 ( .A1(n8847), .A2(n8848), .ZN(n8975) );
  OR2_X1 U8919 ( .A1(n8161), .A2(n8575), .ZN(n8848) );
  OR2_X1 U8920 ( .A1(n8976), .A2(n8977), .ZN(n8847) );
  AND2_X1 U8921 ( .A1(n8844), .A2(n8843), .ZN(n8977) );
  AND2_X1 U8922 ( .A1(n8841), .A2(n8978), .ZN(n8976) );
  OR2_X1 U8923 ( .A1(n8843), .A2(n8844), .ZN(n8978) );
  OR2_X1 U8924 ( .A1(n8156), .A2(n8575), .ZN(n8844) );
  OR2_X1 U8925 ( .A1(n8979), .A2(n8980), .ZN(n8843) );
  AND2_X1 U8926 ( .A1(n8840), .A2(n8839), .ZN(n8980) );
  AND2_X1 U8927 ( .A1(n8837), .A2(n8981), .ZN(n8979) );
  OR2_X1 U8928 ( .A1(n8839), .A2(n8840), .ZN(n8981) );
  OR2_X1 U8929 ( .A1(n8151), .A2(n8575), .ZN(n8840) );
  OR2_X1 U8930 ( .A1(n8982), .A2(n8983), .ZN(n8839) );
  AND2_X1 U8931 ( .A1(n8836), .A2(n8835), .ZN(n8983) );
  AND2_X1 U8932 ( .A1(n8833), .A2(n8984), .ZN(n8982) );
  OR2_X1 U8933 ( .A1(n8835), .A2(n8836), .ZN(n8984) );
  OR2_X1 U8934 ( .A1(n8146), .A2(n8575), .ZN(n8836) );
  OR2_X1 U8935 ( .A1(n8985), .A2(n8986), .ZN(n8835) );
  AND2_X1 U8936 ( .A1(n8832), .A2(n8831), .ZN(n8986) );
  AND2_X1 U8937 ( .A1(n8829), .A2(n8987), .ZN(n8985) );
  OR2_X1 U8938 ( .A1(n8831), .A2(n8832), .ZN(n8987) );
  OR2_X1 U8939 ( .A1(n8141), .A2(n8575), .ZN(n8832) );
  OR2_X1 U8940 ( .A1(n8988), .A2(n8989), .ZN(n8831) );
  AND2_X1 U8941 ( .A1(n8828), .A2(n8827), .ZN(n8989) );
  AND2_X1 U8942 ( .A1(n8825), .A2(n8990), .ZN(n8988) );
  OR2_X1 U8943 ( .A1(n8827), .A2(n8828), .ZN(n8990) );
  OR2_X1 U8944 ( .A1(n8136), .A2(n8575), .ZN(n8828) );
  OR2_X1 U8945 ( .A1(n8991), .A2(n8992), .ZN(n8827) );
  AND2_X1 U8946 ( .A1(n8824), .A2(n8823), .ZN(n8992) );
  AND2_X1 U8947 ( .A1(n8821), .A2(n8993), .ZN(n8991) );
  OR2_X1 U8948 ( .A1(n8823), .A2(n8824), .ZN(n8993) );
  OR2_X1 U8949 ( .A1(n8131), .A2(n8575), .ZN(n8824) );
  OR2_X1 U8950 ( .A1(n8994), .A2(n8995), .ZN(n8823) );
  AND2_X1 U8951 ( .A1(n8820), .A2(n8819), .ZN(n8995) );
  AND2_X1 U8952 ( .A1(n8817), .A2(n8996), .ZN(n8994) );
  OR2_X1 U8953 ( .A1(n8819), .A2(n8820), .ZN(n8996) );
  OR2_X1 U8954 ( .A1(n8126), .A2(n8575), .ZN(n8820) );
  OR2_X1 U8955 ( .A1(n8997), .A2(n8998), .ZN(n8819) );
  AND2_X1 U8956 ( .A1(n8816), .A2(n8815), .ZN(n8998) );
  AND2_X1 U8957 ( .A1(n8813), .A2(n8999), .ZN(n8997) );
  OR2_X1 U8958 ( .A1(n8815), .A2(n8816), .ZN(n8999) );
  OR2_X1 U8959 ( .A1(n8121), .A2(n8575), .ZN(n8816) );
  OR2_X1 U8960 ( .A1(n9000), .A2(n9001), .ZN(n8815) );
  AND2_X1 U8961 ( .A1(n8810), .A2(n8812), .ZN(n9001) );
  AND2_X1 U8962 ( .A1(n9002), .A2(n8811), .ZN(n9000) );
  OR2_X1 U8963 ( .A1(n8812), .A2(n8810), .ZN(n9002) );
  XOR2_X1 U8964 ( .A(n9003), .B(n9004), .Z(n8810) );
  XOR2_X1 U8965 ( .A(n9005), .B(n9006), .Z(n9004) );
  OR2_X1 U8966 ( .A1(n9007), .A2(n9008), .ZN(n8812) );
  AND2_X1 U8967 ( .A1(n8808), .A2(n8807), .ZN(n9008) );
  AND2_X1 U8968 ( .A1(n8805), .A2(n9009), .ZN(n9007) );
  OR2_X1 U8969 ( .A1(n8807), .A2(n8808), .ZN(n9009) );
  OR2_X1 U8970 ( .A1(n8111), .A2(n8575), .ZN(n8808) );
  OR2_X1 U8971 ( .A1(n9010), .A2(n9011), .ZN(n8807) );
  AND2_X1 U8972 ( .A1(n8790), .A2(n8793), .ZN(n9011) );
  AND2_X1 U8973 ( .A1(n8792), .A2(n9012), .ZN(n9010) );
  OR2_X1 U8974 ( .A1(n8793), .A2(n8790), .ZN(n9012) );
  OR2_X1 U8975 ( .A1(n8102), .A2(n8575), .ZN(n8790) );
  OR3_X1 U8976 ( .A1(n8349), .A2(n8575), .A3(n8802), .ZN(n8793) );
  INV_X1 U8977 ( .A(n9013), .ZN(n8792) );
  OR2_X1 U8978 ( .A1(n9014), .A2(n9015), .ZN(n9013) );
  AND2_X1 U8979 ( .A1(b_26_), .A2(n9016), .ZN(n9015) );
  OR2_X1 U8980 ( .A1(n9017), .A2(n7314), .ZN(n9016) );
  AND2_X1 U8981 ( .A1(a_30_), .A2(n9018), .ZN(n9017) );
  AND2_X1 U8982 ( .A1(b_25_), .A2(n9019), .ZN(n9014) );
  OR2_X1 U8983 ( .A1(n9020), .A2(n7318), .ZN(n9019) );
  AND2_X1 U8984 ( .A1(a_31_), .A2(n8802), .ZN(n9020) );
  XNOR2_X1 U8985 ( .A(n9021), .B(n9022), .ZN(n8805) );
  XNOR2_X1 U8986 ( .A(n9023), .B(n9024), .ZN(n9022) );
  XOR2_X1 U8987 ( .A(n9025), .B(n9026), .Z(n8813) );
  XOR2_X1 U8988 ( .A(n9027), .B(n9028), .Z(n9026) );
  XNOR2_X1 U8989 ( .A(n9029), .B(n9030), .ZN(n8817) );
  XNOR2_X1 U8990 ( .A(n9031), .B(n9032), .ZN(n9029) );
  XOR2_X1 U8991 ( .A(n9033), .B(n9034), .Z(n8821) );
  XOR2_X1 U8992 ( .A(n9035), .B(n9036), .Z(n9034) );
  XOR2_X1 U8993 ( .A(n9037), .B(n9038), .Z(n8825) );
  XOR2_X1 U8994 ( .A(n9039), .B(n9040), .Z(n9038) );
  XOR2_X1 U8995 ( .A(n9041), .B(n9042), .Z(n8829) );
  XOR2_X1 U8996 ( .A(n9043), .B(n9044), .Z(n9042) );
  XOR2_X1 U8997 ( .A(n9045), .B(n9046), .Z(n8833) );
  XOR2_X1 U8998 ( .A(n9047), .B(n9048), .Z(n9046) );
  XOR2_X1 U8999 ( .A(n9049), .B(n9050), .Z(n8837) );
  XOR2_X1 U9000 ( .A(n9051), .B(n9052), .Z(n9050) );
  XOR2_X1 U9001 ( .A(n9053), .B(n9054), .Z(n8841) );
  XOR2_X1 U9002 ( .A(n9055), .B(n9056), .Z(n9054) );
  XOR2_X1 U9003 ( .A(n9057), .B(n9058), .Z(n8845) );
  XOR2_X1 U9004 ( .A(n9059), .B(n9060), .Z(n9058) );
  XOR2_X1 U9005 ( .A(n9061), .B(n9062), .Z(n8849) );
  XOR2_X1 U9006 ( .A(n9063), .B(n9064), .Z(n9062) );
  XOR2_X1 U9007 ( .A(n9065), .B(n9066), .Z(n8853) );
  XOR2_X1 U9008 ( .A(n9067), .B(n9068), .Z(n9066) );
  XOR2_X1 U9009 ( .A(n9069), .B(n9070), .Z(n8857) );
  XOR2_X1 U9010 ( .A(n9071), .B(n9072), .Z(n9070) );
  XOR2_X1 U9011 ( .A(n9073), .B(n9074), .Z(n8861) );
  XOR2_X1 U9012 ( .A(n9075), .B(n9076), .Z(n9074) );
  XOR2_X1 U9013 ( .A(n9077), .B(n9078), .Z(n8865) );
  XOR2_X1 U9014 ( .A(n9079), .B(n9080), .Z(n9078) );
  XOR2_X1 U9015 ( .A(n9081), .B(n9082), .Z(n8869) );
  XOR2_X1 U9016 ( .A(n9083), .B(n9084), .Z(n9082) );
  XOR2_X1 U9017 ( .A(n9085), .B(n9086), .Z(n8873) );
  XOR2_X1 U9018 ( .A(n9087), .B(n9088), .Z(n9086) );
  XOR2_X1 U9019 ( .A(n9089), .B(n9090), .Z(n8877) );
  XOR2_X1 U9020 ( .A(n9091), .B(n9092), .Z(n9090) );
  XOR2_X1 U9021 ( .A(n9093), .B(n9094), .Z(n8881) );
  XOR2_X1 U9022 ( .A(n9095), .B(n9096), .Z(n9094) );
  XOR2_X1 U9023 ( .A(n9097), .B(n9098), .Z(n8885) );
  XOR2_X1 U9024 ( .A(n9099), .B(n9100), .Z(n9098) );
  XOR2_X1 U9025 ( .A(n9101), .B(n9102), .Z(n8889) );
  XOR2_X1 U9026 ( .A(n9103), .B(n9104), .Z(n9102) );
  OR2_X1 U9027 ( .A1(n8221), .A2(n8575), .ZN(n8895) );
  XOR2_X1 U9028 ( .A(n9105), .B(n9106), .Z(n8894) );
  XOR2_X1 U9029 ( .A(n9107), .B(n9108), .Z(n9106) );
  XNOR2_X1 U9030 ( .A(n9109), .B(n9110), .ZN(n8897) );
  XNOR2_X1 U9031 ( .A(n9111), .B(n9112), .ZN(n9109) );
  XOR2_X1 U9032 ( .A(n9113), .B(n9114), .Z(n8901) );
  XOR2_X1 U9033 ( .A(n9115), .B(n9116), .Z(n9114) );
  XOR2_X1 U9034 ( .A(n9117), .B(n9118), .Z(n8905) );
  XOR2_X1 U9035 ( .A(n9119), .B(n9120), .Z(n9118) );
  OR2_X1 U9036 ( .A1(n7689), .A2(n8575), .ZN(n8911) );
  XOR2_X1 U9037 ( .A(n9121), .B(n9122), .Z(n8910) );
  XOR2_X1 U9038 ( .A(n9123), .B(n9124), .Z(n9122) );
  OR2_X1 U9039 ( .A1(n8913), .A2(n8916), .ZN(n8924) );
  OR2_X1 U9040 ( .A1(n7656), .A2(n8575), .ZN(n8916) );
  XOR2_X1 U9041 ( .A(n9125), .B(n9126), .Z(n8913) );
  XOR2_X1 U9042 ( .A(n9127), .B(n9128), .Z(n9126) );
  OR2_X1 U9043 ( .A1(n8699), .A2(n8702), .ZN(n8921) );
  OR2_X1 U9044 ( .A1(n7621), .A2(n8575), .ZN(n8702) );
  XOR2_X1 U9045 ( .A(n9129), .B(n9130), .Z(n8699) );
  XOR2_X1 U9046 ( .A(n9131), .B(n9132), .Z(n9130) );
  XOR2_X1 U9047 ( .A(n9133), .B(n9134), .Z(n8697) );
  XOR2_X1 U9048 ( .A(n9135), .B(n9136), .Z(n9134) );
  OR2_X1 U9049 ( .A1(n9137), .A2(n7989), .ZN(n7491) );
  XOR2_X1 U9050 ( .A(n7964), .B(n7966), .Z(n7989) );
  OR2_X1 U9051 ( .A1(n9138), .A2(n9139), .ZN(n7966) );
  AND2_X1 U9052 ( .A1(n9140), .A2(n9141), .ZN(n9139) );
  AND2_X1 U9053 ( .A1(n9142), .A2(n9143), .ZN(n9138) );
  OR2_X1 U9054 ( .A1(n9140), .A2(n9141), .ZN(n9143) );
  XOR2_X1 U9055 ( .A(n7973), .B(n9144), .Z(n7964) );
  XOR2_X1 U9056 ( .A(n7972), .B(n7971), .Z(n9144) );
  OR2_X1 U9057 ( .A1(n7621), .A2(n9145), .ZN(n7971) );
  OR2_X1 U9058 ( .A1(n9146), .A2(n9147), .ZN(n7972) );
  AND2_X1 U9059 ( .A1(n9148), .A2(n9149), .ZN(n9147) );
  AND2_X1 U9060 ( .A1(n9150), .A2(n9151), .ZN(n9146) );
  OR2_X1 U9061 ( .A1(n9148), .A2(n9149), .ZN(n9151) );
  XOR2_X1 U9062 ( .A(n7981), .B(n9152), .Z(n7973) );
  XOR2_X1 U9063 ( .A(n7980), .B(n7979), .Z(n9152) );
  OR2_X1 U9064 ( .A1(n7656), .A2(n7976), .ZN(n7979) );
  OR2_X1 U9065 ( .A1(n9153), .A2(n9154), .ZN(n7980) );
  AND2_X1 U9066 ( .A1(n9155), .A2(n9156), .ZN(n9154) );
  AND2_X1 U9067 ( .A1(n9157), .A2(n9158), .ZN(n9153) );
  OR2_X1 U9068 ( .A1(n9155), .A2(n9156), .ZN(n9158) );
  XOR2_X1 U9069 ( .A(n9159), .B(n9160), .Z(n7981) );
  XOR2_X1 U9070 ( .A(n9161), .B(n9162), .Z(n9160) );
  AND2_X1 U9071 ( .A1(n7990), .A2(n7988), .ZN(n9137) );
  XNOR2_X1 U9072 ( .A(n9142), .B(n9163), .ZN(n7988) );
  XOR2_X1 U9073 ( .A(n9141), .B(n9140), .Z(n9163) );
  OR2_X1 U9074 ( .A1(n7621), .A2(n9018), .ZN(n9140) );
  OR2_X1 U9075 ( .A1(n9164), .A2(n9165), .ZN(n9141) );
  AND2_X1 U9076 ( .A1(n9166), .A2(n9167), .ZN(n9165) );
  AND2_X1 U9077 ( .A1(n9168), .A2(n9169), .ZN(n9164) );
  OR2_X1 U9078 ( .A1(n9166), .A2(n9167), .ZN(n9169) );
  XNOR2_X1 U9079 ( .A(n9170), .B(n9150), .ZN(n9142) );
  XOR2_X1 U9080 ( .A(n9157), .B(n9171), .Z(n9150) );
  XOR2_X1 U9081 ( .A(n9156), .B(n9155), .Z(n9171) );
  OR2_X1 U9082 ( .A1(n7689), .A2(n7976), .ZN(n9155) );
  OR2_X1 U9083 ( .A1(n9172), .A2(n9173), .ZN(n9156) );
  AND2_X1 U9084 ( .A1(n9174), .A2(n9175), .ZN(n9173) );
  AND2_X1 U9085 ( .A1(n9176), .A2(n9177), .ZN(n9172) );
  OR2_X1 U9086 ( .A1(n9174), .A2(n9175), .ZN(n9177) );
  XOR2_X1 U9087 ( .A(n9178), .B(n9179), .Z(n9157) );
  XOR2_X1 U9088 ( .A(n9180), .B(n9181), .Z(n9179) );
  XNOR2_X1 U9089 ( .A(n9149), .B(n9148), .ZN(n9170) );
  OR2_X1 U9090 ( .A1(n9182), .A2(n9183), .ZN(n9148) );
  AND2_X1 U9091 ( .A1(n9184), .A2(n9185), .ZN(n9183) );
  AND2_X1 U9092 ( .A1(n9186), .A2(n9187), .ZN(n9182) );
  OR2_X1 U9093 ( .A1(n9184), .A2(n9185), .ZN(n9187) );
  OR2_X1 U9094 ( .A1(n7656), .A2(n9145), .ZN(n9149) );
  INV_X1 U9095 ( .A(n8917), .ZN(n7990) );
  OR2_X1 U9096 ( .A1(n9188), .A2(n9189), .ZN(n8917) );
  AND2_X1 U9097 ( .A1(n9136), .A2(n9135), .ZN(n9189) );
  AND2_X1 U9098 ( .A1(n9133), .A2(n9190), .ZN(n9188) );
  OR2_X1 U9099 ( .A1(n9135), .A2(n9136), .ZN(n9190) );
  OR2_X1 U9100 ( .A1(n7621), .A2(n8802), .ZN(n9136) );
  OR2_X1 U9101 ( .A1(n9191), .A2(n9192), .ZN(n9135) );
  AND2_X1 U9102 ( .A1(n9132), .A2(n9131), .ZN(n9192) );
  AND2_X1 U9103 ( .A1(n9129), .A2(n9193), .ZN(n9191) );
  OR2_X1 U9104 ( .A1(n9131), .A2(n9132), .ZN(n9193) );
  OR2_X1 U9105 ( .A1(n7656), .A2(n8802), .ZN(n9132) );
  OR2_X1 U9106 ( .A1(n9194), .A2(n9195), .ZN(n9131) );
  AND2_X1 U9107 ( .A1(n9128), .A2(n9127), .ZN(n9195) );
  AND2_X1 U9108 ( .A1(n9125), .A2(n9196), .ZN(n9194) );
  OR2_X1 U9109 ( .A1(n9127), .A2(n9128), .ZN(n9196) );
  OR2_X1 U9110 ( .A1(n7689), .A2(n8802), .ZN(n9128) );
  OR2_X1 U9111 ( .A1(n9197), .A2(n9198), .ZN(n9127) );
  AND2_X1 U9112 ( .A1(n9124), .A2(n9123), .ZN(n9198) );
  AND2_X1 U9113 ( .A1(n9121), .A2(n9199), .ZN(n9197) );
  OR2_X1 U9114 ( .A1(n9123), .A2(n9124), .ZN(n9199) );
  OR2_X1 U9115 ( .A1(n7777), .A2(n8802), .ZN(n9124) );
  OR2_X1 U9116 ( .A1(n9200), .A2(n9201), .ZN(n9123) );
  AND2_X1 U9117 ( .A1(n9120), .A2(n9119), .ZN(n9201) );
  AND2_X1 U9118 ( .A1(n9117), .A2(n9202), .ZN(n9200) );
  OR2_X1 U9119 ( .A1(n9119), .A2(n9120), .ZN(n9202) );
  OR2_X1 U9120 ( .A1(n7785), .A2(n8802), .ZN(n9120) );
  OR2_X1 U9121 ( .A1(n9203), .A2(n9204), .ZN(n9119) );
  AND2_X1 U9122 ( .A1(n9116), .A2(n9115), .ZN(n9204) );
  AND2_X1 U9123 ( .A1(n9113), .A2(n9205), .ZN(n9203) );
  OR2_X1 U9124 ( .A1(n9115), .A2(n9116), .ZN(n9205) );
  OR2_X1 U9125 ( .A1(n8226), .A2(n8802), .ZN(n9116) );
  OR2_X1 U9126 ( .A1(n9206), .A2(n9207), .ZN(n9115) );
  AND2_X1 U9127 ( .A1(n9112), .A2(n9111), .ZN(n9207) );
  AND2_X1 U9128 ( .A1(n9110), .A2(n9208), .ZN(n9206) );
  OR2_X1 U9129 ( .A1(n9111), .A2(n9112), .ZN(n9208) );
  OR2_X1 U9130 ( .A1(n9209), .A2(n9210), .ZN(n9112) );
  AND2_X1 U9131 ( .A1(n9108), .A2(n9107), .ZN(n9210) );
  AND2_X1 U9132 ( .A1(n9105), .A2(n9211), .ZN(n9209) );
  OR2_X1 U9133 ( .A1(n9107), .A2(n9108), .ZN(n9211) );
  OR2_X1 U9134 ( .A1(n8216), .A2(n8802), .ZN(n9108) );
  OR2_X1 U9135 ( .A1(n9212), .A2(n9213), .ZN(n9107) );
  AND2_X1 U9136 ( .A1(n9104), .A2(n9103), .ZN(n9213) );
  AND2_X1 U9137 ( .A1(n9101), .A2(n9214), .ZN(n9212) );
  OR2_X1 U9138 ( .A1(n9103), .A2(n9104), .ZN(n9214) );
  OR2_X1 U9139 ( .A1(n8211), .A2(n8802), .ZN(n9104) );
  OR2_X1 U9140 ( .A1(n9215), .A2(n9216), .ZN(n9103) );
  AND2_X1 U9141 ( .A1(n9100), .A2(n9099), .ZN(n9216) );
  AND2_X1 U9142 ( .A1(n9097), .A2(n9217), .ZN(n9215) );
  OR2_X1 U9143 ( .A1(n9099), .A2(n9100), .ZN(n9217) );
  OR2_X1 U9144 ( .A1(n8206), .A2(n8802), .ZN(n9100) );
  OR2_X1 U9145 ( .A1(n9218), .A2(n9219), .ZN(n9099) );
  AND2_X1 U9146 ( .A1(n9096), .A2(n9095), .ZN(n9219) );
  AND2_X1 U9147 ( .A1(n9093), .A2(n9220), .ZN(n9218) );
  OR2_X1 U9148 ( .A1(n9095), .A2(n9096), .ZN(n9220) );
  OR2_X1 U9149 ( .A1(n8201), .A2(n8802), .ZN(n9096) );
  OR2_X1 U9150 ( .A1(n9221), .A2(n9222), .ZN(n9095) );
  AND2_X1 U9151 ( .A1(n9092), .A2(n9091), .ZN(n9222) );
  AND2_X1 U9152 ( .A1(n9089), .A2(n9223), .ZN(n9221) );
  OR2_X1 U9153 ( .A1(n9091), .A2(n9092), .ZN(n9223) );
  OR2_X1 U9154 ( .A1(n8196), .A2(n8802), .ZN(n9092) );
  OR2_X1 U9155 ( .A1(n9224), .A2(n9225), .ZN(n9091) );
  AND2_X1 U9156 ( .A1(n9088), .A2(n9087), .ZN(n9225) );
  AND2_X1 U9157 ( .A1(n9085), .A2(n9226), .ZN(n9224) );
  OR2_X1 U9158 ( .A1(n9087), .A2(n9088), .ZN(n9226) );
  OR2_X1 U9159 ( .A1(n8191), .A2(n8802), .ZN(n9088) );
  OR2_X1 U9160 ( .A1(n9227), .A2(n9228), .ZN(n9087) );
  AND2_X1 U9161 ( .A1(n9084), .A2(n9083), .ZN(n9228) );
  AND2_X1 U9162 ( .A1(n9081), .A2(n9229), .ZN(n9227) );
  OR2_X1 U9163 ( .A1(n9083), .A2(n9084), .ZN(n9229) );
  OR2_X1 U9164 ( .A1(n8186), .A2(n8802), .ZN(n9084) );
  OR2_X1 U9165 ( .A1(n9230), .A2(n9231), .ZN(n9083) );
  AND2_X1 U9166 ( .A1(n9080), .A2(n9079), .ZN(n9231) );
  AND2_X1 U9167 ( .A1(n9077), .A2(n9232), .ZN(n9230) );
  OR2_X1 U9168 ( .A1(n9079), .A2(n9080), .ZN(n9232) );
  OR2_X1 U9169 ( .A1(n8181), .A2(n8802), .ZN(n9080) );
  OR2_X1 U9170 ( .A1(n9233), .A2(n9234), .ZN(n9079) );
  AND2_X1 U9171 ( .A1(n9076), .A2(n9075), .ZN(n9234) );
  AND2_X1 U9172 ( .A1(n9073), .A2(n9235), .ZN(n9233) );
  OR2_X1 U9173 ( .A1(n9075), .A2(n9076), .ZN(n9235) );
  OR2_X1 U9174 ( .A1(n8176), .A2(n8802), .ZN(n9076) );
  OR2_X1 U9175 ( .A1(n9236), .A2(n9237), .ZN(n9075) );
  AND2_X1 U9176 ( .A1(n9072), .A2(n9071), .ZN(n9237) );
  AND2_X1 U9177 ( .A1(n9069), .A2(n9238), .ZN(n9236) );
  OR2_X1 U9178 ( .A1(n9071), .A2(n9072), .ZN(n9238) );
  OR2_X1 U9179 ( .A1(n8171), .A2(n8802), .ZN(n9072) );
  OR2_X1 U9180 ( .A1(n9239), .A2(n9240), .ZN(n9071) );
  AND2_X1 U9181 ( .A1(n9068), .A2(n9067), .ZN(n9240) );
  AND2_X1 U9182 ( .A1(n9065), .A2(n9241), .ZN(n9239) );
  OR2_X1 U9183 ( .A1(n9067), .A2(n9068), .ZN(n9241) );
  OR2_X1 U9184 ( .A1(n8166), .A2(n8802), .ZN(n9068) );
  OR2_X1 U9185 ( .A1(n9242), .A2(n9243), .ZN(n9067) );
  AND2_X1 U9186 ( .A1(n9064), .A2(n9063), .ZN(n9243) );
  AND2_X1 U9187 ( .A1(n9061), .A2(n9244), .ZN(n9242) );
  OR2_X1 U9188 ( .A1(n9063), .A2(n9064), .ZN(n9244) );
  OR2_X1 U9189 ( .A1(n8161), .A2(n8802), .ZN(n9064) );
  OR2_X1 U9190 ( .A1(n9245), .A2(n9246), .ZN(n9063) );
  AND2_X1 U9191 ( .A1(n9060), .A2(n9059), .ZN(n9246) );
  AND2_X1 U9192 ( .A1(n9057), .A2(n9247), .ZN(n9245) );
  OR2_X1 U9193 ( .A1(n9059), .A2(n9060), .ZN(n9247) );
  OR2_X1 U9194 ( .A1(n8156), .A2(n8802), .ZN(n9060) );
  OR2_X1 U9195 ( .A1(n9248), .A2(n9249), .ZN(n9059) );
  AND2_X1 U9196 ( .A1(n9056), .A2(n9055), .ZN(n9249) );
  AND2_X1 U9197 ( .A1(n9053), .A2(n9250), .ZN(n9248) );
  OR2_X1 U9198 ( .A1(n9055), .A2(n9056), .ZN(n9250) );
  OR2_X1 U9199 ( .A1(n8151), .A2(n8802), .ZN(n9056) );
  OR2_X1 U9200 ( .A1(n9251), .A2(n9252), .ZN(n9055) );
  AND2_X1 U9201 ( .A1(n9052), .A2(n9051), .ZN(n9252) );
  AND2_X1 U9202 ( .A1(n9049), .A2(n9253), .ZN(n9251) );
  OR2_X1 U9203 ( .A1(n9051), .A2(n9052), .ZN(n9253) );
  OR2_X1 U9204 ( .A1(n8146), .A2(n8802), .ZN(n9052) );
  OR2_X1 U9205 ( .A1(n9254), .A2(n9255), .ZN(n9051) );
  AND2_X1 U9206 ( .A1(n9048), .A2(n9047), .ZN(n9255) );
  AND2_X1 U9207 ( .A1(n9045), .A2(n9256), .ZN(n9254) );
  OR2_X1 U9208 ( .A1(n9047), .A2(n9048), .ZN(n9256) );
  OR2_X1 U9209 ( .A1(n8141), .A2(n8802), .ZN(n9048) );
  OR2_X1 U9210 ( .A1(n9257), .A2(n9258), .ZN(n9047) );
  AND2_X1 U9211 ( .A1(n9044), .A2(n9043), .ZN(n9258) );
  AND2_X1 U9212 ( .A1(n9041), .A2(n9259), .ZN(n9257) );
  OR2_X1 U9213 ( .A1(n9043), .A2(n9044), .ZN(n9259) );
  OR2_X1 U9214 ( .A1(n8136), .A2(n8802), .ZN(n9044) );
  OR2_X1 U9215 ( .A1(n9260), .A2(n9261), .ZN(n9043) );
  AND2_X1 U9216 ( .A1(n9040), .A2(n9039), .ZN(n9261) );
  AND2_X1 U9217 ( .A1(n9037), .A2(n9262), .ZN(n9260) );
  OR2_X1 U9218 ( .A1(n9039), .A2(n9040), .ZN(n9262) );
  OR2_X1 U9219 ( .A1(n8131), .A2(n8802), .ZN(n9040) );
  OR2_X1 U9220 ( .A1(n9263), .A2(n9264), .ZN(n9039) );
  AND2_X1 U9221 ( .A1(n9036), .A2(n9035), .ZN(n9264) );
  AND2_X1 U9222 ( .A1(n9033), .A2(n9265), .ZN(n9263) );
  OR2_X1 U9223 ( .A1(n9035), .A2(n9036), .ZN(n9265) );
  OR2_X1 U9224 ( .A1(n8126), .A2(n8802), .ZN(n9036) );
  OR2_X1 U9225 ( .A1(n9266), .A2(n9267), .ZN(n9035) );
  AND2_X1 U9226 ( .A1(n9030), .A2(n9032), .ZN(n9267) );
  AND2_X1 U9227 ( .A1(n9268), .A2(n9031), .ZN(n9266) );
  OR2_X1 U9228 ( .A1(n9032), .A2(n9030), .ZN(n9268) );
  XOR2_X1 U9229 ( .A(n9269), .B(n9270), .Z(n9030) );
  XOR2_X1 U9230 ( .A(n9271), .B(n9272), .Z(n9270) );
  OR2_X1 U9231 ( .A1(n9273), .A2(n9274), .ZN(n9032) );
  AND2_X1 U9232 ( .A1(n9028), .A2(n9027), .ZN(n9274) );
  AND2_X1 U9233 ( .A1(n9025), .A2(n9275), .ZN(n9273) );
  OR2_X1 U9234 ( .A1(n9027), .A2(n9028), .ZN(n9275) );
  OR2_X1 U9235 ( .A1(n8116), .A2(n8802), .ZN(n9028) );
  OR2_X1 U9236 ( .A1(n9276), .A2(n9277), .ZN(n9027) );
  AND2_X1 U9237 ( .A1(n9006), .A2(n9005), .ZN(n9277) );
  AND2_X1 U9238 ( .A1(n9003), .A2(n9278), .ZN(n9276) );
  OR2_X1 U9239 ( .A1(n9005), .A2(n9006), .ZN(n9278) );
  OR2_X1 U9240 ( .A1(n8111), .A2(n8802), .ZN(n9006) );
  OR2_X1 U9241 ( .A1(n9279), .A2(n9280), .ZN(n9005) );
  AND2_X1 U9242 ( .A1(n9021), .A2(n9024), .ZN(n9280) );
  AND2_X1 U9243 ( .A1(n9023), .A2(n9281), .ZN(n9279) );
  OR2_X1 U9244 ( .A1(n9024), .A2(n9021), .ZN(n9281) );
  OR2_X1 U9245 ( .A1(n8102), .A2(n8802), .ZN(n9021) );
  OR3_X1 U9246 ( .A1(n8349), .A2(n9018), .A3(n8802), .ZN(n9024) );
  INV_X1 U9247 ( .A(n9282), .ZN(n9023) );
  OR2_X1 U9248 ( .A1(n9283), .A2(n9284), .ZN(n9282) );
  AND2_X1 U9249 ( .A1(b_25_), .A2(n9285), .ZN(n9284) );
  OR2_X1 U9250 ( .A1(n9286), .A2(n7314), .ZN(n9285) );
  AND2_X1 U9251 ( .A1(a_30_), .A2(n9145), .ZN(n9286) );
  AND2_X1 U9252 ( .A1(b_24_), .A2(n9287), .ZN(n9283) );
  OR2_X1 U9253 ( .A1(n9288), .A2(n7318), .ZN(n9287) );
  AND2_X1 U9254 ( .A1(a_31_), .A2(n9018), .ZN(n9288) );
  XNOR2_X1 U9255 ( .A(n9289), .B(n9290), .ZN(n9003) );
  XNOR2_X1 U9256 ( .A(n9291), .B(n9292), .ZN(n9290) );
  XOR2_X1 U9257 ( .A(n9293), .B(n9294), .Z(n9025) );
  XOR2_X1 U9258 ( .A(n9295), .B(n9296), .Z(n9294) );
  XOR2_X1 U9259 ( .A(n9297), .B(n9298), .Z(n9033) );
  XOR2_X1 U9260 ( .A(n9299), .B(n9300), .Z(n9298) );
  XNOR2_X1 U9261 ( .A(n9301), .B(n9302), .ZN(n9037) );
  XNOR2_X1 U9262 ( .A(n9303), .B(n9304), .ZN(n9301) );
  XOR2_X1 U9263 ( .A(n9305), .B(n9306), .Z(n9041) );
  XOR2_X1 U9264 ( .A(n9307), .B(n9308), .Z(n9306) );
  XOR2_X1 U9265 ( .A(n9309), .B(n9310), .Z(n9045) );
  XOR2_X1 U9266 ( .A(n9311), .B(n9312), .Z(n9310) );
  XOR2_X1 U9267 ( .A(n9313), .B(n9314), .Z(n9049) );
  XOR2_X1 U9268 ( .A(n9315), .B(n9316), .Z(n9314) );
  XOR2_X1 U9269 ( .A(n9317), .B(n9318), .Z(n9053) );
  XOR2_X1 U9270 ( .A(n9319), .B(n9320), .Z(n9318) );
  XOR2_X1 U9271 ( .A(n9321), .B(n9322), .Z(n9057) );
  XOR2_X1 U9272 ( .A(n9323), .B(n9324), .Z(n9322) );
  XOR2_X1 U9273 ( .A(n9325), .B(n9326), .Z(n9061) );
  XOR2_X1 U9274 ( .A(n9327), .B(n9328), .Z(n9326) );
  XOR2_X1 U9275 ( .A(n9329), .B(n9330), .Z(n9065) );
  XOR2_X1 U9276 ( .A(n9331), .B(n9332), .Z(n9330) );
  XOR2_X1 U9277 ( .A(n9333), .B(n9334), .Z(n9069) );
  XOR2_X1 U9278 ( .A(n9335), .B(n9336), .Z(n9334) );
  XOR2_X1 U9279 ( .A(n9337), .B(n9338), .Z(n9073) );
  XOR2_X1 U9280 ( .A(n9339), .B(n9340), .Z(n9338) );
  XOR2_X1 U9281 ( .A(n9341), .B(n9342), .Z(n9077) );
  XOR2_X1 U9282 ( .A(n9343), .B(n9344), .Z(n9342) );
  XOR2_X1 U9283 ( .A(n9345), .B(n9346), .Z(n9081) );
  XOR2_X1 U9284 ( .A(n9347), .B(n9348), .Z(n9346) );
  XOR2_X1 U9285 ( .A(n9349), .B(n9350), .Z(n9085) );
  XOR2_X1 U9286 ( .A(n9351), .B(n9352), .Z(n9350) );
  XOR2_X1 U9287 ( .A(n9353), .B(n9354), .Z(n9089) );
  XOR2_X1 U9288 ( .A(n9355), .B(n9356), .Z(n9354) );
  XOR2_X1 U9289 ( .A(n9357), .B(n9358), .Z(n9093) );
  XOR2_X1 U9290 ( .A(n9359), .B(n9360), .Z(n9358) );
  XNOR2_X1 U9291 ( .A(n9361), .B(n9362), .ZN(n9097) );
  XNOR2_X1 U9292 ( .A(n9363), .B(n9364), .ZN(n9361) );
  XOR2_X1 U9293 ( .A(n9365), .B(n9366), .Z(n9101) );
  XOR2_X1 U9294 ( .A(n9367), .B(n9368), .Z(n9366) );
  XOR2_X1 U9295 ( .A(n9369), .B(n9370), .Z(n9105) );
  XOR2_X1 U9296 ( .A(n9371), .B(n9372), .Z(n9370) );
  OR2_X1 U9297 ( .A1(n8221), .A2(n8802), .ZN(n9111) );
  XOR2_X1 U9298 ( .A(n9373), .B(n9374), .Z(n9110) );
  XOR2_X1 U9299 ( .A(n9375), .B(n9376), .Z(n9374) );
  XNOR2_X1 U9300 ( .A(n9377), .B(n9378), .ZN(n9113) );
  XNOR2_X1 U9301 ( .A(n9379), .B(n9380), .ZN(n9377) );
  XOR2_X1 U9302 ( .A(n9381), .B(n9382), .Z(n9117) );
  XOR2_X1 U9303 ( .A(n9383), .B(n9384), .Z(n9382) );
  XOR2_X1 U9304 ( .A(n9385), .B(n9386), .Z(n9121) );
  XOR2_X1 U9305 ( .A(n9387), .B(n9388), .Z(n9386) );
  XOR2_X1 U9306 ( .A(n9389), .B(n9390), .Z(n9125) );
  XOR2_X1 U9307 ( .A(n9391), .B(n9392), .Z(n9390) );
  XOR2_X1 U9308 ( .A(n9393), .B(n9394), .Z(n9129) );
  XOR2_X1 U9309 ( .A(n9395), .B(n9396), .Z(n9394) );
  XOR2_X1 U9310 ( .A(n9168), .B(n9397), .Z(n9133) );
  XOR2_X1 U9311 ( .A(n9167), .B(n9166), .Z(n9397) );
  OR2_X1 U9312 ( .A1(n7656), .A2(n9018), .ZN(n9166) );
  OR2_X1 U9313 ( .A1(n9398), .A2(n9399), .ZN(n9167) );
  AND2_X1 U9314 ( .A1(n9396), .A2(n9395), .ZN(n9399) );
  AND2_X1 U9315 ( .A1(n9393), .A2(n9400), .ZN(n9398) );
  OR2_X1 U9316 ( .A1(n9396), .A2(n9395), .ZN(n9400) );
  OR2_X1 U9317 ( .A1(n9401), .A2(n9402), .ZN(n9395) );
  AND2_X1 U9318 ( .A1(n9392), .A2(n9391), .ZN(n9402) );
  AND2_X1 U9319 ( .A1(n9389), .A2(n9403), .ZN(n9401) );
  OR2_X1 U9320 ( .A1(n9392), .A2(n9391), .ZN(n9403) );
  OR2_X1 U9321 ( .A1(n9404), .A2(n9405), .ZN(n9391) );
  AND2_X1 U9322 ( .A1(n9388), .A2(n9387), .ZN(n9405) );
  AND2_X1 U9323 ( .A1(n9385), .A2(n9406), .ZN(n9404) );
  OR2_X1 U9324 ( .A1(n9388), .A2(n9387), .ZN(n9406) );
  OR2_X1 U9325 ( .A1(n9407), .A2(n9408), .ZN(n9387) );
  AND2_X1 U9326 ( .A1(n9384), .A2(n9383), .ZN(n9408) );
  AND2_X1 U9327 ( .A1(n9381), .A2(n9409), .ZN(n9407) );
  OR2_X1 U9328 ( .A1(n9384), .A2(n9383), .ZN(n9409) );
  OR2_X1 U9329 ( .A1(n9410), .A2(n9411), .ZN(n9383) );
  AND2_X1 U9330 ( .A1(n9380), .A2(n9379), .ZN(n9411) );
  AND2_X1 U9331 ( .A1(n9378), .A2(n9412), .ZN(n9410) );
  OR2_X1 U9332 ( .A1(n9380), .A2(n9379), .ZN(n9412) );
  OR2_X1 U9333 ( .A1(n8221), .A2(n9018), .ZN(n9379) );
  OR2_X1 U9334 ( .A1(n9413), .A2(n9414), .ZN(n9380) );
  AND2_X1 U9335 ( .A1(n9376), .A2(n9375), .ZN(n9414) );
  AND2_X1 U9336 ( .A1(n9373), .A2(n9415), .ZN(n9413) );
  OR2_X1 U9337 ( .A1(n9376), .A2(n9375), .ZN(n9415) );
  OR2_X1 U9338 ( .A1(n9416), .A2(n9417), .ZN(n9375) );
  AND2_X1 U9339 ( .A1(n9372), .A2(n9371), .ZN(n9417) );
  AND2_X1 U9340 ( .A1(n9369), .A2(n9418), .ZN(n9416) );
  OR2_X1 U9341 ( .A1(n9372), .A2(n9371), .ZN(n9418) );
  OR2_X1 U9342 ( .A1(n9419), .A2(n9420), .ZN(n9371) );
  AND2_X1 U9343 ( .A1(n9368), .A2(n9367), .ZN(n9420) );
  AND2_X1 U9344 ( .A1(n9365), .A2(n9421), .ZN(n9419) );
  OR2_X1 U9345 ( .A1(n9368), .A2(n9367), .ZN(n9421) );
  OR2_X1 U9346 ( .A1(n9422), .A2(n9423), .ZN(n9367) );
  AND2_X1 U9347 ( .A1(n9364), .A2(n9363), .ZN(n9423) );
  AND2_X1 U9348 ( .A1(n9362), .A2(n9424), .ZN(n9422) );
  OR2_X1 U9349 ( .A1(n9364), .A2(n9363), .ZN(n9424) );
  OR2_X1 U9350 ( .A1(n8201), .A2(n9018), .ZN(n9363) );
  OR2_X1 U9351 ( .A1(n9425), .A2(n9426), .ZN(n9364) );
  AND2_X1 U9352 ( .A1(n9360), .A2(n9359), .ZN(n9426) );
  AND2_X1 U9353 ( .A1(n9357), .A2(n9427), .ZN(n9425) );
  OR2_X1 U9354 ( .A1(n9360), .A2(n9359), .ZN(n9427) );
  OR2_X1 U9355 ( .A1(n9428), .A2(n9429), .ZN(n9359) );
  AND2_X1 U9356 ( .A1(n9356), .A2(n9355), .ZN(n9429) );
  AND2_X1 U9357 ( .A1(n9353), .A2(n9430), .ZN(n9428) );
  OR2_X1 U9358 ( .A1(n9356), .A2(n9355), .ZN(n9430) );
  OR2_X1 U9359 ( .A1(n9431), .A2(n9432), .ZN(n9355) );
  AND2_X1 U9360 ( .A1(n9352), .A2(n9351), .ZN(n9432) );
  AND2_X1 U9361 ( .A1(n9349), .A2(n9433), .ZN(n9431) );
  OR2_X1 U9362 ( .A1(n9352), .A2(n9351), .ZN(n9433) );
  OR2_X1 U9363 ( .A1(n9434), .A2(n9435), .ZN(n9351) );
  AND2_X1 U9364 ( .A1(n9348), .A2(n9347), .ZN(n9435) );
  AND2_X1 U9365 ( .A1(n9345), .A2(n9436), .ZN(n9434) );
  OR2_X1 U9366 ( .A1(n9348), .A2(n9347), .ZN(n9436) );
  OR2_X1 U9367 ( .A1(n9437), .A2(n9438), .ZN(n9347) );
  AND2_X1 U9368 ( .A1(n9344), .A2(n9343), .ZN(n9438) );
  AND2_X1 U9369 ( .A1(n9341), .A2(n9439), .ZN(n9437) );
  OR2_X1 U9370 ( .A1(n9344), .A2(n9343), .ZN(n9439) );
  OR2_X1 U9371 ( .A1(n9440), .A2(n9441), .ZN(n9343) );
  AND2_X1 U9372 ( .A1(n9340), .A2(n9339), .ZN(n9441) );
  AND2_X1 U9373 ( .A1(n9337), .A2(n9442), .ZN(n9440) );
  OR2_X1 U9374 ( .A1(n9340), .A2(n9339), .ZN(n9442) );
  OR2_X1 U9375 ( .A1(n9443), .A2(n9444), .ZN(n9339) );
  AND2_X1 U9376 ( .A1(n9336), .A2(n9335), .ZN(n9444) );
  AND2_X1 U9377 ( .A1(n9333), .A2(n9445), .ZN(n9443) );
  OR2_X1 U9378 ( .A1(n9336), .A2(n9335), .ZN(n9445) );
  OR2_X1 U9379 ( .A1(n9446), .A2(n9447), .ZN(n9335) );
  AND2_X1 U9380 ( .A1(n9332), .A2(n9331), .ZN(n9447) );
  AND2_X1 U9381 ( .A1(n9329), .A2(n9448), .ZN(n9446) );
  OR2_X1 U9382 ( .A1(n9332), .A2(n9331), .ZN(n9448) );
  OR2_X1 U9383 ( .A1(n9449), .A2(n9450), .ZN(n9331) );
  AND2_X1 U9384 ( .A1(n9328), .A2(n9327), .ZN(n9450) );
  AND2_X1 U9385 ( .A1(n9325), .A2(n9451), .ZN(n9449) );
  OR2_X1 U9386 ( .A1(n9328), .A2(n9327), .ZN(n9451) );
  OR2_X1 U9387 ( .A1(n9452), .A2(n9453), .ZN(n9327) );
  AND2_X1 U9388 ( .A1(n9324), .A2(n9323), .ZN(n9453) );
  AND2_X1 U9389 ( .A1(n9321), .A2(n9454), .ZN(n9452) );
  OR2_X1 U9390 ( .A1(n9324), .A2(n9323), .ZN(n9454) );
  OR2_X1 U9391 ( .A1(n9455), .A2(n9456), .ZN(n9323) );
  AND2_X1 U9392 ( .A1(n9320), .A2(n9319), .ZN(n9456) );
  AND2_X1 U9393 ( .A1(n9317), .A2(n9457), .ZN(n9455) );
  OR2_X1 U9394 ( .A1(n9320), .A2(n9319), .ZN(n9457) );
  OR2_X1 U9395 ( .A1(n9458), .A2(n9459), .ZN(n9319) );
  AND2_X1 U9396 ( .A1(n9316), .A2(n9315), .ZN(n9459) );
  AND2_X1 U9397 ( .A1(n9313), .A2(n9460), .ZN(n9458) );
  OR2_X1 U9398 ( .A1(n9316), .A2(n9315), .ZN(n9460) );
  OR2_X1 U9399 ( .A1(n9461), .A2(n9462), .ZN(n9315) );
  AND2_X1 U9400 ( .A1(n9312), .A2(n9311), .ZN(n9462) );
  AND2_X1 U9401 ( .A1(n9309), .A2(n9463), .ZN(n9461) );
  OR2_X1 U9402 ( .A1(n9312), .A2(n9311), .ZN(n9463) );
  OR2_X1 U9403 ( .A1(n9464), .A2(n9465), .ZN(n9311) );
  AND2_X1 U9404 ( .A1(n9308), .A2(n9307), .ZN(n9465) );
  AND2_X1 U9405 ( .A1(n9305), .A2(n9466), .ZN(n9464) );
  OR2_X1 U9406 ( .A1(n9308), .A2(n9307), .ZN(n9466) );
  OR2_X1 U9407 ( .A1(n9467), .A2(n9468), .ZN(n9307) );
  AND2_X1 U9408 ( .A1(n9302), .A2(n9304), .ZN(n9468) );
  AND2_X1 U9409 ( .A1(n9469), .A2(n9303), .ZN(n9467) );
  OR2_X1 U9410 ( .A1(n9302), .A2(n9304), .ZN(n9469) );
  OR2_X1 U9411 ( .A1(n9470), .A2(n9471), .ZN(n9304) );
  AND2_X1 U9412 ( .A1(n9300), .A2(n9299), .ZN(n9471) );
  AND2_X1 U9413 ( .A1(n9297), .A2(n9472), .ZN(n9470) );
  OR2_X1 U9414 ( .A1(n9300), .A2(n9299), .ZN(n9472) );
  OR2_X1 U9415 ( .A1(n9473), .A2(n9474), .ZN(n9299) );
  AND2_X1 U9416 ( .A1(n9272), .A2(n9271), .ZN(n9474) );
  AND2_X1 U9417 ( .A1(n9269), .A2(n9475), .ZN(n9473) );
  OR2_X1 U9418 ( .A1(n9272), .A2(n9271), .ZN(n9475) );
  OR2_X1 U9419 ( .A1(n9476), .A2(n9477), .ZN(n9271) );
  AND2_X1 U9420 ( .A1(n9296), .A2(n9295), .ZN(n9477) );
  AND2_X1 U9421 ( .A1(n9293), .A2(n9478), .ZN(n9476) );
  OR2_X1 U9422 ( .A1(n9296), .A2(n9295), .ZN(n9478) );
  OR2_X1 U9423 ( .A1(n9479), .A2(n9480), .ZN(n9295) );
  AND2_X1 U9424 ( .A1(n9289), .A2(n9292), .ZN(n9480) );
  AND2_X1 U9425 ( .A1(n9291), .A2(n9481), .ZN(n9479) );
  OR2_X1 U9426 ( .A1(n9289), .A2(n9292), .ZN(n9481) );
  OR3_X1 U9427 ( .A1(n8349), .A2(n9145), .A3(n9018), .ZN(n9292) );
  OR2_X1 U9428 ( .A1(n8102), .A2(n9018), .ZN(n9289) );
  INV_X1 U9429 ( .A(n9482), .ZN(n9291) );
  OR2_X1 U9430 ( .A1(n9483), .A2(n9484), .ZN(n9482) );
  AND2_X1 U9431 ( .A1(b_24_), .A2(n9485), .ZN(n9484) );
  OR2_X1 U9432 ( .A1(n9486), .A2(n7314), .ZN(n9485) );
  AND2_X1 U9433 ( .A1(a_30_), .A2(n7976), .ZN(n9486) );
  AND2_X1 U9434 ( .A1(b_23_), .A2(n9487), .ZN(n9483) );
  OR2_X1 U9435 ( .A1(n9488), .A2(n7318), .ZN(n9487) );
  AND2_X1 U9436 ( .A1(a_31_), .A2(n9145), .ZN(n9488) );
  OR2_X1 U9437 ( .A1(n8111), .A2(n9018), .ZN(n9296) );
  XNOR2_X1 U9438 ( .A(n9489), .B(n9490), .ZN(n9293) );
  XNOR2_X1 U9439 ( .A(n9491), .B(n9492), .ZN(n9490) );
  OR2_X1 U9440 ( .A1(n8116), .A2(n9018), .ZN(n9272) );
  XOR2_X1 U9441 ( .A(n9493), .B(n9494), .Z(n9269) );
  XOR2_X1 U9442 ( .A(n9495), .B(n9496), .Z(n9494) );
  OR2_X1 U9443 ( .A1(n8121), .A2(n9018), .ZN(n9300) );
  XOR2_X1 U9444 ( .A(n9497), .B(n9498), .Z(n9297) );
  XOR2_X1 U9445 ( .A(n9499), .B(n9500), .Z(n9498) );
  XOR2_X1 U9446 ( .A(n9501), .B(n9502), .Z(n9302) );
  XOR2_X1 U9447 ( .A(n9503), .B(n9504), .Z(n9502) );
  OR2_X1 U9448 ( .A1(n8131), .A2(n9018), .ZN(n9308) );
  XOR2_X1 U9449 ( .A(n9505), .B(n9506), .Z(n9305) );
  XOR2_X1 U9450 ( .A(n9507), .B(n9508), .Z(n9506) );
  OR2_X1 U9451 ( .A1(n8136), .A2(n9018), .ZN(n9312) );
  XNOR2_X1 U9452 ( .A(n9509), .B(n9510), .ZN(n9309) );
  XNOR2_X1 U9453 ( .A(n9511), .B(n9512), .ZN(n9509) );
  OR2_X1 U9454 ( .A1(n8141), .A2(n9018), .ZN(n9316) );
  XOR2_X1 U9455 ( .A(n9513), .B(n9514), .Z(n9313) );
  XOR2_X1 U9456 ( .A(n9515), .B(n9516), .Z(n9514) );
  OR2_X1 U9457 ( .A1(n8146), .A2(n9018), .ZN(n9320) );
  XOR2_X1 U9458 ( .A(n9517), .B(n9518), .Z(n9317) );
  XOR2_X1 U9459 ( .A(n9519), .B(n9520), .Z(n9518) );
  OR2_X1 U9460 ( .A1(n8151), .A2(n9018), .ZN(n9324) );
  XOR2_X1 U9461 ( .A(n9521), .B(n9522), .Z(n9321) );
  XOR2_X1 U9462 ( .A(n9523), .B(n9524), .Z(n9522) );
  OR2_X1 U9463 ( .A1(n8156), .A2(n9018), .ZN(n9328) );
  XOR2_X1 U9464 ( .A(n9525), .B(n9526), .Z(n9325) );
  XOR2_X1 U9465 ( .A(n9527), .B(n9528), .Z(n9526) );
  OR2_X1 U9466 ( .A1(n8161), .A2(n9018), .ZN(n9332) );
  XOR2_X1 U9467 ( .A(n9529), .B(n9530), .Z(n9329) );
  XOR2_X1 U9468 ( .A(n9531), .B(n9532), .Z(n9530) );
  OR2_X1 U9469 ( .A1(n8166), .A2(n9018), .ZN(n9336) );
  XOR2_X1 U9470 ( .A(n9533), .B(n9534), .Z(n9333) );
  XOR2_X1 U9471 ( .A(n9535), .B(n9536), .Z(n9534) );
  OR2_X1 U9472 ( .A1(n8171), .A2(n9018), .ZN(n9340) );
  XOR2_X1 U9473 ( .A(n9537), .B(n9538), .Z(n9337) );
  XOR2_X1 U9474 ( .A(n9539), .B(n9540), .Z(n9538) );
  OR2_X1 U9475 ( .A1(n8176), .A2(n9018), .ZN(n9344) );
  XOR2_X1 U9476 ( .A(n9541), .B(n9542), .Z(n9341) );
  XOR2_X1 U9477 ( .A(n9543), .B(n9544), .Z(n9542) );
  OR2_X1 U9478 ( .A1(n8181), .A2(n9018), .ZN(n9348) );
  XOR2_X1 U9479 ( .A(n9545), .B(n9546), .Z(n9345) );
  XOR2_X1 U9480 ( .A(n9547), .B(n9548), .Z(n9546) );
  OR2_X1 U9481 ( .A1(n8186), .A2(n9018), .ZN(n9352) );
  XOR2_X1 U9482 ( .A(n9549), .B(n9550), .Z(n9349) );
  XOR2_X1 U9483 ( .A(n9551), .B(n9552), .Z(n9550) );
  OR2_X1 U9484 ( .A1(n8191), .A2(n9018), .ZN(n9356) );
  XOR2_X1 U9485 ( .A(n9553), .B(n9554), .Z(n9353) );
  XOR2_X1 U9486 ( .A(n9555), .B(n9556), .Z(n9554) );
  OR2_X1 U9487 ( .A1(n8196), .A2(n9018), .ZN(n9360) );
  XOR2_X1 U9488 ( .A(n9557), .B(n9558), .Z(n9357) );
  XOR2_X1 U9489 ( .A(n9559), .B(n9560), .Z(n9558) );
  XOR2_X1 U9490 ( .A(n9561), .B(n9562), .Z(n9362) );
  XOR2_X1 U9491 ( .A(n9563), .B(n9564), .Z(n9562) );
  OR2_X1 U9492 ( .A1(n8206), .A2(n9018), .ZN(n9368) );
  XNOR2_X1 U9493 ( .A(n9565), .B(n9566), .ZN(n9365) );
  XNOR2_X1 U9494 ( .A(n9567), .B(n9568), .ZN(n9565) );
  OR2_X1 U9495 ( .A1(n8211), .A2(n9018), .ZN(n9372) );
  XOR2_X1 U9496 ( .A(n9569), .B(n9570), .Z(n9369) );
  XOR2_X1 U9497 ( .A(n9571), .B(n9572), .Z(n9570) );
  OR2_X1 U9498 ( .A1(n8216), .A2(n9018), .ZN(n9376) );
  XOR2_X1 U9499 ( .A(n9573), .B(n9574), .Z(n9373) );
  XOR2_X1 U9500 ( .A(n9575), .B(n9576), .Z(n9574) );
  XOR2_X1 U9501 ( .A(n9577), .B(n9578), .Z(n9378) );
  XOR2_X1 U9502 ( .A(n9579), .B(n9580), .Z(n9578) );
  OR2_X1 U9503 ( .A1(n8226), .A2(n9018), .ZN(n9384) );
  XNOR2_X1 U9504 ( .A(n9581), .B(n9582), .ZN(n9381) );
  XNOR2_X1 U9505 ( .A(n9583), .B(n9584), .ZN(n9581) );
  OR2_X1 U9506 ( .A1(n7785), .A2(n9018), .ZN(n9388) );
  XOR2_X1 U9507 ( .A(n9585), .B(n9586), .Z(n9385) );
  XOR2_X1 U9508 ( .A(n9587), .B(n9588), .Z(n9586) );
  OR2_X1 U9509 ( .A1(n7777), .A2(n9018), .ZN(n9392) );
  XOR2_X1 U9510 ( .A(n9589), .B(n9590), .Z(n9389) );
  XOR2_X1 U9511 ( .A(n9591), .B(n9592), .Z(n9590) );
  OR2_X1 U9512 ( .A1(n7689), .A2(n9018), .ZN(n9396) );
  XNOR2_X1 U9513 ( .A(n9593), .B(n9594), .ZN(n9393) );
  XNOR2_X1 U9514 ( .A(n9595), .B(n9596), .ZN(n9593) );
  XOR2_X1 U9515 ( .A(n9186), .B(n9597), .Z(n9168) );
  XOR2_X1 U9516 ( .A(n9185), .B(n9184), .Z(n9597) );
  OR2_X1 U9517 ( .A1(n7689), .A2(n9145), .ZN(n9184) );
  OR2_X1 U9518 ( .A1(n9598), .A2(n9599), .ZN(n9185) );
  AND2_X1 U9519 ( .A1(n9596), .A2(n9595), .ZN(n9599) );
  AND2_X1 U9520 ( .A1(n9594), .A2(n9600), .ZN(n9598) );
  OR2_X1 U9521 ( .A1(n9596), .A2(n9595), .ZN(n9600) );
  OR2_X1 U9522 ( .A1(n7777), .A2(n9145), .ZN(n9595) );
  OR2_X1 U9523 ( .A1(n9601), .A2(n9602), .ZN(n9596) );
  AND2_X1 U9524 ( .A1(n9592), .A2(n9591), .ZN(n9602) );
  AND2_X1 U9525 ( .A1(n9589), .A2(n9603), .ZN(n9601) );
  OR2_X1 U9526 ( .A1(n9592), .A2(n9591), .ZN(n9603) );
  OR2_X1 U9527 ( .A1(n9604), .A2(n9605), .ZN(n9591) );
  AND2_X1 U9528 ( .A1(n9588), .A2(n9587), .ZN(n9605) );
  AND2_X1 U9529 ( .A1(n9585), .A2(n9606), .ZN(n9604) );
  OR2_X1 U9530 ( .A1(n9588), .A2(n9587), .ZN(n9606) );
  OR2_X1 U9531 ( .A1(n9607), .A2(n9608), .ZN(n9587) );
  AND2_X1 U9532 ( .A1(n9584), .A2(n9583), .ZN(n9608) );
  AND2_X1 U9533 ( .A1(n9582), .A2(n9609), .ZN(n9607) );
  OR2_X1 U9534 ( .A1(n9584), .A2(n9583), .ZN(n9609) );
  OR2_X1 U9535 ( .A1(n8221), .A2(n9145), .ZN(n9583) );
  OR2_X1 U9536 ( .A1(n9610), .A2(n9611), .ZN(n9584) );
  AND2_X1 U9537 ( .A1(n9580), .A2(n9579), .ZN(n9611) );
  AND2_X1 U9538 ( .A1(n9577), .A2(n9612), .ZN(n9610) );
  OR2_X1 U9539 ( .A1(n9580), .A2(n9579), .ZN(n9612) );
  OR2_X1 U9540 ( .A1(n9613), .A2(n9614), .ZN(n9579) );
  AND2_X1 U9541 ( .A1(n9576), .A2(n9575), .ZN(n9614) );
  AND2_X1 U9542 ( .A1(n9573), .A2(n9615), .ZN(n9613) );
  OR2_X1 U9543 ( .A1(n9576), .A2(n9575), .ZN(n9615) );
  OR2_X1 U9544 ( .A1(n9616), .A2(n9617), .ZN(n9575) );
  AND2_X1 U9545 ( .A1(n9572), .A2(n9571), .ZN(n9617) );
  AND2_X1 U9546 ( .A1(n9569), .A2(n9618), .ZN(n9616) );
  OR2_X1 U9547 ( .A1(n9572), .A2(n9571), .ZN(n9618) );
  OR2_X1 U9548 ( .A1(n9619), .A2(n9620), .ZN(n9571) );
  AND2_X1 U9549 ( .A1(n9568), .A2(n9567), .ZN(n9620) );
  AND2_X1 U9550 ( .A1(n9566), .A2(n9621), .ZN(n9619) );
  OR2_X1 U9551 ( .A1(n9568), .A2(n9567), .ZN(n9621) );
  OR2_X1 U9552 ( .A1(n8201), .A2(n9145), .ZN(n9567) );
  OR2_X1 U9553 ( .A1(n9622), .A2(n9623), .ZN(n9568) );
  AND2_X1 U9554 ( .A1(n9564), .A2(n9563), .ZN(n9623) );
  AND2_X1 U9555 ( .A1(n9561), .A2(n9624), .ZN(n9622) );
  OR2_X1 U9556 ( .A1(n9564), .A2(n9563), .ZN(n9624) );
  OR2_X1 U9557 ( .A1(n9625), .A2(n9626), .ZN(n9563) );
  AND2_X1 U9558 ( .A1(n9560), .A2(n9559), .ZN(n9626) );
  AND2_X1 U9559 ( .A1(n9557), .A2(n9627), .ZN(n9625) );
  OR2_X1 U9560 ( .A1(n9560), .A2(n9559), .ZN(n9627) );
  OR2_X1 U9561 ( .A1(n9628), .A2(n9629), .ZN(n9559) );
  AND2_X1 U9562 ( .A1(n9556), .A2(n9555), .ZN(n9629) );
  AND2_X1 U9563 ( .A1(n9553), .A2(n9630), .ZN(n9628) );
  OR2_X1 U9564 ( .A1(n9556), .A2(n9555), .ZN(n9630) );
  OR2_X1 U9565 ( .A1(n9631), .A2(n9632), .ZN(n9555) );
  AND2_X1 U9566 ( .A1(n9552), .A2(n9551), .ZN(n9632) );
  AND2_X1 U9567 ( .A1(n9549), .A2(n9633), .ZN(n9631) );
  OR2_X1 U9568 ( .A1(n9552), .A2(n9551), .ZN(n9633) );
  OR2_X1 U9569 ( .A1(n9634), .A2(n9635), .ZN(n9551) );
  AND2_X1 U9570 ( .A1(n9548), .A2(n9547), .ZN(n9635) );
  AND2_X1 U9571 ( .A1(n9545), .A2(n9636), .ZN(n9634) );
  OR2_X1 U9572 ( .A1(n9548), .A2(n9547), .ZN(n9636) );
  OR2_X1 U9573 ( .A1(n9637), .A2(n9638), .ZN(n9547) );
  AND2_X1 U9574 ( .A1(n9544), .A2(n9543), .ZN(n9638) );
  AND2_X1 U9575 ( .A1(n9541), .A2(n9639), .ZN(n9637) );
  OR2_X1 U9576 ( .A1(n9544), .A2(n9543), .ZN(n9639) );
  OR2_X1 U9577 ( .A1(n9640), .A2(n9641), .ZN(n9543) );
  AND2_X1 U9578 ( .A1(n9540), .A2(n9539), .ZN(n9641) );
  AND2_X1 U9579 ( .A1(n9537), .A2(n9642), .ZN(n9640) );
  OR2_X1 U9580 ( .A1(n9540), .A2(n9539), .ZN(n9642) );
  OR2_X1 U9581 ( .A1(n9643), .A2(n9644), .ZN(n9539) );
  AND2_X1 U9582 ( .A1(n9536), .A2(n9535), .ZN(n9644) );
  AND2_X1 U9583 ( .A1(n9533), .A2(n9645), .ZN(n9643) );
  OR2_X1 U9584 ( .A1(n9536), .A2(n9535), .ZN(n9645) );
  OR2_X1 U9585 ( .A1(n9646), .A2(n9647), .ZN(n9535) );
  AND2_X1 U9586 ( .A1(n9532), .A2(n9531), .ZN(n9647) );
  AND2_X1 U9587 ( .A1(n9529), .A2(n9648), .ZN(n9646) );
  OR2_X1 U9588 ( .A1(n9532), .A2(n9531), .ZN(n9648) );
  OR2_X1 U9589 ( .A1(n9649), .A2(n9650), .ZN(n9531) );
  AND2_X1 U9590 ( .A1(n9528), .A2(n9527), .ZN(n9650) );
  AND2_X1 U9591 ( .A1(n9525), .A2(n9651), .ZN(n9649) );
  OR2_X1 U9592 ( .A1(n9528), .A2(n9527), .ZN(n9651) );
  OR2_X1 U9593 ( .A1(n9652), .A2(n9653), .ZN(n9527) );
  AND2_X1 U9594 ( .A1(n9524), .A2(n9523), .ZN(n9653) );
  AND2_X1 U9595 ( .A1(n9521), .A2(n9654), .ZN(n9652) );
  OR2_X1 U9596 ( .A1(n9524), .A2(n9523), .ZN(n9654) );
  OR2_X1 U9597 ( .A1(n9655), .A2(n9656), .ZN(n9523) );
  AND2_X1 U9598 ( .A1(n9520), .A2(n9519), .ZN(n9656) );
  AND2_X1 U9599 ( .A1(n9517), .A2(n9657), .ZN(n9655) );
  OR2_X1 U9600 ( .A1(n9520), .A2(n9519), .ZN(n9657) );
  OR2_X1 U9601 ( .A1(n9658), .A2(n9659), .ZN(n9519) );
  AND2_X1 U9602 ( .A1(n9516), .A2(n9515), .ZN(n9659) );
  AND2_X1 U9603 ( .A1(n9513), .A2(n9660), .ZN(n9658) );
  OR2_X1 U9604 ( .A1(n9516), .A2(n9515), .ZN(n9660) );
  OR2_X1 U9605 ( .A1(n9661), .A2(n9662), .ZN(n9515) );
  AND2_X1 U9606 ( .A1(n9510), .A2(n9512), .ZN(n9662) );
  AND2_X1 U9607 ( .A1(n9663), .A2(n9511), .ZN(n9661) );
  OR2_X1 U9608 ( .A1(n9510), .A2(n9512), .ZN(n9663) );
  OR2_X1 U9609 ( .A1(n9664), .A2(n9665), .ZN(n9512) );
  AND2_X1 U9610 ( .A1(n9508), .A2(n9507), .ZN(n9665) );
  AND2_X1 U9611 ( .A1(n9505), .A2(n9666), .ZN(n9664) );
  OR2_X1 U9612 ( .A1(n9508), .A2(n9507), .ZN(n9666) );
  OR2_X1 U9613 ( .A1(n9667), .A2(n9668), .ZN(n9507) );
  AND2_X1 U9614 ( .A1(n9504), .A2(n9503), .ZN(n9668) );
  AND2_X1 U9615 ( .A1(n9501), .A2(n9669), .ZN(n9667) );
  OR2_X1 U9616 ( .A1(n9504), .A2(n9503), .ZN(n9669) );
  OR2_X1 U9617 ( .A1(n9670), .A2(n9671), .ZN(n9503) );
  AND2_X1 U9618 ( .A1(n9500), .A2(n9499), .ZN(n9671) );
  AND2_X1 U9619 ( .A1(n9497), .A2(n9672), .ZN(n9670) );
  OR2_X1 U9620 ( .A1(n9500), .A2(n9499), .ZN(n9672) );
  OR2_X1 U9621 ( .A1(n9673), .A2(n9674), .ZN(n9499) );
  AND2_X1 U9622 ( .A1(n9496), .A2(n9495), .ZN(n9674) );
  AND2_X1 U9623 ( .A1(n9493), .A2(n9675), .ZN(n9673) );
  OR2_X1 U9624 ( .A1(n9496), .A2(n9495), .ZN(n9675) );
  OR2_X1 U9625 ( .A1(n9676), .A2(n9677), .ZN(n9495) );
  AND2_X1 U9626 ( .A1(n9489), .A2(n9492), .ZN(n9677) );
  AND2_X1 U9627 ( .A1(n9491), .A2(n9678), .ZN(n9676) );
  OR2_X1 U9628 ( .A1(n9489), .A2(n9492), .ZN(n9678) );
  OR3_X1 U9629 ( .A1(n8349), .A2(n7976), .A3(n9145), .ZN(n9492) );
  OR2_X1 U9630 ( .A1(n8102), .A2(n9145), .ZN(n9489) );
  INV_X1 U9631 ( .A(n9679), .ZN(n9491) );
  OR2_X1 U9632 ( .A1(n9680), .A2(n9681), .ZN(n9679) );
  AND2_X1 U9633 ( .A1(b_23_), .A2(n9682), .ZN(n9681) );
  OR2_X1 U9634 ( .A1(n9683), .A2(n7314), .ZN(n9682) );
  AND2_X1 U9635 ( .A1(a_30_), .A2(n9684), .ZN(n9683) );
  AND2_X1 U9636 ( .A1(b_22_), .A2(n9685), .ZN(n9680) );
  OR2_X1 U9637 ( .A1(n9686), .A2(n7318), .ZN(n9685) );
  AND2_X1 U9638 ( .A1(a_31_), .A2(n7976), .ZN(n9686) );
  OR2_X1 U9639 ( .A1(n8111), .A2(n9145), .ZN(n9496) );
  XNOR2_X1 U9640 ( .A(n9687), .B(n9688), .ZN(n9493) );
  XNOR2_X1 U9641 ( .A(n9689), .B(n9690), .ZN(n9688) );
  OR2_X1 U9642 ( .A1(n8116), .A2(n9145), .ZN(n9500) );
  XOR2_X1 U9643 ( .A(n9691), .B(n9692), .Z(n9497) );
  XOR2_X1 U9644 ( .A(n9693), .B(n9694), .Z(n9692) );
  OR2_X1 U9645 ( .A1(n8121), .A2(n9145), .ZN(n9504) );
  XOR2_X1 U9646 ( .A(n9695), .B(n9696), .Z(n9501) );
  XOR2_X1 U9647 ( .A(n9697), .B(n9698), .Z(n9696) );
  OR2_X1 U9648 ( .A1(n8126), .A2(n9145), .ZN(n9508) );
  XOR2_X1 U9649 ( .A(n9699), .B(n9700), .Z(n9505) );
  XOR2_X1 U9650 ( .A(n9701), .B(n9702), .Z(n9700) );
  XOR2_X1 U9651 ( .A(n9703), .B(n9704), .Z(n9510) );
  XOR2_X1 U9652 ( .A(n9705), .B(n9706), .Z(n9704) );
  OR2_X1 U9653 ( .A1(n8136), .A2(n9145), .ZN(n9516) );
  XOR2_X1 U9654 ( .A(n9707), .B(n9708), .Z(n9513) );
  XOR2_X1 U9655 ( .A(n9709), .B(n9710), .Z(n9708) );
  OR2_X1 U9656 ( .A1(n8141), .A2(n9145), .ZN(n9520) );
  XNOR2_X1 U9657 ( .A(n9711), .B(n9712), .ZN(n9517) );
  XNOR2_X1 U9658 ( .A(n9713), .B(n9714), .ZN(n9711) );
  OR2_X1 U9659 ( .A1(n8146), .A2(n9145), .ZN(n9524) );
  XOR2_X1 U9660 ( .A(n9715), .B(n9716), .Z(n9521) );
  XOR2_X1 U9661 ( .A(n9717), .B(n9718), .Z(n9716) );
  OR2_X1 U9662 ( .A1(n8151), .A2(n9145), .ZN(n9528) );
  XOR2_X1 U9663 ( .A(n9719), .B(n9720), .Z(n9525) );
  XOR2_X1 U9664 ( .A(n9721), .B(n9722), .Z(n9720) );
  OR2_X1 U9665 ( .A1(n8156), .A2(n9145), .ZN(n9532) );
  XOR2_X1 U9666 ( .A(n9723), .B(n9724), .Z(n9529) );
  XOR2_X1 U9667 ( .A(n9725), .B(n9726), .Z(n9724) );
  OR2_X1 U9668 ( .A1(n8161), .A2(n9145), .ZN(n9536) );
  XOR2_X1 U9669 ( .A(n9727), .B(n9728), .Z(n9533) );
  XOR2_X1 U9670 ( .A(n9729), .B(n9730), .Z(n9728) );
  OR2_X1 U9671 ( .A1(n8166), .A2(n9145), .ZN(n9540) );
  XOR2_X1 U9672 ( .A(n9731), .B(n9732), .Z(n9537) );
  XOR2_X1 U9673 ( .A(n9733), .B(n9734), .Z(n9732) );
  OR2_X1 U9674 ( .A1(n8171), .A2(n9145), .ZN(n9544) );
  XOR2_X1 U9675 ( .A(n9735), .B(n9736), .Z(n9541) );
  XOR2_X1 U9676 ( .A(n9737), .B(n9738), .Z(n9736) );
  OR2_X1 U9677 ( .A1(n8176), .A2(n9145), .ZN(n9548) );
  XOR2_X1 U9678 ( .A(n9739), .B(n9740), .Z(n9545) );
  XOR2_X1 U9679 ( .A(n9741), .B(n9742), .Z(n9740) );
  OR2_X1 U9680 ( .A1(n8181), .A2(n9145), .ZN(n9552) );
  XOR2_X1 U9681 ( .A(n9743), .B(n9744), .Z(n9549) );
  XOR2_X1 U9682 ( .A(n9745), .B(n9746), .Z(n9744) );
  OR2_X1 U9683 ( .A1(n8186), .A2(n9145), .ZN(n9556) );
  XNOR2_X1 U9684 ( .A(n9747), .B(n9748), .ZN(n9553) );
  XNOR2_X1 U9685 ( .A(n9749), .B(n9750), .ZN(n9747) );
  OR2_X1 U9686 ( .A1(n8191), .A2(n9145), .ZN(n9560) );
  XOR2_X1 U9687 ( .A(n9751), .B(n9752), .Z(n9557) );
  XOR2_X1 U9688 ( .A(n9753), .B(n9754), .Z(n9752) );
  OR2_X1 U9689 ( .A1(n8196), .A2(n9145), .ZN(n9564) );
  XOR2_X1 U9690 ( .A(n9755), .B(n9756), .Z(n9561) );
  XOR2_X1 U9691 ( .A(n9757), .B(n9758), .Z(n9756) );
  XOR2_X1 U9692 ( .A(n9759), .B(n9760), .Z(n9566) );
  XOR2_X1 U9693 ( .A(n9761), .B(n9762), .Z(n9760) );
  OR2_X1 U9694 ( .A1(n8206), .A2(n9145), .ZN(n9572) );
  XNOR2_X1 U9695 ( .A(n9763), .B(n9764), .ZN(n9569) );
  XNOR2_X1 U9696 ( .A(n9765), .B(n9766), .ZN(n9763) );
  OR2_X1 U9697 ( .A1(n8211), .A2(n9145), .ZN(n9576) );
  XOR2_X1 U9698 ( .A(n9767), .B(n9768), .Z(n9573) );
  XOR2_X1 U9699 ( .A(n9769), .B(n9770), .Z(n9768) );
  OR2_X1 U9700 ( .A1(n8216), .A2(n9145), .ZN(n9580) );
  XOR2_X1 U9701 ( .A(n9771), .B(n9772), .Z(n9577) );
  XOR2_X1 U9702 ( .A(n9773), .B(n9774), .Z(n9772) );
  XOR2_X1 U9703 ( .A(n9775), .B(n9776), .Z(n9582) );
  XOR2_X1 U9704 ( .A(n9777), .B(n9778), .Z(n9776) );
  OR2_X1 U9705 ( .A1(n8226), .A2(n9145), .ZN(n9588) );
  XNOR2_X1 U9706 ( .A(n9779), .B(n9780), .ZN(n9585) );
  XNOR2_X1 U9707 ( .A(n9781), .B(n9782), .ZN(n9779) );
  OR2_X1 U9708 ( .A1(n7785), .A2(n9145), .ZN(n9592) );
  XOR2_X1 U9709 ( .A(n9783), .B(n9784), .Z(n9589) );
  XOR2_X1 U9710 ( .A(n9785), .B(n9786), .Z(n9784) );
  XOR2_X1 U9711 ( .A(n9787), .B(n9788), .Z(n9594) );
  XOR2_X1 U9712 ( .A(n9789), .B(n9790), .Z(n9788) );
  XOR2_X1 U9713 ( .A(n9176), .B(n9791), .Z(n9186) );
  XOR2_X1 U9714 ( .A(n9175), .B(n9174), .Z(n9791) );
  OR2_X1 U9715 ( .A1(n7777), .A2(n7976), .ZN(n9174) );
  OR2_X1 U9716 ( .A1(n9792), .A2(n9793), .ZN(n9175) );
  AND2_X1 U9717 ( .A1(n9790), .A2(n9789), .ZN(n9793) );
  AND2_X1 U9718 ( .A1(n9787), .A2(n9794), .ZN(n9792) );
  OR2_X1 U9719 ( .A1(n9790), .A2(n9789), .ZN(n9794) );
  OR2_X1 U9720 ( .A1(n9795), .A2(n9796), .ZN(n9789) );
  AND2_X1 U9721 ( .A1(n9786), .A2(n9785), .ZN(n9796) );
  AND2_X1 U9722 ( .A1(n9783), .A2(n9797), .ZN(n9795) );
  OR2_X1 U9723 ( .A1(n9786), .A2(n9785), .ZN(n9797) );
  OR2_X1 U9724 ( .A1(n9798), .A2(n9799), .ZN(n9785) );
  AND2_X1 U9725 ( .A1(n9782), .A2(n9781), .ZN(n9799) );
  AND2_X1 U9726 ( .A1(n9780), .A2(n9800), .ZN(n9798) );
  OR2_X1 U9727 ( .A1(n9782), .A2(n9781), .ZN(n9800) );
  OR2_X1 U9728 ( .A1(n8221), .A2(n7976), .ZN(n9781) );
  OR2_X1 U9729 ( .A1(n9801), .A2(n9802), .ZN(n9782) );
  AND2_X1 U9730 ( .A1(n9778), .A2(n9777), .ZN(n9802) );
  AND2_X1 U9731 ( .A1(n9775), .A2(n9803), .ZN(n9801) );
  OR2_X1 U9732 ( .A1(n9778), .A2(n9777), .ZN(n9803) );
  OR2_X1 U9733 ( .A1(n9804), .A2(n9805), .ZN(n9777) );
  AND2_X1 U9734 ( .A1(n9774), .A2(n9773), .ZN(n9805) );
  AND2_X1 U9735 ( .A1(n9771), .A2(n9806), .ZN(n9804) );
  OR2_X1 U9736 ( .A1(n9774), .A2(n9773), .ZN(n9806) );
  OR2_X1 U9737 ( .A1(n9807), .A2(n9808), .ZN(n9773) );
  AND2_X1 U9738 ( .A1(n9770), .A2(n9769), .ZN(n9808) );
  AND2_X1 U9739 ( .A1(n9767), .A2(n9809), .ZN(n9807) );
  OR2_X1 U9740 ( .A1(n9770), .A2(n9769), .ZN(n9809) );
  OR2_X1 U9741 ( .A1(n9810), .A2(n9811), .ZN(n9769) );
  AND2_X1 U9742 ( .A1(n9766), .A2(n9765), .ZN(n9811) );
  AND2_X1 U9743 ( .A1(n9764), .A2(n9812), .ZN(n9810) );
  OR2_X1 U9744 ( .A1(n9766), .A2(n9765), .ZN(n9812) );
  OR2_X1 U9745 ( .A1(n8201), .A2(n7976), .ZN(n9765) );
  OR2_X1 U9746 ( .A1(n9813), .A2(n9814), .ZN(n9766) );
  AND2_X1 U9747 ( .A1(n9762), .A2(n9761), .ZN(n9814) );
  AND2_X1 U9748 ( .A1(n9759), .A2(n9815), .ZN(n9813) );
  OR2_X1 U9749 ( .A1(n9762), .A2(n9761), .ZN(n9815) );
  OR2_X1 U9750 ( .A1(n9816), .A2(n9817), .ZN(n9761) );
  AND2_X1 U9751 ( .A1(n9758), .A2(n9757), .ZN(n9817) );
  AND2_X1 U9752 ( .A1(n9755), .A2(n9818), .ZN(n9816) );
  OR2_X1 U9753 ( .A1(n9758), .A2(n9757), .ZN(n9818) );
  OR2_X1 U9754 ( .A1(n9819), .A2(n9820), .ZN(n9757) );
  AND2_X1 U9755 ( .A1(n9754), .A2(n9753), .ZN(n9820) );
  AND2_X1 U9756 ( .A1(n9751), .A2(n9821), .ZN(n9819) );
  OR2_X1 U9757 ( .A1(n9754), .A2(n9753), .ZN(n9821) );
  OR2_X1 U9758 ( .A1(n9822), .A2(n9823), .ZN(n9753) );
  AND2_X1 U9759 ( .A1(n9750), .A2(n9749), .ZN(n9823) );
  AND2_X1 U9760 ( .A1(n9748), .A2(n9824), .ZN(n9822) );
  OR2_X1 U9761 ( .A1(n9750), .A2(n9749), .ZN(n9824) );
  OR2_X1 U9762 ( .A1(n8181), .A2(n7976), .ZN(n9749) );
  OR2_X1 U9763 ( .A1(n9825), .A2(n9826), .ZN(n9750) );
  AND2_X1 U9764 ( .A1(n9746), .A2(n9745), .ZN(n9826) );
  AND2_X1 U9765 ( .A1(n9743), .A2(n9827), .ZN(n9825) );
  OR2_X1 U9766 ( .A1(n9746), .A2(n9745), .ZN(n9827) );
  OR2_X1 U9767 ( .A1(n9828), .A2(n9829), .ZN(n9745) );
  AND2_X1 U9768 ( .A1(n9742), .A2(n9741), .ZN(n9829) );
  AND2_X1 U9769 ( .A1(n9739), .A2(n9830), .ZN(n9828) );
  OR2_X1 U9770 ( .A1(n9742), .A2(n9741), .ZN(n9830) );
  OR2_X1 U9771 ( .A1(n9831), .A2(n9832), .ZN(n9741) );
  AND2_X1 U9772 ( .A1(n9738), .A2(n9737), .ZN(n9832) );
  AND2_X1 U9773 ( .A1(n9735), .A2(n9833), .ZN(n9831) );
  OR2_X1 U9774 ( .A1(n9738), .A2(n9737), .ZN(n9833) );
  OR2_X1 U9775 ( .A1(n9834), .A2(n9835), .ZN(n9737) );
  AND2_X1 U9776 ( .A1(n9734), .A2(n9733), .ZN(n9835) );
  AND2_X1 U9777 ( .A1(n9731), .A2(n9836), .ZN(n9834) );
  OR2_X1 U9778 ( .A1(n9734), .A2(n9733), .ZN(n9836) );
  OR2_X1 U9779 ( .A1(n9837), .A2(n9838), .ZN(n9733) );
  AND2_X1 U9780 ( .A1(n9730), .A2(n9729), .ZN(n9838) );
  AND2_X1 U9781 ( .A1(n9727), .A2(n9839), .ZN(n9837) );
  OR2_X1 U9782 ( .A1(n9730), .A2(n9729), .ZN(n9839) );
  OR2_X1 U9783 ( .A1(n9840), .A2(n9841), .ZN(n9729) );
  AND2_X1 U9784 ( .A1(n9726), .A2(n9725), .ZN(n9841) );
  AND2_X1 U9785 ( .A1(n9723), .A2(n9842), .ZN(n9840) );
  OR2_X1 U9786 ( .A1(n9726), .A2(n9725), .ZN(n9842) );
  OR2_X1 U9787 ( .A1(n9843), .A2(n9844), .ZN(n9725) );
  AND2_X1 U9788 ( .A1(n9722), .A2(n9721), .ZN(n9844) );
  AND2_X1 U9789 ( .A1(n9719), .A2(n9845), .ZN(n9843) );
  OR2_X1 U9790 ( .A1(n9722), .A2(n9721), .ZN(n9845) );
  OR2_X1 U9791 ( .A1(n9846), .A2(n9847), .ZN(n9721) );
  AND2_X1 U9792 ( .A1(n9718), .A2(n9717), .ZN(n9847) );
  AND2_X1 U9793 ( .A1(n9715), .A2(n9848), .ZN(n9846) );
  OR2_X1 U9794 ( .A1(n9718), .A2(n9717), .ZN(n9848) );
  OR2_X1 U9795 ( .A1(n9849), .A2(n9850), .ZN(n9717) );
  AND2_X1 U9796 ( .A1(n9712), .A2(n9714), .ZN(n9850) );
  AND2_X1 U9797 ( .A1(n9851), .A2(n9713), .ZN(n9849) );
  OR2_X1 U9798 ( .A1(n9712), .A2(n9714), .ZN(n9851) );
  OR2_X1 U9799 ( .A1(n9852), .A2(n9853), .ZN(n9714) );
  AND2_X1 U9800 ( .A1(n9710), .A2(n9709), .ZN(n9853) );
  AND2_X1 U9801 ( .A1(n9707), .A2(n9854), .ZN(n9852) );
  OR2_X1 U9802 ( .A1(n9710), .A2(n9709), .ZN(n9854) );
  OR2_X1 U9803 ( .A1(n9855), .A2(n9856), .ZN(n9709) );
  AND2_X1 U9804 ( .A1(n9706), .A2(n9705), .ZN(n9856) );
  AND2_X1 U9805 ( .A1(n9703), .A2(n9857), .ZN(n9855) );
  OR2_X1 U9806 ( .A1(n9706), .A2(n9705), .ZN(n9857) );
  OR2_X1 U9807 ( .A1(n9858), .A2(n9859), .ZN(n9705) );
  AND2_X1 U9808 ( .A1(n9702), .A2(n9701), .ZN(n9859) );
  AND2_X1 U9809 ( .A1(n9699), .A2(n9860), .ZN(n9858) );
  OR2_X1 U9810 ( .A1(n9702), .A2(n9701), .ZN(n9860) );
  OR2_X1 U9811 ( .A1(n9861), .A2(n9862), .ZN(n9701) );
  AND2_X1 U9812 ( .A1(n9698), .A2(n9697), .ZN(n9862) );
  AND2_X1 U9813 ( .A1(n9695), .A2(n9863), .ZN(n9861) );
  OR2_X1 U9814 ( .A1(n9698), .A2(n9697), .ZN(n9863) );
  OR2_X1 U9815 ( .A1(n9864), .A2(n9865), .ZN(n9697) );
  AND2_X1 U9816 ( .A1(n9694), .A2(n9693), .ZN(n9865) );
  AND2_X1 U9817 ( .A1(n9691), .A2(n9866), .ZN(n9864) );
  OR2_X1 U9818 ( .A1(n9694), .A2(n9693), .ZN(n9866) );
  OR2_X1 U9819 ( .A1(n9867), .A2(n9868), .ZN(n9693) );
  AND2_X1 U9820 ( .A1(n9687), .A2(n9690), .ZN(n9868) );
  AND2_X1 U9821 ( .A1(n9689), .A2(n9869), .ZN(n9867) );
  OR2_X1 U9822 ( .A1(n9687), .A2(n9690), .ZN(n9869) );
  OR3_X1 U9823 ( .A1(n8349), .A2(n7976), .A3(n9684), .ZN(n9690) );
  OR2_X1 U9824 ( .A1(n8102), .A2(n7976), .ZN(n9687) );
  INV_X1 U9825 ( .A(n9870), .ZN(n9689) );
  OR2_X1 U9826 ( .A1(n9871), .A2(n9872), .ZN(n9870) );
  AND2_X1 U9827 ( .A1(b_22_), .A2(n9873), .ZN(n9872) );
  OR2_X1 U9828 ( .A1(n9874), .A2(n7314), .ZN(n9873) );
  AND2_X1 U9829 ( .A1(a_30_), .A2(n9875), .ZN(n9874) );
  AND2_X1 U9830 ( .A1(b_21_), .A2(n9876), .ZN(n9871) );
  OR2_X1 U9831 ( .A1(n9877), .A2(n7318), .ZN(n9876) );
  AND2_X1 U9832 ( .A1(a_31_), .A2(n9684), .ZN(n9877) );
  OR2_X1 U9833 ( .A1(n8111), .A2(n7976), .ZN(n9694) );
  XNOR2_X1 U9834 ( .A(n9878), .B(n9879), .ZN(n9691) );
  XNOR2_X1 U9835 ( .A(n9880), .B(n9881), .ZN(n9879) );
  OR2_X1 U9836 ( .A1(n8116), .A2(n7976), .ZN(n9698) );
  XOR2_X1 U9837 ( .A(n9882), .B(n9883), .Z(n9695) );
  XOR2_X1 U9838 ( .A(n9884), .B(n9885), .Z(n9883) );
  OR2_X1 U9839 ( .A1(n8121), .A2(n7976), .ZN(n9702) );
  XOR2_X1 U9840 ( .A(n9886), .B(n9887), .Z(n9699) );
  XOR2_X1 U9841 ( .A(n9888), .B(n9889), .Z(n9887) );
  OR2_X1 U9842 ( .A1(n8126), .A2(n7976), .ZN(n9706) );
  XOR2_X1 U9843 ( .A(n9890), .B(n9891), .Z(n9703) );
  XOR2_X1 U9844 ( .A(n9892), .B(n9893), .Z(n9891) );
  OR2_X1 U9845 ( .A1(n8131), .A2(n7976), .ZN(n9710) );
  XOR2_X1 U9846 ( .A(n9894), .B(n9895), .Z(n9707) );
  XOR2_X1 U9847 ( .A(n9896), .B(n9897), .Z(n9895) );
  XOR2_X1 U9848 ( .A(n9898), .B(n9899), .Z(n9712) );
  XOR2_X1 U9849 ( .A(n9900), .B(n9901), .Z(n9899) );
  OR2_X1 U9850 ( .A1(n8141), .A2(n7976), .ZN(n9718) );
  XOR2_X1 U9851 ( .A(n9902), .B(n9903), .Z(n9715) );
  XOR2_X1 U9852 ( .A(n9904), .B(n9905), .Z(n9903) );
  OR2_X1 U9853 ( .A1(n8146), .A2(n7976), .ZN(n9722) );
  XNOR2_X1 U9854 ( .A(n9906), .B(n9907), .ZN(n9719) );
  XNOR2_X1 U9855 ( .A(n9908), .B(n9909), .ZN(n9906) );
  OR2_X1 U9856 ( .A1(n8151), .A2(n7976), .ZN(n9726) );
  XOR2_X1 U9857 ( .A(n9910), .B(n9911), .Z(n9723) );
  XOR2_X1 U9858 ( .A(n9912), .B(n9913), .Z(n9911) );
  OR2_X1 U9859 ( .A1(n8156), .A2(n7976), .ZN(n9730) );
  XOR2_X1 U9860 ( .A(n9914), .B(n9915), .Z(n9727) );
  XOR2_X1 U9861 ( .A(n9916), .B(n9917), .Z(n9915) );
  OR2_X1 U9862 ( .A1(n8161), .A2(n7976), .ZN(n9734) );
  XOR2_X1 U9863 ( .A(n9918), .B(n9919), .Z(n9731) );
  XOR2_X1 U9864 ( .A(n9920), .B(n9921), .Z(n9919) );
  OR2_X1 U9865 ( .A1(n8166), .A2(n7976), .ZN(n9738) );
  XOR2_X1 U9866 ( .A(n9922), .B(n9923), .Z(n9735) );
  XOR2_X1 U9867 ( .A(n9924), .B(n9925), .Z(n9923) );
  OR2_X1 U9868 ( .A1(n8171), .A2(n7976), .ZN(n9742) );
  XOR2_X1 U9869 ( .A(n9926), .B(n9927), .Z(n9739) );
  XOR2_X1 U9870 ( .A(n9928), .B(n9929), .Z(n9927) );
  OR2_X1 U9871 ( .A1(n8176), .A2(n7976), .ZN(n9746) );
  XOR2_X1 U9872 ( .A(n9930), .B(n9931), .Z(n9743) );
  XOR2_X1 U9873 ( .A(n9932), .B(n9933), .Z(n9931) );
  XOR2_X1 U9874 ( .A(n9934), .B(n9935), .Z(n9748) );
  XOR2_X1 U9875 ( .A(n9936), .B(n9937), .Z(n9935) );
  OR2_X1 U9876 ( .A1(n8186), .A2(n7976), .ZN(n9754) );
  XOR2_X1 U9877 ( .A(n9938), .B(n9939), .Z(n9751) );
  XOR2_X1 U9878 ( .A(n9940), .B(n9941), .Z(n9939) );
  OR2_X1 U9879 ( .A1(n8191), .A2(n7976), .ZN(n9758) );
  XOR2_X1 U9880 ( .A(n9942), .B(n9943), .Z(n9755) );
  XOR2_X1 U9881 ( .A(n9944), .B(n9945), .Z(n9943) );
  OR2_X1 U9882 ( .A1(n8196), .A2(n7976), .ZN(n9762) );
  XOR2_X1 U9883 ( .A(n9946), .B(n9947), .Z(n9759) );
  XOR2_X1 U9884 ( .A(n9948), .B(n9949), .Z(n9947) );
  XOR2_X1 U9885 ( .A(n9950), .B(n9951), .Z(n9764) );
  XOR2_X1 U9886 ( .A(n9952), .B(n9953), .Z(n9951) );
  OR2_X1 U9887 ( .A1(n8206), .A2(n7976), .ZN(n9770) );
  XOR2_X1 U9888 ( .A(n9954), .B(n9955), .Z(n9767) );
  XOR2_X1 U9889 ( .A(n9956), .B(n9957), .Z(n9955) );
  OR2_X1 U9890 ( .A1(n8211), .A2(n7976), .ZN(n9774) );
  XOR2_X1 U9891 ( .A(n9958), .B(n9959), .Z(n9771) );
  XOR2_X1 U9892 ( .A(n9960), .B(n9961), .Z(n9959) );
  OR2_X1 U9893 ( .A1(n8216), .A2(n7976), .ZN(n9778) );
  XOR2_X1 U9894 ( .A(n9962), .B(n9963), .Z(n9775) );
  XOR2_X1 U9895 ( .A(n9964), .B(n9965), .Z(n9963) );
  XOR2_X1 U9896 ( .A(n9966), .B(n9967), .Z(n9780) );
  XOR2_X1 U9897 ( .A(n9968), .B(n9969), .Z(n9967) );
  OR2_X1 U9898 ( .A1(n8226), .A2(n7976), .ZN(n9786) );
  XOR2_X1 U9899 ( .A(n9970), .B(n9971), .Z(n9783) );
  XOR2_X1 U9900 ( .A(n9972), .B(n9973), .Z(n9971) );
  OR2_X1 U9901 ( .A1(n7785), .A2(n7976), .ZN(n9790) );
  XOR2_X1 U9902 ( .A(n9974), .B(n9975), .Z(n9787) );
  XOR2_X1 U9903 ( .A(n9976), .B(n9977), .Z(n9975) );
  XOR2_X1 U9904 ( .A(n9978), .B(n9979), .Z(n9176) );
  XOR2_X1 U9905 ( .A(n9980), .B(n9981), .Z(n9979) );
  OR2_X1 U9906 ( .A1(n9982), .A2(n7936), .ZN(n7508) );
  XOR2_X1 U9907 ( .A(n7897), .B(n7899), .Z(n7936) );
  OR2_X1 U9908 ( .A1(n9983), .A2(n9984), .ZN(n7899) );
  AND2_X1 U9909 ( .A1(n9985), .A2(n9986), .ZN(n9984) );
  AND2_X1 U9910 ( .A1(n9987), .A2(n9988), .ZN(n9983) );
  OR2_X1 U9911 ( .A1(n9985), .A2(n9986), .ZN(n9988) );
  XOR2_X1 U9912 ( .A(n7906), .B(n9989), .Z(n7897) );
  XOR2_X1 U9913 ( .A(n7905), .B(n7904), .Z(n9989) );
  OR2_X1 U9914 ( .A1(n7621), .A2(n9990), .ZN(n7904) );
  OR2_X1 U9915 ( .A1(n9991), .A2(n9992), .ZN(n7905) );
  AND2_X1 U9916 ( .A1(n9993), .A2(n9994), .ZN(n9992) );
  AND2_X1 U9917 ( .A1(n9995), .A2(n9996), .ZN(n9991) );
  OR2_X1 U9918 ( .A1(n9993), .A2(n9994), .ZN(n9996) );
  XOR2_X1 U9919 ( .A(n7914), .B(n9997), .Z(n7906) );
  XOR2_X1 U9920 ( .A(n7913), .B(n7912), .Z(n9997) );
  OR2_X1 U9921 ( .A1(n7656), .A2(n7909), .ZN(n7912) );
  OR2_X1 U9922 ( .A1(n9998), .A2(n9999), .ZN(n7913) );
  AND2_X1 U9923 ( .A1(n10000), .A2(n10001), .ZN(n9999) );
  AND2_X1 U9924 ( .A1(n10002), .A2(n10003), .ZN(n9998) );
  OR2_X1 U9925 ( .A1(n10000), .A2(n10001), .ZN(n10003) );
  XOR2_X1 U9926 ( .A(n7921), .B(n10004), .Z(n7914) );
  XOR2_X1 U9927 ( .A(n7920), .B(n7919), .Z(n10004) );
  OR2_X1 U9928 ( .A1(n7689), .A2(n7877), .ZN(n7919) );
  OR2_X1 U9929 ( .A1(n10005), .A2(n10006), .ZN(n7920) );
  AND2_X1 U9930 ( .A1(n10007), .A2(n10008), .ZN(n10006) );
  AND2_X1 U9931 ( .A1(n10009), .A2(n10010), .ZN(n10005) );
  OR2_X1 U9932 ( .A1(n10007), .A2(n10008), .ZN(n10010) );
  XOR2_X1 U9933 ( .A(n7928), .B(n10011), .Z(n7921) );
  XOR2_X1 U9934 ( .A(n7927), .B(n7926), .Z(n10011) );
  OR2_X1 U9935 ( .A1(n7852), .A2(n7777), .ZN(n7926) );
  OR2_X1 U9936 ( .A1(n10012), .A2(n10013), .ZN(n7927) );
  AND2_X1 U9937 ( .A1(n10014), .A2(n10015), .ZN(n10013) );
  AND2_X1 U9938 ( .A1(n10016), .A2(n10017), .ZN(n10012) );
  OR2_X1 U9939 ( .A1(n10014), .A2(n10015), .ZN(n10017) );
  XOR2_X1 U9940 ( .A(n10018), .B(n10019), .Z(n7928) );
  XOR2_X1 U9941 ( .A(n10020), .B(n10021), .Z(n10019) );
  AND2_X1 U9942 ( .A1(n7937), .A2(n7935), .ZN(n9982) );
  XNOR2_X1 U9943 ( .A(n9987), .B(n10022), .ZN(n7935) );
  XOR2_X1 U9944 ( .A(n9986), .B(n9985), .Z(n10022) );
  OR2_X1 U9945 ( .A1(n7621), .A2(n9875), .ZN(n9985) );
  OR2_X1 U9946 ( .A1(n10023), .A2(n10024), .ZN(n9986) );
  AND2_X1 U9947 ( .A1(n10025), .A2(n10026), .ZN(n10024) );
  AND2_X1 U9948 ( .A1(n10027), .A2(n10028), .ZN(n10023) );
  OR2_X1 U9949 ( .A1(n10025), .A2(n10026), .ZN(n10028) );
  XOR2_X1 U9950 ( .A(n9995), .B(n10029), .Z(n9987) );
  XOR2_X1 U9951 ( .A(n9994), .B(n9993), .Z(n10029) );
  OR2_X1 U9952 ( .A1(n7656), .A2(n9990), .ZN(n9993) );
  OR2_X1 U9953 ( .A1(n10030), .A2(n10031), .ZN(n9994) );
  AND2_X1 U9954 ( .A1(n10032), .A2(n10033), .ZN(n10031) );
  AND2_X1 U9955 ( .A1(n10034), .A2(n10035), .ZN(n10030) );
  OR2_X1 U9956 ( .A1(n10032), .A2(n10033), .ZN(n10035) );
  XOR2_X1 U9957 ( .A(n10002), .B(n10036), .Z(n9995) );
  XOR2_X1 U9958 ( .A(n10001), .B(n10000), .Z(n10036) );
  OR2_X1 U9959 ( .A1(n7689), .A2(n7909), .ZN(n10000) );
  OR2_X1 U9960 ( .A1(n10037), .A2(n10038), .ZN(n10001) );
  AND2_X1 U9961 ( .A1(n10039), .A2(n10040), .ZN(n10038) );
  AND2_X1 U9962 ( .A1(n10041), .A2(n10042), .ZN(n10037) );
  OR2_X1 U9963 ( .A1(n10039), .A2(n10040), .ZN(n10042) );
  XOR2_X1 U9964 ( .A(n10009), .B(n10043), .Z(n10002) );
  XOR2_X1 U9965 ( .A(n10008), .B(n10007), .Z(n10043) );
  OR2_X1 U9966 ( .A1(n7777), .A2(n7877), .ZN(n10007) );
  OR2_X1 U9967 ( .A1(n10044), .A2(n10045), .ZN(n10008) );
  AND2_X1 U9968 ( .A1(n10046), .A2(n10047), .ZN(n10045) );
  AND2_X1 U9969 ( .A1(n10048), .A2(n10049), .ZN(n10044) );
  OR2_X1 U9970 ( .A1(n10046), .A2(n10047), .ZN(n10049) );
  XOR2_X1 U9971 ( .A(n10016), .B(n10050), .Z(n10009) );
  XOR2_X1 U9972 ( .A(n10015), .B(n10014), .Z(n10050) );
  OR2_X1 U9973 ( .A1(n7852), .A2(n7785), .ZN(n10014) );
  OR2_X1 U9974 ( .A1(n10051), .A2(n10052), .ZN(n10015) );
  AND2_X1 U9975 ( .A1(n10053), .A2(n10054), .ZN(n10052) );
  AND2_X1 U9976 ( .A1(n10055), .A2(n10056), .ZN(n10051) );
  OR2_X1 U9977 ( .A1(n10053), .A2(n10054), .ZN(n10056) );
  XOR2_X1 U9978 ( .A(n10057), .B(n10058), .Z(n10016) );
  XOR2_X1 U9979 ( .A(n10059), .B(n10060), .Z(n10058) );
  INV_X1 U9980 ( .A(n10061), .ZN(n7937) );
  OR2_X1 U9981 ( .A1(n10062), .A2(n10063), .ZN(n10061) );
  AND2_X1 U9982 ( .A1(n7961), .A2(n7960), .ZN(n10063) );
  AND2_X1 U9983 ( .A1(n7958), .A2(n10064), .ZN(n10062) );
  OR2_X1 U9984 ( .A1(n7960), .A2(n7961), .ZN(n10064) );
  OR2_X1 U9985 ( .A1(n7621), .A2(n9684), .ZN(n7961) );
  OR2_X1 U9986 ( .A1(n10065), .A2(n10066), .ZN(n7960) );
  AND2_X1 U9987 ( .A1(n7986), .A2(n7985), .ZN(n10066) );
  AND2_X1 U9988 ( .A1(n7983), .A2(n10067), .ZN(n10065) );
  OR2_X1 U9989 ( .A1(n7985), .A2(n7986), .ZN(n10067) );
  OR2_X1 U9990 ( .A1(n7656), .A2(n9684), .ZN(n7986) );
  OR2_X1 U9991 ( .A1(n10068), .A2(n10069), .ZN(n7985) );
  AND2_X1 U9992 ( .A1(n9162), .A2(n9161), .ZN(n10069) );
  AND2_X1 U9993 ( .A1(n9159), .A2(n10070), .ZN(n10068) );
  OR2_X1 U9994 ( .A1(n9161), .A2(n9162), .ZN(n10070) );
  OR2_X1 U9995 ( .A1(n7689), .A2(n9684), .ZN(n9162) );
  OR2_X1 U9996 ( .A1(n10071), .A2(n10072), .ZN(n9161) );
  AND2_X1 U9997 ( .A1(n9181), .A2(n9180), .ZN(n10072) );
  AND2_X1 U9998 ( .A1(n9178), .A2(n10073), .ZN(n10071) );
  OR2_X1 U9999 ( .A1(n9180), .A2(n9181), .ZN(n10073) );
  OR2_X1 U10000 ( .A1(n7777), .A2(n9684), .ZN(n9181) );
  OR2_X1 U10001 ( .A1(n10074), .A2(n10075), .ZN(n9180) );
  AND2_X1 U10002 ( .A1(n9981), .A2(n9980), .ZN(n10075) );
  AND2_X1 U10003 ( .A1(n9978), .A2(n10076), .ZN(n10074) );
  OR2_X1 U10004 ( .A1(n9980), .A2(n9981), .ZN(n10076) );
  OR2_X1 U10005 ( .A1(n7785), .A2(n9684), .ZN(n9981) );
  OR2_X1 U10006 ( .A1(n10077), .A2(n10078), .ZN(n9980) );
  AND2_X1 U10007 ( .A1(n9977), .A2(n9976), .ZN(n10078) );
  AND2_X1 U10008 ( .A1(n9974), .A2(n10079), .ZN(n10077) );
  OR2_X1 U10009 ( .A1(n9976), .A2(n9977), .ZN(n10079) );
  OR2_X1 U10010 ( .A1(n8226), .A2(n9684), .ZN(n9977) );
  OR2_X1 U10011 ( .A1(n10080), .A2(n10081), .ZN(n9976) );
  AND2_X1 U10012 ( .A1(n9973), .A2(n9972), .ZN(n10081) );
  AND2_X1 U10013 ( .A1(n9970), .A2(n10082), .ZN(n10080) );
  OR2_X1 U10014 ( .A1(n9972), .A2(n9973), .ZN(n10082) );
  OR2_X1 U10015 ( .A1(n8221), .A2(n9684), .ZN(n9973) );
  OR2_X1 U10016 ( .A1(n10083), .A2(n10084), .ZN(n9972) );
  AND2_X1 U10017 ( .A1(n9969), .A2(n9968), .ZN(n10084) );
  AND2_X1 U10018 ( .A1(n9966), .A2(n10085), .ZN(n10083) );
  OR2_X1 U10019 ( .A1(n9968), .A2(n9969), .ZN(n10085) );
  OR2_X1 U10020 ( .A1(n8216), .A2(n9684), .ZN(n9969) );
  OR2_X1 U10021 ( .A1(n10086), .A2(n10087), .ZN(n9968) );
  AND2_X1 U10022 ( .A1(n9965), .A2(n9964), .ZN(n10087) );
  AND2_X1 U10023 ( .A1(n9962), .A2(n10088), .ZN(n10086) );
  OR2_X1 U10024 ( .A1(n9964), .A2(n9965), .ZN(n10088) );
  OR2_X1 U10025 ( .A1(n8211), .A2(n9684), .ZN(n9965) );
  OR2_X1 U10026 ( .A1(n10089), .A2(n10090), .ZN(n9964) );
  AND2_X1 U10027 ( .A1(n9961), .A2(n9960), .ZN(n10090) );
  AND2_X1 U10028 ( .A1(n9958), .A2(n10091), .ZN(n10089) );
  OR2_X1 U10029 ( .A1(n9960), .A2(n9961), .ZN(n10091) );
  OR2_X1 U10030 ( .A1(n8206), .A2(n9684), .ZN(n9961) );
  OR2_X1 U10031 ( .A1(n10092), .A2(n10093), .ZN(n9960) );
  AND2_X1 U10032 ( .A1(n9957), .A2(n9956), .ZN(n10093) );
  AND2_X1 U10033 ( .A1(n9954), .A2(n10094), .ZN(n10092) );
  OR2_X1 U10034 ( .A1(n9956), .A2(n9957), .ZN(n10094) );
  OR2_X1 U10035 ( .A1(n8201), .A2(n9684), .ZN(n9957) );
  OR2_X1 U10036 ( .A1(n10095), .A2(n10096), .ZN(n9956) );
  AND2_X1 U10037 ( .A1(n9953), .A2(n9952), .ZN(n10096) );
  AND2_X1 U10038 ( .A1(n9950), .A2(n10097), .ZN(n10095) );
  OR2_X1 U10039 ( .A1(n9952), .A2(n9953), .ZN(n10097) );
  OR2_X1 U10040 ( .A1(n8196), .A2(n9684), .ZN(n9953) );
  OR2_X1 U10041 ( .A1(n10098), .A2(n10099), .ZN(n9952) );
  AND2_X1 U10042 ( .A1(n9949), .A2(n9948), .ZN(n10099) );
  AND2_X1 U10043 ( .A1(n9946), .A2(n10100), .ZN(n10098) );
  OR2_X1 U10044 ( .A1(n9948), .A2(n9949), .ZN(n10100) );
  OR2_X1 U10045 ( .A1(n8191), .A2(n9684), .ZN(n9949) );
  OR2_X1 U10046 ( .A1(n10101), .A2(n10102), .ZN(n9948) );
  AND2_X1 U10047 ( .A1(n9945), .A2(n9944), .ZN(n10102) );
  AND2_X1 U10048 ( .A1(n9942), .A2(n10103), .ZN(n10101) );
  OR2_X1 U10049 ( .A1(n9944), .A2(n9945), .ZN(n10103) );
  OR2_X1 U10050 ( .A1(n8186), .A2(n9684), .ZN(n9945) );
  OR2_X1 U10051 ( .A1(n10104), .A2(n10105), .ZN(n9944) );
  AND2_X1 U10052 ( .A1(n9941), .A2(n9940), .ZN(n10105) );
  AND2_X1 U10053 ( .A1(n9938), .A2(n10106), .ZN(n10104) );
  OR2_X1 U10054 ( .A1(n9940), .A2(n9941), .ZN(n10106) );
  OR2_X1 U10055 ( .A1(n8181), .A2(n9684), .ZN(n9941) );
  OR2_X1 U10056 ( .A1(n10107), .A2(n10108), .ZN(n9940) );
  AND2_X1 U10057 ( .A1(n9937), .A2(n9936), .ZN(n10108) );
  AND2_X1 U10058 ( .A1(n9934), .A2(n10109), .ZN(n10107) );
  OR2_X1 U10059 ( .A1(n9936), .A2(n9937), .ZN(n10109) );
  OR2_X1 U10060 ( .A1(n8176), .A2(n9684), .ZN(n9937) );
  OR2_X1 U10061 ( .A1(n10110), .A2(n10111), .ZN(n9936) );
  AND2_X1 U10062 ( .A1(n9933), .A2(n9932), .ZN(n10111) );
  AND2_X1 U10063 ( .A1(n9930), .A2(n10112), .ZN(n10110) );
  OR2_X1 U10064 ( .A1(n9932), .A2(n9933), .ZN(n10112) );
  OR2_X1 U10065 ( .A1(n8171), .A2(n9684), .ZN(n9933) );
  OR2_X1 U10066 ( .A1(n10113), .A2(n10114), .ZN(n9932) );
  AND2_X1 U10067 ( .A1(n9929), .A2(n9928), .ZN(n10114) );
  AND2_X1 U10068 ( .A1(n9926), .A2(n10115), .ZN(n10113) );
  OR2_X1 U10069 ( .A1(n9928), .A2(n9929), .ZN(n10115) );
  OR2_X1 U10070 ( .A1(n8166), .A2(n9684), .ZN(n9929) );
  OR2_X1 U10071 ( .A1(n10116), .A2(n10117), .ZN(n9928) );
  AND2_X1 U10072 ( .A1(n9925), .A2(n9924), .ZN(n10117) );
  AND2_X1 U10073 ( .A1(n9922), .A2(n10118), .ZN(n10116) );
  OR2_X1 U10074 ( .A1(n9924), .A2(n9925), .ZN(n10118) );
  OR2_X1 U10075 ( .A1(n8161), .A2(n9684), .ZN(n9925) );
  OR2_X1 U10076 ( .A1(n10119), .A2(n10120), .ZN(n9924) );
  AND2_X1 U10077 ( .A1(n9921), .A2(n9920), .ZN(n10120) );
  AND2_X1 U10078 ( .A1(n9918), .A2(n10121), .ZN(n10119) );
  OR2_X1 U10079 ( .A1(n9920), .A2(n9921), .ZN(n10121) );
  OR2_X1 U10080 ( .A1(n8156), .A2(n9684), .ZN(n9921) );
  OR2_X1 U10081 ( .A1(n10122), .A2(n10123), .ZN(n9920) );
  AND2_X1 U10082 ( .A1(n9917), .A2(n9916), .ZN(n10123) );
  AND2_X1 U10083 ( .A1(n9914), .A2(n10124), .ZN(n10122) );
  OR2_X1 U10084 ( .A1(n9916), .A2(n9917), .ZN(n10124) );
  OR2_X1 U10085 ( .A1(n8151), .A2(n9684), .ZN(n9917) );
  OR2_X1 U10086 ( .A1(n10125), .A2(n10126), .ZN(n9916) );
  AND2_X1 U10087 ( .A1(n9913), .A2(n9912), .ZN(n10126) );
  AND2_X1 U10088 ( .A1(n9910), .A2(n10127), .ZN(n10125) );
  OR2_X1 U10089 ( .A1(n9912), .A2(n9913), .ZN(n10127) );
  OR2_X1 U10090 ( .A1(n8146), .A2(n9684), .ZN(n9913) );
  OR2_X1 U10091 ( .A1(n10128), .A2(n10129), .ZN(n9912) );
  AND2_X1 U10092 ( .A1(n9907), .A2(n9909), .ZN(n10129) );
  AND2_X1 U10093 ( .A1(n10130), .A2(n9908), .ZN(n10128) );
  OR2_X1 U10094 ( .A1(n9909), .A2(n9907), .ZN(n10130) );
  XOR2_X1 U10095 ( .A(n10131), .B(n10132), .Z(n9907) );
  XOR2_X1 U10096 ( .A(n10133), .B(n10134), .Z(n10132) );
  OR2_X1 U10097 ( .A1(n10135), .A2(n10136), .ZN(n9909) );
  AND2_X1 U10098 ( .A1(n9905), .A2(n9904), .ZN(n10136) );
  AND2_X1 U10099 ( .A1(n9902), .A2(n10137), .ZN(n10135) );
  OR2_X1 U10100 ( .A1(n9904), .A2(n9905), .ZN(n10137) );
  OR2_X1 U10101 ( .A1(n8136), .A2(n9684), .ZN(n9905) );
  OR2_X1 U10102 ( .A1(n10138), .A2(n10139), .ZN(n9904) );
  AND2_X1 U10103 ( .A1(n9901), .A2(n9900), .ZN(n10139) );
  AND2_X1 U10104 ( .A1(n9898), .A2(n10140), .ZN(n10138) );
  OR2_X1 U10105 ( .A1(n9900), .A2(n9901), .ZN(n10140) );
  OR2_X1 U10106 ( .A1(n8131), .A2(n9684), .ZN(n9901) );
  OR2_X1 U10107 ( .A1(n10141), .A2(n10142), .ZN(n9900) );
  AND2_X1 U10108 ( .A1(n9897), .A2(n9896), .ZN(n10142) );
  AND2_X1 U10109 ( .A1(n9894), .A2(n10143), .ZN(n10141) );
  OR2_X1 U10110 ( .A1(n9896), .A2(n9897), .ZN(n10143) );
  OR2_X1 U10111 ( .A1(n8126), .A2(n9684), .ZN(n9897) );
  OR2_X1 U10112 ( .A1(n10144), .A2(n10145), .ZN(n9896) );
  AND2_X1 U10113 ( .A1(n9893), .A2(n9892), .ZN(n10145) );
  AND2_X1 U10114 ( .A1(n9890), .A2(n10146), .ZN(n10144) );
  OR2_X1 U10115 ( .A1(n9892), .A2(n9893), .ZN(n10146) );
  OR2_X1 U10116 ( .A1(n8121), .A2(n9684), .ZN(n9893) );
  OR2_X1 U10117 ( .A1(n10147), .A2(n10148), .ZN(n9892) );
  AND2_X1 U10118 ( .A1(n9889), .A2(n9888), .ZN(n10148) );
  AND2_X1 U10119 ( .A1(n9886), .A2(n10149), .ZN(n10147) );
  OR2_X1 U10120 ( .A1(n9888), .A2(n9889), .ZN(n10149) );
  OR2_X1 U10121 ( .A1(n8116), .A2(n9684), .ZN(n9889) );
  OR2_X1 U10122 ( .A1(n10150), .A2(n10151), .ZN(n9888) );
  AND2_X1 U10123 ( .A1(n9885), .A2(n9884), .ZN(n10151) );
  AND2_X1 U10124 ( .A1(n9882), .A2(n10152), .ZN(n10150) );
  OR2_X1 U10125 ( .A1(n9884), .A2(n9885), .ZN(n10152) );
  OR2_X1 U10126 ( .A1(n8111), .A2(n9684), .ZN(n9885) );
  OR2_X1 U10127 ( .A1(n10153), .A2(n10154), .ZN(n9884) );
  AND2_X1 U10128 ( .A1(n9878), .A2(n9881), .ZN(n10154) );
  AND2_X1 U10129 ( .A1(n9880), .A2(n10155), .ZN(n10153) );
  OR2_X1 U10130 ( .A1(n9881), .A2(n9878), .ZN(n10155) );
  OR2_X1 U10131 ( .A1(n8102), .A2(n9684), .ZN(n9878) );
  OR3_X1 U10132 ( .A1(n8349), .A2(n9875), .A3(n9684), .ZN(n9881) );
  INV_X1 U10133 ( .A(n10156), .ZN(n9880) );
  OR2_X1 U10134 ( .A1(n10157), .A2(n10158), .ZN(n10156) );
  AND2_X1 U10135 ( .A1(b_21_), .A2(n10159), .ZN(n10158) );
  OR2_X1 U10136 ( .A1(n10160), .A2(n7314), .ZN(n10159) );
  AND2_X1 U10137 ( .A1(a_30_), .A2(n9990), .ZN(n10160) );
  AND2_X1 U10138 ( .A1(b_20_), .A2(n10161), .ZN(n10157) );
  OR2_X1 U10139 ( .A1(n10162), .A2(n7318), .ZN(n10161) );
  AND2_X1 U10140 ( .A1(a_31_), .A2(n9875), .ZN(n10162) );
  XNOR2_X1 U10141 ( .A(n10163), .B(n10164), .ZN(n9882) );
  XNOR2_X1 U10142 ( .A(n10165), .B(n10166), .ZN(n10164) );
  XOR2_X1 U10143 ( .A(n10167), .B(n10168), .Z(n9886) );
  XOR2_X1 U10144 ( .A(n10169), .B(n10170), .Z(n10168) );
  XOR2_X1 U10145 ( .A(n10171), .B(n10172), .Z(n9890) );
  XOR2_X1 U10146 ( .A(n10173), .B(n10174), .Z(n10172) );
  XOR2_X1 U10147 ( .A(n10175), .B(n10176), .Z(n9894) );
  XOR2_X1 U10148 ( .A(n10177), .B(n10178), .Z(n10176) );
  XOR2_X1 U10149 ( .A(n10179), .B(n10180), .Z(n9898) );
  XOR2_X1 U10150 ( .A(n10181), .B(n10182), .Z(n10180) );
  XOR2_X1 U10151 ( .A(n10183), .B(n10184), .Z(n9902) );
  XOR2_X1 U10152 ( .A(n10185), .B(n10186), .Z(n10184) );
  XOR2_X1 U10153 ( .A(n10187), .B(n10188), .Z(n9910) );
  XOR2_X1 U10154 ( .A(n10189), .B(n10190), .Z(n10188) );
  XNOR2_X1 U10155 ( .A(n10191), .B(n10192), .ZN(n9914) );
  XNOR2_X1 U10156 ( .A(n10193), .B(n10194), .ZN(n10191) );
  XOR2_X1 U10157 ( .A(n10195), .B(n10196), .Z(n9918) );
  XOR2_X1 U10158 ( .A(n10197), .B(n10198), .Z(n10196) );
  XOR2_X1 U10159 ( .A(n10199), .B(n10200), .Z(n9922) );
  XOR2_X1 U10160 ( .A(n10201), .B(n10202), .Z(n10200) );
  XOR2_X1 U10161 ( .A(n10203), .B(n10204), .Z(n9926) );
  XOR2_X1 U10162 ( .A(n10205), .B(n10206), .Z(n10204) );
  XOR2_X1 U10163 ( .A(n10207), .B(n10208), .Z(n9930) );
  XOR2_X1 U10164 ( .A(n10209), .B(n10210), .Z(n10208) );
  XOR2_X1 U10165 ( .A(n10211), .B(n10212), .Z(n9934) );
  XOR2_X1 U10166 ( .A(n10213), .B(n10214), .Z(n10212) );
  XOR2_X1 U10167 ( .A(n10215), .B(n10216), .Z(n9938) );
  XOR2_X1 U10168 ( .A(n10217), .B(n10218), .Z(n10216) );
  XOR2_X1 U10169 ( .A(n10219), .B(n10220), .Z(n9942) );
  XOR2_X1 U10170 ( .A(n10221), .B(n10222), .Z(n10220) );
  XOR2_X1 U10171 ( .A(n10223), .B(n10224), .Z(n9946) );
  XOR2_X1 U10172 ( .A(n10225), .B(n10226), .Z(n10224) );
  XOR2_X1 U10173 ( .A(n10227), .B(n10228), .Z(n9950) );
  XOR2_X1 U10174 ( .A(n10229), .B(n10230), .Z(n10228) );
  XOR2_X1 U10175 ( .A(n10231), .B(n10232), .Z(n9954) );
  XOR2_X1 U10176 ( .A(n10233), .B(n10234), .Z(n10232) );
  XOR2_X1 U10177 ( .A(n10235), .B(n10236), .Z(n9958) );
  XOR2_X1 U10178 ( .A(n10237), .B(n10238), .Z(n10236) );
  XOR2_X1 U10179 ( .A(n10239), .B(n10240), .Z(n9962) );
  XOR2_X1 U10180 ( .A(n10241), .B(n10242), .Z(n10240) );
  XOR2_X1 U10181 ( .A(n10243), .B(n10244), .Z(n9966) );
  XOR2_X1 U10182 ( .A(n10245), .B(n10246), .Z(n10244) );
  XOR2_X1 U10183 ( .A(n10247), .B(n10248), .Z(n9970) );
  XOR2_X1 U10184 ( .A(n10249), .B(n10250), .Z(n10248) );
  XOR2_X1 U10185 ( .A(n10251), .B(n10252), .Z(n9974) );
  XOR2_X1 U10186 ( .A(n10253), .B(n10254), .Z(n10252) );
  XOR2_X1 U10187 ( .A(n10255), .B(n10256), .Z(n9978) );
  XOR2_X1 U10188 ( .A(n10257), .B(n10258), .Z(n10256) );
  XOR2_X1 U10189 ( .A(n10259), .B(n10260), .Z(n9178) );
  XOR2_X1 U10190 ( .A(n10261), .B(n10262), .Z(n10260) );
  XOR2_X1 U10191 ( .A(n10263), .B(n10264), .Z(n9159) );
  XOR2_X1 U10192 ( .A(n10265), .B(n10266), .Z(n10264) );
  XOR2_X1 U10193 ( .A(n10267), .B(n10268), .Z(n7983) );
  XOR2_X1 U10194 ( .A(n10269), .B(n10270), .Z(n10268) );
  XOR2_X1 U10195 ( .A(n10027), .B(n10271), .Z(n7958) );
  XOR2_X1 U10196 ( .A(n10026), .B(n10025), .Z(n10271) );
  OR2_X1 U10197 ( .A1(n7656), .A2(n9875), .ZN(n10025) );
  OR2_X1 U10198 ( .A1(n10272), .A2(n10273), .ZN(n10026) );
  AND2_X1 U10199 ( .A1(n10270), .A2(n10269), .ZN(n10273) );
  AND2_X1 U10200 ( .A1(n10267), .A2(n10274), .ZN(n10272) );
  OR2_X1 U10201 ( .A1(n10270), .A2(n10269), .ZN(n10274) );
  OR2_X1 U10202 ( .A1(n10275), .A2(n10276), .ZN(n10269) );
  AND2_X1 U10203 ( .A1(n10266), .A2(n10265), .ZN(n10276) );
  AND2_X1 U10204 ( .A1(n10263), .A2(n10277), .ZN(n10275) );
  OR2_X1 U10205 ( .A1(n10266), .A2(n10265), .ZN(n10277) );
  OR2_X1 U10206 ( .A1(n10278), .A2(n10279), .ZN(n10265) );
  AND2_X1 U10207 ( .A1(n10262), .A2(n10261), .ZN(n10279) );
  AND2_X1 U10208 ( .A1(n10259), .A2(n10280), .ZN(n10278) );
  OR2_X1 U10209 ( .A1(n10262), .A2(n10261), .ZN(n10280) );
  OR2_X1 U10210 ( .A1(n10281), .A2(n10282), .ZN(n10261) );
  AND2_X1 U10211 ( .A1(n10258), .A2(n10257), .ZN(n10282) );
  AND2_X1 U10212 ( .A1(n10255), .A2(n10283), .ZN(n10281) );
  OR2_X1 U10213 ( .A1(n10258), .A2(n10257), .ZN(n10283) );
  OR2_X1 U10214 ( .A1(n10284), .A2(n10285), .ZN(n10257) );
  AND2_X1 U10215 ( .A1(n10254), .A2(n10253), .ZN(n10285) );
  AND2_X1 U10216 ( .A1(n10251), .A2(n10286), .ZN(n10284) );
  OR2_X1 U10217 ( .A1(n10254), .A2(n10253), .ZN(n10286) );
  OR2_X1 U10218 ( .A1(n10287), .A2(n10288), .ZN(n10253) );
  AND2_X1 U10219 ( .A1(n10250), .A2(n10249), .ZN(n10288) );
  AND2_X1 U10220 ( .A1(n10247), .A2(n10289), .ZN(n10287) );
  OR2_X1 U10221 ( .A1(n10250), .A2(n10249), .ZN(n10289) );
  OR2_X1 U10222 ( .A1(n10290), .A2(n10291), .ZN(n10249) );
  AND2_X1 U10223 ( .A1(n10246), .A2(n10245), .ZN(n10291) );
  AND2_X1 U10224 ( .A1(n10243), .A2(n10292), .ZN(n10290) );
  OR2_X1 U10225 ( .A1(n10246), .A2(n10245), .ZN(n10292) );
  OR2_X1 U10226 ( .A1(n10293), .A2(n10294), .ZN(n10245) );
  AND2_X1 U10227 ( .A1(n10242), .A2(n10241), .ZN(n10294) );
  AND2_X1 U10228 ( .A1(n10239), .A2(n10295), .ZN(n10293) );
  OR2_X1 U10229 ( .A1(n10242), .A2(n10241), .ZN(n10295) );
  OR2_X1 U10230 ( .A1(n10296), .A2(n10297), .ZN(n10241) );
  AND2_X1 U10231 ( .A1(n10238), .A2(n10237), .ZN(n10297) );
  AND2_X1 U10232 ( .A1(n10235), .A2(n10298), .ZN(n10296) );
  OR2_X1 U10233 ( .A1(n10238), .A2(n10237), .ZN(n10298) );
  OR2_X1 U10234 ( .A1(n10299), .A2(n10300), .ZN(n10237) );
  AND2_X1 U10235 ( .A1(n10234), .A2(n10233), .ZN(n10300) );
  AND2_X1 U10236 ( .A1(n10231), .A2(n10301), .ZN(n10299) );
  OR2_X1 U10237 ( .A1(n10234), .A2(n10233), .ZN(n10301) );
  OR2_X1 U10238 ( .A1(n10302), .A2(n10303), .ZN(n10233) );
  AND2_X1 U10239 ( .A1(n10230), .A2(n10229), .ZN(n10303) );
  AND2_X1 U10240 ( .A1(n10227), .A2(n10304), .ZN(n10302) );
  OR2_X1 U10241 ( .A1(n10230), .A2(n10229), .ZN(n10304) );
  OR2_X1 U10242 ( .A1(n10305), .A2(n10306), .ZN(n10229) );
  AND2_X1 U10243 ( .A1(n10226), .A2(n10225), .ZN(n10306) );
  AND2_X1 U10244 ( .A1(n10223), .A2(n10307), .ZN(n10305) );
  OR2_X1 U10245 ( .A1(n10226), .A2(n10225), .ZN(n10307) );
  OR2_X1 U10246 ( .A1(n10308), .A2(n10309), .ZN(n10225) );
  AND2_X1 U10247 ( .A1(n10222), .A2(n10221), .ZN(n10309) );
  AND2_X1 U10248 ( .A1(n10219), .A2(n10310), .ZN(n10308) );
  OR2_X1 U10249 ( .A1(n10222), .A2(n10221), .ZN(n10310) );
  OR2_X1 U10250 ( .A1(n10311), .A2(n10312), .ZN(n10221) );
  AND2_X1 U10251 ( .A1(n10218), .A2(n10217), .ZN(n10312) );
  AND2_X1 U10252 ( .A1(n10215), .A2(n10313), .ZN(n10311) );
  OR2_X1 U10253 ( .A1(n10218), .A2(n10217), .ZN(n10313) );
  OR2_X1 U10254 ( .A1(n10314), .A2(n10315), .ZN(n10217) );
  AND2_X1 U10255 ( .A1(n10214), .A2(n10213), .ZN(n10315) );
  AND2_X1 U10256 ( .A1(n10211), .A2(n10316), .ZN(n10314) );
  OR2_X1 U10257 ( .A1(n10214), .A2(n10213), .ZN(n10316) );
  OR2_X1 U10258 ( .A1(n10317), .A2(n10318), .ZN(n10213) );
  AND2_X1 U10259 ( .A1(n10210), .A2(n10209), .ZN(n10318) );
  AND2_X1 U10260 ( .A1(n10207), .A2(n10319), .ZN(n10317) );
  OR2_X1 U10261 ( .A1(n10210), .A2(n10209), .ZN(n10319) );
  OR2_X1 U10262 ( .A1(n10320), .A2(n10321), .ZN(n10209) );
  AND2_X1 U10263 ( .A1(n10206), .A2(n10205), .ZN(n10321) );
  AND2_X1 U10264 ( .A1(n10203), .A2(n10322), .ZN(n10320) );
  OR2_X1 U10265 ( .A1(n10206), .A2(n10205), .ZN(n10322) );
  OR2_X1 U10266 ( .A1(n10323), .A2(n10324), .ZN(n10205) );
  AND2_X1 U10267 ( .A1(n10202), .A2(n10201), .ZN(n10324) );
  AND2_X1 U10268 ( .A1(n10199), .A2(n10325), .ZN(n10323) );
  OR2_X1 U10269 ( .A1(n10202), .A2(n10201), .ZN(n10325) );
  OR2_X1 U10270 ( .A1(n10326), .A2(n10327), .ZN(n10201) );
  AND2_X1 U10271 ( .A1(n10198), .A2(n10197), .ZN(n10327) );
  AND2_X1 U10272 ( .A1(n10195), .A2(n10328), .ZN(n10326) );
  OR2_X1 U10273 ( .A1(n10198), .A2(n10197), .ZN(n10328) );
  OR2_X1 U10274 ( .A1(n10329), .A2(n10330), .ZN(n10197) );
  AND2_X1 U10275 ( .A1(n10192), .A2(n10194), .ZN(n10330) );
  AND2_X1 U10276 ( .A1(n10331), .A2(n10193), .ZN(n10329) );
  OR2_X1 U10277 ( .A1(n10192), .A2(n10194), .ZN(n10331) );
  OR2_X1 U10278 ( .A1(n10332), .A2(n10333), .ZN(n10194) );
  AND2_X1 U10279 ( .A1(n10190), .A2(n10189), .ZN(n10333) );
  AND2_X1 U10280 ( .A1(n10187), .A2(n10334), .ZN(n10332) );
  OR2_X1 U10281 ( .A1(n10190), .A2(n10189), .ZN(n10334) );
  OR2_X1 U10282 ( .A1(n10335), .A2(n10336), .ZN(n10189) );
  AND2_X1 U10283 ( .A1(n10134), .A2(n10133), .ZN(n10336) );
  AND2_X1 U10284 ( .A1(n10131), .A2(n10337), .ZN(n10335) );
  OR2_X1 U10285 ( .A1(n10134), .A2(n10133), .ZN(n10337) );
  OR2_X1 U10286 ( .A1(n10338), .A2(n10339), .ZN(n10133) );
  AND2_X1 U10287 ( .A1(n10186), .A2(n10185), .ZN(n10339) );
  AND2_X1 U10288 ( .A1(n10183), .A2(n10340), .ZN(n10338) );
  OR2_X1 U10289 ( .A1(n10186), .A2(n10185), .ZN(n10340) );
  OR2_X1 U10290 ( .A1(n10341), .A2(n10342), .ZN(n10185) );
  AND2_X1 U10291 ( .A1(n10182), .A2(n10181), .ZN(n10342) );
  AND2_X1 U10292 ( .A1(n10179), .A2(n10343), .ZN(n10341) );
  OR2_X1 U10293 ( .A1(n10182), .A2(n10181), .ZN(n10343) );
  OR2_X1 U10294 ( .A1(n10344), .A2(n10345), .ZN(n10181) );
  AND2_X1 U10295 ( .A1(n10178), .A2(n10177), .ZN(n10345) );
  AND2_X1 U10296 ( .A1(n10175), .A2(n10346), .ZN(n10344) );
  OR2_X1 U10297 ( .A1(n10178), .A2(n10177), .ZN(n10346) );
  OR2_X1 U10298 ( .A1(n10347), .A2(n10348), .ZN(n10177) );
  AND2_X1 U10299 ( .A1(n10174), .A2(n10173), .ZN(n10348) );
  AND2_X1 U10300 ( .A1(n10171), .A2(n10349), .ZN(n10347) );
  OR2_X1 U10301 ( .A1(n10174), .A2(n10173), .ZN(n10349) );
  OR2_X1 U10302 ( .A1(n10350), .A2(n10351), .ZN(n10173) );
  AND2_X1 U10303 ( .A1(n10170), .A2(n10169), .ZN(n10351) );
  AND2_X1 U10304 ( .A1(n10167), .A2(n10352), .ZN(n10350) );
  OR2_X1 U10305 ( .A1(n10170), .A2(n10169), .ZN(n10352) );
  OR2_X1 U10306 ( .A1(n10353), .A2(n10354), .ZN(n10169) );
  AND2_X1 U10307 ( .A1(n10163), .A2(n10166), .ZN(n10354) );
  AND2_X1 U10308 ( .A1(n10165), .A2(n10355), .ZN(n10353) );
  OR2_X1 U10309 ( .A1(n10163), .A2(n10166), .ZN(n10355) );
  OR3_X1 U10310 ( .A1(n8349), .A2(n9990), .A3(n9875), .ZN(n10166) );
  OR2_X1 U10311 ( .A1(n8102), .A2(n9875), .ZN(n10163) );
  INV_X1 U10312 ( .A(n10356), .ZN(n10165) );
  OR2_X1 U10313 ( .A1(n10357), .A2(n10358), .ZN(n10356) );
  AND2_X1 U10314 ( .A1(b_20_), .A2(n10359), .ZN(n10358) );
  OR2_X1 U10315 ( .A1(n10360), .A2(n7314), .ZN(n10359) );
  AND2_X1 U10316 ( .A1(a_30_), .A2(n7909), .ZN(n10360) );
  AND2_X1 U10317 ( .A1(b_19_), .A2(n10361), .ZN(n10357) );
  OR2_X1 U10318 ( .A1(n10362), .A2(n7318), .ZN(n10361) );
  AND2_X1 U10319 ( .A1(a_31_), .A2(n9990), .ZN(n10362) );
  OR2_X1 U10320 ( .A1(n8111), .A2(n9875), .ZN(n10170) );
  XNOR2_X1 U10321 ( .A(n10363), .B(n10364), .ZN(n10167) );
  XNOR2_X1 U10322 ( .A(n10365), .B(n10366), .ZN(n10364) );
  OR2_X1 U10323 ( .A1(n8116), .A2(n9875), .ZN(n10174) );
  XOR2_X1 U10324 ( .A(n10367), .B(n10368), .Z(n10171) );
  XOR2_X1 U10325 ( .A(n10369), .B(n10370), .Z(n10368) );
  OR2_X1 U10326 ( .A1(n8121), .A2(n9875), .ZN(n10178) );
  XOR2_X1 U10327 ( .A(n10371), .B(n10372), .Z(n10175) );
  XOR2_X1 U10328 ( .A(n10373), .B(n10374), .Z(n10372) );
  OR2_X1 U10329 ( .A1(n8126), .A2(n9875), .ZN(n10182) );
  XOR2_X1 U10330 ( .A(n10375), .B(n10376), .Z(n10179) );
  XOR2_X1 U10331 ( .A(n10377), .B(n10378), .Z(n10376) );
  OR2_X1 U10332 ( .A1(n8131), .A2(n9875), .ZN(n10186) );
  XOR2_X1 U10333 ( .A(n10379), .B(n10380), .Z(n10183) );
  XOR2_X1 U10334 ( .A(n10381), .B(n10382), .Z(n10380) );
  OR2_X1 U10335 ( .A1(n8136), .A2(n9875), .ZN(n10134) );
  XOR2_X1 U10336 ( .A(n10383), .B(n10384), .Z(n10131) );
  XOR2_X1 U10337 ( .A(n10385), .B(n10386), .Z(n10384) );
  OR2_X1 U10338 ( .A1(n8141), .A2(n9875), .ZN(n10190) );
  XOR2_X1 U10339 ( .A(n10387), .B(n10388), .Z(n10187) );
  XOR2_X1 U10340 ( .A(n10389), .B(n10390), .Z(n10388) );
  XOR2_X1 U10341 ( .A(n10391), .B(n10392), .Z(n10192) );
  XOR2_X1 U10342 ( .A(n10393), .B(n10394), .Z(n10392) );
  OR2_X1 U10343 ( .A1(n8151), .A2(n9875), .ZN(n10198) );
  XOR2_X1 U10344 ( .A(n10395), .B(n10396), .Z(n10195) );
  XOR2_X1 U10345 ( .A(n10397), .B(n10398), .Z(n10396) );
  OR2_X1 U10346 ( .A1(n8156), .A2(n9875), .ZN(n10202) );
  XNOR2_X1 U10347 ( .A(n10399), .B(n10400), .ZN(n10199) );
  XNOR2_X1 U10348 ( .A(n10401), .B(n10402), .ZN(n10399) );
  OR2_X1 U10349 ( .A1(n8161), .A2(n9875), .ZN(n10206) );
  XOR2_X1 U10350 ( .A(n10403), .B(n10404), .Z(n10203) );
  XOR2_X1 U10351 ( .A(n10405), .B(n10406), .Z(n10404) );
  OR2_X1 U10352 ( .A1(n8166), .A2(n9875), .ZN(n10210) );
  XOR2_X1 U10353 ( .A(n10407), .B(n10408), .Z(n10207) );
  XOR2_X1 U10354 ( .A(n10409), .B(n10410), .Z(n10408) );
  OR2_X1 U10355 ( .A1(n8171), .A2(n9875), .ZN(n10214) );
  XOR2_X1 U10356 ( .A(n10411), .B(n10412), .Z(n10211) );
  XOR2_X1 U10357 ( .A(n10413), .B(n10414), .Z(n10412) );
  OR2_X1 U10358 ( .A1(n8176), .A2(n9875), .ZN(n10218) );
  XOR2_X1 U10359 ( .A(n10415), .B(n10416), .Z(n10215) );
  XOR2_X1 U10360 ( .A(n10417), .B(n10418), .Z(n10416) );
  OR2_X1 U10361 ( .A1(n8181), .A2(n9875), .ZN(n10222) );
  XOR2_X1 U10362 ( .A(n10419), .B(n10420), .Z(n10219) );
  XOR2_X1 U10363 ( .A(n10421), .B(n10422), .Z(n10420) );
  OR2_X1 U10364 ( .A1(n8186), .A2(n9875), .ZN(n10226) );
  XOR2_X1 U10365 ( .A(n10423), .B(n10424), .Z(n10223) );
  XOR2_X1 U10366 ( .A(n10425), .B(n10426), .Z(n10424) );
  OR2_X1 U10367 ( .A1(n8191), .A2(n9875), .ZN(n10230) );
  XOR2_X1 U10368 ( .A(n10427), .B(n10428), .Z(n10227) );
  XOR2_X1 U10369 ( .A(n10429), .B(n10430), .Z(n10428) );
  OR2_X1 U10370 ( .A1(n8196), .A2(n9875), .ZN(n10234) );
  XOR2_X1 U10371 ( .A(n10431), .B(n10432), .Z(n10231) );
  XOR2_X1 U10372 ( .A(n10433), .B(n10434), .Z(n10432) );
  OR2_X1 U10373 ( .A1(n8201), .A2(n9875), .ZN(n10238) );
  XOR2_X1 U10374 ( .A(n10435), .B(n10436), .Z(n10235) );
  XOR2_X1 U10375 ( .A(n10437), .B(n10438), .Z(n10436) );
  OR2_X1 U10376 ( .A1(n8206), .A2(n9875), .ZN(n10242) );
  XOR2_X1 U10377 ( .A(n10439), .B(n10440), .Z(n10239) );
  XOR2_X1 U10378 ( .A(n10441), .B(n10442), .Z(n10440) );
  OR2_X1 U10379 ( .A1(n8211), .A2(n9875), .ZN(n10246) );
  XOR2_X1 U10380 ( .A(n10443), .B(n10444), .Z(n10243) );
  XOR2_X1 U10381 ( .A(n10445), .B(n10446), .Z(n10444) );
  OR2_X1 U10382 ( .A1(n8216), .A2(n9875), .ZN(n10250) );
  XOR2_X1 U10383 ( .A(n10447), .B(n10448), .Z(n10247) );
  XOR2_X1 U10384 ( .A(n10449), .B(n10450), .Z(n10448) );
  OR2_X1 U10385 ( .A1(n8221), .A2(n9875), .ZN(n10254) );
  XOR2_X1 U10386 ( .A(n10451), .B(n10452), .Z(n10251) );
  XOR2_X1 U10387 ( .A(n10453), .B(n10454), .Z(n10452) );
  OR2_X1 U10388 ( .A1(n8226), .A2(n9875), .ZN(n10258) );
  XOR2_X1 U10389 ( .A(n10455), .B(n10456), .Z(n10255) );
  XOR2_X1 U10390 ( .A(n10457), .B(n10458), .Z(n10456) );
  OR2_X1 U10391 ( .A1(n7785), .A2(n9875), .ZN(n10262) );
  XOR2_X1 U10392 ( .A(n10459), .B(n10460), .Z(n10259) );
  XOR2_X1 U10393 ( .A(n10461), .B(n10462), .Z(n10460) );
  OR2_X1 U10394 ( .A1(n7777), .A2(n9875), .ZN(n10266) );
  XOR2_X1 U10395 ( .A(n10463), .B(n10464), .Z(n10263) );
  XOR2_X1 U10396 ( .A(n10465), .B(n10466), .Z(n10464) );
  OR2_X1 U10397 ( .A1(n7689), .A2(n9875), .ZN(n10270) );
  XOR2_X1 U10398 ( .A(n10467), .B(n10468), .Z(n10267) );
  XOR2_X1 U10399 ( .A(n10469), .B(n10470), .Z(n10468) );
  XOR2_X1 U10400 ( .A(n10034), .B(n10471), .Z(n10027) );
  XOR2_X1 U10401 ( .A(n10033), .B(n10032), .Z(n10471) );
  OR2_X1 U10402 ( .A1(n7689), .A2(n9990), .ZN(n10032) );
  OR2_X1 U10403 ( .A1(n10472), .A2(n10473), .ZN(n10033) );
  AND2_X1 U10404 ( .A1(n10470), .A2(n10469), .ZN(n10473) );
  AND2_X1 U10405 ( .A1(n10467), .A2(n10474), .ZN(n10472) );
  OR2_X1 U10406 ( .A1(n10470), .A2(n10469), .ZN(n10474) );
  OR2_X1 U10407 ( .A1(n10475), .A2(n10476), .ZN(n10469) );
  AND2_X1 U10408 ( .A1(n10466), .A2(n10465), .ZN(n10476) );
  AND2_X1 U10409 ( .A1(n10463), .A2(n10477), .ZN(n10475) );
  OR2_X1 U10410 ( .A1(n10466), .A2(n10465), .ZN(n10477) );
  OR2_X1 U10411 ( .A1(n10478), .A2(n10479), .ZN(n10465) );
  AND2_X1 U10412 ( .A1(n10462), .A2(n10461), .ZN(n10479) );
  AND2_X1 U10413 ( .A1(n10459), .A2(n10480), .ZN(n10478) );
  OR2_X1 U10414 ( .A1(n10462), .A2(n10461), .ZN(n10480) );
  OR2_X1 U10415 ( .A1(n10481), .A2(n10482), .ZN(n10461) );
  AND2_X1 U10416 ( .A1(n10458), .A2(n10457), .ZN(n10482) );
  AND2_X1 U10417 ( .A1(n10455), .A2(n10483), .ZN(n10481) );
  OR2_X1 U10418 ( .A1(n10458), .A2(n10457), .ZN(n10483) );
  OR2_X1 U10419 ( .A1(n10484), .A2(n10485), .ZN(n10457) );
  AND2_X1 U10420 ( .A1(n10454), .A2(n10453), .ZN(n10485) );
  AND2_X1 U10421 ( .A1(n10451), .A2(n10486), .ZN(n10484) );
  OR2_X1 U10422 ( .A1(n10454), .A2(n10453), .ZN(n10486) );
  OR2_X1 U10423 ( .A1(n10487), .A2(n10488), .ZN(n10453) );
  AND2_X1 U10424 ( .A1(n10450), .A2(n10449), .ZN(n10488) );
  AND2_X1 U10425 ( .A1(n10447), .A2(n10489), .ZN(n10487) );
  OR2_X1 U10426 ( .A1(n10450), .A2(n10449), .ZN(n10489) );
  OR2_X1 U10427 ( .A1(n10490), .A2(n10491), .ZN(n10449) );
  AND2_X1 U10428 ( .A1(n10446), .A2(n10445), .ZN(n10491) );
  AND2_X1 U10429 ( .A1(n10443), .A2(n10492), .ZN(n10490) );
  OR2_X1 U10430 ( .A1(n10446), .A2(n10445), .ZN(n10492) );
  OR2_X1 U10431 ( .A1(n10493), .A2(n10494), .ZN(n10445) );
  AND2_X1 U10432 ( .A1(n10442), .A2(n10441), .ZN(n10494) );
  AND2_X1 U10433 ( .A1(n10439), .A2(n10495), .ZN(n10493) );
  OR2_X1 U10434 ( .A1(n10442), .A2(n10441), .ZN(n10495) );
  OR2_X1 U10435 ( .A1(n10496), .A2(n10497), .ZN(n10441) );
  AND2_X1 U10436 ( .A1(n10438), .A2(n10437), .ZN(n10497) );
  AND2_X1 U10437 ( .A1(n10435), .A2(n10498), .ZN(n10496) );
  OR2_X1 U10438 ( .A1(n10438), .A2(n10437), .ZN(n10498) );
  OR2_X1 U10439 ( .A1(n10499), .A2(n10500), .ZN(n10437) );
  AND2_X1 U10440 ( .A1(n10434), .A2(n10433), .ZN(n10500) );
  AND2_X1 U10441 ( .A1(n10431), .A2(n10501), .ZN(n10499) );
  OR2_X1 U10442 ( .A1(n10434), .A2(n10433), .ZN(n10501) );
  OR2_X1 U10443 ( .A1(n10502), .A2(n10503), .ZN(n10433) );
  AND2_X1 U10444 ( .A1(n10430), .A2(n10429), .ZN(n10503) );
  AND2_X1 U10445 ( .A1(n10427), .A2(n10504), .ZN(n10502) );
  OR2_X1 U10446 ( .A1(n10430), .A2(n10429), .ZN(n10504) );
  OR2_X1 U10447 ( .A1(n10505), .A2(n10506), .ZN(n10429) );
  AND2_X1 U10448 ( .A1(n10426), .A2(n10425), .ZN(n10506) );
  AND2_X1 U10449 ( .A1(n10423), .A2(n10507), .ZN(n10505) );
  OR2_X1 U10450 ( .A1(n10426), .A2(n10425), .ZN(n10507) );
  OR2_X1 U10451 ( .A1(n10508), .A2(n10509), .ZN(n10425) );
  AND2_X1 U10452 ( .A1(n10422), .A2(n10421), .ZN(n10509) );
  AND2_X1 U10453 ( .A1(n10419), .A2(n10510), .ZN(n10508) );
  OR2_X1 U10454 ( .A1(n10422), .A2(n10421), .ZN(n10510) );
  OR2_X1 U10455 ( .A1(n10511), .A2(n10512), .ZN(n10421) );
  AND2_X1 U10456 ( .A1(n10418), .A2(n10417), .ZN(n10512) );
  AND2_X1 U10457 ( .A1(n10415), .A2(n10513), .ZN(n10511) );
  OR2_X1 U10458 ( .A1(n10418), .A2(n10417), .ZN(n10513) );
  OR2_X1 U10459 ( .A1(n10514), .A2(n10515), .ZN(n10417) );
  AND2_X1 U10460 ( .A1(n10414), .A2(n10413), .ZN(n10515) );
  AND2_X1 U10461 ( .A1(n10411), .A2(n10516), .ZN(n10514) );
  OR2_X1 U10462 ( .A1(n10414), .A2(n10413), .ZN(n10516) );
  OR2_X1 U10463 ( .A1(n10517), .A2(n10518), .ZN(n10413) );
  AND2_X1 U10464 ( .A1(n10410), .A2(n10409), .ZN(n10518) );
  AND2_X1 U10465 ( .A1(n10407), .A2(n10519), .ZN(n10517) );
  OR2_X1 U10466 ( .A1(n10410), .A2(n10409), .ZN(n10519) );
  OR2_X1 U10467 ( .A1(n10520), .A2(n10521), .ZN(n10409) );
  AND2_X1 U10468 ( .A1(n10406), .A2(n10405), .ZN(n10521) );
  AND2_X1 U10469 ( .A1(n10403), .A2(n10522), .ZN(n10520) );
  OR2_X1 U10470 ( .A1(n10406), .A2(n10405), .ZN(n10522) );
  OR2_X1 U10471 ( .A1(n10523), .A2(n10524), .ZN(n10405) );
  AND2_X1 U10472 ( .A1(n10400), .A2(n10402), .ZN(n10524) );
  AND2_X1 U10473 ( .A1(n10525), .A2(n10401), .ZN(n10523) );
  OR2_X1 U10474 ( .A1(n10400), .A2(n10402), .ZN(n10525) );
  OR2_X1 U10475 ( .A1(n10526), .A2(n10527), .ZN(n10402) );
  AND2_X1 U10476 ( .A1(n10398), .A2(n10397), .ZN(n10527) );
  AND2_X1 U10477 ( .A1(n10395), .A2(n10528), .ZN(n10526) );
  OR2_X1 U10478 ( .A1(n10398), .A2(n10397), .ZN(n10528) );
  OR2_X1 U10479 ( .A1(n10529), .A2(n10530), .ZN(n10397) );
  AND2_X1 U10480 ( .A1(n10394), .A2(n10393), .ZN(n10530) );
  AND2_X1 U10481 ( .A1(n10391), .A2(n10531), .ZN(n10529) );
  OR2_X1 U10482 ( .A1(n10394), .A2(n10393), .ZN(n10531) );
  OR2_X1 U10483 ( .A1(n10532), .A2(n10533), .ZN(n10393) );
  AND2_X1 U10484 ( .A1(n10390), .A2(n10389), .ZN(n10533) );
  AND2_X1 U10485 ( .A1(n10387), .A2(n10534), .ZN(n10532) );
  OR2_X1 U10486 ( .A1(n10390), .A2(n10389), .ZN(n10534) );
  OR2_X1 U10487 ( .A1(n10535), .A2(n10536), .ZN(n10389) );
  AND2_X1 U10488 ( .A1(n10386), .A2(n10385), .ZN(n10536) );
  AND2_X1 U10489 ( .A1(n10383), .A2(n10537), .ZN(n10535) );
  OR2_X1 U10490 ( .A1(n10386), .A2(n10385), .ZN(n10537) );
  OR2_X1 U10491 ( .A1(n10538), .A2(n10539), .ZN(n10385) );
  AND2_X1 U10492 ( .A1(n10382), .A2(n10381), .ZN(n10539) );
  AND2_X1 U10493 ( .A1(n10379), .A2(n10540), .ZN(n10538) );
  OR2_X1 U10494 ( .A1(n10382), .A2(n10381), .ZN(n10540) );
  OR2_X1 U10495 ( .A1(n10541), .A2(n10542), .ZN(n10381) );
  AND2_X1 U10496 ( .A1(n10378), .A2(n10377), .ZN(n10542) );
  AND2_X1 U10497 ( .A1(n10375), .A2(n10543), .ZN(n10541) );
  OR2_X1 U10498 ( .A1(n10378), .A2(n10377), .ZN(n10543) );
  OR2_X1 U10499 ( .A1(n10544), .A2(n10545), .ZN(n10377) );
  AND2_X1 U10500 ( .A1(n10374), .A2(n10373), .ZN(n10545) );
  AND2_X1 U10501 ( .A1(n10371), .A2(n10546), .ZN(n10544) );
  OR2_X1 U10502 ( .A1(n10374), .A2(n10373), .ZN(n10546) );
  OR2_X1 U10503 ( .A1(n10547), .A2(n10548), .ZN(n10373) );
  AND2_X1 U10504 ( .A1(n10370), .A2(n10369), .ZN(n10548) );
  AND2_X1 U10505 ( .A1(n10367), .A2(n10549), .ZN(n10547) );
  OR2_X1 U10506 ( .A1(n10370), .A2(n10369), .ZN(n10549) );
  OR2_X1 U10507 ( .A1(n10550), .A2(n10551), .ZN(n10369) );
  AND2_X1 U10508 ( .A1(n10363), .A2(n10366), .ZN(n10551) );
  AND2_X1 U10509 ( .A1(n10365), .A2(n10552), .ZN(n10550) );
  OR2_X1 U10510 ( .A1(n10363), .A2(n10366), .ZN(n10552) );
  OR3_X1 U10511 ( .A1(n8349), .A2(n7909), .A3(n9990), .ZN(n10366) );
  OR2_X1 U10512 ( .A1(n8102), .A2(n9990), .ZN(n10363) );
  INV_X1 U10513 ( .A(n10553), .ZN(n10365) );
  OR2_X1 U10514 ( .A1(n10554), .A2(n10555), .ZN(n10553) );
  AND2_X1 U10515 ( .A1(b_19_), .A2(n10556), .ZN(n10555) );
  OR2_X1 U10516 ( .A1(n10557), .A2(n7314), .ZN(n10556) );
  AND2_X1 U10517 ( .A1(a_30_), .A2(n7877), .ZN(n10557) );
  AND2_X1 U10518 ( .A1(b_18_), .A2(n10558), .ZN(n10554) );
  OR2_X1 U10519 ( .A1(n10559), .A2(n7318), .ZN(n10558) );
  AND2_X1 U10520 ( .A1(a_31_), .A2(n7909), .ZN(n10559) );
  OR2_X1 U10521 ( .A1(n8111), .A2(n9990), .ZN(n10370) );
  XNOR2_X1 U10522 ( .A(n10560), .B(n10561), .ZN(n10367) );
  XNOR2_X1 U10523 ( .A(n10562), .B(n10563), .ZN(n10561) );
  OR2_X1 U10524 ( .A1(n8116), .A2(n9990), .ZN(n10374) );
  XOR2_X1 U10525 ( .A(n10564), .B(n10565), .Z(n10371) );
  XOR2_X1 U10526 ( .A(n10566), .B(n10567), .Z(n10565) );
  OR2_X1 U10527 ( .A1(n8121), .A2(n9990), .ZN(n10378) );
  XOR2_X1 U10528 ( .A(n10568), .B(n10569), .Z(n10375) );
  XOR2_X1 U10529 ( .A(n10570), .B(n10571), .Z(n10569) );
  OR2_X1 U10530 ( .A1(n8126), .A2(n9990), .ZN(n10382) );
  XOR2_X1 U10531 ( .A(n10572), .B(n10573), .Z(n10379) );
  XOR2_X1 U10532 ( .A(n10574), .B(n10575), .Z(n10573) );
  OR2_X1 U10533 ( .A1(n8131), .A2(n9990), .ZN(n10386) );
  XOR2_X1 U10534 ( .A(n10576), .B(n10577), .Z(n10383) );
  XOR2_X1 U10535 ( .A(n10578), .B(n10579), .Z(n10577) );
  OR2_X1 U10536 ( .A1(n8136), .A2(n9990), .ZN(n10390) );
  XOR2_X1 U10537 ( .A(n10580), .B(n10581), .Z(n10387) );
  XOR2_X1 U10538 ( .A(n10582), .B(n10583), .Z(n10581) );
  OR2_X1 U10539 ( .A1(n8141), .A2(n9990), .ZN(n10394) );
  XOR2_X1 U10540 ( .A(n10584), .B(n10585), .Z(n10391) );
  XOR2_X1 U10541 ( .A(n10586), .B(n10587), .Z(n10585) );
  OR2_X1 U10542 ( .A1(n8146), .A2(n9990), .ZN(n10398) );
  XOR2_X1 U10543 ( .A(n10588), .B(n10589), .Z(n10395) );
  XOR2_X1 U10544 ( .A(n10590), .B(n10591), .Z(n10589) );
  XOR2_X1 U10545 ( .A(n10592), .B(n10593), .Z(n10400) );
  XOR2_X1 U10546 ( .A(n10594), .B(n10595), .Z(n10593) );
  OR2_X1 U10547 ( .A1(n8156), .A2(n9990), .ZN(n10406) );
  XOR2_X1 U10548 ( .A(n10596), .B(n10597), .Z(n10403) );
  XOR2_X1 U10549 ( .A(n10598), .B(n10599), .Z(n10597) );
  OR2_X1 U10550 ( .A1(n8161), .A2(n9990), .ZN(n10410) );
  XNOR2_X1 U10551 ( .A(n10600), .B(n10601), .ZN(n10407) );
  XNOR2_X1 U10552 ( .A(n10602), .B(n10603), .ZN(n10600) );
  OR2_X1 U10553 ( .A1(n8166), .A2(n9990), .ZN(n10414) );
  XOR2_X1 U10554 ( .A(n10604), .B(n10605), .Z(n10411) );
  XOR2_X1 U10555 ( .A(n10606), .B(n10607), .Z(n10605) );
  OR2_X1 U10556 ( .A1(n8171), .A2(n9990), .ZN(n10418) );
  XOR2_X1 U10557 ( .A(n10608), .B(n10609), .Z(n10415) );
  XOR2_X1 U10558 ( .A(n10610), .B(n10611), .Z(n10609) );
  OR2_X1 U10559 ( .A1(n8176), .A2(n9990), .ZN(n10422) );
  XOR2_X1 U10560 ( .A(n10612), .B(n10613), .Z(n10419) );
  XOR2_X1 U10561 ( .A(n10614), .B(n10615), .Z(n10613) );
  OR2_X1 U10562 ( .A1(n8181), .A2(n9990), .ZN(n10426) );
  XOR2_X1 U10563 ( .A(n10616), .B(n10617), .Z(n10423) );
  XOR2_X1 U10564 ( .A(n10618), .B(n10619), .Z(n10617) );
  OR2_X1 U10565 ( .A1(n8186), .A2(n9990), .ZN(n10430) );
  XOR2_X1 U10566 ( .A(n10620), .B(n10621), .Z(n10427) );
  XOR2_X1 U10567 ( .A(n10622), .B(n10623), .Z(n10621) );
  OR2_X1 U10568 ( .A1(n8191), .A2(n9990), .ZN(n10434) );
  XOR2_X1 U10569 ( .A(n10624), .B(n10625), .Z(n10431) );
  XOR2_X1 U10570 ( .A(n10626), .B(n10627), .Z(n10625) );
  OR2_X1 U10571 ( .A1(n8196), .A2(n9990), .ZN(n10438) );
  XOR2_X1 U10572 ( .A(n10628), .B(n10629), .Z(n10435) );
  XOR2_X1 U10573 ( .A(n10630), .B(n10631), .Z(n10629) );
  OR2_X1 U10574 ( .A1(n8201), .A2(n9990), .ZN(n10442) );
  XOR2_X1 U10575 ( .A(n10632), .B(n10633), .Z(n10439) );
  XOR2_X1 U10576 ( .A(n10634), .B(n10635), .Z(n10633) );
  OR2_X1 U10577 ( .A1(n8206), .A2(n9990), .ZN(n10446) );
  XOR2_X1 U10578 ( .A(n10636), .B(n10637), .Z(n10443) );
  XOR2_X1 U10579 ( .A(n10638), .B(n10639), .Z(n10637) );
  OR2_X1 U10580 ( .A1(n8211), .A2(n9990), .ZN(n10450) );
  XOR2_X1 U10581 ( .A(n10640), .B(n10641), .Z(n10447) );
  XOR2_X1 U10582 ( .A(n10642), .B(n10643), .Z(n10641) );
  OR2_X1 U10583 ( .A1(n8216), .A2(n9990), .ZN(n10454) );
  XOR2_X1 U10584 ( .A(n10644), .B(n10645), .Z(n10451) );
  XOR2_X1 U10585 ( .A(n10646), .B(n10647), .Z(n10645) );
  OR2_X1 U10586 ( .A1(n8221), .A2(n9990), .ZN(n10458) );
  XOR2_X1 U10587 ( .A(n10648), .B(n10649), .Z(n10455) );
  XOR2_X1 U10588 ( .A(n10650), .B(n10651), .Z(n10649) );
  OR2_X1 U10589 ( .A1(n8226), .A2(n9990), .ZN(n10462) );
  XOR2_X1 U10590 ( .A(n10652), .B(n10653), .Z(n10459) );
  XOR2_X1 U10591 ( .A(n10654), .B(n10655), .Z(n10653) );
  OR2_X1 U10592 ( .A1(n7785), .A2(n9990), .ZN(n10466) );
  XOR2_X1 U10593 ( .A(n10656), .B(n10657), .Z(n10463) );
  XOR2_X1 U10594 ( .A(n10658), .B(n10659), .Z(n10657) );
  OR2_X1 U10595 ( .A1(n7777), .A2(n9990), .ZN(n10470) );
  XOR2_X1 U10596 ( .A(n10660), .B(n10661), .Z(n10467) );
  XOR2_X1 U10597 ( .A(n10662), .B(n10663), .Z(n10661) );
  XOR2_X1 U10598 ( .A(n10041), .B(n10664), .Z(n10034) );
  XOR2_X1 U10599 ( .A(n10040), .B(n10039), .Z(n10664) );
  OR2_X1 U10600 ( .A1(n7777), .A2(n7909), .ZN(n10039) );
  OR2_X1 U10601 ( .A1(n10665), .A2(n10666), .ZN(n10040) );
  AND2_X1 U10602 ( .A1(n10663), .A2(n10662), .ZN(n10666) );
  AND2_X1 U10603 ( .A1(n10660), .A2(n10667), .ZN(n10665) );
  OR2_X1 U10604 ( .A1(n10663), .A2(n10662), .ZN(n10667) );
  OR2_X1 U10605 ( .A1(n10668), .A2(n10669), .ZN(n10662) );
  AND2_X1 U10606 ( .A1(n10659), .A2(n10658), .ZN(n10669) );
  AND2_X1 U10607 ( .A1(n10656), .A2(n10670), .ZN(n10668) );
  OR2_X1 U10608 ( .A1(n10659), .A2(n10658), .ZN(n10670) );
  OR2_X1 U10609 ( .A1(n10671), .A2(n10672), .ZN(n10658) );
  AND2_X1 U10610 ( .A1(n10655), .A2(n10654), .ZN(n10672) );
  AND2_X1 U10611 ( .A1(n10652), .A2(n10673), .ZN(n10671) );
  OR2_X1 U10612 ( .A1(n10655), .A2(n10654), .ZN(n10673) );
  OR2_X1 U10613 ( .A1(n10674), .A2(n10675), .ZN(n10654) );
  AND2_X1 U10614 ( .A1(n10651), .A2(n10650), .ZN(n10675) );
  AND2_X1 U10615 ( .A1(n10648), .A2(n10676), .ZN(n10674) );
  OR2_X1 U10616 ( .A1(n10651), .A2(n10650), .ZN(n10676) );
  OR2_X1 U10617 ( .A1(n10677), .A2(n10678), .ZN(n10650) );
  AND2_X1 U10618 ( .A1(n10647), .A2(n10646), .ZN(n10678) );
  AND2_X1 U10619 ( .A1(n10644), .A2(n10679), .ZN(n10677) );
  OR2_X1 U10620 ( .A1(n10647), .A2(n10646), .ZN(n10679) );
  OR2_X1 U10621 ( .A1(n10680), .A2(n10681), .ZN(n10646) );
  AND2_X1 U10622 ( .A1(n10643), .A2(n10642), .ZN(n10681) );
  AND2_X1 U10623 ( .A1(n10640), .A2(n10682), .ZN(n10680) );
  OR2_X1 U10624 ( .A1(n10643), .A2(n10642), .ZN(n10682) );
  OR2_X1 U10625 ( .A1(n10683), .A2(n10684), .ZN(n10642) );
  AND2_X1 U10626 ( .A1(n10639), .A2(n10638), .ZN(n10684) );
  AND2_X1 U10627 ( .A1(n10636), .A2(n10685), .ZN(n10683) );
  OR2_X1 U10628 ( .A1(n10639), .A2(n10638), .ZN(n10685) );
  OR2_X1 U10629 ( .A1(n10686), .A2(n10687), .ZN(n10638) );
  AND2_X1 U10630 ( .A1(n10635), .A2(n10634), .ZN(n10687) );
  AND2_X1 U10631 ( .A1(n10632), .A2(n10688), .ZN(n10686) );
  OR2_X1 U10632 ( .A1(n10635), .A2(n10634), .ZN(n10688) );
  OR2_X1 U10633 ( .A1(n10689), .A2(n10690), .ZN(n10634) );
  AND2_X1 U10634 ( .A1(n10631), .A2(n10630), .ZN(n10690) );
  AND2_X1 U10635 ( .A1(n10628), .A2(n10691), .ZN(n10689) );
  OR2_X1 U10636 ( .A1(n10631), .A2(n10630), .ZN(n10691) );
  OR2_X1 U10637 ( .A1(n10692), .A2(n10693), .ZN(n10630) );
  AND2_X1 U10638 ( .A1(n10627), .A2(n10626), .ZN(n10693) );
  AND2_X1 U10639 ( .A1(n10624), .A2(n10694), .ZN(n10692) );
  OR2_X1 U10640 ( .A1(n10627), .A2(n10626), .ZN(n10694) );
  OR2_X1 U10641 ( .A1(n10695), .A2(n10696), .ZN(n10626) );
  AND2_X1 U10642 ( .A1(n10623), .A2(n10622), .ZN(n10696) );
  AND2_X1 U10643 ( .A1(n10620), .A2(n10697), .ZN(n10695) );
  OR2_X1 U10644 ( .A1(n10623), .A2(n10622), .ZN(n10697) );
  OR2_X1 U10645 ( .A1(n10698), .A2(n10699), .ZN(n10622) );
  AND2_X1 U10646 ( .A1(n10619), .A2(n10618), .ZN(n10699) );
  AND2_X1 U10647 ( .A1(n10616), .A2(n10700), .ZN(n10698) );
  OR2_X1 U10648 ( .A1(n10619), .A2(n10618), .ZN(n10700) );
  OR2_X1 U10649 ( .A1(n10701), .A2(n10702), .ZN(n10618) );
  AND2_X1 U10650 ( .A1(n10615), .A2(n10614), .ZN(n10702) );
  AND2_X1 U10651 ( .A1(n10612), .A2(n10703), .ZN(n10701) );
  OR2_X1 U10652 ( .A1(n10615), .A2(n10614), .ZN(n10703) );
  OR2_X1 U10653 ( .A1(n10704), .A2(n10705), .ZN(n10614) );
  AND2_X1 U10654 ( .A1(n10611), .A2(n10610), .ZN(n10705) );
  AND2_X1 U10655 ( .A1(n10608), .A2(n10706), .ZN(n10704) );
  OR2_X1 U10656 ( .A1(n10611), .A2(n10610), .ZN(n10706) );
  OR2_X1 U10657 ( .A1(n10707), .A2(n10708), .ZN(n10610) );
  AND2_X1 U10658 ( .A1(n10607), .A2(n10606), .ZN(n10708) );
  AND2_X1 U10659 ( .A1(n10604), .A2(n10709), .ZN(n10707) );
  OR2_X1 U10660 ( .A1(n10607), .A2(n10606), .ZN(n10709) );
  OR2_X1 U10661 ( .A1(n10710), .A2(n10711), .ZN(n10606) );
  AND2_X1 U10662 ( .A1(n10601), .A2(n10603), .ZN(n10711) );
  AND2_X1 U10663 ( .A1(n10712), .A2(n10602), .ZN(n10710) );
  OR2_X1 U10664 ( .A1(n10601), .A2(n10603), .ZN(n10712) );
  OR2_X1 U10665 ( .A1(n10713), .A2(n10714), .ZN(n10603) );
  AND2_X1 U10666 ( .A1(n10599), .A2(n10598), .ZN(n10714) );
  AND2_X1 U10667 ( .A1(n10596), .A2(n10715), .ZN(n10713) );
  OR2_X1 U10668 ( .A1(n10599), .A2(n10598), .ZN(n10715) );
  OR2_X1 U10669 ( .A1(n10716), .A2(n10717), .ZN(n10598) );
  AND2_X1 U10670 ( .A1(n10595), .A2(n10594), .ZN(n10717) );
  AND2_X1 U10671 ( .A1(n10592), .A2(n10718), .ZN(n10716) );
  OR2_X1 U10672 ( .A1(n10595), .A2(n10594), .ZN(n10718) );
  OR2_X1 U10673 ( .A1(n10719), .A2(n10720), .ZN(n10594) );
  AND2_X1 U10674 ( .A1(n10591), .A2(n10590), .ZN(n10720) );
  AND2_X1 U10675 ( .A1(n10588), .A2(n10721), .ZN(n10719) );
  OR2_X1 U10676 ( .A1(n10591), .A2(n10590), .ZN(n10721) );
  OR2_X1 U10677 ( .A1(n10722), .A2(n10723), .ZN(n10590) );
  AND2_X1 U10678 ( .A1(n10587), .A2(n10586), .ZN(n10723) );
  AND2_X1 U10679 ( .A1(n10584), .A2(n10724), .ZN(n10722) );
  OR2_X1 U10680 ( .A1(n10587), .A2(n10586), .ZN(n10724) );
  OR2_X1 U10681 ( .A1(n10725), .A2(n10726), .ZN(n10586) );
  AND2_X1 U10682 ( .A1(n10583), .A2(n10582), .ZN(n10726) );
  AND2_X1 U10683 ( .A1(n10580), .A2(n10727), .ZN(n10725) );
  OR2_X1 U10684 ( .A1(n10583), .A2(n10582), .ZN(n10727) );
  OR2_X1 U10685 ( .A1(n10728), .A2(n10729), .ZN(n10582) );
  AND2_X1 U10686 ( .A1(n10579), .A2(n10578), .ZN(n10729) );
  AND2_X1 U10687 ( .A1(n10576), .A2(n10730), .ZN(n10728) );
  OR2_X1 U10688 ( .A1(n10579), .A2(n10578), .ZN(n10730) );
  OR2_X1 U10689 ( .A1(n10731), .A2(n10732), .ZN(n10578) );
  AND2_X1 U10690 ( .A1(n10575), .A2(n10574), .ZN(n10732) );
  AND2_X1 U10691 ( .A1(n10572), .A2(n10733), .ZN(n10731) );
  OR2_X1 U10692 ( .A1(n10575), .A2(n10574), .ZN(n10733) );
  OR2_X1 U10693 ( .A1(n10734), .A2(n10735), .ZN(n10574) );
  AND2_X1 U10694 ( .A1(n10571), .A2(n10570), .ZN(n10735) );
  AND2_X1 U10695 ( .A1(n10568), .A2(n10736), .ZN(n10734) );
  OR2_X1 U10696 ( .A1(n10571), .A2(n10570), .ZN(n10736) );
  OR2_X1 U10697 ( .A1(n10737), .A2(n10738), .ZN(n10570) );
  AND2_X1 U10698 ( .A1(n10567), .A2(n10566), .ZN(n10738) );
  AND2_X1 U10699 ( .A1(n10564), .A2(n10739), .ZN(n10737) );
  OR2_X1 U10700 ( .A1(n10567), .A2(n10566), .ZN(n10739) );
  OR2_X1 U10701 ( .A1(n10740), .A2(n10741), .ZN(n10566) );
  AND2_X1 U10702 ( .A1(n10560), .A2(n10563), .ZN(n10741) );
  AND2_X1 U10703 ( .A1(n10562), .A2(n10742), .ZN(n10740) );
  OR2_X1 U10704 ( .A1(n10560), .A2(n10563), .ZN(n10742) );
  OR3_X1 U10705 ( .A1(n8349), .A2(n7877), .A3(n7909), .ZN(n10563) );
  OR2_X1 U10706 ( .A1(n8102), .A2(n7909), .ZN(n10560) );
  INV_X1 U10707 ( .A(n10743), .ZN(n10562) );
  OR2_X1 U10708 ( .A1(n10744), .A2(n10745), .ZN(n10743) );
  AND2_X1 U10709 ( .A1(b_18_), .A2(n10746), .ZN(n10745) );
  OR2_X1 U10710 ( .A1(n10747), .A2(n7314), .ZN(n10746) );
  AND2_X1 U10711 ( .A1(a_30_), .A2(n7852), .ZN(n10747) );
  AND2_X1 U10712 ( .A1(b_17_), .A2(n10748), .ZN(n10744) );
  OR2_X1 U10713 ( .A1(n10749), .A2(n7318), .ZN(n10748) );
  AND2_X1 U10714 ( .A1(a_31_), .A2(n7877), .ZN(n10749) );
  OR2_X1 U10715 ( .A1(n8111), .A2(n7909), .ZN(n10567) );
  XNOR2_X1 U10716 ( .A(n10750), .B(n10751), .ZN(n10564) );
  XNOR2_X1 U10717 ( .A(n10752), .B(n10753), .ZN(n10751) );
  OR2_X1 U10718 ( .A1(n8116), .A2(n7909), .ZN(n10571) );
  XOR2_X1 U10719 ( .A(n10754), .B(n10755), .Z(n10568) );
  XOR2_X1 U10720 ( .A(n10756), .B(n10757), .Z(n10755) );
  OR2_X1 U10721 ( .A1(n8121), .A2(n7909), .ZN(n10575) );
  XOR2_X1 U10722 ( .A(n10758), .B(n10759), .Z(n10572) );
  XOR2_X1 U10723 ( .A(n10760), .B(n10761), .Z(n10759) );
  OR2_X1 U10724 ( .A1(n8126), .A2(n7909), .ZN(n10579) );
  XOR2_X1 U10725 ( .A(n10762), .B(n10763), .Z(n10576) );
  XOR2_X1 U10726 ( .A(n10764), .B(n10765), .Z(n10763) );
  OR2_X1 U10727 ( .A1(n8131), .A2(n7909), .ZN(n10583) );
  XOR2_X1 U10728 ( .A(n10766), .B(n10767), .Z(n10580) );
  XOR2_X1 U10729 ( .A(n10768), .B(n10769), .Z(n10767) );
  OR2_X1 U10730 ( .A1(n8136), .A2(n7909), .ZN(n10587) );
  XOR2_X1 U10731 ( .A(n10770), .B(n10771), .Z(n10584) );
  XOR2_X1 U10732 ( .A(n10772), .B(n10773), .Z(n10771) );
  OR2_X1 U10733 ( .A1(n8141), .A2(n7909), .ZN(n10591) );
  XOR2_X1 U10734 ( .A(n10774), .B(n10775), .Z(n10588) );
  XOR2_X1 U10735 ( .A(n10776), .B(n10777), .Z(n10775) );
  OR2_X1 U10736 ( .A1(n8146), .A2(n7909), .ZN(n10595) );
  XOR2_X1 U10737 ( .A(n10778), .B(n10779), .Z(n10592) );
  XOR2_X1 U10738 ( .A(n10780), .B(n10781), .Z(n10779) );
  OR2_X1 U10739 ( .A1(n8151), .A2(n7909), .ZN(n10599) );
  XOR2_X1 U10740 ( .A(n10782), .B(n10783), .Z(n10596) );
  XOR2_X1 U10741 ( .A(n10784), .B(n10785), .Z(n10783) );
  XOR2_X1 U10742 ( .A(n10786), .B(n10787), .Z(n10601) );
  XOR2_X1 U10743 ( .A(n10788), .B(n10789), .Z(n10787) );
  OR2_X1 U10744 ( .A1(n8161), .A2(n7909), .ZN(n10607) );
  XOR2_X1 U10745 ( .A(n10790), .B(n10791), .Z(n10604) );
  XOR2_X1 U10746 ( .A(n10792), .B(n10793), .Z(n10791) );
  OR2_X1 U10747 ( .A1(n8166), .A2(n7909), .ZN(n10611) );
  XNOR2_X1 U10748 ( .A(n10794), .B(n10795), .ZN(n10608) );
  XNOR2_X1 U10749 ( .A(n10796), .B(n10797), .ZN(n10794) );
  OR2_X1 U10750 ( .A1(n8171), .A2(n7909), .ZN(n10615) );
  XOR2_X1 U10751 ( .A(n10798), .B(n10799), .Z(n10612) );
  XOR2_X1 U10752 ( .A(n10800), .B(n10801), .Z(n10799) );
  OR2_X1 U10753 ( .A1(n8176), .A2(n7909), .ZN(n10619) );
  XOR2_X1 U10754 ( .A(n10802), .B(n10803), .Z(n10616) );
  XOR2_X1 U10755 ( .A(n10804), .B(n10805), .Z(n10803) );
  OR2_X1 U10756 ( .A1(n8181), .A2(n7909), .ZN(n10623) );
  XOR2_X1 U10757 ( .A(n10806), .B(n10807), .Z(n10620) );
  XOR2_X1 U10758 ( .A(n10808), .B(n10809), .Z(n10807) );
  OR2_X1 U10759 ( .A1(n8186), .A2(n7909), .ZN(n10627) );
  XOR2_X1 U10760 ( .A(n10810), .B(n10811), .Z(n10624) );
  XOR2_X1 U10761 ( .A(n10812), .B(n10813), .Z(n10811) );
  OR2_X1 U10762 ( .A1(n8191), .A2(n7909), .ZN(n10631) );
  XOR2_X1 U10763 ( .A(n10814), .B(n10815), .Z(n10628) );
  XOR2_X1 U10764 ( .A(n10816), .B(n10817), .Z(n10815) );
  OR2_X1 U10765 ( .A1(n8196), .A2(n7909), .ZN(n10635) );
  XOR2_X1 U10766 ( .A(n10818), .B(n10819), .Z(n10632) );
  XOR2_X1 U10767 ( .A(n10820), .B(n10821), .Z(n10819) );
  OR2_X1 U10768 ( .A1(n8201), .A2(n7909), .ZN(n10639) );
  XOR2_X1 U10769 ( .A(n10822), .B(n10823), .Z(n10636) );
  XOR2_X1 U10770 ( .A(n10824), .B(n10825), .Z(n10823) );
  OR2_X1 U10771 ( .A1(n8206), .A2(n7909), .ZN(n10643) );
  XOR2_X1 U10772 ( .A(n10826), .B(n10827), .Z(n10640) );
  XOR2_X1 U10773 ( .A(n10828), .B(n10829), .Z(n10827) );
  OR2_X1 U10774 ( .A1(n8211), .A2(n7909), .ZN(n10647) );
  XOR2_X1 U10775 ( .A(n10830), .B(n10831), .Z(n10644) );
  XOR2_X1 U10776 ( .A(n10832), .B(n10833), .Z(n10831) );
  OR2_X1 U10777 ( .A1(n8216), .A2(n7909), .ZN(n10651) );
  XOR2_X1 U10778 ( .A(n10834), .B(n10835), .Z(n10648) );
  XOR2_X1 U10779 ( .A(n10836), .B(n10837), .Z(n10835) );
  OR2_X1 U10780 ( .A1(n8221), .A2(n7909), .ZN(n10655) );
  XOR2_X1 U10781 ( .A(n10838), .B(n10839), .Z(n10652) );
  XOR2_X1 U10782 ( .A(n10840), .B(n10841), .Z(n10839) );
  OR2_X1 U10783 ( .A1(n8226), .A2(n7909), .ZN(n10659) );
  XOR2_X1 U10784 ( .A(n10842), .B(n10843), .Z(n10656) );
  XOR2_X1 U10785 ( .A(n10844), .B(n10845), .Z(n10843) );
  OR2_X1 U10786 ( .A1(n7785), .A2(n7909), .ZN(n10663) );
  XOR2_X1 U10787 ( .A(n10846), .B(n10847), .Z(n10660) );
  XOR2_X1 U10788 ( .A(n10848), .B(n10849), .Z(n10847) );
  XOR2_X1 U10789 ( .A(n10048), .B(n10850), .Z(n10041) );
  XOR2_X1 U10790 ( .A(n10047), .B(n10046), .Z(n10850) );
  OR2_X1 U10791 ( .A1(n7785), .A2(n7877), .ZN(n10046) );
  OR2_X1 U10792 ( .A1(n10851), .A2(n10852), .ZN(n10047) );
  AND2_X1 U10793 ( .A1(n10849), .A2(n10848), .ZN(n10852) );
  AND2_X1 U10794 ( .A1(n10846), .A2(n10853), .ZN(n10851) );
  OR2_X1 U10795 ( .A1(n10849), .A2(n10848), .ZN(n10853) );
  OR2_X1 U10796 ( .A1(n10854), .A2(n10855), .ZN(n10848) );
  AND2_X1 U10797 ( .A1(n10845), .A2(n10844), .ZN(n10855) );
  AND2_X1 U10798 ( .A1(n10842), .A2(n10856), .ZN(n10854) );
  OR2_X1 U10799 ( .A1(n10845), .A2(n10844), .ZN(n10856) );
  OR2_X1 U10800 ( .A1(n10857), .A2(n10858), .ZN(n10844) );
  AND2_X1 U10801 ( .A1(n10841), .A2(n10840), .ZN(n10858) );
  AND2_X1 U10802 ( .A1(n10838), .A2(n10859), .ZN(n10857) );
  OR2_X1 U10803 ( .A1(n10841), .A2(n10840), .ZN(n10859) );
  OR2_X1 U10804 ( .A1(n10860), .A2(n10861), .ZN(n10840) );
  AND2_X1 U10805 ( .A1(n10837), .A2(n10836), .ZN(n10861) );
  AND2_X1 U10806 ( .A1(n10834), .A2(n10862), .ZN(n10860) );
  OR2_X1 U10807 ( .A1(n10837), .A2(n10836), .ZN(n10862) );
  OR2_X1 U10808 ( .A1(n10863), .A2(n10864), .ZN(n10836) );
  AND2_X1 U10809 ( .A1(n10833), .A2(n10832), .ZN(n10864) );
  AND2_X1 U10810 ( .A1(n10830), .A2(n10865), .ZN(n10863) );
  OR2_X1 U10811 ( .A1(n10833), .A2(n10832), .ZN(n10865) );
  OR2_X1 U10812 ( .A1(n10866), .A2(n10867), .ZN(n10832) );
  AND2_X1 U10813 ( .A1(n10829), .A2(n10828), .ZN(n10867) );
  AND2_X1 U10814 ( .A1(n10826), .A2(n10868), .ZN(n10866) );
  OR2_X1 U10815 ( .A1(n10829), .A2(n10828), .ZN(n10868) );
  OR2_X1 U10816 ( .A1(n10869), .A2(n10870), .ZN(n10828) );
  AND2_X1 U10817 ( .A1(n10825), .A2(n10824), .ZN(n10870) );
  AND2_X1 U10818 ( .A1(n10822), .A2(n10871), .ZN(n10869) );
  OR2_X1 U10819 ( .A1(n10825), .A2(n10824), .ZN(n10871) );
  OR2_X1 U10820 ( .A1(n10872), .A2(n10873), .ZN(n10824) );
  AND2_X1 U10821 ( .A1(n10821), .A2(n10820), .ZN(n10873) );
  AND2_X1 U10822 ( .A1(n10818), .A2(n10874), .ZN(n10872) );
  OR2_X1 U10823 ( .A1(n10821), .A2(n10820), .ZN(n10874) );
  OR2_X1 U10824 ( .A1(n10875), .A2(n10876), .ZN(n10820) );
  AND2_X1 U10825 ( .A1(n10817), .A2(n10816), .ZN(n10876) );
  AND2_X1 U10826 ( .A1(n10814), .A2(n10877), .ZN(n10875) );
  OR2_X1 U10827 ( .A1(n10817), .A2(n10816), .ZN(n10877) );
  OR2_X1 U10828 ( .A1(n10878), .A2(n10879), .ZN(n10816) );
  AND2_X1 U10829 ( .A1(n10813), .A2(n10812), .ZN(n10879) );
  AND2_X1 U10830 ( .A1(n10810), .A2(n10880), .ZN(n10878) );
  OR2_X1 U10831 ( .A1(n10813), .A2(n10812), .ZN(n10880) );
  OR2_X1 U10832 ( .A1(n10881), .A2(n10882), .ZN(n10812) );
  AND2_X1 U10833 ( .A1(n10809), .A2(n10808), .ZN(n10882) );
  AND2_X1 U10834 ( .A1(n10806), .A2(n10883), .ZN(n10881) );
  OR2_X1 U10835 ( .A1(n10809), .A2(n10808), .ZN(n10883) );
  OR2_X1 U10836 ( .A1(n10884), .A2(n10885), .ZN(n10808) );
  AND2_X1 U10837 ( .A1(n10805), .A2(n10804), .ZN(n10885) );
  AND2_X1 U10838 ( .A1(n10802), .A2(n10886), .ZN(n10884) );
  OR2_X1 U10839 ( .A1(n10805), .A2(n10804), .ZN(n10886) );
  OR2_X1 U10840 ( .A1(n10887), .A2(n10888), .ZN(n10804) );
  AND2_X1 U10841 ( .A1(n10801), .A2(n10800), .ZN(n10888) );
  AND2_X1 U10842 ( .A1(n10798), .A2(n10889), .ZN(n10887) );
  OR2_X1 U10843 ( .A1(n10801), .A2(n10800), .ZN(n10889) );
  OR2_X1 U10844 ( .A1(n10890), .A2(n10891), .ZN(n10800) );
  AND2_X1 U10845 ( .A1(n10795), .A2(n10797), .ZN(n10891) );
  AND2_X1 U10846 ( .A1(n10892), .A2(n10796), .ZN(n10890) );
  OR2_X1 U10847 ( .A1(n10795), .A2(n10797), .ZN(n10892) );
  OR2_X1 U10848 ( .A1(n10893), .A2(n10894), .ZN(n10797) );
  AND2_X1 U10849 ( .A1(n10793), .A2(n10792), .ZN(n10894) );
  AND2_X1 U10850 ( .A1(n10790), .A2(n10895), .ZN(n10893) );
  OR2_X1 U10851 ( .A1(n10793), .A2(n10792), .ZN(n10895) );
  OR2_X1 U10852 ( .A1(n10896), .A2(n10897), .ZN(n10792) );
  AND2_X1 U10853 ( .A1(n10789), .A2(n10788), .ZN(n10897) );
  AND2_X1 U10854 ( .A1(n10786), .A2(n10898), .ZN(n10896) );
  OR2_X1 U10855 ( .A1(n10789), .A2(n10788), .ZN(n10898) );
  OR2_X1 U10856 ( .A1(n10899), .A2(n10900), .ZN(n10788) );
  AND2_X1 U10857 ( .A1(n10785), .A2(n10784), .ZN(n10900) );
  AND2_X1 U10858 ( .A1(n10782), .A2(n10901), .ZN(n10899) );
  OR2_X1 U10859 ( .A1(n10785), .A2(n10784), .ZN(n10901) );
  OR2_X1 U10860 ( .A1(n10902), .A2(n10903), .ZN(n10784) );
  AND2_X1 U10861 ( .A1(n10781), .A2(n10780), .ZN(n10903) );
  AND2_X1 U10862 ( .A1(n10778), .A2(n10904), .ZN(n10902) );
  OR2_X1 U10863 ( .A1(n10781), .A2(n10780), .ZN(n10904) );
  OR2_X1 U10864 ( .A1(n10905), .A2(n10906), .ZN(n10780) );
  AND2_X1 U10865 ( .A1(n10777), .A2(n10776), .ZN(n10906) );
  AND2_X1 U10866 ( .A1(n10774), .A2(n10907), .ZN(n10905) );
  OR2_X1 U10867 ( .A1(n10777), .A2(n10776), .ZN(n10907) );
  OR2_X1 U10868 ( .A1(n10908), .A2(n10909), .ZN(n10776) );
  AND2_X1 U10869 ( .A1(n10773), .A2(n10772), .ZN(n10909) );
  AND2_X1 U10870 ( .A1(n10770), .A2(n10910), .ZN(n10908) );
  OR2_X1 U10871 ( .A1(n10773), .A2(n10772), .ZN(n10910) );
  OR2_X1 U10872 ( .A1(n10911), .A2(n10912), .ZN(n10772) );
  AND2_X1 U10873 ( .A1(n10769), .A2(n10768), .ZN(n10912) );
  AND2_X1 U10874 ( .A1(n10766), .A2(n10913), .ZN(n10911) );
  OR2_X1 U10875 ( .A1(n10769), .A2(n10768), .ZN(n10913) );
  OR2_X1 U10876 ( .A1(n10914), .A2(n10915), .ZN(n10768) );
  AND2_X1 U10877 ( .A1(n10765), .A2(n10764), .ZN(n10915) );
  AND2_X1 U10878 ( .A1(n10762), .A2(n10916), .ZN(n10914) );
  OR2_X1 U10879 ( .A1(n10765), .A2(n10764), .ZN(n10916) );
  OR2_X1 U10880 ( .A1(n10917), .A2(n10918), .ZN(n10764) );
  AND2_X1 U10881 ( .A1(n10761), .A2(n10760), .ZN(n10918) );
  AND2_X1 U10882 ( .A1(n10758), .A2(n10919), .ZN(n10917) );
  OR2_X1 U10883 ( .A1(n10761), .A2(n10760), .ZN(n10919) );
  OR2_X1 U10884 ( .A1(n10920), .A2(n10921), .ZN(n10760) );
  AND2_X1 U10885 ( .A1(n10757), .A2(n10756), .ZN(n10921) );
  AND2_X1 U10886 ( .A1(n10754), .A2(n10922), .ZN(n10920) );
  OR2_X1 U10887 ( .A1(n10757), .A2(n10756), .ZN(n10922) );
  OR2_X1 U10888 ( .A1(n10923), .A2(n10924), .ZN(n10756) );
  AND2_X1 U10889 ( .A1(n10750), .A2(n10753), .ZN(n10924) );
  AND2_X1 U10890 ( .A1(n10752), .A2(n10925), .ZN(n10923) );
  OR2_X1 U10891 ( .A1(n10750), .A2(n10753), .ZN(n10925) );
  OR3_X1 U10892 ( .A1(n7852), .A2(n8349), .A3(n7877), .ZN(n10753) );
  OR2_X1 U10893 ( .A1(n8102), .A2(n7877), .ZN(n10750) );
  INV_X1 U10894 ( .A(n10926), .ZN(n10752) );
  OR2_X1 U10895 ( .A1(n10927), .A2(n10928), .ZN(n10926) );
  AND2_X1 U10896 ( .A1(b_17_), .A2(n10929), .ZN(n10928) );
  OR2_X1 U10897 ( .A1(n10930), .A2(n7314), .ZN(n10929) );
  AND2_X1 U10898 ( .A1(a_30_), .A2(n10931), .ZN(n10930) );
  AND2_X1 U10899 ( .A1(b_16_), .A2(n10932), .ZN(n10927) );
  OR2_X1 U10900 ( .A1(n10933), .A2(n7318), .ZN(n10932) );
  AND2_X1 U10901 ( .A1(a_31_), .A2(n7852), .ZN(n10933) );
  OR2_X1 U10902 ( .A1(n8111), .A2(n7877), .ZN(n10757) );
  XNOR2_X1 U10903 ( .A(n10934), .B(n10935), .ZN(n10754) );
  XNOR2_X1 U10904 ( .A(n10936), .B(n10937), .ZN(n10935) );
  OR2_X1 U10905 ( .A1(n8116), .A2(n7877), .ZN(n10761) );
  XOR2_X1 U10906 ( .A(n10938), .B(n10939), .Z(n10758) );
  XOR2_X1 U10907 ( .A(n10940), .B(n10941), .Z(n10939) );
  OR2_X1 U10908 ( .A1(n8121), .A2(n7877), .ZN(n10765) );
  XOR2_X1 U10909 ( .A(n10942), .B(n10943), .Z(n10762) );
  XOR2_X1 U10910 ( .A(n10944), .B(n10945), .Z(n10943) );
  OR2_X1 U10911 ( .A1(n8126), .A2(n7877), .ZN(n10769) );
  XOR2_X1 U10912 ( .A(n10946), .B(n10947), .Z(n10766) );
  XOR2_X1 U10913 ( .A(n10948), .B(n10949), .Z(n10947) );
  OR2_X1 U10914 ( .A1(n8131), .A2(n7877), .ZN(n10773) );
  XOR2_X1 U10915 ( .A(n10950), .B(n10951), .Z(n10770) );
  XOR2_X1 U10916 ( .A(n10952), .B(n10953), .Z(n10951) );
  OR2_X1 U10917 ( .A1(n8136), .A2(n7877), .ZN(n10777) );
  XOR2_X1 U10918 ( .A(n10954), .B(n10955), .Z(n10774) );
  XOR2_X1 U10919 ( .A(n10956), .B(n10957), .Z(n10955) );
  OR2_X1 U10920 ( .A1(n8141), .A2(n7877), .ZN(n10781) );
  XOR2_X1 U10921 ( .A(n10958), .B(n10959), .Z(n10778) );
  XOR2_X1 U10922 ( .A(n10960), .B(n10961), .Z(n10959) );
  OR2_X1 U10923 ( .A1(n8146), .A2(n7877), .ZN(n10785) );
  XOR2_X1 U10924 ( .A(n10962), .B(n10963), .Z(n10782) );
  XOR2_X1 U10925 ( .A(n10964), .B(n10965), .Z(n10963) );
  OR2_X1 U10926 ( .A1(n8151), .A2(n7877), .ZN(n10789) );
  XOR2_X1 U10927 ( .A(n10966), .B(n10967), .Z(n10786) );
  XOR2_X1 U10928 ( .A(n10968), .B(n10969), .Z(n10967) );
  OR2_X1 U10929 ( .A1(n8156), .A2(n7877), .ZN(n10793) );
  XOR2_X1 U10930 ( .A(n10970), .B(n10971), .Z(n10790) );
  XOR2_X1 U10931 ( .A(n10972), .B(n10973), .Z(n10971) );
  XOR2_X1 U10932 ( .A(n10974), .B(n10975), .Z(n10795) );
  XOR2_X1 U10933 ( .A(n10976), .B(n10977), .Z(n10975) );
  OR2_X1 U10934 ( .A1(n8166), .A2(n7877), .ZN(n10801) );
  XOR2_X1 U10935 ( .A(n10978), .B(n10979), .Z(n10798) );
  XOR2_X1 U10936 ( .A(n10980), .B(n10981), .Z(n10979) );
  OR2_X1 U10937 ( .A1(n8171), .A2(n7877), .ZN(n10805) );
  XNOR2_X1 U10938 ( .A(n10982), .B(n10983), .ZN(n10802) );
  XNOR2_X1 U10939 ( .A(n10984), .B(n10985), .ZN(n10982) );
  OR2_X1 U10940 ( .A1(n8176), .A2(n7877), .ZN(n10809) );
  XOR2_X1 U10941 ( .A(n10986), .B(n10987), .Z(n10806) );
  XOR2_X1 U10942 ( .A(n10988), .B(n10989), .Z(n10987) );
  OR2_X1 U10943 ( .A1(n8181), .A2(n7877), .ZN(n10813) );
  XOR2_X1 U10944 ( .A(n10990), .B(n10991), .Z(n10810) );
  XOR2_X1 U10945 ( .A(n10992), .B(n10993), .Z(n10991) );
  OR2_X1 U10946 ( .A1(n8186), .A2(n7877), .ZN(n10817) );
  XOR2_X1 U10947 ( .A(n10994), .B(n10995), .Z(n10814) );
  XOR2_X1 U10948 ( .A(n10996), .B(n10997), .Z(n10995) );
  OR2_X1 U10949 ( .A1(n8191), .A2(n7877), .ZN(n10821) );
  XOR2_X1 U10950 ( .A(n10998), .B(n10999), .Z(n10818) );
  XOR2_X1 U10951 ( .A(n11000), .B(n11001), .Z(n10999) );
  OR2_X1 U10952 ( .A1(n8196), .A2(n7877), .ZN(n10825) );
  XOR2_X1 U10953 ( .A(n11002), .B(n11003), .Z(n10822) );
  XOR2_X1 U10954 ( .A(n11004), .B(n11005), .Z(n11003) );
  OR2_X1 U10955 ( .A1(n8201), .A2(n7877), .ZN(n10829) );
  XOR2_X1 U10956 ( .A(n11006), .B(n11007), .Z(n10826) );
  XOR2_X1 U10957 ( .A(n11008), .B(n11009), .Z(n11007) );
  OR2_X1 U10958 ( .A1(n8206), .A2(n7877), .ZN(n10833) );
  XOR2_X1 U10959 ( .A(n11010), .B(n11011), .Z(n10830) );
  XOR2_X1 U10960 ( .A(n11012), .B(n11013), .Z(n11011) );
  OR2_X1 U10961 ( .A1(n8211), .A2(n7877), .ZN(n10837) );
  XOR2_X1 U10962 ( .A(n11014), .B(n11015), .Z(n10834) );
  XOR2_X1 U10963 ( .A(n11016), .B(n11017), .Z(n11015) );
  OR2_X1 U10964 ( .A1(n8216), .A2(n7877), .ZN(n10841) );
  XOR2_X1 U10965 ( .A(n11018), .B(n11019), .Z(n10838) );
  XOR2_X1 U10966 ( .A(n11020), .B(n11021), .Z(n11019) );
  OR2_X1 U10967 ( .A1(n8221), .A2(n7877), .ZN(n10845) );
  XOR2_X1 U10968 ( .A(n11022), .B(n11023), .Z(n10842) );
  XOR2_X1 U10969 ( .A(n11024), .B(n11025), .Z(n11023) );
  OR2_X1 U10970 ( .A1(n8226), .A2(n7877), .ZN(n10849) );
  XOR2_X1 U10971 ( .A(n11026), .B(n11027), .Z(n10846) );
  XOR2_X1 U10972 ( .A(n11028), .B(n11029), .Z(n11027) );
  XOR2_X1 U10973 ( .A(n10055), .B(n11030), .Z(n10048) );
  XOR2_X1 U10974 ( .A(n10054), .B(n10053), .Z(n11030) );
  OR2_X1 U10975 ( .A1(n7852), .A2(n8226), .ZN(n10053) );
  OR2_X1 U10976 ( .A1(n11031), .A2(n11032), .ZN(n10054) );
  AND2_X1 U10977 ( .A1(n11029), .A2(n11028), .ZN(n11032) );
  AND2_X1 U10978 ( .A1(n11026), .A2(n11033), .ZN(n11031) );
  OR2_X1 U10979 ( .A1(n11029), .A2(n11028), .ZN(n11033) );
  OR2_X1 U10980 ( .A1(n11034), .A2(n11035), .ZN(n11028) );
  AND2_X1 U10981 ( .A1(n11025), .A2(n11024), .ZN(n11035) );
  AND2_X1 U10982 ( .A1(n11022), .A2(n11036), .ZN(n11034) );
  OR2_X1 U10983 ( .A1(n11025), .A2(n11024), .ZN(n11036) );
  OR2_X1 U10984 ( .A1(n11037), .A2(n11038), .ZN(n11024) );
  AND2_X1 U10985 ( .A1(n11021), .A2(n11020), .ZN(n11038) );
  AND2_X1 U10986 ( .A1(n11018), .A2(n11039), .ZN(n11037) );
  OR2_X1 U10987 ( .A1(n11021), .A2(n11020), .ZN(n11039) );
  OR2_X1 U10988 ( .A1(n11040), .A2(n11041), .ZN(n11020) );
  AND2_X1 U10989 ( .A1(n11017), .A2(n11016), .ZN(n11041) );
  AND2_X1 U10990 ( .A1(n11014), .A2(n11042), .ZN(n11040) );
  OR2_X1 U10991 ( .A1(n11017), .A2(n11016), .ZN(n11042) );
  OR2_X1 U10992 ( .A1(n11043), .A2(n11044), .ZN(n11016) );
  AND2_X1 U10993 ( .A1(n11013), .A2(n11012), .ZN(n11044) );
  AND2_X1 U10994 ( .A1(n11010), .A2(n11045), .ZN(n11043) );
  OR2_X1 U10995 ( .A1(n11013), .A2(n11012), .ZN(n11045) );
  OR2_X1 U10996 ( .A1(n11046), .A2(n11047), .ZN(n11012) );
  AND2_X1 U10997 ( .A1(n11009), .A2(n11008), .ZN(n11047) );
  AND2_X1 U10998 ( .A1(n11006), .A2(n11048), .ZN(n11046) );
  OR2_X1 U10999 ( .A1(n11009), .A2(n11008), .ZN(n11048) );
  OR2_X1 U11000 ( .A1(n11049), .A2(n11050), .ZN(n11008) );
  AND2_X1 U11001 ( .A1(n11005), .A2(n11004), .ZN(n11050) );
  AND2_X1 U11002 ( .A1(n11002), .A2(n11051), .ZN(n11049) );
  OR2_X1 U11003 ( .A1(n11005), .A2(n11004), .ZN(n11051) );
  OR2_X1 U11004 ( .A1(n11052), .A2(n11053), .ZN(n11004) );
  AND2_X1 U11005 ( .A1(n11001), .A2(n11000), .ZN(n11053) );
  AND2_X1 U11006 ( .A1(n10998), .A2(n11054), .ZN(n11052) );
  OR2_X1 U11007 ( .A1(n11001), .A2(n11000), .ZN(n11054) );
  OR2_X1 U11008 ( .A1(n11055), .A2(n11056), .ZN(n11000) );
  AND2_X1 U11009 ( .A1(n10997), .A2(n10996), .ZN(n11056) );
  AND2_X1 U11010 ( .A1(n10994), .A2(n11057), .ZN(n11055) );
  OR2_X1 U11011 ( .A1(n10997), .A2(n10996), .ZN(n11057) );
  OR2_X1 U11012 ( .A1(n11058), .A2(n11059), .ZN(n10996) );
  AND2_X1 U11013 ( .A1(n10993), .A2(n10992), .ZN(n11059) );
  AND2_X1 U11014 ( .A1(n10990), .A2(n11060), .ZN(n11058) );
  OR2_X1 U11015 ( .A1(n10993), .A2(n10992), .ZN(n11060) );
  OR2_X1 U11016 ( .A1(n11061), .A2(n11062), .ZN(n10992) );
  AND2_X1 U11017 ( .A1(n10989), .A2(n10988), .ZN(n11062) );
  AND2_X1 U11018 ( .A1(n10986), .A2(n11063), .ZN(n11061) );
  OR2_X1 U11019 ( .A1(n10989), .A2(n10988), .ZN(n11063) );
  OR2_X1 U11020 ( .A1(n11064), .A2(n11065), .ZN(n10988) );
  AND2_X1 U11021 ( .A1(n10983), .A2(n10985), .ZN(n11065) );
  AND2_X1 U11022 ( .A1(n11066), .A2(n10984), .ZN(n11064) );
  OR2_X1 U11023 ( .A1(n10983), .A2(n10985), .ZN(n11066) );
  OR2_X1 U11024 ( .A1(n11067), .A2(n11068), .ZN(n10985) );
  AND2_X1 U11025 ( .A1(n10981), .A2(n10980), .ZN(n11068) );
  AND2_X1 U11026 ( .A1(n10978), .A2(n11069), .ZN(n11067) );
  OR2_X1 U11027 ( .A1(n10981), .A2(n10980), .ZN(n11069) );
  OR2_X1 U11028 ( .A1(n11070), .A2(n11071), .ZN(n10980) );
  AND2_X1 U11029 ( .A1(n10977), .A2(n10976), .ZN(n11071) );
  AND2_X1 U11030 ( .A1(n10974), .A2(n11072), .ZN(n11070) );
  OR2_X1 U11031 ( .A1(n10977), .A2(n10976), .ZN(n11072) );
  OR2_X1 U11032 ( .A1(n11073), .A2(n11074), .ZN(n10976) );
  AND2_X1 U11033 ( .A1(n10973), .A2(n10972), .ZN(n11074) );
  AND2_X1 U11034 ( .A1(n10970), .A2(n11075), .ZN(n11073) );
  OR2_X1 U11035 ( .A1(n10973), .A2(n10972), .ZN(n11075) );
  OR2_X1 U11036 ( .A1(n11076), .A2(n11077), .ZN(n10972) );
  AND2_X1 U11037 ( .A1(n10969), .A2(n10968), .ZN(n11077) );
  AND2_X1 U11038 ( .A1(n10966), .A2(n11078), .ZN(n11076) );
  OR2_X1 U11039 ( .A1(n10969), .A2(n10968), .ZN(n11078) );
  OR2_X1 U11040 ( .A1(n11079), .A2(n11080), .ZN(n10968) );
  AND2_X1 U11041 ( .A1(n10965), .A2(n10964), .ZN(n11080) );
  AND2_X1 U11042 ( .A1(n10962), .A2(n11081), .ZN(n11079) );
  OR2_X1 U11043 ( .A1(n10965), .A2(n10964), .ZN(n11081) );
  OR2_X1 U11044 ( .A1(n11082), .A2(n11083), .ZN(n10964) );
  AND2_X1 U11045 ( .A1(n10961), .A2(n10960), .ZN(n11083) );
  AND2_X1 U11046 ( .A1(n10958), .A2(n11084), .ZN(n11082) );
  OR2_X1 U11047 ( .A1(n10961), .A2(n10960), .ZN(n11084) );
  OR2_X1 U11048 ( .A1(n11085), .A2(n11086), .ZN(n10960) );
  AND2_X1 U11049 ( .A1(n10957), .A2(n10956), .ZN(n11086) );
  AND2_X1 U11050 ( .A1(n10954), .A2(n11087), .ZN(n11085) );
  OR2_X1 U11051 ( .A1(n10957), .A2(n10956), .ZN(n11087) );
  OR2_X1 U11052 ( .A1(n11088), .A2(n11089), .ZN(n10956) );
  AND2_X1 U11053 ( .A1(n10953), .A2(n10952), .ZN(n11089) );
  AND2_X1 U11054 ( .A1(n10950), .A2(n11090), .ZN(n11088) );
  OR2_X1 U11055 ( .A1(n10953), .A2(n10952), .ZN(n11090) );
  OR2_X1 U11056 ( .A1(n11091), .A2(n11092), .ZN(n10952) );
  AND2_X1 U11057 ( .A1(n10949), .A2(n10948), .ZN(n11092) );
  AND2_X1 U11058 ( .A1(n10946), .A2(n11093), .ZN(n11091) );
  OR2_X1 U11059 ( .A1(n10949), .A2(n10948), .ZN(n11093) );
  OR2_X1 U11060 ( .A1(n11094), .A2(n11095), .ZN(n10948) );
  AND2_X1 U11061 ( .A1(n10945), .A2(n10944), .ZN(n11095) );
  AND2_X1 U11062 ( .A1(n10942), .A2(n11096), .ZN(n11094) );
  OR2_X1 U11063 ( .A1(n10945), .A2(n10944), .ZN(n11096) );
  OR2_X1 U11064 ( .A1(n11097), .A2(n11098), .ZN(n10944) );
  AND2_X1 U11065 ( .A1(n10941), .A2(n10940), .ZN(n11098) );
  AND2_X1 U11066 ( .A1(n10938), .A2(n11099), .ZN(n11097) );
  OR2_X1 U11067 ( .A1(n10941), .A2(n10940), .ZN(n11099) );
  OR2_X1 U11068 ( .A1(n11100), .A2(n11101), .ZN(n10940) );
  AND2_X1 U11069 ( .A1(n10934), .A2(n10937), .ZN(n11101) );
  AND2_X1 U11070 ( .A1(n10936), .A2(n11102), .ZN(n11100) );
  OR2_X1 U11071 ( .A1(n10934), .A2(n10937), .ZN(n11102) );
  OR3_X1 U11072 ( .A1(n7852), .A2(n10931), .A3(n8349), .ZN(n10937) );
  OR2_X1 U11073 ( .A1(n7852), .A2(n8102), .ZN(n10934) );
  INV_X1 U11074 ( .A(n11103), .ZN(n10936) );
  OR2_X1 U11075 ( .A1(n11104), .A2(n11105), .ZN(n11103) );
  AND2_X1 U11076 ( .A1(b_16_), .A2(n11106), .ZN(n11105) );
  OR2_X1 U11077 ( .A1(n11107), .A2(n7314), .ZN(n11106) );
  AND2_X1 U11078 ( .A1(a_30_), .A2(n11108), .ZN(n11107) );
  AND2_X1 U11079 ( .A1(b_15_), .A2(n11109), .ZN(n11104) );
  OR2_X1 U11080 ( .A1(n11110), .A2(n7318), .ZN(n11109) );
  AND2_X1 U11081 ( .A1(a_31_), .A2(n10931), .ZN(n11110) );
  OR2_X1 U11082 ( .A1(n7852), .A2(n8111), .ZN(n10941) );
  XNOR2_X1 U11083 ( .A(n11111), .B(n11112), .ZN(n10938) );
  XNOR2_X1 U11084 ( .A(n11113), .B(n11114), .ZN(n11112) );
  OR2_X1 U11085 ( .A1(n7852), .A2(n8116), .ZN(n10945) );
  XOR2_X1 U11086 ( .A(n11115), .B(n11116), .Z(n10942) );
  XOR2_X1 U11087 ( .A(n11117), .B(n11118), .Z(n11116) );
  OR2_X1 U11088 ( .A1(n7852), .A2(n8121), .ZN(n10949) );
  XOR2_X1 U11089 ( .A(n11119), .B(n11120), .Z(n10946) );
  XOR2_X1 U11090 ( .A(n11121), .B(n11122), .Z(n11120) );
  OR2_X1 U11091 ( .A1(n7852), .A2(n8126), .ZN(n10953) );
  XOR2_X1 U11092 ( .A(n11123), .B(n11124), .Z(n10950) );
  XOR2_X1 U11093 ( .A(n11125), .B(n11126), .Z(n11124) );
  OR2_X1 U11094 ( .A1(n7852), .A2(n8131), .ZN(n10957) );
  XOR2_X1 U11095 ( .A(n11127), .B(n11128), .Z(n10954) );
  XOR2_X1 U11096 ( .A(n11129), .B(n11130), .Z(n11128) );
  OR2_X1 U11097 ( .A1(n7852), .A2(n8136), .ZN(n10961) );
  XOR2_X1 U11098 ( .A(n11131), .B(n11132), .Z(n10958) );
  XOR2_X1 U11099 ( .A(n11133), .B(n11134), .Z(n11132) );
  OR2_X1 U11100 ( .A1(n7852), .A2(n8141), .ZN(n10965) );
  XOR2_X1 U11101 ( .A(n11135), .B(n11136), .Z(n10962) );
  XOR2_X1 U11102 ( .A(n11137), .B(n11138), .Z(n11136) );
  OR2_X1 U11103 ( .A1(n7852), .A2(n8146), .ZN(n10969) );
  XOR2_X1 U11104 ( .A(n11139), .B(n11140), .Z(n10966) );
  XOR2_X1 U11105 ( .A(n11141), .B(n11142), .Z(n11140) );
  OR2_X1 U11106 ( .A1(n7852), .A2(n8151), .ZN(n10973) );
  XOR2_X1 U11107 ( .A(n11143), .B(n11144), .Z(n10970) );
  XOR2_X1 U11108 ( .A(n11145), .B(n11146), .Z(n11144) );
  OR2_X1 U11109 ( .A1(n7852), .A2(n8156), .ZN(n10977) );
  XOR2_X1 U11110 ( .A(n11147), .B(n11148), .Z(n10974) );
  XOR2_X1 U11111 ( .A(n11149), .B(n11150), .Z(n11148) );
  OR2_X1 U11112 ( .A1(n7852), .A2(n8161), .ZN(n10981) );
  XOR2_X1 U11113 ( .A(n11151), .B(n11152), .Z(n10978) );
  XOR2_X1 U11114 ( .A(n11153), .B(n11154), .Z(n11152) );
  XOR2_X1 U11115 ( .A(n11155), .B(n11156), .Z(n10983) );
  XOR2_X1 U11116 ( .A(n11157), .B(n11158), .Z(n11156) );
  OR2_X1 U11117 ( .A1(n7852), .A2(n8171), .ZN(n10989) );
  XOR2_X1 U11118 ( .A(n11159), .B(n11160), .Z(n10986) );
  XOR2_X1 U11119 ( .A(n11161), .B(n11162), .Z(n11160) );
  OR2_X1 U11120 ( .A1(n7852), .A2(n8176), .ZN(n10993) );
  XNOR2_X1 U11121 ( .A(n11163), .B(n11164), .ZN(n10990) );
  XNOR2_X1 U11122 ( .A(n11165), .B(n11166), .ZN(n11163) );
  OR2_X1 U11123 ( .A1(n7852), .A2(n8181), .ZN(n10997) );
  XOR2_X1 U11124 ( .A(n11167), .B(n11168), .Z(n10994) );
  XOR2_X1 U11125 ( .A(n11169), .B(n11170), .Z(n11168) );
  OR2_X1 U11126 ( .A1(n7852), .A2(n8186), .ZN(n11001) );
  XOR2_X1 U11127 ( .A(n11171), .B(n11172), .Z(n10998) );
  XOR2_X1 U11128 ( .A(n11173), .B(n11174), .Z(n11172) );
  OR2_X1 U11129 ( .A1(n7852), .A2(n8191), .ZN(n11005) );
  XOR2_X1 U11130 ( .A(n11175), .B(n11176), .Z(n11002) );
  XOR2_X1 U11131 ( .A(n11177), .B(n11178), .Z(n11176) );
  OR2_X1 U11132 ( .A1(n7852), .A2(n8196), .ZN(n11009) );
  XOR2_X1 U11133 ( .A(n11179), .B(n11180), .Z(n11006) );
  XOR2_X1 U11134 ( .A(n11181), .B(n11182), .Z(n11180) );
  OR2_X1 U11135 ( .A1(n7852), .A2(n8201), .ZN(n11013) );
  XOR2_X1 U11136 ( .A(n11183), .B(n11184), .Z(n11010) );
  XOR2_X1 U11137 ( .A(n11185), .B(n11186), .Z(n11184) );
  OR2_X1 U11138 ( .A1(n7852), .A2(n8206), .ZN(n11017) );
  XOR2_X1 U11139 ( .A(n11187), .B(n11188), .Z(n11014) );
  XOR2_X1 U11140 ( .A(n11189), .B(n11190), .Z(n11188) );
  OR2_X1 U11141 ( .A1(n7852), .A2(n8211), .ZN(n11021) );
  XOR2_X1 U11142 ( .A(n11191), .B(n11192), .Z(n11018) );
  XOR2_X1 U11143 ( .A(n11193), .B(n11194), .Z(n11192) );
  OR2_X1 U11144 ( .A1(n7852), .A2(n8216), .ZN(n11025) );
  XOR2_X1 U11145 ( .A(n11195), .B(n11196), .Z(n11022) );
  XOR2_X1 U11146 ( .A(n11197), .B(n11198), .Z(n11196) );
  OR2_X1 U11147 ( .A1(n7852), .A2(n8221), .ZN(n11029) );
  XOR2_X1 U11148 ( .A(n11199), .B(n11200), .Z(n11026) );
  XOR2_X1 U11149 ( .A(n11201), .B(n11202), .Z(n11200) );
  XOR2_X1 U11150 ( .A(n11203), .B(n11204), .Z(n10055) );
  XOR2_X1 U11151 ( .A(n11205), .B(n11206), .Z(n11204) );
  OR2_X1 U11152 ( .A1(n11207), .A2(n7812), .ZN(n7541) );
  XNOR2_X1 U11153 ( .A(n7552), .B(n7809), .ZN(n7812) );
  OR2_X1 U11154 ( .A1(n11208), .A2(n11209), .ZN(n7809) );
  AND2_X1 U11155 ( .A1(n11210), .A2(n11211), .ZN(n11209) );
  AND2_X1 U11156 ( .A1(n11212), .A2(n11213), .ZN(n11208) );
  OR2_X1 U11157 ( .A1(n11211), .A2(n11210), .ZN(n11213) );
  XNOR2_X1 U11158 ( .A(n11214), .B(n11215), .ZN(n7552) );
  XOR2_X1 U11159 ( .A(n11216), .B(n11217), .Z(n11215) );
  AND2_X1 U11160 ( .A1(n7813), .A2(n7811), .ZN(n11207) );
  XNOR2_X1 U11161 ( .A(n11212), .B(n11218), .ZN(n7811) );
  XOR2_X1 U11162 ( .A(n11211), .B(n11210), .Z(n11218) );
  OR2_X1 U11163 ( .A1(n11108), .A2(n7621), .ZN(n11210) );
  OR2_X1 U11164 ( .A1(n11219), .A2(n11220), .ZN(n11211) );
  AND2_X1 U11165 ( .A1(n11221), .A2(n11222), .ZN(n11220) );
  AND2_X1 U11166 ( .A1(n11223), .A2(n11224), .ZN(n11219) );
  OR2_X1 U11167 ( .A1(n11222), .A2(n11221), .ZN(n11224) );
  XOR2_X1 U11168 ( .A(n11225), .B(n11226), .Z(n11212) );
  XOR2_X1 U11169 ( .A(n11227), .B(n11228), .Z(n11226) );
  INV_X1 U11170 ( .A(n11229), .ZN(n7813) );
  OR2_X1 U11171 ( .A1(n11230), .A2(n11231), .ZN(n11229) );
  AND2_X1 U11172 ( .A1(n7837), .A2(n7836), .ZN(n11231) );
  AND2_X1 U11173 ( .A1(n7834), .A2(n11232), .ZN(n11230) );
  OR2_X1 U11174 ( .A1(n7836), .A2(n7837), .ZN(n11232) );
  OR2_X1 U11175 ( .A1(n10931), .A2(n7621), .ZN(n7837) );
  OR2_X1 U11176 ( .A1(n11233), .A2(n11234), .ZN(n7836) );
  AND2_X1 U11177 ( .A1(n7862), .A2(n7861), .ZN(n11234) );
  AND2_X1 U11178 ( .A1(n7859), .A2(n11235), .ZN(n11233) );
  OR2_X1 U11179 ( .A1(n7861), .A2(n7862), .ZN(n11235) );
  OR2_X1 U11180 ( .A1(n10931), .A2(n7656), .ZN(n7862) );
  OR2_X1 U11181 ( .A1(n11236), .A2(n11237), .ZN(n7861) );
  AND2_X1 U11182 ( .A1(n7894), .A2(n7893), .ZN(n11237) );
  AND2_X1 U11183 ( .A1(n7891), .A2(n11238), .ZN(n11236) );
  OR2_X1 U11184 ( .A1(n7893), .A2(n7894), .ZN(n11238) );
  OR2_X1 U11185 ( .A1(n10931), .A2(n7689), .ZN(n7894) );
  OR2_X1 U11186 ( .A1(n11239), .A2(n11240), .ZN(n7893) );
  AND2_X1 U11187 ( .A1(n7933), .A2(n7932), .ZN(n11240) );
  AND2_X1 U11188 ( .A1(n7930), .A2(n11241), .ZN(n11239) );
  OR2_X1 U11189 ( .A1(n7932), .A2(n7933), .ZN(n11241) );
  OR2_X1 U11190 ( .A1(n10931), .A2(n7777), .ZN(n7933) );
  OR2_X1 U11191 ( .A1(n11242), .A2(n11243), .ZN(n7932) );
  AND2_X1 U11192 ( .A1(n10021), .A2(n10020), .ZN(n11243) );
  AND2_X1 U11193 ( .A1(n10018), .A2(n11244), .ZN(n11242) );
  OR2_X1 U11194 ( .A1(n10020), .A2(n10021), .ZN(n11244) );
  OR2_X1 U11195 ( .A1(n10931), .A2(n7785), .ZN(n10021) );
  OR2_X1 U11196 ( .A1(n11245), .A2(n11246), .ZN(n10020) );
  AND2_X1 U11197 ( .A1(n10060), .A2(n10059), .ZN(n11246) );
  AND2_X1 U11198 ( .A1(n10057), .A2(n11247), .ZN(n11245) );
  OR2_X1 U11199 ( .A1(n10059), .A2(n10060), .ZN(n11247) );
  OR2_X1 U11200 ( .A1(n10931), .A2(n8226), .ZN(n10060) );
  OR2_X1 U11201 ( .A1(n11248), .A2(n11249), .ZN(n10059) );
  AND2_X1 U11202 ( .A1(n11206), .A2(n11205), .ZN(n11249) );
  AND2_X1 U11203 ( .A1(n11203), .A2(n11250), .ZN(n11248) );
  OR2_X1 U11204 ( .A1(n11205), .A2(n11206), .ZN(n11250) );
  OR2_X1 U11205 ( .A1(n10931), .A2(n8221), .ZN(n11206) );
  OR2_X1 U11206 ( .A1(n11251), .A2(n11252), .ZN(n11205) );
  AND2_X1 U11207 ( .A1(n11202), .A2(n11201), .ZN(n11252) );
  AND2_X1 U11208 ( .A1(n11199), .A2(n11253), .ZN(n11251) );
  OR2_X1 U11209 ( .A1(n11201), .A2(n11202), .ZN(n11253) );
  OR2_X1 U11210 ( .A1(n10931), .A2(n8216), .ZN(n11202) );
  OR2_X1 U11211 ( .A1(n11254), .A2(n11255), .ZN(n11201) );
  AND2_X1 U11212 ( .A1(n11198), .A2(n11197), .ZN(n11255) );
  AND2_X1 U11213 ( .A1(n11195), .A2(n11256), .ZN(n11254) );
  OR2_X1 U11214 ( .A1(n11197), .A2(n11198), .ZN(n11256) );
  OR2_X1 U11215 ( .A1(n10931), .A2(n8211), .ZN(n11198) );
  OR2_X1 U11216 ( .A1(n11257), .A2(n11258), .ZN(n11197) );
  AND2_X1 U11217 ( .A1(n11194), .A2(n11193), .ZN(n11258) );
  AND2_X1 U11218 ( .A1(n11191), .A2(n11259), .ZN(n11257) );
  OR2_X1 U11219 ( .A1(n11193), .A2(n11194), .ZN(n11259) );
  OR2_X1 U11220 ( .A1(n10931), .A2(n8206), .ZN(n11194) );
  OR2_X1 U11221 ( .A1(n11260), .A2(n11261), .ZN(n11193) );
  AND2_X1 U11222 ( .A1(n11190), .A2(n11189), .ZN(n11261) );
  AND2_X1 U11223 ( .A1(n11187), .A2(n11262), .ZN(n11260) );
  OR2_X1 U11224 ( .A1(n11189), .A2(n11190), .ZN(n11262) );
  OR2_X1 U11225 ( .A1(n10931), .A2(n8201), .ZN(n11190) );
  OR2_X1 U11226 ( .A1(n11263), .A2(n11264), .ZN(n11189) );
  AND2_X1 U11227 ( .A1(n11186), .A2(n11185), .ZN(n11264) );
  AND2_X1 U11228 ( .A1(n11183), .A2(n11265), .ZN(n11263) );
  OR2_X1 U11229 ( .A1(n11185), .A2(n11186), .ZN(n11265) );
  OR2_X1 U11230 ( .A1(n10931), .A2(n8196), .ZN(n11186) );
  OR2_X1 U11231 ( .A1(n11266), .A2(n11267), .ZN(n11185) );
  AND2_X1 U11232 ( .A1(n11182), .A2(n11181), .ZN(n11267) );
  AND2_X1 U11233 ( .A1(n11179), .A2(n11268), .ZN(n11266) );
  OR2_X1 U11234 ( .A1(n11181), .A2(n11182), .ZN(n11268) );
  OR2_X1 U11235 ( .A1(n10931), .A2(n8191), .ZN(n11182) );
  OR2_X1 U11236 ( .A1(n11269), .A2(n11270), .ZN(n11181) );
  AND2_X1 U11237 ( .A1(n11178), .A2(n11177), .ZN(n11270) );
  AND2_X1 U11238 ( .A1(n11175), .A2(n11271), .ZN(n11269) );
  OR2_X1 U11239 ( .A1(n11177), .A2(n11178), .ZN(n11271) );
  OR2_X1 U11240 ( .A1(n10931), .A2(n8186), .ZN(n11178) );
  OR2_X1 U11241 ( .A1(n11272), .A2(n11273), .ZN(n11177) );
  AND2_X1 U11242 ( .A1(n11174), .A2(n11173), .ZN(n11273) );
  AND2_X1 U11243 ( .A1(n11171), .A2(n11274), .ZN(n11272) );
  OR2_X1 U11244 ( .A1(n11173), .A2(n11174), .ZN(n11274) );
  OR2_X1 U11245 ( .A1(n10931), .A2(n8181), .ZN(n11174) );
  OR2_X1 U11246 ( .A1(n11275), .A2(n11276), .ZN(n11173) );
  AND2_X1 U11247 ( .A1(n11170), .A2(n11169), .ZN(n11276) );
  AND2_X1 U11248 ( .A1(n11167), .A2(n11277), .ZN(n11275) );
  OR2_X1 U11249 ( .A1(n11169), .A2(n11170), .ZN(n11277) );
  OR2_X1 U11250 ( .A1(n10931), .A2(n8176), .ZN(n11170) );
  OR2_X1 U11251 ( .A1(n11278), .A2(n11279), .ZN(n11169) );
  AND2_X1 U11252 ( .A1(n11164), .A2(n11166), .ZN(n11279) );
  AND2_X1 U11253 ( .A1(n11280), .A2(n11165), .ZN(n11278) );
  OR2_X1 U11254 ( .A1(n11166), .A2(n11164), .ZN(n11280) );
  XOR2_X1 U11255 ( .A(n11281), .B(n11282), .Z(n11164) );
  XOR2_X1 U11256 ( .A(n11283), .B(n11284), .Z(n11282) );
  OR2_X1 U11257 ( .A1(n11285), .A2(n11286), .ZN(n11166) );
  AND2_X1 U11258 ( .A1(n11162), .A2(n11161), .ZN(n11286) );
  AND2_X1 U11259 ( .A1(n11159), .A2(n11287), .ZN(n11285) );
  OR2_X1 U11260 ( .A1(n11161), .A2(n11162), .ZN(n11287) );
  OR2_X1 U11261 ( .A1(n8166), .A2(n10931), .ZN(n11162) );
  OR2_X1 U11262 ( .A1(n11288), .A2(n11289), .ZN(n11161) );
  AND2_X1 U11263 ( .A1(n11158), .A2(n11157), .ZN(n11289) );
  AND2_X1 U11264 ( .A1(n11155), .A2(n11290), .ZN(n11288) );
  OR2_X1 U11265 ( .A1(n11157), .A2(n11158), .ZN(n11290) );
  OR2_X1 U11266 ( .A1(n10931), .A2(n8161), .ZN(n11158) );
  OR2_X1 U11267 ( .A1(n11291), .A2(n11292), .ZN(n11157) );
  AND2_X1 U11268 ( .A1(n11154), .A2(n11153), .ZN(n11292) );
  AND2_X1 U11269 ( .A1(n11151), .A2(n11293), .ZN(n11291) );
  OR2_X1 U11270 ( .A1(n11153), .A2(n11154), .ZN(n11293) );
  OR2_X1 U11271 ( .A1(n10931), .A2(n8156), .ZN(n11154) );
  OR2_X1 U11272 ( .A1(n11294), .A2(n11295), .ZN(n11153) );
  AND2_X1 U11273 ( .A1(n11150), .A2(n11149), .ZN(n11295) );
  AND2_X1 U11274 ( .A1(n11147), .A2(n11296), .ZN(n11294) );
  OR2_X1 U11275 ( .A1(n11149), .A2(n11150), .ZN(n11296) );
  OR2_X1 U11276 ( .A1(n10931), .A2(n8151), .ZN(n11150) );
  OR2_X1 U11277 ( .A1(n11297), .A2(n11298), .ZN(n11149) );
  AND2_X1 U11278 ( .A1(n11146), .A2(n11145), .ZN(n11298) );
  AND2_X1 U11279 ( .A1(n11143), .A2(n11299), .ZN(n11297) );
  OR2_X1 U11280 ( .A1(n11145), .A2(n11146), .ZN(n11299) );
  OR2_X1 U11281 ( .A1(n10931), .A2(n8146), .ZN(n11146) );
  OR2_X1 U11282 ( .A1(n11300), .A2(n11301), .ZN(n11145) );
  AND2_X1 U11283 ( .A1(n11142), .A2(n11141), .ZN(n11301) );
  AND2_X1 U11284 ( .A1(n11139), .A2(n11302), .ZN(n11300) );
  OR2_X1 U11285 ( .A1(n11141), .A2(n11142), .ZN(n11302) );
  OR2_X1 U11286 ( .A1(n10931), .A2(n8141), .ZN(n11142) );
  OR2_X1 U11287 ( .A1(n11303), .A2(n11304), .ZN(n11141) );
  AND2_X1 U11288 ( .A1(n11138), .A2(n11137), .ZN(n11304) );
  AND2_X1 U11289 ( .A1(n11135), .A2(n11305), .ZN(n11303) );
  OR2_X1 U11290 ( .A1(n11137), .A2(n11138), .ZN(n11305) );
  OR2_X1 U11291 ( .A1(n10931), .A2(n8136), .ZN(n11138) );
  OR2_X1 U11292 ( .A1(n11306), .A2(n11307), .ZN(n11137) );
  AND2_X1 U11293 ( .A1(n11134), .A2(n11133), .ZN(n11307) );
  AND2_X1 U11294 ( .A1(n11131), .A2(n11308), .ZN(n11306) );
  OR2_X1 U11295 ( .A1(n11133), .A2(n11134), .ZN(n11308) );
  OR2_X1 U11296 ( .A1(n10931), .A2(n8131), .ZN(n11134) );
  OR2_X1 U11297 ( .A1(n11309), .A2(n11310), .ZN(n11133) );
  AND2_X1 U11298 ( .A1(n11130), .A2(n11129), .ZN(n11310) );
  AND2_X1 U11299 ( .A1(n11127), .A2(n11311), .ZN(n11309) );
  OR2_X1 U11300 ( .A1(n11129), .A2(n11130), .ZN(n11311) );
  OR2_X1 U11301 ( .A1(n10931), .A2(n8126), .ZN(n11130) );
  OR2_X1 U11302 ( .A1(n11312), .A2(n11313), .ZN(n11129) );
  AND2_X1 U11303 ( .A1(n11126), .A2(n11125), .ZN(n11313) );
  AND2_X1 U11304 ( .A1(n11123), .A2(n11314), .ZN(n11312) );
  OR2_X1 U11305 ( .A1(n11125), .A2(n11126), .ZN(n11314) );
  OR2_X1 U11306 ( .A1(n10931), .A2(n8121), .ZN(n11126) );
  OR2_X1 U11307 ( .A1(n11315), .A2(n11316), .ZN(n11125) );
  AND2_X1 U11308 ( .A1(n11122), .A2(n11121), .ZN(n11316) );
  AND2_X1 U11309 ( .A1(n11119), .A2(n11317), .ZN(n11315) );
  OR2_X1 U11310 ( .A1(n11121), .A2(n11122), .ZN(n11317) );
  OR2_X1 U11311 ( .A1(n10931), .A2(n8116), .ZN(n11122) );
  OR2_X1 U11312 ( .A1(n11318), .A2(n11319), .ZN(n11121) );
  AND2_X1 U11313 ( .A1(n11118), .A2(n11117), .ZN(n11319) );
  AND2_X1 U11314 ( .A1(n11115), .A2(n11320), .ZN(n11318) );
  OR2_X1 U11315 ( .A1(n11117), .A2(n11118), .ZN(n11320) );
  OR2_X1 U11316 ( .A1(n10931), .A2(n8111), .ZN(n11118) );
  OR2_X1 U11317 ( .A1(n11321), .A2(n11322), .ZN(n11117) );
  AND2_X1 U11318 ( .A1(n11111), .A2(n11114), .ZN(n11322) );
  AND2_X1 U11319 ( .A1(n11113), .A2(n11323), .ZN(n11321) );
  OR2_X1 U11320 ( .A1(n11114), .A2(n11111), .ZN(n11323) );
  OR2_X1 U11321 ( .A1(n10931), .A2(n8102), .ZN(n11111) );
  OR3_X1 U11322 ( .A1(n11108), .A2(n10931), .A3(n8349), .ZN(n11114) );
  INV_X1 U11323 ( .A(n11324), .ZN(n11113) );
  OR2_X1 U11324 ( .A1(n11325), .A2(n11326), .ZN(n11324) );
  AND2_X1 U11325 ( .A1(b_15_), .A2(n11327), .ZN(n11326) );
  OR2_X1 U11326 ( .A1(n11328), .A2(n7314), .ZN(n11327) );
  AND2_X1 U11327 ( .A1(a_30_), .A2(n11329), .ZN(n11328) );
  AND2_X1 U11328 ( .A1(b_14_), .A2(n11330), .ZN(n11325) );
  OR2_X1 U11329 ( .A1(n11331), .A2(n7318), .ZN(n11330) );
  AND2_X1 U11330 ( .A1(a_31_), .A2(n11108), .ZN(n11331) );
  XNOR2_X1 U11331 ( .A(n11332), .B(n11333), .ZN(n11115) );
  XNOR2_X1 U11332 ( .A(n11334), .B(n11335), .ZN(n11333) );
  XOR2_X1 U11333 ( .A(n11336), .B(n11337), .Z(n11119) );
  XOR2_X1 U11334 ( .A(n11338), .B(n11339), .Z(n11337) );
  XOR2_X1 U11335 ( .A(n11340), .B(n11341), .Z(n11123) );
  XOR2_X1 U11336 ( .A(n11342), .B(n11343), .Z(n11341) );
  XOR2_X1 U11337 ( .A(n11344), .B(n11345), .Z(n11127) );
  XOR2_X1 U11338 ( .A(n11346), .B(n11347), .Z(n11345) );
  XOR2_X1 U11339 ( .A(n11348), .B(n11349), .Z(n11131) );
  XOR2_X1 U11340 ( .A(n11350), .B(n11351), .Z(n11349) );
  XOR2_X1 U11341 ( .A(n11352), .B(n11353), .Z(n11135) );
  XOR2_X1 U11342 ( .A(n11354), .B(n11355), .Z(n11353) );
  XOR2_X1 U11343 ( .A(n11356), .B(n11357), .Z(n11139) );
  XOR2_X1 U11344 ( .A(n11358), .B(n11359), .Z(n11357) );
  XOR2_X1 U11345 ( .A(n11360), .B(n11361), .Z(n11143) );
  XOR2_X1 U11346 ( .A(n11362), .B(n11363), .Z(n11361) );
  XOR2_X1 U11347 ( .A(n11364), .B(n11365), .Z(n11147) );
  XOR2_X1 U11348 ( .A(n11366), .B(n11367), .Z(n11365) );
  XOR2_X1 U11349 ( .A(n11368), .B(n11369), .Z(n11151) );
  XOR2_X1 U11350 ( .A(n11370), .B(n11371), .Z(n11369) );
  XOR2_X1 U11351 ( .A(n11372), .B(n11373), .Z(n11155) );
  XOR2_X1 U11352 ( .A(n11374), .B(n11375), .Z(n11373) );
  XOR2_X1 U11353 ( .A(n11376), .B(n11377), .Z(n11159) );
  XOR2_X1 U11354 ( .A(n11378), .B(n11379), .Z(n11377) );
  XOR2_X1 U11355 ( .A(n11380), .B(n11381), .Z(n11167) );
  XOR2_X1 U11356 ( .A(n11382), .B(n11383), .Z(n11381) );
  XNOR2_X1 U11357 ( .A(n11384), .B(n11385), .ZN(n11171) );
  XNOR2_X1 U11358 ( .A(n11386), .B(n11387), .ZN(n11384) );
  XOR2_X1 U11359 ( .A(n11388), .B(n11389), .Z(n11175) );
  XOR2_X1 U11360 ( .A(n11390), .B(n11391), .Z(n11389) );
  XOR2_X1 U11361 ( .A(n11392), .B(n11393), .Z(n11179) );
  XOR2_X1 U11362 ( .A(n11394), .B(n11395), .Z(n11393) );
  XOR2_X1 U11363 ( .A(n11396), .B(n11397), .Z(n11183) );
  XOR2_X1 U11364 ( .A(n11398), .B(n11399), .Z(n11397) );
  XOR2_X1 U11365 ( .A(n11400), .B(n11401), .Z(n11187) );
  XOR2_X1 U11366 ( .A(n11402), .B(n11403), .Z(n11401) );
  XOR2_X1 U11367 ( .A(n11404), .B(n11405), .Z(n11191) );
  XOR2_X1 U11368 ( .A(n11406), .B(n11407), .Z(n11405) );
  XOR2_X1 U11369 ( .A(n11408), .B(n11409), .Z(n11195) );
  XOR2_X1 U11370 ( .A(n11410), .B(n11411), .Z(n11409) );
  XOR2_X1 U11371 ( .A(n11412), .B(n11413), .Z(n11199) );
  XOR2_X1 U11372 ( .A(n11414), .B(n11415), .Z(n11413) );
  XOR2_X1 U11373 ( .A(n11416), .B(n11417), .Z(n11203) );
  XOR2_X1 U11374 ( .A(n11418), .B(n11419), .Z(n11417) );
  XOR2_X1 U11375 ( .A(n11420), .B(n11421), .Z(n10057) );
  XOR2_X1 U11376 ( .A(n11422), .B(n11423), .Z(n11421) );
  XOR2_X1 U11377 ( .A(n11424), .B(n11425), .Z(n10018) );
  XOR2_X1 U11378 ( .A(n11426), .B(n11427), .Z(n11425) );
  XOR2_X1 U11379 ( .A(n11428), .B(n11429), .Z(n7930) );
  XOR2_X1 U11380 ( .A(n11430), .B(n11431), .Z(n11429) );
  XOR2_X1 U11381 ( .A(n11432), .B(n11433), .Z(n7891) );
  XOR2_X1 U11382 ( .A(n11434), .B(n11435), .Z(n11433) );
  XOR2_X1 U11383 ( .A(n11436), .B(n11437), .Z(n7859) );
  XOR2_X1 U11384 ( .A(n11438), .B(n11439), .Z(n11437) );
  XOR2_X1 U11385 ( .A(n11223), .B(n11440), .Z(n7834) );
  XOR2_X1 U11386 ( .A(n11222), .B(n11221), .Z(n11440) );
  OR2_X1 U11387 ( .A1(n11108), .A2(n7656), .ZN(n11221) );
  OR2_X1 U11388 ( .A1(n11441), .A2(n11442), .ZN(n11222) );
  AND2_X1 U11389 ( .A1(n11439), .A2(n11438), .ZN(n11442) );
  AND2_X1 U11390 ( .A1(n11436), .A2(n11443), .ZN(n11441) );
  OR2_X1 U11391 ( .A1(n11438), .A2(n11439), .ZN(n11443) );
  OR2_X1 U11392 ( .A1(n11108), .A2(n7689), .ZN(n11439) );
  OR2_X1 U11393 ( .A1(n11444), .A2(n11445), .ZN(n11438) );
  AND2_X1 U11394 ( .A1(n11435), .A2(n11434), .ZN(n11445) );
  AND2_X1 U11395 ( .A1(n11432), .A2(n11446), .ZN(n11444) );
  OR2_X1 U11396 ( .A1(n11434), .A2(n11435), .ZN(n11446) );
  OR2_X1 U11397 ( .A1(n11108), .A2(n7777), .ZN(n11435) );
  OR2_X1 U11398 ( .A1(n11447), .A2(n11448), .ZN(n11434) );
  AND2_X1 U11399 ( .A1(n11431), .A2(n11430), .ZN(n11448) );
  AND2_X1 U11400 ( .A1(n11428), .A2(n11449), .ZN(n11447) );
  OR2_X1 U11401 ( .A1(n11430), .A2(n11431), .ZN(n11449) );
  OR2_X1 U11402 ( .A1(n11108), .A2(n7785), .ZN(n11431) );
  OR2_X1 U11403 ( .A1(n11450), .A2(n11451), .ZN(n11430) );
  AND2_X1 U11404 ( .A1(n11427), .A2(n11426), .ZN(n11451) );
  AND2_X1 U11405 ( .A1(n11424), .A2(n11452), .ZN(n11450) );
  OR2_X1 U11406 ( .A1(n11426), .A2(n11427), .ZN(n11452) );
  OR2_X1 U11407 ( .A1(n11108), .A2(n8226), .ZN(n11427) );
  OR2_X1 U11408 ( .A1(n11453), .A2(n11454), .ZN(n11426) );
  AND2_X1 U11409 ( .A1(n11423), .A2(n11422), .ZN(n11454) );
  AND2_X1 U11410 ( .A1(n11420), .A2(n11455), .ZN(n11453) );
  OR2_X1 U11411 ( .A1(n11422), .A2(n11423), .ZN(n11455) );
  OR2_X1 U11412 ( .A1(n11108), .A2(n8221), .ZN(n11423) );
  OR2_X1 U11413 ( .A1(n11456), .A2(n11457), .ZN(n11422) );
  AND2_X1 U11414 ( .A1(n11419), .A2(n11418), .ZN(n11457) );
  AND2_X1 U11415 ( .A1(n11416), .A2(n11458), .ZN(n11456) );
  OR2_X1 U11416 ( .A1(n11418), .A2(n11419), .ZN(n11458) );
  OR2_X1 U11417 ( .A1(n11108), .A2(n8216), .ZN(n11419) );
  OR2_X1 U11418 ( .A1(n11459), .A2(n11460), .ZN(n11418) );
  AND2_X1 U11419 ( .A1(n11415), .A2(n11414), .ZN(n11460) );
  AND2_X1 U11420 ( .A1(n11412), .A2(n11461), .ZN(n11459) );
  OR2_X1 U11421 ( .A1(n11414), .A2(n11415), .ZN(n11461) );
  OR2_X1 U11422 ( .A1(n11108), .A2(n8211), .ZN(n11415) );
  OR2_X1 U11423 ( .A1(n11462), .A2(n11463), .ZN(n11414) );
  AND2_X1 U11424 ( .A1(n11411), .A2(n11410), .ZN(n11463) );
  AND2_X1 U11425 ( .A1(n11408), .A2(n11464), .ZN(n11462) );
  OR2_X1 U11426 ( .A1(n11410), .A2(n11411), .ZN(n11464) );
  OR2_X1 U11427 ( .A1(n11108), .A2(n8206), .ZN(n11411) );
  OR2_X1 U11428 ( .A1(n11465), .A2(n11466), .ZN(n11410) );
  AND2_X1 U11429 ( .A1(n11407), .A2(n11406), .ZN(n11466) );
  AND2_X1 U11430 ( .A1(n11404), .A2(n11467), .ZN(n11465) );
  OR2_X1 U11431 ( .A1(n11406), .A2(n11407), .ZN(n11467) );
  OR2_X1 U11432 ( .A1(n11108), .A2(n8201), .ZN(n11407) );
  OR2_X1 U11433 ( .A1(n11468), .A2(n11469), .ZN(n11406) );
  AND2_X1 U11434 ( .A1(n11403), .A2(n11402), .ZN(n11469) );
  AND2_X1 U11435 ( .A1(n11400), .A2(n11470), .ZN(n11468) );
  OR2_X1 U11436 ( .A1(n11402), .A2(n11403), .ZN(n11470) );
  OR2_X1 U11437 ( .A1(n11108), .A2(n8196), .ZN(n11403) );
  OR2_X1 U11438 ( .A1(n11471), .A2(n11472), .ZN(n11402) );
  AND2_X1 U11439 ( .A1(n11399), .A2(n11398), .ZN(n11472) );
  AND2_X1 U11440 ( .A1(n11396), .A2(n11473), .ZN(n11471) );
  OR2_X1 U11441 ( .A1(n11398), .A2(n11399), .ZN(n11473) );
  OR2_X1 U11442 ( .A1(n11108), .A2(n8191), .ZN(n11399) );
  OR2_X1 U11443 ( .A1(n11474), .A2(n11475), .ZN(n11398) );
  AND2_X1 U11444 ( .A1(n11395), .A2(n11394), .ZN(n11475) );
  AND2_X1 U11445 ( .A1(n11392), .A2(n11476), .ZN(n11474) );
  OR2_X1 U11446 ( .A1(n11394), .A2(n11395), .ZN(n11476) );
  OR2_X1 U11447 ( .A1(n11108), .A2(n8186), .ZN(n11395) );
  OR2_X1 U11448 ( .A1(n11477), .A2(n11478), .ZN(n11394) );
  AND2_X1 U11449 ( .A1(n11391), .A2(n11390), .ZN(n11478) );
  AND2_X1 U11450 ( .A1(n11388), .A2(n11479), .ZN(n11477) );
  OR2_X1 U11451 ( .A1(n11390), .A2(n11391), .ZN(n11479) );
  OR2_X1 U11452 ( .A1(n11108), .A2(n8181), .ZN(n11391) );
  OR2_X1 U11453 ( .A1(n11480), .A2(n11481), .ZN(n11390) );
  AND2_X1 U11454 ( .A1(n11385), .A2(n11387), .ZN(n11481) );
  AND2_X1 U11455 ( .A1(n11482), .A2(n11386), .ZN(n11480) );
  OR2_X1 U11456 ( .A1(n11385), .A2(n11387), .ZN(n11482) );
  OR2_X1 U11457 ( .A1(n11483), .A2(n11484), .ZN(n11387) );
  AND2_X1 U11458 ( .A1(n11383), .A2(n11382), .ZN(n11484) );
  AND2_X1 U11459 ( .A1(n11380), .A2(n11485), .ZN(n11483) );
  OR2_X1 U11460 ( .A1(n11382), .A2(n11383), .ZN(n11485) );
  OR2_X1 U11461 ( .A1(n11108), .A2(n8171), .ZN(n11383) );
  OR2_X1 U11462 ( .A1(n11486), .A2(n11487), .ZN(n11382) );
  AND2_X1 U11463 ( .A1(n11284), .A2(n11283), .ZN(n11487) );
  AND2_X1 U11464 ( .A1(n11281), .A2(n11488), .ZN(n11486) );
  OR2_X1 U11465 ( .A1(n11283), .A2(n11284), .ZN(n11488) );
  OR2_X1 U11466 ( .A1(n8166), .A2(n11108), .ZN(n11284) );
  OR2_X1 U11467 ( .A1(n11489), .A2(n11490), .ZN(n11283) );
  AND2_X1 U11468 ( .A1(n11379), .A2(n11378), .ZN(n11490) );
  AND2_X1 U11469 ( .A1(n11376), .A2(n11491), .ZN(n11489) );
  OR2_X1 U11470 ( .A1(n11378), .A2(n11379), .ZN(n11491) );
  OR2_X1 U11471 ( .A1(n11108), .A2(n8161), .ZN(n11379) );
  OR2_X1 U11472 ( .A1(n11492), .A2(n11493), .ZN(n11378) );
  AND2_X1 U11473 ( .A1(n11375), .A2(n11374), .ZN(n11493) );
  AND2_X1 U11474 ( .A1(n11372), .A2(n11494), .ZN(n11492) );
  OR2_X1 U11475 ( .A1(n11374), .A2(n11375), .ZN(n11494) );
  OR2_X1 U11476 ( .A1(n11108), .A2(n8156), .ZN(n11375) );
  OR2_X1 U11477 ( .A1(n11495), .A2(n11496), .ZN(n11374) );
  AND2_X1 U11478 ( .A1(n11371), .A2(n11370), .ZN(n11496) );
  AND2_X1 U11479 ( .A1(n11368), .A2(n11497), .ZN(n11495) );
  OR2_X1 U11480 ( .A1(n11370), .A2(n11371), .ZN(n11497) );
  OR2_X1 U11481 ( .A1(n11108), .A2(n8151), .ZN(n11371) );
  OR2_X1 U11482 ( .A1(n11498), .A2(n11499), .ZN(n11370) );
  AND2_X1 U11483 ( .A1(n11367), .A2(n11366), .ZN(n11499) );
  AND2_X1 U11484 ( .A1(n11364), .A2(n11500), .ZN(n11498) );
  OR2_X1 U11485 ( .A1(n11366), .A2(n11367), .ZN(n11500) );
  OR2_X1 U11486 ( .A1(n11108), .A2(n8146), .ZN(n11367) );
  OR2_X1 U11487 ( .A1(n11501), .A2(n11502), .ZN(n11366) );
  AND2_X1 U11488 ( .A1(n11363), .A2(n11362), .ZN(n11502) );
  AND2_X1 U11489 ( .A1(n11360), .A2(n11503), .ZN(n11501) );
  OR2_X1 U11490 ( .A1(n11362), .A2(n11363), .ZN(n11503) );
  OR2_X1 U11491 ( .A1(n11108), .A2(n8141), .ZN(n11363) );
  OR2_X1 U11492 ( .A1(n11504), .A2(n11505), .ZN(n11362) );
  AND2_X1 U11493 ( .A1(n11359), .A2(n11358), .ZN(n11505) );
  AND2_X1 U11494 ( .A1(n11356), .A2(n11506), .ZN(n11504) );
  OR2_X1 U11495 ( .A1(n11358), .A2(n11359), .ZN(n11506) );
  OR2_X1 U11496 ( .A1(n11108), .A2(n8136), .ZN(n11359) );
  OR2_X1 U11497 ( .A1(n11507), .A2(n11508), .ZN(n11358) );
  AND2_X1 U11498 ( .A1(n11355), .A2(n11354), .ZN(n11508) );
  AND2_X1 U11499 ( .A1(n11352), .A2(n11509), .ZN(n11507) );
  OR2_X1 U11500 ( .A1(n11354), .A2(n11355), .ZN(n11509) );
  OR2_X1 U11501 ( .A1(n11108), .A2(n8131), .ZN(n11355) );
  OR2_X1 U11502 ( .A1(n11510), .A2(n11511), .ZN(n11354) );
  AND2_X1 U11503 ( .A1(n11351), .A2(n11350), .ZN(n11511) );
  AND2_X1 U11504 ( .A1(n11348), .A2(n11512), .ZN(n11510) );
  OR2_X1 U11505 ( .A1(n11350), .A2(n11351), .ZN(n11512) );
  OR2_X1 U11506 ( .A1(n11108), .A2(n8126), .ZN(n11351) );
  OR2_X1 U11507 ( .A1(n11513), .A2(n11514), .ZN(n11350) );
  AND2_X1 U11508 ( .A1(n11347), .A2(n11346), .ZN(n11514) );
  AND2_X1 U11509 ( .A1(n11344), .A2(n11515), .ZN(n11513) );
  OR2_X1 U11510 ( .A1(n11346), .A2(n11347), .ZN(n11515) );
  OR2_X1 U11511 ( .A1(n11108), .A2(n8121), .ZN(n11347) );
  OR2_X1 U11512 ( .A1(n11516), .A2(n11517), .ZN(n11346) );
  AND2_X1 U11513 ( .A1(n11343), .A2(n11342), .ZN(n11517) );
  AND2_X1 U11514 ( .A1(n11340), .A2(n11518), .ZN(n11516) );
  OR2_X1 U11515 ( .A1(n11342), .A2(n11343), .ZN(n11518) );
  OR2_X1 U11516 ( .A1(n11108), .A2(n8116), .ZN(n11343) );
  OR2_X1 U11517 ( .A1(n11519), .A2(n11520), .ZN(n11342) );
  AND2_X1 U11518 ( .A1(n11339), .A2(n11338), .ZN(n11520) );
  AND2_X1 U11519 ( .A1(n11336), .A2(n11521), .ZN(n11519) );
  OR2_X1 U11520 ( .A1(n11338), .A2(n11339), .ZN(n11521) );
  OR2_X1 U11521 ( .A1(n11108), .A2(n8111), .ZN(n11339) );
  OR2_X1 U11522 ( .A1(n11522), .A2(n11523), .ZN(n11338) );
  AND2_X1 U11523 ( .A1(n11332), .A2(n11335), .ZN(n11523) );
  AND2_X1 U11524 ( .A1(n11334), .A2(n11524), .ZN(n11522) );
  OR2_X1 U11525 ( .A1(n11335), .A2(n11332), .ZN(n11524) );
  OR2_X1 U11526 ( .A1(n11108), .A2(n8102), .ZN(n11332) );
  OR3_X1 U11527 ( .A1(n11108), .A2(n8349), .A3(n11329), .ZN(n11335) );
  INV_X1 U11528 ( .A(n11525), .ZN(n11334) );
  OR2_X1 U11529 ( .A1(n11526), .A2(n11527), .ZN(n11525) );
  AND2_X1 U11530 ( .A1(b_14_), .A2(n11528), .ZN(n11527) );
  OR2_X1 U11531 ( .A1(n11529), .A2(n7314), .ZN(n11528) );
  AND2_X1 U11532 ( .A1(a_30_), .A2(n11530), .ZN(n11529) );
  AND2_X1 U11533 ( .A1(b_13_), .A2(n11531), .ZN(n11526) );
  OR2_X1 U11534 ( .A1(n11532), .A2(n7318), .ZN(n11531) );
  AND2_X1 U11535 ( .A1(a_31_), .A2(n11329), .ZN(n11532) );
  XNOR2_X1 U11536 ( .A(n11533), .B(n11534), .ZN(n11336) );
  XNOR2_X1 U11537 ( .A(n11535), .B(n11536), .ZN(n11534) );
  XOR2_X1 U11538 ( .A(n11537), .B(n11538), .Z(n11340) );
  XOR2_X1 U11539 ( .A(n11539), .B(n11540), .Z(n11538) );
  XOR2_X1 U11540 ( .A(n11541), .B(n11542), .Z(n11344) );
  XOR2_X1 U11541 ( .A(n11543), .B(n11544), .Z(n11542) );
  XOR2_X1 U11542 ( .A(n11545), .B(n11546), .Z(n11348) );
  XOR2_X1 U11543 ( .A(n11547), .B(n11548), .Z(n11546) );
  XOR2_X1 U11544 ( .A(n11549), .B(n11550), .Z(n11352) );
  XOR2_X1 U11545 ( .A(n11551), .B(n11552), .Z(n11550) );
  XOR2_X1 U11546 ( .A(n11553), .B(n11554), .Z(n11356) );
  XOR2_X1 U11547 ( .A(n11555), .B(n11556), .Z(n11554) );
  XOR2_X1 U11548 ( .A(n11557), .B(n11558), .Z(n11360) );
  XOR2_X1 U11549 ( .A(n11559), .B(n11560), .Z(n11558) );
  XOR2_X1 U11550 ( .A(n11561), .B(n11562), .Z(n11364) );
  XOR2_X1 U11551 ( .A(n11563), .B(n11564), .Z(n11562) );
  XOR2_X1 U11552 ( .A(n11565), .B(n11566), .Z(n11368) );
  XOR2_X1 U11553 ( .A(n11567), .B(n11568), .Z(n11566) );
  XOR2_X1 U11554 ( .A(n11569), .B(n11570), .Z(n11372) );
  XOR2_X1 U11555 ( .A(n11571), .B(n11572), .Z(n11570) );
  XOR2_X1 U11556 ( .A(n11573), .B(n11574), .Z(n11376) );
  XOR2_X1 U11557 ( .A(n11575), .B(n11576), .Z(n11574) );
  XOR2_X1 U11558 ( .A(n11577), .B(n11578), .Z(n11281) );
  XOR2_X1 U11559 ( .A(n11579), .B(n11580), .Z(n11578) );
  XOR2_X1 U11560 ( .A(n11581), .B(n11582), .Z(n11380) );
  XOR2_X1 U11561 ( .A(n11583), .B(n11584), .Z(n11582) );
  XOR2_X1 U11562 ( .A(n11585), .B(n11586), .Z(n11385) );
  XOR2_X1 U11563 ( .A(n11587), .B(n11588), .Z(n11586) );
  XOR2_X1 U11564 ( .A(n11589), .B(n11590), .Z(n11388) );
  XOR2_X1 U11565 ( .A(n11591), .B(n11592), .Z(n11590) );
  XNOR2_X1 U11566 ( .A(n11593), .B(n11594), .ZN(n11392) );
  XNOR2_X1 U11567 ( .A(n11595), .B(n11596), .ZN(n11593) );
  XOR2_X1 U11568 ( .A(n11597), .B(n11598), .Z(n11396) );
  XOR2_X1 U11569 ( .A(n11599), .B(n11600), .Z(n11598) );
  XOR2_X1 U11570 ( .A(n11601), .B(n11602), .Z(n11400) );
  XOR2_X1 U11571 ( .A(n11603), .B(n11604), .Z(n11602) );
  XOR2_X1 U11572 ( .A(n11605), .B(n11606), .Z(n11404) );
  XOR2_X1 U11573 ( .A(n11607), .B(n11608), .Z(n11606) );
  XOR2_X1 U11574 ( .A(n11609), .B(n11610), .Z(n11408) );
  XOR2_X1 U11575 ( .A(n11611), .B(n11612), .Z(n11610) );
  XOR2_X1 U11576 ( .A(n11613), .B(n11614), .Z(n11412) );
  XOR2_X1 U11577 ( .A(n11615), .B(n11616), .Z(n11614) );
  XOR2_X1 U11578 ( .A(n11617), .B(n11618), .Z(n11416) );
  XOR2_X1 U11579 ( .A(n11619), .B(n11620), .Z(n11618) );
  XOR2_X1 U11580 ( .A(n11621), .B(n11622), .Z(n11420) );
  XOR2_X1 U11581 ( .A(n11623), .B(n11624), .Z(n11622) );
  XOR2_X1 U11582 ( .A(n11625), .B(n11626), .Z(n11424) );
  XOR2_X1 U11583 ( .A(n11627), .B(n11628), .Z(n11626) );
  XOR2_X1 U11584 ( .A(n11629), .B(n11630), .Z(n11428) );
  XOR2_X1 U11585 ( .A(n11631), .B(n11632), .Z(n11630) );
  XOR2_X1 U11586 ( .A(n11633), .B(n11634), .Z(n11432) );
  XOR2_X1 U11587 ( .A(n11635), .B(n11636), .Z(n11634) );
  XOR2_X1 U11588 ( .A(n11637), .B(n11638), .Z(n11436) );
  XOR2_X1 U11589 ( .A(n11639), .B(n11640), .Z(n11638) );
  XOR2_X1 U11590 ( .A(n11641), .B(n11642), .Z(n11223) );
  XOR2_X1 U11591 ( .A(n11643), .B(n11644), .Z(n11642) );
  XNOR2_X1 U11592 ( .A(n7561), .B(n7807), .ZN(n7550) );
  OR2_X1 U11593 ( .A1(n11645), .A2(n11646), .ZN(n7807) );
  AND2_X1 U11594 ( .A1(n11217), .A2(n11216), .ZN(n11646) );
  AND2_X1 U11595 ( .A1(n11214), .A2(n11647), .ZN(n11645) );
  OR2_X1 U11596 ( .A1(n11216), .A2(n11217), .ZN(n11647) );
  OR2_X1 U11597 ( .A1(n11329), .A2(n7621), .ZN(n11217) );
  OR2_X1 U11598 ( .A1(n11648), .A2(n11649), .ZN(n11216) );
  AND2_X1 U11599 ( .A1(n11228), .A2(n11227), .ZN(n11649) );
  AND2_X1 U11600 ( .A1(n11225), .A2(n11650), .ZN(n11648) );
  OR2_X1 U11601 ( .A1(n11227), .A2(n11228), .ZN(n11650) );
  OR2_X1 U11602 ( .A1(n11329), .A2(n7656), .ZN(n11228) );
  OR2_X1 U11603 ( .A1(n11651), .A2(n11652), .ZN(n11227) );
  AND2_X1 U11604 ( .A1(n11644), .A2(n11643), .ZN(n11652) );
  AND2_X1 U11605 ( .A1(n11641), .A2(n11653), .ZN(n11651) );
  OR2_X1 U11606 ( .A1(n11643), .A2(n11644), .ZN(n11653) );
  OR2_X1 U11607 ( .A1(n11329), .A2(n7689), .ZN(n11644) );
  OR2_X1 U11608 ( .A1(n11654), .A2(n11655), .ZN(n11643) );
  AND2_X1 U11609 ( .A1(n11640), .A2(n11639), .ZN(n11655) );
  AND2_X1 U11610 ( .A1(n11637), .A2(n11656), .ZN(n11654) );
  OR2_X1 U11611 ( .A1(n11639), .A2(n11640), .ZN(n11656) );
  OR2_X1 U11612 ( .A1(n11329), .A2(n7777), .ZN(n11640) );
  OR2_X1 U11613 ( .A1(n11657), .A2(n11658), .ZN(n11639) );
  AND2_X1 U11614 ( .A1(n11636), .A2(n11635), .ZN(n11658) );
  AND2_X1 U11615 ( .A1(n11633), .A2(n11659), .ZN(n11657) );
  OR2_X1 U11616 ( .A1(n11635), .A2(n11636), .ZN(n11659) );
  OR2_X1 U11617 ( .A1(n11329), .A2(n7785), .ZN(n11636) );
  OR2_X1 U11618 ( .A1(n11660), .A2(n11661), .ZN(n11635) );
  AND2_X1 U11619 ( .A1(n11632), .A2(n11631), .ZN(n11661) );
  AND2_X1 U11620 ( .A1(n11629), .A2(n11662), .ZN(n11660) );
  OR2_X1 U11621 ( .A1(n11631), .A2(n11632), .ZN(n11662) );
  OR2_X1 U11622 ( .A1(n11329), .A2(n8226), .ZN(n11632) );
  OR2_X1 U11623 ( .A1(n11663), .A2(n11664), .ZN(n11631) );
  AND2_X1 U11624 ( .A1(n11628), .A2(n11627), .ZN(n11664) );
  AND2_X1 U11625 ( .A1(n11625), .A2(n11665), .ZN(n11663) );
  OR2_X1 U11626 ( .A1(n11627), .A2(n11628), .ZN(n11665) );
  OR2_X1 U11627 ( .A1(n11329), .A2(n8221), .ZN(n11628) );
  OR2_X1 U11628 ( .A1(n11666), .A2(n11667), .ZN(n11627) );
  AND2_X1 U11629 ( .A1(n11624), .A2(n11623), .ZN(n11667) );
  AND2_X1 U11630 ( .A1(n11621), .A2(n11668), .ZN(n11666) );
  OR2_X1 U11631 ( .A1(n11623), .A2(n11624), .ZN(n11668) );
  OR2_X1 U11632 ( .A1(n11329), .A2(n8216), .ZN(n11624) );
  OR2_X1 U11633 ( .A1(n11669), .A2(n11670), .ZN(n11623) );
  AND2_X1 U11634 ( .A1(n11620), .A2(n11619), .ZN(n11670) );
  AND2_X1 U11635 ( .A1(n11617), .A2(n11671), .ZN(n11669) );
  OR2_X1 U11636 ( .A1(n11619), .A2(n11620), .ZN(n11671) );
  OR2_X1 U11637 ( .A1(n11329), .A2(n8211), .ZN(n11620) );
  OR2_X1 U11638 ( .A1(n11672), .A2(n11673), .ZN(n11619) );
  AND2_X1 U11639 ( .A1(n11616), .A2(n11615), .ZN(n11673) );
  AND2_X1 U11640 ( .A1(n11613), .A2(n11674), .ZN(n11672) );
  OR2_X1 U11641 ( .A1(n11615), .A2(n11616), .ZN(n11674) );
  OR2_X1 U11642 ( .A1(n11329), .A2(n8206), .ZN(n11616) );
  OR2_X1 U11643 ( .A1(n11675), .A2(n11676), .ZN(n11615) );
  AND2_X1 U11644 ( .A1(n11612), .A2(n11611), .ZN(n11676) );
  AND2_X1 U11645 ( .A1(n11609), .A2(n11677), .ZN(n11675) );
  OR2_X1 U11646 ( .A1(n11611), .A2(n11612), .ZN(n11677) );
  OR2_X1 U11647 ( .A1(n11329), .A2(n8201), .ZN(n11612) );
  OR2_X1 U11648 ( .A1(n11678), .A2(n11679), .ZN(n11611) );
  AND2_X1 U11649 ( .A1(n11608), .A2(n11607), .ZN(n11679) );
  AND2_X1 U11650 ( .A1(n11605), .A2(n11680), .ZN(n11678) );
  OR2_X1 U11651 ( .A1(n11607), .A2(n11608), .ZN(n11680) );
  OR2_X1 U11652 ( .A1(n11329), .A2(n8196), .ZN(n11608) );
  OR2_X1 U11653 ( .A1(n11681), .A2(n11682), .ZN(n11607) );
  AND2_X1 U11654 ( .A1(n11604), .A2(n11603), .ZN(n11682) );
  AND2_X1 U11655 ( .A1(n11601), .A2(n11683), .ZN(n11681) );
  OR2_X1 U11656 ( .A1(n11603), .A2(n11604), .ZN(n11683) );
  OR2_X1 U11657 ( .A1(n11329), .A2(n8191), .ZN(n11604) );
  OR2_X1 U11658 ( .A1(n11684), .A2(n11685), .ZN(n11603) );
  AND2_X1 U11659 ( .A1(n11600), .A2(n11599), .ZN(n11685) );
  AND2_X1 U11660 ( .A1(n11597), .A2(n11686), .ZN(n11684) );
  OR2_X1 U11661 ( .A1(n11599), .A2(n11600), .ZN(n11686) );
  OR2_X1 U11662 ( .A1(n11329), .A2(n8186), .ZN(n11600) );
  OR2_X1 U11663 ( .A1(n11687), .A2(n11688), .ZN(n11599) );
  AND2_X1 U11664 ( .A1(n11594), .A2(n11596), .ZN(n11688) );
  AND2_X1 U11665 ( .A1(n11689), .A2(n11595), .ZN(n11687) );
  OR2_X1 U11666 ( .A1(n11594), .A2(n11596), .ZN(n11689) );
  OR2_X1 U11667 ( .A1(n11690), .A2(n11691), .ZN(n11596) );
  AND2_X1 U11668 ( .A1(n11592), .A2(n11591), .ZN(n11691) );
  AND2_X1 U11669 ( .A1(n11589), .A2(n11692), .ZN(n11690) );
  OR2_X1 U11670 ( .A1(n11591), .A2(n11592), .ZN(n11692) );
  OR2_X1 U11671 ( .A1(n11329), .A2(n8176), .ZN(n11592) );
  OR2_X1 U11672 ( .A1(n11693), .A2(n11694), .ZN(n11591) );
  AND2_X1 U11673 ( .A1(n11588), .A2(n11587), .ZN(n11694) );
  AND2_X1 U11674 ( .A1(n11585), .A2(n11695), .ZN(n11693) );
  OR2_X1 U11675 ( .A1(n11587), .A2(n11588), .ZN(n11695) );
  OR2_X1 U11676 ( .A1(n11329), .A2(n8171), .ZN(n11588) );
  OR2_X1 U11677 ( .A1(n11696), .A2(n11697), .ZN(n11587) );
  AND2_X1 U11678 ( .A1(n11584), .A2(n11583), .ZN(n11697) );
  AND2_X1 U11679 ( .A1(n11581), .A2(n11698), .ZN(n11696) );
  OR2_X1 U11680 ( .A1(n11583), .A2(n11584), .ZN(n11698) );
  OR2_X1 U11681 ( .A1(n8166), .A2(n11329), .ZN(n11584) );
  OR2_X1 U11682 ( .A1(n11699), .A2(n11700), .ZN(n11583) );
  AND2_X1 U11683 ( .A1(n11580), .A2(n11579), .ZN(n11700) );
  AND2_X1 U11684 ( .A1(n11577), .A2(n11701), .ZN(n11699) );
  OR2_X1 U11685 ( .A1(n11579), .A2(n11580), .ZN(n11701) );
  OR2_X1 U11686 ( .A1(n11329), .A2(n8161), .ZN(n11580) );
  OR2_X1 U11687 ( .A1(n11702), .A2(n11703), .ZN(n11579) );
  AND2_X1 U11688 ( .A1(n11576), .A2(n11575), .ZN(n11703) );
  AND2_X1 U11689 ( .A1(n11573), .A2(n11704), .ZN(n11702) );
  OR2_X1 U11690 ( .A1(n11575), .A2(n11576), .ZN(n11704) );
  OR2_X1 U11691 ( .A1(n11329), .A2(n8156), .ZN(n11576) );
  OR2_X1 U11692 ( .A1(n11705), .A2(n11706), .ZN(n11575) );
  AND2_X1 U11693 ( .A1(n11572), .A2(n11571), .ZN(n11706) );
  AND2_X1 U11694 ( .A1(n11569), .A2(n11707), .ZN(n11705) );
  OR2_X1 U11695 ( .A1(n11571), .A2(n11572), .ZN(n11707) );
  OR2_X1 U11696 ( .A1(n11329), .A2(n8151), .ZN(n11572) );
  OR2_X1 U11697 ( .A1(n11708), .A2(n11709), .ZN(n11571) );
  AND2_X1 U11698 ( .A1(n11568), .A2(n11567), .ZN(n11709) );
  AND2_X1 U11699 ( .A1(n11565), .A2(n11710), .ZN(n11708) );
  OR2_X1 U11700 ( .A1(n11567), .A2(n11568), .ZN(n11710) );
  OR2_X1 U11701 ( .A1(n11329), .A2(n8146), .ZN(n11568) );
  OR2_X1 U11702 ( .A1(n11711), .A2(n11712), .ZN(n11567) );
  AND2_X1 U11703 ( .A1(n11564), .A2(n11563), .ZN(n11712) );
  AND2_X1 U11704 ( .A1(n11561), .A2(n11713), .ZN(n11711) );
  OR2_X1 U11705 ( .A1(n11563), .A2(n11564), .ZN(n11713) );
  OR2_X1 U11706 ( .A1(n11329), .A2(n8141), .ZN(n11564) );
  OR2_X1 U11707 ( .A1(n11714), .A2(n11715), .ZN(n11563) );
  AND2_X1 U11708 ( .A1(n11560), .A2(n11559), .ZN(n11715) );
  AND2_X1 U11709 ( .A1(n11557), .A2(n11716), .ZN(n11714) );
  OR2_X1 U11710 ( .A1(n11559), .A2(n11560), .ZN(n11716) );
  OR2_X1 U11711 ( .A1(n11329), .A2(n8136), .ZN(n11560) );
  OR2_X1 U11712 ( .A1(n11717), .A2(n11718), .ZN(n11559) );
  AND2_X1 U11713 ( .A1(n11556), .A2(n11555), .ZN(n11718) );
  AND2_X1 U11714 ( .A1(n11553), .A2(n11719), .ZN(n11717) );
  OR2_X1 U11715 ( .A1(n11555), .A2(n11556), .ZN(n11719) );
  OR2_X1 U11716 ( .A1(n11329), .A2(n8131), .ZN(n11556) );
  OR2_X1 U11717 ( .A1(n11720), .A2(n11721), .ZN(n11555) );
  AND2_X1 U11718 ( .A1(n11552), .A2(n11551), .ZN(n11721) );
  AND2_X1 U11719 ( .A1(n11549), .A2(n11722), .ZN(n11720) );
  OR2_X1 U11720 ( .A1(n11551), .A2(n11552), .ZN(n11722) );
  OR2_X1 U11721 ( .A1(n11329), .A2(n8126), .ZN(n11552) );
  OR2_X1 U11722 ( .A1(n11723), .A2(n11724), .ZN(n11551) );
  AND2_X1 U11723 ( .A1(n11548), .A2(n11547), .ZN(n11724) );
  AND2_X1 U11724 ( .A1(n11545), .A2(n11725), .ZN(n11723) );
  OR2_X1 U11725 ( .A1(n11547), .A2(n11548), .ZN(n11725) );
  OR2_X1 U11726 ( .A1(n11329), .A2(n8121), .ZN(n11548) );
  OR2_X1 U11727 ( .A1(n11726), .A2(n11727), .ZN(n11547) );
  AND2_X1 U11728 ( .A1(n11544), .A2(n11543), .ZN(n11727) );
  AND2_X1 U11729 ( .A1(n11541), .A2(n11728), .ZN(n11726) );
  OR2_X1 U11730 ( .A1(n11543), .A2(n11544), .ZN(n11728) );
  OR2_X1 U11731 ( .A1(n11329), .A2(n8116), .ZN(n11544) );
  OR2_X1 U11732 ( .A1(n11729), .A2(n11730), .ZN(n11543) );
  AND2_X1 U11733 ( .A1(n11540), .A2(n11539), .ZN(n11730) );
  AND2_X1 U11734 ( .A1(n11537), .A2(n11731), .ZN(n11729) );
  OR2_X1 U11735 ( .A1(n11539), .A2(n11540), .ZN(n11731) );
  OR2_X1 U11736 ( .A1(n8111), .A2(n11329), .ZN(n11540) );
  OR2_X1 U11737 ( .A1(n11732), .A2(n11733), .ZN(n11539) );
  AND2_X1 U11738 ( .A1(n11533), .A2(n11536), .ZN(n11733) );
  AND2_X1 U11739 ( .A1(n11535), .A2(n11734), .ZN(n11732) );
  OR2_X1 U11740 ( .A1(n11536), .A2(n11533), .ZN(n11734) );
  OR2_X1 U11741 ( .A1(n8102), .A2(n11329), .ZN(n11533) );
  OR3_X1 U11742 ( .A1(n8349), .A2(n11329), .A3(n11530), .ZN(n11536) );
  INV_X1 U11743 ( .A(n11735), .ZN(n11535) );
  OR2_X1 U11744 ( .A1(n11736), .A2(n11737), .ZN(n11735) );
  AND2_X1 U11745 ( .A1(b_13_), .A2(n11738), .ZN(n11737) );
  OR2_X1 U11746 ( .A1(n11739), .A2(n7314), .ZN(n11738) );
  AND2_X1 U11747 ( .A1(a_30_), .A2(n11740), .ZN(n11739) );
  AND2_X1 U11748 ( .A1(b_12_), .A2(n11741), .ZN(n11736) );
  OR2_X1 U11749 ( .A1(n11742), .A2(n7318), .ZN(n11741) );
  AND2_X1 U11750 ( .A1(a_31_), .A2(n11530), .ZN(n11742) );
  XNOR2_X1 U11751 ( .A(n11743), .B(n11744), .ZN(n11537) );
  XNOR2_X1 U11752 ( .A(n11745), .B(n11746), .ZN(n11744) );
  XOR2_X1 U11753 ( .A(n11747), .B(n11748), .Z(n11541) );
  XOR2_X1 U11754 ( .A(n11749), .B(n11750), .Z(n11748) );
  XOR2_X1 U11755 ( .A(n11751), .B(n11752), .Z(n11545) );
  XOR2_X1 U11756 ( .A(n11753), .B(n11754), .Z(n11752) );
  XOR2_X1 U11757 ( .A(n11755), .B(n11756), .Z(n11549) );
  XOR2_X1 U11758 ( .A(n11757), .B(n11758), .Z(n11756) );
  XOR2_X1 U11759 ( .A(n11759), .B(n11760), .Z(n11553) );
  XOR2_X1 U11760 ( .A(n11761), .B(n11762), .Z(n11760) );
  XOR2_X1 U11761 ( .A(n11763), .B(n11764), .Z(n11557) );
  XOR2_X1 U11762 ( .A(n11765), .B(n11766), .Z(n11764) );
  XOR2_X1 U11763 ( .A(n11767), .B(n11768), .Z(n11561) );
  XOR2_X1 U11764 ( .A(n11769), .B(n11770), .Z(n11768) );
  XOR2_X1 U11765 ( .A(n11771), .B(n11772), .Z(n11565) );
  XOR2_X1 U11766 ( .A(n11773), .B(n11774), .Z(n11772) );
  XOR2_X1 U11767 ( .A(n11775), .B(n11776), .Z(n11569) );
  XOR2_X1 U11768 ( .A(n11777), .B(n11778), .Z(n11776) );
  XOR2_X1 U11769 ( .A(n11779), .B(n11780), .Z(n11573) );
  XOR2_X1 U11770 ( .A(n11781), .B(n11782), .Z(n11780) );
  XOR2_X1 U11771 ( .A(n11783), .B(n11784), .Z(n11577) );
  XOR2_X1 U11772 ( .A(n11785), .B(n11786), .Z(n11784) );
  XOR2_X1 U11773 ( .A(n11787), .B(n11788), .Z(n11581) );
  XOR2_X1 U11774 ( .A(n11789), .B(n11790), .Z(n11788) );
  XOR2_X1 U11775 ( .A(n11791), .B(n11792), .Z(n11585) );
  XOR2_X1 U11776 ( .A(n11793), .B(n11794), .Z(n11792) );
  XOR2_X1 U11777 ( .A(n11795), .B(n11796), .Z(n11589) );
  XOR2_X1 U11778 ( .A(n11797), .B(n11798), .Z(n11796) );
  XOR2_X1 U11779 ( .A(n11799), .B(n11800), .Z(n11594) );
  XOR2_X1 U11780 ( .A(n11801), .B(n11802), .Z(n11800) );
  XOR2_X1 U11781 ( .A(n11803), .B(n11804), .Z(n11597) );
  XOR2_X1 U11782 ( .A(n11805), .B(n11806), .Z(n11804) );
  XNOR2_X1 U11783 ( .A(n11807), .B(n11808), .ZN(n11601) );
  XNOR2_X1 U11784 ( .A(n11809), .B(n11810), .ZN(n11807) );
  XOR2_X1 U11785 ( .A(n11811), .B(n11812), .Z(n11605) );
  XOR2_X1 U11786 ( .A(n11813), .B(n11814), .Z(n11812) );
  XOR2_X1 U11787 ( .A(n11815), .B(n11816), .Z(n11609) );
  XOR2_X1 U11788 ( .A(n11817), .B(n11818), .Z(n11816) );
  XOR2_X1 U11789 ( .A(n11819), .B(n11820), .Z(n11613) );
  XOR2_X1 U11790 ( .A(n11821), .B(n11822), .Z(n11820) );
  XOR2_X1 U11791 ( .A(n11823), .B(n11824), .Z(n11617) );
  XOR2_X1 U11792 ( .A(n11825), .B(n11826), .Z(n11824) );
  XOR2_X1 U11793 ( .A(n11827), .B(n11828), .Z(n11621) );
  XOR2_X1 U11794 ( .A(n11829), .B(n11830), .Z(n11828) );
  XOR2_X1 U11795 ( .A(n11831), .B(n11832), .Z(n11625) );
  XOR2_X1 U11796 ( .A(n11833), .B(n11834), .Z(n11832) );
  XOR2_X1 U11797 ( .A(n11835), .B(n11836), .Z(n11629) );
  XOR2_X1 U11798 ( .A(n11837), .B(n11838), .Z(n11836) );
  XOR2_X1 U11799 ( .A(n11839), .B(n11840), .Z(n11633) );
  XOR2_X1 U11800 ( .A(n11841), .B(n11842), .Z(n11840) );
  XOR2_X1 U11801 ( .A(n11843), .B(n11844), .Z(n11637) );
  XOR2_X1 U11802 ( .A(n11845), .B(n11846), .Z(n11844) );
  XOR2_X1 U11803 ( .A(n11847), .B(n11848), .Z(n11641) );
  XOR2_X1 U11804 ( .A(n11849), .B(n11850), .Z(n11848) );
  XOR2_X1 U11805 ( .A(n11851), .B(n11852), .Z(n11225) );
  XOR2_X1 U11806 ( .A(n11853), .B(n11854), .Z(n11852) );
  XOR2_X1 U11807 ( .A(n11855), .B(n11856), .Z(n11214) );
  XOR2_X1 U11808 ( .A(n11857), .B(n11858), .Z(n11856) );
  XNOR2_X1 U11809 ( .A(n11859), .B(n11860), .ZN(n7561) );
  XOR2_X1 U11810 ( .A(n11861), .B(n11862), .Z(n11860) );
  XNOR2_X1 U11811 ( .A(n7570), .B(n7805), .ZN(n7559) );
  OR2_X1 U11812 ( .A1(n11863), .A2(n11864), .ZN(n7805) );
  AND2_X1 U11813 ( .A1(n11862), .A2(n11861), .ZN(n11864) );
  AND2_X1 U11814 ( .A1(n11859), .A2(n11865), .ZN(n11863) );
  OR2_X1 U11815 ( .A1(n11861), .A2(n11862), .ZN(n11865) );
  OR2_X1 U11816 ( .A1(n11530), .A2(n7621), .ZN(n11862) );
  OR2_X1 U11817 ( .A1(n11866), .A2(n11867), .ZN(n11861) );
  AND2_X1 U11818 ( .A1(n11858), .A2(n11857), .ZN(n11867) );
  AND2_X1 U11819 ( .A1(n11855), .A2(n11868), .ZN(n11866) );
  OR2_X1 U11820 ( .A1(n11857), .A2(n11858), .ZN(n11868) );
  OR2_X1 U11821 ( .A1(n11530), .A2(n7656), .ZN(n11858) );
  OR2_X1 U11822 ( .A1(n11869), .A2(n11870), .ZN(n11857) );
  AND2_X1 U11823 ( .A1(n11854), .A2(n11853), .ZN(n11870) );
  AND2_X1 U11824 ( .A1(n11851), .A2(n11871), .ZN(n11869) );
  OR2_X1 U11825 ( .A1(n11853), .A2(n11854), .ZN(n11871) );
  OR2_X1 U11826 ( .A1(n11530), .A2(n7689), .ZN(n11854) );
  OR2_X1 U11827 ( .A1(n11872), .A2(n11873), .ZN(n11853) );
  AND2_X1 U11828 ( .A1(n11850), .A2(n11849), .ZN(n11873) );
  AND2_X1 U11829 ( .A1(n11847), .A2(n11874), .ZN(n11872) );
  OR2_X1 U11830 ( .A1(n11849), .A2(n11850), .ZN(n11874) );
  OR2_X1 U11831 ( .A1(n11530), .A2(n7777), .ZN(n11850) );
  OR2_X1 U11832 ( .A1(n11875), .A2(n11876), .ZN(n11849) );
  AND2_X1 U11833 ( .A1(n11846), .A2(n11845), .ZN(n11876) );
  AND2_X1 U11834 ( .A1(n11843), .A2(n11877), .ZN(n11875) );
  OR2_X1 U11835 ( .A1(n11845), .A2(n11846), .ZN(n11877) );
  OR2_X1 U11836 ( .A1(n11530), .A2(n7785), .ZN(n11846) );
  OR2_X1 U11837 ( .A1(n11878), .A2(n11879), .ZN(n11845) );
  AND2_X1 U11838 ( .A1(n11842), .A2(n11841), .ZN(n11879) );
  AND2_X1 U11839 ( .A1(n11839), .A2(n11880), .ZN(n11878) );
  OR2_X1 U11840 ( .A1(n11841), .A2(n11842), .ZN(n11880) );
  OR2_X1 U11841 ( .A1(n11530), .A2(n8226), .ZN(n11842) );
  OR2_X1 U11842 ( .A1(n11881), .A2(n11882), .ZN(n11841) );
  AND2_X1 U11843 ( .A1(n11838), .A2(n11837), .ZN(n11882) );
  AND2_X1 U11844 ( .A1(n11835), .A2(n11883), .ZN(n11881) );
  OR2_X1 U11845 ( .A1(n11837), .A2(n11838), .ZN(n11883) );
  OR2_X1 U11846 ( .A1(n11530), .A2(n8221), .ZN(n11838) );
  OR2_X1 U11847 ( .A1(n11884), .A2(n11885), .ZN(n11837) );
  AND2_X1 U11848 ( .A1(n11834), .A2(n11833), .ZN(n11885) );
  AND2_X1 U11849 ( .A1(n11831), .A2(n11886), .ZN(n11884) );
  OR2_X1 U11850 ( .A1(n11833), .A2(n11834), .ZN(n11886) );
  OR2_X1 U11851 ( .A1(n11530), .A2(n8216), .ZN(n11834) );
  OR2_X1 U11852 ( .A1(n11887), .A2(n11888), .ZN(n11833) );
  AND2_X1 U11853 ( .A1(n11830), .A2(n11829), .ZN(n11888) );
  AND2_X1 U11854 ( .A1(n11827), .A2(n11889), .ZN(n11887) );
  OR2_X1 U11855 ( .A1(n11829), .A2(n11830), .ZN(n11889) );
  OR2_X1 U11856 ( .A1(n11530), .A2(n8211), .ZN(n11830) );
  OR2_X1 U11857 ( .A1(n11890), .A2(n11891), .ZN(n11829) );
  AND2_X1 U11858 ( .A1(n11826), .A2(n11825), .ZN(n11891) );
  AND2_X1 U11859 ( .A1(n11823), .A2(n11892), .ZN(n11890) );
  OR2_X1 U11860 ( .A1(n11825), .A2(n11826), .ZN(n11892) );
  OR2_X1 U11861 ( .A1(n11530), .A2(n8206), .ZN(n11826) );
  OR2_X1 U11862 ( .A1(n11893), .A2(n11894), .ZN(n11825) );
  AND2_X1 U11863 ( .A1(n11822), .A2(n11821), .ZN(n11894) );
  AND2_X1 U11864 ( .A1(n11819), .A2(n11895), .ZN(n11893) );
  OR2_X1 U11865 ( .A1(n11821), .A2(n11822), .ZN(n11895) );
  OR2_X1 U11866 ( .A1(n11530), .A2(n8201), .ZN(n11822) );
  OR2_X1 U11867 ( .A1(n11896), .A2(n11897), .ZN(n11821) );
  AND2_X1 U11868 ( .A1(n11818), .A2(n11817), .ZN(n11897) );
  AND2_X1 U11869 ( .A1(n11815), .A2(n11898), .ZN(n11896) );
  OR2_X1 U11870 ( .A1(n11817), .A2(n11818), .ZN(n11898) );
  OR2_X1 U11871 ( .A1(n11530), .A2(n8196), .ZN(n11818) );
  OR2_X1 U11872 ( .A1(n11899), .A2(n11900), .ZN(n11817) );
  AND2_X1 U11873 ( .A1(n11814), .A2(n11813), .ZN(n11900) );
  AND2_X1 U11874 ( .A1(n11811), .A2(n11901), .ZN(n11899) );
  OR2_X1 U11875 ( .A1(n11813), .A2(n11814), .ZN(n11901) );
  OR2_X1 U11876 ( .A1(n11530), .A2(n8191), .ZN(n11814) );
  OR2_X1 U11877 ( .A1(n11902), .A2(n11903), .ZN(n11813) );
  AND2_X1 U11878 ( .A1(n11808), .A2(n11810), .ZN(n11903) );
  AND2_X1 U11879 ( .A1(n11904), .A2(n11809), .ZN(n11902) );
  OR2_X1 U11880 ( .A1(n11808), .A2(n11810), .ZN(n11904) );
  OR2_X1 U11881 ( .A1(n11905), .A2(n11906), .ZN(n11810) );
  AND2_X1 U11882 ( .A1(n11806), .A2(n11805), .ZN(n11906) );
  AND2_X1 U11883 ( .A1(n11803), .A2(n11907), .ZN(n11905) );
  OR2_X1 U11884 ( .A1(n11805), .A2(n11806), .ZN(n11907) );
  OR2_X1 U11885 ( .A1(n11530), .A2(n8181), .ZN(n11806) );
  OR2_X1 U11886 ( .A1(n11908), .A2(n11909), .ZN(n11805) );
  AND2_X1 U11887 ( .A1(n11802), .A2(n11801), .ZN(n11909) );
  AND2_X1 U11888 ( .A1(n11799), .A2(n11910), .ZN(n11908) );
  OR2_X1 U11889 ( .A1(n11801), .A2(n11802), .ZN(n11910) );
  OR2_X1 U11890 ( .A1(n11530), .A2(n8176), .ZN(n11802) );
  OR2_X1 U11891 ( .A1(n11911), .A2(n11912), .ZN(n11801) );
  AND2_X1 U11892 ( .A1(n11798), .A2(n11797), .ZN(n11912) );
  AND2_X1 U11893 ( .A1(n11795), .A2(n11913), .ZN(n11911) );
  OR2_X1 U11894 ( .A1(n11797), .A2(n11798), .ZN(n11913) );
  OR2_X1 U11895 ( .A1(n11530), .A2(n8171), .ZN(n11798) );
  OR2_X1 U11896 ( .A1(n11914), .A2(n11915), .ZN(n11797) );
  AND2_X1 U11897 ( .A1(n11794), .A2(n11793), .ZN(n11915) );
  AND2_X1 U11898 ( .A1(n11791), .A2(n11916), .ZN(n11914) );
  OR2_X1 U11899 ( .A1(n11793), .A2(n11794), .ZN(n11916) );
  OR2_X1 U11900 ( .A1(n8166), .A2(n11530), .ZN(n11794) );
  OR2_X1 U11901 ( .A1(n11917), .A2(n11918), .ZN(n11793) );
  AND2_X1 U11902 ( .A1(n11790), .A2(n11789), .ZN(n11918) );
  AND2_X1 U11903 ( .A1(n11787), .A2(n11919), .ZN(n11917) );
  OR2_X1 U11904 ( .A1(n11789), .A2(n11790), .ZN(n11919) );
  OR2_X1 U11905 ( .A1(n11530), .A2(n8161), .ZN(n11790) );
  OR2_X1 U11906 ( .A1(n11920), .A2(n11921), .ZN(n11789) );
  AND2_X1 U11907 ( .A1(n11786), .A2(n11785), .ZN(n11921) );
  AND2_X1 U11908 ( .A1(n11783), .A2(n11922), .ZN(n11920) );
  OR2_X1 U11909 ( .A1(n11785), .A2(n11786), .ZN(n11922) );
  OR2_X1 U11910 ( .A1(n11530), .A2(n8156), .ZN(n11786) );
  OR2_X1 U11911 ( .A1(n11923), .A2(n11924), .ZN(n11785) );
  AND2_X1 U11912 ( .A1(n11782), .A2(n11781), .ZN(n11924) );
  AND2_X1 U11913 ( .A1(n11779), .A2(n11925), .ZN(n11923) );
  OR2_X1 U11914 ( .A1(n11781), .A2(n11782), .ZN(n11925) );
  OR2_X1 U11915 ( .A1(n11530), .A2(n8151), .ZN(n11782) );
  OR2_X1 U11916 ( .A1(n11926), .A2(n11927), .ZN(n11781) );
  AND2_X1 U11917 ( .A1(n11778), .A2(n11777), .ZN(n11927) );
  AND2_X1 U11918 ( .A1(n11775), .A2(n11928), .ZN(n11926) );
  OR2_X1 U11919 ( .A1(n11777), .A2(n11778), .ZN(n11928) );
  OR2_X1 U11920 ( .A1(n11530), .A2(n8146), .ZN(n11778) );
  OR2_X1 U11921 ( .A1(n11929), .A2(n11930), .ZN(n11777) );
  AND2_X1 U11922 ( .A1(n11774), .A2(n11773), .ZN(n11930) );
  AND2_X1 U11923 ( .A1(n11771), .A2(n11931), .ZN(n11929) );
  OR2_X1 U11924 ( .A1(n11773), .A2(n11774), .ZN(n11931) );
  OR2_X1 U11925 ( .A1(n11530), .A2(n8141), .ZN(n11774) );
  OR2_X1 U11926 ( .A1(n11932), .A2(n11933), .ZN(n11773) );
  AND2_X1 U11927 ( .A1(n11770), .A2(n11769), .ZN(n11933) );
  AND2_X1 U11928 ( .A1(n11767), .A2(n11934), .ZN(n11932) );
  OR2_X1 U11929 ( .A1(n11769), .A2(n11770), .ZN(n11934) );
  OR2_X1 U11930 ( .A1(n11530), .A2(n8136), .ZN(n11770) );
  OR2_X1 U11931 ( .A1(n11935), .A2(n11936), .ZN(n11769) );
  AND2_X1 U11932 ( .A1(n11766), .A2(n11765), .ZN(n11936) );
  AND2_X1 U11933 ( .A1(n11763), .A2(n11937), .ZN(n11935) );
  OR2_X1 U11934 ( .A1(n11765), .A2(n11766), .ZN(n11937) );
  OR2_X1 U11935 ( .A1(n11530), .A2(n8131), .ZN(n11766) );
  OR2_X1 U11936 ( .A1(n11938), .A2(n11939), .ZN(n11765) );
  AND2_X1 U11937 ( .A1(n11762), .A2(n11761), .ZN(n11939) );
  AND2_X1 U11938 ( .A1(n11759), .A2(n11940), .ZN(n11938) );
  OR2_X1 U11939 ( .A1(n11761), .A2(n11762), .ZN(n11940) );
  OR2_X1 U11940 ( .A1(n11530), .A2(n8126), .ZN(n11762) );
  OR2_X1 U11941 ( .A1(n11941), .A2(n11942), .ZN(n11761) );
  AND2_X1 U11942 ( .A1(n11758), .A2(n11757), .ZN(n11942) );
  AND2_X1 U11943 ( .A1(n11755), .A2(n11943), .ZN(n11941) );
  OR2_X1 U11944 ( .A1(n11757), .A2(n11758), .ZN(n11943) );
  OR2_X1 U11945 ( .A1(n11530), .A2(n8121), .ZN(n11758) );
  OR2_X1 U11946 ( .A1(n11944), .A2(n11945), .ZN(n11757) );
  AND2_X1 U11947 ( .A1(n11754), .A2(n11753), .ZN(n11945) );
  AND2_X1 U11948 ( .A1(n11751), .A2(n11946), .ZN(n11944) );
  OR2_X1 U11949 ( .A1(n11753), .A2(n11754), .ZN(n11946) );
  OR2_X1 U11950 ( .A1(n8116), .A2(n11530), .ZN(n11754) );
  OR2_X1 U11951 ( .A1(n11947), .A2(n11948), .ZN(n11753) );
  AND2_X1 U11952 ( .A1(n11750), .A2(n11749), .ZN(n11948) );
  AND2_X1 U11953 ( .A1(n11747), .A2(n11949), .ZN(n11947) );
  OR2_X1 U11954 ( .A1(n11749), .A2(n11750), .ZN(n11949) );
  OR2_X1 U11955 ( .A1(n8111), .A2(n11530), .ZN(n11750) );
  OR2_X1 U11956 ( .A1(n11950), .A2(n11951), .ZN(n11749) );
  AND2_X1 U11957 ( .A1(n11743), .A2(n11746), .ZN(n11951) );
  AND2_X1 U11958 ( .A1(n11745), .A2(n11952), .ZN(n11950) );
  OR2_X1 U11959 ( .A1(n11746), .A2(n11743), .ZN(n11952) );
  OR2_X1 U11960 ( .A1(n8102), .A2(n11530), .ZN(n11743) );
  OR3_X1 U11961 ( .A1(n8349), .A2(n11530), .A3(n11740), .ZN(n11746) );
  INV_X1 U11962 ( .A(n11953), .ZN(n11745) );
  OR2_X1 U11963 ( .A1(n11954), .A2(n11955), .ZN(n11953) );
  AND2_X1 U11964 ( .A1(b_12_), .A2(n11956), .ZN(n11955) );
  OR2_X1 U11965 ( .A1(n11957), .A2(n7314), .ZN(n11956) );
  AND2_X1 U11966 ( .A1(a_30_), .A2(n11958), .ZN(n11957) );
  AND2_X1 U11967 ( .A1(b_11_), .A2(n11959), .ZN(n11954) );
  OR2_X1 U11968 ( .A1(n11960), .A2(n7318), .ZN(n11959) );
  AND2_X1 U11969 ( .A1(a_31_), .A2(n11740), .ZN(n11960) );
  XNOR2_X1 U11970 ( .A(n11961), .B(n11962), .ZN(n11747) );
  XNOR2_X1 U11971 ( .A(n11963), .B(n11964), .ZN(n11962) );
  XOR2_X1 U11972 ( .A(n11965), .B(n11966), .Z(n11751) );
  XOR2_X1 U11973 ( .A(n11967), .B(n11968), .Z(n11966) );
  XOR2_X1 U11974 ( .A(n11969), .B(n11970), .Z(n11755) );
  XOR2_X1 U11975 ( .A(n11971), .B(n11972), .Z(n11970) );
  XOR2_X1 U11976 ( .A(n11973), .B(n11974), .Z(n11759) );
  XOR2_X1 U11977 ( .A(n11975), .B(n11976), .Z(n11974) );
  XOR2_X1 U11978 ( .A(n11977), .B(n11978), .Z(n11763) );
  XOR2_X1 U11979 ( .A(n11979), .B(n11980), .Z(n11978) );
  XOR2_X1 U11980 ( .A(n11981), .B(n11982), .Z(n11767) );
  XOR2_X1 U11981 ( .A(n11983), .B(n11984), .Z(n11982) );
  XOR2_X1 U11982 ( .A(n11985), .B(n11986), .Z(n11771) );
  XOR2_X1 U11983 ( .A(n11987), .B(n11988), .Z(n11986) );
  XOR2_X1 U11984 ( .A(n11989), .B(n11990), .Z(n11775) );
  XOR2_X1 U11985 ( .A(n11991), .B(n11992), .Z(n11990) );
  XOR2_X1 U11986 ( .A(n11993), .B(n11994), .Z(n11779) );
  XOR2_X1 U11987 ( .A(n11995), .B(n11996), .Z(n11994) );
  XOR2_X1 U11988 ( .A(n11997), .B(n11998), .Z(n11783) );
  XOR2_X1 U11989 ( .A(n11999), .B(n12000), .Z(n11998) );
  XOR2_X1 U11990 ( .A(n12001), .B(n12002), .Z(n11787) );
  XOR2_X1 U11991 ( .A(n12003), .B(n12004), .Z(n12002) );
  XOR2_X1 U11992 ( .A(n12005), .B(n12006), .Z(n11791) );
  XOR2_X1 U11993 ( .A(n12007), .B(n12008), .Z(n12006) );
  XOR2_X1 U11994 ( .A(n12009), .B(n12010), .Z(n11795) );
  XOR2_X1 U11995 ( .A(n12011), .B(n12012), .Z(n12010) );
  XOR2_X1 U11996 ( .A(n12013), .B(n12014), .Z(n11799) );
  XOR2_X1 U11997 ( .A(n12015), .B(n12016), .Z(n12014) );
  XOR2_X1 U11998 ( .A(n12017), .B(n12018), .Z(n11803) );
  XOR2_X1 U11999 ( .A(n12019), .B(n12020), .Z(n12018) );
  XOR2_X1 U12000 ( .A(n12021), .B(n12022), .Z(n11808) );
  XOR2_X1 U12001 ( .A(n12023), .B(n12024), .Z(n12022) );
  XOR2_X1 U12002 ( .A(n12025), .B(n12026), .Z(n11811) );
  XOR2_X1 U12003 ( .A(n12027), .B(n12028), .Z(n12026) );
  XNOR2_X1 U12004 ( .A(n12029), .B(n12030), .ZN(n11815) );
  XNOR2_X1 U12005 ( .A(n12031), .B(n12032), .ZN(n12029) );
  XOR2_X1 U12006 ( .A(n12033), .B(n12034), .Z(n11819) );
  XOR2_X1 U12007 ( .A(n12035), .B(n12036), .Z(n12034) );
  XOR2_X1 U12008 ( .A(n12037), .B(n12038), .Z(n11823) );
  XOR2_X1 U12009 ( .A(n12039), .B(n12040), .Z(n12038) );
  XOR2_X1 U12010 ( .A(n12041), .B(n12042), .Z(n11827) );
  XOR2_X1 U12011 ( .A(n12043), .B(n12044), .Z(n12042) );
  XOR2_X1 U12012 ( .A(n12045), .B(n12046), .Z(n11831) );
  XOR2_X1 U12013 ( .A(n12047), .B(n12048), .Z(n12046) );
  XOR2_X1 U12014 ( .A(n12049), .B(n12050), .Z(n11835) );
  XOR2_X1 U12015 ( .A(n12051), .B(n12052), .Z(n12050) );
  XOR2_X1 U12016 ( .A(n12053), .B(n12054), .Z(n11839) );
  XOR2_X1 U12017 ( .A(n12055), .B(n12056), .Z(n12054) );
  XOR2_X1 U12018 ( .A(n12057), .B(n12058), .Z(n11843) );
  XOR2_X1 U12019 ( .A(n12059), .B(n12060), .Z(n12058) );
  XOR2_X1 U12020 ( .A(n12061), .B(n12062), .Z(n11847) );
  XOR2_X1 U12021 ( .A(n12063), .B(n12064), .Z(n12062) );
  XOR2_X1 U12022 ( .A(n12065), .B(n12066), .Z(n11851) );
  XOR2_X1 U12023 ( .A(n12067), .B(n12068), .Z(n12066) );
  XOR2_X1 U12024 ( .A(n12069), .B(n12070), .Z(n11855) );
  XOR2_X1 U12025 ( .A(n12071), .B(n12072), .Z(n12070) );
  XOR2_X1 U12026 ( .A(n12073), .B(n12074), .Z(n11859) );
  XOR2_X1 U12027 ( .A(n12075), .B(n12076), .Z(n12074) );
  XNOR2_X1 U12028 ( .A(n12077), .B(n12078), .ZN(n7570) );
  XOR2_X1 U12029 ( .A(n12079), .B(n12080), .Z(n12078) );
  XNOR2_X1 U12030 ( .A(n7579), .B(n7803), .ZN(n7568) );
  OR2_X1 U12031 ( .A1(n12081), .A2(n12082), .ZN(n7803) );
  AND2_X1 U12032 ( .A1(n12080), .A2(n12079), .ZN(n12082) );
  AND2_X1 U12033 ( .A1(n12077), .A2(n12083), .ZN(n12081) );
  OR2_X1 U12034 ( .A1(n12079), .A2(n12080), .ZN(n12083) );
  OR2_X1 U12035 ( .A1(n11740), .A2(n7621), .ZN(n12080) );
  OR2_X1 U12036 ( .A1(n12084), .A2(n12085), .ZN(n12079) );
  AND2_X1 U12037 ( .A1(n12076), .A2(n12075), .ZN(n12085) );
  AND2_X1 U12038 ( .A1(n12073), .A2(n12086), .ZN(n12084) );
  OR2_X1 U12039 ( .A1(n12075), .A2(n12076), .ZN(n12086) );
  OR2_X1 U12040 ( .A1(n11740), .A2(n7656), .ZN(n12076) );
  OR2_X1 U12041 ( .A1(n12087), .A2(n12088), .ZN(n12075) );
  AND2_X1 U12042 ( .A1(n12072), .A2(n12071), .ZN(n12088) );
  AND2_X1 U12043 ( .A1(n12069), .A2(n12089), .ZN(n12087) );
  OR2_X1 U12044 ( .A1(n12071), .A2(n12072), .ZN(n12089) );
  OR2_X1 U12045 ( .A1(n11740), .A2(n7689), .ZN(n12072) );
  OR2_X1 U12046 ( .A1(n12090), .A2(n12091), .ZN(n12071) );
  AND2_X1 U12047 ( .A1(n12068), .A2(n12067), .ZN(n12091) );
  AND2_X1 U12048 ( .A1(n12065), .A2(n12092), .ZN(n12090) );
  OR2_X1 U12049 ( .A1(n12067), .A2(n12068), .ZN(n12092) );
  OR2_X1 U12050 ( .A1(n11740), .A2(n7777), .ZN(n12068) );
  OR2_X1 U12051 ( .A1(n12093), .A2(n12094), .ZN(n12067) );
  AND2_X1 U12052 ( .A1(n12064), .A2(n12063), .ZN(n12094) );
  AND2_X1 U12053 ( .A1(n12061), .A2(n12095), .ZN(n12093) );
  OR2_X1 U12054 ( .A1(n12063), .A2(n12064), .ZN(n12095) );
  OR2_X1 U12055 ( .A1(n11740), .A2(n7785), .ZN(n12064) );
  OR2_X1 U12056 ( .A1(n12096), .A2(n12097), .ZN(n12063) );
  AND2_X1 U12057 ( .A1(n12060), .A2(n12059), .ZN(n12097) );
  AND2_X1 U12058 ( .A1(n12057), .A2(n12098), .ZN(n12096) );
  OR2_X1 U12059 ( .A1(n12059), .A2(n12060), .ZN(n12098) );
  OR2_X1 U12060 ( .A1(n11740), .A2(n8226), .ZN(n12060) );
  OR2_X1 U12061 ( .A1(n12099), .A2(n12100), .ZN(n12059) );
  AND2_X1 U12062 ( .A1(n12056), .A2(n12055), .ZN(n12100) );
  AND2_X1 U12063 ( .A1(n12053), .A2(n12101), .ZN(n12099) );
  OR2_X1 U12064 ( .A1(n12055), .A2(n12056), .ZN(n12101) );
  OR2_X1 U12065 ( .A1(n11740), .A2(n8221), .ZN(n12056) );
  OR2_X1 U12066 ( .A1(n12102), .A2(n12103), .ZN(n12055) );
  AND2_X1 U12067 ( .A1(n12052), .A2(n12051), .ZN(n12103) );
  AND2_X1 U12068 ( .A1(n12049), .A2(n12104), .ZN(n12102) );
  OR2_X1 U12069 ( .A1(n12051), .A2(n12052), .ZN(n12104) );
  OR2_X1 U12070 ( .A1(n11740), .A2(n8216), .ZN(n12052) );
  OR2_X1 U12071 ( .A1(n12105), .A2(n12106), .ZN(n12051) );
  AND2_X1 U12072 ( .A1(n12048), .A2(n12047), .ZN(n12106) );
  AND2_X1 U12073 ( .A1(n12045), .A2(n12107), .ZN(n12105) );
  OR2_X1 U12074 ( .A1(n12047), .A2(n12048), .ZN(n12107) );
  OR2_X1 U12075 ( .A1(n11740), .A2(n8211), .ZN(n12048) );
  OR2_X1 U12076 ( .A1(n12108), .A2(n12109), .ZN(n12047) );
  AND2_X1 U12077 ( .A1(n12044), .A2(n12043), .ZN(n12109) );
  AND2_X1 U12078 ( .A1(n12041), .A2(n12110), .ZN(n12108) );
  OR2_X1 U12079 ( .A1(n12043), .A2(n12044), .ZN(n12110) );
  OR2_X1 U12080 ( .A1(n11740), .A2(n8206), .ZN(n12044) );
  OR2_X1 U12081 ( .A1(n12111), .A2(n12112), .ZN(n12043) );
  AND2_X1 U12082 ( .A1(n12040), .A2(n12039), .ZN(n12112) );
  AND2_X1 U12083 ( .A1(n12037), .A2(n12113), .ZN(n12111) );
  OR2_X1 U12084 ( .A1(n12039), .A2(n12040), .ZN(n12113) );
  OR2_X1 U12085 ( .A1(n11740), .A2(n8201), .ZN(n12040) );
  OR2_X1 U12086 ( .A1(n12114), .A2(n12115), .ZN(n12039) );
  AND2_X1 U12087 ( .A1(n12036), .A2(n12035), .ZN(n12115) );
  AND2_X1 U12088 ( .A1(n12033), .A2(n12116), .ZN(n12114) );
  OR2_X1 U12089 ( .A1(n12035), .A2(n12036), .ZN(n12116) );
  OR2_X1 U12090 ( .A1(n11740), .A2(n8196), .ZN(n12036) );
  OR2_X1 U12091 ( .A1(n12117), .A2(n12118), .ZN(n12035) );
  AND2_X1 U12092 ( .A1(n12030), .A2(n12032), .ZN(n12118) );
  AND2_X1 U12093 ( .A1(n12119), .A2(n12031), .ZN(n12117) );
  OR2_X1 U12094 ( .A1(n12030), .A2(n12032), .ZN(n12119) );
  OR2_X1 U12095 ( .A1(n12120), .A2(n12121), .ZN(n12032) );
  AND2_X1 U12096 ( .A1(n12028), .A2(n12027), .ZN(n12121) );
  AND2_X1 U12097 ( .A1(n12025), .A2(n12122), .ZN(n12120) );
  OR2_X1 U12098 ( .A1(n12027), .A2(n12028), .ZN(n12122) );
  OR2_X1 U12099 ( .A1(n11740), .A2(n8186), .ZN(n12028) );
  OR2_X1 U12100 ( .A1(n12123), .A2(n12124), .ZN(n12027) );
  AND2_X1 U12101 ( .A1(n12024), .A2(n12023), .ZN(n12124) );
  AND2_X1 U12102 ( .A1(n12021), .A2(n12125), .ZN(n12123) );
  OR2_X1 U12103 ( .A1(n12023), .A2(n12024), .ZN(n12125) );
  OR2_X1 U12104 ( .A1(n11740), .A2(n8181), .ZN(n12024) );
  OR2_X1 U12105 ( .A1(n12126), .A2(n12127), .ZN(n12023) );
  AND2_X1 U12106 ( .A1(n12020), .A2(n12019), .ZN(n12127) );
  AND2_X1 U12107 ( .A1(n12017), .A2(n12128), .ZN(n12126) );
  OR2_X1 U12108 ( .A1(n12019), .A2(n12020), .ZN(n12128) );
  OR2_X1 U12109 ( .A1(n11740), .A2(n8176), .ZN(n12020) );
  OR2_X1 U12110 ( .A1(n12129), .A2(n12130), .ZN(n12019) );
  AND2_X1 U12111 ( .A1(n12016), .A2(n12015), .ZN(n12130) );
  AND2_X1 U12112 ( .A1(n12013), .A2(n12131), .ZN(n12129) );
  OR2_X1 U12113 ( .A1(n12015), .A2(n12016), .ZN(n12131) );
  OR2_X1 U12114 ( .A1(n11740), .A2(n8171), .ZN(n12016) );
  OR2_X1 U12115 ( .A1(n12132), .A2(n12133), .ZN(n12015) );
  AND2_X1 U12116 ( .A1(n12012), .A2(n12011), .ZN(n12133) );
  AND2_X1 U12117 ( .A1(n12009), .A2(n12134), .ZN(n12132) );
  OR2_X1 U12118 ( .A1(n12011), .A2(n12012), .ZN(n12134) );
  OR2_X1 U12119 ( .A1(n8166), .A2(n11740), .ZN(n12012) );
  OR2_X1 U12120 ( .A1(n12135), .A2(n12136), .ZN(n12011) );
  AND2_X1 U12121 ( .A1(n12008), .A2(n12007), .ZN(n12136) );
  AND2_X1 U12122 ( .A1(n12005), .A2(n12137), .ZN(n12135) );
  OR2_X1 U12123 ( .A1(n12007), .A2(n12008), .ZN(n12137) );
  OR2_X1 U12124 ( .A1(n11740), .A2(n8161), .ZN(n12008) );
  OR2_X1 U12125 ( .A1(n12138), .A2(n12139), .ZN(n12007) );
  AND2_X1 U12126 ( .A1(n12004), .A2(n12003), .ZN(n12139) );
  AND2_X1 U12127 ( .A1(n12001), .A2(n12140), .ZN(n12138) );
  OR2_X1 U12128 ( .A1(n12003), .A2(n12004), .ZN(n12140) );
  OR2_X1 U12129 ( .A1(n11740), .A2(n8156), .ZN(n12004) );
  OR2_X1 U12130 ( .A1(n12141), .A2(n12142), .ZN(n12003) );
  AND2_X1 U12131 ( .A1(n12000), .A2(n11999), .ZN(n12142) );
  AND2_X1 U12132 ( .A1(n11997), .A2(n12143), .ZN(n12141) );
  OR2_X1 U12133 ( .A1(n11999), .A2(n12000), .ZN(n12143) );
  OR2_X1 U12134 ( .A1(n11740), .A2(n8151), .ZN(n12000) );
  OR2_X1 U12135 ( .A1(n12144), .A2(n12145), .ZN(n11999) );
  AND2_X1 U12136 ( .A1(n11996), .A2(n11995), .ZN(n12145) );
  AND2_X1 U12137 ( .A1(n11993), .A2(n12146), .ZN(n12144) );
  OR2_X1 U12138 ( .A1(n11995), .A2(n11996), .ZN(n12146) );
  OR2_X1 U12139 ( .A1(n11740), .A2(n8146), .ZN(n11996) );
  OR2_X1 U12140 ( .A1(n12147), .A2(n12148), .ZN(n11995) );
  AND2_X1 U12141 ( .A1(n11992), .A2(n11991), .ZN(n12148) );
  AND2_X1 U12142 ( .A1(n11989), .A2(n12149), .ZN(n12147) );
  OR2_X1 U12143 ( .A1(n11991), .A2(n11992), .ZN(n12149) );
  OR2_X1 U12144 ( .A1(n11740), .A2(n8141), .ZN(n11992) );
  OR2_X1 U12145 ( .A1(n12150), .A2(n12151), .ZN(n11991) );
  AND2_X1 U12146 ( .A1(n11988), .A2(n11987), .ZN(n12151) );
  AND2_X1 U12147 ( .A1(n11985), .A2(n12152), .ZN(n12150) );
  OR2_X1 U12148 ( .A1(n11987), .A2(n11988), .ZN(n12152) );
  OR2_X1 U12149 ( .A1(n11740), .A2(n8136), .ZN(n11988) );
  OR2_X1 U12150 ( .A1(n12153), .A2(n12154), .ZN(n11987) );
  AND2_X1 U12151 ( .A1(n11984), .A2(n11983), .ZN(n12154) );
  AND2_X1 U12152 ( .A1(n11981), .A2(n12155), .ZN(n12153) );
  OR2_X1 U12153 ( .A1(n11983), .A2(n11984), .ZN(n12155) );
  OR2_X1 U12154 ( .A1(n11740), .A2(n8131), .ZN(n11984) );
  OR2_X1 U12155 ( .A1(n12156), .A2(n12157), .ZN(n11983) );
  AND2_X1 U12156 ( .A1(n11980), .A2(n11979), .ZN(n12157) );
  AND2_X1 U12157 ( .A1(n11977), .A2(n12158), .ZN(n12156) );
  OR2_X1 U12158 ( .A1(n11979), .A2(n11980), .ZN(n12158) );
  OR2_X1 U12159 ( .A1(n11740), .A2(n8126), .ZN(n11980) );
  OR2_X1 U12160 ( .A1(n12159), .A2(n12160), .ZN(n11979) );
  AND2_X1 U12161 ( .A1(n11976), .A2(n11975), .ZN(n12160) );
  AND2_X1 U12162 ( .A1(n11973), .A2(n12161), .ZN(n12159) );
  OR2_X1 U12163 ( .A1(n11975), .A2(n11976), .ZN(n12161) );
  OR2_X1 U12164 ( .A1(n8121), .A2(n11740), .ZN(n11976) );
  OR2_X1 U12165 ( .A1(n12162), .A2(n12163), .ZN(n11975) );
  AND2_X1 U12166 ( .A1(n11972), .A2(n11971), .ZN(n12163) );
  AND2_X1 U12167 ( .A1(n11969), .A2(n12164), .ZN(n12162) );
  OR2_X1 U12168 ( .A1(n11971), .A2(n11972), .ZN(n12164) );
  OR2_X1 U12169 ( .A1(n8116), .A2(n11740), .ZN(n11972) );
  OR2_X1 U12170 ( .A1(n12165), .A2(n12166), .ZN(n11971) );
  AND2_X1 U12171 ( .A1(n11968), .A2(n11967), .ZN(n12166) );
  AND2_X1 U12172 ( .A1(n11965), .A2(n12167), .ZN(n12165) );
  OR2_X1 U12173 ( .A1(n11967), .A2(n11968), .ZN(n12167) );
  OR2_X1 U12174 ( .A1(n8111), .A2(n11740), .ZN(n11968) );
  OR2_X1 U12175 ( .A1(n12168), .A2(n12169), .ZN(n11967) );
  AND2_X1 U12176 ( .A1(n11961), .A2(n11964), .ZN(n12169) );
  AND2_X1 U12177 ( .A1(n11963), .A2(n12170), .ZN(n12168) );
  OR2_X1 U12178 ( .A1(n11964), .A2(n11961), .ZN(n12170) );
  OR2_X1 U12179 ( .A1(n8102), .A2(n11740), .ZN(n11961) );
  OR3_X1 U12180 ( .A1(n8349), .A2(n11740), .A3(n11958), .ZN(n11964) );
  INV_X1 U12181 ( .A(n12171), .ZN(n11963) );
  OR2_X1 U12182 ( .A1(n12172), .A2(n12173), .ZN(n12171) );
  AND2_X1 U12183 ( .A1(b_11_), .A2(n12174), .ZN(n12173) );
  OR2_X1 U12184 ( .A1(n12175), .A2(n7314), .ZN(n12174) );
  AND2_X1 U12185 ( .A1(a_30_), .A2(n12176), .ZN(n12175) );
  AND2_X1 U12186 ( .A1(b_10_), .A2(n12177), .ZN(n12172) );
  OR2_X1 U12187 ( .A1(n12178), .A2(n7318), .ZN(n12177) );
  AND2_X1 U12188 ( .A1(a_31_), .A2(n11958), .ZN(n12178) );
  XNOR2_X1 U12189 ( .A(n12179), .B(n12180), .ZN(n11965) );
  XNOR2_X1 U12190 ( .A(n12181), .B(n12182), .ZN(n12180) );
  XNOR2_X1 U12191 ( .A(n12183), .B(n12184), .ZN(n11969) );
  XNOR2_X1 U12192 ( .A(n12185), .B(n12186), .ZN(n12183) );
  XOR2_X1 U12193 ( .A(n12187), .B(n12188), .Z(n11973) );
  XOR2_X1 U12194 ( .A(n12189), .B(n12190), .Z(n12188) );
  XOR2_X1 U12195 ( .A(n12191), .B(n12192), .Z(n11977) );
  XOR2_X1 U12196 ( .A(n12193), .B(n12194), .Z(n12192) );
  XOR2_X1 U12197 ( .A(n12195), .B(n12196), .Z(n11981) );
  XOR2_X1 U12198 ( .A(n12197), .B(n12198), .Z(n12196) );
  XOR2_X1 U12199 ( .A(n12199), .B(n12200), .Z(n11985) );
  XOR2_X1 U12200 ( .A(n12201), .B(n12202), .Z(n12200) );
  XOR2_X1 U12201 ( .A(n12203), .B(n12204), .Z(n11989) );
  XOR2_X1 U12202 ( .A(n12205), .B(n12206), .Z(n12204) );
  XOR2_X1 U12203 ( .A(n12207), .B(n12208), .Z(n11993) );
  XOR2_X1 U12204 ( .A(n12209), .B(n12210), .Z(n12208) );
  XOR2_X1 U12205 ( .A(n12211), .B(n12212), .Z(n11997) );
  XOR2_X1 U12206 ( .A(n12213), .B(n12214), .Z(n12212) );
  XOR2_X1 U12207 ( .A(n12215), .B(n12216), .Z(n12001) );
  XOR2_X1 U12208 ( .A(n12217), .B(n12218), .Z(n12216) );
  XOR2_X1 U12209 ( .A(n12219), .B(n12220), .Z(n12005) );
  XOR2_X1 U12210 ( .A(n12221), .B(n12222), .Z(n12220) );
  XOR2_X1 U12211 ( .A(n12223), .B(n12224), .Z(n12009) );
  XOR2_X1 U12212 ( .A(n12225), .B(n12226), .Z(n12224) );
  XOR2_X1 U12213 ( .A(n12227), .B(n12228), .Z(n12013) );
  XOR2_X1 U12214 ( .A(n12229), .B(n12230), .Z(n12228) );
  XOR2_X1 U12215 ( .A(n12231), .B(n12232), .Z(n12017) );
  XOR2_X1 U12216 ( .A(n12233), .B(n12234), .Z(n12232) );
  XOR2_X1 U12217 ( .A(n12235), .B(n12236), .Z(n12021) );
  XOR2_X1 U12218 ( .A(n12237), .B(n12238), .Z(n12236) );
  XOR2_X1 U12219 ( .A(n12239), .B(n12240), .Z(n12025) );
  XOR2_X1 U12220 ( .A(n12241), .B(n12242), .Z(n12240) );
  XOR2_X1 U12221 ( .A(n12243), .B(n12244), .Z(n12030) );
  XOR2_X1 U12222 ( .A(n12245), .B(n12246), .Z(n12244) );
  XOR2_X1 U12223 ( .A(n12247), .B(n12248), .Z(n12033) );
  XOR2_X1 U12224 ( .A(n12249), .B(n12250), .Z(n12248) );
  XNOR2_X1 U12225 ( .A(n12251), .B(n12252), .ZN(n12037) );
  XNOR2_X1 U12226 ( .A(n12253), .B(n12254), .ZN(n12251) );
  XOR2_X1 U12227 ( .A(n12255), .B(n12256), .Z(n12041) );
  XOR2_X1 U12228 ( .A(n12257), .B(n12258), .Z(n12256) );
  XOR2_X1 U12229 ( .A(n12259), .B(n12260), .Z(n12045) );
  XOR2_X1 U12230 ( .A(n12261), .B(n12262), .Z(n12260) );
  XOR2_X1 U12231 ( .A(n12263), .B(n12264), .Z(n12049) );
  XOR2_X1 U12232 ( .A(n12265), .B(n12266), .Z(n12264) );
  XOR2_X1 U12233 ( .A(n12267), .B(n12268), .Z(n12053) );
  XOR2_X1 U12234 ( .A(n12269), .B(n12270), .Z(n12268) );
  XOR2_X1 U12235 ( .A(n12271), .B(n12272), .Z(n12057) );
  XOR2_X1 U12236 ( .A(n12273), .B(n12274), .Z(n12272) );
  XOR2_X1 U12237 ( .A(n12275), .B(n12276), .Z(n12061) );
  XOR2_X1 U12238 ( .A(n12277), .B(n12278), .Z(n12276) );
  XOR2_X1 U12239 ( .A(n12279), .B(n12280), .Z(n12065) );
  XOR2_X1 U12240 ( .A(n12281), .B(n12282), .Z(n12280) );
  XOR2_X1 U12241 ( .A(n12283), .B(n12284), .Z(n12069) );
  XOR2_X1 U12242 ( .A(n12285), .B(n12286), .Z(n12284) );
  XOR2_X1 U12243 ( .A(n12287), .B(n12288), .Z(n12073) );
  XOR2_X1 U12244 ( .A(n12289), .B(n12290), .Z(n12288) );
  XOR2_X1 U12245 ( .A(n12291), .B(n12292), .Z(n12077) );
  XOR2_X1 U12246 ( .A(n12293), .B(n12294), .Z(n12292) );
  XNOR2_X1 U12247 ( .A(n12295), .B(n12296), .ZN(n7579) );
  XOR2_X1 U12248 ( .A(n12297), .B(n12298), .Z(n12296) );
  XNOR2_X1 U12249 ( .A(n7588), .B(n7801), .ZN(n7577) );
  OR2_X1 U12250 ( .A1(n12299), .A2(n12300), .ZN(n7801) );
  AND2_X1 U12251 ( .A1(n12298), .A2(n12297), .ZN(n12300) );
  AND2_X1 U12252 ( .A1(n12295), .A2(n12301), .ZN(n12299) );
  OR2_X1 U12253 ( .A1(n12297), .A2(n12298), .ZN(n12301) );
  OR2_X1 U12254 ( .A1(n11958), .A2(n7621), .ZN(n12298) );
  OR2_X1 U12255 ( .A1(n12302), .A2(n12303), .ZN(n12297) );
  AND2_X1 U12256 ( .A1(n12294), .A2(n12293), .ZN(n12303) );
  AND2_X1 U12257 ( .A1(n12291), .A2(n12304), .ZN(n12302) );
  OR2_X1 U12258 ( .A1(n12293), .A2(n12294), .ZN(n12304) );
  OR2_X1 U12259 ( .A1(n11958), .A2(n7656), .ZN(n12294) );
  OR2_X1 U12260 ( .A1(n12305), .A2(n12306), .ZN(n12293) );
  AND2_X1 U12261 ( .A1(n12290), .A2(n12289), .ZN(n12306) );
  AND2_X1 U12262 ( .A1(n12287), .A2(n12307), .ZN(n12305) );
  OR2_X1 U12263 ( .A1(n12289), .A2(n12290), .ZN(n12307) );
  OR2_X1 U12264 ( .A1(n11958), .A2(n7689), .ZN(n12290) );
  OR2_X1 U12265 ( .A1(n12308), .A2(n12309), .ZN(n12289) );
  AND2_X1 U12266 ( .A1(n12286), .A2(n12285), .ZN(n12309) );
  AND2_X1 U12267 ( .A1(n12283), .A2(n12310), .ZN(n12308) );
  OR2_X1 U12268 ( .A1(n12285), .A2(n12286), .ZN(n12310) );
  OR2_X1 U12269 ( .A1(n11958), .A2(n7777), .ZN(n12286) );
  OR2_X1 U12270 ( .A1(n12311), .A2(n12312), .ZN(n12285) );
  AND2_X1 U12271 ( .A1(n12282), .A2(n12281), .ZN(n12312) );
  AND2_X1 U12272 ( .A1(n12279), .A2(n12313), .ZN(n12311) );
  OR2_X1 U12273 ( .A1(n12281), .A2(n12282), .ZN(n12313) );
  OR2_X1 U12274 ( .A1(n11958), .A2(n7785), .ZN(n12282) );
  OR2_X1 U12275 ( .A1(n12314), .A2(n12315), .ZN(n12281) );
  AND2_X1 U12276 ( .A1(n12278), .A2(n12277), .ZN(n12315) );
  AND2_X1 U12277 ( .A1(n12275), .A2(n12316), .ZN(n12314) );
  OR2_X1 U12278 ( .A1(n12277), .A2(n12278), .ZN(n12316) );
  OR2_X1 U12279 ( .A1(n11958), .A2(n8226), .ZN(n12278) );
  OR2_X1 U12280 ( .A1(n12317), .A2(n12318), .ZN(n12277) );
  AND2_X1 U12281 ( .A1(n12274), .A2(n12273), .ZN(n12318) );
  AND2_X1 U12282 ( .A1(n12271), .A2(n12319), .ZN(n12317) );
  OR2_X1 U12283 ( .A1(n12273), .A2(n12274), .ZN(n12319) );
  OR2_X1 U12284 ( .A1(n11958), .A2(n8221), .ZN(n12274) );
  OR2_X1 U12285 ( .A1(n12320), .A2(n12321), .ZN(n12273) );
  AND2_X1 U12286 ( .A1(n12270), .A2(n12269), .ZN(n12321) );
  AND2_X1 U12287 ( .A1(n12267), .A2(n12322), .ZN(n12320) );
  OR2_X1 U12288 ( .A1(n12269), .A2(n12270), .ZN(n12322) );
  OR2_X1 U12289 ( .A1(n11958), .A2(n8216), .ZN(n12270) );
  OR2_X1 U12290 ( .A1(n12323), .A2(n12324), .ZN(n12269) );
  AND2_X1 U12291 ( .A1(n12266), .A2(n12265), .ZN(n12324) );
  AND2_X1 U12292 ( .A1(n12263), .A2(n12325), .ZN(n12323) );
  OR2_X1 U12293 ( .A1(n12265), .A2(n12266), .ZN(n12325) );
  OR2_X1 U12294 ( .A1(n11958), .A2(n8211), .ZN(n12266) );
  OR2_X1 U12295 ( .A1(n12326), .A2(n12327), .ZN(n12265) );
  AND2_X1 U12296 ( .A1(n12262), .A2(n12261), .ZN(n12327) );
  AND2_X1 U12297 ( .A1(n12259), .A2(n12328), .ZN(n12326) );
  OR2_X1 U12298 ( .A1(n12261), .A2(n12262), .ZN(n12328) );
  OR2_X1 U12299 ( .A1(n11958), .A2(n8206), .ZN(n12262) );
  OR2_X1 U12300 ( .A1(n12329), .A2(n12330), .ZN(n12261) );
  AND2_X1 U12301 ( .A1(n12258), .A2(n12257), .ZN(n12330) );
  AND2_X1 U12302 ( .A1(n12255), .A2(n12331), .ZN(n12329) );
  OR2_X1 U12303 ( .A1(n12257), .A2(n12258), .ZN(n12331) );
  OR2_X1 U12304 ( .A1(n11958), .A2(n8201), .ZN(n12258) );
  OR2_X1 U12305 ( .A1(n12332), .A2(n12333), .ZN(n12257) );
  AND2_X1 U12306 ( .A1(n12252), .A2(n12254), .ZN(n12333) );
  AND2_X1 U12307 ( .A1(n12334), .A2(n12253), .ZN(n12332) );
  OR2_X1 U12308 ( .A1(n12252), .A2(n12254), .ZN(n12334) );
  OR2_X1 U12309 ( .A1(n12335), .A2(n12336), .ZN(n12254) );
  AND2_X1 U12310 ( .A1(n12250), .A2(n12249), .ZN(n12336) );
  AND2_X1 U12311 ( .A1(n12247), .A2(n12337), .ZN(n12335) );
  OR2_X1 U12312 ( .A1(n12249), .A2(n12250), .ZN(n12337) );
  OR2_X1 U12313 ( .A1(n11958), .A2(n8191), .ZN(n12250) );
  OR2_X1 U12314 ( .A1(n12338), .A2(n12339), .ZN(n12249) );
  AND2_X1 U12315 ( .A1(n12246), .A2(n12245), .ZN(n12339) );
  AND2_X1 U12316 ( .A1(n12243), .A2(n12340), .ZN(n12338) );
  OR2_X1 U12317 ( .A1(n12245), .A2(n12246), .ZN(n12340) );
  OR2_X1 U12318 ( .A1(n11958), .A2(n8186), .ZN(n12246) );
  OR2_X1 U12319 ( .A1(n12341), .A2(n12342), .ZN(n12245) );
  AND2_X1 U12320 ( .A1(n12242), .A2(n12241), .ZN(n12342) );
  AND2_X1 U12321 ( .A1(n12239), .A2(n12343), .ZN(n12341) );
  OR2_X1 U12322 ( .A1(n12241), .A2(n12242), .ZN(n12343) );
  OR2_X1 U12323 ( .A1(n11958), .A2(n8181), .ZN(n12242) );
  OR2_X1 U12324 ( .A1(n12344), .A2(n12345), .ZN(n12241) );
  AND2_X1 U12325 ( .A1(n12238), .A2(n12237), .ZN(n12345) );
  AND2_X1 U12326 ( .A1(n12235), .A2(n12346), .ZN(n12344) );
  OR2_X1 U12327 ( .A1(n12237), .A2(n12238), .ZN(n12346) );
  OR2_X1 U12328 ( .A1(n11958), .A2(n8176), .ZN(n12238) );
  OR2_X1 U12329 ( .A1(n12347), .A2(n12348), .ZN(n12237) );
  AND2_X1 U12330 ( .A1(n12234), .A2(n12233), .ZN(n12348) );
  AND2_X1 U12331 ( .A1(n12231), .A2(n12349), .ZN(n12347) );
  OR2_X1 U12332 ( .A1(n12233), .A2(n12234), .ZN(n12349) );
  OR2_X1 U12333 ( .A1(n11958), .A2(n8171), .ZN(n12234) );
  OR2_X1 U12334 ( .A1(n12350), .A2(n12351), .ZN(n12233) );
  AND2_X1 U12335 ( .A1(n12230), .A2(n12229), .ZN(n12351) );
  AND2_X1 U12336 ( .A1(n12227), .A2(n12352), .ZN(n12350) );
  OR2_X1 U12337 ( .A1(n12229), .A2(n12230), .ZN(n12352) );
  OR2_X1 U12338 ( .A1(n8166), .A2(n11958), .ZN(n12230) );
  OR2_X1 U12339 ( .A1(n12353), .A2(n12354), .ZN(n12229) );
  AND2_X1 U12340 ( .A1(n12226), .A2(n12225), .ZN(n12354) );
  AND2_X1 U12341 ( .A1(n12223), .A2(n12355), .ZN(n12353) );
  OR2_X1 U12342 ( .A1(n12225), .A2(n12226), .ZN(n12355) );
  OR2_X1 U12343 ( .A1(n11958), .A2(n8161), .ZN(n12226) );
  OR2_X1 U12344 ( .A1(n12356), .A2(n12357), .ZN(n12225) );
  AND2_X1 U12345 ( .A1(n12222), .A2(n12221), .ZN(n12357) );
  AND2_X1 U12346 ( .A1(n12219), .A2(n12358), .ZN(n12356) );
  OR2_X1 U12347 ( .A1(n12221), .A2(n12222), .ZN(n12358) );
  OR2_X1 U12348 ( .A1(n11958), .A2(n8156), .ZN(n12222) );
  OR2_X1 U12349 ( .A1(n12359), .A2(n12360), .ZN(n12221) );
  AND2_X1 U12350 ( .A1(n12218), .A2(n12217), .ZN(n12360) );
  AND2_X1 U12351 ( .A1(n12215), .A2(n12361), .ZN(n12359) );
  OR2_X1 U12352 ( .A1(n12217), .A2(n12218), .ZN(n12361) );
  OR2_X1 U12353 ( .A1(n11958), .A2(n8151), .ZN(n12218) );
  OR2_X1 U12354 ( .A1(n12362), .A2(n12363), .ZN(n12217) );
  AND2_X1 U12355 ( .A1(n12214), .A2(n12213), .ZN(n12363) );
  AND2_X1 U12356 ( .A1(n12211), .A2(n12364), .ZN(n12362) );
  OR2_X1 U12357 ( .A1(n12213), .A2(n12214), .ZN(n12364) );
  OR2_X1 U12358 ( .A1(n11958), .A2(n8146), .ZN(n12214) );
  OR2_X1 U12359 ( .A1(n12365), .A2(n12366), .ZN(n12213) );
  AND2_X1 U12360 ( .A1(n12210), .A2(n12209), .ZN(n12366) );
  AND2_X1 U12361 ( .A1(n12207), .A2(n12367), .ZN(n12365) );
  OR2_X1 U12362 ( .A1(n12209), .A2(n12210), .ZN(n12367) );
  OR2_X1 U12363 ( .A1(n11958), .A2(n8141), .ZN(n12210) );
  OR2_X1 U12364 ( .A1(n12368), .A2(n12369), .ZN(n12209) );
  AND2_X1 U12365 ( .A1(n12206), .A2(n12205), .ZN(n12369) );
  AND2_X1 U12366 ( .A1(n12203), .A2(n12370), .ZN(n12368) );
  OR2_X1 U12367 ( .A1(n12205), .A2(n12206), .ZN(n12370) );
  OR2_X1 U12368 ( .A1(n11958), .A2(n8136), .ZN(n12206) );
  OR2_X1 U12369 ( .A1(n12371), .A2(n12372), .ZN(n12205) );
  AND2_X1 U12370 ( .A1(n12202), .A2(n12201), .ZN(n12372) );
  AND2_X1 U12371 ( .A1(n12199), .A2(n12373), .ZN(n12371) );
  OR2_X1 U12372 ( .A1(n12201), .A2(n12202), .ZN(n12373) );
  OR2_X1 U12373 ( .A1(n11958), .A2(n8131), .ZN(n12202) );
  OR2_X1 U12374 ( .A1(n12374), .A2(n12375), .ZN(n12201) );
  AND2_X1 U12375 ( .A1(n12198), .A2(n12197), .ZN(n12375) );
  AND2_X1 U12376 ( .A1(n12195), .A2(n12376), .ZN(n12374) );
  OR2_X1 U12377 ( .A1(n12197), .A2(n12198), .ZN(n12376) );
  OR2_X1 U12378 ( .A1(n8126), .A2(n11958), .ZN(n12198) );
  OR2_X1 U12379 ( .A1(n12377), .A2(n12378), .ZN(n12197) );
  AND2_X1 U12380 ( .A1(n12194), .A2(n12193), .ZN(n12378) );
  AND2_X1 U12381 ( .A1(n12191), .A2(n12379), .ZN(n12377) );
  OR2_X1 U12382 ( .A1(n12193), .A2(n12194), .ZN(n12379) );
  OR2_X1 U12383 ( .A1(n8121), .A2(n11958), .ZN(n12194) );
  OR2_X1 U12384 ( .A1(n12380), .A2(n12381), .ZN(n12193) );
  AND2_X1 U12385 ( .A1(n12190), .A2(n12189), .ZN(n12381) );
  AND2_X1 U12386 ( .A1(n12187), .A2(n12382), .ZN(n12380) );
  OR2_X1 U12387 ( .A1(n12189), .A2(n12190), .ZN(n12382) );
  OR2_X1 U12388 ( .A1(n8116), .A2(n11958), .ZN(n12190) );
  OR2_X1 U12389 ( .A1(n12383), .A2(n12384), .ZN(n12189) );
  AND2_X1 U12390 ( .A1(n12186), .A2(n12185), .ZN(n12384) );
  AND2_X1 U12391 ( .A1(n12184), .A2(n12385), .ZN(n12383) );
  OR2_X1 U12392 ( .A1(n12185), .A2(n12186), .ZN(n12385) );
  OR2_X1 U12393 ( .A1(n8111), .A2(n11958), .ZN(n12186) );
  OR2_X1 U12394 ( .A1(n12386), .A2(n12387), .ZN(n12185) );
  AND2_X1 U12395 ( .A1(n12179), .A2(n12182), .ZN(n12387) );
  AND2_X1 U12396 ( .A1(n12181), .A2(n12388), .ZN(n12386) );
  OR2_X1 U12397 ( .A1(n12182), .A2(n12179), .ZN(n12388) );
  OR2_X1 U12398 ( .A1(n8102), .A2(n11958), .ZN(n12179) );
  OR3_X1 U12399 ( .A1(n8349), .A2(n11958), .A3(n12176), .ZN(n12182) );
  INV_X1 U12400 ( .A(n12389), .ZN(n12181) );
  OR2_X1 U12401 ( .A1(n12390), .A2(n12391), .ZN(n12389) );
  AND2_X1 U12402 ( .A1(b_9_), .A2(n12392), .ZN(n12391) );
  OR2_X1 U12403 ( .A1(n12393), .A2(n7318), .ZN(n12392) );
  AND2_X1 U12404 ( .A1(a_31_), .A2(n12176), .ZN(n12393) );
  AND2_X1 U12405 ( .A1(b_10_), .A2(n12394), .ZN(n12390) );
  OR2_X1 U12406 ( .A1(n12395), .A2(n7314), .ZN(n12394) );
  AND2_X1 U12407 ( .A1(a_30_), .A2(n12396), .ZN(n12395) );
  XNOR2_X1 U12408 ( .A(n12397), .B(n12398), .ZN(n12184) );
  XNOR2_X1 U12409 ( .A(n12399), .B(n12400), .ZN(n12398) );
  XOR2_X1 U12410 ( .A(n12401), .B(n12402), .Z(n12187) );
  XOR2_X1 U12411 ( .A(n12403), .B(n12404), .Z(n12402) );
  XOR2_X1 U12412 ( .A(n12405), .B(n12406), .Z(n12191) );
  XOR2_X1 U12413 ( .A(n12407), .B(n12408), .Z(n12406) );
  XOR2_X1 U12414 ( .A(n12409), .B(n12410), .Z(n12195) );
  XOR2_X1 U12415 ( .A(n12411), .B(n12412), .Z(n12410) );
  XOR2_X1 U12416 ( .A(n12413), .B(n12414), .Z(n12199) );
  XOR2_X1 U12417 ( .A(n12415), .B(n12416), .Z(n12414) );
  XOR2_X1 U12418 ( .A(n12417), .B(n12418), .Z(n12203) );
  XOR2_X1 U12419 ( .A(n12419), .B(n12420), .Z(n12418) );
  XOR2_X1 U12420 ( .A(n12421), .B(n12422), .Z(n12207) );
  XOR2_X1 U12421 ( .A(n12423), .B(n12424), .Z(n12422) );
  XOR2_X1 U12422 ( .A(n12425), .B(n12426), .Z(n12211) );
  XOR2_X1 U12423 ( .A(n12427), .B(n12428), .Z(n12426) );
  XOR2_X1 U12424 ( .A(n12429), .B(n12430), .Z(n12215) );
  XOR2_X1 U12425 ( .A(n12431), .B(n12432), .Z(n12430) );
  XOR2_X1 U12426 ( .A(n12433), .B(n12434), .Z(n12219) );
  XOR2_X1 U12427 ( .A(n12435), .B(n12436), .Z(n12434) );
  XOR2_X1 U12428 ( .A(n12437), .B(n12438), .Z(n12223) );
  XOR2_X1 U12429 ( .A(n12439), .B(n12440), .Z(n12438) );
  XOR2_X1 U12430 ( .A(n12441), .B(n12442), .Z(n12227) );
  XOR2_X1 U12431 ( .A(n12443), .B(n12444), .Z(n12442) );
  XOR2_X1 U12432 ( .A(n12445), .B(n12446), .Z(n12231) );
  XOR2_X1 U12433 ( .A(n12447), .B(n12448), .Z(n12446) );
  XOR2_X1 U12434 ( .A(n12449), .B(n12450), .Z(n12235) );
  XOR2_X1 U12435 ( .A(n12451), .B(n12452), .Z(n12450) );
  XOR2_X1 U12436 ( .A(n12453), .B(n12454), .Z(n12239) );
  XOR2_X1 U12437 ( .A(n12455), .B(n12456), .Z(n12454) );
  XOR2_X1 U12438 ( .A(n12457), .B(n12458), .Z(n12243) );
  XOR2_X1 U12439 ( .A(n12459), .B(n12460), .Z(n12458) );
  XOR2_X1 U12440 ( .A(n12461), .B(n12462), .Z(n12247) );
  XOR2_X1 U12441 ( .A(n12463), .B(n12464), .Z(n12462) );
  XOR2_X1 U12442 ( .A(n12465), .B(n12466), .Z(n12252) );
  XOR2_X1 U12443 ( .A(n12467), .B(n12468), .Z(n12466) );
  XOR2_X1 U12444 ( .A(n12469), .B(n12470), .Z(n12255) );
  XOR2_X1 U12445 ( .A(n12471), .B(n12472), .Z(n12470) );
  XNOR2_X1 U12446 ( .A(n12473), .B(n12474), .ZN(n12259) );
  XNOR2_X1 U12447 ( .A(n12475), .B(n12476), .ZN(n12473) );
  XOR2_X1 U12448 ( .A(n12477), .B(n12478), .Z(n12263) );
  XOR2_X1 U12449 ( .A(n12479), .B(n12480), .Z(n12478) );
  XOR2_X1 U12450 ( .A(n12481), .B(n12482), .Z(n12267) );
  XOR2_X1 U12451 ( .A(n12483), .B(n12484), .Z(n12482) );
  XOR2_X1 U12452 ( .A(n12485), .B(n12486), .Z(n12271) );
  XOR2_X1 U12453 ( .A(n12487), .B(n12488), .Z(n12486) );
  XOR2_X1 U12454 ( .A(n12489), .B(n12490), .Z(n12275) );
  XOR2_X1 U12455 ( .A(n12491), .B(n12492), .Z(n12490) );
  XOR2_X1 U12456 ( .A(n12493), .B(n12494), .Z(n12279) );
  XOR2_X1 U12457 ( .A(n12495), .B(n12496), .Z(n12494) );
  XOR2_X1 U12458 ( .A(n12497), .B(n12498), .Z(n12283) );
  XOR2_X1 U12459 ( .A(n12499), .B(n12500), .Z(n12498) );
  XOR2_X1 U12460 ( .A(n12501), .B(n12502), .Z(n12287) );
  XOR2_X1 U12461 ( .A(n12503), .B(n12504), .Z(n12502) );
  XOR2_X1 U12462 ( .A(n12505), .B(n12506), .Z(n12291) );
  XOR2_X1 U12463 ( .A(n12507), .B(n12508), .Z(n12506) );
  XOR2_X1 U12464 ( .A(n12509), .B(n12510), .Z(n12295) );
  XOR2_X1 U12465 ( .A(n12511), .B(n12512), .Z(n12510) );
  XNOR2_X1 U12466 ( .A(n12513), .B(n12514), .ZN(n7588) );
  XOR2_X1 U12467 ( .A(n12515), .B(n12516), .Z(n12514) );
  XNOR2_X1 U12468 ( .A(n7295), .B(n7799), .ZN(n7586) );
  OR2_X1 U12469 ( .A1(n12517), .A2(n12518), .ZN(n7799) );
  AND2_X1 U12470 ( .A1(n12516), .A2(n12515), .ZN(n12518) );
  AND2_X1 U12471 ( .A1(n12513), .A2(n12519), .ZN(n12517) );
  OR2_X1 U12472 ( .A1(n12515), .A2(n12516), .ZN(n12519) );
  OR2_X1 U12473 ( .A1(n12176), .A2(n7621), .ZN(n12516) );
  OR2_X1 U12474 ( .A1(n12520), .A2(n12521), .ZN(n12515) );
  AND2_X1 U12475 ( .A1(n12512), .A2(n12511), .ZN(n12521) );
  AND2_X1 U12476 ( .A1(n12509), .A2(n12522), .ZN(n12520) );
  OR2_X1 U12477 ( .A1(n12511), .A2(n12512), .ZN(n12522) );
  OR2_X1 U12478 ( .A1(n12176), .A2(n7656), .ZN(n12512) );
  OR2_X1 U12479 ( .A1(n12523), .A2(n12524), .ZN(n12511) );
  AND2_X1 U12480 ( .A1(n12508), .A2(n12507), .ZN(n12524) );
  AND2_X1 U12481 ( .A1(n12505), .A2(n12525), .ZN(n12523) );
  OR2_X1 U12482 ( .A1(n12507), .A2(n12508), .ZN(n12525) );
  OR2_X1 U12483 ( .A1(n12176), .A2(n7689), .ZN(n12508) );
  OR2_X1 U12484 ( .A1(n12526), .A2(n12527), .ZN(n12507) );
  AND2_X1 U12485 ( .A1(n12504), .A2(n12503), .ZN(n12527) );
  AND2_X1 U12486 ( .A1(n12501), .A2(n12528), .ZN(n12526) );
  OR2_X1 U12487 ( .A1(n12503), .A2(n12504), .ZN(n12528) );
  OR2_X1 U12488 ( .A1(n12176), .A2(n7777), .ZN(n12504) );
  OR2_X1 U12489 ( .A1(n12529), .A2(n12530), .ZN(n12503) );
  AND2_X1 U12490 ( .A1(n12500), .A2(n12499), .ZN(n12530) );
  AND2_X1 U12491 ( .A1(n12497), .A2(n12531), .ZN(n12529) );
  OR2_X1 U12492 ( .A1(n12499), .A2(n12500), .ZN(n12531) );
  OR2_X1 U12493 ( .A1(n12176), .A2(n7785), .ZN(n12500) );
  OR2_X1 U12494 ( .A1(n12532), .A2(n12533), .ZN(n12499) );
  AND2_X1 U12495 ( .A1(n12496), .A2(n12495), .ZN(n12533) );
  AND2_X1 U12496 ( .A1(n12493), .A2(n12534), .ZN(n12532) );
  OR2_X1 U12497 ( .A1(n12495), .A2(n12496), .ZN(n12534) );
  OR2_X1 U12498 ( .A1(n12176), .A2(n8226), .ZN(n12496) );
  OR2_X1 U12499 ( .A1(n12535), .A2(n12536), .ZN(n12495) );
  AND2_X1 U12500 ( .A1(n12492), .A2(n12491), .ZN(n12536) );
  AND2_X1 U12501 ( .A1(n12489), .A2(n12537), .ZN(n12535) );
  OR2_X1 U12502 ( .A1(n12491), .A2(n12492), .ZN(n12537) );
  OR2_X1 U12503 ( .A1(n12176), .A2(n8221), .ZN(n12492) );
  OR2_X1 U12504 ( .A1(n12538), .A2(n12539), .ZN(n12491) );
  AND2_X1 U12505 ( .A1(n12488), .A2(n12487), .ZN(n12539) );
  AND2_X1 U12506 ( .A1(n12485), .A2(n12540), .ZN(n12538) );
  OR2_X1 U12507 ( .A1(n12487), .A2(n12488), .ZN(n12540) );
  OR2_X1 U12508 ( .A1(n12176), .A2(n8216), .ZN(n12488) );
  OR2_X1 U12509 ( .A1(n12541), .A2(n12542), .ZN(n12487) );
  AND2_X1 U12510 ( .A1(n12484), .A2(n12483), .ZN(n12542) );
  AND2_X1 U12511 ( .A1(n12481), .A2(n12543), .ZN(n12541) );
  OR2_X1 U12512 ( .A1(n12483), .A2(n12484), .ZN(n12543) );
  OR2_X1 U12513 ( .A1(n12176), .A2(n8211), .ZN(n12484) );
  OR2_X1 U12514 ( .A1(n12544), .A2(n12545), .ZN(n12483) );
  AND2_X1 U12515 ( .A1(n12480), .A2(n12479), .ZN(n12545) );
  AND2_X1 U12516 ( .A1(n12477), .A2(n12546), .ZN(n12544) );
  OR2_X1 U12517 ( .A1(n12479), .A2(n12480), .ZN(n12546) );
  OR2_X1 U12518 ( .A1(n12176), .A2(n8206), .ZN(n12480) );
  OR2_X1 U12519 ( .A1(n12547), .A2(n12548), .ZN(n12479) );
  AND2_X1 U12520 ( .A1(n12474), .A2(n12476), .ZN(n12548) );
  AND2_X1 U12521 ( .A1(n12549), .A2(n12475), .ZN(n12547) );
  OR2_X1 U12522 ( .A1(n12474), .A2(n12476), .ZN(n12549) );
  OR2_X1 U12523 ( .A1(n12550), .A2(n12551), .ZN(n12476) );
  AND2_X1 U12524 ( .A1(n12472), .A2(n12471), .ZN(n12551) );
  AND2_X1 U12525 ( .A1(n12469), .A2(n12552), .ZN(n12550) );
  OR2_X1 U12526 ( .A1(n12471), .A2(n12472), .ZN(n12552) );
  OR2_X1 U12527 ( .A1(n12176), .A2(n8196), .ZN(n12472) );
  OR2_X1 U12528 ( .A1(n12553), .A2(n12554), .ZN(n12471) );
  AND2_X1 U12529 ( .A1(n12468), .A2(n12467), .ZN(n12554) );
  AND2_X1 U12530 ( .A1(n12465), .A2(n12555), .ZN(n12553) );
  OR2_X1 U12531 ( .A1(n12467), .A2(n12468), .ZN(n12555) );
  OR2_X1 U12532 ( .A1(n12176), .A2(n8191), .ZN(n12468) );
  OR2_X1 U12533 ( .A1(n12556), .A2(n12557), .ZN(n12467) );
  AND2_X1 U12534 ( .A1(n12464), .A2(n12463), .ZN(n12557) );
  AND2_X1 U12535 ( .A1(n12461), .A2(n12558), .ZN(n12556) );
  OR2_X1 U12536 ( .A1(n12463), .A2(n12464), .ZN(n12558) );
  OR2_X1 U12537 ( .A1(n12176), .A2(n8186), .ZN(n12464) );
  OR2_X1 U12538 ( .A1(n12559), .A2(n12560), .ZN(n12463) );
  AND2_X1 U12539 ( .A1(n12460), .A2(n12459), .ZN(n12560) );
  AND2_X1 U12540 ( .A1(n12457), .A2(n12561), .ZN(n12559) );
  OR2_X1 U12541 ( .A1(n12459), .A2(n12460), .ZN(n12561) );
  OR2_X1 U12542 ( .A1(n12176), .A2(n8181), .ZN(n12460) );
  OR2_X1 U12543 ( .A1(n12562), .A2(n12563), .ZN(n12459) );
  AND2_X1 U12544 ( .A1(n12456), .A2(n12455), .ZN(n12563) );
  AND2_X1 U12545 ( .A1(n12453), .A2(n12564), .ZN(n12562) );
  OR2_X1 U12546 ( .A1(n12455), .A2(n12456), .ZN(n12564) );
  OR2_X1 U12547 ( .A1(n12176), .A2(n8176), .ZN(n12456) );
  OR2_X1 U12548 ( .A1(n12565), .A2(n12566), .ZN(n12455) );
  AND2_X1 U12549 ( .A1(n12452), .A2(n12451), .ZN(n12566) );
  AND2_X1 U12550 ( .A1(n12449), .A2(n12567), .ZN(n12565) );
  OR2_X1 U12551 ( .A1(n12451), .A2(n12452), .ZN(n12567) );
  OR2_X1 U12552 ( .A1(n12176), .A2(n8171), .ZN(n12452) );
  OR2_X1 U12553 ( .A1(n12568), .A2(n12569), .ZN(n12451) );
  AND2_X1 U12554 ( .A1(n12448), .A2(n12447), .ZN(n12569) );
  AND2_X1 U12555 ( .A1(n12445), .A2(n12570), .ZN(n12568) );
  OR2_X1 U12556 ( .A1(n12447), .A2(n12448), .ZN(n12570) );
  OR2_X1 U12557 ( .A1(n8166), .A2(n12176), .ZN(n12448) );
  OR2_X1 U12558 ( .A1(n12571), .A2(n12572), .ZN(n12447) );
  AND2_X1 U12559 ( .A1(n12444), .A2(n12443), .ZN(n12572) );
  AND2_X1 U12560 ( .A1(n12441), .A2(n12573), .ZN(n12571) );
  OR2_X1 U12561 ( .A1(n12443), .A2(n12444), .ZN(n12573) );
  OR2_X1 U12562 ( .A1(n12176), .A2(n8161), .ZN(n12444) );
  OR2_X1 U12563 ( .A1(n12574), .A2(n12575), .ZN(n12443) );
  AND2_X1 U12564 ( .A1(n12437), .A2(n12440), .ZN(n12575) );
  AND2_X1 U12565 ( .A1(n12576), .A2(n12439), .ZN(n12574) );
  OR2_X1 U12566 ( .A1(n12577), .A2(n12578), .ZN(n12439) );
  AND2_X1 U12567 ( .A1(n12436), .A2(n12435), .ZN(n12578) );
  AND2_X1 U12568 ( .A1(n12433), .A2(n12579), .ZN(n12577) );
  OR2_X1 U12569 ( .A1(n12435), .A2(n12436), .ZN(n12579) );
  OR2_X1 U12570 ( .A1(n12176), .A2(n8151), .ZN(n12436) );
  OR2_X1 U12571 ( .A1(n12580), .A2(n12581), .ZN(n12435) );
  AND2_X1 U12572 ( .A1(n12429), .A2(n12432), .ZN(n12581) );
  AND2_X1 U12573 ( .A1(n12582), .A2(n12431), .ZN(n12580) );
  OR2_X1 U12574 ( .A1(n12583), .A2(n12584), .ZN(n12431) );
  AND2_X1 U12575 ( .A1(n12425), .A2(n12428), .ZN(n12584) );
  AND2_X1 U12576 ( .A1(n12585), .A2(n12427), .ZN(n12583) );
  OR2_X1 U12577 ( .A1(n12586), .A2(n12587), .ZN(n12427) );
  AND2_X1 U12578 ( .A1(n12421), .A2(n12424), .ZN(n12587) );
  AND2_X1 U12579 ( .A1(n12588), .A2(n12423), .ZN(n12586) );
  OR2_X1 U12580 ( .A1(n12589), .A2(n12590), .ZN(n12423) );
  AND2_X1 U12581 ( .A1(n12417), .A2(n12420), .ZN(n12590) );
  AND2_X1 U12582 ( .A1(n12591), .A2(n12419), .ZN(n12589) );
  OR2_X1 U12583 ( .A1(n12592), .A2(n12593), .ZN(n12419) );
  AND2_X1 U12584 ( .A1(n12413), .A2(n12416), .ZN(n12593) );
  AND2_X1 U12585 ( .A1(n12594), .A2(n12415), .ZN(n12592) );
  OR2_X1 U12586 ( .A1(n12595), .A2(n12596), .ZN(n12415) );
  AND2_X1 U12587 ( .A1(n12409), .A2(n12412), .ZN(n12596) );
  AND2_X1 U12588 ( .A1(n12597), .A2(n12411), .ZN(n12595) );
  OR2_X1 U12589 ( .A1(n12598), .A2(n12599), .ZN(n12411) );
  AND2_X1 U12590 ( .A1(n12405), .A2(n12408), .ZN(n12599) );
  AND2_X1 U12591 ( .A1(n12600), .A2(n12407), .ZN(n12598) );
  OR2_X1 U12592 ( .A1(n12601), .A2(n12602), .ZN(n12407) );
  AND2_X1 U12593 ( .A1(n12401), .A2(n12404), .ZN(n12602) );
  AND2_X1 U12594 ( .A1(n12603), .A2(n12403), .ZN(n12601) );
  OR2_X1 U12595 ( .A1(n12604), .A2(n12605), .ZN(n12403) );
  AND2_X1 U12596 ( .A1(n12397), .A2(n12400), .ZN(n12605) );
  AND2_X1 U12597 ( .A1(n12399), .A2(n12606), .ZN(n12604) );
  OR2_X1 U12598 ( .A1(n12400), .A2(n12397), .ZN(n12606) );
  OR2_X1 U12599 ( .A1(n8102), .A2(n12176), .ZN(n12397) );
  OR3_X1 U12600 ( .A1(n8349), .A2(n12176), .A3(n12396), .ZN(n12400) );
  INV_X1 U12601 ( .A(n12607), .ZN(n12399) );
  OR2_X1 U12602 ( .A1(n12608), .A2(n12609), .ZN(n12607) );
  AND2_X1 U12603 ( .A1(b_9_), .A2(n12610), .ZN(n12609) );
  OR2_X1 U12604 ( .A1(n12611), .A2(n7314), .ZN(n12610) );
  AND2_X1 U12605 ( .A1(a_30_), .A2(n12612), .ZN(n12611) );
  AND2_X1 U12606 ( .A1(b_8_), .A2(n12613), .ZN(n12608) );
  OR2_X1 U12607 ( .A1(n12614), .A2(n7318), .ZN(n12613) );
  AND2_X1 U12608 ( .A1(a_31_), .A2(n12396), .ZN(n12614) );
  OR2_X1 U12609 ( .A1(n12404), .A2(n12401), .ZN(n12603) );
  XNOR2_X1 U12610 ( .A(n12615), .B(n12616), .ZN(n12401) );
  XNOR2_X1 U12611 ( .A(n12617), .B(n12618), .ZN(n12616) );
  OR2_X1 U12612 ( .A1(n8111), .A2(n12176), .ZN(n12404) );
  OR2_X1 U12613 ( .A1(n12408), .A2(n12405), .ZN(n12600) );
  XOR2_X1 U12614 ( .A(n12619), .B(n12620), .Z(n12405) );
  XOR2_X1 U12615 ( .A(n12621), .B(n12622), .Z(n12620) );
  OR2_X1 U12616 ( .A1(n8116), .A2(n12176), .ZN(n12408) );
  OR2_X1 U12617 ( .A1(n12412), .A2(n12409), .ZN(n12597) );
  XOR2_X1 U12618 ( .A(n12623), .B(n12624), .Z(n12409) );
  XOR2_X1 U12619 ( .A(n12625), .B(n12626), .Z(n12624) );
  OR2_X1 U12620 ( .A1(n8121), .A2(n12176), .ZN(n12412) );
  OR2_X1 U12621 ( .A1(n12416), .A2(n12413), .ZN(n12594) );
  XOR2_X1 U12622 ( .A(n12627), .B(n12628), .Z(n12413) );
  XOR2_X1 U12623 ( .A(n12629), .B(n12630), .Z(n12628) );
  OR2_X1 U12624 ( .A1(n8126), .A2(n12176), .ZN(n12416) );
  OR2_X1 U12625 ( .A1(n12420), .A2(n12417), .ZN(n12591) );
  XOR2_X1 U12626 ( .A(n12631), .B(n12632), .Z(n12417) );
  XOR2_X1 U12627 ( .A(n12633), .B(n12634), .Z(n12632) );
  OR2_X1 U12628 ( .A1(n8131), .A2(n12176), .ZN(n12420) );
  OR2_X1 U12629 ( .A1(n12424), .A2(n12421), .ZN(n12588) );
  XOR2_X1 U12630 ( .A(n12635), .B(n12636), .Z(n12421) );
  XOR2_X1 U12631 ( .A(n12637), .B(n12638), .Z(n12636) );
  OR2_X1 U12632 ( .A1(n12176), .A2(n8136), .ZN(n12424) );
  OR2_X1 U12633 ( .A1(n12428), .A2(n12425), .ZN(n12585) );
  XOR2_X1 U12634 ( .A(n12639), .B(n12640), .Z(n12425) );
  XOR2_X1 U12635 ( .A(n12641), .B(n12642), .Z(n12640) );
  OR2_X1 U12636 ( .A1(n12176), .A2(n8141), .ZN(n12428) );
  OR2_X1 U12637 ( .A1(n12432), .A2(n12429), .ZN(n12582) );
  XOR2_X1 U12638 ( .A(n12643), .B(n12644), .Z(n12429) );
  XOR2_X1 U12639 ( .A(n12645), .B(n12646), .Z(n12644) );
  OR2_X1 U12640 ( .A1(n12176), .A2(n8146), .ZN(n12432) );
  XOR2_X1 U12641 ( .A(n12647), .B(n12648), .Z(n12433) );
  XOR2_X1 U12642 ( .A(n12649), .B(n12650), .Z(n12648) );
  OR2_X1 U12643 ( .A1(n12440), .A2(n12437), .ZN(n12576) );
  XOR2_X1 U12644 ( .A(n12651), .B(n12652), .Z(n12437) );
  XOR2_X1 U12645 ( .A(n12653), .B(n12654), .Z(n12652) );
  OR2_X1 U12646 ( .A1(n12176), .A2(n8156), .ZN(n12440) );
  XOR2_X1 U12647 ( .A(n12655), .B(n12656), .Z(n12441) );
  XOR2_X1 U12648 ( .A(n12657), .B(n12658), .Z(n12656) );
  XOR2_X1 U12649 ( .A(n12659), .B(n12660), .Z(n12445) );
  XOR2_X1 U12650 ( .A(n12661), .B(n12662), .Z(n12660) );
  XOR2_X1 U12651 ( .A(n12663), .B(n12664), .Z(n12449) );
  XOR2_X1 U12652 ( .A(n12665), .B(n12666), .Z(n12664) );
  XOR2_X1 U12653 ( .A(n12667), .B(n12668), .Z(n12453) );
  XOR2_X1 U12654 ( .A(n12669), .B(n12670), .Z(n12668) );
  XOR2_X1 U12655 ( .A(n12671), .B(n12672), .Z(n12457) );
  XOR2_X1 U12656 ( .A(n12673), .B(n12674), .Z(n12672) );
  XOR2_X1 U12657 ( .A(n12675), .B(n12676), .Z(n12461) );
  XOR2_X1 U12658 ( .A(n12677), .B(n12678), .Z(n12676) );
  XOR2_X1 U12659 ( .A(n12679), .B(n12680), .Z(n12465) );
  XOR2_X1 U12660 ( .A(n12681), .B(n12682), .Z(n12680) );
  XOR2_X1 U12661 ( .A(n12683), .B(n12684), .Z(n12469) );
  XOR2_X1 U12662 ( .A(n12685), .B(n12686), .Z(n12684) );
  XOR2_X1 U12663 ( .A(n12687), .B(n12688), .Z(n12474) );
  XOR2_X1 U12664 ( .A(n12689), .B(n12690), .Z(n12688) );
  XOR2_X1 U12665 ( .A(n12691), .B(n12692), .Z(n12477) );
  XOR2_X1 U12666 ( .A(n12693), .B(n12694), .Z(n12692) );
  XNOR2_X1 U12667 ( .A(n12695), .B(n12696), .ZN(n12481) );
  XNOR2_X1 U12668 ( .A(n12697), .B(n12698), .ZN(n12695) );
  XOR2_X1 U12669 ( .A(n12699), .B(n12700), .Z(n12485) );
  XOR2_X1 U12670 ( .A(n12701), .B(n12702), .Z(n12700) );
  XOR2_X1 U12671 ( .A(n12703), .B(n12704), .Z(n12489) );
  XOR2_X1 U12672 ( .A(n12705), .B(n12706), .Z(n12704) );
  XOR2_X1 U12673 ( .A(n12707), .B(n12708), .Z(n12493) );
  XOR2_X1 U12674 ( .A(n12709), .B(n12710), .Z(n12708) );
  XOR2_X1 U12675 ( .A(n12711), .B(n12712), .Z(n12497) );
  XOR2_X1 U12676 ( .A(n12713), .B(n12714), .Z(n12712) );
  XOR2_X1 U12677 ( .A(n12715), .B(n12716), .Z(n12501) );
  XOR2_X1 U12678 ( .A(n12717), .B(n12718), .Z(n12716) );
  XOR2_X1 U12679 ( .A(n12719), .B(n12720), .Z(n12505) );
  XOR2_X1 U12680 ( .A(n12721), .B(n12722), .Z(n12720) );
  XOR2_X1 U12681 ( .A(n12723), .B(n12724), .Z(n12509) );
  XOR2_X1 U12682 ( .A(n12725), .B(n12726), .Z(n12724) );
  XOR2_X1 U12683 ( .A(n12727), .B(n12728), .Z(n12513) );
  XOR2_X1 U12684 ( .A(n12729), .B(n12730), .Z(n12728) );
  XNOR2_X1 U12685 ( .A(n12731), .B(n12732), .ZN(n7295) );
  XOR2_X1 U12686 ( .A(n12733), .B(n12734), .Z(n12732) );
  INV_X1 U12687 ( .A(n12735), .ZN(n7292) );
  OR2_X1 U12688 ( .A1(n12736), .A2(n7797), .ZN(n12735) );
  INV_X1 U12689 ( .A(n12737), .ZN(n7797) );
  OR2_X1 U12690 ( .A1(n12738), .A2(n12739), .ZN(n12737) );
  AND2_X1 U12691 ( .A1(n12738), .A2(n12739), .ZN(n12736) );
  OR2_X1 U12692 ( .A1(n12740), .A2(n12741), .ZN(n12739) );
  AND2_X1 U12693 ( .A1(n12734), .A2(n12733), .ZN(n12741) );
  AND2_X1 U12694 ( .A1(n12731), .A2(n12742), .ZN(n12740) );
  OR2_X1 U12695 ( .A1(n12733), .A2(n12734), .ZN(n12742) );
  OR2_X1 U12696 ( .A1(n12396), .A2(n7621), .ZN(n12734) );
  OR2_X1 U12697 ( .A1(n12743), .A2(n12744), .ZN(n12733) );
  AND2_X1 U12698 ( .A1(n12730), .A2(n12729), .ZN(n12744) );
  AND2_X1 U12699 ( .A1(n12727), .A2(n12745), .ZN(n12743) );
  OR2_X1 U12700 ( .A1(n12729), .A2(n12730), .ZN(n12745) );
  OR2_X1 U12701 ( .A1(n12396), .A2(n7656), .ZN(n12730) );
  OR2_X1 U12702 ( .A1(n12746), .A2(n12747), .ZN(n12729) );
  AND2_X1 U12703 ( .A1(n12726), .A2(n12725), .ZN(n12747) );
  AND2_X1 U12704 ( .A1(n12723), .A2(n12748), .ZN(n12746) );
  OR2_X1 U12705 ( .A1(n12725), .A2(n12726), .ZN(n12748) );
  OR2_X1 U12706 ( .A1(n12396), .A2(n7689), .ZN(n12726) );
  OR2_X1 U12707 ( .A1(n12749), .A2(n12750), .ZN(n12725) );
  AND2_X1 U12708 ( .A1(n12722), .A2(n12721), .ZN(n12750) );
  AND2_X1 U12709 ( .A1(n12719), .A2(n12751), .ZN(n12749) );
  OR2_X1 U12710 ( .A1(n12721), .A2(n12722), .ZN(n12751) );
  OR2_X1 U12711 ( .A1(n12396), .A2(n7777), .ZN(n12722) );
  OR2_X1 U12712 ( .A1(n12752), .A2(n12753), .ZN(n12721) );
  AND2_X1 U12713 ( .A1(n12718), .A2(n12717), .ZN(n12753) );
  AND2_X1 U12714 ( .A1(n12715), .A2(n12754), .ZN(n12752) );
  OR2_X1 U12715 ( .A1(n12717), .A2(n12718), .ZN(n12754) );
  OR2_X1 U12716 ( .A1(n12396), .A2(n7785), .ZN(n12718) );
  OR2_X1 U12717 ( .A1(n12755), .A2(n12756), .ZN(n12717) );
  AND2_X1 U12718 ( .A1(n12714), .A2(n12713), .ZN(n12756) );
  AND2_X1 U12719 ( .A1(n12711), .A2(n12757), .ZN(n12755) );
  OR2_X1 U12720 ( .A1(n12713), .A2(n12714), .ZN(n12757) );
  OR2_X1 U12721 ( .A1(n12396), .A2(n8226), .ZN(n12714) );
  OR2_X1 U12722 ( .A1(n12758), .A2(n12759), .ZN(n12713) );
  AND2_X1 U12723 ( .A1(n12710), .A2(n12709), .ZN(n12759) );
  AND2_X1 U12724 ( .A1(n12707), .A2(n12760), .ZN(n12758) );
  OR2_X1 U12725 ( .A1(n12709), .A2(n12710), .ZN(n12760) );
  OR2_X1 U12726 ( .A1(n12396), .A2(n8221), .ZN(n12710) );
  OR2_X1 U12727 ( .A1(n12761), .A2(n12762), .ZN(n12709) );
  AND2_X1 U12728 ( .A1(n12706), .A2(n12705), .ZN(n12762) );
  AND2_X1 U12729 ( .A1(n12703), .A2(n12763), .ZN(n12761) );
  OR2_X1 U12730 ( .A1(n12705), .A2(n12706), .ZN(n12763) );
  OR2_X1 U12731 ( .A1(n12396), .A2(n8216), .ZN(n12706) );
  OR2_X1 U12732 ( .A1(n12764), .A2(n12765), .ZN(n12705) );
  AND2_X1 U12733 ( .A1(n12702), .A2(n12701), .ZN(n12765) );
  AND2_X1 U12734 ( .A1(n12699), .A2(n12766), .ZN(n12764) );
  OR2_X1 U12735 ( .A1(n12701), .A2(n12702), .ZN(n12766) );
  OR2_X1 U12736 ( .A1(n12396), .A2(n8211), .ZN(n12702) );
  OR2_X1 U12737 ( .A1(n12767), .A2(n12768), .ZN(n12701) );
  AND2_X1 U12738 ( .A1(n12696), .A2(n12698), .ZN(n12768) );
  AND2_X1 U12739 ( .A1(n12769), .A2(n12697), .ZN(n12767) );
  OR2_X1 U12740 ( .A1(n12696), .A2(n12698), .ZN(n12769) );
  OR2_X1 U12741 ( .A1(n12770), .A2(n12771), .ZN(n12698) );
  AND2_X1 U12742 ( .A1(n12694), .A2(n12693), .ZN(n12771) );
  AND2_X1 U12743 ( .A1(n12691), .A2(n12772), .ZN(n12770) );
  OR2_X1 U12744 ( .A1(n12693), .A2(n12694), .ZN(n12772) );
  OR2_X1 U12745 ( .A1(n12396), .A2(n8201), .ZN(n12694) );
  OR2_X1 U12746 ( .A1(n12773), .A2(n12774), .ZN(n12693) );
  AND2_X1 U12747 ( .A1(n12690), .A2(n12689), .ZN(n12774) );
  AND2_X1 U12748 ( .A1(n12687), .A2(n12775), .ZN(n12773) );
  OR2_X1 U12749 ( .A1(n12689), .A2(n12690), .ZN(n12775) );
  OR2_X1 U12750 ( .A1(n12396), .A2(n8196), .ZN(n12690) );
  OR2_X1 U12751 ( .A1(n12776), .A2(n12777), .ZN(n12689) );
  AND2_X1 U12752 ( .A1(n12686), .A2(n12685), .ZN(n12777) );
  AND2_X1 U12753 ( .A1(n12683), .A2(n12778), .ZN(n12776) );
  OR2_X1 U12754 ( .A1(n12685), .A2(n12686), .ZN(n12778) );
  OR2_X1 U12755 ( .A1(n12396), .A2(n8191), .ZN(n12686) );
  OR2_X1 U12756 ( .A1(n12779), .A2(n12780), .ZN(n12685) );
  AND2_X1 U12757 ( .A1(n12682), .A2(n12681), .ZN(n12780) );
  AND2_X1 U12758 ( .A1(n12679), .A2(n12781), .ZN(n12779) );
  OR2_X1 U12759 ( .A1(n12681), .A2(n12682), .ZN(n12781) );
  OR2_X1 U12760 ( .A1(n12396), .A2(n8186), .ZN(n12682) );
  OR2_X1 U12761 ( .A1(n12782), .A2(n12783), .ZN(n12681) );
  AND2_X1 U12762 ( .A1(n12678), .A2(n12677), .ZN(n12783) );
  AND2_X1 U12763 ( .A1(n12675), .A2(n12784), .ZN(n12782) );
  OR2_X1 U12764 ( .A1(n12677), .A2(n12678), .ZN(n12784) );
  OR2_X1 U12765 ( .A1(n12396), .A2(n8181), .ZN(n12678) );
  OR2_X1 U12766 ( .A1(n12785), .A2(n12786), .ZN(n12677) );
  AND2_X1 U12767 ( .A1(n12674), .A2(n12673), .ZN(n12786) );
  AND2_X1 U12768 ( .A1(n12671), .A2(n12787), .ZN(n12785) );
  OR2_X1 U12769 ( .A1(n12673), .A2(n12674), .ZN(n12787) );
  OR2_X1 U12770 ( .A1(n12396), .A2(n8176), .ZN(n12674) );
  OR2_X1 U12771 ( .A1(n12788), .A2(n12789), .ZN(n12673) );
  AND2_X1 U12772 ( .A1(n12670), .A2(n12669), .ZN(n12789) );
  AND2_X1 U12773 ( .A1(n12667), .A2(n12790), .ZN(n12788) );
  OR2_X1 U12774 ( .A1(n12669), .A2(n12670), .ZN(n12790) );
  OR2_X1 U12775 ( .A1(n12396), .A2(n8171), .ZN(n12670) );
  OR2_X1 U12776 ( .A1(n12791), .A2(n12792), .ZN(n12669) );
  AND2_X1 U12777 ( .A1(n12666), .A2(n12665), .ZN(n12792) );
  AND2_X1 U12778 ( .A1(n12663), .A2(n12793), .ZN(n12791) );
  OR2_X1 U12779 ( .A1(n12665), .A2(n12666), .ZN(n12793) );
  OR2_X1 U12780 ( .A1(n8166), .A2(n12396), .ZN(n12666) );
  OR2_X1 U12781 ( .A1(n12794), .A2(n12795), .ZN(n12665) );
  AND2_X1 U12782 ( .A1(n12662), .A2(n12661), .ZN(n12795) );
  AND2_X1 U12783 ( .A1(n12659), .A2(n12796), .ZN(n12794) );
  OR2_X1 U12784 ( .A1(n12661), .A2(n12662), .ZN(n12796) );
  OR2_X1 U12785 ( .A1(n12396), .A2(n8161), .ZN(n12662) );
  OR2_X1 U12786 ( .A1(n12797), .A2(n12798), .ZN(n12661) );
  AND2_X1 U12787 ( .A1(n12658), .A2(n12657), .ZN(n12798) );
  AND2_X1 U12788 ( .A1(n12655), .A2(n12799), .ZN(n12797) );
  OR2_X1 U12789 ( .A1(n12657), .A2(n12658), .ZN(n12799) );
  OR2_X1 U12790 ( .A1(n12396), .A2(n8156), .ZN(n12658) );
  OR2_X1 U12791 ( .A1(n12800), .A2(n12801), .ZN(n12657) );
  AND2_X1 U12792 ( .A1(n12651), .A2(n12654), .ZN(n12801) );
  AND2_X1 U12793 ( .A1(n12802), .A2(n12653), .ZN(n12800) );
  OR2_X1 U12794 ( .A1(n12803), .A2(n12804), .ZN(n12653) );
  AND2_X1 U12795 ( .A1(n12650), .A2(n12649), .ZN(n12804) );
  AND2_X1 U12796 ( .A1(n12647), .A2(n12805), .ZN(n12803) );
  OR2_X1 U12797 ( .A1(n12649), .A2(n12650), .ZN(n12805) );
  OR2_X1 U12798 ( .A1(n12396), .A2(n8146), .ZN(n12650) );
  OR2_X1 U12799 ( .A1(n12806), .A2(n12807), .ZN(n12649) );
  AND2_X1 U12800 ( .A1(n12643), .A2(n12646), .ZN(n12807) );
  AND2_X1 U12801 ( .A1(n12808), .A2(n12645), .ZN(n12806) );
  OR2_X1 U12802 ( .A1(n12809), .A2(n12810), .ZN(n12645) );
  AND2_X1 U12803 ( .A1(n12639), .A2(n12642), .ZN(n12810) );
  AND2_X1 U12804 ( .A1(n12811), .A2(n12641), .ZN(n12809) );
  OR2_X1 U12805 ( .A1(n12812), .A2(n12813), .ZN(n12641) );
  AND2_X1 U12806 ( .A1(n12635), .A2(n12638), .ZN(n12813) );
  AND2_X1 U12807 ( .A1(n12814), .A2(n12637), .ZN(n12812) );
  OR2_X1 U12808 ( .A1(n12815), .A2(n12816), .ZN(n12637) );
  AND2_X1 U12809 ( .A1(n12631), .A2(n12634), .ZN(n12816) );
  AND2_X1 U12810 ( .A1(n12817), .A2(n12633), .ZN(n12815) );
  OR2_X1 U12811 ( .A1(n12818), .A2(n12819), .ZN(n12633) );
  AND2_X1 U12812 ( .A1(n12627), .A2(n12630), .ZN(n12819) );
  AND2_X1 U12813 ( .A1(n12820), .A2(n12629), .ZN(n12818) );
  OR2_X1 U12814 ( .A1(n12821), .A2(n12822), .ZN(n12629) );
  AND2_X1 U12815 ( .A1(n12623), .A2(n12626), .ZN(n12822) );
  AND2_X1 U12816 ( .A1(n12823), .A2(n12625), .ZN(n12821) );
  OR2_X1 U12817 ( .A1(n12824), .A2(n12825), .ZN(n12625) );
  AND2_X1 U12818 ( .A1(n12619), .A2(n12622), .ZN(n12825) );
  AND2_X1 U12819 ( .A1(n12826), .A2(n12621), .ZN(n12824) );
  OR2_X1 U12820 ( .A1(n12827), .A2(n12828), .ZN(n12621) );
  AND2_X1 U12821 ( .A1(n12615), .A2(n12618), .ZN(n12828) );
  AND2_X1 U12822 ( .A1(n12617), .A2(n12829), .ZN(n12827) );
  OR2_X1 U12823 ( .A1(n12618), .A2(n12615), .ZN(n12829) );
  OR2_X1 U12824 ( .A1(n8102), .A2(n12396), .ZN(n12615) );
  OR3_X1 U12825 ( .A1(n8349), .A2(n12396), .A3(n12612), .ZN(n12618) );
  INV_X1 U12826 ( .A(n12830), .ZN(n12617) );
  OR2_X1 U12827 ( .A1(n12831), .A2(n12832), .ZN(n12830) );
  AND2_X1 U12828 ( .A1(b_8_), .A2(n12833), .ZN(n12832) );
  OR2_X1 U12829 ( .A1(n12834), .A2(n7314), .ZN(n12833) );
  AND2_X1 U12830 ( .A1(a_30_), .A2(n7755), .ZN(n12834) );
  AND2_X1 U12831 ( .A1(b_7_), .A2(n12835), .ZN(n12831) );
  OR2_X1 U12832 ( .A1(n12836), .A2(n7318), .ZN(n12835) );
  AND2_X1 U12833 ( .A1(a_31_), .A2(n12612), .ZN(n12836) );
  OR2_X1 U12834 ( .A1(n12622), .A2(n12619), .ZN(n12826) );
  XNOR2_X1 U12835 ( .A(n12837), .B(n12838), .ZN(n12619) );
  XNOR2_X1 U12836 ( .A(n12839), .B(n12840), .ZN(n12838) );
  OR2_X1 U12837 ( .A1(n8111), .A2(n12396), .ZN(n12622) );
  OR2_X1 U12838 ( .A1(n12626), .A2(n12623), .ZN(n12823) );
  XOR2_X1 U12839 ( .A(n12841), .B(n12842), .Z(n12623) );
  XOR2_X1 U12840 ( .A(n12843), .B(n12844), .Z(n12842) );
  OR2_X1 U12841 ( .A1(n8116), .A2(n12396), .ZN(n12626) );
  OR2_X1 U12842 ( .A1(n12630), .A2(n12627), .ZN(n12820) );
  XOR2_X1 U12843 ( .A(n12845), .B(n12846), .Z(n12627) );
  XOR2_X1 U12844 ( .A(n12847), .B(n12848), .Z(n12846) );
  OR2_X1 U12845 ( .A1(n8121), .A2(n12396), .ZN(n12630) );
  OR2_X1 U12846 ( .A1(n12634), .A2(n12631), .ZN(n12817) );
  XOR2_X1 U12847 ( .A(n12849), .B(n12850), .Z(n12631) );
  XOR2_X1 U12848 ( .A(n12851), .B(n12852), .Z(n12850) );
  OR2_X1 U12849 ( .A1(n8126), .A2(n12396), .ZN(n12634) );
  OR2_X1 U12850 ( .A1(n12638), .A2(n12635), .ZN(n12814) );
  XOR2_X1 U12851 ( .A(n12853), .B(n12854), .Z(n12635) );
  XOR2_X1 U12852 ( .A(n12855), .B(n12856), .Z(n12854) );
  OR2_X1 U12853 ( .A1(n8131), .A2(n12396), .ZN(n12638) );
  OR2_X1 U12854 ( .A1(n12642), .A2(n12639), .ZN(n12811) );
  XOR2_X1 U12855 ( .A(n12857), .B(n12858), .Z(n12639) );
  XOR2_X1 U12856 ( .A(n12859), .B(n12860), .Z(n12858) );
  OR2_X1 U12857 ( .A1(n8136), .A2(n12396), .ZN(n12642) );
  OR2_X1 U12858 ( .A1(n12646), .A2(n12643), .ZN(n12808) );
  XOR2_X1 U12859 ( .A(n12861), .B(n12862), .Z(n12643) );
  XOR2_X1 U12860 ( .A(n12863), .B(n12864), .Z(n12862) );
  OR2_X1 U12861 ( .A1(n12396), .A2(n8141), .ZN(n12646) );
  XOR2_X1 U12862 ( .A(n12865), .B(n12866), .Z(n12647) );
  XOR2_X1 U12863 ( .A(n12867), .B(n12868), .Z(n12866) );
  OR2_X1 U12864 ( .A1(n12654), .A2(n12651), .ZN(n12802) );
  XOR2_X1 U12865 ( .A(n12869), .B(n12870), .Z(n12651) );
  XOR2_X1 U12866 ( .A(n12871), .B(n12872), .Z(n12870) );
  OR2_X1 U12867 ( .A1(n12396), .A2(n8151), .ZN(n12654) );
  XOR2_X1 U12868 ( .A(n12873), .B(n12874), .Z(n12655) );
  XOR2_X1 U12869 ( .A(n12875), .B(n12876), .Z(n12874) );
  XOR2_X1 U12870 ( .A(n12877), .B(n12878), .Z(n12659) );
  XOR2_X1 U12871 ( .A(n12879), .B(n12880), .Z(n12878) );
  XOR2_X1 U12872 ( .A(n12881), .B(n12882), .Z(n12663) );
  XOR2_X1 U12873 ( .A(n12883), .B(n12884), .Z(n12882) );
  XOR2_X1 U12874 ( .A(n12885), .B(n12886), .Z(n12667) );
  XOR2_X1 U12875 ( .A(n12887), .B(n12888), .Z(n12886) );
  XOR2_X1 U12876 ( .A(n12889), .B(n12890), .Z(n12671) );
  XOR2_X1 U12877 ( .A(n12891), .B(n12892), .Z(n12890) );
  XOR2_X1 U12878 ( .A(n12893), .B(n12894), .Z(n12675) );
  XOR2_X1 U12879 ( .A(n12895), .B(n12896), .Z(n12894) );
  XOR2_X1 U12880 ( .A(n12897), .B(n12898), .Z(n12679) );
  XOR2_X1 U12881 ( .A(n12899), .B(n12900), .Z(n12898) );
  XOR2_X1 U12882 ( .A(n12901), .B(n12902), .Z(n12683) );
  XOR2_X1 U12883 ( .A(n12903), .B(n12904), .Z(n12902) );
  XOR2_X1 U12884 ( .A(n12905), .B(n12906), .Z(n12687) );
  XOR2_X1 U12885 ( .A(n12907), .B(n12908), .Z(n12906) );
  XOR2_X1 U12886 ( .A(n12909), .B(n12910), .Z(n12691) );
  XOR2_X1 U12887 ( .A(n12911), .B(n12912), .Z(n12910) );
  XOR2_X1 U12888 ( .A(n12913), .B(n12914), .Z(n12696) );
  XOR2_X1 U12889 ( .A(n12915), .B(n12916), .Z(n12914) );
  XOR2_X1 U12890 ( .A(n12917), .B(n12918), .Z(n12699) );
  XOR2_X1 U12891 ( .A(n12919), .B(n12920), .Z(n12918) );
  XNOR2_X1 U12892 ( .A(n12921), .B(n12922), .ZN(n12703) );
  XNOR2_X1 U12893 ( .A(n12923), .B(n12924), .ZN(n12921) );
  XOR2_X1 U12894 ( .A(n12925), .B(n12926), .Z(n12707) );
  XOR2_X1 U12895 ( .A(n12927), .B(n12928), .Z(n12926) );
  XOR2_X1 U12896 ( .A(n12929), .B(n12930), .Z(n12711) );
  XOR2_X1 U12897 ( .A(n12931), .B(n12932), .Z(n12930) );
  XOR2_X1 U12898 ( .A(n12933), .B(n12934), .Z(n12715) );
  XOR2_X1 U12899 ( .A(n12935), .B(n12936), .Z(n12934) );
  XOR2_X1 U12900 ( .A(n12937), .B(n12938), .Z(n12719) );
  XOR2_X1 U12901 ( .A(n12939), .B(n12940), .Z(n12938) );
  XOR2_X1 U12902 ( .A(n12941), .B(n12942), .Z(n12723) );
  XOR2_X1 U12903 ( .A(n12943), .B(n12944), .Z(n12942) );
  XOR2_X1 U12904 ( .A(n12945), .B(n12946), .Z(n12727) );
  XOR2_X1 U12905 ( .A(n12947), .B(n12948), .Z(n12946) );
  XOR2_X1 U12906 ( .A(n12949), .B(n12950), .Z(n12731) );
  XOR2_X1 U12907 ( .A(n12951), .B(n12952), .Z(n12950) );
  XOR2_X1 U12908 ( .A(n7752), .B(n12953), .Z(n12738) );
  XOR2_X1 U12909 ( .A(n7751), .B(n7750), .Z(n12953) );
  OR2_X1 U12910 ( .A1(n12612), .A2(n7621), .ZN(n7750) );
  OR2_X1 U12911 ( .A1(n12954), .A2(n12955), .ZN(n7751) );
  AND2_X1 U12912 ( .A1(n12952), .A2(n12951), .ZN(n12955) );
  AND2_X1 U12913 ( .A1(n12949), .A2(n12956), .ZN(n12954) );
  OR2_X1 U12914 ( .A1(n12951), .A2(n12952), .ZN(n12956) );
  OR2_X1 U12915 ( .A1(n12612), .A2(n7656), .ZN(n12952) );
  OR2_X1 U12916 ( .A1(n12957), .A2(n12958), .ZN(n12951) );
  AND2_X1 U12917 ( .A1(n12948), .A2(n12947), .ZN(n12958) );
  AND2_X1 U12918 ( .A1(n12945), .A2(n12959), .ZN(n12957) );
  OR2_X1 U12919 ( .A1(n12947), .A2(n12948), .ZN(n12959) );
  OR2_X1 U12920 ( .A1(n12612), .A2(n7689), .ZN(n12948) );
  OR2_X1 U12921 ( .A1(n12960), .A2(n12961), .ZN(n12947) );
  AND2_X1 U12922 ( .A1(n12944), .A2(n12943), .ZN(n12961) );
  AND2_X1 U12923 ( .A1(n12941), .A2(n12962), .ZN(n12960) );
  OR2_X1 U12924 ( .A1(n12943), .A2(n12944), .ZN(n12962) );
  OR2_X1 U12925 ( .A1(n12612), .A2(n7777), .ZN(n12944) );
  OR2_X1 U12926 ( .A1(n12963), .A2(n12964), .ZN(n12943) );
  AND2_X1 U12927 ( .A1(n12940), .A2(n12939), .ZN(n12964) );
  AND2_X1 U12928 ( .A1(n12937), .A2(n12965), .ZN(n12963) );
  OR2_X1 U12929 ( .A1(n12939), .A2(n12940), .ZN(n12965) );
  OR2_X1 U12930 ( .A1(n12612), .A2(n7785), .ZN(n12940) );
  OR2_X1 U12931 ( .A1(n12966), .A2(n12967), .ZN(n12939) );
  AND2_X1 U12932 ( .A1(n12936), .A2(n12935), .ZN(n12967) );
  AND2_X1 U12933 ( .A1(n12933), .A2(n12968), .ZN(n12966) );
  OR2_X1 U12934 ( .A1(n12935), .A2(n12936), .ZN(n12968) );
  OR2_X1 U12935 ( .A1(n12612), .A2(n8226), .ZN(n12936) );
  OR2_X1 U12936 ( .A1(n12969), .A2(n12970), .ZN(n12935) );
  AND2_X1 U12937 ( .A1(n12932), .A2(n12931), .ZN(n12970) );
  AND2_X1 U12938 ( .A1(n12929), .A2(n12971), .ZN(n12969) );
  OR2_X1 U12939 ( .A1(n12931), .A2(n12932), .ZN(n12971) );
  OR2_X1 U12940 ( .A1(n12612), .A2(n8221), .ZN(n12932) );
  OR2_X1 U12941 ( .A1(n12972), .A2(n12973), .ZN(n12931) );
  AND2_X1 U12942 ( .A1(n12928), .A2(n12927), .ZN(n12973) );
  AND2_X1 U12943 ( .A1(n12925), .A2(n12974), .ZN(n12972) );
  OR2_X1 U12944 ( .A1(n12927), .A2(n12928), .ZN(n12974) );
  OR2_X1 U12945 ( .A1(n12612), .A2(n8216), .ZN(n12928) );
  OR2_X1 U12946 ( .A1(n12975), .A2(n12976), .ZN(n12927) );
  AND2_X1 U12947 ( .A1(n12922), .A2(n12924), .ZN(n12976) );
  AND2_X1 U12948 ( .A1(n12977), .A2(n12923), .ZN(n12975) );
  OR2_X1 U12949 ( .A1(n12922), .A2(n12924), .ZN(n12977) );
  OR2_X1 U12950 ( .A1(n12978), .A2(n12979), .ZN(n12924) );
  AND2_X1 U12951 ( .A1(n12920), .A2(n12919), .ZN(n12979) );
  AND2_X1 U12952 ( .A1(n12917), .A2(n12980), .ZN(n12978) );
  OR2_X1 U12953 ( .A1(n12919), .A2(n12920), .ZN(n12980) );
  OR2_X1 U12954 ( .A1(n12612), .A2(n8206), .ZN(n12920) );
  OR2_X1 U12955 ( .A1(n12981), .A2(n12982), .ZN(n12919) );
  AND2_X1 U12956 ( .A1(n12916), .A2(n12915), .ZN(n12982) );
  AND2_X1 U12957 ( .A1(n12913), .A2(n12983), .ZN(n12981) );
  OR2_X1 U12958 ( .A1(n12915), .A2(n12916), .ZN(n12983) );
  OR2_X1 U12959 ( .A1(n12612), .A2(n8201), .ZN(n12916) );
  OR2_X1 U12960 ( .A1(n12984), .A2(n12985), .ZN(n12915) );
  AND2_X1 U12961 ( .A1(n12912), .A2(n12911), .ZN(n12985) );
  AND2_X1 U12962 ( .A1(n12909), .A2(n12986), .ZN(n12984) );
  OR2_X1 U12963 ( .A1(n12911), .A2(n12912), .ZN(n12986) );
  OR2_X1 U12964 ( .A1(n12612), .A2(n8196), .ZN(n12912) );
  OR2_X1 U12965 ( .A1(n12987), .A2(n12988), .ZN(n12911) );
  AND2_X1 U12966 ( .A1(n12908), .A2(n12907), .ZN(n12988) );
  AND2_X1 U12967 ( .A1(n12905), .A2(n12989), .ZN(n12987) );
  OR2_X1 U12968 ( .A1(n12907), .A2(n12908), .ZN(n12989) );
  OR2_X1 U12969 ( .A1(n12612), .A2(n8191), .ZN(n12908) );
  OR2_X1 U12970 ( .A1(n12990), .A2(n12991), .ZN(n12907) );
  AND2_X1 U12971 ( .A1(n12904), .A2(n12903), .ZN(n12991) );
  AND2_X1 U12972 ( .A1(n12901), .A2(n12992), .ZN(n12990) );
  OR2_X1 U12973 ( .A1(n12903), .A2(n12904), .ZN(n12992) );
  OR2_X1 U12974 ( .A1(n12612), .A2(n8186), .ZN(n12904) );
  OR2_X1 U12975 ( .A1(n12993), .A2(n12994), .ZN(n12903) );
  AND2_X1 U12976 ( .A1(n12900), .A2(n12899), .ZN(n12994) );
  AND2_X1 U12977 ( .A1(n12897), .A2(n12995), .ZN(n12993) );
  OR2_X1 U12978 ( .A1(n12899), .A2(n12900), .ZN(n12995) );
  OR2_X1 U12979 ( .A1(n12612), .A2(n8181), .ZN(n12900) );
  OR2_X1 U12980 ( .A1(n12996), .A2(n12997), .ZN(n12899) );
  AND2_X1 U12981 ( .A1(n12896), .A2(n12895), .ZN(n12997) );
  AND2_X1 U12982 ( .A1(n12893), .A2(n12998), .ZN(n12996) );
  OR2_X1 U12983 ( .A1(n12895), .A2(n12896), .ZN(n12998) );
  OR2_X1 U12984 ( .A1(n12612), .A2(n8176), .ZN(n12896) );
  OR2_X1 U12985 ( .A1(n12999), .A2(n13000), .ZN(n12895) );
  AND2_X1 U12986 ( .A1(n12892), .A2(n12891), .ZN(n13000) );
  AND2_X1 U12987 ( .A1(n12889), .A2(n13001), .ZN(n12999) );
  OR2_X1 U12988 ( .A1(n12891), .A2(n12892), .ZN(n13001) );
  OR2_X1 U12989 ( .A1(n12612), .A2(n8171), .ZN(n12892) );
  OR2_X1 U12990 ( .A1(n13002), .A2(n13003), .ZN(n12891) );
  AND2_X1 U12991 ( .A1(n12888), .A2(n12887), .ZN(n13003) );
  AND2_X1 U12992 ( .A1(n12885), .A2(n13004), .ZN(n13002) );
  OR2_X1 U12993 ( .A1(n12887), .A2(n12888), .ZN(n13004) );
  OR2_X1 U12994 ( .A1(n8166), .A2(n12612), .ZN(n12888) );
  OR2_X1 U12995 ( .A1(n13005), .A2(n13006), .ZN(n12887) );
  AND2_X1 U12996 ( .A1(n12884), .A2(n12883), .ZN(n13006) );
  AND2_X1 U12997 ( .A1(n12881), .A2(n13007), .ZN(n13005) );
  OR2_X1 U12998 ( .A1(n12883), .A2(n12884), .ZN(n13007) );
  OR2_X1 U12999 ( .A1(n12612), .A2(n8161), .ZN(n12884) );
  OR2_X1 U13000 ( .A1(n13008), .A2(n13009), .ZN(n12883) );
  AND2_X1 U13001 ( .A1(n12880), .A2(n12879), .ZN(n13009) );
  AND2_X1 U13002 ( .A1(n12877), .A2(n13010), .ZN(n13008) );
  OR2_X1 U13003 ( .A1(n12879), .A2(n12880), .ZN(n13010) );
  OR2_X1 U13004 ( .A1(n12612), .A2(n8156), .ZN(n12880) );
  OR2_X1 U13005 ( .A1(n13011), .A2(n13012), .ZN(n12879) );
  AND2_X1 U13006 ( .A1(n12876), .A2(n12875), .ZN(n13012) );
  AND2_X1 U13007 ( .A1(n12873), .A2(n13013), .ZN(n13011) );
  OR2_X1 U13008 ( .A1(n12875), .A2(n12876), .ZN(n13013) );
  OR2_X1 U13009 ( .A1(n12612), .A2(n8151), .ZN(n12876) );
  OR2_X1 U13010 ( .A1(n13014), .A2(n13015), .ZN(n12875) );
  AND2_X1 U13011 ( .A1(n12869), .A2(n12872), .ZN(n13015) );
  AND2_X1 U13012 ( .A1(n13016), .A2(n12871), .ZN(n13014) );
  OR2_X1 U13013 ( .A1(n13017), .A2(n13018), .ZN(n12871) );
  AND2_X1 U13014 ( .A1(n12868), .A2(n12867), .ZN(n13018) );
  AND2_X1 U13015 ( .A1(n12865), .A2(n13019), .ZN(n13017) );
  OR2_X1 U13016 ( .A1(n12867), .A2(n12868), .ZN(n13019) );
  OR2_X1 U13017 ( .A1(n8141), .A2(n12612), .ZN(n12868) );
  OR2_X1 U13018 ( .A1(n13020), .A2(n13021), .ZN(n12867) );
  AND2_X1 U13019 ( .A1(n12861), .A2(n12864), .ZN(n13021) );
  AND2_X1 U13020 ( .A1(n13022), .A2(n12863), .ZN(n13020) );
  OR2_X1 U13021 ( .A1(n13023), .A2(n13024), .ZN(n12863) );
  AND2_X1 U13022 ( .A1(n12857), .A2(n12860), .ZN(n13024) );
  AND2_X1 U13023 ( .A1(n13025), .A2(n12859), .ZN(n13023) );
  OR2_X1 U13024 ( .A1(n13026), .A2(n13027), .ZN(n12859) );
  AND2_X1 U13025 ( .A1(n12853), .A2(n12856), .ZN(n13027) );
  AND2_X1 U13026 ( .A1(n13028), .A2(n12855), .ZN(n13026) );
  OR2_X1 U13027 ( .A1(n13029), .A2(n13030), .ZN(n12855) );
  AND2_X1 U13028 ( .A1(n12849), .A2(n12852), .ZN(n13030) );
  AND2_X1 U13029 ( .A1(n13031), .A2(n12851), .ZN(n13029) );
  OR2_X1 U13030 ( .A1(n13032), .A2(n13033), .ZN(n12851) );
  AND2_X1 U13031 ( .A1(n12845), .A2(n12848), .ZN(n13033) );
  AND2_X1 U13032 ( .A1(n13034), .A2(n12847), .ZN(n13032) );
  OR2_X1 U13033 ( .A1(n13035), .A2(n13036), .ZN(n12847) );
  AND2_X1 U13034 ( .A1(n12841), .A2(n12844), .ZN(n13036) );
  AND2_X1 U13035 ( .A1(n13037), .A2(n12843), .ZN(n13035) );
  OR2_X1 U13036 ( .A1(n13038), .A2(n13039), .ZN(n12843) );
  AND2_X1 U13037 ( .A1(n12837), .A2(n12840), .ZN(n13039) );
  AND2_X1 U13038 ( .A1(n12839), .A2(n13040), .ZN(n13038) );
  OR2_X1 U13039 ( .A1(n12840), .A2(n12837), .ZN(n13040) );
  OR2_X1 U13040 ( .A1(n8102), .A2(n12612), .ZN(n12837) );
  OR3_X1 U13041 ( .A1(n8349), .A2(n12612), .A3(n7755), .ZN(n12840) );
  INV_X1 U13042 ( .A(n13041), .ZN(n12839) );
  OR2_X1 U13043 ( .A1(n13042), .A2(n13043), .ZN(n13041) );
  AND2_X1 U13044 ( .A1(b_7_), .A2(n13044), .ZN(n13043) );
  OR2_X1 U13045 ( .A1(n13045), .A2(n7314), .ZN(n13044) );
  AND2_X1 U13046 ( .A1(a_30_), .A2(n7716), .ZN(n13045) );
  AND2_X1 U13047 ( .A1(b_6_), .A2(n13046), .ZN(n13042) );
  OR2_X1 U13048 ( .A1(n13047), .A2(n7318), .ZN(n13046) );
  AND2_X1 U13049 ( .A1(a_31_), .A2(n7755), .ZN(n13047) );
  OR2_X1 U13050 ( .A1(n12844), .A2(n12841), .ZN(n13037) );
  XNOR2_X1 U13051 ( .A(n13048), .B(n13049), .ZN(n12841) );
  XNOR2_X1 U13052 ( .A(n13050), .B(n13051), .ZN(n13049) );
  OR2_X1 U13053 ( .A1(n8111), .A2(n12612), .ZN(n12844) );
  OR2_X1 U13054 ( .A1(n12848), .A2(n12845), .ZN(n13034) );
  XOR2_X1 U13055 ( .A(n13052), .B(n13053), .Z(n12845) );
  XOR2_X1 U13056 ( .A(n13054), .B(n13055), .Z(n13053) );
  OR2_X1 U13057 ( .A1(n8116), .A2(n12612), .ZN(n12848) );
  OR2_X1 U13058 ( .A1(n12852), .A2(n12849), .ZN(n13031) );
  XOR2_X1 U13059 ( .A(n13056), .B(n13057), .Z(n12849) );
  XOR2_X1 U13060 ( .A(n13058), .B(n13059), .Z(n13057) );
  OR2_X1 U13061 ( .A1(n8121), .A2(n12612), .ZN(n12852) );
  OR2_X1 U13062 ( .A1(n12856), .A2(n12853), .ZN(n13028) );
  XOR2_X1 U13063 ( .A(n13060), .B(n13061), .Z(n12853) );
  XOR2_X1 U13064 ( .A(n13062), .B(n13063), .Z(n13061) );
  OR2_X1 U13065 ( .A1(n8126), .A2(n12612), .ZN(n12856) );
  OR2_X1 U13066 ( .A1(n12860), .A2(n12857), .ZN(n13025) );
  XOR2_X1 U13067 ( .A(n13064), .B(n13065), .Z(n12857) );
  XOR2_X1 U13068 ( .A(n13066), .B(n13067), .Z(n13065) );
  OR2_X1 U13069 ( .A1(n8131), .A2(n12612), .ZN(n12860) );
  OR2_X1 U13070 ( .A1(n12864), .A2(n12861), .ZN(n13022) );
  XOR2_X1 U13071 ( .A(n13068), .B(n13069), .Z(n12861) );
  XOR2_X1 U13072 ( .A(n13070), .B(n13071), .Z(n13069) );
  OR2_X1 U13073 ( .A1(n8136), .A2(n12612), .ZN(n12864) );
  XOR2_X1 U13074 ( .A(n13072), .B(n13073), .Z(n12865) );
  XOR2_X1 U13075 ( .A(n13074), .B(n13075), .Z(n13073) );
  OR2_X1 U13076 ( .A1(n12872), .A2(n12869), .ZN(n13016) );
  XOR2_X1 U13077 ( .A(n13076), .B(n13077), .Z(n12869) );
  XOR2_X1 U13078 ( .A(n13078), .B(n13079), .Z(n13077) );
  OR2_X1 U13079 ( .A1(n12612), .A2(n8146), .ZN(n12872) );
  XOR2_X1 U13080 ( .A(n13080), .B(n13081), .Z(n12873) );
  XOR2_X1 U13081 ( .A(n13082), .B(n13083), .Z(n13081) );
  XOR2_X1 U13082 ( .A(n13084), .B(n13085), .Z(n12877) );
  XOR2_X1 U13083 ( .A(n13086), .B(n13087), .Z(n13085) );
  XOR2_X1 U13084 ( .A(n13088), .B(n13089), .Z(n12881) );
  XOR2_X1 U13085 ( .A(n13090), .B(n13091), .Z(n13089) );
  XOR2_X1 U13086 ( .A(n13092), .B(n13093), .Z(n12885) );
  XOR2_X1 U13087 ( .A(n13094), .B(n13095), .Z(n13093) );
  XOR2_X1 U13088 ( .A(n13096), .B(n13097), .Z(n12889) );
  XOR2_X1 U13089 ( .A(n13098), .B(n13099), .Z(n13097) );
  XOR2_X1 U13090 ( .A(n13100), .B(n13101), .Z(n12893) );
  XOR2_X1 U13091 ( .A(n13102), .B(n13103), .Z(n13101) );
  XOR2_X1 U13092 ( .A(n13104), .B(n13105), .Z(n12897) );
  XOR2_X1 U13093 ( .A(n13106), .B(n13107), .Z(n13105) );
  XOR2_X1 U13094 ( .A(n13108), .B(n13109), .Z(n12901) );
  XOR2_X1 U13095 ( .A(n13110), .B(n13111), .Z(n13109) );
  XOR2_X1 U13096 ( .A(n13112), .B(n13113), .Z(n12905) );
  XOR2_X1 U13097 ( .A(n13114), .B(n13115), .Z(n13113) );
  XOR2_X1 U13098 ( .A(n13116), .B(n13117), .Z(n12909) );
  XOR2_X1 U13099 ( .A(n13118), .B(n13119), .Z(n13117) );
  XOR2_X1 U13100 ( .A(n13120), .B(n13121), .Z(n12913) );
  XOR2_X1 U13101 ( .A(n13122), .B(n13123), .Z(n13121) );
  XOR2_X1 U13102 ( .A(n13124), .B(n13125), .Z(n12917) );
  XOR2_X1 U13103 ( .A(n13126), .B(n13127), .Z(n13125) );
  XOR2_X1 U13104 ( .A(n13128), .B(n13129), .Z(n12922) );
  XOR2_X1 U13105 ( .A(n13130), .B(n13131), .Z(n13129) );
  XOR2_X1 U13106 ( .A(n13132), .B(n13133), .Z(n12925) );
  XOR2_X1 U13107 ( .A(n13134), .B(n13135), .Z(n13133) );
  XNOR2_X1 U13108 ( .A(n13136), .B(n13137), .ZN(n12929) );
  XNOR2_X1 U13109 ( .A(n13138), .B(n13139), .ZN(n13136) );
  XOR2_X1 U13110 ( .A(n13140), .B(n13141), .Z(n12933) );
  XOR2_X1 U13111 ( .A(n13142), .B(n13143), .Z(n13141) );
  XOR2_X1 U13112 ( .A(n13144), .B(n13145), .Z(n12937) );
  XOR2_X1 U13113 ( .A(n13146), .B(n13147), .Z(n13145) );
  XOR2_X1 U13114 ( .A(n13148), .B(n13149), .Z(n12941) );
  XOR2_X1 U13115 ( .A(n13150), .B(n13151), .Z(n13149) );
  XOR2_X1 U13116 ( .A(n13152), .B(n13153), .Z(n12945) );
  XOR2_X1 U13117 ( .A(n13154), .B(n13155), .Z(n13153) );
  XOR2_X1 U13118 ( .A(n13156), .B(n13157), .Z(n12949) );
  XOR2_X1 U13119 ( .A(n13158), .B(n13159), .Z(n13157) );
  XOR2_X1 U13120 ( .A(n7760), .B(n13160), .Z(n7752) );
  XOR2_X1 U13121 ( .A(n7759), .B(n7758), .Z(n13160) );
  OR2_X1 U13122 ( .A1(n7755), .A2(n7656), .ZN(n7758) );
  OR2_X1 U13123 ( .A1(n13161), .A2(n13162), .ZN(n7759) );
  AND2_X1 U13124 ( .A1(n13159), .A2(n13158), .ZN(n13162) );
  AND2_X1 U13125 ( .A1(n13156), .A2(n13163), .ZN(n13161) );
  OR2_X1 U13126 ( .A1(n13158), .A2(n13159), .ZN(n13163) );
  OR2_X1 U13127 ( .A1(n7755), .A2(n7689), .ZN(n13159) );
  OR2_X1 U13128 ( .A1(n13164), .A2(n13165), .ZN(n13158) );
  AND2_X1 U13129 ( .A1(n13155), .A2(n13154), .ZN(n13165) );
  AND2_X1 U13130 ( .A1(n13152), .A2(n13166), .ZN(n13164) );
  OR2_X1 U13131 ( .A1(n13154), .A2(n13155), .ZN(n13166) );
  OR2_X1 U13132 ( .A1(n7755), .A2(n7777), .ZN(n13155) );
  OR2_X1 U13133 ( .A1(n13167), .A2(n13168), .ZN(n13154) );
  AND2_X1 U13134 ( .A1(n13151), .A2(n13150), .ZN(n13168) );
  AND2_X1 U13135 ( .A1(n13148), .A2(n13169), .ZN(n13167) );
  OR2_X1 U13136 ( .A1(n13150), .A2(n13151), .ZN(n13169) );
  OR2_X1 U13137 ( .A1(n7755), .A2(n7785), .ZN(n13151) );
  OR2_X1 U13138 ( .A1(n13170), .A2(n13171), .ZN(n13150) );
  AND2_X1 U13139 ( .A1(n13147), .A2(n13146), .ZN(n13171) );
  AND2_X1 U13140 ( .A1(n13144), .A2(n13172), .ZN(n13170) );
  OR2_X1 U13141 ( .A1(n13146), .A2(n13147), .ZN(n13172) );
  OR2_X1 U13142 ( .A1(n7755), .A2(n8226), .ZN(n13147) );
  OR2_X1 U13143 ( .A1(n13173), .A2(n13174), .ZN(n13146) );
  AND2_X1 U13144 ( .A1(n13143), .A2(n13142), .ZN(n13174) );
  AND2_X1 U13145 ( .A1(n13140), .A2(n13175), .ZN(n13173) );
  OR2_X1 U13146 ( .A1(n13142), .A2(n13143), .ZN(n13175) );
  OR2_X1 U13147 ( .A1(n7755), .A2(n8221), .ZN(n13143) );
  OR2_X1 U13148 ( .A1(n13176), .A2(n13177), .ZN(n13142) );
  AND2_X1 U13149 ( .A1(n13137), .A2(n13139), .ZN(n13177) );
  AND2_X1 U13150 ( .A1(n13178), .A2(n13138), .ZN(n13176) );
  OR2_X1 U13151 ( .A1(n13137), .A2(n13139), .ZN(n13178) );
  OR2_X1 U13152 ( .A1(n13179), .A2(n13180), .ZN(n13139) );
  AND2_X1 U13153 ( .A1(n13135), .A2(n13134), .ZN(n13180) );
  AND2_X1 U13154 ( .A1(n13132), .A2(n13181), .ZN(n13179) );
  OR2_X1 U13155 ( .A1(n13134), .A2(n13135), .ZN(n13181) );
  OR2_X1 U13156 ( .A1(n7755), .A2(n8211), .ZN(n13135) );
  OR2_X1 U13157 ( .A1(n13182), .A2(n13183), .ZN(n13134) );
  AND2_X1 U13158 ( .A1(n13131), .A2(n13130), .ZN(n13183) );
  AND2_X1 U13159 ( .A1(n13128), .A2(n13184), .ZN(n13182) );
  OR2_X1 U13160 ( .A1(n13130), .A2(n13131), .ZN(n13184) );
  OR2_X1 U13161 ( .A1(n7755), .A2(n8206), .ZN(n13131) );
  OR2_X1 U13162 ( .A1(n13185), .A2(n13186), .ZN(n13130) );
  AND2_X1 U13163 ( .A1(n13127), .A2(n13126), .ZN(n13186) );
  AND2_X1 U13164 ( .A1(n13124), .A2(n13187), .ZN(n13185) );
  OR2_X1 U13165 ( .A1(n13126), .A2(n13127), .ZN(n13187) );
  OR2_X1 U13166 ( .A1(n7755), .A2(n8201), .ZN(n13127) );
  OR2_X1 U13167 ( .A1(n13188), .A2(n13189), .ZN(n13126) );
  AND2_X1 U13168 ( .A1(n13123), .A2(n13122), .ZN(n13189) );
  AND2_X1 U13169 ( .A1(n13120), .A2(n13190), .ZN(n13188) );
  OR2_X1 U13170 ( .A1(n13122), .A2(n13123), .ZN(n13190) );
  OR2_X1 U13171 ( .A1(n7755), .A2(n8196), .ZN(n13123) );
  OR2_X1 U13172 ( .A1(n13191), .A2(n13192), .ZN(n13122) );
  AND2_X1 U13173 ( .A1(n13119), .A2(n13118), .ZN(n13192) );
  AND2_X1 U13174 ( .A1(n13116), .A2(n13193), .ZN(n13191) );
  OR2_X1 U13175 ( .A1(n13118), .A2(n13119), .ZN(n13193) );
  OR2_X1 U13176 ( .A1(n7755), .A2(n8191), .ZN(n13119) );
  OR2_X1 U13177 ( .A1(n13194), .A2(n13195), .ZN(n13118) );
  AND2_X1 U13178 ( .A1(n13115), .A2(n13114), .ZN(n13195) );
  AND2_X1 U13179 ( .A1(n13112), .A2(n13196), .ZN(n13194) );
  OR2_X1 U13180 ( .A1(n13114), .A2(n13115), .ZN(n13196) );
  OR2_X1 U13181 ( .A1(n7755), .A2(n8186), .ZN(n13115) );
  OR2_X1 U13182 ( .A1(n13197), .A2(n13198), .ZN(n13114) );
  AND2_X1 U13183 ( .A1(n13111), .A2(n13110), .ZN(n13198) );
  AND2_X1 U13184 ( .A1(n13108), .A2(n13199), .ZN(n13197) );
  OR2_X1 U13185 ( .A1(n13110), .A2(n13111), .ZN(n13199) );
  OR2_X1 U13186 ( .A1(n7755), .A2(n8181), .ZN(n13111) );
  OR2_X1 U13187 ( .A1(n13200), .A2(n13201), .ZN(n13110) );
  AND2_X1 U13188 ( .A1(n13107), .A2(n13106), .ZN(n13201) );
  AND2_X1 U13189 ( .A1(n13104), .A2(n13202), .ZN(n13200) );
  OR2_X1 U13190 ( .A1(n13106), .A2(n13107), .ZN(n13202) );
  OR2_X1 U13191 ( .A1(n7755), .A2(n8176), .ZN(n13107) );
  OR2_X1 U13192 ( .A1(n13203), .A2(n13204), .ZN(n13106) );
  AND2_X1 U13193 ( .A1(n13103), .A2(n13102), .ZN(n13204) );
  AND2_X1 U13194 ( .A1(n13100), .A2(n13205), .ZN(n13203) );
  OR2_X1 U13195 ( .A1(n13102), .A2(n13103), .ZN(n13205) );
  OR2_X1 U13196 ( .A1(n7755), .A2(n8171), .ZN(n13103) );
  OR2_X1 U13197 ( .A1(n13206), .A2(n13207), .ZN(n13102) );
  AND2_X1 U13198 ( .A1(n13099), .A2(n13098), .ZN(n13207) );
  AND2_X1 U13199 ( .A1(n13096), .A2(n13208), .ZN(n13206) );
  OR2_X1 U13200 ( .A1(n13098), .A2(n13099), .ZN(n13208) );
  OR2_X1 U13201 ( .A1(n8166), .A2(n7755), .ZN(n13099) );
  OR2_X1 U13202 ( .A1(n13209), .A2(n13210), .ZN(n13098) );
  AND2_X1 U13203 ( .A1(n13095), .A2(n13094), .ZN(n13210) );
  AND2_X1 U13204 ( .A1(n13092), .A2(n13211), .ZN(n13209) );
  OR2_X1 U13205 ( .A1(n13094), .A2(n13095), .ZN(n13211) );
  OR2_X1 U13206 ( .A1(n7755), .A2(n8161), .ZN(n13095) );
  OR2_X1 U13207 ( .A1(n13212), .A2(n13213), .ZN(n13094) );
  AND2_X1 U13208 ( .A1(n13091), .A2(n13090), .ZN(n13213) );
  AND2_X1 U13209 ( .A1(n13088), .A2(n13214), .ZN(n13212) );
  OR2_X1 U13210 ( .A1(n13090), .A2(n13091), .ZN(n13214) );
  OR2_X1 U13211 ( .A1(n7755), .A2(n8156), .ZN(n13091) );
  OR2_X1 U13212 ( .A1(n13215), .A2(n13216), .ZN(n13090) );
  AND2_X1 U13213 ( .A1(n13087), .A2(n13086), .ZN(n13216) );
  AND2_X1 U13214 ( .A1(n13084), .A2(n13217), .ZN(n13215) );
  OR2_X1 U13215 ( .A1(n13086), .A2(n13087), .ZN(n13217) );
  OR2_X1 U13216 ( .A1(n7755), .A2(n8151), .ZN(n13087) );
  OR2_X1 U13217 ( .A1(n13218), .A2(n13219), .ZN(n13086) );
  AND2_X1 U13218 ( .A1(n13083), .A2(n13082), .ZN(n13219) );
  AND2_X1 U13219 ( .A1(n13080), .A2(n13220), .ZN(n13218) );
  OR2_X1 U13220 ( .A1(n13082), .A2(n13083), .ZN(n13220) );
  OR2_X1 U13221 ( .A1(n8146), .A2(n7755), .ZN(n13083) );
  OR2_X1 U13222 ( .A1(n13221), .A2(n13222), .ZN(n13082) );
  AND2_X1 U13223 ( .A1(n13076), .A2(n13079), .ZN(n13222) );
  AND2_X1 U13224 ( .A1(n13223), .A2(n13078), .ZN(n13221) );
  OR2_X1 U13225 ( .A1(n13224), .A2(n13225), .ZN(n13078) );
  AND2_X1 U13226 ( .A1(n13075), .A2(n13074), .ZN(n13225) );
  AND2_X1 U13227 ( .A1(n13072), .A2(n13226), .ZN(n13224) );
  OR2_X1 U13228 ( .A1(n13074), .A2(n13075), .ZN(n13226) );
  OR2_X1 U13229 ( .A1(n8136), .A2(n7755), .ZN(n13075) );
  OR2_X1 U13230 ( .A1(n13227), .A2(n13228), .ZN(n13074) );
  AND2_X1 U13231 ( .A1(n13068), .A2(n13071), .ZN(n13228) );
  AND2_X1 U13232 ( .A1(n13229), .A2(n13070), .ZN(n13227) );
  OR2_X1 U13233 ( .A1(n13230), .A2(n13231), .ZN(n13070) );
  AND2_X1 U13234 ( .A1(n13064), .A2(n13067), .ZN(n13231) );
  AND2_X1 U13235 ( .A1(n13232), .A2(n13066), .ZN(n13230) );
  OR2_X1 U13236 ( .A1(n13233), .A2(n13234), .ZN(n13066) );
  AND2_X1 U13237 ( .A1(n13060), .A2(n13063), .ZN(n13234) );
  AND2_X1 U13238 ( .A1(n13235), .A2(n13062), .ZN(n13233) );
  OR2_X1 U13239 ( .A1(n13236), .A2(n13237), .ZN(n13062) );
  AND2_X1 U13240 ( .A1(n13056), .A2(n13059), .ZN(n13237) );
  AND2_X1 U13241 ( .A1(n13238), .A2(n13058), .ZN(n13236) );
  OR2_X1 U13242 ( .A1(n13239), .A2(n13240), .ZN(n13058) );
  AND2_X1 U13243 ( .A1(n13052), .A2(n13055), .ZN(n13240) );
  AND2_X1 U13244 ( .A1(n13241), .A2(n13054), .ZN(n13239) );
  OR2_X1 U13245 ( .A1(n13242), .A2(n13243), .ZN(n13054) );
  AND2_X1 U13246 ( .A1(n13048), .A2(n13051), .ZN(n13243) );
  AND2_X1 U13247 ( .A1(n13050), .A2(n13244), .ZN(n13242) );
  OR2_X1 U13248 ( .A1(n13051), .A2(n13048), .ZN(n13244) );
  OR2_X1 U13249 ( .A1(n8102), .A2(n7755), .ZN(n13048) );
  OR3_X1 U13250 ( .A1(n8349), .A2(n7755), .A3(n7716), .ZN(n13051) );
  INV_X1 U13251 ( .A(n13245), .ZN(n13050) );
  OR2_X1 U13252 ( .A1(n13246), .A2(n13247), .ZN(n13245) );
  AND2_X1 U13253 ( .A1(b_6_), .A2(n13248), .ZN(n13247) );
  OR2_X1 U13254 ( .A1(n13249), .A2(n7314), .ZN(n13248) );
  AND2_X1 U13255 ( .A1(a_30_), .A2(n7674), .ZN(n13249) );
  AND2_X1 U13256 ( .A1(b_5_), .A2(n13250), .ZN(n13246) );
  OR2_X1 U13257 ( .A1(n13251), .A2(n7318), .ZN(n13250) );
  AND2_X1 U13258 ( .A1(a_31_), .A2(n7716), .ZN(n13251) );
  OR2_X1 U13259 ( .A1(n13055), .A2(n13052), .ZN(n13241) );
  XNOR2_X1 U13260 ( .A(n13252), .B(n13253), .ZN(n13052) );
  XNOR2_X1 U13261 ( .A(n13254), .B(n13255), .ZN(n13253) );
  OR2_X1 U13262 ( .A1(n8111), .A2(n7755), .ZN(n13055) );
  OR2_X1 U13263 ( .A1(n13059), .A2(n13056), .ZN(n13238) );
  XOR2_X1 U13264 ( .A(n13256), .B(n13257), .Z(n13056) );
  XOR2_X1 U13265 ( .A(n13258), .B(n13259), .Z(n13257) );
  OR2_X1 U13266 ( .A1(n8116), .A2(n7755), .ZN(n13059) );
  OR2_X1 U13267 ( .A1(n13063), .A2(n13060), .ZN(n13235) );
  XOR2_X1 U13268 ( .A(n13260), .B(n13261), .Z(n13060) );
  XOR2_X1 U13269 ( .A(n13262), .B(n13263), .Z(n13261) );
  OR2_X1 U13270 ( .A1(n8121), .A2(n7755), .ZN(n13063) );
  OR2_X1 U13271 ( .A1(n13067), .A2(n13064), .ZN(n13232) );
  XOR2_X1 U13272 ( .A(n13264), .B(n13265), .Z(n13064) );
  XOR2_X1 U13273 ( .A(n13266), .B(n13267), .Z(n13265) );
  OR2_X1 U13274 ( .A1(n8126), .A2(n7755), .ZN(n13067) );
  OR2_X1 U13275 ( .A1(n13071), .A2(n13068), .ZN(n13229) );
  XOR2_X1 U13276 ( .A(n13268), .B(n13269), .Z(n13068) );
  XOR2_X1 U13277 ( .A(n13270), .B(n13271), .Z(n13269) );
  OR2_X1 U13278 ( .A1(n8131), .A2(n7755), .ZN(n13071) );
  XOR2_X1 U13279 ( .A(n13272), .B(n13273), .Z(n13072) );
  XOR2_X1 U13280 ( .A(n13274), .B(n13275), .Z(n13273) );
  OR2_X1 U13281 ( .A1(n13079), .A2(n13076), .ZN(n13223) );
  XOR2_X1 U13282 ( .A(n13276), .B(n13277), .Z(n13076) );
  XOR2_X1 U13283 ( .A(n13278), .B(n13279), .Z(n13277) );
  OR2_X1 U13284 ( .A1(n8141), .A2(n7755), .ZN(n13079) );
  XOR2_X1 U13285 ( .A(n13280), .B(n13281), .Z(n13080) );
  XOR2_X1 U13286 ( .A(n13282), .B(n13283), .Z(n13281) );
  XOR2_X1 U13287 ( .A(n13284), .B(n13285), .Z(n13084) );
  XOR2_X1 U13288 ( .A(n13286), .B(n13287), .Z(n13285) );
  XOR2_X1 U13289 ( .A(n13288), .B(n13289), .Z(n13088) );
  XOR2_X1 U13290 ( .A(n13290), .B(n13291), .Z(n13289) );
  XOR2_X1 U13291 ( .A(n13292), .B(n13293), .Z(n13092) );
  XOR2_X1 U13292 ( .A(n13294), .B(n13295), .Z(n13293) );
  XOR2_X1 U13293 ( .A(n13296), .B(n13297), .Z(n13096) );
  XOR2_X1 U13294 ( .A(n13298), .B(n13299), .Z(n13297) );
  XOR2_X1 U13295 ( .A(n13300), .B(n13301), .Z(n13100) );
  XOR2_X1 U13296 ( .A(n13302), .B(n13303), .Z(n13301) );
  XOR2_X1 U13297 ( .A(n13304), .B(n13305), .Z(n13104) );
  XOR2_X1 U13298 ( .A(n13306), .B(n13307), .Z(n13305) );
  XOR2_X1 U13299 ( .A(n13308), .B(n13309), .Z(n13108) );
  XOR2_X1 U13300 ( .A(n13310), .B(n13311), .Z(n13309) );
  XOR2_X1 U13301 ( .A(n13312), .B(n13313), .Z(n13112) );
  XOR2_X1 U13302 ( .A(n13314), .B(n13315), .Z(n13313) );
  XOR2_X1 U13303 ( .A(n13316), .B(n13317), .Z(n13116) );
  XOR2_X1 U13304 ( .A(n13318), .B(n13319), .Z(n13317) );
  XOR2_X1 U13305 ( .A(n13320), .B(n13321), .Z(n13120) );
  XOR2_X1 U13306 ( .A(n13322), .B(n13323), .Z(n13321) );
  XOR2_X1 U13307 ( .A(n13324), .B(n13325), .Z(n13124) );
  XOR2_X1 U13308 ( .A(n13326), .B(n13327), .Z(n13325) );
  XOR2_X1 U13309 ( .A(n13328), .B(n13329), .Z(n13128) );
  XOR2_X1 U13310 ( .A(n13330), .B(n13331), .Z(n13329) );
  XOR2_X1 U13311 ( .A(n13332), .B(n13333), .Z(n13132) );
  XOR2_X1 U13312 ( .A(n13334), .B(n13335), .Z(n13333) );
  XOR2_X1 U13313 ( .A(n13336), .B(n13337), .Z(n13137) );
  XOR2_X1 U13314 ( .A(n13338), .B(n13339), .Z(n13337) );
  XOR2_X1 U13315 ( .A(n13340), .B(n13341), .Z(n13140) );
  XOR2_X1 U13316 ( .A(n13342), .B(n13343), .Z(n13341) );
  XNOR2_X1 U13317 ( .A(n13344), .B(n13345), .ZN(n13144) );
  XNOR2_X1 U13318 ( .A(n13346), .B(n13347), .ZN(n13344) );
  XOR2_X1 U13319 ( .A(n13348), .B(n13349), .Z(n13148) );
  XOR2_X1 U13320 ( .A(n13350), .B(n13351), .Z(n13349) );
  XOR2_X1 U13321 ( .A(n13352), .B(n13353), .Z(n13152) );
  XOR2_X1 U13322 ( .A(n13354), .B(n13355), .Z(n13353) );
  XOR2_X1 U13323 ( .A(n13356), .B(n13357), .Z(n13156) );
  XOR2_X1 U13324 ( .A(n13358), .B(n13359), .Z(n13357) );
  XOR2_X1 U13325 ( .A(n7767), .B(n13360), .Z(n7760) );
  XOR2_X1 U13326 ( .A(n7766), .B(n7765), .Z(n13360) );
  OR2_X1 U13327 ( .A1(n7716), .A2(n7689), .ZN(n7765) );
  OR2_X1 U13328 ( .A1(n13361), .A2(n13362), .ZN(n7766) );
  AND2_X1 U13329 ( .A1(n13359), .A2(n13358), .ZN(n13362) );
  AND2_X1 U13330 ( .A1(n13356), .A2(n13363), .ZN(n13361) );
  OR2_X1 U13331 ( .A1(n13358), .A2(n13359), .ZN(n13363) );
  OR2_X1 U13332 ( .A1(n7716), .A2(n7777), .ZN(n13359) );
  OR2_X1 U13333 ( .A1(n13364), .A2(n13365), .ZN(n13358) );
  AND2_X1 U13334 ( .A1(n13355), .A2(n13354), .ZN(n13365) );
  AND2_X1 U13335 ( .A1(n13352), .A2(n13366), .ZN(n13364) );
  OR2_X1 U13336 ( .A1(n13354), .A2(n13355), .ZN(n13366) );
  OR2_X1 U13337 ( .A1(n7716), .A2(n7785), .ZN(n13355) );
  OR2_X1 U13338 ( .A1(n13367), .A2(n13368), .ZN(n13354) );
  AND2_X1 U13339 ( .A1(n13351), .A2(n13350), .ZN(n13368) );
  AND2_X1 U13340 ( .A1(n13348), .A2(n13369), .ZN(n13367) );
  OR2_X1 U13341 ( .A1(n13350), .A2(n13351), .ZN(n13369) );
  OR2_X1 U13342 ( .A1(n7716), .A2(n8226), .ZN(n13351) );
  OR2_X1 U13343 ( .A1(n13370), .A2(n13371), .ZN(n13350) );
  AND2_X1 U13344 ( .A1(n13345), .A2(n13347), .ZN(n13371) );
  AND2_X1 U13345 ( .A1(n13372), .A2(n13346), .ZN(n13370) );
  OR2_X1 U13346 ( .A1(n13345), .A2(n13347), .ZN(n13372) );
  OR2_X1 U13347 ( .A1(n13373), .A2(n13374), .ZN(n13347) );
  AND2_X1 U13348 ( .A1(n13343), .A2(n13342), .ZN(n13374) );
  AND2_X1 U13349 ( .A1(n13340), .A2(n13375), .ZN(n13373) );
  OR2_X1 U13350 ( .A1(n13342), .A2(n13343), .ZN(n13375) );
  OR2_X1 U13351 ( .A1(n7716), .A2(n8216), .ZN(n13343) );
  OR2_X1 U13352 ( .A1(n13376), .A2(n13377), .ZN(n13342) );
  AND2_X1 U13353 ( .A1(n13339), .A2(n13338), .ZN(n13377) );
  AND2_X1 U13354 ( .A1(n13336), .A2(n13378), .ZN(n13376) );
  OR2_X1 U13355 ( .A1(n13338), .A2(n13339), .ZN(n13378) );
  OR2_X1 U13356 ( .A1(n7716), .A2(n8211), .ZN(n13339) );
  OR2_X1 U13357 ( .A1(n13379), .A2(n13380), .ZN(n13338) );
  AND2_X1 U13358 ( .A1(n13335), .A2(n13334), .ZN(n13380) );
  AND2_X1 U13359 ( .A1(n13332), .A2(n13381), .ZN(n13379) );
  OR2_X1 U13360 ( .A1(n13334), .A2(n13335), .ZN(n13381) );
  OR2_X1 U13361 ( .A1(n7716), .A2(n8206), .ZN(n13335) );
  OR2_X1 U13362 ( .A1(n13382), .A2(n13383), .ZN(n13334) );
  AND2_X1 U13363 ( .A1(n13331), .A2(n13330), .ZN(n13383) );
  AND2_X1 U13364 ( .A1(n13328), .A2(n13384), .ZN(n13382) );
  OR2_X1 U13365 ( .A1(n13330), .A2(n13331), .ZN(n13384) );
  OR2_X1 U13366 ( .A1(n7716), .A2(n8201), .ZN(n13331) );
  OR2_X1 U13367 ( .A1(n13385), .A2(n13386), .ZN(n13330) );
  AND2_X1 U13368 ( .A1(n13327), .A2(n13326), .ZN(n13386) );
  AND2_X1 U13369 ( .A1(n13324), .A2(n13387), .ZN(n13385) );
  OR2_X1 U13370 ( .A1(n13326), .A2(n13327), .ZN(n13387) );
  OR2_X1 U13371 ( .A1(n7716), .A2(n8196), .ZN(n13327) );
  OR2_X1 U13372 ( .A1(n13388), .A2(n13389), .ZN(n13326) );
  AND2_X1 U13373 ( .A1(n13323), .A2(n13322), .ZN(n13389) );
  AND2_X1 U13374 ( .A1(n13320), .A2(n13390), .ZN(n13388) );
  OR2_X1 U13375 ( .A1(n13322), .A2(n13323), .ZN(n13390) );
  OR2_X1 U13376 ( .A1(n7716), .A2(n8191), .ZN(n13323) );
  OR2_X1 U13377 ( .A1(n13391), .A2(n13392), .ZN(n13322) );
  AND2_X1 U13378 ( .A1(n13319), .A2(n13318), .ZN(n13392) );
  AND2_X1 U13379 ( .A1(n13316), .A2(n13393), .ZN(n13391) );
  OR2_X1 U13380 ( .A1(n13318), .A2(n13319), .ZN(n13393) );
  OR2_X1 U13381 ( .A1(n7716), .A2(n8186), .ZN(n13319) );
  OR2_X1 U13382 ( .A1(n13394), .A2(n13395), .ZN(n13318) );
  AND2_X1 U13383 ( .A1(n13315), .A2(n13314), .ZN(n13395) );
  AND2_X1 U13384 ( .A1(n13312), .A2(n13396), .ZN(n13394) );
  OR2_X1 U13385 ( .A1(n13314), .A2(n13315), .ZN(n13396) );
  OR2_X1 U13386 ( .A1(n7716), .A2(n8181), .ZN(n13315) );
  OR2_X1 U13387 ( .A1(n13397), .A2(n13398), .ZN(n13314) );
  AND2_X1 U13388 ( .A1(n13311), .A2(n13310), .ZN(n13398) );
  AND2_X1 U13389 ( .A1(n13308), .A2(n13399), .ZN(n13397) );
  OR2_X1 U13390 ( .A1(n13310), .A2(n13311), .ZN(n13399) );
  OR2_X1 U13391 ( .A1(n7716), .A2(n8176), .ZN(n13311) );
  OR2_X1 U13392 ( .A1(n13400), .A2(n13401), .ZN(n13310) );
  AND2_X1 U13393 ( .A1(n13307), .A2(n13306), .ZN(n13401) );
  AND2_X1 U13394 ( .A1(n13304), .A2(n13402), .ZN(n13400) );
  OR2_X1 U13395 ( .A1(n13306), .A2(n13307), .ZN(n13402) );
  OR2_X1 U13396 ( .A1(n7716), .A2(n8171), .ZN(n13307) );
  OR2_X1 U13397 ( .A1(n13403), .A2(n13404), .ZN(n13306) );
  AND2_X1 U13398 ( .A1(n13303), .A2(n13302), .ZN(n13404) );
  AND2_X1 U13399 ( .A1(n13300), .A2(n13405), .ZN(n13403) );
  OR2_X1 U13400 ( .A1(n13302), .A2(n13303), .ZN(n13405) );
  OR2_X1 U13401 ( .A1(n8166), .A2(n7716), .ZN(n13303) );
  OR2_X1 U13402 ( .A1(n13406), .A2(n13407), .ZN(n13302) );
  AND2_X1 U13403 ( .A1(n13299), .A2(n13298), .ZN(n13407) );
  AND2_X1 U13404 ( .A1(n13296), .A2(n13408), .ZN(n13406) );
  OR2_X1 U13405 ( .A1(n13298), .A2(n13299), .ZN(n13408) );
  OR2_X1 U13406 ( .A1(n7716), .A2(n8161), .ZN(n13299) );
  OR2_X1 U13407 ( .A1(n13409), .A2(n13410), .ZN(n13298) );
  AND2_X1 U13408 ( .A1(n13295), .A2(n13294), .ZN(n13410) );
  AND2_X1 U13409 ( .A1(n13292), .A2(n13411), .ZN(n13409) );
  OR2_X1 U13410 ( .A1(n13294), .A2(n13295), .ZN(n13411) );
  OR2_X1 U13411 ( .A1(n7716), .A2(n8156), .ZN(n13295) );
  OR2_X1 U13412 ( .A1(n13412), .A2(n13413), .ZN(n13294) );
  AND2_X1 U13413 ( .A1(n13291), .A2(n13290), .ZN(n13413) );
  AND2_X1 U13414 ( .A1(n13288), .A2(n13414), .ZN(n13412) );
  OR2_X1 U13415 ( .A1(n13290), .A2(n13291), .ZN(n13414) );
  OR2_X1 U13416 ( .A1(n8151), .A2(n7716), .ZN(n13291) );
  OR2_X1 U13417 ( .A1(n13415), .A2(n13416), .ZN(n13290) );
  AND2_X1 U13418 ( .A1(n13287), .A2(n13286), .ZN(n13416) );
  AND2_X1 U13419 ( .A1(n13284), .A2(n13417), .ZN(n13415) );
  OR2_X1 U13420 ( .A1(n13286), .A2(n13287), .ZN(n13417) );
  OR2_X1 U13421 ( .A1(n8146), .A2(n7716), .ZN(n13287) );
  OR2_X1 U13422 ( .A1(n13418), .A2(n13419), .ZN(n13286) );
  AND2_X1 U13423 ( .A1(n13283), .A2(n13282), .ZN(n13419) );
  AND2_X1 U13424 ( .A1(n13280), .A2(n13420), .ZN(n13418) );
  OR2_X1 U13425 ( .A1(n13282), .A2(n13283), .ZN(n13420) );
  OR2_X1 U13426 ( .A1(n8141), .A2(n7716), .ZN(n13283) );
  OR2_X1 U13427 ( .A1(n13421), .A2(n13422), .ZN(n13282) );
  AND2_X1 U13428 ( .A1(n13276), .A2(n13279), .ZN(n13422) );
  AND2_X1 U13429 ( .A1(n13423), .A2(n13278), .ZN(n13421) );
  OR2_X1 U13430 ( .A1(n13424), .A2(n13425), .ZN(n13278) );
  AND2_X1 U13431 ( .A1(n13275), .A2(n13274), .ZN(n13425) );
  AND2_X1 U13432 ( .A1(n13272), .A2(n13426), .ZN(n13424) );
  OR2_X1 U13433 ( .A1(n13274), .A2(n13275), .ZN(n13426) );
  OR2_X1 U13434 ( .A1(n8131), .A2(n7716), .ZN(n13275) );
  OR2_X1 U13435 ( .A1(n13427), .A2(n13428), .ZN(n13274) );
  AND2_X1 U13436 ( .A1(n13268), .A2(n13271), .ZN(n13428) );
  AND2_X1 U13437 ( .A1(n13429), .A2(n13270), .ZN(n13427) );
  OR2_X1 U13438 ( .A1(n13430), .A2(n13431), .ZN(n13270) );
  AND2_X1 U13439 ( .A1(n13264), .A2(n13267), .ZN(n13431) );
  AND2_X1 U13440 ( .A1(n13432), .A2(n13266), .ZN(n13430) );
  OR2_X1 U13441 ( .A1(n13433), .A2(n13434), .ZN(n13266) );
  AND2_X1 U13442 ( .A1(n13260), .A2(n13263), .ZN(n13434) );
  AND2_X1 U13443 ( .A1(n13435), .A2(n13262), .ZN(n13433) );
  OR2_X1 U13444 ( .A1(n13436), .A2(n13437), .ZN(n13262) );
  AND2_X1 U13445 ( .A1(n13256), .A2(n13259), .ZN(n13437) );
  AND2_X1 U13446 ( .A1(n13438), .A2(n13258), .ZN(n13436) );
  OR2_X1 U13447 ( .A1(n13439), .A2(n13440), .ZN(n13258) );
  AND2_X1 U13448 ( .A1(n13252), .A2(n13255), .ZN(n13440) );
  AND2_X1 U13449 ( .A1(n13254), .A2(n13441), .ZN(n13439) );
  OR2_X1 U13450 ( .A1(n13255), .A2(n13252), .ZN(n13441) );
  OR2_X1 U13451 ( .A1(n8102), .A2(n7716), .ZN(n13252) );
  OR3_X1 U13452 ( .A1(n8349), .A2(n7716), .A3(n7674), .ZN(n13255) );
  INV_X1 U13453 ( .A(n13442), .ZN(n13254) );
  OR2_X1 U13454 ( .A1(n13443), .A2(n13444), .ZN(n13442) );
  AND2_X1 U13455 ( .A1(b_5_), .A2(n13445), .ZN(n13444) );
  OR2_X1 U13456 ( .A1(n13446), .A2(n7314), .ZN(n13445) );
  AND2_X1 U13457 ( .A1(a_30_), .A2(n7648), .ZN(n13446) );
  AND2_X1 U13458 ( .A1(b_4_), .A2(n13447), .ZN(n13443) );
  OR2_X1 U13459 ( .A1(n13448), .A2(n7318), .ZN(n13447) );
  AND2_X1 U13460 ( .A1(a_31_), .A2(n7674), .ZN(n13448) );
  OR2_X1 U13461 ( .A1(n13259), .A2(n13256), .ZN(n13438) );
  XNOR2_X1 U13462 ( .A(n13449), .B(n13450), .ZN(n13256) );
  XNOR2_X1 U13463 ( .A(n13451), .B(n13452), .ZN(n13450) );
  OR2_X1 U13464 ( .A1(n8111), .A2(n7716), .ZN(n13259) );
  OR2_X1 U13465 ( .A1(n13263), .A2(n13260), .ZN(n13435) );
  XOR2_X1 U13466 ( .A(n13453), .B(n13454), .Z(n13260) );
  XOR2_X1 U13467 ( .A(n13455), .B(n13456), .Z(n13454) );
  OR2_X1 U13468 ( .A1(n8116), .A2(n7716), .ZN(n13263) );
  OR2_X1 U13469 ( .A1(n13267), .A2(n13264), .ZN(n13432) );
  XOR2_X1 U13470 ( .A(n13457), .B(n13458), .Z(n13264) );
  XOR2_X1 U13471 ( .A(n13459), .B(n13460), .Z(n13458) );
  OR2_X1 U13472 ( .A1(n8121), .A2(n7716), .ZN(n13267) );
  OR2_X1 U13473 ( .A1(n13271), .A2(n13268), .ZN(n13429) );
  XOR2_X1 U13474 ( .A(n13461), .B(n13462), .Z(n13268) );
  XOR2_X1 U13475 ( .A(n13463), .B(n13464), .Z(n13462) );
  OR2_X1 U13476 ( .A1(n8126), .A2(n7716), .ZN(n13271) );
  XOR2_X1 U13477 ( .A(n13465), .B(n13466), .Z(n13272) );
  XOR2_X1 U13478 ( .A(n13467), .B(n13468), .Z(n13466) );
  OR2_X1 U13479 ( .A1(n13279), .A2(n13276), .ZN(n13423) );
  XOR2_X1 U13480 ( .A(n13469), .B(n13470), .Z(n13276) );
  XOR2_X1 U13481 ( .A(n13471), .B(n13472), .Z(n13470) );
  OR2_X1 U13482 ( .A1(n8136), .A2(n7716), .ZN(n13279) );
  XOR2_X1 U13483 ( .A(n13473), .B(n13474), .Z(n13280) );
  XOR2_X1 U13484 ( .A(n13475), .B(n13476), .Z(n13474) );
  XOR2_X1 U13485 ( .A(n13477), .B(n13478), .Z(n13284) );
  XOR2_X1 U13486 ( .A(n13479), .B(n13480), .Z(n13478) );
  XOR2_X1 U13487 ( .A(n13481), .B(n13482), .Z(n13288) );
  XOR2_X1 U13488 ( .A(n13483), .B(n13484), .Z(n13482) );
  XOR2_X1 U13489 ( .A(n13485), .B(n13486), .Z(n13292) );
  XOR2_X1 U13490 ( .A(n13487), .B(n13488), .Z(n13486) );
  XOR2_X1 U13491 ( .A(n13489), .B(n13490), .Z(n13296) );
  XOR2_X1 U13492 ( .A(n13491), .B(n13492), .Z(n13490) );
  XOR2_X1 U13493 ( .A(n13493), .B(n13494), .Z(n13300) );
  XOR2_X1 U13494 ( .A(n13495), .B(n13496), .Z(n13494) );
  XOR2_X1 U13495 ( .A(n13497), .B(n13498), .Z(n13304) );
  XOR2_X1 U13496 ( .A(n13499), .B(n13500), .Z(n13498) );
  XOR2_X1 U13497 ( .A(n13501), .B(n13502), .Z(n13308) );
  XOR2_X1 U13498 ( .A(n13503), .B(n13504), .Z(n13502) );
  XOR2_X1 U13499 ( .A(n13505), .B(n13506), .Z(n13312) );
  XOR2_X1 U13500 ( .A(n13507), .B(n13508), .Z(n13506) );
  XOR2_X1 U13501 ( .A(n13509), .B(n13510), .Z(n13316) );
  XOR2_X1 U13502 ( .A(n13511), .B(n13512), .Z(n13510) );
  XOR2_X1 U13503 ( .A(n13513), .B(n13514), .Z(n13320) );
  XOR2_X1 U13504 ( .A(n13515), .B(n13516), .Z(n13514) );
  XOR2_X1 U13505 ( .A(n13517), .B(n13518), .Z(n13324) );
  XOR2_X1 U13506 ( .A(n13519), .B(n13520), .Z(n13518) );
  XOR2_X1 U13507 ( .A(n13521), .B(n13522), .Z(n13328) );
  XOR2_X1 U13508 ( .A(n13523), .B(n13524), .Z(n13522) );
  XOR2_X1 U13509 ( .A(n13525), .B(n13526), .Z(n13332) );
  XOR2_X1 U13510 ( .A(n13527), .B(n13528), .Z(n13526) );
  XOR2_X1 U13511 ( .A(n13529), .B(n13530), .Z(n13336) );
  XOR2_X1 U13512 ( .A(n13531), .B(n13532), .Z(n13530) );
  XOR2_X1 U13513 ( .A(n13533), .B(n13534), .Z(n13340) );
  XOR2_X1 U13514 ( .A(n13535), .B(n13536), .Z(n13534) );
  XOR2_X1 U13515 ( .A(n13537), .B(n13538), .Z(n13345) );
  XOR2_X1 U13516 ( .A(n13539), .B(n13540), .Z(n13538) );
  XOR2_X1 U13517 ( .A(n13541), .B(n13542), .Z(n13348) );
  XOR2_X1 U13518 ( .A(n13543), .B(n13544), .Z(n13542) );
  XNOR2_X1 U13519 ( .A(n13545), .B(n13546), .ZN(n13352) );
  XNOR2_X1 U13520 ( .A(n13547), .B(n13548), .ZN(n13545) );
  XOR2_X1 U13521 ( .A(n13549), .B(n13550), .Z(n13356) );
  XOR2_X1 U13522 ( .A(n13551), .B(n13552), .Z(n13550) );
  XOR2_X1 U13523 ( .A(n7774), .B(n13553), .Z(n7767) );
  XOR2_X1 U13524 ( .A(n7773), .B(n7772), .Z(n13553) );
  OR2_X1 U13525 ( .A1(n7674), .A2(n7777), .ZN(n7772) );
  OR2_X1 U13526 ( .A1(n13554), .A2(n13555), .ZN(n7773) );
  AND2_X1 U13527 ( .A1(n13552), .A2(n13551), .ZN(n13555) );
  AND2_X1 U13528 ( .A1(n13549), .A2(n13556), .ZN(n13554) );
  OR2_X1 U13529 ( .A1(n13551), .A2(n13552), .ZN(n13556) );
  OR2_X1 U13530 ( .A1(n7674), .A2(n7785), .ZN(n13552) );
  OR2_X1 U13531 ( .A1(n13557), .A2(n13558), .ZN(n13551) );
  AND2_X1 U13532 ( .A1(n13546), .A2(n13548), .ZN(n13558) );
  AND2_X1 U13533 ( .A1(n13559), .A2(n13547), .ZN(n13557) );
  OR2_X1 U13534 ( .A1(n13546), .A2(n13548), .ZN(n13559) );
  OR2_X1 U13535 ( .A1(n13560), .A2(n13561), .ZN(n13548) );
  AND2_X1 U13536 ( .A1(n13544), .A2(n13543), .ZN(n13561) );
  AND2_X1 U13537 ( .A1(n13541), .A2(n13562), .ZN(n13560) );
  OR2_X1 U13538 ( .A1(n13543), .A2(n13544), .ZN(n13562) );
  OR2_X1 U13539 ( .A1(n7674), .A2(n8221), .ZN(n13544) );
  OR2_X1 U13540 ( .A1(n13563), .A2(n13564), .ZN(n13543) );
  AND2_X1 U13541 ( .A1(n13540), .A2(n13539), .ZN(n13564) );
  AND2_X1 U13542 ( .A1(n13537), .A2(n13565), .ZN(n13563) );
  OR2_X1 U13543 ( .A1(n13539), .A2(n13540), .ZN(n13565) );
  OR2_X1 U13544 ( .A1(n7674), .A2(n8216), .ZN(n13540) );
  OR2_X1 U13545 ( .A1(n13566), .A2(n13567), .ZN(n13539) );
  AND2_X1 U13546 ( .A1(n13536), .A2(n13535), .ZN(n13567) );
  AND2_X1 U13547 ( .A1(n13533), .A2(n13568), .ZN(n13566) );
  OR2_X1 U13548 ( .A1(n13535), .A2(n13536), .ZN(n13568) );
  OR2_X1 U13549 ( .A1(n7674), .A2(n8211), .ZN(n13536) );
  OR2_X1 U13550 ( .A1(n13569), .A2(n13570), .ZN(n13535) );
  AND2_X1 U13551 ( .A1(n13532), .A2(n13531), .ZN(n13570) );
  AND2_X1 U13552 ( .A1(n13529), .A2(n13571), .ZN(n13569) );
  OR2_X1 U13553 ( .A1(n13531), .A2(n13532), .ZN(n13571) );
  OR2_X1 U13554 ( .A1(n7674), .A2(n8206), .ZN(n13532) );
  OR2_X1 U13555 ( .A1(n13572), .A2(n13573), .ZN(n13531) );
  AND2_X1 U13556 ( .A1(n13528), .A2(n13527), .ZN(n13573) );
  AND2_X1 U13557 ( .A1(n13525), .A2(n13574), .ZN(n13572) );
  OR2_X1 U13558 ( .A1(n13527), .A2(n13528), .ZN(n13574) );
  OR2_X1 U13559 ( .A1(n7674), .A2(n8201), .ZN(n13528) );
  OR2_X1 U13560 ( .A1(n13575), .A2(n13576), .ZN(n13527) );
  AND2_X1 U13561 ( .A1(n13524), .A2(n13523), .ZN(n13576) );
  AND2_X1 U13562 ( .A1(n13521), .A2(n13577), .ZN(n13575) );
  OR2_X1 U13563 ( .A1(n13523), .A2(n13524), .ZN(n13577) );
  OR2_X1 U13564 ( .A1(n7674), .A2(n8196), .ZN(n13524) );
  OR2_X1 U13565 ( .A1(n13578), .A2(n13579), .ZN(n13523) );
  AND2_X1 U13566 ( .A1(n13520), .A2(n13519), .ZN(n13579) );
  AND2_X1 U13567 ( .A1(n13517), .A2(n13580), .ZN(n13578) );
  OR2_X1 U13568 ( .A1(n13519), .A2(n13520), .ZN(n13580) );
  OR2_X1 U13569 ( .A1(n7674), .A2(n8191), .ZN(n13520) );
  OR2_X1 U13570 ( .A1(n13581), .A2(n13582), .ZN(n13519) );
  AND2_X1 U13571 ( .A1(n13516), .A2(n13515), .ZN(n13582) );
  AND2_X1 U13572 ( .A1(n13513), .A2(n13583), .ZN(n13581) );
  OR2_X1 U13573 ( .A1(n13515), .A2(n13516), .ZN(n13583) );
  OR2_X1 U13574 ( .A1(n7674), .A2(n8186), .ZN(n13516) );
  OR2_X1 U13575 ( .A1(n13584), .A2(n13585), .ZN(n13515) );
  AND2_X1 U13576 ( .A1(n13512), .A2(n13511), .ZN(n13585) );
  AND2_X1 U13577 ( .A1(n13509), .A2(n13586), .ZN(n13584) );
  OR2_X1 U13578 ( .A1(n13511), .A2(n13512), .ZN(n13586) );
  OR2_X1 U13579 ( .A1(n7674), .A2(n8181), .ZN(n13512) );
  OR2_X1 U13580 ( .A1(n13587), .A2(n13588), .ZN(n13511) );
  AND2_X1 U13581 ( .A1(n13508), .A2(n13507), .ZN(n13588) );
  AND2_X1 U13582 ( .A1(n13505), .A2(n13589), .ZN(n13587) );
  OR2_X1 U13583 ( .A1(n13507), .A2(n13508), .ZN(n13589) );
  OR2_X1 U13584 ( .A1(n7674), .A2(n8176), .ZN(n13508) );
  OR2_X1 U13585 ( .A1(n13590), .A2(n13591), .ZN(n13507) );
  AND2_X1 U13586 ( .A1(n13504), .A2(n13503), .ZN(n13591) );
  AND2_X1 U13587 ( .A1(n13501), .A2(n13592), .ZN(n13590) );
  OR2_X1 U13588 ( .A1(n13503), .A2(n13504), .ZN(n13592) );
  OR2_X1 U13589 ( .A1(n7674), .A2(n8171), .ZN(n13504) );
  OR2_X1 U13590 ( .A1(n13593), .A2(n13594), .ZN(n13503) );
  AND2_X1 U13591 ( .A1(n13500), .A2(n13499), .ZN(n13594) );
  AND2_X1 U13592 ( .A1(n13497), .A2(n13595), .ZN(n13593) );
  OR2_X1 U13593 ( .A1(n13499), .A2(n13500), .ZN(n13595) );
  OR2_X1 U13594 ( .A1(n8166), .A2(n7674), .ZN(n13500) );
  OR2_X1 U13595 ( .A1(n13596), .A2(n13597), .ZN(n13499) );
  AND2_X1 U13596 ( .A1(n13496), .A2(n13495), .ZN(n13597) );
  AND2_X1 U13597 ( .A1(n13493), .A2(n13598), .ZN(n13596) );
  OR2_X1 U13598 ( .A1(n13495), .A2(n13496), .ZN(n13598) );
  OR2_X1 U13599 ( .A1(n7674), .A2(n8161), .ZN(n13496) );
  OR2_X1 U13600 ( .A1(n13599), .A2(n13600), .ZN(n13495) );
  AND2_X1 U13601 ( .A1(n13492), .A2(n13491), .ZN(n13600) );
  AND2_X1 U13602 ( .A1(n13489), .A2(n13601), .ZN(n13599) );
  OR2_X1 U13603 ( .A1(n13491), .A2(n13492), .ZN(n13601) );
  OR2_X1 U13604 ( .A1(n8156), .A2(n7674), .ZN(n13492) );
  OR2_X1 U13605 ( .A1(n13602), .A2(n13603), .ZN(n13491) );
  AND2_X1 U13606 ( .A1(n13488), .A2(n13487), .ZN(n13603) );
  AND2_X1 U13607 ( .A1(n13485), .A2(n13604), .ZN(n13602) );
  OR2_X1 U13608 ( .A1(n13487), .A2(n13488), .ZN(n13604) );
  OR2_X1 U13609 ( .A1(n8151), .A2(n7674), .ZN(n13488) );
  OR2_X1 U13610 ( .A1(n13605), .A2(n13606), .ZN(n13487) );
  AND2_X1 U13611 ( .A1(n13484), .A2(n13483), .ZN(n13606) );
  AND2_X1 U13612 ( .A1(n13481), .A2(n13607), .ZN(n13605) );
  OR2_X1 U13613 ( .A1(n13483), .A2(n13484), .ZN(n13607) );
  OR2_X1 U13614 ( .A1(n8146), .A2(n7674), .ZN(n13484) );
  OR2_X1 U13615 ( .A1(n13608), .A2(n13609), .ZN(n13483) );
  AND2_X1 U13616 ( .A1(n13480), .A2(n13479), .ZN(n13609) );
  AND2_X1 U13617 ( .A1(n13477), .A2(n13610), .ZN(n13608) );
  OR2_X1 U13618 ( .A1(n13479), .A2(n13480), .ZN(n13610) );
  OR2_X1 U13619 ( .A1(n8141), .A2(n7674), .ZN(n13480) );
  OR2_X1 U13620 ( .A1(n13611), .A2(n13612), .ZN(n13479) );
  AND2_X1 U13621 ( .A1(n13476), .A2(n13475), .ZN(n13612) );
  AND2_X1 U13622 ( .A1(n13473), .A2(n13613), .ZN(n13611) );
  OR2_X1 U13623 ( .A1(n13475), .A2(n13476), .ZN(n13613) );
  OR2_X1 U13624 ( .A1(n8136), .A2(n7674), .ZN(n13476) );
  OR2_X1 U13625 ( .A1(n13614), .A2(n13615), .ZN(n13475) );
  AND2_X1 U13626 ( .A1(n13469), .A2(n13472), .ZN(n13615) );
  AND2_X1 U13627 ( .A1(n13616), .A2(n13471), .ZN(n13614) );
  OR2_X1 U13628 ( .A1(n13617), .A2(n13618), .ZN(n13471) );
  AND2_X1 U13629 ( .A1(n13468), .A2(n13467), .ZN(n13618) );
  AND2_X1 U13630 ( .A1(n13465), .A2(n13619), .ZN(n13617) );
  OR2_X1 U13631 ( .A1(n13467), .A2(n13468), .ZN(n13619) );
  OR2_X1 U13632 ( .A1(n8126), .A2(n7674), .ZN(n13468) );
  OR2_X1 U13633 ( .A1(n13620), .A2(n13621), .ZN(n13467) );
  AND2_X1 U13634 ( .A1(n13461), .A2(n13464), .ZN(n13621) );
  AND2_X1 U13635 ( .A1(n13622), .A2(n13463), .ZN(n13620) );
  OR2_X1 U13636 ( .A1(n13623), .A2(n13624), .ZN(n13463) );
  AND2_X1 U13637 ( .A1(n13457), .A2(n13460), .ZN(n13624) );
  AND2_X1 U13638 ( .A1(n13625), .A2(n13459), .ZN(n13623) );
  OR2_X1 U13639 ( .A1(n13626), .A2(n13627), .ZN(n13459) );
  AND2_X1 U13640 ( .A1(n13453), .A2(n13456), .ZN(n13627) );
  AND2_X1 U13641 ( .A1(n13628), .A2(n13455), .ZN(n13626) );
  OR2_X1 U13642 ( .A1(n13629), .A2(n13630), .ZN(n13455) );
  AND2_X1 U13643 ( .A1(n13449), .A2(n13452), .ZN(n13630) );
  AND2_X1 U13644 ( .A1(n13451), .A2(n13631), .ZN(n13629) );
  OR2_X1 U13645 ( .A1(n13452), .A2(n13449), .ZN(n13631) );
  OR2_X1 U13646 ( .A1(n8102), .A2(n7674), .ZN(n13449) );
  OR3_X1 U13647 ( .A1(n8349), .A2(n7674), .A3(n7648), .ZN(n13452) );
  INV_X1 U13648 ( .A(n13632), .ZN(n13451) );
  OR2_X1 U13649 ( .A1(n13633), .A2(n13634), .ZN(n13632) );
  AND2_X1 U13650 ( .A1(b_4_), .A2(n13635), .ZN(n13634) );
  OR2_X1 U13651 ( .A1(n13636), .A2(n7314), .ZN(n13635) );
  AND2_X1 U13652 ( .A1(a_30_), .A2(n7620), .ZN(n13636) );
  AND2_X1 U13653 ( .A1(b_3_), .A2(n13637), .ZN(n13633) );
  OR2_X1 U13654 ( .A1(n13638), .A2(n7318), .ZN(n13637) );
  AND2_X1 U13655 ( .A1(a_31_), .A2(n7648), .ZN(n13638) );
  OR2_X1 U13656 ( .A1(n13456), .A2(n13453), .ZN(n13628) );
  XNOR2_X1 U13657 ( .A(n13639), .B(n13640), .ZN(n13453) );
  XNOR2_X1 U13658 ( .A(n13641), .B(n13642), .ZN(n13640) );
  OR2_X1 U13659 ( .A1(n8111), .A2(n7674), .ZN(n13456) );
  OR2_X1 U13660 ( .A1(n13460), .A2(n13457), .ZN(n13625) );
  XOR2_X1 U13661 ( .A(n13643), .B(n13644), .Z(n13457) );
  XOR2_X1 U13662 ( .A(n13645), .B(n13646), .Z(n13644) );
  OR2_X1 U13663 ( .A1(n8116), .A2(n7674), .ZN(n13460) );
  OR2_X1 U13664 ( .A1(n13464), .A2(n13461), .ZN(n13622) );
  XOR2_X1 U13665 ( .A(n13647), .B(n13648), .Z(n13461) );
  XOR2_X1 U13666 ( .A(n13649), .B(n13650), .Z(n13648) );
  OR2_X1 U13667 ( .A1(n8121), .A2(n7674), .ZN(n13464) );
  XOR2_X1 U13668 ( .A(n13651), .B(n13652), .Z(n13465) );
  XOR2_X1 U13669 ( .A(n13653), .B(n13654), .Z(n13652) );
  OR2_X1 U13670 ( .A1(n13472), .A2(n13469), .ZN(n13616) );
  XOR2_X1 U13671 ( .A(n13655), .B(n13656), .Z(n13469) );
  XOR2_X1 U13672 ( .A(n13657), .B(n13658), .Z(n13656) );
  OR2_X1 U13673 ( .A1(n8131), .A2(n7674), .ZN(n13472) );
  XOR2_X1 U13674 ( .A(n13659), .B(n13660), .Z(n13473) );
  XOR2_X1 U13675 ( .A(n13661), .B(n13662), .Z(n13660) );
  XOR2_X1 U13676 ( .A(n13663), .B(n13664), .Z(n13477) );
  XOR2_X1 U13677 ( .A(n13665), .B(n13666), .Z(n13664) );
  XOR2_X1 U13678 ( .A(n13667), .B(n13668), .Z(n13481) );
  XOR2_X1 U13679 ( .A(n13669), .B(n13670), .Z(n13668) );
  XOR2_X1 U13680 ( .A(n13671), .B(n13672), .Z(n13485) );
  XOR2_X1 U13681 ( .A(n13673), .B(n13674), .Z(n13672) );
  XOR2_X1 U13682 ( .A(n13675), .B(n13676), .Z(n13489) );
  XOR2_X1 U13683 ( .A(n13677), .B(n13678), .Z(n13676) );
  XOR2_X1 U13684 ( .A(n13679), .B(n13680), .Z(n13493) );
  XOR2_X1 U13685 ( .A(n13681), .B(n13682), .Z(n13680) );
  XOR2_X1 U13686 ( .A(n13683), .B(n13684), .Z(n13497) );
  XOR2_X1 U13687 ( .A(n13685), .B(n13686), .Z(n13684) );
  XOR2_X1 U13688 ( .A(n13687), .B(n13688), .Z(n13501) );
  XOR2_X1 U13689 ( .A(n13689), .B(n13690), .Z(n13688) );
  XOR2_X1 U13690 ( .A(n13691), .B(n13692), .Z(n13505) );
  XOR2_X1 U13691 ( .A(n13693), .B(n13694), .Z(n13692) );
  XOR2_X1 U13692 ( .A(n13695), .B(n13696), .Z(n13509) );
  XOR2_X1 U13693 ( .A(n13697), .B(n13698), .Z(n13696) );
  XOR2_X1 U13694 ( .A(n13699), .B(n13700), .Z(n13513) );
  XOR2_X1 U13695 ( .A(n13701), .B(n13702), .Z(n13700) );
  XOR2_X1 U13696 ( .A(n13703), .B(n13704), .Z(n13517) );
  XOR2_X1 U13697 ( .A(n13705), .B(n13706), .Z(n13704) );
  XOR2_X1 U13698 ( .A(n13707), .B(n13708), .Z(n13521) );
  XOR2_X1 U13699 ( .A(n13709), .B(n13710), .Z(n13708) );
  XOR2_X1 U13700 ( .A(n13711), .B(n13712), .Z(n13525) );
  XOR2_X1 U13701 ( .A(n13713), .B(n13714), .Z(n13712) );
  XOR2_X1 U13702 ( .A(n13715), .B(n13716), .Z(n13529) );
  XOR2_X1 U13703 ( .A(n13717), .B(n13718), .Z(n13716) );
  XOR2_X1 U13704 ( .A(n13719), .B(n13720), .Z(n13533) );
  XOR2_X1 U13705 ( .A(n13721), .B(n13722), .Z(n13720) );
  XOR2_X1 U13706 ( .A(n13723), .B(n13724), .Z(n13537) );
  XOR2_X1 U13707 ( .A(n13725), .B(n13726), .Z(n13724) );
  XOR2_X1 U13708 ( .A(n13727), .B(n13728), .Z(n13541) );
  XOR2_X1 U13709 ( .A(n13729), .B(n13730), .Z(n13728) );
  XOR2_X1 U13710 ( .A(n13731), .B(n13732), .Z(n13546) );
  XOR2_X1 U13711 ( .A(n13733), .B(n13734), .Z(n13732) );
  XOR2_X1 U13712 ( .A(n13735), .B(n13736), .Z(n13549) );
  XOR2_X1 U13713 ( .A(n13737), .B(n13738), .Z(n13736) );
  XNOR2_X1 U13714 ( .A(n13739), .B(n7780), .ZN(n7774) );
  XOR2_X1 U13715 ( .A(n7790), .B(n13740), .Z(n7780) );
  XOR2_X1 U13716 ( .A(n7789), .B(n7788), .Z(n13740) );
  OR2_X1 U13717 ( .A1(n7620), .A2(n8226), .ZN(n7788) );
  OR2_X1 U13718 ( .A1(n13741), .A2(n13742), .ZN(n7789) );
  AND2_X1 U13719 ( .A1(n13743), .A2(n13744), .ZN(n13742) );
  AND2_X1 U13720 ( .A1(n13745), .A2(n13746), .ZN(n13741) );
  OR2_X1 U13721 ( .A1(n13744), .A2(n13743), .ZN(n13746) );
  XOR2_X1 U13722 ( .A(n13747), .B(n13748), .Z(n7790) );
  XOR2_X1 U13723 ( .A(n13749), .B(n13750), .Z(n13748) );
  XNOR2_X1 U13724 ( .A(n7783), .B(n7781), .ZN(n13739) );
  OR2_X1 U13725 ( .A1(n13751), .A2(n13752), .ZN(n7781) );
  AND2_X1 U13726 ( .A1(n13738), .A2(n13737), .ZN(n13752) );
  AND2_X1 U13727 ( .A1(n13735), .A2(n13753), .ZN(n13751) );
  OR2_X1 U13728 ( .A1(n13737), .A2(n13738), .ZN(n13753) );
  OR2_X1 U13729 ( .A1(n7648), .A2(n8226), .ZN(n13738) );
  OR2_X1 U13730 ( .A1(n13754), .A2(n13755), .ZN(n13737) );
  AND2_X1 U13731 ( .A1(n13734), .A2(n13733), .ZN(n13755) );
  AND2_X1 U13732 ( .A1(n13731), .A2(n13756), .ZN(n13754) );
  OR2_X1 U13733 ( .A1(n13733), .A2(n13734), .ZN(n13756) );
  OR2_X1 U13734 ( .A1(n7648), .A2(n8221), .ZN(n13734) );
  OR2_X1 U13735 ( .A1(n13757), .A2(n13758), .ZN(n13733) );
  AND2_X1 U13736 ( .A1(n13730), .A2(n13729), .ZN(n13758) );
  AND2_X1 U13737 ( .A1(n13727), .A2(n13759), .ZN(n13757) );
  OR2_X1 U13738 ( .A1(n13729), .A2(n13730), .ZN(n13759) );
  OR2_X1 U13739 ( .A1(n7648), .A2(n8216), .ZN(n13730) );
  OR2_X1 U13740 ( .A1(n13760), .A2(n13761), .ZN(n13729) );
  AND2_X1 U13741 ( .A1(n13726), .A2(n13725), .ZN(n13761) );
  AND2_X1 U13742 ( .A1(n13723), .A2(n13762), .ZN(n13760) );
  OR2_X1 U13743 ( .A1(n13725), .A2(n13726), .ZN(n13762) );
  OR2_X1 U13744 ( .A1(n7648), .A2(n8211), .ZN(n13726) );
  OR2_X1 U13745 ( .A1(n13763), .A2(n13764), .ZN(n13725) );
  AND2_X1 U13746 ( .A1(n13722), .A2(n13721), .ZN(n13764) );
  AND2_X1 U13747 ( .A1(n13719), .A2(n13765), .ZN(n13763) );
  OR2_X1 U13748 ( .A1(n13721), .A2(n13722), .ZN(n13765) );
  OR2_X1 U13749 ( .A1(n7648), .A2(n8206), .ZN(n13722) );
  OR2_X1 U13750 ( .A1(n13766), .A2(n13767), .ZN(n13721) );
  AND2_X1 U13751 ( .A1(n13718), .A2(n13717), .ZN(n13767) );
  AND2_X1 U13752 ( .A1(n13715), .A2(n13768), .ZN(n13766) );
  OR2_X1 U13753 ( .A1(n13717), .A2(n13718), .ZN(n13768) );
  OR2_X1 U13754 ( .A1(n7648), .A2(n8201), .ZN(n13718) );
  OR2_X1 U13755 ( .A1(n13769), .A2(n13770), .ZN(n13717) );
  AND2_X1 U13756 ( .A1(n13714), .A2(n13713), .ZN(n13770) );
  AND2_X1 U13757 ( .A1(n13711), .A2(n13771), .ZN(n13769) );
  OR2_X1 U13758 ( .A1(n13713), .A2(n13714), .ZN(n13771) );
  OR2_X1 U13759 ( .A1(n7648), .A2(n8196), .ZN(n13714) );
  OR2_X1 U13760 ( .A1(n13772), .A2(n13773), .ZN(n13713) );
  AND2_X1 U13761 ( .A1(n13710), .A2(n13709), .ZN(n13773) );
  AND2_X1 U13762 ( .A1(n13707), .A2(n13774), .ZN(n13772) );
  OR2_X1 U13763 ( .A1(n13709), .A2(n13710), .ZN(n13774) );
  OR2_X1 U13764 ( .A1(n7648), .A2(n8191), .ZN(n13710) );
  OR2_X1 U13765 ( .A1(n13775), .A2(n13776), .ZN(n13709) );
  AND2_X1 U13766 ( .A1(n13706), .A2(n13705), .ZN(n13776) );
  AND2_X1 U13767 ( .A1(n13703), .A2(n13777), .ZN(n13775) );
  OR2_X1 U13768 ( .A1(n13705), .A2(n13706), .ZN(n13777) );
  OR2_X1 U13769 ( .A1(n7648), .A2(n8186), .ZN(n13706) );
  OR2_X1 U13770 ( .A1(n13778), .A2(n13779), .ZN(n13705) );
  AND2_X1 U13771 ( .A1(n13702), .A2(n13701), .ZN(n13779) );
  AND2_X1 U13772 ( .A1(n13699), .A2(n13780), .ZN(n13778) );
  OR2_X1 U13773 ( .A1(n13701), .A2(n13702), .ZN(n13780) );
  OR2_X1 U13774 ( .A1(n7648), .A2(n8181), .ZN(n13702) );
  OR2_X1 U13775 ( .A1(n13781), .A2(n13782), .ZN(n13701) );
  AND2_X1 U13776 ( .A1(n13698), .A2(n13697), .ZN(n13782) );
  AND2_X1 U13777 ( .A1(n13695), .A2(n13783), .ZN(n13781) );
  OR2_X1 U13778 ( .A1(n13697), .A2(n13698), .ZN(n13783) );
  OR2_X1 U13779 ( .A1(n7648), .A2(n8176), .ZN(n13698) );
  OR2_X1 U13780 ( .A1(n13784), .A2(n13785), .ZN(n13697) );
  AND2_X1 U13781 ( .A1(n13694), .A2(n13693), .ZN(n13785) );
  AND2_X1 U13782 ( .A1(n13691), .A2(n13786), .ZN(n13784) );
  OR2_X1 U13783 ( .A1(n13693), .A2(n13694), .ZN(n13786) );
  OR2_X1 U13784 ( .A1(n7648), .A2(n8171), .ZN(n13694) );
  OR2_X1 U13785 ( .A1(n13787), .A2(n13788), .ZN(n13693) );
  AND2_X1 U13786 ( .A1(n13690), .A2(n13689), .ZN(n13788) );
  AND2_X1 U13787 ( .A1(n13687), .A2(n13789), .ZN(n13787) );
  OR2_X1 U13788 ( .A1(n13689), .A2(n13690), .ZN(n13789) );
  OR2_X1 U13789 ( .A1(n8166), .A2(n7648), .ZN(n13690) );
  OR2_X1 U13790 ( .A1(n13790), .A2(n13791), .ZN(n13689) );
  AND2_X1 U13791 ( .A1(n13686), .A2(n13685), .ZN(n13791) );
  AND2_X1 U13792 ( .A1(n13683), .A2(n13792), .ZN(n13790) );
  OR2_X1 U13793 ( .A1(n13685), .A2(n13686), .ZN(n13792) );
  OR2_X1 U13794 ( .A1(n8161), .A2(n7648), .ZN(n13686) );
  OR2_X1 U13795 ( .A1(n13793), .A2(n13794), .ZN(n13685) );
  AND2_X1 U13796 ( .A1(n13682), .A2(n13681), .ZN(n13794) );
  AND2_X1 U13797 ( .A1(n13679), .A2(n13795), .ZN(n13793) );
  OR2_X1 U13798 ( .A1(n13681), .A2(n13682), .ZN(n13795) );
  OR2_X1 U13799 ( .A1(n8156), .A2(n7648), .ZN(n13682) );
  OR2_X1 U13800 ( .A1(n13796), .A2(n13797), .ZN(n13681) );
  AND2_X1 U13801 ( .A1(n13678), .A2(n13677), .ZN(n13797) );
  AND2_X1 U13802 ( .A1(n13675), .A2(n13798), .ZN(n13796) );
  OR2_X1 U13803 ( .A1(n13677), .A2(n13678), .ZN(n13798) );
  OR2_X1 U13804 ( .A1(n8151), .A2(n7648), .ZN(n13678) );
  OR2_X1 U13805 ( .A1(n13799), .A2(n13800), .ZN(n13677) );
  AND2_X1 U13806 ( .A1(n13674), .A2(n13673), .ZN(n13800) );
  AND2_X1 U13807 ( .A1(n13671), .A2(n13801), .ZN(n13799) );
  OR2_X1 U13808 ( .A1(n13673), .A2(n13674), .ZN(n13801) );
  OR2_X1 U13809 ( .A1(n8146), .A2(n7648), .ZN(n13674) );
  OR2_X1 U13810 ( .A1(n13802), .A2(n13803), .ZN(n13673) );
  AND2_X1 U13811 ( .A1(n13670), .A2(n13669), .ZN(n13803) );
  AND2_X1 U13812 ( .A1(n13667), .A2(n13804), .ZN(n13802) );
  OR2_X1 U13813 ( .A1(n13669), .A2(n13670), .ZN(n13804) );
  OR2_X1 U13814 ( .A1(n8141), .A2(n7648), .ZN(n13670) );
  OR2_X1 U13815 ( .A1(n13805), .A2(n13806), .ZN(n13669) );
  AND2_X1 U13816 ( .A1(n13666), .A2(n13665), .ZN(n13806) );
  AND2_X1 U13817 ( .A1(n13663), .A2(n13807), .ZN(n13805) );
  OR2_X1 U13818 ( .A1(n13665), .A2(n13666), .ZN(n13807) );
  OR2_X1 U13819 ( .A1(n8136), .A2(n7648), .ZN(n13666) );
  OR2_X1 U13820 ( .A1(n13808), .A2(n13809), .ZN(n13665) );
  AND2_X1 U13821 ( .A1(n13662), .A2(n13661), .ZN(n13809) );
  AND2_X1 U13822 ( .A1(n13659), .A2(n13810), .ZN(n13808) );
  OR2_X1 U13823 ( .A1(n13661), .A2(n13662), .ZN(n13810) );
  OR2_X1 U13824 ( .A1(n8131), .A2(n7648), .ZN(n13662) );
  OR2_X1 U13825 ( .A1(n13811), .A2(n13812), .ZN(n13661) );
  AND2_X1 U13826 ( .A1(n13655), .A2(n13658), .ZN(n13812) );
  AND2_X1 U13827 ( .A1(n13813), .A2(n13657), .ZN(n13811) );
  OR2_X1 U13828 ( .A1(n13814), .A2(n13815), .ZN(n13657) );
  AND2_X1 U13829 ( .A1(n13654), .A2(n13653), .ZN(n13815) );
  AND2_X1 U13830 ( .A1(n13651), .A2(n13816), .ZN(n13814) );
  OR2_X1 U13831 ( .A1(n13653), .A2(n13654), .ZN(n13816) );
  OR2_X1 U13832 ( .A1(n8121), .A2(n7648), .ZN(n13654) );
  OR2_X1 U13833 ( .A1(n13817), .A2(n13818), .ZN(n13653) );
  AND2_X1 U13834 ( .A1(n13647), .A2(n13650), .ZN(n13818) );
  AND2_X1 U13835 ( .A1(n13819), .A2(n13649), .ZN(n13817) );
  OR2_X1 U13836 ( .A1(n13820), .A2(n13821), .ZN(n13649) );
  AND2_X1 U13837 ( .A1(n13643), .A2(n13646), .ZN(n13821) );
  AND2_X1 U13838 ( .A1(n13822), .A2(n13645), .ZN(n13820) );
  OR2_X1 U13839 ( .A1(n13823), .A2(n13824), .ZN(n13645) );
  AND2_X1 U13840 ( .A1(n13639), .A2(n13642), .ZN(n13824) );
  AND2_X1 U13841 ( .A1(n13641), .A2(n13825), .ZN(n13823) );
  OR2_X1 U13842 ( .A1(n13642), .A2(n13639), .ZN(n13825) );
  OR2_X1 U13843 ( .A1(n8102), .A2(n7648), .ZN(n13639) );
  OR3_X1 U13844 ( .A1(n8349), .A2(n7648), .A3(n7620), .ZN(n13642) );
  INV_X1 U13845 ( .A(n13826), .ZN(n13641) );
  OR2_X1 U13846 ( .A1(n13827), .A2(n13828), .ZN(n13826) );
  AND2_X1 U13847 ( .A1(b_3_), .A2(n13829), .ZN(n13828) );
  OR2_X1 U13848 ( .A1(n13830), .A2(n7314), .ZN(n13829) );
  AND2_X1 U13849 ( .A1(a_30_), .A2(n13831), .ZN(n13830) );
  AND2_X1 U13850 ( .A1(b_2_), .A2(n13832), .ZN(n13827) );
  OR2_X1 U13851 ( .A1(n13833), .A2(n7318), .ZN(n13832) );
  AND2_X1 U13852 ( .A1(a_31_), .A2(n7620), .ZN(n13833) );
  OR2_X1 U13853 ( .A1(n13646), .A2(n13643), .ZN(n13822) );
  XNOR2_X1 U13854 ( .A(n13834), .B(n13835), .ZN(n13643) );
  XNOR2_X1 U13855 ( .A(n13836), .B(n13837), .ZN(n13835) );
  OR2_X1 U13856 ( .A1(n8111), .A2(n7648), .ZN(n13646) );
  OR2_X1 U13857 ( .A1(n13650), .A2(n13647), .ZN(n13819) );
  XOR2_X1 U13858 ( .A(n13838), .B(n13839), .Z(n13647) );
  XOR2_X1 U13859 ( .A(n13840), .B(n13841), .Z(n13839) );
  OR2_X1 U13860 ( .A1(n8116), .A2(n7648), .ZN(n13650) );
  XOR2_X1 U13861 ( .A(n13842), .B(n13843), .Z(n13651) );
  XOR2_X1 U13862 ( .A(n13844), .B(n13845), .Z(n13843) );
  OR2_X1 U13863 ( .A1(n13658), .A2(n13655), .ZN(n13813) );
  XOR2_X1 U13864 ( .A(n13846), .B(n13847), .Z(n13655) );
  XOR2_X1 U13865 ( .A(n13848), .B(n13849), .Z(n13847) );
  OR2_X1 U13866 ( .A1(n8126), .A2(n7648), .ZN(n13658) );
  XOR2_X1 U13867 ( .A(n13850), .B(n13851), .Z(n13659) );
  XOR2_X1 U13868 ( .A(n13852), .B(n13853), .Z(n13851) );
  XOR2_X1 U13869 ( .A(n13854), .B(n13855), .Z(n13663) );
  XOR2_X1 U13870 ( .A(n13856), .B(n13857), .Z(n13855) );
  XOR2_X1 U13871 ( .A(n13858), .B(n13859), .Z(n13667) );
  XOR2_X1 U13872 ( .A(n13860), .B(n13861), .Z(n13859) );
  XOR2_X1 U13873 ( .A(n13862), .B(n13863), .Z(n13671) );
  XOR2_X1 U13874 ( .A(n13864), .B(n13865), .Z(n13863) );
  XOR2_X1 U13875 ( .A(n13866), .B(n13867), .Z(n13675) );
  XOR2_X1 U13876 ( .A(n13868), .B(n13869), .Z(n13867) );
  XOR2_X1 U13877 ( .A(n13870), .B(n13871), .Z(n13679) );
  XOR2_X1 U13878 ( .A(n13872), .B(n13873), .Z(n13871) );
  XOR2_X1 U13879 ( .A(n13874), .B(n13875), .Z(n13683) );
  XOR2_X1 U13880 ( .A(n13876), .B(n13877), .Z(n13875) );
  XOR2_X1 U13881 ( .A(n13878), .B(n13879), .Z(n13687) );
  XOR2_X1 U13882 ( .A(n13880), .B(n13881), .Z(n13879) );
  XOR2_X1 U13883 ( .A(n13882), .B(n13883), .Z(n13691) );
  XOR2_X1 U13884 ( .A(n13884), .B(n13885), .Z(n13883) );
  XOR2_X1 U13885 ( .A(n13886), .B(n13887), .Z(n13695) );
  XOR2_X1 U13886 ( .A(n13888), .B(n13889), .Z(n13887) );
  XOR2_X1 U13887 ( .A(n13890), .B(n13891), .Z(n13699) );
  XOR2_X1 U13888 ( .A(n13892), .B(n13893), .Z(n13891) );
  XOR2_X1 U13889 ( .A(n13894), .B(n13895), .Z(n13703) );
  XOR2_X1 U13890 ( .A(n13896), .B(n13897), .Z(n13895) );
  XOR2_X1 U13891 ( .A(n13898), .B(n13899), .Z(n13707) );
  XOR2_X1 U13892 ( .A(n13900), .B(n13901), .Z(n13899) );
  XOR2_X1 U13893 ( .A(n13902), .B(n13903), .Z(n13711) );
  XOR2_X1 U13894 ( .A(n13904), .B(n13905), .Z(n13903) );
  XOR2_X1 U13895 ( .A(n13906), .B(n13907), .Z(n13715) );
  XOR2_X1 U13896 ( .A(n13908), .B(n13909), .Z(n13907) );
  XOR2_X1 U13897 ( .A(n13910), .B(n13911), .Z(n13719) );
  XOR2_X1 U13898 ( .A(n13912), .B(n13913), .Z(n13911) );
  XOR2_X1 U13899 ( .A(n13914), .B(n13915), .Z(n13723) );
  XOR2_X1 U13900 ( .A(n13916), .B(n13917), .Z(n13915) );
  XOR2_X1 U13901 ( .A(n13918), .B(n13919), .Z(n13727) );
  XOR2_X1 U13902 ( .A(n13920), .B(n13921), .Z(n13919) );
  XOR2_X1 U13903 ( .A(n13922), .B(n13923), .Z(n13731) );
  XOR2_X1 U13904 ( .A(n13924), .B(n13925), .Z(n13923) );
  XOR2_X1 U13905 ( .A(n13745), .B(n13926), .Z(n13735) );
  XOR2_X1 U13906 ( .A(n13744), .B(n13743), .Z(n13926) );
  OR2_X1 U13907 ( .A1(n7620), .A2(n8221), .ZN(n13743) );
  OR2_X1 U13908 ( .A1(n13927), .A2(n13928), .ZN(n13744) );
  AND2_X1 U13909 ( .A1(n13925), .A2(n13924), .ZN(n13928) );
  AND2_X1 U13910 ( .A1(n13922), .A2(n13929), .ZN(n13927) );
  OR2_X1 U13911 ( .A1(n13924), .A2(n13925), .ZN(n13929) );
  OR2_X1 U13912 ( .A1(n7620), .A2(n8216), .ZN(n13925) );
  OR2_X1 U13913 ( .A1(n13930), .A2(n13931), .ZN(n13924) );
  AND2_X1 U13914 ( .A1(n13921), .A2(n13920), .ZN(n13931) );
  AND2_X1 U13915 ( .A1(n13918), .A2(n13932), .ZN(n13930) );
  OR2_X1 U13916 ( .A1(n13920), .A2(n13921), .ZN(n13932) );
  OR2_X1 U13917 ( .A1(n7620), .A2(n8211), .ZN(n13921) );
  OR2_X1 U13918 ( .A1(n13933), .A2(n13934), .ZN(n13920) );
  AND2_X1 U13919 ( .A1(n13917), .A2(n13916), .ZN(n13934) );
  AND2_X1 U13920 ( .A1(n13914), .A2(n13935), .ZN(n13933) );
  OR2_X1 U13921 ( .A1(n13916), .A2(n13917), .ZN(n13935) );
  OR2_X1 U13922 ( .A1(n7620), .A2(n8206), .ZN(n13917) );
  OR2_X1 U13923 ( .A1(n13936), .A2(n13937), .ZN(n13916) );
  AND2_X1 U13924 ( .A1(n13913), .A2(n13912), .ZN(n13937) );
  AND2_X1 U13925 ( .A1(n13910), .A2(n13938), .ZN(n13936) );
  OR2_X1 U13926 ( .A1(n13912), .A2(n13913), .ZN(n13938) );
  OR2_X1 U13927 ( .A1(n7620), .A2(n8201), .ZN(n13913) );
  OR2_X1 U13928 ( .A1(n13939), .A2(n13940), .ZN(n13912) );
  AND2_X1 U13929 ( .A1(n13909), .A2(n13908), .ZN(n13940) );
  AND2_X1 U13930 ( .A1(n13906), .A2(n13941), .ZN(n13939) );
  OR2_X1 U13931 ( .A1(n13908), .A2(n13909), .ZN(n13941) );
  OR2_X1 U13932 ( .A1(n7620), .A2(n8196), .ZN(n13909) );
  OR2_X1 U13933 ( .A1(n13942), .A2(n13943), .ZN(n13908) );
  AND2_X1 U13934 ( .A1(n13905), .A2(n13904), .ZN(n13943) );
  AND2_X1 U13935 ( .A1(n13902), .A2(n13944), .ZN(n13942) );
  OR2_X1 U13936 ( .A1(n13904), .A2(n13905), .ZN(n13944) );
  OR2_X1 U13937 ( .A1(n7620), .A2(n8191), .ZN(n13905) );
  OR2_X1 U13938 ( .A1(n13945), .A2(n13946), .ZN(n13904) );
  AND2_X1 U13939 ( .A1(n13901), .A2(n13900), .ZN(n13946) );
  AND2_X1 U13940 ( .A1(n13898), .A2(n13947), .ZN(n13945) );
  OR2_X1 U13941 ( .A1(n13900), .A2(n13901), .ZN(n13947) );
  OR2_X1 U13942 ( .A1(n7620), .A2(n8186), .ZN(n13901) );
  OR2_X1 U13943 ( .A1(n13948), .A2(n13949), .ZN(n13900) );
  AND2_X1 U13944 ( .A1(n13897), .A2(n13896), .ZN(n13949) );
  AND2_X1 U13945 ( .A1(n13894), .A2(n13950), .ZN(n13948) );
  OR2_X1 U13946 ( .A1(n13896), .A2(n13897), .ZN(n13950) );
  OR2_X1 U13947 ( .A1(n7620), .A2(n8181), .ZN(n13897) );
  OR2_X1 U13948 ( .A1(n13951), .A2(n13952), .ZN(n13896) );
  AND2_X1 U13949 ( .A1(n13893), .A2(n13892), .ZN(n13952) );
  AND2_X1 U13950 ( .A1(n13890), .A2(n13953), .ZN(n13951) );
  OR2_X1 U13951 ( .A1(n13892), .A2(n13893), .ZN(n13953) );
  OR2_X1 U13952 ( .A1(n7620), .A2(n8176), .ZN(n13893) );
  OR2_X1 U13953 ( .A1(n13954), .A2(n13955), .ZN(n13892) );
  AND2_X1 U13954 ( .A1(n13889), .A2(n13888), .ZN(n13955) );
  AND2_X1 U13955 ( .A1(n13886), .A2(n13956), .ZN(n13954) );
  OR2_X1 U13956 ( .A1(n13888), .A2(n13889), .ZN(n13956) );
  OR2_X1 U13957 ( .A1(n7620), .A2(n8171), .ZN(n13889) );
  OR2_X1 U13958 ( .A1(n13957), .A2(n13958), .ZN(n13888) );
  AND2_X1 U13959 ( .A1(n13885), .A2(n13884), .ZN(n13958) );
  AND2_X1 U13960 ( .A1(n13882), .A2(n13959), .ZN(n13957) );
  OR2_X1 U13961 ( .A1(n13884), .A2(n13885), .ZN(n13959) );
  OR2_X1 U13962 ( .A1(n8166), .A2(n7620), .ZN(n13885) );
  OR2_X1 U13963 ( .A1(n13960), .A2(n13961), .ZN(n13884) );
  AND2_X1 U13964 ( .A1(n13881), .A2(n13880), .ZN(n13961) );
  AND2_X1 U13965 ( .A1(n13878), .A2(n13962), .ZN(n13960) );
  OR2_X1 U13966 ( .A1(n13880), .A2(n13881), .ZN(n13962) );
  OR2_X1 U13967 ( .A1(n8161), .A2(n7620), .ZN(n13881) );
  OR2_X1 U13968 ( .A1(n13963), .A2(n13964), .ZN(n13880) );
  AND2_X1 U13969 ( .A1(n13877), .A2(n13876), .ZN(n13964) );
  AND2_X1 U13970 ( .A1(n13874), .A2(n13965), .ZN(n13963) );
  OR2_X1 U13971 ( .A1(n13876), .A2(n13877), .ZN(n13965) );
  OR2_X1 U13972 ( .A1(n8156), .A2(n7620), .ZN(n13877) );
  OR2_X1 U13973 ( .A1(n13966), .A2(n13967), .ZN(n13876) );
  AND2_X1 U13974 ( .A1(n13873), .A2(n13872), .ZN(n13967) );
  AND2_X1 U13975 ( .A1(n13870), .A2(n13968), .ZN(n13966) );
  OR2_X1 U13976 ( .A1(n13872), .A2(n13873), .ZN(n13968) );
  OR2_X1 U13977 ( .A1(n8151), .A2(n7620), .ZN(n13873) );
  OR2_X1 U13978 ( .A1(n13969), .A2(n13970), .ZN(n13872) );
  AND2_X1 U13979 ( .A1(n13869), .A2(n13868), .ZN(n13970) );
  AND2_X1 U13980 ( .A1(n13866), .A2(n13971), .ZN(n13969) );
  OR2_X1 U13981 ( .A1(n13868), .A2(n13869), .ZN(n13971) );
  OR2_X1 U13982 ( .A1(n8146), .A2(n7620), .ZN(n13869) );
  OR2_X1 U13983 ( .A1(n13972), .A2(n13973), .ZN(n13868) );
  AND2_X1 U13984 ( .A1(n13865), .A2(n13864), .ZN(n13973) );
  AND2_X1 U13985 ( .A1(n13862), .A2(n13974), .ZN(n13972) );
  OR2_X1 U13986 ( .A1(n13864), .A2(n13865), .ZN(n13974) );
  OR2_X1 U13987 ( .A1(n8141), .A2(n7620), .ZN(n13865) );
  OR2_X1 U13988 ( .A1(n13975), .A2(n13976), .ZN(n13864) );
  AND2_X1 U13989 ( .A1(n13861), .A2(n13860), .ZN(n13976) );
  AND2_X1 U13990 ( .A1(n13858), .A2(n13977), .ZN(n13975) );
  OR2_X1 U13991 ( .A1(n13860), .A2(n13861), .ZN(n13977) );
  OR2_X1 U13992 ( .A1(n8136), .A2(n7620), .ZN(n13861) );
  OR2_X1 U13993 ( .A1(n13978), .A2(n13979), .ZN(n13860) );
  AND2_X1 U13994 ( .A1(n13857), .A2(n13856), .ZN(n13979) );
  AND2_X1 U13995 ( .A1(n13854), .A2(n13980), .ZN(n13978) );
  OR2_X1 U13996 ( .A1(n13856), .A2(n13857), .ZN(n13980) );
  OR2_X1 U13997 ( .A1(n8131), .A2(n7620), .ZN(n13857) );
  OR2_X1 U13998 ( .A1(n13981), .A2(n13982), .ZN(n13856) );
  AND2_X1 U13999 ( .A1(n13853), .A2(n13852), .ZN(n13982) );
  AND2_X1 U14000 ( .A1(n13850), .A2(n13983), .ZN(n13981) );
  OR2_X1 U14001 ( .A1(n13852), .A2(n13853), .ZN(n13983) );
  OR2_X1 U14002 ( .A1(n8126), .A2(n7620), .ZN(n13853) );
  OR2_X1 U14003 ( .A1(n13984), .A2(n13985), .ZN(n13852) );
  AND2_X1 U14004 ( .A1(n13846), .A2(n13849), .ZN(n13985) );
  AND2_X1 U14005 ( .A1(n13986), .A2(n13848), .ZN(n13984) );
  OR2_X1 U14006 ( .A1(n13987), .A2(n13988), .ZN(n13848) );
  AND2_X1 U14007 ( .A1(n13845), .A2(n13844), .ZN(n13988) );
  AND2_X1 U14008 ( .A1(n13842), .A2(n13989), .ZN(n13987) );
  OR2_X1 U14009 ( .A1(n13844), .A2(n13845), .ZN(n13989) );
  OR2_X1 U14010 ( .A1(n8116), .A2(n7620), .ZN(n13845) );
  OR2_X1 U14011 ( .A1(n13990), .A2(n13991), .ZN(n13844) );
  AND2_X1 U14012 ( .A1(n13838), .A2(n13841), .ZN(n13991) );
  AND2_X1 U14013 ( .A1(n13992), .A2(n13840), .ZN(n13990) );
  OR2_X1 U14014 ( .A1(n13993), .A2(n13994), .ZN(n13840) );
  AND2_X1 U14015 ( .A1(n13834), .A2(n13837), .ZN(n13994) );
  AND2_X1 U14016 ( .A1(n13836), .A2(n13995), .ZN(n13993) );
  OR2_X1 U14017 ( .A1(n13837), .A2(n13834), .ZN(n13995) );
  OR2_X1 U14018 ( .A1(n8102), .A2(n7620), .ZN(n13834) );
  OR3_X1 U14019 ( .A1(n8349), .A2(n7620), .A3(n13831), .ZN(n13837) );
  INV_X1 U14020 ( .A(n13996), .ZN(n13836) );
  OR2_X1 U14021 ( .A1(n13997), .A2(n13998), .ZN(n13996) );
  AND2_X1 U14022 ( .A1(b_2_), .A2(n13999), .ZN(n13998) );
  OR2_X1 U14023 ( .A1(n14000), .A2(n7314), .ZN(n13999) );
  AND2_X1 U14024 ( .A1(a_30_), .A2(n14001), .ZN(n14000) );
  AND2_X1 U14025 ( .A1(b_1_), .A2(n14002), .ZN(n13997) );
  OR2_X1 U14026 ( .A1(n14003), .A2(n7318), .ZN(n14002) );
  AND2_X1 U14027 ( .A1(a_31_), .A2(n13831), .ZN(n14003) );
  OR2_X1 U14028 ( .A1(n13841), .A2(n13838), .ZN(n13992) );
  XNOR2_X1 U14029 ( .A(n14004), .B(n14005), .ZN(n13838) );
  XNOR2_X1 U14030 ( .A(n14006), .B(n14007), .ZN(n14005) );
  OR2_X1 U14031 ( .A1(n8111), .A2(n7620), .ZN(n13841) );
  XOR2_X1 U14032 ( .A(n14008), .B(n14009), .Z(n13842) );
  XOR2_X1 U14033 ( .A(n14010), .B(n14011), .Z(n14009) );
  OR2_X1 U14034 ( .A1(n13849), .A2(n13846), .ZN(n13986) );
  XOR2_X1 U14035 ( .A(n14012), .B(n14013), .Z(n13846) );
  XOR2_X1 U14036 ( .A(n14014), .B(n14015), .Z(n14013) );
  OR2_X1 U14037 ( .A1(n8121), .A2(n7620), .ZN(n13849) );
  XOR2_X1 U14038 ( .A(n14016), .B(n14017), .Z(n13850) );
  XOR2_X1 U14039 ( .A(n14018), .B(n14019), .Z(n14017) );
  XOR2_X1 U14040 ( .A(n14020), .B(n14021), .Z(n13854) );
  XOR2_X1 U14041 ( .A(n14022), .B(n14023), .Z(n14021) );
  XOR2_X1 U14042 ( .A(n14024), .B(n14025), .Z(n13858) );
  XOR2_X1 U14043 ( .A(n14026), .B(n14027), .Z(n14025) );
  XOR2_X1 U14044 ( .A(n14028), .B(n14029), .Z(n13862) );
  XOR2_X1 U14045 ( .A(n14030), .B(n14031), .Z(n14029) );
  XOR2_X1 U14046 ( .A(n14032), .B(n14033), .Z(n13866) );
  XOR2_X1 U14047 ( .A(n14034), .B(n14035), .Z(n14033) );
  XOR2_X1 U14048 ( .A(n14036), .B(n14037), .Z(n13870) );
  XOR2_X1 U14049 ( .A(n14038), .B(n14039), .Z(n14037) );
  XOR2_X1 U14050 ( .A(n14040), .B(n14041), .Z(n13874) );
  XOR2_X1 U14051 ( .A(n14042), .B(n14043), .Z(n14041) );
  XOR2_X1 U14052 ( .A(n14044), .B(n14045), .Z(n13878) );
  XOR2_X1 U14053 ( .A(n14046), .B(n14047), .Z(n14045) );
  XOR2_X1 U14054 ( .A(n14048), .B(n14049), .Z(n13882) );
  XOR2_X1 U14055 ( .A(n14050), .B(n14051), .Z(n14049) );
  XOR2_X1 U14056 ( .A(n14052), .B(n14053), .Z(n13886) );
  XOR2_X1 U14057 ( .A(n14054), .B(n14055), .Z(n14053) );
  XOR2_X1 U14058 ( .A(n14056), .B(n14057), .Z(n13890) );
  XOR2_X1 U14059 ( .A(n14058), .B(n14059), .Z(n14057) );
  XOR2_X1 U14060 ( .A(n14060), .B(n14061), .Z(n13894) );
  XOR2_X1 U14061 ( .A(n14062), .B(n14063), .Z(n14061) );
  XOR2_X1 U14062 ( .A(n14064), .B(n14065), .Z(n13898) );
  XOR2_X1 U14063 ( .A(n14066), .B(n14067), .Z(n14065) );
  XOR2_X1 U14064 ( .A(n14068), .B(n14069), .Z(n13902) );
  XOR2_X1 U14065 ( .A(n14070), .B(n14071), .Z(n14069) );
  XOR2_X1 U14066 ( .A(n14072), .B(n14073), .Z(n13906) );
  XOR2_X1 U14067 ( .A(n14074), .B(n14075), .Z(n14073) );
  XOR2_X1 U14068 ( .A(n14076), .B(n14077), .Z(n13910) );
  XOR2_X1 U14069 ( .A(n14078), .B(n14079), .Z(n14077) );
  XOR2_X1 U14070 ( .A(n14080), .B(n14081), .Z(n13914) );
  XOR2_X1 U14071 ( .A(n14082), .B(n14083), .Z(n14081) );
  XOR2_X1 U14072 ( .A(n14084), .B(n14085), .Z(n13918) );
  XOR2_X1 U14073 ( .A(n14086), .B(n14087), .Z(n14085) );
  XOR2_X1 U14074 ( .A(n14088), .B(n14089), .Z(n13922) );
  XOR2_X1 U14075 ( .A(n14090), .B(n14091), .Z(n14089) );
  XOR2_X1 U14076 ( .A(n14092), .B(n14093), .Z(n13745) );
  XOR2_X1 U14077 ( .A(n14094), .B(n14095), .Z(n14093) );
  AND3_X1 U14078 ( .A1(n7521), .A2(n7519), .A3(n7520), .ZN(n7522) );
  INV_X1 U14079 ( .A(n7593), .ZN(n7520) );
  OR2_X1 U14080 ( .A1(n14096), .A2(n14097), .ZN(n7593) );
  AND2_X1 U14081 ( .A1(n7612), .A2(n7611), .ZN(n14097) );
  AND2_X1 U14082 ( .A1(n7609), .A2(n14098), .ZN(n14096) );
  OR2_X1 U14083 ( .A1(n7611), .A2(n7612), .ZN(n14098) );
  OR2_X1 U14084 ( .A1(n13831), .A2(n7621), .ZN(n7612) );
  OR2_X1 U14085 ( .A1(n14099), .A2(n14100), .ZN(n7611) );
  AND2_X1 U14086 ( .A1(n7631), .A2(n7630), .ZN(n14100) );
  AND2_X1 U14087 ( .A1(n7628), .A2(n14101), .ZN(n14099) );
  OR2_X1 U14088 ( .A1(n7630), .A2(n7631), .ZN(n14101) );
  OR2_X1 U14089 ( .A1(n13831), .A2(n7656), .ZN(n7631) );
  OR2_X1 U14090 ( .A1(n14102), .A2(n14103), .ZN(n7630) );
  AND2_X1 U14091 ( .A1(n7664), .A2(n7666), .ZN(n14103) );
  AND2_X1 U14092 ( .A1(n14104), .A2(n7665), .ZN(n14102) );
  OR2_X1 U14093 ( .A1(n7664), .A2(n7666), .ZN(n14104) );
  OR2_X1 U14094 ( .A1(n14105), .A2(n14106), .ZN(n7666) );
  AND2_X1 U14095 ( .A1(n7699), .A2(n7698), .ZN(n14106) );
  AND2_X1 U14096 ( .A1(n7696), .A2(n14107), .ZN(n14105) );
  OR2_X1 U14097 ( .A1(n7698), .A2(n7699), .ZN(n14107) );
  OR2_X1 U14098 ( .A1(n13831), .A2(n7777), .ZN(n7699) );
  OR2_X1 U14099 ( .A1(n14108), .A2(n14109), .ZN(n7698) );
  AND2_X1 U14100 ( .A1(n7741), .A2(n7740), .ZN(n14109) );
  AND2_X1 U14101 ( .A1(n7738), .A2(n14110), .ZN(n14108) );
  OR2_X1 U14102 ( .A1(n7740), .A2(n7741), .ZN(n14110) );
  OR2_X1 U14103 ( .A1(n13831), .A2(n7785), .ZN(n7741) );
  OR2_X1 U14104 ( .A1(n14111), .A2(n14112), .ZN(n7740) );
  AND2_X1 U14105 ( .A1(n7795), .A2(n7794), .ZN(n14112) );
  AND2_X1 U14106 ( .A1(n7792), .A2(n14113), .ZN(n14111) );
  OR2_X1 U14107 ( .A1(n7794), .A2(n7795), .ZN(n14113) );
  OR2_X1 U14108 ( .A1(n13831), .A2(n8226), .ZN(n7795) );
  OR2_X1 U14109 ( .A1(n14114), .A2(n14115), .ZN(n7794) );
  AND2_X1 U14110 ( .A1(n13750), .A2(n13749), .ZN(n14115) );
  AND2_X1 U14111 ( .A1(n13747), .A2(n14116), .ZN(n14114) );
  OR2_X1 U14112 ( .A1(n13749), .A2(n13750), .ZN(n14116) );
  OR2_X1 U14113 ( .A1(n13831), .A2(n8221), .ZN(n13750) );
  OR2_X1 U14114 ( .A1(n14117), .A2(n14118), .ZN(n13749) );
  AND2_X1 U14115 ( .A1(n14095), .A2(n14094), .ZN(n14118) );
  AND2_X1 U14116 ( .A1(n14092), .A2(n14119), .ZN(n14117) );
  OR2_X1 U14117 ( .A1(n14094), .A2(n14095), .ZN(n14119) );
  OR2_X1 U14118 ( .A1(n13831), .A2(n8216), .ZN(n14095) );
  OR2_X1 U14119 ( .A1(n14120), .A2(n14121), .ZN(n14094) );
  AND2_X1 U14120 ( .A1(n14091), .A2(n14090), .ZN(n14121) );
  AND2_X1 U14121 ( .A1(n14088), .A2(n14122), .ZN(n14120) );
  OR2_X1 U14122 ( .A1(n14090), .A2(n14091), .ZN(n14122) );
  OR2_X1 U14123 ( .A1(n13831), .A2(n8211), .ZN(n14091) );
  OR2_X1 U14124 ( .A1(n14123), .A2(n14124), .ZN(n14090) );
  AND2_X1 U14125 ( .A1(n14087), .A2(n14086), .ZN(n14124) );
  AND2_X1 U14126 ( .A1(n14084), .A2(n14125), .ZN(n14123) );
  OR2_X1 U14127 ( .A1(n14086), .A2(n14087), .ZN(n14125) );
  OR2_X1 U14128 ( .A1(n13831), .A2(n8206), .ZN(n14087) );
  OR2_X1 U14129 ( .A1(n14126), .A2(n14127), .ZN(n14086) );
  AND2_X1 U14130 ( .A1(n14083), .A2(n14082), .ZN(n14127) );
  AND2_X1 U14131 ( .A1(n14080), .A2(n14128), .ZN(n14126) );
  OR2_X1 U14132 ( .A1(n14082), .A2(n14083), .ZN(n14128) );
  OR2_X1 U14133 ( .A1(n13831), .A2(n8201), .ZN(n14083) );
  OR2_X1 U14134 ( .A1(n14129), .A2(n14130), .ZN(n14082) );
  AND2_X1 U14135 ( .A1(n14079), .A2(n14078), .ZN(n14130) );
  AND2_X1 U14136 ( .A1(n14076), .A2(n14131), .ZN(n14129) );
  OR2_X1 U14137 ( .A1(n14078), .A2(n14079), .ZN(n14131) );
  OR2_X1 U14138 ( .A1(n13831), .A2(n8196), .ZN(n14079) );
  OR2_X1 U14139 ( .A1(n14132), .A2(n14133), .ZN(n14078) );
  AND2_X1 U14140 ( .A1(n14075), .A2(n14074), .ZN(n14133) );
  AND2_X1 U14141 ( .A1(n14072), .A2(n14134), .ZN(n14132) );
  OR2_X1 U14142 ( .A1(n14074), .A2(n14075), .ZN(n14134) );
  OR2_X1 U14143 ( .A1(n13831), .A2(n8191), .ZN(n14075) );
  OR2_X1 U14144 ( .A1(n14135), .A2(n14136), .ZN(n14074) );
  AND2_X1 U14145 ( .A1(n14071), .A2(n14070), .ZN(n14136) );
  AND2_X1 U14146 ( .A1(n14068), .A2(n14137), .ZN(n14135) );
  OR2_X1 U14147 ( .A1(n14070), .A2(n14071), .ZN(n14137) );
  OR2_X1 U14148 ( .A1(n13831), .A2(n8186), .ZN(n14071) );
  OR2_X1 U14149 ( .A1(n14138), .A2(n14139), .ZN(n14070) );
  AND2_X1 U14150 ( .A1(n14067), .A2(n14066), .ZN(n14139) );
  AND2_X1 U14151 ( .A1(n14064), .A2(n14140), .ZN(n14138) );
  OR2_X1 U14152 ( .A1(n14066), .A2(n14067), .ZN(n14140) );
  OR2_X1 U14153 ( .A1(n13831), .A2(n8181), .ZN(n14067) );
  OR2_X1 U14154 ( .A1(n14141), .A2(n14142), .ZN(n14066) );
  AND2_X1 U14155 ( .A1(n14063), .A2(n14062), .ZN(n14142) );
  AND2_X1 U14156 ( .A1(n14060), .A2(n14143), .ZN(n14141) );
  OR2_X1 U14157 ( .A1(n14062), .A2(n14063), .ZN(n14143) );
  OR2_X1 U14158 ( .A1(n13831), .A2(n8176), .ZN(n14063) );
  OR2_X1 U14159 ( .A1(n14144), .A2(n14145), .ZN(n14062) );
  AND2_X1 U14160 ( .A1(n14059), .A2(n14058), .ZN(n14145) );
  AND2_X1 U14161 ( .A1(n14056), .A2(n14146), .ZN(n14144) );
  OR2_X1 U14162 ( .A1(n14058), .A2(n14059), .ZN(n14146) );
  OR2_X1 U14163 ( .A1(n8171), .A2(n13831), .ZN(n14059) );
  OR2_X1 U14164 ( .A1(n14147), .A2(n14148), .ZN(n14058) );
  AND2_X1 U14165 ( .A1(n14055), .A2(n14054), .ZN(n14148) );
  AND2_X1 U14166 ( .A1(n14052), .A2(n14149), .ZN(n14147) );
  OR2_X1 U14167 ( .A1(n14054), .A2(n14055), .ZN(n14149) );
  OR2_X1 U14168 ( .A1(n8166), .A2(n13831), .ZN(n14055) );
  OR2_X1 U14169 ( .A1(n14150), .A2(n14151), .ZN(n14054) );
  AND2_X1 U14170 ( .A1(n14051), .A2(n14050), .ZN(n14151) );
  AND2_X1 U14171 ( .A1(n14048), .A2(n14152), .ZN(n14150) );
  OR2_X1 U14172 ( .A1(n14050), .A2(n14051), .ZN(n14152) );
  OR2_X1 U14173 ( .A1(n8161), .A2(n13831), .ZN(n14051) );
  OR2_X1 U14174 ( .A1(n14153), .A2(n14154), .ZN(n14050) );
  AND2_X1 U14175 ( .A1(n14047), .A2(n14046), .ZN(n14154) );
  AND2_X1 U14176 ( .A1(n14044), .A2(n14155), .ZN(n14153) );
  OR2_X1 U14177 ( .A1(n14046), .A2(n14047), .ZN(n14155) );
  OR2_X1 U14178 ( .A1(n8156), .A2(n13831), .ZN(n14047) );
  OR2_X1 U14179 ( .A1(n14156), .A2(n14157), .ZN(n14046) );
  AND2_X1 U14180 ( .A1(n14043), .A2(n14042), .ZN(n14157) );
  AND2_X1 U14181 ( .A1(n14040), .A2(n14158), .ZN(n14156) );
  OR2_X1 U14182 ( .A1(n14042), .A2(n14043), .ZN(n14158) );
  OR2_X1 U14183 ( .A1(n8151), .A2(n13831), .ZN(n14043) );
  OR2_X1 U14184 ( .A1(n14159), .A2(n14160), .ZN(n14042) );
  AND2_X1 U14185 ( .A1(n14039), .A2(n14038), .ZN(n14160) );
  AND2_X1 U14186 ( .A1(n14036), .A2(n14161), .ZN(n14159) );
  OR2_X1 U14187 ( .A1(n14038), .A2(n14039), .ZN(n14161) );
  OR2_X1 U14188 ( .A1(n8146), .A2(n13831), .ZN(n14039) );
  OR2_X1 U14189 ( .A1(n14162), .A2(n14163), .ZN(n14038) );
  AND2_X1 U14190 ( .A1(n14035), .A2(n14034), .ZN(n14163) );
  AND2_X1 U14191 ( .A1(n14032), .A2(n14164), .ZN(n14162) );
  OR2_X1 U14192 ( .A1(n14034), .A2(n14035), .ZN(n14164) );
  OR2_X1 U14193 ( .A1(n8141), .A2(n13831), .ZN(n14035) );
  OR2_X1 U14194 ( .A1(n14165), .A2(n14166), .ZN(n14034) );
  AND2_X1 U14195 ( .A1(n14031), .A2(n14030), .ZN(n14166) );
  AND2_X1 U14196 ( .A1(n14028), .A2(n14167), .ZN(n14165) );
  OR2_X1 U14197 ( .A1(n14030), .A2(n14031), .ZN(n14167) );
  OR2_X1 U14198 ( .A1(n8136), .A2(n13831), .ZN(n14031) );
  OR2_X1 U14199 ( .A1(n14168), .A2(n14169), .ZN(n14030) );
  AND2_X1 U14200 ( .A1(n14027), .A2(n14026), .ZN(n14169) );
  AND2_X1 U14201 ( .A1(n14024), .A2(n14170), .ZN(n14168) );
  OR2_X1 U14202 ( .A1(n14026), .A2(n14027), .ZN(n14170) );
  OR2_X1 U14203 ( .A1(n8131), .A2(n13831), .ZN(n14027) );
  OR2_X1 U14204 ( .A1(n14171), .A2(n14172), .ZN(n14026) );
  AND2_X1 U14205 ( .A1(n14023), .A2(n14022), .ZN(n14172) );
  AND2_X1 U14206 ( .A1(n14020), .A2(n14173), .ZN(n14171) );
  OR2_X1 U14207 ( .A1(n14022), .A2(n14023), .ZN(n14173) );
  OR2_X1 U14208 ( .A1(n8126), .A2(n13831), .ZN(n14023) );
  OR2_X1 U14209 ( .A1(n14174), .A2(n14175), .ZN(n14022) );
  AND2_X1 U14210 ( .A1(n14019), .A2(n14018), .ZN(n14175) );
  AND2_X1 U14211 ( .A1(n14016), .A2(n14176), .ZN(n14174) );
  OR2_X1 U14212 ( .A1(n14018), .A2(n14019), .ZN(n14176) );
  OR2_X1 U14213 ( .A1(n8121), .A2(n13831), .ZN(n14019) );
  OR2_X1 U14214 ( .A1(n14177), .A2(n14178), .ZN(n14018) );
  AND2_X1 U14215 ( .A1(n14012), .A2(n14015), .ZN(n14178) );
  AND2_X1 U14216 ( .A1(n14179), .A2(n14014), .ZN(n14177) );
  OR2_X1 U14217 ( .A1(n14180), .A2(n14181), .ZN(n14014) );
  AND2_X1 U14218 ( .A1(n14011), .A2(n14010), .ZN(n14181) );
  AND2_X1 U14219 ( .A1(n14008), .A2(n14182), .ZN(n14180) );
  OR2_X1 U14220 ( .A1(n14010), .A2(n14011), .ZN(n14182) );
  OR2_X1 U14221 ( .A1(n8111), .A2(n13831), .ZN(n14011) );
  OR2_X1 U14222 ( .A1(n14183), .A2(n14184), .ZN(n14010) );
  AND2_X1 U14223 ( .A1(n14004), .A2(n14007), .ZN(n14184) );
  AND2_X1 U14224 ( .A1(n14006), .A2(n14185), .ZN(n14183) );
  OR2_X1 U14225 ( .A1(n14007), .A2(n14004), .ZN(n14185) );
  OR2_X1 U14226 ( .A1(n8102), .A2(n13831), .ZN(n14004) );
  OR3_X1 U14227 ( .A1(n8349), .A2(n13831), .A3(n14001), .ZN(n14007) );
  INV_X1 U14228 ( .A(n14186), .ZN(n14006) );
  OR2_X1 U14229 ( .A1(n14187), .A2(n14188), .ZN(n14186) );
  AND2_X1 U14230 ( .A1(b_1_), .A2(n14189), .ZN(n14188) );
  OR2_X1 U14231 ( .A1(n14190), .A2(n7314), .ZN(n14189) );
  AND2_X1 U14232 ( .A1(n14191), .A2(a_30_), .ZN(n7314) );
  AND2_X1 U14233 ( .A1(a_30_), .A2(n14192), .ZN(n14190) );
  AND2_X1 U14234 ( .A1(b_0_), .A2(n14193), .ZN(n14187) );
  OR2_X1 U14235 ( .A1(n14194), .A2(n7318), .ZN(n14193) );
  AND2_X1 U14236 ( .A1(n14195), .A2(a_31_), .ZN(n7318) );
  AND2_X1 U14237 ( .A1(a_31_), .A2(n14001), .ZN(n14194) );
  XNOR2_X1 U14238 ( .A(n14196), .B(n14197), .ZN(n14008) );
  OR2_X1 U14239 ( .A1(n14198), .A2(n14199), .ZN(n14196) );
  AND2_X1 U14240 ( .A1(n14200), .A2(n14201), .ZN(n14198) );
  INV_X1 U14241 ( .A(n14202), .ZN(n14201) );
  OR2_X1 U14242 ( .A1(n14195), .A2(n14192), .ZN(n14200) );
  OR2_X1 U14243 ( .A1(n14015), .A2(n14012), .ZN(n14179) );
  XNOR2_X1 U14244 ( .A(n14203), .B(n14204), .ZN(n14012) );
  XNOR2_X1 U14245 ( .A(n14205), .B(n14206), .ZN(n14204) );
  OR2_X1 U14246 ( .A1(n8116), .A2(n13831), .ZN(n14015) );
  XNOR2_X1 U14247 ( .A(n14207), .B(n14208), .ZN(n14016) );
  XNOR2_X1 U14248 ( .A(n14209), .B(n14210), .ZN(n14207) );
  XNOR2_X1 U14249 ( .A(n14211), .B(n14212), .ZN(n14020) );
  XNOR2_X1 U14250 ( .A(n14213), .B(n14214), .ZN(n14211) );
  XNOR2_X1 U14251 ( .A(n14215), .B(n14216), .ZN(n14024) );
  XNOR2_X1 U14252 ( .A(n14217), .B(n14218), .ZN(n14215) );
  XNOR2_X1 U14253 ( .A(n14219), .B(n14220), .ZN(n14028) );
  XNOR2_X1 U14254 ( .A(n14221), .B(n14222), .ZN(n14219) );
  XNOR2_X1 U14255 ( .A(n14223), .B(n14224), .ZN(n14032) );
  XNOR2_X1 U14256 ( .A(n14225), .B(n14226), .ZN(n14223) );
  XNOR2_X1 U14257 ( .A(n14227), .B(n14228), .ZN(n14036) );
  XNOR2_X1 U14258 ( .A(n14229), .B(n14230), .ZN(n14227) );
  XNOR2_X1 U14259 ( .A(n14231), .B(n14232), .ZN(n14040) );
  XNOR2_X1 U14260 ( .A(n14233), .B(n14234), .ZN(n14231) );
  XNOR2_X1 U14261 ( .A(n14235), .B(n14236), .ZN(n14044) );
  XNOR2_X1 U14262 ( .A(n14237), .B(n14238), .ZN(n14235) );
  XNOR2_X1 U14263 ( .A(n14239), .B(n14240), .ZN(n14048) );
  XNOR2_X1 U14264 ( .A(n14241), .B(n14242), .ZN(n14239) );
  XNOR2_X1 U14265 ( .A(n14243), .B(n14244), .ZN(n14052) );
  XNOR2_X1 U14266 ( .A(n14245), .B(n14246), .ZN(n14243) );
  XNOR2_X1 U14267 ( .A(n14247), .B(n14248), .ZN(n14056) );
  XNOR2_X1 U14268 ( .A(n14249), .B(n14250), .ZN(n14247) );
  XNOR2_X1 U14269 ( .A(n14251), .B(n14252), .ZN(n14060) );
  XNOR2_X1 U14270 ( .A(n14253), .B(n14254), .ZN(n14251) );
  XNOR2_X1 U14271 ( .A(n14255), .B(n14256), .ZN(n14064) );
  XNOR2_X1 U14272 ( .A(n14257), .B(n14258), .ZN(n14255) );
  XNOR2_X1 U14273 ( .A(n14259), .B(n14260), .ZN(n14068) );
  XNOR2_X1 U14274 ( .A(n14261), .B(n14262), .ZN(n14259) );
  XNOR2_X1 U14275 ( .A(n14263), .B(n14264), .ZN(n14072) );
  XNOR2_X1 U14276 ( .A(n14265), .B(n14266), .ZN(n14263) );
  XNOR2_X1 U14277 ( .A(n14267), .B(n14268), .ZN(n14076) );
  XNOR2_X1 U14278 ( .A(n14269), .B(n14270), .ZN(n14267) );
  XNOR2_X1 U14279 ( .A(n14271), .B(n14272), .ZN(n14080) );
  XNOR2_X1 U14280 ( .A(n14273), .B(n14274), .ZN(n14271) );
  XNOR2_X1 U14281 ( .A(n14275), .B(n14276), .ZN(n14084) );
  XNOR2_X1 U14282 ( .A(n14277), .B(n14278), .ZN(n14275) );
  XNOR2_X1 U14283 ( .A(n14279), .B(n14280), .ZN(n14088) );
  XNOR2_X1 U14284 ( .A(n14281), .B(n14282), .ZN(n14279) );
  XOR2_X1 U14285 ( .A(n14283), .B(n14284), .Z(n14092) );
  XOR2_X1 U14286 ( .A(n14285), .B(n14286), .Z(n14284) );
  XOR2_X1 U14287 ( .A(n14287), .B(n14288), .Z(n13747) );
  XOR2_X1 U14288 ( .A(n14289), .B(n14290), .Z(n14288) );
  XOR2_X1 U14289 ( .A(n14291), .B(n14292), .Z(n7792) );
  XOR2_X1 U14290 ( .A(n14293), .B(n14294), .Z(n14292) );
  XOR2_X1 U14291 ( .A(n14295), .B(n14296), .Z(n7738) );
  XOR2_X1 U14292 ( .A(n14297), .B(n14298), .Z(n14296) );
  XOR2_X1 U14293 ( .A(n14299), .B(n14300), .Z(n7696) );
  XOR2_X1 U14294 ( .A(n14301), .B(n14302), .Z(n14300) );
  XOR2_X1 U14295 ( .A(n14303), .B(n14304), .Z(n7664) );
  XOR2_X1 U14296 ( .A(n14305), .B(n14306), .Z(n14304) );
  XOR2_X1 U14297 ( .A(n14307), .B(n14308), .Z(n7628) );
  XOR2_X1 U14298 ( .A(n14309), .B(n14310), .Z(n14308) );
  XOR2_X1 U14299 ( .A(n14311), .B(n14312), .Z(n7609) );
  XOR2_X1 U14300 ( .A(n14313), .B(n14314), .Z(n14312) );
  XOR2_X1 U14301 ( .A(n14315), .B(n7592), .Z(n7519) );
  OR2_X1 U14302 ( .A1(n14316), .A2(n14317), .ZN(n7592) );
  AND2_X1 U14303 ( .A1(n14318), .A2(n14319), .ZN(n14317) );
  AND2_X1 U14304 ( .A1(n14320), .A2(n14321), .ZN(n14316) );
  OR2_X1 U14305 ( .A1(n14319), .A2(n14318), .ZN(n14320) );
  OR2_X1 U14306 ( .A1(n14192), .A2(n7621), .ZN(n14315) );
  XOR2_X1 U14307 ( .A(n14322), .B(n14318), .Z(n7521) );
  OR2_X1 U14308 ( .A1(n14323), .A2(n14324), .ZN(n14318) );
  AND2_X1 U14309 ( .A1(n14311), .A2(n14313), .ZN(n14324) );
  AND2_X1 U14310 ( .A1(n14325), .A2(n14314), .ZN(n14323) );
  OR2_X1 U14311 ( .A1(n14313), .A2(n14311), .ZN(n14325) );
  OR2_X1 U14312 ( .A1(n14192), .A2(n7689), .ZN(n14311) );
  OR2_X1 U14313 ( .A1(n14326), .A2(n14327), .ZN(n14313) );
  AND2_X1 U14314 ( .A1(n14307), .A2(n14309), .ZN(n14327) );
  AND2_X1 U14315 ( .A1(n14328), .A2(n14310), .ZN(n14326) );
  OR2_X1 U14316 ( .A1(n14192), .A2(n7777), .ZN(n14310) );
  OR2_X1 U14317 ( .A1(n14309), .A2(n14307), .ZN(n14328) );
  OR2_X1 U14318 ( .A1(n14001), .A2(n7689), .ZN(n14307) );
  OR2_X1 U14319 ( .A1(n14329), .A2(n14330), .ZN(n14309) );
  AND2_X1 U14320 ( .A1(n14303), .A2(n14305), .ZN(n14330) );
  AND2_X1 U14321 ( .A1(n14331), .A2(n14306), .ZN(n14329) );
  OR2_X1 U14322 ( .A1(n14192), .A2(n7785), .ZN(n14306) );
  OR2_X1 U14323 ( .A1(n14305), .A2(n14303), .ZN(n14331) );
  OR2_X1 U14324 ( .A1(n14001), .A2(n7777), .ZN(n14303) );
  OR2_X1 U14325 ( .A1(n14332), .A2(n14333), .ZN(n14305) );
  AND2_X1 U14326 ( .A1(n14299), .A2(n14301), .ZN(n14333) );
  AND2_X1 U14327 ( .A1(n14334), .A2(n14302), .ZN(n14332) );
  OR2_X1 U14328 ( .A1(n14192), .A2(n8226), .ZN(n14302) );
  OR2_X1 U14329 ( .A1(n14301), .A2(n14299), .ZN(n14334) );
  OR2_X1 U14330 ( .A1(n14001), .A2(n7785), .ZN(n14299) );
  OR2_X1 U14331 ( .A1(n14335), .A2(n14336), .ZN(n14301) );
  AND2_X1 U14332 ( .A1(n14295), .A2(n14297), .ZN(n14336) );
  AND2_X1 U14333 ( .A1(n14337), .A2(n14298), .ZN(n14335) );
  OR2_X1 U14334 ( .A1(n14192), .A2(n8221), .ZN(n14298) );
  OR2_X1 U14335 ( .A1(n14297), .A2(n14295), .ZN(n14337) );
  OR2_X1 U14336 ( .A1(n14001), .A2(n8226), .ZN(n14295) );
  OR2_X1 U14337 ( .A1(n14338), .A2(n14339), .ZN(n14297) );
  AND2_X1 U14338 ( .A1(n14291), .A2(n14293), .ZN(n14339) );
  AND2_X1 U14339 ( .A1(n14340), .A2(n14294), .ZN(n14338) );
  OR2_X1 U14340 ( .A1(n14192), .A2(n8216), .ZN(n14294) );
  OR2_X1 U14341 ( .A1(n14293), .A2(n14291), .ZN(n14340) );
  OR2_X1 U14342 ( .A1(n14001), .A2(n8221), .ZN(n14291) );
  OR2_X1 U14343 ( .A1(n14341), .A2(n14342), .ZN(n14293) );
  AND2_X1 U14344 ( .A1(n14287), .A2(n14289), .ZN(n14342) );
  AND2_X1 U14345 ( .A1(n14343), .A2(n14290), .ZN(n14341) );
  OR2_X1 U14346 ( .A1(n14192), .A2(n8211), .ZN(n14290) );
  OR2_X1 U14347 ( .A1(n14289), .A2(n14287), .ZN(n14343) );
  OR2_X1 U14348 ( .A1(n14001), .A2(n8216), .ZN(n14287) );
  OR2_X1 U14349 ( .A1(n14344), .A2(n14345), .ZN(n14289) );
  AND2_X1 U14350 ( .A1(n14283), .A2(n14285), .ZN(n14345) );
  AND2_X1 U14351 ( .A1(n14346), .A2(n14286), .ZN(n14344) );
  OR2_X1 U14352 ( .A1(n14192), .A2(n8206), .ZN(n14286) );
  OR2_X1 U14353 ( .A1(n14285), .A2(n14283), .ZN(n14346) );
  OR2_X1 U14354 ( .A1(n14001), .A2(n8211), .ZN(n14283) );
  OR2_X1 U14355 ( .A1(n14347), .A2(n14348), .ZN(n14285) );
  AND2_X1 U14356 ( .A1(n14280), .A2(n14282), .ZN(n14348) );
  AND2_X1 U14357 ( .A1(n14349), .A2(n14281), .ZN(n14347) );
  OR2_X1 U14358 ( .A1(n14192), .A2(n8201), .ZN(n14281) );
  OR2_X1 U14359 ( .A1(n14282), .A2(n14280), .ZN(n14349) );
  OR2_X1 U14360 ( .A1(n14001), .A2(n8206), .ZN(n14280) );
  OR2_X1 U14361 ( .A1(n14350), .A2(n14351), .ZN(n14282) );
  AND2_X1 U14362 ( .A1(n14276), .A2(n14278), .ZN(n14351) );
  AND2_X1 U14363 ( .A1(n14352), .A2(n14277), .ZN(n14350) );
  OR2_X1 U14364 ( .A1(n14192), .A2(n8196), .ZN(n14277) );
  OR2_X1 U14365 ( .A1(n14278), .A2(n14276), .ZN(n14352) );
  OR2_X1 U14366 ( .A1(n14001), .A2(n8201), .ZN(n14276) );
  OR2_X1 U14367 ( .A1(n14353), .A2(n14354), .ZN(n14278) );
  AND2_X1 U14368 ( .A1(n14272), .A2(n14274), .ZN(n14354) );
  AND2_X1 U14369 ( .A1(n14355), .A2(n14273), .ZN(n14353) );
  OR2_X1 U14370 ( .A1(n14192), .A2(n8191), .ZN(n14273) );
  OR2_X1 U14371 ( .A1(n14274), .A2(n14272), .ZN(n14355) );
  OR2_X1 U14372 ( .A1(n14001), .A2(n8196), .ZN(n14272) );
  OR2_X1 U14373 ( .A1(n14356), .A2(n14357), .ZN(n14274) );
  AND2_X1 U14374 ( .A1(n14268), .A2(n14270), .ZN(n14357) );
  AND2_X1 U14375 ( .A1(n14358), .A2(n14269), .ZN(n14356) );
  OR2_X1 U14376 ( .A1(n14192), .A2(n8186), .ZN(n14269) );
  OR2_X1 U14377 ( .A1(n14270), .A2(n14268), .ZN(n14358) );
  OR2_X1 U14378 ( .A1(n14001), .A2(n8191), .ZN(n14268) );
  OR2_X1 U14379 ( .A1(n14359), .A2(n14360), .ZN(n14270) );
  AND2_X1 U14380 ( .A1(n14264), .A2(n14266), .ZN(n14360) );
  AND2_X1 U14381 ( .A1(n14361), .A2(n14265), .ZN(n14359) );
  OR2_X1 U14382 ( .A1(n8181), .A2(n14192), .ZN(n14265) );
  OR2_X1 U14383 ( .A1(n14266), .A2(n14264), .ZN(n14361) );
  OR2_X1 U14384 ( .A1(n14001), .A2(n8186), .ZN(n14264) );
  OR2_X1 U14385 ( .A1(n14362), .A2(n14363), .ZN(n14266) );
  AND2_X1 U14386 ( .A1(n14260), .A2(n14262), .ZN(n14363) );
  AND2_X1 U14387 ( .A1(n14364), .A2(n14261), .ZN(n14362) );
  OR2_X1 U14388 ( .A1(n8176), .A2(n14192), .ZN(n14261) );
  OR2_X1 U14389 ( .A1(n14262), .A2(n14260), .ZN(n14364) );
  OR2_X1 U14390 ( .A1(n14001), .A2(n8181), .ZN(n14260) );
  OR2_X1 U14391 ( .A1(n14365), .A2(n14366), .ZN(n14262) );
  AND2_X1 U14392 ( .A1(n14256), .A2(n14258), .ZN(n14366) );
  AND2_X1 U14393 ( .A1(n14367), .A2(n14257), .ZN(n14365) );
  OR2_X1 U14394 ( .A1(n8171), .A2(n14192), .ZN(n14257) );
  OR2_X1 U14395 ( .A1(n14258), .A2(n14256), .ZN(n14367) );
  OR2_X1 U14396 ( .A1(n8176), .A2(n14001), .ZN(n14256) );
  OR2_X1 U14397 ( .A1(n14368), .A2(n14369), .ZN(n14258) );
  AND2_X1 U14398 ( .A1(n14252), .A2(n14254), .ZN(n14369) );
  AND2_X1 U14399 ( .A1(n14370), .A2(n14253), .ZN(n14368) );
  OR2_X1 U14400 ( .A1(n8166), .A2(n14192), .ZN(n14253) );
  OR2_X1 U14401 ( .A1(n14254), .A2(n14252), .ZN(n14370) );
  OR2_X1 U14402 ( .A1(n8171), .A2(n14001), .ZN(n14252) );
  OR2_X1 U14403 ( .A1(n14371), .A2(n14372), .ZN(n14254) );
  AND2_X1 U14404 ( .A1(n14248), .A2(n14250), .ZN(n14372) );
  AND2_X1 U14405 ( .A1(n14373), .A2(n14249), .ZN(n14371) );
  OR2_X1 U14406 ( .A1(n8161), .A2(n14192), .ZN(n14249) );
  OR2_X1 U14407 ( .A1(n14250), .A2(n14248), .ZN(n14373) );
  OR2_X1 U14408 ( .A1(n8166), .A2(n14001), .ZN(n14248) );
  OR2_X1 U14409 ( .A1(n14374), .A2(n14375), .ZN(n14250) );
  AND2_X1 U14410 ( .A1(n14244), .A2(n14246), .ZN(n14375) );
  AND2_X1 U14411 ( .A1(n14376), .A2(n14245), .ZN(n14374) );
  OR2_X1 U14412 ( .A1(n8156), .A2(n14192), .ZN(n14245) );
  OR2_X1 U14413 ( .A1(n14246), .A2(n14244), .ZN(n14376) );
  OR2_X1 U14414 ( .A1(n8161), .A2(n14001), .ZN(n14244) );
  OR2_X1 U14415 ( .A1(n14377), .A2(n14378), .ZN(n14246) );
  AND2_X1 U14416 ( .A1(n14240), .A2(n14242), .ZN(n14378) );
  AND2_X1 U14417 ( .A1(n14379), .A2(n14241), .ZN(n14377) );
  OR2_X1 U14418 ( .A1(n8151), .A2(n14192), .ZN(n14241) );
  OR2_X1 U14419 ( .A1(n14242), .A2(n14240), .ZN(n14379) );
  OR2_X1 U14420 ( .A1(n8156), .A2(n14001), .ZN(n14240) );
  OR2_X1 U14421 ( .A1(n14380), .A2(n14381), .ZN(n14242) );
  AND2_X1 U14422 ( .A1(n14236), .A2(n14238), .ZN(n14381) );
  AND2_X1 U14423 ( .A1(n14382), .A2(n14237), .ZN(n14380) );
  OR2_X1 U14424 ( .A1(n8146), .A2(n14192), .ZN(n14237) );
  OR2_X1 U14425 ( .A1(n14238), .A2(n14236), .ZN(n14382) );
  OR2_X1 U14426 ( .A1(n8151), .A2(n14001), .ZN(n14236) );
  OR2_X1 U14427 ( .A1(n14383), .A2(n14384), .ZN(n14238) );
  AND2_X1 U14428 ( .A1(n14232), .A2(n14234), .ZN(n14384) );
  AND2_X1 U14429 ( .A1(n14385), .A2(n14233), .ZN(n14383) );
  OR2_X1 U14430 ( .A1(n8141), .A2(n14192), .ZN(n14233) );
  OR2_X1 U14431 ( .A1(n14234), .A2(n14232), .ZN(n14385) );
  OR2_X1 U14432 ( .A1(n8146), .A2(n14001), .ZN(n14232) );
  OR2_X1 U14433 ( .A1(n14386), .A2(n14387), .ZN(n14234) );
  AND2_X1 U14434 ( .A1(n14228), .A2(n14230), .ZN(n14387) );
  AND2_X1 U14435 ( .A1(n14388), .A2(n14229), .ZN(n14386) );
  OR2_X1 U14436 ( .A1(n8136), .A2(n14192), .ZN(n14229) );
  OR2_X1 U14437 ( .A1(n14230), .A2(n14228), .ZN(n14388) );
  OR2_X1 U14438 ( .A1(n8141), .A2(n14001), .ZN(n14228) );
  OR2_X1 U14439 ( .A1(n14389), .A2(n14390), .ZN(n14230) );
  AND2_X1 U14440 ( .A1(n14224), .A2(n14226), .ZN(n14390) );
  AND2_X1 U14441 ( .A1(n14391), .A2(n14225), .ZN(n14389) );
  OR2_X1 U14442 ( .A1(n8131), .A2(n14192), .ZN(n14225) );
  OR2_X1 U14443 ( .A1(n14226), .A2(n14224), .ZN(n14391) );
  OR2_X1 U14444 ( .A1(n8136), .A2(n14001), .ZN(n14224) );
  OR2_X1 U14445 ( .A1(n14392), .A2(n14393), .ZN(n14226) );
  AND2_X1 U14446 ( .A1(n14220), .A2(n14222), .ZN(n14393) );
  AND2_X1 U14447 ( .A1(n14394), .A2(n14221), .ZN(n14392) );
  OR2_X1 U14448 ( .A1(n8126), .A2(n14192), .ZN(n14221) );
  OR2_X1 U14449 ( .A1(n14222), .A2(n14220), .ZN(n14394) );
  OR2_X1 U14450 ( .A1(n8131), .A2(n14001), .ZN(n14220) );
  OR2_X1 U14451 ( .A1(n14395), .A2(n14396), .ZN(n14222) );
  AND2_X1 U14452 ( .A1(n14216), .A2(n14218), .ZN(n14396) );
  AND2_X1 U14453 ( .A1(n14397), .A2(n14217), .ZN(n14395) );
  OR2_X1 U14454 ( .A1(n8121), .A2(n14192), .ZN(n14217) );
  OR2_X1 U14455 ( .A1(n14218), .A2(n14216), .ZN(n14397) );
  OR2_X1 U14456 ( .A1(n8126), .A2(n14001), .ZN(n14216) );
  OR2_X1 U14457 ( .A1(n14398), .A2(n14399), .ZN(n14218) );
  AND2_X1 U14458 ( .A1(n14212), .A2(n14214), .ZN(n14399) );
  AND2_X1 U14459 ( .A1(n14400), .A2(n14213), .ZN(n14398) );
  OR2_X1 U14460 ( .A1(n8116), .A2(n14192), .ZN(n14213) );
  OR2_X1 U14461 ( .A1(n14214), .A2(n14212), .ZN(n14400) );
  OR2_X1 U14462 ( .A1(n8121), .A2(n14001), .ZN(n14212) );
  OR2_X1 U14463 ( .A1(n14401), .A2(n14402), .ZN(n14214) );
  AND2_X1 U14464 ( .A1(n14208), .A2(n14210), .ZN(n14402) );
  AND2_X1 U14465 ( .A1(n14403), .A2(n14209), .ZN(n14401) );
  OR2_X1 U14466 ( .A1(n8111), .A2(n14192), .ZN(n14209) );
  OR2_X1 U14467 ( .A1(n14210), .A2(n14208), .ZN(n14403) );
  OR2_X1 U14468 ( .A1(n8116), .A2(n14001), .ZN(n14208) );
  OR2_X1 U14469 ( .A1(n14404), .A2(n14405), .ZN(n14210) );
  AND2_X1 U14470 ( .A1(n14203), .A2(n14206), .ZN(n14405) );
  AND2_X1 U14471 ( .A1(n14205), .A2(n14406), .ZN(n14404) );
  OR2_X1 U14472 ( .A1(n14206), .A2(n14203), .ZN(n14406) );
  OR2_X1 U14473 ( .A1(n8111), .A2(n14001), .ZN(n14203) );
  OR2_X1 U14474 ( .A1(n8102), .A2(n14192), .ZN(n14206) );
  INV_X1 U14475 ( .A(n14407), .ZN(n14205) );
  OR2_X1 U14476 ( .A1(n14199), .A2(n14408), .ZN(n14407) );
  INV_X1 U14477 ( .A(n14197), .ZN(n14408) );
  OR3_X1 U14478 ( .A1(n8349), .A2(n14001), .A3(n14192), .ZN(n14197) );
  OR2_X1 U14479 ( .A1(n14191), .A2(n14195), .ZN(n8349) );
  AND3_X1 U14480 ( .A1(a_30_), .A2(b_0_), .A3(n14202), .ZN(n14199) );
  AND2_X1 U14481 ( .A1(a_29_), .A2(b_1_), .ZN(n14202) );
  XNOR2_X1 U14482 ( .A(n14319), .B(n14321), .ZN(n14322) );
  OR2_X1 U14483 ( .A1(n14001), .A2(n7621), .ZN(n14321) );
  INV_X1 U14484 ( .A(a_0_), .ZN(n7621) );
  OR2_X1 U14485 ( .A1(n14192), .A2(n7656), .ZN(n14319) );
  INV_X1 U14486 ( .A(b_0_), .ZN(n14192) );
  OR3_X1 U14487 ( .A1(n14409), .A2(n14410), .A3(n14411), .ZN(Result_add_9_) );
  INV_X1 U14488 ( .A(n14412), .ZN(n14411) );
  OR2_X1 U14489 ( .A1(n14413), .A2(n12697), .ZN(n14412) );
  AND2_X1 U14490 ( .A1(n14414), .A2(n12396), .ZN(n14410) );
  XNOR2_X1 U14491 ( .A(a_9_), .B(n14413), .ZN(n14414) );
  AND3_X1 U14492 ( .A1(n14413), .A2(n8206), .A3(b_9_), .ZN(n14409) );
  XOR2_X1 U14493 ( .A(n14415), .B(n14416), .Z(Result_add_8_) );
  OR2_X1 U14494 ( .A1(n14417), .A2(n14418), .ZN(n14416) );
  OR3_X1 U14495 ( .A1(n14419), .A2(n14420), .A3(n14421), .ZN(Result_add_7_) );
  INV_X1 U14496 ( .A(n14422), .ZN(n14421) );
  OR2_X1 U14497 ( .A1(n14423), .A2(n13138), .ZN(n14422) );
  AND2_X1 U14498 ( .A1(n14424), .A2(n7755), .ZN(n14420) );
  XNOR2_X1 U14499 ( .A(a_7_), .B(n14423), .ZN(n14424) );
  AND3_X1 U14500 ( .A1(n14423), .A2(n8216), .A3(b_7_), .ZN(n14419) );
  XOR2_X1 U14501 ( .A(n14425), .B(n14426), .Z(Result_add_6_) );
  OR2_X1 U14502 ( .A1(n14427), .A2(n14428), .ZN(n14426) );
  OR3_X1 U14503 ( .A1(n14429), .A2(n14430), .A3(n14431), .ZN(Result_add_5_) );
  INV_X1 U14504 ( .A(n14432), .ZN(n14431) );
  OR2_X1 U14505 ( .A1(n14433), .A2(n13547), .ZN(n14432) );
  AND2_X1 U14506 ( .A1(n14434), .A2(n7674), .ZN(n14430) );
  XNOR2_X1 U14507 ( .A(a_5_), .B(n14433), .ZN(n14434) );
  AND3_X1 U14508 ( .A1(n14433), .A2(n8226), .A3(b_5_), .ZN(n14429) );
  XOR2_X1 U14509 ( .A(n14435), .B(n14436), .Z(Result_add_4_) );
  OR2_X1 U14510 ( .A1(n14437), .A2(n14438), .ZN(n14436) );
  OR3_X1 U14511 ( .A1(n14439), .A2(n14440), .A3(n14441), .ZN(Result_add_3_) );
  INV_X1 U14512 ( .A(n14442), .ZN(n14441) );
  OR2_X1 U14513 ( .A1(n14443), .A2(n7695), .ZN(n14442) );
  AND2_X1 U14514 ( .A1(n14444), .A2(n7620), .ZN(n14440) );
  XNOR2_X1 U14515 ( .A(a_3_), .B(n14443), .ZN(n14444) );
  AND3_X1 U14516 ( .A1(n14443), .A2(n7777), .A3(b_3_), .ZN(n14439) );
  XNOR2_X1 U14517 ( .A(b_31_), .B(n14191), .ZN(Result_add_31_) );
  INV_X1 U14518 ( .A(a_31_), .ZN(n14191) );
  OR3_X1 U14519 ( .A1(n14445), .A2(n14446), .A3(n7322), .ZN(Result_add_30_) );
  AND2_X1 U14520 ( .A1(n8109), .A2(Result_mul_63_), .ZN(n7322) );
  AND3_X1 U14521 ( .A1(n14447), .A2(n14195), .A3(b_30_), .ZN(n14446) );
  INV_X1 U14522 ( .A(Result_mul_63_), .ZN(n14447) );
  AND2_X1 U14523 ( .A1(n14448), .A2(n7315), .ZN(n14445) );
  INV_X1 U14524 ( .A(b_30_), .ZN(n7315) );
  XNOR2_X1 U14525 ( .A(n14195), .B(Result_mul_63_), .ZN(n14448) );
  INV_X1 U14526 ( .A(a_30_), .ZN(n14195) );
  XOR2_X1 U14527 ( .A(n14449), .B(n14450), .Z(Result_add_2_) );
  OR2_X1 U14528 ( .A1(n14451), .A2(n14452), .ZN(n14450) );
  OR3_X1 U14529 ( .A1(n14453), .A2(n14454), .A3(n14455), .ZN(Result_add_29_)
         );
  INV_X1 U14530 ( .A(n14456), .ZN(n14455) );
  OR2_X1 U14531 ( .A1(n8360), .A2(n14457), .ZN(n14456) );
  AND2_X1 U14532 ( .A1(n14458), .A2(n8110), .ZN(n14454) );
  XNOR2_X1 U14533 ( .A(n14457), .B(a_29_), .ZN(n14458) );
  AND3_X1 U14534 ( .A1(n14457), .A2(n8102), .A3(b_29_), .ZN(n14453) );
  XNOR2_X1 U14535 ( .A(n14459), .B(n14460), .ZN(Result_add_28_) );
  AND2_X1 U14536 ( .A1(n8584), .A2(n14461), .ZN(n14460) );
  OR3_X1 U14537 ( .A1(n14462), .A2(n14463), .A3(n14464), .ZN(Result_add_27_)
         );
  AND2_X1 U14538 ( .A1(n14465), .A2(n14466), .ZN(n14464) );
  AND2_X1 U14539 ( .A1(n14467), .A2(n8575), .ZN(n14463) );
  XNOR2_X1 U14540 ( .A(n8116), .B(n14465), .ZN(n14467) );
  AND3_X1 U14541 ( .A1(n14468), .A2(n8116), .A3(b_27_), .ZN(n14462) );
  XNOR2_X1 U14542 ( .A(n14469), .B(n14470), .ZN(Result_add_26_) );
  AND2_X1 U14543 ( .A1(n9031), .A2(n14471), .ZN(n14470) );
  OR3_X1 U14544 ( .A1(n14472), .A2(n14473), .A3(n14474), .ZN(Result_add_25_)
         );
  AND2_X1 U14545 ( .A1(n14475), .A2(n14476), .ZN(n14474) );
  AND2_X1 U14546 ( .A1(n14477), .A2(n9018), .ZN(n14473) );
  XNOR2_X1 U14547 ( .A(n8126), .B(n14475), .ZN(n14477) );
  AND3_X1 U14548 ( .A1(n14478), .A2(n8126), .A3(b_25_), .ZN(n14472) );
  XNOR2_X1 U14549 ( .A(n14479), .B(n14480), .ZN(Result_add_24_) );
  AND2_X1 U14550 ( .A1(n9511), .A2(n14481), .ZN(n14480) );
  OR3_X1 U14551 ( .A1(n14482), .A2(n14483), .A3(n14484), .ZN(Result_add_23_)
         );
  AND2_X1 U14552 ( .A1(n14485), .A2(n14486), .ZN(n14484) );
  AND2_X1 U14553 ( .A1(n14487), .A2(n7976), .ZN(n14483) );
  XNOR2_X1 U14554 ( .A(n8136), .B(n14485), .ZN(n14487) );
  AND3_X1 U14555 ( .A1(n14488), .A2(n8136), .A3(b_23_), .ZN(n14482) );
  XNOR2_X1 U14556 ( .A(n14489), .B(n14490), .ZN(Result_add_22_) );
  AND2_X1 U14557 ( .A1(n9908), .A2(n14491), .ZN(n14490) );
  INV_X1 U14558 ( .A(n14492), .ZN(n14491) );
  OR3_X1 U14559 ( .A1(n14493), .A2(n14494), .A3(n14495), .ZN(Result_add_21_)
         );
  INV_X1 U14560 ( .A(n14496), .ZN(n14495) );
  OR2_X1 U14561 ( .A1(n14497), .A2(n10193), .ZN(n14496) );
  AND2_X1 U14562 ( .A1(n14498), .A2(n9875), .ZN(n14494) );
  XNOR2_X1 U14563 ( .A(a_21_), .B(n14497), .ZN(n14498) );
  AND3_X1 U14564 ( .A1(n14497), .A2(n8146), .A3(b_21_), .ZN(n14493) );
  XOR2_X1 U14565 ( .A(n14499), .B(n14500), .Z(Result_add_20_) );
  OR2_X1 U14566 ( .A1(n14501), .A2(n14502), .ZN(n14500) );
  OR3_X1 U14567 ( .A1(n14503), .A2(n14504), .A3(n14505), .ZN(Result_add_1_) );
  INV_X1 U14568 ( .A(n14506), .ZN(n14505) );
  OR2_X1 U14569 ( .A1(n14507), .A2(n14314), .ZN(n14506) );
  AND2_X1 U14570 ( .A1(n14508), .A2(n14001), .ZN(n14504) );
  XNOR2_X1 U14571 ( .A(a_1_), .B(n14507), .ZN(n14508) );
  AND3_X1 U14572 ( .A1(n14507), .A2(n7656), .A3(b_1_), .ZN(n14503) );
  OR3_X1 U14573 ( .A1(n14509), .A2(n14510), .A3(n14511), .ZN(Result_add_19_)
         );
  INV_X1 U14574 ( .A(n14512), .ZN(n14511) );
  OR2_X1 U14575 ( .A1(n14513), .A2(n10602), .ZN(n14512) );
  AND2_X1 U14576 ( .A1(n14514), .A2(n7909), .ZN(n14510) );
  XNOR2_X1 U14577 ( .A(a_19_), .B(n14513), .ZN(n14514) );
  AND3_X1 U14578 ( .A1(n14513), .A2(n8156), .A3(b_19_), .ZN(n14509) );
  XOR2_X1 U14579 ( .A(n14515), .B(n14516), .Z(Result_add_18_) );
  OR2_X1 U14580 ( .A1(n14517), .A2(n14518), .ZN(n14516) );
  OR3_X1 U14581 ( .A1(n14519), .A2(n14520), .A3(n14521), .ZN(Result_add_17_)
         );
  INV_X1 U14582 ( .A(n14522), .ZN(n14521) );
  OR2_X1 U14583 ( .A1(n14523), .A2(n10984), .ZN(n14522) );
  AND2_X1 U14584 ( .A1(n14524), .A2(n7852), .ZN(n14520) );
  XNOR2_X1 U14585 ( .A(a_17_), .B(n14523), .ZN(n14524) );
  AND3_X1 U14586 ( .A1(n14523), .A2(n8166), .A3(b_17_), .ZN(n14519) );
  XOR2_X1 U14587 ( .A(n14525), .B(n14526), .Z(Result_add_16_) );
  OR2_X1 U14588 ( .A1(n14527), .A2(n14528), .ZN(n14526) );
  OR3_X1 U14589 ( .A1(n14529), .A2(n14530), .A3(n14531), .ZN(Result_add_15_)
         );
  INV_X1 U14590 ( .A(n14532), .ZN(n14531) );
  OR2_X1 U14591 ( .A1(n14533), .A2(n11386), .ZN(n14532) );
  AND2_X1 U14592 ( .A1(n14534), .A2(n11108), .ZN(n14530) );
  XNOR2_X1 U14593 ( .A(a_15_), .B(n14533), .ZN(n14534) );
  AND3_X1 U14594 ( .A1(n14533), .A2(n8176), .A3(b_15_), .ZN(n14529) );
  XOR2_X1 U14595 ( .A(n14535), .B(n14536), .Z(Result_add_14_) );
  OR2_X1 U14596 ( .A1(n14537), .A2(n14538), .ZN(n14536) );
  OR3_X1 U14597 ( .A1(n14539), .A2(n14540), .A3(n14541), .ZN(Result_add_13_)
         );
  INV_X1 U14598 ( .A(n14542), .ZN(n14541) );
  OR2_X1 U14599 ( .A1(n14543), .A2(n11809), .ZN(n14542) );
  AND2_X1 U14600 ( .A1(n14544), .A2(n11530), .ZN(n14540) );
  XNOR2_X1 U14601 ( .A(a_13_), .B(n14543), .ZN(n14544) );
  AND3_X1 U14602 ( .A1(n14543), .A2(n8186), .A3(b_13_), .ZN(n14539) );
  XOR2_X1 U14603 ( .A(n14545), .B(n14546), .Z(Result_add_12_) );
  OR2_X1 U14604 ( .A1(n14547), .A2(n14548), .ZN(n14546) );
  OR3_X1 U14605 ( .A1(n14549), .A2(n14550), .A3(n14551), .ZN(Result_add_11_)
         );
  INV_X1 U14606 ( .A(n14552), .ZN(n14551) );
  OR2_X1 U14607 ( .A1(n14553), .A2(n12253), .ZN(n14552) );
  AND2_X1 U14608 ( .A1(n14554), .A2(n11958), .ZN(n14550) );
  XNOR2_X1 U14609 ( .A(a_11_), .B(n14553), .ZN(n14554) );
  AND3_X1 U14610 ( .A1(n14553), .A2(n8196), .A3(b_11_), .ZN(n14549) );
  XOR2_X1 U14611 ( .A(n14555), .B(n14556), .Z(Result_add_10_) );
  OR2_X1 U14612 ( .A1(n14557), .A2(n14558), .ZN(n14556) );
  XOR2_X1 U14613 ( .A(n14559), .B(n14560), .Z(Result_add_0_) );
  XNOR2_X1 U14614 ( .A(a_0_), .B(b_0_), .ZN(n14560) );
  OR2_X1 U14615 ( .A1(n14561), .A2(n14562), .ZN(n14559) );
  AND2_X1 U14616 ( .A1(n7656), .A2(n14001), .ZN(n14562) );
  AND2_X1 U14617 ( .A1(n14507), .A2(n14314), .ZN(n14561) );
  OR2_X1 U14618 ( .A1(n14001), .A2(n7656), .ZN(n14314) );
  INV_X1 U14619 ( .A(a_1_), .ZN(n7656) );
  INV_X1 U14620 ( .A(b_1_), .ZN(n14001) );
  OR2_X1 U14621 ( .A1(n14563), .A2(n14451), .ZN(n14507) );
  AND2_X1 U14622 ( .A1(n7689), .A2(n13831), .ZN(n14451) );
  INV_X1 U14623 ( .A(b_2_), .ZN(n13831) );
  INV_X1 U14624 ( .A(a_2_), .ZN(n7689) );
  AND2_X1 U14625 ( .A1(n14449), .A2(n7665), .ZN(n14563) );
  INV_X1 U14626 ( .A(n14452), .ZN(n7665) );
  AND2_X1 U14627 ( .A1(b_2_), .A2(a_2_), .ZN(n14452) );
  OR2_X1 U14628 ( .A1(n14564), .A2(n14565), .ZN(n14449) );
  AND2_X1 U14629 ( .A1(n7777), .A2(n7620), .ZN(n14565) );
  AND2_X1 U14630 ( .A1(n14443), .A2(n7695), .ZN(n14564) );
  OR2_X1 U14631 ( .A1(n7620), .A2(n7777), .ZN(n7695) );
  INV_X1 U14632 ( .A(a_3_), .ZN(n7777) );
  OR2_X1 U14633 ( .A1(n14566), .A2(n14437), .ZN(n14443) );
  AND2_X1 U14634 ( .A1(n7785), .A2(n7648), .ZN(n14437) );
  INV_X1 U14635 ( .A(b_4_), .ZN(n7648) );
  INV_X1 U14636 ( .A(a_4_), .ZN(n7785) );
  AND2_X1 U14637 ( .A1(n14435), .A2(n7783), .ZN(n14566) );
  INV_X1 U14638 ( .A(n14438), .ZN(n7783) );
  AND2_X1 U14639 ( .A1(b_4_), .A2(a_4_), .ZN(n14438) );
  OR2_X1 U14640 ( .A1(n14567), .A2(n14568), .ZN(n14435) );
  AND2_X1 U14641 ( .A1(n8226), .A2(n7674), .ZN(n14568) );
  AND2_X1 U14642 ( .A1(n14433), .A2(n13547), .ZN(n14567) );
  OR2_X1 U14643 ( .A1(n7674), .A2(n8226), .ZN(n13547) );
  INV_X1 U14644 ( .A(a_5_), .ZN(n8226) );
  OR2_X1 U14645 ( .A1(n14569), .A2(n14427), .ZN(n14433) );
  AND2_X1 U14646 ( .A1(n8221), .A2(n7716), .ZN(n14427) );
  INV_X1 U14647 ( .A(b_6_), .ZN(n7716) );
  INV_X1 U14648 ( .A(a_6_), .ZN(n8221) );
  AND2_X1 U14649 ( .A1(n14425), .A2(n13346), .ZN(n14569) );
  INV_X1 U14650 ( .A(n14428), .ZN(n13346) );
  AND2_X1 U14651 ( .A1(b_6_), .A2(a_6_), .ZN(n14428) );
  OR2_X1 U14652 ( .A1(n14570), .A2(n14571), .ZN(n14425) );
  AND2_X1 U14653 ( .A1(n8216), .A2(n7755), .ZN(n14571) );
  AND2_X1 U14654 ( .A1(n14423), .A2(n13138), .ZN(n14570) );
  OR2_X1 U14655 ( .A1(n7755), .A2(n8216), .ZN(n13138) );
  INV_X1 U14656 ( .A(a_7_), .ZN(n8216) );
  OR2_X1 U14657 ( .A1(n14572), .A2(n14417), .ZN(n14423) );
  AND2_X1 U14658 ( .A1(n8211), .A2(n12612), .ZN(n14417) );
  INV_X1 U14659 ( .A(b_8_), .ZN(n12612) );
  INV_X1 U14660 ( .A(a_8_), .ZN(n8211) );
  AND2_X1 U14661 ( .A1(n14415), .A2(n12923), .ZN(n14572) );
  INV_X1 U14662 ( .A(n14418), .ZN(n12923) );
  AND2_X1 U14663 ( .A1(b_8_), .A2(a_8_), .ZN(n14418) );
  OR2_X1 U14664 ( .A1(n14573), .A2(n14574), .ZN(n14415) );
  AND2_X1 U14665 ( .A1(n8206), .A2(n12396), .ZN(n14574) );
  AND2_X1 U14666 ( .A1(n14413), .A2(n12697), .ZN(n14573) );
  OR2_X1 U14667 ( .A1(n12396), .A2(n8206), .ZN(n12697) );
  INV_X1 U14668 ( .A(a_9_), .ZN(n8206) );
  OR2_X1 U14669 ( .A1(n14575), .A2(n14557), .ZN(n14413) );
  AND2_X1 U14670 ( .A1(n8201), .A2(n12176), .ZN(n14557) );
  INV_X1 U14671 ( .A(b_10_), .ZN(n12176) );
  INV_X1 U14672 ( .A(a_10_), .ZN(n8201) );
  AND2_X1 U14673 ( .A1(n14555), .A2(n12475), .ZN(n14575) );
  INV_X1 U14674 ( .A(n14558), .ZN(n12475) );
  AND2_X1 U14675 ( .A1(b_10_), .A2(a_10_), .ZN(n14558) );
  OR2_X1 U14676 ( .A1(n14576), .A2(n14577), .ZN(n14555) );
  AND2_X1 U14677 ( .A1(n8196), .A2(n11958), .ZN(n14577) );
  AND2_X1 U14678 ( .A1(n14553), .A2(n12253), .ZN(n14576) );
  OR2_X1 U14679 ( .A1(n11958), .A2(n8196), .ZN(n12253) );
  INV_X1 U14680 ( .A(a_11_), .ZN(n8196) );
  OR2_X1 U14681 ( .A1(n14578), .A2(n14547), .ZN(n14553) );
  AND2_X1 U14682 ( .A1(n8191), .A2(n11740), .ZN(n14547) );
  INV_X1 U14683 ( .A(b_12_), .ZN(n11740) );
  INV_X1 U14684 ( .A(a_12_), .ZN(n8191) );
  AND2_X1 U14685 ( .A1(n14545), .A2(n12031), .ZN(n14578) );
  INV_X1 U14686 ( .A(n14548), .ZN(n12031) );
  AND2_X1 U14687 ( .A1(b_12_), .A2(a_12_), .ZN(n14548) );
  OR2_X1 U14688 ( .A1(n14579), .A2(n14580), .ZN(n14545) );
  AND2_X1 U14689 ( .A1(n8186), .A2(n11530), .ZN(n14580) );
  AND2_X1 U14690 ( .A1(n14543), .A2(n11809), .ZN(n14579) );
  OR2_X1 U14691 ( .A1(n11530), .A2(n8186), .ZN(n11809) );
  INV_X1 U14692 ( .A(a_13_), .ZN(n8186) );
  OR2_X1 U14693 ( .A1(n14581), .A2(n14537), .ZN(n14543) );
  AND2_X1 U14694 ( .A1(n8181), .A2(n11329), .ZN(n14537) );
  INV_X1 U14695 ( .A(b_14_), .ZN(n11329) );
  INV_X1 U14696 ( .A(a_14_), .ZN(n8181) );
  AND2_X1 U14697 ( .A1(n14535), .A2(n11595), .ZN(n14581) );
  INV_X1 U14698 ( .A(n14538), .ZN(n11595) );
  AND2_X1 U14699 ( .A1(b_14_), .A2(a_14_), .ZN(n14538) );
  OR2_X1 U14700 ( .A1(n14582), .A2(n14583), .ZN(n14535) );
  AND2_X1 U14701 ( .A1(n8176), .A2(n11108), .ZN(n14583) );
  AND2_X1 U14702 ( .A1(n14533), .A2(n11386), .ZN(n14582) );
  OR2_X1 U14703 ( .A1(n11108), .A2(n8176), .ZN(n11386) );
  INV_X1 U14704 ( .A(a_15_), .ZN(n8176) );
  OR2_X1 U14705 ( .A1(n14584), .A2(n14527), .ZN(n14533) );
  AND2_X1 U14706 ( .A1(n8171), .A2(n10931), .ZN(n14527) );
  INV_X1 U14707 ( .A(b_16_), .ZN(n10931) );
  INV_X1 U14708 ( .A(a_16_), .ZN(n8171) );
  AND2_X1 U14709 ( .A1(n14525), .A2(n11165), .ZN(n14584) );
  INV_X1 U14710 ( .A(n14528), .ZN(n11165) );
  AND2_X1 U14711 ( .A1(b_16_), .A2(a_16_), .ZN(n14528) );
  OR2_X1 U14712 ( .A1(n14585), .A2(n14586), .ZN(n14525) );
  AND2_X1 U14713 ( .A1(n8166), .A2(n7852), .ZN(n14586) );
  AND2_X1 U14714 ( .A1(n14523), .A2(n10984), .ZN(n14585) );
  OR2_X1 U14715 ( .A1(n8166), .A2(n7852), .ZN(n10984) );
  INV_X1 U14716 ( .A(a_17_), .ZN(n8166) );
  OR2_X1 U14717 ( .A1(n14587), .A2(n14517), .ZN(n14523) );
  AND2_X1 U14718 ( .A1(n8161), .A2(n7877), .ZN(n14517) );
  INV_X1 U14719 ( .A(b_18_), .ZN(n7877) );
  INV_X1 U14720 ( .A(a_18_), .ZN(n8161) );
  AND2_X1 U14721 ( .A1(n14515), .A2(n10796), .ZN(n14587) );
  INV_X1 U14722 ( .A(n14518), .ZN(n10796) );
  AND2_X1 U14723 ( .A1(a_18_), .A2(b_18_), .ZN(n14518) );
  OR2_X1 U14724 ( .A1(n14588), .A2(n14589), .ZN(n14515) );
  AND2_X1 U14725 ( .A1(n8156), .A2(n7909), .ZN(n14589) );
  AND2_X1 U14726 ( .A1(n14513), .A2(n10602), .ZN(n14588) );
  OR2_X1 U14727 ( .A1(n8156), .A2(n7909), .ZN(n10602) );
  INV_X1 U14728 ( .A(a_19_), .ZN(n8156) );
  OR2_X1 U14729 ( .A1(n14590), .A2(n14501), .ZN(n14513) );
  AND2_X1 U14730 ( .A1(n8151), .A2(n9990), .ZN(n14501) );
  INV_X1 U14731 ( .A(b_20_), .ZN(n9990) );
  INV_X1 U14732 ( .A(a_20_), .ZN(n8151) );
  AND2_X1 U14733 ( .A1(n14499), .A2(n10401), .ZN(n14590) );
  INV_X1 U14734 ( .A(n14502), .ZN(n10401) );
  AND2_X1 U14735 ( .A1(a_20_), .A2(b_20_), .ZN(n14502) );
  OR2_X1 U14736 ( .A1(n14591), .A2(n14592), .ZN(n14499) );
  AND2_X1 U14737 ( .A1(n8146), .A2(n9875), .ZN(n14592) );
  AND2_X1 U14738 ( .A1(n14497), .A2(n10193), .ZN(n14591) );
  OR2_X1 U14739 ( .A1(n8146), .A2(n9875), .ZN(n10193) );
  INV_X1 U14740 ( .A(a_21_), .ZN(n8146) );
  OR2_X1 U14741 ( .A1(n14593), .A2(n14492), .ZN(n14497) );
  AND2_X1 U14742 ( .A1(n8141), .A2(n9684), .ZN(n14492) );
  AND2_X1 U14743 ( .A1(n14489), .A2(n9908), .ZN(n14593) );
  OR2_X1 U14744 ( .A1(n8141), .A2(n9684), .ZN(n9908) );
  INV_X1 U14745 ( .A(b_22_), .ZN(n9684) );
  INV_X1 U14746 ( .A(a_22_), .ZN(n8141) );
  OR2_X1 U14747 ( .A1(n14594), .A2(n14595), .ZN(n14489) );
  AND2_X1 U14748 ( .A1(n8136), .A2(n7976), .ZN(n14595) );
  INV_X1 U14749 ( .A(b_23_), .ZN(n7976) );
  INV_X1 U14750 ( .A(a_23_), .ZN(n8136) );
  AND2_X1 U14751 ( .A1(n14488), .A2(n9713), .ZN(n14594) );
  INV_X1 U14752 ( .A(n14486), .ZN(n9713) );
  AND2_X1 U14753 ( .A1(a_23_), .A2(b_23_), .ZN(n14486) );
  INV_X1 U14754 ( .A(n14485), .ZN(n14488) );
  AND2_X1 U14755 ( .A1(n14596), .A2(n14481), .ZN(n14485) );
  OR2_X1 U14756 ( .A1(a_24_), .A2(b_24_), .ZN(n14481) );
  INV_X1 U14757 ( .A(n14597), .ZN(n14596) );
  AND2_X1 U14758 ( .A1(n14479), .A2(n9511), .ZN(n14597) );
  OR2_X1 U14759 ( .A1(n8131), .A2(n9145), .ZN(n9511) );
  INV_X1 U14760 ( .A(b_24_), .ZN(n9145) );
  INV_X1 U14761 ( .A(a_24_), .ZN(n8131) );
  OR2_X1 U14762 ( .A1(n14598), .A2(n14599), .ZN(n14479) );
  AND2_X1 U14763 ( .A1(n8126), .A2(n9018), .ZN(n14599) );
  INV_X1 U14764 ( .A(b_25_), .ZN(n9018) );
  INV_X1 U14765 ( .A(a_25_), .ZN(n8126) );
  AND2_X1 U14766 ( .A1(n14478), .A2(n9303), .ZN(n14598) );
  INV_X1 U14767 ( .A(n14476), .ZN(n9303) );
  AND2_X1 U14768 ( .A1(a_25_), .A2(b_25_), .ZN(n14476) );
  INV_X1 U14769 ( .A(n14475), .ZN(n14478) );
  AND2_X1 U14770 ( .A1(n14600), .A2(n14471), .ZN(n14475) );
  OR2_X1 U14771 ( .A1(a_26_), .A2(b_26_), .ZN(n14471) );
  INV_X1 U14772 ( .A(n14601), .ZN(n14600) );
  AND2_X1 U14773 ( .A1(n14469), .A2(n9031), .ZN(n14601) );
  OR2_X1 U14774 ( .A1(n8121), .A2(n8802), .ZN(n9031) );
  INV_X1 U14775 ( .A(b_26_), .ZN(n8802) );
  INV_X1 U14776 ( .A(a_26_), .ZN(n8121) );
  OR2_X1 U14777 ( .A1(n14602), .A2(n14603), .ZN(n14469) );
  AND2_X1 U14778 ( .A1(n8116), .A2(n8575), .ZN(n14603) );
  INV_X1 U14779 ( .A(b_27_), .ZN(n8575) );
  INV_X1 U14780 ( .A(a_27_), .ZN(n8116) );
  AND2_X1 U14781 ( .A1(n14468), .A2(n8811), .ZN(n14602) );
  INV_X1 U14782 ( .A(n14466), .ZN(n8811) );
  AND2_X1 U14783 ( .A1(a_27_), .A2(b_27_), .ZN(n14466) );
  INV_X1 U14784 ( .A(n14465), .ZN(n14468) );
  AND2_X1 U14785 ( .A1(n14604), .A2(n14461), .ZN(n14465) );
  OR2_X1 U14786 ( .A1(a_28_), .A2(b_28_), .ZN(n14461) );
  INV_X1 U14787 ( .A(n14605), .ZN(n14604) );
  AND2_X1 U14788 ( .A1(n14459), .A2(n8584), .ZN(n14605) );
  OR2_X1 U14789 ( .A1(n8111), .A2(n8355), .ZN(n8584) );
  INV_X1 U14790 ( .A(b_28_), .ZN(n8355) );
  INV_X1 U14791 ( .A(a_28_), .ZN(n8111) );
  OR2_X1 U14792 ( .A1(n14606), .A2(n14607), .ZN(n14459) );
  AND2_X1 U14793 ( .A1(n8102), .A2(n8110), .ZN(n14607) );
  AND2_X1 U14794 ( .A1(n14457), .A2(n8360), .ZN(n14606) );
  OR2_X1 U14795 ( .A1(n8102), .A2(n8110), .ZN(n8360) );
  INV_X1 U14796 ( .A(a_29_), .ZN(n8102) );
  INV_X1 U14797 ( .A(n14608), .ZN(n14457) );
  OR2_X1 U14798 ( .A1(n14609), .A2(n8109), .ZN(n14608) );
  AND2_X1 U14799 ( .A1(a_30_), .A2(b_30_), .ZN(n8109) );
  AND2_X1 U14800 ( .A1(Result_mul_63_), .A2(n14610), .ZN(n14609) );
  OR2_X1 U14801 ( .A1(a_30_), .A2(b_30_), .ZN(n14610) );
  AND2_X1 U14802 ( .A1(a_31_), .A2(b_31_), .ZN(Result_mul_63_) );
endmodule

