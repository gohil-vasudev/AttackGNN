module add_mul_comp_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, 
        a_17_, a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, 
        a_27_, a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, 
        b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, 
        b_16_, b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, 
        b_26_, b_27_, b_28_, b_29_, b_30_, b_31_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, 
        Result_32_, Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, 
        Result_38_, Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, 
        Result_44_, Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, 
        Result_50_, Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, 
        Result_56_, Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, 
        Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   Result_9_, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_31_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_28_ = Result_9_;
  assign Result_26_ = Result_9_;
  assign Result_24_ = Result_9_;
  assign Result_22_ = Result_9_;
  assign Result_20_ = Result_9_;
  assign Result_19_ = Result_9_;
  assign Result_17_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_16_ = Result_9_;
  assign Result_18_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_21_ = Result_9_;
  assign Result_23_ = Result_9_;
  assign Result_25_ = Result_9_;
  assign Result_27_ = Result_9_;
  assign Result_29_ = Result_9_;
  assign Result_30_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  NAND2_X2 U564 ( .A1(n930), .A2(n931), .ZN(Result_9_) );
  INV_X2 U565 ( .A(n544), .ZN(n539) );
  XNOR2_X1 U566 ( .A(n531), .B(a_31_), .ZN(Result_63_) );
  NAND2_X1 U567 ( .A1(n532), .A2(n533), .ZN(Result_62_) );
  NAND4_X1 U568 ( .A1(n534), .A2(a_31_), .A3(n535), .A4(n536), .ZN(n533) );
  NOR2_X1 U569 ( .A1(n537), .A2(n538), .ZN(n534) );
  NOR2_X1 U570 ( .A1(b_31_), .A2(Result_9_), .ZN(n538) );
  NOR2_X1 U571 ( .A1(n539), .A2(n531), .ZN(n537) );
  NAND3_X1 U572 ( .A1(n540), .A2(n541), .A3(n542), .ZN(n532) );
  XNOR2_X1 U573 ( .A(b_30_), .B(n543), .ZN(n542) );
  NAND3_X1 U574 ( .A1(n544), .A2(n531), .A3(a_31_), .ZN(n541) );
  NAND2_X1 U575 ( .A1(n545), .A2(n546), .ZN(n540) );
  NAND2_X1 U576 ( .A1(n547), .A2(n548), .ZN(Result_61_) );
  NAND2_X1 U577 ( .A1(n539), .A2(n549), .ZN(n548) );
  XOR2_X1 U578 ( .A(n550), .B(n551), .Z(n549) );
  NAND2_X1 U579 ( .A1(n552), .A2(Result_9_), .ZN(n547) );
  XNOR2_X1 U580 ( .A(n553), .B(n550), .ZN(n552) );
  NAND2_X1 U581 ( .A1(n554), .A2(n555), .ZN(n550) );
  NAND2_X1 U582 ( .A1(n556), .A2(n557), .ZN(Result_60_) );
  NAND2_X1 U583 ( .A1(n539), .A2(n558), .ZN(n557) );
  XNOR2_X1 U584 ( .A(n559), .B(n560), .ZN(n558) );
  NAND2_X1 U585 ( .A1(n561), .A2(Result_9_), .ZN(n556) );
  XOR2_X1 U586 ( .A(n562), .B(n559), .Z(n561) );
  AND2_X1 U587 ( .A1(n563), .A2(n564), .ZN(n559) );
  NAND2_X1 U588 ( .A1(n565), .A2(n566), .ZN(Result_59_) );
  NAND2_X1 U589 ( .A1(n539), .A2(n567), .ZN(n566) );
  XOR2_X1 U590 ( .A(n568), .B(n569), .Z(n567) );
  NAND2_X1 U591 ( .A1(n570), .A2(Result_9_), .ZN(n565) );
  XNOR2_X1 U592 ( .A(n571), .B(n568), .ZN(n570) );
  NAND2_X1 U593 ( .A1(n572), .A2(n573), .ZN(n568) );
  NAND2_X1 U594 ( .A1(n574), .A2(n575), .ZN(Result_58_) );
  NAND2_X1 U595 ( .A1(n539), .A2(n576), .ZN(n575) );
  XNOR2_X1 U596 ( .A(n577), .B(n578), .ZN(n576) );
  NAND2_X1 U597 ( .A1(n579), .A2(Result_9_), .ZN(n574) );
  XOR2_X1 U598 ( .A(n580), .B(n577), .Z(n579) );
  AND2_X1 U599 ( .A1(n581), .A2(n582), .ZN(n577) );
  NAND2_X1 U600 ( .A1(n583), .A2(n584), .ZN(Result_57_) );
  NAND2_X1 U601 ( .A1(n539), .A2(n585), .ZN(n584) );
  XOR2_X1 U602 ( .A(n586), .B(n587), .Z(n585) );
  NAND2_X1 U603 ( .A1(n588), .A2(Result_9_), .ZN(n583) );
  XNOR2_X1 U604 ( .A(n589), .B(n586), .ZN(n588) );
  NAND2_X1 U605 ( .A1(n590), .A2(n591), .ZN(n586) );
  NAND2_X1 U606 ( .A1(n592), .A2(n593), .ZN(Result_56_) );
  NAND2_X1 U607 ( .A1(n539), .A2(n594), .ZN(n593) );
  XNOR2_X1 U608 ( .A(n595), .B(n596), .ZN(n594) );
  NAND2_X1 U609 ( .A1(n597), .A2(Result_9_), .ZN(n592) );
  XOR2_X1 U610 ( .A(n598), .B(n595), .Z(n597) );
  AND2_X1 U611 ( .A1(n599), .A2(n600), .ZN(n595) );
  NAND2_X1 U612 ( .A1(n601), .A2(n602), .ZN(Result_55_) );
  NAND2_X1 U613 ( .A1(n539), .A2(n603), .ZN(n602) );
  XOR2_X1 U614 ( .A(n604), .B(n605), .Z(n603) );
  NAND2_X1 U615 ( .A1(n606), .A2(Result_9_), .ZN(n601) );
  XNOR2_X1 U616 ( .A(n607), .B(n604), .ZN(n606) );
  NAND2_X1 U617 ( .A1(n608), .A2(n609), .ZN(n604) );
  NAND2_X1 U618 ( .A1(n610), .A2(n611), .ZN(Result_54_) );
  NAND2_X1 U619 ( .A1(n539), .A2(n612), .ZN(n611) );
  XNOR2_X1 U620 ( .A(n613), .B(n614), .ZN(n612) );
  NAND2_X1 U621 ( .A1(n615), .A2(Result_9_), .ZN(n610) );
  XOR2_X1 U622 ( .A(n616), .B(n613), .Z(n615) );
  AND2_X1 U623 ( .A1(n617), .A2(n618), .ZN(n613) );
  NAND2_X1 U624 ( .A1(n619), .A2(n620), .ZN(Result_53_) );
  NAND2_X1 U625 ( .A1(n539), .A2(n621), .ZN(n620) );
  XOR2_X1 U626 ( .A(n622), .B(n623), .Z(n621) );
  NAND2_X1 U627 ( .A1(n624), .A2(Result_9_), .ZN(n619) );
  XNOR2_X1 U628 ( .A(n625), .B(n622), .ZN(n624) );
  NAND2_X1 U629 ( .A1(n626), .A2(n627), .ZN(n622) );
  NAND2_X1 U630 ( .A1(n628), .A2(n629), .ZN(Result_52_) );
  NAND2_X1 U631 ( .A1(n539), .A2(n630), .ZN(n629) );
  XNOR2_X1 U632 ( .A(n631), .B(n632), .ZN(n630) );
  NAND2_X1 U633 ( .A1(n633), .A2(Result_9_), .ZN(n628) );
  XOR2_X1 U634 ( .A(n634), .B(n631), .Z(n633) );
  AND2_X1 U635 ( .A1(n635), .A2(n636), .ZN(n631) );
  NAND2_X1 U636 ( .A1(n637), .A2(n638), .ZN(Result_51_) );
  NAND2_X1 U637 ( .A1(n539), .A2(n639), .ZN(n638) );
  XOR2_X1 U638 ( .A(n640), .B(n641), .Z(n639) );
  NAND2_X1 U639 ( .A1(n642), .A2(Result_9_), .ZN(n637) );
  XNOR2_X1 U640 ( .A(n643), .B(n640), .ZN(n642) );
  NAND2_X1 U641 ( .A1(n644), .A2(n645), .ZN(n640) );
  NAND2_X1 U642 ( .A1(n646), .A2(n647), .ZN(Result_50_) );
  NAND2_X1 U643 ( .A1(n539), .A2(n648), .ZN(n647) );
  XNOR2_X1 U644 ( .A(n649), .B(n650), .ZN(n648) );
  NAND2_X1 U645 ( .A1(n651), .A2(Result_9_), .ZN(n646) );
  XOR2_X1 U646 ( .A(n652), .B(n649), .Z(n651) );
  AND2_X1 U647 ( .A1(n653), .A2(n654), .ZN(n649) );
  NAND2_X1 U648 ( .A1(n655), .A2(n656), .ZN(Result_49_) );
  NAND2_X1 U649 ( .A1(n539), .A2(n657), .ZN(n656) );
  XOR2_X1 U650 ( .A(n658), .B(n659), .Z(n657) );
  NAND2_X1 U651 ( .A1(n660), .A2(Result_9_), .ZN(n655) );
  XNOR2_X1 U652 ( .A(n661), .B(n658), .ZN(n660) );
  NAND2_X1 U653 ( .A1(n662), .A2(n663), .ZN(n658) );
  NAND2_X1 U654 ( .A1(n664), .A2(n665), .ZN(Result_48_) );
  NAND2_X1 U655 ( .A1(n539), .A2(n666), .ZN(n665) );
  XNOR2_X1 U656 ( .A(n667), .B(n668), .ZN(n666) );
  NAND2_X1 U657 ( .A1(n669), .A2(Result_9_), .ZN(n664) );
  XOR2_X1 U658 ( .A(n670), .B(n667), .Z(n669) );
  AND2_X1 U659 ( .A1(n671), .A2(n672), .ZN(n667) );
  NAND2_X1 U660 ( .A1(n673), .A2(n674), .ZN(Result_47_) );
  NAND2_X1 U661 ( .A1(n539), .A2(n675), .ZN(n674) );
  XOR2_X1 U662 ( .A(n676), .B(n677), .Z(n675) );
  NAND2_X1 U663 ( .A1(n678), .A2(Result_9_), .ZN(n673) );
  XNOR2_X1 U664 ( .A(n679), .B(n676), .ZN(n678) );
  NAND2_X1 U665 ( .A1(n680), .A2(n681), .ZN(n676) );
  NAND2_X1 U666 ( .A1(n682), .A2(n683), .ZN(Result_46_) );
  NAND2_X1 U667 ( .A1(n539), .A2(n684), .ZN(n683) );
  XNOR2_X1 U668 ( .A(n685), .B(n686), .ZN(n684) );
  NAND2_X1 U669 ( .A1(n687), .A2(Result_9_), .ZN(n682) );
  XOR2_X1 U670 ( .A(n688), .B(n685), .Z(n687) );
  AND2_X1 U671 ( .A1(n689), .A2(n690), .ZN(n685) );
  NAND2_X1 U672 ( .A1(n691), .A2(n692), .ZN(Result_45_) );
  NAND2_X1 U673 ( .A1(n539), .A2(n693), .ZN(n692) );
  XOR2_X1 U674 ( .A(n694), .B(n695), .Z(n693) );
  NAND2_X1 U675 ( .A1(n696), .A2(Result_9_), .ZN(n691) );
  XNOR2_X1 U676 ( .A(n697), .B(n694), .ZN(n696) );
  NAND2_X1 U677 ( .A1(n698), .A2(n699), .ZN(n694) );
  NAND2_X1 U678 ( .A1(n700), .A2(n701), .ZN(Result_44_) );
  NAND2_X1 U679 ( .A1(n539), .A2(n702), .ZN(n701) );
  XNOR2_X1 U680 ( .A(n703), .B(n704), .ZN(n702) );
  NAND2_X1 U681 ( .A1(n705), .A2(Result_9_), .ZN(n700) );
  XOR2_X1 U682 ( .A(n706), .B(n703), .Z(n705) );
  AND2_X1 U683 ( .A1(n707), .A2(n708), .ZN(n703) );
  NAND2_X1 U684 ( .A1(n709), .A2(n710), .ZN(Result_43_) );
  NAND2_X1 U685 ( .A1(n539), .A2(n711), .ZN(n710) );
  XOR2_X1 U686 ( .A(n712), .B(n713), .Z(n711) );
  NAND2_X1 U687 ( .A1(n714), .A2(Result_9_), .ZN(n709) );
  XNOR2_X1 U688 ( .A(n715), .B(n712), .ZN(n714) );
  NAND2_X1 U689 ( .A1(n716), .A2(n717), .ZN(n712) );
  NAND2_X1 U690 ( .A1(n718), .A2(n719), .ZN(Result_42_) );
  NAND2_X1 U691 ( .A1(n539), .A2(n720), .ZN(n719) );
  XNOR2_X1 U692 ( .A(n721), .B(n722), .ZN(n720) );
  NAND2_X1 U693 ( .A1(n723), .A2(Result_9_), .ZN(n718) );
  XOR2_X1 U694 ( .A(n724), .B(n721), .Z(n723) );
  AND2_X1 U695 ( .A1(n725), .A2(n726), .ZN(n721) );
  NAND2_X1 U696 ( .A1(n727), .A2(n728), .ZN(Result_41_) );
  NAND2_X1 U697 ( .A1(n539), .A2(n729), .ZN(n728) );
  XOR2_X1 U698 ( .A(n730), .B(n731), .Z(n729) );
  NAND2_X1 U699 ( .A1(n732), .A2(Result_9_), .ZN(n727) );
  XNOR2_X1 U700 ( .A(n733), .B(n730), .ZN(n732) );
  NAND2_X1 U701 ( .A1(n734), .A2(n735), .ZN(n730) );
  NAND2_X1 U702 ( .A1(n736), .A2(n737), .ZN(Result_40_) );
  NAND2_X1 U703 ( .A1(n539), .A2(n738), .ZN(n737) );
  XNOR2_X1 U704 ( .A(n739), .B(n740), .ZN(n738) );
  NAND2_X1 U705 ( .A1(n741), .A2(Result_9_), .ZN(n736) );
  XOR2_X1 U706 ( .A(n742), .B(n739), .Z(n741) );
  AND2_X1 U707 ( .A1(n743), .A2(n744), .ZN(n739) );
  NAND2_X1 U708 ( .A1(n745), .A2(n746), .ZN(Result_39_) );
  NAND2_X1 U709 ( .A1(n539), .A2(n747), .ZN(n746) );
  XOR2_X1 U710 ( .A(n748), .B(n749), .Z(n747) );
  NAND2_X1 U711 ( .A1(n750), .A2(Result_9_), .ZN(n745) );
  XNOR2_X1 U712 ( .A(n751), .B(n748), .ZN(n750) );
  NAND2_X1 U713 ( .A1(n752), .A2(n753), .ZN(n748) );
  NAND2_X1 U714 ( .A1(n754), .A2(n755), .ZN(Result_38_) );
  NAND2_X1 U715 ( .A1(n539), .A2(n756), .ZN(n755) );
  XNOR2_X1 U716 ( .A(n757), .B(n758), .ZN(n756) );
  NAND2_X1 U717 ( .A1(n759), .A2(Result_9_), .ZN(n754) );
  XOR2_X1 U718 ( .A(n760), .B(n757), .Z(n759) );
  AND2_X1 U719 ( .A1(n761), .A2(n762), .ZN(n757) );
  NAND2_X1 U720 ( .A1(n763), .A2(n764), .ZN(Result_37_) );
  NAND2_X1 U721 ( .A1(n539), .A2(n765), .ZN(n764) );
  XOR2_X1 U722 ( .A(n766), .B(n767), .Z(n765) );
  NAND2_X1 U723 ( .A1(n768), .A2(Result_9_), .ZN(n763) );
  XNOR2_X1 U724 ( .A(n769), .B(n766), .ZN(n768) );
  NAND2_X1 U725 ( .A1(n770), .A2(n771), .ZN(n766) );
  NAND2_X1 U726 ( .A1(n772), .A2(n773), .ZN(Result_36_) );
  NAND2_X1 U727 ( .A1(n539), .A2(n774), .ZN(n773) );
  XNOR2_X1 U728 ( .A(n775), .B(n776), .ZN(n774) );
  NAND2_X1 U729 ( .A1(n777), .A2(Result_9_), .ZN(n772) );
  XOR2_X1 U730 ( .A(n778), .B(n775), .Z(n777) );
  AND2_X1 U731 ( .A1(n779), .A2(n780), .ZN(n775) );
  NAND2_X1 U732 ( .A1(n781), .A2(n782), .ZN(Result_35_) );
  NAND2_X1 U733 ( .A1(n539), .A2(n783), .ZN(n782) );
  XOR2_X1 U734 ( .A(n784), .B(n785), .Z(n783) );
  NAND2_X1 U735 ( .A1(n786), .A2(Result_9_), .ZN(n781) );
  XNOR2_X1 U736 ( .A(n787), .B(n784), .ZN(n786) );
  NAND2_X1 U737 ( .A1(n788), .A2(n789), .ZN(n784) );
  NAND2_X1 U738 ( .A1(n790), .A2(n791), .ZN(Result_34_) );
  NAND2_X1 U739 ( .A1(n539), .A2(n792), .ZN(n791) );
  XNOR2_X1 U740 ( .A(n793), .B(n794), .ZN(n792) );
  NAND2_X1 U741 ( .A1(n795), .A2(Result_9_), .ZN(n790) );
  XOR2_X1 U742 ( .A(n796), .B(n793), .Z(n795) );
  AND2_X1 U743 ( .A1(n797), .A2(n798), .ZN(n793) );
  NAND2_X1 U744 ( .A1(n799), .A2(n800), .ZN(Result_33_) );
  NAND2_X1 U745 ( .A1(n539), .A2(n801), .ZN(n800) );
  XOR2_X1 U746 ( .A(n802), .B(n803), .Z(n801) );
  NAND2_X1 U747 ( .A1(n804), .A2(Result_9_), .ZN(n799) );
  XNOR2_X1 U748 ( .A(n805), .B(n802), .ZN(n804) );
  NAND2_X1 U749 ( .A1(n806), .A2(n807), .ZN(n802) );
  NAND2_X1 U750 ( .A1(n808), .A2(n809), .ZN(Result_32_) );
  NAND2_X1 U751 ( .A1(n539), .A2(n810), .ZN(n809) );
  XNOR2_X1 U752 ( .A(n811), .B(n812), .ZN(n810) );
  NOR2_X1 U753 ( .A1(n813), .A2(n814), .ZN(n812) );
  AND2_X1 U754 ( .A1(n803), .A2(a_1_), .ZN(n814) );
  NOR2_X1 U755 ( .A1(n815), .A2(n816), .ZN(n813) );
  NOR2_X1 U756 ( .A1(a_1_), .A2(n803), .ZN(n815) );
  NAND2_X1 U757 ( .A1(n817), .A2(n818), .ZN(n803) );
  NAND2_X1 U758 ( .A1(b_2_), .A2(n819), .ZN(n818) );
  OR2_X1 U759 ( .A1(n794), .A2(a_2_), .ZN(n819) );
  NAND2_X1 U760 ( .A1(a_2_), .A2(n794), .ZN(n817) );
  NAND2_X1 U761 ( .A1(n820), .A2(n821), .ZN(n794) );
  NAND2_X1 U762 ( .A1(b_3_), .A2(n822), .ZN(n821) );
  OR2_X1 U763 ( .A1(n785), .A2(a_3_), .ZN(n822) );
  NAND2_X1 U764 ( .A1(a_3_), .A2(n785), .ZN(n820) );
  NAND2_X1 U765 ( .A1(n823), .A2(n824), .ZN(n785) );
  NAND2_X1 U766 ( .A1(b_4_), .A2(n825), .ZN(n824) );
  OR2_X1 U767 ( .A1(n776), .A2(a_4_), .ZN(n825) );
  NAND2_X1 U768 ( .A1(a_4_), .A2(n776), .ZN(n823) );
  NAND2_X1 U769 ( .A1(n826), .A2(n827), .ZN(n776) );
  NAND2_X1 U770 ( .A1(b_5_), .A2(n828), .ZN(n827) );
  OR2_X1 U771 ( .A1(n767), .A2(a_5_), .ZN(n828) );
  NAND2_X1 U772 ( .A1(a_5_), .A2(n767), .ZN(n826) );
  NAND2_X1 U773 ( .A1(n829), .A2(n830), .ZN(n767) );
  NAND2_X1 U774 ( .A1(b_6_), .A2(n831), .ZN(n830) );
  OR2_X1 U775 ( .A1(n758), .A2(a_6_), .ZN(n831) );
  NAND2_X1 U776 ( .A1(a_6_), .A2(n758), .ZN(n829) );
  NAND2_X1 U777 ( .A1(n832), .A2(n833), .ZN(n758) );
  NAND2_X1 U778 ( .A1(b_7_), .A2(n834), .ZN(n833) );
  OR2_X1 U779 ( .A1(n749), .A2(a_7_), .ZN(n834) );
  NAND2_X1 U780 ( .A1(a_7_), .A2(n749), .ZN(n832) );
  NAND2_X1 U781 ( .A1(n835), .A2(n836), .ZN(n749) );
  NAND2_X1 U782 ( .A1(b_8_), .A2(n837), .ZN(n836) );
  OR2_X1 U783 ( .A1(n740), .A2(a_8_), .ZN(n837) );
  NAND2_X1 U784 ( .A1(a_8_), .A2(n740), .ZN(n835) );
  NAND2_X1 U785 ( .A1(n838), .A2(n839), .ZN(n740) );
  NAND2_X1 U786 ( .A1(b_9_), .A2(n840), .ZN(n839) );
  OR2_X1 U787 ( .A1(n731), .A2(a_9_), .ZN(n840) );
  NAND2_X1 U788 ( .A1(a_9_), .A2(n731), .ZN(n838) );
  NAND2_X1 U789 ( .A1(n841), .A2(n842), .ZN(n731) );
  NAND2_X1 U790 ( .A1(b_10_), .A2(n843), .ZN(n842) );
  OR2_X1 U791 ( .A1(n722), .A2(a_10_), .ZN(n843) );
  NAND2_X1 U792 ( .A1(a_10_), .A2(n722), .ZN(n841) );
  NAND2_X1 U793 ( .A1(n844), .A2(n845), .ZN(n722) );
  NAND2_X1 U794 ( .A1(b_11_), .A2(n846), .ZN(n845) );
  OR2_X1 U795 ( .A1(n713), .A2(a_11_), .ZN(n846) );
  NAND2_X1 U796 ( .A1(a_11_), .A2(n713), .ZN(n844) );
  NAND2_X1 U797 ( .A1(n847), .A2(n848), .ZN(n713) );
  NAND2_X1 U798 ( .A1(b_12_), .A2(n849), .ZN(n848) );
  OR2_X1 U799 ( .A1(n704), .A2(a_12_), .ZN(n849) );
  NAND2_X1 U800 ( .A1(a_12_), .A2(n704), .ZN(n847) );
  NAND2_X1 U801 ( .A1(n850), .A2(n851), .ZN(n704) );
  NAND2_X1 U802 ( .A1(b_13_), .A2(n852), .ZN(n851) );
  OR2_X1 U803 ( .A1(n695), .A2(a_13_), .ZN(n852) );
  NAND2_X1 U804 ( .A1(a_13_), .A2(n695), .ZN(n850) );
  NAND2_X1 U805 ( .A1(n853), .A2(n854), .ZN(n695) );
  NAND2_X1 U806 ( .A1(b_14_), .A2(n855), .ZN(n854) );
  OR2_X1 U807 ( .A1(n686), .A2(a_14_), .ZN(n855) );
  NAND2_X1 U808 ( .A1(a_14_), .A2(n686), .ZN(n853) );
  NAND2_X1 U809 ( .A1(n856), .A2(n857), .ZN(n686) );
  NAND2_X1 U810 ( .A1(b_15_), .A2(n858), .ZN(n857) );
  OR2_X1 U811 ( .A1(n677), .A2(a_15_), .ZN(n858) );
  NAND2_X1 U812 ( .A1(a_15_), .A2(n677), .ZN(n856) );
  NAND2_X1 U813 ( .A1(n859), .A2(n860), .ZN(n677) );
  NAND2_X1 U814 ( .A1(b_16_), .A2(n861), .ZN(n860) );
  OR2_X1 U815 ( .A1(n668), .A2(a_16_), .ZN(n861) );
  NAND2_X1 U816 ( .A1(a_16_), .A2(n668), .ZN(n859) );
  NAND2_X1 U817 ( .A1(n862), .A2(n863), .ZN(n668) );
  NAND2_X1 U818 ( .A1(b_17_), .A2(n864), .ZN(n863) );
  OR2_X1 U819 ( .A1(n659), .A2(a_17_), .ZN(n864) );
  NAND2_X1 U820 ( .A1(a_17_), .A2(n659), .ZN(n862) );
  NAND2_X1 U821 ( .A1(n865), .A2(n866), .ZN(n659) );
  NAND2_X1 U822 ( .A1(b_18_), .A2(n867), .ZN(n866) );
  OR2_X1 U823 ( .A1(n650), .A2(a_18_), .ZN(n867) );
  NAND2_X1 U824 ( .A1(a_18_), .A2(n650), .ZN(n865) );
  NAND2_X1 U825 ( .A1(n868), .A2(n869), .ZN(n650) );
  NAND2_X1 U826 ( .A1(b_19_), .A2(n870), .ZN(n869) );
  OR2_X1 U827 ( .A1(n641), .A2(a_19_), .ZN(n870) );
  NAND2_X1 U828 ( .A1(a_19_), .A2(n641), .ZN(n868) );
  NAND2_X1 U829 ( .A1(n871), .A2(n872), .ZN(n641) );
  NAND2_X1 U830 ( .A1(b_20_), .A2(n873), .ZN(n872) );
  OR2_X1 U831 ( .A1(n632), .A2(a_20_), .ZN(n873) );
  NAND2_X1 U832 ( .A1(a_20_), .A2(n632), .ZN(n871) );
  NAND2_X1 U833 ( .A1(n874), .A2(n875), .ZN(n632) );
  NAND2_X1 U834 ( .A1(b_21_), .A2(n876), .ZN(n875) );
  OR2_X1 U835 ( .A1(n623), .A2(a_21_), .ZN(n876) );
  NAND2_X1 U836 ( .A1(a_21_), .A2(n623), .ZN(n874) );
  NAND2_X1 U837 ( .A1(n877), .A2(n878), .ZN(n623) );
  NAND2_X1 U838 ( .A1(b_22_), .A2(n879), .ZN(n878) );
  OR2_X1 U839 ( .A1(n614), .A2(a_22_), .ZN(n879) );
  NAND2_X1 U840 ( .A1(a_22_), .A2(n614), .ZN(n877) );
  NAND2_X1 U841 ( .A1(n880), .A2(n881), .ZN(n614) );
  NAND2_X1 U842 ( .A1(b_23_), .A2(n882), .ZN(n881) );
  OR2_X1 U843 ( .A1(n605), .A2(a_23_), .ZN(n882) );
  NAND2_X1 U844 ( .A1(a_23_), .A2(n605), .ZN(n880) );
  NAND2_X1 U845 ( .A1(n883), .A2(n884), .ZN(n605) );
  NAND2_X1 U846 ( .A1(b_24_), .A2(n885), .ZN(n884) );
  OR2_X1 U847 ( .A1(n596), .A2(a_24_), .ZN(n885) );
  NAND2_X1 U848 ( .A1(a_24_), .A2(n596), .ZN(n883) );
  NAND2_X1 U849 ( .A1(n886), .A2(n887), .ZN(n596) );
  NAND2_X1 U850 ( .A1(b_25_), .A2(n888), .ZN(n887) );
  OR2_X1 U851 ( .A1(n587), .A2(a_25_), .ZN(n888) );
  NAND2_X1 U852 ( .A1(a_25_), .A2(n587), .ZN(n886) );
  NAND2_X1 U853 ( .A1(n889), .A2(n890), .ZN(n587) );
  NAND2_X1 U854 ( .A1(b_26_), .A2(n891), .ZN(n890) );
  OR2_X1 U855 ( .A1(n578), .A2(a_26_), .ZN(n891) );
  NAND2_X1 U856 ( .A1(a_26_), .A2(n578), .ZN(n889) );
  NAND2_X1 U857 ( .A1(n892), .A2(n893), .ZN(n578) );
  NAND2_X1 U858 ( .A1(b_27_), .A2(n894), .ZN(n893) );
  OR2_X1 U859 ( .A1(n569), .A2(a_27_), .ZN(n894) );
  NAND2_X1 U860 ( .A1(a_27_), .A2(n569), .ZN(n892) );
  NAND2_X1 U861 ( .A1(n895), .A2(n896), .ZN(n569) );
  NAND2_X1 U862 ( .A1(b_28_), .A2(n897), .ZN(n896) );
  OR2_X1 U863 ( .A1(n560), .A2(a_28_), .ZN(n897) );
  NAND2_X1 U864 ( .A1(a_28_), .A2(n560), .ZN(n895) );
  NAND2_X1 U865 ( .A1(n898), .A2(n899), .ZN(n560) );
  NAND2_X1 U866 ( .A1(b_29_), .A2(n900), .ZN(n899) );
  OR2_X1 U867 ( .A1(n551), .A2(a_29_), .ZN(n900) );
  NAND2_X1 U868 ( .A1(a_29_), .A2(n551), .ZN(n898) );
  NAND2_X1 U869 ( .A1(n901), .A2(n902), .ZN(n551) );
  NAND2_X1 U870 ( .A1(b_30_), .A2(n903), .ZN(n902) );
  NAND2_X1 U871 ( .A1(n543), .A2(n904), .ZN(n903) );
  NAND2_X1 U872 ( .A1(n545), .A2(a_30_), .ZN(n901) );
  INV_X1 U873 ( .A(n904), .ZN(n545) );
  NAND2_X1 U874 ( .A1(b_31_), .A2(a_31_), .ZN(n904) );
  NAND2_X1 U875 ( .A1(n905), .A2(n546), .ZN(n544) );
  INV_X1 U876 ( .A(Result_9_), .ZN(n546) );
  NAND4_X1 U877 ( .A1(n906), .A2(n907), .A3(n908), .A4(n909), .ZN(n905) );
  NOR4_X1 U878 ( .A1(n910), .A2(n911), .A3(n912), .A4(n913), .ZN(n909) );
  NAND4_X1 U879 ( .A1(n536), .A2(n807), .A3(n671), .A4(n680), .ZN(n910) );
  NOR4_X1 U880 ( .A1(n914), .A2(n915), .A3(n916), .A4(n917), .ZN(n908) );
  NAND3_X1 U881 ( .A1(n734), .A2(n752), .A3(n716), .ZN(n914) );
  NOR4_X1 U882 ( .A1(n918), .A2(n919), .A3(n920), .A4(n921), .ZN(n907) );
  NOR2_X1 U883 ( .A1(a_31_), .A2(n531), .ZN(n919) );
  NAND4_X1 U884 ( .A1(n707), .A2(n635), .A3(n617), .A4(n599), .ZN(n918) );
  NOR4_X1 U885 ( .A1(n922), .A2(n923), .A3(n924), .A4(n925), .ZN(n906) );
  NAND3_X1 U886 ( .A1(n926), .A2(n927), .A3(n928), .ZN(n922) );
  NAND2_X1 U887 ( .A1(n929), .A2(Result_9_), .ZN(n808) );
  NAND3_X1 U888 ( .A1(n932), .A2(n807), .A3(n933), .ZN(n930) );
  NAND3_X1 U889 ( .A1(n798), .A2(n934), .A3(n806), .ZN(n933) );
  NAND2_X1 U890 ( .A1(n935), .A2(n797), .ZN(n934) );
  NAND2_X1 U891 ( .A1(n789), .A2(n936), .ZN(n935) );
  NAND2_X1 U892 ( .A1(n937), .A2(n938), .ZN(n936) );
  NAND3_X1 U893 ( .A1(n780), .A2(n939), .A3(n771), .ZN(n938) );
  NAND2_X1 U894 ( .A1(n940), .A2(n941), .ZN(n939) );
  NAND3_X1 U895 ( .A1(n762), .A2(n942), .A3(n753), .ZN(n941) );
  NAND3_X1 U896 ( .A1(n943), .A2(n752), .A3(n743), .ZN(n942) );
  NAND3_X1 U897 ( .A1(n744), .A2(n944), .A3(n735), .ZN(n943) );
  NAND3_X1 U898 ( .A1(n945), .A2(n734), .A3(n725), .ZN(n944) );
  NAND3_X1 U899 ( .A1(n726), .A2(n946), .A3(n717), .ZN(n945) );
  NAND3_X1 U900 ( .A1(n947), .A2(n716), .A3(n707), .ZN(n946) );
  NAND3_X1 U901 ( .A1(n708), .A2(n948), .A3(n699), .ZN(n947) );
  NAND2_X1 U902 ( .A1(n949), .A2(n950), .ZN(n948) );
  NAND3_X1 U903 ( .A1(n690), .A2(n951), .A3(n681), .ZN(n950) );
  NAND3_X1 U904 ( .A1(n671), .A2(n680), .A3(n952), .ZN(n951) );
  NAND3_X1 U905 ( .A1(n672), .A2(n953), .A3(n663), .ZN(n952) );
  NAND2_X1 U906 ( .A1(n928), .A2(n954), .ZN(n953) );
  NAND3_X1 U907 ( .A1(n654), .A2(n955), .A3(n645), .ZN(n954) );
  NAND3_X1 U908 ( .A1(n956), .A2(n644), .A3(n635), .ZN(n955) );
  NAND3_X1 U909 ( .A1(n636), .A2(n957), .A3(n627), .ZN(n956) );
  NAND3_X1 U910 ( .A1(n958), .A2(n626), .A3(n617), .ZN(n957) );
  NAND3_X1 U911 ( .A1(n618), .A2(n959), .A3(n609), .ZN(n958) );
  NAND3_X1 U912 ( .A1(n960), .A2(n608), .A3(n599), .ZN(n959) );
  NAND3_X1 U913 ( .A1(n600), .A2(n961), .A3(n591), .ZN(n960) );
  NAND2_X1 U914 ( .A1(n926), .A2(n962), .ZN(n961) );
  NAND3_X1 U915 ( .A1(n582), .A2(n963), .A3(n573), .ZN(n962) );
  NAND2_X1 U916 ( .A1(n927), .A2(n964), .ZN(n963) );
  AND2_X1 U917 ( .A1(n563), .A2(n572), .ZN(n927) );
  AND2_X1 U918 ( .A1(n581), .A2(n590), .ZN(n926) );
  AND2_X1 U919 ( .A1(n653), .A2(n662), .ZN(n928) );
  INV_X1 U920 ( .A(n924), .ZN(n949) );
  NAND2_X1 U921 ( .A1(n689), .A2(n698), .ZN(n924) );
  INV_X1 U922 ( .A(n925), .ZN(n940) );
  NAND2_X1 U923 ( .A1(n761), .A2(n770), .ZN(n925) );
  INV_X1 U924 ( .A(n923), .ZN(n937) );
  NAND2_X1 U925 ( .A1(n779), .A2(n788), .ZN(n923) );
  NAND3_X1 U926 ( .A1(n811), .A2(n807), .A3(n965), .ZN(n929) );
  NAND2_X1 U927 ( .A1(n805), .A2(n806), .ZN(n965) );
  NAND2_X1 U928 ( .A1(a_1_), .A2(n816), .ZN(n806) );
  NAND2_X1 U929 ( .A1(n797), .A2(n966), .ZN(n805) );
  NAND2_X1 U930 ( .A1(n798), .A2(n796), .ZN(n966) );
  NAND2_X1 U931 ( .A1(n788), .A2(n967), .ZN(n796) );
  NAND2_X1 U932 ( .A1(n789), .A2(n787), .ZN(n967) );
  NAND2_X1 U933 ( .A1(n779), .A2(n968), .ZN(n787) );
  NAND2_X1 U934 ( .A1(n780), .A2(n778), .ZN(n968) );
  NAND2_X1 U935 ( .A1(n770), .A2(n969), .ZN(n778) );
  NAND2_X1 U936 ( .A1(n771), .A2(n769), .ZN(n969) );
  NAND2_X1 U937 ( .A1(n761), .A2(n970), .ZN(n769) );
  NAND2_X1 U938 ( .A1(n762), .A2(n760), .ZN(n970) );
  NAND2_X1 U939 ( .A1(n752), .A2(n971), .ZN(n760) );
  NAND2_X1 U940 ( .A1(n753), .A2(n751), .ZN(n971) );
  NAND2_X1 U941 ( .A1(n743), .A2(n972), .ZN(n751) );
  NAND2_X1 U942 ( .A1(n744), .A2(n742), .ZN(n972) );
  NAND2_X1 U943 ( .A1(n734), .A2(n973), .ZN(n742) );
  NAND2_X1 U944 ( .A1(n735), .A2(n733), .ZN(n973) );
  NAND2_X1 U945 ( .A1(n725), .A2(n974), .ZN(n733) );
  NAND2_X1 U946 ( .A1(n726), .A2(n724), .ZN(n974) );
  NAND2_X1 U947 ( .A1(n716), .A2(n975), .ZN(n724) );
  NAND2_X1 U948 ( .A1(n717), .A2(n715), .ZN(n975) );
  NAND2_X1 U949 ( .A1(n707), .A2(n976), .ZN(n715) );
  NAND2_X1 U950 ( .A1(n708), .A2(n706), .ZN(n976) );
  NAND2_X1 U951 ( .A1(n698), .A2(n977), .ZN(n706) );
  NAND2_X1 U952 ( .A1(n699), .A2(n697), .ZN(n977) );
  NAND2_X1 U953 ( .A1(n689), .A2(n978), .ZN(n697) );
  NAND2_X1 U954 ( .A1(n690), .A2(n688), .ZN(n978) );
  NAND2_X1 U955 ( .A1(n680), .A2(n979), .ZN(n688) );
  NAND2_X1 U956 ( .A1(n681), .A2(n679), .ZN(n979) );
  NAND2_X1 U957 ( .A1(n671), .A2(n980), .ZN(n679) );
  NAND2_X1 U958 ( .A1(n672), .A2(n670), .ZN(n980) );
  NAND2_X1 U959 ( .A1(n662), .A2(n981), .ZN(n670) );
  NAND2_X1 U960 ( .A1(n663), .A2(n661), .ZN(n981) );
  NAND2_X1 U961 ( .A1(n653), .A2(n982), .ZN(n661) );
  NAND2_X1 U962 ( .A1(n654), .A2(n652), .ZN(n982) );
  NAND2_X1 U963 ( .A1(n644), .A2(n983), .ZN(n652) );
  NAND2_X1 U964 ( .A1(n645), .A2(n643), .ZN(n983) );
  NAND2_X1 U965 ( .A1(n635), .A2(n984), .ZN(n643) );
  NAND2_X1 U966 ( .A1(n636), .A2(n634), .ZN(n984) );
  NAND2_X1 U967 ( .A1(n626), .A2(n985), .ZN(n634) );
  NAND2_X1 U968 ( .A1(n627), .A2(n625), .ZN(n985) );
  NAND2_X1 U969 ( .A1(n617), .A2(n986), .ZN(n625) );
  NAND2_X1 U970 ( .A1(n618), .A2(n616), .ZN(n986) );
  NAND2_X1 U971 ( .A1(n608), .A2(n987), .ZN(n616) );
  NAND2_X1 U972 ( .A1(n609), .A2(n607), .ZN(n987) );
  NAND2_X1 U973 ( .A1(n599), .A2(n988), .ZN(n607) );
  NAND2_X1 U974 ( .A1(n600), .A2(n598), .ZN(n988) );
  NAND2_X1 U975 ( .A1(n590), .A2(n989), .ZN(n598) );
  NAND2_X1 U976 ( .A1(n591), .A2(n589), .ZN(n989) );
  NAND2_X1 U977 ( .A1(n581), .A2(n990), .ZN(n589) );
  NAND2_X1 U978 ( .A1(n582), .A2(n580), .ZN(n990) );
  NAND2_X1 U979 ( .A1(n572), .A2(n991), .ZN(n580) );
  NAND2_X1 U980 ( .A1(n573), .A2(n571), .ZN(n991) );
  NAND2_X1 U981 ( .A1(n563), .A2(n964), .ZN(n571) );
  NAND2_X1 U982 ( .A1(n562), .A2(n564), .ZN(n964) );
  NAND2_X1 U983 ( .A1(a_28_), .A2(n992), .ZN(n564) );
  NAND2_X1 U984 ( .A1(n554), .A2(n993), .ZN(n562) );
  NAND2_X1 U985 ( .A1(n555), .A2(n553), .ZN(n993) );
  NAND2_X1 U986 ( .A1(n536), .A2(n994), .ZN(n553) );
  NAND2_X1 U987 ( .A1(n995), .A2(n535), .ZN(n994) );
  OR2_X1 U988 ( .A1(n543), .A2(b_30_), .ZN(n535) );
  NAND2_X1 U989 ( .A1(a_31_), .A2(n531), .ZN(n995) );
  INV_X1 U990 ( .A(b_31_), .ZN(n531) );
  NAND2_X1 U991 ( .A1(b_30_), .A2(n543), .ZN(n536) );
  INV_X1 U992 ( .A(a_30_), .ZN(n543) );
  NAND2_X1 U993 ( .A1(a_29_), .A2(n996), .ZN(n555) );
  INV_X1 U994 ( .A(n912), .ZN(n554) );
  NOR2_X1 U995 ( .A1(n996), .A2(a_29_), .ZN(n912) );
  INV_X1 U996 ( .A(b_29_), .ZN(n996) );
  OR2_X1 U997 ( .A1(n992), .A2(a_28_), .ZN(n563) );
  INV_X1 U998 ( .A(b_28_), .ZN(n992) );
  NAND2_X1 U999 ( .A1(a_27_), .A2(n997), .ZN(n573) );
  OR2_X1 U1000 ( .A1(n997), .A2(a_27_), .ZN(n572) );
  INV_X1 U1001 ( .A(b_27_), .ZN(n997) );
  NAND2_X1 U1002 ( .A1(a_26_), .A2(n998), .ZN(n582) );
  OR2_X1 U1003 ( .A1(n998), .A2(a_26_), .ZN(n581) );
  INV_X1 U1004 ( .A(b_26_), .ZN(n998) );
  NAND2_X1 U1005 ( .A1(a_25_), .A2(n999), .ZN(n591) );
  OR2_X1 U1006 ( .A1(n999), .A2(a_25_), .ZN(n590) );
  INV_X1 U1007 ( .A(b_25_), .ZN(n999) );
  NAND2_X1 U1008 ( .A1(a_24_), .A2(n1000), .ZN(n600) );
  OR2_X1 U1009 ( .A1(n1000), .A2(a_24_), .ZN(n599) );
  INV_X1 U1010 ( .A(b_24_), .ZN(n1000) );
  NAND2_X1 U1011 ( .A1(a_23_), .A2(n1001), .ZN(n609) );
  INV_X1 U1012 ( .A(n915), .ZN(n608) );
  NOR2_X1 U1013 ( .A1(n1001), .A2(a_23_), .ZN(n915) );
  INV_X1 U1014 ( .A(b_23_), .ZN(n1001) );
  NAND2_X1 U1015 ( .A1(a_22_), .A2(n1002), .ZN(n618) );
  OR2_X1 U1016 ( .A1(n1002), .A2(a_22_), .ZN(n617) );
  INV_X1 U1017 ( .A(b_22_), .ZN(n1002) );
  NAND2_X1 U1018 ( .A1(a_21_), .A2(n1003), .ZN(n627) );
  INV_X1 U1019 ( .A(n917), .ZN(n626) );
  NOR2_X1 U1020 ( .A1(n1003), .A2(a_21_), .ZN(n917) );
  INV_X1 U1021 ( .A(b_21_), .ZN(n1003) );
  NAND2_X1 U1022 ( .A1(a_20_), .A2(n1004), .ZN(n636) );
  OR2_X1 U1023 ( .A1(n1004), .A2(a_20_), .ZN(n635) );
  INV_X1 U1024 ( .A(b_20_), .ZN(n1004) );
  NAND2_X1 U1025 ( .A1(a_19_), .A2(n1005), .ZN(n645) );
  INV_X1 U1026 ( .A(n916), .ZN(n644) );
  NOR2_X1 U1027 ( .A1(n1005), .A2(a_19_), .ZN(n916) );
  INV_X1 U1028 ( .A(b_19_), .ZN(n1005) );
  NAND2_X1 U1029 ( .A1(a_18_), .A2(n1006), .ZN(n654) );
  OR2_X1 U1030 ( .A1(n1006), .A2(a_18_), .ZN(n653) );
  INV_X1 U1031 ( .A(b_18_), .ZN(n1006) );
  NAND2_X1 U1032 ( .A1(a_17_), .A2(n1007), .ZN(n663) );
  OR2_X1 U1033 ( .A1(n1007), .A2(a_17_), .ZN(n662) );
  INV_X1 U1034 ( .A(b_17_), .ZN(n1007) );
  NAND2_X1 U1035 ( .A1(a_16_), .A2(n1008), .ZN(n672) );
  OR2_X1 U1036 ( .A1(n1008), .A2(a_16_), .ZN(n671) );
  INV_X1 U1037 ( .A(b_16_), .ZN(n1008) );
  NAND2_X1 U1038 ( .A1(a_15_), .A2(n1009), .ZN(n681) );
  OR2_X1 U1039 ( .A1(n1009), .A2(a_15_), .ZN(n680) );
  INV_X1 U1040 ( .A(b_15_), .ZN(n1009) );
  NAND2_X1 U1041 ( .A1(a_14_), .A2(n1010), .ZN(n690) );
  OR2_X1 U1042 ( .A1(n1010), .A2(a_14_), .ZN(n689) );
  INV_X1 U1043 ( .A(b_14_), .ZN(n1010) );
  NAND2_X1 U1044 ( .A1(a_13_), .A2(n1011), .ZN(n699) );
  OR2_X1 U1045 ( .A1(n1011), .A2(a_13_), .ZN(n698) );
  INV_X1 U1046 ( .A(b_13_), .ZN(n1011) );
  NAND2_X1 U1047 ( .A1(a_12_), .A2(n1012), .ZN(n708) );
  OR2_X1 U1048 ( .A1(n1012), .A2(a_12_), .ZN(n707) );
  INV_X1 U1049 ( .A(b_12_), .ZN(n1012) );
  NAND2_X1 U1050 ( .A1(a_11_), .A2(n1013), .ZN(n717) );
  OR2_X1 U1051 ( .A1(n1013), .A2(a_11_), .ZN(n716) );
  INV_X1 U1052 ( .A(b_11_), .ZN(n1013) );
  NAND2_X1 U1053 ( .A1(a_10_), .A2(n1014), .ZN(n726) );
  INV_X1 U1054 ( .A(n920), .ZN(n725) );
  NOR2_X1 U1055 ( .A1(n1014), .A2(a_10_), .ZN(n920) );
  INV_X1 U1056 ( .A(b_10_), .ZN(n1014) );
  NAND2_X1 U1057 ( .A1(a_9_), .A2(n1015), .ZN(n735) );
  OR2_X1 U1058 ( .A1(n1015), .A2(a_9_), .ZN(n734) );
  INV_X1 U1059 ( .A(b_9_), .ZN(n1015) );
  NAND2_X1 U1060 ( .A1(a_8_), .A2(n1016), .ZN(n744) );
  INV_X1 U1061 ( .A(n921), .ZN(n743) );
  NOR2_X1 U1062 ( .A1(n1016), .A2(a_8_), .ZN(n921) );
  INV_X1 U1063 ( .A(b_8_), .ZN(n1016) );
  NAND2_X1 U1064 ( .A1(a_7_), .A2(n1017), .ZN(n753) );
  OR2_X1 U1065 ( .A1(n1017), .A2(a_7_), .ZN(n752) );
  INV_X1 U1066 ( .A(b_7_), .ZN(n1017) );
  NAND2_X1 U1067 ( .A1(a_6_), .A2(n1018), .ZN(n762) );
  OR2_X1 U1068 ( .A1(n1018), .A2(a_6_), .ZN(n761) );
  INV_X1 U1069 ( .A(b_6_), .ZN(n1018) );
  NAND2_X1 U1070 ( .A1(a_5_), .A2(n1019), .ZN(n771) );
  OR2_X1 U1071 ( .A1(n1019), .A2(a_5_), .ZN(n770) );
  INV_X1 U1072 ( .A(b_5_), .ZN(n1019) );
  NAND2_X1 U1073 ( .A1(a_4_), .A2(n1020), .ZN(n780) );
  OR2_X1 U1074 ( .A1(n1020), .A2(a_4_), .ZN(n779) );
  INV_X1 U1075 ( .A(b_4_), .ZN(n1020) );
  NAND2_X1 U1076 ( .A1(a_3_), .A2(n1021), .ZN(n789) );
  OR2_X1 U1077 ( .A1(n1021), .A2(a_3_), .ZN(n788) );
  INV_X1 U1078 ( .A(b_3_), .ZN(n1021) );
  NAND2_X1 U1079 ( .A1(a_2_), .A2(n1022), .ZN(n798) );
  INV_X1 U1080 ( .A(n911), .ZN(n797) );
  NOR2_X1 U1081 ( .A1(n1022), .A2(a_2_), .ZN(n911) );
  INV_X1 U1082 ( .A(b_2_), .ZN(n1022) );
  OR2_X1 U1083 ( .A1(n816), .A2(a_1_), .ZN(n807) );
  INV_X1 U1084 ( .A(b_1_), .ZN(n816) );
  NAND2_X1 U1085 ( .A1(n932), .A2(n931), .ZN(n811) );
  NAND2_X1 U1086 ( .A1(a_0_), .A2(n1023), .ZN(n931) );
  INV_X1 U1087 ( .A(n913), .ZN(n932) );
  NOR2_X1 U1088 ( .A1(n1023), .A2(a_0_), .ZN(n913) );
  INV_X1 U1089 ( .A(b_0_), .ZN(n1023) );
endmodule

