module add_mul_comp_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393;

  NOR2_X2 U2209 ( .A1(n4250), .A2(n2487), .ZN(n2488) );
  INV_X2 U2210 ( .A(n2223), .ZN(n2177) );
  NOR2_X1 U2211 ( .A1(n2177), .A2(n2178), .ZN(Result_9_) );
  XOR2_X1 U2212 ( .A(n2179), .B(n2180), .Z(n2178) );
  NOR2_X1 U2213 ( .A1(n2181), .A2(n2182), .ZN(n2180) );
  NOR2_X1 U2214 ( .A1(n2183), .A2(n2184), .ZN(n2182) );
  NOR2_X1 U2215 ( .A1(n2177), .A2(n2185), .ZN(Result_8_) );
  XNOR2_X1 U2216 ( .A(n2186), .B(n2187), .ZN(n2185) );
  NOR2_X1 U2217 ( .A1(n2177), .A2(n2188), .ZN(Result_7_) );
  XOR2_X1 U2218 ( .A(n2189), .B(n2190), .Z(n2188) );
  NOR2_X1 U2219 ( .A1(n2191), .A2(n2192), .ZN(n2190) );
  NOR2_X1 U2220 ( .A1(n2193), .A2(n2194), .ZN(n2192) );
  NOR2_X1 U2221 ( .A1(n2177), .A2(n2195), .ZN(Result_6_) );
  XOR2_X1 U2222 ( .A(n2196), .B(n2197), .Z(n2195) );
  NOR2_X1 U2223 ( .A1(n2177), .A2(n2198), .ZN(Result_5_) );
  XNOR2_X1 U2224 ( .A(n2199), .B(n2200), .ZN(n2198) );
  NOR2_X1 U2225 ( .A1(n2201), .A2(n2202), .ZN(n2200) );
  NOR2_X1 U2226 ( .A1(n2203), .A2(n2204), .ZN(n2202) );
  NOR2_X1 U2227 ( .A1(n2177), .A2(n2205), .ZN(Result_4_) );
  XOR2_X1 U2228 ( .A(n2206), .B(n2207), .Z(n2205) );
  NOR2_X1 U2229 ( .A1(n2177), .A2(n2208), .ZN(Result_3_) );
  XNOR2_X1 U2230 ( .A(n2209), .B(n2210), .ZN(n2208) );
  NOR2_X1 U2231 ( .A1(n2211), .A2(n2212), .ZN(n2210) );
  NOR2_X1 U2232 ( .A1(n2213), .A2(n2214), .ZN(n2212) );
  NAND2_X1 U2233 ( .A1(n2215), .A2(n2216), .ZN(Result_31_) );
  INV_X1 U2234 ( .A(n2217), .ZN(n2216) );
  NOR2_X1 U2235 ( .A1(n2218), .A2(n2177), .ZN(n2217) );
  NAND2_X1 U2236 ( .A1(n2219), .A2(n2177), .ZN(n2215) );
  XOR2_X1 U2237 ( .A(b_15_), .B(a_15_), .Z(n2219) );
  NAND2_X1 U2238 ( .A1(n2220), .A2(n2221), .ZN(Result_30_) );
  NAND2_X1 U2239 ( .A1(n2222), .A2(n2223), .ZN(n2221) );
  NAND2_X1 U2240 ( .A1(n2224), .A2(n2225), .ZN(n2222) );
  NAND2_X1 U2241 ( .A1(b_14_), .A2(n2226), .ZN(n2225) );
  NAND2_X1 U2242 ( .A1(n2227), .A2(n2228), .ZN(n2226) );
  NAND2_X1 U2243 ( .A1(a_15_), .A2(n2229), .ZN(n2228) );
  NAND2_X1 U2244 ( .A1(b_15_), .A2(n2230), .ZN(n2224) );
  NAND2_X1 U2245 ( .A1(n2231), .A2(n2232), .ZN(n2230) );
  NAND2_X1 U2246 ( .A1(a_14_), .A2(n2233), .ZN(n2232) );
  NAND2_X1 U2247 ( .A1(n2234), .A2(n2177), .ZN(n2220) );
  XNOR2_X1 U2248 ( .A(n2218), .B(n2235), .ZN(n2234) );
  XOR2_X1 U2249 ( .A(b_14_), .B(a_14_), .Z(n2235) );
  NOR2_X1 U2250 ( .A1(n2177), .A2(n2236), .ZN(Result_2_) );
  XOR2_X1 U2251 ( .A(n2237), .B(n2238), .Z(n2236) );
  NAND2_X1 U2252 ( .A1(n2239), .A2(n2240), .ZN(Result_29_) );
  NAND2_X1 U2253 ( .A1(n2177), .A2(n2241), .ZN(n2240) );
  NAND2_X1 U2254 ( .A1(n2242), .A2(n2243), .ZN(n2241) );
  NAND2_X1 U2255 ( .A1(n2244), .A2(n2245), .ZN(n2243) );
  NOR2_X1 U2256 ( .A1(n2246), .A2(n2247), .ZN(n2242) );
  NOR2_X1 U2257 ( .A1(b_13_), .A2(n2248), .ZN(n2247) );
  XOR2_X1 U2258 ( .A(a_13_), .B(n2249), .Z(n2248) );
  NOR2_X1 U2259 ( .A1(n2250), .A2(n2251), .ZN(n2246) );
  NAND2_X1 U2260 ( .A1(n2249), .A2(n2252), .ZN(n2251) );
  NAND2_X1 U2261 ( .A1(n2253), .A2(n2223), .ZN(n2239) );
  XOR2_X1 U2262 ( .A(n2254), .B(n2255), .Z(n2253) );
  XOR2_X1 U2263 ( .A(n2256), .B(n2257), .Z(n2255) );
  NAND2_X1 U2264 ( .A1(n2258), .A2(n2259), .ZN(Result_28_) );
  NAND2_X1 U2265 ( .A1(n2260), .A2(n2223), .ZN(n2259) );
  XOR2_X1 U2266 ( .A(n2261), .B(n2262), .Z(n2260) );
  XOR2_X1 U2267 ( .A(n2263), .B(n2264), .Z(n2261) );
  NAND2_X1 U2268 ( .A1(n2177), .A2(n2265), .ZN(n2258) );
  XOR2_X1 U2269 ( .A(n2266), .B(n2267), .Z(n2265) );
  NAND2_X1 U2270 ( .A1(n2268), .A2(n2269), .ZN(n2266) );
  NAND2_X1 U2271 ( .A1(n2270), .A2(n2271), .ZN(Result_27_) );
  NAND2_X1 U2272 ( .A1(n2177), .A2(n2272), .ZN(n2271) );
  NAND2_X1 U2273 ( .A1(n2273), .A2(n2274), .ZN(n2272) );
  NAND2_X1 U2274 ( .A1(n2275), .A2(n2276), .ZN(n2274) );
  NOR2_X1 U2275 ( .A1(n2277), .A2(n2278), .ZN(n2273) );
  NOR2_X1 U2276 ( .A1(b_11_), .A2(n2279), .ZN(n2278) );
  XOR2_X1 U2277 ( .A(n2280), .B(n2276), .Z(n2279) );
  NOR2_X1 U2278 ( .A1(n2281), .A2(n2282), .ZN(n2277) );
  INV_X1 U2279 ( .A(n2283), .ZN(n2282) );
  NOR2_X1 U2280 ( .A1(n2276), .A2(a_11_), .ZN(n2283) );
  NAND2_X1 U2281 ( .A1(n2284), .A2(n2223), .ZN(n2270) );
  XNOR2_X1 U2282 ( .A(n2285), .B(n2286), .ZN(n2284) );
  NAND2_X1 U2283 ( .A1(n2287), .A2(n2288), .ZN(n2285) );
  NAND2_X1 U2284 ( .A1(n2289), .A2(n2290), .ZN(Result_26_) );
  NAND2_X1 U2285 ( .A1(n2291), .A2(n2223), .ZN(n2290) );
  XOR2_X1 U2286 ( .A(n2292), .B(n2293), .Z(n2291) );
  XNOR2_X1 U2287 ( .A(n2294), .B(n2295), .ZN(n2293) );
  NAND2_X1 U2288 ( .A1(n2177), .A2(n2296), .ZN(n2289) );
  XNOR2_X1 U2289 ( .A(n2297), .B(n2298), .ZN(n2296) );
  NAND2_X1 U2290 ( .A1(n2299), .A2(n2300), .ZN(n2298) );
  NAND2_X1 U2291 ( .A1(n2301), .A2(n2302), .ZN(Result_25_) );
  NAND2_X1 U2292 ( .A1(n2177), .A2(n2303), .ZN(n2302) );
  NAND2_X1 U2293 ( .A1(n2304), .A2(n2305), .ZN(n2303) );
  NAND2_X1 U2294 ( .A1(n2306), .A2(n2307), .ZN(n2305) );
  NOR2_X1 U2295 ( .A1(n2308), .A2(n2309), .ZN(n2304) );
  NOR2_X1 U2296 ( .A1(b_9_), .A2(n2310), .ZN(n2309) );
  XOR2_X1 U2297 ( .A(n2311), .B(n2307), .Z(n2310) );
  NOR2_X1 U2298 ( .A1(n2312), .A2(n2313), .ZN(n2308) );
  INV_X1 U2299 ( .A(n2314), .ZN(n2313) );
  NOR2_X1 U2300 ( .A1(n2307), .A2(a_9_), .ZN(n2314) );
  NAND2_X1 U2301 ( .A1(n2315), .A2(n2223), .ZN(n2301) );
  XNOR2_X1 U2302 ( .A(n2316), .B(n2317), .ZN(n2315) );
  NAND2_X1 U2303 ( .A1(n2318), .A2(n2319), .ZN(n2316) );
  NAND2_X1 U2304 ( .A1(n2320), .A2(n2321), .ZN(Result_24_) );
  NAND2_X1 U2305 ( .A1(n2322), .A2(n2223), .ZN(n2321) );
  XNOR2_X1 U2306 ( .A(n2323), .B(n2324), .ZN(n2322) );
  XOR2_X1 U2307 ( .A(n2325), .B(n2326), .Z(n2324) );
  NAND2_X1 U2308 ( .A1(n2177), .A2(n2327), .ZN(n2320) );
  XOR2_X1 U2309 ( .A(n2328), .B(n2329), .Z(n2327) );
  NOR2_X1 U2310 ( .A1(n2330), .A2(n2331), .ZN(n2329) );
  NAND2_X1 U2311 ( .A1(n2332), .A2(n2333), .ZN(Result_23_) );
  NAND2_X1 U2312 ( .A1(n2177), .A2(n2334), .ZN(n2333) );
  NAND2_X1 U2313 ( .A1(n2335), .A2(n2336), .ZN(n2334) );
  NAND2_X1 U2314 ( .A1(n2337), .A2(n2338), .ZN(n2336) );
  NOR2_X1 U2315 ( .A1(n2339), .A2(n2340), .ZN(n2335) );
  NOR2_X1 U2316 ( .A1(b_7_), .A2(n2341), .ZN(n2340) );
  XOR2_X1 U2317 ( .A(n2342), .B(n2338), .Z(n2341) );
  NOR2_X1 U2318 ( .A1(n2343), .A2(n2344), .ZN(n2339) );
  NAND2_X1 U2319 ( .A1(n2345), .A2(n2342), .ZN(n2344) );
  NAND2_X1 U2320 ( .A1(n2346), .A2(n2223), .ZN(n2332) );
  XNOR2_X1 U2321 ( .A(n2347), .B(n2348), .ZN(n2346) );
  NAND2_X1 U2322 ( .A1(n2349), .A2(n2350), .ZN(n2347) );
  NAND2_X1 U2323 ( .A1(n2351), .A2(n2352), .ZN(Result_22_) );
  NAND2_X1 U2324 ( .A1(n2353), .A2(n2223), .ZN(n2352) );
  XNOR2_X1 U2325 ( .A(n2354), .B(n2355), .ZN(n2353) );
  XOR2_X1 U2326 ( .A(n2356), .B(n2357), .Z(n2355) );
  NAND2_X1 U2327 ( .A1(n2177), .A2(n2358), .ZN(n2351) );
  XNOR2_X1 U2328 ( .A(n2359), .B(n2360), .ZN(n2358) );
  NAND2_X1 U2329 ( .A1(n2361), .A2(n2362), .ZN(n2360) );
  NAND2_X1 U2330 ( .A1(n2363), .A2(n2364), .ZN(Result_21_) );
  NAND2_X1 U2331 ( .A1(n2177), .A2(n2365), .ZN(n2364) );
  NAND2_X1 U2332 ( .A1(n2366), .A2(n2367), .ZN(n2365) );
  NAND2_X1 U2333 ( .A1(n2368), .A2(n2369), .ZN(n2367) );
  NOR2_X1 U2334 ( .A1(n2370), .A2(n2371), .ZN(n2366) );
  NOR2_X1 U2335 ( .A1(b_5_), .A2(n2372), .ZN(n2371) );
  XOR2_X1 U2336 ( .A(n2373), .B(n2369), .Z(n2372) );
  NOR2_X1 U2337 ( .A1(n2374), .A2(n2375), .ZN(n2370) );
  INV_X1 U2338 ( .A(n2376), .ZN(n2375) );
  NOR2_X1 U2339 ( .A1(n2369), .A2(a_5_), .ZN(n2376) );
  NAND2_X1 U2340 ( .A1(n2377), .A2(n2223), .ZN(n2363) );
  XNOR2_X1 U2341 ( .A(n2378), .B(n2379), .ZN(n2377) );
  NAND2_X1 U2342 ( .A1(n2380), .A2(n2381), .ZN(n2378) );
  NAND2_X1 U2343 ( .A1(n2382), .A2(n2383), .ZN(Result_20_) );
  NAND2_X1 U2344 ( .A1(n2384), .A2(n2223), .ZN(n2383) );
  XNOR2_X1 U2345 ( .A(n2385), .B(n2386), .ZN(n2384) );
  XOR2_X1 U2346 ( .A(n2387), .B(n2388), .Z(n2386) );
  NAND2_X1 U2347 ( .A1(n2177), .A2(n2389), .ZN(n2382) );
  XNOR2_X1 U2348 ( .A(n2390), .B(n2391), .ZN(n2389) );
  NAND2_X1 U2349 ( .A1(n2392), .A2(n2393), .ZN(n2391) );
  NOR2_X1 U2350 ( .A1(n2177), .A2(n2394), .ZN(Result_1_) );
  XNOR2_X1 U2351 ( .A(n2395), .B(n2396), .ZN(n2394) );
  NAND2_X1 U2352 ( .A1(n2397), .A2(n2398), .ZN(n2396) );
  NAND2_X1 U2353 ( .A1(n2399), .A2(n2237), .ZN(n2395) );
  NAND2_X1 U2354 ( .A1(n2400), .A2(n2401), .ZN(Result_19_) );
  NAND2_X1 U2355 ( .A1(n2177), .A2(n2402), .ZN(n2401) );
  NAND2_X1 U2356 ( .A1(n2403), .A2(n2404), .ZN(n2402) );
  NAND2_X1 U2357 ( .A1(n2405), .A2(n2406), .ZN(n2404) );
  NOR2_X1 U2358 ( .A1(n2407), .A2(n2408), .ZN(n2403) );
  NOR2_X1 U2359 ( .A1(b_3_), .A2(n2409), .ZN(n2408) );
  XOR2_X1 U2360 ( .A(n2410), .B(n2406), .Z(n2409) );
  NOR2_X1 U2361 ( .A1(n2411), .A2(n2412), .ZN(n2407) );
  INV_X1 U2362 ( .A(n2413), .ZN(n2412) );
  NOR2_X1 U2363 ( .A1(n2406), .A2(a_3_), .ZN(n2413) );
  NAND2_X1 U2364 ( .A1(n2414), .A2(n2223), .ZN(n2400) );
  XNOR2_X1 U2365 ( .A(n2415), .B(n2416), .ZN(n2414) );
  NAND2_X1 U2366 ( .A1(n2417), .A2(n2418), .ZN(n2415) );
  NAND2_X1 U2367 ( .A1(n2419), .A2(n2420), .ZN(Result_18_) );
  NAND2_X1 U2368 ( .A1(n2421), .A2(n2223), .ZN(n2420) );
  XOR2_X1 U2369 ( .A(n2422), .B(n2423), .Z(n2421) );
  XOR2_X1 U2370 ( .A(n2424), .B(n2425), .Z(n2422) );
  NOR2_X1 U2371 ( .A1(n2229), .A2(n2426), .ZN(n2425) );
  NAND2_X1 U2372 ( .A1(n2177), .A2(n2427), .ZN(n2419) );
  XNOR2_X1 U2373 ( .A(n2428), .B(n2429), .ZN(n2427) );
  NAND2_X1 U2374 ( .A1(n2430), .A2(n2431), .ZN(n2429) );
  NAND2_X1 U2375 ( .A1(n2432), .A2(n2433), .ZN(Result_17_) );
  NAND2_X1 U2376 ( .A1(n2434), .A2(n2223), .ZN(n2433) );
  XNOR2_X1 U2377 ( .A(n2435), .B(n2436), .ZN(n2434) );
  XOR2_X1 U2378 ( .A(n2437), .B(n2438), .Z(n2436) );
  NAND2_X1 U2379 ( .A1(b_15_), .A2(a_1_), .ZN(n2438) );
  NAND2_X1 U2380 ( .A1(n2439), .A2(n2177), .ZN(n2432) );
  NAND2_X1 U2381 ( .A1(n2440), .A2(n2441), .ZN(n2439) );
  NAND2_X1 U2382 ( .A1(n2442), .A2(n2443), .ZN(n2441) );
  NAND2_X1 U2383 ( .A1(n2444), .A2(n2445), .ZN(n2442) );
  NAND2_X1 U2384 ( .A1(n2446), .A2(n2447), .ZN(n2440) );
  XOR2_X1 U2385 ( .A(b_1_), .B(a_1_), .Z(n2446) );
  NAND2_X1 U2386 ( .A1(n2448), .A2(n2449), .ZN(Result_16_) );
  NAND2_X1 U2387 ( .A1(n2450), .A2(n2223), .ZN(n2449) );
  XNOR2_X1 U2388 ( .A(n2451), .B(n2452), .ZN(n2450) );
  XOR2_X1 U2389 ( .A(n2453), .B(n2454), .Z(n2452) );
  NAND2_X1 U2390 ( .A1(a_0_), .A2(b_15_), .ZN(n2454) );
  NAND2_X1 U2391 ( .A1(n2455), .A2(n2177), .ZN(n2448) );
  XOR2_X1 U2392 ( .A(n2456), .B(n2457), .Z(n2455) );
  NAND2_X1 U2393 ( .A1(n2445), .A2(n2458), .ZN(n2456) );
  NAND2_X1 U2394 ( .A1(n2444), .A2(n2447), .ZN(n2458) );
  INV_X1 U2395 ( .A(n2443), .ZN(n2447) );
  NAND2_X1 U2396 ( .A1(n2431), .A2(n2459), .ZN(n2443) );
  NAND2_X1 U2397 ( .A1(n2430), .A2(n2428), .ZN(n2459) );
  NAND2_X1 U2398 ( .A1(n2460), .A2(n2461), .ZN(n2428) );
  NAND2_X1 U2399 ( .A1(n2462), .A2(n2406), .ZN(n2461) );
  NAND2_X1 U2400 ( .A1(n2393), .A2(n2463), .ZN(n2406) );
  NAND2_X1 U2401 ( .A1(n2392), .A2(n2390), .ZN(n2463) );
  NAND2_X1 U2402 ( .A1(n2464), .A2(n2465), .ZN(n2390) );
  NAND2_X1 U2403 ( .A1(n2466), .A2(n2369), .ZN(n2465) );
  NAND2_X1 U2404 ( .A1(n2362), .A2(n2467), .ZN(n2369) );
  NAND2_X1 U2405 ( .A1(n2361), .A2(n2359), .ZN(n2467) );
  NAND2_X1 U2406 ( .A1(n2468), .A2(n2469), .ZN(n2359) );
  NAND2_X1 U2407 ( .A1(n2470), .A2(n2338), .ZN(n2469) );
  INV_X1 U2408 ( .A(n2345), .ZN(n2338) );
  NOR2_X1 U2409 ( .A1(n2331), .A2(n2471), .ZN(n2345) );
  NOR2_X1 U2410 ( .A1(n2330), .A2(n2472), .ZN(n2471) );
  INV_X1 U2411 ( .A(n2328), .ZN(n2472) );
  NAND2_X1 U2412 ( .A1(n2473), .A2(n2474), .ZN(n2328) );
  NAND2_X1 U2413 ( .A1(n2475), .A2(n2307), .ZN(n2474) );
  NAND2_X1 U2414 ( .A1(n2300), .A2(n2476), .ZN(n2307) );
  NAND2_X1 U2415 ( .A1(n2299), .A2(n2297), .ZN(n2476) );
  NAND2_X1 U2416 ( .A1(n2477), .A2(n2478), .ZN(n2297) );
  NAND2_X1 U2417 ( .A1(n2479), .A2(n2276), .ZN(n2478) );
  NAND2_X1 U2418 ( .A1(n2268), .A2(n2480), .ZN(n2276) );
  NAND2_X1 U2419 ( .A1(n2269), .A2(n2481), .ZN(n2480) );
  INV_X1 U2420 ( .A(n2267), .ZN(n2481) );
  NOR2_X1 U2421 ( .A1(n2244), .A2(n2482), .ZN(n2267) );
  NOR2_X1 U2422 ( .A1(n2483), .A2(n2249), .ZN(n2482) );
  INV_X1 U2423 ( .A(n2245), .ZN(n2249) );
  NAND2_X1 U2424 ( .A1(n2484), .A2(n2485), .ZN(n2245) );
  NAND2_X1 U2425 ( .A1(b_14_), .A2(n2486), .ZN(n2485) );
  NAND2_X1 U2426 ( .A1(n2487), .A2(n2218), .ZN(n2486) );
  NAND2_X1 U2427 ( .A1(a_15_), .A2(b_15_), .ZN(n2218) );
  NAND2_X1 U2428 ( .A1(n2488), .A2(b_15_), .ZN(n2484) );
  NOR2_X1 U2429 ( .A1(b_13_), .A2(a_13_), .ZN(n2483) );
  NAND2_X1 U2430 ( .A1(n2489), .A2(n2490), .ZN(n2269) );
  NAND2_X1 U2431 ( .A1(n2281), .A2(n2280), .ZN(n2479) );
  NAND2_X1 U2432 ( .A1(n2491), .A2(n2492), .ZN(n2299) );
  INV_X1 U2433 ( .A(n2493), .ZN(n2300) );
  NAND2_X1 U2434 ( .A1(n2312), .A2(n2311), .ZN(n2475) );
  NOR2_X1 U2435 ( .A1(b_8_), .A2(a_8_), .ZN(n2330) );
  NAND2_X1 U2436 ( .A1(n2343), .A2(n2342), .ZN(n2470) );
  NAND2_X1 U2437 ( .A1(n2494), .A2(n2495), .ZN(n2361) );
  NAND2_X1 U2438 ( .A1(n2374), .A2(n2373), .ZN(n2466) );
  NAND2_X1 U2439 ( .A1(n2496), .A2(n2497), .ZN(n2392) );
  NAND2_X1 U2440 ( .A1(n2411), .A2(n2410), .ZN(n2462) );
  NAND2_X1 U2441 ( .A1(n2498), .A2(n2426), .ZN(n2430) );
  NAND2_X1 U2442 ( .A1(n2499), .A2(n2500), .ZN(n2445) );
  NOR2_X1 U2443 ( .A1(n2177), .A2(n2501), .ZN(Result_15_) );
  XOR2_X1 U2444 ( .A(n2502), .B(n2503), .Z(n2501) );
  NOR2_X1 U2445 ( .A1(n2504), .A2(n2505), .ZN(Result_14_) );
  NAND2_X1 U2446 ( .A1(n2223), .A2(n2506), .ZN(n2505) );
  NOR2_X1 U2447 ( .A1(n2507), .A2(n2508), .ZN(n2504) );
  NOR2_X1 U2448 ( .A1(n2509), .A2(n2503), .ZN(n2507) );
  INV_X1 U2449 ( .A(n2502), .ZN(n2509) );
  NOR2_X1 U2450 ( .A1(n2177), .A2(n2510), .ZN(Result_13_) );
  XNOR2_X1 U2451 ( .A(n2511), .B(n2506), .ZN(n2510) );
  INV_X1 U2452 ( .A(n2512), .ZN(n2506) );
  NAND2_X1 U2453 ( .A1(n2513), .A2(n2514), .ZN(n2511) );
  INV_X1 U2454 ( .A(n2515), .ZN(n2514) );
  NAND2_X1 U2455 ( .A1(n2516), .A2(n2517), .ZN(n2513) );
  NOR2_X1 U2456 ( .A1(n2177), .A2(n2518), .ZN(Result_12_) );
  XNOR2_X1 U2457 ( .A(n2519), .B(n2520), .ZN(n2518) );
  NOR2_X1 U2458 ( .A1(n2177), .A2(n2521), .ZN(Result_11_) );
  XOR2_X1 U2459 ( .A(n2522), .B(n2523), .Z(n2521) );
  NOR2_X1 U2460 ( .A1(n2524), .A2(n2525), .ZN(n2523) );
  NOR2_X1 U2461 ( .A1(n2526), .A2(n2527), .ZN(n2525) );
  NOR2_X1 U2462 ( .A1(n2177), .A2(n2528), .ZN(Result_10_) );
  XNOR2_X1 U2463 ( .A(n2529), .B(n2530), .ZN(n2528) );
  NOR2_X1 U2464 ( .A1(n2177), .A2(n2531), .ZN(Result_0_) );
  NOR2_X1 U2465 ( .A1(n2532), .A2(n2533), .ZN(n2531) );
  NAND2_X1 U2466 ( .A1(n2398), .A2(n2534), .ZN(n2533) );
  INV_X1 U2467 ( .A(n2535), .ZN(n2398) );
  NOR2_X1 U2468 ( .A1(n2536), .A2(n2537), .ZN(n2535) );
  NOR2_X1 U2469 ( .A1(n2238), .A2(n2538), .ZN(n2532) );
  NAND2_X1 U2470 ( .A1(n2397), .A2(n2237), .ZN(n2538) );
  NAND2_X1 U2471 ( .A1(n2539), .A2(n2540), .ZN(n2237) );
  NAND2_X1 U2472 ( .A1(n2209), .A2(n2214), .ZN(n2540) );
  NOR2_X1 U2473 ( .A1(n2541), .A2(n2206), .ZN(n2209) );
  XNOR2_X1 U2474 ( .A(n2542), .B(n2543), .ZN(n2206) );
  INV_X1 U2475 ( .A(n2207), .ZN(n2541) );
  NAND2_X1 U2476 ( .A1(n2544), .A2(n2545), .ZN(n2207) );
  NAND2_X1 U2477 ( .A1(n2199), .A2(n2204), .ZN(n2545) );
  NOR2_X1 U2478 ( .A1(n2546), .A2(n2197), .ZN(n2199) );
  XOR2_X1 U2479 ( .A(n2547), .B(n2548), .Z(n2197) );
  INV_X1 U2480 ( .A(n2196), .ZN(n2546) );
  NAND2_X1 U2481 ( .A1(n2549), .A2(n2550), .ZN(n2196) );
  NAND2_X1 U2482 ( .A1(n2551), .A2(n2194), .ZN(n2550) );
  INV_X1 U2483 ( .A(n2189), .ZN(n2551) );
  NAND2_X1 U2484 ( .A1(n2186), .A2(n2187), .ZN(n2189) );
  XNOR2_X1 U2485 ( .A(n2552), .B(n2553), .ZN(n2187) );
  NAND2_X1 U2486 ( .A1(n2554), .A2(n2555), .ZN(n2186) );
  NAND2_X1 U2487 ( .A1(n2556), .A2(n2184), .ZN(n2555) );
  INV_X1 U2488 ( .A(n2179), .ZN(n2556) );
  NAND2_X1 U2489 ( .A1(n2529), .A2(n2530), .ZN(n2179) );
  XOR2_X1 U2490 ( .A(n2557), .B(n2558), .Z(n2530) );
  NAND2_X1 U2491 ( .A1(n2559), .A2(n2560), .ZN(n2529) );
  NAND2_X1 U2492 ( .A1(n2561), .A2(n2527), .ZN(n2560) );
  INV_X1 U2493 ( .A(n2522), .ZN(n2561) );
  NAND2_X1 U2494 ( .A1(n2520), .A2(n2519), .ZN(n2522) );
  NAND2_X1 U2495 ( .A1(n2562), .A2(n2563), .ZN(n2519) );
  NAND2_X1 U2496 ( .A1(n2512), .A2(n2564), .ZN(n2563) );
  NOR2_X1 U2497 ( .A1(n2565), .A2(n2503), .ZN(n2512) );
  XOR2_X1 U2498 ( .A(n2566), .B(n2567), .Z(n2503) );
  XOR2_X1 U2499 ( .A(n2568), .B(n2569), .Z(n2567) );
  NAND2_X1 U2500 ( .A1(a_0_), .A2(b_14_), .ZN(n2569) );
  NAND2_X1 U2501 ( .A1(n2502), .A2(n2508), .ZN(n2565) );
  XOR2_X1 U2502 ( .A(n2570), .B(n2571), .Z(n2508) );
  NAND2_X1 U2503 ( .A1(n2572), .A2(n2573), .ZN(n2502) );
  NAND2_X1 U2504 ( .A1(n2574), .A2(a_0_), .ZN(n2573) );
  NOR2_X1 U2505 ( .A1(n2575), .A2(n2229), .ZN(n2574) );
  NOR2_X1 U2506 ( .A1(n2451), .A2(n2453), .ZN(n2575) );
  NAND2_X1 U2507 ( .A1(n2451), .A2(n2453), .ZN(n2572) );
  NAND2_X1 U2508 ( .A1(n2576), .A2(n2577), .ZN(n2453) );
  NAND2_X1 U2509 ( .A1(n2578), .A2(b_15_), .ZN(n2577) );
  NOR2_X1 U2510 ( .A1(n2579), .A2(n2500), .ZN(n2578) );
  NOR2_X1 U2511 ( .A1(n2435), .A2(n2437), .ZN(n2579) );
  NAND2_X1 U2512 ( .A1(n2435), .A2(n2437), .ZN(n2576) );
  NAND2_X1 U2513 ( .A1(n2580), .A2(n2581), .ZN(n2437) );
  NAND2_X1 U2514 ( .A1(n2582), .A2(a_2_), .ZN(n2581) );
  NOR2_X1 U2515 ( .A1(n2583), .A2(n2229), .ZN(n2582) );
  NOR2_X1 U2516 ( .A1(n2423), .A2(n2424), .ZN(n2583) );
  NAND2_X1 U2517 ( .A1(n2423), .A2(n2424), .ZN(n2580) );
  NAND2_X1 U2518 ( .A1(n2417), .A2(n2584), .ZN(n2424) );
  NAND2_X1 U2519 ( .A1(n2416), .A2(n2418), .ZN(n2584) );
  NAND2_X1 U2520 ( .A1(n2585), .A2(n2586), .ZN(n2418) );
  NAND2_X1 U2521 ( .A1(a_3_), .A2(b_15_), .ZN(n2585) );
  XNOR2_X1 U2522 ( .A(n2587), .B(n2588), .ZN(n2416) );
  XOR2_X1 U2523 ( .A(n2589), .B(n2590), .Z(n2588) );
  NAND2_X1 U2524 ( .A1(a_4_), .A2(b_14_), .ZN(n2590) );
  INV_X1 U2525 ( .A(n2591), .ZN(n2417) );
  NOR2_X1 U2526 ( .A1(n2586), .A2(n2410), .ZN(n2591) );
  NAND2_X1 U2527 ( .A1(n2592), .A2(n2593), .ZN(n2586) );
  NAND2_X1 U2528 ( .A1(n2594), .A2(n2387), .ZN(n2593) );
  NAND2_X1 U2529 ( .A1(a_4_), .A2(b_15_), .ZN(n2387) );
  NAND2_X1 U2530 ( .A1(n2385), .A2(n2388), .ZN(n2594) );
  INV_X1 U2531 ( .A(n2595), .ZN(n2592) );
  NOR2_X1 U2532 ( .A1(n2388), .A2(n2385), .ZN(n2595) );
  XNOR2_X1 U2533 ( .A(n2596), .B(n2597), .ZN(n2385) );
  XOR2_X1 U2534 ( .A(n2598), .B(n2599), .Z(n2597) );
  NAND2_X1 U2535 ( .A1(a_5_), .A2(b_14_), .ZN(n2599) );
  NAND2_X1 U2536 ( .A1(n2380), .A2(n2600), .ZN(n2388) );
  NAND2_X1 U2537 ( .A1(n2379), .A2(n2381), .ZN(n2600) );
  NAND2_X1 U2538 ( .A1(n2601), .A2(n2602), .ZN(n2381) );
  NAND2_X1 U2539 ( .A1(a_5_), .A2(b_15_), .ZN(n2601) );
  XNOR2_X1 U2540 ( .A(n2603), .B(n2604), .ZN(n2379) );
  XOR2_X1 U2541 ( .A(n2605), .B(n2606), .Z(n2604) );
  NAND2_X1 U2542 ( .A1(a_6_), .A2(b_14_), .ZN(n2606) );
  INV_X1 U2543 ( .A(n2607), .ZN(n2380) );
  NOR2_X1 U2544 ( .A1(n2602), .A2(n2373), .ZN(n2607) );
  NAND2_X1 U2545 ( .A1(n2608), .A2(n2609), .ZN(n2602) );
  NAND2_X1 U2546 ( .A1(n2610), .A2(n2356), .ZN(n2609) );
  NAND2_X1 U2547 ( .A1(a_6_), .A2(b_15_), .ZN(n2356) );
  NAND2_X1 U2548 ( .A1(n2354), .A2(n2357), .ZN(n2610) );
  INV_X1 U2549 ( .A(n2611), .ZN(n2608) );
  NOR2_X1 U2550 ( .A1(n2357), .A2(n2354), .ZN(n2611) );
  XNOR2_X1 U2551 ( .A(n2612), .B(n2613), .ZN(n2354) );
  XOR2_X1 U2552 ( .A(n2614), .B(n2615), .Z(n2613) );
  NAND2_X1 U2553 ( .A1(a_7_), .A2(b_14_), .ZN(n2615) );
  NAND2_X1 U2554 ( .A1(n2349), .A2(n2616), .ZN(n2357) );
  NAND2_X1 U2555 ( .A1(n2348), .A2(n2350), .ZN(n2616) );
  NAND2_X1 U2556 ( .A1(n2617), .A2(n2618), .ZN(n2350) );
  NAND2_X1 U2557 ( .A1(a_7_), .A2(b_15_), .ZN(n2617) );
  XNOR2_X1 U2558 ( .A(n2619), .B(n2620), .ZN(n2348) );
  XOR2_X1 U2559 ( .A(n2621), .B(n2622), .Z(n2620) );
  INV_X1 U2560 ( .A(n2623), .ZN(n2349) );
  NOR2_X1 U2561 ( .A1(n2618), .A2(n2342), .ZN(n2623) );
  NAND2_X1 U2562 ( .A1(n2624), .A2(n2625), .ZN(n2618) );
  NAND2_X1 U2563 ( .A1(n2626), .A2(n2325), .ZN(n2625) );
  NAND2_X1 U2564 ( .A1(a_8_), .A2(b_15_), .ZN(n2325) );
  NAND2_X1 U2565 ( .A1(n2323), .A2(n2326), .ZN(n2626) );
  INV_X1 U2566 ( .A(n2627), .ZN(n2624) );
  NOR2_X1 U2567 ( .A1(n2326), .A2(n2323), .ZN(n2627) );
  XNOR2_X1 U2568 ( .A(n2628), .B(n2629), .ZN(n2323) );
  XNOR2_X1 U2569 ( .A(n2630), .B(n2631), .ZN(n2629) );
  NAND2_X1 U2570 ( .A1(n2318), .A2(n2632), .ZN(n2326) );
  NAND2_X1 U2571 ( .A1(n2317), .A2(n2319), .ZN(n2632) );
  NAND2_X1 U2572 ( .A1(n2633), .A2(n2634), .ZN(n2319) );
  NAND2_X1 U2573 ( .A1(a_9_), .A2(b_15_), .ZN(n2633) );
  XNOR2_X1 U2574 ( .A(n2635), .B(n2636), .ZN(n2317) );
  XOR2_X1 U2575 ( .A(n2637), .B(n2638), .Z(n2635) );
  INV_X1 U2576 ( .A(n2639), .ZN(n2318) );
  NOR2_X1 U2577 ( .A1(n2634), .A2(n2311), .ZN(n2639) );
  NAND2_X1 U2578 ( .A1(n2640), .A2(n2641), .ZN(n2634) );
  NAND2_X1 U2579 ( .A1(n2642), .A2(n2295), .ZN(n2641) );
  NAND2_X1 U2580 ( .A1(a_10_), .A2(b_15_), .ZN(n2295) );
  NAND2_X1 U2581 ( .A1(n2292), .A2(n2294), .ZN(n2642) );
  INV_X1 U2582 ( .A(n2643), .ZN(n2640) );
  NOR2_X1 U2583 ( .A1(n2294), .A2(n2292), .ZN(n2643) );
  XNOR2_X1 U2584 ( .A(n2644), .B(n2645), .ZN(n2292) );
  NAND2_X1 U2585 ( .A1(n2646), .A2(n2647), .ZN(n2644) );
  NAND2_X1 U2586 ( .A1(n2287), .A2(n2648), .ZN(n2294) );
  NAND2_X1 U2587 ( .A1(n2286), .A2(n2288), .ZN(n2648) );
  NAND2_X1 U2588 ( .A1(n2649), .A2(n2650), .ZN(n2288) );
  NAND2_X1 U2589 ( .A1(a_11_), .A2(b_15_), .ZN(n2650) );
  XNOR2_X1 U2590 ( .A(n2651), .B(n2652), .ZN(n2286) );
  XOR2_X1 U2591 ( .A(n2653), .B(n2654), .Z(n2652) );
  NAND2_X1 U2592 ( .A1(a_12_), .A2(b_14_), .ZN(n2654) );
  NAND2_X1 U2593 ( .A1(a_11_), .A2(n2655), .ZN(n2287) );
  INV_X1 U2594 ( .A(n2649), .ZN(n2655) );
  NOR2_X1 U2595 ( .A1(n2656), .A2(n2657), .ZN(n2649) );
  INV_X1 U2596 ( .A(n2658), .ZN(n2657) );
  NAND2_X1 U2597 ( .A1(n2264), .A2(n2659), .ZN(n2658) );
  NAND2_X1 U2598 ( .A1(n2262), .A2(n2263), .ZN(n2659) );
  NOR2_X1 U2599 ( .A1(n2490), .A2(n2229), .ZN(n2264) );
  NOR2_X1 U2600 ( .A1(n2263), .A2(n2262), .ZN(n2656) );
  XNOR2_X1 U2601 ( .A(n2660), .B(n2661), .ZN(n2262) );
  XOR2_X1 U2602 ( .A(n2662), .B(n2663), .Z(n2661) );
  NAND2_X1 U2603 ( .A1(a_13_), .A2(b_14_), .ZN(n2660) );
  NAND2_X1 U2604 ( .A1(n2664), .A2(n2665), .ZN(n2263) );
  NAND2_X1 U2605 ( .A1(n2666), .A2(n2256), .ZN(n2665) );
  NAND2_X1 U2606 ( .A1(a_13_), .A2(b_15_), .ZN(n2256) );
  NAND2_X1 U2607 ( .A1(n2667), .A2(n2257), .ZN(n2666) );
  INV_X1 U2608 ( .A(n2668), .ZN(n2664) );
  NOR2_X1 U2609 ( .A1(n2257), .A2(n2667), .ZN(n2668) );
  INV_X1 U2610 ( .A(n2254), .ZN(n2667) );
  NAND2_X1 U2611 ( .A1(n2669), .A2(n2488), .ZN(n2254) );
  NOR2_X1 U2612 ( .A1(n2229), .A2(n2233), .ZN(n2669) );
  NAND2_X1 U2613 ( .A1(n2670), .A2(n2671), .ZN(n2257) );
  NAND2_X1 U2614 ( .A1(b_13_), .A2(n2672), .ZN(n2671) );
  NAND2_X1 U2615 ( .A1(n2227), .A2(n2673), .ZN(n2672) );
  NAND2_X1 U2616 ( .A1(a_15_), .A2(n2233), .ZN(n2673) );
  NAND2_X1 U2617 ( .A1(b_14_), .A2(n2674), .ZN(n2670) );
  NAND2_X1 U2618 ( .A1(n2231), .A2(n2675), .ZN(n2674) );
  NAND2_X1 U2619 ( .A1(a_14_), .A2(n2250), .ZN(n2675) );
  XNOR2_X1 U2620 ( .A(n2676), .B(n2677), .ZN(n2423) );
  XOR2_X1 U2621 ( .A(n2678), .B(n2679), .Z(n2677) );
  NAND2_X1 U2622 ( .A1(a_3_), .A2(b_14_), .ZN(n2679) );
  XNOR2_X1 U2623 ( .A(n2680), .B(n2681), .ZN(n2435) );
  XOR2_X1 U2624 ( .A(n2682), .B(n2683), .Z(n2681) );
  NAND2_X1 U2625 ( .A1(a_2_), .A2(b_14_), .ZN(n2683) );
  XNOR2_X1 U2626 ( .A(n2684), .B(n2685), .ZN(n2451) );
  XOR2_X1 U2627 ( .A(n2686), .B(n2687), .Z(n2685) );
  NAND2_X1 U2628 ( .A1(b_14_), .A2(a_1_), .ZN(n2687) );
  NOR2_X1 U2629 ( .A1(n2515), .A2(n2688), .ZN(n2562) );
  NOR2_X1 U2630 ( .A1(n2517), .A2(n2516), .ZN(n2515) );
  INV_X1 U2631 ( .A(n2564), .ZN(n2516) );
  NOR2_X1 U2632 ( .A1(n2688), .A2(n2689), .ZN(n2564) );
  NOR2_X1 U2633 ( .A1(n2690), .A2(n2691), .ZN(n2689) );
  INV_X1 U2634 ( .A(n2692), .ZN(n2688) );
  NAND2_X1 U2635 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  NAND2_X1 U2636 ( .A1(n2693), .A2(n2694), .ZN(n2690) );
  NAND2_X1 U2637 ( .A1(n2695), .A2(n2696), .ZN(n2694) );
  XNOR2_X1 U2638 ( .A(n2697), .B(n2698), .ZN(n2691) );
  NAND2_X1 U2639 ( .A1(n2699), .A2(n2700), .ZN(n2697) );
  NAND2_X1 U2640 ( .A1(n2571), .A2(n2570), .ZN(n2517) );
  NAND2_X1 U2641 ( .A1(n2701), .A2(n2702), .ZN(n2570) );
  NAND2_X1 U2642 ( .A1(n2703), .A2(a_0_), .ZN(n2702) );
  NOR2_X1 U2643 ( .A1(n2704), .A2(n2233), .ZN(n2703) );
  NOR2_X1 U2644 ( .A1(n2566), .A2(n2568), .ZN(n2704) );
  NAND2_X1 U2645 ( .A1(n2566), .A2(n2568), .ZN(n2701) );
  NAND2_X1 U2646 ( .A1(n2705), .A2(n2706), .ZN(n2568) );
  NAND2_X1 U2647 ( .A1(n2707), .A2(b_14_), .ZN(n2706) );
  NOR2_X1 U2648 ( .A1(n2708), .A2(n2500), .ZN(n2707) );
  NOR2_X1 U2649 ( .A1(n2684), .A2(n2686), .ZN(n2708) );
  NAND2_X1 U2650 ( .A1(n2684), .A2(n2686), .ZN(n2705) );
  NAND2_X1 U2651 ( .A1(n2709), .A2(n2710), .ZN(n2686) );
  NAND2_X1 U2652 ( .A1(n2711), .A2(a_2_), .ZN(n2710) );
  NOR2_X1 U2653 ( .A1(n2712), .A2(n2233), .ZN(n2711) );
  NOR2_X1 U2654 ( .A1(n2680), .A2(n2682), .ZN(n2712) );
  NAND2_X1 U2655 ( .A1(n2680), .A2(n2682), .ZN(n2709) );
  NAND2_X1 U2656 ( .A1(n2713), .A2(n2714), .ZN(n2682) );
  NAND2_X1 U2657 ( .A1(n2715), .A2(a_3_), .ZN(n2714) );
  NOR2_X1 U2658 ( .A1(n2716), .A2(n2233), .ZN(n2715) );
  NOR2_X1 U2659 ( .A1(n2676), .A2(n2678), .ZN(n2716) );
  NAND2_X1 U2660 ( .A1(n2676), .A2(n2678), .ZN(n2713) );
  NAND2_X1 U2661 ( .A1(n2717), .A2(n2718), .ZN(n2678) );
  NAND2_X1 U2662 ( .A1(n2719), .A2(a_4_), .ZN(n2718) );
  NOR2_X1 U2663 ( .A1(n2720), .A2(n2233), .ZN(n2719) );
  NOR2_X1 U2664 ( .A1(n2587), .A2(n2589), .ZN(n2720) );
  NAND2_X1 U2665 ( .A1(n2587), .A2(n2589), .ZN(n2717) );
  NAND2_X1 U2666 ( .A1(n2721), .A2(n2722), .ZN(n2589) );
  NAND2_X1 U2667 ( .A1(n2723), .A2(a_5_), .ZN(n2722) );
  NOR2_X1 U2668 ( .A1(n2724), .A2(n2233), .ZN(n2723) );
  NOR2_X1 U2669 ( .A1(n2596), .A2(n2598), .ZN(n2724) );
  NAND2_X1 U2670 ( .A1(n2596), .A2(n2598), .ZN(n2721) );
  NAND2_X1 U2671 ( .A1(n2725), .A2(n2726), .ZN(n2598) );
  NAND2_X1 U2672 ( .A1(n2727), .A2(a_6_), .ZN(n2726) );
  NOR2_X1 U2673 ( .A1(n2728), .A2(n2233), .ZN(n2727) );
  NOR2_X1 U2674 ( .A1(n2603), .A2(n2605), .ZN(n2728) );
  NAND2_X1 U2675 ( .A1(n2603), .A2(n2605), .ZN(n2725) );
  NAND2_X1 U2676 ( .A1(n2729), .A2(n2730), .ZN(n2605) );
  NAND2_X1 U2677 ( .A1(n2731), .A2(a_7_), .ZN(n2730) );
  NOR2_X1 U2678 ( .A1(n2732), .A2(n2233), .ZN(n2731) );
  NOR2_X1 U2679 ( .A1(n2612), .A2(n2614), .ZN(n2732) );
  NAND2_X1 U2680 ( .A1(n2612), .A2(n2614), .ZN(n2729) );
  NAND2_X1 U2681 ( .A1(n2733), .A2(n2734), .ZN(n2614) );
  NAND2_X1 U2682 ( .A1(n2735), .A2(n2736), .ZN(n2734) );
  INV_X1 U2683 ( .A(n2737), .ZN(n2736) );
  NOR2_X1 U2684 ( .A1(n2621), .A2(n2619), .ZN(n2737) );
  INV_X1 U2685 ( .A(n2622), .ZN(n2735) );
  NAND2_X1 U2686 ( .A1(a_8_), .A2(b_14_), .ZN(n2622) );
  NAND2_X1 U2687 ( .A1(n2619), .A2(n2621), .ZN(n2733) );
  NAND2_X1 U2688 ( .A1(n2738), .A2(n2739), .ZN(n2621) );
  NAND2_X1 U2689 ( .A1(n2631), .A2(n2740), .ZN(n2739) );
  NAND2_X1 U2690 ( .A1(n2628), .A2(n2630), .ZN(n2740) );
  NOR2_X1 U2691 ( .A1(n2311), .A2(n2233), .ZN(n2631) );
  INV_X1 U2692 ( .A(n2741), .ZN(n2738) );
  NOR2_X1 U2693 ( .A1(n2630), .A2(n2628), .ZN(n2741) );
  XOR2_X1 U2694 ( .A(n2742), .B(n2743), .Z(n2628) );
  XOR2_X1 U2695 ( .A(n2744), .B(n2745), .Z(n2742) );
  NAND2_X1 U2696 ( .A1(n2746), .A2(n2747), .ZN(n2630) );
  NAND2_X1 U2697 ( .A1(n2636), .A2(n2748), .ZN(n2747) );
  NAND2_X1 U2698 ( .A1(n2638), .A2(n2637), .ZN(n2748) );
  XOR2_X1 U2699 ( .A(n2749), .B(n2750), .Z(n2636) );
  XNOR2_X1 U2700 ( .A(n2751), .B(n2752), .ZN(n2749) );
  INV_X1 U2701 ( .A(n2753), .ZN(n2746) );
  NOR2_X1 U2702 ( .A1(n2637), .A2(n2638), .ZN(n2753) );
  NOR2_X1 U2703 ( .A1(n2492), .A2(n2233), .ZN(n2638) );
  NAND2_X1 U2704 ( .A1(n2646), .A2(n2754), .ZN(n2637) );
  NAND2_X1 U2705 ( .A1(n2645), .A2(n2647), .ZN(n2754) );
  NAND2_X1 U2706 ( .A1(n2755), .A2(n2756), .ZN(n2647) );
  NAND2_X1 U2707 ( .A1(a_11_), .A2(b_14_), .ZN(n2756) );
  INV_X1 U2708 ( .A(n2757), .ZN(n2755) );
  XOR2_X1 U2709 ( .A(n2758), .B(n2759), .Z(n2645) );
  XOR2_X1 U2710 ( .A(n2760), .B(n2761), .Z(n2758) );
  NAND2_X1 U2711 ( .A1(a_11_), .A2(n2757), .ZN(n2646) );
  NAND2_X1 U2712 ( .A1(n2762), .A2(n2763), .ZN(n2757) );
  NAND2_X1 U2713 ( .A1(n2764), .A2(a_12_), .ZN(n2763) );
  NOR2_X1 U2714 ( .A1(n2765), .A2(n2233), .ZN(n2764) );
  NOR2_X1 U2715 ( .A1(n2651), .A2(n2653), .ZN(n2765) );
  NAND2_X1 U2716 ( .A1(n2651), .A2(n2653), .ZN(n2762) );
  NAND2_X1 U2717 ( .A1(n2766), .A2(n2767), .ZN(n2653) );
  NAND2_X1 U2718 ( .A1(n2768), .A2(a_13_), .ZN(n2767) );
  NOR2_X1 U2719 ( .A1(n2769), .A2(n2233), .ZN(n2768) );
  NOR2_X1 U2720 ( .A1(n2770), .A2(n2663), .ZN(n2769) );
  NAND2_X1 U2721 ( .A1(n2770), .A2(n2663), .ZN(n2766) );
  NAND2_X1 U2722 ( .A1(n2771), .A2(n2772), .ZN(n2663) );
  NAND2_X1 U2723 ( .A1(b_12_), .A2(n2773), .ZN(n2772) );
  NAND2_X1 U2724 ( .A1(n2227), .A2(n2774), .ZN(n2773) );
  NAND2_X1 U2725 ( .A1(a_15_), .A2(n2250), .ZN(n2774) );
  NAND2_X1 U2726 ( .A1(b_13_), .A2(n2775), .ZN(n2771) );
  NAND2_X1 U2727 ( .A1(n2231), .A2(n2776), .ZN(n2775) );
  NAND2_X1 U2728 ( .A1(a_14_), .A2(n2489), .ZN(n2776) );
  INV_X1 U2729 ( .A(n2662), .ZN(n2770) );
  NAND2_X1 U2730 ( .A1(n2777), .A2(n2488), .ZN(n2662) );
  NOR2_X1 U2731 ( .A1(n2233), .A2(n2250), .ZN(n2777) );
  XNOR2_X1 U2732 ( .A(n2244), .B(n2778), .ZN(n2651) );
  XOR2_X1 U2733 ( .A(n2779), .B(n2780), .Z(n2778) );
  XNOR2_X1 U2734 ( .A(n2781), .B(n2782), .ZN(n2619) );
  NAND2_X1 U2735 ( .A1(n2783), .A2(n2784), .ZN(n2781) );
  XNOR2_X1 U2736 ( .A(n2785), .B(n2786), .ZN(n2612) );
  NAND2_X1 U2737 ( .A1(n2787), .A2(n2788), .ZN(n2785) );
  XNOR2_X1 U2738 ( .A(n2789), .B(n2790), .ZN(n2603) );
  NAND2_X1 U2739 ( .A1(n2791), .A2(n2792), .ZN(n2789) );
  XNOR2_X1 U2740 ( .A(n2793), .B(n2794), .ZN(n2596) );
  XOR2_X1 U2741 ( .A(n2795), .B(n2796), .Z(n2794) );
  NAND2_X1 U2742 ( .A1(a_6_), .A2(b_13_), .ZN(n2796) );
  XNOR2_X1 U2743 ( .A(n2797), .B(n2798), .ZN(n2587) );
  NAND2_X1 U2744 ( .A1(n2799), .A2(n2800), .ZN(n2797) );
  XOR2_X1 U2745 ( .A(n2801), .B(n2802), .Z(n2676) );
  XOR2_X1 U2746 ( .A(n2803), .B(n2804), .Z(n2801) );
  NOR2_X1 U2747 ( .A1(n2250), .A2(n2497), .ZN(n2804) );
  XNOR2_X1 U2748 ( .A(n2805), .B(n2806), .ZN(n2680) );
  NAND2_X1 U2749 ( .A1(n2807), .A2(n2808), .ZN(n2805) );
  XNOR2_X1 U2750 ( .A(n2809), .B(n2810), .ZN(n2684) );
  XOR2_X1 U2751 ( .A(n2811), .B(n2812), .Z(n2809) );
  XNOR2_X1 U2752 ( .A(n2813), .B(n2814), .ZN(n2566) );
  NAND2_X1 U2753 ( .A1(n2815), .A2(n2816), .ZN(n2813) );
  XNOR2_X1 U2754 ( .A(n2817), .B(n2695), .ZN(n2571) );
  XNOR2_X1 U2755 ( .A(n2818), .B(n2819), .ZN(n2695) );
  XOR2_X1 U2756 ( .A(n2820), .B(n2821), .Z(n2819) );
  NAND2_X1 U2757 ( .A1(b_12_), .A2(a_1_), .ZN(n2821) );
  NAND2_X1 U2758 ( .A1(n2693), .A2(n2696), .ZN(n2817) );
  NAND2_X1 U2759 ( .A1(n2822), .A2(n2823), .ZN(n2696) );
  NAND2_X1 U2760 ( .A1(a_0_), .A2(b_13_), .ZN(n2823) );
  INV_X1 U2761 ( .A(n2824), .ZN(n2822) );
  NAND2_X1 U2762 ( .A1(a_0_), .A2(n2824), .ZN(n2693) );
  NAND2_X1 U2763 ( .A1(n2815), .A2(n2825), .ZN(n2824) );
  NAND2_X1 U2764 ( .A1(n2814), .A2(n2816), .ZN(n2825) );
  NAND2_X1 U2765 ( .A1(n2826), .A2(n2827), .ZN(n2816) );
  NAND2_X1 U2766 ( .A1(b_13_), .A2(a_1_), .ZN(n2827) );
  XNOR2_X1 U2767 ( .A(n2828), .B(n2829), .ZN(n2814) );
  XOR2_X1 U2768 ( .A(n2830), .B(n2831), .Z(n2829) );
  NAND2_X1 U2769 ( .A1(a_2_), .A2(b_12_), .ZN(n2831) );
  INV_X1 U2770 ( .A(n2832), .ZN(n2815) );
  NOR2_X1 U2771 ( .A1(n2826), .A2(n2500), .ZN(n2832) );
  NAND2_X1 U2772 ( .A1(n2833), .A2(n2834), .ZN(n2826) );
  NAND2_X1 U2773 ( .A1(n2810), .A2(n2835), .ZN(n2834) );
  NAND2_X1 U2774 ( .A1(n2812), .A2(n2811), .ZN(n2835) );
  XOR2_X1 U2775 ( .A(n2836), .B(n2837), .Z(n2810) );
  XOR2_X1 U2776 ( .A(n2838), .B(n2839), .Z(n2837) );
  NAND2_X1 U2777 ( .A1(a_3_), .A2(b_12_), .ZN(n2839) );
  INV_X1 U2778 ( .A(n2840), .ZN(n2833) );
  NOR2_X1 U2779 ( .A1(n2811), .A2(n2812), .ZN(n2840) );
  NOR2_X1 U2780 ( .A1(n2426), .A2(n2250), .ZN(n2812) );
  NAND2_X1 U2781 ( .A1(n2807), .A2(n2841), .ZN(n2811) );
  NAND2_X1 U2782 ( .A1(n2806), .A2(n2808), .ZN(n2841) );
  NAND2_X1 U2783 ( .A1(n2842), .A2(n2843), .ZN(n2808) );
  NAND2_X1 U2784 ( .A1(a_3_), .A2(b_13_), .ZN(n2843) );
  INV_X1 U2785 ( .A(n2844), .ZN(n2842) );
  XNOR2_X1 U2786 ( .A(n2845), .B(n2846), .ZN(n2806) );
  XOR2_X1 U2787 ( .A(n2847), .B(n2848), .Z(n2846) );
  NAND2_X1 U2788 ( .A1(a_4_), .A2(b_12_), .ZN(n2848) );
  NAND2_X1 U2789 ( .A1(a_3_), .A2(n2844), .ZN(n2807) );
  NAND2_X1 U2790 ( .A1(n2849), .A2(n2850), .ZN(n2844) );
  NAND2_X1 U2791 ( .A1(n2851), .A2(a_4_), .ZN(n2850) );
  NOR2_X1 U2792 ( .A1(n2852), .A2(n2250), .ZN(n2851) );
  NOR2_X1 U2793 ( .A1(n2802), .A2(n2803), .ZN(n2852) );
  NAND2_X1 U2794 ( .A1(n2802), .A2(n2803), .ZN(n2849) );
  NAND2_X1 U2795 ( .A1(n2799), .A2(n2853), .ZN(n2803) );
  NAND2_X1 U2796 ( .A1(n2798), .A2(n2800), .ZN(n2853) );
  NAND2_X1 U2797 ( .A1(n2854), .A2(n2855), .ZN(n2800) );
  NAND2_X1 U2798 ( .A1(a_5_), .A2(b_13_), .ZN(n2855) );
  INV_X1 U2799 ( .A(n2856), .ZN(n2854) );
  XOR2_X1 U2800 ( .A(n2857), .B(n2858), .Z(n2798) );
  XOR2_X1 U2801 ( .A(n2859), .B(n2860), .Z(n2857) );
  NOR2_X1 U2802 ( .A1(n2489), .A2(n2495), .ZN(n2860) );
  NAND2_X1 U2803 ( .A1(a_5_), .A2(n2856), .ZN(n2799) );
  NAND2_X1 U2804 ( .A1(n2861), .A2(n2862), .ZN(n2856) );
  NAND2_X1 U2805 ( .A1(n2863), .A2(a_6_), .ZN(n2862) );
  NOR2_X1 U2806 ( .A1(n2864), .A2(n2250), .ZN(n2863) );
  NOR2_X1 U2807 ( .A1(n2793), .A2(n2795), .ZN(n2864) );
  NAND2_X1 U2808 ( .A1(n2793), .A2(n2795), .ZN(n2861) );
  NAND2_X1 U2809 ( .A1(n2791), .A2(n2865), .ZN(n2795) );
  NAND2_X1 U2810 ( .A1(n2790), .A2(n2792), .ZN(n2865) );
  NAND2_X1 U2811 ( .A1(n2866), .A2(n2867), .ZN(n2792) );
  NAND2_X1 U2812 ( .A1(a_7_), .A2(b_13_), .ZN(n2867) );
  INV_X1 U2813 ( .A(n2868), .ZN(n2866) );
  XNOR2_X1 U2814 ( .A(n2869), .B(n2870), .ZN(n2790) );
  XOR2_X1 U2815 ( .A(n2871), .B(n2872), .Z(n2870) );
  NAND2_X1 U2816 ( .A1(a_7_), .A2(n2868), .ZN(n2791) );
  NAND2_X1 U2817 ( .A1(n2787), .A2(n2873), .ZN(n2868) );
  NAND2_X1 U2818 ( .A1(n2786), .A2(n2788), .ZN(n2873) );
  NAND2_X1 U2819 ( .A1(n2874), .A2(n2875), .ZN(n2788) );
  NAND2_X1 U2820 ( .A1(a_8_), .A2(b_13_), .ZN(n2875) );
  INV_X1 U2821 ( .A(n2876), .ZN(n2874) );
  XNOR2_X1 U2822 ( .A(n2877), .B(n2878), .ZN(n2786) );
  XNOR2_X1 U2823 ( .A(n2879), .B(n2880), .ZN(n2878) );
  NAND2_X1 U2824 ( .A1(a_8_), .A2(n2876), .ZN(n2787) );
  NAND2_X1 U2825 ( .A1(n2783), .A2(n2881), .ZN(n2876) );
  NAND2_X1 U2826 ( .A1(n2782), .A2(n2784), .ZN(n2881) );
  NAND2_X1 U2827 ( .A1(n2882), .A2(n2883), .ZN(n2784) );
  NAND2_X1 U2828 ( .A1(a_9_), .A2(b_13_), .ZN(n2882) );
  XNOR2_X1 U2829 ( .A(n2884), .B(n2885), .ZN(n2782) );
  XOR2_X1 U2830 ( .A(n2886), .B(n2887), .Z(n2884) );
  INV_X1 U2831 ( .A(n2888), .ZN(n2783) );
  NOR2_X1 U2832 ( .A1(n2883), .A2(n2311), .ZN(n2888) );
  NAND2_X1 U2833 ( .A1(n2889), .A2(n2890), .ZN(n2883) );
  NAND2_X1 U2834 ( .A1(n2743), .A2(n2891), .ZN(n2890) );
  NAND2_X1 U2835 ( .A1(n2745), .A2(n2744), .ZN(n2891) );
  XOR2_X1 U2836 ( .A(n2892), .B(n2893), .Z(n2743) );
  NAND2_X1 U2837 ( .A1(n2894), .A2(n2895), .ZN(n2892) );
  INV_X1 U2838 ( .A(n2896), .ZN(n2889) );
  NOR2_X1 U2839 ( .A1(n2744), .A2(n2745), .ZN(n2896) );
  NOR2_X1 U2840 ( .A1(n2492), .A2(n2250), .ZN(n2745) );
  NAND2_X1 U2841 ( .A1(n2897), .A2(n2898), .ZN(n2744) );
  NAND2_X1 U2842 ( .A1(n2752), .A2(n2899), .ZN(n2898) );
  NAND2_X1 U2843 ( .A1(n2751), .A2(n2750), .ZN(n2899) );
  NOR2_X1 U2844 ( .A1(n2280), .A2(n2250), .ZN(n2752) );
  INV_X1 U2845 ( .A(n2900), .ZN(n2897) );
  NOR2_X1 U2846 ( .A1(n2750), .A2(n2751), .ZN(n2900) );
  NOR2_X1 U2847 ( .A1(n2901), .A2(n2902), .ZN(n2751) );
  INV_X1 U2848 ( .A(n2903), .ZN(n2902) );
  NAND2_X1 U2849 ( .A1(n2761), .A2(n2904), .ZN(n2903) );
  NAND2_X1 U2850 ( .A1(n2759), .A2(n2760), .ZN(n2904) );
  NOR2_X1 U2851 ( .A1(n2490), .A2(n2250), .ZN(n2761) );
  NOR2_X1 U2852 ( .A1(n2760), .A2(n2759), .ZN(n2901) );
  XOR2_X1 U2853 ( .A(n2905), .B(n2906), .Z(n2759) );
  XOR2_X1 U2854 ( .A(n2907), .B(n2908), .Z(n2906) );
  NAND2_X1 U2855 ( .A1(n2909), .A2(n2910), .ZN(n2760) );
  NAND2_X1 U2856 ( .A1(n2911), .A2(n2779), .ZN(n2910) );
  NAND2_X1 U2857 ( .A1(n2912), .A2(n2488), .ZN(n2779) );
  NOR2_X1 U2858 ( .A1(n2250), .A2(n2489), .ZN(n2912) );
  NAND2_X1 U2859 ( .A1(n2244), .A2(n2780), .ZN(n2911) );
  INV_X1 U2860 ( .A(n2913), .ZN(n2909) );
  NOR2_X1 U2861 ( .A1(n2780), .A2(n2244), .ZN(n2913) );
  NOR2_X1 U2862 ( .A1(n2252), .A2(n2250), .ZN(n2244) );
  NAND2_X1 U2863 ( .A1(n2914), .A2(n2915), .ZN(n2780) );
  NAND2_X1 U2864 ( .A1(b_11_), .A2(n2916), .ZN(n2915) );
  NAND2_X1 U2865 ( .A1(n2227), .A2(n2917), .ZN(n2916) );
  NAND2_X1 U2866 ( .A1(a_15_), .A2(n2489), .ZN(n2917) );
  NAND2_X1 U2867 ( .A1(b_12_), .A2(n2918), .ZN(n2914) );
  NAND2_X1 U2868 ( .A1(n2231), .A2(n2919), .ZN(n2918) );
  NAND2_X1 U2869 ( .A1(a_14_), .A2(n2281), .ZN(n2919) );
  XOR2_X1 U2870 ( .A(n2920), .B(n2921), .Z(n2750) );
  XOR2_X1 U2871 ( .A(n2268), .B(n2922), .Z(n2920) );
  XOR2_X1 U2872 ( .A(n2923), .B(n2924), .Z(n2793) );
  XNOR2_X1 U2873 ( .A(n2925), .B(n2926), .ZN(n2923) );
  NAND2_X1 U2874 ( .A1(a_7_), .A2(b_12_), .ZN(n2925) );
  XNOR2_X1 U2875 ( .A(n2927), .B(n2928), .ZN(n2802) );
  XOR2_X1 U2876 ( .A(n2929), .B(n2930), .Z(n2928) );
  NAND2_X1 U2877 ( .A1(a_5_), .A2(b_12_), .ZN(n2930) );
  XNOR2_X1 U2878 ( .A(n2931), .B(n2932), .ZN(n2520) );
  NOR2_X1 U2879 ( .A1(n2524), .A2(n2933), .ZN(n2559) );
  INV_X1 U2880 ( .A(n2934), .ZN(n2524) );
  NAND2_X1 U2881 ( .A1(n2526), .A2(n2527), .ZN(n2934) );
  NOR2_X1 U2882 ( .A1(n2933), .A2(n2935), .ZN(n2527) );
  NOR2_X1 U2883 ( .A1(n2936), .A2(n2937), .ZN(n2935) );
  INV_X1 U2884 ( .A(n2938), .ZN(n2933) );
  NAND2_X1 U2885 ( .A1(n2937), .A2(n2936), .ZN(n2938) );
  NAND2_X1 U2886 ( .A1(n2939), .A2(n2940), .ZN(n2936) );
  NAND2_X1 U2887 ( .A1(n2941), .A2(n2942), .ZN(n2940) );
  XNOR2_X1 U2888 ( .A(n2943), .B(n2944), .ZN(n2937) );
  XNOR2_X1 U2889 ( .A(n2945), .B(n2946), .ZN(n2944) );
  NOR2_X1 U2890 ( .A1(n2947), .A2(n2932), .ZN(n2526) );
  XOR2_X1 U2891 ( .A(n2948), .B(n2941), .Z(n2932) );
  XNOR2_X1 U2892 ( .A(n2949), .B(n2950), .ZN(n2941) );
  XOR2_X1 U2893 ( .A(n2951), .B(n2952), .Z(n2949) );
  NAND2_X1 U2894 ( .A1(n2939), .A2(n2942), .ZN(n2948) );
  NAND2_X1 U2895 ( .A1(n2953), .A2(n2954), .ZN(n2942) );
  NAND2_X1 U2896 ( .A1(a_0_), .A2(b_11_), .ZN(n2954) );
  INV_X1 U2897 ( .A(n2955), .ZN(n2953) );
  NAND2_X1 U2898 ( .A1(a_0_), .A2(n2955), .ZN(n2939) );
  NAND2_X1 U2899 ( .A1(n2956), .A2(n2957), .ZN(n2955) );
  NAND2_X1 U2900 ( .A1(n2958), .A2(n2959), .ZN(n2957) );
  INV_X1 U2901 ( .A(n2931), .ZN(n2947) );
  NAND2_X1 U2902 ( .A1(n2699), .A2(n2960), .ZN(n2931) );
  NAND2_X1 U2903 ( .A1(n2698), .A2(n2700), .ZN(n2960) );
  NAND2_X1 U2904 ( .A1(n2961), .A2(n2962), .ZN(n2700) );
  NAND2_X1 U2905 ( .A1(a_0_), .A2(b_12_), .ZN(n2962) );
  INV_X1 U2906 ( .A(n2963), .ZN(n2961) );
  XNOR2_X1 U2907 ( .A(n2964), .B(n2958), .ZN(n2698) );
  XNOR2_X1 U2908 ( .A(n2965), .B(n2966), .ZN(n2958) );
  NAND2_X1 U2909 ( .A1(n2967), .A2(n2968), .ZN(n2965) );
  NAND2_X1 U2910 ( .A1(n2956), .A2(n2959), .ZN(n2964) );
  NAND2_X1 U2911 ( .A1(n2969), .A2(n2970), .ZN(n2959) );
  NAND2_X1 U2912 ( .A1(b_11_), .A2(a_1_), .ZN(n2970) );
  INV_X1 U2913 ( .A(n2971), .ZN(n2969) );
  NAND2_X1 U2914 ( .A1(a_1_), .A2(n2971), .ZN(n2956) );
  NAND2_X1 U2915 ( .A1(n2972), .A2(n2973), .ZN(n2971) );
  NAND2_X1 U2916 ( .A1(n2974), .A2(a_2_), .ZN(n2973) );
  NOR2_X1 U2917 ( .A1(n2975), .A2(n2281), .ZN(n2974) );
  NOR2_X1 U2918 ( .A1(n2976), .A2(n2977), .ZN(n2975) );
  NAND2_X1 U2919 ( .A1(n2976), .A2(n2977), .ZN(n2972) );
  NAND2_X1 U2920 ( .A1(a_0_), .A2(n2963), .ZN(n2699) );
  NAND2_X1 U2921 ( .A1(n2978), .A2(n2979), .ZN(n2963) );
  NAND2_X1 U2922 ( .A1(n2980), .A2(b_12_), .ZN(n2979) );
  NOR2_X1 U2923 ( .A1(n2981), .A2(n2500), .ZN(n2980) );
  NOR2_X1 U2924 ( .A1(n2818), .A2(n2820), .ZN(n2981) );
  NAND2_X1 U2925 ( .A1(n2818), .A2(n2820), .ZN(n2978) );
  NAND2_X1 U2926 ( .A1(n2982), .A2(n2983), .ZN(n2820) );
  NAND2_X1 U2927 ( .A1(n2984), .A2(a_2_), .ZN(n2983) );
  NOR2_X1 U2928 ( .A1(n2985), .A2(n2489), .ZN(n2984) );
  NOR2_X1 U2929 ( .A1(n2828), .A2(n2830), .ZN(n2985) );
  NAND2_X1 U2930 ( .A1(n2828), .A2(n2830), .ZN(n2982) );
  NAND2_X1 U2931 ( .A1(n2986), .A2(n2987), .ZN(n2830) );
  NAND2_X1 U2932 ( .A1(n2988), .A2(a_3_), .ZN(n2987) );
  NOR2_X1 U2933 ( .A1(n2989), .A2(n2489), .ZN(n2988) );
  NOR2_X1 U2934 ( .A1(n2836), .A2(n2838), .ZN(n2989) );
  NAND2_X1 U2935 ( .A1(n2836), .A2(n2838), .ZN(n2986) );
  NAND2_X1 U2936 ( .A1(n2990), .A2(n2991), .ZN(n2838) );
  NAND2_X1 U2937 ( .A1(n2992), .A2(a_4_), .ZN(n2991) );
  NOR2_X1 U2938 ( .A1(n2993), .A2(n2489), .ZN(n2992) );
  NOR2_X1 U2939 ( .A1(n2845), .A2(n2847), .ZN(n2993) );
  NAND2_X1 U2940 ( .A1(n2845), .A2(n2847), .ZN(n2990) );
  NAND2_X1 U2941 ( .A1(n2994), .A2(n2995), .ZN(n2847) );
  NAND2_X1 U2942 ( .A1(n2996), .A2(a_5_), .ZN(n2995) );
  NOR2_X1 U2943 ( .A1(n2997), .A2(n2489), .ZN(n2996) );
  NOR2_X1 U2944 ( .A1(n2927), .A2(n2929), .ZN(n2997) );
  NAND2_X1 U2945 ( .A1(n2927), .A2(n2929), .ZN(n2994) );
  NAND2_X1 U2946 ( .A1(n2998), .A2(n2999), .ZN(n2929) );
  NAND2_X1 U2947 ( .A1(n3000), .A2(a_6_), .ZN(n2999) );
  NOR2_X1 U2948 ( .A1(n3001), .A2(n2489), .ZN(n3000) );
  NOR2_X1 U2949 ( .A1(n2858), .A2(n2859), .ZN(n3001) );
  NAND2_X1 U2950 ( .A1(n2858), .A2(n2859), .ZN(n2998) );
  NAND2_X1 U2951 ( .A1(n3002), .A2(n3003), .ZN(n2859) );
  NAND2_X1 U2952 ( .A1(n3004), .A2(a_7_), .ZN(n3003) );
  NOR2_X1 U2953 ( .A1(n3005), .A2(n2489), .ZN(n3004) );
  NOR2_X1 U2954 ( .A1(n2924), .A2(n2926), .ZN(n3005) );
  NAND2_X1 U2955 ( .A1(n2924), .A2(n2926), .ZN(n3002) );
  NAND2_X1 U2956 ( .A1(n3006), .A2(n3007), .ZN(n2926) );
  INV_X1 U2957 ( .A(n3008), .ZN(n3007) );
  NOR2_X1 U2958 ( .A1(n2872), .A2(n3009), .ZN(n3008) );
  NOR2_X1 U2959 ( .A1(n2871), .A2(n2869), .ZN(n3009) );
  NAND2_X1 U2960 ( .A1(a_8_), .A2(b_12_), .ZN(n2872) );
  NAND2_X1 U2961 ( .A1(n2869), .A2(n2871), .ZN(n3006) );
  NAND2_X1 U2962 ( .A1(n3010), .A2(n3011), .ZN(n2871) );
  NAND2_X1 U2963 ( .A1(n2880), .A2(n3012), .ZN(n3011) );
  NAND2_X1 U2964 ( .A1(n2877), .A2(n2879), .ZN(n3012) );
  NOR2_X1 U2965 ( .A1(n2311), .A2(n2489), .ZN(n2880) );
  INV_X1 U2966 ( .A(n3013), .ZN(n3010) );
  NOR2_X1 U2967 ( .A1(n2879), .A2(n2877), .ZN(n3013) );
  XOR2_X1 U2968 ( .A(n3014), .B(n3015), .Z(n2877) );
  XOR2_X1 U2969 ( .A(n3016), .B(n3017), .Z(n3014) );
  NAND2_X1 U2970 ( .A1(n3018), .A2(n3019), .ZN(n2879) );
  NAND2_X1 U2971 ( .A1(n2885), .A2(n3020), .ZN(n3019) );
  NAND2_X1 U2972 ( .A1(n2887), .A2(n2886), .ZN(n3020) );
  XNOR2_X1 U2973 ( .A(n3021), .B(n3022), .ZN(n2885) );
  XOR2_X1 U2974 ( .A(n2477), .B(n3023), .Z(n3022) );
  INV_X1 U2975 ( .A(n3024), .ZN(n3018) );
  NOR2_X1 U2976 ( .A1(n2886), .A2(n2887), .ZN(n3024) );
  NOR2_X1 U2977 ( .A1(n2492), .A2(n2489), .ZN(n2887) );
  NAND2_X1 U2978 ( .A1(n2894), .A2(n3025), .ZN(n2886) );
  NAND2_X1 U2979 ( .A1(n2893), .A2(n2895), .ZN(n3025) );
  NAND2_X1 U2980 ( .A1(n3026), .A2(n3027), .ZN(n2895) );
  NAND2_X1 U2981 ( .A1(a_11_), .A2(b_12_), .ZN(n3026) );
  XNOR2_X1 U2982 ( .A(n3028), .B(n3029), .ZN(n2893) );
  XOR2_X1 U2983 ( .A(n3030), .B(n3031), .Z(n3029) );
  NAND2_X1 U2984 ( .A1(b_11_), .A2(a_12_), .ZN(n3031) );
  NAND2_X1 U2985 ( .A1(n3032), .A2(a_11_), .ZN(n2894) );
  INV_X1 U2986 ( .A(n3027), .ZN(n3032) );
  NAND2_X1 U2987 ( .A1(n3033), .A2(n3034), .ZN(n3027) );
  NAND2_X1 U2988 ( .A1(n2921), .A2(n3035), .ZN(n3034) );
  INV_X1 U2989 ( .A(n3036), .ZN(n3035) );
  NOR2_X1 U2990 ( .A1(n2268), .A2(n2922), .ZN(n3036) );
  XNOR2_X1 U2991 ( .A(n3037), .B(n3038), .ZN(n2921) );
  XOR2_X1 U2992 ( .A(n3039), .B(n3040), .Z(n3038) );
  NAND2_X1 U2993 ( .A1(b_11_), .A2(a_13_), .ZN(n3037) );
  NAND2_X1 U2994 ( .A1(n2922), .A2(n2268), .ZN(n3033) );
  NAND2_X1 U2995 ( .A1(b_12_), .A2(a_12_), .ZN(n2268) );
  NOR2_X1 U2996 ( .A1(n3041), .A2(n3042), .ZN(n2922) );
  INV_X1 U2997 ( .A(n3043), .ZN(n3042) );
  NAND2_X1 U2998 ( .A1(n2905), .A2(n3044), .ZN(n3043) );
  NAND2_X1 U2999 ( .A1(n3045), .A2(n2907), .ZN(n3044) );
  NOR2_X1 U3000 ( .A1(n2489), .A2(n2252), .ZN(n2905) );
  NOR2_X1 U3001 ( .A1(n2907), .A2(n3045), .ZN(n3041) );
  INV_X1 U3002 ( .A(n2908), .ZN(n3045) );
  NAND2_X1 U3003 ( .A1(n3046), .A2(n3047), .ZN(n2908) );
  NAND2_X1 U3004 ( .A1(b_10_), .A2(n3048), .ZN(n3047) );
  NAND2_X1 U3005 ( .A1(n2227), .A2(n3049), .ZN(n3048) );
  NAND2_X1 U3006 ( .A1(a_15_), .A2(n2281), .ZN(n3049) );
  NAND2_X1 U3007 ( .A1(b_11_), .A2(n3050), .ZN(n3046) );
  NAND2_X1 U3008 ( .A1(n2231), .A2(n3051), .ZN(n3050) );
  NAND2_X1 U3009 ( .A1(a_14_), .A2(n2491), .ZN(n3051) );
  NAND2_X1 U3010 ( .A1(n3052), .A2(n2488), .ZN(n2907) );
  NOR2_X1 U3011 ( .A1(n2281), .A2(n2489), .ZN(n3052) );
  XNOR2_X1 U3012 ( .A(n3053), .B(n3054), .ZN(n2869) );
  NAND2_X1 U3013 ( .A1(n3055), .A2(n3056), .ZN(n3053) );
  XNOR2_X1 U3014 ( .A(n3057), .B(n3058), .ZN(n2924) );
  NAND2_X1 U3015 ( .A1(n3059), .A2(n3060), .ZN(n3057) );
  XNOR2_X1 U3016 ( .A(n3061), .B(n3062), .ZN(n2858) );
  NAND2_X1 U3017 ( .A1(n3063), .A2(n3064), .ZN(n3061) );
  XNOR2_X1 U3018 ( .A(n3065), .B(n3066), .ZN(n2927) );
  XOR2_X1 U3019 ( .A(n3067), .B(n3068), .Z(n3066) );
  NAND2_X1 U3020 ( .A1(a_6_), .A2(b_11_), .ZN(n3068) );
  XNOR2_X1 U3021 ( .A(n3069), .B(n3070), .ZN(n2845) );
  NAND2_X1 U3022 ( .A1(n3071), .A2(n3072), .ZN(n3069) );
  XOR2_X1 U3023 ( .A(n3073), .B(n3074), .Z(n2836) );
  XOR2_X1 U3024 ( .A(n3075), .B(n3076), .Z(n3073) );
  XOR2_X1 U3025 ( .A(n3077), .B(n3078), .Z(n2828) );
  XOR2_X1 U3026 ( .A(n3079), .B(n3080), .Z(n3077) );
  XNOR2_X1 U3027 ( .A(n2976), .B(n3081), .ZN(n2818) );
  XOR2_X1 U3028 ( .A(n2977), .B(n3082), .Z(n3081) );
  NAND2_X1 U3029 ( .A1(a_2_), .A2(b_11_), .ZN(n3082) );
  NAND2_X1 U3030 ( .A1(n3083), .A2(n3084), .ZN(n2977) );
  NAND2_X1 U3031 ( .A1(n3080), .A2(n3085), .ZN(n3084) );
  INV_X1 U3032 ( .A(n3086), .ZN(n3085) );
  NOR2_X1 U3033 ( .A1(n3079), .A2(n3078), .ZN(n3086) );
  NOR2_X1 U3034 ( .A1(n2410), .A2(n2281), .ZN(n3080) );
  NAND2_X1 U3035 ( .A1(n3078), .A2(n3079), .ZN(n3083) );
  NAND2_X1 U3036 ( .A1(n3087), .A2(n3088), .ZN(n3079) );
  NAND2_X1 U3037 ( .A1(n3076), .A2(n3089), .ZN(n3088) );
  INV_X1 U3038 ( .A(n3090), .ZN(n3089) );
  NOR2_X1 U3039 ( .A1(n3075), .A2(n3074), .ZN(n3090) );
  NOR2_X1 U3040 ( .A1(n2497), .A2(n2281), .ZN(n3076) );
  NAND2_X1 U3041 ( .A1(n3074), .A2(n3075), .ZN(n3087) );
  NAND2_X1 U3042 ( .A1(n3071), .A2(n3091), .ZN(n3075) );
  NAND2_X1 U3043 ( .A1(n3070), .A2(n3072), .ZN(n3091) );
  NAND2_X1 U3044 ( .A1(n3092), .A2(n3093), .ZN(n3072) );
  NAND2_X1 U3045 ( .A1(a_5_), .A2(b_11_), .ZN(n3093) );
  INV_X1 U3046 ( .A(n3094), .ZN(n3092) );
  XOR2_X1 U3047 ( .A(n3095), .B(n3096), .Z(n3070) );
  XOR2_X1 U3048 ( .A(n3097), .B(n3098), .Z(n3096) );
  NAND2_X1 U3049 ( .A1(a_5_), .A2(n3094), .ZN(n3071) );
  NAND2_X1 U3050 ( .A1(n3099), .A2(n3100), .ZN(n3094) );
  NAND2_X1 U3051 ( .A1(n3101), .A2(a_6_), .ZN(n3100) );
  NOR2_X1 U3052 ( .A1(n3102), .A2(n2281), .ZN(n3101) );
  NOR2_X1 U3053 ( .A1(n3065), .A2(n3067), .ZN(n3102) );
  NAND2_X1 U3054 ( .A1(n3065), .A2(n3067), .ZN(n3099) );
  NAND2_X1 U3055 ( .A1(n3063), .A2(n3103), .ZN(n3067) );
  NAND2_X1 U3056 ( .A1(n3062), .A2(n3064), .ZN(n3103) );
  NAND2_X1 U3057 ( .A1(n3104), .A2(n3105), .ZN(n3064) );
  NAND2_X1 U3058 ( .A1(a_7_), .A2(b_11_), .ZN(n3105) );
  INV_X1 U3059 ( .A(n3106), .ZN(n3104) );
  XNOR2_X1 U3060 ( .A(n3107), .B(n3108), .ZN(n3062) );
  XOR2_X1 U3061 ( .A(n3109), .B(n3110), .Z(n3108) );
  NAND2_X1 U3062 ( .A1(a_7_), .A2(n3106), .ZN(n3063) );
  NAND2_X1 U3063 ( .A1(n3059), .A2(n3111), .ZN(n3106) );
  NAND2_X1 U3064 ( .A1(n3058), .A2(n3060), .ZN(n3111) );
  NAND2_X1 U3065 ( .A1(n3112), .A2(n3113), .ZN(n3060) );
  NAND2_X1 U3066 ( .A1(a_8_), .A2(b_11_), .ZN(n3113) );
  INV_X1 U3067 ( .A(n3114), .ZN(n3112) );
  XNOR2_X1 U3068 ( .A(n3115), .B(n3116), .ZN(n3058) );
  XNOR2_X1 U3069 ( .A(n3117), .B(n3118), .ZN(n3116) );
  NAND2_X1 U3070 ( .A1(a_8_), .A2(n3114), .ZN(n3059) );
  NAND2_X1 U3071 ( .A1(n3055), .A2(n3119), .ZN(n3114) );
  NAND2_X1 U3072 ( .A1(n3054), .A2(n3056), .ZN(n3119) );
  NAND2_X1 U3073 ( .A1(n3120), .A2(n3121), .ZN(n3056) );
  NAND2_X1 U3074 ( .A1(a_9_), .A2(b_11_), .ZN(n3120) );
  XNOR2_X1 U3075 ( .A(n3122), .B(n3123), .ZN(n3054) );
  XOR2_X1 U3076 ( .A(n3124), .B(n2493), .Z(n3122) );
  INV_X1 U3077 ( .A(n3125), .ZN(n3055) );
  NOR2_X1 U3078 ( .A1(n3121), .A2(n2311), .ZN(n3125) );
  NAND2_X1 U3079 ( .A1(n3126), .A2(n3127), .ZN(n3121) );
  NAND2_X1 U3080 ( .A1(n3015), .A2(n3128), .ZN(n3127) );
  NAND2_X1 U3081 ( .A1(n3017), .A2(n3016), .ZN(n3128) );
  XOR2_X1 U3082 ( .A(n3129), .B(n3130), .Z(n3015) );
  NAND2_X1 U3083 ( .A1(n3131), .A2(n3132), .ZN(n3129) );
  INV_X1 U3084 ( .A(n3133), .ZN(n3126) );
  NOR2_X1 U3085 ( .A1(n3016), .A2(n3017), .ZN(n3133) );
  NOR2_X1 U3086 ( .A1(n2492), .A2(n2281), .ZN(n3017) );
  NAND2_X1 U3087 ( .A1(n3134), .A2(n3135), .ZN(n3016) );
  INV_X1 U3088 ( .A(n3136), .ZN(n3135) );
  NOR2_X1 U3089 ( .A1(n3021), .A2(n3137), .ZN(n3136) );
  NOR2_X1 U3090 ( .A1(n3023), .A2(n2275), .ZN(n3137) );
  XOR2_X1 U3091 ( .A(n3138), .B(n3139), .Z(n3021) );
  XOR2_X1 U3092 ( .A(n3140), .B(n3141), .Z(n3139) );
  NAND2_X1 U3093 ( .A1(b_10_), .A2(a_12_), .ZN(n3141) );
  NAND2_X1 U3094 ( .A1(n2275), .A2(n3023), .ZN(n3134) );
  NAND2_X1 U3095 ( .A1(n3142), .A2(n3143), .ZN(n3023) );
  NAND2_X1 U3096 ( .A1(n3144), .A2(b_11_), .ZN(n3143) );
  NOR2_X1 U3097 ( .A1(n3145), .A2(n2490), .ZN(n3144) );
  NOR2_X1 U3098 ( .A1(n3028), .A2(n3030), .ZN(n3145) );
  NAND2_X1 U3099 ( .A1(n3028), .A2(n3030), .ZN(n3142) );
  NAND2_X1 U3100 ( .A1(n3146), .A2(n3147), .ZN(n3030) );
  NAND2_X1 U3101 ( .A1(n3148), .A2(b_11_), .ZN(n3147) );
  NOR2_X1 U3102 ( .A1(n3149), .A2(n2252), .ZN(n3148) );
  NOR2_X1 U3103 ( .A1(n3150), .A2(n3040), .ZN(n3149) );
  NAND2_X1 U3104 ( .A1(n3150), .A2(n3040), .ZN(n3146) );
  NAND2_X1 U3105 ( .A1(n3151), .A2(n3152), .ZN(n3040) );
  NAND2_X1 U3106 ( .A1(b_10_), .A2(n3153), .ZN(n3152) );
  NAND2_X1 U3107 ( .A1(n2231), .A2(n3154), .ZN(n3153) );
  NAND2_X1 U3108 ( .A1(a_14_), .A2(n2312), .ZN(n3154) );
  NAND2_X1 U3109 ( .A1(b_9_), .A2(n3155), .ZN(n3151) );
  NAND2_X1 U3110 ( .A1(n2227), .A2(n3156), .ZN(n3155) );
  NAND2_X1 U3111 ( .A1(a_15_), .A2(n2491), .ZN(n3156) );
  INV_X1 U3112 ( .A(n3039), .ZN(n3150) );
  NAND2_X1 U3113 ( .A1(n3157), .A2(n2488), .ZN(n3039) );
  NOR2_X1 U3114 ( .A1(n2281), .A2(n2491), .ZN(n3157) );
  XOR2_X1 U3115 ( .A(n3158), .B(n3159), .Z(n3028) );
  XOR2_X1 U3116 ( .A(n3160), .B(n3161), .Z(n3159) );
  NAND2_X1 U3117 ( .A1(b_10_), .A2(a_13_), .ZN(n3158) );
  INV_X1 U3118 ( .A(n2477), .ZN(n2275) );
  NAND2_X1 U3119 ( .A1(a_11_), .A2(b_11_), .ZN(n2477) );
  XNOR2_X1 U3120 ( .A(n3162), .B(n3163), .ZN(n3065) );
  XNOR2_X1 U3121 ( .A(n3164), .B(n3165), .ZN(n3162) );
  XNOR2_X1 U3122 ( .A(n3166), .B(n3167), .ZN(n3074) );
  NAND2_X1 U3123 ( .A1(n3168), .A2(n3169), .ZN(n3166) );
  XOR2_X1 U3124 ( .A(n3170), .B(n3171), .Z(n3078) );
  XOR2_X1 U3125 ( .A(n3172), .B(n3173), .Z(n3170) );
  NOR2_X1 U3126 ( .A1(n2491), .A2(n2497), .ZN(n3173) );
  XOR2_X1 U3127 ( .A(n3174), .B(n3175), .Z(n2976) );
  XNOR2_X1 U3128 ( .A(n3176), .B(n3177), .ZN(n3175) );
  NOR2_X1 U3129 ( .A1(n3178), .A2(n2181), .ZN(n2554) );
  INV_X1 U3130 ( .A(n3179), .ZN(n2181) );
  NAND2_X1 U3131 ( .A1(n2183), .A2(n2184), .ZN(n3179) );
  NOR2_X1 U3132 ( .A1(n3180), .A2(n3178), .ZN(n2184) );
  NOR2_X1 U3133 ( .A1(n3181), .A2(n3182), .ZN(n3180) );
  NOR2_X1 U3134 ( .A1(n2557), .A2(n2558), .ZN(n2183) );
  XOR2_X1 U3135 ( .A(n3183), .B(n3184), .Z(n2558) );
  XOR2_X1 U3136 ( .A(n3185), .B(n3186), .Z(n3184) );
  NAND2_X1 U3137 ( .A1(a_0_), .A2(b_9_), .ZN(n3186) );
  NOR2_X1 U3138 ( .A1(n3187), .A2(n3188), .ZN(n2557) );
  INV_X1 U3139 ( .A(n3189), .ZN(n3188) );
  NAND2_X1 U3140 ( .A1(n2946), .A2(n3190), .ZN(n3189) );
  NAND2_X1 U3141 ( .A1(n2943), .A2(n2945), .ZN(n3190) );
  NOR2_X1 U3142 ( .A1(n3191), .A2(n2491), .ZN(n2946) );
  NOR2_X1 U3143 ( .A1(n2945), .A2(n2943), .ZN(n3187) );
  XOR2_X1 U3144 ( .A(n3192), .B(n3193), .Z(n2943) );
  XOR2_X1 U3145 ( .A(n3194), .B(n3195), .Z(n3193) );
  NAND2_X1 U3146 ( .A1(b_9_), .A2(a_1_), .ZN(n3195) );
  NAND2_X1 U3147 ( .A1(n3196), .A2(n3197), .ZN(n2945) );
  NAND2_X1 U3148 ( .A1(n2950), .A2(n3198), .ZN(n3197) );
  NAND2_X1 U3149 ( .A1(n2952), .A2(n2951), .ZN(n3198) );
  XOR2_X1 U3150 ( .A(n3199), .B(n3200), .Z(n2950) );
  XOR2_X1 U3151 ( .A(n3201), .B(n3202), .Z(n3200) );
  NAND2_X1 U3152 ( .A1(a_2_), .A2(b_9_), .ZN(n3202) );
  INV_X1 U3153 ( .A(n3203), .ZN(n3196) );
  NOR2_X1 U3154 ( .A1(n2951), .A2(n2952), .ZN(n3203) );
  NOR2_X1 U3155 ( .A1(n2491), .A2(n2500), .ZN(n2952) );
  NAND2_X1 U3156 ( .A1(n2967), .A2(n3204), .ZN(n2951) );
  NAND2_X1 U3157 ( .A1(n2966), .A2(n2968), .ZN(n3204) );
  NAND2_X1 U3158 ( .A1(n3205), .A2(n3206), .ZN(n2968) );
  NAND2_X1 U3159 ( .A1(a_2_), .A2(b_10_), .ZN(n3205) );
  XOR2_X1 U3160 ( .A(n3207), .B(n3208), .Z(n2966) );
  XNOR2_X1 U3161 ( .A(n3209), .B(n3210), .ZN(n3208) );
  NAND2_X1 U3162 ( .A1(a_3_), .A2(b_9_), .ZN(n3210) );
  INV_X1 U3163 ( .A(n3211), .ZN(n2967) );
  NOR2_X1 U3164 ( .A1(n3206), .A2(n2426), .ZN(n3211) );
  NAND2_X1 U3165 ( .A1(n3212), .A2(n3213), .ZN(n3206) );
  NAND2_X1 U3166 ( .A1(n3174), .A2(n3214), .ZN(n3213) );
  NAND2_X1 U3167 ( .A1(n3177), .A2(n3176), .ZN(n3214) );
  XOR2_X1 U3168 ( .A(n3215), .B(n3216), .Z(n3174) );
  XOR2_X1 U3169 ( .A(n3217), .B(n3218), .Z(n3215) );
  INV_X1 U3170 ( .A(n3219), .ZN(n3212) );
  NOR2_X1 U3171 ( .A1(n3176), .A2(n3177), .ZN(n3219) );
  NOR2_X1 U3172 ( .A1(n2410), .A2(n2491), .ZN(n3177) );
  NAND2_X1 U3173 ( .A1(n3220), .A2(n3221), .ZN(n3176) );
  NAND2_X1 U3174 ( .A1(n3222), .A2(a_4_), .ZN(n3221) );
  NOR2_X1 U3175 ( .A1(n3223), .A2(n2491), .ZN(n3222) );
  NOR2_X1 U3176 ( .A1(n3171), .A2(n3172), .ZN(n3223) );
  NAND2_X1 U3177 ( .A1(n3171), .A2(n3172), .ZN(n3220) );
  NAND2_X1 U3178 ( .A1(n3168), .A2(n3224), .ZN(n3172) );
  NAND2_X1 U3179 ( .A1(n3167), .A2(n3169), .ZN(n3224) );
  NAND2_X1 U3180 ( .A1(n3225), .A2(n3226), .ZN(n3169) );
  NAND2_X1 U3181 ( .A1(a_5_), .A2(b_10_), .ZN(n3226) );
  XOR2_X1 U3182 ( .A(n3227), .B(n3228), .Z(n3167) );
  XOR2_X1 U3183 ( .A(n3229), .B(n3230), .Z(n3227) );
  NAND2_X1 U3184 ( .A1(a_5_), .A2(n3231), .ZN(n3168) );
  INV_X1 U3185 ( .A(n3225), .ZN(n3231) );
  NOR2_X1 U3186 ( .A1(n3232), .A2(n3233), .ZN(n3225) );
  INV_X1 U3187 ( .A(n3234), .ZN(n3233) );
  NAND2_X1 U3188 ( .A1(n3098), .A2(n3235), .ZN(n3234) );
  NAND2_X1 U3189 ( .A1(n3097), .A2(n3095), .ZN(n3235) );
  NOR2_X1 U3190 ( .A1(n2495), .A2(n2491), .ZN(n3098) );
  NOR2_X1 U3191 ( .A1(n3095), .A2(n3097), .ZN(n3232) );
  NOR2_X1 U3192 ( .A1(n3236), .A2(n3237), .ZN(n3097) );
  INV_X1 U3193 ( .A(n3238), .ZN(n3237) );
  NAND2_X1 U3194 ( .A1(n3164), .A2(n3239), .ZN(n3238) );
  NAND2_X1 U3195 ( .A1(n3165), .A2(n3163), .ZN(n3239) );
  NOR2_X1 U3196 ( .A1(n2342), .A2(n2491), .ZN(n3164) );
  NOR2_X1 U3197 ( .A1(n3163), .A2(n3165), .ZN(n3236) );
  NOR2_X1 U3198 ( .A1(n3240), .A2(n3241), .ZN(n3165) );
  NOR2_X1 U3199 ( .A1(n3110), .A2(n3242), .ZN(n3241) );
  NOR2_X1 U3200 ( .A1(n3109), .A2(n3107), .ZN(n3242) );
  NAND2_X1 U3201 ( .A1(a_8_), .A2(b_10_), .ZN(n3110) );
  INV_X1 U3202 ( .A(n3243), .ZN(n3240) );
  NAND2_X1 U3203 ( .A1(n3107), .A2(n3109), .ZN(n3243) );
  NAND2_X1 U3204 ( .A1(n3244), .A2(n3245), .ZN(n3109) );
  NAND2_X1 U3205 ( .A1(n3118), .A2(n3246), .ZN(n3245) );
  NAND2_X1 U3206 ( .A1(n3115), .A2(n3117), .ZN(n3246) );
  NOR2_X1 U3207 ( .A1(n2311), .A2(n2491), .ZN(n3118) );
  INV_X1 U3208 ( .A(n3247), .ZN(n3244) );
  NOR2_X1 U3209 ( .A1(n3117), .A2(n3115), .ZN(n3247) );
  XOR2_X1 U3210 ( .A(n3248), .B(n3249), .Z(n3115) );
  XOR2_X1 U3211 ( .A(n3250), .B(n3251), .Z(n3248) );
  NAND2_X1 U3212 ( .A1(n3252), .A2(n3253), .ZN(n3117) );
  NAND2_X1 U3213 ( .A1(n3123), .A2(n3254), .ZN(n3253) );
  NAND2_X1 U3214 ( .A1(n2493), .A2(n3124), .ZN(n3254) );
  XOR2_X1 U3215 ( .A(n3255), .B(n3256), .Z(n3123) );
  NAND2_X1 U3216 ( .A1(n3257), .A2(n3258), .ZN(n3255) );
  INV_X1 U3217 ( .A(n3259), .ZN(n3252) );
  NOR2_X1 U3218 ( .A1(n3124), .A2(n2493), .ZN(n3259) );
  NOR2_X1 U3219 ( .A1(n2491), .A2(n2492), .ZN(n2493) );
  NAND2_X1 U3220 ( .A1(n3131), .A2(n3260), .ZN(n3124) );
  NAND2_X1 U3221 ( .A1(n3130), .A2(n3132), .ZN(n3260) );
  NAND2_X1 U3222 ( .A1(n3261), .A2(n3262), .ZN(n3132) );
  NAND2_X1 U3223 ( .A1(b_10_), .A2(a_11_), .ZN(n3262) );
  INV_X1 U3224 ( .A(n3263), .ZN(n3261) );
  XNOR2_X1 U3225 ( .A(n3264), .B(n3265), .ZN(n3130) );
  XOR2_X1 U3226 ( .A(n3266), .B(n3267), .Z(n3265) );
  NAND2_X1 U3227 ( .A1(b_9_), .A2(a_12_), .ZN(n3267) );
  NAND2_X1 U3228 ( .A1(a_11_), .A2(n3263), .ZN(n3131) );
  NAND2_X1 U3229 ( .A1(n3268), .A2(n3269), .ZN(n3263) );
  NAND2_X1 U3230 ( .A1(n3270), .A2(b_10_), .ZN(n3269) );
  NOR2_X1 U3231 ( .A1(n3271), .A2(n2490), .ZN(n3270) );
  NOR2_X1 U3232 ( .A1(n3138), .A2(n3140), .ZN(n3271) );
  NAND2_X1 U3233 ( .A1(n3138), .A2(n3140), .ZN(n3268) );
  NAND2_X1 U3234 ( .A1(n3272), .A2(n3273), .ZN(n3140) );
  NAND2_X1 U3235 ( .A1(n3274), .A2(b_10_), .ZN(n3273) );
  NOR2_X1 U3236 ( .A1(n3275), .A2(n2252), .ZN(n3274) );
  NOR2_X1 U3237 ( .A1(n3276), .A2(n3161), .ZN(n3275) );
  NAND2_X1 U3238 ( .A1(n3276), .A2(n3161), .ZN(n3272) );
  NAND2_X1 U3239 ( .A1(n3277), .A2(n3278), .ZN(n3161) );
  NAND2_X1 U3240 ( .A1(b_8_), .A2(n3279), .ZN(n3278) );
  NAND2_X1 U3241 ( .A1(n2227), .A2(n3280), .ZN(n3279) );
  NAND2_X1 U3242 ( .A1(a_15_), .A2(n2312), .ZN(n3280) );
  NAND2_X1 U3243 ( .A1(b_9_), .A2(n3281), .ZN(n3277) );
  NAND2_X1 U3244 ( .A1(n2231), .A2(n3282), .ZN(n3281) );
  NAND2_X1 U3245 ( .A1(a_14_), .A2(n3283), .ZN(n3282) );
  INV_X1 U3246 ( .A(n3160), .ZN(n3276) );
  NAND2_X1 U3247 ( .A1(n3284), .A2(n2488), .ZN(n3160) );
  NOR2_X1 U3248 ( .A1(n2491), .A2(n2312), .ZN(n3284) );
  XOR2_X1 U3249 ( .A(n3285), .B(n3286), .Z(n3138) );
  XOR2_X1 U3250 ( .A(n3287), .B(n3288), .Z(n3286) );
  NAND2_X1 U3251 ( .A1(b_9_), .A2(a_13_), .ZN(n3285) );
  XNOR2_X1 U3252 ( .A(n3289), .B(n3290), .ZN(n3107) );
  XOR2_X1 U3253 ( .A(n3291), .B(n2473), .Z(n3290) );
  XNOR2_X1 U3254 ( .A(n3292), .B(n3293), .ZN(n3163) );
  XOR2_X1 U3255 ( .A(n3294), .B(n3295), .Z(n3292) );
  XOR2_X1 U3256 ( .A(n3296), .B(n3297), .Z(n3095) );
  XNOR2_X1 U3257 ( .A(n3298), .B(n3299), .ZN(n3296) );
  XNOR2_X1 U3258 ( .A(n3300), .B(n3301), .ZN(n3171) );
  NAND2_X1 U3259 ( .A1(n3302), .A2(n3303), .ZN(n3300) );
  INV_X1 U3260 ( .A(n3304), .ZN(n3178) );
  NAND2_X1 U3261 ( .A1(n3181), .A2(n3182), .ZN(n3304) );
  NAND2_X1 U3262 ( .A1(n3305), .A2(n3306), .ZN(n3182) );
  NAND2_X1 U3263 ( .A1(n3307), .A2(a_0_), .ZN(n3306) );
  NOR2_X1 U3264 ( .A1(n3308), .A2(n2312), .ZN(n3307) );
  NOR2_X1 U3265 ( .A1(n3183), .A2(n3185), .ZN(n3308) );
  NAND2_X1 U3266 ( .A1(n3183), .A2(n3185), .ZN(n3305) );
  NAND2_X1 U3267 ( .A1(n3309), .A2(n3310), .ZN(n3185) );
  NAND2_X1 U3268 ( .A1(n3311), .A2(b_9_), .ZN(n3310) );
  NOR2_X1 U3269 ( .A1(n3312), .A2(n2500), .ZN(n3311) );
  NOR2_X1 U3270 ( .A1(n3194), .A2(n3192), .ZN(n3312) );
  NAND2_X1 U3271 ( .A1(n3192), .A2(n3194), .ZN(n3309) );
  NAND2_X1 U3272 ( .A1(n3313), .A2(n3314), .ZN(n3194) );
  NAND2_X1 U3273 ( .A1(n3315), .A2(a_2_), .ZN(n3314) );
  NOR2_X1 U3274 ( .A1(n3316), .A2(n2312), .ZN(n3315) );
  NOR2_X1 U3275 ( .A1(n3199), .A2(n3201), .ZN(n3316) );
  NAND2_X1 U3276 ( .A1(n3199), .A2(n3201), .ZN(n3313) );
  NAND2_X1 U3277 ( .A1(n3317), .A2(n3318), .ZN(n3201) );
  NAND2_X1 U3278 ( .A1(n3319), .A2(a_3_), .ZN(n3318) );
  NOR2_X1 U3279 ( .A1(n3320), .A2(n2312), .ZN(n3319) );
  NOR2_X1 U3280 ( .A1(n3209), .A2(n3207), .ZN(n3320) );
  NAND2_X1 U3281 ( .A1(n3207), .A2(n3209), .ZN(n3317) );
  NOR2_X1 U3282 ( .A1(n3321), .A2(n3322), .ZN(n3209) );
  INV_X1 U3283 ( .A(n3323), .ZN(n3322) );
  NAND2_X1 U3284 ( .A1(n3216), .A2(n3324), .ZN(n3323) );
  NAND2_X1 U3285 ( .A1(n3218), .A2(n3217), .ZN(n3324) );
  XOR2_X1 U3286 ( .A(n3325), .B(n3326), .Z(n3216) );
  XOR2_X1 U3287 ( .A(n3327), .B(n3328), .Z(n3326) );
  NAND2_X1 U3288 ( .A1(a_5_), .A2(b_8_), .ZN(n3328) );
  NOR2_X1 U3289 ( .A1(n3217), .A2(n3218), .ZN(n3321) );
  NOR2_X1 U3290 ( .A1(n2497), .A2(n2312), .ZN(n3218) );
  NAND2_X1 U3291 ( .A1(n3302), .A2(n3329), .ZN(n3217) );
  NAND2_X1 U3292 ( .A1(n3301), .A2(n3303), .ZN(n3329) );
  NAND2_X1 U3293 ( .A1(n3330), .A2(n3331), .ZN(n3303) );
  NAND2_X1 U3294 ( .A1(a_5_), .A2(b_9_), .ZN(n3331) );
  INV_X1 U3295 ( .A(n3332), .ZN(n3330) );
  XOR2_X1 U3296 ( .A(n3333), .B(n3334), .Z(n3301) );
  XOR2_X1 U3297 ( .A(n3335), .B(n3336), .Z(n3333) );
  NOR2_X1 U3298 ( .A1(n3283), .A2(n2495), .ZN(n3336) );
  NAND2_X1 U3299 ( .A1(a_5_), .A2(n3332), .ZN(n3302) );
  NAND2_X1 U3300 ( .A1(n3337), .A2(n3338), .ZN(n3332) );
  NAND2_X1 U3301 ( .A1(n3230), .A2(n3339), .ZN(n3338) );
  INV_X1 U3302 ( .A(n3340), .ZN(n3339) );
  NOR2_X1 U3303 ( .A1(n3228), .A2(n3229), .ZN(n3340) );
  NOR2_X1 U3304 ( .A1(n2495), .A2(n2312), .ZN(n3230) );
  NAND2_X1 U3305 ( .A1(n3228), .A2(n3229), .ZN(n3337) );
  NAND2_X1 U3306 ( .A1(n3341), .A2(n3342), .ZN(n3229) );
  NAND2_X1 U3307 ( .A1(n3299), .A2(n3343), .ZN(n3342) );
  NAND2_X1 U3308 ( .A1(n3297), .A2(n3298), .ZN(n3343) );
  NOR2_X1 U3309 ( .A1(n2342), .A2(n2312), .ZN(n3299) );
  INV_X1 U3310 ( .A(n3344), .ZN(n3341) );
  NOR2_X1 U3311 ( .A1(n3297), .A2(n3298), .ZN(n3344) );
  NOR2_X1 U3312 ( .A1(n3345), .A2(n3346), .ZN(n3298) );
  INV_X1 U3313 ( .A(n3347), .ZN(n3346) );
  NAND2_X1 U3314 ( .A1(n3295), .A2(n3348), .ZN(n3347) );
  NAND2_X1 U3315 ( .A1(n3293), .A2(n3294), .ZN(n3348) );
  NOR2_X1 U3316 ( .A1(n3349), .A2(n2312), .ZN(n3295) );
  NOR2_X1 U3317 ( .A1(n3293), .A2(n3294), .ZN(n3345) );
  NAND2_X1 U3318 ( .A1(n3350), .A2(n3351), .ZN(n3294) );
  NAND2_X1 U3319 ( .A1(n3289), .A2(n3352), .ZN(n3351) );
  NAND2_X1 U3320 ( .A1(n2306), .A2(n3353), .ZN(n3352) );
  INV_X1 U3321 ( .A(n3291), .ZN(n3353) );
  INV_X1 U3322 ( .A(n2473), .ZN(n2306) );
  XOR2_X1 U3323 ( .A(n3354), .B(n3355), .Z(n3289) );
  XOR2_X1 U3324 ( .A(n3356), .B(n3357), .Z(n3354) );
  NAND2_X1 U3325 ( .A1(n2473), .A2(n3291), .ZN(n3350) );
  NAND2_X1 U3326 ( .A1(n3358), .A2(n3359), .ZN(n3291) );
  NAND2_X1 U3327 ( .A1(n3249), .A2(n3360), .ZN(n3359) );
  NAND2_X1 U3328 ( .A1(n3251), .A2(n3250), .ZN(n3360) );
  XOR2_X1 U3329 ( .A(n3361), .B(n3362), .Z(n3249) );
  NAND2_X1 U3330 ( .A1(n3363), .A2(n3364), .ZN(n3361) );
  INV_X1 U3331 ( .A(n3365), .ZN(n3358) );
  NOR2_X1 U3332 ( .A1(n3250), .A2(n3251), .ZN(n3365) );
  NOR2_X1 U3333 ( .A1(n2312), .A2(n2492), .ZN(n3251) );
  NAND2_X1 U3334 ( .A1(n3257), .A2(n3366), .ZN(n3250) );
  NAND2_X1 U3335 ( .A1(n3256), .A2(n3258), .ZN(n3366) );
  NAND2_X1 U3336 ( .A1(n3367), .A2(n3368), .ZN(n3258) );
  NAND2_X1 U3337 ( .A1(b_9_), .A2(a_11_), .ZN(n3368) );
  INV_X1 U3338 ( .A(n3369), .ZN(n3367) );
  XNOR2_X1 U3339 ( .A(n3370), .B(n3371), .ZN(n3256) );
  XOR2_X1 U3340 ( .A(n3372), .B(n3373), .Z(n3371) );
  NAND2_X1 U3341 ( .A1(b_8_), .A2(a_12_), .ZN(n3373) );
  NAND2_X1 U3342 ( .A1(a_11_), .A2(n3369), .ZN(n3257) );
  NAND2_X1 U3343 ( .A1(n3374), .A2(n3375), .ZN(n3369) );
  NAND2_X1 U3344 ( .A1(n3376), .A2(b_9_), .ZN(n3375) );
  NOR2_X1 U3345 ( .A1(n3377), .A2(n2490), .ZN(n3376) );
  NOR2_X1 U3346 ( .A1(n3264), .A2(n3266), .ZN(n3377) );
  NAND2_X1 U3347 ( .A1(n3264), .A2(n3266), .ZN(n3374) );
  NAND2_X1 U3348 ( .A1(n3378), .A2(n3379), .ZN(n3266) );
  NAND2_X1 U3349 ( .A1(n3380), .A2(b_9_), .ZN(n3379) );
  NOR2_X1 U3350 ( .A1(n3381), .A2(n2252), .ZN(n3380) );
  NOR2_X1 U3351 ( .A1(n3382), .A2(n3288), .ZN(n3381) );
  NAND2_X1 U3352 ( .A1(n3382), .A2(n3288), .ZN(n3378) );
  NAND2_X1 U3353 ( .A1(n3383), .A2(n3384), .ZN(n3288) );
  NAND2_X1 U3354 ( .A1(b_7_), .A2(n3385), .ZN(n3384) );
  NAND2_X1 U3355 ( .A1(n2227), .A2(n3386), .ZN(n3385) );
  NAND2_X1 U3356 ( .A1(a_15_), .A2(n3283), .ZN(n3386) );
  NAND2_X1 U3357 ( .A1(b_8_), .A2(n3387), .ZN(n3383) );
  NAND2_X1 U3358 ( .A1(n2231), .A2(n3388), .ZN(n3387) );
  NAND2_X1 U3359 ( .A1(a_14_), .A2(n2343), .ZN(n3388) );
  INV_X1 U3360 ( .A(n3287), .ZN(n3382) );
  NAND2_X1 U3361 ( .A1(n3389), .A2(n2488), .ZN(n3287) );
  NOR2_X1 U3362 ( .A1(n2312), .A2(n3283), .ZN(n3389) );
  INV_X1 U3363 ( .A(b_9_), .ZN(n2312) );
  XOR2_X1 U3364 ( .A(n3390), .B(n3391), .Z(n3264) );
  XOR2_X1 U3365 ( .A(n3392), .B(n3393), .Z(n3391) );
  NAND2_X1 U3366 ( .A1(b_8_), .A2(a_13_), .ZN(n3390) );
  NAND2_X1 U3367 ( .A1(a_9_), .A2(b_9_), .ZN(n2473) );
  XNOR2_X1 U3368 ( .A(n3394), .B(n3395), .ZN(n3293) );
  XOR2_X1 U3369 ( .A(n3396), .B(n3397), .Z(n3395) );
  XNOR2_X1 U3370 ( .A(n3398), .B(n3399), .ZN(n3297) );
  XNOR2_X1 U3371 ( .A(n3400), .B(n2331), .ZN(n3399) );
  XNOR2_X1 U3372 ( .A(n3401), .B(n3402), .ZN(n3228) );
  XNOR2_X1 U3373 ( .A(n3403), .B(n3404), .ZN(n3402) );
  XNOR2_X1 U3374 ( .A(n3405), .B(n3406), .ZN(n3207) );
  NAND2_X1 U3375 ( .A1(n3407), .A2(n3408), .ZN(n3405) );
  XOR2_X1 U3376 ( .A(n3409), .B(n3410), .Z(n3199) );
  XOR2_X1 U3377 ( .A(n3411), .B(n3412), .Z(n3409) );
  NOR2_X1 U3378 ( .A1(n3283), .A2(n2410), .ZN(n3412) );
  XNOR2_X1 U3379 ( .A(n3413), .B(n3414), .ZN(n3192) );
  NAND2_X1 U3380 ( .A1(n3415), .A2(n3416), .ZN(n3413) );
  XNOR2_X1 U3381 ( .A(n3417), .B(n3418), .ZN(n3183) );
  NAND2_X1 U3382 ( .A1(n3419), .A2(n3420), .ZN(n3417) );
  XNOR2_X1 U3383 ( .A(n3421), .B(n3422), .ZN(n3181) );
  XNOR2_X1 U3384 ( .A(n3423), .B(n3424), .ZN(n3421) );
  NOR2_X1 U3385 ( .A1(n3425), .A2(n2191), .ZN(n2549) );
  INV_X1 U3386 ( .A(n3426), .ZN(n2191) );
  NAND2_X1 U3387 ( .A1(n2193), .A2(n2194), .ZN(n3426) );
  NOR2_X1 U3388 ( .A1(n3427), .A2(n3425), .ZN(n2194) );
  NOR2_X1 U3389 ( .A1(n3428), .A2(n3429), .ZN(n3427) );
  NOR2_X1 U3390 ( .A1(n3430), .A2(n2553), .ZN(n2193) );
  XOR2_X1 U3391 ( .A(n3431), .B(n3432), .Z(n2553) );
  NAND2_X1 U3392 ( .A1(n3433), .A2(n3434), .ZN(n3431) );
  INV_X1 U3393 ( .A(n2552), .ZN(n3430) );
  NAND2_X1 U3394 ( .A1(n3435), .A2(n3436), .ZN(n2552) );
  NAND2_X1 U3395 ( .A1(n3424), .A2(n3437), .ZN(n3436) );
  INV_X1 U3396 ( .A(n3438), .ZN(n3437) );
  NOR2_X1 U3397 ( .A1(n3423), .A2(n3422), .ZN(n3438) );
  NOR2_X1 U3398 ( .A1(n3191), .A2(n3283), .ZN(n3424) );
  NAND2_X1 U3399 ( .A1(n3422), .A2(n3423), .ZN(n3435) );
  NAND2_X1 U3400 ( .A1(n3419), .A2(n3439), .ZN(n3423) );
  NAND2_X1 U3401 ( .A1(n3418), .A2(n3420), .ZN(n3439) );
  NAND2_X1 U3402 ( .A1(n3440), .A2(n3441), .ZN(n3420) );
  NAND2_X1 U3403 ( .A1(b_8_), .A2(a_1_), .ZN(n3441) );
  INV_X1 U3404 ( .A(n3442), .ZN(n3440) );
  XNOR2_X1 U3405 ( .A(n3443), .B(n3444), .ZN(n3418) );
  XOR2_X1 U3406 ( .A(n3445), .B(n3446), .Z(n3444) );
  NAND2_X1 U3407 ( .A1(a_2_), .A2(b_7_), .ZN(n3446) );
  NAND2_X1 U3408 ( .A1(a_1_), .A2(n3442), .ZN(n3419) );
  NAND2_X1 U3409 ( .A1(n3415), .A2(n3447), .ZN(n3442) );
  NAND2_X1 U3410 ( .A1(n3414), .A2(n3416), .ZN(n3447) );
  NAND2_X1 U3411 ( .A1(n3448), .A2(n3449), .ZN(n3416) );
  NAND2_X1 U3412 ( .A1(a_2_), .A2(b_8_), .ZN(n3449) );
  INV_X1 U3413 ( .A(n3450), .ZN(n3448) );
  XNOR2_X1 U3414 ( .A(n3451), .B(n3452), .ZN(n3414) );
  XOR2_X1 U3415 ( .A(n3453), .B(n3454), .Z(n3452) );
  NAND2_X1 U3416 ( .A1(a_3_), .A2(b_7_), .ZN(n3454) );
  NAND2_X1 U3417 ( .A1(a_2_), .A2(n3450), .ZN(n3415) );
  NAND2_X1 U3418 ( .A1(n3455), .A2(n3456), .ZN(n3450) );
  NAND2_X1 U3419 ( .A1(n3457), .A2(a_3_), .ZN(n3456) );
  NOR2_X1 U3420 ( .A1(n3458), .A2(n3283), .ZN(n3457) );
  NOR2_X1 U3421 ( .A1(n3411), .A2(n3410), .ZN(n3458) );
  NAND2_X1 U3422 ( .A1(n3410), .A2(n3411), .ZN(n3455) );
  NAND2_X1 U3423 ( .A1(n3407), .A2(n3459), .ZN(n3411) );
  NAND2_X1 U3424 ( .A1(n3406), .A2(n3408), .ZN(n3459) );
  NAND2_X1 U3425 ( .A1(n3460), .A2(n3461), .ZN(n3408) );
  NAND2_X1 U3426 ( .A1(a_4_), .A2(b_8_), .ZN(n3461) );
  INV_X1 U3427 ( .A(n3462), .ZN(n3460) );
  XNOR2_X1 U3428 ( .A(n3463), .B(n3464), .ZN(n3406) );
  NAND2_X1 U3429 ( .A1(n3465), .A2(n3466), .ZN(n3463) );
  NAND2_X1 U3430 ( .A1(a_4_), .A2(n3462), .ZN(n3407) );
  NAND2_X1 U3431 ( .A1(n3467), .A2(n3468), .ZN(n3462) );
  NAND2_X1 U3432 ( .A1(n3469), .A2(a_5_), .ZN(n3468) );
  NOR2_X1 U3433 ( .A1(n3470), .A2(n3283), .ZN(n3469) );
  NOR2_X1 U3434 ( .A1(n3327), .A2(n3325), .ZN(n3470) );
  NAND2_X1 U3435 ( .A1(n3325), .A2(n3327), .ZN(n3467) );
  NAND2_X1 U3436 ( .A1(n3471), .A2(n3472), .ZN(n3327) );
  NAND2_X1 U3437 ( .A1(n3473), .A2(a_6_), .ZN(n3472) );
  NOR2_X1 U3438 ( .A1(n3474), .A2(n3283), .ZN(n3473) );
  NOR2_X1 U3439 ( .A1(n3335), .A2(n3334), .ZN(n3474) );
  NAND2_X1 U3440 ( .A1(n3334), .A2(n3335), .ZN(n3471) );
  NAND2_X1 U3441 ( .A1(n3475), .A2(n3476), .ZN(n3335) );
  NAND2_X1 U3442 ( .A1(n3404), .A2(n3477), .ZN(n3476) );
  NAND2_X1 U3443 ( .A1(n3401), .A2(n3403), .ZN(n3477) );
  NOR2_X1 U3444 ( .A1(n2342), .A2(n3283), .ZN(n3404) );
  INV_X1 U3445 ( .A(n3478), .ZN(n3475) );
  NOR2_X1 U3446 ( .A1(n3403), .A2(n3401), .ZN(n3478) );
  XNOR2_X1 U3447 ( .A(n3479), .B(n3480), .ZN(n3401) );
  XOR2_X1 U3448 ( .A(n3481), .B(n3482), .Z(n3480) );
  NAND2_X1 U3449 ( .A1(n3483), .A2(n3484), .ZN(n3403) );
  NAND2_X1 U3450 ( .A1(n3398), .A2(n3485), .ZN(n3484) );
  NAND2_X1 U3451 ( .A1(n2331), .A2(n3400), .ZN(n3485) );
  XOR2_X1 U3452 ( .A(n3486), .B(n3487), .Z(n3398) );
  XNOR2_X1 U3453 ( .A(n3488), .B(n3489), .ZN(n3487) );
  INV_X1 U3454 ( .A(n3490), .ZN(n3483) );
  NOR2_X1 U3455 ( .A1(n3400), .A2(n2331), .ZN(n3490) );
  NOR2_X1 U3456 ( .A1(n3283), .A2(n3349), .ZN(n2331) );
  NAND2_X1 U3457 ( .A1(n3491), .A2(n3492), .ZN(n3400) );
  NAND2_X1 U3458 ( .A1(n3397), .A2(n3493), .ZN(n3492) );
  INV_X1 U3459 ( .A(n3494), .ZN(n3493) );
  NOR2_X1 U3460 ( .A1(n3394), .A2(n3396), .ZN(n3494) );
  NOR2_X1 U3461 ( .A1(n3283), .A2(n2311), .ZN(n3397) );
  NAND2_X1 U3462 ( .A1(n3394), .A2(n3396), .ZN(n3491) );
  NOR2_X1 U3463 ( .A1(n3495), .A2(n3496), .ZN(n3396) );
  INV_X1 U3464 ( .A(n3497), .ZN(n3496) );
  NAND2_X1 U3465 ( .A1(n3355), .A2(n3498), .ZN(n3497) );
  NAND2_X1 U3466 ( .A1(n3357), .A2(n3356), .ZN(n3498) );
  XOR2_X1 U3467 ( .A(n3499), .B(n3500), .Z(n3355) );
  NAND2_X1 U3468 ( .A1(n3501), .A2(n3502), .ZN(n3499) );
  NOR2_X1 U3469 ( .A1(n3356), .A2(n3357), .ZN(n3495) );
  NOR2_X1 U3470 ( .A1(n3283), .A2(n2492), .ZN(n3357) );
  NAND2_X1 U3471 ( .A1(n3363), .A2(n3503), .ZN(n3356) );
  NAND2_X1 U3472 ( .A1(n3362), .A2(n3364), .ZN(n3503) );
  NAND2_X1 U3473 ( .A1(n3504), .A2(n3505), .ZN(n3364) );
  NAND2_X1 U3474 ( .A1(b_8_), .A2(a_11_), .ZN(n3505) );
  INV_X1 U3475 ( .A(n3506), .ZN(n3504) );
  XNOR2_X1 U3476 ( .A(n3507), .B(n3508), .ZN(n3362) );
  XOR2_X1 U3477 ( .A(n3509), .B(n3510), .Z(n3508) );
  NAND2_X1 U3478 ( .A1(b_7_), .A2(a_12_), .ZN(n3510) );
  NAND2_X1 U3479 ( .A1(a_11_), .A2(n3506), .ZN(n3363) );
  NAND2_X1 U3480 ( .A1(n3511), .A2(n3512), .ZN(n3506) );
  NAND2_X1 U3481 ( .A1(n3513), .A2(b_8_), .ZN(n3512) );
  NOR2_X1 U3482 ( .A1(n3514), .A2(n2490), .ZN(n3513) );
  NOR2_X1 U3483 ( .A1(n3370), .A2(n3372), .ZN(n3514) );
  NAND2_X1 U3484 ( .A1(n3370), .A2(n3372), .ZN(n3511) );
  NAND2_X1 U3485 ( .A1(n3515), .A2(n3516), .ZN(n3372) );
  NAND2_X1 U3486 ( .A1(n3517), .A2(b_8_), .ZN(n3516) );
  NOR2_X1 U3487 ( .A1(n3518), .A2(n2252), .ZN(n3517) );
  NOR2_X1 U3488 ( .A1(n3519), .A2(n3393), .ZN(n3518) );
  NAND2_X1 U3489 ( .A1(n3519), .A2(n3393), .ZN(n3515) );
  NAND2_X1 U3490 ( .A1(n3520), .A2(n3521), .ZN(n3393) );
  NAND2_X1 U3491 ( .A1(b_6_), .A2(n3522), .ZN(n3521) );
  NAND2_X1 U3492 ( .A1(n2227), .A2(n3523), .ZN(n3522) );
  NAND2_X1 U3493 ( .A1(a_15_), .A2(n2343), .ZN(n3523) );
  NAND2_X1 U3494 ( .A1(b_7_), .A2(n3524), .ZN(n3520) );
  NAND2_X1 U3495 ( .A1(n2231), .A2(n3525), .ZN(n3524) );
  NAND2_X1 U3496 ( .A1(a_14_), .A2(n2494), .ZN(n3525) );
  INV_X1 U3497 ( .A(n3392), .ZN(n3519) );
  NAND2_X1 U3498 ( .A1(n3526), .A2(n2488), .ZN(n3392) );
  NOR2_X1 U3499 ( .A1(n2343), .A2(n3283), .ZN(n3526) );
  XOR2_X1 U3500 ( .A(n3527), .B(n3528), .Z(n3370) );
  XOR2_X1 U3501 ( .A(n3529), .B(n3530), .Z(n3528) );
  NAND2_X1 U3502 ( .A1(b_7_), .A2(a_13_), .ZN(n3527) );
  XNOR2_X1 U3503 ( .A(n3531), .B(n3532), .ZN(n3394) );
  XOR2_X1 U3504 ( .A(n3533), .B(n3534), .Z(n3531) );
  XNOR2_X1 U3505 ( .A(n3535), .B(n3536), .ZN(n3334) );
  XNOR2_X1 U3506 ( .A(n2337), .B(n3537), .ZN(n3535) );
  XNOR2_X1 U3507 ( .A(n3538), .B(n3539), .ZN(n3325) );
  NAND2_X1 U3508 ( .A1(n3540), .A2(n3541), .ZN(n3538) );
  XNOR2_X1 U3509 ( .A(n3542), .B(n3543), .ZN(n3410) );
  XOR2_X1 U3510 ( .A(n3544), .B(n3545), .Z(n3543) );
  NAND2_X1 U3511 ( .A1(a_4_), .A2(b_7_), .ZN(n3545) );
  XNOR2_X1 U3512 ( .A(n3546), .B(n3547), .ZN(n3422) );
  XOR2_X1 U3513 ( .A(n3548), .B(n3549), .Z(n3547) );
  NAND2_X1 U3514 ( .A1(b_7_), .A2(a_1_), .ZN(n3549) );
  INV_X1 U3515 ( .A(n3550), .ZN(n3425) );
  NAND2_X1 U3516 ( .A1(n3428), .A2(n3429), .ZN(n3550) );
  NAND2_X1 U3517 ( .A1(n3433), .A2(n3551), .ZN(n3429) );
  NAND2_X1 U3518 ( .A1(n3432), .A2(n3434), .ZN(n3551) );
  NAND2_X1 U3519 ( .A1(n3552), .A2(n3553), .ZN(n3434) );
  NAND2_X1 U3520 ( .A1(a_0_), .A2(b_7_), .ZN(n3553) );
  INV_X1 U3521 ( .A(n3554), .ZN(n3552) );
  XNOR2_X1 U3522 ( .A(n3555), .B(n3556), .ZN(n3432) );
  XNOR2_X1 U3523 ( .A(n3557), .B(n3558), .ZN(n3556) );
  NAND2_X1 U3524 ( .A1(a_0_), .A2(n3554), .ZN(n3433) );
  NAND2_X1 U3525 ( .A1(n3559), .A2(n3560), .ZN(n3554) );
  NAND2_X1 U3526 ( .A1(n3561), .A2(b_7_), .ZN(n3560) );
  NOR2_X1 U3527 ( .A1(n3562), .A2(n2500), .ZN(n3561) );
  NOR2_X1 U3528 ( .A1(n3548), .A2(n3546), .ZN(n3562) );
  NAND2_X1 U3529 ( .A1(n3546), .A2(n3548), .ZN(n3559) );
  NAND2_X1 U3530 ( .A1(n3563), .A2(n3564), .ZN(n3548) );
  NAND2_X1 U3531 ( .A1(n3565), .A2(a_2_), .ZN(n3564) );
  NOR2_X1 U3532 ( .A1(n3566), .A2(n2343), .ZN(n3565) );
  NOR2_X1 U3533 ( .A1(n3443), .A2(n3445), .ZN(n3566) );
  NAND2_X1 U3534 ( .A1(n3443), .A2(n3445), .ZN(n3563) );
  NAND2_X1 U3535 ( .A1(n3567), .A2(n3568), .ZN(n3445) );
  NAND2_X1 U3536 ( .A1(n3569), .A2(a_3_), .ZN(n3568) );
  NOR2_X1 U3537 ( .A1(n3570), .A2(n2343), .ZN(n3569) );
  NOR2_X1 U3538 ( .A1(n3451), .A2(n3453), .ZN(n3570) );
  NAND2_X1 U3539 ( .A1(n3451), .A2(n3453), .ZN(n3567) );
  NAND2_X1 U3540 ( .A1(n3571), .A2(n3572), .ZN(n3453) );
  NAND2_X1 U3541 ( .A1(n3573), .A2(a_4_), .ZN(n3572) );
  NOR2_X1 U3542 ( .A1(n3574), .A2(n2343), .ZN(n3573) );
  NOR2_X1 U3543 ( .A1(n3542), .A2(n3544), .ZN(n3574) );
  NAND2_X1 U3544 ( .A1(n3542), .A2(n3544), .ZN(n3571) );
  NAND2_X1 U3545 ( .A1(n3465), .A2(n3575), .ZN(n3544) );
  NAND2_X1 U3546 ( .A1(n3464), .A2(n3466), .ZN(n3575) );
  NAND2_X1 U3547 ( .A1(n3576), .A2(n3577), .ZN(n3466) );
  NAND2_X1 U3548 ( .A1(a_5_), .A2(b_7_), .ZN(n3577) );
  INV_X1 U3549 ( .A(n3578), .ZN(n3576) );
  XOR2_X1 U3550 ( .A(n3579), .B(n3580), .Z(n3464) );
  XOR2_X1 U3551 ( .A(n3581), .B(n3582), .Z(n3580) );
  NAND2_X1 U3552 ( .A1(a_5_), .A2(n3578), .ZN(n3465) );
  NAND2_X1 U3553 ( .A1(n3540), .A2(n3583), .ZN(n3578) );
  NAND2_X1 U3554 ( .A1(n3539), .A2(n3541), .ZN(n3583) );
  NAND2_X1 U3555 ( .A1(n3584), .A2(n3585), .ZN(n3541) );
  NAND2_X1 U3556 ( .A1(a_6_), .A2(b_7_), .ZN(n3585) );
  XNOR2_X1 U3557 ( .A(n3586), .B(n3587), .ZN(n3539) );
  XOR2_X1 U3558 ( .A(n3588), .B(n3589), .Z(n3587) );
  NAND2_X1 U3559 ( .A1(b_6_), .A2(a_7_), .ZN(n3589) );
  NAND2_X1 U3560 ( .A1(n3590), .A2(a_6_), .ZN(n3540) );
  INV_X1 U3561 ( .A(n3584), .ZN(n3590) );
  NAND2_X1 U3562 ( .A1(n3591), .A2(n3592), .ZN(n3584) );
  NAND2_X1 U3563 ( .A1(n3536), .A2(n3593), .ZN(n3592) );
  INV_X1 U3564 ( .A(n3594), .ZN(n3593) );
  NOR2_X1 U3565 ( .A1(n2468), .A2(n3537), .ZN(n3594) );
  XOR2_X1 U3566 ( .A(n3595), .B(n3596), .Z(n3536) );
  XOR2_X1 U3567 ( .A(n3597), .B(n3598), .Z(n3596) );
  NAND2_X1 U3568 ( .A1(b_6_), .A2(a_8_), .ZN(n3598) );
  NAND2_X1 U3569 ( .A1(n3537), .A2(n2468), .ZN(n3591) );
  INV_X1 U3570 ( .A(n2337), .ZN(n2468) );
  NOR2_X1 U3571 ( .A1(n2342), .A2(n2343), .ZN(n2337) );
  NOR2_X1 U3572 ( .A1(n3599), .A2(n3600), .ZN(n3537) );
  INV_X1 U3573 ( .A(n3601), .ZN(n3600) );
  NAND2_X1 U3574 ( .A1(n3482), .A2(n3602), .ZN(n3601) );
  NAND2_X1 U3575 ( .A1(n3481), .A2(n3479), .ZN(n3602) );
  NOR2_X1 U3576 ( .A1(n2343), .A2(n3349), .ZN(n3482) );
  NOR2_X1 U3577 ( .A1(n3479), .A2(n3481), .ZN(n3599) );
  NOR2_X1 U3578 ( .A1(n3603), .A2(n3604), .ZN(n3481) );
  INV_X1 U3579 ( .A(n3605), .ZN(n3604) );
  NAND2_X1 U3580 ( .A1(n3489), .A2(n3606), .ZN(n3605) );
  NAND2_X1 U3581 ( .A1(n3486), .A2(n3488), .ZN(n3606) );
  NOR2_X1 U3582 ( .A1(n2343), .A2(n2311), .ZN(n3489) );
  NOR2_X1 U3583 ( .A1(n3486), .A2(n3488), .ZN(n3603) );
  NAND2_X1 U3584 ( .A1(n3607), .A2(n3608), .ZN(n3488) );
  NAND2_X1 U3585 ( .A1(n3532), .A2(n3609), .ZN(n3608) );
  NAND2_X1 U3586 ( .A1(n3534), .A2(n3533), .ZN(n3609) );
  XOR2_X1 U3587 ( .A(n3610), .B(n3611), .Z(n3532) );
  NAND2_X1 U3588 ( .A1(n3612), .A2(n3613), .ZN(n3610) );
  INV_X1 U3589 ( .A(n3614), .ZN(n3607) );
  NOR2_X1 U3590 ( .A1(n3533), .A2(n3534), .ZN(n3614) );
  NOR2_X1 U3591 ( .A1(n2343), .A2(n2492), .ZN(n3534) );
  NAND2_X1 U3592 ( .A1(n3501), .A2(n3615), .ZN(n3533) );
  NAND2_X1 U3593 ( .A1(n3500), .A2(n3502), .ZN(n3615) );
  NAND2_X1 U3594 ( .A1(n3616), .A2(n3617), .ZN(n3502) );
  NAND2_X1 U3595 ( .A1(b_7_), .A2(a_11_), .ZN(n3617) );
  INV_X1 U3596 ( .A(n3618), .ZN(n3616) );
  XNOR2_X1 U3597 ( .A(n3619), .B(n3620), .ZN(n3500) );
  XOR2_X1 U3598 ( .A(n3621), .B(n3622), .Z(n3620) );
  NAND2_X1 U3599 ( .A1(b_6_), .A2(a_12_), .ZN(n3622) );
  NAND2_X1 U3600 ( .A1(a_11_), .A2(n3618), .ZN(n3501) );
  NAND2_X1 U3601 ( .A1(n3623), .A2(n3624), .ZN(n3618) );
  NAND2_X1 U3602 ( .A1(n3625), .A2(b_7_), .ZN(n3624) );
  NOR2_X1 U3603 ( .A1(n3626), .A2(n2490), .ZN(n3625) );
  NOR2_X1 U3604 ( .A1(n3507), .A2(n3509), .ZN(n3626) );
  NAND2_X1 U3605 ( .A1(n3507), .A2(n3509), .ZN(n3623) );
  NAND2_X1 U3606 ( .A1(n3627), .A2(n3628), .ZN(n3509) );
  NAND2_X1 U3607 ( .A1(n3629), .A2(b_7_), .ZN(n3628) );
  NOR2_X1 U3608 ( .A1(n3630), .A2(n2252), .ZN(n3629) );
  NOR2_X1 U3609 ( .A1(n3631), .A2(n3530), .ZN(n3630) );
  NAND2_X1 U3610 ( .A1(n3631), .A2(n3530), .ZN(n3627) );
  NAND2_X1 U3611 ( .A1(n3632), .A2(n3633), .ZN(n3530) );
  NAND2_X1 U3612 ( .A1(b_5_), .A2(n3634), .ZN(n3633) );
  NAND2_X1 U3613 ( .A1(n2227), .A2(n3635), .ZN(n3634) );
  NAND2_X1 U3614 ( .A1(a_15_), .A2(n2494), .ZN(n3635) );
  NAND2_X1 U3615 ( .A1(b_6_), .A2(n3636), .ZN(n3632) );
  NAND2_X1 U3616 ( .A1(n2231), .A2(n3637), .ZN(n3636) );
  NAND2_X1 U3617 ( .A1(a_14_), .A2(n2374), .ZN(n3637) );
  INV_X1 U3618 ( .A(n3529), .ZN(n3631) );
  NAND2_X1 U3619 ( .A1(n3638), .A2(n2488), .ZN(n3529) );
  NOR2_X1 U3620 ( .A1(n2343), .A2(n2494), .ZN(n3638) );
  XOR2_X1 U3621 ( .A(n3639), .B(n3640), .Z(n3507) );
  XOR2_X1 U3622 ( .A(n3641), .B(n3642), .Z(n3640) );
  NAND2_X1 U3623 ( .A1(b_6_), .A2(a_13_), .ZN(n3639) );
  XOR2_X1 U3624 ( .A(n3643), .B(n3644), .Z(n3486) );
  XOR2_X1 U3625 ( .A(n3645), .B(n3646), .Z(n3643) );
  XOR2_X1 U3626 ( .A(n3647), .B(n3648), .Z(n3479) );
  XNOR2_X1 U3627 ( .A(n3649), .B(n3650), .ZN(n3648) );
  XOR2_X1 U3628 ( .A(n3651), .B(n3652), .Z(n3542) );
  XOR2_X1 U3629 ( .A(n3653), .B(n3654), .Z(n3651) );
  XNOR2_X1 U3630 ( .A(n3655), .B(n3656), .ZN(n3451) );
  XNOR2_X1 U3631 ( .A(n3657), .B(n3658), .ZN(n3656) );
  XNOR2_X1 U3632 ( .A(n3659), .B(n3660), .ZN(n3443) );
  XNOR2_X1 U3633 ( .A(n3661), .B(n3662), .ZN(n3660) );
  XOR2_X1 U3634 ( .A(n3663), .B(n3664), .Z(n3546) );
  XOR2_X1 U3635 ( .A(n3665), .B(n3666), .Z(n3663) );
  XNOR2_X1 U3636 ( .A(n3667), .B(n3668), .ZN(n3428) );
  XNOR2_X1 U3637 ( .A(n3669), .B(n3670), .ZN(n3667) );
  NOR2_X1 U3638 ( .A1(n3671), .A2(n2201), .ZN(n2544) );
  INV_X1 U3639 ( .A(n3672), .ZN(n2201) );
  NAND2_X1 U3640 ( .A1(n2203), .A2(n2204), .ZN(n3672) );
  NOR2_X1 U3641 ( .A1(n3673), .A2(n3671), .ZN(n2204) );
  NOR2_X1 U3642 ( .A1(n3674), .A2(n3675), .ZN(n3673) );
  NOR2_X1 U3643 ( .A1(n3676), .A2(n2548), .ZN(n2203) );
  XOR2_X1 U3644 ( .A(n3677), .B(n3678), .Z(n2548) );
  XOR2_X1 U3645 ( .A(n3679), .B(n3680), .Z(n3678) );
  NAND2_X1 U3646 ( .A1(a_0_), .A2(b_5_), .ZN(n3680) );
  INV_X1 U3647 ( .A(n2547), .ZN(n3676) );
  NAND2_X1 U3648 ( .A1(n3681), .A2(n3682), .ZN(n2547) );
  NAND2_X1 U3649 ( .A1(n3670), .A2(n3683), .ZN(n3682) );
  INV_X1 U3650 ( .A(n3684), .ZN(n3683) );
  NOR2_X1 U3651 ( .A1(n3669), .A2(n3668), .ZN(n3684) );
  NOR2_X1 U3652 ( .A1(n3191), .A2(n2494), .ZN(n3670) );
  NAND2_X1 U3653 ( .A1(n3668), .A2(n3669), .ZN(n3681) );
  NAND2_X1 U3654 ( .A1(n3685), .A2(n3686), .ZN(n3669) );
  NAND2_X1 U3655 ( .A1(n3558), .A2(n3687), .ZN(n3686) );
  INV_X1 U3656 ( .A(n3688), .ZN(n3687) );
  NOR2_X1 U3657 ( .A1(n3555), .A2(n3557), .ZN(n3688) );
  NOR2_X1 U3658 ( .A1(n2494), .A2(n2500), .ZN(n3558) );
  NAND2_X1 U3659 ( .A1(n3555), .A2(n3557), .ZN(n3685) );
  NAND2_X1 U3660 ( .A1(n3689), .A2(n3690), .ZN(n3557) );
  NAND2_X1 U3661 ( .A1(n3665), .A2(n3691), .ZN(n3690) );
  INV_X1 U3662 ( .A(n3692), .ZN(n3691) );
  NOR2_X1 U3663 ( .A1(n3666), .A2(n3664), .ZN(n3692) );
  NOR2_X1 U3664 ( .A1(n2426), .A2(n2494), .ZN(n3665) );
  NAND2_X1 U3665 ( .A1(n3664), .A2(n3666), .ZN(n3689) );
  NAND2_X1 U3666 ( .A1(n3693), .A2(n3694), .ZN(n3666) );
  NAND2_X1 U3667 ( .A1(n3662), .A2(n3695), .ZN(n3694) );
  INV_X1 U3668 ( .A(n3696), .ZN(n3695) );
  NOR2_X1 U3669 ( .A1(n3659), .A2(n3661), .ZN(n3696) );
  NOR2_X1 U3670 ( .A1(n2410), .A2(n2494), .ZN(n3662) );
  NAND2_X1 U3671 ( .A1(n3659), .A2(n3661), .ZN(n3693) );
  NAND2_X1 U3672 ( .A1(n3697), .A2(n3698), .ZN(n3661) );
  NAND2_X1 U3673 ( .A1(n3658), .A2(n3699), .ZN(n3698) );
  INV_X1 U3674 ( .A(n3700), .ZN(n3699) );
  NOR2_X1 U3675 ( .A1(n3655), .A2(n3657), .ZN(n3700) );
  NOR2_X1 U3676 ( .A1(n2497), .A2(n2494), .ZN(n3658) );
  NAND2_X1 U3677 ( .A1(n3655), .A2(n3657), .ZN(n3697) );
  NAND2_X1 U3678 ( .A1(n3701), .A2(n3702), .ZN(n3657) );
  NAND2_X1 U3679 ( .A1(n3654), .A2(n3703), .ZN(n3702) );
  NAND2_X1 U3680 ( .A1(n3652), .A2(n3653), .ZN(n3703) );
  NOR2_X1 U3681 ( .A1(n2373), .A2(n2494), .ZN(n3654) );
  INV_X1 U3682 ( .A(n3704), .ZN(n3701) );
  NOR2_X1 U3683 ( .A1(n3652), .A2(n3653), .ZN(n3704) );
  NAND2_X1 U3684 ( .A1(n3705), .A2(n3706), .ZN(n3653) );
  NAND2_X1 U3685 ( .A1(n3579), .A2(n3707), .ZN(n3706) );
  NAND2_X1 U3686 ( .A1(n3582), .A2(n3708), .ZN(n3707) );
  XOR2_X1 U3687 ( .A(n3709), .B(n3710), .Z(n3579) );
  XOR2_X1 U3688 ( .A(n3711), .B(n3712), .Z(n3710) );
  NAND2_X1 U3689 ( .A1(b_5_), .A2(a_7_), .ZN(n3712) );
  NAND2_X1 U3690 ( .A1(n3581), .A2(n2362), .ZN(n3705) );
  INV_X1 U3691 ( .A(n3582), .ZN(n2362) );
  NOR2_X1 U3692 ( .A1(n2494), .A2(n2495), .ZN(n3582) );
  INV_X1 U3693 ( .A(n3708), .ZN(n3581) );
  NAND2_X1 U3694 ( .A1(n3713), .A2(n3714), .ZN(n3708) );
  NAND2_X1 U3695 ( .A1(n3715), .A2(b_6_), .ZN(n3714) );
  NOR2_X1 U3696 ( .A1(n3716), .A2(n2342), .ZN(n3715) );
  NOR2_X1 U3697 ( .A1(n3586), .A2(n3588), .ZN(n3716) );
  NAND2_X1 U3698 ( .A1(n3586), .A2(n3588), .ZN(n3713) );
  NAND2_X1 U3699 ( .A1(n3717), .A2(n3718), .ZN(n3588) );
  NAND2_X1 U3700 ( .A1(n3719), .A2(b_6_), .ZN(n3718) );
  NOR2_X1 U3701 ( .A1(n3720), .A2(n3349), .ZN(n3719) );
  NOR2_X1 U3702 ( .A1(n3597), .A2(n3595), .ZN(n3720) );
  NAND2_X1 U3703 ( .A1(n3595), .A2(n3597), .ZN(n3717) );
  NAND2_X1 U3704 ( .A1(n3721), .A2(n3722), .ZN(n3597) );
  NAND2_X1 U3705 ( .A1(n3650), .A2(n3723), .ZN(n3722) );
  NAND2_X1 U3706 ( .A1(n3647), .A2(n3649), .ZN(n3723) );
  NOR2_X1 U3707 ( .A1(n2494), .A2(n2311), .ZN(n3650) );
  INV_X1 U3708 ( .A(n3724), .ZN(n3721) );
  NOR2_X1 U3709 ( .A1(n3647), .A2(n3649), .ZN(n3724) );
  NAND2_X1 U3710 ( .A1(n3725), .A2(n3726), .ZN(n3649) );
  NAND2_X1 U3711 ( .A1(n3644), .A2(n3727), .ZN(n3726) );
  NAND2_X1 U3712 ( .A1(n3646), .A2(n3645), .ZN(n3727) );
  XOR2_X1 U3713 ( .A(n3728), .B(n3729), .Z(n3644) );
  NAND2_X1 U3714 ( .A1(n3730), .A2(n3731), .ZN(n3728) );
  INV_X1 U3715 ( .A(n3732), .ZN(n3725) );
  NOR2_X1 U3716 ( .A1(n3645), .A2(n3646), .ZN(n3732) );
  NOR2_X1 U3717 ( .A1(n2494), .A2(n2492), .ZN(n3646) );
  NAND2_X1 U3718 ( .A1(n3612), .A2(n3733), .ZN(n3645) );
  NAND2_X1 U3719 ( .A1(n3611), .A2(n3613), .ZN(n3733) );
  NAND2_X1 U3720 ( .A1(n3734), .A2(n3735), .ZN(n3613) );
  NAND2_X1 U3721 ( .A1(b_6_), .A2(a_11_), .ZN(n3735) );
  INV_X1 U3722 ( .A(n3736), .ZN(n3734) );
  XNOR2_X1 U3723 ( .A(n3737), .B(n3738), .ZN(n3611) );
  XOR2_X1 U3724 ( .A(n3739), .B(n3740), .Z(n3738) );
  NAND2_X1 U3725 ( .A1(b_5_), .A2(a_12_), .ZN(n3740) );
  NAND2_X1 U3726 ( .A1(a_11_), .A2(n3736), .ZN(n3612) );
  NAND2_X1 U3727 ( .A1(n3741), .A2(n3742), .ZN(n3736) );
  NAND2_X1 U3728 ( .A1(n3743), .A2(b_6_), .ZN(n3742) );
  NOR2_X1 U3729 ( .A1(n3744), .A2(n2490), .ZN(n3743) );
  NOR2_X1 U3730 ( .A1(n3619), .A2(n3621), .ZN(n3744) );
  NAND2_X1 U3731 ( .A1(n3619), .A2(n3621), .ZN(n3741) );
  NAND2_X1 U3732 ( .A1(n3745), .A2(n3746), .ZN(n3621) );
  NAND2_X1 U3733 ( .A1(n3747), .A2(b_6_), .ZN(n3746) );
  NOR2_X1 U3734 ( .A1(n3748), .A2(n2252), .ZN(n3747) );
  NOR2_X1 U3735 ( .A1(n3749), .A2(n3642), .ZN(n3748) );
  NAND2_X1 U3736 ( .A1(n3749), .A2(n3642), .ZN(n3745) );
  NAND2_X1 U3737 ( .A1(n3750), .A2(n3751), .ZN(n3642) );
  NAND2_X1 U3738 ( .A1(b_4_), .A2(n3752), .ZN(n3751) );
  NAND2_X1 U3739 ( .A1(n2227), .A2(n3753), .ZN(n3752) );
  NAND2_X1 U3740 ( .A1(a_15_), .A2(n2374), .ZN(n3753) );
  NAND2_X1 U3741 ( .A1(b_5_), .A2(n3754), .ZN(n3750) );
  NAND2_X1 U3742 ( .A1(n2231), .A2(n3755), .ZN(n3754) );
  NAND2_X1 U3743 ( .A1(a_14_), .A2(n2496), .ZN(n3755) );
  INV_X1 U3744 ( .A(n3641), .ZN(n3749) );
  NAND2_X1 U3745 ( .A1(n3756), .A2(n2488), .ZN(n3641) );
  NOR2_X1 U3746 ( .A1(n2374), .A2(n2494), .ZN(n3756) );
  XOR2_X1 U3747 ( .A(n3757), .B(n3758), .Z(n3619) );
  XOR2_X1 U3748 ( .A(n3759), .B(n3760), .Z(n3758) );
  NAND2_X1 U3749 ( .A1(b_5_), .A2(a_13_), .ZN(n3757) );
  XOR2_X1 U3750 ( .A(n3761), .B(n3762), .Z(n3647) );
  XOR2_X1 U3751 ( .A(n3763), .B(n3764), .Z(n3761) );
  XNOR2_X1 U3752 ( .A(n3765), .B(n3766), .ZN(n3595) );
  XNOR2_X1 U3753 ( .A(n3767), .B(n3768), .ZN(n3766) );
  XNOR2_X1 U3754 ( .A(n3769), .B(n3770), .ZN(n3586) );
  NAND2_X1 U3755 ( .A1(n3771), .A2(n3772), .ZN(n3769) );
  XNOR2_X1 U3756 ( .A(n3773), .B(n3774), .ZN(n3652) );
  XOR2_X1 U3757 ( .A(n3775), .B(n3776), .Z(n3773) );
  NOR2_X1 U3758 ( .A1(n2495), .A2(n2374), .ZN(n3776) );
  XNOR2_X1 U3759 ( .A(n3777), .B(n3778), .ZN(n3655) );
  XOR2_X1 U3760 ( .A(n3779), .B(n2368), .Z(n3777) );
  XOR2_X1 U3761 ( .A(n3780), .B(n3781), .Z(n3659) );
  XNOR2_X1 U3762 ( .A(n3782), .B(n3783), .ZN(n3781) );
  NAND2_X1 U3763 ( .A1(a_4_), .A2(b_5_), .ZN(n3783) );
  XOR2_X1 U3764 ( .A(n3784), .B(n3785), .Z(n3664) );
  XNOR2_X1 U3765 ( .A(n3786), .B(n3787), .ZN(n3784) );
  NAND2_X1 U3766 ( .A1(a_3_), .A2(b_5_), .ZN(n3786) );
  XOR2_X1 U3767 ( .A(n3788), .B(n3789), .Z(n3555) );
  XNOR2_X1 U3768 ( .A(n3790), .B(n3791), .ZN(n3788) );
  NAND2_X1 U3769 ( .A1(a_2_), .A2(b_5_), .ZN(n3790) );
  XNOR2_X1 U3770 ( .A(n3792), .B(n3793), .ZN(n3668) );
  XOR2_X1 U3771 ( .A(n3794), .B(n3795), .Z(n3793) );
  NAND2_X1 U3772 ( .A1(b_5_), .A2(a_1_), .ZN(n3795) );
  INV_X1 U3773 ( .A(n3796), .ZN(n3671) );
  NAND2_X1 U3774 ( .A1(n3674), .A2(n3675), .ZN(n3796) );
  NAND2_X1 U3775 ( .A1(n3797), .A2(n3798), .ZN(n3675) );
  NAND2_X1 U3776 ( .A1(n3799), .A2(a_0_), .ZN(n3798) );
  NOR2_X1 U3777 ( .A1(n3800), .A2(n2374), .ZN(n3799) );
  NOR2_X1 U3778 ( .A1(n3677), .A2(n3679), .ZN(n3800) );
  NAND2_X1 U3779 ( .A1(n3677), .A2(n3679), .ZN(n3797) );
  NAND2_X1 U3780 ( .A1(n3801), .A2(n3802), .ZN(n3679) );
  NAND2_X1 U3781 ( .A1(n3803), .A2(b_5_), .ZN(n3802) );
  NOR2_X1 U3782 ( .A1(n3804), .A2(n2500), .ZN(n3803) );
  NOR2_X1 U3783 ( .A1(n3794), .A2(n3792), .ZN(n3804) );
  NAND2_X1 U3784 ( .A1(n3792), .A2(n3794), .ZN(n3801) );
  NAND2_X1 U3785 ( .A1(n3805), .A2(n3806), .ZN(n3794) );
  NAND2_X1 U3786 ( .A1(n3807), .A2(a_2_), .ZN(n3806) );
  NOR2_X1 U3787 ( .A1(n3808), .A2(n2374), .ZN(n3807) );
  NOR2_X1 U3788 ( .A1(n3789), .A2(n3791), .ZN(n3808) );
  NAND2_X1 U3789 ( .A1(n3789), .A2(n3791), .ZN(n3805) );
  NAND2_X1 U3790 ( .A1(n3809), .A2(n3810), .ZN(n3791) );
  NAND2_X1 U3791 ( .A1(n3811), .A2(a_3_), .ZN(n3810) );
  NOR2_X1 U3792 ( .A1(n3812), .A2(n2374), .ZN(n3811) );
  NOR2_X1 U3793 ( .A1(n3787), .A2(n3785), .ZN(n3812) );
  NAND2_X1 U3794 ( .A1(n3785), .A2(n3787), .ZN(n3809) );
  NAND2_X1 U3795 ( .A1(n3813), .A2(n3814), .ZN(n3787) );
  NAND2_X1 U3796 ( .A1(n3815), .A2(a_4_), .ZN(n3814) );
  NOR2_X1 U3797 ( .A1(n3816), .A2(n2374), .ZN(n3815) );
  NOR2_X1 U3798 ( .A1(n3782), .A2(n3780), .ZN(n3816) );
  NAND2_X1 U3799 ( .A1(n3782), .A2(n3780), .ZN(n3813) );
  XOR2_X1 U3800 ( .A(n3817), .B(n3818), .Z(n3780) );
  XOR2_X1 U3801 ( .A(n3819), .B(n3820), .Z(n3817) );
  NOR2_X1 U3802 ( .A1(n3821), .A2(n3822), .ZN(n3782) );
  INV_X1 U3803 ( .A(n3823), .ZN(n3822) );
  NAND2_X1 U3804 ( .A1(n3778), .A2(n3824), .ZN(n3823) );
  NAND2_X1 U3805 ( .A1(n2368), .A2(n3779), .ZN(n3824) );
  XOR2_X1 U3806 ( .A(n3825), .B(n3826), .Z(n3778) );
  XOR2_X1 U3807 ( .A(n3827), .B(n3828), .Z(n3826) );
  NOR2_X1 U3808 ( .A1(n3779), .A2(n2368), .ZN(n3821) );
  INV_X1 U3809 ( .A(n2464), .ZN(n2368) );
  NAND2_X1 U3810 ( .A1(a_5_), .A2(b_5_), .ZN(n2464) );
  NAND2_X1 U3811 ( .A1(n3829), .A2(n3830), .ZN(n3779) );
  NAND2_X1 U3812 ( .A1(n3831), .A2(b_5_), .ZN(n3830) );
  NOR2_X1 U3813 ( .A1(n3832), .A2(n2495), .ZN(n3831) );
  NOR2_X1 U3814 ( .A1(n3775), .A2(n3774), .ZN(n3832) );
  NAND2_X1 U3815 ( .A1(n3774), .A2(n3775), .ZN(n3829) );
  NAND2_X1 U3816 ( .A1(n3833), .A2(n3834), .ZN(n3775) );
  NAND2_X1 U3817 ( .A1(n3835), .A2(b_5_), .ZN(n3834) );
  NOR2_X1 U3818 ( .A1(n3836), .A2(n2342), .ZN(n3835) );
  NOR2_X1 U3819 ( .A1(n3709), .A2(n3711), .ZN(n3836) );
  NAND2_X1 U3820 ( .A1(n3709), .A2(n3711), .ZN(n3833) );
  NAND2_X1 U3821 ( .A1(n3771), .A2(n3837), .ZN(n3711) );
  NAND2_X1 U3822 ( .A1(n3770), .A2(n3772), .ZN(n3837) );
  NAND2_X1 U3823 ( .A1(n3838), .A2(n3839), .ZN(n3772) );
  NAND2_X1 U3824 ( .A1(b_5_), .A2(a_8_), .ZN(n3839) );
  INV_X1 U3825 ( .A(n3840), .ZN(n3838) );
  XNOR2_X1 U3826 ( .A(n3841), .B(n3842), .ZN(n3770) );
  XNOR2_X1 U3827 ( .A(n3843), .B(n3844), .ZN(n3842) );
  NAND2_X1 U3828 ( .A1(a_8_), .A2(n3840), .ZN(n3771) );
  NAND2_X1 U3829 ( .A1(n3845), .A2(n3846), .ZN(n3840) );
  NAND2_X1 U3830 ( .A1(n3768), .A2(n3847), .ZN(n3846) );
  NAND2_X1 U3831 ( .A1(n3765), .A2(n3767), .ZN(n3847) );
  NOR2_X1 U3832 ( .A1(n2374), .A2(n2311), .ZN(n3768) );
  INV_X1 U3833 ( .A(n3848), .ZN(n3845) );
  NOR2_X1 U3834 ( .A1(n3767), .A2(n3765), .ZN(n3848) );
  XOR2_X1 U3835 ( .A(n3849), .B(n3850), .Z(n3765) );
  XOR2_X1 U3836 ( .A(n3851), .B(n3852), .Z(n3849) );
  NAND2_X1 U3837 ( .A1(n3853), .A2(n3854), .ZN(n3767) );
  NAND2_X1 U3838 ( .A1(n3762), .A2(n3855), .ZN(n3854) );
  NAND2_X1 U3839 ( .A1(n3764), .A2(n3763), .ZN(n3855) );
  XOR2_X1 U3840 ( .A(n3856), .B(n3857), .Z(n3762) );
  NAND2_X1 U3841 ( .A1(n3858), .A2(n3859), .ZN(n3856) );
  INV_X1 U3842 ( .A(n3860), .ZN(n3853) );
  NOR2_X1 U3843 ( .A1(n3763), .A2(n3764), .ZN(n3860) );
  NOR2_X1 U3844 ( .A1(n2374), .A2(n2492), .ZN(n3764) );
  NAND2_X1 U3845 ( .A1(n3730), .A2(n3861), .ZN(n3763) );
  NAND2_X1 U3846 ( .A1(n3729), .A2(n3731), .ZN(n3861) );
  NAND2_X1 U3847 ( .A1(n3862), .A2(n3863), .ZN(n3731) );
  NAND2_X1 U3848 ( .A1(b_5_), .A2(a_11_), .ZN(n3863) );
  INV_X1 U3849 ( .A(n3864), .ZN(n3862) );
  XNOR2_X1 U3850 ( .A(n3865), .B(n3866), .ZN(n3729) );
  XOR2_X1 U3851 ( .A(n3867), .B(n3868), .Z(n3866) );
  NAND2_X1 U3852 ( .A1(b_4_), .A2(a_12_), .ZN(n3868) );
  NAND2_X1 U3853 ( .A1(a_11_), .A2(n3864), .ZN(n3730) );
  NAND2_X1 U3854 ( .A1(n3869), .A2(n3870), .ZN(n3864) );
  NAND2_X1 U3855 ( .A1(n3871), .A2(b_5_), .ZN(n3870) );
  NOR2_X1 U3856 ( .A1(n3872), .A2(n2490), .ZN(n3871) );
  NOR2_X1 U3857 ( .A1(n3737), .A2(n3739), .ZN(n3872) );
  NAND2_X1 U3858 ( .A1(n3737), .A2(n3739), .ZN(n3869) );
  NAND2_X1 U3859 ( .A1(n3873), .A2(n3874), .ZN(n3739) );
  NAND2_X1 U3860 ( .A1(n3875), .A2(b_5_), .ZN(n3874) );
  NOR2_X1 U3861 ( .A1(n3876), .A2(n2252), .ZN(n3875) );
  NOR2_X1 U3862 ( .A1(n3877), .A2(n3760), .ZN(n3876) );
  NAND2_X1 U3863 ( .A1(n3877), .A2(n3760), .ZN(n3873) );
  NAND2_X1 U3864 ( .A1(n3878), .A2(n3879), .ZN(n3760) );
  NAND2_X1 U3865 ( .A1(b_3_), .A2(n3880), .ZN(n3879) );
  NAND2_X1 U3866 ( .A1(n2227), .A2(n3881), .ZN(n3880) );
  NAND2_X1 U3867 ( .A1(a_15_), .A2(n2496), .ZN(n3881) );
  NAND2_X1 U3868 ( .A1(b_4_), .A2(n3882), .ZN(n3878) );
  NAND2_X1 U3869 ( .A1(n2231), .A2(n3883), .ZN(n3882) );
  NAND2_X1 U3870 ( .A1(a_14_), .A2(n2411), .ZN(n3883) );
  INV_X1 U3871 ( .A(n3759), .ZN(n3877) );
  NAND2_X1 U3872 ( .A1(n3884), .A2(n2488), .ZN(n3759) );
  NOR2_X1 U3873 ( .A1(n2374), .A2(n2496), .ZN(n3884) );
  XOR2_X1 U3874 ( .A(n3885), .B(n3886), .Z(n3737) );
  XOR2_X1 U3875 ( .A(n3887), .B(n3888), .Z(n3886) );
  NAND2_X1 U3876 ( .A1(b_4_), .A2(a_13_), .ZN(n3885) );
  XNOR2_X1 U3877 ( .A(n3889), .B(n3890), .ZN(n3709) );
  XNOR2_X1 U3878 ( .A(n3891), .B(n3892), .ZN(n3889) );
  XNOR2_X1 U3879 ( .A(n3893), .B(n3894), .ZN(n3774) );
  XNOR2_X1 U3880 ( .A(n3895), .B(n3896), .ZN(n3893) );
  XOR2_X1 U3881 ( .A(n3897), .B(n3898), .Z(n3785) );
  XOR2_X1 U3882 ( .A(n3899), .B(n2393), .Z(n3898) );
  INV_X1 U3883 ( .A(n3900), .ZN(n2393) );
  XNOR2_X1 U3884 ( .A(n3901), .B(n3902), .ZN(n3789) );
  XNOR2_X1 U3885 ( .A(n3903), .B(n3904), .ZN(n3902) );
  XOR2_X1 U3886 ( .A(n3905), .B(n3906), .Z(n3792) );
  XOR2_X1 U3887 ( .A(n3907), .B(n3908), .Z(n3906) );
  XNOR2_X1 U3888 ( .A(n3909), .B(n3910), .ZN(n3677) );
  XNOR2_X1 U3889 ( .A(n3911), .B(n3912), .ZN(n3910) );
  XNOR2_X1 U3890 ( .A(n3913), .B(n3914), .ZN(n3674) );
  XNOR2_X1 U3891 ( .A(n3915), .B(n3916), .ZN(n3914) );
  NOR2_X1 U3892 ( .A1(n3917), .A2(n2211), .ZN(n2539) );
  INV_X1 U3893 ( .A(n3918), .ZN(n2211) );
  NAND2_X1 U3894 ( .A1(n2213), .A2(n2214), .ZN(n3918) );
  NOR2_X1 U3895 ( .A1(n3919), .A2(n3917), .ZN(n2214) );
  NOR2_X1 U3896 ( .A1(n3920), .A2(n3921), .ZN(n3919) );
  NOR2_X1 U3897 ( .A1(n2543), .A2(n2542), .ZN(n2213) );
  XNOR2_X1 U3898 ( .A(n3922), .B(n3923), .ZN(n2542) );
  XOR2_X1 U3899 ( .A(n3924), .B(n3925), .Z(n3922) );
  NOR2_X1 U3900 ( .A1(n2411), .A2(n3191), .ZN(n3925) );
  INV_X1 U3901 ( .A(n3926), .ZN(n2543) );
  NAND2_X1 U3902 ( .A1(n3927), .A2(n3928), .ZN(n3926) );
  NAND2_X1 U3903 ( .A1(n3916), .A2(n3929), .ZN(n3928) );
  INV_X1 U3904 ( .A(n3930), .ZN(n3929) );
  NOR2_X1 U3905 ( .A1(n3915), .A2(n3913), .ZN(n3930) );
  NOR2_X1 U3906 ( .A1(n3191), .A2(n2496), .ZN(n3916) );
  NAND2_X1 U3907 ( .A1(n3913), .A2(n3915), .ZN(n3927) );
  NAND2_X1 U3908 ( .A1(n3931), .A2(n3932), .ZN(n3915) );
  NAND2_X1 U3909 ( .A1(n3912), .A2(n3933), .ZN(n3932) );
  INV_X1 U3910 ( .A(n3934), .ZN(n3933) );
  NOR2_X1 U3911 ( .A1(n3909), .A2(n3911), .ZN(n3934) );
  NOR2_X1 U3912 ( .A1(n2496), .A2(n2500), .ZN(n3912) );
  NAND2_X1 U3913 ( .A1(n3909), .A2(n3911), .ZN(n3931) );
  NAND2_X1 U3914 ( .A1(n3935), .A2(n3936), .ZN(n3911) );
  NAND2_X1 U3915 ( .A1(n3908), .A2(n3937), .ZN(n3936) );
  NAND2_X1 U3916 ( .A1(n3907), .A2(n3905), .ZN(n3937) );
  NOR2_X1 U3917 ( .A1(n2426), .A2(n2496), .ZN(n3908) );
  INV_X1 U3918 ( .A(n3938), .ZN(n3935) );
  NOR2_X1 U3919 ( .A1(n3905), .A2(n3907), .ZN(n3938) );
  NOR2_X1 U3920 ( .A1(n3939), .A2(n3940), .ZN(n3907) );
  INV_X1 U3921 ( .A(n3941), .ZN(n3940) );
  NAND2_X1 U3922 ( .A1(n3904), .A2(n3942), .ZN(n3941) );
  NAND2_X1 U3923 ( .A1(n3901), .A2(n3903), .ZN(n3942) );
  NOR2_X1 U3924 ( .A1(n2410), .A2(n2496), .ZN(n3904) );
  NOR2_X1 U3925 ( .A1(n3901), .A2(n3903), .ZN(n3939) );
  NAND2_X1 U3926 ( .A1(n3943), .A2(n3944), .ZN(n3903) );
  NAND2_X1 U3927 ( .A1(n3897), .A2(n3945), .ZN(n3944) );
  NAND2_X1 U3928 ( .A1(n3900), .A2(n3899), .ZN(n3945) );
  XNOR2_X1 U3929 ( .A(n3946), .B(n3947), .ZN(n3897) );
  XOR2_X1 U3930 ( .A(n3948), .B(n3949), .Z(n3946) );
  NOR2_X1 U3931 ( .A1(n2373), .A2(n2411), .ZN(n3949) );
  INV_X1 U3932 ( .A(n3950), .ZN(n3943) );
  NOR2_X1 U3933 ( .A1(n3899), .A2(n3900), .ZN(n3950) );
  NOR2_X1 U3934 ( .A1(n2496), .A2(n2497), .ZN(n3900) );
  NAND2_X1 U3935 ( .A1(n3951), .A2(n3952), .ZN(n3899) );
  NAND2_X1 U3936 ( .A1(n3820), .A2(n3953), .ZN(n3952) );
  INV_X1 U3937 ( .A(n3954), .ZN(n3953) );
  NOR2_X1 U3938 ( .A1(n3819), .A2(n3818), .ZN(n3954) );
  NOR2_X1 U3939 ( .A1(n2496), .A2(n2373), .ZN(n3820) );
  NAND2_X1 U3940 ( .A1(n3818), .A2(n3819), .ZN(n3951) );
  NAND2_X1 U3941 ( .A1(n3955), .A2(n3956), .ZN(n3819) );
  NAND2_X1 U3942 ( .A1(n3828), .A2(n3957), .ZN(n3956) );
  NAND2_X1 U3943 ( .A1(n3958), .A2(n3827), .ZN(n3957) );
  INV_X1 U3944 ( .A(n3959), .ZN(n3827) );
  NOR2_X1 U3945 ( .A1(n2496), .A2(n2495), .ZN(n3828) );
  NAND2_X1 U3946 ( .A1(n3825), .A2(n3959), .ZN(n3955) );
  NAND2_X1 U3947 ( .A1(n3960), .A2(n3961), .ZN(n3959) );
  NAND2_X1 U3948 ( .A1(n3896), .A2(n3962), .ZN(n3961) );
  NAND2_X1 U3949 ( .A1(n3895), .A2(n3894), .ZN(n3962) );
  NOR2_X1 U3950 ( .A1(n2496), .A2(n2342), .ZN(n3896) );
  INV_X1 U3951 ( .A(n3963), .ZN(n3960) );
  NOR2_X1 U3952 ( .A1(n3894), .A2(n3895), .ZN(n3963) );
  NOR2_X1 U3953 ( .A1(n3964), .A2(n3965), .ZN(n3895) );
  INV_X1 U3954 ( .A(n3966), .ZN(n3965) );
  NAND2_X1 U3955 ( .A1(n3892), .A2(n3967), .ZN(n3966) );
  NAND2_X1 U3956 ( .A1(n3890), .A2(n3891), .ZN(n3967) );
  NOR2_X1 U3957 ( .A1(n2496), .A2(n3349), .ZN(n3892) );
  NOR2_X1 U3958 ( .A1(n3890), .A2(n3891), .ZN(n3964) );
  NOR2_X1 U3959 ( .A1(n3968), .A2(n3969), .ZN(n3891) );
  INV_X1 U3960 ( .A(n3970), .ZN(n3969) );
  NAND2_X1 U3961 ( .A1(n3844), .A2(n3971), .ZN(n3970) );
  NAND2_X1 U3962 ( .A1(n3841), .A2(n3843), .ZN(n3971) );
  NOR2_X1 U3963 ( .A1(n2496), .A2(n2311), .ZN(n3844) );
  NOR2_X1 U3964 ( .A1(n3841), .A2(n3843), .ZN(n3968) );
  NAND2_X1 U3965 ( .A1(n3972), .A2(n3973), .ZN(n3843) );
  NAND2_X1 U3966 ( .A1(n3850), .A2(n3974), .ZN(n3973) );
  NAND2_X1 U3967 ( .A1(n3852), .A2(n3851), .ZN(n3974) );
  XOR2_X1 U3968 ( .A(n3975), .B(n3976), .Z(n3850) );
  NAND2_X1 U3969 ( .A1(n3977), .A2(n3978), .ZN(n3975) );
  INV_X1 U3970 ( .A(n3979), .ZN(n3972) );
  NOR2_X1 U3971 ( .A1(n3851), .A2(n3852), .ZN(n3979) );
  NOR2_X1 U3972 ( .A1(n2496), .A2(n2492), .ZN(n3852) );
  NAND2_X1 U3973 ( .A1(n3858), .A2(n3980), .ZN(n3851) );
  NAND2_X1 U3974 ( .A1(n3857), .A2(n3859), .ZN(n3980) );
  NAND2_X1 U3975 ( .A1(n3981), .A2(n3982), .ZN(n3859) );
  NAND2_X1 U3976 ( .A1(b_4_), .A2(a_11_), .ZN(n3982) );
  INV_X1 U3977 ( .A(n3983), .ZN(n3981) );
  XNOR2_X1 U3978 ( .A(n3984), .B(n3985), .ZN(n3857) );
  XOR2_X1 U3979 ( .A(n3986), .B(n3987), .Z(n3985) );
  NAND2_X1 U3980 ( .A1(b_3_), .A2(a_12_), .ZN(n3987) );
  NAND2_X1 U3981 ( .A1(a_11_), .A2(n3983), .ZN(n3858) );
  NAND2_X1 U3982 ( .A1(n3988), .A2(n3989), .ZN(n3983) );
  NAND2_X1 U3983 ( .A1(n3990), .A2(b_4_), .ZN(n3989) );
  NOR2_X1 U3984 ( .A1(n3991), .A2(n2490), .ZN(n3990) );
  NOR2_X1 U3985 ( .A1(n3865), .A2(n3867), .ZN(n3991) );
  NAND2_X1 U3986 ( .A1(n3865), .A2(n3867), .ZN(n3988) );
  NAND2_X1 U3987 ( .A1(n3992), .A2(n3993), .ZN(n3867) );
  NAND2_X1 U3988 ( .A1(n3994), .A2(b_4_), .ZN(n3993) );
  NOR2_X1 U3989 ( .A1(n3995), .A2(n2252), .ZN(n3994) );
  NOR2_X1 U3990 ( .A1(n3996), .A2(n3888), .ZN(n3995) );
  NAND2_X1 U3991 ( .A1(n3996), .A2(n3888), .ZN(n3992) );
  NAND2_X1 U3992 ( .A1(n3997), .A2(n3998), .ZN(n3888) );
  NAND2_X1 U3993 ( .A1(b_2_), .A2(n3999), .ZN(n3998) );
  NAND2_X1 U3994 ( .A1(n2227), .A2(n4000), .ZN(n3999) );
  NAND2_X1 U3995 ( .A1(a_15_), .A2(n2411), .ZN(n4000) );
  NAND2_X1 U3996 ( .A1(b_3_), .A2(n4001), .ZN(n3997) );
  NAND2_X1 U3997 ( .A1(n2231), .A2(n4002), .ZN(n4001) );
  NAND2_X1 U3998 ( .A1(a_14_), .A2(n2498), .ZN(n4002) );
  INV_X1 U3999 ( .A(n3887), .ZN(n3996) );
  NAND2_X1 U4000 ( .A1(n4003), .A2(n2488), .ZN(n3887) );
  NOR2_X1 U4001 ( .A1(n2411), .A2(n2496), .ZN(n4003) );
  XOR2_X1 U4002 ( .A(n4004), .B(n4005), .Z(n3865) );
  XOR2_X1 U4003 ( .A(n4006), .B(n4007), .Z(n4005) );
  NAND2_X1 U4004 ( .A1(b_3_), .A2(a_13_), .ZN(n4004) );
  XOR2_X1 U4005 ( .A(n4008), .B(n4009), .Z(n3841) );
  NAND2_X1 U4006 ( .A1(n4010), .A2(n4011), .ZN(n4008) );
  XOR2_X1 U4007 ( .A(n4012), .B(n4013), .Z(n3890) );
  NAND2_X1 U4008 ( .A1(n4014), .A2(n4015), .ZN(n4012) );
  XNOR2_X1 U4009 ( .A(n4016), .B(n4017), .ZN(n3894) );
  XOR2_X1 U4010 ( .A(n4018), .B(n4019), .Z(n4016) );
  NOR2_X1 U4011 ( .A1(n3349), .A2(n2411), .ZN(n4019) );
  INV_X1 U4012 ( .A(n3958), .ZN(n3825) );
  XOR2_X1 U4013 ( .A(n4020), .B(n4021), .Z(n3958) );
  NAND2_X1 U4014 ( .A1(n4022), .A2(n4023), .ZN(n4020) );
  XOR2_X1 U4015 ( .A(n4024), .B(n4025), .Z(n3818) );
  XOR2_X1 U4016 ( .A(n4026), .B(n4027), .Z(n4024) );
  NOR2_X1 U4017 ( .A1(n2495), .A2(n2411), .ZN(n4027) );
  XNOR2_X1 U4018 ( .A(n4028), .B(n4029), .ZN(n3901) );
  XOR2_X1 U4019 ( .A(n4030), .B(n4031), .Z(n4028) );
  NOR2_X1 U4020 ( .A1(n2497), .A2(n2411), .ZN(n4031) );
  XOR2_X1 U4021 ( .A(n4032), .B(n4033), .Z(n3905) );
  XOR2_X1 U4022 ( .A(n4034), .B(n2405), .Z(n4032) );
  XOR2_X1 U4023 ( .A(n4035), .B(n4036), .Z(n3909) );
  XNOR2_X1 U4024 ( .A(n4037), .B(n4038), .ZN(n4036) );
  NAND2_X1 U4025 ( .A1(a_2_), .A2(b_3_), .ZN(n4038) );
  XOR2_X1 U4026 ( .A(n4039), .B(n4040), .Z(n3913) );
  XNOR2_X1 U4027 ( .A(n4041), .B(n4042), .ZN(n4039) );
  NAND2_X1 U4028 ( .A1(b_3_), .A2(a_1_), .ZN(n4041) );
  INV_X1 U4029 ( .A(n4043), .ZN(n3917) );
  NAND2_X1 U4030 ( .A1(n3920), .A2(n3921), .ZN(n4043) );
  NAND2_X1 U4031 ( .A1(n4044), .A2(n4045), .ZN(n3921) );
  NAND2_X1 U4032 ( .A1(n4046), .A2(a_0_), .ZN(n4045) );
  NOR2_X1 U4033 ( .A1(n4047), .A2(n2411), .ZN(n4046) );
  NOR2_X1 U4034 ( .A1(n3923), .A2(n3924), .ZN(n4047) );
  NAND2_X1 U4035 ( .A1(n3923), .A2(n3924), .ZN(n4044) );
  NAND2_X1 U4036 ( .A1(n4048), .A2(n4049), .ZN(n3924) );
  NAND2_X1 U4037 ( .A1(n4050), .A2(b_3_), .ZN(n4049) );
  NOR2_X1 U4038 ( .A1(n4051), .A2(n2500), .ZN(n4050) );
  NOR2_X1 U4039 ( .A1(n4042), .A2(n4040), .ZN(n4051) );
  NAND2_X1 U4040 ( .A1(n4040), .A2(n4042), .ZN(n4048) );
  NAND2_X1 U4041 ( .A1(n4052), .A2(n4053), .ZN(n4042) );
  NAND2_X1 U4042 ( .A1(n4054), .A2(a_2_), .ZN(n4053) );
  NOR2_X1 U4043 ( .A1(n4055), .A2(n2411), .ZN(n4054) );
  NOR2_X1 U4044 ( .A1(n4037), .A2(n4035), .ZN(n4055) );
  NAND2_X1 U4045 ( .A1(n4037), .A2(n4035), .ZN(n4052) );
  XNOR2_X1 U4046 ( .A(n4056), .B(n4057), .ZN(n4035) );
  XNOR2_X1 U4047 ( .A(n4058), .B(n4059), .ZN(n4056) );
  NOR2_X1 U4048 ( .A1(n4060), .A2(n4061), .ZN(n4037) );
  INV_X1 U4049 ( .A(n4062), .ZN(n4061) );
  NAND2_X1 U4050 ( .A1(n4033), .A2(n4063), .ZN(n4062) );
  NAND2_X1 U4051 ( .A1(n2405), .A2(n4034), .ZN(n4063) );
  XOR2_X1 U4052 ( .A(n4064), .B(n4065), .Z(n4033) );
  XNOR2_X1 U4053 ( .A(n4066), .B(n4067), .ZN(n4064) );
  NOR2_X1 U4054 ( .A1(n4034), .A2(n2405), .ZN(n4060) );
  INV_X1 U4055 ( .A(n2460), .ZN(n2405) );
  NAND2_X1 U4056 ( .A1(a_3_), .A2(b_3_), .ZN(n2460) );
  NAND2_X1 U4057 ( .A1(n4068), .A2(n4069), .ZN(n4034) );
  NAND2_X1 U4058 ( .A1(n4070), .A2(b_3_), .ZN(n4069) );
  NOR2_X1 U4059 ( .A1(n4071), .A2(n2497), .ZN(n4070) );
  NOR2_X1 U4060 ( .A1(n4030), .A2(n4029), .ZN(n4071) );
  NAND2_X1 U4061 ( .A1(n4029), .A2(n4030), .ZN(n4068) );
  NAND2_X1 U4062 ( .A1(n4072), .A2(n4073), .ZN(n4030) );
  NAND2_X1 U4063 ( .A1(n4074), .A2(b_3_), .ZN(n4073) );
  NOR2_X1 U4064 ( .A1(n4075), .A2(n2373), .ZN(n4074) );
  NOR2_X1 U4065 ( .A1(n3948), .A2(n3947), .ZN(n4075) );
  NAND2_X1 U4066 ( .A1(n3947), .A2(n3948), .ZN(n4072) );
  NAND2_X1 U4067 ( .A1(n4076), .A2(n4077), .ZN(n3948) );
  NAND2_X1 U4068 ( .A1(n4078), .A2(b_3_), .ZN(n4077) );
  NOR2_X1 U4069 ( .A1(n4079), .A2(n2495), .ZN(n4078) );
  NOR2_X1 U4070 ( .A1(n4026), .A2(n4025), .ZN(n4079) );
  NAND2_X1 U4071 ( .A1(n4025), .A2(n4026), .ZN(n4076) );
  NAND2_X1 U4072 ( .A1(n4022), .A2(n4080), .ZN(n4026) );
  NAND2_X1 U4073 ( .A1(n4021), .A2(n4023), .ZN(n4080) );
  NAND2_X1 U4074 ( .A1(n4081), .A2(n4082), .ZN(n4023) );
  NAND2_X1 U4075 ( .A1(b_3_), .A2(a_7_), .ZN(n4082) );
  INV_X1 U4076 ( .A(n4083), .ZN(n4081) );
  XNOR2_X1 U4077 ( .A(n4084), .B(n4085), .ZN(n4021) );
  XNOR2_X1 U4078 ( .A(n4086), .B(n4087), .ZN(n4084) );
  NAND2_X1 U4079 ( .A1(a_7_), .A2(n4083), .ZN(n4022) );
  NAND2_X1 U4080 ( .A1(n4088), .A2(n4089), .ZN(n4083) );
  NAND2_X1 U4081 ( .A1(n4090), .A2(b_3_), .ZN(n4089) );
  NOR2_X1 U4082 ( .A1(n4091), .A2(n3349), .ZN(n4090) );
  NOR2_X1 U4083 ( .A1(n4018), .A2(n4017), .ZN(n4091) );
  NAND2_X1 U4084 ( .A1(n4017), .A2(n4018), .ZN(n4088) );
  NAND2_X1 U4085 ( .A1(n4014), .A2(n4092), .ZN(n4018) );
  NAND2_X1 U4086 ( .A1(n4013), .A2(n4015), .ZN(n4092) );
  NAND2_X1 U4087 ( .A1(n4093), .A2(n4094), .ZN(n4015) );
  NAND2_X1 U4088 ( .A1(b_3_), .A2(a_9_), .ZN(n4094) );
  INV_X1 U4089 ( .A(n4095), .ZN(n4093) );
  XOR2_X1 U4090 ( .A(n4096), .B(n4097), .Z(n4013) );
  XOR2_X1 U4091 ( .A(n4098), .B(n4099), .Z(n4097) );
  NAND2_X1 U4092 ( .A1(a_9_), .A2(n4095), .ZN(n4014) );
  NAND2_X1 U4093 ( .A1(n4010), .A2(n4100), .ZN(n4095) );
  NAND2_X1 U4094 ( .A1(n4009), .A2(n4011), .ZN(n4100) );
  NAND2_X1 U4095 ( .A1(n4101), .A2(n4102), .ZN(n4011) );
  NAND2_X1 U4096 ( .A1(b_3_), .A2(a_10_), .ZN(n4102) );
  INV_X1 U4097 ( .A(n4103), .ZN(n4101) );
  XNOR2_X1 U4098 ( .A(n4104), .B(n4105), .ZN(n4009) );
  XNOR2_X1 U4099 ( .A(n4106), .B(n4107), .ZN(n4105) );
  NAND2_X1 U4100 ( .A1(a_10_), .A2(n4103), .ZN(n4010) );
  NAND2_X1 U4101 ( .A1(n3977), .A2(n4108), .ZN(n4103) );
  NAND2_X1 U4102 ( .A1(n3976), .A2(n3978), .ZN(n4108) );
  NAND2_X1 U4103 ( .A1(n4109), .A2(n4110), .ZN(n3978) );
  NAND2_X1 U4104 ( .A1(b_3_), .A2(a_11_), .ZN(n4110) );
  INV_X1 U4105 ( .A(n4111), .ZN(n4109) );
  XOR2_X1 U4106 ( .A(n4112), .B(n4113), .Z(n3976) );
  XNOR2_X1 U4107 ( .A(n4114), .B(n4115), .ZN(n4113) );
  NAND2_X1 U4108 ( .A1(a_11_), .A2(n4111), .ZN(n3977) );
  NAND2_X1 U4109 ( .A1(n4116), .A2(n4117), .ZN(n4111) );
  NAND2_X1 U4110 ( .A1(n4118), .A2(b_3_), .ZN(n4117) );
  NOR2_X1 U4111 ( .A1(n4119), .A2(n2490), .ZN(n4118) );
  NOR2_X1 U4112 ( .A1(n3984), .A2(n3986), .ZN(n4119) );
  NAND2_X1 U4113 ( .A1(n3984), .A2(n3986), .ZN(n4116) );
  NAND2_X1 U4114 ( .A1(n4120), .A2(n4121), .ZN(n3986) );
  NAND2_X1 U4115 ( .A1(n4122), .A2(b_3_), .ZN(n4121) );
  NOR2_X1 U4116 ( .A1(n4123), .A2(n2252), .ZN(n4122) );
  NOR2_X1 U4117 ( .A1(n4124), .A2(n4007), .ZN(n4123) );
  NAND2_X1 U4118 ( .A1(n4124), .A2(n4007), .ZN(n4120) );
  NAND2_X1 U4119 ( .A1(n4125), .A2(n4126), .ZN(n4007) );
  NAND2_X1 U4120 ( .A1(b_1_), .A2(n4127), .ZN(n4126) );
  NAND2_X1 U4121 ( .A1(n2227), .A2(n4128), .ZN(n4127) );
  NAND2_X1 U4122 ( .A1(a_15_), .A2(n2498), .ZN(n4128) );
  NAND2_X1 U4123 ( .A1(b_2_), .A2(n4129), .ZN(n4125) );
  NAND2_X1 U4124 ( .A1(n2231), .A2(n4130), .ZN(n4129) );
  NAND2_X1 U4125 ( .A1(a_14_), .A2(n2499), .ZN(n4130) );
  INV_X1 U4126 ( .A(n4006), .ZN(n4124) );
  NAND2_X1 U4127 ( .A1(n4131), .A2(n2488), .ZN(n4006) );
  NOR2_X1 U4128 ( .A1(n2411), .A2(n2498), .ZN(n4131) );
  XOR2_X1 U4129 ( .A(n4132), .B(n4133), .Z(n3984) );
  XOR2_X1 U4130 ( .A(n4134), .B(n4135), .Z(n4133) );
  NAND2_X1 U4131 ( .A1(b_2_), .A2(a_13_), .ZN(n4132) );
  XNOR2_X1 U4132 ( .A(n4136), .B(n4137), .ZN(n4017) );
  XOR2_X1 U4133 ( .A(n4138), .B(n4139), .Z(n4136) );
  XNOR2_X1 U4134 ( .A(n4140), .B(n4141), .ZN(n4025) );
  XNOR2_X1 U4135 ( .A(n4142), .B(n4143), .ZN(n4140) );
  XNOR2_X1 U4136 ( .A(n4144), .B(n4145), .ZN(n3947) );
  XNOR2_X1 U4137 ( .A(n4146), .B(n4147), .ZN(n4144) );
  XNOR2_X1 U4138 ( .A(n4148), .B(n4149), .ZN(n4029) );
  XNOR2_X1 U4139 ( .A(n4150), .B(n4151), .ZN(n4148) );
  XNOR2_X1 U4140 ( .A(n4152), .B(n4153), .ZN(n4040) );
  XOR2_X1 U4141 ( .A(n4154), .B(n2431), .Z(n4152) );
  XNOR2_X1 U4142 ( .A(n4155), .B(n4156), .ZN(n3923) );
  XNOR2_X1 U4143 ( .A(n4157), .B(n4158), .ZN(n4156) );
  XNOR2_X1 U4144 ( .A(n4159), .B(n4160), .ZN(n3920) );
  XOR2_X1 U4145 ( .A(n4161), .B(n4162), .Z(n4159) );
  NOR2_X1 U4146 ( .A1(n2498), .A2(n3191), .ZN(n4162) );
  NAND2_X1 U4147 ( .A1(n2537), .A2(n2536), .ZN(n2397) );
  NAND2_X1 U4148 ( .A1(n2534), .A2(b_0_), .ZN(n2536) );
  NAND2_X1 U4149 ( .A1(n4163), .A2(b_1_), .ZN(n2534) );
  NAND2_X1 U4150 ( .A1(n4164), .A2(n4165), .ZN(n2537) );
  INV_X1 U4151 ( .A(n2399), .ZN(n2238) );
  XOR2_X1 U4152 ( .A(n4165), .B(n4164), .Z(n2399) );
  NAND2_X1 U4153 ( .A1(n4166), .A2(n4167), .ZN(n4164) );
  XOR2_X1 U4154 ( .A(n4168), .B(n4163), .Z(n4167) );
  NOR2_X1 U4155 ( .A1(n2500), .A2(n4169), .ZN(n4163) );
  NAND2_X1 U4156 ( .A1(a_0_), .A2(b_1_), .ZN(n4168) );
  NOR2_X1 U4157 ( .A1(n4170), .A2(n4171), .ZN(n4166) );
  NOR2_X1 U4158 ( .A1(n2444), .A2(n4172), .ZN(n4170) );
  NAND2_X1 U4159 ( .A1(n4161), .A2(n4173), .ZN(n4165) );
  NAND2_X1 U4160 ( .A1(n4160), .A2(b_2_), .ZN(n4173) );
  XNOR2_X1 U4161 ( .A(n4172), .B(n4174), .ZN(n4160) );
  NOR2_X1 U4162 ( .A1(n2444), .A2(n4171), .ZN(n4174) );
  NAND2_X1 U4163 ( .A1(n4175), .A2(n4176), .ZN(n4171) );
  NAND2_X1 U4164 ( .A1(n4177), .A2(b_1_), .ZN(n4176) );
  NOR2_X1 U4165 ( .A1(n4178), .A2(n2426), .ZN(n4177) );
  NOR2_X1 U4166 ( .A1(n4179), .A2(n4180), .ZN(n4178) );
  NAND2_X1 U4167 ( .A1(n4179), .A2(n4180), .ZN(n4175) );
  NAND2_X1 U4168 ( .A1(b_1_), .A2(a_1_), .ZN(n2444) );
  NAND2_X1 U4169 ( .A1(a_2_), .A2(b_0_), .ZN(n4172) );
  NOR2_X1 U4170 ( .A1(n4181), .A2(n4182), .ZN(n4161) );
  INV_X1 U4171 ( .A(n4183), .ZN(n4182) );
  NAND2_X1 U4172 ( .A1(n4158), .A2(n4184), .ZN(n4183) );
  NAND2_X1 U4173 ( .A1(n4155), .A2(n4157), .ZN(n4184) );
  NOR2_X1 U4174 ( .A1(n2498), .A2(n2500), .ZN(n4158) );
  INV_X1 U4175 ( .A(a_1_), .ZN(n2500) );
  NOR2_X1 U4176 ( .A1(n4155), .A2(n4157), .ZN(n4181) );
  NAND2_X1 U4177 ( .A1(n4185), .A2(n4186), .ZN(n4157) );
  NAND2_X1 U4178 ( .A1(n4153), .A2(n4187), .ZN(n4186) );
  INV_X1 U4179 ( .A(n4188), .ZN(n4187) );
  NOR2_X1 U4180 ( .A1(n2431), .A2(n4154), .ZN(n4188) );
  XNOR2_X1 U4181 ( .A(n4189), .B(n4190), .ZN(n4153) );
  XNOR2_X1 U4182 ( .A(n4191), .B(n4192), .ZN(n4190) );
  NAND2_X1 U4183 ( .A1(b_1_), .A2(a_3_), .ZN(n4189) );
  NAND2_X1 U4184 ( .A1(n4154), .A2(n2431), .ZN(n4185) );
  NAND2_X1 U4185 ( .A1(b_2_), .A2(a_2_), .ZN(n2431) );
  NOR2_X1 U4186 ( .A1(n4193), .A2(n4194), .ZN(n4154) );
  INV_X1 U4187 ( .A(n4195), .ZN(n4194) );
  NAND2_X1 U4188 ( .A1(n4058), .A2(n4196), .ZN(n4195) );
  NAND2_X1 U4189 ( .A1(n4059), .A2(n4057), .ZN(n4196) );
  NOR2_X1 U4190 ( .A1(n2498), .A2(n2410), .ZN(n4058) );
  NOR2_X1 U4191 ( .A1(n4057), .A2(n4059), .ZN(n4193) );
  NOR2_X1 U4192 ( .A1(n4197), .A2(n4198), .ZN(n4059) );
  INV_X1 U4193 ( .A(n4199), .ZN(n4198) );
  NAND2_X1 U4194 ( .A1(n4067), .A2(n4200), .ZN(n4199) );
  NAND2_X1 U4195 ( .A1(n4066), .A2(n4065), .ZN(n4200) );
  NOR2_X1 U4196 ( .A1(n2498), .A2(n2497), .ZN(n4067) );
  NOR2_X1 U4197 ( .A1(n4065), .A2(n4066), .ZN(n4197) );
  NOR2_X1 U4198 ( .A1(n4201), .A2(n4202), .ZN(n4066) );
  INV_X1 U4199 ( .A(n4203), .ZN(n4202) );
  NAND2_X1 U4200 ( .A1(n4150), .A2(n4204), .ZN(n4203) );
  NAND2_X1 U4201 ( .A1(n4151), .A2(n4149), .ZN(n4204) );
  NOR2_X1 U4202 ( .A1(n2498), .A2(n2373), .ZN(n4150) );
  NOR2_X1 U4203 ( .A1(n4149), .A2(n4151), .ZN(n4201) );
  NOR2_X1 U4204 ( .A1(n4205), .A2(n4206), .ZN(n4151) );
  INV_X1 U4205 ( .A(n4207), .ZN(n4206) );
  NAND2_X1 U4206 ( .A1(n4147), .A2(n4208), .ZN(n4207) );
  NAND2_X1 U4207 ( .A1(n4146), .A2(n4145), .ZN(n4208) );
  NOR2_X1 U4208 ( .A1(n2498), .A2(n2495), .ZN(n4147) );
  NOR2_X1 U4209 ( .A1(n4145), .A2(n4146), .ZN(n4205) );
  NOR2_X1 U4210 ( .A1(n4209), .A2(n4210), .ZN(n4146) );
  INV_X1 U4211 ( .A(n4211), .ZN(n4210) );
  NAND2_X1 U4212 ( .A1(n4142), .A2(n4212), .ZN(n4211) );
  NAND2_X1 U4213 ( .A1(n4143), .A2(n4141), .ZN(n4212) );
  NOR2_X1 U4214 ( .A1(n2498), .A2(n2342), .ZN(n4142) );
  NOR2_X1 U4215 ( .A1(n4141), .A2(n4143), .ZN(n4209) );
  NOR2_X1 U4216 ( .A1(n4213), .A2(n4214), .ZN(n4143) );
  INV_X1 U4217 ( .A(n4215), .ZN(n4214) );
  NAND2_X1 U4218 ( .A1(n4087), .A2(n4216), .ZN(n4215) );
  NAND2_X1 U4219 ( .A1(n4086), .A2(n4085), .ZN(n4216) );
  NOR2_X1 U4220 ( .A1(n2498), .A2(n3349), .ZN(n4087) );
  NOR2_X1 U4221 ( .A1(n4085), .A2(n4086), .ZN(n4213) );
  NOR2_X1 U4222 ( .A1(n4217), .A2(n4218), .ZN(n4086) );
  INV_X1 U4223 ( .A(n4219), .ZN(n4218) );
  NAND2_X1 U4224 ( .A1(n4138), .A2(n4220), .ZN(n4219) );
  NAND2_X1 U4225 ( .A1(n4221), .A2(n4137), .ZN(n4220) );
  NOR2_X1 U4226 ( .A1(n2498), .A2(n2311), .ZN(n4138) );
  NOR2_X1 U4227 ( .A1(n4137), .A2(n4221), .ZN(n4217) );
  INV_X1 U4228 ( .A(n4139), .ZN(n4221) );
  NAND2_X1 U4229 ( .A1(n4222), .A2(n4223), .ZN(n4139) );
  NAND2_X1 U4230 ( .A1(n4099), .A2(n4224), .ZN(n4223) );
  NAND2_X1 U4231 ( .A1(n4098), .A2(n4096), .ZN(n4224) );
  INV_X1 U4232 ( .A(n4225), .ZN(n4096) );
  INV_X1 U4233 ( .A(n4226), .ZN(n4098) );
  NOR2_X1 U4234 ( .A1(n2498), .A2(n2492), .ZN(n4099) );
  NAND2_X1 U4235 ( .A1(n4225), .A2(n4226), .ZN(n4222) );
  NAND2_X1 U4236 ( .A1(n4227), .A2(n4228), .ZN(n4226) );
  NAND2_X1 U4237 ( .A1(n4107), .A2(n4229), .ZN(n4228) );
  NAND2_X1 U4238 ( .A1(n4104), .A2(n4106), .ZN(n4229) );
  NOR2_X1 U4239 ( .A1(n2498), .A2(n2280), .ZN(n4107) );
  INV_X1 U4240 ( .A(n4230), .ZN(n4227) );
  NOR2_X1 U4241 ( .A1(n4104), .A2(n4106), .ZN(n4230) );
  NAND2_X1 U4242 ( .A1(n4231), .A2(n4232), .ZN(n4106) );
  NAND2_X1 U4243 ( .A1(n4112), .A2(n4233), .ZN(n4232) );
  NAND2_X1 U4244 ( .A1(n4115), .A2(n4114), .ZN(n4233) );
  XOR2_X1 U4245 ( .A(n4234), .B(n4235), .Z(n4112) );
  XOR2_X1 U4246 ( .A(n4236), .B(n4237), .Z(n4234) );
  INV_X1 U4247 ( .A(n4238), .ZN(n4231) );
  NOR2_X1 U4248 ( .A1(n4114), .A2(n4115), .ZN(n4238) );
  NOR2_X1 U4249 ( .A1(n2498), .A2(n2490), .ZN(n4115) );
  NAND2_X1 U4250 ( .A1(n4239), .A2(n4240), .ZN(n4114) );
  NAND2_X1 U4251 ( .A1(n4241), .A2(b_2_), .ZN(n4240) );
  NOR2_X1 U4252 ( .A1(n4242), .A2(n2252), .ZN(n4241) );
  NOR2_X1 U4253 ( .A1(n4243), .A2(n4135), .ZN(n4242) );
  NAND2_X1 U4254 ( .A1(n4243), .A2(n4135), .ZN(n4239) );
  NAND2_X1 U4255 ( .A1(n4244), .A2(n4245), .ZN(n4135) );
  NAND2_X1 U4256 ( .A1(b_0_), .A2(n4246), .ZN(n4245) );
  NAND2_X1 U4257 ( .A1(n2227), .A2(n4247), .ZN(n4246) );
  NAND2_X1 U4258 ( .A1(a_15_), .A2(n2499), .ZN(n4247) );
  NAND2_X1 U4259 ( .A1(a_15_), .A2(n2487), .ZN(n2227) );
  NAND2_X1 U4260 ( .A1(b_1_), .A2(n4248), .ZN(n4244) );
  NAND2_X1 U4261 ( .A1(n2231), .A2(n4249), .ZN(n4248) );
  NAND2_X1 U4262 ( .A1(a_14_), .A2(n4169), .ZN(n4249) );
  NAND2_X1 U4263 ( .A1(a_14_), .A2(n4250), .ZN(n2231) );
  INV_X1 U4264 ( .A(n4134), .ZN(n4243) );
  NAND2_X1 U4265 ( .A1(n4251), .A2(n2488), .ZN(n4134) );
  NOR2_X1 U4266 ( .A1(n2499), .A2(n2498), .ZN(n4251) );
  XOR2_X1 U4267 ( .A(n4252), .B(n4253), .Z(n4104) );
  NAND2_X1 U4268 ( .A1(n4254), .A2(n4255), .ZN(n4252) );
  NAND2_X1 U4269 ( .A1(n4256), .A2(n4257), .ZN(n4255) );
  NAND2_X1 U4270 ( .A1(b_1_), .A2(a_12_), .ZN(n4256) );
  XOR2_X1 U4271 ( .A(n4258), .B(n4259), .Z(n4225) );
  XNOR2_X1 U4272 ( .A(n4260), .B(n4261), .ZN(n4259) );
  NAND2_X1 U4273 ( .A1(b_1_), .A2(a_11_), .ZN(n4258) );
  XNOR2_X1 U4274 ( .A(n4262), .B(n4263), .ZN(n4137) );
  XNOR2_X1 U4275 ( .A(n4264), .B(n4265), .ZN(n4263) );
  NAND2_X1 U4276 ( .A1(b_1_), .A2(a_10_), .ZN(n4262) );
  XNOR2_X1 U4277 ( .A(n4266), .B(n4267), .ZN(n4085) );
  XNOR2_X1 U4278 ( .A(n4268), .B(n4269), .ZN(n4267) );
  NAND2_X1 U4279 ( .A1(b_1_), .A2(a_9_), .ZN(n4266) );
  XNOR2_X1 U4280 ( .A(n4270), .B(n4271), .ZN(n4141) );
  XNOR2_X1 U4281 ( .A(n4272), .B(n4273), .ZN(n4271) );
  NAND2_X1 U4282 ( .A1(b_1_), .A2(a_8_), .ZN(n4270) );
  XNOR2_X1 U4283 ( .A(n4274), .B(n4275), .ZN(n4145) );
  XNOR2_X1 U4284 ( .A(n4276), .B(n4277), .ZN(n4275) );
  NAND2_X1 U4285 ( .A1(b_1_), .A2(a_7_), .ZN(n4274) );
  XNOR2_X1 U4286 ( .A(n4278), .B(n4279), .ZN(n4149) );
  XNOR2_X1 U4287 ( .A(n4280), .B(n4281), .ZN(n4279) );
  NAND2_X1 U4288 ( .A1(b_1_), .A2(a_6_), .ZN(n4278) );
  XNOR2_X1 U4289 ( .A(n4282), .B(n4283), .ZN(n4065) );
  XNOR2_X1 U4290 ( .A(n4284), .B(n4285), .ZN(n4283) );
  NAND2_X1 U4291 ( .A1(b_1_), .A2(a_5_), .ZN(n4282) );
  XNOR2_X1 U4292 ( .A(n4286), .B(n4287), .ZN(n4057) );
  XNOR2_X1 U4293 ( .A(n4288), .B(n4289), .ZN(n4287) );
  NAND2_X1 U4294 ( .A1(b_1_), .A2(a_4_), .ZN(n4286) );
  XNOR2_X1 U4295 ( .A(n4290), .B(n4291), .ZN(n4155) );
  XNOR2_X1 U4296 ( .A(n4179), .B(n4180), .ZN(n4291) );
  NAND2_X1 U4297 ( .A1(n4292), .A2(n4293), .ZN(n4180) );
  NAND2_X1 U4298 ( .A1(n4294), .A2(b_1_), .ZN(n4293) );
  NOR2_X1 U4299 ( .A1(n4295), .A2(n2410), .ZN(n4294) );
  NOR2_X1 U4300 ( .A1(n4191), .A2(n4192), .ZN(n4295) );
  NAND2_X1 U4301 ( .A1(n4191), .A2(n4192), .ZN(n4292) );
  NAND2_X1 U4302 ( .A1(n4296), .A2(n4297), .ZN(n4192) );
  NAND2_X1 U4303 ( .A1(n4298), .A2(b_1_), .ZN(n4297) );
  NOR2_X1 U4304 ( .A1(n4299), .A2(n2497), .ZN(n4298) );
  NOR2_X1 U4305 ( .A1(n4288), .A2(n4289), .ZN(n4299) );
  NAND2_X1 U4306 ( .A1(n4288), .A2(n4289), .ZN(n4296) );
  NAND2_X1 U4307 ( .A1(n4300), .A2(n4301), .ZN(n4289) );
  NAND2_X1 U4308 ( .A1(n4302), .A2(b_1_), .ZN(n4301) );
  NOR2_X1 U4309 ( .A1(n4303), .A2(n2373), .ZN(n4302) );
  NOR2_X1 U4310 ( .A1(n4284), .A2(n4285), .ZN(n4303) );
  NAND2_X1 U4311 ( .A1(n4284), .A2(n4285), .ZN(n4300) );
  NAND2_X1 U4312 ( .A1(n4304), .A2(n4305), .ZN(n4285) );
  NAND2_X1 U4313 ( .A1(n4306), .A2(b_1_), .ZN(n4305) );
  NOR2_X1 U4314 ( .A1(n4307), .A2(n2495), .ZN(n4306) );
  NOR2_X1 U4315 ( .A1(n4280), .A2(n4281), .ZN(n4307) );
  NAND2_X1 U4316 ( .A1(n4280), .A2(n4281), .ZN(n4304) );
  NAND2_X1 U4317 ( .A1(n4308), .A2(n4309), .ZN(n4281) );
  NAND2_X1 U4318 ( .A1(n4310), .A2(b_1_), .ZN(n4309) );
  NOR2_X1 U4319 ( .A1(n4311), .A2(n2342), .ZN(n4310) );
  NOR2_X1 U4320 ( .A1(n4276), .A2(n4277), .ZN(n4311) );
  NAND2_X1 U4321 ( .A1(n4276), .A2(n4277), .ZN(n4308) );
  NAND2_X1 U4322 ( .A1(n4312), .A2(n4313), .ZN(n4277) );
  NAND2_X1 U4323 ( .A1(n4314), .A2(b_1_), .ZN(n4313) );
  NOR2_X1 U4324 ( .A1(n4315), .A2(n3349), .ZN(n4314) );
  NOR2_X1 U4325 ( .A1(n4272), .A2(n4273), .ZN(n4315) );
  NAND2_X1 U4326 ( .A1(n4272), .A2(n4273), .ZN(n4312) );
  NAND2_X1 U4327 ( .A1(n4316), .A2(n4317), .ZN(n4273) );
  NAND2_X1 U4328 ( .A1(n4318), .A2(b_1_), .ZN(n4317) );
  NOR2_X1 U4329 ( .A1(n4319), .A2(n2311), .ZN(n4318) );
  NOR2_X1 U4330 ( .A1(n4268), .A2(n4269), .ZN(n4319) );
  NAND2_X1 U4331 ( .A1(n4268), .A2(n4269), .ZN(n4316) );
  NAND2_X1 U4332 ( .A1(n4320), .A2(n4321), .ZN(n4269) );
  NAND2_X1 U4333 ( .A1(n4322), .A2(b_1_), .ZN(n4321) );
  NOR2_X1 U4334 ( .A1(n4323), .A2(n2492), .ZN(n4322) );
  NOR2_X1 U4335 ( .A1(n4264), .A2(n4265), .ZN(n4323) );
  NAND2_X1 U4336 ( .A1(n4264), .A2(n4265), .ZN(n4320) );
  NAND2_X1 U4337 ( .A1(n4324), .A2(n4325), .ZN(n4265) );
  NAND2_X1 U4338 ( .A1(n4326), .A2(b_1_), .ZN(n4325) );
  NOR2_X1 U4339 ( .A1(n4327), .A2(n2280), .ZN(n4326) );
  NOR2_X1 U4340 ( .A1(n4260), .A2(n4261), .ZN(n4327) );
  NAND2_X1 U4341 ( .A1(n4260), .A2(n4261), .ZN(n4324) );
  NAND2_X1 U4342 ( .A1(n4254), .A2(n4328), .ZN(n4261) );
  NAND2_X1 U4343 ( .A1(n4329), .A2(n4253), .ZN(n4328) );
  NAND2_X1 U4344 ( .A1(n4237), .A2(n4330), .ZN(n4253) );
  NAND2_X1 U4345 ( .A1(n4235), .A2(n4236), .ZN(n4330) );
  NOR2_X1 U4346 ( .A1(n2499), .A2(n2252), .ZN(n4236) );
  NOR2_X1 U4347 ( .A1(n4169), .A2(n2487), .ZN(n4235) );
  NAND2_X1 U4348 ( .A1(n4331), .A2(n2488), .ZN(n4237) );
  NOR2_X1 U4349 ( .A1(n4169), .A2(n2499), .ZN(n4331) );
  NAND2_X1 U4350 ( .A1(n4257), .A2(n2490), .ZN(n4329) );
  NAND2_X1 U4351 ( .A1(n4332), .A2(n4333), .ZN(n4254) );
  INV_X1 U4352 ( .A(n4257), .ZN(n4333) );
  NAND2_X1 U4353 ( .A1(a_13_), .A2(b_0_), .ZN(n4257) );
  NOR2_X1 U4354 ( .A1(n2490), .A2(n2499), .ZN(n4332) );
  NOR2_X1 U4355 ( .A1(n2490), .A2(n4169), .ZN(n4260) );
  NOR2_X1 U4356 ( .A1(n2280), .A2(n4169), .ZN(n4264) );
  NOR2_X1 U4357 ( .A1(n2492), .A2(n4169), .ZN(n4268) );
  INV_X1 U4358 ( .A(a_10_), .ZN(n2492) );
  NOR2_X1 U4359 ( .A1(n2311), .A2(n4169), .ZN(n4272) );
  NOR2_X1 U4360 ( .A1(n3349), .A2(n4169), .ZN(n4276) );
  NOR2_X1 U4361 ( .A1(n2342), .A2(n4169), .ZN(n4280) );
  NOR2_X1 U4362 ( .A1(n2495), .A2(n4169), .ZN(n4284) );
  NOR2_X1 U4363 ( .A1(n2373), .A2(n4169), .ZN(n4288) );
  NOR2_X1 U4364 ( .A1(n2497), .A2(n4169), .ZN(n4191) );
  NOR2_X1 U4365 ( .A1(n2410), .A2(n4169), .ZN(n4179) );
  NAND2_X1 U4366 ( .A1(b_1_), .A2(a_2_), .ZN(n4290) );
  NAND2_X1 U4367 ( .A1(n4334), .A2(n4335), .ZN(n2223) );
  NAND2_X1 U4368 ( .A1(n4336), .A2(n2457), .ZN(n4335) );
  NAND2_X1 U4369 ( .A1(b_0_), .A2(n3191), .ZN(n2457) );
  INV_X1 U4370 ( .A(a_0_), .ZN(n3191) );
  NAND2_X1 U4371 ( .A1(n4337), .A2(n4338), .ZN(n4336) );
  NAND2_X1 U4372 ( .A1(a_1_), .A2(n2499), .ZN(n4338) );
  NAND2_X1 U4373 ( .A1(n4339), .A2(n4340), .ZN(n4337) );
  NAND2_X1 U4374 ( .A1(b_2_), .A2(n2426), .ZN(n4340) );
  INV_X1 U4375 ( .A(a_2_), .ZN(n2426) );
  NOR2_X1 U4376 ( .A1(n4341), .A2(n4342), .ZN(n4339) );
  NOR2_X1 U4377 ( .A1(a_1_), .A2(n2499), .ZN(n4342) );
  INV_X1 U4378 ( .A(b_1_), .ZN(n2499) );
  NOR2_X1 U4379 ( .A1(n4343), .A2(n4344), .ZN(n4341) );
  NAND2_X1 U4380 ( .A1(n4345), .A2(n4346), .ZN(n4344) );
  NAND2_X1 U4381 ( .A1(n4347), .A2(n4348), .ZN(n4346) );
  NAND2_X1 U4382 ( .A1(b_4_), .A2(n2497), .ZN(n4348) );
  INV_X1 U4383 ( .A(a_4_), .ZN(n2497) );
  NOR2_X1 U4384 ( .A1(n4349), .A2(n4350), .ZN(n4347) );
  NOR2_X1 U4385 ( .A1(a_3_), .A2(n2411), .ZN(n4350) );
  INV_X1 U4386 ( .A(b_3_), .ZN(n2411) );
  NOR2_X1 U4387 ( .A1(n4351), .A2(n4352), .ZN(n4349) );
  NAND2_X1 U4388 ( .A1(n4353), .A2(n4354), .ZN(n4352) );
  NAND2_X1 U4389 ( .A1(n4355), .A2(n4356), .ZN(n4354) );
  NAND2_X1 U4390 ( .A1(b_6_), .A2(n2495), .ZN(n4356) );
  INV_X1 U4391 ( .A(a_6_), .ZN(n2495) );
  NOR2_X1 U4392 ( .A1(n4357), .A2(n4358), .ZN(n4355) );
  NOR2_X1 U4393 ( .A1(a_5_), .A2(n2374), .ZN(n4358) );
  INV_X1 U4394 ( .A(b_5_), .ZN(n2374) );
  NOR2_X1 U4395 ( .A1(n4359), .A2(n4360), .ZN(n4357) );
  NAND2_X1 U4396 ( .A1(n4361), .A2(n4362), .ZN(n4360) );
  NAND2_X1 U4397 ( .A1(n4363), .A2(n4364), .ZN(n4362) );
  NAND2_X1 U4398 ( .A1(b_8_), .A2(n3349), .ZN(n4364) );
  INV_X1 U4399 ( .A(a_8_), .ZN(n3349) );
  NOR2_X1 U4400 ( .A1(n4365), .A2(n4366), .ZN(n4363) );
  NOR2_X1 U4401 ( .A1(a_7_), .A2(n2343), .ZN(n4366) );
  INV_X1 U4402 ( .A(b_7_), .ZN(n2343) );
  NOR2_X1 U4403 ( .A1(n4367), .A2(n4368), .ZN(n4365) );
  NAND2_X1 U4404 ( .A1(n4369), .A2(n4370), .ZN(n4368) );
  NAND2_X1 U4405 ( .A1(n4371), .A2(n4372), .ZN(n4370) );
  NAND2_X1 U4406 ( .A1(b_9_), .A2(n2311), .ZN(n4372) );
  NOR2_X1 U4407 ( .A1(n4373), .A2(n4374), .ZN(n4371) );
  NOR2_X1 U4408 ( .A1(a_10_), .A2(n2491), .ZN(n4374) );
  NOR2_X1 U4409 ( .A1(n4375), .A2(n4376), .ZN(n4373) );
  NAND2_X1 U4410 ( .A1(n4377), .A2(n4378), .ZN(n4376) );
  NAND2_X1 U4411 ( .A1(n4379), .A2(n4380), .ZN(n4378) );
  NAND2_X1 U4412 ( .A1(b_12_), .A2(n2490), .ZN(n4380) );
  INV_X1 U4413 ( .A(a_12_), .ZN(n2490) );
  NOR2_X1 U4414 ( .A1(n4381), .A2(n4382), .ZN(n4379) );
  NOR2_X1 U4415 ( .A1(a_11_), .A2(n2281), .ZN(n4382) );
  INV_X1 U4416 ( .A(b_11_), .ZN(n2281) );
  NOR2_X1 U4417 ( .A1(n4383), .A2(n4384), .ZN(n4381) );
  NAND2_X1 U4418 ( .A1(n4385), .A2(n4386), .ZN(n4384) );
  NAND2_X1 U4419 ( .A1(n4387), .A2(n4388), .ZN(n4386) );
  NOR2_X1 U4420 ( .A1(n4389), .A2(n4390), .ZN(n4388) );
  NOR2_X1 U4421 ( .A1(n2488), .A2(n2233), .ZN(n4390) );
  INV_X1 U4422 ( .A(b_14_), .ZN(n2233) );
  INV_X1 U4423 ( .A(a_15_), .ZN(n4250) );
  NOR2_X1 U4424 ( .A1(n4391), .A2(n2229), .ZN(n4389) );
  INV_X1 U4425 ( .A(b_15_), .ZN(n2229) );
  NOR2_X1 U4426 ( .A1(b_14_), .A2(n2487), .ZN(n4391) );
  INV_X1 U4427 ( .A(a_14_), .ZN(n2487) );
  NOR2_X1 U4428 ( .A1(n4392), .A2(n4393), .ZN(n4387) );
  NOR2_X1 U4429 ( .A1(a_15_), .A2(a_14_), .ZN(n4393) );
  NOR2_X1 U4430 ( .A1(a_13_), .A2(n2250), .ZN(n4392) );
  INV_X1 U4431 ( .A(b_13_), .ZN(n2250) );
  NAND2_X1 U4432 ( .A1(a_12_), .A2(n2489), .ZN(n4385) );
  INV_X1 U4433 ( .A(b_12_), .ZN(n2489) );
  NOR2_X1 U4434 ( .A1(b_13_), .A2(n2252), .ZN(n4383) );
  INV_X1 U4435 ( .A(a_13_), .ZN(n2252) );
  NAND2_X1 U4436 ( .A1(a_10_), .A2(n2491), .ZN(n4377) );
  INV_X1 U4437 ( .A(b_10_), .ZN(n2491) );
  NOR2_X1 U4438 ( .A1(b_11_), .A2(n2280), .ZN(n4375) );
  INV_X1 U4439 ( .A(a_11_), .ZN(n2280) );
  NAND2_X1 U4440 ( .A1(a_8_), .A2(n3283), .ZN(n4369) );
  INV_X1 U4441 ( .A(b_8_), .ZN(n3283) );
  NOR2_X1 U4442 ( .A1(b_9_), .A2(n2311), .ZN(n4367) );
  INV_X1 U4443 ( .A(a_9_), .ZN(n2311) );
  NAND2_X1 U4444 ( .A1(a_6_), .A2(n2494), .ZN(n4361) );
  INV_X1 U4445 ( .A(b_6_), .ZN(n2494) );
  NOR2_X1 U4446 ( .A1(b_7_), .A2(n2342), .ZN(n4359) );
  INV_X1 U4447 ( .A(a_7_), .ZN(n2342) );
  NAND2_X1 U4448 ( .A1(a_4_), .A2(n2496), .ZN(n4353) );
  INV_X1 U4449 ( .A(b_4_), .ZN(n2496) );
  NOR2_X1 U4450 ( .A1(b_5_), .A2(n2373), .ZN(n4351) );
  INV_X1 U4451 ( .A(a_5_), .ZN(n2373) );
  NAND2_X1 U4452 ( .A1(a_2_), .A2(n2498), .ZN(n4345) );
  INV_X1 U4453 ( .A(b_2_), .ZN(n2498) );
  NOR2_X1 U4454 ( .A1(b_3_), .A2(n2410), .ZN(n4343) );
  INV_X1 U4455 ( .A(a_3_), .ZN(n2410) );
  NAND2_X1 U4456 ( .A1(a_0_), .A2(n4169), .ZN(n4334) );
  INV_X1 U4457 ( .A(b_0_), .ZN(n4169) );
endmodule

