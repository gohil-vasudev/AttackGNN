module add_mul_mix_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, 
        c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_,
         c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817;

  OR2_X1 U939 ( .A1(n924), .A2(n925), .ZN(Result_9_) );
  AND2_X1 U940 ( .A1(n926), .A2(n927), .ZN(n925) );
  INV_X1 U941 ( .A(n928), .ZN(n924) );
  OR2_X1 U942 ( .A1(n927), .A2(n926), .ZN(n928) );
  OR2_X1 U943 ( .A1(n929), .A2(n930), .ZN(n926) );
  AND2_X1 U944 ( .A1(n931), .A2(n932), .ZN(n930) );
  INV_X1 U945 ( .A(n933), .ZN(n931) );
  AND2_X1 U946 ( .A1(n934), .A2(n933), .ZN(n929) );
  INV_X1 U947 ( .A(n932), .ZN(n934) );
  OR2_X1 U948 ( .A1(n935), .A2(n936), .ZN(Result_8_) );
  AND2_X1 U949 ( .A1(n937), .A2(n938), .ZN(n936) );
  INV_X1 U950 ( .A(n939), .ZN(n935) );
  OR2_X1 U951 ( .A1(n938), .A2(n937), .ZN(n939) );
  OR2_X1 U952 ( .A1(n940), .A2(n941), .ZN(n937) );
  AND2_X1 U953 ( .A1(n942), .A2(n943), .ZN(n941) );
  INV_X1 U954 ( .A(n944), .ZN(n942) );
  AND2_X1 U955 ( .A1(n945), .A2(n944), .ZN(n940) );
  INV_X1 U956 ( .A(n943), .ZN(n945) );
  OR2_X1 U957 ( .A1(n946), .A2(n947), .ZN(Result_7_) );
  AND2_X1 U958 ( .A1(n948), .A2(n949), .ZN(n947) );
  AND2_X1 U959 ( .A1(n950), .A2(n951), .ZN(n946) );
  AND2_X1 U960 ( .A1(n952), .A2(n953), .ZN(Result_6_) );
  OR2_X1 U961 ( .A1(n954), .A2(n955), .ZN(n952) );
  AND2_X1 U962 ( .A1(n951), .A2(n948), .ZN(n954) );
  INV_X1 U963 ( .A(n950), .ZN(n948) );
  INV_X1 U964 ( .A(n949), .ZN(n951) );
  AND2_X1 U965 ( .A1(n956), .A2(n957), .ZN(Result_5_) );
  INV_X1 U966 ( .A(n958), .ZN(n956) );
  AND2_X1 U967 ( .A1(n959), .A2(n960), .ZN(n958) );
  AND2_X1 U968 ( .A1(n961), .A2(n962), .ZN(Result_4_) );
  INV_X1 U969 ( .A(n963), .ZN(n961) );
  AND2_X1 U970 ( .A1(n964), .A2(n965), .ZN(n963) );
  AND2_X1 U971 ( .A1(n966), .A2(n967), .ZN(Result_3_) );
  INV_X1 U972 ( .A(n968), .ZN(n966) );
  AND2_X1 U973 ( .A1(n969), .A2(n970), .ZN(n968) );
  OR2_X1 U974 ( .A1(n971), .A2(n972), .ZN(Result_2_) );
  AND2_X1 U975 ( .A1(n973), .A2(n974), .ZN(n972) );
  AND2_X1 U976 ( .A1(n975), .A2(n967), .ZN(n971) );
  OR2_X1 U977 ( .A1(n976), .A2(n977), .ZN(n975) );
  AND2_X1 U978 ( .A1(n978), .A2(n979), .ZN(n977) );
  AND2_X1 U979 ( .A1(n980), .A2(n974), .ZN(n976) );
  OR2_X1 U980 ( .A1(n981), .A2(n982), .ZN(Result_1_) );
  INV_X1 U981 ( .A(n983), .ZN(n982) );
  OR2_X1 U982 ( .A1(n984), .A2(n985), .ZN(n983) );
  AND2_X1 U983 ( .A1(n985), .A2(n984), .ZN(n981) );
  OR2_X1 U984 ( .A1(n986), .A2(n987), .ZN(n984) );
  AND2_X1 U985 ( .A1(n988), .A2(n989), .ZN(n987) );
  OR2_X1 U986 ( .A1(n990), .A2(n991), .ZN(n989) );
  OR2_X1 U987 ( .A1(n992), .A2(n993), .ZN(Result_14_) );
  AND2_X1 U988 ( .A1(n994), .A2(n995), .ZN(n993) );
  INV_X1 U989 ( .A(n996), .ZN(n992) );
  OR2_X1 U990 ( .A1(n995), .A2(n994), .ZN(n996) );
  AND2_X1 U991 ( .A1(n997), .A2(n998), .ZN(n994) );
  OR2_X1 U992 ( .A1(n999), .A2(n1000), .ZN(n995) );
  OR2_X1 U993 ( .A1(n1001), .A2(n1002), .ZN(Result_13_) );
  AND2_X1 U994 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
  INV_X1 U995 ( .A(n1005), .ZN(n1001) );
  OR2_X1 U996 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  OR2_X1 U997 ( .A1(n1006), .A2(n1007), .ZN(n1003) );
  INV_X1 U998 ( .A(n1008), .ZN(n1007) );
  OR2_X1 U999 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
  AND2_X1 U1000 ( .A1(n1010), .A2(n1009), .ZN(n1006) );
  OR2_X1 U1001 ( .A1(n1011), .A2(n1012), .ZN(Result_12_) );
  AND2_X1 U1002 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
  INV_X1 U1003 ( .A(n1015), .ZN(n1011) );
  OR2_X1 U1004 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  OR2_X1 U1005 ( .A1(n1016), .A2(n1017), .ZN(n1013) );
  AND2_X1 U1006 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
  INV_X1 U1007 ( .A(n1020), .ZN(n1018) );
  AND2_X1 U1008 ( .A1(n1021), .A2(n1020), .ZN(n1016) );
  INV_X1 U1009 ( .A(n1019), .ZN(n1021) );
  OR2_X1 U1010 ( .A1(n1022), .A2(n1023), .ZN(Result_11_) );
  AND2_X1 U1011 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
  INV_X1 U1012 ( .A(n1026), .ZN(n1022) );
  OR2_X1 U1013 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  OR2_X1 U1014 ( .A1(n1027), .A2(n1028), .ZN(n1024) );
  AND2_X1 U1015 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
  INV_X1 U1016 ( .A(n1031), .ZN(n1029) );
  AND2_X1 U1017 ( .A1(n1032), .A2(n1031), .ZN(n1027) );
  INV_X1 U1018 ( .A(n1030), .ZN(n1032) );
  OR2_X1 U1019 ( .A1(n1033), .A2(n1034), .ZN(Result_10_) );
  AND2_X1 U1020 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
  INV_X1 U1021 ( .A(n1037), .ZN(n1033) );
  OR2_X1 U1022 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  OR2_X1 U1023 ( .A1(n1038), .A2(n1039), .ZN(n1035) );
  AND2_X1 U1024 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
  INV_X1 U1025 ( .A(n1042), .ZN(n1040) );
  AND2_X1 U1026 ( .A1(n1043), .A2(n1042), .ZN(n1038) );
  INV_X1 U1027 ( .A(n1041), .ZN(n1043) );
  OR3_X1 U1028 ( .A1(n986), .A2(n1044), .A3(n1045), .ZN(Result_0_) );
  AND2_X1 U1029 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
  AND2_X1 U1030 ( .A1(n985), .A2(n1048), .ZN(n1044) );
  AND2_X1 U1031 ( .A1(n1049), .A2(n978), .ZN(n985) );
  INV_X1 U1032 ( .A(n974), .ZN(n978) );
  AND2_X1 U1033 ( .A1(n1050), .A2(n1051), .ZN(n974) );
  OR2_X1 U1034 ( .A1(n990), .A2(n1052), .ZN(n1051) );
  INV_X1 U1035 ( .A(n1053), .ZN(n990) );
  OR2_X1 U1036 ( .A1(n1053), .A2(n991), .ZN(n1050) );
  OR2_X1 U1037 ( .A1(n980), .A2(n973), .ZN(n1049) );
  INV_X1 U1038 ( .A(n967), .ZN(n973) );
  OR2_X1 U1039 ( .A1(n970), .A2(n969), .ZN(n967) );
  OR2_X1 U1040 ( .A1(n1054), .A2(n980), .ZN(n969) );
  AND2_X1 U1041 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
  AND2_X1 U1042 ( .A1(n962), .A2(n1057), .ZN(n970) );
  OR2_X1 U1043 ( .A1(n965), .A2(n964), .ZN(n962) );
  OR2_X1 U1044 ( .A1(n1058), .A2(n1059), .ZN(n964) );
  INV_X1 U1045 ( .A(n1057), .ZN(n1059) );
  OR2_X1 U1046 ( .A1(n1060), .A2(n1061), .ZN(n1057) );
  AND2_X1 U1047 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
  OR2_X1 U1048 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
  AND2_X1 U1049 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
  AND2_X1 U1050 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
  OR2_X1 U1051 ( .A1(n1065), .A2(n1064), .ZN(n1067) );
  AND2_X1 U1052 ( .A1(n1068), .A2(n1069), .ZN(n1060) );
  INV_X1 U1053 ( .A(n1070), .ZN(n1069) );
  AND2_X1 U1054 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
  OR2_X1 U1055 ( .A1(n1072), .A2(n1071), .ZN(n1068) );
  OR2_X1 U1056 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
  INV_X1 U1057 ( .A(n1075), .ZN(n1074) );
  OR2_X1 U1058 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
  AND2_X1 U1059 ( .A1(n1077), .A2(n1076), .ZN(n1073) );
  INV_X1 U1060 ( .A(n1078), .ZN(n1077) );
  AND2_X1 U1061 ( .A1(n957), .A2(n1079), .ZN(n965) );
  OR2_X1 U1062 ( .A1(n960), .A2(n959), .ZN(n957) );
  OR2_X1 U1063 ( .A1(n1080), .A2(n1081), .ZN(n959) );
  INV_X1 U1064 ( .A(n1079), .ZN(n1081) );
  OR2_X1 U1065 ( .A1(n1082), .A2(n1083), .ZN(n1079) );
  AND2_X1 U1066 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
  OR2_X1 U1067 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
  AND2_X1 U1068 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
  AND2_X1 U1069 ( .A1(n1088), .A2(n1089), .ZN(n1084) );
  OR2_X1 U1070 ( .A1(n1087), .A2(n1086), .ZN(n1088) );
  AND2_X1 U1071 ( .A1(n1090), .A2(n1091), .ZN(n1082) );
  INV_X1 U1072 ( .A(n1092), .ZN(n1091) );
  AND2_X1 U1073 ( .A1(n1093), .A2(n1066), .ZN(n1092) );
  OR2_X1 U1074 ( .A1(n1066), .A2(n1093), .ZN(n1090) );
  OR2_X1 U1075 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
  INV_X1 U1076 ( .A(n1096), .ZN(n1095) );
  OR2_X1 U1077 ( .A1(n1064), .A2(n1097), .ZN(n1096) );
  AND2_X1 U1078 ( .A1(n1097), .A2(n1064), .ZN(n1094) );
  OR2_X1 U1079 ( .A1(n1098), .A2(n1099), .ZN(n1064) );
  INV_X1 U1080 ( .A(n1065), .ZN(n1097) );
  OR2_X1 U1081 ( .A1(n1100), .A2(n1101), .ZN(n1065) );
  AND2_X1 U1082 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
  AND2_X1 U1083 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
  OR2_X1 U1084 ( .A1(n1103), .A2(n1102), .ZN(n1104) );
  AND2_X1 U1085 ( .A1(n1106), .A2(n1107), .ZN(n1066) );
  INV_X1 U1086 ( .A(n1108), .ZN(n1107) );
  AND2_X1 U1087 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
  OR2_X1 U1088 ( .A1(n1110), .A2(n1109), .ZN(n1106) );
  OR2_X1 U1089 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
  INV_X1 U1090 ( .A(n1113), .ZN(n1112) );
  OR2_X1 U1091 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
  AND2_X1 U1092 ( .A1(n1115), .A2(n1114), .ZN(n1111) );
  INV_X1 U1093 ( .A(n1116), .ZN(n1115) );
  AND2_X1 U1094 ( .A1(n1117), .A2(n953), .ZN(n960) );
  OR3_X1 U1095 ( .A1(n950), .A2(n949), .A3(n1118), .ZN(n953) );
  INV_X1 U1096 ( .A(n955), .ZN(n1118) );
  AND2_X1 U1097 ( .A1(n1117), .A2(n1119), .ZN(n955) );
  INV_X1 U1098 ( .A(n1120), .ZN(n1119) );
  AND2_X1 U1099 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
  OR2_X1 U1100 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
  OR2_X1 U1101 ( .A1(n1125), .A2(n1126), .ZN(n949) );
  AND2_X1 U1102 ( .A1(n944), .A2(n943), .ZN(n1126) );
  AND2_X1 U1103 ( .A1(n938), .A2(n1127), .ZN(n1125) );
  OR2_X1 U1104 ( .A1(n943), .A2(n944), .ZN(n1127) );
  OR2_X1 U1105 ( .A1(n1099), .A2(n1000), .ZN(n944) );
  OR2_X1 U1106 ( .A1(n1128), .A2(n1129), .ZN(n943) );
  AND2_X1 U1107 ( .A1(n933), .A2(n932), .ZN(n1129) );
  AND2_X1 U1108 ( .A1(n927), .A2(n1130), .ZN(n1128) );
  OR2_X1 U1109 ( .A1(n932), .A2(n933), .ZN(n1130) );
  OR2_X1 U1110 ( .A1(n1131), .A2(n1000), .ZN(n933) );
  OR2_X1 U1111 ( .A1(n1132), .A2(n1133), .ZN(n932) );
  AND2_X1 U1112 ( .A1(n1042), .A2(n1041), .ZN(n1133) );
  AND2_X1 U1113 ( .A1(n1036), .A2(n1134), .ZN(n1132) );
  OR2_X1 U1114 ( .A1(n1042), .A2(n1041), .ZN(n1134) );
  OR2_X1 U1115 ( .A1(n1135), .A2(n1136), .ZN(n1041) );
  AND2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1136) );
  AND2_X1 U1117 ( .A1(n1025), .A2(n1137), .ZN(n1135) );
  OR2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1137) );
  OR2_X1 U1119 ( .A1(n1138), .A2(n1139), .ZN(n1030) );
  AND2_X1 U1120 ( .A1(n1020), .A2(n1019), .ZN(n1139) );
  AND2_X1 U1121 ( .A1(n1014), .A2(n1140), .ZN(n1138) );
  OR2_X1 U1122 ( .A1(n1020), .A2(n1019), .ZN(n1140) );
  OR2_X1 U1123 ( .A1(n1141), .A2(n1142), .ZN(n1019) );
  AND2_X1 U1124 ( .A1(n1009), .A2(n1143), .ZN(n1142) );
  AND2_X1 U1125 ( .A1(n1004), .A2(n1144), .ZN(n1141) );
  OR2_X1 U1126 ( .A1(n1009), .A2(n1143), .ZN(n1144) );
  INV_X1 U1127 ( .A(n1010), .ZN(n1143) );
  AND2_X1 U1128 ( .A1(n1145), .A2(Result_15_), .ZN(n1010) );
  AND2_X1 U1129 ( .A1(n998), .A2(n1146), .ZN(Result_15_) );
  OR2_X1 U1130 ( .A1(n1147), .A2(n1000), .ZN(n1009) );
  AND2_X1 U1131 ( .A1(n1148), .A2(n1149), .ZN(n1004) );
  OR2_X1 U1132 ( .A1(n1150), .A2(n1145), .ZN(n1149) );
  INV_X1 U1133 ( .A(n1151), .ZN(n1148) );
  AND2_X1 U1134 ( .A1(n1145), .A2(n1150), .ZN(n1151) );
  OR2_X1 U1135 ( .A1(n1152), .A2(n1000), .ZN(n1020) );
  AND2_X1 U1136 ( .A1(n1153), .A2(n1154), .ZN(n1014) );
  INV_X1 U1137 ( .A(n1155), .ZN(n1154) );
  AND2_X1 U1138 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
  OR2_X1 U1139 ( .A1(n1157), .A2(n1156), .ZN(n1153) );
  OR2_X1 U1140 ( .A1(n1158), .A2(n1159), .ZN(n1156) );
  INV_X1 U1141 ( .A(n1160), .ZN(n1159) );
  OR2_X1 U1142 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
  AND2_X1 U1143 ( .A1(n1162), .A2(n1161), .ZN(n1158) );
  OR2_X1 U1144 ( .A1(n1163), .A2(n1000), .ZN(n1031) );
  AND2_X1 U1145 ( .A1(n1164), .A2(n1165), .ZN(n1025) );
  INV_X1 U1146 ( .A(n1166), .ZN(n1165) );
  AND2_X1 U1147 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
  OR2_X1 U1148 ( .A1(n1168), .A2(n1167), .ZN(n1164) );
  OR2_X1 U1149 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
  INV_X1 U1150 ( .A(n1171), .ZN(n1170) );
  OR2_X1 U1151 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
  AND2_X1 U1152 ( .A1(n1173), .A2(n1172), .ZN(n1169) );
  INV_X1 U1153 ( .A(n1174), .ZN(n1173) );
  OR2_X1 U1154 ( .A1(n1175), .A2(n1000), .ZN(n1042) );
  INV_X1 U1155 ( .A(n1146), .ZN(n1000) );
  AND2_X1 U1156 ( .A1(n1176), .A2(n1177), .ZN(n1146) );
  OR2_X1 U1157 ( .A1(c_7_), .A2(d_7_), .ZN(n1176) );
  AND2_X1 U1158 ( .A1(n1178), .A2(n1179), .ZN(n1036) );
  INV_X1 U1159 ( .A(n1180), .ZN(n1179) );
  AND2_X1 U1160 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
  OR2_X1 U1161 ( .A1(n1182), .A2(n1181), .ZN(n1178) );
  OR2_X1 U1162 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
  AND2_X1 U1163 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
  INV_X1 U1164 ( .A(n1187), .ZN(n1183) );
  OR2_X1 U1165 ( .A1(n1186), .A2(n1185), .ZN(n1187) );
  INV_X1 U1166 ( .A(n1188), .ZN(n1185) );
  AND2_X1 U1167 ( .A1(n1189), .A2(n1190), .ZN(n927) );
  INV_X1 U1168 ( .A(n1191), .ZN(n1190) );
  AND2_X1 U1169 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
  OR2_X1 U1170 ( .A1(n1193), .A2(n1192), .ZN(n1189) );
  OR2_X1 U1171 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
  INV_X1 U1172 ( .A(n1196), .ZN(n1195) );
  OR2_X1 U1173 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
  AND2_X1 U1174 ( .A1(n1198), .A2(n1197), .ZN(n1194) );
  INV_X1 U1175 ( .A(n1199), .ZN(n1198) );
  AND2_X1 U1176 ( .A1(n1200), .A2(n1201), .ZN(n938) );
  INV_X1 U1177 ( .A(n1202), .ZN(n1201) );
  AND2_X1 U1178 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
  OR2_X1 U1179 ( .A1(n1204), .A2(n1203), .ZN(n1200) );
  OR2_X1 U1180 ( .A1(n1205), .A2(n1206), .ZN(n1203) );
  INV_X1 U1181 ( .A(n1207), .ZN(n1206) );
  OR2_X1 U1182 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
  AND2_X1 U1183 ( .A1(n1209), .A2(n1208), .ZN(n1205) );
  INV_X1 U1184 ( .A(n1210), .ZN(n1209) );
  AND2_X1 U1185 ( .A1(n1211), .A2(n1212), .ZN(n950) );
  INV_X1 U1186 ( .A(n1213), .ZN(n1212) );
  AND2_X1 U1187 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
  OR2_X1 U1188 ( .A1(n1215), .A2(n1214), .ZN(n1211) );
  OR2_X1 U1189 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
  AND2_X1 U1190 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
  AND2_X1 U1191 ( .A1(n1220), .A2(n1221), .ZN(n1216) );
  INV_X1 U1192 ( .A(n1219), .ZN(n1220) );
  OR3_X1 U1193 ( .A1(n1123), .A2(n1124), .A3(n1122), .ZN(n1117) );
  OR2_X1 U1194 ( .A1(n1222), .A2(n1223), .ZN(n1122) );
  AND2_X1 U1195 ( .A1(n1221), .A2(n1219), .ZN(n1223) );
  AND2_X1 U1196 ( .A1(n1215), .A2(n1224), .ZN(n1222) );
  OR2_X1 U1197 ( .A1(n1219), .A2(n1221), .ZN(n1224) );
  INV_X1 U1198 ( .A(n1218), .ZN(n1221) );
  AND2_X1 U1199 ( .A1(n997), .A2(n1047), .ZN(n1218) );
  OR2_X1 U1200 ( .A1(n1225), .A2(n1226), .ZN(n1219) );
  AND2_X1 U1201 ( .A1(n1208), .A2(n1210), .ZN(n1226) );
  AND2_X1 U1202 ( .A1(n1204), .A2(n1227), .ZN(n1225) );
  OR2_X1 U1203 ( .A1(n1210), .A2(n1208), .ZN(n1227) );
  OR2_X1 U1204 ( .A1(n1228), .A2(n1131), .ZN(n1208) );
  OR2_X1 U1205 ( .A1(n1229), .A2(n1230), .ZN(n1210) );
  AND2_X1 U1206 ( .A1(n1197), .A2(n1199), .ZN(n1230) );
  AND2_X1 U1207 ( .A1(n1193), .A2(n1231), .ZN(n1229) );
  OR2_X1 U1208 ( .A1(n1199), .A2(n1197), .ZN(n1231) );
  OR2_X1 U1209 ( .A1(n1228), .A2(n1175), .ZN(n1197) );
  OR2_X1 U1210 ( .A1(n1232), .A2(n1233), .ZN(n1199) );
  AND2_X1 U1211 ( .A1(n1188), .A2(n1186), .ZN(n1233) );
  AND2_X1 U1212 ( .A1(n1182), .A2(n1234), .ZN(n1232) );
  OR2_X1 U1213 ( .A1(n1188), .A2(n1186), .ZN(n1234) );
  OR2_X1 U1214 ( .A1(n1235), .A2(n1236), .ZN(n1186) );
  AND2_X1 U1215 ( .A1(n1172), .A2(n1174), .ZN(n1236) );
  AND2_X1 U1216 ( .A1(n1168), .A2(n1237), .ZN(n1235) );
  OR2_X1 U1217 ( .A1(n1172), .A2(n1174), .ZN(n1237) );
  OR2_X1 U1218 ( .A1(n1238), .A2(n1239), .ZN(n1174) );
  AND2_X1 U1219 ( .A1(n1161), .A2(n1240), .ZN(n1239) );
  AND2_X1 U1220 ( .A1(n1157), .A2(n1241), .ZN(n1238) );
  OR2_X1 U1221 ( .A1(n1161), .A2(n1240), .ZN(n1241) );
  INV_X1 U1222 ( .A(n1162), .ZN(n1240) );
  AND2_X1 U1223 ( .A1(n1242), .A2(n1145), .ZN(n1162) );
  AND2_X1 U1224 ( .A1(n1243), .A2(n997), .ZN(n1145) );
  INV_X1 U1225 ( .A(n1150), .ZN(n1242) );
  OR2_X1 U1226 ( .A1(n1244), .A2(n1245), .ZN(n1150) );
  OR2_X1 U1227 ( .A1(n1228), .A2(n1147), .ZN(n1161) );
  AND2_X1 U1228 ( .A1(n1246), .A2(n1247), .ZN(n1157) );
  OR3_X1 U1229 ( .A1(n999), .A2(n1245), .A3(n1248), .ZN(n1247) );
  OR2_X1 U1230 ( .A1(n1249), .A2(n1250), .ZN(n1246) );
  INV_X1 U1231 ( .A(n1251), .ZN(n1250) );
  OR2_X1 U1232 ( .A1(n999), .A2(n1245), .ZN(n1251) );
  OR2_X1 U1233 ( .A1(n1152), .A2(n1228), .ZN(n1172) );
  AND2_X1 U1234 ( .A1(n1252), .A2(n1253), .ZN(n1168) );
  INV_X1 U1235 ( .A(n1254), .ZN(n1253) );
  AND2_X1 U1236 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
  OR2_X1 U1237 ( .A1(n1256), .A2(n1255), .ZN(n1252) );
  OR2_X1 U1238 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
  INV_X1 U1239 ( .A(n1259), .ZN(n1258) );
  OR2_X1 U1240 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
  AND2_X1 U1241 ( .A1(n1261), .A2(n1260), .ZN(n1257) );
  INV_X1 U1242 ( .A(n1262), .ZN(n1261) );
  OR2_X1 U1243 ( .A1(n1163), .A2(n1228), .ZN(n1188) );
  INV_X1 U1244 ( .A(n997), .ZN(n1228) );
  OR2_X1 U1245 ( .A1(n1263), .A2(n1264), .ZN(n997) );
  AND3_X1 U1246 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1264) );
  OR2_X1 U1247 ( .A1(c_6_), .A2(n1268), .ZN(n1266) );
  OR2_X1 U1248 ( .A1(d_6_), .A2(n1269), .ZN(n1265) );
  AND2_X1 U1249 ( .A1(n1270), .A2(n1177), .ZN(n1263) );
  INV_X1 U1250 ( .A(n1267), .ZN(n1177) );
  OR2_X1 U1251 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
  AND2_X1 U1252 ( .A1(c_6_), .A2(n1268), .ZN(n1272) );
  INV_X1 U1253 ( .A(d_6_), .ZN(n1268) );
  AND2_X1 U1254 ( .A1(d_6_), .A2(n1269), .ZN(n1271) );
  INV_X1 U1255 ( .A(c_6_), .ZN(n1269) );
  AND2_X1 U1256 ( .A1(n1273), .A2(n1274), .ZN(n1182) );
  INV_X1 U1257 ( .A(n1275), .ZN(n1274) );
  AND2_X1 U1258 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
  OR2_X1 U1259 ( .A1(n1277), .A2(n1276), .ZN(n1273) );
  OR2_X1 U1260 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
  AND2_X1 U1261 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
  INV_X1 U1262 ( .A(n1282), .ZN(n1278) );
  OR2_X1 U1263 ( .A1(n1281), .A2(n1280), .ZN(n1282) );
  INV_X1 U1264 ( .A(n1283), .ZN(n1280) );
  AND2_X1 U1265 ( .A1(n1284), .A2(n1285), .ZN(n1193) );
  INV_X1 U1266 ( .A(n1286), .ZN(n1285) );
  AND2_X1 U1267 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
  OR2_X1 U1268 ( .A1(n1288), .A2(n1287), .ZN(n1284) );
  OR2_X1 U1269 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
  INV_X1 U1270 ( .A(n1291), .ZN(n1290) );
  OR2_X1 U1271 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
  AND2_X1 U1272 ( .A1(n1293), .A2(n1292), .ZN(n1289) );
  INV_X1 U1273 ( .A(n1294), .ZN(n1293) );
  AND2_X1 U1274 ( .A1(n1295), .A2(n1296), .ZN(n1204) );
  INV_X1 U1275 ( .A(n1297), .ZN(n1296) );
  AND2_X1 U1276 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
  OR2_X1 U1277 ( .A1(n1299), .A2(n1298), .ZN(n1295) );
  OR2_X1 U1278 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
  INV_X1 U1279 ( .A(n1302), .ZN(n1301) );
  OR2_X1 U1280 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
  AND2_X1 U1281 ( .A1(n1304), .A2(n1303), .ZN(n1300) );
  INV_X1 U1282 ( .A(n1305), .ZN(n1304) );
  AND2_X1 U1283 ( .A1(n1306), .A2(n1307), .ZN(n1215) );
  INV_X1 U1284 ( .A(n1308), .ZN(n1307) );
  AND2_X1 U1285 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
  OR2_X1 U1286 ( .A1(n1310), .A2(n1309), .ZN(n1306) );
  OR2_X1 U1287 ( .A1(n1311), .A2(n1312), .ZN(n1309) );
  INV_X1 U1288 ( .A(n1313), .ZN(n1312) );
  OR2_X1 U1289 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
  AND2_X1 U1290 ( .A1(n1315), .A2(n1314), .ZN(n1311) );
  INV_X1 U1291 ( .A(n1316), .ZN(n1315) );
  AND2_X1 U1292 ( .A1(n1317), .A2(n1318), .ZN(n1124) );
  AND2_X1 U1293 ( .A1(n1086), .A2(n1319), .ZN(n1123) );
  INV_X1 U1294 ( .A(n1317), .ZN(n1319) );
  OR2_X1 U1295 ( .A1(n1320), .A2(n1321), .ZN(n1317) );
  AND2_X1 U1296 ( .A1(n1322), .A2(n1089), .ZN(n1321) );
  INV_X1 U1297 ( .A(n1323), .ZN(n1320) );
  OR2_X1 U1298 ( .A1(n1089), .A2(n1322), .ZN(n1323) );
  INV_X1 U1299 ( .A(n1087), .ZN(n1322) );
  OR2_X1 U1300 ( .A1(n1099), .A2(n1245), .ZN(n1087) );
  OR2_X1 U1301 ( .A1(n1324), .A2(n1325), .ZN(n1089) );
  AND2_X1 U1302 ( .A1(n1314), .A2(n1316), .ZN(n1325) );
  AND2_X1 U1303 ( .A1(n1310), .A2(n1326), .ZN(n1324) );
  OR2_X1 U1304 ( .A1(n1316), .A2(n1314), .ZN(n1326) );
  OR2_X1 U1305 ( .A1(n1131), .A2(n1245), .ZN(n1314) );
  OR2_X1 U1306 ( .A1(n1327), .A2(n1328), .ZN(n1316) );
  AND2_X1 U1307 ( .A1(n1303), .A2(n1305), .ZN(n1328) );
  AND2_X1 U1308 ( .A1(n1299), .A2(n1329), .ZN(n1327) );
  OR2_X1 U1309 ( .A1(n1305), .A2(n1303), .ZN(n1329) );
  OR2_X1 U1310 ( .A1(n1175), .A2(n1245), .ZN(n1303) );
  OR2_X1 U1311 ( .A1(n1330), .A2(n1331), .ZN(n1305) );
  AND2_X1 U1312 ( .A1(n1292), .A2(n1294), .ZN(n1331) );
  AND2_X1 U1313 ( .A1(n1288), .A2(n1332), .ZN(n1330) );
  OR2_X1 U1314 ( .A1(n1294), .A2(n1292), .ZN(n1332) );
  OR2_X1 U1315 ( .A1(n1163), .A2(n1245), .ZN(n1292) );
  OR2_X1 U1316 ( .A1(n1333), .A2(n1334), .ZN(n1294) );
  AND2_X1 U1317 ( .A1(n1283), .A2(n1281), .ZN(n1334) );
  AND2_X1 U1318 ( .A1(n1277), .A2(n1335), .ZN(n1333) );
  OR2_X1 U1319 ( .A1(n1283), .A2(n1281), .ZN(n1335) );
  OR2_X1 U1320 ( .A1(n1336), .A2(n1337), .ZN(n1281) );
  AND2_X1 U1321 ( .A1(n1260), .A2(n1262), .ZN(n1337) );
  AND2_X1 U1322 ( .A1(n1256), .A2(n1338), .ZN(n1336) );
  OR2_X1 U1323 ( .A1(n1260), .A2(n1262), .ZN(n1338) );
  OR3_X1 U1324 ( .A1(n999), .A2(n1249), .A3(n1245), .ZN(n1262) );
  OR2_X1 U1325 ( .A1(n1147), .A2(n1245), .ZN(n1260) );
  AND2_X1 U1326 ( .A1(n1339), .A2(n1340), .ZN(n1256) );
  OR2_X1 U1327 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
  INV_X1 U1328 ( .A(n1343), .ZN(n1339) );
  AND2_X1 U1329 ( .A1(n1342), .A2(n1341), .ZN(n1343) );
  OR2_X1 U1330 ( .A1(n1344), .A2(n1244), .ZN(n1341) );
  AND2_X1 U1331 ( .A1(n1243), .A2(n1345), .ZN(n1342) );
  OR2_X1 U1332 ( .A1(n1152), .A2(n1245), .ZN(n1283) );
  OR2_X1 U1333 ( .A1(n1346), .A2(n1347), .ZN(n1245) );
  AND2_X1 U1334 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
  INV_X1 U1335 ( .A(n1350), .ZN(n1346) );
  OR2_X1 U1336 ( .A1(n1348), .A2(n1349), .ZN(n1350) );
  OR2_X1 U1337 ( .A1(n1351), .A2(n1352), .ZN(n1348) );
  AND2_X1 U1338 ( .A1(c_5_), .A2(n1353), .ZN(n1352) );
  AND2_X1 U1339 ( .A1(d_5_), .A2(n1354), .ZN(n1351) );
  AND2_X1 U1340 ( .A1(n1355), .A2(n1356), .ZN(n1277) );
  INV_X1 U1341 ( .A(n1357), .ZN(n1356) );
  AND2_X1 U1342 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
  OR2_X1 U1343 ( .A1(n1359), .A2(n1358), .ZN(n1355) );
  OR2_X1 U1344 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
  INV_X1 U1345 ( .A(n1362), .ZN(n1361) );
  OR2_X1 U1346 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
  AND2_X1 U1347 ( .A1(n1364), .A2(n1363), .ZN(n1360) );
  INV_X1 U1348 ( .A(n1365), .ZN(n1364) );
  AND2_X1 U1349 ( .A1(n1366), .A2(n1367), .ZN(n1288) );
  INV_X1 U1350 ( .A(n1368), .ZN(n1367) );
  AND2_X1 U1351 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
  OR2_X1 U1352 ( .A1(n1370), .A2(n1369), .ZN(n1366) );
  OR2_X1 U1353 ( .A1(n1371), .A2(n1372), .ZN(n1369) );
  INV_X1 U1354 ( .A(n1373), .ZN(n1372) );
  OR2_X1 U1355 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
  AND2_X1 U1356 ( .A1(n1375), .A2(n1374), .ZN(n1371) );
  INV_X1 U1357 ( .A(n1376), .ZN(n1375) );
  AND2_X1 U1358 ( .A1(n1377), .A2(n1378), .ZN(n1299) );
  INV_X1 U1359 ( .A(n1379), .ZN(n1378) );
  AND2_X1 U1360 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
  OR2_X1 U1361 ( .A1(n1381), .A2(n1380), .ZN(n1377) );
  OR2_X1 U1362 ( .A1(n1382), .A2(n1383), .ZN(n1380) );
  INV_X1 U1363 ( .A(n1384), .ZN(n1383) );
  OR2_X1 U1364 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
  AND2_X1 U1365 ( .A1(n1386), .A2(n1385), .ZN(n1382) );
  INV_X1 U1366 ( .A(n1387), .ZN(n1386) );
  AND2_X1 U1367 ( .A1(n1388), .A2(n1389), .ZN(n1310) );
  INV_X1 U1368 ( .A(n1390), .ZN(n1389) );
  AND2_X1 U1369 ( .A1(n1391), .A2(n1392), .ZN(n1390) );
  OR2_X1 U1370 ( .A1(n1392), .A2(n1391), .ZN(n1388) );
  OR2_X1 U1371 ( .A1(n1393), .A2(n1394), .ZN(n1391) );
  INV_X1 U1372 ( .A(n1395), .ZN(n1394) );
  OR2_X1 U1373 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
  AND2_X1 U1374 ( .A1(n1397), .A2(n1396), .ZN(n1393) );
  INV_X1 U1375 ( .A(n1398), .ZN(n1397) );
  INV_X1 U1376 ( .A(n1318), .ZN(n1086) );
  AND2_X1 U1377 ( .A1(n1399), .A2(n1400), .ZN(n1318) );
  OR2_X1 U1378 ( .A1(n1401), .A2(n1102), .ZN(n1400) );
  INV_X1 U1379 ( .A(n1402), .ZN(n1399) );
  AND2_X1 U1380 ( .A1(n1102), .A2(n1401), .ZN(n1402) );
  AND2_X1 U1381 ( .A1(n1403), .A2(n1404), .ZN(n1401) );
  OR2_X1 U1382 ( .A1(n1103), .A2(n1405), .ZN(n1404) );
  INV_X1 U1383 ( .A(n1406), .ZN(n1403) );
  AND2_X1 U1384 ( .A1(n1405), .A2(n1103), .ZN(n1406) );
  OR2_X1 U1385 ( .A1(n1098), .A2(n1131), .ZN(n1103) );
  INV_X1 U1386 ( .A(n1105), .ZN(n1405) );
  OR2_X1 U1387 ( .A1(n1407), .A2(n1408), .ZN(n1105) );
  AND2_X1 U1388 ( .A1(n1396), .A2(n1398), .ZN(n1408) );
  AND2_X1 U1389 ( .A1(n1392), .A2(n1409), .ZN(n1407) );
  OR2_X1 U1390 ( .A1(n1398), .A2(n1396), .ZN(n1409) );
  OR2_X1 U1391 ( .A1(n1098), .A2(n1175), .ZN(n1396) );
  OR2_X1 U1392 ( .A1(n1410), .A2(n1411), .ZN(n1398) );
  AND2_X1 U1393 ( .A1(n1385), .A2(n1387), .ZN(n1411) );
  AND2_X1 U1394 ( .A1(n1381), .A2(n1412), .ZN(n1410) );
  OR2_X1 U1395 ( .A1(n1387), .A2(n1385), .ZN(n1412) );
  OR2_X1 U1396 ( .A1(n1098), .A2(n1163), .ZN(n1385) );
  OR2_X1 U1397 ( .A1(n1413), .A2(n1414), .ZN(n1387) );
  AND2_X1 U1398 ( .A1(n1374), .A2(n1376), .ZN(n1414) );
  AND2_X1 U1399 ( .A1(n1370), .A2(n1415), .ZN(n1413) );
  OR2_X1 U1400 ( .A1(n1376), .A2(n1374), .ZN(n1415) );
  OR2_X1 U1401 ( .A1(n1098), .A2(n1152), .ZN(n1374) );
  OR2_X1 U1402 ( .A1(n1416), .A2(n1417), .ZN(n1376) );
  AND2_X1 U1403 ( .A1(n1363), .A2(n1365), .ZN(n1417) );
  AND2_X1 U1404 ( .A1(n1359), .A2(n1418), .ZN(n1416) );
  OR2_X1 U1405 ( .A1(n1363), .A2(n1365), .ZN(n1418) );
  OR2_X1 U1406 ( .A1(n1419), .A2(n1249), .ZN(n1365) );
  INV_X1 U1407 ( .A(n1248), .ZN(n1249) );
  AND2_X1 U1408 ( .A1(n1345), .A2(n998), .ZN(n1248) );
  OR2_X1 U1409 ( .A1(n1098), .A2(n1147), .ZN(n1363) );
  INV_X1 U1410 ( .A(n1345), .ZN(n1098) );
  OR2_X1 U1411 ( .A1(n1420), .A2(n1421), .ZN(n1345) );
  AND2_X1 U1412 ( .A1(n1422), .A2(n1423), .ZN(n1421) );
  INV_X1 U1413 ( .A(n1424), .ZN(n1420) );
  OR2_X1 U1414 ( .A1(n1422), .A2(n1423), .ZN(n1424) );
  OR2_X1 U1415 ( .A1(n1425), .A2(n1426), .ZN(n1422) );
  AND2_X1 U1416 ( .A1(c_4_), .A2(n1427), .ZN(n1426) );
  AND2_X1 U1417 ( .A1(d_4_), .A2(n1428), .ZN(n1425) );
  AND2_X1 U1418 ( .A1(n1429), .A2(n1430), .ZN(n1359) );
  INV_X1 U1419 ( .A(n1431), .ZN(n1430) );
  AND3_X1 U1420 ( .A1(n998), .A2(n1432), .A3(n1419), .ZN(n1431) );
  OR2_X1 U1421 ( .A1(n1419), .A2(n1433), .ZN(n1429) );
  AND2_X1 U1422 ( .A1(n1432), .A2(n998), .ZN(n1433) );
  INV_X1 U1423 ( .A(n1434), .ZN(n1432) );
  AND2_X1 U1424 ( .A1(n1435), .A2(n1436), .ZN(n1370) );
  INV_X1 U1425 ( .A(n1437), .ZN(n1436) );
  AND2_X1 U1426 ( .A1(n1438), .A2(n1439), .ZN(n1437) );
  OR2_X1 U1427 ( .A1(n1439), .A2(n1438), .ZN(n1435) );
  OR2_X1 U1428 ( .A1(n1440), .A2(n1441), .ZN(n1438) );
  AND2_X1 U1429 ( .A1(n1442), .A2(n1443), .ZN(n1441) );
  INV_X1 U1430 ( .A(n1444), .ZN(n1442) );
  AND2_X1 U1431 ( .A1(n1445), .A2(n1444), .ZN(n1440) );
  INV_X1 U1432 ( .A(n1443), .ZN(n1445) );
  AND2_X1 U1433 ( .A1(n1446), .A2(n1447), .ZN(n1381) );
  INV_X1 U1434 ( .A(n1448), .ZN(n1447) );
  AND2_X1 U1435 ( .A1(n1449), .A2(n1450), .ZN(n1448) );
  OR2_X1 U1436 ( .A1(n1450), .A2(n1449), .ZN(n1446) );
  OR2_X1 U1437 ( .A1(n1451), .A2(n1452), .ZN(n1449) );
  INV_X1 U1438 ( .A(n1453), .ZN(n1452) );
  OR2_X1 U1439 ( .A1(n1454), .A2(n1455), .ZN(n1453) );
  AND2_X1 U1440 ( .A1(n1455), .A2(n1454), .ZN(n1451) );
  INV_X1 U1441 ( .A(n1456), .ZN(n1455) );
  AND2_X1 U1442 ( .A1(n1457), .A2(n1458), .ZN(n1392) );
  INV_X1 U1443 ( .A(n1459), .ZN(n1458) );
  AND2_X1 U1444 ( .A1(n1460), .A2(n1461), .ZN(n1459) );
  OR2_X1 U1445 ( .A1(n1461), .A2(n1460), .ZN(n1457) );
  OR2_X1 U1446 ( .A1(n1462), .A2(n1463), .ZN(n1460) );
  INV_X1 U1447 ( .A(n1464), .ZN(n1463) );
  OR2_X1 U1448 ( .A1(n1465), .A2(n1466), .ZN(n1464) );
  AND2_X1 U1449 ( .A1(n1466), .A2(n1465), .ZN(n1462) );
  INV_X1 U1450 ( .A(n1467), .ZN(n1466) );
  OR2_X1 U1451 ( .A1(n1468), .A2(n1469), .ZN(n1102) );
  INV_X1 U1452 ( .A(n1470), .ZN(n1469) );
  OR2_X1 U1453 ( .A1(n1471), .A2(n1472), .ZN(n1470) );
  AND2_X1 U1454 ( .A1(n1472), .A2(n1471), .ZN(n1468) );
  AND2_X1 U1455 ( .A1(n1473), .A2(n1474), .ZN(n1471) );
  OR2_X1 U1456 ( .A1(n1475), .A2(n1476), .ZN(n1474) );
  INV_X1 U1457 ( .A(n1477), .ZN(n1473) );
  AND2_X1 U1458 ( .A1(n1476), .A2(n1475), .ZN(n1477) );
  INV_X1 U1459 ( .A(n1478), .ZN(n1476) );
  INV_X1 U1460 ( .A(n979), .ZN(n980) );
  OR2_X1 U1461 ( .A1(n1055), .A2(n1056), .ZN(n979) );
  OR2_X1 U1462 ( .A1(n1479), .A2(n1480), .ZN(n1056) );
  AND2_X1 U1463 ( .A1(n1076), .A2(n1078), .ZN(n1480) );
  AND2_X1 U1464 ( .A1(n1072), .A2(n1481), .ZN(n1479) );
  OR2_X1 U1465 ( .A1(n1078), .A2(n1076), .ZN(n1481) );
  OR2_X1 U1466 ( .A1(n1482), .A2(n1483), .ZN(n1076) );
  AND2_X1 U1467 ( .A1(n1114), .A2(n1116), .ZN(n1483) );
  AND2_X1 U1468 ( .A1(n1110), .A2(n1484), .ZN(n1482) );
  OR2_X1 U1469 ( .A1(n1116), .A2(n1114), .ZN(n1484) );
  OR2_X1 U1470 ( .A1(n1485), .A2(n1486), .ZN(n1114) );
  AND2_X1 U1471 ( .A1(n1475), .A2(n1478), .ZN(n1486) );
  AND2_X1 U1472 ( .A1(n1472), .A2(n1487), .ZN(n1485) );
  OR2_X1 U1473 ( .A1(n1478), .A2(n1475), .ZN(n1487) );
  OR2_X1 U1474 ( .A1(n1488), .A2(n1489), .ZN(n1475) );
  AND2_X1 U1475 ( .A1(n1465), .A2(n1467), .ZN(n1489) );
  AND2_X1 U1476 ( .A1(n1461), .A2(n1490), .ZN(n1488) );
  OR2_X1 U1477 ( .A1(n1467), .A2(n1465), .ZN(n1490) );
  OR2_X1 U1478 ( .A1(n1491), .A2(n1492), .ZN(n1465) );
  AND2_X1 U1479 ( .A1(n1454), .A2(n1456), .ZN(n1492) );
  AND2_X1 U1480 ( .A1(n1450), .A2(n1493), .ZN(n1491) );
  OR2_X1 U1481 ( .A1(n1456), .A2(n1454), .ZN(n1493) );
  OR2_X1 U1482 ( .A1(n1344), .A2(n1152), .ZN(n1454) );
  OR2_X1 U1483 ( .A1(n1494), .A2(n1495), .ZN(n1456) );
  AND2_X1 U1484 ( .A1(n1444), .A2(n1443), .ZN(n1495) );
  AND2_X1 U1485 ( .A1(n1439), .A2(n1496), .ZN(n1494) );
  OR2_X1 U1486 ( .A1(n1443), .A2(n1444), .ZN(n1496) );
  OR2_X1 U1487 ( .A1(n1344), .A2(n1147), .ZN(n1444) );
  OR3_X1 U1488 ( .A1(n1434), .A2(n1244), .A3(n1419), .ZN(n1443) );
  OR2_X1 U1489 ( .A1(n999), .A2(n1344), .ZN(n1419) );
  AND2_X1 U1490 ( .A1(n1497), .A2(n1498), .ZN(n1439) );
  OR2_X1 U1491 ( .A1(n1499), .A2(n1500), .ZN(n1498) );
  INV_X1 U1492 ( .A(n1501), .ZN(n1500) );
  OR2_X1 U1493 ( .A1(n1501), .A2(n1502), .ZN(n1497) );
  INV_X1 U1494 ( .A(n1499), .ZN(n1502) );
  AND2_X1 U1495 ( .A1(n1503), .A2(n1504), .ZN(n1450) );
  INV_X1 U1496 ( .A(n1505), .ZN(n1504) );
  AND2_X1 U1497 ( .A1(n1506), .A2(n1507), .ZN(n1505) );
  OR2_X1 U1498 ( .A1(n1507), .A2(n1506), .ZN(n1503) );
  OR2_X1 U1499 ( .A1(n1508), .A2(n1509), .ZN(n1506) );
  AND2_X1 U1500 ( .A1(n1510), .A2(n1511), .ZN(n1509) );
  INV_X1 U1501 ( .A(n1512), .ZN(n1510) );
  AND2_X1 U1502 ( .A1(n1513), .A2(n1512), .ZN(n1508) );
  INV_X1 U1503 ( .A(n1511), .ZN(n1513) );
  OR2_X1 U1504 ( .A1(n1344), .A2(n1163), .ZN(n1467) );
  AND2_X1 U1505 ( .A1(n1514), .A2(n1515), .ZN(n1461) );
  INV_X1 U1506 ( .A(n1516), .ZN(n1515) );
  AND2_X1 U1507 ( .A1(n1517), .A2(n1518), .ZN(n1516) );
  OR2_X1 U1508 ( .A1(n1518), .A2(n1517), .ZN(n1514) );
  OR2_X1 U1509 ( .A1(n1519), .A2(n1520), .ZN(n1517) );
  INV_X1 U1510 ( .A(n1521), .ZN(n1520) );
  OR2_X1 U1511 ( .A1(n1522), .A2(n1523), .ZN(n1521) );
  AND2_X1 U1512 ( .A1(n1523), .A2(n1522), .ZN(n1519) );
  INV_X1 U1513 ( .A(n1524), .ZN(n1523) );
  OR2_X1 U1514 ( .A1(n1344), .A2(n1175), .ZN(n1478) );
  OR2_X1 U1515 ( .A1(n1525), .A2(n1526), .ZN(n1472) );
  INV_X1 U1516 ( .A(n1527), .ZN(n1526) );
  OR2_X1 U1517 ( .A1(n1528), .A2(n1529), .ZN(n1527) );
  AND2_X1 U1518 ( .A1(n1529), .A2(n1528), .ZN(n1525) );
  AND2_X1 U1519 ( .A1(n1530), .A2(n1531), .ZN(n1528) );
  OR2_X1 U1520 ( .A1(n1532), .A2(n1533), .ZN(n1531) );
  INV_X1 U1521 ( .A(n1534), .ZN(n1530) );
  AND2_X1 U1522 ( .A1(n1533), .A2(n1532), .ZN(n1534) );
  INV_X1 U1523 ( .A(n1535), .ZN(n1533) );
  OR2_X1 U1524 ( .A1(n1344), .A2(n1131), .ZN(n1116) );
  AND2_X1 U1525 ( .A1(n1536), .A2(n1537), .ZN(n1110) );
  INV_X1 U1526 ( .A(n1538), .ZN(n1537) );
  AND2_X1 U1527 ( .A1(n1539), .A2(n1540), .ZN(n1538) );
  OR2_X1 U1528 ( .A1(n1540), .A2(n1539), .ZN(n1536) );
  OR2_X1 U1529 ( .A1(n1541), .A2(n1542), .ZN(n1539) );
  INV_X1 U1530 ( .A(n1543), .ZN(n1542) );
  OR2_X1 U1531 ( .A1(n1544), .A2(n1545), .ZN(n1543) );
  AND2_X1 U1532 ( .A1(n1545), .A2(n1544), .ZN(n1541) );
  INV_X1 U1533 ( .A(n1546), .ZN(n1545) );
  OR2_X1 U1534 ( .A1(n1344), .A2(n1099), .ZN(n1078) );
  AND2_X1 U1535 ( .A1(n1547), .A2(n1548), .ZN(n1344) );
  INV_X1 U1536 ( .A(n1549), .ZN(n1548) );
  AND2_X1 U1537 ( .A1(n1550), .A2(n1551), .ZN(n1549) );
  OR2_X1 U1538 ( .A1(n1550), .A2(n1551), .ZN(n1547) );
  OR2_X1 U1539 ( .A1(n1552), .A2(n1553), .ZN(n1550) );
  AND2_X1 U1540 ( .A1(c_3_), .A2(n1554), .ZN(n1553) );
  AND2_X1 U1541 ( .A1(d_3_), .A2(n1555), .ZN(n1552) );
  AND2_X1 U1542 ( .A1(n1556), .A2(n1557), .ZN(n1072) );
  INV_X1 U1543 ( .A(n1558), .ZN(n1557) );
  AND2_X1 U1544 ( .A1(n1559), .A2(n1560), .ZN(n1558) );
  OR2_X1 U1545 ( .A1(n1560), .A2(n1559), .ZN(n1556) );
  OR2_X1 U1546 ( .A1(n1561), .A2(n1562), .ZN(n1559) );
  INV_X1 U1547 ( .A(n1563), .ZN(n1562) );
  OR2_X1 U1548 ( .A1(n1564), .A2(n1565), .ZN(n1563) );
  AND2_X1 U1549 ( .A1(n1565), .A2(n1564), .ZN(n1561) );
  INV_X1 U1550 ( .A(n1566), .ZN(n1565) );
  AND2_X1 U1551 ( .A1(n1567), .A2(n1568), .ZN(n1055) );
  INV_X1 U1552 ( .A(n1569), .ZN(n1568) );
  AND2_X1 U1553 ( .A1(n1570), .A2(n1571), .ZN(n1569) );
  OR2_X1 U1554 ( .A1(n1571), .A2(n1570), .ZN(n1567) );
  OR2_X1 U1555 ( .A1(n1572), .A2(n1573), .ZN(n1570) );
  INV_X1 U1556 ( .A(n1574), .ZN(n1573) );
  OR2_X1 U1557 ( .A1(n1575), .A2(n1576), .ZN(n1574) );
  AND2_X1 U1558 ( .A1(n1576), .A2(n1575), .ZN(n1572) );
  INV_X1 U1559 ( .A(n1577), .ZN(n1576) );
  AND3_X1 U1560 ( .A1(n1053), .A2(n1048), .A3(n1052), .ZN(n986) );
  INV_X1 U1561 ( .A(n991), .ZN(n1052) );
  OR2_X1 U1562 ( .A1(n1578), .A2(n1579), .ZN(n991) );
  AND2_X1 U1563 ( .A1(n1575), .A2(n1577), .ZN(n1579) );
  AND2_X1 U1564 ( .A1(n1571), .A2(n1580), .ZN(n1578) );
  OR2_X1 U1565 ( .A1(n1577), .A2(n1575), .ZN(n1580) );
  OR2_X1 U1566 ( .A1(n1434), .A2(n1099), .ZN(n1575) );
  OR2_X1 U1567 ( .A1(n1581), .A2(n1582), .ZN(n1577) );
  AND2_X1 U1568 ( .A1(n1564), .A2(n1566), .ZN(n1582) );
  AND2_X1 U1569 ( .A1(n1560), .A2(n1583), .ZN(n1581) );
  OR2_X1 U1570 ( .A1(n1566), .A2(n1564), .ZN(n1583) );
  OR2_X1 U1571 ( .A1(n1434), .A2(n1131), .ZN(n1564) );
  OR2_X1 U1572 ( .A1(n1584), .A2(n1585), .ZN(n1566) );
  AND2_X1 U1573 ( .A1(n1544), .A2(n1546), .ZN(n1585) );
  AND2_X1 U1574 ( .A1(n1540), .A2(n1586), .ZN(n1584) );
  OR2_X1 U1575 ( .A1(n1546), .A2(n1544), .ZN(n1586) );
  OR2_X1 U1576 ( .A1(n1587), .A2(n1588), .ZN(n1544) );
  AND2_X1 U1577 ( .A1(n1532), .A2(n1535), .ZN(n1588) );
  AND2_X1 U1578 ( .A1(n1529), .A2(n1589), .ZN(n1587) );
  OR2_X1 U1579 ( .A1(n1535), .A2(n1532), .ZN(n1589) );
  OR2_X1 U1580 ( .A1(n1590), .A2(n1591), .ZN(n1532) );
  AND2_X1 U1581 ( .A1(n1522), .A2(n1524), .ZN(n1591) );
  AND2_X1 U1582 ( .A1(n1518), .A2(n1592), .ZN(n1590) );
  OR2_X1 U1583 ( .A1(n1524), .A2(n1522), .ZN(n1592) );
  OR2_X1 U1584 ( .A1(n1434), .A2(n1152), .ZN(n1522) );
  OR2_X1 U1585 ( .A1(n1593), .A2(n1594), .ZN(n1524) );
  AND2_X1 U1586 ( .A1(n1512), .A2(n1511), .ZN(n1594) );
  AND2_X1 U1587 ( .A1(n1507), .A2(n1595), .ZN(n1593) );
  OR2_X1 U1588 ( .A1(n1511), .A2(n1512), .ZN(n1595) );
  OR2_X1 U1589 ( .A1(n1434), .A2(n1147), .ZN(n1512) );
  OR2_X1 U1590 ( .A1(n1501), .A2(n1499), .ZN(n1511) );
  OR2_X1 U1591 ( .A1(n1434), .A2(n999), .ZN(n1501) );
  AND2_X1 U1592 ( .A1(n1596), .A2(n1597), .ZN(n1507) );
  INV_X1 U1593 ( .A(n1598), .ZN(n1597) );
  AND3_X1 U1594 ( .A1(n998), .A2(n1599), .A3(n1600), .ZN(n1598) );
  OR2_X1 U1595 ( .A1(n1600), .A2(n1601), .ZN(n1596) );
  AND2_X1 U1596 ( .A1(n1599), .A2(n998), .ZN(n1601) );
  AND2_X1 U1597 ( .A1(n1602), .A2(n1603), .ZN(n1518) );
  INV_X1 U1598 ( .A(n1604), .ZN(n1603) );
  AND2_X1 U1599 ( .A1(n1605), .A2(n1606), .ZN(n1604) );
  OR2_X1 U1600 ( .A1(n1606), .A2(n1605), .ZN(n1602) );
  AND2_X1 U1601 ( .A1(n1607), .A2(n1608), .ZN(n1605) );
  OR2_X1 U1602 ( .A1(n1609), .A2(n1147), .ZN(n1606) );
  OR2_X1 U1603 ( .A1(n1434), .A2(n1163), .ZN(n1535) );
  OR2_X1 U1604 ( .A1(n1610), .A2(n1611), .ZN(n1529) );
  AND2_X1 U1605 ( .A1(n1612), .A2(n1613), .ZN(n1611) );
  INV_X1 U1606 ( .A(n1614), .ZN(n1610) );
  OR2_X1 U1607 ( .A1(n1612), .A2(n1613), .ZN(n1614) );
  OR2_X1 U1608 ( .A1(n1615), .A2(n1616), .ZN(n1612) );
  INV_X1 U1609 ( .A(n1617), .ZN(n1616) );
  OR2_X1 U1610 ( .A1(n1618), .A2(n1619), .ZN(n1617) );
  AND2_X1 U1611 ( .A1(n1619), .A2(n1618), .ZN(n1615) );
  OR2_X1 U1612 ( .A1(n1434), .A2(n1175), .ZN(n1546) );
  AND2_X1 U1613 ( .A1(n1620), .A2(n1621), .ZN(n1434) );
  INV_X1 U1614 ( .A(n1622), .ZN(n1621) );
  AND2_X1 U1615 ( .A1(n1623), .A2(n1624), .ZN(n1622) );
  OR2_X1 U1616 ( .A1(n1623), .A2(n1624), .ZN(n1620) );
  OR2_X1 U1617 ( .A1(n1625), .A2(n1626), .ZN(n1623) );
  AND2_X1 U1618 ( .A1(c_2_), .A2(n1627), .ZN(n1626) );
  AND2_X1 U1619 ( .A1(d_2_), .A2(n1628), .ZN(n1625) );
  AND2_X1 U1620 ( .A1(n1629), .A2(n1630), .ZN(n1540) );
  INV_X1 U1621 ( .A(n1631), .ZN(n1630) );
  AND2_X1 U1622 ( .A1(n1632), .A2(n1633), .ZN(n1631) );
  OR2_X1 U1623 ( .A1(n1632), .A2(n1633), .ZN(n1629) );
  OR2_X1 U1624 ( .A1(n1634), .A2(n1635), .ZN(n1632) );
  INV_X1 U1625 ( .A(n1636), .ZN(n1635) );
  OR2_X1 U1626 ( .A1(n1637), .A2(n1638), .ZN(n1636) );
  AND2_X1 U1627 ( .A1(n1638), .A2(n1637), .ZN(n1634) );
  INV_X1 U1628 ( .A(n1639), .ZN(n1638) );
  AND2_X1 U1629 ( .A1(n1640), .A2(n1641), .ZN(n1560) );
  INV_X1 U1630 ( .A(n1642), .ZN(n1641) );
  AND2_X1 U1631 ( .A1(n1643), .A2(n1644), .ZN(n1642) );
  OR2_X1 U1632 ( .A1(n1643), .A2(n1644), .ZN(n1640) );
  OR2_X1 U1633 ( .A1(n1645), .A2(n1646), .ZN(n1643) );
  INV_X1 U1634 ( .A(n1647), .ZN(n1646) );
  OR2_X1 U1635 ( .A1(n1648), .A2(n1649), .ZN(n1647) );
  AND2_X1 U1636 ( .A1(n1649), .A2(n1648), .ZN(n1645) );
  INV_X1 U1637 ( .A(n1650), .ZN(n1649) );
  AND2_X1 U1638 ( .A1(n1651), .A2(n1652), .ZN(n1571) );
  INV_X1 U1639 ( .A(n1653), .ZN(n1652) );
  AND2_X1 U1640 ( .A1(n1654), .A2(n1655), .ZN(n1653) );
  OR2_X1 U1641 ( .A1(n1654), .A2(n1655), .ZN(n1651) );
  OR2_X1 U1642 ( .A1(n1656), .A2(n1657), .ZN(n1654) );
  INV_X1 U1643 ( .A(n1658), .ZN(n1657) );
  OR2_X1 U1644 ( .A1(n1659), .A2(n1660), .ZN(n1658) );
  AND2_X1 U1645 ( .A1(n1660), .A2(n1659), .ZN(n1656) );
  INV_X1 U1646 ( .A(n1661), .ZN(n1660) );
  INV_X1 U1647 ( .A(n988), .ZN(n1048) );
  AND2_X1 U1648 ( .A1(n1662), .A2(n1663), .ZN(n988) );
  OR2_X1 U1649 ( .A1(n1664), .A2(n1046), .ZN(n1663) );
  INV_X1 U1650 ( .A(n1665), .ZN(n1046) );
  OR2_X1 U1651 ( .A1(n1665), .A2(n1666), .ZN(n1662) );
  INV_X1 U1652 ( .A(n1664), .ZN(n1666) );
  OR2_X1 U1653 ( .A1(n1667), .A2(n1099), .ZN(n1664) );
  OR2_X1 U1654 ( .A1(n1668), .A2(n1669), .ZN(n1665) );
  AND2_X1 U1655 ( .A1(n1670), .A2(n1671), .ZN(n1669) );
  AND2_X1 U1656 ( .A1(n1672), .A2(n1673), .ZN(n1668) );
  OR2_X1 U1657 ( .A1(n1671), .A2(n1670), .ZN(n1672) );
  OR2_X1 U1658 ( .A1(n1674), .A2(n1675), .ZN(n1053) );
  AND2_X1 U1659 ( .A1(n1676), .A2(n1670), .ZN(n1675) );
  INV_X1 U1660 ( .A(n1677), .ZN(n1674) );
  OR2_X1 U1661 ( .A1(n1676), .A2(n1670), .ZN(n1677) );
  OR2_X1 U1662 ( .A1(n1131), .A2(n1667), .ZN(n1670) );
  OR2_X1 U1663 ( .A1(n1678), .A2(n1679), .ZN(n1676) );
  INV_X1 U1664 ( .A(n1680), .ZN(n1679) );
  OR2_X1 U1665 ( .A1(n1673), .A2(n1681), .ZN(n1680) );
  AND2_X1 U1666 ( .A1(n1681), .A2(n1673), .ZN(n1678) );
  OR2_X1 U1667 ( .A1(n1609), .A2(n1099), .ZN(n1673) );
  INV_X1 U1668 ( .A(n1047), .ZN(n1099) );
  OR2_X1 U1669 ( .A1(n1682), .A2(n1683), .ZN(n1047) );
  AND2_X1 U1670 ( .A1(n1684), .A2(n1685), .ZN(n1683) );
  INV_X1 U1671 ( .A(n1686), .ZN(n1682) );
  OR2_X1 U1672 ( .A1(n1685), .A2(n1684), .ZN(n1686) );
  OR2_X1 U1673 ( .A1(n1687), .A2(n1688), .ZN(n1684) );
  INV_X1 U1674 ( .A(n1689), .ZN(n1688) );
  OR2_X1 U1675 ( .A1(n1690), .A2(b_0_), .ZN(n1689) );
  AND2_X1 U1676 ( .A1(b_0_), .A2(n1690), .ZN(n1687) );
  INV_X1 U1677 ( .A(a_0_), .ZN(n1690) );
  OR2_X1 U1678 ( .A1(n1691), .A2(n1692), .ZN(n1685) );
  AND2_X1 U1679 ( .A1(n1693), .A2(n1694), .ZN(n1692) );
  AND2_X1 U1680 ( .A1(n1695), .A2(n1696), .ZN(n1691) );
  OR2_X1 U1681 ( .A1(n1694), .A2(n1693), .ZN(n1695) );
  INV_X1 U1682 ( .A(n1671), .ZN(n1681) );
  OR2_X1 U1683 ( .A1(n1697), .A2(n1698), .ZN(n1671) );
  AND2_X1 U1684 ( .A1(n1655), .A2(n1661), .ZN(n1698) );
  AND2_X1 U1685 ( .A1(n1699), .A2(n1659), .ZN(n1697) );
  OR2_X1 U1686 ( .A1(n1609), .A2(n1131), .ZN(n1659) );
  AND2_X1 U1687 ( .A1(n1700), .A2(n1701), .ZN(n1131) );
  INV_X1 U1688 ( .A(n1702), .ZN(n1701) );
  AND2_X1 U1689 ( .A1(n1703), .A2(n1693), .ZN(n1702) );
  OR2_X1 U1690 ( .A1(n1703), .A2(n1693), .ZN(n1700) );
  OR2_X1 U1691 ( .A1(n1704), .A2(n1705), .ZN(n1693) );
  AND2_X1 U1692 ( .A1(n1706), .A2(n1707), .ZN(n1705) );
  AND2_X1 U1693 ( .A1(n1708), .A2(n1709), .ZN(n1704) );
  OR2_X1 U1694 ( .A1(n1707), .A2(n1706), .ZN(n1708) );
  OR2_X1 U1695 ( .A1(n1710), .A2(n1711), .ZN(n1703) );
  AND2_X1 U1696 ( .A1(a_1_), .A2(n1696), .ZN(n1711) );
  INV_X1 U1697 ( .A(b_1_), .ZN(n1696) );
  AND2_X1 U1698 ( .A1(b_1_), .A2(n1694), .ZN(n1710) );
  INV_X1 U1699 ( .A(a_1_), .ZN(n1694) );
  OR2_X1 U1700 ( .A1(n1661), .A2(n1655), .ZN(n1699) );
  OR2_X1 U1701 ( .A1(n1175), .A2(n1667), .ZN(n1655) );
  OR2_X1 U1702 ( .A1(n1712), .A2(n1713), .ZN(n1661) );
  AND2_X1 U1703 ( .A1(n1644), .A2(n1650), .ZN(n1713) );
  AND2_X1 U1704 ( .A1(n1714), .A2(n1648), .ZN(n1712) );
  OR2_X1 U1705 ( .A1(n1163), .A2(n1667), .ZN(n1648) );
  OR2_X1 U1706 ( .A1(n1650), .A2(n1644), .ZN(n1714) );
  OR2_X1 U1707 ( .A1(n1609), .A2(n1175), .ZN(n1644) );
  AND2_X1 U1708 ( .A1(n1715), .A2(n1716), .ZN(n1175) );
  INV_X1 U1709 ( .A(n1717), .ZN(n1716) );
  AND2_X1 U1710 ( .A1(n1718), .A2(n1706), .ZN(n1717) );
  OR2_X1 U1711 ( .A1(n1718), .A2(n1706), .ZN(n1715) );
  OR2_X1 U1712 ( .A1(n1719), .A2(n1720), .ZN(n1706) );
  AND2_X1 U1713 ( .A1(n1721), .A2(n1722), .ZN(n1720) );
  AND2_X1 U1714 ( .A1(n1723), .A2(n1724), .ZN(n1719) );
  OR2_X1 U1715 ( .A1(n1722), .A2(n1721), .ZN(n1723) );
  OR2_X1 U1716 ( .A1(n1725), .A2(n1726), .ZN(n1718) );
  AND2_X1 U1717 ( .A1(a_2_), .A2(n1709), .ZN(n1726) );
  INV_X1 U1718 ( .A(b_2_), .ZN(n1709) );
  AND2_X1 U1719 ( .A1(b_2_), .A2(n1707), .ZN(n1725) );
  INV_X1 U1720 ( .A(a_2_), .ZN(n1707) );
  OR2_X1 U1721 ( .A1(n1727), .A2(n1728), .ZN(n1650) );
  AND2_X1 U1722 ( .A1(n1633), .A2(n1639), .ZN(n1728) );
  AND2_X1 U1723 ( .A1(n1729), .A2(n1637), .ZN(n1727) );
  OR2_X1 U1724 ( .A1(n1609), .A2(n1163), .ZN(n1637) );
  AND2_X1 U1725 ( .A1(n1730), .A2(n1731), .ZN(n1163) );
  INV_X1 U1726 ( .A(n1732), .ZN(n1731) );
  AND2_X1 U1727 ( .A1(n1733), .A2(n1721), .ZN(n1732) );
  OR2_X1 U1728 ( .A1(n1733), .A2(n1721), .ZN(n1730) );
  OR2_X1 U1729 ( .A1(n1734), .A2(n1735), .ZN(n1721) );
  AND2_X1 U1730 ( .A1(n1736), .A2(n1737), .ZN(n1735) );
  AND2_X1 U1731 ( .A1(n1738), .A2(n1739), .ZN(n1734) );
  OR2_X1 U1732 ( .A1(n1737), .A2(n1736), .ZN(n1738) );
  OR2_X1 U1733 ( .A1(n1740), .A2(n1741), .ZN(n1733) );
  AND2_X1 U1734 ( .A1(a_3_), .A2(n1724), .ZN(n1741) );
  INV_X1 U1735 ( .A(b_3_), .ZN(n1724) );
  AND2_X1 U1736 ( .A1(b_3_), .A2(n1722), .ZN(n1740) );
  INV_X1 U1737 ( .A(a_3_), .ZN(n1722) );
  OR2_X1 U1738 ( .A1(n1639), .A2(n1633), .ZN(n1729) );
  OR2_X1 U1739 ( .A1(n1152), .A2(n1667), .ZN(n1633) );
  OR2_X1 U1740 ( .A1(n1742), .A2(n1743), .ZN(n1639) );
  AND2_X1 U1741 ( .A1(n1613), .A2(n1618), .ZN(n1743) );
  AND2_X1 U1742 ( .A1(n1619), .A2(n1744), .ZN(n1742) );
  OR2_X1 U1743 ( .A1(n1618), .A2(n1613), .ZN(n1744) );
  OR2_X1 U1744 ( .A1(n1609), .A2(n1152), .ZN(n1613) );
  AND2_X1 U1745 ( .A1(n1745), .A2(n1746), .ZN(n1152) );
  INV_X1 U1746 ( .A(n1747), .ZN(n1746) );
  AND2_X1 U1747 ( .A1(n1748), .A2(n1736), .ZN(n1747) );
  OR2_X1 U1748 ( .A1(n1748), .A2(n1736), .ZN(n1745) );
  OR2_X1 U1749 ( .A1(n1749), .A2(n1750), .ZN(n1736) );
  AND2_X1 U1750 ( .A1(n1751), .A2(n1752), .ZN(n1750) );
  AND2_X1 U1751 ( .A1(n1753), .A2(n1754), .ZN(n1749) );
  OR2_X1 U1752 ( .A1(n1751), .A2(n1752), .ZN(n1753) );
  INV_X1 U1753 ( .A(n1755), .ZN(n1751) );
  OR2_X1 U1754 ( .A1(n1756), .A2(n1757), .ZN(n1748) );
  AND2_X1 U1755 ( .A1(a_4_), .A2(n1739), .ZN(n1757) );
  INV_X1 U1756 ( .A(b_4_), .ZN(n1739) );
  AND2_X1 U1757 ( .A1(b_4_), .A2(n1737), .ZN(n1756) );
  INV_X1 U1758 ( .A(a_4_), .ZN(n1737) );
  AND2_X1 U1759 ( .A1(n1607), .A2(n1758), .ZN(n1619) );
  OR2_X1 U1760 ( .A1(n1618), .A2(n1600), .ZN(n1758) );
  OR2_X1 U1761 ( .A1(n999), .A2(n1609), .ZN(n1600) );
  INV_X1 U1762 ( .A(n1243), .ZN(n999) );
  OR2_X1 U1763 ( .A1(n1667), .A2(n1147), .ZN(n1618) );
  OR2_X1 U1764 ( .A1(n1759), .A2(n1760), .ZN(n1147) );
  AND2_X1 U1765 ( .A1(n1761), .A2(n1755), .ZN(n1760) );
  INV_X1 U1766 ( .A(n1762), .ZN(n1759) );
  OR2_X1 U1767 ( .A1(n1761), .A2(n1755), .ZN(n1762) );
  OR2_X1 U1768 ( .A1(n1763), .A2(n1764), .ZN(n1755) );
  AND2_X1 U1769 ( .A1(n1765), .A2(a_6_), .ZN(n1764) );
  AND2_X1 U1770 ( .A1(b_6_), .A2(n1766), .ZN(n1763) );
  OR2_X1 U1771 ( .A1(n1765), .A2(a_6_), .ZN(n1766) );
  OR2_X1 U1772 ( .A1(n1767), .A2(n1768), .ZN(n1761) );
  AND2_X1 U1773 ( .A1(a_5_), .A2(n1754), .ZN(n1768) );
  INV_X1 U1774 ( .A(b_5_), .ZN(n1754) );
  AND2_X1 U1775 ( .A1(b_5_), .A2(n1752), .ZN(n1767) );
  INV_X1 U1776 ( .A(a_5_), .ZN(n1752) );
  OR2_X1 U1777 ( .A1(n1499), .A2(n1769), .ZN(n1607) );
  INV_X1 U1778 ( .A(n1608), .ZN(n1769) );
  AND2_X1 U1779 ( .A1(n1243), .A2(n1599), .ZN(n1608) );
  INV_X1 U1780 ( .A(n1667), .ZN(n1599) );
  AND2_X1 U1781 ( .A1(n1770), .A2(n1771), .ZN(n1667) );
  INV_X1 U1782 ( .A(n1772), .ZN(n1771) );
  AND2_X1 U1783 ( .A1(n1773), .A2(n1774), .ZN(n1772) );
  OR2_X1 U1784 ( .A1(n1774), .A2(n1773), .ZN(n1770) );
  OR2_X1 U1785 ( .A1(n1775), .A2(n1776), .ZN(n1773) );
  INV_X1 U1786 ( .A(n1777), .ZN(n1776) );
  OR2_X1 U1787 ( .A1(n1778), .A2(d_0_), .ZN(n1777) );
  AND2_X1 U1788 ( .A1(d_0_), .A2(n1778), .ZN(n1775) );
  INV_X1 U1789 ( .A(c_0_), .ZN(n1778) );
  OR2_X1 U1790 ( .A1(n1779), .A2(n1780), .ZN(n1774) );
  AND2_X1 U1791 ( .A1(n1781), .A2(n1782), .ZN(n1780) );
  AND2_X1 U1792 ( .A1(n1783), .A2(n1784), .ZN(n1779) );
  OR2_X1 U1793 ( .A1(n1782), .A2(n1781), .ZN(n1783) );
  OR2_X1 U1794 ( .A1(n1785), .A2(n1786), .ZN(n1243) );
  AND3_X1 U1795 ( .A1(n1787), .A2(n1788), .A3(n1765), .ZN(n1786) );
  OR2_X1 U1796 ( .A1(a_6_), .A2(n1789), .ZN(n1788) );
  OR2_X1 U1797 ( .A1(b_6_), .A2(n1790), .ZN(n1787) );
  AND2_X1 U1798 ( .A1(n1791), .A2(n1792), .ZN(n1785) );
  OR2_X1 U1799 ( .A1(n1793), .A2(n1794), .ZN(n1791) );
  AND2_X1 U1800 ( .A1(a_6_), .A2(n1789), .ZN(n1794) );
  INV_X1 U1801 ( .A(b_6_), .ZN(n1789) );
  AND2_X1 U1802 ( .A1(b_6_), .A2(n1790), .ZN(n1793) );
  INV_X1 U1803 ( .A(a_6_), .ZN(n1790) );
  OR2_X1 U1804 ( .A1(n1609), .A2(n1244), .ZN(n1499) );
  INV_X1 U1805 ( .A(n998), .ZN(n1244) );
  AND2_X1 U1806 ( .A1(n1795), .A2(n1792), .ZN(n998) );
  INV_X1 U1807 ( .A(n1765), .ZN(n1792) );
  AND2_X1 U1808 ( .A1(a_7_), .A2(b_7_), .ZN(n1765) );
  OR2_X1 U1809 ( .A1(a_7_), .A2(b_7_), .ZN(n1795) );
  AND2_X1 U1810 ( .A1(n1796), .A2(n1797), .ZN(n1609) );
  INV_X1 U1811 ( .A(n1798), .ZN(n1797) );
  AND2_X1 U1812 ( .A1(n1799), .A2(n1781), .ZN(n1798) );
  OR2_X1 U1813 ( .A1(n1799), .A2(n1781), .ZN(n1796) );
  OR2_X1 U1814 ( .A1(n1800), .A2(n1801), .ZN(n1781) );
  AND2_X1 U1815 ( .A1(n1624), .A2(n1628), .ZN(n1801) );
  AND2_X1 U1816 ( .A1(n1802), .A2(n1627), .ZN(n1800) );
  INV_X1 U1817 ( .A(d_2_), .ZN(n1627) );
  OR2_X1 U1818 ( .A1(n1628), .A2(n1624), .ZN(n1802) );
  OR2_X1 U1819 ( .A1(n1803), .A2(n1804), .ZN(n1624) );
  AND2_X1 U1820 ( .A1(n1551), .A2(n1555), .ZN(n1804) );
  AND2_X1 U1821 ( .A1(n1805), .A2(n1554), .ZN(n1803) );
  INV_X1 U1822 ( .A(d_3_), .ZN(n1554) );
  OR2_X1 U1823 ( .A1(n1551), .A2(n1555), .ZN(n1805) );
  INV_X1 U1824 ( .A(c_3_), .ZN(n1555) );
  OR2_X1 U1825 ( .A1(n1806), .A2(n1807), .ZN(n1551) );
  AND2_X1 U1826 ( .A1(n1423), .A2(n1428), .ZN(n1807) );
  AND2_X1 U1827 ( .A1(n1808), .A2(n1427), .ZN(n1806) );
  INV_X1 U1828 ( .A(d_4_), .ZN(n1427) );
  OR2_X1 U1829 ( .A1(n1423), .A2(n1428), .ZN(n1808) );
  INV_X1 U1830 ( .A(c_4_), .ZN(n1428) );
  OR2_X1 U1831 ( .A1(n1809), .A2(n1810), .ZN(n1423) );
  AND2_X1 U1832 ( .A1(n1811), .A2(n1354), .ZN(n1810) );
  AND2_X1 U1833 ( .A1(n1812), .A2(n1353), .ZN(n1809) );
  INV_X1 U1834 ( .A(d_5_), .ZN(n1353) );
  OR2_X1 U1835 ( .A1(n1811), .A2(n1354), .ZN(n1812) );
  INV_X1 U1836 ( .A(c_5_), .ZN(n1354) );
  INV_X1 U1837 ( .A(n1349), .ZN(n1811) );
  OR2_X1 U1838 ( .A1(n1813), .A2(n1814), .ZN(n1349) );
  AND2_X1 U1839 ( .A1(c_6_), .A2(n1267), .ZN(n1814) );
  AND2_X1 U1840 ( .A1(d_6_), .A2(n1815), .ZN(n1813) );
  OR2_X1 U1841 ( .A1(n1267), .A2(c_6_), .ZN(n1815) );
  AND2_X1 U1842 ( .A1(c_7_), .A2(d_7_), .ZN(n1267) );
  INV_X1 U1843 ( .A(c_2_), .ZN(n1628) );
  OR2_X1 U1844 ( .A1(n1816), .A2(n1817), .ZN(n1799) );
  AND2_X1 U1845 ( .A1(c_1_), .A2(n1784), .ZN(n1817) );
  INV_X1 U1846 ( .A(d_1_), .ZN(n1784) );
  AND2_X1 U1847 ( .A1(d_1_), .A2(n1782), .ZN(n1816) );
  INV_X1 U1848 ( .A(c_1_), .ZN(n1782) );
endmodule

