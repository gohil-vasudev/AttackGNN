module add_mul_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, 
        b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, 
        b_15_, operation, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823;

  INV_X2 U1914 ( .A(operation), .ZN(n1882) );
  NOR2_X1 U1915 ( .A1(n1882), .A2(n1883), .ZN(Result_9_) );
  XOR2_X1 U1916 ( .A(n1884), .B(n1885), .Z(n1883) );
  NAND2_X1 U1917 ( .A1(n1886), .A2(n1887), .ZN(n1885) );
  NOR2_X1 U1918 ( .A1(n1882), .A2(n1888), .ZN(Result_8_) );
  XOR2_X1 U1919 ( .A(n1889), .B(n1890), .Z(n1888) );
  NAND2_X1 U1920 ( .A1(n1891), .A2(n1892), .ZN(n1890) );
  NOR2_X1 U1921 ( .A1(n1882), .A2(n1893), .ZN(Result_7_) );
  XOR2_X1 U1922 ( .A(n1894), .B(n1895), .Z(n1893) );
  NAND2_X1 U1923 ( .A1(n1896), .A2(n1897), .ZN(n1895) );
  NOR2_X1 U1924 ( .A1(n1882), .A2(n1898), .ZN(Result_6_) );
  XOR2_X1 U1925 ( .A(n1899), .B(n1900), .Z(n1898) );
  NAND2_X1 U1926 ( .A1(n1901), .A2(n1902), .ZN(n1900) );
  NOR2_X1 U1927 ( .A1(n1882), .A2(n1903), .ZN(Result_5_) );
  XOR2_X1 U1928 ( .A(n1904), .B(n1905), .Z(n1903) );
  NAND2_X1 U1929 ( .A1(n1906), .A2(n1907), .ZN(n1905) );
  NOR2_X1 U1930 ( .A1(n1882), .A2(n1908), .ZN(Result_4_) );
  XOR2_X1 U1931 ( .A(n1909), .B(n1910), .Z(n1908) );
  NAND2_X1 U1932 ( .A1(n1911), .A2(n1912), .ZN(n1910) );
  NOR2_X1 U1933 ( .A1(n1882), .A2(n1913), .ZN(Result_3_) );
  XOR2_X1 U1934 ( .A(n1914), .B(n1915), .Z(n1913) );
  NAND2_X1 U1935 ( .A1(n1916), .A2(n1917), .ZN(n1915) );
  NAND2_X1 U1936 ( .A1(n1918), .A2(n1919), .ZN(Result_31_) );
  NAND2_X1 U1937 ( .A1(n1920), .A2(n1882), .ZN(n1919) );
  XNOR2_X1 U1938 ( .A(n1921), .B(a_15_), .ZN(n1920) );
  OR2_X1 U1939 ( .A1(n1922), .A2(n1882), .ZN(n1918) );
  NAND2_X1 U1940 ( .A1(n1923), .A2(n1924), .ZN(Result_30_) );
  NAND2_X1 U1941 ( .A1(operation), .A2(n1925), .ZN(n1924) );
  NAND2_X1 U1942 ( .A1(n1926), .A2(n1927), .ZN(n1925) );
  NAND2_X1 U1943 ( .A1(b_14_), .A2(n1928), .ZN(n1927) );
  NAND2_X1 U1944 ( .A1(n1929), .A2(n1930), .ZN(n1928) );
  NAND2_X1 U1945 ( .A1(a_15_), .A2(n1921), .ZN(n1930) );
  NAND2_X1 U1946 ( .A1(b_15_), .A2(n1931), .ZN(n1926) );
  NAND2_X1 U1947 ( .A1(n1932), .A2(n1933), .ZN(n1931) );
  NAND2_X1 U1948 ( .A1(a_14_), .A2(n1934), .ZN(n1933) );
  NAND2_X1 U1949 ( .A1(n1935), .A2(n1882), .ZN(n1923) );
  XNOR2_X1 U1950 ( .A(n1922), .B(n1936), .ZN(n1935) );
  XNOR2_X1 U1951 ( .A(n1934), .B(a_14_), .ZN(n1936) );
  NOR2_X1 U1952 ( .A1(n1882), .A2(n1937), .ZN(Result_2_) );
  XOR2_X1 U1953 ( .A(n1938), .B(n1939), .Z(n1937) );
  NAND2_X1 U1954 ( .A1(n1940), .A2(n1941), .ZN(n1939) );
  NAND2_X1 U1955 ( .A1(n1942), .A2(n1943), .ZN(Result_29_) );
  NAND2_X1 U1956 ( .A1(n1944), .A2(n1882), .ZN(n1943) );
  NAND3_X1 U1957 ( .A1(n1945), .A2(n1946), .A3(n1947), .ZN(n1944) );
  NAND2_X1 U1958 ( .A1(n1948), .A2(n1949), .ZN(n1947) );
  OR3_X1 U1959 ( .A1(n1949), .A2(a_13_), .A3(n1950), .ZN(n1946) );
  NAND2_X1 U1960 ( .A1(n1951), .A2(n1950), .ZN(n1945) );
  XNOR2_X1 U1961 ( .A(n1949), .B(n1952), .ZN(n1951) );
  NAND2_X1 U1962 ( .A1(n1953), .A2(operation), .ZN(n1942) );
  XOR2_X1 U1963 ( .A(n1954), .B(n1955), .Z(n1953) );
  NOR2_X1 U1964 ( .A1(n1952), .A2(n1921), .ZN(n1955) );
  XOR2_X1 U1965 ( .A(n1956), .B(n1957), .Z(n1954) );
  NAND2_X1 U1966 ( .A1(n1958), .A2(n1959), .ZN(Result_28_) );
  NAND2_X1 U1967 ( .A1(n1960), .A2(n1882), .ZN(n1959) );
  XOR2_X1 U1968 ( .A(n1961), .B(n1962), .Z(n1960) );
  AND2_X1 U1969 ( .A1(n1963), .A2(n1964), .ZN(n1962) );
  NAND2_X1 U1970 ( .A1(n1965), .A2(operation), .ZN(n1958) );
  XOR2_X1 U1971 ( .A(n1966), .B(n1967), .Z(n1965) );
  XOR2_X1 U1972 ( .A(n1968), .B(n1969), .Z(n1967) );
  NOR2_X1 U1973 ( .A1(n1970), .A2(n1921), .ZN(n1969) );
  NAND2_X1 U1974 ( .A1(n1971), .A2(n1972), .ZN(Result_27_) );
  NAND2_X1 U1975 ( .A1(n1973), .A2(n1882), .ZN(n1972) );
  NAND3_X1 U1976 ( .A1(n1974), .A2(n1975), .A3(n1976), .ZN(n1973) );
  NAND2_X1 U1977 ( .A1(n1977), .A2(n1978), .ZN(n1976) );
  OR3_X1 U1978 ( .A1(n1978), .A2(a_11_), .A3(n1979), .ZN(n1975) );
  NAND2_X1 U1979 ( .A1(n1980), .A2(n1979), .ZN(n1974) );
  XNOR2_X1 U1980 ( .A(n1978), .B(n1981), .ZN(n1980) );
  NAND2_X1 U1981 ( .A1(n1982), .A2(operation), .ZN(n1971) );
  XNOR2_X1 U1982 ( .A(n1983), .B(n1984), .ZN(n1982) );
  NAND2_X1 U1983 ( .A1(n1985), .A2(n1986), .ZN(n1983) );
  NAND2_X1 U1984 ( .A1(n1987), .A2(n1988), .ZN(Result_26_) );
  NAND2_X1 U1985 ( .A1(n1989), .A2(n1882), .ZN(n1988) );
  XNOR2_X1 U1986 ( .A(n1990), .B(n1991), .ZN(n1989) );
  NOR2_X1 U1987 ( .A1(n1992), .A2(n1993), .ZN(n1991) );
  NAND2_X1 U1988 ( .A1(n1994), .A2(operation), .ZN(n1987) );
  XNOR2_X1 U1989 ( .A(n1995), .B(n1996), .ZN(n1994) );
  XOR2_X1 U1990 ( .A(n1997), .B(n1998), .Z(n1996) );
  NAND2_X1 U1991 ( .A1(b_15_), .A2(a_10_), .ZN(n1998) );
  NAND2_X1 U1992 ( .A1(n1999), .A2(n2000), .ZN(Result_25_) );
  NAND2_X1 U1993 ( .A1(n2001), .A2(n1882), .ZN(n2000) );
  NAND3_X1 U1994 ( .A1(n2002), .A2(n2003), .A3(n2004), .ZN(n2001) );
  NAND2_X1 U1995 ( .A1(n2005), .A2(n2006), .ZN(n2004) );
  NAND3_X1 U1996 ( .A1(n2007), .A2(n2008), .A3(b_9_), .ZN(n2003) );
  NAND2_X1 U1997 ( .A1(n2009), .A2(n2010), .ZN(n2002) );
  XNOR2_X1 U1998 ( .A(n2007), .B(a_9_), .ZN(n2009) );
  NAND2_X1 U1999 ( .A1(n2011), .A2(operation), .ZN(n1999) );
  XNOR2_X1 U2000 ( .A(n2012), .B(n2013), .ZN(n2011) );
  NAND2_X1 U2001 ( .A1(n2014), .A2(n2015), .ZN(n2012) );
  NAND2_X1 U2002 ( .A1(n2016), .A2(n2017), .ZN(Result_24_) );
  NAND2_X1 U2003 ( .A1(n2018), .A2(n1882), .ZN(n2017) );
  XOR2_X1 U2004 ( .A(n2019), .B(n2020), .Z(n2018) );
  AND2_X1 U2005 ( .A1(n2021), .A2(n2022), .ZN(n2020) );
  NAND2_X1 U2006 ( .A1(n2023), .A2(operation), .ZN(n2016) );
  XOR2_X1 U2007 ( .A(n2024), .B(n2025), .Z(n2023) );
  XNOR2_X1 U2008 ( .A(n2026), .B(n2027), .ZN(n2025) );
  NAND2_X1 U2009 ( .A1(b_15_), .A2(a_8_), .ZN(n2026) );
  NAND2_X1 U2010 ( .A1(n2028), .A2(n2029), .ZN(Result_23_) );
  NAND2_X1 U2011 ( .A1(n2030), .A2(n1882), .ZN(n2029) );
  NAND3_X1 U2012 ( .A1(n2031), .A2(n2032), .A3(n2033), .ZN(n2030) );
  NAND2_X1 U2013 ( .A1(n2034), .A2(n2035), .ZN(n2033) );
  OR3_X1 U2014 ( .A1(n2035), .A2(a_7_), .A3(n2036), .ZN(n2032) );
  NAND2_X1 U2015 ( .A1(n2037), .A2(n2036), .ZN(n2031) );
  XNOR2_X1 U2016 ( .A(n2035), .B(n2038), .ZN(n2037) );
  NAND2_X1 U2017 ( .A1(n2039), .A2(operation), .ZN(n2028) );
  XNOR2_X1 U2018 ( .A(n2040), .B(n2041), .ZN(n2039) );
  NAND2_X1 U2019 ( .A1(n2042), .A2(n2043), .ZN(n2040) );
  NAND2_X1 U2020 ( .A1(n2044), .A2(n2045), .ZN(Result_22_) );
  NAND2_X1 U2021 ( .A1(n2046), .A2(n1882), .ZN(n2045) );
  XNOR2_X1 U2022 ( .A(n2047), .B(n2048), .ZN(n2046) );
  NOR2_X1 U2023 ( .A1(n2049), .A2(n2050), .ZN(n2048) );
  NAND2_X1 U2024 ( .A1(n2051), .A2(operation), .ZN(n2044) );
  XOR2_X1 U2025 ( .A(n2052), .B(n2053), .Z(n2051) );
  XOR2_X1 U2026 ( .A(n2054), .B(n2055), .Z(n2053) );
  NOR2_X1 U2027 ( .A1(n2056), .A2(n1921), .ZN(n2055) );
  INV_X1 U2028 ( .A(b_15_), .ZN(n1921) );
  NAND2_X1 U2029 ( .A1(n2057), .A2(n2058), .ZN(Result_21_) );
  NAND2_X1 U2030 ( .A1(n2059), .A2(n1882), .ZN(n2058) );
  NAND3_X1 U2031 ( .A1(n2060), .A2(n2061), .A3(n2062), .ZN(n2059) );
  NAND2_X1 U2032 ( .A1(n2063), .A2(n2064), .ZN(n2062) );
  NAND3_X1 U2033 ( .A1(n2065), .A2(n2066), .A3(b_5_), .ZN(n2061) );
  NAND2_X1 U2034 ( .A1(n2067), .A2(n2068), .ZN(n2060) );
  XNOR2_X1 U2035 ( .A(n2065), .B(a_5_), .ZN(n2067) );
  NAND2_X1 U2036 ( .A1(n2069), .A2(operation), .ZN(n2057) );
  XOR2_X1 U2037 ( .A(n2070), .B(n2071), .Z(n2069) );
  XNOR2_X1 U2038 ( .A(n2072), .B(n2073), .ZN(n2071) );
  NAND2_X1 U2039 ( .A1(b_15_), .A2(a_5_), .ZN(n2073) );
  NAND2_X1 U2040 ( .A1(n2074), .A2(n2075), .ZN(Result_20_) );
  NAND2_X1 U2041 ( .A1(n2076), .A2(n1882), .ZN(n2075) );
  XNOR2_X1 U2042 ( .A(n2077), .B(n2078), .ZN(n2076) );
  NOR2_X1 U2043 ( .A1(n2079), .A2(n2080), .ZN(n2078) );
  NAND2_X1 U2044 ( .A1(n2081), .A2(operation), .ZN(n2074) );
  XOR2_X1 U2045 ( .A(n2082), .B(n2083), .Z(n2081) );
  XNOR2_X1 U2046 ( .A(n2084), .B(n2085), .ZN(n2083) );
  NAND2_X1 U2047 ( .A1(b_15_), .A2(a_4_), .ZN(n2085) );
  NOR2_X1 U2048 ( .A1(n1882), .A2(n2086), .ZN(Result_1_) );
  XOR2_X1 U2049 ( .A(n2087), .B(n2088), .Z(n2086) );
  NAND2_X1 U2050 ( .A1(n2089), .A2(n2090), .ZN(n2088) );
  NAND2_X1 U2051 ( .A1(n2091), .A2(n2092), .ZN(Result_19_) );
  NAND2_X1 U2052 ( .A1(n2093), .A2(n1882), .ZN(n2092) );
  NAND3_X1 U2053 ( .A1(n2094), .A2(n2095), .A3(n2096), .ZN(n2093) );
  NAND2_X1 U2054 ( .A1(n2097), .A2(n2098), .ZN(n2096) );
  NAND3_X1 U2055 ( .A1(n2099), .A2(n2100), .A3(b_3_), .ZN(n2095) );
  NAND2_X1 U2056 ( .A1(n2101), .A2(n2102), .ZN(n2094) );
  XNOR2_X1 U2057 ( .A(n2099), .B(a_3_), .ZN(n2101) );
  NAND2_X1 U2058 ( .A1(n2103), .A2(operation), .ZN(n2091) );
  XNOR2_X1 U2059 ( .A(n2104), .B(n2105), .ZN(n2103) );
  XOR2_X1 U2060 ( .A(n2106), .B(n2107), .Z(n2105) );
  NAND2_X1 U2061 ( .A1(b_15_), .A2(a_3_), .ZN(n2107) );
  NAND2_X1 U2062 ( .A1(n2108), .A2(n2109), .ZN(Result_18_) );
  NAND2_X1 U2063 ( .A1(n2110), .A2(n1882), .ZN(n2109) );
  XOR2_X1 U2064 ( .A(n2111), .B(n2112), .Z(n2110) );
  AND2_X1 U2065 ( .A1(n2113), .A2(n2114), .ZN(n2112) );
  NAND2_X1 U2066 ( .A1(n2115), .A2(operation), .ZN(n2108) );
  XOR2_X1 U2067 ( .A(n2116), .B(n2117), .Z(n2115) );
  XNOR2_X1 U2068 ( .A(n2118), .B(n2119), .ZN(n2117) );
  NAND2_X1 U2069 ( .A1(b_15_), .A2(a_2_), .ZN(n2119) );
  NAND2_X1 U2070 ( .A1(n2120), .A2(n2121), .ZN(Result_17_) );
  NAND2_X1 U2071 ( .A1(n2122), .A2(n1882), .ZN(n2121) );
  NAND2_X1 U2072 ( .A1(n2123), .A2(n2124), .ZN(n2122) );
  NAND2_X1 U2073 ( .A1(n2125), .A2(n2126), .ZN(n2124) );
  OR2_X1 U2074 ( .A1(n2127), .A2(n2128), .ZN(n2125) );
  NAND2_X1 U2075 ( .A1(n2129), .A2(n2130), .ZN(n2123) );
  INV_X1 U2076 ( .A(n2126), .ZN(n2130) );
  XNOR2_X1 U2077 ( .A(n2131), .B(a_1_), .ZN(n2129) );
  NAND2_X1 U2078 ( .A1(n2132), .A2(operation), .ZN(n2120) );
  XOR2_X1 U2079 ( .A(n2133), .B(n2134), .Z(n2132) );
  XNOR2_X1 U2080 ( .A(n2135), .B(n2136), .ZN(n2134) );
  NAND2_X1 U2081 ( .A1(b_15_), .A2(a_1_), .ZN(n2136) );
  NAND2_X1 U2082 ( .A1(n2137), .A2(n2138), .ZN(Result_16_) );
  NAND2_X1 U2083 ( .A1(n2139), .A2(n1882), .ZN(n2138) );
  XOR2_X1 U2084 ( .A(n2140), .B(n2141), .Z(n2139) );
  NOR2_X1 U2085 ( .A1(n2142), .A2(n2143), .ZN(n2141) );
  NOR2_X1 U2086 ( .A1(b_0_), .A2(a_0_), .ZN(n2142) );
  NOR2_X1 U2087 ( .A1(n2128), .A2(n2144), .ZN(n2140) );
  NOR2_X1 U2088 ( .A1(n2127), .A2(n2126), .ZN(n2144) );
  NAND2_X1 U2089 ( .A1(n2114), .A2(n2145), .ZN(n2126) );
  NAND2_X1 U2090 ( .A1(n2113), .A2(n2111), .ZN(n2145) );
  NAND2_X1 U2091 ( .A1(n2146), .A2(n2147), .ZN(n2111) );
  NAND2_X1 U2092 ( .A1(n2148), .A2(n2098), .ZN(n2147) );
  INV_X1 U2093 ( .A(n2099), .ZN(n2098) );
  NOR2_X1 U2094 ( .A1(n2080), .A2(n2149), .ZN(n2099) );
  NOR2_X1 U2095 ( .A1(n2079), .A2(n2077), .ZN(n2149) );
  AND2_X1 U2096 ( .A1(n2150), .A2(n2151), .ZN(n2077) );
  NAND2_X1 U2097 ( .A1(n2152), .A2(n2064), .ZN(n2151) );
  INV_X1 U2098 ( .A(n2065), .ZN(n2064) );
  NOR2_X1 U2099 ( .A1(n2050), .A2(n2153), .ZN(n2065) );
  NOR2_X1 U2100 ( .A1(n2049), .A2(n2047), .ZN(n2153) );
  AND2_X1 U2101 ( .A1(n2154), .A2(n2155), .ZN(n2047) );
  NAND2_X1 U2102 ( .A1(n2156), .A2(n2035), .ZN(n2155) );
  NAND2_X1 U2103 ( .A1(n2022), .A2(n2157), .ZN(n2035) );
  NAND2_X1 U2104 ( .A1(n2021), .A2(n2019), .ZN(n2157) );
  NAND2_X1 U2105 ( .A1(n2158), .A2(n2159), .ZN(n2019) );
  NAND2_X1 U2106 ( .A1(n2160), .A2(n2006), .ZN(n2159) );
  INV_X1 U2107 ( .A(n2007), .ZN(n2006) );
  NOR2_X1 U2108 ( .A1(n1993), .A2(n2161), .ZN(n2007) );
  NOR2_X1 U2109 ( .A1(n1992), .A2(n1990), .ZN(n2161) );
  AND2_X1 U2110 ( .A1(n2162), .A2(n2163), .ZN(n1990) );
  NAND2_X1 U2111 ( .A1(n2164), .A2(n1978), .ZN(n2163) );
  NAND2_X1 U2112 ( .A1(n1964), .A2(n2165), .ZN(n1978) );
  NAND2_X1 U2113 ( .A1(n1963), .A2(n1961), .ZN(n2165) );
  NAND2_X1 U2114 ( .A1(n2166), .A2(n2167), .ZN(n1961) );
  NAND2_X1 U2115 ( .A1(n2168), .A2(n1949), .ZN(n2167) );
  NAND2_X1 U2116 ( .A1(n2169), .A2(n2170), .ZN(n1949) );
  NAND2_X1 U2117 ( .A1(b_14_), .A2(n2171), .ZN(n2170) );
  NAND2_X1 U2118 ( .A1(n2172), .A2(n1922), .ZN(n2171) );
  NAND2_X1 U2119 ( .A1(b_15_), .A2(a_15_), .ZN(n1922) );
  NAND2_X1 U2120 ( .A1(b_15_), .A2(n2173), .ZN(n2169) );
  NAND2_X1 U2121 ( .A1(n1950), .A2(n1952), .ZN(n2168) );
  NAND2_X1 U2122 ( .A1(n2174), .A2(n1970), .ZN(n1963) );
  NAND2_X1 U2123 ( .A1(n1979), .A2(n1981), .ZN(n2164) );
  NOR2_X1 U2124 ( .A1(b_10_), .A2(a_10_), .ZN(n1992) );
  NAND2_X1 U2125 ( .A1(n2010), .A2(n2008), .ZN(n2160) );
  NAND2_X1 U2126 ( .A1(n2175), .A2(n2176), .ZN(n2021) );
  NAND2_X1 U2127 ( .A1(n2036), .A2(n2038), .ZN(n2156) );
  NOR2_X1 U2128 ( .A1(b_6_), .A2(a_6_), .ZN(n2049) );
  NAND2_X1 U2129 ( .A1(n2068), .A2(n2066), .ZN(n2152) );
  NOR2_X1 U2130 ( .A1(b_4_), .A2(a_4_), .ZN(n2079) );
  NAND2_X1 U2131 ( .A1(n2102), .A2(n2100), .ZN(n2148) );
  NAND2_X1 U2132 ( .A1(n2177), .A2(n2178), .ZN(n2113) );
  NOR2_X1 U2133 ( .A1(b_1_), .A2(a_1_), .ZN(n2128) );
  NAND2_X1 U2134 ( .A1(n2179), .A2(operation), .ZN(n2137) );
  XOR2_X1 U2135 ( .A(n2180), .B(n2181), .Z(n2179) );
  XNOR2_X1 U2136 ( .A(n2182), .B(n2183), .ZN(n2181) );
  NAND2_X1 U2137 ( .A1(b_15_), .A2(a_0_), .ZN(n2183) );
  NOR2_X1 U2138 ( .A1(n2184), .A2(n1882), .ZN(Result_15_) );
  XNOR2_X1 U2139 ( .A(n2185), .B(n2186), .ZN(n2184) );
  NOR3_X1 U2140 ( .A1(n1882), .A2(n2187), .A3(n2188), .ZN(Result_14_) );
  NOR2_X1 U2141 ( .A1(n2189), .A2(n2190), .ZN(n2188) );
  AND2_X1 U2142 ( .A1(n2186), .A2(n2185), .ZN(n2189) );
  NOR2_X1 U2143 ( .A1(n2191), .A2(n1882), .ZN(Result_13_) );
  XOR2_X1 U2144 ( .A(n2192), .B(n2187), .Z(n2191) );
  NAND2_X1 U2145 ( .A1(n2193), .A2(n2194), .ZN(n2192) );
  NAND2_X1 U2146 ( .A1(n2195), .A2(n2196), .ZN(n2193) );
  NAND2_X1 U2147 ( .A1(n2197), .A2(n2198), .ZN(n2196) );
  NOR2_X1 U2148 ( .A1(n2199), .A2(n1882), .ZN(Result_12_) );
  XNOR2_X1 U2149 ( .A(n2200), .B(n2201), .ZN(n2199) );
  NOR2_X1 U2150 ( .A1(n2202), .A2(n1882), .ZN(Result_11_) );
  XOR2_X1 U2151 ( .A(n2203), .B(n2204), .Z(n2202) );
  NAND2_X1 U2152 ( .A1(n2205), .A2(n2206), .ZN(n2203) );
  NAND2_X1 U2153 ( .A1(n2207), .A2(n2208), .ZN(n2205) );
  NOR2_X1 U2154 ( .A1(n1882), .A2(n2209), .ZN(Result_10_) );
  XOR2_X1 U2155 ( .A(n2210), .B(n2211), .Z(n2209) );
  NAND2_X1 U2156 ( .A1(n2212), .A2(n2213), .ZN(n2211) );
  NOR2_X1 U2157 ( .A1(n2214), .A2(n1882), .ZN(Result_0_) );
  NOR3_X1 U2158 ( .A1(n2215), .A2(n2216), .A3(n2217), .ZN(n2214) );
  AND2_X1 U2159 ( .A1(n2087), .A2(n2089), .ZN(n2217) );
  NAND2_X1 U2160 ( .A1(n2218), .A2(n2219), .ZN(n2089) );
  NAND2_X1 U2161 ( .A1(n2220), .A2(n2221), .ZN(n2219) );
  XOR2_X1 U2162 ( .A(n2143), .B(n2222), .Z(n2218) );
  NAND2_X1 U2163 ( .A1(n1940), .A2(n2223), .ZN(n2087) );
  NAND2_X1 U2164 ( .A1(n1941), .A2(n1938), .ZN(n2223) );
  NAND2_X1 U2165 ( .A1(n1916), .A2(n2224), .ZN(n1938) );
  NAND2_X1 U2166 ( .A1(n1917), .A2(n1914), .ZN(n2224) );
  NAND2_X1 U2167 ( .A1(n1911), .A2(n2225), .ZN(n1914) );
  NAND2_X1 U2168 ( .A1(n1912), .A2(n1909), .ZN(n2225) );
  NAND2_X1 U2169 ( .A1(n1906), .A2(n2226), .ZN(n1909) );
  NAND2_X1 U2170 ( .A1(n1907), .A2(n1904), .ZN(n2226) );
  NAND2_X1 U2171 ( .A1(n1901), .A2(n2227), .ZN(n1904) );
  NAND2_X1 U2172 ( .A1(n1902), .A2(n1899), .ZN(n2227) );
  NAND2_X1 U2173 ( .A1(n1896), .A2(n2228), .ZN(n1899) );
  NAND2_X1 U2174 ( .A1(n1897), .A2(n1894), .ZN(n2228) );
  NAND2_X1 U2175 ( .A1(n1891), .A2(n2229), .ZN(n1894) );
  NAND2_X1 U2176 ( .A1(n1892), .A2(n1889), .ZN(n2229) );
  NAND2_X1 U2177 ( .A1(n1886), .A2(n2230), .ZN(n1889) );
  NAND2_X1 U2178 ( .A1(n1887), .A2(n1884), .ZN(n2230) );
  NAND2_X1 U2179 ( .A1(n2231), .A2(n2212), .ZN(n1884) );
  NAND2_X1 U2180 ( .A1(n2232), .A2(n2233), .ZN(n2212) );
  NAND2_X1 U2181 ( .A1(n2210), .A2(n2213), .ZN(n2231) );
  OR2_X1 U2182 ( .A1(n2233), .A2(n2232), .ZN(n2213) );
  XOR2_X1 U2183 ( .A(n2234), .B(n2235), .Z(n2233) );
  NAND2_X1 U2184 ( .A1(n2236), .A2(n2206), .ZN(n2210) );
  OR2_X1 U2185 ( .A1(n2207), .A2(n2208), .ZN(n2206) );
  NAND2_X1 U2186 ( .A1(n2237), .A2(n2238), .ZN(n2208) );
  INV_X1 U2187 ( .A(n2239), .ZN(n2207) );
  NAND2_X1 U2188 ( .A1(n2204), .A2(n2239), .ZN(n2236) );
  NOR2_X1 U2189 ( .A1(n2232), .A2(n2240), .ZN(n2239) );
  AND2_X1 U2190 ( .A1(n2241), .A2(n2242), .ZN(n2240) );
  NOR2_X1 U2191 ( .A1(n2242), .A2(n2241), .ZN(n2232) );
  XOR2_X1 U2192 ( .A(n2243), .B(n2244), .Z(n2241) );
  NAND2_X1 U2193 ( .A1(n2245), .A2(n2246), .ZN(n2243) );
  NAND2_X1 U2194 ( .A1(n2247), .A2(n2248), .ZN(n2242) );
  NAND2_X1 U2195 ( .A1(n2249), .A2(n2250), .ZN(n2248) );
  NAND2_X1 U2196 ( .A1(n2251), .A2(n2252), .ZN(n2250) );
  OR2_X1 U2197 ( .A1(n2252), .A2(n2251), .ZN(n2247) );
  AND2_X1 U2198 ( .A1(n2200), .A2(n2201), .ZN(n2204) );
  NAND3_X1 U2199 ( .A1(n2253), .A2(n2194), .A3(n2254), .ZN(n2201) );
  NAND2_X1 U2200 ( .A1(n2187), .A2(n2255), .ZN(n2254) );
  AND3_X1 U2201 ( .A1(n2185), .A2(n2186), .A3(n2190), .ZN(n2187) );
  XOR2_X1 U2202 ( .A(n2198), .B(n2197), .Z(n2190) );
  NAND2_X1 U2203 ( .A1(n2256), .A2(n2257), .ZN(n2186) );
  NAND3_X1 U2204 ( .A1(a_0_), .A2(n2258), .A3(b_15_), .ZN(n2257) );
  NAND2_X1 U2205 ( .A1(n2182), .A2(n2180), .ZN(n2258) );
  OR2_X1 U2206 ( .A1(n2180), .A2(n2182), .ZN(n2256) );
  AND2_X1 U2207 ( .A1(n2259), .A2(n2260), .ZN(n2182) );
  NAND3_X1 U2208 ( .A1(a_1_), .A2(n2261), .A3(b_15_), .ZN(n2260) );
  NAND2_X1 U2209 ( .A1(n2135), .A2(n2133), .ZN(n2261) );
  OR2_X1 U2210 ( .A1(n2133), .A2(n2135), .ZN(n2259) );
  AND2_X1 U2211 ( .A1(n2262), .A2(n2263), .ZN(n2135) );
  NAND3_X1 U2212 ( .A1(a_2_), .A2(n2264), .A3(b_15_), .ZN(n2263) );
  NAND2_X1 U2213 ( .A1(n2118), .A2(n2116), .ZN(n2264) );
  OR2_X1 U2214 ( .A1(n2116), .A2(n2118), .ZN(n2262) );
  AND2_X1 U2215 ( .A1(n2265), .A2(n2266), .ZN(n2118) );
  NAND3_X1 U2216 ( .A1(a_3_), .A2(n2267), .A3(b_15_), .ZN(n2266) );
  OR2_X1 U2217 ( .A1(n2106), .A2(n2104), .ZN(n2267) );
  NAND2_X1 U2218 ( .A1(n2104), .A2(n2106), .ZN(n2265) );
  NAND2_X1 U2219 ( .A1(n2268), .A2(n2269), .ZN(n2106) );
  NAND3_X1 U2220 ( .A1(a_4_), .A2(n2270), .A3(b_15_), .ZN(n2269) );
  NAND2_X1 U2221 ( .A1(n2084), .A2(n2082), .ZN(n2270) );
  OR2_X1 U2222 ( .A1(n2082), .A2(n2084), .ZN(n2268) );
  AND2_X1 U2223 ( .A1(n2271), .A2(n2272), .ZN(n2084) );
  NAND3_X1 U2224 ( .A1(a_5_), .A2(n2273), .A3(b_15_), .ZN(n2272) );
  NAND2_X1 U2225 ( .A1(n2072), .A2(n2070), .ZN(n2273) );
  OR2_X1 U2226 ( .A1(n2070), .A2(n2072), .ZN(n2271) );
  AND2_X1 U2227 ( .A1(n2274), .A2(n2275), .ZN(n2072) );
  NAND3_X1 U2228 ( .A1(a_6_), .A2(n2276), .A3(b_15_), .ZN(n2275) );
  NAND2_X1 U2229 ( .A1(n2054), .A2(n2052), .ZN(n2276) );
  OR2_X1 U2230 ( .A1(n2052), .A2(n2054), .ZN(n2274) );
  AND2_X1 U2231 ( .A1(n2042), .A2(n2277), .ZN(n2054) );
  NAND2_X1 U2232 ( .A1(n2041), .A2(n2043), .ZN(n2277) );
  NAND2_X1 U2233 ( .A1(n2278), .A2(n2279), .ZN(n2043) );
  NAND2_X1 U2234 ( .A1(b_15_), .A2(a_7_), .ZN(n2279) );
  INV_X1 U2235 ( .A(n2280), .ZN(n2278) );
  XOR2_X1 U2236 ( .A(n2281), .B(n2282), .Z(n2041) );
  XNOR2_X1 U2237 ( .A(n2283), .B(n2284), .ZN(n2281) );
  NAND2_X1 U2238 ( .A1(b_14_), .A2(a_8_), .ZN(n2283) );
  NAND2_X1 U2239 ( .A1(a_7_), .A2(n2280), .ZN(n2042) );
  NAND2_X1 U2240 ( .A1(n2285), .A2(n2286), .ZN(n2280) );
  NAND3_X1 U2241 ( .A1(a_8_), .A2(n2287), .A3(b_15_), .ZN(n2286) );
  OR2_X1 U2242 ( .A1(n2027), .A2(n2024), .ZN(n2287) );
  NAND2_X1 U2243 ( .A1(n2024), .A2(n2027), .ZN(n2285) );
  NAND2_X1 U2244 ( .A1(n2014), .A2(n2288), .ZN(n2027) );
  NAND2_X1 U2245 ( .A1(n2013), .A2(n2015), .ZN(n2288) );
  NAND2_X1 U2246 ( .A1(n2289), .A2(n2290), .ZN(n2015) );
  NAND2_X1 U2247 ( .A1(b_15_), .A2(a_9_), .ZN(n2290) );
  INV_X1 U2248 ( .A(n2291), .ZN(n2289) );
  XNOR2_X1 U2249 ( .A(n2292), .B(n2293), .ZN(n2013) );
  NAND2_X1 U2250 ( .A1(n2294), .A2(n2295), .ZN(n2292) );
  NAND2_X1 U2251 ( .A1(a_9_), .A2(n2291), .ZN(n2014) );
  NAND2_X1 U2252 ( .A1(n2296), .A2(n2297), .ZN(n2291) );
  NAND3_X1 U2253 ( .A1(a_10_), .A2(n2298), .A3(b_15_), .ZN(n2297) );
  OR2_X1 U2254 ( .A1(n1997), .A2(n1995), .ZN(n2298) );
  NAND2_X1 U2255 ( .A1(n1995), .A2(n1997), .ZN(n2296) );
  NAND2_X1 U2256 ( .A1(n1985), .A2(n2299), .ZN(n1997) );
  NAND2_X1 U2257 ( .A1(n1984), .A2(n1986), .ZN(n2299) );
  NAND2_X1 U2258 ( .A1(n2300), .A2(n2301), .ZN(n1986) );
  NAND2_X1 U2259 ( .A1(b_15_), .A2(a_11_), .ZN(n2301) );
  INV_X1 U2260 ( .A(n2302), .ZN(n2300) );
  XNOR2_X1 U2261 ( .A(n2303), .B(n2304), .ZN(n1984) );
  XOR2_X1 U2262 ( .A(n2305), .B(n2306), .Z(n2303) );
  NAND2_X1 U2263 ( .A1(b_14_), .A2(a_12_), .ZN(n2305) );
  NAND2_X1 U2264 ( .A1(a_11_), .A2(n2302), .ZN(n1985) );
  NAND2_X1 U2265 ( .A1(n2307), .A2(n2308), .ZN(n2302) );
  NAND3_X1 U2266 ( .A1(a_12_), .A2(n2309), .A3(b_15_), .ZN(n2308) );
  NAND2_X1 U2267 ( .A1(n1968), .A2(n1966), .ZN(n2309) );
  OR2_X1 U2268 ( .A1(n1966), .A2(n1968), .ZN(n2307) );
  AND2_X1 U2269 ( .A1(n2310), .A2(n2311), .ZN(n1968) );
  NAND3_X1 U2270 ( .A1(a_13_), .A2(n2312), .A3(b_15_), .ZN(n2311) );
  OR2_X1 U2271 ( .A1(n1956), .A2(n1957), .ZN(n2312) );
  NAND2_X1 U2272 ( .A1(n1957), .A2(n1956), .ZN(n2310) );
  NAND2_X1 U2273 ( .A1(n2313), .A2(n2314), .ZN(n1956) );
  NAND2_X1 U2274 ( .A1(b_13_), .A2(n2315), .ZN(n2314) );
  NAND2_X1 U2275 ( .A1(n1929), .A2(n2316), .ZN(n2315) );
  NAND2_X1 U2276 ( .A1(a_15_), .A2(n1934), .ZN(n2316) );
  NAND2_X1 U2277 ( .A1(b_14_), .A2(n2317), .ZN(n2313) );
  NAND2_X1 U2278 ( .A1(n1932), .A2(n2318), .ZN(n2317) );
  NAND2_X1 U2279 ( .A1(a_14_), .A2(n1950), .ZN(n2318) );
  AND3_X1 U2280 ( .A1(b_14_), .A2(n2173), .A3(b_15_), .ZN(n1957) );
  XNOR2_X1 U2281 ( .A(n2319), .B(n2320), .ZN(n1966) );
  XOR2_X1 U2282 ( .A(n2321), .B(n2322), .Z(n2319) );
  XNOR2_X1 U2283 ( .A(n2323), .B(n2324), .ZN(n1995) );
  NAND2_X1 U2284 ( .A1(n2325), .A2(n2326), .ZN(n2323) );
  XOR2_X1 U2285 ( .A(n2327), .B(n2328), .Z(n2024) );
  XOR2_X1 U2286 ( .A(n2329), .B(n2330), .Z(n2327) );
  XOR2_X1 U2287 ( .A(n2331), .B(n2332), .Z(n2052) );
  XNOR2_X1 U2288 ( .A(n2333), .B(n2334), .ZN(n2332) );
  XNOR2_X1 U2289 ( .A(n2335), .B(n2336), .ZN(n2070) );
  XOR2_X1 U2290 ( .A(n2337), .B(n2338), .Z(n2335) );
  NOR2_X1 U2291 ( .A1(n2056), .A2(n1934), .ZN(n2338) );
  XNOR2_X1 U2292 ( .A(n2339), .B(n2340), .ZN(n2082) );
  XOR2_X1 U2293 ( .A(n2341), .B(n2342), .Z(n2339) );
  XNOR2_X1 U2294 ( .A(n2343), .B(n2344), .ZN(n2104) );
  XNOR2_X1 U2295 ( .A(n2345), .B(n2346), .ZN(n2343) );
  NOR2_X1 U2296 ( .A1(n2347), .A2(n1934), .ZN(n2346) );
  XOR2_X1 U2297 ( .A(n2348), .B(n2349), .Z(n2116) );
  XNOR2_X1 U2298 ( .A(n2350), .B(n2351), .ZN(n2349) );
  XOR2_X1 U2299 ( .A(n2352), .B(n2353), .Z(n2133) );
  XOR2_X1 U2300 ( .A(n2354), .B(n2355), .Z(n2353) );
  NAND2_X1 U2301 ( .A1(b_14_), .A2(a_2_), .ZN(n2355) );
  XNOR2_X1 U2302 ( .A(n2356), .B(n2357), .ZN(n2180) );
  XOR2_X1 U2303 ( .A(n2358), .B(n2359), .Z(n2356) );
  NOR2_X1 U2304 ( .A1(n2360), .A2(n1934), .ZN(n2359) );
  XNOR2_X1 U2305 ( .A(n2361), .B(n2362), .ZN(n2185) );
  XNOR2_X1 U2306 ( .A(n2363), .B(n2364), .ZN(n2362) );
  NAND3_X1 U2307 ( .A1(n2197), .A2(n2198), .A3(n2255), .ZN(n2194) );
  INV_X1 U2308 ( .A(n2195), .ZN(n2255) );
  NAND2_X1 U2309 ( .A1(n2253), .A2(n2365), .ZN(n2195) );
  NAND2_X1 U2310 ( .A1(n2366), .A2(n2367), .ZN(n2365) );
  NAND2_X1 U2311 ( .A1(n2368), .A2(n2369), .ZN(n2198) );
  NAND2_X1 U2312 ( .A1(n2364), .A2(n2370), .ZN(n2369) );
  OR2_X1 U2313 ( .A1(n2363), .A2(n2361), .ZN(n2370) );
  NOR2_X1 U2314 ( .A1(n1934), .A2(n2371), .ZN(n2364) );
  NAND2_X1 U2315 ( .A1(n2361), .A2(n2363), .ZN(n2368) );
  NAND2_X1 U2316 ( .A1(n2372), .A2(n2373), .ZN(n2363) );
  NAND3_X1 U2317 ( .A1(a_1_), .A2(n2374), .A3(b_14_), .ZN(n2373) );
  OR2_X1 U2318 ( .A1(n2358), .A2(n2357), .ZN(n2374) );
  NAND2_X1 U2319 ( .A1(n2357), .A2(n2358), .ZN(n2372) );
  NAND2_X1 U2320 ( .A1(n2375), .A2(n2376), .ZN(n2358) );
  NAND3_X1 U2321 ( .A1(a_2_), .A2(n2377), .A3(b_14_), .ZN(n2376) );
  OR2_X1 U2322 ( .A1(n2354), .A2(n2352), .ZN(n2377) );
  NAND2_X1 U2323 ( .A1(n2352), .A2(n2354), .ZN(n2375) );
  NAND2_X1 U2324 ( .A1(n2378), .A2(n2379), .ZN(n2354) );
  NAND2_X1 U2325 ( .A1(n2351), .A2(n2380), .ZN(n2379) );
  OR2_X1 U2326 ( .A1(n2350), .A2(n2348), .ZN(n2380) );
  NOR2_X1 U2327 ( .A1(n1934), .A2(n2100), .ZN(n2351) );
  NAND2_X1 U2328 ( .A1(n2348), .A2(n2350), .ZN(n2378) );
  NAND2_X1 U2329 ( .A1(n2381), .A2(n2382), .ZN(n2350) );
  NAND3_X1 U2330 ( .A1(a_4_), .A2(n2383), .A3(b_14_), .ZN(n2382) );
  NAND2_X1 U2331 ( .A1(n2345), .A2(n2344), .ZN(n2383) );
  OR2_X1 U2332 ( .A1(n2344), .A2(n2345), .ZN(n2381) );
  AND2_X1 U2333 ( .A1(n2384), .A2(n2385), .ZN(n2345) );
  NAND2_X1 U2334 ( .A1(n2342), .A2(n2386), .ZN(n2385) );
  OR2_X1 U2335 ( .A1(n2341), .A2(n2340), .ZN(n2386) );
  NOR2_X1 U2336 ( .A1(n1934), .A2(n2066), .ZN(n2342) );
  NAND2_X1 U2337 ( .A1(n2340), .A2(n2341), .ZN(n2384) );
  NAND2_X1 U2338 ( .A1(n2387), .A2(n2388), .ZN(n2341) );
  NAND3_X1 U2339 ( .A1(a_6_), .A2(n2389), .A3(b_14_), .ZN(n2388) );
  OR2_X1 U2340 ( .A1(n2337), .A2(n2336), .ZN(n2389) );
  NAND2_X1 U2341 ( .A1(n2336), .A2(n2337), .ZN(n2387) );
  NAND2_X1 U2342 ( .A1(n2390), .A2(n2391), .ZN(n2337) );
  NAND2_X1 U2343 ( .A1(n2334), .A2(n2392), .ZN(n2391) );
  OR2_X1 U2344 ( .A1(n2333), .A2(n2331), .ZN(n2392) );
  NOR2_X1 U2345 ( .A1(n1934), .A2(n2038), .ZN(n2334) );
  NAND2_X1 U2346 ( .A1(n2331), .A2(n2333), .ZN(n2390) );
  NAND2_X1 U2347 ( .A1(n2393), .A2(n2394), .ZN(n2333) );
  NAND3_X1 U2348 ( .A1(a_8_), .A2(n2395), .A3(b_14_), .ZN(n2394) );
  OR2_X1 U2349 ( .A1(n2284), .A2(n2282), .ZN(n2395) );
  NAND2_X1 U2350 ( .A1(n2282), .A2(n2284), .ZN(n2393) );
  NAND2_X1 U2351 ( .A1(n2396), .A2(n2397), .ZN(n2284) );
  NAND2_X1 U2352 ( .A1(n2330), .A2(n2398), .ZN(n2397) );
  OR2_X1 U2353 ( .A1(n2329), .A2(n2328), .ZN(n2398) );
  NOR2_X1 U2354 ( .A1(n1934), .A2(n2008), .ZN(n2330) );
  NAND2_X1 U2355 ( .A1(n2328), .A2(n2329), .ZN(n2396) );
  NAND2_X1 U2356 ( .A1(n2294), .A2(n2399), .ZN(n2329) );
  NAND2_X1 U2357 ( .A1(n2293), .A2(n2295), .ZN(n2399) );
  NAND2_X1 U2358 ( .A1(n2400), .A2(n2401), .ZN(n2295) );
  NAND2_X1 U2359 ( .A1(b_14_), .A2(a_10_), .ZN(n2401) );
  INV_X1 U2360 ( .A(n2402), .ZN(n2400) );
  XNOR2_X1 U2361 ( .A(n2403), .B(n2404), .ZN(n2293) );
  NAND2_X1 U2362 ( .A1(n2405), .A2(n2406), .ZN(n2403) );
  NAND2_X1 U2363 ( .A1(a_10_), .A2(n2402), .ZN(n2294) );
  NAND2_X1 U2364 ( .A1(n2325), .A2(n2407), .ZN(n2402) );
  NAND2_X1 U2365 ( .A1(n2324), .A2(n2326), .ZN(n2407) );
  NAND2_X1 U2366 ( .A1(n2408), .A2(n2409), .ZN(n2326) );
  NAND2_X1 U2367 ( .A1(b_14_), .A2(a_11_), .ZN(n2409) );
  INV_X1 U2368 ( .A(n2410), .ZN(n2408) );
  XNOR2_X1 U2369 ( .A(n2411), .B(n2412), .ZN(n2324) );
  XOR2_X1 U2370 ( .A(n2413), .B(n2414), .Z(n2411) );
  NAND2_X1 U2371 ( .A1(b_13_), .A2(a_12_), .ZN(n2413) );
  NAND2_X1 U2372 ( .A1(a_11_), .A2(n2410), .ZN(n2325) );
  NAND2_X1 U2373 ( .A1(n2415), .A2(n2416), .ZN(n2410) );
  NAND3_X1 U2374 ( .A1(a_12_), .A2(n2417), .A3(b_14_), .ZN(n2416) );
  NAND2_X1 U2375 ( .A1(n2306), .A2(n2304), .ZN(n2417) );
  OR2_X1 U2376 ( .A1(n2304), .A2(n2306), .ZN(n2415) );
  AND2_X1 U2377 ( .A1(n2418), .A2(n2419), .ZN(n2306) );
  NAND2_X1 U2378 ( .A1(n2320), .A2(n2420), .ZN(n2419) );
  OR2_X1 U2379 ( .A1(n2321), .A2(n2322), .ZN(n2420) );
  NOR2_X1 U2380 ( .A1(n1934), .A2(n1952), .ZN(n2320) );
  INV_X1 U2381 ( .A(b_14_), .ZN(n1934) );
  NAND2_X1 U2382 ( .A1(n2322), .A2(n2321), .ZN(n2418) );
  NAND2_X1 U2383 ( .A1(n2421), .A2(n2422), .ZN(n2321) );
  NAND2_X1 U2384 ( .A1(b_12_), .A2(n2423), .ZN(n2422) );
  NAND2_X1 U2385 ( .A1(n1929), .A2(n2424), .ZN(n2423) );
  NAND2_X1 U2386 ( .A1(a_15_), .A2(n1950), .ZN(n2424) );
  NAND2_X1 U2387 ( .A1(b_13_), .A2(n2425), .ZN(n2421) );
  NAND2_X1 U2388 ( .A1(n1932), .A2(n2426), .ZN(n2425) );
  NAND2_X1 U2389 ( .A1(a_14_), .A2(n2174), .ZN(n2426) );
  AND3_X1 U2390 ( .A1(b_14_), .A2(n2173), .A3(b_13_), .ZN(n2322) );
  XOR2_X1 U2391 ( .A(n2427), .B(n2166), .Z(n2304) );
  INV_X1 U2392 ( .A(n1948), .ZN(n2166) );
  XOR2_X1 U2393 ( .A(n2428), .B(n2429), .Z(n2427) );
  XNOR2_X1 U2394 ( .A(n2430), .B(n2431), .ZN(n2328) );
  NAND2_X1 U2395 ( .A1(n2432), .A2(n2433), .ZN(n2430) );
  XNOR2_X1 U2396 ( .A(n2434), .B(n2435), .ZN(n2282) );
  XNOR2_X1 U2397 ( .A(n2436), .B(n2437), .ZN(n2434) );
  XNOR2_X1 U2398 ( .A(n2438), .B(n2439), .ZN(n2331) );
  XOR2_X1 U2399 ( .A(n2440), .B(n2441), .Z(n2439) );
  NAND2_X1 U2400 ( .A1(b_13_), .A2(a_8_), .ZN(n2441) );
  XNOR2_X1 U2401 ( .A(n2442), .B(n2443), .ZN(n2336) );
  XNOR2_X1 U2402 ( .A(n2444), .B(n2445), .ZN(n2443) );
  XNOR2_X1 U2403 ( .A(n2446), .B(n2447), .ZN(n2340) );
  XOR2_X1 U2404 ( .A(n2448), .B(n2449), .Z(n2447) );
  NAND2_X1 U2405 ( .A1(b_13_), .A2(a_6_), .ZN(n2449) );
  XNOR2_X1 U2406 ( .A(n2450), .B(n2451), .ZN(n2344) );
  XOR2_X1 U2407 ( .A(n2452), .B(n2453), .Z(n2450) );
  XNOR2_X1 U2408 ( .A(n2454), .B(n2455), .ZN(n2348) );
  XNOR2_X1 U2409 ( .A(n2456), .B(n2457), .ZN(n2454) );
  NOR2_X1 U2410 ( .A1(n2347), .A2(n1950), .ZN(n2457) );
  XNOR2_X1 U2411 ( .A(n2458), .B(n2459), .ZN(n2352) );
  XNOR2_X1 U2412 ( .A(n2460), .B(n2461), .ZN(n2459) );
  XNOR2_X1 U2413 ( .A(n2462), .B(n2463), .ZN(n2357) );
  XNOR2_X1 U2414 ( .A(n2464), .B(n2465), .ZN(n2462) );
  XNOR2_X1 U2415 ( .A(n2466), .B(n2467), .ZN(n2361) );
  XNOR2_X1 U2416 ( .A(n2468), .B(n2469), .ZN(n2466) );
  NOR2_X1 U2417 ( .A1(n2360), .A2(n1950), .ZN(n2469) );
  XOR2_X1 U2418 ( .A(n2470), .B(n2471), .Z(n2197) );
  XNOR2_X1 U2419 ( .A(n2472), .B(n2473), .ZN(n2471) );
  OR2_X1 U2420 ( .A1(n2367), .A2(n2366), .ZN(n2253) );
  XOR2_X1 U2421 ( .A(n2474), .B(n2475), .Z(n2366) );
  XNOR2_X1 U2422 ( .A(n2476), .B(n2477), .ZN(n2474) );
  NOR2_X1 U2423 ( .A1(n2371), .A2(n2174), .ZN(n2477) );
  NAND2_X1 U2424 ( .A1(n2478), .A2(n2479), .ZN(n2367) );
  NAND2_X1 U2425 ( .A1(n2470), .A2(n2480), .ZN(n2479) );
  NAND2_X1 U2426 ( .A1(n2473), .A2(n2472), .ZN(n2480) );
  XNOR2_X1 U2427 ( .A(n2481), .B(n2482), .ZN(n2470) );
  XOR2_X1 U2428 ( .A(n2483), .B(n2484), .Z(n2481) );
  OR2_X1 U2429 ( .A1(n2472), .A2(n2473), .ZN(n2478) );
  NOR2_X1 U2430 ( .A1(n1950), .A2(n2371), .ZN(n2473) );
  NAND2_X1 U2431 ( .A1(n2485), .A2(n2486), .ZN(n2472) );
  NAND3_X1 U2432 ( .A1(a_1_), .A2(n2487), .A3(b_13_), .ZN(n2486) );
  NAND2_X1 U2433 ( .A1(n2468), .A2(n2467), .ZN(n2487) );
  OR2_X1 U2434 ( .A1(n2467), .A2(n2468), .ZN(n2485) );
  AND2_X1 U2435 ( .A1(n2488), .A2(n2489), .ZN(n2468) );
  NAND2_X1 U2436 ( .A1(n2465), .A2(n2490), .ZN(n2489) );
  NAND2_X1 U2437 ( .A1(n2464), .A2(n2463), .ZN(n2490) );
  NOR2_X1 U2438 ( .A1(n1950), .A2(n2178), .ZN(n2465) );
  OR2_X1 U2439 ( .A1(n2463), .A2(n2464), .ZN(n2488) );
  AND2_X1 U2440 ( .A1(n2491), .A2(n2492), .ZN(n2464) );
  NAND2_X1 U2441 ( .A1(n2461), .A2(n2493), .ZN(n2492) );
  OR2_X1 U2442 ( .A1(n2460), .A2(n2458), .ZN(n2493) );
  NOR2_X1 U2443 ( .A1(n1950), .A2(n2100), .ZN(n2461) );
  NAND2_X1 U2444 ( .A1(n2458), .A2(n2460), .ZN(n2491) );
  NAND2_X1 U2445 ( .A1(n2494), .A2(n2495), .ZN(n2460) );
  NAND3_X1 U2446 ( .A1(a_4_), .A2(n2496), .A3(b_13_), .ZN(n2495) );
  NAND2_X1 U2447 ( .A1(n2456), .A2(n2455), .ZN(n2496) );
  OR2_X1 U2448 ( .A1(n2455), .A2(n2456), .ZN(n2494) );
  AND2_X1 U2449 ( .A1(n2497), .A2(n2498), .ZN(n2456) );
  NAND2_X1 U2450 ( .A1(n2453), .A2(n2499), .ZN(n2498) );
  OR2_X1 U2451 ( .A1(n2451), .A2(n2452), .ZN(n2499) );
  NOR2_X1 U2452 ( .A1(n1950), .A2(n2066), .ZN(n2453) );
  NAND2_X1 U2453 ( .A1(n2451), .A2(n2452), .ZN(n2497) );
  NAND2_X1 U2454 ( .A1(n2500), .A2(n2501), .ZN(n2452) );
  NAND3_X1 U2455 ( .A1(a_6_), .A2(n2502), .A3(b_13_), .ZN(n2501) );
  OR2_X1 U2456 ( .A1(n2448), .A2(n2446), .ZN(n2502) );
  NAND2_X1 U2457 ( .A1(n2446), .A2(n2448), .ZN(n2500) );
  NAND2_X1 U2458 ( .A1(n2503), .A2(n2504), .ZN(n2448) );
  NAND2_X1 U2459 ( .A1(n2445), .A2(n2505), .ZN(n2504) );
  OR2_X1 U2460 ( .A1(n2444), .A2(n2442), .ZN(n2505) );
  NOR2_X1 U2461 ( .A1(n1950), .A2(n2038), .ZN(n2445) );
  NAND2_X1 U2462 ( .A1(n2442), .A2(n2444), .ZN(n2503) );
  NAND2_X1 U2463 ( .A1(n2506), .A2(n2507), .ZN(n2444) );
  NAND3_X1 U2464 ( .A1(a_8_), .A2(n2508), .A3(b_13_), .ZN(n2507) );
  OR2_X1 U2465 ( .A1(n2440), .A2(n2438), .ZN(n2508) );
  NAND2_X1 U2466 ( .A1(n2438), .A2(n2440), .ZN(n2506) );
  NAND2_X1 U2467 ( .A1(n2509), .A2(n2510), .ZN(n2440) );
  NAND2_X1 U2468 ( .A1(n2437), .A2(n2511), .ZN(n2510) );
  NAND2_X1 U2469 ( .A1(n2436), .A2(n2435), .ZN(n2511) );
  NOR2_X1 U2470 ( .A1(n1950), .A2(n2008), .ZN(n2437) );
  OR2_X1 U2471 ( .A1(n2435), .A2(n2436), .ZN(n2509) );
  AND2_X1 U2472 ( .A1(n2432), .A2(n2512), .ZN(n2436) );
  NAND2_X1 U2473 ( .A1(n2431), .A2(n2433), .ZN(n2512) );
  NAND2_X1 U2474 ( .A1(n2513), .A2(n2514), .ZN(n2433) );
  NAND2_X1 U2475 ( .A1(b_13_), .A2(a_10_), .ZN(n2514) );
  INV_X1 U2476 ( .A(n2515), .ZN(n2513) );
  XNOR2_X1 U2477 ( .A(n2516), .B(n2517), .ZN(n2431) );
  NAND2_X1 U2478 ( .A1(n2518), .A2(n2519), .ZN(n2516) );
  NAND2_X1 U2479 ( .A1(a_10_), .A2(n2515), .ZN(n2432) );
  NAND2_X1 U2480 ( .A1(n2405), .A2(n2520), .ZN(n2515) );
  NAND2_X1 U2481 ( .A1(n2404), .A2(n2406), .ZN(n2520) );
  NAND2_X1 U2482 ( .A1(n2521), .A2(n2522), .ZN(n2406) );
  NAND2_X1 U2483 ( .A1(b_13_), .A2(a_11_), .ZN(n2522) );
  INV_X1 U2484 ( .A(n2523), .ZN(n2521) );
  XOR2_X1 U2485 ( .A(n2524), .B(n2525), .Z(n2404) );
  XNOR2_X1 U2486 ( .A(n2526), .B(n2527), .ZN(n2524) );
  NAND2_X1 U2487 ( .A1(a_11_), .A2(n2523), .ZN(n2405) );
  NAND2_X1 U2488 ( .A1(n2528), .A2(n2529), .ZN(n2523) );
  NAND3_X1 U2489 ( .A1(a_12_), .A2(n2530), .A3(b_13_), .ZN(n2529) );
  NAND2_X1 U2490 ( .A1(n2414), .A2(n2412), .ZN(n2530) );
  OR2_X1 U2491 ( .A1(n2412), .A2(n2414), .ZN(n2528) );
  AND2_X1 U2492 ( .A1(n2531), .A2(n2532), .ZN(n2414) );
  NAND2_X1 U2493 ( .A1(n1948), .A2(n2533), .ZN(n2532) );
  OR2_X1 U2494 ( .A1(n2428), .A2(n2429), .ZN(n2533) );
  NOR2_X1 U2495 ( .A1(n1950), .A2(n1952), .ZN(n1948) );
  INV_X1 U2496 ( .A(b_13_), .ZN(n1950) );
  NAND2_X1 U2497 ( .A1(n2429), .A2(n2428), .ZN(n2531) );
  NAND2_X1 U2498 ( .A1(n2534), .A2(n2535), .ZN(n2428) );
  NAND2_X1 U2499 ( .A1(b_11_), .A2(n2536), .ZN(n2535) );
  NAND2_X1 U2500 ( .A1(n1929), .A2(n2537), .ZN(n2536) );
  NAND2_X1 U2501 ( .A1(a_15_), .A2(n2174), .ZN(n2537) );
  NAND2_X1 U2502 ( .A1(b_12_), .A2(n2538), .ZN(n2534) );
  NAND2_X1 U2503 ( .A1(n1932), .A2(n2539), .ZN(n2538) );
  NAND2_X1 U2504 ( .A1(a_14_), .A2(n1979), .ZN(n2539) );
  AND3_X1 U2505 ( .A1(b_12_), .A2(n2173), .A3(b_13_), .ZN(n2429) );
  XNOR2_X1 U2506 ( .A(n2540), .B(n2541), .ZN(n2412) );
  XOR2_X1 U2507 ( .A(n2542), .B(n2543), .Z(n2540) );
  XNOR2_X1 U2508 ( .A(n2544), .B(n2545), .ZN(n2435) );
  NOR2_X1 U2509 ( .A1(n2546), .A2(n2547), .ZN(n2545) );
  NOR2_X1 U2510 ( .A1(n2548), .A2(n2549), .ZN(n2546) );
  NOR2_X1 U2511 ( .A1(n2550), .A2(n2174), .ZN(n2548) );
  XOR2_X1 U2512 ( .A(n2551), .B(n2552), .Z(n2438) );
  XOR2_X1 U2513 ( .A(n2553), .B(n2554), .Z(n2551) );
  XOR2_X1 U2514 ( .A(n2555), .B(n2556), .Z(n2442) );
  XOR2_X1 U2515 ( .A(n2557), .B(n2558), .Z(n2555) );
  NOR2_X1 U2516 ( .A1(n2176), .A2(n2174), .ZN(n2558) );
  XNOR2_X1 U2517 ( .A(n2559), .B(n2560), .ZN(n2446) );
  XNOR2_X1 U2518 ( .A(n2561), .B(n2562), .ZN(n2560) );
  XNOR2_X1 U2519 ( .A(n2563), .B(n2564), .ZN(n2451) );
  XNOR2_X1 U2520 ( .A(n2565), .B(n2566), .ZN(n2563) );
  NOR2_X1 U2521 ( .A1(n2056), .A2(n2174), .ZN(n2566) );
  XNOR2_X1 U2522 ( .A(n2567), .B(n2568), .ZN(n2455) );
  XOR2_X1 U2523 ( .A(n2569), .B(n2570), .Z(n2567) );
  XOR2_X1 U2524 ( .A(n2571), .B(n2572), .Z(n2458) );
  XOR2_X1 U2525 ( .A(n2573), .B(n2574), .Z(n2571) );
  NOR2_X1 U2526 ( .A1(n2347), .A2(n2174), .ZN(n2574) );
  XOR2_X1 U2527 ( .A(n2575), .B(n2576), .Z(n2463) );
  XOR2_X1 U2528 ( .A(n2577), .B(n2578), .Z(n2576) );
  NAND2_X1 U2529 ( .A1(b_12_), .A2(a_3_), .ZN(n2578) );
  XNOR2_X1 U2530 ( .A(n2579), .B(n2580), .ZN(n2467) );
  XOR2_X1 U2531 ( .A(n2581), .B(n2582), .Z(n2579) );
  XOR2_X1 U2532 ( .A(n2238), .B(n2237), .Z(n2200) );
  XOR2_X1 U2533 ( .A(n2249), .B(n2583), .Z(n2237) );
  XNOR2_X1 U2534 ( .A(n2252), .B(n2251), .ZN(n2583) );
  NOR2_X1 U2535 ( .A1(n2371), .A2(n1979), .ZN(n2251) );
  NAND2_X1 U2536 ( .A1(n2584), .A2(n2585), .ZN(n2252) );
  NAND3_X1 U2537 ( .A1(b_11_), .A2(n2586), .A3(a_1_), .ZN(n2585) );
  OR2_X1 U2538 ( .A1(n2587), .A2(n2588), .ZN(n2586) );
  NAND2_X1 U2539 ( .A1(n2588), .A2(n2587), .ZN(n2584) );
  XOR2_X1 U2540 ( .A(n2589), .B(n2590), .Z(n2249) );
  XNOR2_X1 U2541 ( .A(n2591), .B(n2592), .ZN(n2590) );
  NAND2_X1 U2542 ( .A1(n2593), .A2(n2594), .ZN(n2238) );
  NAND3_X1 U2543 ( .A1(a_0_), .A2(n2595), .A3(b_12_), .ZN(n2594) );
  NAND2_X1 U2544 ( .A1(n2476), .A2(n2475), .ZN(n2595) );
  OR2_X1 U2545 ( .A1(n2475), .A2(n2476), .ZN(n2593) );
  AND2_X1 U2546 ( .A1(n2596), .A2(n2597), .ZN(n2476) );
  NAND2_X1 U2547 ( .A1(n2484), .A2(n2598), .ZN(n2597) );
  OR2_X1 U2548 ( .A1(n2483), .A2(n2482), .ZN(n2598) );
  NOR2_X1 U2549 ( .A1(n2174), .A2(n2360), .ZN(n2484) );
  NAND2_X1 U2550 ( .A1(n2482), .A2(n2483), .ZN(n2596) );
  NAND2_X1 U2551 ( .A1(n2599), .A2(n2600), .ZN(n2483) );
  NAND2_X1 U2552 ( .A1(n2582), .A2(n2601), .ZN(n2600) );
  OR2_X1 U2553 ( .A1(n2581), .A2(n2580), .ZN(n2601) );
  NOR2_X1 U2554 ( .A1(n2174), .A2(n2178), .ZN(n2582) );
  NAND2_X1 U2555 ( .A1(n2580), .A2(n2581), .ZN(n2599) );
  NAND2_X1 U2556 ( .A1(n2602), .A2(n2603), .ZN(n2581) );
  NAND3_X1 U2557 ( .A1(a_3_), .A2(n2604), .A3(b_12_), .ZN(n2603) );
  OR2_X1 U2558 ( .A1(n2577), .A2(n2575), .ZN(n2604) );
  NAND2_X1 U2559 ( .A1(n2575), .A2(n2577), .ZN(n2602) );
  NAND2_X1 U2560 ( .A1(n2605), .A2(n2606), .ZN(n2577) );
  NAND3_X1 U2561 ( .A1(a_4_), .A2(n2607), .A3(b_12_), .ZN(n2606) );
  OR2_X1 U2562 ( .A1(n2573), .A2(n2572), .ZN(n2607) );
  NAND2_X1 U2563 ( .A1(n2572), .A2(n2573), .ZN(n2605) );
  NAND2_X1 U2564 ( .A1(n2608), .A2(n2609), .ZN(n2573) );
  NAND2_X1 U2565 ( .A1(n2570), .A2(n2610), .ZN(n2609) );
  OR2_X1 U2566 ( .A1(n2569), .A2(n2568), .ZN(n2610) );
  NOR2_X1 U2567 ( .A1(n2174), .A2(n2066), .ZN(n2570) );
  NAND2_X1 U2568 ( .A1(n2568), .A2(n2569), .ZN(n2608) );
  NAND2_X1 U2569 ( .A1(n2611), .A2(n2612), .ZN(n2569) );
  NAND3_X1 U2570 ( .A1(a_6_), .A2(n2613), .A3(b_12_), .ZN(n2612) );
  NAND2_X1 U2571 ( .A1(n2565), .A2(n2564), .ZN(n2613) );
  OR2_X1 U2572 ( .A1(n2564), .A2(n2565), .ZN(n2611) );
  AND2_X1 U2573 ( .A1(n2614), .A2(n2615), .ZN(n2565) );
  NAND2_X1 U2574 ( .A1(n2562), .A2(n2616), .ZN(n2615) );
  OR2_X1 U2575 ( .A1(n2561), .A2(n2559), .ZN(n2616) );
  NOR2_X1 U2576 ( .A1(n2174), .A2(n2038), .ZN(n2562) );
  NAND2_X1 U2577 ( .A1(n2559), .A2(n2561), .ZN(n2614) );
  NAND2_X1 U2578 ( .A1(n2617), .A2(n2618), .ZN(n2561) );
  NAND3_X1 U2579 ( .A1(a_8_), .A2(n2619), .A3(b_12_), .ZN(n2618) );
  OR2_X1 U2580 ( .A1(n2557), .A2(n2556), .ZN(n2619) );
  NAND2_X1 U2581 ( .A1(n2556), .A2(n2557), .ZN(n2617) );
  NAND2_X1 U2582 ( .A1(n2620), .A2(n2621), .ZN(n2557) );
  NAND2_X1 U2583 ( .A1(n2554), .A2(n2622), .ZN(n2621) );
  OR2_X1 U2584 ( .A1(n2553), .A2(n2552), .ZN(n2622) );
  NOR2_X1 U2585 ( .A1(n2174), .A2(n2008), .ZN(n2554) );
  NAND2_X1 U2586 ( .A1(n2552), .A2(n2553), .ZN(n2620) );
  OR2_X1 U2587 ( .A1(n2547), .A2(n2623), .ZN(n2553) );
  AND2_X1 U2588 ( .A1(n2544), .A2(n2624), .ZN(n2623) );
  NAND2_X1 U2589 ( .A1(n2625), .A2(n2626), .ZN(n2624) );
  NAND2_X1 U2590 ( .A1(b_12_), .A2(a_10_), .ZN(n2626) );
  XOR2_X1 U2591 ( .A(n2627), .B(n2628), .Z(n2544) );
  XNOR2_X1 U2592 ( .A(n2629), .B(n2162), .ZN(n2627) );
  INV_X1 U2593 ( .A(n1977), .ZN(n2162) );
  NOR2_X1 U2594 ( .A1(n2550), .A2(n2625), .ZN(n2547) );
  INV_X1 U2595 ( .A(n2549), .ZN(n2625) );
  NAND2_X1 U2596 ( .A1(n2518), .A2(n2630), .ZN(n2549) );
  NAND2_X1 U2597 ( .A1(n2517), .A2(n2519), .ZN(n2630) );
  NAND2_X1 U2598 ( .A1(n2631), .A2(n2632), .ZN(n2519) );
  NAND2_X1 U2599 ( .A1(b_12_), .A2(a_11_), .ZN(n2632) );
  INV_X1 U2600 ( .A(n2633), .ZN(n2631) );
  XNOR2_X1 U2601 ( .A(n2634), .B(n2635), .ZN(n2517) );
  XOR2_X1 U2602 ( .A(n2636), .B(n2637), .Z(n2634) );
  NAND2_X1 U2603 ( .A1(a_12_), .A2(b_11_), .ZN(n2636) );
  NAND2_X1 U2604 ( .A1(a_11_), .A2(n2633), .ZN(n2518) );
  NAND2_X1 U2605 ( .A1(n2638), .A2(n2639), .ZN(n2633) );
  NAND2_X1 U2606 ( .A1(n2525), .A2(n2640), .ZN(n2639) );
  NAND2_X1 U2607 ( .A1(n2527), .A2(n1964), .ZN(n2640) );
  INV_X1 U2608 ( .A(n2526), .ZN(n1964) );
  INV_X1 U2609 ( .A(n2641), .ZN(n2527) );
  XOR2_X1 U2610 ( .A(n2642), .B(n2643), .Z(n2525) );
  XOR2_X1 U2611 ( .A(n2644), .B(n2645), .Z(n2642) );
  NAND2_X1 U2612 ( .A1(n2526), .A2(n2641), .ZN(n2638) );
  NAND2_X1 U2613 ( .A1(n2646), .A2(n2647), .ZN(n2641) );
  NAND2_X1 U2614 ( .A1(n2541), .A2(n2648), .ZN(n2647) );
  OR2_X1 U2615 ( .A1(n2542), .A2(n2543), .ZN(n2648) );
  NOR2_X1 U2616 ( .A1(n2174), .A2(n1952), .ZN(n2541) );
  NAND2_X1 U2617 ( .A1(n2543), .A2(n2542), .ZN(n2646) );
  NAND2_X1 U2618 ( .A1(n2649), .A2(n2650), .ZN(n2542) );
  NAND2_X1 U2619 ( .A1(b_10_), .A2(n2651), .ZN(n2650) );
  NAND2_X1 U2620 ( .A1(n1929), .A2(n2652), .ZN(n2651) );
  NAND2_X1 U2621 ( .A1(a_15_), .A2(n1979), .ZN(n2652) );
  NAND2_X1 U2622 ( .A1(b_11_), .A2(n2653), .ZN(n2649) );
  NAND2_X1 U2623 ( .A1(n1932), .A2(n2654), .ZN(n2653) );
  NAND2_X1 U2624 ( .A1(a_14_), .A2(n2655), .ZN(n2654) );
  AND3_X1 U2625 ( .A1(n2173), .A2(b_11_), .A3(b_12_), .ZN(n2543) );
  NOR2_X1 U2626 ( .A1(n2174), .A2(n1970), .ZN(n2526) );
  INV_X1 U2627 ( .A(b_12_), .ZN(n2174) );
  XNOR2_X1 U2628 ( .A(n2656), .B(n2657), .ZN(n2552) );
  NAND2_X1 U2629 ( .A1(n2658), .A2(n2659), .ZN(n2656) );
  XNOR2_X1 U2630 ( .A(n2660), .B(n2661), .ZN(n2556) );
  XNOR2_X1 U2631 ( .A(n2662), .B(n2663), .ZN(n2660) );
  XNOR2_X1 U2632 ( .A(n2664), .B(n2665), .ZN(n2559) );
  XNOR2_X1 U2633 ( .A(n2666), .B(n2667), .ZN(n2664) );
  NOR2_X1 U2634 ( .A1(n1979), .A2(n2176), .ZN(n2667) );
  XOR2_X1 U2635 ( .A(n2668), .B(n2669), .Z(n2564) );
  XNOR2_X1 U2636 ( .A(n2670), .B(n2671), .ZN(n2669) );
  XNOR2_X1 U2637 ( .A(n2672), .B(n2673), .ZN(n2568) );
  XOR2_X1 U2638 ( .A(n2674), .B(n2675), .Z(n2673) );
  NAND2_X1 U2639 ( .A1(a_6_), .A2(b_11_), .ZN(n2675) );
  XNOR2_X1 U2640 ( .A(n2676), .B(n2677), .ZN(n2572) );
  XNOR2_X1 U2641 ( .A(n2678), .B(n2679), .ZN(n2676) );
  XNOR2_X1 U2642 ( .A(n2680), .B(n2681), .ZN(n2575) );
  XNOR2_X1 U2643 ( .A(n2682), .B(n2683), .ZN(n2680) );
  XNOR2_X1 U2644 ( .A(n2684), .B(n2685), .ZN(n2580) );
  XOR2_X1 U2645 ( .A(n2686), .B(n2687), .Z(n2685) );
  NAND2_X1 U2646 ( .A1(a_3_), .A2(b_11_), .ZN(n2687) );
  XNOR2_X1 U2647 ( .A(n2688), .B(n2689), .ZN(n2482) );
  XOR2_X1 U2648 ( .A(n2690), .B(n2691), .Z(n2689) );
  NAND2_X1 U2649 ( .A1(a_2_), .A2(b_11_), .ZN(n2691) );
  XOR2_X1 U2650 ( .A(n2588), .B(n2692), .Z(n2475) );
  XOR2_X1 U2651 ( .A(n2587), .B(n2693), .Z(n2692) );
  NAND2_X1 U2652 ( .A1(a_1_), .A2(b_11_), .ZN(n2693) );
  NAND2_X1 U2653 ( .A1(n2694), .A2(n2695), .ZN(n2587) );
  NAND3_X1 U2654 ( .A1(b_11_), .A2(n2696), .A3(a_2_), .ZN(n2695) );
  OR2_X1 U2655 ( .A1(n2690), .A2(n2688), .ZN(n2696) );
  NAND2_X1 U2656 ( .A1(n2688), .A2(n2690), .ZN(n2694) );
  NAND2_X1 U2657 ( .A1(n2697), .A2(n2698), .ZN(n2690) );
  NAND3_X1 U2658 ( .A1(b_11_), .A2(n2699), .A3(a_3_), .ZN(n2698) );
  OR2_X1 U2659 ( .A1(n2686), .A2(n2684), .ZN(n2699) );
  NAND2_X1 U2660 ( .A1(n2684), .A2(n2686), .ZN(n2697) );
  NAND2_X1 U2661 ( .A1(n2700), .A2(n2701), .ZN(n2686) );
  NAND2_X1 U2662 ( .A1(n2683), .A2(n2702), .ZN(n2701) );
  NAND2_X1 U2663 ( .A1(n2682), .A2(n2681), .ZN(n2702) );
  NOR2_X1 U2664 ( .A1(n1979), .A2(n2347), .ZN(n2683) );
  OR2_X1 U2665 ( .A1(n2681), .A2(n2682), .ZN(n2700) );
  AND2_X1 U2666 ( .A1(n2703), .A2(n2704), .ZN(n2682) );
  NAND2_X1 U2667 ( .A1(n2679), .A2(n2705), .ZN(n2704) );
  NAND2_X1 U2668 ( .A1(n2678), .A2(n2677), .ZN(n2705) );
  NOR2_X1 U2669 ( .A1(n2066), .A2(n1979), .ZN(n2679) );
  OR2_X1 U2670 ( .A1(n2677), .A2(n2678), .ZN(n2703) );
  AND2_X1 U2671 ( .A1(n2706), .A2(n2707), .ZN(n2678) );
  NAND3_X1 U2672 ( .A1(b_11_), .A2(n2708), .A3(a_6_), .ZN(n2707) );
  OR2_X1 U2673 ( .A1(n2674), .A2(n2672), .ZN(n2708) );
  NAND2_X1 U2674 ( .A1(n2672), .A2(n2674), .ZN(n2706) );
  NAND2_X1 U2675 ( .A1(n2709), .A2(n2710), .ZN(n2674) );
  NAND2_X1 U2676 ( .A1(n2671), .A2(n2711), .ZN(n2710) );
  OR2_X1 U2677 ( .A1(n2670), .A2(n2668), .ZN(n2711) );
  NOR2_X1 U2678 ( .A1(n2038), .A2(n1979), .ZN(n2671) );
  NAND2_X1 U2679 ( .A1(n2668), .A2(n2670), .ZN(n2709) );
  NAND2_X1 U2680 ( .A1(n2712), .A2(n2713), .ZN(n2670) );
  NAND3_X1 U2681 ( .A1(b_11_), .A2(n2714), .A3(a_8_), .ZN(n2713) );
  NAND2_X1 U2682 ( .A1(n2666), .A2(n2665), .ZN(n2714) );
  OR2_X1 U2683 ( .A1(n2665), .A2(n2666), .ZN(n2712) );
  AND2_X1 U2684 ( .A1(n2715), .A2(n2716), .ZN(n2666) );
  NAND2_X1 U2685 ( .A1(n2663), .A2(n2717), .ZN(n2716) );
  NAND2_X1 U2686 ( .A1(n2662), .A2(n2661), .ZN(n2717) );
  NOR2_X1 U2687 ( .A1(n2008), .A2(n1979), .ZN(n2663) );
  OR2_X1 U2688 ( .A1(n2661), .A2(n2662), .ZN(n2715) );
  AND2_X1 U2689 ( .A1(n2658), .A2(n2718), .ZN(n2662) );
  NAND2_X1 U2690 ( .A1(n2657), .A2(n2659), .ZN(n2718) );
  NAND2_X1 U2691 ( .A1(n2719), .A2(n2720), .ZN(n2659) );
  NAND2_X1 U2692 ( .A1(a_10_), .A2(b_11_), .ZN(n2720) );
  INV_X1 U2693 ( .A(n2721), .ZN(n2719) );
  XNOR2_X1 U2694 ( .A(n2722), .B(n2723), .ZN(n2657) );
  NAND2_X1 U2695 ( .A1(n2724), .A2(n2725), .ZN(n2722) );
  NAND2_X1 U2696 ( .A1(a_10_), .A2(n2721), .ZN(n2658) );
  NAND2_X1 U2697 ( .A1(n2726), .A2(n2727), .ZN(n2721) );
  NAND2_X1 U2698 ( .A1(n2628), .A2(n2728), .ZN(n2727) );
  OR2_X1 U2699 ( .A1(n2629), .A2(n1977), .ZN(n2728) );
  XNOR2_X1 U2700 ( .A(n2729), .B(n2730), .ZN(n2628) );
  XOR2_X1 U2701 ( .A(n2731), .B(n2732), .Z(n2729) );
  NAND2_X1 U2702 ( .A1(a_12_), .A2(b_10_), .ZN(n2731) );
  NAND2_X1 U2703 ( .A1(n1977), .A2(n2629), .ZN(n2726) );
  NAND2_X1 U2704 ( .A1(n2733), .A2(n2734), .ZN(n2629) );
  NAND3_X1 U2705 ( .A1(b_11_), .A2(n2735), .A3(a_12_), .ZN(n2734) );
  NAND2_X1 U2706 ( .A1(n2637), .A2(n2635), .ZN(n2735) );
  OR2_X1 U2707 ( .A1(n2635), .A2(n2637), .ZN(n2733) );
  AND2_X1 U2708 ( .A1(n2736), .A2(n2737), .ZN(n2637) );
  NAND2_X1 U2709 ( .A1(n2643), .A2(n2738), .ZN(n2737) );
  OR2_X1 U2710 ( .A1(n2644), .A2(n2645), .ZN(n2738) );
  NOR2_X1 U2711 ( .A1(n1952), .A2(n1979), .ZN(n2643) );
  NAND2_X1 U2712 ( .A1(n2645), .A2(n2644), .ZN(n2736) );
  NAND2_X1 U2713 ( .A1(n2739), .A2(n2740), .ZN(n2644) );
  NAND2_X1 U2714 ( .A1(b_10_), .A2(n2741), .ZN(n2740) );
  NAND2_X1 U2715 ( .A1(n1932), .A2(n2742), .ZN(n2741) );
  NAND2_X1 U2716 ( .A1(a_14_), .A2(n2010), .ZN(n2742) );
  NAND2_X1 U2717 ( .A1(b_9_), .A2(n2743), .ZN(n2739) );
  NAND2_X1 U2718 ( .A1(n1929), .A2(n2744), .ZN(n2743) );
  NAND2_X1 U2719 ( .A1(a_15_), .A2(n2655), .ZN(n2744) );
  AND3_X1 U2720 ( .A1(n2173), .A2(b_11_), .A3(b_10_), .ZN(n2645) );
  XNOR2_X1 U2721 ( .A(n2745), .B(n2746), .ZN(n2635) );
  XOR2_X1 U2722 ( .A(n2747), .B(n2748), .Z(n2745) );
  NOR2_X1 U2723 ( .A1(n1981), .A2(n1979), .ZN(n1977) );
  INV_X1 U2724 ( .A(b_11_), .ZN(n1979) );
  XOR2_X1 U2725 ( .A(n2749), .B(n2750), .Z(n2661) );
  XNOR2_X1 U2726 ( .A(n1993), .B(n2751), .ZN(n2750) );
  XNOR2_X1 U2727 ( .A(n2752), .B(n2753), .ZN(n2665) );
  XOR2_X1 U2728 ( .A(n2754), .B(n2755), .Z(n2752) );
  XNOR2_X1 U2729 ( .A(n2756), .B(n2757), .ZN(n2668) );
  XNOR2_X1 U2730 ( .A(n2758), .B(n2759), .ZN(n2756) );
  NOR2_X1 U2731 ( .A1(n2655), .A2(n2176), .ZN(n2759) );
  XNOR2_X1 U2732 ( .A(n2760), .B(n2761), .ZN(n2672) );
  XNOR2_X1 U2733 ( .A(n2762), .B(n2763), .ZN(n2761) );
  XOR2_X1 U2734 ( .A(n2764), .B(n2765), .Z(n2677) );
  XOR2_X1 U2735 ( .A(n2766), .B(n2767), .Z(n2765) );
  NAND2_X1 U2736 ( .A1(a_6_), .A2(b_10_), .ZN(n2767) );
  XNOR2_X1 U2737 ( .A(n2768), .B(n2769), .ZN(n2681) );
  XOR2_X1 U2738 ( .A(n2770), .B(n2771), .Z(n2768) );
  NOR2_X1 U2739 ( .A1(n2066), .A2(n2655), .ZN(n2771) );
  XNOR2_X1 U2740 ( .A(n2772), .B(n2773), .ZN(n2684) );
  XNOR2_X1 U2741 ( .A(n2774), .B(n2775), .ZN(n2773) );
  XOR2_X1 U2742 ( .A(n2776), .B(n2777), .Z(n2688) );
  XOR2_X1 U2743 ( .A(n2778), .B(n2779), .Z(n2776) );
  XOR2_X1 U2744 ( .A(n2780), .B(n2781), .Z(n2588) );
  XOR2_X1 U2745 ( .A(n2782), .B(n2783), .Z(n2780) );
  NOR2_X1 U2746 ( .A1(n2655), .A2(n2178), .ZN(n2783) );
  NAND2_X1 U2747 ( .A1(n2784), .A2(n2785), .ZN(n1887) );
  NAND2_X1 U2748 ( .A1(n2234), .A2(n2235), .ZN(n2785) );
  XNOR2_X1 U2749 ( .A(n2786), .B(n2787), .ZN(n2784) );
  NAND3_X1 U2750 ( .A1(n2234), .A2(n2235), .A3(n2788), .ZN(n1886) );
  XOR2_X1 U2751 ( .A(n2786), .B(n2787), .Z(n2788) );
  NAND2_X1 U2752 ( .A1(n2245), .A2(n2789), .ZN(n2235) );
  NAND2_X1 U2753 ( .A1(n2244), .A2(n2246), .ZN(n2789) );
  NAND2_X1 U2754 ( .A1(n2790), .A2(n2791), .ZN(n2246) );
  NAND2_X1 U2755 ( .A1(a_0_), .A2(b_10_), .ZN(n2791) );
  INV_X1 U2756 ( .A(n2792), .ZN(n2790) );
  XNOR2_X1 U2757 ( .A(n2793), .B(n2794), .ZN(n2244) );
  XOR2_X1 U2758 ( .A(n2795), .B(n2796), .Z(n2794) );
  NAND2_X1 U2759 ( .A1(a_1_), .A2(b_9_), .ZN(n2796) );
  NAND2_X1 U2760 ( .A1(a_0_), .A2(n2792), .ZN(n2245) );
  NAND2_X1 U2761 ( .A1(n2797), .A2(n2798), .ZN(n2792) );
  NAND2_X1 U2762 ( .A1(n2592), .A2(n2799), .ZN(n2798) );
  OR2_X1 U2763 ( .A1(n2589), .A2(n2591), .ZN(n2799) );
  NOR2_X1 U2764 ( .A1(n2360), .A2(n2655), .ZN(n2592) );
  NAND2_X1 U2765 ( .A1(n2589), .A2(n2591), .ZN(n2797) );
  NAND2_X1 U2766 ( .A1(n2800), .A2(n2801), .ZN(n2591) );
  NAND3_X1 U2767 ( .A1(b_10_), .A2(n2802), .A3(a_2_), .ZN(n2801) );
  OR2_X1 U2768 ( .A1(n2782), .A2(n2781), .ZN(n2802) );
  NAND2_X1 U2769 ( .A1(n2781), .A2(n2782), .ZN(n2800) );
  NAND2_X1 U2770 ( .A1(n2803), .A2(n2804), .ZN(n2782) );
  NAND2_X1 U2771 ( .A1(n2779), .A2(n2805), .ZN(n2804) );
  OR2_X1 U2772 ( .A1(n2777), .A2(n2778), .ZN(n2805) );
  NOR2_X1 U2773 ( .A1(n2100), .A2(n2655), .ZN(n2779) );
  NAND2_X1 U2774 ( .A1(n2777), .A2(n2778), .ZN(n2803) );
  NAND2_X1 U2775 ( .A1(n2806), .A2(n2807), .ZN(n2778) );
  NAND2_X1 U2776 ( .A1(n2775), .A2(n2808), .ZN(n2807) );
  OR2_X1 U2777 ( .A1(n2772), .A2(n2774), .ZN(n2808) );
  NOR2_X1 U2778 ( .A1(n2655), .A2(n2347), .ZN(n2775) );
  NAND2_X1 U2779 ( .A1(n2772), .A2(n2774), .ZN(n2806) );
  NAND2_X1 U2780 ( .A1(n2809), .A2(n2810), .ZN(n2774) );
  NAND3_X1 U2781 ( .A1(a_5_), .A2(n2811), .A3(b_10_), .ZN(n2810) );
  OR2_X1 U2782 ( .A1(n2769), .A2(n2770), .ZN(n2811) );
  NAND2_X1 U2783 ( .A1(n2769), .A2(n2770), .ZN(n2809) );
  NAND2_X1 U2784 ( .A1(n2812), .A2(n2813), .ZN(n2770) );
  NAND3_X1 U2785 ( .A1(b_10_), .A2(n2814), .A3(a_6_), .ZN(n2813) );
  OR2_X1 U2786 ( .A1(n2764), .A2(n2766), .ZN(n2814) );
  NAND2_X1 U2787 ( .A1(n2764), .A2(n2766), .ZN(n2812) );
  NAND2_X1 U2788 ( .A1(n2815), .A2(n2816), .ZN(n2766) );
  NAND2_X1 U2789 ( .A1(n2763), .A2(n2817), .ZN(n2816) );
  OR2_X1 U2790 ( .A1(n2760), .A2(n2762), .ZN(n2817) );
  NOR2_X1 U2791 ( .A1(n2655), .A2(n2038), .ZN(n2763) );
  NAND2_X1 U2792 ( .A1(n2760), .A2(n2762), .ZN(n2815) );
  NAND2_X1 U2793 ( .A1(n2818), .A2(n2819), .ZN(n2762) );
  NAND3_X1 U2794 ( .A1(b_10_), .A2(n2820), .A3(a_8_), .ZN(n2819) );
  NAND2_X1 U2795 ( .A1(n2758), .A2(n2757), .ZN(n2820) );
  OR2_X1 U2796 ( .A1(n2757), .A2(n2758), .ZN(n2818) );
  AND2_X1 U2797 ( .A1(n2821), .A2(n2822), .ZN(n2758) );
  NAND2_X1 U2798 ( .A1(n2755), .A2(n2823), .ZN(n2822) );
  OR2_X1 U2799 ( .A1(n2753), .A2(n2754), .ZN(n2823) );
  NOR2_X1 U2800 ( .A1(n2655), .A2(n2008), .ZN(n2755) );
  NAND2_X1 U2801 ( .A1(n2753), .A2(n2754), .ZN(n2821) );
  NAND2_X1 U2802 ( .A1(n2824), .A2(n2825), .ZN(n2754) );
  NAND2_X1 U2803 ( .A1(n2749), .A2(n2826), .ZN(n2825) );
  OR2_X1 U2804 ( .A1(n2751), .A2(n1993), .ZN(n2826) );
  XNOR2_X1 U2805 ( .A(n2827), .B(n2828), .ZN(n2749) );
  NAND2_X1 U2806 ( .A1(n2829), .A2(n2830), .ZN(n2827) );
  NAND2_X1 U2807 ( .A1(n1993), .A2(n2751), .ZN(n2824) );
  NAND2_X1 U2808 ( .A1(n2724), .A2(n2831), .ZN(n2751) );
  NAND2_X1 U2809 ( .A1(n2723), .A2(n2725), .ZN(n2831) );
  NAND2_X1 U2810 ( .A1(n2832), .A2(n2833), .ZN(n2725) );
  NAND2_X1 U2811 ( .A1(b_10_), .A2(a_11_), .ZN(n2833) );
  INV_X1 U2812 ( .A(n2834), .ZN(n2832) );
  XNOR2_X1 U2813 ( .A(n2835), .B(n2836), .ZN(n2723) );
  XOR2_X1 U2814 ( .A(n2837), .B(n2838), .Z(n2835) );
  NAND2_X1 U2815 ( .A1(a_12_), .A2(b_9_), .ZN(n2837) );
  NAND2_X1 U2816 ( .A1(a_11_), .A2(n2834), .ZN(n2724) );
  NAND2_X1 U2817 ( .A1(n2839), .A2(n2840), .ZN(n2834) );
  NAND3_X1 U2818 ( .A1(b_10_), .A2(n2841), .A3(a_12_), .ZN(n2840) );
  NAND2_X1 U2819 ( .A1(n2732), .A2(n2730), .ZN(n2841) );
  OR2_X1 U2820 ( .A1(n2730), .A2(n2732), .ZN(n2839) );
  AND2_X1 U2821 ( .A1(n2842), .A2(n2843), .ZN(n2732) );
  NAND2_X1 U2822 ( .A1(n2746), .A2(n2844), .ZN(n2843) );
  OR2_X1 U2823 ( .A1(n2747), .A2(n2748), .ZN(n2844) );
  NOR2_X1 U2824 ( .A1(n2655), .A2(n1952), .ZN(n2746) );
  NAND2_X1 U2825 ( .A1(n2748), .A2(n2747), .ZN(n2842) );
  NAND2_X1 U2826 ( .A1(n2845), .A2(n2846), .ZN(n2747) );
  NAND2_X1 U2827 ( .A1(b_8_), .A2(n2847), .ZN(n2846) );
  NAND2_X1 U2828 ( .A1(n1929), .A2(n2848), .ZN(n2847) );
  NAND2_X1 U2829 ( .A1(a_15_), .A2(n2010), .ZN(n2848) );
  NAND2_X1 U2830 ( .A1(b_9_), .A2(n2849), .ZN(n2845) );
  NAND2_X1 U2831 ( .A1(n1932), .A2(n2850), .ZN(n2849) );
  NAND2_X1 U2832 ( .A1(a_14_), .A2(n2175), .ZN(n2850) );
  AND3_X1 U2833 ( .A1(b_10_), .A2(n2173), .A3(b_9_), .ZN(n2748) );
  XNOR2_X1 U2834 ( .A(n2851), .B(n2852), .ZN(n2730) );
  XOR2_X1 U2835 ( .A(n2853), .B(n2854), .Z(n2851) );
  NOR2_X1 U2836 ( .A1(n2550), .A2(n2655), .ZN(n1993) );
  INV_X1 U2837 ( .A(b_10_), .ZN(n2655) );
  XNOR2_X1 U2838 ( .A(n2855), .B(n2856), .ZN(n2753) );
  NAND2_X1 U2839 ( .A1(n2857), .A2(n2858), .ZN(n2855) );
  XNOR2_X1 U2840 ( .A(n2859), .B(n2860), .ZN(n2757) );
  XNOR2_X1 U2841 ( .A(n2861), .B(n2158), .ZN(n2859) );
  INV_X1 U2842 ( .A(n2005), .ZN(n2158) );
  XNOR2_X1 U2843 ( .A(n2862), .B(n2863), .ZN(n2760) );
  XNOR2_X1 U2844 ( .A(n2864), .B(n2865), .ZN(n2862) );
  NOR2_X1 U2845 ( .A1(n2010), .A2(n2176), .ZN(n2865) );
  XNOR2_X1 U2846 ( .A(n2866), .B(n2867), .ZN(n2764) );
  XNOR2_X1 U2847 ( .A(n2868), .B(n2869), .ZN(n2867) );
  XNOR2_X1 U2848 ( .A(n2870), .B(n2871), .ZN(n2769) );
  XNOR2_X1 U2849 ( .A(n2872), .B(n2873), .ZN(n2871) );
  XNOR2_X1 U2850 ( .A(n2874), .B(n2875), .ZN(n2772) );
  XNOR2_X1 U2851 ( .A(n2876), .B(n2877), .ZN(n2874) );
  NOR2_X1 U2852 ( .A1(n2066), .A2(n2010), .ZN(n2877) );
  XNOR2_X1 U2853 ( .A(n2878), .B(n2879), .ZN(n2777) );
  NAND2_X1 U2854 ( .A1(n2880), .A2(n2881), .ZN(n2878) );
  XOR2_X1 U2855 ( .A(n2882), .B(n2883), .Z(n2781) );
  XNOR2_X1 U2856 ( .A(n2884), .B(n2885), .ZN(n2882) );
  NAND2_X1 U2857 ( .A1(a_3_), .A2(b_9_), .ZN(n2884) );
  XOR2_X1 U2858 ( .A(n2886), .B(n2887), .Z(n2589) );
  XNOR2_X1 U2859 ( .A(n2888), .B(n2889), .ZN(n2887) );
  NAND2_X1 U2860 ( .A1(a_2_), .A2(b_9_), .ZN(n2889) );
  XOR2_X1 U2861 ( .A(n2890), .B(n2891), .Z(n2234) );
  XNOR2_X1 U2862 ( .A(n2892), .B(n2893), .ZN(n2891) );
  NAND2_X1 U2863 ( .A1(a_0_), .A2(b_9_), .ZN(n2893) );
  NAND2_X1 U2864 ( .A1(n2894), .A2(n2895), .ZN(n1892) );
  NAND2_X1 U2865 ( .A1(n2787), .A2(n2786), .ZN(n2895) );
  XNOR2_X1 U2866 ( .A(n2896), .B(n2897), .ZN(n2894) );
  NAND3_X1 U2867 ( .A1(n2898), .A2(n2786), .A3(n2787), .ZN(n1891) );
  XNOR2_X1 U2868 ( .A(n2899), .B(n2900), .ZN(n2787) );
  NAND2_X1 U2869 ( .A1(n2901), .A2(n2902), .ZN(n2899) );
  NAND2_X1 U2870 ( .A1(n2903), .A2(n2904), .ZN(n2786) );
  NAND3_X1 U2871 ( .A1(b_9_), .A2(n2905), .A3(a_0_), .ZN(n2904) );
  NAND2_X1 U2872 ( .A1(n2892), .A2(n2890), .ZN(n2905) );
  OR2_X1 U2873 ( .A1(n2890), .A2(n2892), .ZN(n2903) );
  AND2_X1 U2874 ( .A1(n2906), .A2(n2907), .ZN(n2892) );
  NAND3_X1 U2875 ( .A1(b_9_), .A2(n2908), .A3(a_1_), .ZN(n2907) );
  OR2_X1 U2876 ( .A1(n2793), .A2(n2795), .ZN(n2908) );
  NAND2_X1 U2877 ( .A1(n2793), .A2(n2795), .ZN(n2906) );
  NAND2_X1 U2878 ( .A1(n2909), .A2(n2910), .ZN(n2795) );
  NAND3_X1 U2879 ( .A1(b_9_), .A2(n2911), .A3(a_2_), .ZN(n2910) );
  NAND2_X1 U2880 ( .A1(n2888), .A2(n2886), .ZN(n2911) );
  OR2_X1 U2881 ( .A1(n2886), .A2(n2888), .ZN(n2909) );
  AND2_X1 U2882 ( .A1(n2912), .A2(n2913), .ZN(n2888) );
  NAND3_X1 U2883 ( .A1(b_9_), .A2(n2914), .A3(a_3_), .ZN(n2913) );
  OR2_X1 U2884 ( .A1(n2883), .A2(n2885), .ZN(n2914) );
  NAND2_X1 U2885 ( .A1(n2883), .A2(n2885), .ZN(n2912) );
  NAND2_X1 U2886 ( .A1(n2880), .A2(n2915), .ZN(n2885) );
  NAND2_X1 U2887 ( .A1(n2879), .A2(n2881), .ZN(n2915) );
  NAND2_X1 U2888 ( .A1(n2916), .A2(n2917), .ZN(n2881) );
  NAND2_X1 U2889 ( .A1(b_9_), .A2(a_4_), .ZN(n2917) );
  INV_X1 U2890 ( .A(n2918), .ZN(n2916) );
  XNOR2_X1 U2891 ( .A(n2919), .B(n2920), .ZN(n2879) );
  XNOR2_X1 U2892 ( .A(n2921), .B(n2922), .ZN(n2919) );
  NOR2_X1 U2893 ( .A1(n2066), .A2(n2175), .ZN(n2922) );
  NAND2_X1 U2894 ( .A1(a_4_), .A2(n2918), .ZN(n2880) );
  NAND2_X1 U2895 ( .A1(n2923), .A2(n2924), .ZN(n2918) );
  NAND3_X1 U2896 ( .A1(a_5_), .A2(n2925), .A3(b_9_), .ZN(n2924) );
  NAND2_X1 U2897 ( .A1(n2876), .A2(n2875), .ZN(n2925) );
  OR2_X1 U2898 ( .A1(n2875), .A2(n2876), .ZN(n2923) );
  AND2_X1 U2899 ( .A1(n2926), .A2(n2927), .ZN(n2876) );
  NAND2_X1 U2900 ( .A1(n2873), .A2(n2928), .ZN(n2927) );
  OR2_X1 U2901 ( .A1(n2872), .A2(n2870), .ZN(n2928) );
  NOR2_X1 U2902 ( .A1(n2056), .A2(n2010), .ZN(n2873) );
  NAND2_X1 U2903 ( .A1(n2870), .A2(n2872), .ZN(n2926) );
  NAND2_X1 U2904 ( .A1(n2929), .A2(n2930), .ZN(n2872) );
  NAND2_X1 U2905 ( .A1(n2869), .A2(n2931), .ZN(n2930) );
  OR2_X1 U2906 ( .A1(n2868), .A2(n2866), .ZN(n2931) );
  NOR2_X1 U2907 ( .A1(n2010), .A2(n2038), .ZN(n2869) );
  NAND2_X1 U2908 ( .A1(n2866), .A2(n2868), .ZN(n2929) );
  NAND2_X1 U2909 ( .A1(n2932), .A2(n2933), .ZN(n2868) );
  NAND3_X1 U2910 ( .A1(b_9_), .A2(n2934), .A3(a_8_), .ZN(n2933) );
  NAND2_X1 U2911 ( .A1(n2864), .A2(n2863), .ZN(n2934) );
  OR2_X1 U2912 ( .A1(n2863), .A2(n2864), .ZN(n2932) );
  AND2_X1 U2913 ( .A1(n2935), .A2(n2936), .ZN(n2864) );
  NAND2_X1 U2914 ( .A1(n2005), .A2(n2937), .ZN(n2936) );
  OR2_X1 U2915 ( .A1(n2860), .A2(n2861), .ZN(n2937) );
  NOR2_X1 U2916 ( .A1(n2010), .A2(n2008), .ZN(n2005) );
  NAND2_X1 U2917 ( .A1(n2860), .A2(n2861), .ZN(n2935) );
  NAND2_X1 U2918 ( .A1(n2857), .A2(n2938), .ZN(n2861) );
  NAND2_X1 U2919 ( .A1(n2856), .A2(n2858), .ZN(n2938) );
  NAND2_X1 U2920 ( .A1(n2939), .A2(n2940), .ZN(n2858) );
  NAND2_X1 U2921 ( .A1(a_10_), .A2(b_9_), .ZN(n2940) );
  INV_X1 U2922 ( .A(n2941), .ZN(n2939) );
  XNOR2_X1 U2923 ( .A(n2942), .B(n2943), .ZN(n2856) );
  NAND2_X1 U2924 ( .A1(n2944), .A2(n2945), .ZN(n2942) );
  NAND2_X1 U2925 ( .A1(a_10_), .A2(n2941), .ZN(n2857) );
  NAND2_X1 U2926 ( .A1(n2829), .A2(n2946), .ZN(n2941) );
  NAND2_X1 U2927 ( .A1(n2828), .A2(n2830), .ZN(n2946) );
  NAND2_X1 U2928 ( .A1(n2947), .A2(n2948), .ZN(n2830) );
  NAND2_X1 U2929 ( .A1(b_9_), .A2(a_11_), .ZN(n2948) );
  INV_X1 U2930 ( .A(n2949), .ZN(n2947) );
  XNOR2_X1 U2931 ( .A(n2950), .B(n2951), .ZN(n2828) );
  XOR2_X1 U2932 ( .A(n2952), .B(n2953), .Z(n2950) );
  NAND2_X1 U2933 ( .A1(a_12_), .A2(b_8_), .ZN(n2952) );
  NAND2_X1 U2934 ( .A1(a_11_), .A2(n2949), .ZN(n2829) );
  NAND2_X1 U2935 ( .A1(n2954), .A2(n2955), .ZN(n2949) );
  NAND3_X1 U2936 ( .A1(b_9_), .A2(n2956), .A3(a_12_), .ZN(n2955) );
  NAND2_X1 U2937 ( .A1(n2838), .A2(n2836), .ZN(n2956) );
  OR2_X1 U2938 ( .A1(n2836), .A2(n2838), .ZN(n2954) );
  AND2_X1 U2939 ( .A1(n2957), .A2(n2958), .ZN(n2838) );
  NAND2_X1 U2940 ( .A1(n2852), .A2(n2959), .ZN(n2958) );
  OR2_X1 U2941 ( .A1(n2853), .A2(n2854), .ZN(n2959) );
  NOR2_X1 U2942 ( .A1(n2010), .A2(n1952), .ZN(n2852) );
  INV_X1 U2943 ( .A(b_9_), .ZN(n2010) );
  NAND2_X1 U2944 ( .A1(n2854), .A2(n2853), .ZN(n2957) );
  NAND2_X1 U2945 ( .A1(n2960), .A2(n2961), .ZN(n2853) );
  NAND2_X1 U2946 ( .A1(b_7_), .A2(n2962), .ZN(n2961) );
  NAND2_X1 U2947 ( .A1(n1929), .A2(n2963), .ZN(n2962) );
  NAND2_X1 U2948 ( .A1(a_15_), .A2(n2175), .ZN(n2963) );
  NAND2_X1 U2949 ( .A1(b_8_), .A2(n2964), .ZN(n2960) );
  NAND2_X1 U2950 ( .A1(n1932), .A2(n2965), .ZN(n2964) );
  NAND2_X1 U2951 ( .A1(a_14_), .A2(n2036), .ZN(n2965) );
  AND3_X1 U2952 ( .A1(b_9_), .A2(n2173), .A3(b_8_), .ZN(n2854) );
  XNOR2_X1 U2953 ( .A(n2966), .B(n2967), .ZN(n2836) );
  XOR2_X1 U2954 ( .A(n2968), .B(n2969), .Z(n2966) );
  XNOR2_X1 U2955 ( .A(n2970), .B(n2971), .ZN(n2860) );
  NAND2_X1 U2956 ( .A1(n2972), .A2(n2973), .ZN(n2970) );
  XNOR2_X1 U2957 ( .A(n2974), .B(n2975), .ZN(n2863) );
  XOR2_X1 U2958 ( .A(n2976), .B(n2977), .Z(n2974) );
  XOR2_X1 U2959 ( .A(n2978), .B(n2979), .Z(n2866) );
  XNOR2_X1 U2960 ( .A(n2980), .B(n2022), .ZN(n2978) );
  INV_X1 U2961 ( .A(n2981), .ZN(n2022) );
  XOR2_X1 U2962 ( .A(n2982), .B(n2983), .Z(n2870) );
  XOR2_X1 U2963 ( .A(n2984), .B(n2985), .Z(n2982) );
  NOR2_X1 U2964 ( .A1(n2038), .A2(n2175), .ZN(n2985) );
  XOR2_X1 U2965 ( .A(n2986), .B(n2987), .Z(n2875) );
  XOR2_X1 U2966 ( .A(n2988), .B(n2989), .Z(n2987) );
  NAND2_X1 U2967 ( .A1(a_6_), .A2(b_8_), .ZN(n2989) );
  XOR2_X1 U2968 ( .A(n2990), .B(n2991), .Z(n2883) );
  XNOR2_X1 U2969 ( .A(n2992), .B(n2993), .ZN(n2991) );
  NAND2_X1 U2970 ( .A1(b_8_), .A2(a_4_), .ZN(n2993) );
  XNOR2_X1 U2971 ( .A(n2994), .B(n2995), .ZN(n2886) );
  XOR2_X1 U2972 ( .A(n2996), .B(n2997), .Z(n2994) );
  XOR2_X1 U2973 ( .A(n2998), .B(n2999), .Z(n2793) );
  XOR2_X1 U2974 ( .A(n3000), .B(n3001), .Z(n2999) );
  XNOR2_X1 U2975 ( .A(n3002), .B(n3003), .ZN(n2890) );
  XOR2_X1 U2976 ( .A(n3004), .B(n3005), .Z(n3002) );
  XOR2_X1 U2977 ( .A(n2896), .B(n2897), .Z(n2898) );
  NAND2_X1 U2978 ( .A1(n3006), .A2(n3007), .ZN(n1897) );
  NAND2_X1 U2979 ( .A1(n2897), .A2(n2896), .ZN(n3007) );
  XNOR2_X1 U2980 ( .A(n3008), .B(n3009), .ZN(n3006) );
  NAND3_X1 U2981 ( .A1(n3010), .A2(n2896), .A3(n2897), .ZN(n1896) );
  XNOR2_X1 U2982 ( .A(n3011), .B(n3012), .ZN(n2897) );
  XOR2_X1 U2983 ( .A(n3013), .B(n3014), .Z(n3012) );
  NAND2_X1 U2984 ( .A1(a_0_), .A2(b_7_), .ZN(n3014) );
  NAND2_X1 U2985 ( .A1(n2901), .A2(n3015), .ZN(n2896) );
  NAND2_X1 U2986 ( .A1(n2900), .A2(n2902), .ZN(n3015) );
  NAND2_X1 U2987 ( .A1(n3016), .A2(n3017), .ZN(n2902) );
  NAND2_X1 U2988 ( .A1(a_0_), .A2(b_8_), .ZN(n3017) );
  INV_X1 U2989 ( .A(n3018), .ZN(n3016) );
  XNOR2_X1 U2990 ( .A(n3019), .B(n3020), .ZN(n2900) );
  XNOR2_X1 U2991 ( .A(n3021), .B(n3022), .ZN(n3019) );
  NOR2_X1 U2992 ( .A1(n2036), .A2(n2360), .ZN(n3022) );
  NAND2_X1 U2993 ( .A1(a_0_), .A2(n3018), .ZN(n2901) );
  NAND2_X1 U2994 ( .A1(n3023), .A2(n3024), .ZN(n3018) );
  NAND2_X1 U2995 ( .A1(n3005), .A2(n3025), .ZN(n3024) );
  OR2_X1 U2996 ( .A1(n3003), .A2(n3004), .ZN(n3025) );
  NOR2_X1 U2997 ( .A1(n2360), .A2(n2175), .ZN(n3005) );
  NAND2_X1 U2998 ( .A1(n3003), .A2(n3004), .ZN(n3023) );
  NAND2_X1 U2999 ( .A1(n3026), .A2(n3027), .ZN(n3004) );
  NAND2_X1 U3000 ( .A1(n3001), .A2(n3028), .ZN(n3027) );
  NAND2_X1 U3001 ( .A1(n3000), .A2(n2998), .ZN(n3028) );
  NOR2_X1 U3002 ( .A1(n2178), .A2(n2175), .ZN(n3001) );
  OR2_X1 U3003 ( .A1(n2998), .A2(n3000), .ZN(n3026) );
  AND2_X1 U3004 ( .A1(n3029), .A2(n3030), .ZN(n3000) );
  NAND2_X1 U3005 ( .A1(n2997), .A2(n3031), .ZN(n3030) );
  OR2_X1 U3006 ( .A1(n2995), .A2(n2996), .ZN(n3031) );
  NOR2_X1 U3007 ( .A1(n2100), .A2(n2175), .ZN(n2997) );
  NAND2_X1 U3008 ( .A1(n2995), .A2(n2996), .ZN(n3029) );
  NAND2_X1 U3009 ( .A1(n3032), .A2(n3033), .ZN(n2996) );
  NAND3_X1 U3010 ( .A1(a_4_), .A2(n3034), .A3(b_8_), .ZN(n3033) );
  NAND2_X1 U3011 ( .A1(n2992), .A2(n2990), .ZN(n3034) );
  OR2_X1 U3012 ( .A1(n2990), .A2(n2992), .ZN(n3032) );
  AND2_X1 U3013 ( .A1(n3035), .A2(n3036), .ZN(n2992) );
  NAND3_X1 U3014 ( .A1(a_5_), .A2(n3037), .A3(b_8_), .ZN(n3036) );
  NAND2_X1 U3015 ( .A1(n2921), .A2(n2920), .ZN(n3037) );
  OR2_X1 U3016 ( .A1(n2920), .A2(n2921), .ZN(n3035) );
  AND2_X1 U3017 ( .A1(n3038), .A2(n3039), .ZN(n2921) );
  NAND3_X1 U3018 ( .A1(b_8_), .A2(n3040), .A3(a_6_), .ZN(n3039) );
  OR2_X1 U3019 ( .A1(n2986), .A2(n2988), .ZN(n3040) );
  NAND2_X1 U3020 ( .A1(n2986), .A2(n2988), .ZN(n3038) );
  NAND2_X1 U3021 ( .A1(n3041), .A2(n3042), .ZN(n2988) );
  NAND3_X1 U3022 ( .A1(a_7_), .A2(n3043), .A3(b_8_), .ZN(n3042) );
  OR2_X1 U3023 ( .A1(n2983), .A2(n2984), .ZN(n3043) );
  NAND2_X1 U3024 ( .A1(n2983), .A2(n2984), .ZN(n3041) );
  NAND2_X1 U3025 ( .A1(n3044), .A2(n3045), .ZN(n2984) );
  NAND2_X1 U3026 ( .A1(n2979), .A2(n3046), .ZN(n3045) );
  OR2_X1 U3027 ( .A1(n2980), .A2(n2981), .ZN(n3046) );
  XNOR2_X1 U3028 ( .A(n3047), .B(n3048), .ZN(n2979) );
  XNOR2_X1 U3029 ( .A(n3049), .B(n3050), .ZN(n3047) );
  NAND2_X1 U3030 ( .A1(n2981), .A2(n2980), .ZN(n3044) );
  NAND2_X1 U3031 ( .A1(n3051), .A2(n3052), .ZN(n2980) );
  NAND2_X1 U3032 ( .A1(n2977), .A2(n3053), .ZN(n3052) );
  OR2_X1 U3033 ( .A1(n2975), .A2(n2976), .ZN(n3053) );
  NOR2_X1 U3034 ( .A1(n2175), .A2(n2008), .ZN(n2977) );
  NAND2_X1 U3035 ( .A1(n2975), .A2(n2976), .ZN(n3051) );
  NAND2_X1 U3036 ( .A1(n2972), .A2(n3054), .ZN(n2976) );
  NAND2_X1 U3037 ( .A1(n2971), .A2(n2973), .ZN(n3054) );
  NAND2_X1 U3038 ( .A1(n3055), .A2(n3056), .ZN(n2973) );
  NAND2_X1 U3039 ( .A1(a_10_), .A2(b_8_), .ZN(n3056) );
  INV_X1 U3040 ( .A(n3057), .ZN(n3055) );
  XNOR2_X1 U3041 ( .A(n3058), .B(n3059), .ZN(n2971) );
  NAND2_X1 U3042 ( .A1(n3060), .A2(n3061), .ZN(n3058) );
  NAND2_X1 U3043 ( .A1(a_10_), .A2(n3057), .ZN(n2972) );
  NAND2_X1 U3044 ( .A1(n2944), .A2(n3062), .ZN(n3057) );
  NAND2_X1 U3045 ( .A1(n2943), .A2(n2945), .ZN(n3062) );
  NAND2_X1 U3046 ( .A1(n3063), .A2(n3064), .ZN(n2945) );
  NAND2_X1 U3047 ( .A1(b_8_), .A2(a_11_), .ZN(n3064) );
  INV_X1 U3048 ( .A(n3065), .ZN(n3063) );
  XNOR2_X1 U3049 ( .A(n3066), .B(n3067), .ZN(n2943) );
  XOR2_X1 U3050 ( .A(n3068), .B(n3069), .Z(n3066) );
  NAND2_X1 U3051 ( .A1(b_7_), .A2(a_12_), .ZN(n3068) );
  NAND2_X1 U3052 ( .A1(a_11_), .A2(n3065), .ZN(n2944) );
  NAND2_X1 U3053 ( .A1(n3070), .A2(n3071), .ZN(n3065) );
  NAND3_X1 U3054 ( .A1(b_8_), .A2(n3072), .A3(a_12_), .ZN(n3071) );
  NAND2_X1 U3055 ( .A1(n2953), .A2(n2951), .ZN(n3072) );
  OR2_X1 U3056 ( .A1(n2951), .A2(n2953), .ZN(n3070) );
  AND2_X1 U3057 ( .A1(n3073), .A2(n3074), .ZN(n2953) );
  NAND2_X1 U3058 ( .A1(n2967), .A2(n3075), .ZN(n3074) );
  OR2_X1 U3059 ( .A1(n2968), .A2(n2969), .ZN(n3075) );
  NOR2_X1 U3060 ( .A1(n2175), .A2(n1952), .ZN(n2967) );
  NAND2_X1 U3061 ( .A1(n2969), .A2(n2968), .ZN(n3073) );
  NAND2_X1 U3062 ( .A1(n3076), .A2(n3077), .ZN(n2968) );
  NAND2_X1 U3063 ( .A1(b_6_), .A2(n3078), .ZN(n3077) );
  NAND2_X1 U3064 ( .A1(n1929), .A2(n3079), .ZN(n3078) );
  NAND2_X1 U3065 ( .A1(a_15_), .A2(n2036), .ZN(n3079) );
  NAND2_X1 U3066 ( .A1(b_7_), .A2(n3080), .ZN(n3076) );
  NAND2_X1 U3067 ( .A1(n1932), .A2(n3081), .ZN(n3080) );
  NAND2_X1 U3068 ( .A1(a_14_), .A2(n3082), .ZN(n3081) );
  AND3_X1 U3069 ( .A1(b_8_), .A2(n2173), .A3(b_7_), .ZN(n2969) );
  XNOR2_X1 U3070 ( .A(n3083), .B(n3084), .ZN(n2951) );
  XOR2_X1 U3071 ( .A(n3085), .B(n3086), .Z(n3083) );
  XNOR2_X1 U3072 ( .A(n3087), .B(n3088), .ZN(n2975) );
  NAND2_X1 U3073 ( .A1(n3089), .A2(n3090), .ZN(n3087) );
  NOR2_X1 U3074 ( .A1(n2176), .A2(n2175), .ZN(n2981) );
  INV_X1 U3075 ( .A(b_8_), .ZN(n2175) );
  XNOR2_X1 U3076 ( .A(n3091), .B(n3092), .ZN(n2983) );
  XNOR2_X1 U3077 ( .A(n3093), .B(n3094), .ZN(n3091) );
  NOR2_X1 U3078 ( .A1(n2036), .A2(n2176), .ZN(n3094) );
  XOR2_X1 U3079 ( .A(n3095), .B(n3096), .Z(n2986) );
  XNOR2_X1 U3080 ( .A(n3097), .B(n2154), .ZN(n3095) );
  INV_X1 U3081 ( .A(n2034), .ZN(n2154) );
  XOR2_X1 U3082 ( .A(n3098), .B(n3099), .Z(n2920) );
  XOR2_X1 U3083 ( .A(n3100), .B(n3101), .Z(n3099) );
  NAND2_X1 U3084 ( .A1(a_6_), .A2(b_7_), .ZN(n3101) );
  XOR2_X1 U3085 ( .A(n3102), .B(n3103), .Z(n2990) );
  XOR2_X1 U3086 ( .A(n3104), .B(n3105), .Z(n3103) );
  NAND2_X1 U3087 ( .A1(b_7_), .A2(a_5_), .ZN(n3105) );
  XOR2_X1 U3088 ( .A(n3106), .B(n3107), .Z(n2995) );
  XOR2_X1 U3089 ( .A(n3108), .B(n3109), .Z(n3106) );
  NOR2_X1 U3090 ( .A1(n2347), .A2(n2036), .ZN(n3109) );
  XOR2_X1 U3091 ( .A(n3110), .B(n3111), .Z(n2998) );
  XOR2_X1 U3092 ( .A(n3112), .B(n3113), .Z(n3111) );
  NAND2_X1 U3093 ( .A1(a_3_), .A2(b_7_), .ZN(n3113) );
  XOR2_X1 U3094 ( .A(n3114), .B(n3115), .Z(n3003) );
  XOR2_X1 U3095 ( .A(n3116), .B(n3117), .Z(n3114) );
  NOR2_X1 U3096 ( .A1(n2036), .A2(n2178), .ZN(n3117) );
  XOR2_X1 U3097 ( .A(n3008), .B(n3009), .Z(n3010) );
  NAND2_X1 U3098 ( .A1(n3118), .A2(n3119), .ZN(n1902) );
  NAND2_X1 U3099 ( .A1(n3009), .A2(n3008), .ZN(n3119) );
  XNOR2_X1 U3100 ( .A(n3120), .B(n3121), .ZN(n3118) );
  NAND3_X1 U3101 ( .A1(n3122), .A2(n3008), .A3(n3009), .ZN(n1901) );
  XNOR2_X1 U3102 ( .A(n3123), .B(n3124), .ZN(n3009) );
  XOR2_X1 U3103 ( .A(n3125), .B(n3126), .Z(n3124) );
  NAND2_X1 U3104 ( .A1(a_0_), .A2(b_6_), .ZN(n3126) );
  NAND2_X1 U3105 ( .A1(n3127), .A2(n3128), .ZN(n3008) );
  NAND3_X1 U3106 ( .A1(b_7_), .A2(n3129), .A3(a_0_), .ZN(n3128) );
  OR2_X1 U3107 ( .A1(n3011), .A2(n3013), .ZN(n3129) );
  NAND2_X1 U3108 ( .A1(n3011), .A2(n3013), .ZN(n3127) );
  NAND2_X1 U3109 ( .A1(n3130), .A2(n3131), .ZN(n3013) );
  NAND3_X1 U3110 ( .A1(b_7_), .A2(n3132), .A3(a_1_), .ZN(n3131) );
  NAND2_X1 U3111 ( .A1(n3020), .A2(n3021), .ZN(n3132) );
  OR2_X1 U3112 ( .A1(n3020), .A2(n3021), .ZN(n3130) );
  AND2_X1 U3113 ( .A1(n3133), .A2(n3134), .ZN(n3021) );
  NAND3_X1 U3114 ( .A1(b_7_), .A2(n3135), .A3(a_2_), .ZN(n3134) );
  OR2_X1 U3115 ( .A1(n3116), .A2(n3115), .ZN(n3135) );
  NAND2_X1 U3116 ( .A1(n3115), .A2(n3116), .ZN(n3133) );
  NAND2_X1 U3117 ( .A1(n3136), .A2(n3137), .ZN(n3116) );
  NAND3_X1 U3118 ( .A1(b_7_), .A2(n3138), .A3(a_3_), .ZN(n3137) );
  OR2_X1 U3119 ( .A1(n3110), .A2(n3112), .ZN(n3138) );
  NAND2_X1 U3120 ( .A1(n3110), .A2(n3112), .ZN(n3136) );
  NAND2_X1 U3121 ( .A1(n3139), .A2(n3140), .ZN(n3112) );
  NAND3_X1 U3122 ( .A1(a_4_), .A2(n3141), .A3(b_7_), .ZN(n3140) );
  OR2_X1 U3123 ( .A1(n3108), .A2(n3107), .ZN(n3141) );
  NAND2_X1 U3124 ( .A1(n3107), .A2(n3108), .ZN(n3139) );
  NAND2_X1 U3125 ( .A1(n3142), .A2(n3143), .ZN(n3108) );
  NAND3_X1 U3126 ( .A1(a_5_), .A2(n3144), .A3(b_7_), .ZN(n3143) );
  OR2_X1 U3127 ( .A1(n3102), .A2(n3104), .ZN(n3144) );
  NAND2_X1 U3128 ( .A1(n3102), .A2(n3104), .ZN(n3142) );
  NAND2_X1 U3129 ( .A1(n3145), .A2(n3146), .ZN(n3104) );
  NAND3_X1 U3130 ( .A1(b_7_), .A2(n3147), .A3(a_6_), .ZN(n3146) );
  OR2_X1 U3131 ( .A1(n3098), .A2(n3100), .ZN(n3147) );
  NAND2_X1 U3132 ( .A1(n3098), .A2(n3100), .ZN(n3145) );
  NAND2_X1 U3133 ( .A1(n3148), .A2(n3149), .ZN(n3100) );
  NAND2_X1 U3134 ( .A1(n3096), .A2(n3150), .ZN(n3149) );
  OR2_X1 U3135 ( .A1(n3097), .A2(n2034), .ZN(n3150) );
  XNOR2_X1 U3136 ( .A(n3151), .B(n3152), .ZN(n3096) );
  XNOR2_X1 U3137 ( .A(n3153), .B(n3154), .ZN(n3151) );
  NOR2_X1 U3138 ( .A1(n3082), .A2(n2176), .ZN(n3154) );
  NAND2_X1 U3139 ( .A1(n2034), .A2(n3097), .ZN(n3148) );
  NAND2_X1 U3140 ( .A1(n3155), .A2(n3156), .ZN(n3097) );
  NAND3_X1 U3141 ( .A1(b_7_), .A2(n3157), .A3(a_8_), .ZN(n3156) );
  NAND2_X1 U3142 ( .A1(n3093), .A2(n3092), .ZN(n3157) );
  OR2_X1 U3143 ( .A1(n3092), .A2(n3093), .ZN(n3155) );
  AND2_X1 U3144 ( .A1(n3158), .A2(n3159), .ZN(n3093) );
  NAND2_X1 U3145 ( .A1(n3050), .A2(n3160), .ZN(n3159) );
  NAND2_X1 U3146 ( .A1(n3049), .A2(n3048), .ZN(n3160) );
  NOR2_X1 U3147 ( .A1(n2036), .A2(n2008), .ZN(n3050) );
  OR2_X1 U3148 ( .A1(n3048), .A2(n3049), .ZN(n3158) );
  AND2_X1 U3149 ( .A1(n3089), .A2(n3161), .ZN(n3049) );
  NAND2_X1 U3150 ( .A1(n3088), .A2(n3090), .ZN(n3161) );
  NAND2_X1 U3151 ( .A1(n3162), .A2(n3163), .ZN(n3090) );
  NAND2_X1 U3152 ( .A1(a_10_), .A2(b_7_), .ZN(n3163) );
  INV_X1 U3153 ( .A(n3164), .ZN(n3162) );
  XNOR2_X1 U3154 ( .A(n3165), .B(n3166), .ZN(n3088) );
  NAND2_X1 U3155 ( .A1(n3167), .A2(n3168), .ZN(n3165) );
  NAND2_X1 U3156 ( .A1(a_10_), .A2(n3164), .ZN(n3089) );
  NAND2_X1 U3157 ( .A1(n3060), .A2(n3169), .ZN(n3164) );
  NAND2_X1 U3158 ( .A1(n3059), .A2(n3061), .ZN(n3169) );
  NAND2_X1 U3159 ( .A1(n3170), .A2(n3171), .ZN(n3061) );
  NAND2_X1 U3160 ( .A1(b_7_), .A2(a_11_), .ZN(n3171) );
  INV_X1 U3161 ( .A(n3172), .ZN(n3170) );
  XNOR2_X1 U3162 ( .A(n3173), .B(n3174), .ZN(n3059) );
  XOR2_X1 U3163 ( .A(n3175), .B(n3176), .Z(n3173) );
  NAND2_X1 U3164 ( .A1(b_6_), .A2(a_12_), .ZN(n3175) );
  NAND2_X1 U3165 ( .A1(a_11_), .A2(n3172), .ZN(n3060) );
  NAND2_X1 U3166 ( .A1(n3177), .A2(n3178), .ZN(n3172) );
  NAND3_X1 U3167 ( .A1(a_12_), .A2(n3179), .A3(b_7_), .ZN(n3178) );
  NAND2_X1 U3168 ( .A1(n3069), .A2(n3067), .ZN(n3179) );
  OR2_X1 U3169 ( .A1(n3067), .A2(n3069), .ZN(n3177) );
  AND2_X1 U3170 ( .A1(n3180), .A2(n3181), .ZN(n3069) );
  NAND2_X1 U3171 ( .A1(n3084), .A2(n3182), .ZN(n3181) );
  OR2_X1 U3172 ( .A1(n3085), .A2(n3086), .ZN(n3182) );
  NOR2_X1 U3173 ( .A1(n2036), .A2(n1952), .ZN(n3084) );
  NAND2_X1 U3174 ( .A1(n3086), .A2(n3085), .ZN(n3180) );
  NAND2_X1 U3175 ( .A1(n3183), .A2(n3184), .ZN(n3085) );
  NAND2_X1 U3176 ( .A1(b_5_), .A2(n3185), .ZN(n3184) );
  NAND2_X1 U3177 ( .A1(n1929), .A2(n3186), .ZN(n3185) );
  NAND2_X1 U3178 ( .A1(a_15_), .A2(n3082), .ZN(n3186) );
  NAND2_X1 U3179 ( .A1(b_6_), .A2(n3187), .ZN(n3183) );
  NAND2_X1 U3180 ( .A1(n1932), .A2(n3188), .ZN(n3187) );
  NAND2_X1 U3181 ( .A1(a_14_), .A2(n2068), .ZN(n3188) );
  AND3_X1 U3182 ( .A1(b_7_), .A2(n2173), .A3(b_6_), .ZN(n3086) );
  XNOR2_X1 U3183 ( .A(n3189), .B(n3190), .ZN(n3067) );
  XOR2_X1 U3184 ( .A(n3191), .B(n3192), .Z(n3189) );
  XOR2_X1 U3185 ( .A(n3193), .B(n3194), .Z(n3048) );
  NAND2_X1 U3186 ( .A1(n3195), .A2(n3196), .ZN(n3193) );
  XOR2_X1 U3187 ( .A(n3197), .B(n3198), .Z(n3092) );
  NAND2_X1 U3188 ( .A1(n3199), .A2(n3200), .ZN(n3197) );
  NOR2_X1 U3189 ( .A1(n2036), .A2(n2038), .ZN(n2034) );
  INV_X1 U3190 ( .A(b_7_), .ZN(n2036) );
  XOR2_X1 U3191 ( .A(n3201), .B(n3202), .Z(n3098) );
  XOR2_X1 U3192 ( .A(n3203), .B(n3204), .Z(n3201) );
  NOR2_X1 U3193 ( .A1(n2038), .A2(n3082), .ZN(n3204) );
  XOR2_X1 U3194 ( .A(n3205), .B(n3206), .Z(n3102) );
  XNOR2_X1 U3195 ( .A(n2050), .B(n3207), .ZN(n3206) );
  XOR2_X1 U3196 ( .A(n3208), .B(n3209), .Z(n3107) );
  NOR2_X1 U3197 ( .A1(n3210), .A2(n3211), .ZN(n3209) );
  NOR2_X1 U3198 ( .A1(n3212), .A2(n3213), .ZN(n3210) );
  NOR2_X1 U3199 ( .A1(n2066), .A2(n3082), .ZN(n3213) );
  INV_X1 U3200 ( .A(n3214), .ZN(n3212) );
  XOR2_X1 U3201 ( .A(n3215), .B(n3216), .Z(n3110) );
  XOR2_X1 U3202 ( .A(n3217), .B(n3218), .Z(n3216) );
  XNOR2_X1 U3203 ( .A(n3219), .B(n3220), .ZN(n3115) );
  NAND2_X1 U3204 ( .A1(n3221), .A2(n3222), .ZN(n3219) );
  XNOR2_X1 U3205 ( .A(n3223), .B(n3224), .ZN(n3020) );
  XNOR2_X1 U3206 ( .A(n3225), .B(n3226), .ZN(n3223) );
  NAND2_X1 U3207 ( .A1(a_2_), .A2(b_6_), .ZN(n3225) );
  XOR2_X1 U3208 ( .A(n3227), .B(n3228), .Z(n3011) );
  XOR2_X1 U3209 ( .A(n3229), .B(n3230), .Z(n3228) );
  XOR2_X1 U3210 ( .A(n3120), .B(n3121), .Z(n3122) );
  NAND2_X1 U3211 ( .A1(n3231), .A2(n3232), .ZN(n1907) );
  NAND2_X1 U3212 ( .A1(n3121), .A2(n3120), .ZN(n3232) );
  XNOR2_X1 U3213 ( .A(n3233), .B(n3234), .ZN(n3231) );
  NAND3_X1 U3214 ( .A1(n3121), .A2(n3120), .A3(n3235), .ZN(n1906) );
  XNOR2_X1 U3215 ( .A(n3233), .B(n3236), .ZN(n3235) );
  INV_X1 U3216 ( .A(n3234), .ZN(n3236) );
  NAND2_X1 U3217 ( .A1(n3237), .A2(n3238), .ZN(n3120) );
  NAND3_X1 U3218 ( .A1(b_6_), .A2(n3239), .A3(a_0_), .ZN(n3238) );
  OR2_X1 U3219 ( .A1(n3123), .A2(n3125), .ZN(n3239) );
  NAND2_X1 U3220 ( .A1(n3123), .A2(n3125), .ZN(n3237) );
  NAND2_X1 U3221 ( .A1(n3240), .A2(n3241), .ZN(n3125) );
  NAND2_X1 U3222 ( .A1(n3230), .A2(n3242), .ZN(n3241) );
  NAND2_X1 U3223 ( .A1(n3229), .A2(n3227), .ZN(n3242) );
  NOR2_X1 U3224 ( .A1(n2360), .A2(n3082), .ZN(n3230) );
  OR2_X1 U3225 ( .A1(n3227), .A2(n3229), .ZN(n3240) );
  AND2_X1 U3226 ( .A1(n3243), .A2(n3244), .ZN(n3229) );
  NAND3_X1 U3227 ( .A1(b_6_), .A2(n3245), .A3(a_2_), .ZN(n3244) );
  OR2_X1 U3228 ( .A1(n3226), .A2(n3224), .ZN(n3245) );
  NAND2_X1 U3229 ( .A1(n3224), .A2(n3226), .ZN(n3243) );
  NAND2_X1 U3230 ( .A1(n3221), .A2(n3246), .ZN(n3226) );
  NAND2_X1 U3231 ( .A1(n3220), .A2(n3222), .ZN(n3246) );
  NAND2_X1 U3232 ( .A1(n3247), .A2(n3248), .ZN(n3222) );
  NAND2_X1 U3233 ( .A1(a_3_), .A2(b_6_), .ZN(n3248) );
  INV_X1 U3234 ( .A(n3249), .ZN(n3247) );
  XNOR2_X1 U3235 ( .A(n3250), .B(n3251), .ZN(n3220) );
  XNOR2_X1 U3236 ( .A(n3252), .B(n3253), .ZN(n3250) );
  NOR2_X1 U3237 ( .A1(n2347), .A2(n2068), .ZN(n3253) );
  NAND2_X1 U3238 ( .A1(a_3_), .A2(n3249), .ZN(n3221) );
  NAND2_X1 U3239 ( .A1(n3254), .A2(n3255), .ZN(n3249) );
  NAND2_X1 U3240 ( .A1(n3218), .A2(n3256), .ZN(n3255) );
  NAND2_X1 U3241 ( .A1(n3217), .A2(n3215), .ZN(n3256) );
  NOR2_X1 U3242 ( .A1(n3082), .A2(n2347), .ZN(n3218) );
  OR2_X1 U3243 ( .A1(n3215), .A2(n3217), .ZN(n3254) );
  NOR2_X1 U3244 ( .A1(n3211), .A2(n3257), .ZN(n3217) );
  AND2_X1 U3245 ( .A1(n3208), .A2(n3258), .ZN(n3257) );
  NAND2_X1 U3246 ( .A1(n3214), .A2(n3259), .ZN(n3258) );
  NAND2_X1 U3247 ( .A1(b_6_), .A2(a_5_), .ZN(n3259) );
  XNOR2_X1 U3248 ( .A(n3260), .B(n3261), .ZN(n3208) );
  XOR2_X1 U3249 ( .A(n3262), .B(n3263), .Z(n3261) );
  NAND2_X1 U3250 ( .A1(a_6_), .A2(b_5_), .ZN(n3263) );
  NOR2_X1 U3251 ( .A1(n3214), .A2(n2066), .ZN(n3211) );
  NAND2_X1 U3252 ( .A1(n3264), .A2(n3265), .ZN(n3214) );
  NAND2_X1 U3253 ( .A1(n3205), .A2(n3266), .ZN(n3265) );
  NAND2_X1 U3254 ( .A1(n2050), .A2(n3207), .ZN(n3266) );
  XNOR2_X1 U3255 ( .A(n3267), .B(n3268), .ZN(n3205) );
  XOR2_X1 U3256 ( .A(n3269), .B(n3270), .Z(n3267) );
  NOR2_X1 U3257 ( .A1(n2038), .A2(n2068), .ZN(n3270) );
  OR2_X1 U3258 ( .A1(n3207), .A2(n2050), .ZN(n3264) );
  NOR2_X1 U3259 ( .A1(n2056), .A2(n3082), .ZN(n2050) );
  NAND2_X1 U3260 ( .A1(n3271), .A2(n3272), .ZN(n3207) );
  NAND3_X1 U3261 ( .A1(a_7_), .A2(n3273), .A3(b_6_), .ZN(n3272) );
  OR2_X1 U3262 ( .A1(n3203), .A2(n3202), .ZN(n3273) );
  NAND2_X1 U3263 ( .A1(n3202), .A2(n3203), .ZN(n3271) );
  NAND2_X1 U3264 ( .A1(n3274), .A2(n3275), .ZN(n3203) );
  NAND3_X1 U3265 ( .A1(b_6_), .A2(n3276), .A3(a_8_), .ZN(n3275) );
  NAND2_X1 U3266 ( .A1(n3152), .A2(n3153), .ZN(n3276) );
  OR2_X1 U3267 ( .A1(n3152), .A2(n3153), .ZN(n3274) );
  AND2_X1 U3268 ( .A1(n3199), .A2(n3277), .ZN(n3153) );
  NAND2_X1 U3269 ( .A1(n3198), .A2(n3200), .ZN(n3277) );
  NAND2_X1 U3270 ( .A1(n3278), .A2(n3279), .ZN(n3200) );
  NAND2_X1 U3271 ( .A1(b_6_), .A2(a_9_), .ZN(n3279) );
  INV_X1 U3272 ( .A(n3280), .ZN(n3278) );
  XNOR2_X1 U3273 ( .A(n3281), .B(n3282), .ZN(n3198) );
  XNOR2_X1 U3274 ( .A(n3283), .B(n3284), .ZN(n3282) );
  NAND2_X1 U3275 ( .A1(a_9_), .A2(n3280), .ZN(n3199) );
  NAND2_X1 U3276 ( .A1(n3195), .A2(n3285), .ZN(n3280) );
  NAND2_X1 U3277 ( .A1(n3194), .A2(n3196), .ZN(n3285) );
  NAND2_X1 U3278 ( .A1(n3286), .A2(n3287), .ZN(n3196) );
  NAND2_X1 U3279 ( .A1(b_6_), .A2(a_10_), .ZN(n3287) );
  INV_X1 U3280 ( .A(n3288), .ZN(n3286) );
  XNOR2_X1 U3281 ( .A(n3289), .B(n3290), .ZN(n3194) );
  XNOR2_X1 U3282 ( .A(n3291), .B(n3292), .ZN(n3289) );
  NAND2_X1 U3283 ( .A1(a_10_), .A2(n3288), .ZN(n3195) );
  NAND2_X1 U3284 ( .A1(n3167), .A2(n3293), .ZN(n3288) );
  NAND2_X1 U3285 ( .A1(n3166), .A2(n3168), .ZN(n3293) );
  NAND2_X1 U3286 ( .A1(n3294), .A2(n3295), .ZN(n3168) );
  NAND2_X1 U3287 ( .A1(b_6_), .A2(a_11_), .ZN(n3295) );
  INV_X1 U3288 ( .A(n3296), .ZN(n3294) );
  XNOR2_X1 U3289 ( .A(n3297), .B(n3298), .ZN(n3166) );
  XOR2_X1 U3290 ( .A(n3299), .B(n3300), .Z(n3297) );
  NAND2_X1 U3291 ( .A1(b_5_), .A2(a_12_), .ZN(n3299) );
  NAND2_X1 U3292 ( .A1(a_11_), .A2(n3296), .ZN(n3167) );
  NAND2_X1 U3293 ( .A1(n3301), .A2(n3302), .ZN(n3296) );
  NAND3_X1 U3294 ( .A1(a_12_), .A2(n3303), .A3(b_6_), .ZN(n3302) );
  NAND2_X1 U3295 ( .A1(n3176), .A2(n3174), .ZN(n3303) );
  OR2_X1 U3296 ( .A1(n3174), .A2(n3176), .ZN(n3301) );
  AND2_X1 U3297 ( .A1(n3304), .A2(n3305), .ZN(n3176) );
  NAND2_X1 U3298 ( .A1(n3190), .A2(n3306), .ZN(n3305) );
  OR2_X1 U3299 ( .A1(n3191), .A2(n3192), .ZN(n3306) );
  NOR2_X1 U3300 ( .A1(n3082), .A2(n1952), .ZN(n3190) );
  INV_X1 U3301 ( .A(b_6_), .ZN(n3082) );
  NAND2_X1 U3302 ( .A1(n3192), .A2(n3191), .ZN(n3304) );
  NAND2_X1 U3303 ( .A1(n3307), .A2(n3308), .ZN(n3191) );
  NAND2_X1 U3304 ( .A1(b_4_), .A2(n3309), .ZN(n3308) );
  NAND2_X1 U3305 ( .A1(n1929), .A2(n3310), .ZN(n3309) );
  NAND2_X1 U3306 ( .A1(a_15_), .A2(n2068), .ZN(n3310) );
  NAND2_X1 U3307 ( .A1(b_5_), .A2(n3311), .ZN(n3307) );
  NAND2_X1 U3308 ( .A1(n1932), .A2(n3312), .ZN(n3311) );
  NAND2_X1 U3309 ( .A1(a_14_), .A2(n3313), .ZN(n3312) );
  AND3_X1 U3310 ( .A1(b_6_), .A2(n2173), .A3(b_5_), .ZN(n3192) );
  XNOR2_X1 U3311 ( .A(n3314), .B(n3315), .ZN(n3174) );
  XOR2_X1 U3312 ( .A(n3316), .B(n3317), .Z(n3314) );
  XOR2_X1 U3313 ( .A(n3318), .B(n3319), .Z(n3152) );
  NAND2_X1 U3314 ( .A1(n3320), .A2(n3321), .ZN(n3318) );
  XOR2_X1 U3315 ( .A(n3322), .B(n3323), .Z(n3202) );
  XNOR2_X1 U3316 ( .A(n3324), .B(n3325), .ZN(n3322) );
  NAND2_X1 U3317 ( .A1(a_8_), .A2(b_5_), .ZN(n3324) );
  XNOR2_X1 U3318 ( .A(n3326), .B(n3327), .ZN(n3215) );
  XNOR2_X1 U3319 ( .A(n3328), .B(n2150), .ZN(n3326) );
  INV_X1 U3320 ( .A(n2063), .ZN(n2150) );
  XNOR2_X1 U3321 ( .A(n3329), .B(n3330), .ZN(n3224) );
  XNOR2_X1 U3322 ( .A(n3331), .B(n3332), .ZN(n3329) );
  NOR2_X1 U3323 ( .A1(n2068), .A2(n2100), .ZN(n3332) );
  XNOR2_X1 U3324 ( .A(n3333), .B(n3334), .ZN(n3227) );
  XOR2_X1 U3325 ( .A(n3335), .B(n3336), .Z(n3333) );
  NOR2_X1 U3326 ( .A1(n2068), .A2(n2178), .ZN(n3336) );
  XOR2_X1 U3327 ( .A(n3337), .B(n3338), .Z(n3123) );
  XNOR2_X1 U3328 ( .A(n3339), .B(n3340), .ZN(n3338) );
  NAND2_X1 U3329 ( .A1(a_1_), .A2(b_5_), .ZN(n3340) );
  XOR2_X1 U3330 ( .A(n3341), .B(n3342), .Z(n3121) );
  XOR2_X1 U3331 ( .A(n3343), .B(n3344), .Z(n3341) );
  NOR2_X1 U3332 ( .A1(n2068), .A2(n2371), .ZN(n3344) );
  NAND2_X1 U3333 ( .A1(n3345), .A2(n3346), .ZN(n1912) );
  NAND2_X1 U3334 ( .A1(n3234), .A2(n3233), .ZN(n3346) );
  XNOR2_X1 U3335 ( .A(n3347), .B(n3348), .ZN(n3345) );
  NAND3_X1 U3336 ( .A1(n3234), .A2(n3233), .A3(n3349), .ZN(n1911) );
  XOR2_X1 U3337 ( .A(n3347), .B(n3348), .Z(n3349) );
  NAND2_X1 U3338 ( .A1(n3350), .A2(n3351), .ZN(n3233) );
  NAND3_X1 U3339 ( .A1(b_5_), .A2(n3352), .A3(a_0_), .ZN(n3351) );
  OR2_X1 U3340 ( .A1(n3342), .A2(n3343), .ZN(n3352) );
  NAND2_X1 U3341 ( .A1(n3342), .A2(n3343), .ZN(n3350) );
  NAND2_X1 U3342 ( .A1(n3353), .A2(n3354), .ZN(n3343) );
  NAND3_X1 U3343 ( .A1(b_5_), .A2(n3355), .A3(a_1_), .ZN(n3354) );
  NAND2_X1 U3344 ( .A1(n3339), .A2(n3337), .ZN(n3355) );
  OR2_X1 U3345 ( .A1(n3337), .A2(n3339), .ZN(n3353) );
  AND2_X1 U3346 ( .A1(n3356), .A2(n3357), .ZN(n3339) );
  NAND3_X1 U3347 ( .A1(b_5_), .A2(n3358), .A3(a_2_), .ZN(n3357) );
  OR2_X1 U3348 ( .A1(n3334), .A2(n3335), .ZN(n3358) );
  NAND2_X1 U3349 ( .A1(n3334), .A2(n3335), .ZN(n3356) );
  NAND2_X1 U3350 ( .A1(n3359), .A2(n3360), .ZN(n3335) );
  NAND3_X1 U3351 ( .A1(b_5_), .A2(n3361), .A3(a_3_), .ZN(n3360) );
  NAND2_X1 U3352 ( .A1(n3330), .A2(n3331), .ZN(n3361) );
  OR2_X1 U3353 ( .A1(n3330), .A2(n3331), .ZN(n3359) );
  AND2_X1 U3354 ( .A1(n3362), .A2(n3363), .ZN(n3331) );
  NAND3_X1 U3355 ( .A1(a_4_), .A2(n3364), .A3(b_5_), .ZN(n3363) );
  NAND2_X1 U3356 ( .A1(n3251), .A2(n3252), .ZN(n3364) );
  OR2_X1 U3357 ( .A1(n3251), .A2(n3252), .ZN(n3362) );
  AND2_X1 U3358 ( .A1(n3365), .A2(n3366), .ZN(n3252) );
  NAND2_X1 U3359 ( .A1(n3327), .A2(n3367), .ZN(n3366) );
  OR2_X1 U3360 ( .A1(n3328), .A2(n2063), .ZN(n3367) );
  XNOR2_X1 U3361 ( .A(n3368), .B(n3369), .ZN(n3327) );
  XOR2_X1 U3362 ( .A(n3370), .B(n3371), .Z(n3369) );
  NAND2_X1 U3363 ( .A1(a_6_), .A2(b_4_), .ZN(n3371) );
  NAND2_X1 U3364 ( .A1(n2063), .A2(n3328), .ZN(n3365) );
  NAND2_X1 U3365 ( .A1(n3372), .A2(n3373), .ZN(n3328) );
  NAND3_X1 U3366 ( .A1(b_5_), .A2(n3374), .A3(a_6_), .ZN(n3373) );
  OR2_X1 U3367 ( .A1(n3260), .A2(n3262), .ZN(n3374) );
  NAND2_X1 U3368 ( .A1(n3260), .A2(n3262), .ZN(n3372) );
  NAND2_X1 U3369 ( .A1(n3375), .A2(n3376), .ZN(n3262) );
  NAND3_X1 U3370 ( .A1(a_7_), .A2(n3377), .A3(b_5_), .ZN(n3376) );
  OR2_X1 U3371 ( .A1(n3268), .A2(n3269), .ZN(n3377) );
  NAND2_X1 U3372 ( .A1(n3268), .A2(n3269), .ZN(n3375) );
  NAND2_X1 U3373 ( .A1(n3378), .A2(n3379), .ZN(n3269) );
  NAND3_X1 U3374 ( .A1(b_5_), .A2(n3380), .A3(a_8_), .ZN(n3379) );
  OR2_X1 U3375 ( .A1(n3323), .A2(n3325), .ZN(n3380) );
  NAND2_X1 U3376 ( .A1(n3323), .A2(n3325), .ZN(n3378) );
  NAND2_X1 U3377 ( .A1(n3320), .A2(n3381), .ZN(n3325) );
  NAND2_X1 U3378 ( .A1(n3319), .A2(n3321), .ZN(n3381) );
  NAND2_X1 U3379 ( .A1(n3382), .A2(n3383), .ZN(n3321) );
  NAND2_X1 U3380 ( .A1(b_5_), .A2(a_9_), .ZN(n3383) );
  INV_X1 U3381 ( .A(n3384), .ZN(n3382) );
  XNOR2_X1 U3382 ( .A(n3385), .B(n3386), .ZN(n3319) );
  XNOR2_X1 U3383 ( .A(n3387), .B(n3388), .ZN(n3386) );
  NAND2_X1 U3384 ( .A1(a_9_), .A2(n3384), .ZN(n3320) );
  NAND2_X1 U3385 ( .A1(n3389), .A2(n3390), .ZN(n3384) );
  NAND2_X1 U3386 ( .A1(n3284), .A2(n3391), .ZN(n3390) );
  OR2_X1 U3387 ( .A1(n3281), .A2(n3283), .ZN(n3391) );
  NOR2_X1 U3388 ( .A1(n2068), .A2(n2550), .ZN(n3284) );
  NAND2_X1 U3389 ( .A1(n3281), .A2(n3283), .ZN(n3389) );
  NAND2_X1 U3390 ( .A1(n3392), .A2(n3393), .ZN(n3283) );
  NAND2_X1 U3391 ( .A1(n3292), .A2(n3394), .ZN(n3393) );
  NAND2_X1 U3392 ( .A1(n3290), .A2(n3291), .ZN(n3394) );
  NOR2_X1 U3393 ( .A1(n2068), .A2(n1981), .ZN(n3292) );
  OR2_X1 U3394 ( .A1(n3290), .A2(n3291), .ZN(n3392) );
  AND2_X1 U3395 ( .A1(n3395), .A2(n3396), .ZN(n3291) );
  NAND3_X1 U3396 ( .A1(a_12_), .A2(n3397), .A3(b_5_), .ZN(n3396) );
  NAND2_X1 U3397 ( .A1(n3300), .A2(n3298), .ZN(n3397) );
  OR2_X1 U3398 ( .A1(n3298), .A2(n3300), .ZN(n3395) );
  AND2_X1 U3399 ( .A1(n3398), .A2(n3399), .ZN(n3300) );
  NAND2_X1 U3400 ( .A1(n3315), .A2(n3400), .ZN(n3399) );
  OR2_X1 U3401 ( .A1(n3316), .A2(n3317), .ZN(n3400) );
  NOR2_X1 U3402 ( .A1(n2068), .A2(n1952), .ZN(n3315) );
  NAND2_X1 U3403 ( .A1(n3317), .A2(n3316), .ZN(n3398) );
  NAND2_X1 U3404 ( .A1(n3401), .A2(n3402), .ZN(n3316) );
  NAND2_X1 U3405 ( .A1(b_3_), .A2(n3403), .ZN(n3402) );
  NAND2_X1 U3406 ( .A1(n1929), .A2(n3404), .ZN(n3403) );
  NAND2_X1 U3407 ( .A1(a_15_), .A2(n3313), .ZN(n3404) );
  NAND2_X1 U3408 ( .A1(b_4_), .A2(n3405), .ZN(n3401) );
  NAND2_X1 U3409 ( .A1(n1932), .A2(n3406), .ZN(n3405) );
  NAND2_X1 U3410 ( .A1(a_14_), .A2(n2102), .ZN(n3406) );
  AND3_X1 U3411 ( .A1(b_5_), .A2(n2173), .A3(b_4_), .ZN(n3317) );
  XNOR2_X1 U3412 ( .A(n3407), .B(n3408), .ZN(n3298) );
  XOR2_X1 U3413 ( .A(n3409), .B(n3410), .Z(n3407) );
  XNOR2_X1 U3414 ( .A(n3411), .B(n3412), .ZN(n3290) );
  XNOR2_X1 U3415 ( .A(n3413), .B(n3414), .ZN(n3411) );
  NAND2_X1 U3416 ( .A1(b_4_), .A2(a_12_), .ZN(n3413) );
  XNOR2_X1 U3417 ( .A(n3415), .B(n3416), .ZN(n3281) );
  NAND2_X1 U3418 ( .A1(n3417), .A2(n3418), .ZN(n3415) );
  XNOR2_X1 U3419 ( .A(n3419), .B(n3420), .ZN(n3323) );
  NAND2_X1 U3420 ( .A1(n3421), .A2(n3422), .ZN(n3419) );
  XOR2_X1 U3421 ( .A(n3423), .B(n3424), .Z(n3268) );
  XOR2_X1 U3422 ( .A(n3425), .B(n3426), .Z(n3423) );
  NOR2_X1 U3423 ( .A1(n3313), .A2(n2176), .ZN(n3426) );
  XOR2_X1 U3424 ( .A(n3427), .B(n3428), .Z(n3260) );
  XNOR2_X1 U3425 ( .A(n3429), .B(n3430), .ZN(n3428) );
  NAND2_X1 U3426 ( .A1(b_4_), .A2(a_7_), .ZN(n3430) );
  NOR2_X1 U3427 ( .A1(n2068), .A2(n2066), .ZN(n2063) );
  INV_X1 U3428 ( .A(b_5_), .ZN(n2068) );
  XNOR2_X1 U3429 ( .A(n3431), .B(n3432), .ZN(n3251) );
  XOR2_X1 U3430 ( .A(n3433), .B(n3434), .Z(n3431) );
  NOR2_X1 U3431 ( .A1(n2066), .A2(n3313), .ZN(n3434) );
  XOR2_X1 U3432 ( .A(n3435), .B(n3436), .Z(n3330) );
  XNOR2_X1 U3433 ( .A(n2080), .B(n3437), .ZN(n3436) );
  XOR2_X1 U3434 ( .A(n3438), .B(n3439), .Z(n3334) );
  XNOR2_X1 U3435 ( .A(n3440), .B(n3441), .ZN(n3438) );
  NAND2_X1 U3436 ( .A1(a_3_), .A2(b_4_), .ZN(n3440) );
  XOR2_X1 U3437 ( .A(n3442), .B(n3443), .Z(n3337) );
  XOR2_X1 U3438 ( .A(n3444), .B(n3445), .Z(n3443) );
  NAND2_X1 U3439 ( .A1(a_2_), .A2(b_4_), .ZN(n3445) );
  XOR2_X1 U3440 ( .A(n3446), .B(n3447), .Z(n3342) );
  XOR2_X1 U3441 ( .A(n3448), .B(n3449), .Z(n3446) );
  XOR2_X1 U3442 ( .A(n3450), .B(n3451), .Z(n3234) );
  XOR2_X1 U3443 ( .A(n3452), .B(n3453), .Z(n3450) );
  NOR2_X1 U3444 ( .A1(n3313), .A2(n2371), .ZN(n3453) );
  NAND2_X1 U3445 ( .A1(n3454), .A2(n3455), .ZN(n1917) );
  NAND2_X1 U3446 ( .A1(n3348), .A2(n3347), .ZN(n3455) );
  XNOR2_X1 U3447 ( .A(n3456), .B(n3457), .ZN(n3454) );
  NAND3_X1 U3448 ( .A1(n3458), .A2(n3347), .A3(n3348), .ZN(n1916) );
  XOR2_X1 U3449 ( .A(n3459), .B(n3460), .Z(n3348) );
  XOR2_X1 U3450 ( .A(n3461), .B(n3462), .Z(n3459) );
  NOR2_X1 U3451 ( .A1(n2102), .A2(n2371), .ZN(n3462) );
  NAND2_X1 U3452 ( .A1(n3463), .A2(n3464), .ZN(n3347) );
  NAND3_X1 U3453 ( .A1(b_4_), .A2(n3465), .A3(a_0_), .ZN(n3464) );
  OR2_X1 U3454 ( .A1(n3452), .A2(n3451), .ZN(n3465) );
  NAND2_X1 U3455 ( .A1(n3451), .A2(n3452), .ZN(n3463) );
  NAND2_X1 U3456 ( .A1(n3466), .A2(n3467), .ZN(n3452) );
  NAND2_X1 U3457 ( .A1(n3449), .A2(n3468), .ZN(n3467) );
  OR2_X1 U3458 ( .A1(n3448), .A2(n3447), .ZN(n3468) );
  NOR2_X1 U3459 ( .A1(n2360), .A2(n3313), .ZN(n3449) );
  NAND2_X1 U3460 ( .A1(n3447), .A2(n3448), .ZN(n3466) );
  NAND2_X1 U3461 ( .A1(n3469), .A2(n3470), .ZN(n3448) );
  NAND3_X1 U3462 ( .A1(b_4_), .A2(n3471), .A3(a_2_), .ZN(n3470) );
  OR2_X1 U3463 ( .A1(n3442), .A2(n3444), .ZN(n3471) );
  NAND2_X1 U3464 ( .A1(n3442), .A2(n3444), .ZN(n3469) );
  NAND2_X1 U3465 ( .A1(n3472), .A2(n3473), .ZN(n3444) );
  NAND3_X1 U3466 ( .A1(b_4_), .A2(n3474), .A3(a_3_), .ZN(n3473) );
  OR2_X1 U3467 ( .A1(n3441), .A2(n3439), .ZN(n3474) );
  NAND2_X1 U3468 ( .A1(n3439), .A2(n3441), .ZN(n3472) );
  NAND2_X1 U3469 ( .A1(n3475), .A2(n3476), .ZN(n3441) );
  NAND2_X1 U3470 ( .A1(n3435), .A2(n3477), .ZN(n3476) );
  OR2_X1 U3471 ( .A1(n3437), .A2(n2080), .ZN(n3477) );
  XNOR2_X1 U3472 ( .A(n3478), .B(n3479), .ZN(n3435) );
  NAND2_X1 U3473 ( .A1(n3480), .A2(n3481), .ZN(n3478) );
  NAND2_X1 U3474 ( .A1(n2080), .A2(n3437), .ZN(n3475) );
  NAND2_X1 U3475 ( .A1(n3482), .A2(n3483), .ZN(n3437) );
  NAND3_X1 U3476 ( .A1(a_5_), .A2(n3484), .A3(b_4_), .ZN(n3483) );
  OR2_X1 U3477 ( .A1(n3433), .A2(n3432), .ZN(n3484) );
  NAND2_X1 U3478 ( .A1(n3432), .A2(n3433), .ZN(n3482) );
  NAND2_X1 U3479 ( .A1(n3485), .A2(n3486), .ZN(n3433) );
  NAND3_X1 U3480 ( .A1(b_4_), .A2(n3487), .A3(a_6_), .ZN(n3486) );
  OR2_X1 U3481 ( .A1(n3370), .A2(n3368), .ZN(n3487) );
  NAND2_X1 U3482 ( .A1(n3368), .A2(n3370), .ZN(n3485) );
  NAND2_X1 U3483 ( .A1(n3488), .A2(n3489), .ZN(n3370) );
  NAND3_X1 U3484 ( .A1(a_7_), .A2(n3490), .A3(b_4_), .ZN(n3489) );
  NAND2_X1 U3485 ( .A1(n3429), .A2(n3427), .ZN(n3490) );
  OR2_X1 U3486 ( .A1(n3427), .A2(n3429), .ZN(n3488) );
  AND2_X1 U3487 ( .A1(n3491), .A2(n3492), .ZN(n3429) );
  NAND3_X1 U3488 ( .A1(b_4_), .A2(n3493), .A3(a_8_), .ZN(n3492) );
  OR2_X1 U3489 ( .A1(n3425), .A2(n3424), .ZN(n3493) );
  NAND2_X1 U3490 ( .A1(n3424), .A2(n3425), .ZN(n3491) );
  NAND2_X1 U3491 ( .A1(n3421), .A2(n3494), .ZN(n3425) );
  NAND2_X1 U3492 ( .A1(n3420), .A2(n3422), .ZN(n3494) );
  NAND2_X1 U3493 ( .A1(n3495), .A2(n3496), .ZN(n3422) );
  NAND2_X1 U3494 ( .A1(b_4_), .A2(a_9_), .ZN(n3496) );
  INV_X1 U3495 ( .A(n3497), .ZN(n3495) );
  XNOR2_X1 U3496 ( .A(n3498), .B(n3499), .ZN(n3420) );
  NAND2_X1 U3497 ( .A1(n3500), .A2(n3501), .ZN(n3498) );
  NAND2_X1 U3498 ( .A1(a_9_), .A2(n3497), .ZN(n3421) );
  NAND2_X1 U3499 ( .A1(n3502), .A2(n3503), .ZN(n3497) );
  NAND2_X1 U3500 ( .A1(n3388), .A2(n3504), .ZN(n3503) );
  OR2_X1 U3501 ( .A1(n3387), .A2(n3385), .ZN(n3504) );
  NOR2_X1 U3502 ( .A1(n3313), .A2(n2550), .ZN(n3388) );
  NAND2_X1 U3503 ( .A1(n3385), .A2(n3387), .ZN(n3502) );
  NAND2_X1 U3504 ( .A1(n3417), .A2(n3505), .ZN(n3387) );
  NAND2_X1 U3505 ( .A1(n3416), .A2(n3418), .ZN(n3505) );
  NAND2_X1 U3506 ( .A1(n3506), .A2(n3507), .ZN(n3418) );
  NAND2_X1 U3507 ( .A1(b_4_), .A2(a_11_), .ZN(n3507) );
  INV_X1 U3508 ( .A(n3508), .ZN(n3506) );
  XNOR2_X1 U3509 ( .A(n3509), .B(n3510), .ZN(n3416) );
  XNOR2_X1 U3510 ( .A(n3511), .B(n3512), .ZN(n3509) );
  NAND2_X1 U3511 ( .A1(a_11_), .A2(n3508), .ZN(n3417) );
  NAND2_X1 U3512 ( .A1(n3513), .A2(n3514), .ZN(n3508) );
  NAND3_X1 U3513 ( .A1(a_12_), .A2(n3515), .A3(b_4_), .ZN(n3514) );
  OR2_X1 U3514 ( .A1(n3414), .A2(n3412), .ZN(n3515) );
  NAND2_X1 U3515 ( .A1(n3412), .A2(n3414), .ZN(n3513) );
  NAND2_X1 U3516 ( .A1(n3516), .A2(n3517), .ZN(n3414) );
  NAND2_X1 U3517 ( .A1(n3408), .A2(n3518), .ZN(n3517) );
  OR2_X1 U3518 ( .A1(n3409), .A2(n3410), .ZN(n3518) );
  NOR2_X1 U3519 ( .A1(n3313), .A2(n1952), .ZN(n3408) );
  NAND2_X1 U3520 ( .A1(n3410), .A2(n3409), .ZN(n3516) );
  NAND2_X1 U3521 ( .A1(n3519), .A2(n3520), .ZN(n3409) );
  NAND2_X1 U3522 ( .A1(b_2_), .A2(n3521), .ZN(n3520) );
  NAND2_X1 U3523 ( .A1(n1929), .A2(n3522), .ZN(n3521) );
  NAND2_X1 U3524 ( .A1(a_15_), .A2(n2102), .ZN(n3522) );
  NAND2_X1 U3525 ( .A1(b_3_), .A2(n3523), .ZN(n3519) );
  NAND2_X1 U3526 ( .A1(n1932), .A2(n3524), .ZN(n3523) );
  NAND2_X1 U3527 ( .A1(a_14_), .A2(n2177), .ZN(n3524) );
  AND3_X1 U3528 ( .A1(b_4_), .A2(n2173), .A3(b_3_), .ZN(n3410) );
  XOR2_X1 U3529 ( .A(n3525), .B(n3526), .Z(n3412) );
  NOR2_X1 U3530 ( .A1(n1952), .A2(n2102), .ZN(n3526) );
  XOR2_X1 U3531 ( .A(n3527), .B(n3528), .Z(n3525) );
  XNOR2_X1 U3532 ( .A(n3529), .B(n3530), .ZN(n3385) );
  NAND2_X1 U3533 ( .A1(n3531), .A2(n3532), .ZN(n3529) );
  XNOR2_X1 U3534 ( .A(n3533), .B(n3534), .ZN(n3424) );
  NAND2_X1 U3535 ( .A1(n3535), .A2(n3536), .ZN(n3533) );
  XNOR2_X1 U3536 ( .A(n3537), .B(n3538), .ZN(n3427) );
  XOR2_X1 U3537 ( .A(n3539), .B(n3540), .Z(n3537) );
  NOR2_X1 U3538 ( .A1(n2176), .A2(n2102), .ZN(n3540) );
  XNOR2_X1 U3539 ( .A(n3541), .B(n3542), .ZN(n3368) );
  NAND2_X1 U3540 ( .A1(n3543), .A2(n3544), .ZN(n3541) );
  XOR2_X1 U3541 ( .A(n3545), .B(n3546), .Z(n3432) );
  XOR2_X1 U3542 ( .A(n3547), .B(n3548), .Z(n3545) );
  NOR2_X1 U3543 ( .A1(n2102), .A2(n2056), .ZN(n3548) );
  NOR2_X1 U3544 ( .A1(n3313), .A2(n2347), .ZN(n2080) );
  INV_X1 U3545 ( .A(b_4_), .ZN(n3313) );
  XNOR2_X1 U3546 ( .A(n3549), .B(n3550), .ZN(n3439) );
  XNOR2_X1 U3547 ( .A(n3551), .B(n3552), .ZN(n3549) );
  NOR2_X1 U3548 ( .A1(n2347), .A2(n2102), .ZN(n3552) );
  XOR2_X1 U3549 ( .A(n3553), .B(n3554), .Z(n3442) );
  XNOR2_X1 U3550 ( .A(n3555), .B(n2146), .ZN(n3553) );
  INV_X1 U3551 ( .A(n2097), .ZN(n2146) );
  XOR2_X1 U3552 ( .A(n3556), .B(n3557), .Z(n3447) );
  XOR2_X1 U3553 ( .A(n3558), .B(n3559), .Z(n3556) );
  NOR2_X1 U3554 ( .A1(n2102), .A2(n2178), .ZN(n3559) );
  XOR2_X1 U3555 ( .A(n3560), .B(n3561), .Z(n3451) );
  XOR2_X1 U3556 ( .A(n3562), .B(n3563), .Z(n3560) );
  XOR2_X1 U3557 ( .A(n3456), .B(n3457), .Z(n3458) );
  NAND2_X1 U3558 ( .A1(n3564), .A2(n3565), .ZN(n1941) );
  NAND2_X1 U3559 ( .A1(n3457), .A2(n3456), .ZN(n3565) );
  XNOR2_X1 U3560 ( .A(n2221), .B(n2220), .ZN(n3564) );
  NAND3_X1 U3561 ( .A1(n3566), .A2(n3456), .A3(n3457), .ZN(n1940) );
  XNOR2_X1 U3562 ( .A(n3567), .B(n3568), .ZN(n3457) );
  NAND2_X1 U3563 ( .A1(n3569), .A2(n3570), .ZN(n3567) );
  NAND2_X1 U3564 ( .A1(n3571), .A2(n3572), .ZN(n3456) );
  NAND3_X1 U3565 ( .A1(b_3_), .A2(n3573), .A3(a_0_), .ZN(n3572) );
  OR2_X1 U3566 ( .A1(n3460), .A2(n3461), .ZN(n3573) );
  NAND2_X1 U3567 ( .A1(n3460), .A2(n3461), .ZN(n3571) );
  NAND2_X1 U3568 ( .A1(n3574), .A2(n3575), .ZN(n3461) );
  NAND2_X1 U3569 ( .A1(n3563), .A2(n3576), .ZN(n3575) );
  OR2_X1 U3570 ( .A1(n3561), .A2(n3562), .ZN(n3576) );
  NOR2_X1 U3571 ( .A1(n2360), .A2(n2102), .ZN(n3563) );
  NAND2_X1 U3572 ( .A1(n3561), .A2(n3562), .ZN(n3574) );
  NAND2_X1 U3573 ( .A1(n3577), .A2(n3578), .ZN(n3562) );
  NAND3_X1 U3574 ( .A1(b_3_), .A2(n3579), .A3(a_2_), .ZN(n3578) );
  OR2_X1 U3575 ( .A1(n3557), .A2(n3558), .ZN(n3579) );
  NAND2_X1 U3576 ( .A1(n3557), .A2(n3558), .ZN(n3577) );
  NAND2_X1 U3577 ( .A1(n3580), .A2(n3581), .ZN(n3558) );
  NAND2_X1 U3578 ( .A1(n3554), .A2(n3582), .ZN(n3581) );
  OR2_X1 U3579 ( .A1(n3555), .A2(n2097), .ZN(n3582) );
  XNOR2_X1 U3580 ( .A(n3583), .B(n3584), .ZN(n3554) );
  NAND2_X1 U3581 ( .A1(n3585), .A2(n3586), .ZN(n3583) );
  NAND2_X1 U3582 ( .A1(n2097), .A2(n3555), .ZN(n3580) );
  NAND2_X1 U3583 ( .A1(n3587), .A2(n3588), .ZN(n3555) );
  NAND3_X1 U3584 ( .A1(a_4_), .A2(n3589), .A3(b_3_), .ZN(n3588) );
  NAND2_X1 U3585 ( .A1(n3550), .A2(n3551), .ZN(n3589) );
  OR2_X1 U3586 ( .A1(n3550), .A2(n3551), .ZN(n3587) );
  AND2_X1 U3587 ( .A1(n3480), .A2(n3590), .ZN(n3551) );
  NAND2_X1 U3588 ( .A1(n3479), .A2(n3481), .ZN(n3590) );
  NAND2_X1 U3589 ( .A1(n3591), .A2(n3592), .ZN(n3481) );
  NAND2_X1 U3590 ( .A1(b_3_), .A2(a_5_), .ZN(n3592) );
  INV_X1 U3591 ( .A(n3593), .ZN(n3591) );
  XNOR2_X1 U3592 ( .A(n3594), .B(n3595), .ZN(n3479) );
  NAND2_X1 U3593 ( .A1(n3596), .A2(n3597), .ZN(n3594) );
  NAND2_X1 U3594 ( .A1(a_5_), .A2(n3593), .ZN(n3480) );
  NAND2_X1 U3595 ( .A1(n3598), .A2(n3599), .ZN(n3593) );
  NAND3_X1 U3596 ( .A1(b_3_), .A2(n3600), .A3(a_6_), .ZN(n3599) );
  OR2_X1 U3597 ( .A1(n3546), .A2(n3547), .ZN(n3600) );
  NAND2_X1 U3598 ( .A1(n3546), .A2(n3547), .ZN(n3598) );
  NAND2_X1 U3599 ( .A1(n3543), .A2(n3601), .ZN(n3547) );
  NAND2_X1 U3600 ( .A1(n3542), .A2(n3544), .ZN(n3601) );
  NAND2_X1 U3601 ( .A1(n3602), .A2(n3603), .ZN(n3544) );
  NAND2_X1 U3602 ( .A1(b_3_), .A2(a_7_), .ZN(n3603) );
  INV_X1 U3603 ( .A(n3604), .ZN(n3602) );
  XNOR2_X1 U3604 ( .A(n3605), .B(n3606), .ZN(n3542) );
  NAND2_X1 U3605 ( .A1(n3607), .A2(n3608), .ZN(n3605) );
  NAND2_X1 U3606 ( .A1(a_7_), .A2(n3604), .ZN(n3543) );
  NAND2_X1 U3607 ( .A1(n3609), .A2(n3610), .ZN(n3604) );
  NAND3_X1 U3608 ( .A1(a_8_), .A2(n3611), .A3(b_3_), .ZN(n3610) );
  OR2_X1 U3609 ( .A1(n3538), .A2(n3539), .ZN(n3611) );
  NAND2_X1 U3610 ( .A1(n3538), .A2(n3539), .ZN(n3609) );
  NAND2_X1 U3611 ( .A1(n3535), .A2(n3612), .ZN(n3539) );
  NAND2_X1 U3612 ( .A1(n3534), .A2(n3536), .ZN(n3612) );
  NAND2_X1 U3613 ( .A1(n3613), .A2(n3614), .ZN(n3536) );
  NAND2_X1 U3614 ( .A1(b_3_), .A2(a_9_), .ZN(n3614) );
  INV_X1 U3615 ( .A(n3615), .ZN(n3613) );
  XNOR2_X1 U3616 ( .A(n3616), .B(n3617), .ZN(n3534) );
  NAND2_X1 U3617 ( .A1(n3618), .A2(n3619), .ZN(n3616) );
  NAND2_X1 U3618 ( .A1(a_9_), .A2(n3615), .ZN(n3535) );
  NAND2_X1 U3619 ( .A1(n3500), .A2(n3620), .ZN(n3615) );
  NAND2_X1 U3620 ( .A1(n3499), .A2(n3501), .ZN(n3620) );
  NAND2_X1 U3621 ( .A1(n3621), .A2(n3622), .ZN(n3501) );
  NAND2_X1 U3622 ( .A1(b_3_), .A2(a_10_), .ZN(n3622) );
  INV_X1 U3623 ( .A(n3623), .ZN(n3621) );
  XNOR2_X1 U3624 ( .A(n3624), .B(n3625), .ZN(n3499) );
  XNOR2_X1 U3625 ( .A(n3626), .B(n3627), .ZN(n3625) );
  NAND2_X1 U3626 ( .A1(a_10_), .A2(n3623), .ZN(n3500) );
  NAND2_X1 U3627 ( .A1(n3531), .A2(n3628), .ZN(n3623) );
  NAND2_X1 U3628 ( .A1(n3530), .A2(n3532), .ZN(n3628) );
  NAND2_X1 U3629 ( .A1(n3629), .A2(n3630), .ZN(n3532) );
  NAND2_X1 U3630 ( .A1(b_3_), .A2(a_11_), .ZN(n3630) );
  INV_X1 U3631 ( .A(n3631), .ZN(n3629) );
  XNOR2_X1 U3632 ( .A(n3632), .B(n3633), .ZN(n3530) );
  XNOR2_X1 U3633 ( .A(n3634), .B(n3635), .ZN(n3632) );
  NOR2_X1 U3634 ( .A1(n1970), .A2(n2177), .ZN(n3635) );
  NAND2_X1 U3635 ( .A1(a_11_), .A2(n3631), .ZN(n3531) );
  NAND2_X1 U3636 ( .A1(n3636), .A2(n3637), .ZN(n3631) );
  NAND2_X1 U3637 ( .A1(n3511), .A2(n3638), .ZN(n3637) );
  NAND2_X1 U3638 ( .A1(n3512), .A2(n3510), .ZN(n3638) );
  NOR2_X1 U3639 ( .A1(n2102), .A2(n1970), .ZN(n3511) );
  OR2_X1 U3640 ( .A1(n3510), .A2(n3512), .ZN(n3636) );
  AND2_X1 U3641 ( .A1(n3639), .A2(n3640), .ZN(n3512) );
  NAND3_X1 U3642 ( .A1(a_13_), .A2(n3641), .A3(b_3_), .ZN(n3640) );
  OR2_X1 U3643 ( .A1(n3527), .A2(n3528), .ZN(n3641) );
  NAND2_X1 U3644 ( .A1(n3528), .A2(n3527), .ZN(n3639) );
  NAND2_X1 U3645 ( .A1(n3642), .A2(n3643), .ZN(n3527) );
  NAND2_X1 U3646 ( .A1(b_1_), .A2(n3644), .ZN(n3643) );
  NAND2_X1 U3647 ( .A1(n1929), .A2(n3645), .ZN(n3644) );
  NAND2_X1 U3648 ( .A1(a_15_), .A2(n2177), .ZN(n3645) );
  NAND2_X1 U3649 ( .A1(b_2_), .A2(n3646), .ZN(n3642) );
  NAND2_X1 U3650 ( .A1(n1932), .A2(n3647), .ZN(n3646) );
  NAND2_X1 U3651 ( .A1(a_14_), .A2(n2131), .ZN(n3647) );
  AND3_X1 U3652 ( .A1(b_3_), .A2(n2173), .A3(b_2_), .ZN(n3528) );
  XNOR2_X1 U3653 ( .A(n3648), .B(n3649), .ZN(n3510) );
  NOR2_X1 U3654 ( .A1(n1952), .A2(n2177), .ZN(n3649) );
  XOR2_X1 U3655 ( .A(n3650), .B(n3651), .Z(n3648) );
  XOR2_X1 U3656 ( .A(n3652), .B(n3653), .Z(n3538) );
  XOR2_X1 U3657 ( .A(n3654), .B(n3655), .Z(n3652) );
  XOR2_X1 U3658 ( .A(n3656), .B(n3657), .Z(n3546) );
  XOR2_X1 U3659 ( .A(n3658), .B(n3659), .Z(n3656) );
  XNOR2_X1 U3660 ( .A(n3660), .B(n3661), .ZN(n3550) );
  XOR2_X1 U3661 ( .A(n3662), .B(n3663), .Z(n3660) );
  NOR2_X1 U3662 ( .A1(n2100), .A2(n2102), .ZN(n2097) );
  INV_X1 U3663 ( .A(b_3_), .ZN(n2102) );
  XOR2_X1 U3664 ( .A(n3664), .B(n3665), .Z(n3557) );
  XOR2_X1 U3665 ( .A(n3666), .B(n3667), .Z(n3664) );
  XOR2_X1 U3666 ( .A(n3668), .B(n3669), .Z(n3561) );
  XOR2_X1 U3667 ( .A(n2114), .B(n3670), .Z(n3668) );
  XOR2_X1 U3668 ( .A(n3671), .B(n3672), .Z(n3460) );
  XOR2_X1 U3669 ( .A(n3673), .B(n3674), .Z(n3671) );
  NOR2_X1 U3670 ( .A1(n2177), .A2(n2360), .ZN(n3674) );
  XOR2_X1 U3671 ( .A(n2221), .B(n2220), .Z(n3566) );
  INV_X1 U3672 ( .A(n2090), .ZN(n2216) );
  NAND4_X1 U3673 ( .A1(n2143), .A2(n2222), .A3(n2220), .A4(n2221), .ZN(n2090)
         );
  NAND2_X1 U3674 ( .A1(n3569), .A2(n3675), .ZN(n2221) );
  NAND2_X1 U3675 ( .A1(n3568), .A2(n3570), .ZN(n3675) );
  NAND2_X1 U3676 ( .A1(n3676), .A2(n3677), .ZN(n3570) );
  NAND2_X1 U3677 ( .A1(a_0_), .A2(b_2_), .ZN(n3677) );
  INV_X1 U3678 ( .A(n3678), .ZN(n3676) );
  XOR2_X1 U3679 ( .A(n3679), .B(n3680), .Z(n3568) );
  XOR2_X1 U3680 ( .A(n3681), .B(n2127), .Z(n3679) );
  NAND2_X1 U3681 ( .A1(a_0_), .A2(n3678), .ZN(n3569) );
  NAND2_X1 U3682 ( .A1(n3682), .A2(n3683), .ZN(n3678) );
  NAND3_X1 U3683 ( .A1(b_2_), .A2(n3684), .A3(a_1_), .ZN(n3683) );
  OR2_X1 U3684 ( .A1(n3673), .A2(n3672), .ZN(n3684) );
  NAND2_X1 U3685 ( .A1(n3672), .A2(n3673), .ZN(n3682) );
  NAND2_X1 U3686 ( .A1(n3685), .A2(n3686), .ZN(n3673) );
  NAND2_X1 U3687 ( .A1(n3669), .A2(n3687), .ZN(n3686) );
  NAND2_X1 U3688 ( .A1(n3670), .A2(n2114), .ZN(n3687) );
  XOR2_X1 U3689 ( .A(n3688), .B(n3689), .Z(n3669) );
  XOR2_X1 U3690 ( .A(n3690), .B(n3691), .Z(n3688) );
  OR2_X1 U3691 ( .A1(n2114), .A2(n3670), .ZN(n3685) );
  AND2_X1 U3692 ( .A1(n3692), .A2(n3693), .ZN(n3670) );
  NAND2_X1 U3693 ( .A1(n3667), .A2(n3694), .ZN(n3693) );
  OR2_X1 U3694 ( .A1(n3666), .A2(n3665), .ZN(n3694) );
  NOR2_X1 U3695 ( .A1(n2100), .A2(n2177), .ZN(n3667) );
  NAND2_X1 U3696 ( .A1(n3665), .A2(n3666), .ZN(n3692) );
  NAND2_X1 U3697 ( .A1(n3585), .A2(n3695), .ZN(n3666) );
  NAND2_X1 U3698 ( .A1(n3584), .A2(n3586), .ZN(n3695) );
  NAND2_X1 U3699 ( .A1(n3696), .A2(n3697), .ZN(n3586) );
  NAND2_X1 U3700 ( .A1(b_2_), .A2(a_4_), .ZN(n3697) );
  INV_X1 U3701 ( .A(n3698), .ZN(n3696) );
  XOR2_X1 U3702 ( .A(n3699), .B(n3700), .Z(n3584) );
  XOR2_X1 U3703 ( .A(n3701), .B(n3702), .Z(n3699) );
  NAND2_X1 U3704 ( .A1(a_4_), .A2(n3698), .ZN(n3585) );
  NAND2_X1 U3705 ( .A1(n3703), .A2(n3704), .ZN(n3698) );
  NAND2_X1 U3706 ( .A1(n3663), .A2(n3705), .ZN(n3704) );
  OR2_X1 U3707 ( .A1(n3662), .A2(n3661), .ZN(n3705) );
  NOR2_X1 U3708 ( .A1(n2177), .A2(n2066), .ZN(n3663) );
  NAND2_X1 U3709 ( .A1(n3661), .A2(n3662), .ZN(n3703) );
  NAND2_X1 U3710 ( .A1(n3596), .A2(n3706), .ZN(n3662) );
  NAND2_X1 U3711 ( .A1(n3595), .A2(n3597), .ZN(n3706) );
  NAND2_X1 U3712 ( .A1(n3707), .A2(n3708), .ZN(n3597) );
  NAND2_X1 U3713 ( .A1(a_6_), .A2(b_2_), .ZN(n3708) );
  INV_X1 U3714 ( .A(n3709), .ZN(n3707) );
  XOR2_X1 U3715 ( .A(n3710), .B(n3711), .Z(n3595) );
  XOR2_X1 U3716 ( .A(n3712), .B(n3713), .Z(n3710) );
  NAND2_X1 U3717 ( .A1(a_6_), .A2(n3709), .ZN(n3596) );
  NAND2_X1 U3718 ( .A1(n3714), .A2(n3715), .ZN(n3709) );
  NAND2_X1 U3719 ( .A1(n3659), .A2(n3716), .ZN(n3715) );
  OR2_X1 U3720 ( .A1(n3658), .A2(n3657), .ZN(n3716) );
  NOR2_X1 U3721 ( .A1(n2177), .A2(n2038), .ZN(n3659) );
  NAND2_X1 U3722 ( .A1(n3657), .A2(n3658), .ZN(n3714) );
  NAND2_X1 U3723 ( .A1(n3607), .A2(n3717), .ZN(n3658) );
  NAND2_X1 U3724 ( .A1(n3606), .A2(n3608), .ZN(n3717) );
  NAND2_X1 U3725 ( .A1(n3718), .A2(n3719), .ZN(n3608) );
  NAND2_X1 U3726 ( .A1(b_2_), .A2(a_8_), .ZN(n3719) );
  INV_X1 U3727 ( .A(n3720), .ZN(n3718) );
  XNOR2_X1 U3728 ( .A(n3721), .B(n3722), .ZN(n3606) );
  XNOR2_X1 U3729 ( .A(n3723), .B(n3724), .ZN(n3722) );
  NAND2_X1 U3730 ( .A1(a_8_), .A2(n3720), .ZN(n3607) );
  NAND2_X1 U3731 ( .A1(n3725), .A2(n3726), .ZN(n3720) );
  NAND2_X1 U3732 ( .A1(n3655), .A2(n3727), .ZN(n3726) );
  OR2_X1 U3733 ( .A1(n3654), .A2(n3653), .ZN(n3727) );
  NOR2_X1 U3734 ( .A1(n2177), .A2(n2008), .ZN(n3655) );
  NAND2_X1 U3735 ( .A1(n3653), .A2(n3654), .ZN(n3725) );
  NAND2_X1 U3736 ( .A1(n3618), .A2(n3728), .ZN(n3654) );
  NAND2_X1 U3737 ( .A1(n3617), .A2(n3619), .ZN(n3728) );
  NAND2_X1 U3738 ( .A1(n3729), .A2(n3730), .ZN(n3619) );
  NAND2_X1 U3739 ( .A1(b_2_), .A2(a_10_), .ZN(n3730) );
  INV_X1 U3740 ( .A(n3731), .ZN(n3729) );
  XNOR2_X1 U3741 ( .A(n3732), .B(n3733), .ZN(n3617) );
  XNOR2_X1 U3742 ( .A(n3734), .B(n3735), .ZN(n3733) );
  NAND2_X1 U3743 ( .A1(a_10_), .A2(n3731), .ZN(n3618) );
  NAND2_X1 U3744 ( .A1(n3736), .A2(n3737), .ZN(n3731) );
  NAND2_X1 U3745 ( .A1(n3627), .A2(n3738), .ZN(n3737) );
  OR2_X1 U3746 ( .A1(n3626), .A2(n3624), .ZN(n3738) );
  NOR2_X1 U3747 ( .A1(n2177), .A2(n1981), .ZN(n3627) );
  INV_X1 U3748 ( .A(b_2_), .ZN(n2177) );
  NAND2_X1 U3749 ( .A1(n3624), .A2(n3626), .ZN(n3736) );
  NAND2_X1 U3750 ( .A1(n3739), .A2(n3740), .ZN(n3626) );
  NAND3_X1 U3751 ( .A1(a_12_), .A2(n3741), .A3(b_2_), .ZN(n3740) );
  NAND2_X1 U3752 ( .A1(n3633), .A2(n3634), .ZN(n3741) );
  OR2_X1 U3753 ( .A1(n3633), .A2(n3634), .ZN(n3739) );
  AND2_X1 U3754 ( .A1(n3742), .A2(n3743), .ZN(n3634) );
  NAND3_X1 U3755 ( .A1(a_13_), .A2(n3744), .A3(b_2_), .ZN(n3743) );
  OR2_X1 U3756 ( .A1(n3650), .A2(n3651), .ZN(n3744) );
  NAND2_X1 U3757 ( .A1(n3651), .A2(n3650), .ZN(n3742) );
  NAND2_X1 U3758 ( .A1(n3745), .A2(n3746), .ZN(n3650) );
  NAND2_X1 U3759 ( .A1(b_0_), .A2(n3747), .ZN(n3746) );
  NAND2_X1 U3760 ( .A1(n3748), .A2(n1929), .ZN(n3747) );
  NAND2_X1 U3761 ( .A1(a_15_), .A2(n2172), .ZN(n1929) );
  NAND2_X1 U3762 ( .A1(a_15_), .A2(n2131), .ZN(n3748) );
  NAND2_X1 U3763 ( .A1(b_1_), .A2(n3749), .ZN(n3745) );
  NAND2_X1 U3764 ( .A1(n3750), .A2(n1932), .ZN(n3749) );
  OR2_X1 U3765 ( .A1(n2172), .A2(a_15_), .ZN(n1932) );
  INV_X1 U3766 ( .A(a_14_), .ZN(n2172) );
  NAND2_X1 U3767 ( .A1(a_14_), .A2(n3751), .ZN(n3750) );
  AND3_X1 U3768 ( .A1(b_2_), .A2(n2173), .A3(b_1_), .ZN(n3651) );
  XOR2_X1 U3769 ( .A(n3752), .B(n3753), .Z(n3633) );
  XNOR2_X1 U3770 ( .A(n3754), .B(n3755), .ZN(n3753) );
  NAND2_X1 U3771 ( .A1(b_0_), .A2(a_14_), .ZN(n3752) );
  XOR2_X1 U3772 ( .A(n3756), .B(n3757), .Z(n3624) );
  XOR2_X1 U3773 ( .A(n3758), .B(n3759), .Z(n3756) );
  XOR2_X1 U3774 ( .A(n3760), .B(n3761), .Z(n3653) );
  XOR2_X1 U3775 ( .A(n3762), .B(n3763), .Z(n3760) );
  XOR2_X1 U3776 ( .A(n3764), .B(n3765), .Z(n3657) );
  XOR2_X1 U3777 ( .A(n3766), .B(n3767), .Z(n3764) );
  XOR2_X1 U3778 ( .A(n3768), .B(n3769), .Z(n3661) );
  XOR2_X1 U3779 ( .A(n3770), .B(n3771), .Z(n3768) );
  XOR2_X1 U3780 ( .A(n3772), .B(n3773), .Z(n3665) );
  XOR2_X1 U3781 ( .A(n3774), .B(n3775), .Z(n3772) );
  NAND2_X1 U3782 ( .A1(a_2_), .A2(b_2_), .ZN(n2114) );
  XOR2_X1 U3783 ( .A(n3776), .B(n3777), .Z(n3672) );
  NOR2_X1 U3784 ( .A1(n2131), .A2(n2178), .ZN(n3777) );
  XOR2_X1 U3785 ( .A(n3778), .B(n3779), .Z(n3776) );
  XOR2_X1 U3786 ( .A(n3780), .B(n3781), .Z(n2220) );
  NOR2_X1 U3787 ( .A1(n3751), .A2(n2360), .ZN(n3781) );
  XOR2_X1 U3788 ( .A(n3782), .B(n3783), .Z(n3780) );
  NOR2_X1 U3789 ( .A1(n2371), .A2(n3751), .ZN(n2143) );
  NOR2_X1 U3790 ( .A1(n2222), .A2(n2371), .ZN(n2215) );
  AND2_X1 U3791 ( .A1(n3784), .A2(n3785), .ZN(n2222) );
  NAND3_X1 U3792 ( .A1(b_0_), .A2(n3786), .A3(a_1_), .ZN(n3785) );
  OR2_X1 U3793 ( .A1(n3783), .A2(n3782), .ZN(n3786) );
  NAND2_X1 U3794 ( .A1(n3782), .A2(n3783), .ZN(n3784) );
  NAND2_X1 U3795 ( .A1(n3787), .A2(n3788), .ZN(n3783) );
  NAND2_X1 U3796 ( .A1(n3680), .A2(n3789), .ZN(n3788) );
  OR2_X1 U3797 ( .A1(n3681), .A2(n2127), .ZN(n3789) );
  NOR2_X1 U3798 ( .A1(n2178), .A2(n3751), .ZN(n3680) );
  INV_X1 U3799 ( .A(a_2_), .ZN(n2178) );
  NAND2_X1 U3800 ( .A1(n2127), .A2(n3681), .ZN(n3787) );
  NAND2_X1 U3801 ( .A1(n3790), .A2(n3791), .ZN(n3681) );
  NAND3_X1 U3802 ( .A1(b_1_), .A2(n3792), .A3(a_2_), .ZN(n3791) );
  OR2_X1 U3803 ( .A1(n3779), .A2(n3778), .ZN(n3792) );
  NAND2_X1 U3804 ( .A1(n3778), .A2(n3779), .ZN(n3790) );
  NAND2_X1 U3805 ( .A1(n3793), .A2(n3794), .ZN(n3779) );
  NAND2_X1 U3806 ( .A1(n3689), .A2(n3795), .ZN(n3794) );
  OR2_X1 U3807 ( .A1(n3690), .A2(n3691), .ZN(n3795) );
  NOR2_X1 U3808 ( .A1(n2100), .A2(n2131), .ZN(n3689) );
  NAND2_X1 U3809 ( .A1(n3691), .A2(n3690), .ZN(n3793) );
  NAND2_X1 U3810 ( .A1(n3796), .A2(n3797), .ZN(n3690) );
  NAND2_X1 U3811 ( .A1(n3773), .A2(n3798), .ZN(n3797) );
  OR2_X1 U3812 ( .A1(n3775), .A2(n3774), .ZN(n3798) );
  NOR2_X1 U3813 ( .A1(n2131), .A2(n2347), .ZN(n3773) );
  NAND2_X1 U3814 ( .A1(n3774), .A2(n3775), .ZN(n3796) );
  NAND2_X1 U3815 ( .A1(n3799), .A2(n3800), .ZN(n3775) );
  NAND2_X1 U3816 ( .A1(n3700), .A2(n3801), .ZN(n3800) );
  OR2_X1 U3817 ( .A1(n3701), .A2(n3702), .ZN(n3801) );
  NOR2_X1 U3818 ( .A1(n2131), .A2(n2066), .ZN(n3700) );
  NAND2_X1 U3819 ( .A1(n3702), .A2(n3701), .ZN(n3799) );
  NAND2_X1 U3820 ( .A1(n3802), .A2(n3803), .ZN(n3701) );
  NAND2_X1 U3821 ( .A1(n3769), .A2(n3804), .ZN(n3803) );
  OR2_X1 U3822 ( .A1(n3771), .A2(n3770), .ZN(n3804) );
  NOR2_X1 U3823 ( .A1(n2131), .A2(n2056), .ZN(n3769) );
  NAND2_X1 U3824 ( .A1(n3770), .A2(n3771), .ZN(n3802) );
  NAND2_X1 U3825 ( .A1(n3805), .A2(n3806), .ZN(n3771) );
  NAND2_X1 U3826 ( .A1(n3711), .A2(n3807), .ZN(n3806) );
  OR2_X1 U3827 ( .A1(n3712), .A2(n3713), .ZN(n3807) );
  NOR2_X1 U3828 ( .A1(n2131), .A2(n2038), .ZN(n3711) );
  NAND2_X1 U3829 ( .A1(n3713), .A2(n3712), .ZN(n3805) );
  NAND2_X1 U3830 ( .A1(n3808), .A2(n3809), .ZN(n3712) );
  NAND2_X1 U3831 ( .A1(n3765), .A2(n3810), .ZN(n3809) );
  OR2_X1 U3832 ( .A1(n3767), .A2(n3766), .ZN(n3810) );
  NOR2_X1 U3833 ( .A1(n2131), .A2(n2176), .ZN(n3765) );
  NAND2_X1 U3834 ( .A1(n3766), .A2(n3767), .ZN(n3808) );
  NAND2_X1 U3835 ( .A1(n3811), .A2(n3812), .ZN(n3767) );
  NAND2_X1 U3836 ( .A1(n3721), .A2(n3813), .ZN(n3812) );
  NAND2_X1 U3837 ( .A1(n3723), .A2(n3724), .ZN(n3813) );
  NOR2_X1 U3838 ( .A1(n2131), .A2(n2008), .ZN(n3721) );
  OR2_X1 U3839 ( .A1(n3724), .A2(n3723), .ZN(n3811) );
  AND2_X1 U3840 ( .A1(n3814), .A2(n3815), .ZN(n3723) );
  NAND2_X1 U3841 ( .A1(n3761), .A2(n3816), .ZN(n3815) );
  OR2_X1 U3842 ( .A1(n3763), .A2(n3762), .ZN(n3816) );
  NOR2_X1 U3843 ( .A1(n2131), .A2(n2550), .ZN(n3761) );
  INV_X1 U3844 ( .A(a_10_), .ZN(n2550) );
  NAND2_X1 U3845 ( .A1(n3762), .A2(n3763), .ZN(n3814) );
  NAND2_X1 U3846 ( .A1(n3817), .A2(n3818), .ZN(n3763) );
  NAND2_X1 U3847 ( .A1(n3732), .A2(n3819), .ZN(n3818) );
  NAND2_X1 U3848 ( .A1(n3734), .A2(n3735), .ZN(n3819) );
  NOR2_X1 U3849 ( .A1(n2131), .A2(n1981), .ZN(n3732) );
  OR2_X1 U3850 ( .A1(n3735), .A2(n3734), .ZN(n3817) );
  AND2_X1 U3851 ( .A1(n3820), .A2(n3821), .ZN(n3734) );
  NAND2_X1 U3852 ( .A1(n3757), .A2(n3822), .ZN(n3821) );
  OR2_X1 U3853 ( .A1(n3759), .A2(n3758), .ZN(n3822) );
  NOR2_X1 U3854 ( .A1(n2131), .A2(n1970), .ZN(n3757) );
  INV_X1 U3855 ( .A(a_12_), .ZN(n1970) );
  NAND2_X1 U3856 ( .A1(n3758), .A2(n3759), .ZN(n3820) );
  NAND2_X1 U3857 ( .A1(n3755), .A2(n3823), .ZN(n3759) );
  NAND3_X1 U3858 ( .A1(b_0_), .A2(a_14_), .A3(n3754), .ZN(n3823) );
  NOR2_X1 U3859 ( .A1(n2131), .A2(n1952), .ZN(n3754) );
  NAND3_X1 U3860 ( .A1(b_1_), .A2(n2173), .A3(b_0_), .ZN(n3755) );
  AND2_X1 U3861 ( .A1(a_15_), .A2(a_14_), .ZN(n2173) );
  NOR2_X1 U3862 ( .A1(n3751), .A2(n1952), .ZN(n3758) );
  INV_X1 U3863 ( .A(a_13_), .ZN(n1952) );
  NAND2_X1 U3864 ( .A1(b_0_), .A2(a_12_), .ZN(n3735) );
  NOR2_X1 U3865 ( .A1(n3751), .A2(n1981), .ZN(n3762) );
  INV_X1 U3866 ( .A(a_11_), .ZN(n1981) );
  NAND2_X1 U3867 ( .A1(b_0_), .A2(a_10_), .ZN(n3724) );
  NOR2_X1 U3868 ( .A1(n3751), .A2(n2008), .ZN(n3766) );
  INV_X1 U3869 ( .A(a_9_), .ZN(n2008) );
  NOR2_X1 U3870 ( .A1(n3751), .A2(n2176), .ZN(n3713) );
  INV_X1 U3871 ( .A(a_8_), .ZN(n2176) );
  NOR2_X1 U3872 ( .A1(n3751), .A2(n2038), .ZN(n3770) );
  INV_X1 U3873 ( .A(a_7_), .ZN(n2038) );
  NOR2_X1 U3874 ( .A1(n3751), .A2(n2056), .ZN(n3702) );
  INV_X1 U3875 ( .A(a_6_), .ZN(n2056) );
  NOR2_X1 U3876 ( .A1(n3751), .A2(n2066), .ZN(n3774) );
  INV_X1 U3877 ( .A(a_5_), .ZN(n2066) );
  NOR2_X1 U3878 ( .A1(n3751), .A2(n2347), .ZN(n3691) );
  INV_X1 U3879 ( .A(a_4_), .ZN(n2347) );
  NOR2_X1 U3880 ( .A1(n2100), .A2(n3751), .ZN(n3778) );
  INV_X1 U3881 ( .A(b_0_), .ZN(n3751) );
  INV_X1 U3882 ( .A(a_3_), .ZN(n2100) );
  NOR2_X1 U3883 ( .A1(n2360), .A2(n2131), .ZN(n2127) );
  INV_X1 U3884 ( .A(a_1_), .ZN(n2360) );
  NOR2_X1 U3885 ( .A1(n2371), .A2(n2131), .ZN(n3782) );
  INV_X1 U3886 ( .A(b_1_), .ZN(n2131) );
  INV_X1 U3887 ( .A(a_0_), .ZN(n2371) );
endmodule

