module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n608_, new_n501_, new_n1157_, new_n421_, new_n777_, new_n1048_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n241_, new_n566_, new_n186_, new_n339_, new_n641_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n173_, new_n728_, new_n1071_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n1213_, new_n752_, new_n1045_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n721_, new_n504_, new_n742_, new_n892_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n774_, new_n792_, new_n953_, new_n257_, new_n481_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1212_, new_n1059_, new_n634_, new_n192_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n655_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n694_, new_n461_, new_n297_, new_n565_, new_n1196_, new_n183_, new_n511_, new_n303_, new_n325_, new_n1031_, new_n1216_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n324_, new_n960_, new_n491_, new_n549_, new_n676_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1062_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1198_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n207_, new_n267_, new_n473_, new_n1147_, new_n1229_, new_n187_, new_n969_, new_n334_, new_n331_, new_n835_, new_n378_, new_n621_, new_n244_, new_n172_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n1003_, new_n696_, new_n208_, new_n1039_, new_n528_, new_n952_, new_n179_, new_n1158_, new_n729_, new_n1111_, new_n1218_, new_n559_, new_n1201_, new_n762_, new_n1193_, new_n1187_, new_n1205_, new_n1154_, new_n295_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n1032_, new_n867_, new_n954_, new_n901_, new_n1171_, new_n276_, new_n688_, new_n410_, new_n985_, new_n851_, new_n932_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n724_, new_n1070_, new_n1109_, new_n261_, new_n672_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n604_, new_n1104_, new_n571_, new_n758_, new_n328_, new_n460_, new_n268_, new_n380_, new_n1079_, new_n861_, new_n352_, new_n931_, new_n575_, new_n562_, new_n944_, new_n1064_, new_n1065_, new_n177_, new_n1118_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n993_, new_n1191_, new_n824_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n858_, new_n936_, new_n189_, new_n411_, new_n1016_, new_n673_, new_n1144_, new_n182_, new_n407_, new_n666_, new_n736_, new_n879_, new_n513_, new_n558_, new_n219_, new_n313_, new_n382_, new_n239_, new_n718_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n1040_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n537_, new_n345_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n1122_, new_n1185_, new_n354_, new_n1174_, new_n968_, new_n613_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n591_, new_n837_, new_n801_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n531_, new_n593_, new_n974_, new_n252_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n1052_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1220_, new_n989_, new_n1117_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n196_, new_n818_, new_n881_, new_n640_, new_n684_, new_n754_, new_n653_, new_n377_, new_n905_, new_n375_, new_n962_, new_n760_, new_n627_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n1183_, new_n245_, new_n643_, new_n1194_, new_n1230_, new_n1027_, new_n348_, new_n610_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1165_, new_n175_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n770_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n955_, new_n847_, new_n250_, new_n888_, new_n288_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n827_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n197_, new_n1211_, new_n1207_, new_n1176_, new_n601_, new_n842_, new_n1057_, new_n682_, new_n1075_, new_n812_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n1210_, new_n188_, new_n1060_, new_n240_, new_n413_, new_n442_, new_n677_, new_n642_, new_n211_, new_n462_, new_n603_, new_n564_, new_n761_, new_n840_, new_n735_, new_n898_, new_n799_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n716_, new_n701_, new_n1058_, new_n1162_, new_n212_, new_n902_, new_n364_, new_n832_, new_n201_, new_n414_, new_n1101_, new_n315_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n281_, new_n430_, new_n844_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n829_, new_n988_, new_n478_, new_n1228_, new_n710_, new_n971_, new_n906_, new_n361_, new_n764_, new_n683_, new_n463_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n517_, new_n609_, new_n180_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1051_, new_n899_, new_n1053_, new_n205_, new_n492_, new_n1200_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1219_, new_n920_, new_n1121_, new_n820_, new_n771_, new_n979_, new_n508_, new_n714_, new_n1007_, new_n882_, new_n1145_, new_n929_, new_n986_, new_n314_, new_n1159_, new_n216_, new_n917_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n210_, new_n541_, new_n447_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n341_, new_n996_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n848_, new_n277_, new_n663_, new_n579_, new_n286_, new_n198_, new_n438_, new_n939_, new_n632_, new_n671_, new_n965_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n397_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n948_, new_n1231_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1128_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1161_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n1000_, new_n633_, new_n784_, new_n258_, new_n176_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n747_, new_n749_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n1094_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n578_, new_n918_, new_n940_, new_n810_, new_n808_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1001_, new_n253_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n592_, new_n726_, new_n1123_, new_n231_, new_n583_, new_n617_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n1155_, new_n1186_, new_n191_, new_n225_, new_n922_, new_n387_, new_n476_, new_n987_, new_n949_, new_n221_, new_n243_, new_n450_, new_n1179_, new_n298_, new_n184_, new_n1088_, new_n1148_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n203_, new_n316_, new_n590_, new_n826_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n307_, new_n190_, new_n1181_, new_n597_, new_n1093_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n435_, new_n1010_, new_n776_, new_n687_, new_n370_, new_n1029_, new_n638_, new_n523_, new_n909_, new_n217_, new_n788_, new_n841_, new_n1112_, new_n711_, new_n1156_, new_n731_, new_n599_, new_n930_, new_n973_, new_n412_, new_n607_, new_n645_, new_n1096_, new_n1087_, new_n723_, new_n756_, new_n823_, new_n574_, new_n928_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n294_, new_n1173_, new_n704_, new_n1189_, new_n1197_, new_n474_, new_n1223_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n866_, new_n947_, new_n994_, new_n982_, new_n964_, new_n1078_, new_n551_, new_n279_, new_n455_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n1103_;

not g0000 ( new_n172_, keyIn_0_21 );
or g0001 ( new_n173_, keyIn_0_12, N102 );
not g0002 ( new_n174_, N108 );
and g0003 ( new_n175_, keyIn_0_12, N102 );
or g0004 ( new_n176_, new_n175_, new_n174_ );
not g0005 ( new_n177_, new_n176_ );
and g0006 ( new_n178_, new_n177_, new_n173_ );
and g0007 ( new_n179_, new_n178_, new_n172_ );
not g0008 ( new_n180_, new_n179_ );
or g0009 ( new_n181_, new_n178_, new_n172_ );
and g0010 ( new_n182_, new_n180_, new_n181_ );
not g0011 ( new_n183_, new_n182_ );
not g0012 ( new_n184_, N95 );
not g0013 ( new_n185_, keyIn_0_11 );
or g0014 ( new_n186_, new_n185_, N89 );
not g0015 ( new_n187_, N89 );
or g0016 ( new_n188_, new_n187_, keyIn_0_11 );
and g0017 ( new_n189_, new_n186_, new_n188_ );
or g0018 ( new_n190_, new_n189_, new_n184_ );
and g0019 ( new_n191_, new_n190_, keyIn_0_20 );
not g0020 ( new_n192_, keyIn_0_20 );
and g0021 ( new_n193_, new_n187_, keyIn_0_11 );
and g0022 ( new_n194_, new_n185_, N89 );
or g0023 ( new_n195_, new_n193_, new_n194_ );
and g0024 ( new_n196_, new_n195_, N95 );
and g0025 ( new_n197_, new_n196_, new_n192_ );
or g0026 ( new_n198_, new_n191_, new_n197_ );
not g0027 ( new_n199_, keyIn_0_19 );
or g0028 ( new_n200_, keyIn_0_7, N50 );
not g0029 ( new_n201_, new_n200_ );
not g0030 ( new_n202_, N56 );
and g0031 ( new_n203_, keyIn_0_7, N50 );
or g0032 ( new_n204_, new_n203_, new_n202_ );
or g0033 ( new_n205_, new_n204_, new_n201_ );
and g0034 ( new_n206_, new_n205_, new_n199_ );
not g0035 ( new_n207_, new_n206_ );
or g0036 ( new_n208_, new_n205_, new_n199_ );
and g0037 ( new_n209_, new_n207_, new_n208_ );
or g0038 ( new_n210_, new_n198_, new_n209_ );
or g0039 ( new_n211_, new_n210_, new_n183_ );
not g0040 ( new_n212_, N4 );
and g0041 ( new_n213_, keyIn_0_0, N1 );
not g0042 ( new_n214_, new_n213_ );
or g0043 ( new_n215_, keyIn_0_0, N1 );
and g0044 ( new_n216_, new_n214_, new_n215_ );
or g0045 ( new_n217_, new_n216_, new_n212_ );
and g0046 ( new_n218_, new_n217_, keyIn_0_14 );
not g0047 ( new_n219_, keyIn_0_14 );
not g0048 ( new_n220_, keyIn_0_0 );
not g0049 ( new_n221_, N1 );
and g0050 ( new_n222_, new_n220_, new_n221_ );
or g0051 ( new_n223_, new_n222_, new_n213_ );
and g0052 ( new_n224_, new_n223_, N4 );
and g0053 ( new_n225_, new_n224_, new_n219_ );
or g0054 ( new_n226_, new_n218_, new_n225_ );
not g0055 ( new_n227_, keyIn_0_9 );
and g0056 ( new_n228_, new_n227_, N76 );
not g0057 ( new_n229_, new_n228_ );
or g0058 ( new_n230_, new_n227_, N76 );
and g0059 ( new_n231_, new_n230_, N82 );
and g0060 ( new_n232_, new_n231_, new_n229_ );
not g0061 ( new_n233_, keyIn_0_2 );
not g0062 ( new_n234_, N11 );
and g0063 ( new_n235_, new_n233_, new_n234_ );
and g0064 ( new_n236_, keyIn_0_2, N11 );
or g0065 ( new_n237_, new_n235_, new_n236_ );
and g0066 ( new_n238_, new_n237_, N17 );
not g0067 ( new_n239_, N63 );
and g0068 ( new_n240_, new_n239_, N69 );
or g0069 ( new_n241_, new_n238_, new_n240_ );
or g0070 ( new_n242_, new_n241_, new_n232_ );
or g0071 ( new_n243_, new_n226_, new_n242_ );
not g0072 ( new_n244_, keyIn_0_18 );
not g0073 ( new_n245_, N43 );
not g0074 ( new_n246_, keyIn_0_6 );
or g0075 ( new_n247_, new_n246_, N37 );
not g0076 ( new_n248_, N37 );
or g0077 ( new_n249_, new_n248_, keyIn_0_6 );
and g0078 ( new_n250_, new_n247_, new_n249_ );
or g0079 ( new_n251_, new_n250_, new_n245_ );
or g0080 ( new_n252_, new_n251_, new_n244_ );
and g0081 ( new_n253_, new_n248_, keyIn_0_6 );
and g0082 ( new_n254_, new_n246_, N37 );
or g0083 ( new_n255_, new_n253_, new_n254_ );
and g0084 ( new_n256_, new_n255_, N43 );
or g0085 ( new_n257_, new_n256_, keyIn_0_18 );
and g0086 ( new_n258_, new_n252_, new_n257_ );
not g0087 ( new_n259_, keyIn_0_17 );
or g0088 ( new_n260_, keyIn_0_4, N24 );
not g0089 ( new_n261_, new_n260_ );
not g0090 ( new_n262_, N30 );
and g0091 ( new_n263_, keyIn_0_4, N24 );
or g0092 ( new_n264_, new_n263_, new_n262_ );
or g0093 ( new_n265_, new_n264_, new_n261_ );
and g0094 ( new_n266_, new_n265_, new_n259_ );
not g0095 ( new_n267_, new_n266_ );
or g0096 ( new_n268_, new_n265_, new_n259_ );
and g0097 ( new_n269_, new_n267_, new_n268_ );
or g0098 ( new_n270_, new_n258_, new_n269_ );
or g0099 ( new_n271_, new_n243_, new_n270_ );
or g0100 ( new_n272_, new_n271_, new_n211_ );
and g0101 ( new_n273_, new_n272_, keyIn_0_38 );
not g0102 ( new_n274_, keyIn_0_38 );
or g0103 ( new_n275_, new_n196_, new_n192_ );
or g0104 ( new_n276_, new_n190_, keyIn_0_20 );
and g0105 ( new_n277_, new_n276_, new_n275_ );
not g0106 ( new_n278_, new_n204_ );
and g0107 ( new_n279_, new_n278_, new_n200_ );
and g0108 ( new_n280_, new_n279_, keyIn_0_19 );
or g0109 ( new_n281_, new_n280_, new_n206_ );
and g0110 ( new_n282_, new_n277_, new_n281_ );
and g0111 ( new_n283_, new_n282_, new_n182_ );
or g0112 ( new_n284_, new_n224_, new_n219_ );
or g0113 ( new_n285_, new_n217_, keyIn_0_14 );
and g0114 ( new_n286_, new_n284_, new_n285_ );
not g0115 ( new_n287_, new_n232_ );
not g0116 ( new_n288_, N17 );
or g0117 ( new_n289_, keyIn_0_2, N11 );
not g0118 ( new_n290_, new_n236_ );
and g0119 ( new_n291_, new_n290_, new_n289_ );
or g0120 ( new_n292_, new_n291_, new_n288_ );
not g0121 ( new_n293_, new_n240_ );
and g0122 ( new_n294_, new_n292_, new_n293_ );
and g0123 ( new_n295_, new_n294_, new_n287_ );
and g0124 ( new_n296_, new_n286_, new_n295_ );
and g0125 ( new_n297_, new_n256_, keyIn_0_18 );
and g0126 ( new_n298_, new_n251_, new_n244_ );
or g0127 ( new_n299_, new_n298_, new_n297_ );
not g0128 ( new_n300_, new_n264_ );
and g0129 ( new_n301_, new_n300_, new_n260_ );
and g0130 ( new_n302_, new_n301_, keyIn_0_17 );
or g0131 ( new_n303_, new_n302_, new_n266_ );
and g0132 ( new_n304_, new_n299_, new_n303_ );
and g0133 ( new_n305_, new_n304_, new_n296_ );
and g0134 ( new_n306_, new_n305_, new_n283_ );
and g0135 ( new_n307_, new_n306_, new_n274_ );
or g0136 ( N223, new_n273_, new_n307_ );
not g0137 ( new_n309_, keyIn_0_80 );
not g0138 ( new_n310_, keyIn_0_71 );
not g0139 ( new_n311_, keyIn_0_47 );
and g0140 ( new_n312_, new_n272_, keyIn_0_37 );
not g0141 ( new_n313_, keyIn_0_37 );
and g0142 ( new_n314_, new_n306_, new_n313_ );
or g0143 ( new_n315_, new_n312_, new_n314_ );
and g0144 ( new_n316_, new_n315_, new_n182_ );
and g0145 ( new_n317_, new_n183_, new_n313_ );
or g0146 ( new_n318_, new_n316_, new_n317_ );
and g0147 ( new_n319_, new_n318_, new_n311_ );
not g0148 ( new_n320_, new_n319_ );
or g0149 ( new_n321_, new_n318_, new_n311_ );
and g0150 ( new_n322_, new_n320_, new_n321_ );
not g0151 ( new_n323_, N112 );
and g0152 ( new_n324_, new_n174_, keyIn_0_13 );
not g0153 ( new_n325_, new_n324_ );
or g0154 ( new_n326_, new_n174_, keyIn_0_13 );
and g0155 ( new_n327_, new_n325_, new_n326_ );
and g0156 ( new_n328_, new_n327_, new_n323_ );
not g0157 ( new_n329_, new_n328_ );
and g0158 ( new_n330_, new_n329_, keyIn_0_35 );
not g0159 ( new_n331_, new_n330_ );
or g0160 ( new_n332_, new_n329_, keyIn_0_35 );
and g0161 ( new_n333_, new_n331_, new_n332_ );
not g0162 ( new_n334_, new_n333_ );
or g0163 ( new_n335_, new_n322_, new_n334_ );
and g0164 ( new_n336_, new_n335_, keyIn_0_62 );
not g0165 ( new_n337_, new_n336_ );
or g0166 ( new_n338_, new_n335_, keyIn_0_62 );
and g0167 ( new_n339_, new_n337_, new_n338_ );
not g0168 ( new_n340_, keyIn_0_59 );
and g0169 ( new_n341_, new_n315_, new_n293_ );
or g0170 ( new_n342_, new_n306_, new_n313_ );
not g0171 ( new_n343_, new_n314_ );
and g0172 ( new_n344_, new_n343_, new_n342_ );
and g0173 ( new_n345_, new_n344_, new_n240_ );
or g0174 ( new_n346_, new_n341_, new_n345_ );
or g0175 ( new_n347_, new_n346_, keyIn_0_43 );
not g0176 ( new_n348_, keyIn_0_43 );
or g0177 ( new_n349_, new_n344_, new_n240_ );
or g0178 ( new_n350_, new_n315_, new_n293_ );
and g0179 ( new_n351_, new_n350_, new_n349_ );
or g0180 ( new_n352_, new_n351_, new_n348_ );
and g0181 ( new_n353_, new_n347_, new_n352_ );
not g0182 ( new_n354_, N73 );
and g0183 ( new_n355_, new_n354_, N69 );
not g0184 ( new_n356_, new_n355_ );
and g0185 ( new_n357_, new_n356_, keyIn_0_29 );
not g0186 ( new_n358_, new_n357_ );
or g0187 ( new_n359_, new_n356_, keyIn_0_29 );
and g0188 ( new_n360_, new_n358_, new_n359_ );
not g0189 ( new_n361_, new_n360_ );
or g0190 ( new_n362_, new_n353_, new_n361_ );
or g0191 ( new_n363_, new_n362_, new_n340_ );
and g0192 ( new_n364_, new_n351_, new_n348_ );
and g0193 ( new_n365_, new_n346_, keyIn_0_43 );
or g0194 ( new_n366_, new_n365_, new_n364_ );
and g0195 ( new_n367_, new_n366_, new_n360_ );
or g0196 ( new_n368_, new_n367_, keyIn_0_59 );
and g0197 ( new_n369_, new_n363_, new_n368_ );
not g0198 ( new_n370_, keyIn_0_61 );
and g0199 ( new_n371_, new_n315_, new_n277_ );
and g0200 ( new_n372_, new_n344_, new_n198_ );
or g0201 ( new_n373_, new_n371_, new_n372_ );
or g0202 ( new_n374_, new_n373_, keyIn_0_45 );
not g0203 ( new_n375_, keyIn_0_45 );
or g0204 ( new_n376_, new_n344_, new_n198_ );
or g0205 ( new_n377_, new_n315_, new_n277_ );
and g0206 ( new_n378_, new_n377_, new_n376_ );
or g0207 ( new_n379_, new_n378_, new_n375_ );
and g0208 ( new_n380_, new_n374_, new_n379_ );
not g0209 ( new_n381_, N99 );
and g0210 ( new_n382_, new_n381_, N95 );
not g0211 ( new_n383_, new_n382_ );
and g0212 ( new_n384_, new_n383_, keyIn_0_33 );
not g0213 ( new_n385_, new_n384_ );
or g0214 ( new_n386_, new_n383_, keyIn_0_33 );
and g0215 ( new_n387_, new_n385_, new_n386_ );
or g0216 ( new_n388_, new_n380_, new_n387_ );
or g0217 ( new_n389_, new_n388_, new_n370_ );
and g0218 ( new_n390_, new_n378_, new_n375_ );
and g0219 ( new_n391_, new_n373_, keyIn_0_45 );
or g0220 ( new_n392_, new_n391_, new_n390_ );
not g0221 ( new_n393_, new_n387_ );
and g0222 ( new_n394_, new_n392_, new_n393_ );
or g0223 ( new_n395_, new_n394_, keyIn_0_61 );
and g0224 ( new_n396_, new_n389_, new_n395_ );
or g0225 ( new_n397_, new_n369_, new_n396_ );
or g0226 ( new_n398_, new_n397_, new_n339_ );
not g0227 ( new_n399_, keyIn_0_57 );
and g0228 ( new_n400_, new_n315_, new_n303_ );
and g0229 ( new_n401_, new_n344_, new_n269_ );
or g0230 ( new_n402_, new_n400_, new_n401_ );
and g0231 ( new_n403_, new_n402_, keyIn_0_40 );
not g0232 ( new_n404_, keyIn_0_40 );
or g0233 ( new_n405_, new_n344_, new_n269_ );
or g0234 ( new_n406_, new_n315_, new_n303_ );
and g0235 ( new_n407_, new_n406_, new_n405_ );
and g0236 ( new_n408_, new_n407_, new_n404_ );
or g0237 ( new_n409_, new_n403_, new_n408_ );
not g0238 ( new_n410_, N34 );
and g0239 ( new_n411_, new_n262_, keyIn_0_5 );
not g0240 ( new_n412_, new_n411_ );
or g0241 ( new_n413_, new_n262_, keyIn_0_5 );
and g0242 ( new_n414_, new_n412_, new_n413_ );
not g0243 ( new_n415_, new_n414_ );
and g0244 ( new_n416_, new_n415_, new_n410_ );
and g0245 ( new_n417_, new_n416_, keyIn_0_23 );
not g0246 ( new_n418_, new_n417_ );
or g0247 ( new_n419_, new_n416_, keyIn_0_23 );
and g0248 ( new_n420_, new_n418_, new_n419_ );
not g0249 ( new_n421_, new_n420_ );
or g0250 ( new_n422_, new_n409_, new_n421_ );
or g0251 ( new_n423_, new_n422_, new_n399_ );
or g0252 ( new_n424_, new_n407_, new_n404_ );
or g0253 ( new_n425_, new_n402_, keyIn_0_40 );
and g0254 ( new_n426_, new_n425_, new_n424_ );
and g0255 ( new_n427_, new_n426_, new_n420_ );
or g0256 ( new_n428_, new_n427_, keyIn_0_57 );
and g0257 ( new_n429_, new_n423_, new_n428_ );
and g0258 ( new_n430_, new_n315_, new_n287_ );
and g0259 ( new_n431_, new_n344_, new_n232_ );
or g0260 ( new_n432_, new_n430_, new_n431_ );
not g0261 ( new_n433_, N86 );
not g0262 ( new_n434_, N82 );
and g0263 ( new_n435_, new_n434_, keyIn_0_10 );
not g0264 ( new_n436_, new_n435_ );
or g0265 ( new_n437_, new_n434_, keyIn_0_10 );
and g0266 ( new_n438_, new_n436_, new_n437_ );
and g0267 ( new_n439_, new_n438_, new_n433_ );
not g0268 ( new_n440_, new_n439_ );
and g0269 ( new_n441_, new_n440_, keyIn_0_31 );
not g0270 ( new_n442_, new_n441_ );
or g0271 ( new_n443_, new_n440_, keyIn_0_31 );
and g0272 ( new_n444_, new_n442_, new_n443_ );
and g0273 ( new_n445_, new_n432_, new_n444_ );
and g0274 ( new_n446_, new_n445_, keyIn_0_60 );
not g0275 ( new_n447_, new_n446_ );
or g0276 ( new_n448_, new_n445_, keyIn_0_60 );
and g0277 ( new_n449_, new_n447_, new_n448_ );
not g0278 ( new_n450_, new_n449_ );
or g0279 ( new_n451_, new_n315_, new_n286_ );
or g0280 ( new_n452_, new_n344_, new_n226_ );
and g0281 ( new_n453_, new_n451_, new_n452_ );
not g0282 ( new_n454_, N8 );
and g0283 ( new_n455_, new_n212_, keyIn_0_1 );
not g0284 ( new_n456_, new_n455_ );
or g0285 ( new_n457_, new_n212_, keyIn_0_1 );
and g0286 ( new_n458_, new_n456_, new_n457_ );
and g0287 ( new_n459_, new_n458_, new_n454_ );
not g0288 ( new_n460_, new_n459_ );
and g0289 ( new_n461_, new_n460_, keyIn_0_15 );
not g0290 ( new_n462_, new_n461_ );
or g0291 ( new_n463_, new_n460_, keyIn_0_15 );
and g0292 ( new_n464_, new_n462_, new_n463_ );
or g0293 ( new_n465_, new_n453_, new_n464_ );
and g0294 ( new_n466_, new_n465_, keyIn_0_54 );
not g0295 ( new_n467_, keyIn_0_54 );
and g0296 ( new_n468_, new_n344_, new_n226_ );
and g0297 ( new_n469_, new_n315_, new_n286_ );
or g0298 ( new_n470_, new_n469_, new_n468_ );
not g0299 ( new_n471_, new_n464_ );
and g0300 ( new_n472_, new_n470_, new_n471_ );
and g0301 ( new_n473_, new_n472_, new_n467_ );
or g0302 ( new_n474_, new_n466_, new_n473_ );
not g0303 ( new_n475_, keyIn_0_42 );
and g0304 ( new_n476_, new_n315_, new_n281_ );
and g0305 ( new_n477_, new_n344_, new_n209_ );
or g0306 ( new_n478_, new_n476_, new_n477_ );
or g0307 ( new_n479_, new_n478_, new_n475_ );
or g0308 ( new_n480_, new_n344_, new_n209_ );
or g0309 ( new_n481_, new_n315_, new_n281_ );
and g0310 ( new_n482_, new_n481_, new_n480_ );
or g0311 ( new_n483_, new_n482_, keyIn_0_42 );
and g0312 ( new_n484_, new_n479_, new_n483_ );
not g0313 ( new_n485_, N60 );
and g0314 ( new_n486_, keyIn_0_8, N56 );
not g0315 ( new_n487_, new_n486_ );
or g0316 ( new_n488_, keyIn_0_8, N56 );
and g0317 ( new_n489_, new_n487_, new_n488_ );
not g0318 ( new_n490_, new_n489_ );
and g0319 ( new_n491_, new_n490_, new_n485_ );
and g0320 ( new_n492_, new_n491_, keyIn_0_27 );
not g0321 ( new_n493_, new_n492_ );
or g0322 ( new_n494_, new_n491_, keyIn_0_27 );
and g0323 ( new_n495_, new_n493_, new_n494_ );
and g0324 ( new_n496_, new_n484_, new_n495_ );
or g0325 ( new_n497_, new_n474_, new_n496_ );
or g0326 ( new_n498_, new_n497_, new_n450_ );
or g0327 ( new_n499_, new_n498_, new_n429_ );
not g0328 ( new_n500_, keyIn_0_58 );
and g0329 ( new_n501_, new_n315_, new_n299_ );
and g0330 ( new_n502_, new_n344_, new_n258_ );
or g0331 ( new_n503_, new_n501_, new_n502_ );
and g0332 ( new_n504_, new_n503_, keyIn_0_41 );
not g0333 ( new_n505_, keyIn_0_41 );
or g0334 ( new_n506_, new_n344_, new_n258_ );
or g0335 ( new_n507_, new_n315_, new_n299_ );
and g0336 ( new_n508_, new_n507_, new_n506_ );
and g0337 ( new_n509_, new_n508_, new_n505_ );
or g0338 ( new_n510_, new_n504_, new_n509_ );
not g0339 ( new_n511_, N47 );
and g0340 ( new_n512_, new_n511_, N43 );
not g0341 ( new_n513_, new_n512_ );
and g0342 ( new_n514_, new_n513_, keyIn_0_25 );
not g0343 ( new_n515_, new_n514_ );
or g0344 ( new_n516_, new_n513_, keyIn_0_25 );
and g0345 ( new_n517_, new_n515_, new_n516_ );
not g0346 ( new_n518_, new_n517_ );
or g0347 ( new_n519_, new_n510_, new_n518_ );
and g0348 ( new_n520_, new_n519_, new_n500_ );
or g0349 ( new_n521_, new_n508_, new_n505_ );
or g0350 ( new_n522_, new_n503_, keyIn_0_41 );
and g0351 ( new_n523_, new_n522_, new_n521_ );
and g0352 ( new_n524_, new_n523_, new_n517_ );
and g0353 ( new_n525_, new_n524_, keyIn_0_58 );
or g0354 ( new_n526_, new_n520_, new_n525_ );
not g0355 ( new_n527_, keyIn_0_39 );
and g0356 ( new_n528_, new_n315_, new_n292_ );
and g0357 ( new_n529_, new_n344_, new_n238_ );
or g0358 ( new_n530_, new_n528_, new_n529_ );
or g0359 ( new_n531_, new_n530_, new_n527_ );
or g0360 ( new_n532_, new_n344_, new_n238_ );
or g0361 ( new_n533_, new_n315_, new_n292_ );
and g0362 ( new_n534_, new_n533_, new_n532_ );
or g0363 ( new_n535_, new_n534_, keyIn_0_39 );
and g0364 ( new_n536_, new_n531_, new_n535_ );
not g0365 ( new_n537_, N21 );
and g0366 ( new_n538_, keyIn_0_3, N17 );
not g0367 ( new_n539_, new_n538_ );
or g0368 ( new_n540_, keyIn_0_3, N17 );
and g0369 ( new_n541_, new_n539_, new_n540_ );
and g0370 ( new_n542_, new_n541_, new_n537_ );
not g0371 ( new_n543_, new_n542_ );
and g0372 ( new_n544_, new_n543_, keyIn_0_22 );
not g0373 ( new_n545_, new_n544_ );
or g0374 ( new_n546_, new_n543_, keyIn_0_22 );
and g0375 ( new_n547_, new_n545_, new_n546_ );
or g0376 ( new_n548_, new_n536_, new_n547_ );
or g0377 ( new_n549_, new_n548_, keyIn_0_56 );
not g0378 ( new_n550_, keyIn_0_56 );
and g0379 ( new_n551_, new_n534_, keyIn_0_39 );
and g0380 ( new_n552_, new_n530_, new_n527_ );
or g0381 ( new_n553_, new_n552_, new_n551_ );
not g0382 ( new_n554_, new_n547_ );
and g0383 ( new_n555_, new_n553_, new_n554_ );
or g0384 ( new_n556_, new_n555_, new_n550_ );
and g0385 ( new_n557_, new_n549_, new_n556_ );
or g0386 ( new_n558_, new_n526_, new_n557_ );
or g0387 ( new_n559_, new_n499_, new_n558_ );
or g0388 ( new_n560_, new_n559_, new_n398_ );
and g0389 ( new_n561_, new_n560_, new_n310_ );
not g0390 ( new_n562_, new_n338_ );
or g0391 ( new_n563_, new_n562_, new_n336_ );
and g0392 ( new_n564_, new_n367_, keyIn_0_59 );
and g0393 ( new_n565_, new_n362_, new_n340_ );
or g0394 ( new_n566_, new_n565_, new_n564_ );
and g0395 ( new_n567_, new_n394_, keyIn_0_61 );
and g0396 ( new_n568_, new_n388_, new_n370_ );
or g0397 ( new_n569_, new_n568_, new_n567_ );
and g0398 ( new_n570_, new_n566_, new_n569_ );
and g0399 ( new_n571_, new_n570_, new_n563_ );
and g0400 ( new_n572_, new_n427_, keyIn_0_57 );
and g0401 ( new_n573_, new_n422_, new_n399_ );
or g0402 ( new_n574_, new_n573_, new_n572_ );
or g0403 ( new_n575_, new_n472_, new_n467_ );
or g0404 ( new_n576_, new_n465_, keyIn_0_54 );
and g0405 ( new_n577_, new_n576_, new_n575_ );
and g0406 ( new_n578_, new_n482_, keyIn_0_42 );
and g0407 ( new_n579_, new_n478_, new_n475_ );
or g0408 ( new_n580_, new_n579_, new_n578_ );
not g0409 ( new_n581_, new_n495_ );
or g0410 ( new_n582_, new_n580_, new_n581_ );
and g0411 ( new_n583_, new_n582_, new_n577_ );
and g0412 ( new_n584_, new_n583_, new_n449_ );
and g0413 ( new_n585_, new_n574_, new_n584_ );
or g0414 ( new_n586_, new_n524_, keyIn_0_58 );
or g0415 ( new_n587_, new_n519_, new_n500_ );
and g0416 ( new_n588_, new_n587_, new_n586_ );
and g0417 ( new_n589_, new_n555_, new_n550_ );
and g0418 ( new_n590_, new_n548_, keyIn_0_56 );
or g0419 ( new_n591_, new_n590_, new_n589_ );
and g0420 ( new_n592_, new_n591_, new_n588_ );
and g0421 ( new_n593_, new_n592_, new_n585_ );
and g0422 ( new_n594_, new_n571_, new_n593_ );
and g0423 ( new_n595_, new_n594_, keyIn_0_71 );
or g0424 ( new_n596_, new_n561_, new_n595_ );
and g0425 ( new_n597_, new_n596_, new_n309_ );
or g0426 ( new_n598_, new_n594_, keyIn_0_71 );
not g0427 ( new_n599_, new_n595_ );
and g0428 ( new_n600_, new_n599_, new_n598_ );
and g0429 ( new_n601_, new_n600_, keyIn_0_80 );
or g0430 ( N329, new_n597_, new_n601_ );
not g0431 ( new_n603_, keyIn_0_83 );
and g0432 ( new_n604_, new_n596_, keyIn_0_78 );
not g0433 ( new_n605_, keyIn_0_78 );
and g0434 ( new_n606_, new_n600_, new_n605_ );
or g0435 ( new_n607_, new_n604_, new_n606_ );
and g0436 ( new_n608_, new_n607_, new_n582_ );
or g0437 ( new_n609_, new_n600_, new_n605_ );
or g0438 ( new_n610_, new_n596_, keyIn_0_78 );
and g0439 ( new_n611_, new_n610_, new_n609_ );
and g0440 ( new_n612_, new_n611_, new_n496_ );
or g0441 ( new_n613_, new_n608_, new_n612_ );
and g0442 ( new_n614_, new_n613_, new_n603_ );
not g0443 ( new_n615_, new_n614_ );
or g0444 ( new_n616_, new_n613_, new_n603_ );
and g0445 ( new_n617_, new_n615_, new_n616_ );
not g0446 ( new_n618_, N66 );
and g0447 ( new_n619_, new_n490_, new_n618_ );
and g0448 ( new_n620_, new_n619_, keyIn_0_28 );
not g0449 ( new_n621_, new_n620_ );
or g0450 ( new_n622_, new_n619_, keyIn_0_28 );
and g0451 ( new_n623_, new_n621_, new_n622_ );
or g0452 ( new_n624_, new_n580_, new_n623_ );
not g0453 ( new_n625_, new_n624_ );
and g0454 ( new_n626_, new_n625_, keyIn_0_66 );
not g0455 ( new_n627_, new_n626_ );
or g0456 ( new_n628_, new_n625_, keyIn_0_66 );
and g0457 ( new_n629_, new_n627_, new_n628_ );
or g0458 ( new_n630_, new_n617_, new_n629_ );
and g0459 ( new_n631_, new_n607_, new_n449_ );
and g0460 ( new_n632_, new_n611_, new_n450_ );
or g0461 ( new_n633_, new_n631_, new_n632_ );
and g0462 ( new_n634_, new_n633_, keyIn_0_86 );
not g0463 ( new_n635_, new_n634_ );
or g0464 ( new_n636_, new_n633_, keyIn_0_86 );
and g0465 ( new_n637_, new_n635_, new_n636_ );
not g0466 ( new_n638_, new_n432_ );
not g0467 ( new_n639_, N92 );
and g0468 ( new_n640_, new_n438_, new_n639_ );
and g0469 ( new_n641_, new_n640_, keyIn_0_32 );
not g0470 ( new_n642_, new_n641_ );
or g0471 ( new_n643_, new_n640_, keyIn_0_32 );
and g0472 ( new_n644_, new_n642_, new_n643_ );
or g0473 ( new_n645_, new_n638_, new_n644_ );
not g0474 ( new_n646_, new_n645_ );
and g0475 ( new_n647_, new_n646_, keyIn_0_68 );
not g0476 ( new_n648_, new_n647_ );
or g0477 ( new_n649_, new_n646_, keyIn_0_68 );
and g0478 ( new_n650_, new_n648_, new_n649_ );
and g0479 ( new_n651_, new_n650_, keyIn_0_75 );
not g0480 ( new_n652_, new_n651_ );
or g0481 ( new_n653_, new_n650_, keyIn_0_75 );
and g0482 ( new_n654_, new_n652_, new_n653_ );
or g0483 ( new_n655_, new_n637_, new_n654_ );
and g0484 ( new_n656_, new_n630_, new_n655_ );
not g0485 ( new_n657_, new_n656_ );
and g0486 ( new_n658_, new_n607_, new_n588_ );
and g0487 ( new_n659_, new_n611_, new_n526_ );
or g0488 ( new_n660_, new_n658_, new_n659_ );
not g0489 ( new_n661_, N53 );
and g0490 ( new_n662_, new_n661_, N43 );
and g0491 ( new_n663_, new_n662_, keyIn_0_26 );
not g0492 ( new_n664_, new_n663_ );
or g0493 ( new_n665_, new_n662_, keyIn_0_26 );
and g0494 ( new_n666_, new_n664_, new_n665_ );
and g0495 ( new_n667_, new_n523_, new_n666_ );
and g0496 ( new_n668_, new_n667_, keyIn_0_65 );
not g0497 ( new_n669_, new_n668_ );
or g0498 ( new_n670_, new_n667_, keyIn_0_65 );
and g0499 ( new_n671_, new_n669_, new_n670_ );
and g0500 ( new_n672_, new_n660_, new_n671_ );
not g0501 ( new_n673_, new_n672_ );
and g0502 ( new_n674_, new_n673_, keyIn_0_96 );
not g0503 ( new_n675_, new_n674_ );
or g0504 ( new_n676_, new_n673_, keyIn_0_96 );
and g0505 ( new_n677_, new_n675_, new_n676_ );
and g0506 ( new_n678_, new_n607_, new_n574_ );
and g0507 ( new_n679_, new_n611_, new_n429_ );
or g0508 ( new_n680_, new_n678_, new_n679_ );
not g0509 ( new_n681_, N40 );
and g0510 ( new_n682_, new_n415_, new_n681_ );
not g0511 ( new_n683_, new_n682_ );
and g0512 ( new_n684_, new_n683_, keyIn_0_24 );
not g0513 ( new_n685_, new_n684_ );
or g0514 ( new_n686_, new_n683_, keyIn_0_24 );
and g0515 ( new_n687_, new_n685_, new_n686_ );
or g0516 ( new_n688_, new_n409_, new_n687_ );
and g0517 ( new_n689_, new_n688_, keyIn_0_64 );
not g0518 ( new_n690_, new_n689_ );
or g0519 ( new_n691_, new_n688_, keyIn_0_64 );
and g0520 ( new_n692_, new_n690_, new_n691_ );
not g0521 ( new_n693_, new_n692_ );
and g0522 ( new_n694_, new_n693_, keyIn_0_73 );
not g0523 ( new_n695_, new_n694_ );
or g0524 ( new_n696_, new_n693_, keyIn_0_73 );
and g0525 ( new_n697_, new_n695_, new_n696_ );
not g0526 ( new_n698_, new_n697_ );
and g0527 ( new_n699_, new_n680_, new_n698_ );
and g0528 ( new_n700_, new_n699_, keyIn_0_95 );
not g0529 ( new_n701_, new_n700_ );
or g0530 ( new_n702_, new_n699_, keyIn_0_95 );
and g0531 ( new_n703_, new_n701_, new_n702_ );
or g0532 ( new_n704_, new_n677_, new_n703_ );
or g0533 ( new_n705_, new_n657_, new_n704_ );
not g0534 ( new_n706_, keyIn_0_82 );
and g0535 ( new_n707_, new_n607_, new_n591_ );
and g0536 ( new_n708_, new_n611_, new_n557_ );
or g0537 ( new_n709_, new_n707_, new_n708_ );
and g0538 ( new_n710_, new_n709_, new_n706_ );
not g0539 ( new_n711_, new_n710_ );
or g0540 ( new_n712_, new_n709_, new_n706_ );
not g0541 ( new_n713_, N27 );
and g0542 ( new_n714_, new_n541_, new_n713_ );
and g0543 ( new_n715_, new_n553_, new_n714_ );
and g0544 ( new_n716_, new_n715_, keyIn_0_63 );
not g0545 ( new_n717_, new_n716_ );
or g0546 ( new_n718_, new_n715_, keyIn_0_63 );
and g0547 ( new_n719_, new_n717_, new_n718_ );
not g0548 ( new_n720_, new_n719_ );
and g0549 ( new_n721_, new_n712_, new_n720_ );
and g0550 ( new_n722_, new_n721_, new_n711_ );
and g0551 ( new_n723_, new_n722_, keyIn_0_94 );
not g0552 ( new_n724_, new_n723_ );
or g0553 ( new_n725_, new_n722_, keyIn_0_94 );
and g0554 ( new_n726_, new_n724_, new_n725_ );
not g0555 ( new_n727_, new_n726_ );
or g0556 ( new_n728_, new_n705_, new_n727_ );
not g0557 ( new_n729_, keyIn_0_98 );
and g0558 ( new_n730_, new_n607_, new_n569_ );
and g0559 ( new_n731_, new_n611_, new_n396_ );
or g0560 ( new_n732_, new_n730_, new_n731_ );
or g0561 ( new_n733_, new_n732_, keyIn_0_88 );
not g0562 ( new_n734_, keyIn_0_88 );
or g0563 ( new_n735_, new_n611_, new_n396_ );
or g0564 ( new_n736_, new_n607_, new_n569_ );
and g0565 ( new_n737_, new_n736_, new_n735_ );
or g0566 ( new_n738_, new_n737_, new_n734_ );
and g0567 ( new_n739_, new_n733_, new_n738_ );
not g0568 ( new_n740_, N105 );
and g0569 ( new_n741_, new_n740_, N95 );
and g0570 ( new_n742_, new_n741_, keyIn_0_34 );
not g0571 ( new_n743_, new_n742_ );
or g0572 ( new_n744_, new_n741_, keyIn_0_34 );
and g0573 ( new_n745_, new_n743_, new_n744_ );
or g0574 ( new_n746_, new_n380_, new_n745_ );
and g0575 ( new_n747_, new_n746_, keyIn_0_69 );
not g0576 ( new_n748_, new_n747_ );
or g0577 ( new_n749_, new_n746_, keyIn_0_69 );
and g0578 ( new_n750_, new_n748_, new_n749_ );
and g0579 ( new_n751_, new_n750_, keyIn_0_76 );
not g0580 ( new_n752_, new_n751_ );
or g0581 ( new_n753_, new_n750_, keyIn_0_76 );
and g0582 ( new_n754_, new_n752_, new_n753_ );
not g0583 ( new_n755_, new_n754_ );
or g0584 ( new_n756_, new_n739_, new_n755_ );
or g0585 ( new_n757_, new_n756_, new_n729_ );
and g0586 ( new_n758_, new_n737_, new_n734_ );
and g0587 ( new_n759_, new_n732_, keyIn_0_88 );
or g0588 ( new_n760_, new_n759_, new_n758_ );
and g0589 ( new_n761_, new_n760_, new_n754_ );
or g0590 ( new_n762_, new_n761_, keyIn_0_98 );
and g0591 ( new_n763_, new_n757_, new_n762_ );
not g0592 ( new_n764_, keyIn_0_90 );
and g0593 ( new_n765_, new_n607_, new_n563_ );
and g0594 ( new_n766_, new_n611_, new_n339_ );
or g0595 ( new_n767_, new_n765_, new_n766_ );
or g0596 ( new_n768_, new_n767_, new_n764_ );
or g0597 ( new_n769_, new_n611_, new_n339_ );
or g0598 ( new_n770_, new_n607_, new_n563_ );
and g0599 ( new_n771_, new_n770_, new_n769_ );
or g0600 ( new_n772_, new_n771_, keyIn_0_90 );
and g0601 ( new_n773_, new_n768_, new_n772_ );
not g0602 ( new_n774_, N115 );
and g0603 ( new_n775_, new_n327_, new_n774_ );
not g0604 ( new_n776_, new_n775_ );
and g0605 ( new_n777_, new_n776_, keyIn_0_36 );
not g0606 ( new_n778_, new_n777_ );
or g0607 ( new_n779_, new_n776_, keyIn_0_36 );
and g0608 ( new_n780_, new_n778_, new_n779_ );
or g0609 ( new_n781_, new_n322_, new_n780_ );
not g0610 ( new_n782_, new_n781_ );
and g0611 ( new_n783_, new_n782_, keyIn_0_70 );
not g0612 ( new_n784_, new_n783_ );
or g0613 ( new_n785_, new_n782_, keyIn_0_70 );
and g0614 ( new_n786_, new_n784_, new_n785_ );
not g0615 ( new_n787_, new_n786_ );
and g0616 ( new_n788_, new_n787_, keyIn_0_77 );
not g0617 ( new_n789_, new_n788_ );
or g0618 ( new_n790_, new_n787_, keyIn_0_77 );
and g0619 ( new_n791_, new_n789_, new_n790_ );
or g0620 ( new_n792_, new_n773_, new_n791_ );
or g0621 ( new_n793_, new_n792_, keyIn_0_99 );
not g0622 ( new_n794_, keyIn_0_99 );
and g0623 ( new_n795_, new_n771_, keyIn_0_90 );
and g0624 ( new_n796_, new_n767_, new_n764_ );
or g0625 ( new_n797_, new_n796_, new_n795_ );
not g0626 ( new_n798_, new_n791_ );
and g0627 ( new_n799_, new_n797_, new_n798_ );
or g0628 ( new_n800_, new_n799_, new_n794_ );
and g0629 ( new_n801_, new_n793_, new_n800_ );
or g0630 ( new_n802_, new_n763_, new_n801_ );
not g0631 ( new_n803_, keyIn_0_93 );
not g0632 ( new_n804_, keyIn_0_81 );
and g0633 ( new_n805_, new_n611_, new_n474_ );
and g0634 ( new_n806_, new_n607_, new_n577_ );
or g0635 ( new_n807_, new_n806_, new_n805_ );
and g0636 ( new_n808_, new_n807_, new_n804_ );
or g0637 ( new_n809_, new_n607_, new_n577_ );
or g0638 ( new_n810_, new_n611_, new_n474_ );
and g0639 ( new_n811_, new_n809_, new_n810_ );
and g0640 ( new_n812_, new_n811_, keyIn_0_81 );
not g0641 ( new_n813_, N14 );
and g0642 ( new_n814_, new_n458_, new_n813_ );
not g0643 ( new_n815_, new_n814_ );
and g0644 ( new_n816_, new_n815_, keyIn_0_16 );
not g0645 ( new_n817_, new_n816_ );
or g0646 ( new_n818_, new_n815_, keyIn_0_16 );
and g0647 ( new_n819_, new_n817_, new_n818_ );
or g0648 ( new_n820_, new_n453_, new_n819_ );
and g0649 ( new_n821_, new_n820_, keyIn_0_55 );
not g0650 ( new_n822_, new_n821_ );
or g0651 ( new_n823_, new_n820_, keyIn_0_55 );
and g0652 ( new_n824_, new_n822_, new_n823_ );
and g0653 ( new_n825_, new_n824_, keyIn_0_72 );
not g0654 ( new_n826_, new_n825_ );
or g0655 ( new_n827_, new_n824_, keyIn_0_72 );
and g0656 ( new_n828_, new_n826_, new_n827_ );
not g0657 ( new_n829_, new_n828_ );
or g0658 ( new_n830_, new_n812_, new_n829_ );
or g0659 ( new_n831_, new_n830_, new_n808_ );
or g0660 ( new_n832_, new_n831_, new_n803_ );
not g0661 ( new_n833_, new_n808_ );
or g0662 ( new_n834_, new_n807_, new_n804_ );
and g0663 ( new_n835_, new_n834_, new_n828_ );
and g0664 ( new_n836_, new_n835_, new_n833_ );
or g0665 ( new_n837_, new_n836_, keyIn_0_93 );
and g0666 ( new_n838_, new_n832_, new_n837_ );
not g0667 ( new_n839_, keyIn_0_85 );
and g0668 ( new_n840_, new_n611_, new_n369_ );
and g0669 ( new_n841_, new_n607_, new_n566_ );
or g0670 ( new_n842_, new_n841_, new_n840_ );
and g0671 ( new_n843_, new_n842_, new_n839_ );
or g0672 ( new_n844_, new_n607_, new_n566_ );
or g0673 ( new_n845_, new_n611_, new_n369_ );
and g0674 ( new_n846_, new_n844_, new_n845_ );
and g0675 ( new_n847_, new_n846_, keyIn_0_85 );
not g0676 ( new_n848_, N79 );
and g0677 ( new_n849_, new_n848_, N69 );
and g0678 ( new_n850_, new_n849_, keyIn_0_30 );
not g0679 ( new_n851_, new_n850_ );
or g0680 ( new_n852_, new_n849_, keyIn_0_30 );
and g0681 ( new_n853_, new_n851_, new_n852_ );
or g0682 ( new_n854_, new_n353_, new_n853_ );
not g0683 ( new_n855_, new_n854_ );
and g0684 ( new_n856_, new_n855_, keyIn_0_67 );
not g0685 ( new_n857_, new_n856_ );
or g0686 ( new_n858_, new_n855_, keyIn_0_67 );
and g0687 ( new_n859_, new_n857_, new_n858_ );
not g0688 ( new_n860_, new_n859_ );
and g0689 ( new_n861_, new_n860_, keyIn_0_74 );
not g0690 ( new_n862_, new_n861_ );
or g0691 ( new_n863_, new_n860_, keyIn_0_74 );
and g0692 ( new_n864_, new_n862_, new_n863_ );
or g0693 ( new_n865_, new_n847_, new_n864_ );
or g0694 ( new_n866_, new_n865_, new_n843_ );
or g0695 ( new_n867_, new_n866_, keyIn_0_97 );
not g0696 ( new_n868_, keyIn_0_97 );
not g0697 ( new_n869_, new_n843_ );
or g0698 ( new_n870_, new_n842_, new_n839_ );
not g0699 ( new_n871_, new_n864_ );
and g0700 ( new_n872_, new_n870_, new_n871_ );
and g0701 ( new_n873_, new_n872_, new_n869_ );
or g0702 ( new_n874_, new_n873_, new_n868_ );
and g0703 ( new_n875_, new_n867_, new_n874_ );
or g0704 ( new_n876_, new_n838_, new_n875_ );
or g0705 ( new_n877_, new_n802_, new_n876_ );
or g0706 ( N370, new_n877_, new_n728_ );
not g0707 ( new_n879_, keyIn_0_115 );
not g0708 ( new_n880_, keyIn_0_114 );
not g0709 ( new_n881_, keyIn_0_100 );
not g0710 ( new_n882_, new_n677_ );
not g0711 ( new_n883_, new_n703_ );
and g0712 ( new_n884_, new_n882_, new_n883_ );
and g0713 ( new_n885_, new_n884_, new_n656_ );
and g0714 ( new_n886_, new_n885_, new_n726_ );
and g0715 ( new_n887_, new_n761_, keyIn_0_98 );
and g0716 ( new_n888_, new_n756_, new_n729_ );
or g0717 ( new_n889_, new_n888_, new_n887_ );
and g0718 ( new_n890_, new_n799_, new_n794_ );
and g0719 ( new_n891_, new_n792_, keyIn_0_99 );
or g0720 ( new_n892_, new_n891_, new_n890_ );
and g0721 ( new_n893_, new_n889_, new_n892_ );
and g0722 ( new_n894_, new_n836_, keyIn_0_93 );
and g0723 ( new_n895_, new_n831_, new_n803_ );
or g0724 ( new_n896_, new_n895_, new_n894_ );
and g0725 ( new_n897_, new_n873_, new_n868_ );
and g0726 ( new_n898_, new_n866_, keyIn_0_97 );
or g0727 ( new_n899_, new_n898_, new_n897_ );
and g0728 ( new_n900_, new_n896_, new_n899_ );
and g0729 ( new_n901_, new_n893_, new_n900_ );
and g0730 ( new_n902_, new_n901_, new_n886_ );
and g0731 ( new_n903_, new_n902_, new_n881_ );
and g0732 ( new_n904_, N370, keyIn_0_100 );
or g0733 ( new_n905_, new_n904_, new_n903_ );
or g0734 ( new_n906_, new_n905_, new_n639_ );
or g0735 ( new_n907_, new_n906_, keyIn_0_107 );
not g0736 ( new_n908_, keyIn_0_107 );
not g0737 ( new_n909_, new_n903_ );
or g0738 ( new_n910_, new_n902_, new_n881_ );
and g0739 ( new_n911_, new_n909_, new_n910_ );
and g0740 ( new_n912_, new_n911_, N92 );
or g0741 ( new_n913_, new_n912_, new_n908_ );
and g0742 ( new_n914_, new_n907_, new_n913_ );
and g0743 ( new_n915_, new_n600_, keyIn_0_79 );
not g0744 ( new_n916_, new_n915_ );
or g0745 ( new_n917_, new_n600_, keyIn_0_79 );
and g0746 ( new_n918_, new_n916_, new_n917_ );
and g0747 ( new_n919_, new_n918_, N86 );
and g0748 ( new_n920_, new_n272_, N76 );
not g0749 ( new_n921_, new_n920_ );
and g0750 ( new_n922_, new_n921_, keyIn_0_51 );
not g0751 ( new_n923_, new_n922_ );
or g0752 ( new_n924_, new_n921_, keyIn_0_51 );
and g0753 ( new_n925_, new_n923_, new_n924_ );
or g0754 ( new_n926_, new_n925_, new_n434_ );
or g0755 ( new_n927_, new_n919_, new_n926_ );
or g0756 ( new_n928_, new_n914_, new_n927_ );
and g0757 ( new_n929_, new_n928_, new_n880_ );
and g0758 ( new_n930_, new_n912_, new_n908_ );
and g0759 ( new_n931_, new_n906_, keyIn_0_107 );
or g0760 ( new_n932_, new_n931_, new_n930_ );
not g0761 ( new_n933_, new_n927_ );
and g0762 ( new_n934_, new_n932_, new_n933_ );
and g0763 ( new_n935_, new_n934_, keyIn_0_114 );
or g0764 ( new_n936_, new_n929_, new_n935_ );
and g0765 ( new_n937_, new_n911_, N79 );
and g0766 ( new_n938_, new_n937_, keyIn_0_106 );
not g0767 ( new_n939_, new_n938_ );
or g0768 ( new_n940_, new_n937_, keyIn_0_106 );
and g0769 ( new_n941_, new_n939_, new_n940_ );
and g0770 ( new_n942_, new_n918_, N73 );
not g0771 ( new_n943_, new_n942_ );
and g0772 ( new_n944_, new_n943_, keyIn_0_91 );
not g0773 ( new_n945_, new_n944_ );
or g0774 ( new_n946_, new_n943_, keyIn_0_91 );
and g0775 ( new_n947_, new_n945_, new_n946_ );
not g0776 ( new_n948_, new_n947_ );
and g0777 ( new_n949_, new_n272_, N63 );
not g0778 ( new_n950_, new_n949_ );
and g0779 ( new_n951_, new_n950_, keyIn_0_50 );
not g0780 ( new_n952_, new_n951_ );
or g0781 ( new_n953_, new_n950_, keyIn_0_50 );
and g0782 ( new_n954_, new_n952_, new_n953_ );
not g0783 ( new_n955_, new_n954_ );
and g0784 ( new_n956_, new_n955_, N69 );
and g0785 ( new_n957_, new_n948_, new_n956_ );
not g0786 ( new_n958_, new_n957_ );
or g0787 ( new_n959_, new_n941_, new_n958_ );
and g0788 ( new_n960_, new_n959_, keyIn_0_113 );
not g0789 ( new_n961_, new_n960_ );
or g0790 ( new_n962_, new_n959_, keyIn_0_113 );
and g0791 ( new_n963_, new_n961_, new_n962_ );
and g0792 ( new_n964_, new_n911_, N105 );
and g0793 ( new_n965_, new_n964_, keyIn_0_108 );
not g0794 ( new_n966_, new_n965_ );
or g0795 ( new_n967_, new_n964_, keyIn_0_108 );
and g0796 ( new_n968_, new_n966_, new_n967_ );
not g0797 ( new_n969_, keyIn_0_92 );
and g0798 ( new_n970_, new_n918_, N99 );
not g0799 ( new_n971_, new_n970_ );
and g0800 ( new_n972_, new_n971_, new_n969_ );
and g0801 ( new_n973_, new_n970_, keyIn_0_92 );
and g0802 ( new_n974_, new_n272_, N89 );
and g0803 ( new_n975_, new_n974_, keyIn_0_52 );
not g0804 ( new_n976_, new_n975_ );
or g0805 ( new_n977_, new_n974_, keyIn_0_52 );
and g0806 ( new_n978_, new_n976_, new_n977_ );
or g0807 ( new_n979_, new_n978_, new_n184_ );
or g0808 ( new_n980_, new_n973_, new_n979_ );
or g0809 ( new_n981_, new_n980_, new_n972_ );
or g0810 ( new_n982_, new_n968_, new_n981_ );
and g0811 ( new_n983_, new_n911_, N115 );
and g0812 ( new_n984_, new_n918_, N112 );
and g0813 ( new_n985_, new_n272_, N102 );
and g0814 ( new_n986_, new_n985_, keyIn_0_53 );
not g0815 ( new_n987_, new_n986_ );
or g0816 ( new_n988_, new_n985_, keyIn_0_53 );
and g0817 ( new_n989_, new_n987_, new_n988_ );
or g0818 ( new_n990_, new_n989_, new_n174_ );
or g0819 ( new_n991_, new_n984_, new_n990_ );
or g0820 ( new_n992_, new_n983_, new_n991_ );
and g0821 ( new_n993_, new_n982_, new_n992_ );
and g0822 ( new_n994_, new_n963_, new_n993_ );
and g0823 ( new_n995_, new_n994_, new_n936_ );
not g0824 ( new_n996_, keyIn_0_102 );
and g0825 ( new_n997_, new_n911_, N27 );
and g0826 ( new_n998_, new_n997_, new_n996_ );
not g0827 ( new_n999_, new_n998_ );
or g0828 ( new_n1000_, new_n997_, new_n996_ );
and g0829 ( new_n1001_, new_n999_, new_n1000_ );
not g0830 ( new_n1002_, keyIn_0_84 );
and g0831 ( new_n1003_, new_n918_, N21 );
and g0832 ( new_n1004_, new_n1003_, new_n1002_ );
not g0833 ( new_n1005_, new_n1004_ );
or g0834 ( new_n1006_, new_n1003_, new_n1002_ );
and g0835 ( new_n1007_, new_n272_, N11 );
or g0836 ( new_n1008_, new_n1007_, new_n288_ );
not g0837 ( new_n1009_, new_n1008_ );
and g0838 ( new_n1010_, new_n1006_, new_n1009_ );
and g0839 ( new_n1011_, new_n1010_, new_n1005_ );
not g0840 ( new_n1012_, new_n1011_ );
or g0841 ( new_n1013_, new_n1001_, new_n1012_ );
or g0842 ( new_n1014_, new_n1013_, keyIn_0_110 );
not g0843 ( new_n1015_, new_n1014_ );
and g0844 ( new_n1016_, new_n1013_, keyIn_0_110 );
or g0845 ( new_n1017_, new_n1015_, new_n1016_ );
not g0846 ( new_n1018_, keyIn_0_111 );
and g0847 ( new_n1019_, new_n911_, N40 );
not g0848 ( new_n1020_, new_n1019_ );
and g0849 ( new_n1021_, new_n1020_, keyIn_0_103 );
not g0850 ( new_n1022_, keyIn_0_103 );
and g0851 ( new_n1023_, new_n1019_, new_n1022_ );
or g0852 ( new_n1024_, new_n1021_, new_n1023_ );
and g0853 ( new_n1025_, new_n918_, N34 );
not g0854 ( new_n1026_, new_n1025_ );
not g0855 ( new_n1027_, keyIn_0_46 );
and g0856 ( new_n1028_, new_n272_, N24 );
and g0857 ( new_n1029_, new_n1028_, new_n1027_ );
not g0858 ( new_n1030_, new_n1029_ );
or g0859 ( new_n1031_, new_n1028_, new_n1027_ );
and g0860 ( new_n1032_, new_n1031_, N30 );
and g0861 ( new_n1033_, new_n1032_, new_n1030_ );
and g0862 ( new_n1034_, new_n1026_, new_n1033_ );
and g0863 ( new_n1035_, new_n1024_, new_n1034_ );
and g0864 ( new_n1036_, new_n1035_, new_n1018_ );
not g0865 ( new_n1037_, new_n1036_ );
or g0866 ( new_n1038_, new_n1035_, new_n1018_ );
and g0867 ( new_n1039_, new_n1037_, new_n1038_ );
and g0868 ( new_n1040_, new_n1017_, new_n1039_ );
not g0869 ( new_n1041_, keyIn_0_105 );
and g0870 ( new_n1042_, new_n911_, N66 );
and g0871 ( new_n1043_, new_n1042_, new_n1041_ );
or g0872 ( new_n1044_, new_n905_, new_n618_ );
and g0873 ( new_n1045_, new_n1044_, keyIn_0_105 );
and g0874 ( new_n1046_, new_n918_, N60 );
not g0875 ( new_n1047_, new_n1046_ );
and g0876 ( new_n1048_, new_n1047_, keyIn_0_89 );
not g0877 ( new_n1049_, new_n1048_ );
or g0878 ( new_n1050_, new_n1047_, keyIn_0_89 );
and g0879 ( new_n1051_, new_n1049_, new_n1050_ );
not g0880 ( new_n1052_, keyIn_0_49 );
and g0881 ( new_n1053_, new_n272_, N50 );
not g0882 ( new_n1054_, new_n1053_ );
and g0883 ( new_n1055_, new_n1054_, new_n1052_ );
and g0884 ( new_n1056_, new_n1053_, keyIn_0_49 );
or g0885 ( new_n1057_, new_n1056_, new_n202_ );
or g0886 ( new_n1058_, new_n1057_, new_n1055_ );
or g0887 ( new_n1059_, new_n1051_, new_n1058_ );
or g0888 ( new_n1060_, new_n1045_, new_n1059_ );
or g0889 ( new_n1061_, new_n1060_, new_n1043_ );
and g0890 ( new_n1062_, new_n1061_, keyIn_0_112 );
not g0891 ( new_n1063_, keyIn_0_112 );
not g0892 ( new_n1064_, new_n1043_ );
or g0893 ( new_n1065_, new_n1042_, new_n1041_ );
not g0894 ( new_n1066_, new_n1059_ );
and g0895 ( new_n1067_, new_n1065_, new_n1066_ );
and g0896 ( new_n1068_, new_n1067_, new_n1064_ );
and g0897 ( new_n1069_, new_n1068_, new_n1063_ );
or g0898 ( new_n1070_, new_n1062_, new_n1069_ );
and g0899 ( new_n1071_, new_n911_, N53 );
and g0900 ( new_n1072_, new_n1071_, keyIn_0_104 );
not g0901 ( new_n1073_, new_n1072_ );
or g0902 ( new_n1074_, new_n1071_, keyIn_0_104 );
and g0903 ( new_n1075_, new_n1073_, new_n1074_ );
not g0904 ( new_n1076_, keyIn_0_87 );
and g0905 ( new_n1077_, new_n918_, N47 );
not g0906 ( new_n1078_, new_n1077_ );
and g0907 ( new_n1079_, new_n1078_, new_n1076_ );
not g0908 ( new_n1080_, new_n1079_ );
and g0909 ( new_n1081_, new_n1077_, keyIn_0_87 );
not g0910 ( new_n1082_, new_n1081_ );
not g0911 ( new_n1083_, keyIn_0_48 );
and g0912 ( new_n1084_, new_n272_, N37 );
and g0913 ( new_n1085_, new_n1084_, new_n1083_ );
not g0914 ( new_n1086_, new_n1085_ );
or g0915 ( new_n1087_, new_n1084_, new_n1083_ );
and g0916 ( new_n1088_, new_n1087_, N43 );
and g0917 ( new_n1089_, new_n1088_, new_n1086_ );
and g0918 ( new_n1090_, new_n1082_, new_n1089_ );
and g0919 ( new_n1091_, new_n1090_, new_n1080_ );
not g0920 ( new_n1092_, new_n1091_ );
or g0921 ( new_n1093_, new_n1075_, new_n1092_ );
and g0922 ( new_n1094_, new_n1070_, new_n1093_ );
and g0923 ( new_n1095_, new_n1040_, new_n1094_ );
and g0924 ( new_n1096_, new_n1095_, new_n995_ );
or g0925 ( new_n1097_, new_n1096_, new_n879_ );
not g0926 ( new_n1098_, new_n1097_ );
and g0927 ( new_n1099_, new_n1096_, new_n879_ );
or g0928 ( new_n1100_, new_n1098_, new_n1099_ );
not g0929 ( new_n1101_, keyIn_0_101 );
and g0930 ( new_n1102_, new_n911_, N14 );
not g0931 ( new_n1103_, new_n1102_ );
and g0932 ( new_n1104_, new_n1103_, new_n1101_ );
and g0933 ( new_n1105_, new_n1102_, keyIn_0_101 );
and g0934 ( new_n1106_, new_n918_, N8 );
not g0935 ( new_n1107_, keyIn_0_44 );
and g0936 ( new_n1108_, new_n272_, N1 );
not g0937 ( new_n1109_, new_n1108_ );
and g0938 ( new_n1110_, new_n1109_, new_n1107_ );
and g0939 ( new_n1111_, new_n1108_, keyIn_0_44 );
or g0940 ( new_n1112_, new_n1111_, new_n212_ );
or g0941 ( new_n1113_, new_n1112_, new_n1110_ );
or g0942 ( new_n1114_, new_n1106_, new_n1113_ );
or g0943 ( new_n1115_, new_n1105_, new_n1114_ );
or g0944 ( new_n1116_, new_n1115_, new_n1104_ );
not g0945 ( new_n1117_, new_n1116_ );
and g0946 ( new_n1118_, new_n1117_, keyIn_0_109 );
not g0947 ( new_n1119_, new_n1118_ );
or g0948 ( new_n1120_, new_n1117_, keyIn_0_109 );
and g0949 ( new_n1121_, new_n1119_, new_n1120_ );
and g0950 ( new_n1122_, new_n1100_, new_n1121_ );
or g0951 ( new_n1123_, new_n1122_, keyIn_0_120 );
not g0952 ( new_n1124_, keyIn_0_120 );
not g0953 ( new_n1125_, new_n1099_ );
and g0954 ( new_n1126_, new_n1125_, new_n1097_ );
not g0955 ( new_n1127_, new_n1121_ );
or g0956 ( new_n1128_, new_n1126_, new_n1127_ );
or g0957 ( new_n1129_, new_n1128_, new_n1124_ );
and g0958 ( N421, new_n1123_, new_n1129_ );
not g0959 ( new_n1131_, keyIn_0_125 );
and g0960 ( new_n1132_, new_n1093_, keyIn_0_116 );
not g0961 ( new_n1133_, new_n1132_ );
or g0962 ( new_n1134_, new_n1093_, keyIn_0_116 );
and g0963 ( new_n1135_, new_n1133_, new_n1134_ );
and g0964 ( new_n1136_, new_n1039_, new_n1135_ );
and g0965 ( new_n1137_, new_n1136_, keyIn_0_121 );
not g0966 ( new_n1138_, new_n1137_ );
or g0967 ( new_n1139_, new_n1136_, keyIn_0_121 );
and g0968 ( new_n1140_, new_n1138_, new_n1139_ );
and g0969 ( new_n1141_, new_n1040_, new_n1070_ );
and g0970 ( new_n1142_, new_n1140_, new_n1141_ );
not g0971 ( new_n1143_, new_n1142_ );
and g0972 ( new_n1144_, new_n1143_, new_n1131_ );
and g0973 ( new_n1145_, new_n1142_, keyIn_0_125 );
or g0974 ( N430, new_n1144_, new_n1145_ );
not g0975 ( new_n1147_, keyIn_0_117 );
not g0976 ( new_n1148_, new_n962_ );
or g0977 ( new_n1149_, new_n1148_, new_n960_ );
or g0978 ( new_n1150_, new_n1149_, new_n1147_ );
or g0979 ( new_n1151_, new_n963_, keyIn_0_117 );
and g0980 ( new_n1152_, new_n1150_, new_n1151_ );
and g0981 ( new_n1153_, new_n1039_, new_n1093_ );
and g0982 ( new_n1154_, new_n1153_, new_n1070_ );
not g0983 ( new_n1155_, new_n1154_ );
or g0984 ( new_n1156_, new_n1155_, new_n1152_ );
and g0985 ( new_n1157_, new_n1156_, keyIn_0_122 );
not g0986 ( new_n1158_, keyIn_0_122 );
and g0987 ( new_n1159_, new_n963_, keyIn_0_117 );
and g0988 ( new_n1160_, new_n1149_, new_n1147_ );
or g0989 ( new_n1161_, new_n1160_, new_n1159_ );
and g0990 ( new_n1162_, new_n1161_, new_n1154_ );
and g0991 ( new_n1163_, new_n1162_, new_n1158_ );
or g0992 ( new_n1164_, new_n1157_, new_n1163_ );
not g0993 ( new_n1165_, new_n1016_ );
and g0994 ( new_n1166_, new_n1165_, new_n1014_ );
not g0995 ( new_n1167_, new_n1038_ );
or g0996 ( new_n1168_, new_n1167_, new_n1036_ );
or g0997 ( new_n1169_, new_n1168_, new_n1166_ );
not g0998 ( new_n1170_, keyIn_0_123 );
not g0999 ( new_n1171_, keyIn_0_118 );
and g1000 ( new_n1172_, new_n936_, new_n1171_ );
or g1001 ( new_n1173_, new_n1068_, new_n1063_ );
or g1002 ( new_n1174_, new_n1061_, keyIn_0_112 );
and g1003 ( new_n1175_, new_n1174_, new_n1173_ );
not g1004 ( new_n1176_, new_n1093_ );
or g1005 ( new_n1177_, new_n1175_, new_n1176_ );
or g1006 ( new_n1178_, new_n934_, keyIn_0_114 );
or g1007 ( new_n1179_, new_n928_, new_n880_ );
and g1008 ( new_n1180_, new_n1179_, new_n1178_ );
and g1009 ( new_n1181_, new_n1180_, keyIn_0_118 );
or g1010 ( new_n1182_, new_n1177_, new_n1181_ );
or g1011 ( new_n1183_, new_n1182_, new_n1172_ );
or g1012 ( new_n1184_, new_n1183_, new_n1170_ );
not g1013 ( new_n1185_, new_n1172_ );
or g1014 ( new_n1186_, new_n936_, new_n1171_ );
and g1015 ( new_n1187_, new_n1186_, new_n1094_ );
and g1016 ( new_n1188_, new_n1187_, new_n1185_ );
or g1017 ( new_n1189_, new_n1188_, keyIn_0_123 );
and g1018 ( new_n1190_, new_n1184_, new_n1189_ );
or g1019 ( new_n1191_, new_n1190_, new_n1169_ );
or g1020 ( new_n1192_, new_n1191_, new_n1164_ );
and g1021 ( new_n1193_, new_n1192_, keyIn_0_126 );
not g1022 ( new_n1194_, keyIn_0_126 );
or g1023 ( new_n1195_, new_n1162_, new_n1158_ );
not g1024 ( new_n1196_, new_n1163_ );
and g1025 ( new_n1197_, new_n1196_, new_n1195_ );
and g1026 ( new_n1198_, new_n1188_, keyIn_0_123 );
and g1027 ( new_n1199_, new_n1183_, new_n1170_ );
or g1028 ( new_n1200_, new_n1199_, new_n1198_ );
and g1029 ( new_n1201_, new_n1200_, new_n1040_ );
and g1030 ( new_n1202_, new_n1197_, new_n1201_ );
and g1031 ( new_n1203_, new_n1202_, new_n1194_ );
or g1032 ( N431, new_n1193_, new_n1203_ );
and g1033 ( new_n1205_, new_n982_, keyIn_0_119 );
not g1034 ( new_n1206_, new_n1205_ );
or g1035 ( new_n1207_, new_n982_, keyIn_0_119 );
and g1036 ( new_n1208_, new_n1206_, new_n1207_ );
and g1037 ( new_n1209_, new_n1208_, new_n936_ );
and g1038 ( new_n1210_, new_n1209_, new_n1153_ );
and g1039 ( new_n1211_, new_n1210_, keyIn_0_124 );
not g1040 ( new_n1212_, new_n1211_ );
or g1041 ( new_n1213_, new_n1210_, keyIn_0_124 );
and g1042 ( new_n1214_, new_n1212_, new_n1213_ );
not g1043 ( new_n1215_, keyIn_0_121 );
not g1044 ( new_n1216_, keyIn_0_116 );
and g1045 ( new_n1217_, new_n1176_, new_n1216_ );
or g1046 ( new_n1218_, new_n1217_, new_n1132_ );
or g1047 ( new_n1219_, new_n1168_, new_n1218_ );
and g1048 ( new_n1220_, new_n1219_, new_n1215_ );
or g1049 ( new_n1221_, new_n1220_, new_n1137_ );
or g1050 ( new_n1222_, new_n1221_, new_n1166_ );
or g1051 ( new_n1223_, new_n1222_, new_n1214_ );
or g1052 ( new_n1224_, new_n1223_, new_n1164_ );
and g1053 ( new_n1225_, new_n1224_, keyIn_0_127 );
not g1054 ( new_n1226_, keyIn_0_127 );
not g1055 ( new_n1227_, new_n1213_ );
or g1056 ( new_n1228_, new_n1227_, new_n1211_ );
and g1057 ( new_n1229_, new_n1140_, new_n1017_ );
and g1058 ( new_n1230_, new_n1228_, new_n1229_ );
and g1059 ( new_n1231_, new_n1197_, new_n1230_ );
and g1060 ( new_n1232_, new_n1231_, new_n1226_ );
or g1061 ( N432, new_n1225_, new_n1232_ );
endmodule