module add_mul_combine_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, Result_mul_0_, Result_mul_1_, 
        Result_mul_2_, Result_mul_3_, Result_mul_4_, Result_mul_5_, 
        Result_mul_6_, Result_mul_7_, Result_mul_8_, Result_mul_9_, 
        Result_mul_10_, Result_mul_11_, Result_mul_12_, Result_mul_13_, 
        Result_mul_14_, Result_mul_15_, Result_mul_16_, Result_mul_17_, 
        Result_mul_18_, Result_mul_19_, Result_mul_20_, Result_mul_21_, 
        Result_mul_22_, Result_mul_23_, Result_mul_24_, Result_mul_25_, 
        Result_mul_26_, Result_mul_27_, Result_mul_28_, Result_mul_29_, 
        Result_mul_30_, Result_mul_31_, Result_mul_32_, Result_mul_33_, 
        Result_mul_34_, Result_mul_35_, Result_mul_36_, Result_mul_37_, 
        Result_mul_38_, Result_mul_39_, Result_mul_40_, Result_mul_41_, 
        Result_mul_42_, Result_mul_43_, Result_mul_44_, Result_mul_45_, 
        Result_mul_46_, Result_mul_47_, Result_mul_48_, Result_mul_49_, 
        Result_mul_50_, Result_mul_51_, Result_mul_52_, Result_mul_53_, 
        Result_mul_54_, Result_mul_55_, Result_mul_56_, Result_mul_57_, 
        Result_mul_58_, Result_mul_59_, Result_mul_60_, Result_mul_61_, 
        Result_mul_62_, Result_mul_63_, Result_add_0_, Result_add_1_, 
        Result_add_2_, Result_add_3_, Result_add_4_, Result_add_5_, 
        Result_add_6_, Result_add_7_, Result_add_8_, Result_add_9_, 
        Result_add_10_, Result_add_11_, Result_add_12_, Result_add_13_, 
        Result_add_14_, Result_add_15_, Result_add_16_, Result_add_17_, 
        Result_add_18_, Result_add_19_, Result_add_20_, Result_add_21_, 
        Result_add_22_, Result_add_23_, Result_add_24_, Result_add_25_, 
        Result_add_26_, Result_add_27_, Result_add_28_, Result_add_29_, 
        Result_add_30_, Result_add_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_mul_32_, Result_mul_33_, Result_mul_34_, Result_mul_35_,
         Result_mul_36_, Result_mul_37_, Result_mul_38_, Result_mul_39_,
         Result_mul_40_, Result_mul_41_, Result_mul_42_, Result_mul_43_,
         Result_mul_44_, Result_mul_45_, Result_mul_46_, Result_mul_47_,
         Result_mul_48_, Result_mul_49_, Result_mul_50_, Result_mul_51_,
         Result_mul_52_, Result_mul_53_, Result_mul_54_, Result_mul_55_,
         Result_mul_56_, Result_mul_57_, Result_mul_58_, Result_mul_59_,
         Result_mul_60_, Result_mul_61_, Result_mul_62_, Result_mul_63_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_,
         Result_add_16_, Result_add_17_, Result_add_18_, Result_add_19_,
         Result_add_20_, Result_add_21_, Result_add_22_, Result_add_23_,
         Result_add_24_, Result_add_25_, Result_add_26_, Result_add_27_,
         Result_add_28_, Result_add_29_, Result_add_30_, Result_add_31_;
  wire   n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651;

  INV_X2 U8433 ( .A(b_10_), .ZN(n13725) );
  INV_X2 U8434 ( .A(b_2_), .ZN(n15690) );
  INV_X2 U8435 ( .A(b_8_), .ZN(n14216) );
  INV_X2 U8436 ( .A(b_3_), .ZN(n15446) );
  INV_X2 U8437 ( .A(b_0_), .ZN(n16206) );
  INV_X2 U8438 ( .A(n16207), .ZN(n8362) );
  INV_X2 U8439 ( .A(a_4_), .ZN(n8712) );
  INV_X2 U8440 ( .A(a_1_), .ZN(n8502) );
  INV_X2 U8441 ( .A(a_2_), .ZN(n8497) );
  INV_X2 U8442 ( .A(a_0_), .ZN(n8690) );
  INV_X2 U8443 ( .A(a_20_), .ZN(n10633) );
  INV_X2 U8444 ( .A(a_12_), .ZN(n8750) );
  INV_X2 U8445 ( .A(a_6_), .ZN(n8480) );
  INV_X2 U8446 ( .A(a_27_), .ZN(n8839) );
  INV_X2 U8447 ( .A(a_5_), .ZN(n8717) );
  INV_X2 U8448 ( .A(a_9_), .ZN(n8736) );
  NAND2_X2 U8449 ( .A1(a_31_), .A2(n16203), .ZN(n8358) );
  INV_X2 U8450 ( .A(a_26_), .ZN(n8830) );
  INV_X2 U8451 ( .A(b_4_), .ZN(n15197) );
  INV_X2 U8452 ( .A(a_24_), .ZN(n9131) );
  INV_X2 U8453 ( .A(a_28_), .ZN(n8844) );
  INV_X2 U8454 ( .A(a_29_), .ZN(n9161) );
  INV_X2 U8455 ( .A(a_25_), .ZN(n8825) );
  INV_X2 U8456 ( .A(a_11_), .ZN(n8452) );
  INV_X2 U8457 ( .A(b_1_), .ZN(n15994) );
  INV_X2 U8458 ( .A(a_15_), .ZN(n8763) );
  INV_X2 U8459 ( .A(a_19_), .ZN(n8881) );
  INV_X2 U8460 ( .A(b_11_), .ZN(n13436) );
  INV_X2 U8461 ( .A(b_7_), .ZN(n14438) );
  INV_X2 U8462 ( .A(a_23_), .ZN(n8812) );
  INV_X2 U8463 ( .A(b_5_), .ZN(n14947) );
  INV_X2 U8464 ( .A(b_9_), .ZN(n13926) );
  XOR2_X1 U8465 ( .A(n8337), .B(n8338), .Z(Result_mul_9_) );
  NOR2_X1 U8466 ( .A1(n8339), .A2(n8340), .ZN(n8338) );
  INV_X1 U8467 ( .A(n8341), .ZN(n8340) );
  NOR2_X1 U8468 ( .A1(n8342), .A2(n8343), .ZN(n8339) );
  XOR2_X1 U8469 ( .A(n8344), .B(n8345), .Z(Result_mul_8_) );
  XOR2_X1 U8470 ( .A(n8346), .B(n8347), .Z(Result_mul_7_) );
  NOR2_X1 U8471 ( .A1(n8348), .A2(n8349), .ZN(n8347) );
  INV_X1 U8472 ( .A(n8350), .ZN(n8349) );
  NOR2_X1 U8473 ( .A1(n8351), .A2(n8352), .ZN(n8348) );
  XOR2_X1 U8474 ( .A(n8353), .B(n8354), .Z(Result_mul_6_) );
  NAND2_X1 U8475 ( .A1(n8355), .A2(n8356), .ZN(Result_mul_62_) );
  NAND2_X1 U8476 ( .A1(b_30_), .A2(n8357), .ZN(n8356) );
  NAND2_X1 U8477 ( .A1(n8358), .A2(n8359), .ZN(n8357) );
  NAND2_X1 U8478 ( .A1(a_31_), .A2(n8360), .ZN(n8359) );
  NAND2_X1 U8479 ( .A1(b_31_), .A2(n8361), .ZN(n8355) );
  NAND2_X1 U8480 ( .A1(n8362), .A2(n8363), .ZN(n8361) );
  NAND2_X1 U8481 ( .A1(a_30_), .A2(n8364), .ZN(n8363) );
  XNOR2_X1 U8482 ( .A(n8365), .B(n8366), .ZN(Result_mul_61_) );
  XOR2_X1 U8483 ( .A(n8367), .B(n8368), .Z(n8366) );
  XOR2_X1 U8484 ( .A(n8369), .B(n8370), .Z(Result_mul_60_) );
  XOR2_X1 U8485 ( .A(n8371), .B(n8372), .Z(n8369) );
  XOR2_X1 U8486 ( .A(n8373), .B(n8374), .Z(Result_mul_5_) );
  NOR2_X1 U8487 ( .A1(n8375), .A2(n8376), .ZN(n8374) );
  INV_X1 U8488 ( .A(n8377), .ZN(n8376) );
  NOR2_X1 U8489 ( .A1(n8378), .A2(n8379), .ZN(n8375) );
  XNOR2_X1 U8490 ( .A(n8380), .B(n8381), .ZN(Result_mul_59_) );
  NAND2_X1 U8491 ( .A1(n8382), .A2(n8383), .ZN(n8380) );
  XOR2_X1 U8492 ( .A(n8384), .B(n8385), .Z(Result_mul_58_) );
  XOR2_X1 U8493 ( .A(n8386), .B(n8387), .Z(n8385) );
  XOR2_X1 U8494 ( .A(n8388), .B(n8389), .Z(Result_mul_57_) );
  XOR2_X1 U8495 ( .A(n8390), .B(n8391), .Z(n8389) );
  XOR2_X1 U8496 ( .A(n8392), .B(n8393), .Z(Result_mul_56_) );
  XNOR2_X1 U8497 ( .A(n8394), .B(n8395), .ZN(n8393) );
  XNOR2_X1 U8498 ( .A(n8396), .B(n8397), .ZN(Result_mul_55_) );
  NAND2_X1 U8499 ( .A1(n8398), .A2(n8399), .ZN(n8396) );
  XNOR2_X1 U8500 ( .A(n8400), .B(n8401), .ZN(Result_mul_54_) );
  XNOR2_X1 U8501 ( .A(n8402), .B(n8403), .ZN(n8401) );
  XOR2_X1 U8502 ( .A(n8404), .B(n8405), .Z(Result_mul_53_) );
  XOR2_X1 U8503 ( .A(n8406), .B(n8407), .Z(n8405) );
  XNOR2_X1 U8504 ( .A(n8408), .B(n8409), .ZN(Result_mul_52_) );
  XOR2_X1 U8505 ( .A(n8410), .B(n8411), .Z(n8409) );
  XOR2_X1 U8506 ( .A(n8412), .B(n8413), .Z(Result_mul_51_) );
  XOR2_X1 U8507 ( .A(n8414), .B(n8415), .Z(n8413) );
  XNOR2_X1 U8508 ( .A(n8416), .B(n8417), .ZN(Result_mul_50_) );
  XOR2_X1 U8509 ( .A(n8418), .B(n8419), .Z(n8417) );
  XOR2_X1 U8510 ( .A(n8420), .B(n8421), .Z(Result_mul_4_) );
  XOR2_X1 U8511 ( .A(n8422), .B(n8423), .Z(Result_mul_49_) );
  XOR2_X1 U8512 ( .A(n8424), .B(n8425), .Z(n8423) );
  XOR2_X1 U8513 ( .A(n8426), .B(n8427), .Z(Result_mul_48_) );
  XNOR2_X1 U8514 ( .A(n8428), .B(n8429), .ZN(n8426) );
  NAND2_X1 U8515 ( .A1(b_31_), .A2(a_16_), .ZN(n8428) );
  XNOR2_X1 U8516 ( .A(n8430), .B(n8431), .ZN(Result_mul_47_) );
  XOR2_X1 U8517 ( .A(n8432), .B(n8433), .Z(n8431) );
  NAND2_X1 U8518 ( .A1(b_31_), .A2(a_15_), .ZN(n8433) );
  XOR2_X1 U8519 ( .A(n8434), .B(n8435), .Z(Result_mul_46_) );
  XOR2_X1 U8520 ( .A(n8436), .B(n8437), .Z(n8434) );
  NOR2_X1 U8521 ( .A1(n8438), .A2(n8360), .ZN(n8437) );
  XOR2_X1 U8522 ( .A(n8439), .B(n8440), .Z(Result_mul_45_) );
  XOR2_X1 U8523 ( .A(n8441), .B(n8442), .Z(n8439) );
  NOR2_X1 U8524 ( .A1(n8443), .A2(n8360), .ZN(n8442) );
  XNOR2_X1 U8525 ( .A(n8444), .B(n8445), .ZN(Result_mul_44_) );
  XOR2_X1 U8526 ( .A(n8446), .B(n8447), .Z(n8445) );
  NAND2_X1 U8527 ( .A1(b_31_), .A2(a_12_), .ZN(n8447) );
  XOR2_X1 U8528 ( .A(n8448), .B(n8449), .Z(Result_mul_43_) );
  XOR2_X1 U8529 ( .A(n8450), .B(n8451), .Z(n8448) );
  NOR2_X1 U8530 ( .A1(n8452), .A2(n8360), .ZN(n8451) );
  XNOR2_X1 U8531 ( .A(n8453), .B(n8454), .ZN(Result_mul_42_) );
  XOR2_X1 U8532 ( .A(n8455), .B(n8456), .Z(n8454) );
  NAND2_X1 U8533 ( .A1(b_31_), .A2(a_10_), .ZN(n8456) );
  XNOR2_X1 U8534 ( .A(n8457), .B(n8458), .ZN(Result_mul_41_) );
  XOR2_X1 U8535 ( .A(n8459), .B(n8460), .Z(n8458) );
  NAND2_X1 U8536 ( .A1(b_31_), .A2(a_9_), .ZN(n8460) );
  XNOR2_X1 U8537 ( .A(n8461), .B(n8462), .ZN(Result_mul_40_) );
  XOR2_X1 U8538 ( .A(n8463), .B(n8464), .Z(n8462) );
  NAND2_X1 U8539 ( .A1(b_31_), .A2(a_8_), .ZN(n8464) );
  XOR2_X1 U8540 ( .A(n8465), .B(n8466), .Z(Result_mul_3_) );
  NOR2_X1 U8541 ( .A1(n8467), .A2(n8468), .ZN(n8466) );
  INV_X1 U8542 ( .A(n8469), .ZN(n8468) );
  NOR2_X1 U8543 ( .A1(n8470), .A2(n8471), .ZN(n8467) );
  XNOR2_X1 U8544 ( .A(n8472), .B(n8473), .ZN(Result_mul_39_) );
  XOR2_X1 U8545 ( .A(n8474), .B(n8475), .Z(n8473) );
  NAND2_X1 U8546 ( .A1(b_31_), .A2(a_7_), .ZN(n8475) );
  XOR2_X1 U8547 ( .A(n8476), .B(n8477), .Z(Result_mul_38_) );
  XOR2_X1 U8548 ( .A(n8478), .B(n8479), .Z(n8476) );
  NOR2_X1 U8549 ( .A1(n8480), .A2(n8360), .ZN(n8479) );
  XNOR2_X1 U8550 ( .A(n8481), .B(n8482), .ZN(Result_mul_37_) );
  XOR2_X1 U8551 ( .A(n8483), .B(n8484), .Z(n8482) );
  NAND2_X1 U8552 ( .A1(b_31_), .A2(a_5_), .ZN(n8484) );
  XNOR2_X1 U8553 ( .A(n8485), .B(n8486), .ZN(Result_mul_36_) );
  XOR2_X1 U8554 ( .A(n8487), .B(n8488), .Z(n8486) );
  NAND2_X1 U8555 ( .A1(b_31_), .A2(a_4_), .ZN(n8488) );
  XNOR2_X1 U8556 ( .A(n8489), .B(n8490), .ZN(Result_mul_35_) );
  XOR2_X1 U8557 ( .A(n8491), .B(n8492), .Z(n8490) );
  NAND2_X1 U8558 ( .A1(b_31_), .A2(a_3_), .ZN(n8492) );
  XOR2_X1 U8559 ( .A(n8493), .B(n8494), .Z(Result_mul_34_) );
  XOR2_X1 U8560 ( .A(n8495), .B(n8496), .Z(n8493) );
  NOR2_X1 U8561 ( .A1(n8497), .A2(n8360), .ZN(n8496) );
  XOR2_X1 U8562 ( .A(n8498), .B(n8499), .Z(Result_mul_33_) );
  XOR2_X1 U8563 ( .A(n8500), .B(n8501), .Z(n8498) );
  NOR2_X1 U8564 ( .A1(n8502), .A2(n8360), .ZN(n8501) );
  XNOR2_X1 U8565 ( .A(n8503), .B(n8504), .ZN(Result_mul_32_) );
  XOR2_X1 U8566 ( .A(n8505), .B(n8506), .Z(n8504) );
  NAND2_X1 U8567 ( .A1(b_31_), .A2(a_0_), .ZN(n8506) );
  XOR2_X1 U8568 ( .A(n8507), .B(n8508), .Z(Result_mul_31_) );
  NOR2_X1 U8569 ( .A1(n8509), .A2(n8510), .ZN(Result_mul_30_) );
  NOR2_X1 U8570 ( .A1(n8511), .A2(n8512), .ZN(n8510) );
  NOR2_X1 U8571 ( .A1(n8507), .A2(n8508), .ZN(n8511) );
  INV_X1 U8572 ( .A(n8513), .ZN(n8507) );
  XOR2_X1 U8573 ( .A(n8514), .B(n8515), .Z(Result_mul_2_) );
  XNOR2_X1 U8574 ( .A(n8509), .B(n8516), .ZN(Result_mul_29_) );
  NAND2_X1 U8575 ( .A1(n8517), .A2(n8518), .ZN(n8516) );
  XNOR2_X1 U8576 ( .A(n8519), .B(n8520), .ZN(Result_mul_28_) );
  NAND2_X1 U8577 ( .A1(n8521), .A2(n8522), .ZN(n8519) );
  XNOR2_X1 U8578 ( .A(n8523), .B(n8524), .ZN(Result_mul_27_) );
  NAND2_X1 U8579 ( .A1(n8525), .A2(n8526), .ZN(n8524) );
  XNOR2_X1 U8580 ( .A(n8527), .B(n8528), .ZN(Result_mul_26_) );
  NAND2_X1 U8581 ( .A1(n8529), .A2(n8530), .ZN(n8528) );
  XOR2_X1 U8582 ( .A(n8531), .B(n8532), .Z(Result_mul_25_) );
  NOR2_X1 U8583 ( .A1(n8533), .A2(n8534), .ZN(n8532) );
  NOR2_X1 U8584 ( .A1(n8535), .A2(n8536), .ZN(n8534) );
  INV_X1 U8585 ( .A(n8537), .ZN(n8533) );
  XNOR2_X1 U8586 ( .A(n8538), .B(n8539), .ZN(Result_mul_24_) );
  NAND2_X1 U8587 ( .A1(n8540), .A2(n8541), .ZN(n8539) );
  XNOR2_X1 U8588 ( .A(n8542), .B(n8543), .ZN(Result_mul_23_) );
  NAND2_X1 U8589 ( .A1(n8544), .A2(n8545), .ZN(n8543) );
  XNOR2_X1 U8590 ( .A(n8546), .B(n8547), .ZN(Result_mul_22_) );
  NAND2_X1 U8591 ( .A1(n8548), .A2(n8549), .ZN(n8547) );
  XNOR2_X1 U8592 ( .A(n8550), .B(n8551), .ZN(Result_mul_21_) );
  NAND2_X1 U8593 ( .A1(n8552), .A2(n8553), .ZN(n8551) );
  XNOR2_X1 U8594 ( .A(n8554), .B(n8555), .ZN(Result_mul_20_) );
  NAND2_X1 U8595 ( .A1(n8556), .A2(n8557), .ZN(n8555) );
  XOR2_X1 U8596 ( .A(n8558), .B(n8559), .Z(Result_mul_1_) );
  NOR2_X1 U8597 ( .A1(n8560), .A2(n8561), .ZN(n8559) );
  XNOR2_X1 U8598 ( .A(n8562), .B(n8563), .ZN(Result_mul_19_) );
  NAND2_X1 U8599 ( .A1(n8564), .A2(n8565), .ZN(n8563) );
  XNOR2_X1 U8600 ( .A(n8566), .B(n8567), .ZN(Result_mul_18_) );
  NAND2_X1 U8601 ( .A1(n8568), .A2(n8569), .ZN(n8567) );
  XOR2_X1 U8602 ( .A(n8570), .B(n8571), .Z(Result_mul_17_) );
  NOR2_X1 U8603 ( .A1(n8572), .A2(n8573), .ZN(n8571) );
  INV_X1 U8604 ( .A(n8574), .ZN(n8573) );
  NOR2_X1 U8605 ( .A1(n8575), .A2(n8576), .ZN(n8572) );
  XOR2_X1 U8606 ( .A(n8577), .B(n8578), .Z(Result_mul_16_) );
  NOR2_X1 U8607 ( .A1(n8579), .A2(n8580), .ZN(n8578) );
  INV_X1 U8608 ( .A(n8581), .ZN(n8579) );
  XNOR2_X1 U8609 ( .A(n8582), .B(n8583), .ZN(Result_mul_15_) );
  XOR2_X1 U8610 ( .A(n8584), .B(n8585), .Z(n8583) );
  XOR2_X1 U8611 ( .A(n8586), .B(n8587), .Z(Result_mul_14_) );
  XOR2_X1 U8612 ( .A(n8588), .B(n8589), .Z(Result_mul_13_) );
  NOR2_X1 U8613 ( .A1(n8590), .A2(n8591), .ZN(n8589) );
  INV_X1 U8614 ( .A(n8592), .ZN(n8591) );
  NOR2_X1 U8615 ( .A1(n8593), .A2(n8594), .ZN(n8590) );
  XOR2_X1 U8616 ( .A(n8595), .B(n8596), .Z(Result_mul_12_) );
  XOR2_X1 U8617 ( .A(n8597), .B(n8598), .Z(Result_mul_11_) );
  NOR2_X1 U8618 ( .A1(n8599), .A2(n8600), .ZN(n8598) );
  INV_X1 U8619 ( .A(n8601), .ZN(n8600) );
  NOR2_X1 U8620 ( .A1(n8602), .A2(n8603), .ZN(n8599) );
  XOR2_X1 U8621 ( .A(n8604), .B(n8605), .Z(Result_mul_10_) );
  NAND2_X1 U8622 ( .A1(n8606), .A2(n8607), .ZN(Result_mul_0_) );
  NAND2_X1 U8623 ( .A1(a_0_), .A2(n8608), .ZN(n8607) );
  NOR2_X1 U8624 ( .A1(n8561), .A2(n8609), .ZN(n8606) );
  NOR2_X1 U8625 ( .A1(n8560), .A2(n8610), .ZN(n8609) );
  INV_X1 U8626 ( .A(n8558), .ZN(n8610) );
  NOR2_X1 U8627 ( .A1(n8514), .A2(n8515), .ZN(n8558) );
  NOR2_X1 U8628 ( .A1(n8611), .A2(n8612), .ZN(n8515) );
  NAND2_X1 U8629 ( .A1(n8469), .A2(n8613), .ZN(n8611) );
  NAND2_X1 U8630 ( .A1(n8465), .A2(n8470), .ZN(n8613) );
  NOR2_X1 U8631 ( .A1(n8421), .A2(n8420), .ZN(n8465) );
  NOR2_X1 U8632 ( .A1(n8614), .A2(n8615), .ZN(n8420) );
  NAND2_X1 U8633 ( .A1(n8377), .A2(n8616), .ZN(n8614) );
  NAND2_X1 U8634 ( .A1(n8373), .A2(n8378), .ZN(n8616) );
  NOR2_X1 U8635 ( .A1(n8354), .A2(n8353), .ZN(n8373) );
  NOR2_X1 U8636 ( .A1(n8617), .A2(n8618), .ZN(n8353) );
  NAND2_X1 U8637 ( .A1(n8350), .A2(n8619), .ZN(n8617) );
  NAND2_X1 U8638 ( .A1(n8346), .A2(n8351), .ZN(n8619) );
  NOR2_X1 U8639 ( .A1(n8345), .A2(n8344), .ZN(n8346) );
  NOR2_X1 U8640 ( .A1(n8620), .A2(n8621), .ZN(n8344) );
  NAND2_X1 U8641 ( .A1(n8341), .A2(n8622), .ZN(n8620) );
  NAND2_X1 U8642 ( .A1(n8337), .A2(n8342), .ZN(n8622) );
  NOR2_X1 U8643 ( .A1(n8605), .A2(n8604), .ZN(n8337) );
  NOR2_X1 U8644 ( .A1(n8623), .A2(n8624), .ZN(n8604) );
  NAND2_X1 U8645 ( .A1(n8601), .A2(n8625), .ZN(n8624) );
  NAND2_X1 U8646 ( .A1(n8602), .A2(n8597), .ZN(n8625) );
  NOR2_X1 U8647 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  NOR2_X1 U8648 ( .A1(n8626), .A2(n8627), .ZN(n8595) );
  NAND2_X1 U8649 ( .A1(n8592), .A2(n8628), .ZN(n8627) );
  NAND2_X1 U8650 ( .A1(n8593), .A2(n8588), .ZN(n8628) );
  NOR2_X1 U8651 ( .A1(n8586), .A2(n8587), .ZN(n8588) );
  NOR2_X1 U8652 ( .A1(n8629), .A2(n8630), .ZN(n8587) );
  NOR2_X1 U8653 ( .A1(n8584), .A2(n8631), .ZN(n8630) );
  INV_X1 U8654 ( .A(n8632), .ZN(n8631) );
  NAND2_X1 U8655 ( .A1(n8582), .A2(n8585), .ZN(n8632) );
  NOR2_X1 U8656 ( .A1(n8580), .A2(n8633), .ZN(n8582) );
  INV_X1 U8657 ( .A(n8634), .ZN(n8633) );
  NAND2_X1 U8658 ( .A1(n8581), .A2(n8577), .ZN(n8634) );
  NAND2_X1 U8659 ( .A1(n8574), .A2(n8635), .ZN(n8577) );
  NAND2_X1 U8660 ( .A1(n8575), .A2(n8570), .ZN(n8635) );
  NAND2_X1 U8661 ( .A1(n8636), .A2(n8568), .ZN(n8570) );
  NAND2_X1 U8662 ( .A1(n8637), .A2(n8638), .ZN(n8568) );
  NAND2_X1 U8663 ( .A1(n8566), .A2(n8569), .ZN(n8636) );
  INV_X1 U8664 ( .A(n8639), .ZN(n8569) );
  NOR2_X1 U8665 ( .A1(n8637), .A2(n8638), .ZN(n8639) );
  XOR2_X1 U8666 ( .A(n8640), .B(n8641), .Z(n8637) );
  NAND2_X1 U8667 ( .A1(n8565), .A2(n8642), .ZN(n8566) );
  NAND2_X1 U8668 ( .A1(n8562), .A2(n8564), .ZN(n8642) );
  NAND2_X1 U8669 ( .A1(n8643), .A2(n8644), .ZN(n8564) );
  NAND2_X1 U8670 ( .A1(n8556), .A2(n8645), .ZN(n8562) );
  NAND2_X1 U8671 ( .A1(n8554), .A2(n8557), .ZN(n8645) );
  NAND2_X1 U8672 ( .A1(n8646), .A2(n8647), .ZN(n8557) );
  NAND2_X1 U8673 ( .A1(n8648), .A2(n8649), .ZN(n8647) );
  XNOR2_X1 U8674 ( .A(n8650), .B(n8651), .ZN(n8646) );
  NAND2_X1 U8675 ( .A1(n8552), .A2(n8652), .ZN(n8554) );
  NAND2_X1 U8676 ( .A1(n8553), .A2(n8550), .ZN(n8652) );
  NAND2_X1 U8677 ( .A1(n8653), .A2(n8548), .ZN(n8550) );
  NAND2_X1 U8678 ( .A1(n8654), .A2(n8655), .ZN(n8548) );
  NAND2_X1 U8679 ( .A1(n8546), .A2(n8549), .ZN(n8653) );
  INV_X1 U8680 ( .A(n8656), .ZN(n8549) );
  NOR2_X1 U8681 ( .A1(n8654), .A2(n8655), .ZN(n8656) );
  XOR2_X1 U8682 ( .A(n8657), .B(n8658), .Z(n8654) );
  NAND2_X1 U8683 ( .A1(n8545), .A2(n8659), .ZN(n8546) );
  NAND2_X1 U8684 ( .A1(n8542), .A2(n8544), .ZN(n8659) );
  NAND2_X1 U8685 ( .A1(n8660), .A2(n8661), .ZN(n8544) );
  NAND2_X1 U8686 ( .A1(n8540), .A2(n8662), .ZN(n8542) );
  NAND2_X1 U8687 ( .A1(n8538), .A2(n8541), .ZN(n8662) );
  NAND2_X1 U8688 ( .A1(n8663), .A2(n8664), .ZN(n8541) );
  NAND2_X1 U8689 ( .A1(n8537), .A2(n8665), .ZN(n8538) );
  NAND2_X1 U8690 ( .A1(n8536), .A2(n8531), .ZN(n8665) );
  NAND2_X1 U8691 ( .A1(n8530), .A2(n8666), .ZN(n8531) );
  NAND2_X1 U8692 ( .A1(n8527), .A2(n8529), .ZN(n8666) );
  NAND2_X1 U8693 ( .A1(n8667), .A2(n8668), .ZN(n8529) );
  XOR2_X1 U8694 ( .A(n8669), .B(n8670), .Z(n8667) );
  NAND2_X1 U8695 ( .A1(n8525), .A2(n8671), .ZN(n8527) );
  NAND2_X1 U8696 ( .A1(n8523), .A2(n8526), .ZN(n8671) );
  NAND2_X1 U8697 ( .A1(n8672), .A2(n8673), .ZN(n8526) );
  NAND2_X1 U8698 ( .A1(n8521), .A2(n8674), .ZN(n8523) );
  NAND2_X1 U8699 ( .A1(n8520), .A2(n8522), .ZN(n8674) );
  NAND2_X1 U8700 ( .A1(n8675), .A2(n8676), .ZN(n8522) );
  INV_X1 U8701 ( .A(n8677), .ZN(n8676) );
  XOR2_X1 U8702 ( .A(n8678), .B(n8679), .Z(n8675) );
  NAND2_X1 U8703 ( .A1(n8518), .A2(n8680), .ZN(n8520) );
  NAND2_X1 U8704 ( .A1(n8509), .A2(n8517), .ZN(n8680) );
  NAND2_X1 U8705 ( .A1(n8681), .A2(n8682), .ZN(n8517) );
  NAND2_X1 U8706 ( .A1(n8683), .A2(n8684), .ZN(n8682) );
  NOR2_X1 U8707 ( .A1(n8685), .A2(n8508), .ZN(n8509) );
  XNOR2_X1 U8708 ( .A(n8686), .B(n8687), .ZN(n8508) );
  XOR2_X1 U8709 ( .A(n8688), .B(n8689), .Z(n8686) );
  NOR2_X1 U8710 ( .A1(n8690), .A2(n8364), .ZN(n8689) );
  NAND2_X1 U8711 ( .A1(n8513), .A2(n8512), .ZN(n8685) );
  XOR2_X1 U8712 ( .A(n8684), .B(n8683), .Z(n8512) );
  NAND2_X1 U8713 ( .A1(n8691), .A2(n8692), .ZN(n8513) );
  NAND2_X1 U8714 ( .A1(n8693), .A2(b_31_), .ZN(n8692) );
  NOR2_X1 U8715 ( .A1(n8694), .A2(n8690), .ZN(n8693) );
  NOR2_X1 U8716 ( .A1(n8503), .A2(n8505), .ZN(n8694) );
  NAND2_X1 U8717 ( .A1(n8503), .A2(n8505), .ZN(n8691) );
  NAND2_X1 U8718 ( .A1(n8695), .A2(n8696), .ZN(n8505) );
  NAND2_X1 U8719 ( .A1(n8697), .A2(b_31_), .ZN(n8696) );
  NOR2_X1 U8720 ( .A1(n8698), .A2(n8502), .ZN(n8697) );
  NOR2_X1 U8721 ( .A1(n8499), .A2(n8500), .ZN(n8698) );
  NAND2_X1 U8722 ( .A1(n8499), .A2(n8500), .ZN(n8695) );
  NAND2_X1 U8723 ( .A1(n8699), .A2(n8700), .ZN(n8500) );
  NAND2_X1 U8724 ( .A1(n8701), .A2(b_31_), .ZN(n8700) );
  NOR2_X1 U8725 ( .A1(n8702), .A2(n8497), .ZN(n8701) );
  NOR2_X1 U8726 ( .A1(n8494), .A2(n8495), .ZN(n8702) );
  NAND2_X1 U8727 ( .A1(n8494), .A2(n8495), .ZN(n8699) );
  NAND2_X1 U8728 ( .A1(n8703), .A2(n8704), .ZN(n8495) );
  NAND2_X1 U8729 ( .A1(n8705), .A2(b_31_), .ZN(n8704) );
  NOR2_X1 U8730 ( .A1(n8706), .A2(n8707), .ZN(n8705) );
  NOR2_X1 U8731 ( .A1(n8489), .A2(n8491), .ZN(n8706) );
  NAND2_X1 U8732 ( .A1(n8489), .A2(n8491), .ZN(n8703) );
  NAND2_X1 U8733 ( .A1(n8708), .A2(n8709), .ZN(n8491) );
  NAND2_X1 U8734 ( .A1(n8710), .A2(b_31_), .ZN(n8709) );
  NOR2_X1 U8735 ( .A1(n8711), .A2(n8712), .ZN(n8710) );
  NOR2_X1 U8736 ( .A1(n8485), .A2(n8487), .ZN(n8711) );
  NAND2_X1 U8737 ( .A1(n8485), .A2(n8487), .ZN(n8708) );
  NAND2_X1 U8738 ( .A1(n8713), .A2(n8714), .ZN(n8487) );
  NAND2_X1 U8739 ( .A1(n8715), .A2(b_31_), .ZN(n8714) );
  NOR2_X1 U8740 ( .A1(n8716), .A2(n8717), .ZN(n8715) );
  NOR2_X1 U8741 ( .A1(n8481), .A2(n8483), .ZN(n8716) );
  NAND2_X1 U8742 ( .A1(n8481), .A2(n8483), .ZN(n8713) );
  NAND2_X1 U8743 ( .A1(n8718), .A2(n8719), .ZN(n8483) );
  NAND2_X1 U8744 ( .A1(n8720), .A2(b_31_), .ZN(n8719) );
  NOR2_X1 U8745 ( .A1(n8721), .A2(n8480), .ZN(n8720) );
  NOR2_X1 U8746 ( .A1(n8477), .A2(n8478), .ZN(n8721) );
  NAND2_X1 U8747 ( .A1(n8477), .A2(n8478), .ZN(n8718) );
  NAND2_X1 U8748 ( .A1(n8722), .A2(n8723), .ZN(n8478) );
  NAND2_X1 U8749 ( .A1(n8724), .A2(b_31_), .ZN(n8723) );
  NOR2_X1 U8750 ( .A1(n8725), .A2(n8726), .ZN(n8724) );
  NOR2_X1 U8751 ( .A1(n8472), .A2(n8474), .ZN(n8725) );
  NAND2_X1 U8752 ( .A1(n8472), .A2(n8474), .ZN(n8722) );
  NAND2_X1 U8753 ( .A1(n8727), .A2(n8728), .ZN(n8474) );
  NAND2_X1 U8754 ( .A1(n8729), .A2(b_31_), .ZN(n8728) );
  NOR2_X1 U8755 ( .A1(n8730), .A2(n8731), .ZN(n8729) );
  NOR2_X1 U8756 ( .A1(n8461), .A2(n8463), .ZN(n8730) );
  NAND2_X1 U8757 ( .A1(n8461), .A2(n8463), .ZN(n8727) );
  NAND2_X1 U8758 ( .A1(n8732), .A2(n8733), .ZN(n8463) );
  NAND2_X1 U8759 ( .A1(n8734), .A2(b_31_), .ZN(n8733) );
  NOR2_X1 U8760 ( .A1(n8735), .A2(n8736), .ZN(n8734) );
  NOR2_X1 U8761 ( .A1(n8457), .A2(n8459), .ZN(n8735) );
  NAND2_X1 U8762 ( .A1(n8457), .A2(n8459), .ZN(n8732) );
  NAND2_X1 U8763 ( .A1(n8737), .A2(n8738), .ZN(n8459) );
  NAND2_X1 U8764 ( .A1(n8739), .A2(b_31_), .ZN(n8738) );
  NOR2_X1 U8765 ( .A1(n8740), .A2(n8741), .ZN(n8739) );
  NOR2_X1 U8766 ( .A1(n8453), .A2(n8455), .ZN(n8740) );
  NAND2_X1 U8767 ( .A1(n8453), .A2(n8455), .ZN(n8737) );
  NAND2_X1 U8768 ( .A1(n8742), .A2(n8743), .ZN(n8455) );
  NAND2_X1 U8769 ( .A1(n8744), .A2(b_31_), .ZN(n8743) );
  NOR2_X1 U8770 ( .A1(n8745), .A2(n8452), .ZN(n8744) );
  NOR2_X1 U8771 ( .A1(n8449), .A2(n8450), .ZN(n8745) );
  NAND2_X1 U8772 ( .A1(n8449), .A2(n8450), .ZN(n8742) );
  NAND2_X1 U8773 ( .A1(n8746), .A2(n8747), .ZN(n8450) );
  NAND2_X1 U8774 ( .A1(n8748), .A2(b_31_), .ZN(n8747) );
  NOR2_X1 U8775 ( .A1(n8749), .A2(n8750), .ZN(n8748) );
  NOR2_X1 U8776 ( .A1(n8444), .A2(n8446), .ZN(n8749) );
  NAND2_X1 U8777 ( .A1(n8444), .A2(n8446), .ZN(n8746) );
  NAND2_X1 U8778 ( .A1(n8751), .A2(n8752), .ZN(n8446) );
  NAND2_X1 U8779 ( .A1(n8753), .A2(b_31_), .ZN(n8752) );
  NOR2_X1 U8780 ( .A1(n8754), .A2(n8443), .ZN(n8753) );
  NOR2_X1 U8781 ( .A1(n8440), .A2(n8441), .ZN(n8754) );
  NAND2_X1 U8782 ( .A1(n8440), .A2(n8441), .ZN(n8751) );
  NAND2_X1 U8783 ( .A1(n8755), .A2(n8756), .ZN(n8441) );
  NAND2_X1 U8784 ( .A1(n8757), .A2(b_31_), .ZN(n8756) );
  NOR2_X1 U8785 ( .A1(n8758), .A2(n8438), .ZN(n8757) );
  NOR2_X1 U8786 ( .A1(n8435), .A2(n8436), .ZN(n8758) );
  NAND2_X1 U8787 ( .A1(n8435), .A2(n8436), .ZN(n8755) );
  NAND2_X1 U8788 ( .A1(n8759), .A2(n8760), .ZN(n8436) );
  NAND2_X1 U8789 ( .A1(n8761), .A2(b_31_), .ZN(n8760) );
  NOR2_X1 U8790 ( .A1(n8762), .A2(n8763), .ZN(n8761) );
  NOR2_X1 U8791 ( .A1(n8430), .A2(n8432), .ZN(n8762) );
  NAND2_X1 U8792 ( .A1(n8430), .A2(n8432), .ZN(n8759) );
  NAND2_X1 U8793 ( .A1(n8764), .A2(n8765), .ZN(n8432) );
  NAND2_X1 U8794 ( .A1(n8766), .A2(b_31_), .ZN(n8765) );
  NOR2_X1 U8795 ( .A1(n8767), .A2(n8768), .ZN(n8766) );
  NOR2_X1 U8796 ( .A1(n8427), .A2(n8429), .ZN(n8767) );
  NAND2_X1 U8797 ( .A1(n8427), .A2(n8429), .ZN(n8764) );
  NAND2_X1 U8798 ( .A1(n8769), .A2(n8770), .ZN(n8429) );
  NAND2_X1 U8799 ( .A1(n8425), .A2(n8771), .ZN(n8770) );
  NAND2_X1 U8800 ( .A1(n8424), .A2(n8422), .ZN(n8771) );
  NOR2_X1 U8801 ( .A1(n8360), .A2(n8772), .ZN(n8425) );
  INV_X1 U8802 ( .A(n8773), .ZN(n8769) );
  NOR2_X1 U8803 ( .A1(n8422), .A2(n8424), .ZN(n8773) );
  NOR2_X1 U8804 ( .A1(n8774), .A2(n8775), .ZN(n8424) );
  NOR2_X1 U8805 ( .A1(n8419), .A2(n8776), .ZN(n8775) );
  NOR2_X1 U8806 ( .A1(n8418), .A2(n8416), .ZN(n8776) );
  NAND2_X1 U8807 ( .A1(b_31_), .A2(a_18_), .ZN(n8419) );
  INV_X1 U8808 ( .A(n8777), .ZN(n8774) );
  NAND2_X1 U8809 ( .A1(n8416), .A2(n8418), .ZN(n8777) );
  NAND2_X1 U8810 ( .A1(n8778), .A2(n8779), .ZN(n8418) );
  NAND2_X1 U8811 ( .A1(n8412), .A2(n8780), .ZN(n8779) );
  NAND2_X1 U8812 ( .A1(n8415), .A2(n8414), .ZN(n8780) );
  XNOR2_X1 U8813 ( .A(n8781), .B(n8782), .ZN(n8412) );
  NAND2_X1 U8814 ( .A1(n8783), .A2(n8784), .ZN(n8781) );
  INV_X1 U8815 ( .A(n8785), .ZN(n8778) );
  NOR2_X1 U8816 ( .A1(n8414), .A2(n8415), .ZN(n8785) );
  NAND2_X1 U8817 ( .A1(b_31_), .A2(a_19_), .ZN(n8415) );
  NAND2_X1 U8818 ( .A1(n8786), .A2(n8787), .ZN(n8414) );
  NAND2_X1 U8819 ( .A1(n8788), .A2(n8410), .ZN(n8787) );
  NAND2_X1 U8820 ( .A1(b_31_), .A2(a_20_), .ZN(n8410) );
  NAND2_X1 U8821 ( .A1(n8408), .A2(n8411), .ZN(n8788) );
  INV_X1 U8822 ( .A(n8789), .ZN(n8786) );
  NOR2_X1 U8823 ( .A1(n8411), .A2(n8408), .ZN(n8789) );
  XNOR2_X1 U8824 ( .A(n8790), .B(n8791), .ZN(n8408) );
  NAND2_X1 U8825 ( .A1(n8792), .A2(n8793), .ZN(n8790) );
  NAND2_X1 U8826 ( .A1(n8794), .A2(n8795), .ZN(n8411) );
  NAND2_X1 U8827 ( .A1(n8407), .A2(n8796), .ZN(n8795) );
  INV_X1 U8828 ( .A(n8797), .ZN(n8796) );
  NOR2_X1 U8829 ( .A1(n8406), .A2(n8404), .ZN(n8797) );
  NOR2_X1 U8830 ( .A1(n8360), .A2(n8798), .ZN(n8407) );
  NAND2_X1 U8831 ( .A1(n8404), .A2(n8406), .ZN(n8794) );
  NAND2_X1 U8832 ( .A1(n8799), .A2(n8800), .ZN(n8406) );
  NAND2_X1 U8833 ( .A1(n8402), .A2(n8801), .ZN(n8800) );
  INV_X1 U8834 ( .A(n8802), .ZN(n8801) );
  NOR2_X1 U8835 ( .A1(n8403), .A2(n8400), .ZN(n8802) );
  NOR2_X1 U8836 ( .A1(n8360), .A2(n8803), .ZN(n8402) );
  NAND2_X1 U8837 ( .A1(n8400), .A2(n8403), .ZN(n8799) );
  NAND2_X1 U8838 ( .A1(n8398), .A2(n8804), .ZN(n8403) );
  NAND2_X1 U8839 ( .A1(n8397), .A2(n8399), .ZN(n8804) );
  NAND2_X1 U8840 ( .A1(n8805), .A2(n8806), .ZN(n8399) );
  NAND2_X1 U8841 ( .A1(b_31_), .A2(a_23_), .ZN(n8805) );
  XOR2_X1 U8842 ( .A(n8807), .B(n8808), .Z(n8397) );
  XOR2_X1 U8843 ( .A(n8809), .B(n8810), .Z(n8807) );
  INV_X1 U8844 ( .A(n8811), .ZN(n8398) );
  NOR2_X1 U8845 ( .A1(n8806), .A2(n8812), .ZN(n8811) );
  NAND2_X1 U8846 ( .A1(n8813), .A2(n8814), .ZN(n8806) );
  NAND2_X1 U8847 ( .A1(n8815), .A2(n8394), .ZN(n8814) );
  NAND2_X1 U8848 ( .A1(b_31_), .A2(a_24_), .ZN(n8394) );
  NAND2_X1 U8849 ( .A1(n8392), .A2(n8395), .ZN(n8815) );
  INV_X1 U8850 ( .A(n8816), .ZN(n8813) );
  NOR2_X1 U8851 ( .A1(n8395), .A2(n8392), .ZN(n8816) );
  XOR2_X1 U8852 ( .A(n8817), .B(n8818), .Z(n8392) );
  XOR2_X1 U8853 ( .A(n8819), .B(n8820), .Z(n8818) );
  NAND2_X1 U8854 ( .A1(n8821), .A2(n8822), .ZN(n8395) );
  NAND2_X1 U8855 ( .A1(n8391), .A2(n8823), .ZN(n8822) );
  INV_X1 U8856 ( .A(n8824), .ZN(n8823) );
  NOR2_X1 U8857 ( .A1(n8390), .A2(n8388), .ZN(n8824) );
  NOR2_X1 U8858 ( .A1(n8360), .A2(n8825), .ZN(n8391) );
  NAND2_X1 U8859 ( .A1(n8388), .A2(n8390), .ZN(n8821) );
  NAND2_X1 U8860 ( .A1(n8826), .A2(n8827), .ZN(n8390) );
  NAND2_X1 U8861 ( .A1(n8387), .A2(n8828), .ZN(n8827) );
  INV_X1 U8862 ( .A(n8829), .ZN(n8828) );
  NOR2_X1 U8863 ( .A1(n8386), .A2(n8384), .ZN(n8829) );
  NOR2_X1 U8864 ( .A1(n8360), .A2(n8830), .ZN(n8387) );
  NAND2_X1 U8865 ( .A1(n8384), .A2(n8386), .ZN(n8826) );
  NAND2_X1 U8866 ( .A1(n8382), .A2(n8831), .ZN(n8386) );
  NAND2_X1 U8867 ( .A1(n8381), .A2(n8383), .ZN(n8831) );
  NAND2_X1 U8868 ( .A1(n8832), .A2(n8833), .ZN(n8383) );
  NAND2_X1 U8869 ( .A1(b_31_), .A2(a_27_), .ZN(n8833) );
  XNOR2_X1 U8870 ( .A(n8834), .B(n8835), .ZN(n8381) );
  XNOR2_X1 U8871 ( .A(n8836), .B(n8837), .ZN(n8834) );
  INV_X1 U8872 ( .A(n8838), .ZN(n8382) );
  NOR2_X1 U8873 ( .A1(n8839), .A2(n8832), .ZN(n8838) );
  NOR2_X1 U8874 ( .A1(n8840), .A2(n8841), .ZN(n8832) );
  INV_X1 U8875 ( .A(n8842), .ZN(n8841) );
  NAND2_X1 U8876 ( .A1(n8372), .A2(n8843), .ZN(n8842) );
  NAND2_X1 U8877 ( .A1(n8370), .A2(n8371), .ZN(n8843) );
  NOR2_X1 U8878 ( .A1(n8360), .A2(n8844), .ZN(n8372) );
  INV_X1 U8879 ( .A(b_31_), .ZN(n8360) );
  NOR2_X1 U8880 ( .A1(n8371), .A2(n8370), .ZN(n8840) );
  XOR2_X1 U8881 ( .A(n8845), .B(n8846), .Z(n8370) );
  XOR2_X1 U8882 ( .A(n8847), .B(n8848), .Z(n8846) );
  NAND2_X1 U8883 ( .A1(n8849), .A2(n8850), .ZN(n8371) );
  NAND2_X1 U8884 ( .A1(n8851), .A2(n8367), .ZN(n8850) );
  NAND2_X1 U8885 ( .A1(b_31_), .A2(a_29_), .ZN(n8367) );
  NAND2_X1 U8886 ( .A1(n8365), .A2(n8368), .ZN(n8851) );
  INV_X1 U8887 ( .A(n8852), .ZN(n8365) );
  NAND2_X1 U8888 ( .A1(n8853), .A2(n8852), .ZN(n8849) );
  INV_X1 U8889 ( .A(n8368), .ZN(n8853) );
  NAND2_X1 U8890 ( .A1(n8854), .A2(n8855), .ZN(n8368) );
  NAND2_X1 U8891 ( .A1(b_29_), .A2(n8856), .ZN(n8855) );
  NAND2_X1 U8892 ( .A1(n8358), .A2(n8857), .ZN(n8856) );
  NAND2_X1 U8893 ( .A1(a_31_), .A2(n8364), .ZN(n8857) );
  NAND2_X1 U8894 ( .A1(b_30_), .A2(n8858), .ZN(n8854) );
  NAND2_X1 U8895 ( .A1(n8362), .A2(n8859), .ZN(n8858) );
  NAND2_X1 U8896 ( .A1(a_30_), .A2(n8860), .ZN(n8859) );
  XNOR2_X1 U8897 ( .A(n8861), .B(n8862), .ZN(n8384) );
  NAND2_X1 U8898 ( .A1(n8863), .A2(n8864), .ZN(n8861) );
  XNOR2_X1 U8899 ( .A(n8865), .B(n8866), .ZN(n8388) );
  XOR2_X1 U8900 ( .A(n8867), .B(n8868), .Z(n8865) );
  XOR2_X1 U8901 ( .A(n8869), .B(n8870), .Z(n8400) );
  XOR2_X1 U8902 ( .A(n8871), .B(n8872), .Z(n8869) );
  NOR2_X1 U8903 ( .A1(n8812), .A2(n8364), .ZN(n8872) );
  XNOR2_X1 U8904 ( .A(n8873), .B(n8874), .ZN(n8404) );
  XOR2_X1 U8905 ( .A(n8875), .B(n8876), .Z(n8873) );
  XOR2_X1 U8906 ( .A(n8877), .B(n8878), .Z(n8416) );
  XOR2_X1 U8907 ( .A(n8879), .B(n8880), .Z(n8877) );
  NOR2_X1 U8908 ( .A1(n8881), .A2(n8364), .ZN(n8880) );
  XOR2_X1 U8909 ( .A(n8882), .B(n8883), .Z(n8422) );
  NAND2_X1 U8910 ( .A1(n8884), .A2(n8885), .ZN(n8882) );
  XNOR2_X1 U8911 ( .A(n8886), .B(n8887), .ZN(n8427) );
  NAND2_X1 U8912 ( .A1(n8888), .A2(n8889), .ZN(n8886) );
  XNOR2_X1 U8913 ( .A(n8890), .B(n8891), .ZN(n8430) );
  NAND2_X1 U8914 ( .A1(n8892), .A2(n8893), .ZN(n8890) );
  XOR2_X1 U8915 ( .A(n8894), .B(n8895), .Z(n8435) );
  XOR2_X1 U8916 ( .A(n8896), .B(n8897), .Z(n8894) );
  NOR2_X1 U8917 ( .A1(n8763), .A2(n8364), .ZN(n8897) );
  XNOR2_X1 U8918 ( .A(n8898), .B(n8899), .ZN(n8440) );
  NAND2_X1 U8919 ( .A1(n8900), .A2(n8901), .ZN(n8898) );
  XNOR2_X1 U8920 ( .A(n8902), .B(n8903), .ZN(n8444) );
  NAND2_X1 U8921 ( .A1(n8904), .A2(n8905), .ZN(n8902) );
  XNOR2_X1 U8922 ( .A(n8906), .B(n8907), .ZN(n8449) );
  NAND2_X1 U8923 ( .A1(n8908), .A2(n8909), .ZN(n8906) );
  XOR2_X1 U8924 ( .A(n8910), .B(n8911), .Z(n8453) );
  XOR2_X1 U8925 ( .A(n8912), .B(n8913), .Z(n8910) );
  NOR2_X1 U8926 ( .A1(n8452), .A2(n8364), .ZN(n8913) );
  XOR2_X1 U8927 ( .A(n8914), .B(n8915), .Z(n8457) );
  XNOR2_X1 U8928 ( .A(n8916), .B(n8917), .ZN(n8915) );
  XOR2_X1 U8929 ( .A(n8918), .B(n8919), .Z(n8461) );
  XOR2_X1 U8930 ( .A(n8920), .B(n8921), .Z(n8918) );
  XNOR2_X1 U8931 ( .A(n8922), .B(n8923), .ZN(n8472) );
  NAND2_X1 U8932 ( .A1(n8924), .A2(n8925), .ZN(n8922) );
  XNOR2_X1 U8933 ( .A(n8926), .B(n8927), .ZN(n8477) );
  NAND2_X1 U8934 ( .A1(n8928), .A2(n8929), .ZN(n8926) );
  XOR2_X1 U8935 ( .A(n8930), .B(n8931), .Z(n8481) );
  XNOR2_X1 U8936 ( .A(n8932), .B(n8933), .ZN(n8931) );
  XNOR2_X1 U8937 ( .A(n8934), .B(n8935), .ZN(n8485) );
  NAND2_X1 U8938 ( .A1(n8936), .A2(n8937), .ZN(n8934) );
  XNOR2_X1 U8939 ( .A(n8938), .B(n8939), .ZN(n8489) );
  NAND2_X1 U8940 ( .A1(n8940), .A2(n8941), .ZN(n8938) );
  XNOR2_X1 U8941 ( .A(n8942), .B(n8943), .ZN(n8494) );
  NAND2_X1 U8942 ( .A1(n8944), .A2(n8945), .ZN(n8942) );
  XNOR2_X1 U8943 ( .A(n8946), .B(n8947), .ZN(n8499) );
  XOR2_X1 U8944 ( .A(n8948), .B(n8949), .Z(n8946) );
  XOR2_X1 U8945 ( .A(n8950), .B(n8951), .Z(n8503) );
  XOR2_X1 U8946 ( .A(n8952), .B(n8953), .Z(n8950) );
  NAND2_X1 U8947 ( .A1(n8954), .A2(n8683), .ZN(n8518) );
  XNOR2_X1 U8948 ( .A(n8955), .B(n8956), .ZN(n8683) );
  XNOR2_X1 U8949 ( .A(n8957), .B(n8958), .ZN(n8955) );
  NOR2_X1 U8950 ( .A1(n8959), .A2(n8681), .ZN(n8954) );
  XNOR2_X1 U8951 ( .A(n8960), .B(n8961), .ZN(n8681) );
  INV_X1 U8952 ( .A(n8684), .ZN(n8959) );
  NAND2_X1 U8953 ( .A1(n8962), .A2(n8963), .ZN(n8684) );
  NAND2_X1 U8954 ( .A1(n8964), .A2(b_30_), .ZN(n8963) );
  NOR2_X1 U8955 ( .A1(n8965), .A2(n8690), .ZN(n8964) );
  NOR2_X1 U8956 ( .A1(n8687), .A2(n8688), .ZN(n8965) );
  NAND2_X1 U8957 ( .A1(n8687), .A2(n8688), .ZN(n8962) );
  NAND2_X1 U8958 ( .A1(n8966), .A2(n8967), .ZN(n8688) );
  NAND2_X1 U8959 ( .A1(n8953), .A2(n8968), .ZN(n8967) );
  NAND2_X1 U8960 ( .A1(n8951), .A2(n8952), .ZN(n8968) );
  NOR2_X1 U8961 ( .A1(n8364), .A2(n8502), .ZN(n8953) );
  NAND2_X1 U8962 ( .A1(n8969), .A2(n8970), .ZN(n8966) );
  INV_X1 U8963 ( .A(n8952), .ZN(n8970) );
  NAND2_X1 U8964 ( .A1(n8971), .A2(n8972), .ZN(n8952) );
  NAND2_X1 U8965 ( .A1(n8947), .A2(n8973), .ZN(n8972) );
  NAND2_X1 U8966 ( .A1(n8949), .A2(n8948), .ZN(n8973) );
  XOR2_X1 U8967 ( .A(n8974), .B(n8975), .Z(n8947) );
  NAND2_X1 U8968 ( .A1(n8976), .A2(n8977), .ZN(n8974) );
  INV_X1 U8969 ( .A(n8978), .ZN(n8971) );
  NOR2_X1 U8970 ( .A1(n8948), .A2(n8949), .ZN(n8978) );
  NOR2_X1 U8971 ( .A1(n8364), .A2(n8497), .ZN(n8949) );
  NAND2_X1 U8972 ( .A1(n8944), .A2(n8979), .ZN(n8948) );
  NAND2_X1 U8973 ( .A1(n8943), .A2(n8945), .ZN(n8979) );
  NAND2_X1 U8974 ( .A1(n8980), .A2(n8981), .ZN(n8945) );
  NAND2_X1 U8975 ( .A1(b_30_), .A2(a_3_), .ZN(n8981) );
  INV_X1 U8976 ( .A(n8982), .ZN(n8980) );
  XNOR2_X1 U8977 ( .A(n8983), .B(n8984), .ZN(n8943) );
  NAND2_X1 U8978 ( .A1(n8985), .A2(n8986), .ZN(n8983) );
  NAND2_X1 U8979 ( .A1(a_3_), .A2(n8982), .ZN(n8944) );
  NAND2_X1 U8980 ( .A1(n8940), .A2(n8987), .ZN(n8982) );
  NAND2_X1 U8981 ( .A1(n8939), .A2(n8941), .ZN(n8987) );
  NAND2_X1 U8982 ( .A1(n8988), .A2(n8989), .ZN(n8941) );
  NAND2_X1 U8983 ( .A1(b_30_), .A2(a_4_), .ZN(n8989) );
  INV_X1 U8984 ( .A(n8990), .ZN(n8988) );
  XOR2_X1 U8985 ( .A(n8991), .B(n8992), .Z(n8939) );
  XNOR2_X1 U8986 ( .A(n8993), .B(n8994), .ZN(n8992) );
  NAND2_X1 U8987 ( .A1(b_29_), .A2(a_5_), .ZN(n8994) );
  NAND2_X1 U8988 ( .A1(a_4_), .A2(n8990), .ZN(n8940) );
  NAND2_X1 U8989 ( .A1(n8936), .A2(n8995), .ZN(n8990) );
  NAND2_X1 U8990 ( .A1(n8935), .A2(n8937), .ZN(n8995) );
  NAND2_X1 U8991 ( .A1(n8996), .A2(n8997), .ZN(n8937) );
  INV_X1 U8992 ( .A(n8998), .ZN(n8997) );
  NAND2_X1 U8993 ( .A1(b_30_), .A2(a_5_), .ZN(n8996) );
  XNOR2_X1 U8994 ( .A(n8999), .B(n9000), .ZN(n8935) );
  XOR2_X1 U8995 ( .A(n9001), .B(n9002), .Z(n8999) );
  NAND2_X1 U8996 ( .A1(n8998), .A2(a_5_), .ZN(n8936) );
  NOR2_X1 U8997 ( .A1(n9003), .A2(n9004), .ZN(n8998) );
  INV_X1 U8998 ( .A(n9005), .ZN(n9004) );
  NAND2_X1 U8999 ( .A1(n8930), .A2(n9006), .ZN(n9005) );
  NAND2_X1 U9000 ( .A1(n8933), .A2(n8932), .ZN(n9006) );
  XOR2_X1 U9001 ( .A(n9007), .B(n9008), .Z(n8930) );
  NAND2_X1 U9002 ( .A1(n9009), .A2(n9010), .ZN(n9007) );
  NOR2_X1 U9003 ( .A1(n8932), .A2(n8933), .ZN(n9003) );
  NOR2_X1 U9004 ( .A1(n8364), .A2(n8480), .ZN(n8933) );
  NAND2_X1 U9005 ( .A1(n8928), .A2(n9011), .ZN(n8932) );
  NAND2_X1 U9006 ( .A1(n8927), .A2(n8929), .ZN(n9011) );
  NAND2_X1 U9007 ( .A1(n9012), .A2(n9013), .ZN(n8929) );
  NAND2_X1 U9008 ( .A1(b_30_), .A2(a_7_), .ZN(n9013) );
  INV_X1 U9009 ( .A(n9014), .ZN(n9012) );
  XOR2_X1 U9010 ( .A(n9015), .B(n9016), .Z(n8927) );
  XNOR2_X1 U9011 ( .A(n9017), .B(n9018), .ZN(n9016) );
  NAND2_X1 U9012 ( .A1(a_7_), .A2(n9014), .ZN(n8928) );
  NAND2_X1 U9013 ( .A1(n8924), .A2(n9019), .ZN(n9014) );
  NAND2_X1 U9014 ( .A1(n8923), .A2(n8925), .ZN(n9019) );
  NAND2_X1 U9015 ( .A1(n9020), .A2(n9021), .ZN(n8925) );
  NAND2_X1 U9016 ( .A1(b_30_), .A2(a_8_), .ZN(n9021) );
  XOR2_X1 U9017 ( .A(n9022), .B(n9023), .Z(n8923) );
  XOR2_X1 U9018 ( .A(n9024), .B(n9025), .Z(n9022) );
  NOR2_X1 U9019 ( .A1(n8736), .A2(n8860), .ZN(n9025) );
  INV_X1 U9020 ( .A(n9026), .ZN(n8924) );
  NOR2_X1 U9021 ( .A1(n8731), .A2(n9020), .ZN(n9026) );
  NOR2_X1 U9022 ( .A1(n9027), .A2(n9028), .ZN(n9020) );
  INV_X1 U9023 ( .A(n9029), .ZN(n9028) );
  NAND2_X1 U9024 ( .A1(n8921), .A2(n9030), .ZN(n9029) );
  NAND2_X1 U9025 ( .A1(n8919), .A2(n8920), .ZN(n9030) );
  NOR2_X1 U9026 ( .A1(n8364), .A2(n8736), .ZN(n8921) );
  NOR2_X1 U9027 ( .A1(n8919), .A2(n8920), .ZN(n9027) );
  NAND2_X1 U9028 ( .A1(n9031), .A2(n9032), .ZN(n8920) );
  NAND2_X1 U9029 ( .A1(n8914), .A2(n9033), .ZN(n9032) );
  NAND2_X1 U9030 ( .A1(n8917), .A2(n8916), .ZN(n9033) );
  XNOR2_X1 U9031 ( .A(n9034), .B(n9035), .ZN(n8914) );
  XOR2_X1 U9032 ( .A(n9036), .B(n9037), .Z(n9034) );
  NOR2_X1 U9033 ( .A1(n8452), .A2(n8860), .ZN(n9037) );
  INV_X1 U9034 ( .A(n9038), .ZN(n9031) );
  NOR2_X1 U9035 ( .A1(n8916), .A2(n8917), .ZN(n9038) );
  NOR2_X1 U9036 ( .A1(n8364), .A2(n8741), .ZN(n8917) );
  NAND2_X1 U9037 ( .A1(n9039), .A2(n9040), .ZN(n8916) );
  NAND2_X1 U9038 ( .A1(n9041), .A2(b_30_), .ZN(n9040) );
  NOR2_X1 U9039 ( .A1(n9042), .A2(n8452), .ZN(n9041) );
  NOR2_X1 U9040 ( .A1(n8912), .A2(n8911), .ZN(n9042) );
  NAND2_X1 U9041 ( .A1(n8911), .A2(n8912), .ZN(n9039) );
  NAND2_X1 U9042 ( .A1(n8908), .A2(n9043), .ZN(n8912) );
  NAND2_X1 U9043 ( .A1(n8907), .A2(n8909), .ZN(n9043) );
  NAND2_X1 U9044 ( .A1(n9044), .A2(n9045), .ZN(n8909) );
  NAND2_X1 U9045 ( .A1(b_30_), .A2(a_12_), .ZN(n9045) );
  INV_X1 U9046 ( .A(n9046), .ZN(n9044) );
  XNOR2_X1 U9047 ( .A(n9047), .B(n9048), .ZN(n8907) );
  NAND2_X1 U9048 ( .A1(n9049), .A2(n9050), .ZN(n9047) );
  NAND2_X1 U9049 ( .A1(a_12_), .A2(n9046), .ZN(n8908) );
  NAND2_X1 U9050 ( .A1(n8904), .A2(n9051), .ZN(n9046) );
  NAND2_X1 U9051 ( .A1(n8903), .A2(n8905), .ZN(n9051) );
  NAND2_X1 U9052 ( .A1(n9052), .A2(n9053), .ZN(n8905) );
  NAND2_X1 U9053 ( .A1(b_30_), .A2(a_13_), .ZN(n9053) );
  INV_X1 U9054 ( .A(n9054), .ZN(n9052) );
  XNOR2_X1 U9055 ( .A(n9055), .B(n9056), .ZN(n8903) );
  NAND2_X1 U9056 ( .A1(n9057), .A2(n9058), .ZN(n9055) );
  NAND2_X1 U9057 ( .A1(a_13_), .A2(n9054), .ZN(n8904) );
  NAND2_X1 U9058 ( .A1(n8900), .A2(n9059), .ZN(n9054) );
  NAND2_X1 U9059 ( .A1(n8899), .A2(n8901), .ZN(n9059) );
  NAND2_X1 U9060 ( .A1(n9060), .A2(n9061), .ZN(n8901) );
  NAND2_X1 U9061 ( .A1(b_30_), .A2(a_14_), .ZN(n9061) );
  INV_X1 U9062 ( .A(n9062), .ZN(n9060) );
  XOR2_X1 U9063 ( .A(n9063), .B(n9064), .Z(n8899) );
  XOR2_X1 U9064 ( .A(n9065), .B(n9066), .Z(n9063) );
  NOR2_X1 U9065 ( .A1(n8763), .A2(n8860), .ZN(n9066) );
  NAND2_X1 U9066 ( .A1(a_14_), .A2(n9062), .ZN(n8900) );
  NAND2_X1 U9067 ( .A1(n9067), .A2(n9068), .ZN(n9062) );
  NAND2_X1 U9068 ( .A1(n9069), .A2(b_30_), .ZN(n9068) );
  NOR2_X1 U9069 ( .A1(n9070), .A2(n8763), .ZN(n9069) );
  NOR2_X1 U9070 ( .A1(n8895), .A2(n8896), .ZN(n9070) );
  NAND2_X1 U9071 ( .A1(n8895), .A2(n8896), .ZN(n9067) );
  NAND2_X1 U9072 ( .A1(n8892), .A2(n9071), .ZN(n8896) );
  NAND2_X1 U9073 ( .A1(n8891), .A2(n8893), .ZN(n9071) );
  NAND2_X1 U9074 ( .A1(n9072), .A2(n9073), .ZN(n8893) );
  NAND2_X1 U9075 ( .A1(b_30_), .A2(a_16_), .ZN(n9073) );
  INV_X1 U9076 ( .A(n9074), .ZN(n9072) );
  XNOR2_X1 U9077 ( .A(n9075), .B(n9076), .ZN(n8891) );
  NAND2_X1 U9078 ( .A1(n9077), .A2(n9078), .ZN(n9075) );
  NAND2_X1 U9079 ( .A1(a_16_), .A2(n9074), .ZN(n8892) );
  NAND2_X1 U9080 ( .A1(n8888), .A2(n9079), .ZN(n9074) );
  NAND2_X1 U9081 ( .A1(n8887), .A2(n8889), .ZN(n9079) );
  NAND2_X1 U9082 ( .A1(n9080), .A2(n9081), .ZN(n8889) );
  NAND2_X1 U9083 ( .A1(b_30_), .A2(a_17_), .ZN(n9081) );
  INV_X1 U9084 ( .A(n9082), .ZN(n9080) );
  XNOR2_X1 U9085 ( .A(n9083), .B(n9084), .ZN(n8887) );
  NAND2_X1 U9086 ( .A1(n9085), .A2(n9086), .ZN(n9083) );
  NAND2_X1 U9087 ( .A1(a_17_), .A2(n9082), .ZN(n8888) );
  NAND2_X1 U9088 ( .A1(n8884), .A2(n9087), .ZN(n9082) );
  NAND2_X1 U9089 ( .A1(n8883), .A2(n8885), .ZN(n9087) );
  NAND2_X1 U9090 ( .A1(n9088), .A2(n9089), .ZN(n8885) );
  NAND2_X1 U9091 ( .A1(b_30_), .A2(a_18_), .ZN(n9089) );
  INV_X1 U9092 ( .A(n9090), .ZN(n9088) );
  XOR2_X1 U9093 ( .A(n9091), .B(n9092), .Z(n8883) );
  XOR2_X1 U9094 ( .A(n9093), .B(n9094), .Z(n9091) );
  NOR2_X1 U9095 ( .A1(n8881), .A2(n8860), .ZN(n9094) );
  NAND2_X1 U9096 ( .A1(a_18_), .A2(n9090), .ZN(n8884) );
  NAND2_X1 U9097 ( .A1(n9095), .A2(n9096), .ZN(n9090) );
  NAND2_X1 U9098 ( .A1(n9097), .A2(b_30_), .ZN(n9096) );
  NOR2_X1 U9099 ( .A1(n9098), .A2(n8881), .ZN(n9097) );
  NOR2_X1 U9100 ( .A1(n8878), .A2(n8879), .ZN(n9098) );
  NAND2_X1 U9101 ( .A1(n8878), .A2(n8879), .ZN(n9095) );
  NAND2_X1 U9102 ( .A1(n8783), .A2(n9099), .ZN(n8879) );
  NAND2_X1 U9103 ( .A1(n8782), .A2(n8784), .ZN(n9099) );
  NAND2_X1 U9104 ( .A1(n9100), .A2(n9101), .ZN(n8784) );
  NAND2_X1 U9105 ( .A1(b_30_), .A2(a_20_), .ZN(n9101) );
  INV_X1 U9106 ( .A(n9102), .ZN(n9100) );
  XNOR2_X1 U9107 ( .A(n9103), .B(n9104), .ZN(n8782) );
  NAND2_X1 U9108 ( .A1(n9105), .A2(n9106), .ZN(n9103) );
  NAND2_X1 U9109 ( .A1(a_20_), .A2(n9102), .ZN(n8783) );
  NAND2_X1 U9110 ( .A1(n8792), .A2(n9107), .ZN(n9102) );
  NAND2_X1 U9111 ( .A1(n8791), .A2(n8793), .ZN(n9107) );
  NAND2_X1 U9112 ( .A1(n9108), .A2(n9109), .ZN(n8793) );
  INV_X1 U9113 ( .A(n9110), .ZN(n9109) );
  NAND2_X1 U9114 ( .A1(b_30_), .A2(a_21_), .ZN(n9108) );
  XNOR2_X1 U9115 ( .A(n9111), .B(n9112), .ZN(n8791) );
  NAND2_X1 U9116 ( .A1(n9113), .A2(n9114), .ZN(n9111) );
  NAND2_X1 U9117 ( .A1(n9110), .A2(a_21_), .ZN(n8792) );
  NOR2_X1 U9118 ( .A1(n9115), .A2(n9116), .ZN(n9110) );
  INV_X1 U9119 ( .A(n9117), .ZN(n9116) );
  NAND2_X1 U9120 ( .A1(n8874), .A2(n9118), .ZN(n9117) );
  NAND2_X1 U9121 ( .A1(n8876), .A2(n8875), .ZN(n9118) );
  XOR2_X1 U9122 ( .A(n9119), .B(n9120), .Z(n8874) );
  XOR2_X1 U9123 ( .A(n9121), .B(n9122), .Z(n9120) );
  NAND2_X1 U9124 ( .A1(b_29_), .A2(a_23_), .ZN(n9122) );
  NOR2_X1 U9125 ( .A1(n8875), .A2(n8876), .ZN(n9115) );
  NOR2_X1 U9126 ( .A1(n8364), .A2(n8803), .ZN(n8876) );
  NAND2_X1 U9127 ( .A1(n9123), .A2(n9124), .ZN(n8875) );
  NAND2_X1 U9128 ( .A1(n9125), .A2(b_30_), .ZN(n9124) );
  NOR2_X1 U9129 ( .A1(n9126), .A2(n8812), .ZN(n9125) );
  NOR2_X1 U9130 ( .A1(n8871), .A2(n8870), .ZN(n9126) );
  NAND2_X1 U9131 ( .A1(n8870), .A2(n8871), .ZN(n9123) );
  NAND2_X1 U9132 ( .A1(n9127), .A2(n9128), .ZN(n8871) );
  NAND2_X1 U9133 ( .A1(n8810), .A2(n9129), .ZN(n9128) );
  INV_X1 U9134 ( .A(n9130), .ZN(n9129) );
  NOR2_X1 U9135 ( .A1(n8808), .A2(n8809), .ZN(n9130) );
  NOR2_X1 U9136 ( .A1(n8364), .A2(n9131), .ZN(n8810) );
  NAND2_X1 U9137 ( .A1(n8808), .A2(n8809), .ZN(n9127) );
  NAND2_X1 U9138 ( .A1(n9132), .A2(n9133), .ZN(n8809) );
  NAND2_X1 U9139 ( .A1(n8820), .A2(n9134), .ZN(n9133) );
  INV_X1 U9140 ( .A(n9135), .ZN(n9134) );
  NOR2_X1 U9141 ( .A1(n8817), .A2(n8819), .ZN(n9135) );
  NOR2_X1 U9142 ( .A1(n8364), .A2(n8825), .ZN(n8820) );
  NAND2_X1 U9143 ( .A1(n8817), .A2(n8819), .ZN(n9132) );
  NOR2_X1 U9144 ( .A1(n9136), .A2(n9137), .ZN(n8819) );
  INV_X1 U9145 ( .A(n9138), .ZN(n9137) );
  NAND2_X1 U9146 ( .A1(n8866), .A2(n9139), .ZN(n9138) );
  NAND2_X1 U9147 ( .A1(n8868), .A2(n8867), .ZN(n9139) );
  XOR2_X1 U9148 ( .A(n9140), .B(n9141), .Z(n8866) );
  NAND2_X1 U9149 ( .A1(n9142), .A2(n9143), .ZN(n9140) );
  NOR2_X1 U9150 ( .A1(n8867), .A2(n8868), .ZN(n9136) );
  NOR2_X1 U9151 ( .A1(n8364), .A2(n8830), .ZN(n8868) );
  NAND2_X1 U9152 ( .A1(n8863), .A2(n9144), .ZN(n8867) );
  NAND2_X1 U9153 ( .A1(n8862), .A2(n8864), .ZN(n9144) );
  NAND2_X1 U9154 ( .A1(n9145), .A2(n9146), .ZN(n8864) );
  NAND2_X1 U9155 ( .A1(b_30_), .A2(a_27_), .ZN(n9146) );
  XNOR2_X1 U9156 ( .A(n9147), .B(n9148), .ZN(n8862) );
  XNOR2_X1 U9157 ( .A(n9149), .B(n9150), .ZN(n9147) );
  NOR2_X1 U9158 ( .A1(n8844), .A2(n8860), .ZN(n9150) );
  INV_X1 U9159 ( .A(n9151), .ZN(n8863) );
  NOR2_X1 U9160 ( .A1(n8839), .A2(n9145), .ZN(n9151) );
  NOR2_X1 U9161 ( .A1(n9152), .A2(n9153), .ZN(n9145) );
  INV_X1 U9162 ( .A(n9154), .ZN(n9153) );
  NAND2_X1 U9163 ( .A1(n8836), .A2(n9155), .ZN(n9154) );
  NAND2_X1 U9164 ( .A1(n8837), .A2(n8835), .ZN(n9155) );
  NOR2_X1 U9165 ( .A1(n8364), .A2(n8844), .ZN(n8836) );
  NOR2_X1 U9166 ( .A1(n8835), .A2(n8837), .ZN(n9152) );
  NOR2_X1 U9167 ( .A1(n9156), .A2(n9157), .ZN(n8837) );
  INV_X1 U9168 ( .A(n9158), .ZN(n9157) );
  NAND2_X1 U9169 ( .A1(n8845), .A2(n9159), .ZN(n9158) );
  NAND2_X1 U9170 ( .A1(n9160), .A2(n8847), .ZN(n9159) );
  NOR2_X1 U9171 ( .A1(n8364), .A2(n9161), .ZN(n8845) );
  NOR2_X1 U9172 ( .A1(n8847), .A2(n9160), .ZN(n9156) );
  INV_X1 U9173 ( .A(n8848), .ZN(n9160) );
  NAND2_X1 U9174 ( .A1(n9162), .A2(n9163), .ZN(n8848) );
  NAND2_X1 U9175 ( .A1(b_28_), .A2(n9164), .ZN(n9163) );
  NAND2_X1 U9176 ( .A1(n8358), .A2(n9165), .ZN(n9164) );
  NAND2_X1 U9177 ( .A1(a_31_), .A2(n8860), .ZN(n9165) );
  NAND2_X1 U9178 ( .A1(b_29_), .A2(n9166), .ZN(n9162) );
  NAND2_X1 U9179 ( .A1(n8362), .A2(n9167), .ZN(n9166) );
  NAND2_X1 U9180 ( .A1(a_30_), .A2(n9168), .ZN(n9167) );
  NAND2_X1 U9181 ( .A1(n9169), .A2(b_30_), .ZN(n8847) );
  NOR2_X1 U9182 ( .A1(n9170), .A2(n8860), .ZN(n9169) );
  XOR2_X1 U9183 ( .A(n9171), .B(n9172), .Z(n8835) );
  XOR2_X1 U9184 ( .A(n9173), .B(n9174), .Z(n9172) );
  XOR2_X1 U9185 ( .A(n9175), .B(n9176), .Z(n8817) );
  XNOR2_X1 U9186 ( .A(n9177), .B(n9178), .ZN(n9176) );
  XNOR2_X1 U9187 ( .A(n9179), .B(n9180), .ZN(n8808) );
  XNOR2_X1 U9188 ( .A(n9181), .B(n9182), .ZN(n9179) );
  XOR2_X1 U9189 ( .A(n9183), .B(n9184), .Z(n8870) );
  XOR2_X1 U9190 ( .A(n9185), .B(n9186), .Z(n9183) );
  NOR2_X1 U9191 ( .A1(n9131), .A2(n8860), .ZN(n9186) );
  XNOR2_X1 U9192 ( .A(n9187), .B(n9188), .ZN(n8878) );
  NAND2_X1 U9193 ( .A1(n9189), .A2(n9190), .ZN(n9187) );
  XNOR2_X1 U9194 ( .A(n9191), .B(n9192), .ZN(n8895) );
  NAND2_X1 U9195 ( .A1(n9193), .A2(n9194), .ZN(n9191) );
  XNOR2_X1 U9196 ( .A(n9195), .B(n9196), .ZN(n8911) );
  NAND2_X1 U9197 ( .A1(n9197), .A2(n9198), .ZN(n9195) );
  XOR2_X1 U9198 ( .A(n9199), .B(n9200), .Z(n8919) );
  NAND2_X1 U9199 ( .A1(n9201), .A2(n9202), .ZN(n9199) );
  INV_X1 U9200 ( .A(n8951), .ZN(n8969) );
  XNOR2_X1 U9201 ( .A(n9203), .B(n9204), .ZN(n8951) );
  XOR2_X1 U9202 ( .A(n9205), .B(n9206), .Z(n9203) );
  XNOR2_X1 U9203 ( .A(n9207), .B(n9208), .ZN(n8687) );
  XOR2_X1 U9204 ( .A(n9209), .B(n9210), .Z(n9207) );
  NAND2_X1 U9205 ( .A1(n8677), .A2(n9211), .ZN(n8521) );
  XOR2_X1 U9206 ( .A(n9212), .B(n8679), .Z(n9211) );
  NOR2_X1 U9207 ( .A1(n8961), .A2(n8960), .ZN(n8677) );
  NOR2_X1 U9208 ( .A1(n9213), .A2(n9214), .ZN(n8960) );
  INV_X1 U9209 ( .A(n9215), .ZN(n9214) );
  NAND2_X1 U9210 ( .A1(n8957), .A2(n9216), .ZN(n9215) );
  NAND2_X1 U9211 ( .A1(n8958), .A2(n8956), .ZN(n9216) );
  NOR2_X1 U9212 ( .A1(n8860), .A2(n8690), .ZN(n8957) );
  NOR2_X1 U9213 ( .A1(n8956), .A2(n8958), .ZN(n9213) );
  NOR2_X1 U9214 ( .A1(n9217), .A2(n9218), .ZN(n8958) );
  INV_X1 U9215 ( .A(n9219), .ZN(n9218) );
  NAND2_X1 U9216 ( .A1(n9210), .A2(n9220), .ZN(n9219) );
  NAND2_X1 U9217 ( .A1(n9221), .A2(n9208), .ZN(n9220) );
  NOR2_X1 U9218 ( .A1(n8860), .A2(n8502), .ZN(n9210) );
  NOR2_X1 U9219 ( .A1(n9208), .A2(n9221), .ZN(n9217) );
  INV_X1 U9220 ( .A(n9209), .ZN(n9221) );
  NAND2_X1 U9221 ( .A1(n9222), .A2(n9223), .ZN(n9209) );
  NAND2_X1 U9222 ( .A1(n9205), .A2(n9224), .ZN(n9223) );
  INV_X1 U9223 ( .A(n9225), .ZN(n9224) );
  NOR2_X1 U9224 ( .A1(n9204), .A2(n9206), .ZN(n9225) );
  NAND2_X1 U9225 ( .A1(n8976), .A2(n9226), .ZN(n9205) );
  NAND2_X1 U9226 ( .A1(n8975), .A2(n8977), .ZN(n9226) );
  NAND2_X1 U9227 ( .A1(n9227), .A2(n9228), .ZN(n8977) );
  NAND2_X1 U9228 ( .A1(b_29_), .A2(a_3_), .ZN(n9228) );
  INV_X1 U9229 ( .A(n9229), .ZN(n9227) );
  XNOR2_X1 U9230 ( .A(n9230), .B(n9231), .ZN(n8975) );
  XOR2_X1 U9231 ( .A(n9232), .B(n9233), .Z(n9231) );
  NAND2_X1 U9232 ( .A1(b_28_), .A2(a_4_), .ZN(n9233) );
  NAND2_X1 U9233 ( .A1(a_3_), .A2(n9229), .ZN(n8976) );
  NAND2_X1 U9234 ( .A1(n8985), .A2(n9234), .ZN(n9229) );
  NAND2_X1 U9235 ( .A1(n8984), .A2(n8986), .ZN(n9234) );
  NAND2_X1 U9236 ( .A1(n9235), .A2(n9236), .ZN(n8986) );
  NAND2_X1 U9237 ( .A1(b_29_), .A2(a_4_), .ZN(n9236) );
  INV_X1 U9238 ( .A(n9237), .ZN(n9235) );
  XNOR2_X1 U9239 ( .A(n9238), .B(n9239), .ZN(n8984) );
  XNOR2_X1 U9240 ( .A(n9240), .B(n9241), .ZN(n9238) );
  NOR2_X1 U9241 ( .A1(n8717), .A2(n9168), .ZN(n9241) );
  NAND2_X1 U9242 ( .A1(a_4_), .A2(n9237), .ZN(n8985) );
  NAND2_X1 U9243 ( .A1(n9242), .A2(n9243), .ZN(n9237) );
  NAND2_X1 U9244 ( .A1(n9244), .A2(b_29_), .ZN(n9243) );
  NOR2_X1 U9245 ( .A1(n9245), .A2(n8717), .ZN(n9244) );
  NOR2_X1 U9246 ( .A1(n8993), .A2(n8991), .ZN(n9245) );
  NAND2_X1 U9247 ( .A1(n8993), .A2(n8991), .ZN(n9242) );
  XOR2_X1 U9248 ( .A(n9246), .B(n9247), .Z(n8991) );
  XNOR2_X1 U9249 ( .A(n9248), .B(n9249), .ZN(n9247) );
  NOR2_X1 U9250 ( .A1(n9250), .A2(n9251), .ZN(n8993) );
  INV_X1 U9251 ( .A(n9252), .ZN(n9251) );
  NAND2_X1 U9252 ( .A1(n9000), .A2(n9253), .ZN(n9252) );
  NAND2_X1 U9253 ( .A1(n9002), .A2(n9001), .ZN(n9253) );
  XOR2_X1 U9254 ( .A(n9254), .B(n9255), .Z(n9000) );
  NAND2_X1 U9255 ( .A1(n9256), .A2(n9257), .ZN(n9254) );
  NOR2_X1 U9256 ( .A1(n9001), .A2(n9002), .ZN(n9250) );
  NOR2_X1 U9257 ( .A1(n8860), .A2(n8480), .ZN(n9002) );
  NAND2_X1 U9258 ( .A1(n9009), .A2(n9258), .ZN(n9001) );
  NAND2_X1 U9259 ( .A1(n9008), .A2(n9010), .ZN(n9258) );
  NAND2_X1 U9260 ( .A1(n9259), .A2(n9260), .ZN(n9010) );
  INV_X1 U9261 ( .A(n9261), .ZN(n9260) );
  NAND2_X1 U9262 ( .A1(b_29_), .A2(a_7_), .ZN(n9259) );
  XNOR2_X1 U9263 ( .A(n9262), .B(n9263), .ZN(n9008) );
  NAND2_X1 U9264 ( .A1(n9264), .A2(n9265), .ZN(n9262) );
  NAND2_X1 U9265 ( .A1(n9261), .A2(a_7_), .ZN(n9009) );
  NOR2_X1 U9266 ( .A1(n9266), .A2(n9267), .ZN(n9261) );
  INV_X1 U9267 ( .A(n9268), .ZN(n9267) );
  NAND2_X1 U9268 ( .A1(n9015), .A2(n9269), .ZN(n9268) );
  NAND2_X1 U9269 ( .A1(n9018), .A2(n9017), .ZN(n9269) );
  XOR2_X1 U9270 ( .A(n9270), .B(n9271), .Z(n9015) );
  NAND2_X1 U9271 ( .A1(n9272), .A2(n9273), .ZN(n9270) );
  NOR2_X1 U9272 ( .A1(n9017), .A2(n9018), .ZN(n9266) );
  NOR2_X1 U9273 ( .A1(n8860), .A2(n8731), .ZN(n9018) );
  NAND2_X1 U9274 ( .A1(n9274), .A2(n9275), .ZN(n9017) );
  NAND2_X1 U9275 ( .A1(n9276), .A2(b_29_), .ZN(n9275) );
  NOR2_X1 U9276 ( .A1(n9277), .A2(n8736), .ZN(n9276) );
  NOR2_X1 U9277 ( .A1(n9023), .A2(n9024), .ZN(n9277) );
  NAND2_X1 U9278 ( .A1(n9023), .A2(n9024), .ZN(n9274) );
  NAND2_X1 U9279 ( .A1(n9201), .A2(n9278), .ZN(n9024) );
  NAND2_X1 U9280 ( .A1(n9200), .A2(n9202), .ZN(n9278) );
  NAND2_X1 U9281 ( .A1(n9279), .A2(n9280), .ZN(n9202) );
  NAND2_X1 U9282 ( .A1(b_29_), .A2(a_10_), .ZN(n9280) );
  INV_X1 U9283 ( .A(n9281), .ZN(n9279) );
  XOR2_X1 U9284 ( .A(n9282), .B(n9283), .Z(n9200) );
  XOR2_X1 U9285 ( .A(n9284), .B(n9285), .Z(n9282) );
  NOR2_X1 U9286 ( .A1(n8452), .A2(n9168), .ZN(n9285) );
  NAND2_X1 U9287 ( .A1(a_10_), .A2(n9281), .ZN(n9201) );
  NAND2_X1 U9288 ( .A1(n9286), .A2(n9287), .ZN(n9281) );
  NAND2_X1 U9289 ( .A1(n9288), .A2(b_29_), .ZN(n9287) );
  NOR2_X1 U9290 ( .A1(n9289), .A2(n8452), .ZN(n9288) );
  NOR2_X1 U9291 ( .A1(n9035), .A2(n9036), .ZN(n9289) );
  NAND2_X1 U9292 ( .A1(n9035), .A2(n9036), .ZN(n9286) );
  NAND2_X1 U9293 ( .A1(n9197), .A2(n9290), .ZN(n9036) );
  NAND2_X1 U9294 ( .A1(n9196), .A2(n9198), .ZN(n9290) );
  NAND2_X1 U9295 ( .A1(n9291), .A2(n9292), .ZN(n9198) );
  NAND2_X1 U9296 ( .A1(b_29_), .A2(a_12_), .ZN(n9292) );
  INV_X1 U9297 ( .A(n9293), .ZN(n9291) );
  XNOR2_X1 U9298 ( .A(n9294), .B(n9295), .ZN(n9196) );
  NAND2_X1 U9299 ( .A1(n9296), .A2(n9297), .ZN(n9294) );
  NAND2_X1 U9300 ( .A1(a_12_), .A2(n9293), .ZN(n9197) );
  NAND2_X1 U9301 ( .A1(n9049), .A2(n9298), .ZN(n9293) );
  NAND2_X1 U9302 ( .A1(n9048), .A2(n9050), .ZN(n9298) );
  NAND2_X1 U9303 ( .A1(n9299), .A2(n9300), .ZN(n9050) );
  NAND2_X1 U9304 ( .A1(b_29_), .A2(a_13_), .ZN(n9300) );
  INV_X1 U9305 ( .A(n9301), .ZN(n9299) );
  XNOR2_X1 U9306 ( .A(n9302), .B(n9303), .ZN(n9048) );
  NAND2_X1 U9307 ( .A1(n9304), .A2(n9305), .ZN(n9302) );
  NAND2_X1 U9308 ( .A1(a_13_), .A2(n9301), .ZN(n9049) );
  NAND2_X1 U9309 ( .A1(n9057), .A2(n9306), .ZN(n9301) );
  NAND2_X1 U9310 ( .A1(n9056), .A2(n9058), .ZN(n9306) );
  NAND2_X1 U9311 ( .A1(n9307), .A2(n9308), .ZN(n9058) );
  NAND2_X1 U9312 ( .A1(b_29_), .A2(a_14_), .ZN(n9308) );
  INV_X1 U9313 ( .A(n9309), .ZN(n9307) );
  XOR2_X1 U9314 ( .A(n9310), .B(n9311), .Z(n9056) );
  XOR2_X1 U9315 ( .A(n9312), .B(n9313), .Z(n9310) );
  NOR2_X1 U9316 ( .A1(n8763), .A2(n9168), .ZN(n9313) );
  NAND2_X1 U9317 ( .A1(a_14_), .A2(n9309), .ZN(n9057) );
  NAND2_X1 U9318 ( .A1(n9314), .A2(n9315), .ZN(n9309) );
  NAND2_X1 U9319 ( .A1(n9316), .A2(b_29_), .ZN(n9315) );
  NOR2_X1 U9320 ( .A1(n9317), .A2(n8763), .ZN(n9316) );
  NOR2_X1 U9321 ( .A1(n9064), .A2(n9065), .ZN(n9317) );
  NAND2_X1 U9322 ( .A1(n9064), .A2(n9065), .ZN(n9314) );
  NAND2_X1 U9323 ( .A1(n9193), .A2(n9318), .ZN(n9065) );
  NAND2_X1 U9324 ( .A1(n9192), .A2(n9194), .ZN(n9318) );
  NAND2_X1 U9325 ( .A1(n9319), .A2(n9320), .ZN(n9194) );
  NAND2_X1 U9326 ( .A1(b_29_), .A2(a_16_), .ZN(n9320) );
  INV_X1 U9327 ( .A(n9321), .ZN(n9319) );
  XNOR2_X1 U9328 ( .A(n9322), .B(n9323), .ZN(n9192) );
  NAND2_X1 U9329 ( .A1(n9324), .A2(n9325), .ZN(n9322) );
  NAND2_X1 U9330 ( .A1(a_16_), .A2(n9321), .ZN(n9193) );
  NAND2_X1 U9331 ( .A1(n9077), .A2(n9326), .ZN(n9321) );
  NAND2_X1 U9332 ( .A1(n9076), .A2(n9078), .ZN(n9326) );
  NAND2_X1 U9333 ( .A1(n9327), .A2(n9328), .ZN(n9078) );
  NAND2_X1 U9334 ( .A1(b_29_), .A2(a_17_), .ZN(n9328) );
  INV_X1 U9335 ( .A(n9329), .ZN(n9327) );
  XNOR2_X1 U9336 ( .A(n9330), .B(n9331), .ZN(n9076) );
  NAND2_X1 U9337 ( .A1(n9332), .A2(n9333), .ZN(n9330) );
  NAND2_X1 U9338 ( .A1(a_17_), .A2(n9329), .ZN(n9077) );
  NAND2_X1 U9339 ( .A1(n9085), .A2(n9334), .ZN(n9329) );
  NAND2_X1 U9340 ( .A1(n9084), .A2(n9086), .ZN(n9334) );
  NAND2_X1 U9341 ( .A1(n9335), .A2(n9336), .ZN(n9086) );
  NAND2_X1 U9342 ( .A1(b_29_), .A2(a_18_), .ZN(n9336) );
  INV_X1 U9343 ( .A(n9337), .ZN(n9335) );
  XNOR2_X1 U9344 ( .A(n9338), .B(n9339), .ZN(n9084) );
  XOR2_X1 U9345 ( .A(n9340), .B(n9341), .Z(n9339) );
  NAND2_X1 U9346 ( .A1(b_28_), .A2(a_19_), .ZN(n9341) );
  NAND2_X1 U9347 ( .A1(a_18_), .A2(n9337), .ZN(n9085) );
  NAND2_X1 U9348 ( .A1(n9342), .A2(n9343), .ZN(n9337) );
  NAND2_X1 U9349 ( .A1(n9344), .A2(b_29_), .ZN(n9343) );
  NOR2_X1 U9350 ( .A1(n9345), .A2(n8881), .ZN(n9344) );
  NOR2_X1 U9351 ( .A1(n9092), .A2(n9093), .ZN(n9345) );
  NAND2_X1 U9352 ( .A1(n9092), .A2(n9093), .ZN(n9342) );
  NAND2_X1 U9353 ( .A1(n9189), .A2(n9346), .ZN(n9093) );
  NAND2_X1 U9354 ( .A1(n9188), .A2(n9190), .ZN(n9346) );
  NAND2_X1 U9355 ( .A1(n9347), .A2(n9348), .ZN(n9190) );
  NAND2_X1 U9356 ( .A1(b_29_), .A2(a_20_), .ZN(n9348) );
  INV_X1 U9357 ( .A(n9349), .ZN(n9347) );
  XNOR2_X1 U9358 ( .A(n9350), .B(n9351), .ZN(n9188) );
  NAND2_X1 U9359 ( .A1(n9352), .A2(n9353), .ZN(n9350) );
  NAND2_X1 U9360 ( .A1(a_20_), .A2(n9349), .ZN(n9189) );
  NAND2_X1 U9361 ( .A1(n9105), .A2(n9354), .ZN(n9349) );
  NAND2_X1 U9362 ( .A1(n9104), .A2(n9106), .ZN(n9354) );
  NAND2_X1 U9363 ( .A1(n9355), .A2(n9356), .ZN(n9106) );
  NAND2_X1 U9364 ( .A1(b_29_), .A2(a_21_), .ZN(n9356) );
  INV_X1 U9365 ( .A(n9357), .ZN(n9355) );
  XNOR2_X1 U9366 ( .A(n9358), .B(n9359), .ZN(n9104) );
  NAND2_X1 U9367 ( .A1(n9360), .A2(n9361), .ZN(n9358) );
  NAND2_X1 U9368 ( .A1(a_21_), .A2(n9357), .ZN(n9105) );
  NAND2_X1 U9369 ( .A1(n9113), .A2(n9362), .ZN(n9357) );
  NAND2_X1 U9370 ( .A1(n9112), .A2(n9114), .ZN(n9362) );
  NAND2_X1 U9371 ( .A1(n9363), .A2(n9364), .ZN(n9114) );
  NAND2_X1 U9372 ( .A1(b_29_), .A2(a_22_), .ZN(n9364) );
  INV_X1 U9373 ( .A(n9365), .ZN(n9363) );
  XOR2_X1 U9374 ( .A(n9366), .B(n9367), .Z(n9112) );
  XNOR2_X1 U9375 ( .A(n9368), .B(n9369), .ZN(n9366) );
  NAND2_X1 U9376 ( .A1(b_28_), .A2(a_23_), .ZN(n9368) );
  NAND2_X1 U9377 ( .A1(a_22_), .A2(n9365), .ZN(n9113) );
  NAND2_X1 U9378 ( .A1(n9370), .A2(n9371), .ZN(n9365) );
  NAND2_X1 U9379 ( .A1(n9372), .A2(b_29_), .ZN(n9371) );
  NOR2_X1 U9380 ( .A1(n9373), .A2(n8812), .ZN(n9372) );
  NOR2_X1 U9381 ( .A1(n9119), .A2(n9121), .ZN(n9373) );
  NAND2_X1 U9382 ( .A1(n9119), .A2(n9121), .ZN(n9370) );
  NAND2_X1 U9383 ( .A1(n9374), .A2(n9375), .ZN(n9121) );
  NAND2_X1 U9384 ( .A1(n9376), .A2(b_29_), .ZN(n9375) );
  NOR2_X1 U9385 ( .A1(n9377), .A2(n9131), .ZN(n9376) );
  NOR2_X1 U9386 ( .A1(n9184), .A2(n9185), .ZN(n9377) );
  NAND2_X1 U9387 ( .A1(n9184), .A2(n9185), .ZN(n9374) );
  NAND2_X1 U9388 ( .A1(n9378), .A2(n9379), .ZN(n9185) );
  NAND2_X1 U9389 ( .A1(n9182), .A2(n9380), .ZN(n9379) );
  INV_X1 U9390 ( .A(n9381), .ZN(n9380) );
  NOR2_X1 U9391 ( .A1(n9180), .A2(n9181), .ZN(n9381) );
  NOR2_X1 U9392 ( .A1(n8860), .A2(n8825), .ZN(n9182) );
  NAND2_X1 U9393 ( .A1(n9181), .A2(n9180), .ZN(n9378) );
  XOR2_X1 U9394 ( .A(n9382), .B(n9383), .Z(n9180) );
  XNOR2_X1 U9395 ( .A(n9384), .B(n9385), .ZN(n9383) );
  NOR2_X1 U9396 ( .A1(n9386), .A2(n9387), .ZN(n9181) );
  INV_X1 U9397 ( .A(n9388), .ZN(n9387) );
  NAND2_X1 U9398 ( .A1(n9175), .A2(n9389), .ZN(n9388) );
  NAND2_X1 U9399 ( .A1(n9178), .A2(n9177), .ZN(n9389) );
  XOR2_X1 U9400 ( .A(n9390), .B(n9391), .Z(n9175) );
  XNOR2_X1 U9401 ( .A(n9392), .B(n9393), .ZN(n9390) );
  NOR2_X1 U9402 ( .A1(n9177), .A2(n9178), .ZN(n9386) );
  NOR2_X1 U9403 ( .A1(n8860), .A2(n8830), .ZN(n9178) );
  NAND2_X1 U9404 ( .A1(n9142), .A2(n9394), .ZN(n9177) );
  NAND2_X1 U9405 ( .A1(n9141), .A2(n9143), .ZN(n9394) );
  NAND2_X1 U9406 ( .A1(n9395), .A2(n9396), .ZN(n9143) );
  NAND2_X1 U9407 ( .A1(b_29_), .A2(a_27_), .ZN(n9396) );
  INV_X1 U9408 ( .A(n9397), .ZN(n9395) );
  XNOR2_X1 U9409 ( .A(n9398), .B(n9399), .ZN(n9141) );
  XNOR2_X1 U9410 ( .A(n9400), .B(n9401), .ZN(n9398) );
  NAND2_X1 U9411 ( .A1(a_27_), .A2(n9397), .ZN(n9142) );
  NAND2_X1 U9412 ( .A1(n9402), .A2(n9403), .ZN(n9397) );
  NAND2_X1 U9413 ( .A1(n9404), .A2(b_29_), .ZN(n9403) );
  NOR2_X1 U9414 ( .A1(n9405), .A2(n8844), .ZN(n9404) );
  NOR2_X1 U9415 ( .A1(n9149), .A2(n9148), .ZN(n9405) );
  NAND2_X1 U9416 ( .A1(n9149), .A2(n9148), .ZN(n9402) );
  XNOR2_X1 U9417 ( .A(n9406), .B(n9407), .ZN(n9148) );
  XOR2_X1 U9418 ( .A(n9408), .B(n9409), .Z(n9407) );
  NOR2_X1 U9419 ( .A1(n9410), .A2(n9411), .ZN(n9149) );
  INV_X1 U9420 ( .A(n9412), .ZN(n9411) );
  NAND2_X1 U9421 ( .A1(n9413), .A2(n9173), .ZN(n9412) );
  NAND2_X1 U9422 ( .A1(n9414), .A2(b_29_), .ZN(n9173) );
  NOR2_X1 U9423 ( .A1(n9170), .A2(n9168), .ZN(n9414) );
  NAND2_X1 U9424 ( .A1(n9171), .A2(n9174), .ZN(n9413) );
  NOR2_X1 U9425 ( .A1(n9174), .A2(n9171), .ZN(n9410) );
  NAND2_X1 U9426 ( .A1(n9415), .A2(n9416), .ZN(n9174) );
  NAND2_X1 U9427 ( .A1(b_27_), .A2(n9417), .ZN(n9416) );
  NAND2_X1 U9428 ( .A1(n8358), .A2(n9418), .ZN(n9417) );
  NAND2_X1 U9429 ( .A1(a_31_), .A2(n9168), .ZN(n9418) );
  NAND2_X1 U9430 ( .A1(b_28_), .A2(n9419), .ZN(n9415) );
  NAND2_X1 U9431 ( .A1(n8362), .A2(n9420), .ZN(n9419) );
  NAND2_X1 U9432 ( .A1(a_30_), .A2(n9421), .ZN(n9420) );
  XOR2_X1 U9433 ( .A(n9422), .B(n9423), .Z(n9184) );
  XOR2_X1 U9434 ( .A(n9424), .B(n9425), .Z(n9423) );
  XNOR2_X1 U9435 ( .A(n9426), .B(n9427), .ZN(n9119) );
  XOR2_X1 U9436 ( .A(n9428), .B(n9429), .Z(n9427) );
  XNOR2_X1 U9437 ( .A(n9430), .B(n9431), .ZN(n9092) );
  NAND2_X1 U9438 ( .A1(n9432), .A2(n9433), .ZN(n9430) );
  XNOR2_X1 U9439 ( .A(n9434), .B(n9435), .ZN(n9064) );
  NAND2_X1 U9440 ( .A1(n9436), .A2(n9437), .ZN(n9434) );
  XNOR2_X1 U9441 ( .A(n9438), .B(n9439), .ZN(n9035) );
  NAND2_X1 U9442 ( .A1(n9440), .A2(n9441), .ZN(n9438) );
  XOR2_X1 U9443 ( .A(n9442), .B(n9443), .Z(n9023) );
  XNOR2_X1 U9444 ( .A(n9444), .B(n9445), .ZN(n9443) );
  NAND2_X1 U9445 ( .A1(n9206), .A2(n9204), .ZN(n9222) );
  XNOR2_X1 U9446 ( .A(n9446), .B(n9447), .ZN(n9204) );
  XOR2_X1 U9447 ( .A(n9448), .B(n9449), .Z(n9447) );
  NAND2_X1 U9448 ( .A1(b_28_), .A2(a_3_), .ZN(n9449) );
  NOR2_X1 U9449 ( .A1(n8860), .A2(n8497), .ZN(n9206) );
  XOR2_X1 U9450 ( .A(n9450), .B(n9451), .Z(n9208) );
  NAND2_X1 U9451 ( .A1(n9452), .A2(n9453), .ZN(n9450) );
  XOR2_X1 U9452 ( .A(n9454), .B(n9455), .Z(n8956) );
  XOR2_X1 U9453 ( .A(n9456), .B(n9457), .Z(n9454) );
  XOR2_X1 U9454 ( .A(n9458), .B(n9459), .Z(n8961) );
  XNOR2_X1 U9455 ( .A(n9460), .B(n9461), .ZN(n9459) );
  INV_X1 U9456 ( .A(n9462), .ZN(n8525) );
  NOR2_X1 U9457 ( .A1(n8672), .A2(n8673), .ZN(n9462) );
  NAND2_X1 U9458 ( .A1(n9463), .A2(n8668), .ZN(n8673) );
  NAND2_X1 U9459 ( .A1(n9464), .A2(n9465), .ZN(n9463) );
  XOR2_X1 U9460 ( .A(n9466), .B(n9467), .Z(n9465) );
  INV_X1 U9461 ( .A(n9468), .ZN(n9464) );
  NAND2_X1 U9462 ( .A1(n8679), .A2(n9212), .ZN(n8672) );
  INV_X1 U9463 ( .A(n8678), .ZN(n9212) );
  NOR2_X1 U9464 ( .A1(n9469), .A2(n9470), .ZN(n8678) );
  INV_X1 U9465 ( .A(n9471), .ZN(n9470) );
  NAND2_X1 U9466 ( .A1(n9461), .A2(n9472), .ZN(n9471) );
  NAND2_X1 U9467 ( .A1(n9458), .A2(n9460), .ZN(n9472) );
  NOR2_X1 U9468 ( .A1(n9168), .A2(n8690), .ZN(n9461) );
  NOR2_X1 U9469 ( .A1(n9460), .A2(n9458), .ZN(n9469) );
  XNOR2_X1 U9470 ( .A(n9473), .B(n9474), .ZN(n9458) );
  XOR2_X1 U9471 ( .A(n9475), .B(n9476), .Z(n9473) );
  NOR2_X1 U9472 ( .A1(n8502), .A2(n9421), .ZN(n9476) );
  NAND2_X1 U9473 ( .A1(n9477), .A2(n9478), .ZN(n9460) );
  NAND2_X1 U9474 ( .A1(n9455), .A2(n9479), .ZN(n9478) );
  NAND2_X1 U9475 ( .A1(n9457), .A2(n9456), .ZN(n9479) );
  XOR2_X1 U9476 ( .A(n9480), .B(n9481), .Z(n9455) );
  NAND2_X1 U9477 ( .A1(n9482), .A2(n9483), .ZN(n9480) );
  INV_X1 U9478 ( .A(n9484), .ZN(n9477) );
  NOR2_X1 U9479 ( .A1(n9456), .A2(n9457), .ZN(n9484) );
  NOR2_X1 U9480 ( .A1(n9168), .A2(n8502), .ZN(n9457) );
  NAND2_X1 U9481 ( .A1(n9452), .A2(n9485), .ZN(n9456) );
  NAND2_X1 U9482 ( .A1(n9451), .A2(n9453), .ZN(n9485) );
  NAND2_X1 U9483 ( .A1(n9486), .A2(n9487), .ZN(n9453) );
  NAND2_X1 U9484 ( .A1(b_28_), .A2(a_2_), .ZN(n9487) );
  INV_X1 U9485 ( .A(n9488), .ZN(n9486) );
  XNOR2_X1 U9486 ( .A(n9489), .B(n9490), .ZN(n9451) );
  NAND2_X1 U9487 ( .A1(n9491), .A2(n9492), .ZN(n9489) );
  NAND2_X1 U9488 ( .A1(a_2_), .A2(n9488), .ZN(n9452) );
  NAND2_X1 U9489 ( .A1(n9493), .A2(n9494), .ZN(n9488) );
  NAND2_X1 U9490 ( .A1(n9495), .A2(b_28_), .ZN(n9494) );
  NOR2_X1 U9491 ( .A1(n9496), .A2(n8707), .ZN(n9495) );
  NOR2_X1 U9492 ( .A1(n9446), .A2(n9448), .ZN(n9496) );
  NAND2_X1 U9493 ( .A1(n9446), .A2(n9448), .ZN(n9493) );
  NAND2_X1 U9494 ( .A1(n9497), .A2(n9498), .ZN(n9448) );
  NAND2_X1 U9495 ( .A1(n9499), .A2(b_28_), .ZN(n9498) );
  NOR2_X1 U9496 ( .A1(n9500), .A2(n8712), .ZN(n9499) );
  NOR2_X1 U9497 ( .A1(n9230), .A2(n9232), .ZN(n9500) );
  NAND2_X1 U9498 ( .A1(n9230), .A2(n9232), .ZN(n9497) );
  NAND2_X1 U9499 ( .A1(n9501), .A2(n9502), .ZN(n9232) );
  NAND2_X1 U9500 ( .A1(n9503), .A2(b_28_), .ZN(n9502) );
  NOR2_X1 U9501 ( .A1(n9504), .A2(n8717), .ZN(n9503) );
  NOR2_X1 U9502 ( .A1(n9240), .A2(n9239), .ZN(n9504) );
  NAND2_X1 U9503 ( .A1(n9240), .A2(n9239), .ZN(n9501) );
  XOR2_X1 U9504 ( .A(n9505), .B(n9506), .Z(n9239) );
  XOR2_X1 U9505 ( .A(n9507), .B(n9508), .Z(n9505) );
  NOR2_X1 U9506 ( .A1(n8480), .A2(n9421), .ZN(n9508) );
  NOR2_X1 U9507 ( .A1(n9509), .A2(n9510), .ZN(n9240) );
  INV_X1 U9508 ( .A(n9511), .ZN(n9510) );
  NAND2_X1 U9509 ( .A1(n9246), .A2(n9512), .ZN(n9511) );
  NAND2_X1 U9510 ( .A1(n9249), .A2(n9248), .ZN(n9512) );
  XOR2_X1 U9511 ( .A(n9513), .B(n9514), .Z(n9246) );
  NAND2_X1 U9512 ( .A1(n9515), .A2(n9516), .ZN(n9513) );
  NOR2_X1 U9513 ( .A1(n9248), .A2(n9249), .ZN(n9509) );
  NOR2_X1 U9514 ( .A1(n9168), .A2(n8480), .ZN(n9249) );
  NAND2_X1 U9515 ( .A1(n9256), .A2(n9517), .ZN(n9248) );
  NAND2_X1 U9516 ( .A1(n9255), .A2(n9257), .ZN(n9517) );
  NAND2_X1 U9517 ( .A1(n9518), .A2(n9519), .ZN(n9257) );
  NAND2_X1 U9518 ( .A1(b_28_), .A2(a_7_), .ZN(n9519) );
  INV_X1 U9519 ( .A(n9520), .ZN(n9518) );
  XNOR2_X1 U9520 ( .A(n9521), .B(n9522), .ZN(n9255) );
  NAND2_X1 U9521 ( .A1(n9523), .A2(n9524), .ZN(n9521) );
  NAND2_X1 U9522 ( .A1(a_7_), .A2(n9520), .ZN(n9256) );
  NAND2_X1 U9523 ( .A1(n9264), .A2(n9525), .ZN(n9520) );
  NAND2_X1 U9524 ( .A1(n9263), .A2(n9265), .ZN(n9525) );
  NAND2_X1 U9525 ( .A1(n9526), .A2(n9527), .ZN(n9265) );
  NAND2_X1 U9526 ( .A1(b_28_), .A2(a_8_), .ZN(n9527) );
  INV_X1 U9527 ( .A(n9528), .ZN(n9526) );
  XNOR2_X1 U9528 ( .A(n9529), .B(n9530), .ZN(n9263) );
  XNOR2_X1 U9529 ( .A(n9531), .B(n9532), .ZN(n9529) );
  NOR2_X1 U9530 ( .A1(n8736), .A2(n9421), .ZN(n9532) );
  NAND2_X1 U9531 ( .A1(a_8_), .A2(n9528), .ZN(n9264) );
  NAND2_X1 U9532 ( .A1(n9272), .A2(n9533), .ZN(n9528) );
  NAND2_X1 U9533 ( .A1(n9271), .A2(n9273), .ZN(n9533) );
  NAND2_X1 U9534 ( .A1(n9534), .A2(n9535), .ZN(n9273) );
  INV_X1 U9535 ( .A(n9536), .ZN(n9535) );
  NAND2_X1 U9536 ( .A1(b_28_), .A2(a_9_), .ZN(n9534) );
  XOR2_X1 U9537 ( .A(n9537), .B(n9538), .Z(n9271) );
  XNOR2_X1 U9538 ( .A(n9539), .B(n9540), .ZN(n9538) );
  NAND2_X1 U9539 ( .A1(n9536), .A2(a_9_), .ZN(n9272) );
  NOR2_X1 U9540 ( .A1(n9541), .A2(n9542), .ZN(n9536) );
  INV_X1 U9541 ( .A(n9543), .ZN(n9542) );
  NAND2_X1 U9542 ( .A1(n9442), .A2(n9544), .ZN(n9543) );
  NAND2_X1 U9543 ( .A1(n9445), .A2(n9444), .ZN(n9544) );
  XOR2_X1 U9544 ( .A(n9545), .B(n9546), .Z(n9442) );
  NAND2_X1 U9545 ( .A1(n9547), .A2(n9548), .ZN(n9545) );
  NOR2_X1 U9546 ( .A1(n9444), .A2(n9445), .ZN(n9541) );
  NOR2_X1 U9547 ( .A1(n9168), .A2(n8741), .ZN(n9445) );
  NAND2_X1 U9548 ( .A1(n9549), .A2(n9550), .ZN(n9444) );
  NAND2_X1 U9549 ( .A1(n9551), .A2(b_28_), .ZN(n9550) );
  NOR2_X1 U9550 ( .A1(n9552), .A2(n8452), .ZN(n9551) );
  NOR2_X1 U9551 ( .A1(n9283), .A2(n9284), .ZN(n9552) );
  NAND2_X1 U9552 ( .A1(n9283), .A2(n9284), .ZN(n9549) );
  NAND2_X1 U9553 ( .A1(n9440), .A2(n9553), .ZN(n9284) );
  NAND2_X1 U9554 ( .A1(n9439), .A2(n9441), .ZN(n9553) );
  NAND2_X1 U9555 ( .A1(n9554), .A2(n9555), .ZN(n9441) );
  NAND2_X1 U9556 ( .A1(b_28_), .A2(a_12_), .ZN(n9555) );
  INV_X1 U9557 ( .A(n9556), .ZN(n9554) );
  XNOR2_X1 U9558 ( .A(n9557), .B(n9558), .ZN(n9439) );
  NAND2_X1 U9559 ( .A1(n9559), .A2(n9560), .ZN(n9557) );
  NAND2_X1 U9560 ( .A1(a_12_), .A2(n9556), .ZN(n9440) );
  NAND2_X1 U9561 ( .A1(n9296), .A2(n9561), .ZN(n9556) );
  NAND2_X1 U9562 ( .A1(n9295), .A2(n9297), .ZN(n9561) );
  NAND2_X1 U9563 ( .A1(n9562), .A2(n9563), .ZN(n9297) );
  NAND2_X1 U9564 ( .A1(b_28_), .A2(a_13_), .ZN(n9563) );
  INV_X1 U9565 ( .A(n9564), .ZN(n9562) );
  XNOR2_X1 U9566 ( .A(n9565), .B(n9566), .ZN(n9295) );
  NAND2_X1 U9567 ( .A1(n9567), .A2(n9568), .ZN(n9565) );
  NAND2_X1 U9568 ( .A1(a_13_), .A2(n9564), .ZN(n9296) );
  NAND2_X1 U9569 ( .A1(n9304), .A2(n9569), .ZN(n9564) );
  NAND2_X1 U9570 ( .A1(n9303), .A2(n9305), .ZN(n9569) );
  NAND2_X1 U9571 ( .A1(n9570), .A2(n9571), .ZN(n9305) );
  NAND2_X1 U9572 ( .A1(b_28_), .A2(a_14_), .ZN(n9571) );
  INV_X1 U9573 ( .A(n9572), .ZN(n9570) );
  XOR2_X1 U9574 ( .A(n9573), .B(n9574), .Z(n9303) );
  XOR2_X1 U9575 ( .A(n9575), .B(n9576), .Z(n9573) );
  NOR2_X1 U9576 ( .A1(n8763), .A2(n9421), .ZN(n9576) );
  NAND2_X1 U9577 ( .A1(a_14_), .A2(n9572), .ZN(n9304) );
  NAND2_X1 U9578 ( .A1(n9577), .A2(n9578), .ZN(n9572) );
  NAND2_X1 U9579 ( .A1(n9579), .A2(b_28_), .ZN(n9578) );
  NOR2_X1 U9580 ( .A1(n9580), .A2(n8763), .ZN(n9579) );
  NOR2_X1 U9581 ( .A1(n9311), .A2(n9312), .ZN(n9580) );
  NAND2_X1 U9582 ( .A1(n9311), .A2(n9312), .ZN(n9577) );
  NAND2_X1 U9583 ( .A1(n9436), .A2(n9581), .ZN(n9312) );
  NAND2_X1 U9584 ( .A1(n9435), .A2(n9437), .ZN(n9581) );
  NAND2_X1 U9585 ( .A1(n9582), .A2(n9583), .ZN(n9437) );
  NAND2_X1 U9586 ( .A1(b_28_), .A2(a_16_), .ZN(n9583) );
  INV_X1 U9587 ( .A(n9584), .ZN(n9582) );
  XNOR2_X1 U9588 ( .A(n9585), .B(n9586), .ZN(n9435) );
  NAND2_X1 U9589 ( .A1(n9587), .A2(n9588), .ZN(n9585) );
  NAND2_X1 U9590 ( .A1(a_16_), .A2(n9584), .ZN(n9436) );
  NAND2_X1 U9591 ( .A1(n9324), .A2(n9589), .ZN(n9584) );
  NAND2_X1 U9592 ( .A1(n9323), .A2(n9325), .ZN(n9589) );
  NAND2_X1 U9593 ( .A1(n9590), .A2(n9591), .ZN(n9325) );
  NAND2_X1 U9594 ( .A1(b_28_), .A2(a_17_), .ZN(n9591) );
  INV_X1 U9595 ( .A(n9592), .ZN(n9590) );
  XNOR2_X1 U9596 ( .A(n9593), .B(n9594), .ZN(n9323) );
  NAND2_X1 U9597 ( .A1(n9595), .A2(n9596), .ZN(n9593) );
  NAND2_X1 U9598 ( .A1(a_17_), .A2(n9592), .ZN(n9324) );
  NAND2_X1 U9599 ( .A1(n9332), .A2(n9597), .ZN(n9592) );
  NAND2_X1 U9600 ( .A1(n9331), .A2(n9333), .ZN(n9597) );
  NAND2_X1 U9601 ( .A1(n9598), .A2(n9599), .ZN(n9333) );
  NAND2_X1 U9602 ( .A1(b_28_), .A2(a_18_), .ZN(n9599) );
  INV_X1 U9603 ( .A(n9600), .ZN(n9598) );
  XOR2_X1 U9604 ( .A(n9601), .B(n9602), .Z(n9331) );
  XOR2_X1 U9605 ( .A(n9603), .B(n9604), .Z(n9601) );
  NOR2_X1 U9606 ( .A1(n8881), .A2(n9421), .ZN(n9604) );
  NAND2_X1 U9607 ( .A1(a_18_), .A2(n9600), .ZN(n9332) );
  NAND2_X1 U9608 ( .A1(n9605), .A2(n9606), .ZN(n9600) );
  NAND2_X1 U9609 ( .A1(n9607), .A2(b_28_), .ZN(n9606) );
  NOR2_X1 U9610 ( .A1(n9608), .A2(n8881), .ZN(n9607) );
  NOR2_X1 U9611 ( .A1(n9338), .A2(n9340), .ZN(n9608) );
  NAND2_X1 U9612 ( .A1(n9338), .A2(n9340), .ZN(n9605) );
  NAND2_X1 U9613 ( .A1(n9432), .A2(n9609), .ZN(n9340) );
  NAND2_X1 U9614 ( .A1(n9431), .A2(n9433), .ZN(n9609) );
  NAND2_X1 U9615 ( .A1(n9610), .A2(n9611), .ZN(n9433) );
  NAND2_X1 U9616 ( .A1(b_28_), .A2(a_20_), .ZN(n9611) );
  INV_X1 U9617 ( .A(n9612), .ZN(n9610) );
  XNOR2_X1 U9618 ( .A(n9613), .B(n9614), .ZN(n9431) );
  NAND2_X1 U9619 ( .A1(n9615), .A2(n9616), .ZN(n9613) );
  NAND2_X1 U9620 ( .A1(a_20_), .A2(n9612), .ZN(n9432) );
  NAND2_X1 U9621 ( .A1(n9352), .A2(n9617), .ZN(n9612) );
  NAND2_X1 U9622 ( .A1(n9351), .A2(n9353), .ZN(n9617) );
  NAND2_X1 U9623 ( .A1(n9618), .A2(n9619), .ZN(n9353) );
  NAND2_X1 U9624 ( .A1(b_28_), .A2(a_21_), .ZN(n9619) );
  INV_X1 U9625 ( .A(n9620), .ZN(n9618) );
  XNOR2_X1 U9626 ( .A(n9621), .B(n9622), .ZN(n9351) );
  NAND2_X1 U9627 ( .A1(n9623), .A2(n9624), .ZN(n9621) );
  NAND2_X1 U9628 ( .A1(a_21_), .A2(n9620), .ZN(n9352) );
  NAND2_X1 U9629 ( .A1(n9360), .A2(n9625), .ZN(n9620) );
  NAND2_X1 U9630 ( .A1(n9359), .A2(n9361), .ZN(n9625) );
  NAND2_X1 U9631 ( .A1(n9626), .A2(n9627), .ZN(n9361) );
  NAND2_X1 U9632 ( .A1(b_28_), .A2(a_22_), .ZN(n9627) );
  INV_X1 U9633 ( .A(n9628), .ZN(n9626) );
  XOR2_X1 U9634 ( .A(n9629), .B(n9630), .Z(n9359) );
  XOR2_X1 U9635 ( .A(n9631), .B(n9632), .Z(n9629) );
  NOR2_X1 U9636 ( .A1(n8812), .A2(n9421), .ZN(n9632) );
  NAND2_X1 U9637 ( .A1(a_22_), .A2(n9628), .ZN(n9360) );
  NAND2_X1 U9638 ( .A1(n9633), .A2(n9634), .ZN(n9628) );
  NAND2_X1 U9639 ( .A1(n9635), .A2(b_28_), .ZN(n9634) );
  NOR2_X1 U9640 ( .A1(n9636), .A2(n8812), .ZN(n9635) );
  NOR2_X1 U9641 ( .A1(n9367), .A2(n9369), .ZN(n9636) );
  NAND2_X1 U9642 ( .A1(n9367), .A2(n9369), .ZN(n9633) );
  NAND2_X1 U9643 ( .A1(n9637), .A2(n9638), .ZN(n9369) );
  INV_X1 U9644 ( .A(n9639), .ZN(n9638) );
  NOR2_X1 U9645 ( .A1(n9429), .A2(n9640), .ZN(n9639) );
  NOR2_X1 U9646 ( .A1(n9428), .A2(n9426), .ZN(n9640) );
  NAND2_X1 U9647 ( .A1(b_28_), .A2(a_24_), .ZN(n9429) );
  NAND2_X1 U9648 ( .A1(n9426), .A2(n9428), .ZN(n9637) );
  NAND2_X1 U9649 ( .A1(n9641), .A2(n9642), .ZN(n9428) );
  NAND2_X1 U9650 ( .A1(n9425), .A2(n9643), .ZN(n9642) );
  INV_X1 U9651 ( .A(n9644), .ZN(n9643) );
  NOR2_X1 U9652 ( .A1(n9422), .A2(n9424), .ZN(n9644) );
  NOR2_X1 U9653 ( .A1(n9168), .A2(n8825), .ZN(n9425) );
  NAND2_X1 U9654 ( .A1(n9424), .A2(n9422), .ZN(n9641) );
  XNOR2_X1 U9655 ( .A(n9645), .B(n9646), .ZN(n9422) );
  XOR2_X1 U9656 ( .A(n9647), .B(n9648), .Z(n9645) );
  NOR2_X1 U9657 ( .A1(n9649), .A2(n9650), .ZN(n9424) );
  INV_X1 U9658 ( .A(n9651), .ZN(n9650) );
  NAND2_X1 U9659 ( .A1(n9382), .A2(n9652), .ZN(n9651) );
  NAND2_X1 U9660 ( .A1(n9385), .A2(n9384), .ZN(n9652) );
  XNOR2_X1 U9661 ( .A(n9653), .B(n9654), .ZN(n9382) );
  XOR2_X1 U9662 ( .A(n9655), .B(n9656), .Z(n9654) );
  NOR2_X1 U9663 ( .A1(n9384), .A2(n9385), .ZN(n9649) );
  NOR2_X1 U9664 ( .A1(n9168), .A2(n8830), .ZN(n9385) );
  NAND2_X1 U9665 ( .A1(n9657), .A2(n9658), .ZN(n9384) );
  NAND2_X1 U9666 ( .A1(n9393), .A2(n9659), .ZN(n9658) );
  INV_X1 U9667 ( .A(n9660), .ZN(n9659) );
  NOR2_X1 U9668 ( .A1(n9391), .A2(n9392), .ZN(n9660) );
  NOR2_X1 U9669 ( .A1(n9168), .A2(n8839), .ZN(n9393) );
  NAND2_X1 U9670 ( .A1(n9392), .A2(n9391), .ZN(n9657) );
  XOR2_X1 U9671 ( .A(n9661), .B(n9662), .Z(n9391) );
  XNOR2_X1 U9672 ( .A(n9663), .B(n9664), .ZN(n9661) );
  NAND2_X1 U9673 ( .A1(b_27_), .A2(a_28_), .ZN(n9663) );
  NOR2_X1 U9674 ( .A1(n9665), .A2(n9666), .ZN(n9392) );
  NOR2_X1 U9675 ( .A1(n9667), .A2(n9400), .ZN(n9666) );
  NOR2_X1 U9676 ( .A1(n9399), .A2(n9401), .ZN(n9667) );
  INV_X1 U9677 ( .A(n9668), .ZN(n9665) );
  NAND2_X1 U9678 ( .A1(n9401), .A2(n9399), .ZN(n9668) );
  XOR2_X1 U9679 ( .A(n9669), .B(n9670), .Z(n9399) );
  XNOR2_X1 U9680 ( .A(n9671), .B(n9672), .ZN(n9670) );
  NOR2_X1 U9681 ( .A1(n9673), .A2(n9674), .ZN(n9401) );
  INV_X1 U9682 ( .A(n9675), .ZN(n9674) );
  NAND2_X1 U9683 ( .A1(n9406), .A2(n9676), .ZN(n9675) );
  NAND2_X1 U9684 ( .A1(n9677), .A2(n9408), .ZN(n9676) );
  NOR2_X1 U9685 ( .A1(n9168), .A2(n9161), .ZN(n9406) );
  NOR2_X1 U9686 ( .A1(n9408), .A2(n9677), .ZN(n9673) );
  INV_X1 U9687 ( .A(n9409), .ZN(n9677) );
  NAND2_X1 U9688 ( .A1(n9678), .A2(n9679), .ZN(n9409) );
  NAND2_X1 U9689 ( .A1(b_26_), .A2(n9680), .ZN(n9679) );
  NAND2_X1 U9690 ( .A1(n8358), .A2(n9681), .ZN(n9680) );
  NAND2_X1 U9691 ( .A1(a_31_), .A2(n9421), .ZN(n9681) );
  NAND2_X1 U9692 ( .A1(b_27_), .A2(n9682), .ZN(n9678) );
  NAND2_X1 U9693 ( .A1(n8362), .A2(n9683), .ZN(n9682) );
  NAND2_X1 U9694 ( .A1(a_30_), .A2(n9684), .ZN(n9683) );
  NAND2_X1 U9695 ( .A1(n9685), .A2(b_28_), .ZN(n9408) );
  NOR2_X1 U9696 ( .A1(n9170), .A2(n9421), .ZN(n9685) );
  XNOR2_X1 U9697 ( .A(n9686), .B(n9687), .ZN(n9426) );
  XNOR2_X1 U9698 ( .A(n9688), .B(n9689), .ZN(n9687) );
  XOR2_X1 U9699 ( .A(n9690), .B(n9691), .Z(n9367) );
  XOR2_X1 U9700 ( .A(n9692), .B(n9693), .Z(n9690) );
  XNOR2_X1 U9701 ( .A(n9694), .B(n9695), .ZN(n9338) );
  NAND2_X1 U9702 ( .A1(n9696), .A2(n9697), .ZN(n9694) );
  XNOR2_X1 U9703 ( .A(n9698), .B(n9699), .ZN(n9311) );
  NAND2_X1 U9704 ( .A1(n9700), .A2(n9701), .ZN(n9698) );
  XOR2_X1 U9705 ( .A(n9702), .B(n9703), .Z(n9283) );
  XNOR2_X1 U9706 ( .A(n9704), .B(n9705), .ZN(n9703) );
  XOR2_X1 U9707 ( .A(n9706), .B(n9707), .Z(n9230) );
  XOR2_X1 U9708 ( .A(n9708), .B(n9709), .Z(n9706) );
  NOR2_X1 U9709 ( .A1(n8717), .A2(n9421), .ZN(n9709) );
  XNOR2_X1 U9710 ( .A(n9710), .B(n9711), .ZN(n9446) );
  XOR2_X1 U9711 ( .A(n9712), .B(n9713), .Z(n9711) );
  NAND2_X1 U9712 ( .A1(b_27_), .A2(a_4_), .ZN(n9713) );
  XNOR2_X1 U9713 ( .A(n9714), .B(n9715), .ZN(n8679) );
  XOR2_X1 U9714 ( .A(n9716), .B(n9717), .Z(n9715) );
  NAND2_X1 U9715 ( .A1(b_27_), .A2(a_0_), .ZN(n9717) );
  INV_X1 U9716 ( .A(n9718), .ZN(n8530) );
  NOR2_X1 U9717 ( .A1(n9719), .A2(n8668), .ZN(n9718) );
  NAND2_X1 U9718 ( .A1(n9720), .A2(n9468), .ZN(n8668) );
  NAND2_X1 U9719 ( .A1(n9721), .A2(n9722), .ZN(n9468) );
  NAND2_X1 U9720 ( .A1(n9723), .A2(b_27_), .ZN(n9722) );
  NOR2_X1 U9721 ( .A1(n9724), .A2(n8690), .ZN(n9723) );
  NOR2_X1 U9722 ( .A1(n9714), .A2(n9716), .ZN(n9724) );
  NAND2_X1 U9723 ( .A1(n9714), .A2(n9716), .ZN(n9721) );
  NAND2_X1 U9724 ( .A1(n9725), .A2(n9726), .ZN(n9716) );
  NAND2_X1 U9725 ( .A1(n9727), .A2(b_27_), .ZN(n9726) );
  NOR2_X1 U9726 ( .A1(n9728), .A2(n8502), .ZN(n9727) );
  NOR2_X1 U9727 ( .A1(n9474), .A2(n9475), .ZN(n9728) );
  NAND2_X1 U9728 ( .A1(n9474), .A2(n9475), .ZN(n9725) );
  NAND2_X1 U9729 ( .A1(n9482), .A2(n9729), .ZN(n9475) );
  NAND2_X1 U9730 ( .A1(n9481), .A2(n9483), .ZN(n9729) );
  NAND2_X1 U9731 ( .A1(n9730), .A2(n9731), .ZN(n9483) );
  NAND2_X1 U9732 ( .A1(b_27_), .A2(a_2_), .ZN(n9731) );
  INV_X1 U9733 ( .A(n9732), .ZN(n9730) );
  XNOR2_X1 U9734 ( .A(n9733), .B(n9734), .ZN(n9481) );
  XOR2_X1 U9735 ( .A(n9735), .B(n9736), .Z(n9734) );
  NAND2_X1 U9736 ( .A1(a_2_), .A2(n9732), .ZN(n9482) );
  NAND2_X1 U9737 ( .A1(n9491), .A2(n9737), .ZN(n9732) );
  NAND2_X1 U9738 ( .A1(n9490), .A2(n9492), .ZN(n9737) );
  NAND2_X1 U9739 ( .A1(n9738), .A2(n9739), .ZN(n9492) );
  NAND2_X1 U9740 ( .A1(b_27_), .A2(a_3_), .ZN(n9739) );
  INV_X1 U9741 ( .A(n9740), .ZN(n9738) );
  XNOR2_X1 U9742 ( .A(n9741), .B(n9742), .ZN(n9490) );
  XOR2_X1 U9743 ( .A(n9743), .B(n9744), .Z(n9742) );
  NAND2_X1 U9744 ( .A1(b_26_), .A2(a_4_), .ZN(n9744) );
  NAND2_X1 U9745 ( .A1(a_3_), .A2(n9740), .ZN(n9491) );
  NAND2_X1 U9746 ( .A1(n9745), .A2(n9746), .ZN(n9740) );
  NAND2_X1 U9747 ( .A1(n9747), .A2(b_27_), .ZN(n9746) );
  NOR2_X1 U9748 ( .A1(n9748), .A2(n8712), .ZN(n9747) );
  NOR2_X1 U9749 ( .A1(n9710), .A2(n9712), .ZN(n9748) );
  NAND2_X1 U9750 ( .A1(n9710), .A2(n9712), .ZN(n9745) );
  NAND2_X1 U9751 ( .A1(n9749), .A2(n9750), .ZN(n9712) );
  NAND2_X1 U9752 ( .A1(n9751), .A2(b_27_), .ZN(n9750) );
  NOR2_X1 U9753 ( .A1(n9752), .A2(n8717), .ZN(n9751) );
  NOR2_X1 U9754 ( .A1(n9707), .A2(n9708), .ZN(n9752) );
  NAND2_X1 U9755 ( .A1(n9707), .A2(n9708), .ZN(n9749) );
  NAND2_X1 U9756 ( .A1(n9753), .A2(n9754), .ZN(n9708) );
  NAND2_X1 U9757 ( .A1(n9755), .A2(b_27_), .ZN(n9754) );
  NOR2_X1 U9758 ( .A1(n9756), .A2(n8480), .ZN(n9755) );
  NOR2_X1 U9759 ( .A1(n9506), .A2(n9507), .ZN(n9756) );
  NAND2_X1 U9760 ( .A1(n9506), .A2(n9507), .ZN(n9753) );
  NAND2_X1 U9761 ( .A1(n9515), .A2(n9757), .ZN(n9507) );
  NAND2_X1 U9762 ( .A1(n9514), .A2(n9516), .ZN(n9757) );
  NAND2_X1 U9763 ( .A1(n9758), .A2(n9759), .ZN(n9516) );
  NAND2_X1 U9764 ( .A1(b_27_), .A2(a_7_), .ZN(n9759) );
  INV_X1 U9765 ( .A(n9760), .ZN(n9758) );
  XNOR2_X1 U9766 ( .A(n9761), .B(n9762), .ZN(n9514) );
  XOR2_X1 U9767 ( .A(n9763), .B(n9764), .Z(n9762) );
  NAND2_X1 U9768 ( .A1(b_26_), .A2(a_8_), .ZN(n9764) );
  NAND2_X1 U9769 ( .A1(a_7_), .A2(n9760), .ZN(n9515) );
  NAND2_X1 U9770 ( .A1(n9523), .A2(n9765), .ZN(n9760) );
  NAND2_X1 U9771 ( .A1(n9522), .A2(n9524), .ZN(n9765) );
  NAND2_X1 U9772 ( .A1(n9766), .A2(n9767), .ZN(n9524) );
  NAND2_X1 U9773 ( .A1(b_27_), .A2(a_8_), .ZN(n9767) );
  INV_X1 U9774 ( .A(n9768), .ZN(n9766) );
  XNOR2_X1 U9775 ( .A(n9769), .B(n9770), .ZN(n9522) );
  XNOR2_X1 U9776 ( .A(n9771), .B(n9772), .ZN(n9769) );
  NOR2_X1 U9777 ( .A1(n8736), .A2(n9684), .ZN(n9772) );
  NAND2_X1 U9778 ( .A1(a_8_), .A2(n9768), .ZN(n9523) );
  NAND2_X1 U9779 ( .A1(n9773), .A2(n9774), .ZN(n9768) );
  NAND2_X1 U9780 ( .A1(n9775), .A2(b_27_), .ZN(n9774) );
  NOR2_X1 U9781 ( .A1(n9776), .A2(n8736), .ZN(n9775) );
  NOR2_X1 U9782 ( .A1(n9531), .A2(n9530), .ZN(n9776) );
  NAND2_X1 U9783 ( .A1(n9531), .A2(n9530), .ZN(n9773) );
  XOR2_X1 U9784 ( .A(n9777), .B(n9778), .Z(n9530) );
  XNOR2_X1 U9785 ( .A(n9779), .B(n9780), .ZN(n9778) );
  NOR2_X1 U9786 ( .A1(n9781), .A2(n9782), .ZN(n9531) );
  INV_X1 U9787 ( .A(n9783), .ZN(n9782) );
  NAND2_X1 U9788 ( .A1(n9537), .A2(n9784), .ZN(n9783) );
  NAND2_X1 U9789 ( .A1(n9540), .A2(n9539), .ZN(n9784) );
  XOR2_X1 U9790 ( .A(n9785), .B(n9786), .Z(n9537) );
  XNOR2_X1 U9791 ( .A(n9787), .B(n9788), .ZN(n9785) );
  NOR2_X1 U9792 ( .A1(n8452), .A2(n9684), .ZN(n9788) );
  NOR2_X1 U9793 ( .A1(n9539), .A2(n9540), .ZN(n9781) );
  NOR2_X1 U9794 ( .A1(n9421), .A2(n8741), .ZN(n9540) );
  NAND2_X1 U9795 ( .A1(n9547), .A2(n9789), .ZN(n9539) );
  NAND2_X1 U9796 ( .A1(n9546), .A2(n9548), .ZN(n9789) );
  NAND2_X1 U9797 ( .A1(n9790), .A2(n9791), .ZN(n9548) );
  INV_X1 U9798 ( .A(n9792), .ZN(n9791) );
  NAND2_X1 U9799 ( .A1(b_27_), .A2(a_11_), .ZN(n9790) );
  XOR2_X1 U9800 ( .A(n9793), .B(n9794), .Z(n9546) );
  XNOR2_X1 U9801 ( .A(n9795), .B(n9796), .ZN(n9794) );
  NAND2_X1 U9802 ( .A1(n9792), .A2(a_11_), .ZN(n9547) );
  NOR2_X1 U9803 ( .A1(n9797), .A2(n9798), .ZN(n9792) );
  INV_X1 U9804 ( .A(n9799), .ZN(n9798) );
  NAND2_X1 U9805 ( .A1(n9702), .A2(n9800), .ZN(n9799) );
  NAND2_X1 U9806 ( .A1(n9705), .A2(n9704), .ZN(n9800) );
  XOR2_X1 U9807 ( .A(n9801), .B(n9802), .Z(n9702) );
  NAND2_X1 U9808 ( .A1(n9803), .A2(n9804), .ZN(n9801) );
  NOR2_X1 U9809 ( .A1(n9704), .A2(n9705), .ZN(n9797) );
  NOR2_X1 U9810 ( .A1(n9421), .A2(n8750), .ZN(n9705) );
  NAND2_X1 U9811 ( .A1(n9559), .A2(n9805), .ZN(n9704) );
  NAND2_X1 U9812 ( .A1(n9558), .A2(n9560), .ZN(n9805) );
  NAND2_X1 U9813 ( .A1(n9806), .A2(n9807), .ZN(n9560) );
  NAND2_X1 U9814 ( .A1(b_27_), .A2(a_13_), .ZN(n9807) );
  INV_X1 U9815 ( .A(n9808), .ZN(n9806) );
  XOR2_X1 U9816 ( .A(n9809), .B(n9810), .Z(n9558) );
  XNOR2_X1 U9817 ( .A(n9811), .B(n9812), .ZN(n9810) );
  NAND2_X1 U9818 ( .A1(a_13_), .A2(n9808), .ZN(n9559) );
  NAND2_X1 U9819 ( .A1(n9567), .A2(n9813), .ZN(n9808) );
  NAND2_X1 U9820 ( .A1(n9566), .A2(n9568), .ZN(n9813) );
  NAND2_X1 U9821 ( .A1(n9814), .A2(n9815), .ZN(n9568) );
  NAND2_X1 U9822 ( .A1(b_27_), .A2(a_14_), .ZN(n9815) );
  INV_X1 U9823 ( .A(n9816), .ZN(n9814) );
  XNOR2_X1 U9824 ( .A(n9817), .B(n9818), .ZN(n9566) );
  XOR2_X1 U9825 ( .A(n9819), .B(n9820), .Z(n9818) );
  NAND2_X1 U9826 ( .A1(b_26_), .A2(a_15_), .ZN(n9820) );
  NAND2_X1 U9827 ( .A1(a_14_), .A2(n9816), .ZN(n9567) );
  NAND2_X1 U9828 ( .A1(n9821), .A2(n9822), .ZN(n9816) );
  NAND2_X1 U9829 ( .A1(n9823), .A2(b_27_), .ZN(n9822) );
  NOR2_X1 U9830 ( .A1(n9824), .A2(n8763), .ZN(n9823) );
  NOR2_X1 U9831 ( .A1(n9574), .A2(n9575), .ZN(n9824) );
  NAND2_X1 U9832 ( .A1(n9574), .A2(n9575), .ZN(n9821) );
  NAND2_X1 U9833 ( .A1(n9700), .A2(n9825), .ZN(n9575) );
  NAND2_X1 U9834 ( .A1(n9699), .A2(n9701), .ZN(n9825) );
  NAND2_X1 U9835 ( .A1(n9826), .A2(n9827), .ZN(n9701) );
  NAND2_X1 U9836 ( .A1(b_27_), .A2(a_16_), .ZN(n9827) );
  INV_X1 U9837 ( .A(n9828), .ZN(n9826) );
  XNOR2_X1 U9838 ( .A(n9829), .B(n9830), .ZN(n9699) );
  NAND2_X1 U9839 ( .A1(n9831), .A2(n9832), .ZN(n9829) );
  NAND2_X1 U9840 ( .A1(a_16_), .A2(n9828), .ZN(n9700) );
  NAND2_X1 U9841 ( .A1(n9587), .A2(n9833), .ZN(n9828) );
  NAND2_X1 U9842 ( .A1(n9586), .A2(n9588), .ZN(n9833) );
  NAND2_X1 U9843 ( .A1(n9834), .A2(n9835), .ZN(n9588) );
  NAND2_X1 U9844 ( .A1(b_27_), .A2(a_17_), .ZN(n9835) );
  INV_X1 U9845 ( .A(n9836), .ZN(n9834) );
  XNOR2_X1 U9846 ( .A(n9837), .B(n9838), .ZN(n9586) );
  NAND2_X1 U9847 ( .A1(n9839), .A2(n9840), .ZN(n9837) );
  NAND2_X1 U9848 ( .A1(a_17_), .A2(n9836), .ZN(n9587) );
  NAND2_X1 U9849 ( .A1(n9595), .A2(n9841), .ZN(n9836) );
  NAND2_X1 U9850 ( .A1(n9594), .A2(n9596), .ZN(n9841) );
  NAND2_X1 U9851 ( .A1(n9842), .A2(n9843), .ZN(n9596) );
  NAND2_X1 U9852 ( .A1(b_27_), .A2(a_18_), .ZN(n9843) );
  INV_X1 U9853 ( .A(n9844), .ZN(n9842) );
  XNOR2_X1 U9854 ( .A(n9845), .B(n9846), .ZN(n9594) );
  XOR2_X1 U9855 ( .A(n9847), .B(n9848), .Z(n9846) );
  NAND2_X1 U9856 ( .A1(b_26_), .A2(a_19_), .ZN(n9848) );
  NAND2_X1 U9857 ( .A1(a_18_), .A2(n9844), .ZN(n9595) );
  NAND2_X1 U9858 ( .A1(n9849), .A2(n9850), .ZN(n9844) );
  NAND2_X1 U9859 ( .A1(n9851), .A2(b_27_), .ZN(n9850) );
  NOR2_X1 U9860 ( .A1(n9852), .A2(n8881), .ZN(n9851) );
  NOR2_X1 U9861 ( .A1(n9602), .A2(n9603), .ZN(n9852) );
  NAND2_X1 U9862 ( .A1(n9602), .A2(n9603), .ZN(n9849) );
  NAND2_X1 U9863 ( .A1(n9696), .A2(n9853), .ZN(n9603) );
  NAND2_X1 U9864 ( .A1(n9695), .A2(n9697), .ZN(n9853) );
  NAND2_X1 U9865 ( .A1(n9854), .A2(n9855), .ZN(n9697) );
  NAND2_X1 U9866 ( .A1(b_27_), .A2(a_20_), .ZN(n9855) );
  INV_X1 U9867 ( .A(n9856), .ZN(n9854) );
  XNOR2_X1 U9868 ( .A(n9857), .B(n9858), .ZN(n9695) );
  NAND2_X1 U9869 ( .A1(n9859), .A2(n9860), .ZN(n9857) );
  NAND2_X1 U9870 ( .A1(a_20_), .A2(n9856), .ZN(n9696) );
  NAND2_X1 U9871 ( .A1(n9615), .A2(n9861), .ZN(n9856) );
  NAND2_X1 U9872 ( .A1(n9614), .A2(n9616), .ZN(n9861) );
  NAND2_X1 U9873 ( .A1(n9862), .A2(n9863), .ZN(n9616) );
  NAND2_X1 U9874 ( .A1(b_27_), .A2(a_21_), .ZN(n9863) );
  INV_X1 U9875 ( .A(n9864), .ZN(n9862) );
  XNOR2_X1 U9876 ( .A(n9865), .B(n9866), .ZN(n9614) );
  NAND2_X1 U9877 ( .A1(n9867), .A2(n9868), .ZN(n9865) );
  NAND2_X1 U9878 ( .A1(a_21_), .A2(n9864), .ZN(n9615) );
  NAND2_X1 U9879 ( .A1(n9623), .A2(n9869), .ZN(n9864) );
  NAND2_X1 U9880 ( .A1(n9622), .A2(n9624), .ZN(n9869) );
  NAND2_X1 U9881 ( .A1(n9870), .A2(n9871), .ZN(n9624) );
  NAND2_X1 U9882 ( .A1(b_27_), .A2(a_22_), .ZN(n9871) );
  INV_X1 U9883 ( .A(n9872), .ZN(n9870) );
  XOR2_X1 U9884 ( .A(n9873), .B(n9874), .Z(n9622) );
  XOR2_X1 U9885 ( .A(n9875), .B(n9876), .Z(n9873) );
  NOR2_X1 U9886 ( .A1(n8812), .A2(n9684), .ZN(n9876) );
  NAND2_X1 U9887 ( .A1(a_22_), .A2(n9872), .ZN(n9623) );
  NAND2_X1 U9888 ( .A1(n9877), .A2(n9878), .ZN(n9872) );
  NAND2_X1 U9889 ( .A1(n9879), .A2(b_27_), .ZN(n9878) );
  NOR2_X1 U9890 ( .A1(n9880), .A2(n8812), .ZN(n9879) );
  NOR2_X1 U9891 ( .A1(n9630), .A2(n9631), .ZN(n9880) );
  NAND2_X1 U9892 ( .A1(n9630), .A2(n9631), .ZN(n9877) );
  NAND2_X1 U9893 ( .A1(n9881), .A2(n9882), .ZN(n9631) );
  NAND2_X1 U9894 ( .A1(n9693), .A2(n9883), .ZN(n9882) );
  INV_X1 U9895 ( .A(n9884), .ZN(n9883) );
  NOR2_X1 U9896 ( .A1(n9692), .A2(n9691), .ZN(n9884) );
  NOR2_X1 U9897 ( .A1(n9421), .A2(n9131), .ZN(n9693) );
  NAND2_X1 U9898 ( .A1(n9691), .A2(n9692), .ZN(n9881) );
  NAND2_X1 U9899 ( .A1(n9885), .A2(n9886), .ZN(n9692) );
  NAND2_X1 U9900 ( .A1(n9689), .A2(n9887), .ZN(n9886) );
  NAND2_X1 U9901 ( .A1(n9686), .A2(n9688), .ZN(n9887) );
  NOR2_X1 U9902 ( .A1(n9421), .A2(n8825), .ZN(n9689) );
  INV_X1 U9903 ( .A(n9888), .ZN(n9885) );
  NOR2_X1 U9904 ( .A1(n9688), .A2(n9686), .ZN(n9888) );
  XNOR2_X1 U9905 ( .A(n9889), .B(n9890), .ZN(n9686) );
  XNOR2_X1 U9906 ( .A(n9891), .B(n9892), .ZN(n9889) );
  NAND2_X1 U9907 ( .A1(n9893), .A2(n9894), .ZN(n9688) );
  NAND2_X1 U9908 ( .A1(n9646), .A2(n9895), .ZN(n9894) );
  NAND2_X1 U9909 ( .A1(n9648), .A2(n9647), .ZN(n9895) );
  XOR2_X1 U9910 ( .A(n9896), .B(n9897), .Z(n9646) );
  NAND2_X1 U9911 ( .A1(n9898), .A2(n9899), .ZN(n9896) );
  INV_X1 U9912 ( .A(n9900), .ZN(n9893) );
  NOR2_X1 U9913 ( .A1(n9647), .A2(n9648), .ZN(n9900) );
  NOR2_X1 U9914 ( .A1(n9421), .A2(n8830), .ZN(n9648) );
  NAND2_X1 U9915 ( .A1(n9901), .A2(n9902), .ZN(n9647) );
  INV_X1 U9916 ( .A(n9903), .ZN(n9902) );
  NOR2_X1 U9917 ( .A1(n9653), .A2(n9904), .ZN(n9903) );
  NOR2_X1 U9918 ( .A1(n9656), .A2(n9905), .ZN(n9904) );
  XOR2_X1 U9919 ( .A(n9906), .B(n9907), .Z(n9653) );
  XNOR2_X1 U9920 ( .A(n9908), .B(n9909), .ZN(n9906) );
  NAND2_X1 U9921 ( .A1(n9905), .A2(n9656), .ZN(n9901) );
  NAND2_X1 U9922 ( .A1(n9910), .A2(n9911), .ZN(n9656) );
  NAND2_X1 U9923 ( .A1(n9912), .A2(b_27_), .ZN(n9911) );
  NOR2_X1 U9924 ( .A1(n9913), .A2(n8844), .ZN(n9912) );
  NOR2_X1 U9925 ( .A1(n9662), .A2(n9664), .ZN(n9913) );
  NAND2_X1 U9926 ( .A1(n9662), .A2(n9664), .ZN(n9910) );
  NAND2_X1 U9927 ( .A1(n9914), .A2(n9915), .ZN(n9664) );
  NAND2_X1 U9928 ( .A1(n9669), .A2(n9916), .ZN(n9915) );
  INV_X1 U9929 ( .A(n9917), .ZN(n9916) );
  NOR2_X1 U9930 ( .A1(n9672), .A2(n9671), .ZN(n9917) );
  NOR2_X1 U9931 ( .A1(n9421), .A2(n9161), .ZN(n9669) );
  NAND2_X1 U9932 ( .A1(n9671), .A2(n9672), .ZN(n9914) );
  NAND2_X1 U9933 ( .A1(n9918), .A2(n9919), .ZN(n9672) );
  NAND2_X1 U9934 ( .A1(b_25_), .A2(n9920), .ZN(n9919) );
  NAND2_X1 U9935 ( .A1(n8358), .A2(n9921), .ZN(n9920) );
  NAND2_X1 U9936 ( .A1(a_31_), .A2(n9684), .ZN(n9921) );
  NAND2_X1 U9937 ( .A1(b_26_), .A2(n9922), .ZN(n9918) );
  NAND2_X1 U9938 ( .A1(n8362), .A2(n9923), .ZN(n9922) );
  NAND2_X1 U9939 ( .A1(a_30_), .A2(n9924), .ZN(n9923) );
  NOR2_X1 U9940 ( .A1(n9925), .A2(n9684), .ZN(n9671) );
  NAND2_X1 U9941 ( .A1(n9926), .A2(b_27_), .ZN(n9925) );
  XNOR2_X1 U9942 ( .A(n9927), .B(n9928), .ZN(n9662) );
  XOR2_X1 U9943 ( .A(n9929), .B(n9930), .Z(n9928) );
  XNOR2_X1 U9944 ( .A(n9931), .B(n9932), .ZN(n9691) );
  XNOR2_X1 U9945 ( .A(n9933), .B(n9934), .ZN(n9931) );
  XOR2_X1 U9946 ( .A(n9935), .B(n9936), .Z(n9630) );
  XOR2_X1 U9947 ( .A(n9937), .B(n9938), .Z(n9935) );
  XNOR2_X1 U9948 ( .A(n9939), .B(n9940), .ZN(n9602) );
  NAND2_X1 U9949 ( .A1(n9941), .A2(n9942), .ZN(n9939) );
  XNOR2_X1 U9950 ( .A(n9943), .B(n9944), .ZN(n9574) );
  NAND2_X1 U9951 ( .A1(n9945), .A2(n9946), .ZN(n9943) );
  XNOR2_X1 U9952 ( .A(n9947), .B(n9948), .ZN(n9506) );
  XOR2_X1 U9953 ( .A(n9949), .B(n9950), .Z(n9948) );
  NAND2_X1 U9954 ( .A1(b_26_), .A2(a_7_), .ZN(n9950) );
  XNOR2_X1 U9955 ( .A(n9951), .B(n9952), .ZN(n9707) );
  NAND2_X1 U9956 ( .A1(n9953), .A2(n9954), .ZN(n9951) );
  XOR2_X1 U9957 ( .A(n9955), .B(n9956), .Z(n9710) );
  XOR2_X1 U9958 ( .A(n9957), .B(n9958), .Z(n9955) );
  NOR2_X1 U9959 ( .A1(n8717), .A2(n9684), .ZN(n9958) );
  XNOR2_X1 U9960 ( .A(n9959), .B(n9960), .ZN(n9474) );
  XNOR2_X1 U9961 ( .A(n9961), .B(n9962), .ZN(n9959) );
  XOR2_X1 U9962 ( .A(n9963), .B(n9964), .Z(n9714) );
  XOR2_X1 U9963 ( .A(n9965), .B(n9966), .Z(n9964) );
  XNOR2_X1 U9964 ( .A(n9466), .B(n9467), .ZN(n9720) );
  XNOR2_X1 U9965 ( .A(n9967), .B(n9968), .ZN(n9466) );
  NAND2_X1 U9966 ( .A1(n9969), .A2(n9970), .ZN(n9719) );
  NAND2_X1 U9967 ( .A1(n8670), .A2(n9971), .ZN(n9970) );
  INV_X1 U9968 ( .A(n8535), .ZN(n9969) );
  NAND2_X1 U9969 ( .A1(n8535), .A2(n8536), .ZN(n8537) );
  INV_X1 U9970 ( .A(n9972), .ZN(n8536) );
  NAND2_X1 U9971 ( .A1(n9973), .A2(n8664), .ZN(n9972) );
  NAND2_X1 U9972 ( .A1(n9974), .A2(n9975), .ZN(n9973) );
  INV_X1 U9973 ( .A(n9976), .ZN(n9975) );
  XOR2_X1 U9974 ( .A(n9977), .B(n9978), .Z(n9974) );
  NOR2_X1 U9975 ( .A1(n8670), .A2(n9971), .ZN(n8535) );
  INV_X1 U9976 ( .A(n8669), .ZN(n9971) );
  NAND2_X1 U9977 ( .A1(n9979), .A2(n9980), .ZN(n8669) );
  NAND2_X1 U9978 ( .A1(n9968), .A2(n9981), .ZN(n9980) );
  INV_X1 U9979 ( .A(n9982), .ZN(n9981) );
  NOR2_X1 U9980 ( .A1(n9467), .A2(n9967), .ZN(n9982) );
  NOR2_X1 U9981 ( .A1(n9684), .A2(n8690), .ZN(n9968) );
  NAND2_X1 U9982 ( .A1(n9467), .A2(n9967), .ZN(n9979) );
  NAND2_X1 U9983 ( .A1(n9983), .A2(n9984), .ZN(n9967) );
  NAND2_X1 U9984 ( .A1(n9966), .A2(n9985), .ZN(n9984) );
  NAND2_X1 U9985 ( .A1(n9963), .A2(n9965), .ZN(n9985) );
  NOR2_X1 U9986 ( .A1(n9684), .A2(n8502), .ZN(n9966) );
  INV_X1 U9987 ( .A(n9986), .ZN(n9983) );
  NOR2_X1 U9988 ( .A1(n9963), .A2(n9965), .ZN(n9986) );
  NOR2_X1 U9989 ( .A1(n9987), .A2(n9988), .ZN(n9965) );
  INV_X1 U9990 ( .A(n9989), .ZN(n9988) );
  NAND2_X1 U9991 ( .A1(n9961), .A2(n9990), .ZN(n9989) );
  NAND2_X1 U9992 ( .A1(n9962), .A2(n9960), .ZN(n9990) );
  NOR2_X1 U9993 ( .A1(n9684), .A2(n8497), .ZN(n9961) );
  NOR2_X1 U9994 ( .A1(n9960), .A2(n9962), .ZN(n9987) );
  NOR2_X1 U9995 ( .A1(n9991), .A2(n9992), .ZN(n9962) );
  NOR2_X1 U9996 ( .A1(n9736), .A2(n9993), .ZN(n9992) );
  NOR2_X1 U9997 ( .A1(n9733), .A2(n9735), .ZN(n9993) );
  NAND2_X1 U9998 ( .A1(b_26_), .A2(a_3_), .ZN(n9736) );
  INV_X1 U9999 ( .A(n9994), .ZN(n9991) );
  NAND2_X1 U10000 ( .A1(n9733), .A2(n9735), .ZN(n9994) );
  NAND2_X1 U10001 ( .A1(n9995), .A2(n9996), .ZN(n9735) );
  NAND2_X1 U10002 ( .A1(n9997), .A2(b_26_), .ZN(n9996) );
  NOR2_X1 U10003 ( .A1(n9998), .A2(n8712), .ZN(n9997) );
  NOR2_X1 U10004 ( .A1(n9743), .A2(n9741), .ZN(n9998) );
  NAND2_X1 U10005 ( .A1(n9741), .A2(n9743), .ZN(n9995) );
  NAND2_X1 U10006 ( .A1(n9999), .A2(n10000), .ZN(n9743) );
  NAND2_X1 U10007 ( .A1(n10001), .A2(b_26_), .ZN(n10000) );
  NOR2_X1 U10008 ( .A1(n10002), .A2(n8717), .ZN(n10001) );
  NOR2_X1 U10009 ( .A1(n9956), .A2(n9957), .ZN(n10002) );
  NAND2_X1 U10010 ( .A1(n9956), .A2(n9957), .ZN(n9999) );
  NAND2_X1 U10011 ( .A1(n9953), .A2(n10003), .ZN(n9957) );
  NAND2_X1 U10012 ( .A1(n9952), .A2(n9954), .ZN(n10003) );
  NAND2_X1 U10013 ( .A1(n10004), .A2(n10005), .ZN(n9954) );
  NAND2_X1 U10014 ( .A1(b_26_), .A2(a_6_), .ZN(n10005) );
  INV_X1 U10015 ( .A(n10006), .ZN(n10004) );
  XNOR2_X1 U10016 ( .A(n10007), .B(n10008), .ZN(n9952) );
  NAND2_X1 U10017 ( .A1(n10009), .A2(n10010), .ZN(n10007) );
  NAND2_X1 U10018 ( .A1(a_6_), .A2(n10006), .ZN(n9953) );
  NAND2_X1 U10019 ( .A1(n10011), .A2(n10012), .ZN(n10006) );
  NAND2_X1 U10020 ( .A1(n10013), .A2(b_26_), .ZN(n10012) );
  NOR2_X1 U10021 ( .A1(n10014), .A2(n8726), .ZN(n10013) );
  NOR2_X1 U10022 ( .A1(n9949), .A2(n9947), .ZN(n10014) );
  NAND2_X1 U10023 ( .A1(n9947), .A2(n9949), .ZN(n10011) );
  NAND2_X1 U10024 ( .A1(n10015), .A2(n10016), .ZN(n9949) );
  NAND2_X1 U10025 ( .A1(n10017), .A2(b_26_), .ZN(n10016) );
  NOR2_X1 U10026 ( .A1(n10018), .A2(n8731), .ZN(n10017) );
  NOR2_X1 U10027 ( .A1(n9761), .A2(n9763), .ZN(n10018) );
  NAND2_X1 U10028 ( .A1(n9761), .A2(n9763), .ZN(n10015) );
  NAND2_X1 U10029 ( .A1(n10019), .A2(n10020), .ZN(n9763) );
  NAND2_X1 U10030 ( .A1(n10021), .A2(b_26_), .ZN(n10020) );
  NOR2_X1 U10031 ( .A1(n10022), .A2(n8736), .ZN(n10021) );
  NOR2_X1 U10032 ( .A1(n9771), .A2(n9770), .ZN(n10022) );
  NAND2_X1 U10033 ( .A1(n9771), .A2(n9770), .ZN(n10019) );
  XOR2_X1 U10034 ( .A(n10023), .B(n10024), .Z(n9770) );
  XOR2_X1 U10035 ( .A(n10025), .B(n10026), .Z(n10024) );
  NOR2_X1 U10036 ( .A1(n10027), .A2(n10028), .ZN(n9771) );
  INV_X1 U10037 ( .A(n10029), .ZN(n10028) );
  NAND2_X1 U10038 ( .A1(n9777), .A2(n10030), .ZN(n10029) );
  NAND2_X1 U10039 ( .A1(n9780), .A2(n9779), .ZN(n10030) );
  XNOR2_X1 U10040 ( .A(n10031), .B(n10032), .ZN(n9777) );
  XOR2_X1 U10041 ( .A(n10033), .B(n10034), .Z(n10031) );
  NOR2_X1 U10042 ( .A1(n8452), .A2(n9924), .ZN(n10034) );
  NOR2_X1 U10043 ( .A1(n9779), .A2(n9780), .ZN(n10027) );
  NOR2_X1 U10044 ( .A1(n9684), .A2(n8741), .ZN(n9780) );
  NAND2_X1 U10045 ( .A1(n10035), .A2(n10036), .ZN(n9779) );
  NAND2_X1 U10046 ( .A1(n10037), .A2(b_26_), .ZN(n10036) );
  NOR2_X1 U10047 ( .A1(n10038), .A2(n8452), .ZN(n10037) );
  NOR2_X1 U10048 ( .A1(n9787), .A2(n9786), .ZN(n10038) );
  NAND2_X1 U10049 ( .A1(n9787), .A2(n9786), .ZN(n10035) );
  XNOR2_X1 U10050 ( .A(n10039), .B(n10040), .ZN(n9786) );
  NAND2_X1 U10051 ( .A1(n10041), .A2(n10042), .ZN(n10039) );
  NOR2_X1 U10052 ( .A1(n10043), .A2(n10044), .ZN(n9787) );
  INV_X1 U10053 ( .A(n10045), .ZN(n10044) );
  NAND2_X1 U10054 ( .A1(n9793), .A2(n10046), .ZN(n10045) );
  NAND2_X1 U10055 ( .A1(n9796), .A2(n9795), .ZN(n10046) );
  XOR2_X1 U10056 ( .A(n10047), .B(n10048), .Z(n9793) );
  NAND2_X1 U10057 ( .A1(n10049), .A2(n10050), .ZN(n10047) );
  NOR2_X1 U10058 ( .A1(n9795), .A2(n9796), .ZN(n10043) );
  NOR2_X1 U10059 ( .A1(n9684), .A2(n8750), .ZN(n9796) );
  NAND2_X1 U10060 ( .A1(n9803), .A2(n10051), .ZN(n9795) );
  NAND2_X1 U10061 ( .A1(n9802), .A2(n9804), .ZN(n10051) );
  NAND2_X1 U10062 ( .A1(n10052), .A2(n10053), .ZN(n9804) );
  INV_X1 U10063 ( .A(n10054), .ZN(n10053) );
  NAND2_X1 U10064 ( .A1(b_26_), .A2(a_13_), .ZN(n10052) );
  XNOR2_X1 U10065 ( .A(n10055), .B(n10056), .ZN(n9802) );
  NAND2_X1 U10066 ( .A1(n10057), .A2(n10058), .ZN(n10055) );
  NAND2_X1 U10067 ( .A1(n10054), .A2(a_13_), .ZN(n9803) );
  NOR2_X1 U10068 ( .A1(n10059), .A2(n10060), .ZN(n10054) );
  INV_X1 U10069 ( .A(n10061), .ZN(n10060) );
  NAND2_X1 U10070 ( .A1(n9809), .A2(n10062), .ZN(n10061) );
  NAND2_X1 U10071 ( .A1(n9812), .A2(n9811), .ZN(n10062) );
  XOR2_X1 U10072 ( .A(n10063), .B(n10064), .Z(n9809) );
  NAND2_X1 U10073 ( .A1(n10065), .A2(n10066), .ZN(n10063) );
  NOR2_X1 U10074 ( .A1(n9811), .A2(n9812), .ZN(n10059) );
  NOR2_X1 U10075 ( .A1(n9684), .A2(n8438), .ZN(n9812) );
  NAND2_X1 U10076 ( .A1(n10067), .A2(n10068), .ZN(n9811) );
  NAND2_X1 U10077 ( .A1(n10069), .A2(b_26_), .ZN(n10068) );
  NOR2_X1 U10078 ( .A1(n10070), .A2(n8763), .ZN(n10069) );
  NOR2_X1 U10079 ( .A1(n9817), .A2(n9819), .ZN(n10070) );
  NAND2_X1 U10080 ( .A1(n9817), .A2(n9819), .ZN(n10067) );
  NAND2_X1 U10081 ( .A1(n9945), .A2(n10071), .ZN(n9819) );
  NAND2_X1 U10082 ( .A1(n9944), .A2(n9946), .ZN(n10071) );
  NAND2_X1 U10083 ( .A1(n10072), .A2(n10073), .ZN(n9946) );
  NAND2_X1 U10084 ( .A1(b_26_), .A2(a_16_), .ZN(n10073) );
  INV_X1 U10085 ( .A(n10074), .ZN(n10072) );
  XNOR2_X1 U10086 ( .A(n10075), .B(n10076), .ZN(n9944) );
  NAND2_X1 U10087 ( .A1(n10077), .A2(n10078), .ZN(n10075) );
  NAND2_X1 U10088 ( .A1(a_16_), .A2(n10074), .ZN(n9945) );
  NAND2_X1 U10089 ( .A1(n9831), .A2(n10079), .ZN(n10074) );
  NAND2_X1 U10090 ( .A1(n9830), .A2(n9832), .ZN(n10079) );
  NAND2_X1 U10091 ( .A1(n10080), .A2(n10081), .ZN(n9832) );
  NAND2_X1 U10092 ( .A1(b_26_), .A2(a_17_), .ZN(n10081) );
  INV_X1 U10093 ( .A(n10082), .ZN(n10080) );
  XNOR2_X1 U10094 ( .A(n10083), .B(n10084), .ZN(n9830) );
  NAND2_X1 U10095 ( .A1(n10085), .A2(n10086), .ZN(n10083) );
  NAND2_X1 U10096 ( .A1(a_17_), .A2(n10082), .ZN(n9831) );
  NAND2_X1 U10097 ( .A1(n9839), .A2(n10087), .ZN(n10082) );
  NAND2_X1 U10098 ( .A1(n9838), .A2(n9840), .ZN(n10087) );
  NAND2_X1 U10099 ( .A1(n10088), .A2(n10089), .ZN(n9840) );
  NAND2_X1 U10100 ( .A1(b_26_), .A2(a_18_), .ZN(n10089) );
  INV_X1 U10101 ( .A(n10090), .ZN(n10088) );
  XNOR2_X1 U10102 ( .A(n10091), .B(n10092), .ZN(n9838) );
  XOR2_X1 U10103 ( .A(n10093), .B(n10094), .Z(n10092) );
  NAND2_X1 U10104 ( .A1(b_25_), .A2(a_19_), .ZN(n10094) );
  NAND2_X1 U10105 ( .A1(a_18_), .A2(n10090), .ZN(n9839) );
  NAND2_X1 U10106 ( .A1(n10095), .A2(n10096), .ZN(n10090) );
  NAND2_X1 U10107 ( .A1(n10097), .A2(b_26_), .ZN(n10096) );
  NOR2_X1 U10108 ( .A1(n10098), .A2(n8881), .ZN(n10097) );
  NOR2_X1 U10109 ( .A1(n9847), .A2(n9845), .ZN(n10098) );
  NAND2_X1 U10110 ( .A1(n9845), .A2(n9847), .ZN(n10095) );
  NAND2_X1 U10111 ( .A1(n9941), .A2(n10099), .ZN(n9847) );
  NAND2_X1 U10112 ( .A1(n9940), .A2(n9942), .ZN(n10099) );
  NAND2_X1 U10113 ( .A1(n10100), .A2(n10101), .ZN(n9942) );
  NAND2_X1 U10114 ( .A1(b_26_), .A2(a_20_), .ZN(n10101) );
  INV_X1 U10115 ( .A(n10102), .ZN(n10100) );
  XNOR2_X1 U10116 ( .A(n10103), .B(n10104), .ZN(n9940) );
  NAND2_X1 U10117 ( .A1(n10105), .A2(n10106), .ZN(n10103) );
  NAND2_X1 U10118 ( .A1(a_20_), .A2(n10102), .ZN(n9941) );
  NAND2_X1 U10119 ( .A1(n9859), .A2(n10107), .ZN(n10102) );
  NAND2_X1 U10120 ( .A1(n9858), .A2(n9860), .ZN(n10107) );
  NAND2_X1 U10121 ( .A1(n10108), .A2(n10109), .ZN(n9860) );
  NAND2_X1 U10122 ( .A1(b_26_), .A2(a_21_), .ZN(n10109) );
  INV_X1 U10123 ( .A(n10110), .ZN(n10108) );
  XNOR2_X1 U10124 ( .A(n10111), .B(n10112), .ZN(n9858) );
  NAND2_X1 U10125 ( .A1(n10113), .A2(n10114), .ZN(n10111) );
  NAND2_X1 U10126 ( .A1(a_21_), .A2(n10110), .ZN(n9859) );
  NAND2_X1 U10127 ( .A1(n9867), .A2(n10115), .ZN(n10110) );
  NAND2_X1 U10128 ( .A1(n9866), .A2(n9868), .ZN(n10115) );
  NAND2_X1 U10129 ( .A1(n10116), .A2(n10117), .ZN(n9868) );
  NAND2_X1 U10130 ( .A1(b_26_), .A2(a_22_), .ZN(n10117) );
  INV_X1 U10131 ( .A(n10118), .ZN(n10116) );
  XOR2_X1 U10132 ( .A(n10119), .B(n10120), .Z(n9866) );
  XOR2_X1 U10133 ( .A(n10121), .B(n10122), .Z(n10119) );
  NOR2_X1 U10134 ( .A1(n8812), .A2(n9924), .ZN(n10122) );
  NAND2_X1 U10135 ( .A1(a_22_), .A2(n10118), .ZN(n9867) );
  NAND2_X1 U10136 ( .A1(n10123), .A2(n10124), .ZN(n10118) );
  NAND2_X1 U10137 ( .A1(n10125), .A2(b_26_), .ZN(n10124) );
  NOR2_X1 U10138 ( .A1(n10126), .A2(n8812), .ZN(n10125) );
  NOR2_X1 U10139 ( .A1(n9875), .A2(n9874), .ZN(n10126) );
  NAND2_X1 U10140 ( .A1(n9874), .A2(n9875), .ZN(n10123) );
  NAND2_X1 U10141 ( .A1(n10127), .A2(n10128), .ZN(n9875) );
  NAND2_X1 U10142 ( .A1(n9938), .A2(n10129), .ZN(n10128) );
  INV_X1 U10143 ( .A(n10130), .ZN(n10129) );
  NOR2_X1 U10144 ( .A1(n9936), .A2(n9937), .ZN(n10130) );
  NOR2_X1 U10145 ( .A1(n9684), .A2(n9131), .ZN(n9938) );
  NAND2_X1 U10146 ( .A1(n9936), .A2(n9937), .ZN(n10127) );
  NAND2_X1 U10147 ( .A1(n10131), .A2(n10132), .ZN(n9937) );
  NAND2_X1 U10148 ( .A1(n9934), .A2(n10133), .ZN(n10132) );
  INV_X1 U10149 ( .A(n10134), .ZN(n10133) );
  NOR2_X1 U10150 ( .A1(n9932), .A2(n9933), .ZN(n10134) );
  NOR2_X1 U10151 ( .A1(n9684), .A2(n8825), .ZN(n9934) );
  NAND2_X1 U10152 ( .A1(n9933), .A2(n9932), .ZN(n10131) );
  XOR2_X1 U10153 ( .A(n10135), .B(n10136), .Z(n9932) );
  XNOR2_X1 U10154 ( .A(n10137), .B(n10138), .ZN(n10136) );
  NOR2_X1 U10155 ( .A1(n10139), .A2(n10140), .ZN(n9933) );
  INV_X1 U10156 ( .A(n10141), .ZN(n10140) );
  NAND2_X1 U10157 ( .A1(n10142), .A2(n9892), .ZN(n10141) );
  NAND2_X1 U10158 ( .A1(n9890), .A2(n9891), .ZN(n10142) );
  NOR2_X1 U10159 ( .A1(n9891), .A2(n9890), .ZN(n10139) );
  XNOR2_X1 U10160 ( .A(n10143), .B(n10144), .ZN(n9890) );
  XNOR2_X1 U10161 ( .A(n10145), .B(n10146), .ZN(n10144) );
  NAND2_X1 U10162 ( .A1(n9898), .A2(n10147), .ZN(n9891) );
  NAND2_X1 U10163 ( .A1(n9897), .A2(n9899), .ZN(n10147) );
  NAND2_X1 U10164 ( .A1(n10148), .A2(n10149), .ZN(n9899) );
  NAND2_X1 U10165 ( .A1(b_26_), .A2(a_27_), .ZN(n10149) );
  XNOR2_X1 U10166 ( .A(n10150), .B(n10151), .ZN(n9897) );
  XNOR2_X1 U10167 ( .A(n10152), .B(n10153), .ZN(n10150) );
  INV_X1 U10168 ( .A(n10154), .ZN(n9898) );
  NOR2_X1 U10169 ( .A1(n8839), .A2(n10148), .ZN(n10154) );
  NOR2_X1 U10170 ( .A1(n10155), .A2(n10156), .ZN(n10148) );
  INV_X1 U10171 ( .A(n10157), .ZN(n10156) );
  NAND2_X1 U10172 ( .A1(n9908), .A2(n10158), .ZN(n10157) );
  NAND2_X1 U10173 ( .A1(n9909), .A2(n9907), .ZN(n10158) );
  NOR2_X1 U10174 ( .A1(n9684), .A2(n8844), .ZN(n9908) );
  NOR2_X1 U10175 ( .A1(n9907), .A2(n9909), .ZN(n10155) );
  NOR2_X1 U10176 ( .A1(n10159), .A2(n10160), .ZN(n9909) );
  INV_X1 U10177 ( .A(n10161), .ZN(n10160) );
  NAND2_X1 U10178 ( .A1(n9927), .A2(n10162), .ZN(n10161) );
  NAND2_X1 U10179 ( .A1(n10163), .A2(n9929), .ZN(n10162) );
  NOR2_X1 U10180 ( .A1(n9684), .A2(n9161), .ZN(n9927) );
  NOR2_X1 U10181 ( .A1(n9929), .A2(n10163), .ZN(n10159) );
  INV_X1 U10182 ( .A(n9930), .ZN(n10163) );
  NAND2_X1 U10183 ( .A1(n10164), .A2(n10165), .ZN(n9930) );
  NAND2_X1 U10184 ( .A1(b_24_), .A2(n10166), .ZN(n10165) );
  NAND2_X1 U10185 ( .A1(n8358), .A2(n10167), .ZN(n10166) );
  NAND2_X1 U10186 ( .A1(a_31_), .A2(n9924), .ZN(n10167) );
  NAND2_X1 U10187 ( .A1(b_25_), .A2(n10168), .ZN(n10164) );
  NAND2_X1 U10188 ( .A1(n8362), .A2(n10169), .ZN(n10168) );
  NAND2_X1 U10189 ( .A1(a_30_), .A2(n10170), .ZN(n10169) );
  NAND2_X1 U10190 ( .A1(n10171), .A2(b_26_), .ZN(n9929) );
  NOR2_X1 U10191 ( .A1(n9170), .A2(n9924), .ZN(n10171) );
  XOR2_X1 U10192 ( .A(n10172), .B(n10173), .Z(n9907) );
  XOR2_X1 U10193 ( .A(n10174), .B(n10175), .Z(n10173) );
  XNOR2_X1 U10194 ( .A(n10176), .B(n10177), .ZN(n9936) );
  XOR2_X1 U10195 ( .A(n10178), .B(n10179), .Z(n10177) );
  XNOR2_X1 U10196 ( .A(n10180), .B(n10181), .ZN(n9874) );
  XNOR2_X1 U10197 ( .A(n10182), .B(n10183), .ZN(n10181) );
  XNOR2_X1 U10198 ( .A(n10184), .B(n10185), .ZN(n9845) );
  NAND2_X1 U10199 ( .A1(n10186), .A2(n10187), .ZN(n10184) );
  XOR2_X1 U10200 ( .A(n10188), .B(n10189), .Z(n9817) );
  XNOR2_X1 U10201 ( .A(n10190), .B(n10191), .ZN(n10189) );
  XOR2_X1 U10202 ( .A(n10192), .B(n10193), .Z(n9761) );
  XOR2_X1 U10203 ( .A(n10194), .B(n10195), .Z(n10192) );
  NOR2_X1 U10204 ( .A1(n8736), .A2(n9924), .ZN(n10195) );
  XNOR2_X1 U10205 ( .A(n10196), .B(n10197), .ZN(n9947) );
  XOR2_X1 U10206 ( .A(n10198), .B(n10199), .Z(n10197) );
  NAND2_X1 U10207 ( .A1(b_25_), .A2(a_8_), .ZN(n10199) );
  XNOR2_X1 U10208 ( .A(n10200), .B(n10201), .ZN(n9956) );
  NAND2_X1 U10209 ( .A1(n10202), .A2(n10203), .ZN(n10200) );
  XNOR2_X1 U10210 ( .A(n10204), .B(n10205), .ZN(n9741) );
  XOR2_X1 U10211 ( .A(n10206), .B(n10207), .Z(n10205) );
  NAND2_X1 U10212 ( .A1(b_25_), .A2(a_5_), .ZN(n10207) );
  XNOR2_X1 U10213 ( .A(n10208), .B(n10209), .ZN(n9733) );
  NAND2_X1 U10214 ( .A1(n10210), .A2(n10211), .ZN(n10208) );
  XNOR2_X1 U10215 ( .A(n10212), .B(n10213), .ZN(n9960) );
  XOR2_X1 U10216 ( .A(n10214), .B(n10215), .Z(n10212) );
  NOR2_X1 U10217 ( .A1(n8707), .A2(n9924), .ZN(n10215) );
  XNOR2_X1 U10218 ( .A(n10216), .B(n10217), .ZN(n9963) );
  XOR2_X1 U10219 ( .A(n10218), .B(n10219), .Z(n10216) );
  NOR2_X1 U10220 ( .A1(n8497), .A2(n9924), .ZN(n10219) );
  XNOR2_X1 U10221 ( .A(n10220), .B(n10221), .ZN(n9467) );
  XOR2_X1 U10222 ( .A(n10222), .B(n10223), .Z(n10221) );
  NAND2_X1 U10223 ( .A1(b_25_), .A2(a_1_), .ZN(n10223) );
  XNOR2_X1 U10224 ( .A(n10224), .B(n10225), .ZN(n8670) );
  XOR2_X1 U10225 ( .A(n10226), .B(n10227), .Z(n10224) );
  NOR2_X1 U10226 ( .A1(n8690), .A2(n9924), .ZN(n10227) );
  INV_X1 U10227 ( .A(n10228), .ZN(n8540) );
  NOR2_X1 U10228 ( .A1(n8664), .A2(n8663), .ZN(n10228) );
  NAND2_X1 U10229 ( .A1(n8661), .A2(n10229), .ZN(n8663) );
  INV_X1 U10230 ( .A(n10230), .ZN(n10229) );
  NOR2_X1 U10231 ( .A1(n10231), .A2(n10232), .ZN(n10230) );
  NAND2_X1 U10232 ( .A1(n10233), .A2(n9976), .ZN(n8664) );
  NAND2_X1 U10233 ( .A1(n10234), .A2(n10235), .ZN(n9976) );
  NAND2_X1 U10234 ( .A1(n10236), .A2(b_25_), .ZN(n10235) );
  NOR2_X1 U10235 ( .A1(n10237), .A2(n8690), .ZN(n10236) );
  NOR2_X1 U10236 ( .A1(n10225), .A2(n10226), .ZN(n10237) );
  NAND2_X1 U10237 ( .A1(n10225), .A2(n10226), .ZN(n10234) );
  NAND2_X1 U10238 ( .A1(n10238), .A2(n10239), .ZN(n10226) );
  NAND2_X1 U10239 ( .A1(n10240), .A2(b_25_), .ZN(n10239) );
  NOR2_X1 U10240 ( .A1(n10241), .A2(n8502), .ZN(n10240) );
  NOR2_X1 U10241 ( .A1(n10220), .A2(n10222), .ZN(n10241) );
  NAND2_X1 U10242 ( .A1(n10220), .A2(n10222), .ZN(n10238) );
  NAND2_X1 U10243 ( .A1(n10242), .A2(n10243), .ZN(n10222) );
  NAND2_X1 U10244 ( .A1(n10244), .A2(b_25_), .ZN(n10243) );
  NOR2_X1 U10245 ( .A1(n10245), .A2(n8497), .ZN(n10244) );
  NOR2_X1 U10246 ( .A1(n10217), .A2(n10218), .ZN(n10245) );
  NAND2_X1 U10247 ( .A1(n10217), .A2(n10218), .ZN(n10242) );
  NAND2_X1 U10248 ( .A1(n10246), .A2(n10247), .ZN(n10218) );
  NAND2_X1 U10249 ( .A1(n10248), .A2(b_25_), .ZN(n10247) );
  NOR2_X1 U10250 ( .A1(n10249), .A2(n8707), .ZN(n10248) );
  NOR2_X1 U10251 ( .A1(n10213), .A2(n10214), .ZN(n10249) );
  NAND2_X1 U10252 ( .A1(n10213), .A2(n10214), .ZN(n10246) );
  NAND2_X1 U10253 ( .A1(n10210), .A2(n10250), .ZN(n10214) );
  NAND2_X1 U10254 ( .A1(n10209), .A2(n10211), .ZN(n10250) );
  NAND2_X1 U10255 ( .A1(n10251), .A2(n10252), .ZN(n10211) );
  NAND2_X1 U10256 ( .A1(b_25_), .A2(a_4_), .ZN(n10252) );
  INV_X1 U10257 ( .A(n10253), .ZN(n10251) );
  XOR2_X1 U10258 ( .A(n10254), .B(n10255), .Z(n10209) );
  XOR2_X1 U10259 ( .A(n10256), .B(n10257), .Z(n10254) );
  NAND2_X1 U10260 ( .A1(a_4_), .A2(n10253), .ZN(n10210) );
  NAND2_X1 U10261 ( .A1(n10258), .A2(n10259), .ZN(n10253) );
  NAND2_X1 U10262 ( .A1(n10260), .A2(b_25_), .ZN(n10259) );
  NOR2_X1 U10263 ( .A1(n10261), .A2(n8717), .ZN(n10260) );
  NOR2_X1 U10264 ( .A1(n10204), .A2(n10206), .ZN(n10261) );
  NAND2_X1 U10265 ( .A1(n10204), .A2(n10206), .ZN(n10258) );
  NAND2_X1 U10266 ( .A1(n10202), .A2(n10262), .ZN(n10206) );
  NAND2_X1 U10267 ( .A1(n10201), .A2(n10203), .ZN(n10262) );
  NAND2_X1 U10268 ( .A1(n10263), .A2(n10264), .ZN(n10203) );
  NAND2_X1 U10269 ( .A1(b_25_), .A2(a_6_), .ZN(n10264) );
  INV_X1 U10270 ( .A(n10265), .ZN(n10263) );
  XNOR2_X1 U10271 ( .A(n10266), .B(n10267), .ZN(n10201) );
  NAND2_X1 U10272 ( .A1(n10268), .A2(n10269), .ZN(n10266) );
  NAND2_X1 U10273 ( .A1(a_6_), .A2(n10265), .ZN(n10202) );
  NAND2_X1 U10274 ( .A1(n10009), .A2(n10270), .ZN(n10265) );
  NAND2_X1 U10275 ( .A1(n10008), .A2(n10010), .ZN(n10270) );
  NAND2_X1 U10276 ( .A1(n10271), .A2(n10272), .ZN(n10010) );
  NAND2_X1 U10277 ( .A1(b_25_), .A2(a_7_), .ZN(n10272) );
  INV_X1 U10278 ( .A(n10273), .ZN(n10271) );
  XNOR2_X1 U10279 ( .A(n10274), .B(n10275), .ZN(n10008) );
  XOR2_X1 U10280 ( .A(n10276), .B(n10277), .Z(n10275) );
  NAND2_X1 U10281 ( .A1(b_24_), .A2(a_8_), .ZN(n10277) );
  NAND2_X1 U10282 ( .A1(a_7_), .A2(n10273), .ZN(n10009) );
  NAND2_X1 U10283 ( .A1(n10278), .A2(n10279), .ZN(n10273) );
  NAND2_X1 U10284 ( .A1(n10280), .A2(b_25_), .ZN(n10279) );
  NOR2_X1 U10285 ( .A1(n10281), .A2(n8731), .ZN(n10280) );
  NOR2_X1 U10286 ( .A1(n10196), .A2(n10198), .ZN(n10281) );
  NAND2_X1 U10287 ( .A1(n10196), .A2(n10198), .ZN(n10278) );
  NAND2_X1 U10288 ( .A1(n10282), .A2(n10283), .ZN(n10198) );
  NAND2_X1 U10289 ( .A1(n10284), .A2(b_25_), .ZN(n10283) );
  NOR2_X1 U10290 ( .A1(n10285), .A2(n8736), .ZN(n10284) );
  NOR2_X1 U10291 ( .A1(n10193), .A2(n10194), .ZN(n10285) );
  NAND2_X1 U10292 ( .A1(n10193), .A2(n10194), .ZN(n10282) );
  NAND2_X1 U10293 ( .A1(n10286), .A2(n10287), .ZN(n10194) );
  NAND2_X1 U10294 ( .A1(n10025), .A2(n10288), .ZN(n10287) );
  NAND2_X1 U10295 ( .A1(n10023), .A2(n10026), .ZN(n10288) );
  NAND2_X1 U10296 ( .A1(n10289), .A2(n10290), .ZN(n10025) );
  NAND2_X1 U10297 ( .A1(n10291), .A2(b_25_), .ZN(n10290) );
  NOR2_X1 U10298 ( .A1(n10292), .A2(n8452), .ZN(n10291) );
  NOR2_X1 U10299 ( .A1(n10032), .A2(n10033), .ZN(n10292) );
  NAND2_X1 U10300 ( .A1(n10032), .A2(n10033), .ZN(n10289) );
  NAND2_X1 U10301 ( .A1(n10041), .A2(n10293), .ZN(n10033) );
  NAND2_X1 U10302 ( .A1(n10040), .A2(n10042), .ZN(n10293) );
  NAND2_X1 U10303 ( .A1(n10294), .A2(n10295), .ZN(n10042) );
  NAND2_X1 U10304 ( .A1(b_25_), .A2(a_12_), .ZN(n10295) );
  INV_X1 U10305 ( .A(n10296), .ZN(n10294) );
  XNOR2_X1 U10306 ( .A(n10297), .B(n10298), .ZN(n10040) );
  NAND2_X1 U10307 ( .A1(n10299), .A2(n10300), .ZN(n10297) );
  NAND2_X1 U10308 ( .A1(a_12_), .A2(n10296), .ZN(n10041) );
  NAND2_X1 U10309 ( .A1(n10049), .A2(n10301), .ZN(n10296) );
  NAND2_X1 U10310 ( .A1(n10048), .A2(n10050), .ZN(n10301) );
  NAND2_X1 U10311 ( .A1(n10302), .A2(n10303), .ZN(n10050) );
  NAND2_X1 U10312 ( .A1(b_25_), .A2(a_13_), .ZN(n10303) );
  INV_X1 U10313 ( .A(n10304), .ZN(n10302) );
  XOR2_X1 U10314 ( .A(n10305), .B(n10306), .Z(n10048) );
  XNOR2_X1 U10315 ( .A(n10307), .B(n10308), .ZN(n10306) );
  NAND2_X1 U10316 ( .A1(a_13_), .A2(n10304), .ZN(n10049) );
  NAND2_X1 U10317 ( .A1(n10057), .A2(n10309), .ZN(n10304) );
  NAND2_X1 U10318 ( .A1(n10056), .A2(n10058), .ZN(n10309) );
  NAND2_X1 U10319 ( .A1(n10310), .A2(n10311), .ZN(n10058) );
  NAND2_X1 U10320 ( .A1(b_25_), .A2(a_14_), .ZN(n10311) );
  INV_X1 U10321 ( .A(n10312), .ZN(n10310) );
  XNOR2_X1 U10322 ( .A(n10313), .B(n10314), .ZN(n10056) );
  XNOR2_X1 U10323 ( .A(n10315), .B(n10316), .ZN(n10313) );
  NOR2_X1 U10324 ( .A1(n8763), .A2(n10170), .ZN(n10316) );
  NAND2_X1 U10325 ( .A1(a_14_), .A2(n10312), .ZN(n10057) );
  NAND2_X1 U10326 ( .A1(n10065), .A2(n10317), .ZN(n10312) );
  NAND2_X1 U10327 ( .A1(n10064), .A2(n10066), .ZN(n10317) );
  NAND2_X1 U10328 ( .A1(n10318), .A2(n10319), .ZN(n10066) );
  INV_X1 U10329 ( .A(n10320), .ZN(n10319) );
  NAND2_X1 U10330 ( .A1(b_25_), .A2(a_15_), .ZN(n10318) );
  XOR2_X1 U10331 ( .A(n10321), .B(n10322), .Z(n10064) );
  XNOR2_X1 U10332 ( .A(n10323), .B(n10324), .ZN(n10322) );
  NAND2_X1 U10333 ( .A1(n10320), .A2(a_15_), .ZN(n10065) );
  NOR2_X1 U10334 ( .A1(n10325), .A2(n10326), .ZN(n10320) );
  INV_X1 U10335 ( .A(n10327), .ZN(n10326) );
  NAND2_X1 U10336 ( .A1(n10188), .A2(n10328), .ZN(n10327) );
  NAND2_X1 U10337 ( .A1(n10191), .A2(n10190), .ZN(n10328) );
  XOR2_X1 U10338 ( .A(n10329), .B(n10330), .Z(n10188) );
  NAND2_X1 U10339 ( .A1(n10331), .A2(n10332), .ZN(n10329) );
  NOR2_X1 U10340 ( .A1(n10190), .A2(n10191), .ZN(n10325) );
  NOR2_X1 U10341 ( .A1(n9924), .A2(n8768), .ZN(n10191) );
  NAND2_X1 U10342 ( .A1(n10077), .A2(n10333), .ZN(n10190) );
  NAND2_X1 U10343 ( .A1(n10076), .A2(n10078), .ZN(n10333) );
  NAND2_X1 U10344 ( .A1(n10334), .A2(n10335), .ZN(n10078) );
  NAND2_X1 U10345 ( .A1(b_25_), .A2(a_17_), .ZN(n10335) );
  INV_X1 U10346 ( .A(n10336), .ZN(n10334) );
  XOR2_X1 U10347 ( .A(n10337), .B(n10338), .Z(n10076) );
  XNOR2_X1 U10348 ( .A(n10339), .B(n10340), .ZN(n10338) );
  NAND2_X1 U10349 ( .A1(a_17_), .A2(n10336), .ZN(n10077) );
  NAND2_X1 U10350 ( .A1(n10085), .A2(n10341), .ZN(n10336) );
  NAND2_X1 U10351 ( .A1(n10084), .A2(n10086), .ZN(n10341) );
  NAND2_X1 U10352 ( .A1(n10342), .A2(n10343), .ZN(n10086) );
  NAND2_X1 U10353 ( .A1(b_25_), .A2(a_18_), .ZN(n10343) );
  INV_X1 U10354 ( .A(n10344), .ZN(n10342) );
  XOR2_X1 U10355 ( .A(n10345), .B(n10346), .Z(n10084) );
  XNOR2_X1 U10356 ( .A(n10347), .B(n10348), .ZN(n10346) );
  NAND2_X1 U10357 ( .A1(b_24_), .A2(a_19_), .ZN(n10348) );
  NAND2_X1 U10358 ( .A1(a_18_), .A2(n10344), .ZN(n10085) );
  NAND2_X1 U10359 ( .A1(n10349), .A2(n10350), .ZN(n10344) );
  NAND2_X1 U10360 ( .A1(n10351), .A2(b_25_), .ZN(n10350) );
  NOR2_X1 U10361 ( .A1(n10352), .A2(n8881), .ZN(n10351) );
  NOR2_X1 U10362 ( .A1(n10091), .A2(n10093), .ZN(n10352) );
  NAND2_X1 U10363 ( .A1(n10091), .A2(n10093), .ZN(n10349) );
  NAND2_X1 U10364 ( .A1(n10186), .A2(n10353), .ZN(n10093) );
  NAND2_X1 U10365 ( .A1(n10185), .A2(n10187), .ZN(n10353) );
  NAND2_X1 U10366 ( .A1(n10354), .A2(n10355), .ZN(n10187) );
  NAND2_X1 U10367 ( .A1(b_25_), .A2(a_20_), .ZN(n10355) );
  INV_X1 U10368 ( .A(n10356), .ZN(n10354) );
  XNOR2_X1 U10369 ( .A(n10357), .B(n10358), .ZN(n10185) );
  NAND2_X1 U10370 ( .A1(n10359), .A2(n10360), .ZN(n10357) );
  NAND2_X1 U10371 ( .A1(a_20_), .A2(n10356), .ZN(n10186) );
  NAND2_X1 U10372 ( .A1(n10105), .A2(n10361), .ZN(n10356) );
  NAND2_X1 U10373 ( .A1(n10104), .A2(n10106), .ZN(n10361) );
  NAND2_X1 U10374 ( .A1(n10362), .A2(n10363), .ZN(n10106) );
  NAND2_X1 U10375 ( .A1(b_25_), .A2(a_21_), .ZN(n10363) );
  INV_X1 U10376 ( .A(n10364), .ZN(n10362) );
  XNOR2_X1 U10377 ( .A(n10365), .B(n10366), .ZN(n10104) );
  NAND2_X1 U10378 ( .A1(n10367), .A2(n10368), .ZN(n10365) );
  NAND2_X1 U10379 ( .A1(a_21_), .A2(n10364), .ZN(n10105) );
  NAND2_X1 U10380 ( .A1(n10113), .A2(n10369), .ZN(n10364) );
  NAND2_X1 U10381 ( .A1(n10112), .A2(n10114), .ZN(n10369) );
  NAND2_X1 U10382 ( .A1(n10370), .A2(n10371), .ZN(n10114) );
  NAND2_X1 U10383 ( .A1(b_25_), .A2(a_22_), .ZN(n10371) );
  INV_X1 U10384 ( .A(n10372), .ZN(n10370) );
  XOR2_X1 U10385 ( .A(n10373), .B(n10374), .Z(n10112) );
  XNOR2_X1 U10386 ( .A(n10375), .B(n10376), .ZN(n10374) );
  NAND2_X1 U10387 ( .A1(b_24_), .A2(a_23_), .ZN(n10376) );
  NAND2_X1 U10388 ( .A1(a_22_), .A2(n10372), .ZN(n10113) );
  NAND2_X1 U10389 ( .A1(n10377), .A2(n10378), .ZN(n10372) );
  NAND2_X1 U10390 ( .A1(n10379), .A2(b_25_), .ZN(n10378) );
  NOR2_X1 U10391 ( .A1(n10380), .A2(n8812), .ZN(n10379) );
  NOR2_X1 U10392 ( .A1(n10120), .A2(n10121), .ZN(n10380) );
  NAND2_X1 U10393 ( .A1(n10120), .A2(n10121), .ZN(n10377) );
  NAND2_X1 U10394 ( .A1(n10381), .A2(n10382), .ZN(n10121) );
  NAND2_X1 U10395 ( .A1(n10183), .A2(n10383), .ZN(n10382) );
  NAND2_X1 U10396 ( .A1(n10180), .A2(n10182), .ZN(n10383) );
  NOR2_X1 U10397 ( .A1(n9924), .A2(n9131), .ZN(n10183) );
  INV_X1 U10398 ( .A(n10384), .ZN(n10381) );
  NOR2_X1 U10399 ( .A1(n10182), .A2(n10180), .ZN(n10384) );
  XOR2_X1 U10400 ( .A(n10385), .B(n10386), .Z(n10180) );
  XNOR2_X1 U10401 ( .A(n10387), .B(n10388), .ZN(n10386) );
  NAND2_X1 U10402 ( .A1(n10389), .A2(n10390), .ZN(n10182) );
  NAND2_X1 U10403 ( .A1(n10176), .A2(n10391), .ZN(n10390) );
  NAND2_X1 U10404 ( .A1(n10392), .A2(n10393), .ZN(n10391) );
  INV_X1 U10405 ( .A(n10178), .ZN(n10392) );
  XNOR2_X1 U10406 ( .A(n10394), .B(n10395), .ZN(n10176) );
  XNOR2_X1 U10407 ( .A(n10396), .B(n10397), .ZN(n10395) );
  NAND2_X1 U10408 ( .A1(n10179), .A2(n10178), .ZN(n10389) );
  NAND2_X1 U10409 ( .A1(n10398), .A2(n10399), .ZN(n10178) );
  NAND2_X1 U10410 ( .A1(n10135), .A2(n10400), .ZN(n10399) );
  NAND2_X1 U10411 ( .A1(n10138), .A2(n10137), .ZN(n10400) );
  XNOR2_X1 U10412 ( .A(n10401), .B(n10402), .ZN(n10135) );
  XOR2_X1 U10413 ( .A(n10403), .B(n10404), .Z(n10402) );
  INV_X1 U10414 ( .A(n10405), .ZN(n10398) );
  NOR2_X1 U10415 ( .A1(n10137), .A2(n10138), .ZN(n10405) );
  NOR2_X1 U10416 ( .A1(n9924), .A2(n8830), .ZN(n10138) );
  NAND2_X1 U10417 ( .A1(n10406), .A2(n10407), .ZN(n10137) );
  NAND2_X1 U10418 ( .A1(n10146), .A2(n10408), .ZN(n10407) );
  INV_X1 U10419 ( .A(n10409), .ZN(n10408) );
  NOR2_X1 U10420 ( .A1(n10145), .A2(n10143), .ZN(n10409) );
  NOR2_X1 U10421 ( .A1(n9924), .A2(n8839), .ZN(n10146) );
  NAND2_X1 U10422 ( .A1(n10143), .A2(n10145), .ZN(n10406) );
  NAND2_X1 U10423 ( .A1(n10410), .A2(n10411), .ZN(n10145) );
  NAND2_X1 U10424 ( .A1(n10152), .A2(n10412), .ZN(n10411) );
  NAND2_X1 U10425 ( .A1(n10153), .A2(n10151), .ZN(n10412) );
  NOR2_X1 U10426 ( .A1(n9924), .A2(n8844), .ZN(n10152) );
  INV_X1 U10427 ( .A(n10413), .ZN(n10410) );
  NOR2_X1 U10428 ( .A1(n10151), .A2(n10153), .ZN(n10413) );
  NOR2_X1 U10429 ( .A1(n10414), .A2(n10415), .ZN(n10153) );
  INV_X1 U10430 ( .A(n10416), .ZN(n10415) );
  NAND2_X1 U10431 ( .A1(n10172), .A2(n10417), .ZN(n10416) );
  NAND2_X1 U10432 ( .A1(n10418), .A2(n10174), .ZN(n10417) );
  NOR2_X1 U10433 ( .A1(n9924), .A2(n9161), .ZN(n10172) );
  NOR2_X1 U10434 ( .A1(n10174), .A2(n10418), .ZN(n10414) );
  INV_X1 U10435 ( .A(n10175), .ZN(n10418) );
  NAND2_X1 U10436 ( .A1(n10419), .A2(n10420), .ZN(n10175) );
  NAND2_X1 U10437 ( .A1(b_23_), .A2(n10421), .ZN(n10420) );
  NAND2_X1 U10438 ( .A1(n8358), .A2(n10422), .ZN(n10421) );
  NAND2_X1 U10439 ( .A1(a_31_), .A2(n10170), .ZN(n10422) );
  NAND2_X1 U10440 ( .A1(b_24_), .A2(n10423), .ZN(n10419) );
  NAND2_X1 U10441 ( .A1(n8362), .A2(n10424), .ZN(n10423) );
  NAND2_X1 U10442 ( .A1(a_30_), .A2(n10425), .ZN(n10424) );
  NAND2_X1 U10443 ( .A1(n10426), .A2(b_25_), .ZN(n10174) );
  NOR2_X1 U10444 ( .A1(n9170), .A2(n10170), .ZN(n10426) );
  XOR2_X1 U10445 ( .A(n10427), .B(n10428), .Z(n10151) );
  XOR2_X1 U10446 ( .A(n10429), .B(n10430), .Z(n10428) );
  XNOR2_X1 U10447 ( .A(n10431), .B(n10432), .ZN(n10143) );
  XNOR2_X1 U10448 ( .A(n10433), .B(n10434), .ZN(n10431) );
  XOR2_X1 U10449 ( .A(n10435), .B(n10436), .Z(n10120) );
  XNOR2_X1 U10450 ( .A(n10437), .B(n10438), .ZN(n10435) );
  XNOR2_X1 U10451 ( .A(n10439), .B(n10440), .ZN(n10091) );
  XOR2_X1 U10452 ( .A(n10441), .B(n10442), .Z(n10439) );
  XOR2_X1 U10453 ( .A(n10443), .B(n10444), .Z(n10032) );
  XOR2_X1 U10454 ( .A(n10445), .B(n10446), .Z(n10443) );
  NOR2_X1 U10455 ( .A1(n8750), .A2(n10170), .ZN(n10446) );
  INV_X1 U10456 ( .A(n10447), .ZN(n10286) );
  NOR2_X1 U10457 ( .A1(n10026), .A2(n10023), .ZN(n10447) );
  XOR2_X1 U10458 ( .A(n10448), .B(n10449), .Z(n10023) );
  XOR2_X1 U10459 ( .A(n10450), .B(n10451), .Z(n10449) );
  NAND2_X1 U10460 ( .A1(b_24_), .A2(a_11_), .ZN(n10451) );
  NAND2_X1 U10461 ( .A1(b_25_), .A2(a_10_), .ZN(n10026) );
  XNOR2_X1 U10462 ( .A(n10452), .B(n10453), .ZN(n10193) );
  NAND2_X1 U10463 ( .A1(n10454), .A2(n10455), .ZN(n10452) );
  XOR2_X1 U10464 ( .A(n10456), .B(n10457), .Z(n10196) );
  XOR2_X1 U10465 ( .A(n10458), .B(n10459), .Z(n10456) );
  NOR2_X1 U10466 ( .A1(n8736), .A2(n10170), .ZN(n10459) );
  XOR2_X1 U10467 ( .A(n10460), .B(n10461), .Z(n10204) );
  XOR2_X1 U10468 ( .A(n10462), .B(n10463), .Z(n10460) );
  XOR2_X1 U10469 ( .A(n10464), .B(n10465), .Z(n10213) );
  XOR2_X1 U10470 ( .A(n10466), .B(n10467), .Z(n10464) );
  NOR2_X1 U10471 ( .A1(n8712), .A2(n10170), .ZN(n10467) );
  XNOR2_X1 U10472 ( .A(n10468), .B(n10469), .ZN(n10217) );
  NAND2_X1 U10473 ( .A1(n10470), .A2(n10471), .ZN(n10468) );
  XNOR2_X1 U10474 ( .A(n10472), .B(n10473), .ZN(n10220) );
  NAND2_X1 U10475 ( .A1(n10474), .A2(n10475), .ZN(n10472) );
  XNOR2_X1 U10476 ( .A(n10476), .B(n10477), .ZN(n10225) );
  XOR2_X1 U10477 ( .A(n10478), .B(n10479), .Z(n10477) );
  NAND2_X1 U10478 ( .A1(b_24_), .A2(a_1_), .ZN(n10479) );
  XNOR2_X1 U10479 ( .A(n9977), .B(n9978), .ZN(n10233) );
  NAND2_X1 U10480 ( .A1(n10480), .A2(n10481), .ZN(n9977) );
  INV_X1 U10481 ( .A(n10482), .ZN(n8545) );
  NOR2_X1 U10482 ( .A1(n8661), .A2(n8660), .ZN(n10482) );
  NAND2_X1 U10483 ( .A1(n10483), .A2(n10484), .ZN(n8660) );
  NAND2_X1 U10484 ( .A1(n10485), .A2(n10486), .ZN(n10484) );
  INV_X1 U10485 ( .A(n8655), .ZN(n10483) );
  NOR2_X1 U10486 ( .A1(n10486), .A2(n10485), .ZN(n8655) );
  INV_X1 U10487 ( .A(n10487), .ZN(n10485) );
  NAND2_X1 U10488 ( .A1(n10488), .A2(n10489), .ZN(n10487) );
  NAND2_X1 U10489 ( .A1(n10490), .A2(n10491), .ZN(n10489) );
  XOR2_X1 U10490 ( .A(n10492), .B(n10493), .Z(n10486) );
  XOR2_X1 U10491 ( .A(n10494), .B(n10495), .Z(n10493) );
  NAND2_X1 U10492 ( .A1(n10232), .A2(n10231), .ZN(n8661) );
  NAND2_X1 U10493 ( .A1(n10480), .A2(n10496), .ZN(n10231) );
  NAND2_X1 U10494 ( .A1(n9978), .A2(n10481), .ZN(n10496) );
  NAND2_X1 U10495 ( .A1(n10497), .A2(n10498), .ZN(n10481) );
  NAND2_X1 U10496 ( .A1(b_24_), .A2(a_0_), .ZN(n10498) );
  INV_X1 U10497 ( .A(n10499), .ZN(n10497) );
  XNOR2_X1 U10498 ( .A(n10500), .B(n10501), .ZN(n9978) );
  NAND2_X1 U10499 ( .A1(n10502), .A2(n10503), .ZN(n10500) );
  NAND2_X1 U10500 ( .A1(a_0_), .A2(n10499), .ZN(n10480) );
  NAND2_X1 U10501 ( .A1(n10504), .A2(n10505), .ZN(n10499) );
  NAND2_X1 U10502 ( .A1(n10506), .A2(b_24_), .ZN(n10505) );
  NOR2_X1 U10503 ( .A1(n10507), .A2(n8502), .ZN(n10506) );
  NOR2_X1 U10504 ( .A1(n10476), .A2(n10478), .ZN(n10507) );
  NAND2_X1 U10505 ( .A1(n10476), .A2(n10478), .ZN(n10504) );
  NAND2_X1 U10506 ( .A1(n10474), .A2(n10508), .ZN(n10478) );
  NAND2_X1 U10507 ( .A1(n10473), .A2(n10475), .ZN(n10508) );
  NAND2_X1 U10508 ( .A1(n10509), .A2(n10510), .ZN(n10475) );
  NAND2_X1 U10509 ( .A1(b_24_), .A2(a_2_), .ZN(n10510) );
  INV_X1 U10510 ( .A(n10511), .ZN(n10509) );
  XOR2_X1 U10511 ( .A(n10512), .B(n10513), .Z(n10473) );
  XNOR2_X1 U10512 ( .A(n10514), .B(n10515), .ZN(n10513) );
  NAND2_X1 U10513 ( .A1(a_2_), .A2(n10511), .ZN(n10474) );
  NAND2_X1 U10514 ( .A1(n10470), .A2(n10516), .ZN(n10511) );
  NAND2_X1 U10515 ( .A1(n10469), .A2(n10471), .ZN(n10516) );
  NAND2_X1 U10516 ( .A1(n10517), .A2(n10518), .ZN(n10471) );
  NAND2_X1 U10517 ( .A1(b_24_), .A2(a_3_), .ZN(n10518) );
  INV_X1 U10518 ( .A(n10519), .ZN(n10517) );
  XOR2_X1 U10519 ( .A(n10520), .B(n10521), .Z(n10469) );
  XOR2_X1 U10520 ( .A(n10522), .B(n10523), .Z(n10520) );
  NOR2_X1 U10521 ( .A1(n8712), .A2(n10425), .ZN(n10523) );
  NAND2_X1 U10522 ( .A1(a_3_), .A2(n10519), .ZN(n10470) );
  NAND2_X1 U10523 ( .A1(n10524), .A2(n10525), .ZN(n10519) );
  NAND2_X1 U10524 ( .A1(n10526), .A2(b_24_), .ZN(n10525) );
  NOR2_X1 U10525 ( .A1(n10527), .A2(n8712), .ZN(n10526) );
  NOR2_X1 U10526 ( .A1(n10465), .A2(n10466), .ZN(n10527) );
  NAND2_X1 U10527 ( .A1(n10465), .A2(n10466), .ZN(n10524) );
  NAND2_X1 U10528 ( .A1(n10528), .A2(n10529), .ZN(n10466) );
  NAND2_X1 U10529 ( .A1(n10257), .A2(n10530), .ZN(n10529) );
  INV_X1 U10530 ( .A(n10531), .ZN(n10530) );
  NOR2_X1 U10531 ( .A1(n10256), .A2(n10255), .ZN(n10531) );
  NOR2_X1 U10532 ( .A1(n10170), .A2(n8717), .ZN(n10257) );
  NAND2_X1 U10533 ( .A1(n10255), .A2(n10256), .ZN(n10528) );
  NAND2_X1 U10534 ( .A1(n10532), .A2(n10533), .ZN(n10256) );
  NAND2_X1 U10535 ( .A1(n10463), .A2(n10534), .ZN(n10533) );
  INV_X1 U10536 ( .A(n10535), .ZN(n10534) );
  NOR2_X1 U10537 ( .A1(n10462), .A2(n10461), .ZN(n10535) );
  NOR2_X1 U10538 ( .A1(n10170), .A2(n8480), .ZN(n10463) );
  NAND2_X1 U10539 ( .A1(n10461), .A2(n10462), .ZN(n10532) );
  NAND2_X1 U10540 ( .A1(n10268), .A2(n10536), .ZN(n10462) );
  NAND2_X1 U10541 ( .A1(n10267), .A2(n10269), .ZN(n10536) );
  NAND2_X1 U10542 ( .A1(n10537), .A2(n10538), .ZN(n10269) );
  NAND2_X1 U10543 ( .A1(b_24_), .A2(a_7_), .ZN(n10538) );
  INV_X1 U10544 ( .A(n10539), .ZN(n10537) );
  XOR2_X1 U10545 ( .A(n10540), .B(n10541), .Z(n10267) );
  XOR2_X1 U10546 ( .A(n10542), .B(n10543), .Z(n10540) );
  NAND2_X1 U10547 ( .A1(a_7_), .A2(n10539), .ZN(n10268) );
  NAND2_X1 U10548 ( .A1(n10544), .A2(n10545), .ZN(n10539) );
  NAND2_X1 U10549 ( .A1(n10546), .A2(b_24_), .ZN(n10545) );
  NOR2_X1 U10550 ( .A1(n10547), .A2(n8731), .ZN(n10546) );
  NOR2_X1 U10551 ( .A1(n10274), .A2(n10276), .ZN(n10547) );
  NAND2_X1 U10552 ( .A1(n10274), .A2(n10276), .ZN(n10544) );
  NAND2_X1 U10553 ( .A1(n10548), .A2(n10549), .ZN(n10276) );
  NAND2_X1 U10554 ( .A1(n10550), .A2(b_24_), .ZN(n10549) );
  NOR2_X1 U10555 ( .A1(n10551), .A2(n8736), .ZN(n10550) );
  NOR2_X1 U10556 ( .A1(n10457), .A2(n10458), .ZN(n10551) );
  NAND2_X1 U10557 ( .A1(n10457), .A2(n10458), .ZN(n10548) );
  NAND2_X1 U10558 ( .A1(n10454), .A2(n10552), .ZN(n10458) );
  NAND2_X1 U10559 ( .A1(n10453), .A2(n10455), .ZN(n10552) );
  NAND2_X1 U10560 ( .A1(n10553), .A2(n10554), .ZN(n10455) );
  NAND2_X1 U10561 ( .A1(b_24_), .A2(a_10_), .ZN(n10554) );
  INV_X1 U10562 ( .A(n10555), .ZN(n10553) );
  XNOR2_X1 U10563 ( .A(n10556), .B(n10557), .ZN(n10453) );
  XOR2_X1 U10564 ( .A(n10558), .B(n10559), .Z(n10557) );
  NAND2_X1 U10565 ( .A1(b_23_), .A2(a_11_), .ZN(n10559) );
  NAND2_X1 U10566 ( .A1(a_10_), .A2(n10555), .ZN(n10454) );
  NAND2_X1 U10567 ( .A1(n10560), .A2(n10561), .ZN(n10555) );
  NAND2_X1 U10568 ( .A1(n10562), .A2(b_24_), .ZN(n10561) );
  NOR2_X1 U10569 ( .A1(n10563), .A2(n8452), .ZN(n10562) );
  NOR2_X1 U10570 ( .A1(n10448), .A2(n10450), .ZN(n10563) );
  NAND2_X1 U10571 ( .A1(n10448), .A2(n10450), .ZN(n10560) );
  NAND2_X1 U10572 ( .A1(n10564), .A2(n10565), .ZN(n10450) );
  NAND2_X1 U10573 ( .A1(n10566), .A2(b_24_), .ZN(n10565) );
  NOR2_X1 U10574 ( .A1(n10567), .A2(n8750), .ZN(n10566) );
  NOR2_X1 U10575 ( .A1(n10444), .A2(n10445), .ZN(n10567) );
  NAND2_X1 U10576 ( .A1(n10444), .A2(n10445), .ZN(n10564) );
  NAND2_X1 U10577 ( .A1(n10299), .A2(n10568), .ZN(n10445) );
  NAND2_X1 U10578 ( .A1(n10298), .A2(n10300), .ZN(n10568) );
  NAND2_X1 U10579 ( .A1(n10569), .A2(n10570), .ZN(n10300) );
  INV_X1 U10580 ( .A(n10571), .ZN(n10570) );
  NAND2_X1 U10581 ( .A1(b_24_), .A2(a_13_), .ZN(n10569) );
  XNOR2_X1 U10582 ( .A(n10572), .B(n10573), .ZN(n10298) );
  NAND2_X1 U10583 ( .A1(n10574), .A2(n10575), .ZN(n10572) );
  NAND2_X1 U10584 ( .A1(n10571), .A2(a_13_), .ZN(n10299) );
  NOR2_X1 U10585 ( .A1(n10576), .A2(n10577), .ZN(n10571) );
  INV_X1 U10586 ( .A(n10578), .ZN(n10577) );
  NAND2_X1 U10587 ( .A1(n10305), .A2(n10579), .ZN(n10578) );
  NAND2_X1 U10588 ( .A1(n10308), .A2(n10307), .ZN(n10579) );
  XOR2_X1 U10589 ( .A(n10580), .B(n10581), .Z(n10305) );
  XOR2_X1 U10590 ( .A(n10582), .B(n10583), .Z(n10581) );
  NAND2_X1 U10591 ( .A1(b_23_), .A2(a_15_), .ZN(n10583) );
  NOR2_X1 U10592 ( .A1(n10307), .A2(n10308), .ZN(n10576) );
  NOR2_X1 U10593 ( .A1(n10170), .A2(n8438), .ZN(n10308) );
  NAND2_X1 U10594 ( .A1(n10584), .A2(n10585), .ZN(n10307) );
  NAND2_X1 U10595 ( .A1(n10586), .A2(b_24_), .ZN(n10585) );
  NOR2_X1 U10596 ( .A1(n10587), .A2(n8763), .ZN(n10586) );
  NOR2_X1 U10597 ( .A1(n10315), .A2(n10314), .ZN(n10587) );
  NAND2_X1 U10598 ( .A1(n10315), .A2(n10314), .ZN(n10584) );
  XNOR2_X1 U10599 ( .A(n10588), .B(n10589), .ZN(n10314) );
  NAND2_X1 U10600 ( .A1(n10590), .A2(n10591), .ZN(n10588) );
  NOR2_X1 U10601 ( .A1(n10592), .A2(n10593), .ZN(n10315) );
  INV_X1 U10602 ( .A(n10594), .ZN(n10593) );
  NAND2_X1 U10603 ( .A1(n10321), .A2(n10595), .ZN(n10594) );
  NAND2_X1 U10604 ( .A1(n10324), .A2(n10323), .ZN(n10595) );
  XOR2_X1 U10605 ( .A(n10596), .B(n10597), .Z(n10321) );
  NAND2_X1 U10606 ( .A1(n10598), .A2(n10599), .ZN(n10596) );
  NOR2_X1 U10607 ( .A1(n10323), .A2(n10324), .ZN(n10592) );
  NOR2_X1 U10608 ( .A1(n10170), .A2(n8768), .ZN(n10324) );
  NAND2_X1 U10609 ( .A1(n10331), .A2(n10600), .ZN(n10323) );
  NAND2_X1 U10610 ( .A1(n10330), .A2(n10332), .ZN(n10600) );
  NAND2_X1 U10611 ( .A1(n10601), .A2(n10602), .ZN(n10332) );
  INV_X1 U10612 ( .A(n10603), .ZN(n10602) );
  NAND2_X1 U10613 ( .A1(b_24_), .A2(a_17_), .ZN(n10601) );
  XNOR2_X1 U10614 ( .A(n10604), .B(n10605), .ZN(n10330) );
  NAND2_X1 U10615 ( .A1(n10606), .A2(n10607), .ZN(n10604) );
  NAND2_X1 U10616 ( .A1(n10603), .A2(a_17_), .ZN(n10331) );
  NOR2_X1 U10617 ( .A1(n10608), .A2(n10609), .ZN(n10603) );
  INV_X1 U10618 ( .A(n10610), .ZN(n10609) );
  NAND2_X1 U10619 ( .A1(n10337), .A2(n10611), .ZN(n10610) );
  NAND2_X1 U10620 ( .A1(n10340), .A2(n10339), .ZN(n10611) );
  XNOR2_X1 U10621 ( .A(n10612), .B(n10613), .ZN(n10337) );
  XNOR2_X1 U10622 ( .A(n10614), .B(n10615), .ZN(n10613) );
  NOR2_X1 U10623 ( .A1(n10339), .A2(n10340), .ZN(n10608) );
  NOR2_X1 U10624 ( .A1(n10170), .A2(n10616), .ZN(n10340) );
  NAND2_X1 U10625 ( .A1(n10617), .A2(n10618), .ZN(n10339) );
  NAND2_X1 U10626 ( .A1(n10619), .A2(b_24_), .ZN(n10618) );
  NOR2_X1 U10627 ( .A1(n10620), .A2(n8881), .ZN(n10619) );
  NOR2_X1 U10628 ( .A1(n10347), .A2(n10345), .ZN(n10620) );
  NAND2_X1 U10629 ( .A1(n10347), .A2(n10345), .ZN(n10617) );
  XNOR2_X1 U10630 ( .A(n10621), .B(n10622), .ZN(n10345) );
  NAND2_X1 U10631 ( .A1(n10623), .A2(n10624), .ZN(n10621) );
  NOR2_X1 U10632 ( .A1(n10625), .A2(n10626), .ZN(n10347) );
  INV_X1 U10633 ( .A(n10627), .ZN(n10626) );
  NAND2_X1 U10634 ( .A1(n10440), .A2(n10628), .ZN(n10627) );
  NAND2_X1 U10635 ( .A1(n10442), .A2(n10441), .ZN(n10628) );
  XOR2_X1 U10636 ( .A(n10629), .B(n10630), .Z(n10440) );
  NAND2_X1 U10637 ( .A1(n10631), .A2(n10632), .ZN(n10629) );
  NOR2_X1 U10638 ( .A1(n10441), .A2(n10442), .ZN(n10625) );
  NOR2_X1 U10639 ( .A1(n10170), .A2(n10633), .ZN(n10442) );
  NAND2_X1 U10640 ( .A1(n10359), .A2(n10634), .ZN(n10441) );
  NAND2_X1 U10641 ( .A1(n10358), .A2(n10360), .ZN(n10634) );
  NAND2_X1 U10642 ( .A1(n10635), .A2(n10636), .ZN(n10360) );
  NAND2_X1 U10643 ( .A1(b_24_), .A2(a_21_), .ZN(n10636) );
  INV_X1 U10644 ( .A(n10637), .ZN(n10635) );
  XNOR2_X1 U10645 ( .A(n10638), .B(n10639), .ZN(n10358) );
  NAND2_X1 U10646 ( .A1(n10640), .A2(n10641), .ZN(n10638) );
  NAND2_X1 U10647 ( .A1(a_21_), .A2(n10637), .ZN(n10359) );
  NAND2_X1 U10648 ( .A1(n10367), .A2(n10642), .ZN(n10637) );
  NAND2_X1 U10649 ( .A1(n10366), .A2(n10368), .ZN(n10642) );
  NAND2_X1 U10650 ( .A1(n10643), .A2(n10644), .ZN(n10368) );
  NAND2_X1 U10651 ( .A1(b_24_), .A2(a_22_), .ZN(n10644) );
  INV_X1 U10652 ( .A(n10645), .ZN(n10643) );
  XNOR2_X1 U10653 ( .A(n10646), .B(n10647), .ZN(n10366) );
  XOR2_X1 U10654 ( .A(n10648), .B(n10649), .Z(n10646) );
  NAND2_X1 U10655 ( .A1(a_22_), .A2(n10645), .ZN(n10367) );
  NAND2_X1 U10656 ( .A1(n10650), .A2(n10651), .ZN(n10645) );
  NAND2_X1 U10657 ( .A1(n10652), .A2(b_24_), .ZN(n10651) );
  NOR2_X1 U10658 ( .A1(n10653), .A2(n8812), .ZN(n10652) );
  NOR2_X1 U10659 ( .A1(n10375), .A2(n10373), .ZN(n10653) );
  NAND2_X1 U10660 ( .A1(n10375), .A2(n10373), .ZN(n10650) );
  XOR2_X1 U10661 ( .A(n10654), .B(n10655), .Z(n10373) );
  XOR2_X1 U10662 ( .A(n10656), .B(n10657), .Z(n10654) );
  NOR2_X1 U10663 ( .A1(n10658), .A2(n10659), .ZN(n10375) );
  INV_X1 U10664 ( .A(n10660), .ZN(n10659) );
  NAND2_X1 U10665 ( .A1(n10661), .A2(n10438), .ZN(n10660) );
  NAND2_X1 U10666 ( .A1(n10436), .A2(n10437), .ZN(n10661) );
  NOR2_X1 U10667 ( .A1(n10437), .A2(n10436), .ZN(n10658) );
  XNOR2_X1 U10668 ( .A(n10662), .B(n10663), .ZN(n10436) );
  XNOR2_X1 U10669 ( .A(n10664), .B(n10665), .ZN(n10663) );
  NAND2_X1 U10670 ( .A1(n10666), .A2(n10667), .ZN(n10437) );
  NAND2_X1 U10671 ( .A1(n10388), .A2(n10668), .ZN(n10667) );
  NAND2_X1 U10672 ( .A1(n10385), .A2(n10387), .ZN(n10668) );
  NOR2_X1 U10673 ( .A1(n10170), .A2(n8825), .ZN(n10388) );
  INV_X1 U10674 ( .A(n10669), .ZN(n10666) );
  NOR2_X1 U10675 ( .A1(n10387), .A2(n10385), .ZN(n10669) );
  XNOR2_X1 U10676 ( .A(n10670), .B(n10671), .ZN(n10385) );
  XNOR2_X1 U10677 ( .A(n10672), .B(n10673), .ZN(n10671) );
  NAND2_X1 U10678 ( .A1(n10674), .A2(n10675), .ZN(n10387) );
  NAND2_X1 U10679 ( .A1(n10394), .A2(n10676), .ZN(n10675) );
  NAND2_X1 U10680 ( .A1(n10397), .A2(n10396), .ZN(n10676) );
  XNOR2_X1 U10681 ( .A(n10677), .B(n10678), .ZN(n10394) );
  XOR2_X1 U10682 ( .A(n10679), .B(n10680), .Z(n10678) );
  INV_X1 U10683 ( .A(n10681), .ZN(n10674) );
  NOR2_X1 U10684 ( .A1(n10396), .A2(n10397), .ZN(n10681) );
  NOR2_X1 U10685 ( .A1(n10170), .A2(n8830), .ZN(n10397) );
  NAND2_X1 U10686 ( .A1(n10682), .A2(n10683), .ZN(n10396) );
  NAND2_X1 U10687 ( .A1(n10404), .A2(n10684), .ZN(n10683) );
  NAND2_X1 U10688 ( .A1(n10403), .A2(n10401), .ZN(n10684) );
  NOR2_X1 U10689 ( .A1(n10170), .A2(n8839), .ZN(n10404) );
  INV_X1 U10690 ( .A(n10685), .ZN(n10682) );
  NOR2_X1 U10691 ( .A1(n10401), .A2(n10403), .ZN(n10685) );
  NOR2_X1 U10692 ( .A1(n10686), .A2(n10687), .ZN(n10403) );
  INV_X1 U10693 ( .A(n10688), .ZN(n10687) );
  NAND2_X1 U10694 ( .A1(n10433), .A2(n10689), .ZN(n10688) );
  NAND2_X1 U10695 ( .A1(n10434), .A2(n10432), .ZN(n10689) );
  NOR2_X1 U10696 ( .A1(n10170), .A2(n8844), .ZN(n10433) );
  NOR2_X1 U10697 ( .A1(n10432), .A2(n10434), .ZN(n10686) );
  NOR2_X1 U10698 ( .A1(n10690), .A2(n10691), .ZN(n10434) );
  INV_X1 U10699 ( .A(n10692), .ZN(n10691) );
  NAND2_X1 U10700 ( .A1(n10427), .A2(n10693), .ZN(n10692) );
  NAND2_X1 U10701 ( .A1(n10694), .A2(n10429), .ZN(n10693) );
  NOR2_X1 U10702 ( .A1(n10170), .A2(n9161), .ZN(n10427) );
  NOR2_X1 U10703 ( .A1(n10429), .A2(n10694), .ZN(n10690) );
  INV_X1 U10704 ( .A(n10430), .ZN(n10694) );
  NAND2_X1 U10705 ( .A1(n10695), .A2(n10696), .ZN(n10430) );
  NAND2_X1 U10706 ( .A1(b_22_), .A2(n10697), .ZN(n10696) );
  NAND2_X1 U10707 ( .A1(n8358), .A2(n10698), .ZN(n10697) );
  NAND2_X1 U10708 ( .A1(a_31_), .A2(n10425), .ZN(n10698) );
  NAND2_X1 U10709 ( .A1(b_23_), .A2(n10699), .ZN(n10695) );
  NAND2_X1 U10710 ( .A1(n8362), .A2(n10700), .ZN(n10699) );
  NAND2_X1 U10711 ( .A1(a_30_), .A2(n10701), .ZN(n10700) );
  NAND2_X1 U10712 ( .A1(n10702), .A2(b_24_), .ZN(n10429) );
  XOR2_X1 U10713 ( .A(n10703), .B(n10704), .Z(n10432) );
  XOR2_X1 U10714 ( .A(n10705), .B(n10706), .Z(n10704) );
  XOR2_X1 U10715 ( .A(n10707), .B(n10708), .Z(n10401) );
  XNOR2_X1 U10716 ( .A(n10709), .B(n10710), .ZN(n10707) );
  XOR2_X1 U10717 ( .A(n10711), .B(n10712), .Z(n10444) );
  XOR2_X1 U10718 ( .A(n10713), .B(n10714), .Z(n10711) );
  NOR2_X1 U10719 ( .A1(n8443), .A2(n10425), .ZN(n10714) );
  XNOR2_X1 U10720 ( .A(n10715), .B(n10716), .ZN(n10448) );
  XOR2_X1 U10721 ( .A(n10717), .B(n10718), .Z(n10716) );
  NAND2_X1 U10722 ( .A1(b_23_), .A2(a_12_), .ZN(n10718) );
  XOR2_X1 U10723 ( .A(n10719), .B(n10720), .Z(n10457) );
  XOR2_X1 U10724 ( .A(n10721), .B(n10722), .Z(n10720) );
  XOR2_X1 U10725 ( .A(n10723), .B(n10724), .Z(n10274) );
  XOR2_X1 U10726 ( .A(n10725), .B(n10726), .Z(n10723) );
  XOR2_X1 U10727 ( .A(n10727), .B(n10728), .Z(n10461) );
  XOR2_X1 U10728 ( .A(n10729), .B(n10730), .Z(n10727) );
  NOR2_X1 U10729 ( .A1(n8726), .A2(n10425), .ZN(n10730) );
  XNOR2_X1 U10730 ( .A(n10731), .B(n10732), .ZN(n10255) );
  XOR2_X1 U10731 ( .A(n10733), .B(n10734), .Z(n10732) );
  XOR2_X1 U10732 ( .A(n10735), .B(n10736), .Z(n10465) );
  XOR2_X1 U10733 ( .A(n10737), .B(n10738), .Z(n10735) );
  NOR2_X1 U10734 ( .A1(n8717), .A2(n10425), .ZN(n10738) );
  XNOR2_X1 U10735 ( .A(n10739), .B(n10740), .ZN(n10476) );
  NAND2_X1 U10736 ( .A1(n10741), .A2(n10742), .ZN(n10739) );
  XNOR2_X1 U10737 ( .A(n10743), .B(n10490), .ZN(n10232) );
  XNOR2_X1 U10738 ( .A(n10744), .B(n10745), .ZN(n10490) );
  XNOR2_X1 U10739 ( .A(n10746), .B(n10747), .ZN(n10745) );
  NAND2_X1 U10740 ( .A1(n10488), .A2(n10491), .ZN(n10743) );
  NAND2_X1 U10741 ( .A1(n10748), .A2(n10749), .ZN(n10491) );
  NAND2_X1 U10742 ( .A1(b_23_), .A2(a_0_), .ZN(n10749) );
  INV_X1 U10743 ( .A(n10750), .ZN(n10748) );
  NAND2_X1 U10744 ( .A1(a_0_), .A2(n10750), .ZN(n10488) );
  NAND2_X1 U10745 ( .A1(n10502), .A2(n10751), .ZN(n10750) );
  NAND2_X1 U10746 ( .A1(n10501), .A2(n10503), .ZN(n10751) );
  NAND2_X1 U10747 ( .A1(n10752), .A2(n10753), .ZN(n10503) );
  NAND2_X1 U10748 ( .A1(b_23_), .A2(a_1_), .ZN(n10753) );
  INV_X1 U10749 ( .A(n10754), .ZN(n10752) );
  XOR2_X1 U10750 ( .A(n10755), .B(n10756), .Z(n10501) );
  XNOR2_X1 U10751 ( .A(n10757), .B(n10758), .ZN(n10756) );
  NAND2_X1 U10752 ( .A1(a_1_), .A2(n10754), .ZN(n10502) );
  NAND2_X1 U10753 ( .A1(n10741), .A2(n10759), .ZN(n10754) );
  NAND2_X1 U10754 ( .A1(n10740), .A2(n10742), .ZN(n10759) );
  NAND2_X1 U10755 ( .A1(n10760), .A2(n10761), .ZN(n10742) );
  INV_X1 U10756 ( .A(n10762), .ZN(n10761) );
  NAND2_X1 U10757 ( .A1(b_23_), .A2(a_2_), .ZN(n10760) );
  XNOR2_X1 U10758 ( .A(n10763), .B(n10764), .ZN(n10740) );
  NAND2_X1 U10759 ( .A1(n10765), .A2(n10766), .ZN(n10763) );
  NAND2_X1 U10760 ( .A1(n10762), .A2(a_2_), .ZN(n10741) );
  NOR2_X1 U10761 ( .A1(n10767), .A2(n10768), .ZN(n10762) );
  INV_X1 U10762 ( .A(n10769), .ZN(n10768) );
  NAND2_X1 U10763 ( .A1(n10512), .A2(n10770), .ZN(n10769) );
  NAND2_X1 U10764 ( .A1(n10515), .A2(n10514), .ZN(n10770) );
  XNOR2_X1 U10765 ( .A(n10771), .B(n10772), .ZN(n10512) );
  XNOR2_X1 U10766 ( .A(n10773), .B(n10774), .ZN(n10772) );
  NOR2_X1 U10767 ( .A1(n10514), .A2(n10515), .ZN(n10767) );
  NOR2_X1 U10768 ( .A1(n10425), .A2(n8707), .ZN(n10515) );
  NAND2_X1 U10769 ( .A1(n10775), .A2(n10776), .ZN(n10514) );
  NAND2_X1 U10770 ( .A1(n10777), .A2(b_23_), .ZN(n10776) );
  NOR2_X1 U10771 ( .A1(n10778), .A2(n8712), .ZN(n10777) );
  NOR2_X1 U10772 ( .A1(n10521), .A2(n10522), .ZN(n10778) );
  NAND2_X1 U10773 ( .A1(n10521), .A2(n10522), .ZN(n10775) );
  NAND2_X1 U10774 ( .A1(n10779), .A2(n10780), .ZN(n10522) );
  NAND2_X1 U10775 ( .A1(n10781), .A2(b_23_), .ZN(n10780) );
  NOR2_X1 U10776 ( .A1(n10782), .A2(n8717), .ZN(n10781) );
  NOR2_X1 U10777 ( .A1(n10736), .A2(n10737), .ZN(n10782) );
  NAND2_X1 U10778 ( .A1(n10736), .A2(n10737), .ZN(n10779) );
  NAND2_X1 U10779 ( .A1(n10783), .A2(n10784), .ZN(n10737) );
  NAND2_X1 U10780 ( .A1(n10785), .A2(n10786), .ZN(n10784) );
  INV_X1 U10781 ( .A(n10787), .ZN(n10786) );
  NOR2_X1 U10782 ( .A1(n10734), .A2(n10731), .ZN(n10787) );
  INV_X1 U10783 ( .A(n10733), .ZN(n10785) );
  NAND2_X1 U10784 ( .A1(b_23_), .A2(a_6_), .ZN(n10733) );
  NAND2_X1 U10785 ( .A1(n10731), .A2(n10734), .ZN(n10783) );
  NAND2_X1 U10786 ( .A1(n10788), .A2(n10789), .ZN(n10734) );
  NAND2_X1 U10787 ( .A1(n10790), .A2(b_23_), .ZN(n10789) );
  NOR2_X1 U10788 ( .A1(n10791), .A2(n8726), .ZN(n10790) );
  NOR2_X1 U10789 ( .A1(n10728), .A2(n10729), .ZN(n10791) );
  NAND2_X1 U10790 ( .A1(n10728), .A2(n10729), .ZN(n10788) );
  NAND2_X1 U10791 ( .A1(n10792), .A2(n10793), .ZN(n10729) );
  NAND2_X1 U10792 ( .A1(n10543), .A2(n10794), .ZN(n10793) );
  INV_X1 U10793 ( .A(n10795), .ZN(n10794) );
  NOR2_X1 U10794 ( .A1(n10542), .A2(n10541), .ZN(n10795) );
  NOR2_X1 U10795 ( .A1(n10425), .A2(n8731), .ZN(n10543) );
  NAND2_X1 U10796 ( .A1(n10541), .A2(n10542), .ZN(n10792) );
  NAND2_X1 U10797 ( .A1(n10796), .A2(n10797), .ZN(n10542) );
  NAND2_X1 U10798 ( .A1(n10726), .A2(n10798), .ZN(n10797) );
  INV_X1 U10799 ( .A(n10799), .ZN(n10798) );
  NOR2_X1 U10800 ( .A1(n10725), .A2(n10724), .ZN(n10799) );
  NOR2_X1 U10801 ( .A1(n10425), .A2(n8736), .ZN(n10726) );
  NAND2_X1 U10802 ( .A1(n10724), .A2(n10725), .ZN(n10796) );
  NAND2_X1 U10803 ( .A1(n10800), .A2(n10801), .ZN(n10725) );
  NAND2_X1 U10804 ( .A1(n10721), .A2(n10802), .ZN(n10801) );
  NAND2_X1 U10805 ( .A1(n10719), .A2(n10722), .ZN(n10802) );
  NAND2_X1 U10806 ( .A1(n10803), .A2(n10804), .ZN(n10721) );
  NAND2_X1 U10807 ( .A1(n10805), .A2(b_23_), .ZN(n10804) );
  NOR2_X1 U10808 ( .A1(n10806), .A2(n8452), .ZN(n10805) );
  NOR2_X1 U10809 ( .A1(n10556), .A2(n10558), .ZN(n10806) );
  NAND2_X1 U10810 ( .A1(n10556), .A2(n10558), .ZN(n10803) );
  NAND2_X1 U10811 ( .A1(n10807), .A2(n10808), .ZN(n10558) );
  NAND2_X1 U10812 ( .A1(n10809), .A2(b_23_), .ZN(n10808) );
  NOR2_X1 U10813 ( .A1(n10810), .A2(n8750), .ZN(n10809) );
  NOR2_X1 U10814 ( .A1(n10715), .A2(n10717), .ZN(n10810) );
  NAND2_X1 U10815 ( .A1(n10715), .A2(n10717), .ZN(n10807) );
  NAND2_X1 U10816 ( .A1(n10811), .A2(n10812), .ZN(n10717) );
  NAND2_X1 U10817 ( .A1(n10813), .A2(b_23_), .ZN(n10812) );
  NOR2_X1 U10818 ( .A1(n10814), .A2(n8443), .ZN(n10813) );
  NOR2_X1 U10819 ( .A1(n10712), .A2(n10713), .ZN(n10814) );
  NAND2_X1 U10820 ( .A1(n10712), .A2(n10713), .ZN(n10811) );
  NAND2_X1 U10821 ( .A1(n10574), .A2(n10815), .ZN(n10713) );
  NAND2_X1 U10822 ( .A1(n10573), .A2(n10575), .ZN(n10815) );
  NAND2_X1 U10823 ( .A1(n10816), .A2(n10817), .ZN(n10575) );
  NAND2_X1 U10824 ( .A1(b_23_), .A2(a_14_), .ZN(n10817) );
  INV_X1 U10825 ( .A(n10818), .ZN(n10816) );
  XOR2_X1 U10826 ( .A(n10819), .B(n10820), .Z(n10573) );
  XOR2_X1 U10827 ( .A(n10821), .B(n10822), .Z(n10819) );
  NOR2_X1 U10828 ( .A1(n8763), .A2(n10701), .ZN(n10822) );
  NAND2_X1 U10829 ( .A1(a_14_), .A2(n10818), .ZN(n10574) );
  NAND2_X1 U10830 ( .A1(n10823), .A2(n10824), .ZN(n10818) );
  NAND2_X1 U10831 ( .A1(n10825), .A2(b_23_), .ZN(n10824) );
  NOR2_X1 U10832 ( .A1(n10826), .A2(n8763), .ZN(n10825) );
  NOR2_X1 U10833 ( .A1(n10580), .A2(n10582), .ZN(n10826) );
  NAND2_X1 U10834 ( .A1(n10580), .A2(n10582), .ZN(n10823) );
  NAND2_X1 U10835 ( .A1(n10590), .A2(n10827), .ZN(n10582) );
  NAND2_X1 U10836 ( .A1(n10589), .A2(n10591), .ZN(n10827) );
  NAND2_X1 U10837 ( .A1(n10828), .A2(n10829), .ZN(n10591) );
  NAND2_X1 U10838 ( .A1(b_23_), .A2(a_16_), .ZN(n10829) );
  INV_X1 U10839 ( .A(n10830), .ZN(n10828) );
  XNOR2_X1 U10840 ( .A(n10831), .B(n10832), .ZN(n10589) );
  NAND2_X1 U10841 ( .A1(n10833), .A2(n10834), .ZN(n10831) );
  NAND2_X1 U10842 ( .A1(a_16_), .A2(n10830), .ZN(n10590) );
  NAND2_X1 U10843 ( .A1(n10598), .A2(n10835), .ZN(n10830) );
  NAND2_X1 U10844 ( .A1(n10597), .A2(n10599), .ZN(n10835) );
  NAND2_X1 U10845 ( .A1(n10836), .A2(n10837), .ZN(n10599) );
  NAND2_X1 U10846 ( .A1(b_23_), .A2(a_17_), .ZN(n10837) );
  INV_X1 U10847 ( .A(n10838), .ZN(n10836) );
  XNOR2_X1 U10848 ( .A(n10839), .B(n10840), .ZN(n10597) );
  NAND2_X1 U10849 ( .A1(n10841), .A2(n10842), .ZN(n10839) );
  NAND2_X1 U10850 ( .A1(a_17_), .A2(n10838), .ZN(n10598) );
  NAND2_X1 U10851 ( .A1(n10606), .A2(n10843), .ZN(n10838) );
  NAND2_X1 U10852 ( .A1(n10605), .A2(n10607), .ZN(n10843) );
  NAND2_X1 U10853 ( .A1(n10844), .A2(n10845), .ZN(n10607) );
  INV_X1 U10854 ( .A(n10846), .ZN(n10845) );
  NAND2_X1 U10855 ( .A1(b_23_), .A2(a_18_), .ZN(n10844) );
  XOR2_X1 U10856 ( .A(n10847), .B(n10848), .Z(n10605) );
  XOR2_X1 U10857 ( .A(n10849), .B(n10850), .Z(n10847) );
  NOR2_X1 U10858 ( .A1(n8881), .A2(n10701), .ZN(n10850) );
  NAND2_X1 U10859 ( .A1(n10846), .A2(a_18_), .ZN(n10606) );
  NOR2_X1 U10860 ( .A1(n10851), .A2(n10852), .ZN(n10846) );
  INV_X1 U10861 ( .A(n10853), .ZN(n10852) );
  NAND2_X1 U10862 ( .A1(n10612), .A2(n10854), .ZN(n10853) );
  NAND2_X1 U10863 ( .A1(n10615), .A2(n10614), .ZN(n10854) );
  XOR2_X1 U10864 ( .A(n10855), .B(n10856), .Z(n10612) );
  NAND2_X1 U10865 ( .A1(n10857), .A2(n10858), .ZN(n10855) );
  NOR2_X1 U10866 ( .A1(n10614), .A2(n10615), .ZN(n10851) );
  NOR2_X1 U10867 ( .A1(n10425), .A2(n8881), .ZN(n10615) );
  NAND2_X1 U10868 ( .A1(n10623), .A2(n10859), .ZN(n10614) );
  NAND2_X1 U10869 ( .A1(n10622), .A2(n10624), .ZN(n10859) );
  NAND2_X1 U10870 ( .A1(n10860), .A2(n10861), .ZN(n10624) );
  NAND2_X1 U10871 ( .A1(b_23_), .A2(a_20_), .ZN(n10861) );
  INV_X1 U10872 ( .A(n10862), .ZN(n10860) );
  XNOR2_X1 U10873 ( .A(n10863), .B(n10864), .ZN(n10622) );
  NAND2_X1 U10874 ( .A1(n10865), .A2(n10866), .ZN(n10863) );
  NAND2_X1 U10875 ( .A1(a_20_), .A2(n10862), .ZN(n10623) );
  NAND2_X1 U10876 ( .A1(n10631), .A2(n10867), .ZN(n10862) );
  NAND2_X1 U10877 ( .A1(n10630), .A2(n10632), .ZN(n10867) );
  NAND2_X1 U10878 ( .A1(n10868), .A2(n10869), .ZN(n10632) );
  NAND2_X1 U10879 ( .A1(b_23_), .A2(a_21_), .ZN(n10869) );
  INV_X1 U10880 ( .A(n10870), .ZN(n10868) );
  XOR2_X1 U10881 ( .A(n10871), .B(n10872), .Z(n10630) );
  XNOR2_X1 U10882 ( .A(n10873), .B(n10874), .ZN(n10871) );
  NAND2_X1 U10883 ( .A1(a_21_), .A2(n10870), .ZN(n10631) );
  NAND2_X1 U10884 ( .A1(n10640), .A2(n10875), .ZN(n10870) );
  NAND2_X1 U10885 ( .A1(n10639), .A2(n10641), .ZN(n10875) );
  NAND2_X1 U10886 ( .A1(n10876), .A2(n10877), .ZN(n10641) );
  NAND2_X1 U10887 ( .A1(b_23_), .A2(a_22_), .ZN(n10876) );
  XOR2_X1 U10888 ( .A(n10878), .B(n10879), .Z(n10639) );
  XOR2_X1 U10889 ( .A(n10880), .B(n10881), .Z(n10878) );
  NOR2_X1 U10890 ( .A1(n8812), .A2(n10701), .ZN(n10881) );
  NAND2_X1 U10891 ( .A1(n10882), .A2(a_22_), .ZN(n10640) );
  INV_X1 U10892 ( .A(n10877), .ZN(n10882) );
  NAND2_X1 U10893 ( .A1(n10883), .A2(n10884), .ZN(n10877) );
  NAND2_X1 U10894 ( .A1(n10647), .A2(n10885), .ZN(n10884) );
  NAND2_X1 U10895 ( .A1(n10886), .A2(n10887), .ZN(n10885) );
  XNOR2_X1 U10896 ( .A(n10888), .B(n10889), .ZN(n10647) );
  XOR2_X1 U10897 ( .A(n10890), .B(n10891), .Z(n10888) );
  NAND2_X1 U10898 ( .A1(n10648), .A2(n10649), .ZN(n10883) );
  INV_X1 U10899 ( .A(n10887), .ZN(n10648) );
  NAND2_X1 U10900 ( .A1(n10892), .A2(n10893), .ZN(n10887) );
  NAND2_X1 U10901 ( .A1(n10657), .A2(n10894), .ZN(n10893) );
  INV_X1 U10902 ( .A(n10895), .ZN(n10894) );
  NOR2_X1 U10903 ( .A1(n10656), .A2(n10655), .ZN(n10895) );
  NOR2_X1 U10904 ( .A1(n10425), .A2(n9131), .ZN(n10657) );
  NAND2_X1 U10905 ( .A1(n10655), .A2(n10656), .ZN(n10892) );
  NAND2_X1 U10906 ( .A1(n10896), .A2(n10897), .ZN(n10656) );
  NAND2_X1 U10907 ( .A1(n10665), .A2(n10898), .ZN(n10897) );
  NAND2_X1 U10908 ( .A1(n10662), .A2(n10664), .ZN(n10898) );
  NOR2_X1 U10909 ( .A1(n10425), .A2(n8825), .ZN(n10665) );
  INV_X1 U10910 ( .A(n10899), .ZN(n10896) );
  NOR2_X1 U10911 ( .A1(n10664), .A2(n10662), .ZN(n10899) );
  XNOR2_X1 U10912 ( .A(n10900), .B(n10901), .ZN(n10662) );
  XNOR2_X1 U10913 ( .A(n10902), .B(n10903), .ZN(n10901) );
  NAND2_X1 U10914 ( .A1(n10904), .A2(n10905), .ZN(n10664) );
  NAND2_X1 U10915 ( .A1(n10670), .A2(n10906), .ZN(n10905) );
  NAND2_X1 U10916 ( .A1(n10673), .A2(n10672), .ZN(n10906) );
  XNOR2_X1 U10917 ( .A(n10907), .B(n10908), .ZN(n10670) );
  XOR2_X1 U10918 ( .A(n10909), .B(n10910), .Z(n10908) );
  INV_X1 U10919 ( .A(n10911), .ZN(n10904) );
  NOR2_X1 U10920 ( .A1(n10672), .A2(n10673), .ZN(n10911) );
  NOR2_X1 U10921 ( .A1(n10425), .A2(n8830), .ZN(n10673) );
  NAND2_X1 U10922 ( .A1(n10912), .A2(n10913), .ZN(n10672) );
  NAND2_X1 U10923 ( .A1(n10680), .A2(n10914), .ZN(n10913) );
  NAND2_X1 U10924 ( .A1(n10679), .A2(n10677), .ZN(n10914) );
  NOR2_X1 U10925 ( .A1(n10425), .A2(n8839), .ZN(n10680) );
  INV_X1 U10926 ( .A(n10915), .ZN(n10912) );
  NOR2_X1 U10927 ( .A1(n10677), .A2(n10679), .ZN(n10915) );
  NOR2_X1 U10928 ( .A1(n10916), .A2(n10917), .ZN(n10679) );
  INV_X1 U10929 ( .A(n10918), .ZN(n10917) );
  NAND2_X1 U10930 ( .A1(n10709), .A2(n10919), .ZN(n10918) );
  NAND2_X1 U10931 ( .A1(n10710), .A2(n10708), .ZN(n10919) );
  NOR2_X1 U10932 ( .A1(n10425), .A2(n8844), .ZN(n10709) );
  NOR2_X1 U10933 ( .A1(n10708), .A2(n10710), .ZN(n10916) );
  NOR2_X1 U10934 ( .A1(n10920), .A2(n10921), .ZN(n10710) );
  INV_X1 U10935 ( .A(n10922), .ZN(n10921) );
  NAND2_X1 U10936 ( .A1(n10703), .A2(n10923), .ZN(n10922) );
  NAND2_X1 U10937 ( .A1(n10924), .A2(n10705), .ZN(n10923) );
  NOR2_X1 U10938 ( .A1(n10425), .A2(n9161), .ZN(n10703) );
  NOR2_X1 U10939 ( .A1(n10705), .A2(n10924), .ZN(n10920) );
  INV_X1 U10940 ( .A(n10706), .ZN(n10924) );
  NAND2_X1 U10941 ( .A1(n10925), .A2(n10926), .ZN(n10706) );
  NAND2_X1 U10942 ( .A1(b_21_), .A2(n10927), .ZN(n10926) );
  NAND2_X1 U10943 ( .A1(n8358), .A2(n10928), .ZN(n10927) );
  NAND2_X1 U10944 ( .A1(a_31_), .A2(n10701), .ZN(n10928) );
  NAND2_X1 U10945 ( .A1(b_22_), .A2(n10929), .ZN(n10925) );
  NAND2_X1 U10946 ( .A1(n8362), .A2(n10930), .ZN(n10929) );
  NAND2_X1 U10947 ( .A1(a_30_), .A2(n10931), .ZN(n10930) );
  NAND2_X1 U10948 ( .A1(n10702), .A2(b_22_), .ZN(n10705) );
  NOR2_X1 U10949 ( .A1(n9170), .A2(n10425), .ZN(n10702) );
  XOR2_X1 U10950 ( .A(n10932), .B(n10933), .Z(n10708) );
  XOR2_X1 U10951 ( .A(n10934), .B(n10935), .Z(n10933) );
  XOR2_X1 U10952 ( .A(n10936), .B(n10937), .Z(n10677) );
  XNOR2_X1 U10953 ( .A(n10938), .B(n10939), .ZN(n10936) );
  XNOR2_X1 U10954 ( .A(n10940), .B(n10941), .ZN(n10655) );
  XNOR2_X1 U10955 ( .A(n10942), .B(n10943), .ZN(n10941) );
  XNOR2_X1 U10956 ( .A(n10944), .B(n10945), .ZN(n10580) );
  NAND2_X1 U10957 ( .A1(n10946), .A2(n10947), .ZN(n10944) );
  XNOR2_X1 U10958 ( .A(n10948), .B(n10949), .ZN(n10712) );
  XOR2_X1 U10959 ( .A(n10950), .B(n10951), .Z(n10949) );
  NAND2_X1 U10960 ( .A1(b_22_), .A2(a_14_), .ZN(n10951) );
  XNOR2_X1 U10961 ( .A(n10952), .B(n10953), .ZN(n10715) );
  NAND2_X1 U10962 ( .A1(n10954), .A2(n10955), .ZN(n10952) );
  XOR2_X1 U10963 ( .A(n10956), .B(n10957), .Z(n10556) );
  XOR2_X1 U10964 ( .A(n10958), .B(n10959), .Z(n10956) );
  NOR2_X1 U10965 ( .A1(n8750), .A2(n10701), .ZN(n10959) );
  INV_X1 U10966 ( .A(n10960), .ZN(n10800) );
  NOR2_X1 U10967 ( .A1(n10722), .A2(n10719), .ZN(n10960) );
  XOR2_X1 U10968 ( .A(n10961), .B(n10962), .Z(n10719) );
  NAND2_X1 U10969 ( .A1(n10963), .A2(n10964), .ZN(n10961) );
  NAND2_X1 U10970 ( .A1(b_23_), .A2(a_10_), .ZN(n10722) );
  XNOR2_X1 U10971 ( .A(n10965), .B(n10966), .ZN(n10724) );
  NAND2_X1 U10972 ( .A1(n10967), .A2(n10968), .ZN(n10965) );
  XNOR2_X1 U10973 ( .A(n10969), .B(n10970), .ZN(n10541) );
  NAND2_X1 U10974 ( .A1(n10971), .A2(n10972), .ZN(n10969) );
  XNOR2_X1 U10975 ( .A(n10973), .B(n10974), .ZN(n10728) );
  NAND2_X1 U10976 ( .A1(n10975), .A2(n10976), .ZN(n10973) );
  XNOR2_X1 U10977 ( .A(n10977), .B(n10978), .ZN(n10731) );
  NAND2_X1 U10978 ( .A1(n10979), .A2(n10980), .ZN(n10977) );
  XOR2_X1 U10979 ( .A(n10981), .B(n10982), .Z(n10736) );
  XOR2_X1 U10980 ( .A(n10983), .B(n10984), .Z(n10981) );
  NOR2_X1 U10981 ( .A1(n8480), .A2(n10701), .ZN(n10984) );
  XNOR2_X1 U10982 ( .A(n10985), .B(n10986), .ZN(n10521) );
  NAND2_X1 U10983 ( .A1(n10987), .A2(n10988), .ZN(n10985) );
  NAND2_X1 U10984 ( .A1(n10989), .A2(n10990), .ZN(n8553) );
  NAND2_X1 U10985 ( .A1(n8658), .A2(n8657), .ZN(n10990) );
  NAND2_X1 U10986 ( .A1(n10991), .A2(n8658), .ZN(n8552) );
  XNOR2_X1 U10987 ( .A(n10992), .B(n10993), .ZN(n8658) );
  NAND2_X1 U10988 ( .A1(n10994), .A2(n10995), .ZN(n10992) );
  NOR2_X1 U10989 ( .A1(n10996), .A2(n10989), .ZN(n10991) );
  XNOR2_X1 U10990 ( .A(n8649), .B(n8648), .ZN(n10989) );
  INV_X1 U10991 ( .A(n8657), .ZN(n10996) );
  NAND2_X1 U10992 ( .A1(n10997), .A2(n10998), .ZN(n8657) );
  INV_X1 U10993 ( .A(n10999), .ZN(n10998) );
  NOR2_X1 U10994 ( .A1(n10495), .A2(n11000), .ZN(n10999) );
  NOR2_X1 U10995 ( .A1(n10492), .A2(n10494), .ZN(n11000) );
  NAND2_X1 U10996 ( .A1(b_22_), .A2(a_0_), .ZN(n10495) );
  NAND2_X1 U10997 ( .A1(n10492), .A2(n10494), .ZN(n10997) );
  NAND2_X1 U10998 ( .A1(n11001), .A2(n11002), .ZN(n10494) );
  NAND2_X1 U10999 ( .A1(n10747), .A2(n11003), .ZN(n11002) );
  NAND2_X1 U11000 ( .A1(n10744), .A2(n10746), .ZN(n11003) );
  NOR2_X1 U11001 ( .A1(n10701), .A2(n8502), .ZN(n10747) );
  INV_X1 U11002 ( .A(n11004), .ZN(n11001) );
  NOR2_X1 U11003 ( .A1(n10744), .A2(n10746), .ZN(n11004) );
  NAND2_X1 U11004 ( .A1(n11005), .A2(n11006), .ZN(n10746) );
  NAND2_X1 U11005 ( .A1(n10755), .A2(n11007), .ZN(n11006) );
  NAND2_X1 U11006 ( .A1(n10758), .A2(n10757), .ZN(n11007) );
  XOR2_X1 U11007 ( .A(n11008), .B(n11009), .Z(n10755) );
  NAND2_X1 U11008 ( .A1(n11010), .A2(n11011), .ZN(n11008) );
  INV_X1 U11009 ( .A(n11012), .ZN(n11005) );
  NOR2_X1 U11010 ( .A1(n10757), .A2(n10758), .ZN(n11012) );
  NOR2_X1 U11011 ( .A1(n10701), .A2(n8497), .ZN(n10758) );
  NAND2_X1 U11012 ( .A1(n10765), .A2(n11013), .ZN(n10757) );
  NAND2_X1 U11013 ( .A1(n10764), .A2(n10766), .ZN(n11013) );
  NAND2_X1 U11014 ( .A1(n11014), .A2(n11015), .ZN(n10766) );
  INV_X1 U11015 ( .A(n11016), .ZN(n11015) );
  NAND2_X1 U11016 ( .A1(b_22_), .A2(a_3_), .ZN(n11014) );
  XOR2_X1 U11017 ( .A(n11017), .B(n11018), .Z(n10764) );
  XNOR2_X1 U11018 ( .A(n11019), .B(n11020), .ZN(n11018) );
  NAND2_X1 U11019 ( .A1(n11016), .A2(a_3_), .ZN(n10765) );
  NOR2_X1 U11020 ( .A1(n11021), .A2(n11022), .ZN(n11016) );
  INV_X1 U11021 ( .A(n11023), .ZN(n11022) );
  NAND2_X1 U11022 ( .A1(n10771), .A2(n11024), .ZN(n11023) );
  NAND2_X1 U11023 ( .A1(n10774), .A2(n10773), .ZN(n11024) );
  XOR2_X1 U11024 ( .A(n11025), .B(n11026), .Z(n10771) );
  NAND2_X1 U11025 ( .A1(n11027), .A2(n11028), .ZN(n11025) );
  NOR2_X1 U11026 ( .A1(n10773), .A2(n10774), .ZN(n11021) );
  NOR2_X1 U11027 ( .A1(n10701), .A2(n8712), .ZN(n10774) );
  NAND2_X1 U11028 ( .A1(n10987), .A2(n11029), .ZN(n10773) );
  NAND2_X1 U11029 ( .A1(n10986), .A2(n10988), .ZN(n11029) );
  NAND2_X1 U11030 ( .A1(n11030), .A2(n11031), .ZN(n10988) );
  NAND2_X1 U11031 ( .A1(b_22_), .A2(a_5_), .ZN(n11031) );
  INV_X1 U11032 ( .A(n11032), .ZN(n11030) );
  XOR2_X1 U11033 ( .A(n11033), .B(n11034), .Z(n10986) );
  XNOR2_X1 U11034 ( .A(n11035), .B(n11036), .ZN(n11034) );
  NAND2_X1 U11035 ( .A1(a_5_), .A2(n11032), .ZN(n10987) );
  NAND2_X1 U11036 ( .A1(n11037), .A2(n11038), .ZN(n11032) );
  NAND2_X1 U11037 ( .A1(n11039), .A2(b_22_), .ZN(n11038) );
  NOR2_X1 U11038 ( .A1(n11040), .A2(n8480), .ZN(n11039) );
  NOR2_X1 U11039 ( .A1(n10982), .A2(n10983), .ZN(n11040) );
  NAND2_X1 U11040 ( .A1(n10982), .A2(n10983), .ZN(n11037) );
  NAND2_X1 U11041 ( .A1(n10979), .A2(n11041), .ZN(n10983) );
  NAND2_X1 U11042 ( .A1(n10978), .A2(n10980), .ZN(n11041) );
  NAND2_X1 U11043 ( .A1(n11042), .A2(n11043), .ZN(n10980) );
  NAND2_X1 U11044 ( .A1(b_22_), .A2(a_7_), .ZN(n11043) );
  INV_X1 U11045 ( .A(n11044), .ZN(n11042) );
  XNOR2_X1 U11046 ( .A(n11045), .B(n11046), .ZN(n10978) );
  XOR2_X1 U11047 ( .A(n11047), .B(n11048), .Z(n11045) );
  NAND2_X1 U11048 ( .A1(a_7_), .A2(n11044), .ZN(n10979) );
  NAND2_X1 U11049 ( .A1(n10975), .A2(n11049), .ZN(n11044) );
  NAND2_X1 U11050 ( .A1(n10974), .A2(n10976), .ZN(n11049) );
  NAND2_X1 U11051 ( .A1(n11050), .A2(n11051), .ZN(n10976) );
  NAND2_X1 U11052 ( .A1(b_22_), .A2(a_8_), .ZN(n11051) );
  INV_X1 U11053 ( .A(n11052), .ZN(n11050) );
  XNOR2_X1 U11054 ( .A(n11053), .B(n11054), .ZN(n10974) );
  NAND2_X1 U11055 ( .A1(n11055), .A2(n11056), .ZN(n11053) );
  NAND2_X1 U11056 ( .A1(a_8_), .A2(n11052), .ZN(n10975) );
  NAND2_X1 U11057 ( .A1(n10971), .A2(n11057), .ZN(n11052) );
  NAND2_X1 U11058 ( .A1(n10970), .A2(n10972), .ZN(n11057) );
  NAND2_X1 U11059 ( .A1(n11058), .A2(n11059), .ZN(n10972) );
  NAND2_X1 U11060 ( .A1(b_22_), .A2(a_9_), .ZN(n11059) );
  INV_X1 U11061 ( .A(n11060), .ZN(n11058) );
  XOR2_X1 U11062 ( .A(n11061), .B(n11062), .Z(n10970) );
  XOR2_X1 U11063 ( .A(n11063), .B(n11064), .Z(n11061) );
  NOR2_X1 U11064 ( .A1(n8741), .A2(n10931), .ZN(n11064) );
  NAND2_X1 U11065 ( .A1(a_9_), .A2(n11060), .ZN(n10971) );
  NAND2_X1 U11066 ( .A1(n10967), .A2(n11065), .ZN(n11060) );
  NAND2_X1 U11067 ( .A1(n10966), .A2(n10968), .ZN(n11065) );
  NAND2_X1 U11068 ( .A1(n11066), .A2(n11067), .ZN(n10968) );
  NAND2_X1 U11069 ( .A1(b_22_), .A2(a_10_), .ZN(n11067) );
  INV_X1 U11070 ( .A(n11068), .ZN(n11066) );
  XOR2_X1 U11071 ( .A(n11069), .B(n11070), .Z(n10966) );
  XOR2_X1 U11072 ( .A(n11071), .B(n11072), .Z(n11069) );
  NOR2_X1 U11073 ( .A1(n8452), .A2(n10931), .ZN(n11072) );
  NAND2_X1 U11074 ( .A1(a_10_), .A2(n11068), .ZN(n10967) );
  NAND2_X1 U11075 ( .A1(n10963), .A2(n11073), .ZN(n11068) );
  NAND2_X1 U11076 ( .A1(n10962), .A2(n10964), .ZN(n11073) );
  NAND2_X1 U11077 ( .A1(n11074), .A2(n11075), .ZN(n10964) );
  NAND2_X1 U11078 ( .A1(b_22_), .A2(a_11_), .ZN(n11075) );
  INV_X1 U11079 ( .A(n11076), .ZN(n11074) );
  XNOR2_X1 U11080 ( .A(n11077), .B(n11078), .ZN(n10962) );
  NAND2_X1 U11081 ( .A1(n11079), .A2(n11080), .ZN(n11077) );
  NAND2_X1 U11082 ( .A1(a_11_), .A2(n11076), .ZN(n10963) );
  NAND2_X1 U11083 ( .A1(n11081), .A2(n11082), .ZN(n11076) );
  NAND2_X1 U11084 ( .A1(n11083), .A2(b_22_), .ZN(n11082) );
  NOR2_X1 U11085 ( .A1(n11084), .A2(n8750), .ZN(n11083) );
  NOR2_X1 U11086 ( .A1(n10957), .A2(n10958), .ZN(n11084) );
  NAND2_X1 U11087 ( .A1(n10957), .A2(n10958), .ZN(n11081) );
  NAND2_X1 U11088 ( .A1(n10954), .A2(n11085), .ZN(n10958) );
  NAND2_X1 U11089 ( .A1(n10953), .A2(n10955), .ZN(n11085) );
  NAND2_X1 U11090 ( .A1(n11086), .A2(n11087), .ZN(n10955) );
  NAND2_X1 U11091 ( .A1(b_22_), .A2(a_13_), .ZN(n11087) );
  INV_X1 U11092 ( .A(n11088), .ZN(n11086) );
  XNOR2_X1 U11093 ( .A(n11089), .B(n11090), .ZN(n10953) );
  XOR2_X1 U11094 ( .A(n11091), .B(n11092), .Z(n11090) );
  NAND2_X1 U11095 ( .A1(b_21_), .A2(a_14_), .ZN(n11092) );
  NAND2_X1 U11096 ( .A1(a_13_), .A2(n11088), .ZN(n10954) );
  NAND2_X1 U11097 ( .A1(n11093), .A2(n11094), .ZN(n11088) );
  NAND2_X1 U11098 ( .A1(n11095), .A2(b_22_), .ZN(n11094) );
  NOR2_X1 U11099 ( .A1(n11096), .A2(n8438), .ZN(n11095) );
  NOR2_X1 U11100 ( .A1(n10948), .A2(n10950), .ZN(n11096) );
  NAND2_X1 U11101 ( .A1(n10948), .A2(n10950), .ZN(n11093) );
  NAND2_X1 U11102 ( .A1(n11097), .A2(n11098), .ZN(n10950) );
  NAND2_X1 U11103 ( .A1(n11099), .A2(b_22_), .ZN(n11098) );
  NOR2_X1 U11104 ( .A1(n11100), .A2(n8763), .ZN(n11099) );
  NOR2_X1 U11105 ( .A1(n10820), .A2(n10821), .ZN(n11100) );
  NAND2_X1 U11106 ( .A1(n10820), .A2(n10821), .ZN(n11097) );
  NAND2_X1 U11107 ( .A1(n10946), .A2(n11101), .ZN(n10821) );
  NAND2_X1 U11108 ( .A1(n10945), .A2(n10947), .ZN(n11101) );
  NAND2_X1 U11109 ( .A1(n11102), .A2(n11103), .ZN(n10947) );
  NAND2_X1 U11110 ( .A1(b_22_), .A2(a_16_), .ZN(n11103) );
  INV_X1 U11111 ( .A(n11104), .ZN(n11102) );
  XOR2_X1 U11112 ( .A(n11105), .B(n11106), .Z(n10945) );
  XNOR2_X1 U11113 ( .A(n11107), .B(n11108), .ZN(n11106) );
  NAND2_X1 U11114 ( .A1(b_21_), .A2(a_17_), .ZN(n11108) );
  NAND2_X1 U11115 ( .A1(a_16_), .A2(n11104), .ZN(n10946) );
  NAND2_X1 U11116 ( .A1(n10833), .A2(n11109), .ZN(n11104) );
  NAND2_X1 U11117 ( .A1(n10832), .A2(n10834), .ZN(n11109) );
  NAND2_X1 U11118 ( .A1(n11110), .A2(n11111), .ZN(n10834) );
  NAND2_X1 U11119 ( .A1(b_22_), .A2(a_17_), .ZN(n11111) );
  INV_X1 U11120 ( .A(n11112), .ZN(n11110) );
  XOR2_X1 U11121 ( .A(n11113), .B(n11114), .Z(n10832) );
  XNOR2_X1 U11122 ( .A(n11115), .B(n11116), .ZN(n11114) );
  NAND2_X1 U11123 ( .A1(a_17_), .A2(n11112), .ZN(n10833) );
  NAND2_X1 U11124 ( .A1(n10841), .A2(n11117), .ZN(n11112) );
  NAND2_X1 U11125 ( .A1(n10840), .A2(n10842), .ZN(n11117) );
  NAND2_X1 U11126 ( .A1(n11118), .A2(n11119), .ZN(n10842) );
  NAND2_X1 U11127 ( .A1(b_22_), .A2(a_18_), .ZN(n11119) );
  INV_X1 U11128 ( .A(n11120), .ZN(n11118) );
  XOR2_X1 U11129 ( .A(n11121), .B(n11122), .Z(n10840) );
  XNOR2_X1 U11130 ( .A(n11123), .B(n11124), .ZN(n11122) );
  NAND2_X1 U11131 ( .A1(b_21_), .A2(a_19_), .ZN(n11124) );
  NAND2_X1 U11132 ( .A1(a_18_), .A2(n11120), .ZN(n10841) );
  NAND2_X1 U11133 ( .A1(n11125), .A2(n11126), .ZN(n11120) );
  NAND2_X1 U11134 ( .A1(n11127), .A2(b_22_), .ZN(n11126) );
  NOR2_X1 U11135 ( .A1(n11128), .A2(n8881), .ZN(n11127) );
  NOR2_X1 U11136 ( .A1(n10848), .A2(n10849), .ZN(n11128) );
  NAND2_X1 U11137 ( .A1(n10848), .A2(n10849), .ZN(n11125) );
  NAND2_X1 U11138 ( .A1(n10857), .A2(n11129), .ZN(n10849) );
  NAND2_X1 U11139 ( .A1(n10856), .A2(n10858), .ZN(n11129) );
  NAND2_X1 U11140 ( .A1(n11130), .A2(n11131), .ZN(n10858) );
  NAND2_X1 U11141 ( .A1(b_22_), .A2(a_20_), .ZN(n11131) );
  INV_X1 U11142 ( .A(n11132), .ZN(n11130) );
  XOR2_X1 U11143 ( .A(n11133), .B(n11134), .Z(n10856) );
  XOR2_X1 U11144 ( .A(n11135), .B(n11136), .Z(n11133) );
  NAND2_X1 U11145 ( .A1(a_20_), .A2(n11132), .ZN(n10857) );
  NAND2_X1 U11146 ( .A1(n10865), .A2(n11137), .ZN(n11132) );
  NAND2_X1 U11147 ( .A1(n10864), .A2(n10866), .ZN(n11137) );
  NAND2_X1 U11148 ( .A1(n11138), .A2(n11139), .ZN(n10866) );
  NAND2_X1 U11149 ( .A1(b_22_), .A2(a_21_), .ZN(n11138) );
  XNOR2_X1 U11150 ( .A(n11140), .B(n11141), .ZN(n10864) );
  NAND2_X1 U11151 ( .A1(n11142), .A2(n11143), .ZN(n11140) );
  NAND2_X1 U11152 ( .A1(n11144), .A2(a_21_), .ZN(n10865) );
  INV_X1 U11153 ( .A(n11139), .ZN(n11144) );
  NAND2_X1 U11154 ( .A1(n11145), .A2(n11146), .ZN(n11139) );
  NAND2_X1 U11155 ( .A1(n11147), .A2(n10874), .ZN(n11146) );
  NAND2_X1 U11156 ( .A1(n10872), .A2(n10873), .ZN(n11147) );
  INV_X1 U11157 ( .A(n11148), .ZN(n11145) );
  NOR2_X1 U11158 ( .A1(n10873), .A2(n10872), .ZN(n11148) );
  XOR2_X1 U11159 ( .A(n11149), .B(n11150), .Z(n10872) );
  XOR2_X1 U11160 ( .A(n11151), .B(n11152), .Z(n11149) );
  NOR2_X1 U11161 ( .A1(n8812), .A2(n10931), .ZN(n11152) );
  NAND2_X1 U11162 ( .A1(n11153), .A2(n11154), .ZN(n10873) );
  NAND2_X1 U11163 ( .A1(n11155), .A2(b_22_), .ZN(n11154) );
  NOR2_X1 U11164 ( .A1(n11156), .A2(n8812), .ZN(n11155) );
  NOR2_X1 U11165 ( .A1(n10879), .A2(n10880), .ZN(n11156) );
  NAND2_X1 U11166 ( .A1(n10879), .A2(n10880), .ZN(n11153) );
  NAND2_X1 U11167 ( .A1(n11157), .A2(n11158), .ZN(n10880) );
  NAND2_X1 U11168 ( .A1(n10891), .A2(n11159), .ZN(n11158) );
  INV_X1 U11169 ( .A(n11160), .ZN(n11159) );
  NOR2_X1 U11170 ( .A1(n10890), .A2(n10889), .ZN(n11160) );
  NOR2_X1 U11171 ( .A1(n10701), .A2(n9131), .ZN(n10891) );
  NAND2_X1 U11172 ( .A1(n10889), .A2(n10890), .ZN(n11157) );
  NAND2_X1 U11173 ( .A1(n11161), .A2(n11162), .ZN(n10890) );
  NAND2_X1 U11174 ( .A1(n10943), .A2(n11163), .ZN(n11162) );
  NAND2_X1 U11175 ( .A1(n10940), .A2(n10942), .ZN(n11163) );
  NOR2_X1 U11176 ( .A1(n10701), .A2(n8825), .ZN(n10943) );
  INV_X1 U11177 ( .A(n11164), .ZN(n11161) );
  NOR2_X1 U11178 ( .A1(n10942), .A2(n10940), .ZN(n11164) );
  XNOR2_X1 U11179 ( .A(n11165), .B(n11166), .ZN(n10940) );
  XNOR2_X1 U11180 ( .A(n11167), .B(n11168), .ZN(n11166) );
  NAND2_X1 U11181 ( .A1(n11169), .A2(n11170), .ZN(n10942) );
  NAND2_X1 U11182 ( .A1(n10900), .A2(n11171), .ZN(n11170) );
  NAND2_X1 U11183 ( .A1(n10903), .A2(n10902), .ZN(n11171) );
  XNOR2_X1 U11184 ( .A(n11172), .B(n11173), .ZN(n10900) );
  XOR2_X1 U11185 ( .A(n11174), .B(n11175), .Z(n11173) );
  INV_X1 U11186 ( .A(n11176), .ZN(n11169) );
  NOR2_X1 U11187 ( .A1(n10902), .A2(n10903), .ZN(n11176) );
  NOR2_X1 U11188 ( .A1(n10701), .A2(n8830), .ZN(n10903) );
  NAND2_X1 U11189 ( .A1(n11177), .A2(n11178), .ZN(n10902) );
  NAND2_X1 U11190 ( .A1(n10910), .A2(n11179), .ZN(n11178) );
  NAND2_X1 U11191 ( .A1(n10909), .A2(n10907), .ZN(n11179) );
  NOR2_X1 U11192 ( .A1(n10701), .A2(n8839), .ZN(n10910) );
  INV_X1 U11193 ( .A(n11180), .ZN(n11177) );
  NOR2_X1 U11194 ( .A1(n10907), .A2(n10909), .ZN(n11180) );
  NOR2_X1 U11195 ( .A1(n11181), .A2(n11182), .ZN(n10909) );
  INV_X1 U11196 ( .A(n11183), .ZN(n11182) );
  NAND2_X1 U11197 ( .A1(n10938), .A2(n11184), .ZN(n11183) );
  NAND2_X1 U11198 ( .A1(n10939), .A2(n10937), .ZN(n11184) );
  NOR2_X1 U11199 ( .A1(n10701), .A2(n8844), .ZN(n10938) );
  NOR2_X1 U11200 ( .A1(n10937), .A2(n10939), .ZN(n11181) );
  NOR2_X1 U11201 ( .A1(n11185), .A2(n11186), .ZN(n10939) );
  INV_X1 U11202 ( .A(n11187), .ZN(n11186) );
  NAND2_X1 U11203 ( .A1(n10932), .A2(n11188), .ZN(n11187) );
  NAND2_X1 U11204 ( .A1(n11189), .A2(n10934), .ZN(n11188) );
  NOR2_X1 U11205 ( .A1(n10701), .A2(n9161), .ZN(n10932) );
  NOR2_X1 U11206 ( .A1(n10934), .A2(n11189), .ZN(n11185) );
  INV_X1 U11207 ( .A(n10935), .ZN(n11189) );
  NAND2_X1 U11208 ( .A1(n11190), .A2(n11191), .ZN(n10935) );
  NAND2_X1 U11209 ( .A1(b_20_), .A2(n11192), .ZN(n11191) );
  NAND2_X1 U11210 ( .A1(n8358), .A2(n11193), .ZN(n11192) );
  NAND2_X1 U11211 ( .A1(a_31_), .A2(n10931), .ZN(n11193) );
  NAND2_X1 U11212 ( .A1(b_21_), .A2(n11194), .ZN(n11190) );
  NAND2_X1 U11213 ( .A1(n8362), .A2(n11195), .ZN(n11194) );
  NAND2_X1 U11214 ( .A1(a_30_), .A2(n11196), .ZN(n11195) );
  NAND2_X1 U11215 ( .A1(n11197), .A2(b_22_), .ZN(n10934) );
  NOR2_X1 U11216 ( .A1(n9170), .A2(n10931), .ZN(n11197) );
  XOR2_X1 U11217 ( .A(n11198), .B(n11199), .Z(n10937) );
  XOR2_X1 U11218 ( .A(n11200), .B(n11201), .Z(n11199) );
  XOR2_X1 U11219 ( .A(n11202), .B(n11203), .Z(n10907) );
  XNOR2_X1 U11220 ( .A(n11204), .B(n11205), .ZN(n11202) );
  XNOR2_X1 U11221 ( .A(n11206), .B(n11207), .ZN(n10889) );
  XNOR2_X1 U11222 ( .A(n11208), .B(n11209), .ZN(n11207) );
  XOR2_X1 U11223 ( .A(n11210), .B(n11211), .Z(n10879) );
  XOR2_X1 U11224 ( .A(n11212), .B(n11213), .Z(n11210) );
  XOR2_X1 U11225 ( .A(n11214), .B(n11215), .Z(n10848) );
  XNOR2_X1 U11226 ( .A(n11216), .B(n11217), .ZN(n11215) );
  XOR2_X1 U11227 ( .A(n11218), .B(n11219), .Z(n10820) );
  XOR2_X1 U11228 ( .A(n11220), .B(n11221), .Z(n11218) );
  NOR2_X1 U11229 ( .A1(n8768), .A2(n10931), .ZN(n11221) );
  XNOR2_X1 U11230 ( .A(n11222), .B(n11223), .ZN(n10948) );
  XOR2_X1 U11231 ( .A(n11224), .B(n11225), .Z(n11223) );
  NAND2_X1 U11232 ( .A1(b_21_), .A2(a_15_), .ZN(n11225) );
  XNOR2_X1 U11233 ( .A(n11226), .B(n11227), .ZN(n10957) );
  NAND2_X1 U11234 ( .A1(n11228), .A2(n11229), .ZN(n11226) );
  XNOR2_X1 U11235 ( .A(n11230), .B(n11231), .ZN(n10982) );
  XNOR2_X1 U11236 ( .A(n11232), .B(n11233), .ZN(n11230) );
  NOR2_X1 U11237 ( .A1(n8726), .A2(n10931), .ZN(n11233) );
  XNOR2_X1 U11238 ( .A(n11234), .B(n11235), .ZN(n10744) );
  XNOR2_X1 U11239 ( .A(n11236), .B(n11237), .ZN(n11235) );
  XNOR2_X1 U11240 ( .A(n11238), .B(n11239), .ZN(n10492) );
  NAND2_X1 U11241 ( .A1(n11240), .A2(n11241), .ZN(n11238) );
  INV_X1 U11242 ( .A(n11242), .ZN(n8556) );
  NOR2_X1 U11243 ( .A1(n11243), .A2(n11244), .ZN(n11242) );
  NAND2_X1 U11244 ( .A1(n8644), .A2(n8649), .ZN(n11244) );
  NAND2_X1 U11245 ( .A1(n10994), .A2(n11245), .ZN(n8649) );
  NAND2_X1 U11246 ( .A1(n10993), .A2(n10995), .ZN(n11245) );
  NAND2_X1 U11247 ( .A1(n11246), .A2(n11247), .ZN(n10995) );
  NAND2_X1 U11248 ( .A1(b_21_), .A2(a_0_), .ZN(n11247) );
  INV_X1 U11249 ( .A(n11248), .ZN(n11246) );
  XNOR2_X1 U11250 ( .A(n11249), .B(n11250), .ZN(n10993) );
  XOR2_X1 U11251 ( .A(n11251), .B(n11252), .Z(n11249) );
  NAND2_X1 U11252 ( .A1(a_0_), .A2(n11248), .ZN(n10994) );
  NAND2_X1 U11253 ( .A1(n11240), .A2(n11253), .ZN(n11248) );
  NAND2_X1 U11254 ( .A1(n11239), .A2(n11241), .ZN(n11253) );
  NAND2_X1 U11255 ( .A1(n11254), .A2(n11255), .ZN(n11241) );
  INV_X1 U11256 ( .A(n11256), .ZN(n11255) );
  NAND2_X1 U11257 ( .A1(b_21_), .A2(a_1_), .ZN(n11254) );
  XNOR2_X1 U11258 ( .A(n11257), .B(n11258), .ZN(n11239) );
  NAND2_X1 U11259 ( .A1(n11259), .A2(n11260), .ZN(n11257) );
  NAND2_X1 U11260 ( .A1(n11256), .A2(a_1_), .ZN(n11240) );
  NOR2_X1 U11261 ( .A1(n11261), .A2(n11262), .ZN(n11256) );
  INV_X1 U11262 ( .A(n11263), .ZN(n11262) );
  NAND2_X1 U11263 ( .A1(n11234), .A2(n11264), .ZN(n11263) );
  NAND2_X1 U11264 ( .A1(n11237), .A2(n11236), .ZN(n11264) );
  XNOR2_X1 U11265 ( .A(n11265), .B(n11266), .ZN(n11234) );
  XNOR2_X1 U11266 ( .A(n11267), .B(n11268), .ZN(n11266) );
  NOR2_X1 U11267 ( .A1(n11236), .A2(n11237), .ZN(n11261) );
  NOR2_X1 U11268 ( .A1(n10931), .A2(n8497), .ZN(n11237) );
  NAND2_X1 U11269 ( .A1(n11010), .A2(n11269), .ZN(n11236) );
  NAND2_X1 U11270 ( .A1(n11009), .A2(n11011), .ZN(n11269) );
  NAND2_X1 U11271 ( .A1(n11270), .A2(n11271), .ZN(n11011) );
  INV_X1 U11272 ( .A(n11272), .ZN(n11271) );
  NAND2_X1 U11273 ( .A1(b_21_), .A2(a_3_), .ZN(n11270) );
  XNOR2_X1 U11274 ( .A(n11273), .B(n11274), .ZN(n11009) );
  NAND2_X1 U11275 ( .A1(n11275), .A2(n11276), .ZN(n11273) );
  NAND2_X1 U11276 ( .A1(n11272), .A2(a_3_), .ZN(n11010) );
  NOR2_X1 U11277 ( .A1(n11277), .A2(n11278), .ZN(n11272) );
  INV_X1 U11278 ( .A(n11279), .ZN(n11278) );
  NAND2_X1 U11279 ( .A1(n11017), .A2(n11280), .ZN(n11279) );
  NAND2_X1 U11280 ( .A1(n11020), .A2(n11019), .ZN(n11280) );
  XNOR2_X1 U11281 ( .A(n11281), .B(n11282), .ZN(n11017) );
  XNOR2_X1 U11282 ( .A(n11283), .B(n11284), .ZN(n11282) );
  NOR2_X1 U11283 ( .A1(n11019), .A2(n11020), .ZN(n11277) );
  NOR2_X1 U11284 ( .A1(n10931), .A2(n8712), .ZN(n11020) );
  NAND2_X1 U11285 ( .A1(n11027), .A2(n11285), .ZN(n11019) );
  NAND2_X1 U11286 ( .A1(n11026), .A2(n11028), .ZN(n11285) );
  NAND2_X1 U11287 ( .A1(n11286), .A2(n11287), .ZN(n11028) );
  INV_X1 U11288 ( .A(n11288), .ZN(n11287) );
  NAND2_X1 U11289 ( .A1(b_21_), .A2(a_5_), .ZN(n11286) );
  XNOR2_X1 U11290 ( .A(n11289), .B(n11290), .ZN(n11026) );
  NAND2_X1 U11291 ( .A1(n11291), .A2(n11292), .ZN(n11289) );
  NAND2_X1 U11292 ( .A1(n11288), .A2(a_5_), .ZN(n11027) );
  NOR2_X1 U11293 ( .A1(n11293), .A2(n11294), .ZN(n11288) );
  INV_X1 U11294 ( .A(n11295), .ZN(n11294) );
  NAND2_X1 U11295 ( .A1(n11033), .A2(n11296), .ZN(n11295) );
  NAND2_X1 U11296 ( .A1(n11036), .A2(n11035), .ZN(n11296) );
  XOR2_X1 U11297 ( .A(n11297), .B(n11298), .Z(n11033) );
  XOR2_X1 U11298 ( .A(n11299), .B(n11300), .Z(n11297) );
  NOR2_X1 U11299 ( .A1(n11035), .A2(n11036), .ZN(n11293) );
  NOR2_X1 U11300 ( .A1(n10931), .A2(n8480), .ZN(n11036) );
  NAND2_X1 U11301 ( .A1(n11301), .A2(n11302), .ZN(n11035) );
  NAND2_X1 U11302 ( .A1(n11303), .A2(b_21_), .ZN(n11302) );
  NOR2_X1 U11303 ( .A1(n11304), .A2(n8726), .ZN(n11303) );
  NOR2_X1 U11304 ( .A1(n11232), .A2(n11231), .ZN(n11304) );
  NAND2_X1 U11305 ( .A1(n11232), .A2(n11231), .ZN(n11301) );
  XNOR2_X1 U11306 ( .A(n11305), .B(n11306), .ZN(n11231) );
  NAND2_X1 U11307 ( .A1(n11307), .A2(n11308), .ZN(n11305) );
  NOR2_X1 U11308 ( .A1(n11309), .A2(n11310), .ZN(n11232) );
  INV_X1 U11309 ( .A(n11311), .ZN(n11310) );
  NAND2_X1 U11310 ( .A1(n11046), .A2(n11312), .ZN(n11311) );
  NAND2_X1 U11311 ( .A1(n11048), .A2(n11047), .ZN(n11312) );
  XOR2_X1 U11312 ( .A(n11313), .B(n11314), .Z(n11046) );
  XOR2_X1 U11313 ( .A(n11315), .B(n11316), .Z(n11314) );
  NAND2_X1 U11314 ( .A1(b_20_), .A2(a_9_), .ZN(n11316) );
  NOR2_X1 U11315 ( .A1(n11047), .A2(n11048), .ZN(n11309) );
  NOR2_X1 U11316 ( .A1(n10931), .A2(n8731), .ZN(n11048) );
  NAND2_X1 U11317 ( .A1(n11055), .A2(n11317), .ZN(n11047) );
  NAND2_X1 U11318 ( .A1(n11054), .A2(n11056), .ZN(n11317) );
  NAND2_X1 U11319 ( .A1(n11318), .A2(n11319), .ZN(n11056) );
  NAND2_X1 U11320 ( .A1(b_21_), .A2(a_9_), .ZN(n11319) );
  INV_X1 U11321 ( .A(n11320), .ZN(n11318) );
  XNOR2_X1 U11322 ( .A(n11321), .B(n11322), .ZN(n11054) );
  XOR2_X1 U11323 ( .A(n11323), .B(n11324), .Z(n11322) );
  NAND2_X1 U11324 ( .A1(b_20_), .A2(a_10_), .ZN(n11324) );
  NAND2_X1 U11325 ( .A1(a_9_), .A2(n11320), .ZN(n11055) );
  NAND2_X1 U11326 ( .A1(n11325), .A2(n11326), .ZN(n11320) );
  NAND2_X1 U11327 ( .A1(n11327), .A2(b_21_), .ZN(n11326) );
  NOR2_X1 U11328 ( .A1(n11328), .A2(n8741), .ZN(n11327) );
  NOR2_X1 U11329 ( .A1(n11062), .A2(n11063), .ZN(n11328) );
  NAND2_X1 U11330 ( .A1(n11062), .A2(n11063), .ZN(n11325) );
  NAND2_X1 U11331 ( .A1(n11329), .A2(n11330), .ZN(n11063) );
  NAND2_X1 U11332 ( .A1(n11331), .A2(b_21_), .ZN(n11330) );
  NOR2_X1 U11333 ( .A1(n11332), .A2(n8452), .ZN(n11331) );
  NOR2_X1 U11334 ( .A1(n11070), .A2(n11071), .ZN(n11332) );
  NAND2_X1 U11335 ( .A1(n11070), .A2(n11071), .ZN(n11329) );
  NAND2_X1 U11336 ( .A1(n11079), .A2(n11333), .ZN(n11071) );
  NAND2_X1 U11337 ( .A1(n11078), .A2(n11080), .ZN(n11333) );
  NAND2_X1 U11338 ( .A1(n11334), .A2(n11335), .ZN(n11080) );
  NAND2_X1 U11339 ( .A1(b_21_), .A2(a_12_), .ZN(n11335) );
  INV_X1 U11340 ( .A(n11336), .ZN(n11334) );
  XNOR2_X1 U11341 ( .A(n11337), .B(n11338), .ZN(n11078) );
  NAND2_X1 U11342 ( .A1(n11339), .A2(n11340), .ZN(n11337) );
  NAND2_X1 U11343 ( .A1(a_12_), .A2(n11336), .ZN(n11079) );
  NAND2_X1 U11344 ( .A1(n11228), .A2(n11341), .ZN(n11336) );
  NAND2_X1 U11345 ( .A1(n11227), .A2(n11229), .ZN(n11341) );
  NAND2_X1 U11346 ( .A1(n11342), .A2(n11343), .ZN(n11229) );
  NAND2_X1 U11347 ( .A1(b_21_), .A2(a_13_), .ZN(n11343) );
  INV_X1 U11348 ( .A(n11344), .ZN(n11342) );
  XNOR2_X1 U11349 ( .A(n11345), .B(n11346), .ZN(n11227) );
  NAND2_X1 U11350 ( .A1(n11347), .A2(n11348), .ZN(n11345) );
  NAND2_X1 U11351 ( .A1(a_13_), .A2(n11344), .ZN(n11228) );
  NAND2_X1 U11352 ( .A1(n11349), .A2(n11350), .ZN(n11344) );
  NAND2_X1 U11353 ( .A1(n11351), .A2(b_21_), .ZN(n11350) );
  NOR2_X1 U11354 ( .A1(n11352), .A2(n8438), .ZN(n11351) );
  NOR2_X1 U11355 ( .A1(n11089), .A2(n11091), .ZN(n11352) );
  NAND2_X1 U11356 ( .A1(n11089), .A2(n11091), .ZN(n11349) );
  NAND2_X1 U11357 ( .A1(n11353), .A2(n11354), .ZN(n11091) );
  NAND2_X1 U11358 ( .A1(n11355), .A2(b_21_), .ZN(n11354) );
  NOR2_X1 U11359 ( .A1(n11356), .A2(n8763), .ZN(n11355) );
  NOR2_X1 U11360 ( .A1(n11222), .A2(n11224), .ZN(n11356) );
  NAND2_X1 U11361 ( .A1(n11222), .A2(n11224), .ZN(n11353) );
  NAND2_X1 U11362 ( .A1(n11357), .A2(n11358), .ZN(n11224) );
  NAND2_X1 U11363 ( .A1(n11359), .A2(b_21_), .ZN(n11358) );
  NOR2_X1 U11364 ( .A1(n11360), .A2(n8768), .ZN(n11359) );
  NOR2_X1 U11365 ( .A1(n11219), .A2(n11220), .ZN(n11360) );
  NAND2_X1 U11366 ( .A1(n11219), .A2(n11220), .ZN(n11357) );
  NAND2_X1 U11367 ( .A1(n11361), .A2(n11362), .ZN(n11220) );
  NAND2_X1 U11368 ( .A1(n11363), .A2(b_21_), .ZN(n11362) );
  NOR2_X1 U11369 ( .A1(n11364), .A2(n8772), .ZN(n11363) );
  NOR2_X1 U11370 ( .A1(n11107), .A2(n11105), .ZN(n11364) );
  NAND2_X1 U11371 ( .A1(n11107), .A2(n11105), .ZN(n11361) );
  XNOR2_X1 U11372 ( .A(n11365), .B(n11366), .ZN(n11105) );
  XOR2_X1 U11373 ( .A(n11367), .B(n11368), .Z(n11366) );
  NAND2_X1 U11374 ( .A1(b_20_), .A2(a_18_), .ZN(n11368) );
  NOR2_X1 U11375 ( .A1(n11369), .A2(n11370), .ZN(n11107) );
  INV_X1 U11376 ( .A(n11371), .ZN(n11370) );
  NAND2_X1 U11377 ( .A1(n11113), .A2(n11372), .ZN(n11371) );
  NAND2_X1 U11378 ( .A1(n11116), .A2(n11115), .ZN(n11372) );
  XNOR2_X1 U11379 ( .A(n11373), .B(n11374), .ZN(n11113) );
  XNOR2_X1 U11380 ( .A(n11375), .B(n11376), .ZN(n11373) );
  NAND2_X1 U11381 ( .A1(b_20_), .A2(a_19_), .ZN(n11375) );
  NOR2_X1 U11382 ( .A1(n11115), .A2(n11116), .ZN(n11369) );
  NOR2_X1 U11383 ( .A1(n10931), .A2(n10616), .ZN(n11116) );
  NAND2_X1 U11384 ( .A1(n11377), .A2(n11378), .ZN(n11115) );
  NAND2_X1 U11385 ( .A1(n11379), .A2(b_21_), .ZN(n11378) );
  NOR2_X1 U11386 ( .A1(n11380), .A2(n8881), .ZN(n11379) );
  NOR2_X1 U11387 ( .A1(n11123), .A2(n11121), .ZN(n11380) );
  NAND2_X1 U11388 ( .A1(n11123), .A2(n11121), .ZN(n11377) );
  XNOR2_X1 U11389 ( .A(n11381), .B(n11382), .ZN(n11121) );
  XOR2_X1 U11390 ( .A(n11383), .B(n11384), .Z(n11382) );
  NOR2_X1 U11391 ( .A1(n11385), .A2(n11386), .ZN(n11123) );
  INV_X1 U11392 ( .A(n11387), .ZN(n11386) );
  NAND2_X1 U11393 ( .A1(n11214), .A2(n11388), .ZN(n11387) );
  NAND2_X1 U11394 ( .A1(n11217), .A2(n11216), .ZN(n11388) );
  XOR2_X1 U11395 ( .A(n11389), .B(n11390), .Z(n11214) );
  NAND2_X1 U11396 ( .A1(n11391), .A2(n11392), .ZN(n11389) );
  NOR2_X1 U11397 ( .A1(n11216), .A2(n11217), .ZN(n11385) );
  NOR2_X1 U11398 ( .A1(n10931), .A2(n10633), .ZN(n11217) );
  NAND2_X1 U11399 ( .A1(n11393), .A2(n11394), .ZN(n11216) );
  NAND2_X1 U11400 ( .A1(n11134), .A2(n11395), .ZN(n11394) );
  INV_X1 U11401 ( .A(n11396), .ZN(n11395) );
  NOR2_X1 U11402 ( .A1(n11135), .A2(n11136), .ZN(n11396) );
  XNOR2_X1 U11403 ( .A(n11397), .B(n11398), .ZN(n11134) );
  NAND2_X1 U11404 ( .A1(n11399), .A2(n11400), .ZN(n11397) );
  NAND2_X1 U11405 ( .A1(n11136), .A2(n11135), .ZN(n11393) );
  NAND2_X1 U11406 ( .A1(n11142), .A2(n11401), .ZN(n11135) );
  NAND2_X1 U11407 ( .A1(n11141), .A2(n11143), .ZN(n11401) );
  NAND2_X1 U11408 ( .A1(n11402), .A2(n11403), .ZN(n11143) );
  NAND2_X1 U11409 ( .A1(b_21_), .A2(a_22_), .ZN(n11403) );
  INV_X1 U11410 ( .A(n11404), .ZN(n11402) );
  XOR2_X1 U11411 ( .A(n11405), .B(n11406), .Z(n11141) );
  XOR2_X1 U11412 ( .A(n11407), .B(n11408), .Z(n11405) );
  NOR2_X1 U11413 ( .A1(n8812), .A2(n11196), .ZN(n11408) );
  NAND2_X1 U11414 ( .A1(a_22_), .A2(n11404), .ZN(n11142) );
  NAND2_X1 U11415 ( .A1(n11409), .A2(n11410), .ZN(n11404) );
  NAND2_X1 U11416 ( .A1(n11411), .A2(b_21_), .ZN(n11410) );
  NOR2_X1 U11417 ( .A1(n11412), .A2(n8812), .ZN(n11411) );
  NOR2_X1 U11418 ( .A1(n11150), .A2(n11151), .ZN(n11412) );
  NAND2_X1 U11419 ( .A1(n11150), .A2(n11151), .ZN(n11409) );
  NAND2_X1 U11420 ( .A1(n11413), .A2(n11414), .ZN(n11151) );
  NAND2_X1 U11421 ( .A1(n11213), .A2(n11415), .ZN(n11414) );
  INV_X1 U11422 ( .A(n11416), .ZN(n11415) );
  NOR2_X1 U11423 ( .A1(n11212), .A2(n11211), .ZN(n11416) );
  NOR2_X1 U11424 ( .A1(n10931), .A2(n9131), .ZN(n11213) );
  NAND2_X1 U11425 ( .A1(n11211), .A2(n11212), .ZN(n11413) );
  NAND2_X1 U11426 ( .A1(n11417), .A2(n11418), .ZN(n11212) );
  NAND2_X1 U11427 ( .A1(n11209), .A2(n11419), .ZN(n11418) );
  NAND2_X1 U11428 ( .A1(n11206), .A2(n11208), .ZN(n11419) );
  NOR2_X1 U11429 ( .A1(n10931), .A2(n8825), .ZN(n11209) );
  INV_X1 U11430 ( .A(n11420), .ZN(n11417) );
  NOR2_X1 U11431 ( .A1(n11208), .A2(n11206), .ZN(n11420) );
  XNOR2_X1 U11432 ( .A(n11421), .B(n11422), .ZN(n11206) );
  XNOR2_X1 U11433 ( .A(n11423), .B(n11424), .ZN(n11422) );
  NAND2_X1 U11434 ( .A1(n11425), .A2(n11426), .ZN(n11208) );
  NAND2_X1 U11435 ( .A1(n11165), .A2(n11427), .ZN(n11426) );
  NAND2_X1 U11436 ( .A1(n11168), .A2(n11167), .ZN(n11427) );
  XNOR2_X1 U11437 ( .A(n11428), .B(n11429), .ZN(n11165) );
  XOR2_X1 U11438 ( .A(n11430), .B(n11431), .Z(n11429) );
  INV_X1 U11439 ( .A(n11432), .ZN(n11425) );
  NOR2_X1 U11440 ( .A1(n11167), .A2(n11168), .ZN(n11432) );
  NOR2_X1 U11441 ( .A1(n10931), .A2(n8830), .ZN(n11168) );
  NAND2_X1 U11442 ( .A1(n11433), .A2(n11434), .ZN(n11167) );
  NAND2_X1 U11443 ( .A1(n11175), .A2(n11435), .ZN(n11434) );
  NAND2_X1 U11444 ( .A1(n11174), .A2(n11172), .ZN(n11435) );
  NOR2_X1 U11445 ( .A1(n10931), .A2(n8839), .ZN(n11175) );
  INV_X1 U11446 ( .A(n11436), .ZN(n11433) );
  NOR2_X1 U11447 ( .A1(n11172), .A2(n11174), .ZN(n11436) );
  NOR2_X1 U11448 ( .A1(n11437), .A2(n11438), .ZN(n11174) );
  INV_X1 U11449 ( .A(n11439), .ZN(n11438) );
  NAND2_X1 U11450 ( .A1(n11204), .A2(n11440), .ZN(n11439) );
  NAND2_X1 U11451 ( .A1(n11205), .A2(n11203), .ZN(n11440) );
  NOR2_X1 U11452 ( .A1(n10931), .A2(n8844), .ZN(n11204) );
  NOR2_X1 U11453 ( .A1(n11203), .A2(n11205), .ZN(n11437) );
  NOR2_X1 U11454 ( .A1(n11441), .A2(n11442), .ZN(n11205) );
  INV_X1 U11455 ( .A(n11443), .ZN(n11442) );
  NAND2_X1 U11456 ( .A1(n11198), .A2(n11444), .ZN(n11443) );
  NAND2_X1 U11457 ( .A1(n11445), .A2(n11200), .ZN(n11444) );
  NOR2_X1 U11458 ( .A1(n10931), .A2(n9161), .ZN(n11198) );
  NOR2_X1 U11459 ( .A1(n11200), .A2(n11445), .ZN(n11441) );
  INV_X1 U11460 ( .A(n11201), .ZN(n11445) );
  NAND2_X1 U11461 ( .A1(n11446), .A2(n11447), .ZN(n11201) );
  NAND2_X1 U11462 ( .A1(b_19_), .A2(n11448), .ZN(n11447) );
  NAND2_X1 U11463 ( .A1(n8358), .A2(n11449), .ZN(n11448) );
  NAND2_X1 U11464 ( .A1(a_31_), .A2(n11196), .ZN(n11449) );
  NAND2_X1 U11465 ( .A1(b_20_), .A2(n11450), .ZN(n11446) );
  NAND2_X1 U11466 ( .A1(n8362), .A2(n11451), .ZN(n11450) );
  NAND2_X1 U11467 ( .A1(a_30_), .A2(n11452), .ZN(n11451) );
  NAND2_X1 U11468 ( .A1(n11453), .A2(b_21_), .ZN(n11200) );
  NOR2_X1 U11469 ( .A1(n9170), .A2(n11196), .ZN(n11453) );
  XOR2_X1 U11470 ( .A(n11454), .B(n11455), .Z(n11203) );
  XOR2_X1 U11471 ( .A(n11456), .B(n11457), .Z(n11455) );
  XOR2_X1 U11472 ( .A(n11458), .B(n11459), .Z(n11172) );
  XNOR2_X1 U11473 ( .A(n11460), .B(n11461), .ZN(n11458) );
  XNOR2_X1 U11474 ( .A(n11462), .B(n11463), .ZN(n11211) );
  XNOR2_X1 U11475 ( .A(n11464), .B(n11465), .ZN(n11463) );
  XOR2_X1 U11476 ( .A(n11466), .B(n11467), .Z(n11150) );
  XOR2_X1 U11477 ( .A(n11468), .B(n11469), .Z(n11466) );
  XNOR2_X1 U11478 ( .A(n11470), .B(n11471), .ZN(n11219) );
  NAND2_X1 U11479 ( .A1(n11472), .A2(n11473), .ZN(n11470) );
  XNOR2_X1 U11480 ( .A(n11474), .B(n11475), .ZN(n11222) );
  NAND2_X1 U11481 ( .A1(n11476), .A2(n11477), .ZN(n11474) );
  XNOR2_X1 U11482 ( .A(n11478), .B(n11479), .ZN(n11089) );
  NAND2_X1 U11483 ( .A1(n11480), .A2(n11481), .ZN(n11478) );
  XOR2_X1 U11484 ( .A(n11482), .B(n11483), .Z(n11070) );
  XOR2_X1 U11485 ( .A(n11484), .B(n11485), .Z(n11482) );
  NOR2_X1 U11486 ( .A1(n8750), .A2(n11196), .ZN(n11485) );
  XNOR2_X1 U11487 ( .A(n11486), .B(n11487), .ZN(n11062) );
  XOR2_X1 U11488 ( .A(n11488), .B(n11489), .Z(n11487) );
  NAND2_X1 U11489 ( .A1(b_20_), .A2(a_11_), .ZN(n11489) );
  NAND2_X1 U11490 ( .A1(n11490), .A2(n8648), .ZN(n11243) );
  XNOR2_X1 U11491 ( .A(n11491), .B(n11492), .ZN(n8648) );
  NAND2_X1 U11492 ( .A1(n11493), .A2(n11494), .ZN(n11491) );
  INV_X1 U11493 ( .A(n11495), .ZN(n11490) );
  NOR2_X1 U11494 ( .A1(n8651), .A2(n8650), .ZN(n11495) );
  INV_X1 U11495 ( .A(n11496), .ZN(n8565) );
  NOR2_X1 U11496 ( .A1(n8644), .A2(n8643), .ZN(n11496) );
  NAND2_X1 U11497 ( .A1(n11497), .A2(n11498), .ZN(n8643) );
  NAND2_X1 U11498 ( .A1(n11499), .A2(n11500), .ZN(n11498) );
  INV_X1 U11499 ( .A(n8638), .ZN(n11497) );
  NOR2_X1 U11500 ( .A1(n11500), .A2(n11499), .ZN(n8638) );
  INV_X1 U11501 ( .A(n11501), .ZN(n11499) );
  NAND2_X1 U11502 ( .A1(n11502), .A2(n11503), .ZN(n11501) );
  NAND2_X1 U11503 ( .A1(n11504), .A2(b_19_), .ZN(n11503) );
  NOR2_X1 U11504 ( .A1(n11505), .A2(n8690), .ZN(n11504) );
  NOR2_X1 U11505 ( .A1(n11506), .A2(n11507), .ZN(n11505) );
  NAND2_X1 U11506 ( .A1(n11506), .A2(n11507), .ZN(n11502) );
  XNOR2_X1 U11507 ( .A(n11508), .B(n11509), .ZN(n11500) );
  XNOR2_X1 U11508 ( .A(n11510), .B(n11511), .ZN(n11509) );
  NAND2_X1 U11509 ( .A1(n8651), .A2(n8650), .ZN(n8644) );
  NAND2_X1 U11510 ( .A1(n11493), .A2(n11512), .ZN(n8650) );
  NAND2_X1 U11511 ( .A1(n11492), .A2(n11494), .ZN(n11512) );
  NAND2_X1 U11512 ( .A1(n11513), .A2(n11514), .ZN(n11494) );
  INV_X1 U11513 ( .A(n11515), .ZN(n11514) );
  NAND2_X1 U11514 ( .A1(b_20_), .A2(a_0_), .ZN(n11513) );
  XNOR2_X1 U11515 ( .A(n11516), .B(n11517), .ZN(n11492) );
  NAND2_X1 U11516 ( .A1(n11518), .A2(n11519), .ZN(n11516) );
  NAND2_X1 U11517 ( .A1(n11515), .A2(a_0_), .ZN(n11493) );
  NOR2_X1 U11518 ( .A1(n11520), .A2(n11521), .ZN(n11515) );
  INV_X1 U11519 ( .A(n11522), .ZN(n11521) );
  NAND2_X1 U11520 ( .A1(n11250), .A2(n11523), .ZN(n11522) );
  NAND2_X1 U11521 ( .A1(n11252), .A2(n11251), .ZN(n11523) );
  XNOR2_X1 U11522 ( .A(n11524), .B(n11525), .ZN(n11250) );
  XNOR2_X1 U11523 ( .A(n11526), .B(n11527), .ZN(n11525) );
  NOR2_X1 U11524 ( .A1(n11251), .A2(n11252), .ZN(n11520) );
  NOR2_X1 U11525 ( .A1(n11196), .A2(n8502), .ZN(n11252) );
  NAND2_X1 U11526 ( .A1(n11259), .A2(n11528), .ZN(n11251) );
  NAND2_X1 U11527 ( .A1(n11258), .A2(n11260), .ZN(n11528) );
  NAND2_X1 U11528 ( .A1(n11529), .A2(n11530), .ZN(n11260) );
  INV_X1 U11529 ( .A(n11531), .ZN(n11530) );
  NAND2_X1 U11530 ( .A1(b_20_), .A2(a_2_), .ZN(n11529) );
  XNOR2_X1 U11531 ( .A(n11532), .B(n11533), .ZN(n11258) );
  XNOR2_X1 U11532 ( .A(n11534), .B(n11535), .ZN(n11532) );
  NOR2_X1 U11533 ( .A1(n8707), .A2(n11452), .ZN(n11535) );
  NAND2_X1 U11534 ( .A1(n11531), .A2(a_2_), .ZN(n11259) );
  NOR2_X1 U11535 ( .A1(n11536), .A2(n11537), .ZN(n11531) );
  INV_X1 U11536 ( .A(n11538), .ZN(n11537) );
  NAND2_X1 U11537 ( .A1(n11265), .A2(n11539), .ZN(n11538) );
  NAND2_X1 U11538 ( .A1(n11268), .A2(n11267), .ZN(n11539) );
  XNOR2_X1 U11539 ( .A(n11540), .B(n11541), .ZN(n11265) );
  XNOR2_X1 U11540 ( .A(n11542), .B(n11543), .ZN(n11541) );
  NOR2_X1 U11541 ( .A1(n11267), .A2(n11268), .ZN(n11536) );
  NOR2_X1 U11542 ( .A1(n11196), .A2(n8707), .ZN(n11268) );
  NAND2_X1 U11543 ( .A1(n11275), .A2(n11544), .ZN(n11267) );
  NAND2_X1 U11544 ( .A1(n11274), .A2(n11276), .ZN(n11544) );
  NAND2_X1 U11545 ( .A1(n11545), .A2(n11546), .ZN(n11276) );
  INV_X1 U11546 ( .A(n11547), .ZN(n11546) );
  NAND2_X1 U11547 ( .A1(b_20_), .A2(a_4_), .ZN(n11545) );
  XNOR2_X1 U11548 ( .A(n11548), .B(n11549), .ZN(n11274) );
  NAND2_X1 U11549 ( .A1(n11550), .A2(n11551), .ZN(n11548) );
  NAND2_X1 U11550 ( .A1(n11547), .A2(a_4_), .ZN(n11275) );
  NOR2_X1 U11551 ( .A1(n11552), .A2(n11553), .ZN(n11547) );
  INV_X1 U11552 ( .A(n11554), .ZN(n11553) );
  NAND2_X1 U11553 ( .A1(n11281), .A2(n11555), .ZN(n11554) );
  NAND2_X1 U11554 ( .A1(n11284), .A2(n11283), .ZN(n11555) );
  XNOR2_X1 U11555 ( .A(n11556), .B(n11557), .ZN(n11281) );
  XNOR2_X1 U11556 ( .A(n11558), .B(n11559), .ZN(n11557) );
  NOR2_X1 U11557 ( .A1(n11283), .A2(n11284), .ZN(n11552) );
  NOR2_X1 U11558 ( .A1(n11196), .A2(n8717), .ZN(n11284) );
  NAND2_X1 U11559 ( .A1(n11291), .A2(n11560), .ZN(n11283) );
  NAND2_X1 U11560 ( .A1(n11290), .A2(n11292), .ZN(n11560) );
  NAND2_X1 U11561 ( .A1(n11561), .A2(n11562), .ZN(n11292) );
  INV_X1 U11562 ( .A(n11563), .ZN(n11562) );
  NAND2_X1 U11563 ( .A1(b_20_), .A2(a_6_), .ZN(n11561) );
  XNOR2_X1 U11564 ( .A(n11564), .B(n11565), .ZN(n11290) );
  NAND2_X1 U11565 ( .A1(n11566), .A2(n11567), .ZN(n11564) );
  NAND2_X1 U11566 ( .A1(n11563), .A2(a_6_), .ZN(n11291) );
  NOR2_X1 U11567 ( .A1(n11568), .A2(n11569), .ZN(n11563) );
  INV_X1 U11568 ( .A(n11570), .ZN(n11569) );
  NAND2_X1 U11569 ( .A1(n11298), .A2(n11571), .ZN(n11570) );
  NAND2_X1 U11570 ( .A1(n11300), .A2(n11299), .ZN(n11571) );
  XNOR2_X1 U11571 ( .A(n11572), .B(n11573), .ZN(n11298) );
  XNOR2_X1 U11572 ( .A(n11574), .B(n11575), .ZN(n11573) );
  NOR2_X1 U11573 ( .A1(n11299), .A2(n11300), .ZN(n11568) );
  NOR2_X1 U11574 ( .A1(n11196), .A2(n8726), .ZN(n11300) );
  NAND2_X1 U11575 ( .A1(n11307), .A2(n11576), .ZN(n11299) );
  NAND2_X1 U11576 ( .A1(n11306), .A2(n11308), .ZN(n11576) );
  NAND2_X1 U11577 ( .A1(n11577), .A2(n11578), .ZN(n11308) );
  NAND2_X1 U11578 ( .A1(b_20_), .A2(a_8_), .ZN(n11578) );
  INV_X1 U11579 ( .A(n11579), .ZN(n11577) );
  XNOR2_X1 U11580 ( .A(n11580), .B(n11581), .ZN(n11306) );
  XOR2_X1 U11581 ( .A(n11582), .B(n11583), .Z(n11581) );
  NAND2_X1 U11582 ( .A1(b_19_), .A2(a_9_), .ZN(n11583) );
  NAND2_X1 U11583 ( .A1(a_8_), .A2(n11579), .ZN(n11307) );
  NAND2_X1 U11584 ( .A1(n11584), .A2(n11585), .ZN(n11579) );
  NAND2_X1 U11585 ( .A1(n11586), .A2(b_20_), .ZN(n11585) );
  NOR2_X1 U11586 ( .A1(n11587), .A2(n8736), .ZN(n11586) );
  NOR2_X1 U11587 ( .A1(n11313), .A2(n11315), .ZN(n11587) );
  NAND2_X1 U11588 ( .A1(n11313), .A2(n11315), .ZN(n11584) );
  NAND2_X1 U11589 ( .A1(n11588), .A2(n11589), .ZN(n11315) );
  NAND2_X1 U11590 ( .A1(n11590), .A2(b_20_), .ZN(n11589) );
  NOR2_X1 U11591 ( .A1(n11591), .A2(n8741), .ZN(n11590) );
  NOR2_X1 U11592 ( .A1(n11321), .A2(n11323), .ZN(n11591) );
  NAND2_X1 U11593 ( .A1(n11321), .A2(n11323), .ZN(n11588) );
  NAND2_X1 U11594 ( .A1(n11592), .A2(n11593), .ZN(n11323) );
  NAND2_X1 U11595 ( .A1(n11594), .A2(b_20_), .ZN(n11593) );
  NOR2_X1 U11596 ( .A1(n11595), .A2(n8452), .ZN(n11594) );
  NOR2_X1 U11597 ( .A1(n11486), .A2(n11488), .ZN(n11595) );
  NAND2_X1 U11598 ( .A1(n11486), .A2(n11488), .ZN(n11592) );
  NAND2_X1 U11599 ( .A1(n11596), .A2(n11597), .ZN(n11488) );
  NAND2_X1 U11600 ( .A1(n11598), .A2(b_20_), .ZN(n11597) );
  NOR2_X1 U11601 ( .A1(n11599), .A2(n8750), .ZN(n11598) );
  NOR2_X1 U11602 ( .A1(n11483), .A2(n11484), .ZN(n11599) );
  NAND2_X1 U11603 ( .A1(n11483), .A2(n11484), .ZN(n11596) );
  NAND2_X1 U11604 ( .A1(n11339), .A2(n11600), .ZN(n11484) );
  NAND2_X1 U11605 ( .A1(n11338), .A2(n11340), .ZN(n11600) );
  NAND2_X1 U11606 ( .A1(n11601), .A2(n11602), .ZN(n11340) );
  NAND2_X1 U11607 ( .A1(b_20_), .A2(a_13_), .ZN(n11602) );
  INV_X1 U11608 ( .A(n11603), .ZN(n11601) );
  XNOR2_X1 U11609 ( .A(n11604), .B(n11605), .ZN(n11338) );
  XOR2_X1 U11610 ( .A(n11606), .B(n11607), .Z(n11605) );
  NAND2_X1 U11611 ( .A1(b_19_), .A2(a_14_), .ZN(n11607) );
  NAND2_X1 U11612 ( .A1(a_13_), .A2(n11603), .ZN(n11339) );
  NAND2_X1 U11613 ( .A1(n11347), .A2(n11608), .ZN(n11603) );
  NAND2_X1 U11614 ( .A1(n11346), .A2(n11348), .ZN(n11608) );
  NAND2_X1 U11615 ( .A1(n11609), .A2(n11610), .ZN(n11348) );
  NAND2_X1 U11616 ( .A1(b_20_), .A2(a_14_), .ZN(n11610) );
  INV_X1 U11617 ( .A(n11611), .ZN(n11609) );
  XOR2_X1 U11618 ( .A(n11612), .B(n11613), .Z(n11346) );
  XOR2_X1 U11619 ( .A(n11614), .B(n11615), .Z(n11612) );
  NOR2_X1 U11620 ( .A1(n8763), .A2(n11452), .ZN(n11615) );
  NAND2_X1 U11621 ( .A1(a_14_), .A2(n11611), .ZN(n11347) );
  NAND2_X1 U11622 ( .A1(n11480), .A2(n11616), .ZN(n11611) );
  NAND2_X1 U11623 ( .A1(n11479), .A2(n11481), .ZN(n11616) );
  NAND2_X1 U11624 ( .A1(n11617), .A2(n11618), .ZN(n11481) );
  NAND2_X1 U11625 ( .A1(b_20_), .A2(a_15_), .ZN(n11618) );
  INV_X1 U11626 ( .A(n11619), .ZN(n11617) );
  XNOR2_X1 U11627 ( .A(n11620), .B(n11621), .ZN(n11479) );
  NAND2_X1 U11628 ( .A1(n11622), .A2(n11623), .ZN(n11620) );
  NAND2_X1 U11629 ( .A1(a_15_), .A2(n11619), .ZN(n11480) );
  NAND2_X1 U11630 ( .A1(n11476), .A2(n11624), .ZN(n11619) );
  NAND2_X1 U11631 ( .A1(n11475), .A2(n11477), .ZN(n11624) );
  NAND2_X1 U11632 ( .A1(n11625), .A2(n11626), .ZN(n11477) );
  NAND2_X1 U11633 ( .A1(b_20_), .A2(a_16_), .ZN(n11626) );
  INV_X1 U11634 ( .A(n11627), .ZN(n11625) );
  XNOR2_X1 U11635 ( .A(n11628), .B(n11629), .ZN(n11475) );
  NAND2_X1 U11636 ( .A1(n11630), .A2(n11631), .ZN(n11628) );
  NAND2_X1 U11637 ( .A1(a_16_), .A2(n11627), .ZN(n11476) );
  NAND2_X1 U11638 ( .A1(n11472), .A2(n11632), .ZN(n11627) );
  NAND2_X1 U11639 ( .A1(n11471), .A2(n11473), .ZN(n11632) );
  NAND2_X1 U11640 ( .A1(n11633), .A2(n11634), .ZN(n11473) );
  NAND2_X1 U11641 ( .A1(b_20_), .A2(a_17_), .ZN(n11634) );
  INV_X1 U11642 ( .A(n11635), .ZN(n11633) );
  XOR2_X1 U11643 ( .A(n11636), .B(n11637), .Z(n11471) );
  XOR2_X1 U11644 ( .A(n11638), .B(n11639), .Z(n11636) );
  NAND2_X1 U11645 ( .A1(a_17_), .A2(n11635), .ZN(n11472) );
  NAND2_X1 U11646 ( .A1(n11640), .A2(n11641), .ZN(n11635) );
  NAND2_X1 U11647 ( .A1(n11642), .A2(b_20_), .ZN(n11641) );
  NOR2_X1 U11648 ( .A1(n11643), .A2(n10616), .ZN(n11642) );
  NOR2_X1 U11649 ( .A1(n11365), .A2(n11367), .ZN(n11643) );
  NAND2_X1 U11650 ( .A1(n11365), .A2(n11367), .ZN(n11640) );
  NAND2_X1 U11651 ( .A1(n11644), .A2(n11645), .ZN(n11367) );
  NAND2_X1 U11652 ( .A1(n11646), .A2(b_20_), .ZN(n11645) );
  NOR2_X1 U11653 ( .A1(n11647), .A2(n8881), .ZN(n11646) );
  NOR2_X1 U11654 ( .A1(n11374), .A2(n11376), .ZN(n11647) );
  NAND2_X1 U11655 ( .A1(n11374), .A2(n11376), .ZN(n11644) );
  NAND2_X1 U11656 ( .A1(n11648), .A2(n11649), .ZN(n11376) );
  INV_X1 U11657 ( .A(n11650), .ZN(n11649) );
  NOR2_X1 U11658 ( .A1(n11383), .A2(n11651), .ZN(n11650) );
  NOR2_X1 U11659 ( .A1(n11384), .A2(n11381), .ZN(n11651) );
  NAND2_X1 U11660 ( .A1(n11381), .A2(n11384), .ZN(n11648) );
  NAND2_X1 U11661 ( .A1(n11391), .A2(n11652), .ZN(n11384) );
  NAND2_X1 U11662 ( .A1(n11390), .A2(n11392), .ZN(n11652) );
  NAND2_X1 U11663 ( .A1(n11653), .A2(n11654), .ZN(n11392) );
  NAND2_X1 U11664 ( .A1(b_20_), .A2(a_21_), .ZN(n11654) );
  INV_X1 U11665 ( .A(n11655), .ZN(n11653) );
  XNOR2_X1 U11666 ( .A(n11656), .B(n11657), .ZN(n11390) );
  NAND2_X1 U11667 ( .A1(n11658), .A2(n11659), .ZN(n11656) );
  NAND2_X1 U11668 ( .A1(a_21_), .A2(n11655), .ZN(n11391) );
  NAND2_X1 U11669 ( .A1(n11399), .A2(n11660), .ZN(n11655) );
  NAND2_X1 U11670 ( .A1(n11398), .A2(n11400), .ZN(n11660) );
  NAND2_X1 U11671 ( .A1(n11661), .A2(n11662), .ZN(n11400) );
  NAND2_X1 U11672 ( .A1(b_20_), .A2(a_22_), .ZN(n11662) );
  INV_X1 U11673 ( .A(n11663), .ZN(n11661) );
  XOR2_X1 U11674 ( .A(n11664), .B(n11665), .Z(n11398) );
  XOR2_X1 U11675 ( .A(n11666), .B(n11667), .Z(n11664) );
  NOR2_X1 U11676 ( .A1(n8812), .A2(n11452), .ZN(n11667) );
  NAND2_X1 U11677 ( .A1(a_22_), .A2(n11663), .ZN(n11399) );
  NAND2_X1 U11678 ( .A1(n11668), .A2(n11669), .ZN(n11663) );
  NAND2_X1 U11679 ( .A1(n11670), .A2(b_20_), .ZN(n11669) );
  NOR2_X1 U11680 ( .A1(n11671), .A2(n8812), .ZN(n11670) );
  NOR2_X1 U11681 ( .A1(n11406), .A2(n11407), .ZN(n11671) );
  NAND2_X1 U11682 ( .A1(n11406), .A2(n11407), .ZN(n11668) );
  NAND2_X1 U11683 ( .A1(n11672), .A2(n11673), .ZN(n11407) );
  NAND2_X1 U11684 ( .A1(n11469), .A2(n11674), .ZN(n11673) );
  INV_X1 U11685 ( .A(n11675), .ZN(n11674) );
  NOR2_X1 U11686 ( .A1(n11468), .A2(n11467), .ZN(n11675) );
  NOR2_X1 U11687 ( .A1(n11196), .A2(n9131), .ZN(n11469) );
  NAND2_X1 U11688 ( .A1(n11467), .A2(n11468), .ZN(n11672) );
  NAND2_X1 U11689 ( .A1(n11676), .A2(n11677), .ZN(n11468) );
  NAND2_X1 U11690 ( .A1(n11465), .A2(n11678), .ZN(n11677) );
  NAND2_X1 U11691 ( .A1(n11462), .A2(n11464), .ZN(n11678) );
  NOR2_X1 U11692 ( .A1(n11196), .A2(n8825), .ZN(n11465) );
  INV_X1 U11693 ( .A(n11679), .ZN(n11676) );
  NOR2_X1 U11694 ( .A1(n11464), .A2(n11462), .ZN(n11679) );
  XNOR2_X1 U11695 ( .A(n11680), .B(n11681), .ZN(n11462) );
  XNOR2_X1 U11696 ( .A(n11682), .B(n11683), .ZN(n11681) );
  NAND2_X1 U11697 ( .A1(n11684), .A2(n11685), .ZN(n11464) );
  NAND2_X1 U11698 ( .A1(n11421), .A2(n11686), .ZN(n11685) );
  NAND2_X1 U11699 ( .A1(n11424), .A2(n11423), .ZN(n11686) );
  XNOR2_X1 U11700 ( .A(n11687), .B(n11688), .ZN(n11421) );
  XOR2_X1 U11701 ( .A(n11689), .B(n11690), .Z(n11688) );
  INV_X1 U11702 ( .A(n11691), .ZN(n11684) );
  NOR2_X1 U11703 ( .A1(n11423), .A2(n11424), .ZN(n11691) );
  NOR2_X1 U11704 ( .A1(n11196), .A2(n8830), .ZN(n11424) );
  NAND2_X1 U11705 ( .A1(n11692), .A2(n11693), .ZN(n11423) );
  NAND2_X1 U11706 ( .A1(n11431), .A2(n11694), .ZN(n11693) );
  NAND2_X1 U11707 ( .A1(n11430), .A2(n11428), .ZN(n11694) );
  NOR2_X1 U11708 ( .A1(n11196), .A2(n8839), .ZN(n11431) );
  INV_X1 U11709 ( .A(n11695), .ZN(n11692) );
  NOR2_X1 U11710 ( .A1(n11428), .A2(n11430), .ZN(n11695) );
  NOR2_X1 U11711 ( .A1(n11696), .A2(n11697), .ZN(n11430) );
  INV_X1 U11712 ( .A(n11698), .ZN(n11697) );
  NAND2_X1 U11713 ( .A1(n11460), .A2(n11699), .ZN(n11698) );
  NAND2_X1 U11714 ( .A1(n11461), .A2(n11459), .ZN(n11699) );
  NOR2_X1 U11715 ( .A1(n11196), .A2(n8844), .ZN(n11460) );
  NOR2_X1 U11716 ( .A1(n11459), .A2(n11461), .ZN(n11696) );
  NOR2_X1 U11717 ( .A1(n11700), .A2(n11701), .ZN(n11461) );
  INV_X1 U11718 ( .A(n11702), .ZN(n11701) );
  NAND2_X1 U11719 ( .A1(n11454), .A2(n11703), .ZN(n11702) );
  NAND2_X1 U11720 ( .A1(n11704), .A2(n11456), .ZN(n11703) );
  NOR2_X1 U11721 ( .A1(n11196), .A2(n9161), .ZN(n11454) );
  NOR2_X1 U11722 ( .A1(n11456), .A2(n11704), .ZN(n11700) );
  INV_X1 U11723 ( .A(n11457), .ZN(n11704) );
  NAND2_X1 U11724 ( .A1(n11705), .A2(n11706), .ZN(n11457) );
  NAND2_X1 U11725 ( .A1(b_18_), .A2(n11707), .ZN(n11706) );
  NAND2_X1 U11726 ( .A1(n8358), .A2(n11708), .ZN(n11707) );
  NAND2_X1 U11727 ( .A1(a_31_), .A2(n11452), .ZN(n11708) );
  NAND2_X1 U11728 ( .A1(b_19_), .A2(n11709), .ZN(n11705) );
  NAND2_X1 U11729 ( .A1(n8362), .A2(n11710), .ZN(n11709) );
  NAND2_X1 U11730 ( .A1(a_30_), .A2(n11711), .ZN(n11710) );
  NAND2_X1 U11731 ( .A1(n11712), .A2(b_20_), .ZN(n11456) );
  XOR2_X1 U11732 ( .A(n11713), .B(n11714), .Z(n11459) );
  XOR2_X1 U11733 ( .A(n11715), .B(n11716), .Z(n11714) );
  XOR2_X1 U11734 ( .A(n11717), .B(n11718), .Z(n11428) );
  XNOR2_X1 U11735 ( .A(n11719), .B(n11720), .ZN(n11717) );
  XNOR2_X1 U11736 ( .A(n11721), .B(n11722), .ZN(n11467) );
  XNOR2_X1 U11737 ( .A(n11723), .B(n11724), .ZN(n11722) );
  XOR2_X1 U11738 ( .A(n11725), .B(n11726), .Z(n11406) );
  XOR2_X1 U11739 ( .A(n11727), .B(n11728), .Z(n11725) );
  XNOR2_X1 U11740 ( .A(n11729), .B(n11730), .ZN(n11381) );
  NAND2_X1 U11741 ( .A1(n11731), .A2(n11732), .ZN(n11729) );
  XOR2_X1 U11742 ( .A(n11733), .B(n11734), .Z(n11374) );
  XNOR2_X1 U11743 ( .A(n11735), .B(n11736), .ZN(n11734) );
  XOR2_X1 U11744 ( .A(n11737), .B(n11738), .Z(n11365) );
  XOR2_X1 U11745 ( .A(n11739), .B(n11740), .Z(n11738) );
  XNOR2_X1 U11746 ( .A(n11741), .B(n11742), .ZN(n11483) );
  NAND2_X1 U11747 ( .A1(n11743), .A2(n11744), .ZN(n11741) );
  XNOR2_X1 U11748 ( .A(n11745), .B(n11746), .ZN(n11486) );
  XOR2_X1 U11749 ( .A(n11747), .B(n11748), .Z(n11745) );
  XNOR2_X1 U11750 ( .A(n11749), .B(n11750), .ZN(n11321) );
  XNOR2_X1 U11751 ( .A(n11751), .B(n11752), .ZN(n11749) );
  XNOR2_X1 U11752 ( .A(n11753), .B(n11754), .ZN(n11313) );
  XOR2_X1 U11753 ( .A(n11755), .B(n11756), .Z(n11754) );
  NAND2_X1 U11754 ( .A1(b_19_), .A2(a_10_), .ZN(n11756) );
  XNOR2_X1 U11755 ( .A(n11506), .B(n11757), .ZN(n8651) );
  XOR2_X1 U11756 ( .A(n11507), .B(n11758), .Z(n11757) );
  NAND2_X1 U11757 ( .A1(b_19_), .A2(a_0_), .ZN(n11758) );
  NAND2_X1 U11758 ( .A1(n11518), .A2(n11759), .ZN(n11507) );
  NAND2_X1 U11759 ( .A1(n11517), .A2(n11519), .ZN(n11759) );
  NAND2_X1 U11760 ( .A1(n11760), .A2(n11761), .ZN(n11519) );
  INV_X1 U11761 ( .A(n11762), .ZN(n11761) );
  NAND2_X1 U11762 ( .A1(b_19_), .A2(a_1_), .ZN(n11760) );
  XOR2_X1 U11763 ( .A(n11763), .B(n11764), .Z(n11517) );
  XOR2_X1 U11764 ( .A(n11765), .B(n11766), .Z(n11763) );
  NAND2_X1 U11765 ( .A1(n11762), .A2(a_1_), .ZN(n11518) );
  NOR2_X1 U11766 ( .A1(n11767), .A2(n11768), .ZN(n11762) );
  INV_X1 U11767 ( .A(n11769), .ZN(n11768) );
  NAND2_X1 U11768 ( .A1(n11524), .A2(n11770), .ZN(n11769) );
  NAND2_X1 U11769 ( .A1(n11527), .A2(n11526), .ZN(n11770) );
  XNOR2_X1 U11770 ( .A(n11771), .B(n11772), .ZN(n11524) );
  XNOR2_X1 U11771 ( .A(n11773), .B(n11774), .ZN(n11772) );
  NOR2_X1 U11772 ( .A1(n11526), .A2(n11527), .ZN(n11767) );
  NOR2_X1 U11773 ( .A1(n11452), .A2(n8497), .ZN(n11527) );
  NAND2_X1 U11774 ( .A1(n11775), .A2(n11776), .ZN(n11526) );
  NAND2_X1 U11775 ( .A1(n11777), .A2(b_19_), .ZN(n11776) );
  NOR2_X1 U11776 ( .A1(n11778), .A2(n8707), .ZN(n11777) );
  NOR2_X1 U11777 ( .A1(n11534), .A2(n11533), .ZN(n11778) );
  NAND2_X1 U11778 ( .A1(n11534), .A2(n11533), .ZN(n11775) );
  XNOR2_X1 U11779 ( .A(n11779), .B(n11780), .ZN(n11533) );
  NAND2_X1 U11780 ( .A1(n11781), .A2(n11782), .ZN(n11779) );
  NOR2_X1 U11781 ( .A1(n11783), .A2(n11784), .ZN(n11534) );
  INV_X1 U11782 ( .A(n11785), .ZN(n11784) );
  NAND2_X1 U11783 ( .A1(n11540), .A2(n11786), .ZN(n11785) );
  NAND2_X1 U11784 ( .A1(n11543), .A2(n11542), .ZN(n11786) );
  XNOR2_X1 U11785 ( .A(n11787), .B(n11788), .ZN(n11540) );
  XOR2_X1 U11786 ( .A(n11789), .B(n11790), .Z(n11787) );
  NOR2_X1 U11787 ( .A1(n8717), .A2(n11711), .ZN(n11790) );
  NOR2_X1 U11788 ( .A1(n11542), .A2(n11543), .ZN(n11783) );
  NOR2_X1 U11789 ( .A1(n11452), .A2(n8712), .ZN(n11543) );
  NAND2_X1 U11790 ( .A1(n11550), .A2(n11791), .ZN(n11542) );
  NAND2_X1 U11791 ( .A1(n11549), .A2(n11551), .ZN(n11791) );
  NAND2_X1 U11792 ( .A1(n11792), .A2(n11793), .ZN(n11551) );
  INV_X1 U11793 ( .A(n11794), .ZN(n11793) );
  NAND2_X1 U11794 ( .A1(b_19_), .A2(a_5_), .ZN(n11792) );
  XNOR2_X1 U11795 ( .A(n11795), .B(n11796), .ZN(n11549) );
  NAND2_X1 U11796 ( .A1(n11797), .A2(n11798), .ZN(n11795) );
  NAND2_X1 U11797 ( .A1(n11794), .A2(a_5_), .ZN(n11550) );
  NOR2_X1 U11798 ( .A1(n11799), .A2(n11800), .ZN(n11794) );
  INV_X1 U11799 ( .A(n11801), .ZN(n11800) );
  NAND2_X1 U11800 ( .A1(n11556), .A2(n11802), .ZN(n11801) );
  NAND2_X1 U11801 ( .A1(n11559), .A2(n11558), .ZN(n11802) );
  XNOR2_X1 U11802 ( .A(n11803), .B(n11804), .ZN(n11556) );
  XNOR2_X1 U11803 ( .A(n11805), .B(n11806), .ZN(n11804) );
  NOR2_X1 U11804 ( .A1(n11558), .A2(n11559), .ZN(n11799) );
  NOR2_X1 U11805 ( .A1(n11452), .A2(n8480), .ZN(n11559) );
  NAND2_X1 U11806 ( .A1(n11566), .A2(n11807), .ZN(n11558) );
  NAND2_X1 U11807 ( .A1(n11565), .A2(n11567), .ZN(n11807) );
  NAND2_X1 U11808 ( .A1(n11808), .A2(n11809), .ZN(n11567) );
  INV_X1 U11809 ( .A(n11810), .ZN(n11809) );
  NAND2_X1 U11810 ( .A1(b_19_), .A2(a_7_), .ZN(n11808) );
  XNOR2_X1 U11811 ( .A(n11811), .B(n11812), .ZN(n11565) );
  NAND2_X1 U11812 ( .A1(n11813), .A2(n11814), .ZN(n11811) );
  NAND2_X1 U11813 ( .A1(n11810), .A2(a_7_), .ZN(n11566) );
  NOR2_X1 U11814 ( .A1(n11815), .A2(n11816), .ZN(n11810) );
  INV_X1 U11815 ( .A(n11817), .ZN(n11816) );
  NAND2_X1 U11816 ( .A1(n11572), .A2(n11818), .ZN(n11817) );
  NAND2_X1 U11817 ( .A1(n11575), .A2(n11574), .ZN(n11818) );
  XOR2_X1 U11818 ( .A(n11819), .B(n11820), .Z(n11572) );
  XOR2_X1 U11819 ( .A(n11821), .B(n11822), .Z(n11819) );
  NOR2_X1 U11820 ( .A1(n11574), .A2(n11575), .ZN(n11815) );
  NOR2_X1 U11821 ( .A1(n11452), .A2(n8731), .ZN(n11575) );
  NAND2_X1 U11822 ( .A1(n11823), .A2(n11824), .ZN(n11574) );
  NAND2_X1 U11823 ( .A1(n11825), .A2(b_19_), .ZN(n11824) );
  NOR2_X1 U11824 ( .A1(n11826), .A2(n8736), .ZN(n11825) );
  NOR2_X1 U11825 ( .A1(n11580), .A2(n11582), .ZN(n11826) );
  NAND2_X1 U11826 ( .A1(n11580), .A2(n11582), .ZN(n11823) );
  NAND2_X1 U11827 ( .A1(n11827), .A2(n11828), .ZN(n11582) );
  NAND2_X1 U11828 ( .A1(n11829), .A2(b_19_), .ZN(n11828) );
  NOR2_X1 U11829 ( .A1(n11830), .A2(n8741), .ZN(n11829) );
  NOR2_X1 U11830 ( .A1(n11753), .A2(n11755), .ZN(n11830) );
  NAND2_X1 U11831 ( .A1(n11753), .A2(n11755), .ZN(n11827) );
  NAND2_X1 U11832 ( .A1(n11831), .A2(n11832), .ZN(n11755) );
  NAND2_X1 U11833 ( .A1(n11752), .A2(n11833), .ZN(n11832) );
  NAND2_X1 U11834 ( .A1(n11751), .A2(n11750), .ZN(n11833) );
  NOR2_X1 U11835 ( .A1(n11452), .A2(n8452), .ZN(n11752) );
  INV_X1 U11836 ( .A(n11834), .ZN(n11831) );
  NOR2_X1 U11837 ( .A1(n11750), .A2(n11751), .ZN(n11834) );
  NOR2_X1 U11838 ( .A1(n11835), .A2(n11836), .ZN(n11751) );
  INV_X1 U11839 ( .A(n11837), .ZN(n11836) );
  NAND2_X1 U11840 ( .A1(n11748), .A2(n11838), .ZN(n11837) );
  NAND2_X1 U11841 ( .A1(n11839), .A2(n11746), .ZN(n11838) );
  NOR2_X1 U11842 ( .A1(n11452), .A2(n8750), .ZN(n11748) );
  NOR2_X1 U11843 ( .A1(n11746), .A2(n11839), .ZN(n11835) );
  INV_X1 U11844 ( .A(n11747), .ZN(n11839) );
  NAND2_X1 U11845 ( .A1(n11743), .A2(n11840), .ZN(n11747) );
  NAND2_X1 U11846 ( .A1(n11742), .A2(n11744), .ZN(n11840) );
  NAND2_X1 U11847 ( .A1(n11841), .A2(n11842), .ZN(n11744) );
  NAND2_X1 U11848 ( .A1(b_19_), .A2(a_13_), .ZN(n11842) );
  INV_X1 U11849 ( .A(n11843), .ZN(n11841) );
  XOR2_X1 U11850 ( .A(n11844), .B(n11845), .Z(n11742) );
  XOR2_X1 U11851 ( .A(n11846), .B(n11847), .Z(n11844) );
  NOR2_X1 U11852 ( .A1(n8438), .A2(n11711), .ZN(n11847) );
  NAND2_X1 U11853 ( .A1(a_13_), .A2(n11843), .ZN(n11743) );
  NAND2_X1 U11854 ( .A1(n11848), .A2(n11849), .ZN(n11843) );
  NAND2_X1 U11855 ( .A1(n11850), .A2(b_19_), .ZN(n11849) );
  NOR2_X1 U11856 ( .A1(n11851), .A2(n8438), .ZN(n11850) );
  NOR2_X1 U11857 ( .A1(n11604), .A2(n11606), .ZN(n11851) );
  NAND2_X1 U11858 ( .A1(n11604), .A2(n11606), .ZN(n11848) );
  NAND2_X1 U11859 ( .A1(n11852), .A2(n11853), .ZN(n11606) );
  NAND2_X1 U11860 ( .A1(n11854), .A2(b_19_), .ZN(n11853) );
  NOR2_X1 U11861 ( .A1(n11855), .A2(n8763), .ZN(n11854) );
  NOR2_X1 U11862 ( .A1(n11613), .A2(n11614), .ZN(n11855) );
  NAND2_X1 U11863 ( .A1(n11613), .A2(n11614), .ZN(n11852) );
  NAND2_X1 U11864 ( .A1(n11622), .A2(n11856), .ZN(n11614) );
  NAND2_X1 U11865 ( .A1(n11621), .A2(n11623), .ZN(n11856) );
  NAND2_X1 U11866 ( .A1(n11857), .A2(n11858), .ZN(n11623) );
  NAND2_X1 U11867 ( .A1(b_19_), .A2(a_16_), .ZN(n11858) );
  INV_X1 U11868 ( .A(n11859), .ZN(n11857) );
  XNOR2_X1 U11869 ( .A(n11860), .B(n11861), .ZN(n11621) );
  NAND2_X1 U11870 ( .A1(n11862), .A2(n11863), .ZN(n11860) );
  NAND2_X1 U11871 ( .A1(a_16_), .A2(n11859), .ZN(n11622) );
  NAND2_X1 U11872 ( .A1(n11630), .A2(n11864), .ZN(n11859) );
  NAND2_X1 U11873 ( .A1(n11629), .A2(n11631), .ZN(n11864) );
  NAND2_X1 U11874 ( .A1(n11865), .A2(n11866), .ZN(n11631) );
  NAND2_X1 U11875 ( .A1(b_19_), .A2(a_17_), .ZN(n11866) );
  INV_X1 U11876 ( .A(n11867), .ZN(n11865) );
  XOR2_X1 U11877 ( .A(n11868), .B(n11869), .Z(n11629) );
  XOR2_X1 U11878 ( .A(n11870), .B(n11871), .Z(n11868) );
  NAND2_X1 U11879 ( .A1(a_17_), .A2(n11867), .ZN(n11630) );
  NAND2_X1 U11880 ( .A1(n11872), .A2(n11873), .ZN(n11867) );
  NAND2_X1 U11881 ( .A1(n11639), .A2(n11874), .ZN(n11873) );
  INV_X1 U11882 ( .A(n11875), .ZN(n11874) );
  NOR2_X1 U11883 ( .A1(n11638), .A2(n11637), .ZN(n11875) );
  NOR2_X1 U11884 ( .A1(n11452), .A2(n10616), .ZN(n11639) );
  NAND2_X1 U11885 ( .A1(n11637), .A2(n11638), .ZN(n11872) );
  NAND2_X1 U11886 ( .A1(n11876), .A2(n11877), .ZN(n11638) );
  NAND2_X1 U11887 ( .A1(n11740), .A2(n11878), .ZN(n11877) );
  INV_X1 U11888 ( .A(n11879), .ZN(n11878) );
  NOR2_X1 U11889 ( .A1(n11737), .A2(n11739), .ZN(n11879) );
  NAND2_X1 U11890 ( .A1(n11739), .A2(n11737), .ZN(n11876) );
  XOR2_X1 U11891 ( .A(n11880), .B(n11881), .Z(n11737) );
  XOR2_X1 U11892 ( .A(n11882), .B(n11883), .Z(n11880) );
  NOR2_X1 U11893 ( .A1(n10633), .A2(n11711), .ZN(n11883) );
  NOR2_X1 U11894 ( .A1(n11884), .A2(n11885), .ZN(n11739) );
  INV_X1 U11895 ( .A(n11886), .ZN(n11885) );
  NAND2_X1 U11896 ( .A1(n11733), .A2(n11887), .ZN(n11886) );
  NAND2_X1 U11897 ( .A1(n11736), .A2(n11735), .ZN(n11887) );
  XOR2_X1 U11898 ( .A(n11888), .B(n11889), .Z(n11733) );
  NAND2_X1 U11899 ( .A1(n11890), .A2(n11891), .ZN(n11888) );
  NOR2_X1 U11900 ( .A1(n11735), .A2(n11736), .ZN(n11884) );
  NOR2_X1 U11901 ( .A1(n11452), .A2(n10633), .ZN(n11736) );
  NAND2_X1 U11902 ( .A1(n11731), .A2(n11892), .ZN(n11735) );
  NAND2_X1 U11903 ( .A1(n11730), .A2(n11732), .ZN(n11892) );
  NAND2_X1 U11904 ( .A1(n11893), .A2(n11894), .ZN(n11732) );
  NAND2_X1 U11905 ( .A1(b_19_), .A2(a_21_), .ZN(n11894) );
  INV_X1 U11906 ( .A(n11895), .ZN(n11893) );
  XNOR2_X1 U11907 ( .A(n11896), .B(n11897), .ZN(n11730) );
  NAND2_X1 U11908 ( .A1(n11898), .A2(n11899), .ZN(n11896) );
  NAND2_X1 U11909 ( .A1(a_21_), .A2(n11895), .ZN(n11731) );
  NAND2_X1 U11910 ( .A1(n11658), .A2(n11900), .ZN(n11895) );
  NAND2_X1 U11911 ( .A1(n11657), .A2(n11659), .ZN(n11900) );
  NAND2_X1 U11912 ( .A1(n11901), .A2(n11902), .ZN(n11659) );
  NAND2_X1 U11913 ( .A1(b_19_), .A2(a_22_), .ZN(n11902) );
  INV_X1 U11914 ( .A(n11903), .ZN(n11901) );
  XOR2_X1 U11915 ( .A(n11904), .B(n11905), .Z(n11657) );
  XOR2_X1 U11916 ( .A(n11906), .B(n11907), .Z(n11904) );
  NOR2_X1 U11917 ( .A1(n8812), .A2(n11711), .ZN(n11907) );
  NAND2_X1 U11918 ( .A1(a_22_), .A2(n11903), .ZN(n11658) );
  NAND2_X1 U11919 ( .A1(n11908), .A2(n11909), .ZN(n11903) );
  NAND2_X1 U11920 ( .A1(n11910), .A2(b_19_), .ZN(n11909) );
  NOR2_X1 U11921 ( .A1(n11911), .A2(n8812), .ZN(n11910) );
  NOR2_X1 U11922 ( .A1(n11665), .A2(n11666), .ZN(n11911) );
  NAND2_X1 U11923 ( .A1(n11665), .A2(n11666), .ZN(n11908) );
  NAND2_X1 U11924 ( .A1(n11912), .A2(n11913), .ZN(n11666) );
  NAND2_X1 U11925 ( .A1(n11728), .A2(n11914), .ZN(n11913) );
  INV_X1 U11926 ( .A(n11915), .ZN(n11914) );
  NOR2_X1 U11927 ( .A1(n11727), .A2(n11726), .ZN(n11915) );
  NOR2_X1 U11928 ( .A1(n11452), .A2(n9131), .ZN(n11728) );
  NAND2_X1 U11929 ( .A1(n11726), .A2(n11727), .ZN(n11912) );
  NAND2_X1 U11930 ( .A1(n11916), .A2(n11917), .ZN(n11727) );
  NAND2_X1 U11931 ( .A1(n11724), .A2(n11918), .ZN(n11917) );
  NAND2_X1 U11932 ( .A1(n11721), .A2(n11723), .ZN(n11918) );
  NOR2_X1 U11933 ( .A1(n11452), .A2(n8825), .ZN(n11724) );
  INV_X1 U11934 ( .A(n11919), .ZN(n11916) );
  NOR2_X1 U11935 ( .A1(n11723), .A2(n11721), .ZN(n11919) );
  XNOR2_X1 U11936 ( .A(n11920), .B(n11921), .ZN(n11721) );
  XNOR2_X1 U11937 ( .A(n11922), .B(n11923), .ZN(n11921) );
  NAND2_X1 U11938 ( .A1(n11924), .A2(n11925), .ZN(n11723) );
  NAND2_X1 U11939 ( .A1(n11680), .A2(n11926), .ZN(n11925) );
  NAND2_X1 U11940 ( .A1(n11683), .A2(n11682), .ZN(n11926) );
  XNOR2_X1 U11941 ( .A(n11927), .B(n11928), .ZN(n11680) );
  XOR2_X1 U11942 ( .A(n11929), .B(n11930), .Z(n11928) );
  INV_X1 U11943 ( .A(n11931), .ZN(n11924) );
  NOR2_X1 U11944 ( .A1(n11682), .A2(n11683), .ZN(n11931) );
  NOR2_X1 U11945 ( .A1(n11452), .A2(n8830), .ZN(n11683) );
  NAND2_X1 U11946 ( .A1(n11932), .A2(n11933), .ZN(n11682) );
  NAND2_X1 U11947 ( .A1(n11690), .A2(n11934), .ZN(n11933) );
  NAND2_X1 U11948 ( .A1(n11689), .A2(n11687), .ZN(n11934) );
  NOR2_X1 U11949 ( .A1(n11452), .A2(n8839), .ZN(n11690) );
  INV_X1 U11950 ( .A(n11935), .ZN(n11932) );
  NOR2_X1 U11951 ( .A1(n11687), .A2(n11689), .ZN(n11935) );
  NOR2_X1 U11952 ( .A1(n11936), .A2(n11937), .ZN(n11689) );
  INV_X1 U11953 ( .A(n11938), .ZN(n11937) );
  NAND2_X1 U11954 ( .A1(n11719), .A2(n11939), .ZN(n11938) );
  NAND2_X1 U11955 ( .A1(n11720), .A2(n11718), .ZN(n11939) );
  NOR2_X1 U11956 ( .A1(n11452), .A2(n8844), .ZN(n11719) );
  NOR2_X1 U11957 ( .A1(n11718), .A2(n11720), .ZN(n11936) );
  NOR2_X1 U11958 ( .A1(n11940), .A2(n11941), .ZN(n11720) );
  INV_X1 U11959 ( .A(n11942), .ZN(n11941) );
  NAND2_X1 U11960 ( .A1(n11713), .A2(n11943), .ZN(n11942) );
  NAND2_X1 U11961 ( .A1(n11944), .A2(n11715), .ZN(n11943) );
  NOR2_X1 U11962 ( .A1(n11452), .A2(n9161), .ZN(n11713) );
  NOR2_X1 U11963 ( .A1(n11715), .A2(n11944), .ZN(n11940) );
  INV_X1 U11964 ( .A(n11716), .ZN(n11944) );
  NAND2_X1 U11965 ( .A1(n11945), .A2(n11946), .ZN(n11716) );
  NAND2_X1 U11966 ( .A1(b_17_), .A2(n11947), .ZN(n11946) );
  NAND2_X1 U11967 ( .A1(n8358), .A2(n11948), .ZN(n11947) );
  NAND2_X1 U11968 ( .A1(a_31_), .A2(n11711), .ZN(n11948) );
  NAND2_X1 U11969 ( .A1(b_18_), .A2(n11949), .ZN(n11945) );
  NAND2_X1 U11970 ( .A1(n8362), .A2(n11950), .ZN(n11949) );
  NAND2_X1 U11971 ( .A1(a_30_), .A2(n11951), .ZN(n11950) );
  NAND2_X1 U11972 ( .A1(n11712), .A2(b_18_), .ZN(n11715) );
  NOR2_X1 U11973 ( .A1(n9170), .A2(n11452), .ZN(n11712) );
  XOR2_X1 U11974 ( .A(n11952), .B(n11953), .Z(n11718) );
  XOR2_X1 U11975 ( .A(n11954), .B(n11955), .Z(n11953) );
  XOR2_X1 U11976 ( .A(n11956), .B(n11957), .Z(n11687) );
  XNOR2_X1 U11977 ( .A(n11958), .B(n11959), .ZN(n11956) );
  XNOR2_X1 U11978 ( .A(n11960), .B(n11961), .ZN(n11726) );
  XNOR2_X1 U11979 ( .A(n11962), .B(n11963), .ZN(n11961) );
  XOR2_X1 U11980 ( .A(n11964), .B(n11965), .Z(n11665) );
  XOR2_X1 U11981 ( .A(n11966), .B(n11967), .Z(n11964) );
  XNOR2_X1 U11982 ( .A(n11968), .B(n11969), .ZN(n11637) );
  NAND2_X1 U11983 ( .A1(n11970), .A2(n11971), .ZN(n11968) );
  XNOR2_X1 U11984 ( .A(n11972), .B(n11973), .ZN(n11613) );
  NAND2_X1 U11985 ( .A1(n11974), .A2(n11975), .ZN(n11972) );
  XNOR2_X1 U11986 ( .A(n11976), .B(n11977), .ZN(n11604) );
  XOR2_X1 U11987 ( .A(n11978), .B(n11979), .Z(n11977) );
  NAND2_X1 U11988 ( .A1(b_18_), .A2(a_15_), .ZN(n11979) );
  XOR2_X1 U11989 ( .A(n11980), .B(n11981), .Z(n11746) );
  NAND2_X1 U11990 ( .A1(n11982), .A2(n11983), .ZN(n11980) );
  XNOR2_X1 U11991 ( .A(n11984), .B(n11985), .ZN(n11750) );
  XOR2_X1 U11992 ( .A(n11986), .B(n11987), .Z(n11984) );
  NOR2_X1 U11993 ( .A1(n8750), .A2(n11711), .ZN(n11987) );
  XNOR2_X1 U11994 ( .A(n11988), .B(n11989), .ZN(n11753) );
  XOR2_X1 U11995 ( .A(n11990), .B(n11991), .Z(n11989) );
  NAND2_X1 U11996 ( .A1(b_18_), .A2(a_11_), .ZN(n11991) );
  XNOR2_X1 U11997 ( .A(n11992), .B(n11993), .ZN(n11580) );
  NAND2_X1 U11998 ( .A1(n11994), .A2(n11995), .ZN(n11992) );
  XNOR2_X1 U11999 ( .A(n11996), .B(n11997), .ZN(n11506) );
  XNOR2_X1 U12000 ( .A(n11998), .B(n11999), .ZN(n11996) );
  NAND2_X1 U12001 ( .A1(n8576), .A2(n8575), .ZN(n8574) );
  INV_X1 U12002 ( .A(n12000), .ZN(n8575) );
  NAND2_X1 U12003 ( .A1(n12001), .A2(n12002), .ZN(n12000) );
  NAND2_X1 U12004 ( .A1(n12003), .A2(n12004), .ZN(n12001) );
  INV_X1 U12005 ( .A(n12005), .ZN(n12004) );
  XOR2_X1 U12006 ( .A(n12006), .B(n12007), .Z(n12003) );
  NOR2_X1 U12007 ( .A1(n8640), .A2(n8641), .ZN(n8576) );
  XNOR2_X1 U12008 ( .A(n12008), .B(n12009), .ZN(n8641) );
  XOR2_X1 U12009 ( .A(n12010), .B(n12011), .Z(n12008) );
  NOR2_X1 U12010 ( .A1(n8690), .A2(n11951), .ZN(n12011) );
  NOR2_X1 U12011 ( .A1(n12012), .A2(n12013), .ZN(n8640) );
  NOR2_X1 U12012 ( .A1(n11511), .A2(n12014), .ZN(n12013) );
  INV_X1 U12013 ( .A(n12015), .ZN(n12014) );
  NAND2_X1 U12014 ( .A1(n11510), .A2(n11508), .ZN(n12015) );
  NAND2_X1 U12015 ( .A1(b_18_), .A2(a_0_), .ZN(n11511) );
  NOR2_X1 U12016 ( .A1(n11508), .A2(n11510), .ZN(n12012) );
  NOR2_X1 U12017 ( .A1(n12016), .A2(n12017), .ZN(n11510) );
  INV_X1 U12018 ( .A(n12018), .ZN(n12017) );
  NAND2_X1 U12019 ( .A1(n11999), .A2(n12019), .ZN(n12018) );
  NAND2_X1 U12020 ( .A1(n11997), .A2(n11998), .ZN(n12019) );
  NOR2_X1 U12021 ( .A1(n11711), .A2(n8502), .ZN(n11999) );
  NOR2_X1 U12022 ( .A1(n11997), .A2(n11998), .ZN(n12016) );
  NOR2_X1 U12023 ( .A1(n12020), .A2(n12021), .ZN(n11998) );
  INV_X1 U12024 ( .A(n12022), .ZN(n12021) );
  NAND2_X1 U12025 ( .A1(n11766), .A2(n12023), .ZN(n12022) );
  NAND2_X1 U12026 ( .A1(n11764), .A2(n11765), .ZN(n12023) );
  NOR2_X1 U12027 ( .A1(n11711), .A2(n8497), .ZN(n11766) );
  NOR2_X1 U12028 ( .A1(n11764), .A2(n11765), .ZN(n12020) );
  NAND2_X1 U12029 ( .A1(n12024), .A2(n12025), .ZN(n11765) );
  NAND2_X1 U12030 ( .A1(n11771), .A2(n12026), .ZN(n12025) );
  NAND2_X1 U12031 ( .A1(n11774), .A2(n11773), .ZN(n12026) );
  XNOR2_X1 U12032 ( .A(n12027), .B(n12028), .ZN(n11771) );
  XNOR2_X1 U12033 ( .A(n12029), .B(n12030), .ZN(n12028) );
  NAND2_X1 U12034 ( .A1(b_17_), .A2(a_4_), .ZN(n12030) );
  INV_X1 U12035 ( .A(n12031), .ZN(n12024) );
  NOR2_X1 U12036 ( .A1(n11773), .A2(n11774), .ZN(n12031) );
  NOR2_X1 U12037 ( .A1(n11711), .A2(n8707), .ZN(n11774) );
  NAND2_X1 U12038 ( .A1(n11781), .A2(n12032), .ZN(n11773) );
  NAND2_X1 U12039 ( .A1(n11780), .A2(n11782), .ZN(n12032) );
  NAND2_X1 U12040 ( .A1(n12033), .A2(n12034), .ZN(n11782) );
  NAND2_X1 U12041 ( .A1(b_18_), .A2(a_4_), .ZN(n12034) );
  INV_X1 U12042 ( .A(n12035), .ZN(n12033) );
  XOR2_X1 U12043 ( .A(n12036), .B(n12037), .Z(n11780) );
  XNOR2_X1 U12044 ( .A(n12038), .B(n12039), .ZN(n12037) );
  NAND2_X1 U12045 ( .A1(a_4_), .A2(n12035), .ZN(n11781) );
  NAND2_X1 U12046 ( .A1(n12040), .A2(n12041), .ZN(n12035) );
  NAND2_X1 U12047 ( .A1(n12042), .A2(b_18_), .ZN(n12041) );
  NOR2_X1 U12048 ( .A1(n12043), .A2(n8717), .ZN(n12042) );
  NOR2_X1 U12049 ( .A1(n11788), .A2(n11789), .ZN(n12043) );
  NAND2_X1 U12050 ( .A1(n11788), .A2(n11789), .ZN(n12040) );
  NAND2_X1 U12051 ( .A1(n11797), .A2(n12044), .ZN(n11789) );
  NAND2_X1 U12052 ( .A1(n11796), .A2(n11798), .ZN(n12044) );
  NAND2_X1 U12053 ( .A1(n12045), .A2(n12046), .ZN(n11798) );
  INV_X1 U12054 ( .A(n12047), .ZN(n12046) );
  NAND2_X1 U12055 ( .A1(b_18_), .A2(a_6_), .ZN(n12045) );
  XNOR2_X1 U12056 ( .A(n12048), .B(n12049), .ZN(n11796) );
  NAND2_X1 U12057 ( .A1(n12050), .A2(n12051), .ZN(n12048) );
  NAND2_X1 U12058 ( .A1(n12047), .A2(a_6_), .ZN(n11797) );
  NOR2_X1 U12059 ( .A1(n12052), .A2(n12053), .ZN(n12047) );
  INV_X1 U12060 ( .A(n12054), .ZN(n12053) );
  NAND2_X1 U12061 ( .A1(n11803), .A2(n12055), .ZN(n12054) );
  NAND2_X1 U12062 ( .A1(n11806), .A2(n11805), .ZN(n12055) );
  XNOR2_X1 U12063 ( .A(n12056), .B(n12057), .ZN(n11803) );
  XNOR2_X1 U12064 ( .A(n12058), .B(n12059), .ZN(n12057) );
  NOR2_X1 U12065 ( .A1(n11805), .A2(n11806), .ZN(n12052) );
  NOR2_X1 U12066 ( .A1(n11711), .A2(n8726), .ZN(n11806) );
  NAND2_X1 U12067 ( .A1(n11813), .A2(n12060), .ZN(n11805) );
  NAND2_X1 U12068 ( .A1(n11812), .A2(n11814), .ZN(n12060) );
  NAND2_X1 U12069 ( .A1(n12061), .A2(n12062), .ZN(n11814) );
  INV_X1 U12070 ( .A(n12063), .ZN(n12062) );
  NAND2_X1 U12071 ( .A1(b_18_), .A2(a_8_), .ZN(n12061) );
  XNOR2_X1 U12072 ( .A(n12064), .B(n12065), .ZN(n11812) );
  NAND2_X1 U12073 ( .A1(n12066), .A2(n12067), .ZN(n12064) );
  NAND2_X1 U12074 ( .A1(n12063), .A2(a_8_), .ZN(n11813) );
  NOR2_X1 U12075 ( .A1(n12068), .A2(n12069), .ZN(n12063) );
  INV_X1 U12076 ( .A(n12070), .ZN(n12069) );
  NAND2_X1 U12077 ( .A1(n11820), .A2(n12071), .ZN(n12070) );
  NAND2_X1 U12078 ( .A1(n11822), .A2(n11821), .ZN(n12071) );
  XNOR2_X1 U12079 ( .A(n12072), .B(n12073), .ZN(n11820) );
  XNOR2_X1 U12080 ( .A(n12074), .B(n12075), .ZN(n12073) );
  NOR2_X1 U12081 ( .A1(n11821), .A2(n11822), .ZN(n12068) );
  NOR2_X1 U12082 ( .A1(n11711), .A2(n8736), .ZN(n11822) );
  NAND2_X1 U12083 ( .A1(n11994), .A2(n12076), .ZN(n11821) );
  NAND2_X1 U12084 ( .A1(n11993), .A2(n11995), .ZN(n12076) );
  NAND2_X1 U12085 ( .A1(n12077), .A2(n12078), .ZN(n11995) );
  NAND2_X1 U12086 ( .A1(b_18_), .A2(a_10_), .ZN(n12078) );
  INV_X1 U12087 ( .A(n12079), .ZN(n12077) );
  XNOR2_X1 U12088 ( .A(n12080), .B(n12081), .ZN(n11993) );
  XOR2_X1 U12089 ( .A(n12082), .B(n12083), .Z(n12081) );
  NAND2_X1 U12090 ( .A1(b_17_), .A2(a_11_), .ZN(n12083) );
  NAND2_X1 U12091 ( .A1(a_10_), .A2(n12079), .ZN(n11994) );
  NAND2_X1 U12092 ( .A1(n12084), .A2(n12085), .ZN(n12079) );
  NAND2_X1 U12093 ( .A1(n12086), .A2(b_18_), .ZN(n12085) );
  NOR2_X1 U12094 ( .A1(n12087), .A2(n8452), .ZN(n12086) );
  NOR2_X1 U12095 ( .A1(n11990), .A2(n11988), .ZN(n12087) );
  NAND2_X1 U12096 ( .A1(n11988), .A2(n11990), .ZN(n12084) );
  NAND2_X1 U12097 ( .A1(n12088), .A2(n12089), .ZN(n11990) );
  NAND2_X1 U12098 ( .A1(n12090), .A2(b_18_), .ZN(n12089) );
  NOR2_X1 U12099 ( .A1(n12091), .A2(n8750), .ZN(n12090) );
  NOR2_X1 U12100 ( .A1(n11986), .A2(n11985), .ZN(n12091) );
  NAND2_X1 U12101 ( .A1(n11985), .A2(n11986), .ZN(n12088) );
  NAND2_X1 U12102 ( .A1(n11982), .A2(n12092), .ZN(n11986) );
  NAND2_X1 U12103 ( .A1(n11981), .A2(n11983), .ZN(n12092) );
  NAND2_X1 U12104 ( .A1(n12093), .A2(n12094), .ZN(n11983) );
  NAND2_X1 U12105 ( .A1(b_18_), .A2(a_13_), .ZN(n12094) );
  INV_X1 U12106 ( .A(n12095), .ZN(n12093) );
  XNOR2_X1 U12107 ( .A(n12096), .B(n12097), .ZN(n11981) );
  XOR2_X1 U12108 ( .A(n12098), .B(n12099), .Z(n12097) );
  NAND2_X1 U12109 ( .A1(a_13_), .A2(n12095), .ZN(n11982) );
  NAND2_X1 U12110 ( .A1(n12100), .A2(n12101), .ZN(n12095) );
  NAND2_X1 U12111 ( .A1(n12102), .A2(b_18_), .ZN(n12101) );
  NOR2_X1 U12112 ( .A1(n12103), .A2(n8438), .ZN(n12102) );
  NOR2_X1 U12113 ( .A1(n11846), .A2(n11845), .ZN(n12103) );
  NAND2_X1 U12114 ( .A1(n11845), .A2(n11846), .ZN(n12100) );
  NAND2_X1 U12115 ( .A1(n12104), .A2(n12105), .ZN(n11846) );
  NAND2_X1 U12116 ( .A1(n12106), .A2(b_18_), .ZN(n12105) );
  NOR2_X1 U12117 ( .A1(n12107), .A2(n8763), .ZN(n12106) );
  NOR2_X1 U12118 ( .A1(n11976), .A2(n11978), .ZN(n12107) );
  NAND2_X1 U12119 ( .A1(n11976), .A2(n11978), .ZN(n12104) );
  NAND2_X1 U12120 ( .A1(n11974), .A2(n12108), .ZN(n11978) );
  NAND2_X1 U12121 ( .A1(n11973), .A2(n11975), .ZN(n12108) );
  NAND2_X1 U12122 ( .A1(n12109), .A2(n12110), .ZN(n11975) );
  NAND2_X1 U12123 ( .A1(b_18_), .A2(a_16_), .ZN(n12110) );
  INV_X1 U12124 ( .A(n12111), .ZN(n12109) );
  XOR2_X1 U12125 ( .A(n12112), .B(n12113), .Z(n11973) );
  XNOR2_X1 U12126 ( .A(n12114), .B(n12115), .ZN(n12113) );
  NAND2_X1 U12127 ( .A1(a_16_), .A2(n12111), .ZN(n11974) );
  NAND2_X1 U12128 ( .A1(n11862), .A2(n12116), .ZN(n12111) );
  NAND2_X1 U12129 ( .A1(n11861), .A2(n11863), .ZN(n12116) );
  NAND2_X1 U12130 ( .A1(n12117), .A2(n12118), .ZN(n11863) );
  NAND2_X1 U12131 ( .A1(b_18_), .A2(a_17_), .ZN(n12118) );
  INV_X1 U12132 ( .A(n12119), .ZN(n12117) );
  XNOR2_X1 U12133 ( .A(n12120), .B(n12121), .ZN(n11861) );
  XOR2_X1 U12134 ( .A(n12122), .B(n12123), .Z(n12121) );
  NAND2_X1 U12135 ( .A1(b_17_), .A2(a_18_), .ZN(n12123) );
  NAND2_X1 U12136 ( .A1(a_17_), .A2(n12119), .ZN(n11862) );
  NAND2_X1 U12137 ( .A1(n12124), .A2(n12125), .ZN(n12119) );
  NAND2_X1 U12138 ( .A1(n11871), .A2(n12126), .ZN(n12125) );
  INV_X1 U12139 ( .A(n12127), .ZN(n12126) );
  NOR2_X1 U12140 ( .A1(n11870), .A2(n11869), .ZN(n12127) );
  NAND2_X1 U12141 ( .A1(n11869), .A2(n11870), .ZN(n12124) );
  NAND2_X1 U12142 ( .A1(n11970), .A2(n12128), .ZN(n11870) );
  NAND2_X1 U12143 ( .A1(n11969), .A2(n11971), .ZN(n12128) );
  NAND2_X1 U12144 ( .A1(n12129), .A2(n12130), .ZN(n11971) );
  NAND2_X1 U12145 ( .A1(b_18_), .A2(a_19_), .ZN(n12130) );
  INV_X1 U12146 ( .A(n12131), .ZN(n12129) );
  XNOR2_X1 U12147 ( .A(n12132), .B(n12133), .ZN(n11969) );
  XOR2_X1 U12148 ( .A(n12134), .B(n12135), .Z(n12132) );
  NAND2_X1 U12149 ( .A1(a_19_), .A2(n12131), .ZN(n11970) );
  NAND2_X1 U12150 ( .A1(n12136), .A2(n12137), .ZN(n12131) );
  NAND2_X1 U12151 ( .A1(n12138), .A2(b_18_), .ZN(n12137) );
  NOR2_X1 U12152 ( .A1(n12139), .A2(n10633), .ZN(n12138) );
  NOR2_X1 U12153 ( .A1(n11882), .A2(n11881), .ZN(n12139) );
  NAND2_X1 U12154 ( .A1(n11881), .A2(n11882), .ZN(n12136) );
  NAND2_X1 U12155 ( .A1(n11890), .A2(n12140), .ZN(n11882) );
  NAND2_X1 U12156 ( .A1(n11889), .A2(n11891), .ZN(n12140) );
  NAND2_X1 U12157 ( .A1(n12141), .A2(n12142), .ZN(n11891) );
  NAND2_X1 U12158 ( .A1(b_18_), .A2(a_21_), .ZN(n12142) );
  INV_X1 U12159 ( .A(n12143), .ZN(n12141) );
  XOR2_X1 U12160 ( .A(n12144), .B(n12145), .Z(n11889) );
  XOR2_X1 U12161 ( .A(n12146), .B(n12147), .Z(n12144) );
  NOR2_X1 U12162 ( .A1(n8803), .A2(n11951), .ZN(n12147) );
  NAND2_X1 U12163 ( .A1(a_21_), .A2(n12143), .ZN(n11890) );
  NAND2_X1 U12164 ( .A1(n11898), .A2(n12148), .ZN(n12143) );
  NAND2_X1 U12165 ( .A1(n11897), .A2(n11899), .ZN(n12148) );
  NAND2_X1 U12166 ( .A1(n12149), .A2(n12150), .ZN(n11899) );
  NAND2_X1 U12167 ( .A1(b_18_), .A2(a_22_), .ZN(n12150) );
  INV_X1 U12168 ( .A(n12151), .ZN(n12149) );
  XOR2_X1 U12169 ( .A(n12152), .B(n12153), .Z(n11897) );
  XOR2_X1 U12170 ( .A(n12154), .B(n12155), .Z(n12152) );
  NOR2_X1 U12171 ( .A1(n8812), .A2(n11951), .ZN(n12155) );
  NAND2_X1 U12172 ( .A1(a_22_), .A2(n12151), .ZN(n11898) );
  NAND2_X1 U12173 ( .A1(n12156), .A2(n12157), .ZN(n12151) );
  NAND2_X1 U12174 ( .A1(n12158), .A2(b_18_), .ZN(n12157) );
  NOR2_X1 U12175 ( .A1(n12159), .A2(n8812), .ZN(n12158) );
  NOR2_X1 U12176 ( .A1(n11905), .A2(n11906), .ZN(n12159) );
  NAND2_X1 U12177 ( .A1(n11905), .A2(n11906), .ZN(n12156) );
  NAND2_X1 U12178 ( .A1(n12160), .A2(n12161), .ZN(n11906) );
  NAND2_X1 U12179 ( .A1(n11967), .A2(n12162), .ZN(n12161) );
  INV_X1 U12180 ( .A(n12163), .ZN(n12162) );
  NOR2_X1 U12181 ( .A1(n11965), .A2(n11966), .ZN(n12163) );
  NOR2_X1 U12182 ( .A1(n11711), .A2(n9131), .ZN(n11967) );
  NAND2_X1 U12183 ( .A1(n11965), .A2(n11966), .ZN(n12160) );
  NAND2_X1 U12184 ( .A1(n12164), .A2(n12165), .ZN(n11966) );
  NAND2_X1 U12185 ( .A1(n11963), .A2(n12166), .ZN(n12165) );
  NAND2_X1 U12186 ( .A1(n11960), .A2(n11962), .ZN(n12166) );
  NOR2_X1 U12187 ( .A1(n11711), .A2(n8825), .ZN(n11963) );
  INV_X1 U12188 ( .A(n12167), .ZN(n12164) );
  NOR2_X1 U12189 ( .A1(n11962), .A2(n11960), .ZN(n12167) );
  XNOR2_X1 U12190 ( .A(n12168), .B(n12169), .ZN(n11960) );
  XNOR2_X1 U12191 ( .A(n12170), .B(n12171), .ZN(n12169) );
  NAND2_X1 U12192 ( .A1(n12172), .A2(n12173), .ZN(n11962) );
  NAND2_X1 U12193 ( .A1(n11920), .A2(n12174), .ZN(n12173) );
  NAND2_X1 U12194 ( .A1(n11923), .A2(n11922), .ZN(n12174) );
  XNOR2_X1 U12195 ( .A(n12175), .B(n12176), .ZN(n11920) );
  XOR2_X1 U12196 ( .A(n12177), .B(n12178), .Z(n12176) );
  INV_X1 U12197 ( .A(n12179), .ZN(n12172) );
  NOR2_X1 U12198 ( .A1(n11922), .A2(n11923), .ZN(n12179) );
  NOR2_X1 U12199 ( .A1(n11711), .A2(n8830), .ZN(n11923) );
  NAND2_X1 U12200 ( .A1(n12180), .A2(n12181), .ZN(n11922) );
  NAND2_X1 U12201 ( .A1(n11930), .A2(n12182), .ZN(n12181) );
  NAND2_X1 U12202 ( .A1(n11927), .A2(n11929), .ZN(n12182) );
  NOR2_X1 U12203 ( .A1(n11711), .A2(n8839), .ZN(n11930) );
  INV_X1 U12204 ( .A(n12183), .ZN(n12180) );
  NOR2_X1 U12205 ( .A1(n11927), .A2(n11929), .ZN(n12183) );
  NOR2_X1 U12206 ( .A1(n12184), .A2(n12185), .ZN(n11929) );
  INV_X1 U12207 ( .A(n12186), .ZN(n12185) );
  NAND2_X1 U12208 ( .A1(n11958), .A2(n12187), .ZN(n12186) );
  NAND2_X1 U12209 ( .A1(n11959), .A2(n11957), .ZN(n12187) );
  NOR2_X1 U12210 ( .A1(n11711), .A2(n8844), .ZN(n11958) );
  NOR2_X1 U12211 ( .A1(n11957), .A2(n11959), .ZN(n12184) );
  NOR2_X1 U12212 ( .A1(n12188), .A2(n12189), .ZN(n11959) );
  INV_X1 U12213 ( .A(n12190), .ZN(n12189) );
  NAND2_X1 U12214 ( .A1(n11952), .A2(n12191), .ZN(n12190) );
  NAND2_X1 U12215 ( .A1(n12192), .A2(n11954), .ZN(n12191) );
  NOR2_X1 U12216 ( .A1(n11711), .A2(n9161), .ZN(n11952) );
  NOR2_X1 U12217 ( .A1(n11954), .A2(n12192), .ZN(n12188) );
  INV_X1 U12218 ( .A(n11955), .ZN(n12192) );
  NAND2_X1 U12219 ( .A1(n12193), .A2(n12194), .ZN(n11955) );
  NAND2_X1 U12220 ( .A1(b_16_), .A2(n12195), .ZN(n12194) );
  NAND2_X1 U12221 ( .A1(n8358), .A2(n12196), .ZN(n12195) );
  NAND2_X1 U12222 ( .A1(a_31_), .A2(n11951), .ZN(n12196) );
  NAND2_X1 U12223 ( .A1(b_17_), .A2(n12197), .ZN(n12193) );
  NAND2_X1 U12224 ( .A1(n8362), .A2(n12198), .ZN(n12197) );
  NAND2_X1 U12225 ( .A1(a_30_), .A2(n12199), .ZN(n12198) );
  NAND2_X1 U12226 ( .A1(n12200), .A2(b_18_), .ZN(n11954) );
  NOR2_X1 U12227 ( .A1(n9170), .A2(n11951), .ZN(n12200) );
  XOR2_X1 U12228 ( .A(n12201), .B(n12202), .Z(n11957) );
  XOR2_X1 U12229 ( .A(n12203), .B(n12204), .Z(n12202) );
  XOR2_X1 U12230 ( .A(n12205), .B(n12206), .Z(n11927) );
  XNOR2_X1 U12231 ( .A(n12207), .B(n12208), .ZN(n12205) );
  XNOR2_X1 U12232 ( .A(n12209), .B(n12210), .ZN(n11965) );
  XNOR2_X1 U12233 ( .A(n12211), .B(n12212), .ZN(n12210) );
  XOR2_X1 U12234 ( .A(n12213), .B(n12214), .Z(n11905) );
  XOR2_X1 U12235 ( .A(n12215), .B(n12216), .Z(n12213) );
  XNOR2_X1 U12236 ( .A(n12217), .B(n12218), .ZN(n11881) );
  NAND2_X1 U12237 ( .A1(n12219), .A2(n12220), .ZN(n12217) );
  XOR2_X1 U12238 ( .A(n12221), .B(n12222), .Z(n11869) );
  XNOR2_X1 U12239 ( .A(n12223), .B(n12224), .ZN(n12222) );
  NAND2_X1 U12240 ( .A1(b_17_), .A2(a_19_), .ZN(n12224) );
  XNOR2_X1 U12241 ( .A(n12225), .B(n12226), .ZN(n11976) );
  XOR2_X1 U12242 ( .A(n12227), .B(n12228), .Z(n12225) );
  XNOR2_X1 U12243 ( .A(n12229), .B(n12230), .ZN(n11845) );
  XNOR2_X1 U12244 ( .A(n12231), .B(n12232), .ZN(n12230) );
  XNOR2_X1 U12245 ( .A(n12233), .B(n12234), .ZN(n11985) );
  XNOR2_X1 U12246 ( .A(n12235), .B(n12236), .ZN(n12234) );
  XOR2_X1 U12247 ( .A(n12237), .B(n12238), .Z(n11988) );
  XOR2_X1 U12248 ( .A(n12239), .B(n12240), .Z(n12237) );
  NOR2_X1 U12249 ( .A1(n8750), .A2(n11951), .ZN(n12240) );
  XOR2_X1 U12250 ( .A(n12241), .B(n12242), .Z(n11788) );
  XOR2_X1 U12251 ( .A(n12243), .B(n12244), .Z(n12241) );
  NOR2_X1 U12252 ( .A1(n8480), .A2(n11951), .ZN(n12244) );
  XOR2_X1 U12253 ( .A(n12245), .B(n12246), .Z(n11764) );
  NAND2_X1 U12254 ( .A1(n12247), .A2(n12248), .ZN(n12245) );
  XNOR2_X1 U12255 ( .A(n12249), .B(n12250), .ZN(n11997) );
  XOR2_X1 U12256 ( .A(n12251), .B(n12252), .Z(n12249) );
  NOR2_X1 U12257 ( .A1(n8497), .A2(n11951), .ZN(n12252) );
  XOR2_X1 U12258 ( .A(n12253), .B(n12254), .Z(n11508) );
  NAND2_X1 U12259 ( .A1(n12255), .A2(n12256), .ZN(n12253) );
  NAND2_X1 U12260 ( .A1(n12257), .A2(n12002), .ZN(n8581) );
  XNOR2_X1 U12261 ( .A(n12258), .B(n12259), .ZN(n12257) );
  NOR2_X1 U12262 ( .A1(n12260), .A2(n12002), .ZN(n8580) );
  NAND2_X1 U12263 ( .A1(n12261), .A2(n12005), .ZN(n12002) );
  NAND2_X1 U12264 ( .A1(n12262), .A2(n12263), .ZN(n12005) );
  NAND2_X1 U12265 ( .A1(n12264), .A2(b_17_), .ZN(n12263) );
  NOR2_X1 U12266 ( .A1(n12265), .A2(n8690), .ZN(n12264) );
  NOR2_X1 U12267 ( .A1(n12009), .A2(n12010), .ZN(n12265) );
  NAND2_X1 U12268 ( .A1(n12009), .A2(n12010), .ZN(n12262) );
  NAND2_X1 U12269 ( .A1(n12255), .A2(n12266), .ZN(n12010) );
  NAND2_X1 U12270 ( .A1(n12254), .A2(n12256), .ZN(n12266) );
  NAND2_X1 U12271 ( .A1(n12267), .A2(n12268), .ZN(n12256) );
  NAND2_X1 U12272 ( .A1(b_17_), .A2(a_1_), .ZN(n12268) );
  INV_X1 U12273 ( .A(n12269), .ZN(n12267) );
  XNOR2_X1 U12274 ( .A(n12270), .B(n12271), .ZN(n12254) );
  XOR2_X1 U12275 ( .A(n12272), .B(n12273), .Z(n12270) );
  NAND2_X1 U12276 ( .A1(a_1_), .A2(n12269), .ZN(n12255) );
  NAND2_X1 U12277 ( .A1(n12274), .A2(n12275), .ZN(n12269) );
  NAND2_X1 U12278 ( .A1(n12276), .A2(b_17_), .ZN(n12275) );
  NOR2_X1 U12279 ( .A1(n12277), .A2(n8497), .ZN(n12276) );
  NOR2_X1 U12280 ( .A1(n12250), .A2(n12251), .ZN(n12277) );
  NAND2_X1 U12281 ( .A1(n12250), .A2(n12251), .ZN(n12274) );
  NAND2_X1 U12282 ( .A1(n12247), .A2(n12278), .ZN(n12251) );
  NAND2_X1 U12283 ( .A1(n12246), .A2(n12248), .ZN(n12278) );
  NAND2_X1 U12284 ( .A1(n12279), .A2(n12280), .ZN(n12248) );
  NAND2_X1 U12285 ( .A1(b_17_), .A2(a_3_), .ZN(n12280) );
  INV_X1 U12286 ( .A(n12281), .ZN(n12279) );
  XNOR2_X1 U12287 ( .A(n12282), .B(n12283), .ZN(n12246) );
  XOR2_X1 U12288 ( .A(n12284), .B(n12285), .Z(n12282) );
  NAND2_X1 U12289 ( .A1(a_3_), .A2(n12281), .ZN(n12247) );
  NAND2_X1 U12290 ( .A1(n12286), .A2(n12287), .ZN(n12281) );
  NAND2_X1 U12291 ( .A1(n12288), .A2(b_17_), .ZN(n12287) );
  NOR2_X1 U12292 ( .A1(n12289), .A2(n8712), .ZN(n12288) );
  NOR2_X1 U12293 ( .A1(n12029), .A2(n12027), .ZN(n12289) );
  NAND2_X1 U12294 ( .A1(n12029), .A2(n12027), .ZN(n12286) );
  XNOR2_X1 U12295 ( .A(n12290), .B(n12291), .ZN(n12027) );
  NAND2_X1 U12296 ( .A1(n12292), .A2(n12293), .ZN(n12290) );
  NOR2_X1 U12297 ( .A1(n12294), .A2(n12295), .ZN(n12029) );
  INV_X1 U12298 ( .A(n12296), .ZN(n12295) );
  NAND2_X1 U12299 ( .A1(n12036), .A2(n12297), .ZN(n12296) );
  NAND2_X1 U12300 ( .A1(n12039), .A2(n12038), .ZN(n12297) );
  XNOR2_X1 U12301 ( .A(n12298), .B(n12299), .ZN(n12036) );
  XOR2_X1 U12302 ( .A(n12300), .B(n12301), .Z(n12298) );
  NOR2_X1 U12303 ( .A1(n8480), .A2(n12199), .ZN(n12301) );
  NOR2_X1 U12304 ( .A1(n12038), .A2(n12039), .ZN(n12294) );
  NOR2_X1 U12305 ( .A1(n11951), .A2(n8717), .ZN(n12039) );
  NAND2_X1 U12306 ( .A1(n12302), .A2(n12303), .ZN(n12038) );
  NAND2_X1 U12307 ( .A1(n12304), .A2(b_17_), .ZN(n12303) );
  NOR2_X1 U12308 ( .A1(n12305), .A2(n8480), .ZN(n12304) );
  NOR2_X1 U12309 ( .A1(n12242), .A2(n12243), .ZN(n12305) );
  NAND2_X1 U12310 ( .A1(n12242), .A2(n12243), .ZN(n12302) );
  NAND2_X1 U12311 ( .A1(n12050), .A2(n12306), .ZN(n12243) );
  NAND2_X1 U12312 ( .A1(n12049), .A2(n12051), .ZN(n12306) );
  NAND2_X1 U12313 ( .A1(n12307), .A2(n12308), .ZN(n12051) );
  INV_X1 U12314 ( .A(n12309), .ZN(n12308) );
  NAND2_X1 U12315 ( .A1(b_17_), .A2(a_7_), .ZN(n12307) );
  XOR2_X1 U12316 ( .A(n12310), .B(n12311), .Z(n12049) );
  XNOR2_X1 U12317 ( .A(n12312), .B(n12313), .ZN(n12311) );
  NAND2_X1 U12318 ( .A1(b_16_), .A2(a_8_), .ZN(n12313) );
  NAND2_X1 U12319 ( .A1(n12309), .A2(a_7_), .ZN(n12050) );
  NOR2_X1 U12320 ( .A1(n12314), .A2(n12315), .ZN(n12309) );
  INV_X1 U12321 ( .A(n12316), .ZN(n12315) );
  NAND2_X1 U12322 ( .A1(n12056), .A2(n12317), .ZN(n12316) );
  NAND2_X1 U12323 ( .A1(n12059), .A2(n12058), .ZN(n12317) );
  XOR2_X1 U12324 ( .A(n12318), .B(n12319), .Z(n12056) );
  XOR2_X1 U12325 ( .A(n12320), .B(n12321), .Z(n12318) );
  NOR2_X1 U12326 ( .A1(n12058), .A2(n12059), .ZN(n12314) );
  NOR2_X1 U12327 ( .A1(n11951), .A2(n8731), .ZN(n12059) );
  NAND2_X1 U12328 ( .A1(n12066), .A2(n12322), .ZN(n12058) );
  NAND2_X1 U12329 ( .A1(n12065), .A2(n12067), .ZN(n12322) );
  NAND2_X1 U12330 ( .A1(n12323), .A2(n12324), .ZN(n12067) );
  INV_X1 U12331 ( .A(n12325), .ZN(n12324) );
  NAND2_X1 U12332 ( .A1(b_17_), .A2(a_9_), .ZN(n12323) );
  XNOR2_X1 U12333 ( .A(n12326), .B(n12327), .ZN(n12065) );
  NAND2_X1 U12334 ( .A1(n12328), .A2(n12329), .ZN(n12326) );
  NAND2_X1 U12335 ( .A1(n12325), .A2(a_9_), .ZN(n12066) );
  NOR2_X1 U12336 ( .A1(n12330), .A2(n12331), .ZN(n12325) );
  INV_X1 U12337 ( .A(n12332), .ZN(n12331) );
  NAND2_X1 U12338 ( .A1(n12072), .A2(n12333), .ZN(n12332) );
  NAND2_X1 U12339 ( .A1(n12075), .A2(n12074), .ZN(n12333) );
  XOR2_X1 U12340 ( .A(n12334), .B(n12335), .Z(n12072) );
  NAND2_X1 U12341 ( .A1(n12336), .A2(n12337), .ZN(n12334) );
  NOR2_X1 U12342 ( .A1(n12074), .A2(n12075), .ZN(n12330) );
  NOR2_X1 U12343 ( .A1(n11951), .A2(n8741), .ZN(n12075) );
  NAND2_X1 U12344 ( .A1(n12338), .A2(n12339), .ZN(n12074) );
  NAND2_X1 U12345 ( .A1(n12340), .A2(b_17_), .ZN(n12339) );
  NOR2_X1 U12346 ( .A1(n12341), .A2(n8452), .ZN(n12340) );
  NOR2_X1 U12347 ( .A1(n12080), .A2(n12082), .ZN(n12341) );
  NAND2_X1 U12348 ( .A1(n12080), .A2(n12082), .ZN(n12338) );
  NAND2_X1 U12349 ( .A1(n12342), .A2(n12343), .ZN(n12082) );
  NAND2_X1 U12350 ( .A1(n12344), .A2(b_17_), .ZN(n12343) );
  NOR2_X1 U12351 ( .A1(n12345), .A2(n8750), .ZN(n12344) );
  NOR2_X1 U12352 ( .A1(n12238), .A2(n12239), .ZN(n12345) );
  NAND2_X1 U12353 ( .A1(n12238), .A2(n12239), .ZN(n12342) );
  NAND2_X1 U12354 ( .A1(n12346), .A2(n12347), .ZN(n12239) );
  NAND2_X1 U12355 ( .A1(n12236), .A2(n12348), .ZN(n12347) );
  INV_X1 U12356 ( .A(n12349), .ZN(n12348) );
  NOR2_X1 U12357 ( .A1(n12235), .A2(n12233), .ZN(n12349) );
  NOR2_X1 U12358 ( .A1(n11951), .A2(n8443), .ZN(n12236) );
  NAND2_X1 U12359 ( .A1(n12233), .A2(n12235), .ZN(n12346) );
  NAND2_X1 U12360 ( .A1(n12350), .A2(n12351), .ZN(n12235) );
  INV_X1 U12361 ( .A(n12352), .ZN(n12351) );
  NOR2_X1 U12362 ( .A1(n12099), .A2(n12353), .ZN(n12352) );
  NOR2_X1 U12363 ( .A1(n12098), .A2(n12096), .ZN(n12353) );
  NAND2_X1 U12364 ( .A1(b_17_), .A2(a_14_), .ZN(n12099) );
  NAND2_X1 U12365 ( .A1(n12096), .A2(n12098), .ZN(n12350) );
  NAND2_X1 U12366 ( .A1(n12354), .A2(n12355), .ZN(n12098) );
  NAND2_X1 U12367 ( .A1(n12232), .A2(n12356), .ZN(n12355) );
  NAND2_X1 U12368 ( .A1(n12229), .A2(n12231), .ZN(n12356) );
  NOR2_X1 U12369 ( .A1(n11951), .A2(n8763), .ZN(n12232) );
  INV_X1 U12370 ( .A(n12357), .ZN(n12354) );
  NOR2_X1 U12371 ( .A1(n12231), .A2(n12229), .ZN(n12357) );
  XNOR2_X1 U12372 ( .A(n12358), .B(n12359), .ZN(n12229) );
  XOR2_X1 U12373 ( .A(n12360), .B(n12361), .Z(n12358) );
  NAND2_X1 U12374 ( .A1(n12362), .A2(n12363), .ZN(n12231) );
  NAND2_X1 U12375 ( .A1(n12226), .A2(n12364), .ZN(n12363) );
  NAND2_X1 U12376 ( .A1(n12228), .A2(n12227), .ZN(n12364) );
  XOR2_X1 U12377 ( .A(n12365), .B(n12366), .Z(n12226) );
  NAND2_X1 U12378 ( .A1(n12367), .A2(n12368), .ZN(n12365) );
  INV_X1 U12379 ( .A(n12369), .ZN(n12362) );
  NOR2_X1 U12380 ( .A1(n12227), .A2(n12228), .ZN(n12369) );
  NOR2_X1 U12381 ( .A1(n11951), .A2(n8768), .ZN(n12228) );
  NAND2_X1 U12382 ( .A1(n12370), .A2(n12371), .ZN(n12227) );
  INV_X1 U12383 ( .A(n12372), .ZN(n12371) );
  NOR2_X1 U12384 ( .A1(n12112), .A2(n12373), .ZN(n12372) );
  NOR2_X1 U12385 ( .A1(n12115), .A2(n12114), .ZN(n12373) );
  XOR2_X1 U12386 ( .A(n12374), .B(n12375), .Z(n12112) );
  XOR2_X1 U12387 ( .A(n12376), .B(n12377), .Z(n12375) );
  NAND2_X1 U12388 ( .A1(b_16_), .A2(a_18_), .ZN(n12377) );
  NAND2_X1 U12389 ( .A1(n12114), .A2(n12115), .ZN(n12370) );
  NAND2_X1 U12390 ( .A1(n12378), .A2(n12379), .ZN(n12115) );
  NAND2_X1 U12391 ( .A1(n12380), .A2(b_17_), .ZN(n12379) );
  NOR2_X1 U12392 ( .A1(n12381), .A2(n10616), .ZN(n12380) );
  NOR2_X1 U12393 ( .A1(n12120), .A2(n12122), .ZN(n12381) );
  NAND2_X1 U12394 ( .A1(n12120), .A2(n12122), .ZN(n12378) );
  NAND2_X1 U12395 ( .A1(n12382), .A2(n12383), .ZN(n12122) );
  NAND2_X1 U12396 ( .A1(n12384), .A2(b_17_), .ZN(n12383) );
  NOR2_X1 U12397 ( .A1(n12385), .A2(n8881), .ZN(n12384) );
  NOR2_X1 U12398 ( .A1(n12223), .A2(n12221), .ZN(n12385) );
  NAND2_X1 U12399 ( .A1(n12223), .A2(n12221), .ZN(n12382) );
  XOR2_X1 U12400 ( .A(n12386), .B(n12387), .Z(n12221) );
  XNOR2_X1 U12401 ( .A(n12388), .B(n12389), .ZN(n12387) );
  NAND2_X1 U12402 ( .A1(b_16_), .A2(a_20_), .ZN(n12389) );
  NOR2_X1 U12403 ( .A1(n12390), .A2(n12391), .ZN(n12223) );
  INV_X1 U12404 ( .A(n12392), .ZN(n12391) );
  NAND2_X1 U12405 ( .A1(n12133), .A2(n12393), .ZN(n12392) );
  NAND2_X1 U12406 ( .A1(n12135), .A2(n12134), .ZN(n12393) );
  XOR2_X1 U12407 ( .A(n12394), .B(n12395), .Z(n12133) );
  XOR2_X1 U12408 ( .A(n12396), .B(n12397), .Z(n12394) );
  NOR2_X1 U12409 ( .A1(n12134), .A2(n12135), .ZN(n12390) );
  NOR2_X1 U12410 ( .A1(n11951), .A2(n10633), .ZN(n12135) );
  NAND2_X1 U12411 ( .A1(n12219), .A2(n12398), .ZN(n12134) );
  NAND2_X1 U12412 ( .A1(n12218), .A2(n12220), .ZN(n12398) );
  NAND2_X1 U12413 ( .A1(n12399), .A2(n12400), .ZN(n12220) );
  NAND2_X1 U12414 ( .A1(b_17_), .A2(a_21_), .ZN(n12400) );
  INV_X1 U12415 ( .A(n12401), .ZN(n12399) );
  XNOR2_X1 U12416 ( .A(n12402), .B(n12403), .ZN(n12218) );
  NAND2_X1 U12417 ( .A1(n12404), .A2(n12405), .ZN(n12402) );
  NAND2_X1 U12418 ( .A1(a_21_), .A2(n12401), .ZN(n12219) );
  NAND2_X1 U12419 ( .A1(n12406), .A2(n12407), .ZN(n12401) );
  NAND2_X1 U12420 ( .A1(n12408), .A2(b_17_), .ZN(n12407) );
  NOR2_X1 U12421 ( .A1(n12409), .A2(n8803), .ZN(n12408) );
  NOR2_X1 U12422 ( .A1(n12145), .A2(n12146), .ZN(n12409) );
  NAND2_X1 U12423 ( .A1(n12145), .A2(n12146), .ZN(n12406) );
  NAND2_X1 U12424 ( .A1(n12410), .A2(n12411), .ZN(n12146) );
  NAND2_X1 U12425 ( .A1(n12412), .A2(b_17_), .ZN(n12411) );
  NOR2_X1 U12426 ( .A1(n12413), .A2(n8812), .ZN(n12412) );
  NOR2_X1 U12427 ( .A1(n12153), .A2(n12154), .ZN(n12413) );
  NAND2_X1 U12428 ( .A1(n12153), .A2(n12154), .ZN(n12410) );
  NAND2_X1 U12429 ( .A1(n12414), .A2(n12415), .ZN(n12154) );
  NAND2_X1 U12430 ( .A1(n12216), .A2(n12416), .ZN(n12415) );
  INV_X1 U12431 ( .A(n12417), .ZN(n12416) );
  NOR2_X1 U12432 ( .A1(n12215), .A2(n12214), .ZN(n12417) );
  NOR2_X1 U12433 ( .A1(n11951), .A2(n9131), .ZN(n12216) );
  NAND2_X1 U12434 ( .A1(n12214), .A2(n12215), .ZN(n12414) );
  NAND2_X1 U12435 ( .A1(n12418), .A2(n12419), .ZN(n12215) );
  NAND2_X1 U12436 ( .A1(n12212), .A2(n12420), .ZN(n12419) );
  NAND2_X1 U12437 ( .A1(n12209), .A2(n12211), .ZN(n12420) );
  NOR2_X1 U12438 ( .A1(n11951), .A2(n8825), .ZN(n12212) );
  INV_X1 U12439 ( .A(n12421), .ZN(n12418) );
  NOR2_X1 U12440 ( .A1(n12211), .A2(n12209), .ZN(n12421) );
  XNOR2_X1 U12441 ( .A(n12422), .B(n12423), .ZN(n12209) );
  XNOR2_X1 U12442 ( .A(n12424), .B(n12425), .ZN(n12423) );
  NAND2_X1 U12443 ( .A1(n12426), .A2(n12427), .ZN(n12211) );
  NAND2_X1 U12444 ( .A1(n12168), .A2(n12428), .ZN(n12427) );
  NAND2_X1 U12445 ( .A1(n12171), .A2(n12170), .ZN(n12428) );
  XNOR2_X1 U12446 ( .A(n12429), .B(n12430), .ZN(n12168) );
  XOR2_X1 U12447 ( .A(n12431), .B(n12432), .Z(n12430) );
  INV_X1 U12448 ( .A(n12433), .ZN(n12426) );
  NOR2_X1 U12449 ( .A1(n12170), .A2(n12171), .ZN(n12433) );
  NOR2_X1 U12450 ( .A1(n11951), .A2(n8830), .ZN(n12171) );
  NAND2_X1 U12451 ( .A1(n12434), .A2(n12435), .ZN(n12170) );
  NAND2_X1 U12452 ( .A1(n12178), .A2(n12436), .ZN(n12435) );
  NAND2_X1 U12453 ( .A1(n12177), .A2(n12175), .ZN(n12436) );
  NOR2_X1 U12454 ( .A1(n11951), .A2(n8839), .ZN(n12178) );
  INV_X1 U12455 ( .A(n12437), .ZN(n12434) );
  NOR2_X1 U12456 ( .A1(n12175), .A2(n12177), .ZN(n12437) );
  NOR2_X1 U12457 ( .A1(n12438), .A2(n12439), .ZN(n12177) );
  INV_X1 U12458 ( .A(n12440), .ZN(n12439) );
  NAND2_X1 U12459 ( .A1(n12207), .A2(n12441), .ZN(n12440) );
  NAND2_X1 U12460 ( .A1(n12208), .A2(n12206), .ZN(n12441) );
  NOR2_X1 U12461 ( .A1(n11951), .A2(n8844), .ZN(n12207) );
  NOR2_X1 U12462 ( .A1(n12206), .A2(n12208), .ZN(n12438) );
  NOR2_X1 U12463 ( .A1(n12442), .A2(n12443), .ZN(n12208) );
  INV_X1 U12464 ( .A(n12444), .ZN(n12443) );
  NAND2_X1 U12465 ( .A1(n12201), .A2(n12445), .ZN(n12444) );
  NAND2_X1 U12466 ( .A1(n12446), .A2(n12203), .ZN(n12445) );
  NOR2_X1 U12467 ( .A1(n11951), .A2(n9161), .ZN(n12201) );
  NOR2_X1 U12468 ( .A1(n12203), .A2(n12446), .ZN(n12442) );
  INV_X1 U12469 ( .A(n12204), .ZN(n12446) );
  NAND2_X1 U12470 ( .A1(n12447), .A2(n12448), .ZN(n12204) );
  NAND2_X1 U12471 ( .A1(b_15_), .A2(n12449), .ZN(n12448) );
  NAND2_X1 U12472 ( .A1(n8358), .A2(n12450), .ZN(n12449) );
  NAND2_X1 U12473 ( .A1(a_31_), .A2(n12199), .ZN(n12450) );
  NAND2_X1 U12474 ( .A1(b_16_), .A2(n12451), .ZN(n12447) );
  NAND2_X1 U12475 ( .A1(n8362), .A2(n12452), .ZN(n12451) );
  NAND2_X1 U12476 ( .A1(a_30_), .A2(n12453), .ZN(n12452) );
  NAND2_X1 U12477 ( .A1(n12454), .A2(b_17_), .ZN(n12203) );
  NOR2_X1 U12478 ( .A1(n9170), .A2(n12199), .ZN(n12454) );
  XOR2_X1 U12479 ( .A(n12455), .B(n12456), .Z(n12206) );
  XOR2_X1 U12480 ( .A(n12457), .B(n12458), .Z(n12456) );
  XOR2_X1 U12481 ( .A(n12459), .B(n12460), .Z(n12175) );
  XNOR2_X1 U12482 ( .A(n12461), .B(n12462), .ZN(n12459) );
  XNOR2_X1 U12483 ( .A(n12463), .B(n12464), .ZN(n12214) );
  XNOR2_X1 U12484 ( .A(n12465), .B(n12466), .ZN(n12464) );
  XOR2_X1 U12485 ( .A(n12467), .B(n12468), .Z(n12153) );
  XOR2_X1 U12486 ( .A(n12469), .B(n12470), .Z(n12467) );
  XNOR2_X1 U12487 ( .A(n12471), .B(n12472), .ZN(n12145) );
  NAND2_X1 U12488 ( .A1(n12473), .A2(n12474), .ZN(n12471) );
  XNOR2_X1 U12489 ( .A(n12475), .B(n12476), .ZN(n12120) );
  XOR2_X1 U12490 ( .A(n12477), .B(n12478), .Z(n12476) );
  NAND2_X1 U12491 ( .A1(b_16_), .A2(a_19_), .ZN(n12478) );
  XNOR2_X1 U12492 ( .A(n12479), .B(n12480), .ZN(n12096) );
  NAND2_X1 U12493 ( .A1(n12481), .A2(n12482), .ZN(n12479) );
  XNOR2_X1 U12494 ( .A(n12483), .B(n12484), .ZN(n12233) );
  XOR2_X1 U12495 ( .A(n12485), .B(n12486), .Z(n12484) );
  NAND2_X1 U12496 ( .A1(b_16_), .A2(a_14_), .ZN(n12486) );
  XNOR2_X1 U12497 ( .A(n12487), .B(n12488), .ZN(n12238) );
  XOR2_X1 U12498 ( .A(n12489), .B(n12490), .Z(n12488) );
  NAND2_X1 U12499 ( .A1(b_16_), .A2(a_13_), .ZN(n12490) );
  XNOR2_X1 U12500 ( .A(n12491), .B(n12492), .ZN(n12080) );
  NAND2_X1 U12501 ( .A1(n12493), .A2(n12494), .ZN(n12491) );
  XNOR2_X1 U12502 ( .A(n12495), .B(n12496), .ZN(n12242) );
  NAND2_X1 U12503 ( .A1(n12497), .A2(n12498), .ZN(n12495) );
  XNOR2_X1 U12504 ( .A(n12499), .B(n12500), .ZN(n12250) );
  NAND2_X1 U12505 ( .A1(n12501), .A2(n12502), .ZN(n12499) );
  XNOR2_X1 U12506 ( .A(n12503), .B(n12504), .ZN(n12009) );
  NAND2_X1 U12507 ( .A1(n12505), .A2(n12506), .ZN(n12503) );
  XOR2_X1 U12508 ( .A(n12507), .B(n12007), .Z(n12261) );
  XNOR2_X1 U12509 ( .A(n12508), .B(n12509), .ZN(n12007) );
  INV_X1 U12510 ( .A(n12006), .ZN(n12507) );
  NAND2_X1 U12511 ( .A1(n8585), .A2(n12510), .ZN(n12260) );
  INV_X1 U12512 ( .A(n12511), .ZN(n12510) );
  NOR2_X1 U12513 ( .A1(n12258), .A2(n12259), .ZN(n12511) );
  NAND2_X1 U12514 ( .A1(n12258), .A2(n12259), .ZN(n8585) );
  XNOR2_X1 U12515 ( .A(n12512), .B(n12513), .ZN(n12259) );
  XOR2_X1 U12516 ( .A(n12514), .B(n12515), .Z(n12513) );
  NAND2_X1 U12517 ( .A1(b_15_), .A2(a_0_), .ZN(n12515) );
  NOR2_X1 U12518 ( .A1(n12516), .A2(n12517), .ZN(n12258) );
  NOR2_X1 U12519 ( .A1(n12006), .A2(n12518), .ZN(n12517) );
  INV_X1 U12520 ( .A(n12519), .ZN(n12518) );
  NAND2_X1 U12521 ( .A1(n12509), .A2(n12508), .ZN(n12519) );
  XNOR2_X1 U12522 ( .A(n12520), .B(n12521), .ZN(n12006) );
  XOR2_X1 U12523 ( .A(n12522), .B(n12523), .Z(n12521) );
  NAND2_X1 U12524 ( .A1(b_15_), .A2(a_1_), .ZN(n12523) );
  NOR2_X1 U12525 ( .A1(n12508), .A2(n12509), .ZN(n12516) );
  NOR2_X1 U12526 ( .A1(n12199), .A2(n8690), .ZN(n12509) );
  NAND2_X1 U12527 ( .A1(n12505), .A2(n12524), .ZN(n12508) );
  NAND2_X1 U12528 ( .A1(n12504), .A2(n12506), .ZN(n12524) );
  NAND2_X1 U12529 ( .A1(n12525), .A2(n12526), .ZN(n12506) );
  INV_X1 U12530 ( .A(n12527), .ZN(n12526) );
  NAND2_X1 U12531 ( .A1(b_16_), .A2(a_1_), .ZN(n12525) );
  XNOR2_X1 U12532 ( .A(n12528), .B(n12529), .ZN(n12504) );
  XOR2_X1 U12533 ( .A(n12530), .B(n12531), .Z(n12529) );
  NAND2_X1 U12534 ( .A1(b_15_), .A2(a_2_), .ZN(n12531) );
  NAND2_X1 U12535 ( .A1(n12527), .A2(a_1_), .ZN(n12505) );
  NOR2_X1 U12536 ( .A1(n12532), .A2(n12533), .ZN(n12527) );
  INV_X1 U12537 ( .A(n12534), .ZN(n12533) );
  NAND2_X1 U12538 ( .A1(n12271), .A2(n12535), .ZN(n12534) );
  NAND2_X1 U12539 ( .A1(n12273), .A2(n12272), .ZN(n12535) );
  XOR2_X1 U12540 ( .A(n12536), .B(n12537), .Z(n12271) );
  XOR2_X1 U12541 ( .A(n12538), .B(n12539), .Z(n12537) );
  NAND2_X1 U12542 ( .A1(b_15_), .A2(a_3_), .ZN(n12539) );
  NOR2_X1 U12543 ( .A1(n12272), .A2(n12273), .ZN(n12532) );
  NOR2_X1 U12544 ( .A1(n12199), .A2(n8497), .ZN(n12273) );
  NAND2_X1 U12545 ( .A1(n12501), .A2(n12540), .ZN(n12272) );
  NAND2_X1 U12546 ( .A1(n12500), .A2(n12502), .ZN(n12540) );
  NAND2_X1 U12547 ( .A1(n12541), .A2(n12542), .ZN(n12502) );
  INV_X1 U12548 ( .A(n12543), .ZN(n12542) );
  NAND2_X1 U12549 ( .A1(b_16_), .A2(a_3_), .ZN(n12541) );
  XNOR2_X1 U12550 ( .A(n12544), .B(n12545), .ZN(n12500) );
  XOR2_X1 U12551 ( .A(n12546), .B(n12547), .Z(n12545) );
  NAND2_X1 U12552 ( .A1(b_15_), .A2(a_4_), .ZN(n12547) );
  NAND2_X1 U12553 ( .A1(n12543), .A2(a_3_), .ZN(n12501) );
  NOR2_X1 U12554 ( .A1(n12548), .A2(n12549), .ZN(n12543) );
  INV_X1 U12555 ( .A(n12550), .ZN(n12549) );
  NAND2_X1 U12556 ( .A1(n12283), .A2(n12551), .ZN(n12550) );
  NAND2_X1 U12557 ( .A1(n12285), .A2(n12284), .ZN(n12551) );
  XOR2_X1 U12558 ( .A(n12552), .B(n12553), .Z(n12283) );
  XOR2_X1 U12559 ( .A(n12554), .B(n12555), .Z(n12553) );
  NAND2_X1 U12560 ( .A1(b_15_), .A2(a_5_), .ZN(n12555) );
  NOR2_X1 U12561 ( .A1(n12284), .A2(n12285), .ZN(n12548) );
  NOR2_X1 U12562 ( .A1(n12199), .A2(n8712), .ZN(n12285) );
  NAND2_X1 U12563 ( .A1(n12292), .A2(n12556), .ZN(n12284) );
  NAND2_X1 U12564 ( .A1(n12291), .A2(n12293), .ZN(n12556) );
  NAND2_X1 U12565 ( .A1(n12557), .A2(n12558), .ZN(n12293) );
  NAND2_X1 U12566 ( .A1(b_16_), .A2(a_5_), .ZN(n12558) );
  INV_X1 U12567 ( .A(n12559), .ZN(n12557) );
  XNOR2_X1 U12568 ( .A(n12560), .B(n12561), .ZN(n12291) );
  XOR2_X1 U12569 ( .A(n12562), .B(n12563), .Z(n12561) );
  NAND2_X1 U12570 ( .A1(b_15_), .A2(a_6_), .ZN(n12563) );
  NAND2_X1 U12571 ( .A1(a_5_), .A2(n12559), .ZN(n12292) );
  NAND2_X1 U12572 ( .A1(n12564), .A2(n12565), .ZN(n12559) );
  NAND2_X1 U12573 ( .A1(n12566), .A2(b_16_), .ZN(n12565) );
  NOR2_X1 U12574 ( .A1(n12567), .A2(n8480), .ZN(n12566) );
  NOR2_X1 U12575 ( .A1(n12299), .A2(n12300), .ZN(n12567) );
  NAND2_X1 U12576 ( .A1(n12299), .A2(n12300), .ZN(n12564) );
  NAND2_X1 U12577 ( .A1(n12497), .A2(n12568), .ZN(n12300) );
  NAND2_X1 U12578 ( .A1(n12496), .A2(n12498), .ZN(n12568) );
  NAND2_X1 U12579 ( .A1(n12569), .A2(n12570), .ZN(n12498) );
  NAND2_X1 U12580 ( .A1(b_16_), .A2(a_7_), .ZN(n12570) );
  INV_X1 U12581 ( .A(n12571), .ZN(n12569) );
  XNOR2_X1 U12582 ( .A(n12572), .B(n12573), .ZN(n12496) );
  NAND2_X1 U12583 ( .A1(n12574), .A2(n12575), .ZN(n12572) );
  NAND2_X1 U12584 ( .A1(a_7_), .A2(n12571), .ZN(n12497) );
  NAND2_X1 U12585 ( .A1(n12576), .A2(n12577), .ZN(n12571) );
  NAND2_X1 U12586 ( .A1(n12578), .A2(b_16_), .ZN(n12577) );
  NOR2_X1 U12587 ( .A1(n12579), .A2(n8731), .ZN(n12578) );
  NOR2_X1 U12588 ( .A1(n12312), .A2(n12310), .ZN(n12579) );
  NAND2_X1 U12589 ( .A1(n12312), .A2(n12310), .ZN(n12576) );
  XOR2_X1 U12590 ( .A(n12580), .B(n12581), .Z(n12310) );
  XOR2_X1 U12591 ( .A(n12582), .B(n12583), .Z(n12580) );
  NOR2_X1 U12592 ( .A1(n8736), .A2(n12453), .ZN(n12583) );
  NOR2_X1 U12593 ( .A1(n12584), .A2(n12585), .ZN(n12312) );
  INV_X1 U12594 ( .A(n12586), .ZN(n12585) );
  NAND2_X1 U12595 ( .A1(n12319), .A2(n12587), .ZN(n12586) );
  NAND2_X1 U12596 ( .A1(n12321), .A2(n12320), .ZN(n12587) );
  XOR2_X1 U12597 ( .A(n12588), .B(n12589), .Z(n12319) );
  NAND2_X1 U12598 ( .A1(n12590), .A2(n12591), .ZN(n12588) );
  NOR2_X1 U12599 ( .A1(n12320), .A2(n12321), .ZN(n12584) );
  NOR2_X1 U12600 ( .A1(n12199), .A2(n8736), .ZN(n12321) );
  NAND2_X1 U12601 ( .A1(n12328), .A2(n12592), .ZN(n12320) );
  NAND2_X1 U12602 ( .A1(n12327), .A2(n12329), .ZN(n12592) );
  NAND2_X1 U12603 ( .A1(n12593), .A2(n12594), .ZN(n12329) );
  NAND2_X1 U12604 ( .A1(b_16_), .A2(a_10_), .ZN(n12594) );
  INV_X1 U12605 ( .A(n12595), .ZN(n12593) );
  XNOR2_X1 U12606 ( .A(n12596), .B(n12597), .ZN(n12327) );
  XOR2_X1 U12607 ( .A(n12598), .B(n12599), .Z(n12597) );
  NAND2_X1 U12608 ( .A1(b_15_), .A2(a_11_), .ZN(n12599) );
  NAND2_X1 U12609 ( .A1(a_10_), .A2(n12595), .ZN(n12328) );
  NAND2_X1 U12610 ( .A1(n12336), .A2(n12600), .ZN(n12595) );
  NAND2_X1 U12611 ( .A1(n12335), .A2(n12337), .ZN(n12600) );
  NAND2_X1 U12612 ( .A1(n12601), .A2(n12602), .ZN(n12337) );
  NAND2_X1 U12613 ( .A1(b_16_), .A2(a_11_), .ZN(n12602) );
  INV_X1 U12614 ( .A(n12603), .ZN(n12601) );
  XNOR2_X1 U12615 ( .A(n12604), .B(n12605), .ZN(n12335) );
  XNOR2_X1 U12616 ( .A(n12606), .B(n12607), .ZN(n12604) );
  NOR2_X1 U12617 ( .A1(n8750), .A2(n12453), .ZN(n12607) );
  NAND2_X1 U12618 ( .A1(a_11_), .A2(n12603), .ZN(n12336) );
  NAND2_X1 U12619 ( .A1(n12493), .A2(n12608), .ZN(n12603) );
  NAND2_X1 U12620 ( .A1(n12492), .A2(n12494), .ZN(n12608) );
  NAND2_X1 U12621 ( .A1(n12609), .A2(n12610), .ZN(n12494) );
  NAND2_X1 U12622 ( .A1(b_16_), .A2(a_12_), .ZN(n12610) );
  INV_X1 U12623 ( .A(n12611), .ZN(n12609) );
  XOR2_X1 U12624 ( .A(n12612), .B(n12613), .Z(n12492) );
  XNOR2_X1 U12625 ( .A(n12614), .B(n12615), .ZN(n12613) );
  NAND2_X1 U12626 ( .A1(a_12_), .A2(n12611), .ZN(n12493) );
  NAND2_X1 U12627 ( .A1(n12616), .A2(n12617), .ZN(n12611) );
  NAND2_X1 U12628 ( .A1(n12618), .A2(b_16_), .ZN(n12617) );
  NOR2_X1 U12629 ( .A1(n12619), .A2(n8443), .ZN(n12618) );
  NOR2_X1 U12630 ( .A1(n12487), .A2(n12489), .ZN(n12619) );
  NAND2_X1 U12631 ( .A1(n12487), .A2(n12489), .ZN(n12616) );
  NAND2_X1 U12632 ( .A1(n12620), .A2(n12621), .ZN(n12489) );
  NAND2_X1 U12633 ( .A1(n12622), .A2(b_16_), .ZN(n12621) );
  NOR2_X1 U12634 ( .A1(n12623), .A2(n8438), .ZN(n12622) );
  NOR2_X1 U12635 ( .A1(n12483), .A2(n12485), .ZN(n12623) );
  NAND2_X1 U12636 ( .A1(n12483), .A2(n12485), .ZN(n12620) );
  NAND2_X1 U12637 ( .A1(n12481), .A2(n12624), .ZN(n12485) );
  NAND2_X1 U12638 ( .A1(n12480), .A2(n12482), .ZN(n12624) );
  NAND2_X1 U12639 ( .A1(n12625), .A2(n12626), .ZN(n12482) );
  NAND2_X1 U12640 ( .A1(b_16_), .A2(a_15_), .ZN(n12626) );
  INV_X1 U12641 ( .A(n12627), .ZN(n12625) );
  XNOR2_X1 U12642 ( .A(n12628), .B(n12629), .ZN(n12480) );
  XOR2_X1 U12643 ( .A(n12630), .B(n12631), .Z(n12628) );
  NAND2_X1 U12644 ( .A1(a_15_), .A2(n12627), .ZN(n12481) );
  NAND2_X1 U12645 ( .A1(n12632), .A2(n12633), .ZN(n12627) );
  NAND2_X1 U12646 ( .A1(n12361), .A2(n12634), .ZN(n12633) );
  INV_X1 U12647 ( .A(n12635), .ZN(n12634) );
  NOR2_X1 U12648 ( .A1(n12360), .A2(n12359), .ZN(n12635) );
  NAND2_X1 U12649 ( .A1(n12359), .A2(n12360), .ZN(n12632) );
  NAND2_X1 U12650 ( .A1(n12367), .A2(n12636), .ZN(n12360) );
  NAND2_X1 U12651 ( .A1(n12366), .A2(n12368), .ZN(n12636) );
  NAND2_X1 U12652 ( .A1(n12637), .A2(n12638), .ZN(n12368) );
  NAND2_X1 U12653 ( .A1(b_16_), .A2(a_17_), .ZN(n12638) );
  INV_X1 U12654 ( .A(n12639), .ZN(n12637) );
  XNOR2_X1 U12655 ( .A(n12640), .B(n12641), .ZN(n12366) );
  XOR2_X1 U12656 ( .A(n12642), .B(n12643), .Z(n12641) );
  NAND2_X1 U12657 ( .A1(b_15_), .A2(a_18_), .ZN(n12643) );
  NAND2_X1 U12658 ( .A1(a_17_), .A2(n12639), .ZN(n12367) );
  NAND2_X1 U12659 ( .A1(n12644), .A2(n12645), .ZN(n12639) );
  NAND2_X1 U12660 ( .A1(n12646), .A2(b_16_), .ZN(n12645) );
  NOR2_X1 U12661 ( .A1(n12647), .A2(n10616), .ZN(n12646) );
  NOR2_X1 U12662 ( .A1(n12374), .A2(n12376), .ZN(n12647) );
  NAND2_X1 U12663 ( .A1(n12374), .A2(n12376), .ZN(n12644) );
  NAND2_X1 U12664 ( .A1(n12648), .A2(n12649), .ZN(n12376) );
  NAND2_X1 U12665 ( .A1(n12650), .A2(b_16_), .ZN(n12649) );
  NOR2_X1 U12666 ( .A1(n12651), .A2(n8881), .ZN(n12650) );
  NOR2_X1 U12667 ( .A1(n12475), .A2(n12477), .ZN(n12651) );
  NAND2_X1 U12668 ( .A1(n12475), .A2(n12477), .ZN(n12648) );
  NAND2_X1 U12669 ( .A1(n12652), .A2(n12653), .ZN(n12477) );
  NAND2_X1 U12670 ( .A1(n12654), .A2(b_16_), .ZN(n12653) );
  NOR2_X1 U12671 ( .A1(n12655), .A2(n10633), .ZN(n12654) );
  NOR2_X1 U12672 ( .A1(n12388), .A2(n12386), .ZN(n12655) );
  NAND2_X1 U12673 ( .A1(n12388), .A2(n12386), .ZN(n12652) );
  XNOR2_X1 U12674 ( .A(n12656), .B(n12657), .ZN(n12386) );
  NAND2_X1 U12675 ( .A1(n12658), .A2(n12659), .ZN(n12656) );
  NOR2_X1 U12676 ( .A1(n12660), .A2(n12661), .ZN(n12388) );
  INV_X1 U12677 ( .A(n12662), .ZN(n12661) );
  NAND2_X1 U12678 ( .A1(n12395), .A2(n12663), .ZN(n12662) );
  NAND2_X1 U12679 ( .A1(n12397), .A2(n12396), .ZN(n12663) );
  XOR2_X1 U12680 ( .A(n12664), .B(n12665), .Z(n12395) );
  XNOR2_X1 U12681 ( .A(n12666), .B(n12667), .ZN(n12665) );
  NOR2_X1 U12682 ( .A1(n12396), .A2(n12397), .ZN(n12660) );
  NOR2_X1 U12683 ( .A1(n12199), .A2(n8798), .ZN(n12397) );
  NAND2_X1 U12684 ( .A1(n12404), .A2(n12668), .ZN(n12396) );
  NAND2_X1 U12685 ( .A1(n12403), .A2(n12405), .ZN(n12668) );
  NAND2_X1 U12686 ( .A1(n12669), .A2(n12670), .ZN(n12405) );
  NAND2_X1 U12687 ( .A1(b_16_), .A2(a_22_), .ZN(n12670) );
  INV_X1 U12688 ( .A(n12671), .ZN(n12669) );
  XOR2_X1 U12689 ( .A(n12672), .B(n12673), .Z(n12403) );
  XOR2_X1 U12690 ( .A(n12674), .B(n12675), .Z(n12672) );
  NAND2_X1 U12691 ( .A1(a_22_), .A2(n12671), .ZN(n12404) );
  NAND2_X1 U12692 ( .A1(n12473), .A2(n12676), .ZN(n12671) );
  NAND2_X1 U12693 ( .A1(n12472), .A2(n12474), .ZN(n12676) );
  NAND2_X1 U12694 ( .A1(n12677), .A2(n12678), .ZN(n12474) );
  NAND2_X1 U12695 ( .A1(b_16_), .A2(a_23_), .ZN(n12678) );
  INV_X1 U12696 ( .A(n12679), .ZN(n12677) );
  XOR2_X1 U12697 ( .A(n12680), .B(n12681), .Z(n12472) );
  XOR2_X1 U12698 ( .A(n12682), .B(n12683), .Z(n12680) );
  NAND2_X1 U12699 ( .A1(a_23_), .A2(n12679), .ZN(n12473) );
  NAND2_X1 U12700 ( .A1(n12684), .A2(n12685), .ZN(n12679) );
  NAND2_X1 U12701 ( .A1(n12470), .A2(n12686), .ZN(n12685) );
  INV_X1 U12702 ( .A(n12687), .ZN(n12686) );
  NOR2_X1 U12703 ( .A1(n12469), .A2(n12468), .ZN(n12687) );
  NOR2_X1 U12704 ( .A1(n12199), .A2(n9131), .ZN(n12470) );
  NAND2_X1 U12705 ( .A1(n12468), .A2(n12469), .ZN(n12684) );
  NAND2_X1 U12706 ( .A1(n12688), .A2(n12689), .ZN(n12469) );
  NAND2_X1 U12707 ( .A1(n12466), .A2(n12690), .ZN(n12689) );
  NAND2_X1 U12708 ( .A1(n12463), .A2(n12465), .ZN(n12690) );
  NOR2_X1 U12709 ( .A1(n12199), .A2(n8825), .ZN(n12466) );
  INV_X1 U12710 ( .A(n12691), .ZN(n12688) );
  NOR2_X1 U12711 ( .A1(n12465), .A2(n12463), .ZN(n12691) );
  XNOR2_X1 U12712 ( .A(n12692), .B(n12693), .ZN(n12463) );
  XNOR2_X1 U12713 ( .A(n12694), .B(n12695), .ZN(n12693) );
  NAND2_X1 U12714 ( .A1(n12696), .A2(n12697), .ZN(n12465) );
  NAND2_X1 U12715 ( .A1(n12422), .A2(n12698), .ZN(n12697) );
  NAND2_X1 U12716 ( .A1(n12425), .A2(n12424), .ZN(n12698) );
  XNOR2_X1 U12717 ( .A(n12699), .B(n12700), .ZN(n12422) );
  XOR2_X1 U12718 ( .A(n12701), .B(n12702), .Z(n12700) );
  INV_X1 U12719 ( .A(n12703), .ZN(n12696) );
  NOR2_X1 U12720 ( .A1(n12424), .A2(n12425), .ZN(n12703) );
  NOR2_X1 U12721 ( .A1(n12199), .A2(n8830), .ZN(n12425) );
  NAND2_X1 U12722 ( .A1(n12704), .A2(n12705), .ZN(n12424) );
  NAND2_X1 U12723 ( .A1(n12432), .A2(n12706), .ZN(n12705) );
  NAND2_X1 U12724 ( .A1(n12431), .A2(n12429), .ZN(n12706) );
  NOR2_X1 U12725 ( .A1(n12199), .A2(n8839), .ZN(n12432) );
  INV_X1 U12726 ( .A(n12707), .ZN(n12704) );
  NOR2_X1 U12727 ( .A1(n12429), .A2(n12431), .ZN(n12707) );
  NOR2_X1 U12728 ( .A1(n12708), .A2(n12709), .ZN(n12431) );
  INV_X1 U12729 ( .A(n12710), .ZN(n12709) );
  NAND2_X1 U12730 ( .A1(n12461), .A2(n12711), .ZN(n12710) );
  NAND2_X1 U12731 ( .A1(n12462), .A2(n12460), .ZN(n12711) );
  NOR2_X1 U12732 ( .A1(n12199), .A2(n8844), .ZN(n12461) );
  NOR2_X1 U12733 ( .A1(n12460), .A2(n12462), .ZN(n12708) );
  NOR2_X1 U12734 ( .A1(n12712), .A2(n12713), .ZN(n12462) );
  INV_X1 U12735 ( .A(n12714), .ZN(n12713) );
  NAND2_X1 U12736 ( .A1(n12455), .A2(n12715), .ZN(n12714) );
  NAND2_X1 U12737 ( .A1(n12716), .A2(n12457), .ZN(n12715) );
  NOR2_X1 U12738 ( .A1(n12199), .A2(n9161), .ZN(n12455) );
  NOR2_X1 U12739 ( .A1(n12457), .A2(n12716), .ZN(n12712) );
  INV_X1 U12740 ( .A(n12458), .ZN(n12716) );
  NAND2_X1 U12741 ( .A1(n12717), .A2(n12718), .ZN(n12458) );
  NAND2_X1 U12742 ( .A1(b_14_), .A2(n12719), .ZN(n12718) );
  NAND2_X1 U12743 ( .A1(n8358), .A2(n12720), .ZN(n12719) );
  NAND2_X1 U12744 ( .A1(a_31_), .A2(n12453), .ZN(n12720) );
  NAND2_X1 U12745 ( .A1(b_15_), .A2(n12721), .ZN(n12717) );
  NAND2_X1 U12746 ( .A1(n8362), .A2(n12722), .ZN(n12721) );
  NAND2_X1 U12747 ( .A1(a_30_), .A2(n12723), .ZN(n12722) );
  NAND2_X1 U12748 ( .A1(n12724), .A2(b_16_), .ZN(n12457) );
  XOR2_X1 U12749 ( .A(n12725), .B(n12726), .Z(n12460) );
  XOR2_X1 U12750 ( .A(n12727), .B(n12728), .Z(n12726) );
  XOR2_X1 U12751 ( .A(n12729), .B(n12730), .Z(n12429) );
  XNOR2_X1 U12752 ( .A(n12731), .B(n12732), .ZN(n12729) );
  XNOR2_X1 U12753 ( .A(n12733), .B(n12734), .ZN(n12468) );
  XNOR2_X1 U12754 ( .A(n12735), .B(n12736), .ZN(n12734) );
  XOR2_X1 U12755 ( .A(n12737), .B(n12738), .Z(n12475) );
  XOR2_X1 U12756 ( .A(n12739), .B(n12740), .Z(n12737) );
  NOR2_X1 U12757 ( .A1(n10633), .A2(n12453), .ZN(n12740) );
  XNOR2_X1 U12758 ( .A(n12741), .B(n12742), .ZN(n12374) );
  XOR2_X1 U12759 ( .A(n12743), .B(n12744), .Z(n12742) );
  NAND2_X1 U12760 ( .A1(b_15_), .A2(a_19_), .ZN(n12744) );
  XNOR2_X1 U12761 ( .A(n12745), .B(n12746), .ZN(n12359) );
  NAND2_X1 U12762 ( .A1(n12747), .A2(n12748), .ZN(n12745) );
  XNOR2_X1 U12763 ( .A(n12749), .B(n12750), .ZN(n12483) );
  XOR2_X1 U12764 ( .A(n12751), .B(n12752), .Z(n12750) );
  XNOR2_X1 U12765 ( .A(n12753), .B(n12754), .ZN(n12487) );
  XOR2_X1 U12766 ( .A(n12755), .B(n12756), .Z(n12753) );
  NOR2_X1 U12767 ( .A1(n8438), .A2(n12453), .ZN(n12756) );
  XOR2_X1 U12768 ( .A(n12757), .B(n12758), .Z(n12299) );
  XOR2_X1 U12769 ( .A(n12759), .B(n12760), .Z(n12757) );
  NOR2_X1 U12770 ( .A1(n8726), .A2(n12453), .ZN(n12760) );
  NAND2_X1 U12771 ( .A1(n12761), .A2(n12762), .ZN(n8584) );
  NAND2_X1 U12772 ( .A1(n12763), .A2(n12764), .ZN(n12761) );
  INV_X1 U12773 ( .A(n12765), .ZN(n12764) );
  XNOR2_X1 U12774 ( .A(n12766), .B(n12767), .ZN(n12763) );
  INV_X1 U12775 ( .A(n12762), .ZN(n8629) );
  NAND2_X1 U12776 ( .A1(n12768), .A2(n12765), .ZN(n12762) );
  NAND2_X1 U12777 ( .A1(n12769), .A2(n12770), .ZN(n12765) );
  NAND2_X1 U12778 ( .A1(n12771), .A2(b_15_), .ZN(n12770) );
  NOR2_X1 U12779 ( .A1(n12772), .A2(n8690), .ZN(n12771) );
  NOR2_X1 U12780 ( .A1(n12512), .A2(n12514), .ZN(n12772) );
  NAND2_X1 U12781 ( .A1(n12512), .A2(n12514), .ZN(n12769) );
  NAND2_X1 U12782 ( .A1(n12773), .A2(n12774), .ZN(n12514) );
  NAND2_X1 U12783 ( .A1(n12775), .A2(b_15_), .ZN(n12774) );
  NOR2_X1 U12784 ( .A1(n12776), .A2(n8502), .ZN(n12775) );
  NOR2_X1 U12785 ( .A1(n12520), .A2(n12522), .ZN(n12776) );
  NAND2_X1 U12786 ( .A1(n12520), .A2(n12522), .ZN(n12773) );
  NAND2_X1 U12787 ( .A1(n12777), .A2(n12778), .ZN(n12522) );
  NAND2_X1 U12788 ( .A1(n12779), .A2(b_15_), .ZN(n12778) );
  NOR2_X1 U12789 ( .A1(n12780), .A2(n8497), .ZN(n12779) );
  NOR2_X1 U12790 ( .A1(n12528), .A2(n12530), .ZN(n12780) );
  NAND2_X1 U12791 ( .A1(n12528), .A2(n12530), .ZN(n12777) );
  NAND2_X1 U12792 ( .A1(n12781), .A2(n12782), .ZN(n12530) );
  NAND2_X1 U12793 ( .A1(n12783), .A2(b_15_), .ZN(n12782) );
  NOR2_X1 U12794 ( .A1(n12784), .A2(n8707), .ZN(n12783) );
  NOR2_X1 U12795 ( .A1(n12536), .A2(n12538), .ZN(n12784) );
  NAND2_X1 U12796 ( .A1(n12536), .A2(n12538), .ZN(n12781) );
  NAND2_X1 U12797 ( .A1(n12785), .A2(n12786), .ZN(n12538) );
  NAND2_X1 U12798 ( .A1(n12787), .A2(b_15_), .ZN(n12786) );
  NOR2_X1 U12799 ( .A1(n12788), .A2(n8712), .ZN(n12787) );
  NOR2_X1 U12800 ( .A1(n12544), .A2(n12546), .ZN(n12788) );
  NAND2_X1 U12801 ( .A1(n12544), .A2(n12546), .ZN(n12785) );
  NAND2_X1 U12802 ( .A1(n12789), .A2(n12790), .ZN(n12546) );
  NAND2_X1 U12803 ( .A1(n12791), .A2(b_15_), .ZN(n12790) );
  NOR2_X1 U12804 ( .A1(n12792), .A2(n8717), .ZN(n12791) );
  NOR2_X1 U12805 ( .A1(n12552), .A2(n12554), .ZN(n12792) );
  NAND2_X1 U12806 ( .A1(n12552), .A2(n12554), .ZN(n12789) );
  NAND2_X1 U12807 ( .A1(n12793), .A2(n12794), .ZN(n12554) );
  NAND2_X1 U12808 ( .A1(n12795), .A2(b_15_), .ZN(n12794) );
  NOR2_X1 U12809 ( .A1(n12796), .A2(n8480), .ZN(n12795) );
  NOR2_X1 U12810 ( .A1(n12560), .A2(n12562), .ZN(n12796) );
  NAND2_X1 U12811 ( .A1(n12560), .A2(n12562), .ZN(n12793) );
  NAND2_X1 U12812 ( .A1(n12797), .A2(n12798), .ZN(n12562) );
  NAND2_X1 U12813 ( .A1(n12799), .A2(b_15_), .ZN(n12798) );
  NOR2_X1 U12814 ( .A1(n12800), .A2(n8726), .ZN(n12799) );
  NOR2_X1 U12815 ( .A1(n12758), .A2(n12759), .ZN(n12800) );
  NAND2_X1 U12816 ( .A1(n12758), .A2(n12759), .ZN(n12797) );
  NAND2_X1 U12817 ( .A1(n12574), .A2(n12801), .ZN(n12759) );
  NAND2_X1 U12818 ( .A1(n12573), .A2(n12575), .ZN(n12801) );
  NAND2_X1 U12819 ( .A1(n12802), .A2(n12803), .ZN(n12575) );
  NAND2_X1 U12820 ( .A1(b_15_), .A2(a_8_), .ZN(n12803) );
  INV_X1 U12821 ( .A(n12804), .ZN(n12802) );
  XNOR2_X1 U12822 ( .A(n12805), .B(n12806), .ZN(n12573) );
  NAND2_X1 U12823 ( .A1(n12807), .A2(n12808), .ZN(n12805) );
  NAND2_X1 U12824 ( .A1(a_8_), .A2(n12804), .ZN(n12574) );
  NAND2_X1 U12825 ( .A1(n12809), .A2(n12810), .ZN(n12804) );
  NAND2_X1 U12826 ( .A1(n12811), .A2(b_15_), .ZN(n12810) );
  NOR2_X1 U12827 ( .A1(n12812), .A2(n8736), .ZN(n12811) );
  NOR2_X1 U12828 ( .A1(n12581), .A2(n12582), .ZN(n12812) );
  NAND2_X1 U12829 ( .A1(n12581), .A2(n12582), .ZN(n12809) );
  NAND2_X1 U12830 ( .A1(n12590), .A2(n12813), .ZN(n12582) );
  NAND2_X1 U12831 ( .A1(n12589), .A2(n12591), .ZN(n12813) );
  NAND2_X1 U12832 ( .A1(n12814), .A2(n12815), .ZN(n12591) );
  NAND2_X1 U12833 ( .A1(b_15_), .A2(a_10_), .ZN(n12815) );
  INV_X1 U12834 ( .A(n12816), .ZN(n12814) );
  XNOR2_X1 U12835 ( .A(n12817), .B(n12818), .ZN(n12589) );
  NAND2_X1 U12836 ( .A1(n12819), .A2(n12820), .ZN(n12817) );
  NAND2_X1 U12837 ( .A1(a_10_), .A2(n12816), .ZN(n12590) );
  NAND2_X1 U12838 ( .A1(n12821), .A2(n12822), .ZN(n12816) );
  NAND2_X1 U12839 ( .A1(n12823), .A2(b_15_), .ZN(n12822) );
  NOR2_X1 U12840 ( .A1(n12824), .A2(n8452), .ZN(n12823) );
  NOR2_X1 U12841 ( .A1(n12596), .A2(n12598), .ZN(n12824) );
  NAND2_X1 U12842 ( .A1(n12596), .A2(n12598), .ZN(n12821) );
  NAND2_X1 U12843 ( .A1(n12825), .A2(n12826), .ZN(n12598) );
  NAND2_X1 U12844 ( .A1(n12827), .A2(b_15_), .ZN(n12826) );
  NOR2_X1 U12845 ( .A1(n12828), .A2(n8750), .ZN(n12827) );
  NOR2_X1 U12846 ( .A1(n12606), .A2(n12605), .ZN(n12828) );
  NAND2_X1 U12847 ( .A1(n12606), .A2(n12605), .ZN(n12825) );
  XNOR2_X1 U12848 ( .A(n12829), .B(n12830), .ZN(n12605) );
  NAND2_X1 U12849 ( .A1(n12831), .A2(n12832), .ZN(n12829) );
  NOR2_X1 U12850 ( .A1(n12833), .A2(n12834), .ZN(n12606) );
  INV_X1 U12851 ( .A(n12835), .ZN(n12834) );
  NAND2_X1 U12852 ( .A1(n12612), .A2(n12836), .ZN(n12835) );
  NAND2_X1 U12853 ( .A1(n12615), .A2(n12614), .ZN(n12836) );
  XNOR2_X1 U12854 ( .A(n12837), .B(n12838), .ZN(n12612) );
  XNOR2_X1 U12855 ( .A(n12839), .B(n12840), .ZN(n12837) );
  NOR2_X1 U12856 ( .A1(n12614), .A2(n12615), .ZN(n12833) );
  NOR2_X1 U12857 ( .A1(n12453), .A2(n8443), .ZN(n12615) );
  NAND2_X1 U12858 ( .A1(n12841), .A2(n12842), .ZN(n12614) );
  NAND2_X1 U12859 ( .A1(n12843), .A2(b_15_), .ZN(n12842) );
  NOR2_X1 U12860 ( .A1(n12844), .A2(n8438), .ZN(n12843) );
  NOR2_X1 U12861 ( .A1(n12845), .A2(n12754), .ZN(n12844) );
  NAND2_X1 U12862 ( .A1(n12845), .A2(n12754), .ZN(n12841) );
  XNOR2_X1 U12863 ( .A(n12846), .B(n12847), .ZN(n12754) );
  NAND2_X1 U12864 ( .A1(n12848), .A2(n12849), .ZN(n12846) );
  INV_X1 U12865 ( .A(n12755), .ZN(n12845) );
  NAND2_X1 U12866 ( .A1(n12850), .A2(n12851), .ZN(n12755) );
  NAND2_X1 U12867 ( .A1(n12749), .A2(n12852), .ZN(n12851) );
  NAND2_X1 U12868 ( .A1(n12853), .A2(n12854), .ZN(n12852) );
  INV_X1 U12869 ( .A(n12751), .ZN(n12853) );
  XOR2_X1 U12870 ( .A(n12855), .B(n12856), .Z(n12749) );
  NAND2_X1 U12871 ( .A1(n12857), .A2(n12858), .ZN(n12855) );
  NAND2_X1 U12872 ( .A1(n12752), .A2(n12751), .ZN(n12850) );
  NAND2_X1 U12873 ( .A1(n12859), .A2(n12860), .ZN(n12751) );
  NAND2_X1 U12874 ( .A1(n12629), .A2(n12861), .ZN(n12860) );
  NAND2_X1 U12875 ( .A1(n12631), .A2(n12630), .ZN(n12861) );
  XOR2_X1 U12876 ( .A(n12862), .B(n12863), .Z(n12629) );
  NAND2_X1 U12877 ( .A1(n12864), .A2(n12865), .ZN(n12862) );
  INV_X1 U12878 ( .A(n12866), .ZN(n12859) );
  NOR2_X1 U12879 ( .A1(n12630), .A2(n12631), .ZN(n12866) );
  NOR2_X1 U12880 ( .A1(n12453), .A2(n8768), .ZN(n12631) );
  NAND2_X1 U12881 ( .A1(n12747), .A2(n12867), .ZN(n12630) );
  NAND2_X1 U12882 ( .A1(n12746), .A2(n12748), .ZN(n12867) );
  NAND2_X1 U12883 ( .A1(n12868), .A2(n12869), .ZN(n12748) );
  NAND2_X1 U12884 ( .A1(b_15_), .A2(a_17_), .ZN(n12869) );
  INV_X1 U12885 ( .A(n12870), .ZN(n12868) );
  XNOR2_X1 U12886 ( .A(n12871), .B(n12872), .ZN(n12746) );
  XOR2_X1 U12887 ( .A(n12873), .B(n12874), .Z(n12872) );
  NAND2_X1 U12888 ( .A1(b_14_), .A2(a_18_), .ZN(n12874) );
  NAND2_X1 U12889 ( .A1(a_17_), .A2(n12870), .ZN(n12747) );
  NAND2_X1 U12890 ( .A1(n12875), .A2(n12876), .ZN(n12870) );
  NAND2_X1 U12891 ( .A1(n12877), .A2(b_15_), .ZN(n12876) );
  NOR2_X1 U12892 ( .A1(n12878), .A2(n10616), .ZN(n12877) );
  NOR2_X1 U12893 ( .A1(n12640), .A2(n12642), .ZN(n12878) );
  NAND2_X1 U12894 ( .A1(n12640), .A2(n12642), .ZN(n12875) );
  NAND2_X1 U12895 ( .A1(n12879), .A2(n12880), .ZN(n12642) );
  NAND2_X1 U12896 ( .A1(n12881), .A2(b_15_), .ZN(n12880) );
  NOR2_X1 U12897 ( .A1(n12882), .A2(n8881), .ZN(n12881) );
  NOR2_X1 U12898 ( .A1(n12741), .A2(n12743), .ZN(n12882) );
  NAND2_X1 U12899 ( .A1(n12741), .A2(n12743), .ZN(n12879) );
  NAND2_X1 U12900 ( .A1(n12883), .A2(n12884), .ZN(n12743) );
  NAND2_X1 U12901 ( .A1(n12885), .A2(b_15_), .ZN(n12884) );
  NOR2_X1 U12902 ( .A1(n12886), .A2(n10633), .ZN(n12885) );
  NOR2_X1 U12903 ( .A1(n12738), .A2(n12739), .ZN(n12886) );
  NAND2_X1 U12904 ( .A1(n12738), .A2(n12739), .ZN(n12883) );
  NAND2_X1 U12905 ( .A1(n12658), .A2(n12887), .ZN(n12739) );
  NAND2_X1 U12906 ( .A1(n12657), .A2(n12659), .ZN(n12887) );
  NAND2_X1 U12907 ( .A1(n12888), .A2(n12889), .ZN(n12659) );
  NAND2_X1 U12908 ( .A1(b_15_), .A2(a_21_), .ZN(n12889) );
  INV_X1 U12909 ( .A(n12890), .ZN(n12888) );
  XOR2_X1 U12910 ( .A(n12891), .B(n12892), .Z(n12657) );
  XOR2_X1 U12911 ( .A(n12893), .B(n12894), .Z(n12891) );
  NAND2_X1 U12912 ( .A1(a_21_), .A2(n12890), .ZN(n12658) );
  NAND2_X1 U12913 ( .A1(n12895), .A2(n12896), .ZN(n12890) );
  NAND2_X1 U12914 ( .A1(n12667), .A2(n12897), .ZN(n12896) );
  INV_X1 U12915 ( .A(n12898), .ZN(n12897) );
  NOR2_X1 U12916 ( .A1(n12666), .A2(n12664), .ZN(n12898) );
  NOR2_X1 U12917 ( .A1(n12453), .A2(n8803), .ZN(n12667) );
  NAND2_X1 U12918 ( .A1(n12664), .A2(n12666), .ZN(n12895) );
  NAND2_X1 U12919 ( .A1(n12899), .A2(n12900), .ZN(n12666) );
  NAND2_X1 U12920 ( .A1(n12675), .A2(n12901), .ZN(n12900) );
  INV_X1 U12921 ( .A(n12902), .ZN(n12901) );
  NOR2_X1 U12922 ( .A1(n12674), .A2(n12673), .ZN(n12902) );
  NOR2_X1 U12923 ( .A1(n12453), .A2(n8812), .ZN(n12675) );
  NAND2_X1 U12924 ( .A1(n12673), .A2(n12674), .ZN(n12899) );
  NAND2_X1 U12925 ( .A1(n12903), .A2(n12904), .ZN(n12674) );
  NAND2_X1 U12926 ( .A1(n12683), .A2(n12905), .ZN(n12904) );
  INV_X1 U12927 ( .A(n12906), .ZN(n12905) );
  NOR2_X1 U12928 ( .A1(n12682), .A2(n12681), .ZN(n12906) );
  NOR2_X1 U12929 ( .A1(n12453), .A2(n9131), .ZN(n12683) );
  NAND2_X1 U12930 ( .A1(n12681), .A2(n12682), .ZN(n12903) );
  NAND2_X1 U12931 ( .A1(n12907), .A2(n12908), .ZN(n12682) );
  NAND2_X1 U12932 ( .A1(n12736), .A2(n12909), .ZN(n12908) );
  NAND2_X1 U12933 ( .A1(n12733), .A2(n12735), .ZN(n12909) );
  NOR2_X1 U12934 ( .A1(n12453), .A2(n8825), .ZN(n12736) );
  INV_X1 U12935 ( .A(n12910), .ZN(n12907) );
  NOR2_X1 U12936 ( .A1(n12735), .A2(n12733), .ZN(n12910) );
  XNOR2_X1 U12937 ( .A(n12911), .B(n12912), .ZN(n12733) );
  XNOR2_X1 U12938 ( .A(n12913), .B(n12914), .ZN(n12912) );
  NAND2_X1 U12939 ( .A1(n12915), .A2(n12916), .ZN(n12735) );
  NAND2_X1 U12940 ( .A1(n12692), .A2(n12917), .ZN(n12916) );
  NAND2_X1 U12941 ( .A1(n12695), .A2(n12694), .ZN(n12917) );
  XNOR2_X1 U12942 ( .A(n12918), .B(n12919), .ZN(n12692) );
  XOR2_X1 U12943 ( .A(n12920), .B(n12921), .Z(n12919) );
  INV_X1 U12944 ( .A(n12922), .ZN(n12915) );
  NOR2_X1 U12945 ( .A1(n12694), .A2(n12695), .ZN(n12922) );
  NOR2_X1 U12946 ( .A1(n12453), .A2(n8830), .ZN(n12695) );
  NAND2_X1 U12947 ( .A1(n12923), .A2(n12924), .ZN(n12694) );
  NAND2_X1 U12948 ( .A1(n12702), .A2(n12925), .ZN(n12924) );
  NAND2_X1 U12949 ( .A1(n12701), .A2(n12699), .ZN(n12925) );
  NOR2_X1 U12950 ( .A1(n12453), .A2(n8839), .ZN(n12702) );
  INV_X1 U12951 ( .A(n12926), .ZN(n12923) );
  NOR2_X1 U12952 ( .A1(n12699), .A2(n12701), .ZN(n12926) );
  NOR2_X1 U12953 ( .A1(n12927), .A2(n12928), .ZN(n12701) );
  INV_X1 U12954 ( .A(n12929), .ZN(n12928) );
  NAND2_X1 U12955 ( .A1(n12731), .A2(n12930), .ZN(n12929) );
  NAND2_X1 U12956 ( .A1(n12732), .A2(n12730), .ZN(n12930) );
  NOR2_X1 U12957 ( .A1(n12453), .A2(n8844), .ZN(n12731) );
  NOR2_X1 U12958 ( .A1(n12730), .A2(n12732), .ZN(n12927) );
  NOR2_X1 U12959 ( .A1(n12931), .A2(n12932), .ZN(n12732) );
  INV_X1 U12960 ( .A(n12933), .ZN(n12932) );
  NAND2_X1 U12961 ( .A1(n12725), .A2(n12934), .ZN(n12933) );
  NAND2_X1 U12962 ( .A1(n12935), .A2(n12727), .ZN(n12934) );
  NOR2_X1 U12963 ( .A1(n12453), .A2(n9161), .ZN(n12725) );
  NOR2_X1 U12964 ( .A1(n12727), .A2(n12935), .ZN(n12931) );
  INV_X1 U12965 ( .A(n12728), .ZN(n12935) );
  NAND2_X1 U12966 ( .A1(n12936), .A2(n12937), .ZN(n12728) );
  NAND2_X1 U12967 ( .A1(b_13_), .A2(n12938), .ZN(n12937) );
  NAND2_X1 U12968 ( .A1(n8358), .A2(n12939), .ZN(n12938) );
  NAND2_X1 U12969 ( .A1(a_31_), .A2(n12723), .ZN(n12939) );
  NAND2_X1 U12970 ( .A1(b_14_), .A2(n12940), .ZN(n12936) );
  NAND2_X1 U12971 ( .A1(n8362), .A2(n12941), .ZN(n12940) );
  NAND2_X1 U12972 ( .A1(a_30_), .A2(n12942), .ZN(n12941) );
  NAND2_X1 U12973 ( .A1(n12724), .A2(b_14_), .ZN(n12727) );
  NOR2_X1 U12974 ( .A1(n9170), .A2(n12453), .ZN(n12724) );
  XOR2_X1 U12975 ( .A(n12943), .B(n12944), .Z(n12730) );
  XOR2_X1 U12976 ( .A(n12945), .B(n12946), .Z(n12944) );
  XOR2_X1 U12977 ( .A(n12947), .B(n12948), .Z(n12699) );
  XNOR2_X1 U12978 ( .A(n12949), .B(n12950), .ZN(n12947) );
  XNOR2_X1 U12979 ( .A(n12951), .B(n12952), .ZN(n12681) );
  XNOR2_X1 U12980 ( .A(n12953), .B(n12954), .ZN(n12952) );
  XOR2_X1 U12981 ( .A(n12955), .B(n12956), .Z(n12673) );
  XOR2_X1 U12982 ( .A(n12957), .B(n12958), .Z(n12955) );
  XOR2_X1 U12983 ( .A(n12959), .B(n12960), .Z(n12664) );
  XOR2_X1 U12984 ( .A(n12961), .B(n12962), .Z(n12959) );
  XNOR2_X1 U12985 ( .A(n12963), .B(n12964), .ZN(n12738) );
  NAND2_X1 U12986 ( .A1(n12965), .A2(n12966), .ZN(n12963) );
  XNOR2_X1 U12987 ( .A(n12967), .B(n12968), .ZN(n12741) );
  XOR2_X1 U12988 ( .A(n12969), .B(n12970), .Z(n12968) );
  NAND2_X1 U12989 ( .A1(b_14_), .A2(a_20_), .ZN(n12970) );
  XNOR2_X1 U12990 ( .A(n12971), .B(n12972), .ZN(n12640) );
  XOR2_X1 U12991 ( .A(n12973), .B(n12974), .Z(n12972) );
  NAND2_X1 U12992 ( .A1(b_14_), .A2(a_19_), .ZN(n12974) );
  XOR2_X1 U12993 ( .A(n12975), .B(n12976), .Z(n12596) );
  XNOR2_X1 U12994 ( .A(n12977), .B(n12978), .ZN(n12976) );
  XOR2_X1 U12995 ( .A(n12979), .B(n12980), .Z(n12581) );
  XNOR2_X1 U12996 ( .A(n12981), .B(n12982), .ZN(n12980) );
  XOR2_X1 U12997 ( .A(n12983), .B(n12984), .Z(n12758) );
  XNOR2_X1 U12998 ( .A(n12985), .B(n12986), .ZN(n12984) );
  XNOR2_X1 U12999 ( .A(n12987), .B(n12988), .ZN(n12560) );
  NAND2_X1 U13000 ( .A1(n12989), .A2(n12990), .ZN(n12987) );
  XNOR2_X1 U13001 ( .A(n12991), .B(n12992), .ZN(n12552) );
  XOR2_X1 U13002 ( .A(n12993), .B(n12994), .Z(n12992) );
  NAND2_X1 U13003 ( .A1(b_14_), .A2(a_6_), .ZN(n12994) );
  XNOR2_X1 U13004 ( .A(n12995), .B(n12996), .ZN(n12544) );
  NAND2_X1 U13005 ( .A1(n12997), .A2(n12998), .ZN(n12995) );
  XNOR2_X1 U13006 ( .A(n12999), .B(n13000), .ZN(n12536) );
  XOR2_X1 U13007 ( .A(n13001), .B(n13002), .Z(n12999) );
  XNOR2_X1 U13008 ( .A(n13003), .B(n13004), .ZN(n12528) );
  NAND2_X1 U13009 ( .A1(n13005), .A2(n13006), .ZN(n13003) );
  XOR2_X1 U13010 ( .A(n13007), .B(n13008), .Z(n12520) );
  XNOR2_X1 U13011 ( .A(n13009), .B(n13010), .ZN(n13008) );
  XNOR2_X1 U13012 ( .A(n13011), .B(n13012), .ZN(n12512) );
  NAND2_X1 U13013 ( .A1(n13013), .A2(n13014), .ZN(n13011) );
  XOR2_X1 U13014 ( .A(n12766), .B(n12767), .Z(n12768) );
  XNOR2_X1 U13015 ( .A(n13015), .B(n13016), .ZN(n12767) );
  XNOR2_X1 U13016 ( .A(n13017), .B(n13018), .ZN(n8586) );
  NAND2_X1 U13017 ( .A1(n8594), .A2(n8593), .ZN(n8592) );
  NOR2_X1 U13018 ( .A1(n13019), .A2(n8626), .ZN(n8593) );
  NOR2_X1 U13019 ( .A1(n13020), .A2(n13021), .ZN(n13019) );
  NOR2_X1 U13020 ( .A1(n13017), .A2(n13018), .ZN(n8594) );
  XOR2_X1 U13021 ( .A(n13022), .B(n13023), .Z(n13018) );
  XOR2_X1 U13022 ( .A(n13024), .B(n13025), .Z(n13023) );
  NAND2_X1 U13023 ( .A1(b_13_), .A2(a_0_), .ZN(n13025) );
  NAND2_X1 U13024 ( .A1(n13026), .A2(n13027), .ZN(n13017) );
  NAND2_X1 U13025 ( .A1(n12766), .A2(n13028), .ZN(n13027) );
  NAND2_X1 U13026 ( .A1(n13016), .A2(n13015), .ZN(n13028) );
  XOR2_X1 U13027 ( .A(n13029), .B(n13030), .Z(n12766) );
  XOR2_X1 U13028 ( .A(n13031), .B(n13032), .Z(n13030) );
  NAND2_X1 U13029 ( .A1(b_13_), .A2(a_1_), .ZN(n13032) );
  INV_X1 U13030 ( .A(n13033), .ZN(n13026) );
  NOR2_X1 U13031 ( .A1(n13015), .A2(n13016), .ZN(n13033) );
  NOR2_X1 U13032 ( .A1(n12723), .A2(n8690), .ZN(n13016) );
  NAND2_X1 U13033 ( .A1(n13013), .A2(n13034), .ZN(n13015) );
  NAND2_X1 U13034 ( .A1(n13012), .A2(n13014), .ZN(n13034) );
  NAND2_X1 U13035 ( .A1(n13035), .A2(n13036), .ZN(n13014) );
  INV_X1 U13036 ( .A(n13037), .ZN(n13036) );
  NAND2_X1 U13037 ( .A1(b_14_), .A2(a_1_), .ZN(n13035) );
  XNOR2_X1 U13038 ( .A(n13038), .B(n13039), .ZN(n13012) );
  XOR2_X1 U13039 ( .A(n13040), .B(n13041), .Z(n13039) );
  NAND2_X1 U13040 ( .A1(b_13_), .A2(a_2_), .ZN(n13041) );
  NAND2_X1 U13041 ( .A1(n13037), .A2(a_1_), .ZN(n13013) );
  NOR2_X1 U13042 ( .A1(n13042), .A2(n13043), .ZN(n13037) );
  INV_X1 U13043 ( .A(n13044), .ZN(n13043) );
  NAND2_X1 U13044 ( .A1(n13007), .A2(n13045), .ZN(n13044) );
  NAND2_X1 U13045 ( .A1(n13010), .A2(n13009), .ZN(n13045) );
  XOR2_X1 U13046 ( .A(n13046), .B(n13047), .Z(n13007) );
  XOR2_X1 U13047 ( .A(n13048), .B(n13049), .Z(n13047) );
  NAND2_X1 U13048 ( .A1(b_13_), .A2(a_3_), .ZN(n13049) );
  NOR2_X1 U13049 ( .A1(n13009), .A2(n13010), .ZN(n13042) );
  NOR2_X1 U13050 ( .A1(n12723), .A2(n8497), .ZN(n13010) );
  NAND2_X1 U13051 ( .A1(n13005), .A2(n13050), .ZN(n13009) );
  NAND2_X1 U13052 ( .A1(n13004), .A2(n13006), .ZN(n13050) );
  NAND2_X1 U13053 ( .A1(n13051), .A2(n13052), .ZN(n13006) );
  INV_X1 U13054 ( .A(n13053), .ZN(n13052) );
  NAND2_X1 U13055 ( .A1(b_14_), .A2(a_3_), .ZN(n13051) );
  XNOR2_X1 U13056 ( .A(n13054), .B(n13055), .ZN(n13004) );
  XOR2_X1 U13057 ( .A(n13056), .B(n13057), .Z(n13055) );
  NAND2_X1 U13058 ( .A1(b_13_), .A2(a_4_), .ZN(n13057) );
  NAND2_X1 U13059 ( .A1(n13053), .A2(a_3_), .ZN(n13005) );
  NOR2_X1 U13060 ( .A1(n13058), .A2(n13059), .ZN(n13053) );
  INV_X1 U13061 ( .A(n13060), .ZN(n13059) );
  NAND2_X1 U13062 ( .A1(n13000), .A2(n13061), .ZN(n13060) );
  NAND2_X1 U13063 ( .A1(n13002), .A2(n13001), .ZN(n13061) );
  XOR2_X1 U13064 ( .A(n13062), .B(n13063), .Z(n13000) );
  XOR2_X1 U13065 ( .A(n13064), .B(n13065), .Z(n13063) );
  NAND2_X1 U13066 ( .A1(b_13_), .A2(a_5_), .ZN(n13065) );
  NOR2_X1 U13067 ( .A1(n13001), .A2(n13002), .ZN(n13058) );
  NOR2_X1 U13068 ( .A1(n12723), .A2(n8712), .ZN(n13002) );
  NAND2_X1 U13069 ( .A1(n12997), .A2(n13066), .ZN(n13001) );
  NAND2_X1 U13070 ( .A1(n12996), .A2(n12998), .ZN(n13066) );
  NAND2_X1 U13071 ( .A1(n13067), .A2(n13068), .ZN(n12998) );
  NAND2_X1 U13072 ( .A1(b_14_), .A2(a_5_), .ZN(n13068) );
  INV_X1 U13073 ( .A(n13069), .ZN(n13067) );
  XNOR2_X1 U13074 ( .A(n13070), .B(n13071), .ZN(n12996) );
  XOR2_X1 U13075 ( .A(n13072), .B(n13073), .Z(n13071) );
  NAND2_X1 U13076 ( .A1(b_13_), .A2(a_6_), .ZN(n13073) );
  NAND2_X1 U13077 ( .A1(a_5_), .A2(n13069), .ZN(n12997) );
  NAND2_X1 U13078 ( .A1(n13074), .A2(n13075), .ZN(n13069) );
  NAND2_X1 U13079 ( .A1(n13076), .A2(b_14_), .ZN(n13075) );
  NOR2_X1 U13080 ( .A1(n13077), .A2(n8480), .ZN(n13076) );
  NOR2_X1 U13081 ( .A1(n12993), .A2(n12991), .ZN(n13077) );
  NAND2_X1 U13082 ( .A1(n12991), .A2(n12993), .ZN(n13074) );
  NAND2_X1 U13083 ( .A1(n12989), .A2(n13078), .ZN(n12993) );
  NAND2_X1 U13084 ( .A1(n12988), .A2(n12990), .ZN(n13078) );
  NAND2_X1 U13085 ( .A1(n13079), .A2(n13080), .ZN(n12990) );
  INV_X1 U13086 ( .A(n13081), .ZN(n13080) );
  NAND2_X1 U13087 ( .A1(b_14_), .A2(a_7_), .ZN(n13079) );
  XNOR2_X1 U13088 ( .A(n13082), .B(n13083), .ZN(n12988) );
  XOR2_X1 U13089 ( .A(n13084), .B(n13085), .Z(n13082) );
  NAND2_X1 U13090 ( .A1(n13081), .A2(a_7_), .ZN(n12989) );
  NOR2_X1 U13091 ( .A1(n13086), .A2(n13087), .ZN(n13081) );
  INV_X1 U13092 ( .A(n13088), .ZN(n13087) );
  NAND2_X1 U13093 ( .A1(n12983), .A2(n13089), .ZN(n13088) );
  NAND2_X1 U13094 ( .A1(n12986), .A2(n12985), .ZN(n13089) );
  XNOR2_X1 U13095 ( .A(n13090), .B(n13091), .ZN(n12983) );
  XOR2_X1 U13096 ( .A(n13092), .B(n13093), .Z(n13090) );
  NOR2_X1 U13097 ( .A1(n8736), .A2(n12942), .ZN(n13093) );
  NOR2_X1 U13098 ( .A1(n12985), .A2(n12986), .ZN(n13086) );
  NOR2_X1 U13099 ( .A1(n12723), .A2(n8731), .ZN(n12986) );
  NAND2_X1 U13100 ( .A1(n12807), .A2(n13094), .ZN(n12985) );
  NAND2_X1 U13101 ( .A1(n12806), .A2(n12808), .ZN(n13094) );
  NAND2_X1 U13102 ( .A1(n13095), .A2(n13096), .ZN(n12808) );
  INV_X1 U13103 ( .A(n13097), .ZN(n13096) );
  NAND2_X1 U13104 ( .A1(b_14_), .A2(a_9_), .ZN(n13095) );
  XOR2_X1 U13105 ( .A(n13098), .B(n13099), .Z(n12806) );
  XOR2_X1 U13106 ( .A(n13100), .B(n13101), .Z(n13098) );
  NOR2_X1 U13107 ( .A1(n8741), .A2(n12942), .ZN(n13101) );
  NAND2_X1 U13108 ( .A1(n13097), .A2(a_9_), .ZN(n12807) );
  NOR2_X1 U13109 ( .A1(n13102), .A2(n13103), .ZN(n13097) );
  INV_X1 U13110 ( .A(n13104), .ZN(n13103) );
  NAND2_X1 U13111 ( .A1(n12979), .A2(n13105), .ZN(n13104) );
  NAND2_X1 U13112 ( .A1(n12982), .A2(n12981), .ZN(n13105) );
  XNOR2_X1 U13113 ( .A(n13106), .B(n13107), .ZN(n12979) );
  XOR2_X1 U13114 ( .A(n13108), .B(n13109), .Z(n13106) );
  NOR2_X1 U13115 ( .A1(n8452), .A2(n12942), .ZN(n13109) );
  NOR2_X1 U13116 ( .A1(n12981), .A2(n12982), .ZN(n13102) );
  NOR2_X1 U13117 ( .A1(n12723), .A2(n8741), .ZN(n12982) );
  NAND2_X1 U13118 ( .A1(n12819), .A2(n13110), .ZN(n12981) );
  NAND2_X1 U13119 ( .A1(n12818), .A2(n12820), .ZN(n13110) );
  NAND2_X1 U13120 ( .A1(n13111), .A2(n13112), .ZN(n12820) );
  INV_X1 U13121 ( .A(n13113), .ZN(n13112) );
  NAND2_X1 U13122 ( .A1(b_14_), .A2(a_11_), .ZN(n13111) );
  XOR2_X1 U13123 ( .A(n13114), .B(n13115), .Z(n12818) );
  XNOR2_X1 U13124 ( .A(n13116), .B(n13117), .ZN(n13114) );
  NAND2_X1 U13125 ( .A1(b_13_), .A2(a_12_), .ZN(n13116) );
  NAND2_X1 U13126 ( .A1(n13113), .A2(a_11_), .ZN(n12819) );
  NOR2_X1 U13127 ( .A1(n13118), .A2(n13119), .ZN(n13113) );
  INV_X1 U13128 ( .A(n13120), .ZN(n13119) );
  NAND2_X1 U13129 ( .A1(n12975), .A2(n13121), .ZN(n13120) );
  NAND2_X1 U13130 ( .A1(n12978), .A2(n12977), .ZN(n13121) );
  XNOR2_X1 U13131 ( .A(n13122), .B(n13123), .ZN(n12975) );
  XOR2_X1 U13132 ( .A(n13124), .B(n13125), .Z(n13123) );
  NOR2_X1 U13133 ( .A1(n12977), .A2(n12978), .ZN(n13118) );
  NOR2_X1 U13134 ( .A1(n12723), .A2(n8750), .ZN(n12978) );
  NAND2_X1 U13135 ( .A1(n12831), .A2(n13126), .ZN(n12977) );
  NAND2_X1 U13136 ( .A1(n12830), .A2(n12832), .ZN(n13126) );
  NAND2_X1 U13137 ( .A1(n13127), .A2(n13128), .ZN(n12832) );
  NAND2_X1 U13138 ( .A1(b_14_), .A2(a_13_), .ZN(n13127) );
  XNOR2_X1 U13139 ( .A(n13129), .B(n13130), .ZN(n12830) );
  XOR2_X1 U13140 ( .A(n13131), .B(n13132), .Z(n13130) );
  NAND2_X1 U13141 ( .A1(b_13_), .A2(a_14_), .ZN(n13132) );
  NAND2_X1 U13142 ( .A1(n13133), .A2(a_13_), .ZN(n12831) );
  INV_X1 U13143 ( .A(n13128), .ZN(n13133) );
  NAND2_X1 U13144 ( .A1(n13134), .A2(n13135), .ZN(n13128) );
  NAND2_X1 U13145 ( .A1(n13136), .A2(n12840), .ZN(n13135) );
  NAND2_X1 U13146 ( .A1(n12838), .A2(n12839), .ZN(n13136) );
  INV_X1 U13147 ( .A(n13137), .ZN(n13134) );
  NOR2_X1 U13148 ( .A1(n12839), .A2(n12838), .ZN(n13137) );
  XNOR2_X1 U13149 ( .A(n13138), .B(n13139), .ZN(n12838) );
  XNOR2_X1 U13150 ( .A(n13140), .B(n13141), .ZN(n13138) );
  NOR2_X1 U13151 ( .A1(n8763), .A2(n12942), .ZN(n13141) );
  NAND2_X1 U13152 ( .A1(n12848), .A2(n13142), .ZN(n12839) );
  NAND2_X1 U13153 ( .A1(n12847), .A2(n12849), .ZN(n13142) );
  NAND2_X1 U13154 ( .A1(n13143), .A2(n13144), .ZN(n12849) );
  NAND2_X1 U13155 ( .A1(b_14_), .A2(a_15_), .ZN(n13144) );
  INV_X1 U13156 ( .A(n13145), .ZN(n13143) );
  XNOR2_X1 U13157 ( .A(n13146), .B(n13147), .ZN(n12847) );
  XOR2_X1 U13158 ( .A(n13148), .B(n13149), .Z(n13146) );
  NAND2_X1 U13159 ( .A1(a_15_), .A2(n13145), .ZN(n12848) );
  NAND2_X1 U13160 ( .A1(n12857), .A2(n13150), .ZN(n13145) );
  NAND2_X1 U13161 ( .A1(n12856), .A2(n12858), .ZN(n13150) );
  NAND2_X1 U13162 ( .A1(n13151), .A2(n13152), .ZN(n12858) );
  NAND2_X1 U13163 ( .A1(b_14_), .A2(a_16_), .ZN(n13152) );
  INV_X1 U13164 ( .A(n13153), .ZN(n13151) );
  XNOR2_X1 U13165 ( .A(n13154), .B(n13155), .ZN(n12856) );
  NAND2_X1 U13166 ( .A1(n13156), .A2(n13157), .ZN(n13154) );
  NAND2_X1 U13167 ( .A1(a_16_), .A2(n13153), .ZN(n12857) );
  NAND2_X1 U13168 ( .A1(n12864), .A2(n13158), .ZN(n13153) );
  NAND2_X1 U13169 ( .A1(n12863), .A2(n12865), .ZN(n13158) );
  NAND2_X1 U13170 ( .A1(n13159), .A2(n13160), .ZN(n12865) );
  NAND2_X1 U13171 ( .A1(b_14_), .A2(a_17_), .ZN(n13160) );
  INV_X1 U13172 ( .A(n13161), .ZN(n13159) );
  XNOR2_X1 U13173 ( .A(n13162), .B(n13163), .ZN(n12863) );
  XOR2_X1 U13174 ( .A(n13164), .B(n13165), .Z(n13163) );
  NAND2_X1 U13175 ( .A1(b_13_), .A2(a_18_), .ZN(n13165) );
  NAND2_X1 U13176 ( .A1(a_17_), .A2(n13161), .ZN(n12864) );
  NAND2_X1 U13177 ( .A1(n13166), .A2(n13167), .ZN(n13161) );
  NAND2_X1 U13178 ( .A1(n13168), .A2(b_14_), .ZN(n13167) );
  NOR2_X1 U13179 ( .A1(n13169), .A2(n10616), .ZN(n13168) );
  NOR2_X1 U13180 ( .A1(n12873), .A2(n12871), .ZN(n13169) );
  NAND2_X1 U13181 ( .A1(n12871), .A2(n12873), .ZN(n13166) );
  NAND2_X1 U13182 ( .A1(n13170), .A2(n13171), .ZN(n12873) );
  NAND2_X1 U13183 ( .A1(n13172), .A2(b_14_), .ZN(n13171) );
  NOR2_X1 U13184 ( .A1(n13173), .A2(n8881), .ZN(n13172) );
  NOR2_X1 U13185 ( .A1(n12973), .A2(n12971), .ZN(n13173) );
  NAND2_X1 U13186 ( .A1(n12971), .A2(n12973), .ZN(n13170) );
  NAND2_X1 U13187 ( .A1(n13174), .A2(n13175), .ZN(n12973) );
  NAND2_X1 U13188 ( .A1(n13176), .A2(b_14_), .ZN(n13175) );
  NOR2_X1 U13189 ( .A1(n13177), .A2(n10633), .ZN(n13176) );
  NOR2_X1 U13190 ( .A1(n12967), .A2(n12969), .ZN(n13177) );
  NAND2_X1 U13191 ( .A1(n12967), .A2(n12969), .ZN(n13174) );
  NAND2_X1 U13192 ( .A1(n12965), .A2(n13178), .ZN(n12969) );
  NAND2_X1 U13193 ( .A1(n12964), .A2(n12966), .ZN(n13178) );
  NAND2_X1 U13194 ( .A1(n13179), .A2(n13180), .ZN(n12966) );
  NAND2_X1 U13195 ( .A1(b_14_), .A2(a_21_), .ZN(n13180) );
  INV_X1 U13196 ( .A(n13181), .ZN(n13179) );
  XNOR2_X1 U13197 ( .A(n13182), .B(n13183), .ZN(n12964) );
  XNOR2_X1 U13198 ( .A(n13184), .B(n13185), .ZN(n13183) );
  NAND2_X1 U13199 ( .A1(a_21_), .A2(n13181), .ZN(n12965) );
  NAND2_X1 U13200 ( .A1(n13186), .A2(n13187), .ZN(n13181) );
  NAND2_X1 U13201 ( .A1(n12894), .A2(n13188), .ZN(n13187) );
  INV_X1 U13202 ( .A(n13189), .ZN(n13188) );
  NOR2_X1 U13203 ( .A1(n12892), .A2(n12893), .ZN(n13189) );
  NOR2_X1 U13204 ( .A1(n12723), .A2(n8803), .ZN(n12894) );
  NAND2_X1 U13205 ( .A1(n12892), .A2(n12893), .ZN(n13186) );
  NAND2_X1 U13206 ( .A1(n13190), .A2(n13191), .ZN(n12893) );
  NAND2_X1 U13207 ( .A1(n12961), .A2(n13192), .ZN(n13191) );
  INV_X1 U13208 ( .A(n13193), .ZN(n13192) );
  NOR2_X1 U13209 ( .A1(n12962), .A2(n12960), .ZN(n13193) );
  NOR2_X1 U13210 ( .A1(n12723), .A2(n8812), .ZN(n12961) );
  NAND2_X1 U13211 ( .A1(n12960), .A2(n12962), .ZN(n13190) );
  NAND2_X1 U13212 ( .A1(n13194), .A2(n13195), .ZN(n12962) );
  NAND2_X1 U13213 ( .A1(n12958), .A2(n13196), .ZN(n13195) );
  INV_X1 U13214 ( .A(n13197), .ZN(n13196) );
  NOR2_X1 U13215 ( .A1(n12956), .A2(n12957), .ZN(n13197) );
  NOR2_X1 U13216 ( .A1(n12723), .A2(n9131), .ZN(n12958) );
  NAND2_X1 U13217 ( .A1(n12956), .A2(n12957), .ZN(n13194) );
  NAND2_X1 U13218 ( .A1(n13198), .A2(n13199), .ZN(n12957) );
  NAND2_X1 U13219 ( .A1(n12954), .A2(n13200), .ZN(n13199) );
  NAND2_X1 U13220 ( .A1(n12951), .A2(n12953), .ZN(n13200) );
  NOR2_X1 U13221 ( .A1(n12723), .A2(n8825), .ZN(n12954) );
  INV_X1 U13222 ( .A(n13201), .ZN(n13198) );
  NOR2_X1 U13223 ( .A1(n12953), .A2(n12951), .ZN(n13201) );
  XOR2_X1 U13224 ( .A(n13202), .B(n13203), .Z(n12951) );
  XOR2_X1 U13225 ( .A(n13204), .B(n13205), .Z(n13202) );
  NAND2_X1 U13226 ( .A1(n13206), .A2(n13207), .ZN(n12953) );
  NAND2_X1 U13227 ( .A1(n12911), .A2(n13208), .ZN(n13207) );
  NAND2_X1 U13228 ( .A1(n12914), .A2(n12913), .ZN(n13208) );
  XOR2_X1 U13229 ( .A(n13209), .B(n13210), .Z(n12911) );
  XNOR2_X1 U13230 ( .A(n13211), .B(n13212), .ZN(n13209) );
  INV_X1 U13231 ( .A(n13213), .ZN(n13206) );
  NOR2_X1 U13232 ( .A1(n12913), .A2(n12914), .ZN(n13213) );
  NOR2_X1 U13233 ( .A1(n12723), .A2(n8830), .ZN(n12914) );
  NAND2_X1 U13234 ( .A1(n13214), .A2(n13215), .ZN(n12913) );
  NAND2_X1 U13235 ( .A1(n12921), .A2(n13216), .ZN(n13215) );
  NAND2_X1 U13236 ( .A1(n12918), .A2(n12920), .ZN(n13216) );
  NOR2_X1 U13237 ( .A1(n12723), .A2(n8839), .ZN(n12921) );
  INV_X1 U13238 ( .A(n13217), .ZN(n13214) );
  NOR2_X1 U13239 ( .A1(n12918), .A2(n12920), .ZN(n13217) );
  NOR2_X1 U13240 ( .A1(n13218), .A2(n13219), .ZN(n12920) );
  INV_X1 U13241 ( .A(n13220), .ZN(n13219) );
  NAND2_X1 U13242 ( .A1(n12949), .A2(n13221), .ZN(n13220) );
  NAND2_X1 U13243 ( .A1(n12950), .A2(n12948), .ZN(n13221) );
  NOR2_X1 U13244 ( .A1(n12723), .A2(n8844), .ZN(n12949) );
  NOR2_X1 U13245 ( .A1(n12948), .A2(n12950), .ZN(n13218) );
  NOR2_X1 U13246 ( .A1(n13222), .A2(n13223), .ZN(n12950) );
  INV_X1 U13247 ( .A(n13224), .ZN(n13223) );
  NAND2_X1 U13248 ( .A1(n12943), .A2(n13225), .ZN(n13224) );
  NAND2_X1 U13249 ( .A1(n13226), .A2(n12945), .ZN(n13225) );
  NOR2_X1 U13250 ( .A1(n12723), .A2(n9161), .ZN(n12943) );
  NOR2_X1 U13251 ( .A1(n12945), .A2(n13226), .ZN(n13222) );
  INV_X1 U13252 ( .A(n12946), .ZN(n13226) );
  NAND2_X1 U13253 ( .A1(n13227), .A2(n13228), .ZN(n12946) );
  NAND2_X1 U13254 ( .A1(b_12_), .A2(n13229), .ZN(n13228) );
  NAND2_X1 U13255 ( .A1(n8358), .A2(n13230), .ZN(n13229) );
  NAND2_X1 U13256 ( .A1(a_31_), .A2(n12942), .ZN(n13230) );
  NAND2_X1 U13257 ( .A1(b_13_), .A2(n13231), .ZN(n13227) );
  NAND2_X1 U13258 ( .A1(n8362), .A2(n13232), .ZN(n13231) );
  NAND2_X1 U13259 ( .A1(a_30_), .A2(n13233), .ZN(n13232) );
  NAND2_X1 U13260 ( .A1(n13234), .A2(b_14_), .ZN(n12945) );
  XOR2_X1 U13261 ( .A(n13235), .B(n13236), .Z(n12948) );
  XOR2_X1 U13262 ( .A(n13237), .B(n13238), .Z(n13236) );
  XOR2_X1 U13263 ( .A(n13239), .B(n13240), .Z(n12918) );
  XNOR2_X1 U13264 ( .A(n13241), .B(n13242), .ZN(n13239) );
  XNOR2_X1 U13265 ( .A(n13243), .B(n13244), .ZN(n12956) );
  XNOR2_X1 U13266 ( .A(n13245), .B(n13246), .ZN(n13244) );
  XOR2_X1 U13267 ( .A(n13247), .B(n13248), .Z(n12960) );
  XOR2_X1 U13268 ( .A(n13249), .B(n13250), .Z(n13248) );
  XOR2_X1 U13269 ( .A(n13251), .B(n13252), .Z(n12892) );
  XOR2_X1 U13270 ( .A(n13253), .B(n13254), .Z(n13251) );
  XNOR2_X1 U13271 ( .A(n13255), .B(n13256), .ZN(n12967) );
  NAND2_X1 U13272 ( .A1(n13257), .A2(n13258), .ZN(n13255) );
  XOR2_X1 U13273 ( .A(n13259), .B(n13260), .Z(n12971) );
  XOR2_X1 U13274 ( .A(n13261), .B(n13262), .Z(n13259) );
  NOR2_X1 U13275 ( .A1(n10633), .A2(n12942), .ZN(n13262) );
  XNOR2_X1 U13276 ( .A(n13263), .B(n13264), .ZN(n12871) );
  XOR2_X1 U13277 ( .A(n13265), .B(n13266), .Z(n13264) );
  NAND2_X1 U13278 ( .A1(b_13_), .A2(a_19_), .ZN(n13266) );
  XOR2_X1 U13279 ( .A(n13267), .B(n13268), .Z(n12991) );
  XNOR2_X1 U13280 ( .A(n13269), .B(n13270), .ZN(n13268) );
  NAND2_X1 U13281 ( .A1(b_13_), .A2(a_7_), .ZN(n13270) );
  INV_X1 U13282 ( .A(n13271), .ZN(n8626) );
  NAND2_X1 U13283 ( .A1(n13020), .A2(n13021), .ZN(n13271) );
  NAND2_X1 U13284 ( .A1(n13272), .A2(n13273), .ZN(n13021) );
  NAND2_X1 U13285 ( .A1(n13274), .A2(b_13_), .ZN(n13273) );
  NOR2_X1 U13286 ( .A1(n13275), .A2(n8690), .ZN(n13274) );
  NOR2_X1 U13287 ( .A1(n13022), .A2(n13024), .ZN(n13275) );
  NAND2_X1 U13288 ( .A1(n13022), .A2(n13024), .ZN(n13272) );
  NAND2_X1 U13289 ( .A1(n13276), .A2(n13277), .ZN(n13024) );
  NAND2_X1 U13290 ( .A1(n13278), .A2(b_13_), .ZN(n13277) );
  NOR2_X1 U13291 ( .A1(n13279), .A2(n8502), .ZN(n13278) );
  NOR2_X1 U13292 ( .A1(n13029), .A2(n13031), .ZN(n13279) );
  NAND2_X1 U13293 ( .A1(n13029), .A2(n13031), .ZN(n13276) );
  NAND2_X1 U13294 ( .A1(n13280), .A2(n13281), .ZN(n13031) );
  NAND2_X1 U13295 ( .A1(n13282), .A2(b_13_), .ZN(n13281) );
  NOR2_X1 U13296 ( .A1(n13283), .A2(n8497), .ZN(n13282) );
  NOR2_X1 U13297 ( .A1(n13038), .A2(n13040), .ZN(n13283) );
  NAND2_X1 U13298 ( .A1(n13038), .A2(n13040), .ZN(n13280) );
  NAND2_X1 U13299 ( .A1(n13284), .A2(n13285), .ZN(n13040) );
  NAND2_X1 U13300 ( .A1(n13286), .A2(b_13_), .ZN(n13285) );
  NOR2_X1 U13301 ( .A1(n13287), .A2(n8707), .ZN(n13286) );
  NOR2_X1 U13302 ( .A1(n13046), .A2(n13048), .ZN(n13287) );
  NAND2_X1 U13303 ( .A1(n13046), .A2(n13048), .ZN(n13284) );
  NAND2_X1 U13304 ( .A1(n13288), .A2(n13289), .ZN(n13048) );
  NAND2_X1 U13305 ( .A1(n13290), .A2(b_13_), .ZN(n13289) );
  NOR2_X1 U13306 ( .A1(n13291), .A2(n8712), .ZN(n13290) );
  NOR2_X1 U13307 ( .A1(n13054), .A2(n13056), .ZN(n13291) );
  NAND2_X1 U13308 ( .A1(n13054), .A2(n13056), .ZN(n13288) );
  NAND2_X1 U13309 ( .A1(n13292), .A2(n13293), .ZN(n13056) );
  NAND2_X1 U13310 ( .A1(n13294), .A2(b_13_), .ZN(n13293) );
  NOR2_X1 U13311 ( .A1(n13295), .A2(n8717), .ZN(n13294) );
  NOR2_X1 U13312 ( .A1(n13062), .A2(n13064), .ZN(n13295) );
  NAND2_X1 U13313 ( .A1(n13062), .A2(n13064), .ZN(n13292) );
  NAND2_X1 U13314 ( .A1(n13296), .A2(n13297), .ZN(n13064) );
  NAND2_X1 U13315 ( .A1(n13298), .A2(b_13_), .ZN(n13297) );
  NOR2_X1 U13316 ( .A1(n13299), .A2(n8480), .ZN(n13298) );
  NOR2_X1 U13317 ( .A1(n13070), .A2(n13072), .ZN(n13299) );
  NAND2_X1 U13318 ( .A1(n13070), .A2(n13072), .ZN(n13296) );
  NAND2_X1 U13319 ( .A1(n13300), .A2(n13301), .ZN(n13072) );
  NAND2_X1 U13320 ( .A1(n13302), .A2(b_13_), .ZN(n13301) );
  NOR2_X1 U13321 ( .A1(n13303), .A2(n8726), .ZN(n13302) );
  NOR2_X1 U13322 ( .A1(n13269), .A2(n13267), .ZN(n13303) );
  NAND2_X1 U13323 ( .A1(n13269), .A2(n13267), .ZN(n13300) );
  XNOR2_X1 U13324 ( .A(n13304), .B(n13305), .ZN(n13267) );
  NAND2_X1 U13325 ( .A1(n13306), .A2(n13307), .ZN(n13304) );
  NOR2_X1 U13326 ( .A1(n13308), .A2(n13309), .ZN(n13269) );
  INV_X1 U13327 ( .A(n13310), .ZN(n13309) );
  NAND2_X1 U13328 ( .A1(n13083), .A2(n13311), .ZN(n13310) );
  NAND2_X1 U13329 ( .A1(n13085), .A2(n13084), .ZN(n13311) );
  XOR2_X1 U13330 ( .A(n13312), .B(n13313), .Z(n13083) );
  NAND2_X1 U13331 ( .A1(n13314), .A2(n13315), .ZN(n13312) );
  NOR2_X1 U13332 ( .A1(n13084), .A2(n13085), .ZN(n13308) );
  NOR2_X1 U13333 ( .A1(n12942), .A2(n8731), .ZN(n13085) );
  NAND2_X1 U13334 ( .A1(n13316), .A2(n13317), .ZN(n13084) );
  NAND2_X1 U13335 ( .A1(n13318), .A2(b_13_), .ZN(n13317) );
  NOR2_X1 U13336 ( .A1(n13319), .A2(n8736), .ZN(n13318) );
  NOR2_X1 U13337 ( .A1(n13091), .A2(n13092), .ZN(n13319) );
  NAND2_X1 U13338 ( .A1(n13091), .A2(n13092), .ZN(n13316) );
  NAND2_X1 U13339 ( .A1(n13320), .A2(n13321), .ZN(n13092) );
  NAND2_X1 U13340 ( .A1(n13322), .A2(b_13_), .ZN(n13321) );
  NOR2_X1 U13341 ( .A1(n13323), .A2(n8741), .ZN(n13322) );
  NOR2_X1 U13342 ( .A1(n13099), .A2(n13100), .ZN(n13323) );
  NAND2_X1 U13343 ( .A1(n13099), .A2(n13100), .ZN(n13320) );
  NAND2_X1 U13344 ( .A1(n13324), .A2(n13325), .ZN(n13100) );
  NAND2_X1 U13345 ( .A1(n13326), .A2(b_13_), .ZN(n13325) );
  NOR2_X1 U13346 ( .A1(n13327), .A2(n8452), .ZN(n13326) );
  NOR2_X1 U13347 ( .A1(n13107), .A2(n13108), .ZN(n13327) );
  NAND2_X1 U13348 ( .A1(n13107), .A2(n13108), .ZN(n13324) );
  NAND2_X1 U13349 ( .A1(n13328), .A2(n13329), .ZN(n13108) );
  NAND2_X1 U13350 ( .A1(n13330), .A2(b_13_), .ZN(n13329) );
  NOR2_X1 U13351 ( .A1(n13331), .A2(n8750), .ZN(n13330) );
  NOR2_X1 U13352 ( .A1(n13115), .A2(n13117), .ZN(n13331) );
  NAND2_X1 U13353 ( .A1(n13115), .A2(n13117), .ZN(n13328) );
  NAND2_X1 U13354 ( .A1(n13332), .A2(n13333), .ZN(n13117) );
  INV_X1 U13355 ( .A(n13334), .ZN(n13333) );
  NOR2_X1 U13356 ( .A1(n13122), .A2(n13335), .ZN(n13334) );
  NOR2_X1 U13357 ( .A1(n13125), .A2(n13336), .ZN(n13335) );
  XOR2_X1 U13358 ( .A(n13337), .B(n13338), .Z(n13122) );
  NAND2_X1 U13359 ( .A1(n13339), .A2(n13340), .ZN(n13337) );
  NAND2_X1 U13360 ( .A1(n13336), .A2(n13125), .ZN(n13332) );
  NAND2_X1 U13361 ( .A1(n13341), .A2(n13342), .ZN(n13125) );
  NAND2_X1 U13362 ( .A1(n13343), .A2(b_13_), .ZN(n13342) );
  NOR2_X1 U13363 ( .A1(n13344), .A2(n8438), .ZN(n13343) );
  NOR2_X1 U13364 ( .A1(n13129), .A2(n13131), .ZN(n13344) );
  NAND2_X1 U13365 ( .A1(n13129), .A2(n13131), .ZN(n13341) );
  NAND2_X1 U13366 ( .A1(n13345), .A2(n13346), .ZN(n13131) );
  NAND2_X1 U13367 ( .A1(n13347), .A2(b_13_), .ZN(n13346) );
  NOR2_X1 U13368 ( .A1(n13348), .A2(n8763), .ZN(n13347) );
  NOR2_X1 U13369 ( .A1(n13140), .A2(n13139), .ZN(n13348) );
  NAND2_X1 U13370 ( .A1(n13140), .A2(n13139), .ZN(n13345) );
  XNOR2_X1 U13371 ( .A(n13349), .B(n13350), .ZN(n13139) );
  NAND2_X1 U13372 ( .A1(n13351), .A2(n13352), .ZN(n13349) );
  NOR2_X1 U13373 ( .A1(n13353), .A2(n13354), .ZN(n13140) );
  INV_X1 U13374 ( .A(n13355), .ZN(n13354) );
  NAND2_X1 U13375 ( .A1(n13147), .A2(n13356), .ZN(n13355) );
  NAND2_X1 U13376 ( .A1(n13149), .A2(n13148), .ZN(n13356) );
  XNOR2_X1 U13377 ( .A(n13357), .B(n13358), .ZN(n13147) );
  XOR2_X1 U13378 ( .A(n13359), .B(n13360), .Z(n13357) );
  NOR2_X1 U13379 ( .A1(n8772), .A2(n13233), .ZN(n13360) );
  NOR2_X1 U13380 ( .A1(n13148), .A2(n13149), .ZN(n13353) );
  NOR2_X1 U13381 ( .A1(n12942), .A2(n8768), .ZN(n13149) );
  NAND2_X1 U13382 ( .A1(n13156), .A2(n13361), .ZN(n13148) );
  NAND2_X1 U13383 ( .A1(n13155), .A2(n13157), .ZN(n13361) );
  NAND2_X1 U13384 ( .A1(n13362), .A2(n13363), .ZN(n13157) );
  NAND2_X1 U13385 ( .A1(b_13_), .A2(a_17_), .ZN(n13363) );
  INV_X1 U13386 ( .A(n13364), .ZN(n13362) );
  XOR2_X1 U13387 ( .A(n13365), .B(n13366), .Z(n13155) );
  XOR2_X1 U13388 ( .A(n13367), .B(n13368), .Z(n13365) );
  NOR2_X1 U13389 ( .A1(n10616), .A2(n13233), .ZN(n13368) );
  NAND2_X1 U13390 ( .A1(a_17_), .A2(n13364), .ZN(n13156) );
  NAND2_X1 U13391 ( .A1(n13369), .A2(n13370), .ZN(n13364) );
  NAND2_X1 U13392 ( .A1(n13371), .A2(b_13_), .ZN(n13370) );
  NOR2_X1 U13393 ( .A1(n13372), .A2(n10616), .ZN(n13371) );
  NOR2_X1 U13394 ( .A1(n13162), .A2(n13164), .ZN(n13372) );
  NAND2_X1 U13395 ( .A1(n13162), .A2(n13164), .ZN(n13369) );
  NAND2_X1 U13396 ( .A1(n13373), .A2(n13374), .ZN(n13164) );
  NAND2_X1 U13397 ( .A1(n13375), .A2(b_13_), .ZN(n13374) );
  NOR2_X1 U13398 ( .A1(n13376), .A2(n8881), .ZN(n13375) );
  NOR2_X1 U13399 ( .A1(n13263), .A2(n13265), .ZN(n13376) );
  NAND2_X1 U13400 ( .A1(n13263), .A2(n13265), .ZN(n13373) );
  NAND2_X1 U13401 ( .A1(n13377), .A2(n13378), .ZN(n13265) );
  NAND2_X1 U13402 ( .A1(n13379), .A2(b_13_), .ZN(n13378) );
  NOR2_X1 U13403 ( .A1(n13380), .A2(n10633), .ZN(n13379) );
  NOR2_X1 U13404 ( .A1(n13260), .A2(n13261), .ZN(n13380) );
  NAND2_X1 U13405 ( .A1(n13260), .A2(n13261), .ZN(n13377) );
  NAND2_X1 U13406 ( .A1(n13257), .A2(n13381), .ZN(n13261) );
  NAND2_X1 U13407 ( .A1(n13256), .A2(n13258), .ZN(n13381) );
  NAND2_X1 U13408 ( .A1(n13382), .A2(n13383), .ZN(n13258) );
  NAND2_X1 U13409 ( .A1(b_13_), .A2(a_21_), .ZN(n13383) );
  INV_X1 U13410 ( .A(n13384), .ZN(n13382) );
  XNOR2_X1 U13411 ( .A(n13385), .B(n13386), .ZN(n13256) );
  XNOR2_X1 U13412 ( .A(n13387), .B(n13388), .ZN(n13386) );
  NAND2_X1 U13413 ( .A1(a_21_), .A2(n13384), .ZN(n13257) );
  NAND2_X1 U13414 ( .A1(n13389), .A2(n13390), .ZN(n13384) );
  NAND2_X1 U13415 ( .A1(n13185), .A2(n13391), .ZN(n13390) );
  INV_X1 U13416 ( .A(n13392), .ZN(n13391) );
  NOR2_X1 U13417 ( .A1(n13184), .A2(n13182), .ZN(n13392) );
  NOR2_X1 U13418 ( .A1(n12942), .A2(n8803), .ZN(n13185) );
  NAND2_X1 U13419 ( .A1(n13182), .A2(n13184), .ZN(n13389) );
  NAND2_X1 U13420 ( .A1(n13393), .A2(n13394), .ZN(n13184) );
  NAND2_X1 U13421 ( .A1(n13253), .A2(n13395), .ZN(n13394) );
  INV_X1 U13422 ( .A(n13396), .ZN(n13395) );
  NOR2_X1 U13423 ( .A1(n13254), .A2(n13252), .ZN(n13396) );
  NOR2_X1 U13424 ( .A1(n12942), .A2(n8812), .ZN(n13253) );
  NAND2_X1 U13425 ( .A1(n13252), .A2(n13254), .ZN(n13393) );
  NAND2_X1 U13426 ( .A1(n13397), .A2(n13398), .ZN(n13254) );
  NAND2_X1 U13427 ( .A1(n13250), .A2(n13399), .ZN(n13398) );
  NAND2_X1 U13428 ( .A1(n13249), .A2(n13247), .ZN(n13399) );
  NOR2_X1 U13429 ( .A1(n12942), .A2(n9131), .ZN(n13250) );
  INV_X1 U13430 ( .A(n13400), .ZN(n13397) );
  NOR2_X1 U13431 ( .A1(n13247), .A2(n13249), .ZN(n13400) );
  NOR2_X1 U13432 ( .A1(n13401), .A2(n13402), .ZN(n13249) );
  INV_X1 U13433 ( .A(n13403), .ZN(n13402) );
  NAND2_X1 U13434 ( .A1(n13246), .A2(n13404), .ZN(n13403) );
  NAND2_X1 U13435 ( .A1(n13243), .A2(n13245), .ZN(n13404) );
  NOR2_X1 U13436 ( .A1(n12942), .A2(n8825), .ZN(n13246) );
  NOR2_X1 U13437 ( .A1(n13245), .A2(n13243), .ZN(n13401) );
  XOR2_X1 U13438 ( .A(n13405), .B(n13406), .Z(n13243) );
  XOR2_X1 U13439 ( .A(n13407), .B(n13408), .Z(n13405) );
  NAND2_X1 U13440 ( .A1(n13409), .A2(n13410), .ZN(n13245) );
  NAND2_X1 U13441 ( .A1(n13203), .A2(n13411), .ZN(n13410) );
  INV_X1 U13442 ( .A(n13412), .ZN(n13411) );
  NOR2_X1 U13443 ( .A1(n13204), .A2(n13205), .ZN(n13412) );
  XNOR2_X1 U13444 ( .A(n13413), .B(n13414), .ZN(n13203) );
  XNOR2_X1 U13445 ( .A(n13415), .B(n13416), .ZN(n13413) );
  NAND2_X1 U13446 ( .A1(n13205), .A2(n13204), .ZN(n13409) );
  NAND2_X1 U13447 ( .A1(b_13_), .A2(a_26_), .ZN(n13204) );
  NOR2_X1 U13448 ( .A1(n13417), .A2(n13418), .ZN(n13205) );
  INV_X1 U13449 ( .A(n13419), .ZN(n13418) );
  NAND2_X1 U13450 ( .A1(n13212), .A2(n13420), .ZN(n13419) );
  NAND2_X1 U13451 ( .A1(n13211), .A2(n13210), .ZN(n13420) );
  NOR2_X1 U13452 ( .A1(n12942), .A2(n8839), .ZN(n13212) );
  NOR2_X1 U13453 ( .A1(n13210), .A2(n13211), .ZN(n13417) );
  NOR2_X1 U13454 ( .A1(n13421), .A2(n13422), .ZN(n13211) );
  INV_X1 U13455 ( .A(n13423), .ZN(n13422) );
  NAND2_X1 U13456 ( .A1(n13241), .A2(n13424), .ZN(n13423) );
  NAND2_X1 U13457 ( .A1(n13242), .A2(n13240), .ZN(n13424) );
  NOR2_X1 U13458 ( .A1(n12942), .A2(n8844), .ZN(n13241) );
  NOR2_X1 U13459 ( .A1(n13240), .A2(n13242), .ZN(n13421) );
  NOR2_X1 U13460 ( .A1(n13425), .A2(n13426), .ZN(n13242) );
  INV_X1 U13461 ( .A(n13427), .ZN(n13426) );
  NAND2_X1 U13462 ( .A1(n13235), .A2(n13428), .ZN(n13427) );
  NAND2_X1 U13463 ( .A1(n13429), .A2(n13237), .ZN(n13428) );
  NOR2_X1 U13464 ( .A1(n12942), .A2(n9161), .ZN(n13235) );
  NOR2_X1 U13465 ( .A1(n13237), .A2(n13429), .ZN(n13425) );
  INV_X1 U13466 ( .A(n13238), .ZN(n13429) );
  NAND2_X1 U13467 ( .A1(n13430), .A2(n13431), .ZN(n13238) );
  NAND2_X1 U13468 ( .A1(b_11_), .A2(n13432), .ZN(n13431) );
  NAND2_X1 U13469 ( .A1(n8358), .A2(n13433), .ZN(n13432) );
  NAND2_X1 U13470 ( .A1(a_31_), .A2(n13233), .ZN(n13433) );
  NAND2_X1 U13471 ( .A1(b_12_), .A2(n13434), .ZN(n13430) );
  NAND2_X1 U13472 ( .A1(n8362), .A2(n13435), .ZN(n13434) );
  NAND2_X1 U13473 ( .A1(a_30_), .A2(n13436), .ZN(n13435) );
  NAND2_X1 U13474 ( .A1(n13234), .A2(b_12_), .ZN(n13237) );
  NOR2_X1 U13475 ( .A1(n9170), .A2(n12942), .ZN(n13234) );
  XOR2_X1 U13476 ( .A(n13437), .B(n13438), .Z(n13240) );
  XNOR2_X1 U13477 ( .A(n13439), .B(n13440), .ZN(n13438) );
  XOR2_X1 U13478 ( .A(n13441), .B(n13442), .Z(n13210) );
  XNOR2_X1 U13479 ( .A(n13443), .B(n13444), .ZN(n13442) );
  XOR2_X1 U13480 ( .A(n13445), .B(n13446), .Z(n13247) );
  XNOR2_X1 U13481 ( .A(n13447), .B(n13448), .ZN(n13446) );
  XOR2_X1 U13482 ( .A(n13449), .B(n13450), .Z(n13252) );
  XOR2_X1 U13483 ( .A(n13451), .B(n13452), .Z(n13449) );
  XOR2_X1 U13484 ( .A(n13453), .B(n13454), .Z(n13182) );
  XOR2_X1 U13485 ( .A(n13455), .B(n13456), .Z(n13453) );
  XNOR2_X1 U13486 ( .A(n13457), .B(n13458), .ZN(n13260) );
  NAND2_X1 U13487 ( .A1(n13459), .A2(n13460), .ZN(n13457) );
  XOR2_X1 U13488 ( .A(n13461), .B(n13462), .Z(n13263) );
  XOR2_X1 U13489 ( .A(n13463), .B(n13464), .Z(n13461) );
  NOR2_X1 U13490 ( .A1(n10633), .A2(n13233), .ZN(n13464) );
  XOR2_X1 U13491 ( .A(n13465), .B(n13466), .Z(n13162) );
  XOR2_X1 U13492 ( .A(n13467), .B(n13468), .Z(n13465) );
  NOR2_X1 U13493 ( .A1(n8881), .A2(n13233), .ZN(n13468) );
  XOR2_X1 U13494 ( .A(n13469), .B(n13470), .Z(n13129) );
  XOR2_X1 U13495 ( .A(n13471), .B(n13472), .Z(n13469) );
  NOR2_X1 U13496 ( .A1(n8763), .A2(n13233), .ZN(n13472) );
  XNOR2_X1 U13497 ( .A(n13473), .B(n13474), .ZN(n13115) );
  NAND2_X1 U13498 ( .A1(n13475), .A2(n13476), .ZN(n13473) );
  XNOR2_X1 U13499 ( .A(n13477), .B(n13478), .ZN(n13107) );
  XOR2_X1 U13500 ( .A(n13479), .B(n13480), .Z(n13478) );
  XOR2_X1 U13501 ( .A(n13481), .B(n13482), .Z(n13099) );
  XNOR2_X1 U13502 ( .A(n13483), .B(n13484), .ZN(n13482) );
  XNOR2_X1 U13503 ( .A(n13485), .B(n13486), .ZN(n13091) );
  NAND2_X1 U13504 ( .A1(n13487), .A2(n13488), .ZN(n13485) );
  XOR2_X1 U13505 ( .A(n13489), .B(n13490), .Z(n13070) );
  XNOR2_X1 U13506 ( .A(n13491), .B(n13492), .ZN(n13490) );
  XNOR2_X1 U13507 ( .A(n13493), .B(n13494), .ZN(n13062) );
  NAND2_X1 U13508 ( .A1(n13495), .A2(n13496), .ZN(n13493) );
  XOR2_X1 U13509 ( .A(n13497), .B(n13498), .Z(n13054) );
  XNOR2_X1 U13510 ( .A(n13499), .B(n13500), .ZN(n13498) );
  XNOR2_X1 U13511 ( .A(n13501), .B(n13502), .ZN(n13046) );
  NAND2_X1 U13512 ( .A1(n13503), .A2(n13504), .ZN(n13501) );
  XOR2_X1 U13513 ( .A(n13505), .B(n13506), .Z(n13038) );
  XNOR2_X1 U13514 ( .A(n13507), .B(n13508), .ZN(n13506) );
  XNOR2_X1 U13515 ( .A(n13509), .B(n13510), .ZN(n13029) );
  NAND2_X1 U13516 ( .A1(n13511), .A2(n13512), .ZN(n13509) );
  XOR2_X1 U13517 ( .A(n13513), .B(n13514), .Z(n13022) );
  XNOR2_X1 U13518 ( .A(n13515), .B(n13516), .ZN(n13514) );
  XNOR2_X1 U13519 ( .A(n13517), .B(n13518), .ZN(n13020) );
  XNOR2_X1 U13520 ( .A(n13519), .B(n13520), .ZN(n13518) );
  XNOR2_X1 U13521 ( .A(n13521), .B(n13522), .ZN(n8596) );
  NAND2_X1 U13522 ( .A1(n8603), .A2(n8602), .ZN(n8601) );
  NOR2_X1 U13523 ( .A1(n13523), .A2(n8623), .ZN(n8602) );
  NOR2_X1 U13524 ( .A1(n13524), .A2(n13525), .ZN(n13523) );
  INV_X1 U13525 ( .A(n13526), .ZN(n8603) );
  NAND2_X1 U13526 ( .A1(n13522), .A2(n13521), .ZN(n13526) );
  NAND2_X1 U13527 ( .A1(n13527), .A2(n13528), .ZN(n13521) );
  NAND2_X1 U13528 ( .A1(n13520), .A2(n13529), .ZN(n13528) );
  NAND2_X1 U13529 ( .A1(n13517), .A2(n13519), .ZN(n13529) );
  NOR2_X1 U13530 ( .A1(n13233), .A2(n8690), .ZN(n13520) );
  INV_X1 U13531 ( .A(n13530), .ZN(n13527) );
  NOR2_X1 U13532 ( .A1(n13519), .A2(n13517), .ZN(n13530) );
  XNOR2_X1 U13533 ( .A(n13531), .B(n13532), .ZN(n13517) );
  XOR2_X1 U13534 ( .A(n13533), .B(n13534), .Z(n13531) );
  NOR2_X1 U13535 ( .A1(n13436), .A2(n8502), .ZN(n13534) );
  NAND2_X1 U13536 ( .A1(n13535), .A2(n13536), .ZN(n13519) );
  NAND2_X1 U13537 ( .A1(n13513), .A2(n13537), .ZN(n13536) );
  NAND2_X1 U13538 ( .A1(n13516), .A2(n13515), .ZN(n13537) );
  XNOR2_X1 U13539 ( .A(n13538), .B(n13539), .ZN(n13513) );
  XOR2_X1 U13540 ( .A(n13540), .B(n13541), .Z(n13538) );
  NOR2_X1 U13541 ( .A1(n13436), .A2(n8497), .ZN(n13541) );
  INV_X1 U13542 ( .A(n13542), .ZN(n13535) );
  NOR2_X1 U13543 ( .A1(n13515), .A2(n13516), .ZN(n13542) );
  NOR2_X1 U13544 ( .A1(n13233), .A2(n8502), .ZN(n13516) );
  NAND2_X1 U13545 ( .A1(n13511), .A2(n13543), .ZN(n13515) );
  NAND2_X1 U13546 ( .A1(n13510), .A2(n13512), .ZN(n13543) );
  NAND2_X1 U13547 ( .A1(n13544), .A2(n13545), .ZN(n13512) );
  INV_X1 U13548 ( .A(n13546), .ZN(n13545) );
  NAND2_X1 U13549 ( .A1(b_12_), .A2(a_2_), .ZN(n13544) );
  XOR2_X1 U13550 ( .A(n13547), .B(n13548), .Z(n13510) );
  XOR2_X1 U13551 ( .A(n13549), .B(n13550), .Z(n13547) );
  NOR2_X1 U13552 ( .A1(n13436), .A2(n8707), .ZN(n13550) );
  NAND2_X1 U13553 ( .A1(n13546), .A2(a_2_), .ZN(n13511) );
  NOR2_X1 U13554 ( .A1(n13551), .A2(n13552), .ZN(n13546) );
  INV_X1 U13555 ( .A(n13553), .ZN(n13552) );
  NAND2_X1 U13556 ( .A1(n13505), .A2(n13554), .ZN(n13553) );
  NAND2_X1 U13557 ( .A1(n13508), .A2(n13507), .ZN(n13554) );
  XNOR2_X1 U13558 ( .A(n13555), .B(n13556), .ZN(n13505) );
  XOR2_X1 U13559 ( .A(n13557), .B(n13558), .Z(n13555) );
  NOR2_X1 U13560 ( .A1(n13436), .A2(n8712), .ZN(n13558) );
  NOR2_X1 U13561 ( .A1(n13507), .A2(n13508), .ZN(n13551) );
  NOR2_X1 U13562 ( .A1(n13233), .A2(n8707), .ZN(n13508) );
  NAND2_X1 U13563 ( .A1(n13503), .A2(n13559), .ZN(n13507) );
  NAND2_X1 U13564 ( .A1(n13502), .A2(n13504), .ZN(n13559) );
  NAND2_X1 U13565 ( .A1(n13560), .A2(n13561), .ZN(n13504) );
  INV_X1 U13566 ( .A(n13562), .ZN(n13561) );
  NAND2_X1 U13567 ( .A1(b_12_), .A2(a_4_), .ZN(n13560) );
  XOR2_X1 U13568 ( .A(n13563), .B(n13564), .Z(n13502) );
  XOR2_X1 U13569 ( .A(n13565), .B(n13566), .Z(n13563) );
  NOR2_X1 U13570 ( .A1(n13436), .A2(n8717), .ZN(n13566) );
  NAND2_X1 U13571 ( .A1(n13562), .A2(a_4_), .ZN(n13503) );
  NOR2_X1 U13572 ( .A1(n13567), .A2(n13568), .ZN(n13562) );
  INV_X1 U13573 ( .A(n13569), .ZN(n13568) );
  NAND2_X1 U13574 ( .A1(n13497), .A2(n13570), .ZN(n13569) );
  NAND2_X1 U13575 ( .A1(n13500), .A2(n13499), .ZN(n13570) );
  XOR2_X1 U13576 ( .A(n13571), .B(n13572), .Z(n13497) );
  XOR2_X1 U13577 ( .A(n13573), .B(n13574), .Z(n13572) );
  NAND2_X1 U13578 ( .A1(a_6_), .A2(b_11_), .ZN(n13574) );
  NOR2_X1 U13579 ( .A1(n13499), .A2(n13500), .ZN(n13567) );
  NOR2_X1 U13580 ( .A1(n13233), .A2(n8717), .ZN(n13500) );
  NAND2_X1 U13581 ( .A1(n13495), .A2(n13575), .ZN(n13499) );
  NAND2_X1 U13582 ( .A1(n13494), .A2(n13496), .ZN(n13575) );
  NAND2_X1 U13583 ( .A1(n13576), .A2(n13577), .ZN(n13496) );
  INV_X1 U13584 ( .A(n13578), .ZN(n13577) );
  NAND2_X1 U13585 ( .A1(b_12_), .A2(a_6_), .ZN(n13576) );
  XNOR2_X1 U13586 ( .A(n13579), .B(n13580), .ZN(n13494) );
  XOR2_X1 U13587 ( .A(n13581), .B(n13582), .Z(n13580) );
  NAND2_X1 U13588 ( .A1(a_7_), .A2(b_11_), .ZN(n13582) );
  NAND2_X1 U13589 ( .A1(n13578), .A2(a_6_), .ZN(n13495) );
  NOR2_X1 U13590 ( .A1(n13583), .A2(n13584), .ZN(n13578) );
  INV_X1 U13591 ( .A(n13585), .ZN(n13584) );
  NAND2_X1 U13592 ( .A1(n13489), .A2(n13586), .ZN(n13585) );
  NAND2_X1 U13593 ( .A1(n13492), .A2(n13491), .ZN(n13586) );
  XNOR2_X1 U13594 ( .A(n13587), .B(n13588), .ZN(n13489) );
  XOR2_X1 U13595 ( .A(n13589), .B(n13590), .Z(n13587) );
  NOR2_X1 U13596 ( .A1(n13436), .A2(n8731), .ZN(n13590) );
  NOR2_X1 U13597 ( .A1(n13491), .A2(n13492), .ZN(n13583) );
  NOR2_X1 U13598 ( .A1(n13233), .A2(n8726), .ZN(n13492) );
  NAND2_X1 U13599 ( .A1(n13306), .A2(n13591), .ZN(n13491) );
  NAND2_X1 U13600 ( .A1(n13305), .A2(n13307), .ZN(n13591) );
  NAND2_X1 U13601 ( .A1(n13592), .A2(n13593), .ZN(n13307) );
  NAND2_X1 U13602 ( .A1(b_12_), .A2(a_8_), .ZN(n13593) );
  INV_X1 U13603 ( .A(n13594), .ZN(n13592) );
  XOR2_X1 U13604 ( .A(n13595), .B(n13596), .Z(n13305) );
  XNOR2_X1 U13605 ( .A(n13597), .B(n13598), .ZN(n13595) );
  NAND2_X1 U13606 ( .A1(a_9_), .A2(b_11_), .ZN(n13597) );
  NAND2_X1 U13607 ( .A1(a_8_), .A2(n13594), .ZN(n13306) );
  NAND2_X1 U13608 ( .A1(n13314), .A2(n13599), .ZN(n13594) );
  NAND2_X1 U13609 ( .A1(n13313), .A2(n13315), .ZN(n13599) );
  NAND2_X1 U13610 ( .A1(n13600), .A2(n13601), .ZN(n13315) );
  NAND2_X1 U13611 ( .A1(b_12_), .A2(a_9_), .ZN(n13601) );
  INV_X1 U13612 ( .A(n13602), .ZN(n13600) );
  XOR2_X1 U13613 ( .A(n13603), .B(n13604), .Z(n13313) );
  XNOR2_X1 U13614 ( .A(n13605), .B(n13606), .ZN(n13604) );
  NAND2_X1 U13615 ( .A1(a_10_), .A2(b_11_), .ZN(n13606) );
  NAND2_X1 U13616 ( .A1(a_9_), .A2(n13602), .ZN(n13314) );
  NAND2_X1 U13617 ( .A1(n13487), .A2(n13607), .ZN(n13602) );
  NAND2_X1 U13618 ( .A1(n13486), .A2(n13488), .ZN(n13607) );
  NAND2_X1 U13619 ( .A1(n13608), .A2(n13609), .ZN(n13488) );
  NAND2_X1 U13620 ( .A1(b_12_), .A2(a_10_), .ZN(n13608) );
  XOR2_X1 U13621 ( .A(n13610), .B(n13611), .Z(n13486) );
  XOR2_X1 U13622 ( .A(n13612), .B(n13613), .Z(n13611) );
  NAND2_X1 U13623 ( .A1(n13614), .A2(a_10_), .ZN(n13487) );
  INV_X1 U13624 ( .A(n13609), .ZN(n13614) );
  NAND2_X1 U13625 ( .A1(n13615), .A2(n13616), .ZN(n13609) );
  NAND2_X1 U13626 ( .A1(n13481), .A2(n13617), .ZN(n13616) );
  INV_X1 U13627 ( .A(n13618), .ZN(n13617) );
  NOR2_X1 U13628 ( .A1(n13484), .A2(n13483), .ZN(n13618) );
  XNOR2_X1 U13629 ( .A(n13619), .B(n13620), .ZN(n13481) );
  XOR2_X1 U13630 ( .A(n13621), .B(n13622), .Z(n13619) );
  NOR2_X1 U13631 ( .A1(n13436), .A2(n8750), .ZN(n13622) );
  NAND2_X1 U13632 ( .A1(n13483), .A2(n13484), .ZN(n13615) );
  NAND2_X1 U13633 ( .A1(b_12_), .A2(a_11_), .ZN(n13484) );
  NOR2_X1 U13634 ( .A1(n13623), .A2(n13624), .ZN(n13483) );
  NOR2_X1 U13635 ( .A1(n13479), .A2(n13625), .ZN(n13624) );
  NOR2_X1 U13636 ( .A1(n13480), .A2(n13477), .ZN(n13625) );
  INV_X1 U13637 ( .A(n13626), .ZN(n13623) );
  NAND2_X1 U13638 ( .A1(n13477), .A2(n13480), .ZN(n13626) );
  NAND2_X1 U13639 ( .A1(n13475), .A2(n13627), .ZN(n13480) );
  NAND2_X1 U13640 ( .A1(n13474), .A2(n13476), .ZN(n13627) );
  NAND2_X1 U13641 ( .A1(n13628), .A2(n13629), .ZN(n13476) );
  NAND2_X1 U13642 ( .A1(b_12_), .A2(a_13_), .ZN(n13629) );
  INV_X1 U13643 ( .A(n13630), .ZN(n13628) );
  XNOR2_X1 U13644 ( .A(n13631), .B(n13632), .ZN(n13474) );
  XOR2_X1 U13645 ( .A(n13633), .B(n13634), .Z(n13632) );
  NAND2_X1 U13646 ( .A1(a_14_), .A2(b_11_), .ZN(n13634) );
  NAND2_X1 U13647 ( .A1(a_13_), .A2(n13630), .ZN(n13475) );
  NAND2_X1 U13648 ( .A1(n13339), .A2(n13635), .ZN(n13630) );
  NAND2_X1 U13649 ( .A1(n13338), .A2(n13340), .ZN(n13635) );
  NAND2_X1 U13650 ( .A1(n13636), .A2(n13637), .ZN(n13340) );
  NAND2_X1 U13651 ( .A1(b_12_), .A2(a_14_), .ZN(n13637) );
  INV_X1 U13652 ( .A(n13638), .ZN(n13636) );
  XNOR2_X1 U13653 ( .A(n13639), .B(n13640), .ZN(n13338) );
  XOR2_X1 U13654 ( .A(n13641), .B(n13642), .Z(n13640) );
  NAND2_X1 U13655 ( .A1(a_15_), .A2(b_11_), .ZN(n13642) );
  NAND2_X1 U13656 ( .A1(a_14_), .A2(n13638), .ZN(n13339) );
  NAND2_X1 U13657 ( .A1(n13643), .A2(n13644), .ZN(n13638) );
  NAND2_X1 U13658 ( .A1(n13645), .A2(b_12_), .ZN(n13644) );
  NOR2_X1 U13659 ( .A1(n13646), .A2(n8763), .ZN(n13645) );
  NOR2_X1 U13660 ( .A1(n13470), .A2(n13471), .ZN(n13646) );
  NAND2_X1 U13661 ( .A1(n13470), .A2(n13471), .ZN(n13643) );
  NAND2_X1 U13662 ( .A1(n13351), .A2(n13647), .ZN(n13471) );
  NAND2_X1 U13663 ( .A1(n13350), .A2(n13352), .ZN(n13647) );
  NAND2_X1 U13664 ( .A1(n13648), .A2(n13649), .ZN(n13352) );
  NAND2_X1 U13665 ( .A1(b_12_), .A2(a_16_), .ZN(n13649) );
  INV_X1 U13666 ( .A(n13650), .ZN(n13648) );
  XOR2_X1 U13667 ( .A(n13651), .B(n13652), .Z(n13350) );
  XNOR2_X1 U13668 ( .A(n13653), .B(n13654), .ZN(n13652) );
  NAND2_X1 U13669 ( .A1(a_16_), .A2(n13650), .ZN(n13351) );
  NAND2_X1 U13670 ( .A1(n13655), .A2(n13656), .ZN(n13650) );
  NAND2_X1 U13671 ( .A1(n13657), .A2(b_12_), .ZN(n13656) );
  NOR2_X1 U13672 ( .A1(n13658), .A2(n8772), .ZN(n13657) );
  NOR2_X1 U13673 ( .A1(n13359), .A2(n13358), .ZN(n13658) );
  NAND2_X1 U13674 ( .A1(n13358), .A2(n13359), .ZN(n13655) );
  NAND2_X1 U13675 ( .A1(n13659), .A2(n13660), .ZN(n13359) );
  NAND2_X1 U13676 ( .A1(n13661), .A2(b_12_), .ZN(n13660) );
  NOR2_X1 U13677 ( .A1(n13662), .A2(n10616), .ZN(n13661) );
  NOR2_X1 U13678 ( .A1(n13366), .A2(n13367), .ZN(n13662) );
  NAND2_X1 U13679 ( .A1(n13366), .A2(n13367), .ZN(n13659) );
  NAND2_X1 U13680 ( .A1(n13663), .A2(n13664), .ZN(n13367) );
  NAND2_X1 U13681 ( .A1(n13665), .A2(b_12_), .ZN(n13664) );
  NOR2_X1 U13682 ( .A1(n13666), .A2(n8881), .ZN(n13665) );
  NOR2_X1 U13683 ( .A1(n13466), .A2(n13467), .ZN(n13666) );
  NAND2_X1 U13684 ( .A1(n13466), .A2(n13467), .ZN(n13663) );
  NAND2_X1 U13685 ( .A1(n13667), .A2(n13668), .ZN(n13467) );
  NAND2_X1 U13686 ( .A1(n13669), .A2(b_12_), .ZN(n13668) );
  NOR2_X1 U13687 ( .A1(n13670), .A2(n10633), .ZN(n13669) );
  NOR2_X1 U13688 ( .A1(n13463), .A2(n13462), .ZN(n13670) );
  NAND2_X1 U13689 ( .A1(n13462), .A2(n13463), .ZN(n13667) );
  NAND2_X1 U13690 ( .A1(n13459), .A2(n13671), .ZN(n13463) );
  NAND2_X1 U13691 ( .A1(n13458), .A2(n13460), .ZN(n13671) );
  NAND2_X1 U13692 ( .A1(n13672), .A2(n13673), .ZN(n13460) );
  NAND2_X1 U13693 ( .A1(b_12_), .A2(a_21_), .ZN(n13673) );
  INV_X1 U13694 ( .A(n13674), .ZN(n13672) );
  XNOR2_X1 U13695 ( .A(n13675), .B(n13676), .ZN(n13458) );
  XNOR2_X1 U13696 ( .A(n13677), .B(n13678), .ZN(n13676) );
  NAND2_X1 U13697 ( .A1(a_21_), .A2(n13674), .ZN(n13459) );
  NAND2_X1 U13698 ( .A1(n13679), .A2(n13680), .ZN(n13674) );
  NAND2_X1 U13699 ( .A1(n13388), .A2(n13681), .ZN(n13680) );
  INV_X1 U13700 ( .A(n13682), .ZN(n13681) );
  NOR2_X1 U13701 ( .A1(n13385), .A2(n13387), .ZN(n13682) );
  NOR2_X1 U13702 ( .A1(n13233), .A2(n8803), .ZN(n13388) );
  NAND2_X1 U13703 ( .A1(n13385), .A2(n13387), .ZN(n13679) );
  NAND2_X1 U13704 ( .A1(n13683), .A2(n13684), .ZN(n13387) );
  NAND2_X1 U13705 ( .A1(n13456), .A2(n13685), .ZN(n13684) );
  INV_X1 U13706 ( .A(n13686), .ZN(n13685) );
  NOR2_X1 U13707 ( .A1(n13455), .A2(n13454), .ZN(n13686) );
  NOR2_X1 U13708 ( .A1(n13233), .A2(n8812), .ZN(n13456) );
  NAND2_X1 U13709 ( .A1(n13454), .A2(n13455), .ZN(n13683) );
  NAND2_X1 U13710 ( .A1(n13687), .A2(n13688), .ZN(n13455) );
  NAND2_X1 U13711 ( .A1(n13452), .A2(n13689), .ZN(n13688) );
  INV_X1 U13712 ( .A(n13690), .ZN(n13689) );
  NOR2_X1 U13713 ( .A1(n13450), .A2(n13451), .ZN(n13690) );
  NOR2_X1 U13714 ( .A1(n13233), .A2(n9131), .ZN(n13452) );
  NAND2_X1 U13715 ( .A1(n13450), .A2(n13451), .ZN(n13687) );
  NAND2_X1 U13716 ( .A1(n13691), .A2(n13692), .ZN(n13451) );
  NAND2_X1 U13717 ( .A1(n13448), .A2(n13693), .ZN(n13692) );
  NAND2_X1 U13718 ( .A1(n13445), .A2(n13447), .ZN(n13693) );
  NOR2_X1 U13719 ( .A1(n13233), .A2(n8825), .ZN(n13448) );
  INV_X1 U13720 ( .A(n13694), .ZN(n13691) );
  NOR2_X1 U13721 ( .A1(n13447), .A2(n13445), .ZN(n13694) );
  XNOR2_X1 U13722 ( .A(n13695), .B(n13696), .ZN(n13445) );
  XNOR2_X1 U13723 ( .A(n13697), .B(n13698), .ZN(n13696) );
  NAND2_X1 U13724 ( .A1(n13699), .A2(n13700), .ZN(n13447) );
  NAND2_X1 U13725 ( .A1(n13406), .A2(n13701), .ZN(n13700) );
  NAND2_X1 U13726 ( .A1(n13408), .A2(n13407), .ZN(n13701) );
  XNOR2_X1 U13727 ( .A(n13702), .B(n13703), .ZN(n13406) );
  XNOR2_X1 U13728 ( .A(n13704), .B(n13705), .ZN(n13702) );
  INV_X1 U13729 ( .A(n13706), .ZN(n13699) );
  NOR2_X1 U13730 ( .A1(n13407), .A2(n13408), .ZN(n13706) );
  NOR2_X1 U13731 ( .A1(n13233), .A2(n8830), .ZN(n13408) );
  NAND2_X1 U13732 ( .A1(n13707), .A2(n13708), .ZN(n13407) );
  INV_X1 U13733 ( .A(n13709), .ZN(n13708) );
  NOR2_X1 U13734 ( .A1(n13415), .A2(n13710), .ZN(n13709) );
  NOR2_X1 U13735 ( .A1(n13414), .A2(n13416), .ZN(n13710) );
  NAND2_X1 U13736 ( .A1(b_12_), .A2(a_27_), .ZN(n13415) );
  NAND2_X1 U13737 ( .A1(n13414), .A2(n13416), .ZN(n13707) );
  NAND2_X1 U13738 ( .A1(n13711), .A2(n13712), .ZN(n13416) );
  NAND2_X1 U13739 ( .A1(n13444), .A2(n13713), .ZN(n13712) );
  INV_X1 U13740 ( .A(n13714), .ZN(n13713) );
  NOR2_X1 U13741 ( .A1(n13443), .A2(n13441), .ZN(n13714) );
  NOR2_X1 U13742 ( .A1(n13233), .A2(n8844), .ZN(n13444) );
  NAND2_X1 U13743 ( .A1(n13441), .A2(n13443), .ZN(n13711) );
  NAND2_X1 U13744 ( .A1(n13715), .A2(n13716), .ZN(n13443) );
  NAND2_X1 U13745 ( .A1(n13437), .A2(n13717), .ZN(n13716) );
  INV_X1 U13746 ( .A(n13718), .ZN(n13717) );
  NOR2_X1 U13747 ( .A1(n13440), .A2(n13439), .ZN(n13718) );
  NOR2_X1 U13748 ( .A1(n13233), .A2(n9161), .ZN(n13437) );
  NAND2_X1 U13749 ( .A1(n13439), .A2(n13440), .ZN(n13715) );
  NAND2_X1 U13750 ( .A1(n13719), .A2(n13720), .ZN(n13440) );
  NAND2_X1 U13751 ( .A1(b_10_), .A2(n13721), .ZN(n13720) );
  NAND2_X1 U13752 ( .A1(n8358), .A2(n13722), .ZN(n13721) );
  NAND2_X1 U13753 ( .A1(a_31_), .A2(n13436), .ZN(n13722) );
  NAND2_X1 U13754 ( .A1(b_11_), .A2(n13723), .ZN(n13719) );
  NAND2_X1 U13755 ( .A1(n8362), .A2(n13724), .ZN(n13723) );
  NAND2_X1 U13756 ( .A1(a_30_), .A2(n13725), .ZN(n13724) );
  NOR2_X1 U13757 ( .A1(n13726), .A2(n13233), .ZN(n13439) );
  XNOR2_X1 U13758 ( .A(n13727), .B(n13728), .ZN(n13441) );
  XNOR2_X1 U13759 ( .A(n13729), .B(n13730), .ZN(n13728) );
  XNOR2_X1 U13760 ( .A(n13731), .B(n13732), .ZN(n13414) );
  XNOR2_X1 U13761 ( .A(n13733), .B(n13734), .ZN(n13732) );
  XNOR2_X1 U13762 ( .A(n13735), .B(n13736), .ZN(n13450) );
  XNOR2_X1 U13763 ( .A(n13737), .B(n13738), .ZN(n13736) );
  XNOR2_X1 U13764 ( .A(n13739), .B(n13740), .ZN(n13454) );
  XNOR2_X1 U13765 ( .A(n13741), .B(n13742), .ZN(n13739) );
  XOR2_X1 U13766 ( .A(n13743), .B(n13744), .Z(n13385) );
  XOR2_X1 U13767 ( .A(n13745), .B(n13746), .Z(n13743) );
  XOR2_X1 U13768 ( .A(n13747), .B(n13748), .Z(n13462) );
  XOR2_X1 U13769 ( .A(n13749), .B(n13750), .Z(n13747) );
  XOR2_X1 U13770 ( .A(n13751), .B(n13752), .Z(n13466) );
  XOR2_X1 U13771 ( .A(n13753), .B(n13754), .Z(n13751) );
  XOR2_X1 U13772 ( .A(n13755), .B(n13756), .Z(n13366) );
  XNOR2_X1 U13773 ( .A(n13757), .B(n13758), .ZN(n13755) );
  XOR2_X1 U13774 ( .A(n13759), .B(n13760), .Z(n13358) );
  XOR2_X1 U13775 ( .A(n13761), .B(n13762), .Z(n13759) );
  NOR2_X1 U13776 ( .A1(n13436), .A2(n10616), .ZN(n13762) );
  XNOR2_X1 U13777 ( .A(n13763), .B(n13764), .ZN(n13470) );
  XNOR2_X1 U13778 ( .A(n13765), .B(n13766), .ZN(n13763) );
  NOR2_X1 U13779 ( .A1(n13436), .A2(n8768), .ZN(n13766) );
  XNOR2_X1 U13780 ( .A(n13767), .B(n13768), .ZN(n13477) );
  XOR2_X1 U13781 ( .A(n13769), .B(n13770), .Z(n13768) );
  NAND2_X1 U13782 ( .A1(a_13_), .A2(b_11_), .ZN(n13770) );
  XNOR2_X1 U13783 ( .A(n13771), .B(n13772), .ZN(n13522) );
  XOR2_X1 U13784 ( .A(n13773), .B(n13774), .Z(n13772) );
  NAND2_X1 U13785 ( .A1(a_0_), .A2(b_11_), .ZN(n13774) );
  INV_X1 U13786 ( .A(n13775), .ZN(n8623) );
  NAND2_X1 U13787 ( .A1(n13525), .A2(n13524), .ZN(n13775) );
  NAND2_X1 U13788 ( .A1(n13776), .A2(n13777), .ZN(n13524) );
  NAND2_X1 U13789 ( .A1(n13778), .A2(a_0_), .ZN(n13777) );
  NOR2_X1 U13790 ( .A1(n13779), .A2(n13436), .ZN(n13778) );
  NOR2_X1 U13791 ( .A1(n13771), .A2(n13773), .ZN(n13779) );
  NAND2_X1 U13792 ( .A1(n13771), .A2(n13773), .ZN(n13776) );
  NAND2_X1 U13793 ( .A1(n13780), .A2(n13781), .ZN(n13773) );
  NAND2_X1 U13794 ( .A1(n13782), .A2(a_1_), .ZN(n13781) );
  NOR2_X1 U13795 ( .A1(n13783), .A2(n13436), .ZN(n13782) );
  NOR2_X1 U13796 ( .A1(n13532), .A2(n13533), .ZN(n13783) );
  NAND2_X1 U13797 ( .A1(n13532), .A2(n13533), .ZN(n13780) );
  NAND2_X1 U13798 ( .A1(n13784), .A2(n13785), .ZN(n13533) );
  NAND2_X1 U13799 ( .A1(n13786), .A2(a_2_), .ZN(n13785) );
  NOR2_X1 U13800 ( .A1(n13787), .A2(n13436), .ZN(n13786) );
  NOR2_X1 U13801 ( .A1(n13539), .A2(n13540), .ZN(n13787) );
  NAND2_X1 U13802 ( .A1(n13539), .A2(n13540), .ZN(n13784) );
  NAND2_X1 U13803 ( .A1(n13788), .A2(n13789), .ZN(n13540) );
  NAND2_X1 U13804 ( .A1(n13790), .A2(a_3_), .ZN(n13789) );
  NOR2_X1 U13805 ( .A1(n13791), .A2(n13436), .ZN(n13790) );
  NOR2_X1 U13806 ( .A1(n13548), .A2(n13549), .ZN(n13791) );
  NAND2_X1 U13807 ( .A1(n13548), .A2(n13549), .ZN(n13788) );
  NAND2_X1 U13808 ( .A1(n13792), .A2(n13793), .ZN(n13549) );
  NAND2_X1 U13809 ( .A1(n13794), .A2(a_4_), .ZN(n13793) );
  NOR2_X1 U13810 ( .A1(n13795), .A2(n13436), .ZN(n13794) );
  NOR2_X1 U13811 ( .A1(n13556), .A2(n13557), .ZN(n13795) );
  NAND2_X1 U13812 ( .A1(n13556), .A2(n13557), .ZN(n13792) );
  NAND2_X1 U13813 ( .A1(n13796), .A2(n13797), .ZN(n13557) );
  NAND2_X1 U13814 ( .A1(n13798), .A2(a_5_), .ZN(n13797) );
  NOR2_X1 U13815 ( .A1(n13799), .A2(n13436), .ZN(n13798) );
  NOR2_X1 U13816 ( .A1(n13564), .A2(n13565), .ZN(n13799) );
  NAND2_X1 U13817 ( .A1(n13564), .A2(n13565), .ZN(n13796) );
  NAND2_X1 U13818 ( .A1(n13800), .A2(n13801), .ZN(n13565) );
  NAND2_X1 U13819 ( .A1(n13802), .A2(a_6_), .ZN(n13801) );
  NOR2_X1 U13820 ( .A1(n13803), .A2(n13436), .ZN(n13802) );
  NOR2_X1 U13821 ( .A1(n13571), .A2(n13573), .ZN(n13803) );
  NAND2_X1 U13822 ( .A1(n13571), .A2(n13573), .ZN(n13800) );
  NAND2_X1 U13823 ( .A1(n13804), .A2(n13805), .ZN(n13573) );
  NAND2_X1 U13824 ( .A1(n13806), .A2(a_7_), .ZN(n13805) );
  NOR2_X1 U13825 ( .A1(n13807), .A2(n13436), .ZN(n13806) );
  NOR2_X1 U13826 ( .A1(n13579), .A2(n13581), .ZN(n13807) );
  NAND2_X1 U13827 ( .A1(n13579), .A2(n13581), .ZN(n13804) );
  NAND2_X1 U13828 ( .A1(n13808), .A2(n13809), .ZN(n13581) );
  NAND2_X1 U13829 ( .A1(n13810), .A2(a_8_), .ZN(n13809) );
  NOR2_X1 U13830 ( .A1(n13811), .A2(n13436), .ZN(n13810) );
  NOR2_X1 U13831 ( .A1(n13588), .A2(n13589), .ZN(n13811) );
  NAND2_X1 U13832 ( .A1(n13588), .A2(n13589), .ZN(n13808) );
  NAND2_X1 U13833 ( .A1(n13812), .A2(n13813), .ZN(n13589) );
  NAND2_X1 U13834 ( .A1(n13814), .A2(a_9_), .ZN(n13813) );
  NOR2_X1 U13835 ( .A1(n13815), .A2(n13436), .ZN(n13814) );
  NOR2_X1 U13836 ( .A1(n13596), .A2(n13598), .ZN(n13815) );
  NAND2_X1 U13837 ( .A1(n13596), .A2(n13598), .ZN(n13812) );
  NAND2_X1 U13838 ( .A1(n13816), .A2(n13817), .ZN(n13598) );
  NAND2_X1 U13839 ( .A1(n13818), .A2(a_10_), .ZN(n13817) );
  NOR2_X1 U13840 ( .A1(n13819), .A2(n13436), .ZN(n13818) );
  NOR2_X1 U13841 ( .A1(n13605), .A2(n13603), .ZN(n13819) );
  NAND2_X1 U13842 ( .A1(n13605), .A2(n13603), .ZN(n13816) );
  XNOR2_X1 U13843 ( .A(n13820), .B(n13821), .ZN(n13603) );
  NAND2_X1 U13844 ( .A1(n13822), .A2(n13823), .ZN(n13820) );
  NOR2_X1 U13845 ( .A1(n13824), .A2(n13825), .ZN(n13605) );
  INV_X1 U13846 ( .A(n13826), .ZN(n13825) );
  NAND2_X1 U13847 ( .A1(n13610), .A2(n13827), .ZN(n13826) );
  NAND2_X1 U13848 ( .A1(n13828), .A2(n13612), .ZN(n13827) );
  XOR2_X1 U13849 ( .A(n13829), .B(n13830), .Z(n13610) );
  NAND2_X1 U13850 ( .A1(n13831), .A2(n13832), .ZN(n13829) );
  NOR2_X1 U13851 ( .A1(n13612), .A2(n13828), .ZN(n13824) );
  NAND2_X1 U13852 ( .A1(n13833), .A2(n13834), .ZN(n13612) );
  NAND2_X1 U13853 ( .A1(n13835), .A2(a_12_), .ZN(n13834) );
  NOR2_X1 U13854 ( .A1(n13836), .A2(n13436), .ZN(n13835) );
  NOR2_X1 U13855 ( .A1(n13620), .A2(n13621), .ZN(n13836) );
  NAND2_X1 U13856 ( .A1(n13620), .A2(n13621), .ZN(n13833) );
  NAND2_X1 U13857 ( .A1(n13837), .A2(n13838), .ZN(n13621) );
  NAND2_X1 U13858 ( .A1(n13839), .A2(a_13_), .ZN(n13838) );
  NOR2_X1 U13859 ( .A1(n13840), .A2(n13436), .ZN(n13839) );
  NOR2_X1 U13860 ( .A1(n13767), .A2(n13769), .ZN(n13840) );
  NAND2_X1 U13861 ( .A1(n13767), .A2(n13769), .ZN(n13837) );
  NAND2_X1 U13862 ( .A1(n13841), .A2(n13842), .ZN(n13769) );
  NAND2_X1 U13863 ( .A1(n13843), .A2(a_14_), .ZN(n13842) );
  NOR2_X1 U13864 ( .A1(n13844), .A2(n13436), .ZN(n13843) );
  NOR2_X1 U13865 ( .A1(n13631), .A2(n13633), .ZN(n13844) );
  NAND2_X1 U13866 ( .A1(n13631), .A2(n13633), .ZN(n13841) );
  NAND2_X1 U13867 ( .A1(n13845), .A2(n13846), .ZN(n13633) );
  NAND2_X1 U13868 ( .A1(n13847), .A2(a_15_), .ZN(n13846) );
  NOR2_X1 U13869 ( .A1(n13848), .A2(n13436), .ZN(n13847) );
  NOR2_X1 U13870 ( .A1(n13639), .A2(n13641), .ZN(n13848) );
  NAND2_X1 U13871 ( .A1(n13639), .A2(n13641), .ZN(n13845) );
  NAND2_X1 U13872 ( .A1(n13849), .A2(n13850), .ZN(n13641) );
  NAND2_X1 U13873 ( .A1(n13851), .A2(a_16_), .ZN(n13850) );
  NOR2_X1 U13874 ( .A1(n13852), .A2(n13436), .ZN(n13851) );
  NOR2_X1 U13875 ( .A1(n13765), .A2(n13764), .ZN(n13852) );
  NAND2_X1 U13876 ( .A1(n13765), .A2(n13764), .ZN(n13849) );
  XNOR2_X1 U13877 ( .A(n13853), .B(n13854), .ZN(n13764) );
  NAND2_X1 U13878 ( .A1(n13855), .A2(n13856), .ZN(n13853) );
  NOR2_X1 U13879 ( .A1(n13857), .A2(n13858), .ZN(n13765) );
  INV_X1 U13880 ( .A(n13859), .ZN(n13858) );
  NAND2_X1 U13881 ( .A1(n13651), .A2(n13860), .ZN(n13859) );
  NAND2_X1 U13882 ( .A1(n13654), .A2(n13653), .ZN(n13860) );
  XOR2_X1 U13883 ( .A(n13861), .B(n13862), .Z(n13651) );
  XNOR2_X1 U13884 ( .A(n13863), .B(n13864), .ZN(n13861) );
  NOR2_X1 U13885 ( .A1(n13725), .A2(n10616), .ZN(n13864) );
  NOR2_X1 U13886 ( .A1(n13653), .A2(n13654), .ZN(n13857) );
  NOR2_X1 U13887 ( .A1(n8772), .A2(n13436), .ZN(n13654) );
  NAND2_X1 U13888 ( .A1(n13865), .A2(n13866), .ZN(n13653) );
  NAND2_X1 U13889 ( .A1(n13867), .A2(a_18_), .ZN(n13866) );
  NOR2_X1 U13890 ( .A1(n13868), .A2(n13436), .ZN(n13867) );
  NOR2_X1 U13891 ( .A1(n13760), .A2(n13761), .ZN(n13868) );
  NAND2_X1 U13892 ( .A1(n13760), .A2(n13761), .ZN(n13865) );
  NAND2_X1 U13893 ( .A1(n13869), .A2(n13870), .ZN(n13761) );
  INV_X1 U13894 ( .A(n13871), .ZN(n13870) );
  NOR2_X1 U13895 ( .A1(n13757), .A2(n13872), .ZN(n13871) );
  NOR2_X1 U13896 ( .A1(n13758), .A2(n13756), .ZN(n13872) );
  NAND2_X1 U13897 ( .A1(b_11_), .A2(a_19_), .ZN(n13757) );
  NAND2_X1 U13898 ( .A1(n13756), .A2(n13758), .ZN(n13869) );
  NAND2_X1 U13899 ( .A1(n13873), .A2(n13874), .ZN(n13758) );
  NAND2_X1 U13900 ( .A1(n13754), .A2(n13875), .ZN(n13874) );
  INV_X1 U13901 ( .A(n13876), .ZN(n13875) );
  NOR2_X1 U13902 ( .A1(n13753), .A2(n13752), .ZN(n13876) );
  NOR2_X1 U13903 ( .A1(n10633), .A2(n13436), .ZN(n13754) );
  NAND2_X1 U13904 ( .A1(n13752), .A2(n13753), .ZN(n13873) );
  NAND2_X1 U13905 ( .A1(n13877), .A2(n13878), .ZN(n13753) );
  NAND2_X1 U13906 ( .A1(n13750), .A2(n13879), .ZN(n13878) );
  INV_X1 U13907 ( .A(n13880), .ZN(n13879) );
  NOR2_X1 U13908 ( .A1(n13749), .A2(n13748), .ZN(n13880) );
  NOR2_X1 U13909 ( .A1(n8798), .A2(n13436), .ZN(n13750) );
  NAND2_X1 U13910 ( .A1(n13748), .A2(n13749), .ZN(n13877) );
  NAND2_X1 U13911 ( .A1(n13881), .A2(n13882), .ZN(n13749) );
  NAND2_X1 U13912 ( .A1(n13678), .A2(n13883), .ZN(n13882) );
  INV_X1 U13913 ( .A(n13884), .ZN(n13883) );
  NOR2_X1 U13914 ( .A1(n13677), .A2(n13675), .ZN(n13884) );
  NOR2_X1 U13915 ( .A1(n8803), .A2(n13436), .ZN(n13678) );
  NAND2_X1 U13916 ( .A1(n13675), .A2(n13677), .ZN(n13881) );
  NAND2_X1 U13917 ( .A1(n13885), .A2(n13886), .ZN(n13677) );
  NAND2_X1 U13918 ( .A1(n13746), .A2(n13887), .ZN(n13886) );
  NAND2_X1 U13919 ( .A1(n13888), .A2(n13889), .ZN(n13887) );
  INV_X1 U13920 ( .A(n13744), .ZN(n13889) );
  INV_X1 U13921 ( .A(n13745), .ZN(n13888) );
  NOR2_X1 U13922 ( .A1(n8812), .A2(n13436), .ZN(n13746) );
  NAND2_X1 U13923 ( .A1(n13744), .A2(n13745), .ZN(n13885) );
  NAND2_X1 U13924 ( .A1(n13890), .A2(n13891), .ZN(n13745) );
  NAND2_X1 U13925 ( .A1(n13742), .A2(n13892), .ZN(n13891) );
  NAND2_X1 U13926 ( .A1(n13741), .A2(n13740), .ZN(n13892) );
  NOR2_X1 U13927 ( .A1(n9131), .A2(n13436), .ZN(n13742) );
  INV_X1 U13928 ( .A(n13893), .ZN(n13890) );
  NOR2_X1 U13929 ( .A1(n13740), .A2(n13741), .ZN(n13893) );
  NOR2_X1 U13930 ( .A1(n13894), .A2(n13895), .ZN(n13741) );
  INV_X1 U13931 ( .A(n13896), .ZN(n13895) );
  NAND2_X1 U13932 ( .A1(n13738), .A2(n13897), .ZN(n13896) );
  NAND2_X1 U13933 ( .A1(n13735), .A2(n13737), .ZN(n13897) );
  NOR2_X1 U13934 ( .A1(n8825), .A2(n13436), .ZN(n13738) );
  NOR2_X1 U13935 ( .A1(n13737), .A2(n13735), .ZN(n13894) );
  XNOR2_X1 U13936 ( .A(n13898), .B(n13899), .ZN(n13735) );
  XNOR2_X1 U13937 ( .A(n13900), .B(n13901), .ZN(n13899) );
  NAND2_X1 U13938 ( .A1(n13902), .A2(n13903), .ZN(n13737) );
  NAND2_X1 U13939 ( .A1(n13695), .A2(n13904), .ZN(n13903) );
  INV_X1 U13940 ( .A(n13905), .ZN(n13904) );
  NOR2_X1 U13941 ( .A1(n13698), .A2(n13697), .ZN(n13905) );
  XNOR2_X1 U13942 ( .A(n13906), .B(n13907), .ZN(n13695) );
  XOR2_X1 U13943 ( .A(n13908), .B(n13909), .Z(n13907) );
  NAND2_X1 U13944 ( .A1(n13697), .A2(n13698), .ZN(n13902) );
  NAND2_X1 U13945 ( .A1(a_26_), .A2(b_11_), .ZN(n13698) );
  NOR2_X1 U13946 ( .A1(n13910), .A2(n13911), .ZN(n13697) );
  NOR2_X1 U13947 ( .A1(n13704), .A2(n13912), .ZN(n13911) );
  NOR2_X1 U13948 ( .A1(n13705), .A2(n13703), .ZN(n13912) );
  NAND2_X1 U13949 ( .A1(a_27_), .A2(b_11_), .ZN(n13704) );
  INV_X1 U13950 ( .A(n13913), .ZN(n13910) );
  NAND2_X1 U13951 ( .A1(n13703), .A2(n13705), .ZN(n13913) );
  NAND2_X1 U13952 ( .A1(n13914), .A2(n13915), .ZN(n13705) );
  NAND2_X1 U13953 ( .A1(n13734), .A2(n13916), .ZN(n13915) );
  INV_X1 U13954 ( .A(n13917), .ZN(n13916) );
  NOR2_X1 U13955 ( .A1(n13733), .A2(n13731), .ZN(n13917) );
  NOR2_X1 U13956 ( .A1(n8844), .A2(n13436), .ZN(n13734) );
  NAND2_X1 U13957 ( .A1(n13731), .A2(n13733), .ZN(n13914) );
  NAND2_X1 U13958 ( .A1(n13918), .A2(n13919), .ZN(n13733) );
  NAND2_X1 U13959 ( .A1(n13727), .A2(n13920), .ZN(n13919) );
  INV_X1 U13960 ( .A(n13921), .ZN(n13920) );
  NOR2_X1 U13961 ( .A1(n13730), .A2(n13729), .ZN(n13921) );
  NOR2_X1 U13962 ( .A1(n9161), .A2(n13436), .ZN(n13727) );
  NAND2_X1 U13963 ( .A1(n13729), .A2(n13730), .ZN(n13918) );
  NAND2_X1 U13964 ( .A1(n13922), .A2(n13923), .ZN(n13730) );
  NAND2_X1 U13965 ( .A1(b_10_), .A2(n13924), .ZN(n13923) );
  NAND2_X1 U13966 ( .A1(n8362), .A2(n13925), .ZN(n13924) );
  NAND2_X1 U13967 ( .A1(a_30_), .A2(n13926), .ZN(n13925) );
  NAND2_X1 U13968 ( .A1(b_9_), .A2(n13927), .ZN(n13922) );
  NAND2_X1 U13969 ( .A1(n8358), .A2(n13928), .ZN(n13927) );
  NAND2_X1 U13970 ( .A1(a_31_), .A2(n13725), .ZN(n13928) );
  NOR2_X1 U13971 ( .A1(n13726), .A2(n13725), .ZN(n13729) );
  NAND2_X1 U13972 ( .A1(b_11_), .A2(n9926), .ZN(n13726) );
  XNOR2_X1 U13973 ( .A(n13929), .B(n13930), .ZN(n13731) );
  XOR2_X1 U13974 ( .A(n13931), .B(n13932), .Z(n13930) );
  XNOR2_X1 U13975 ( .A(n13933), .B(n13934), .ZN(n13703) );
  XNOR2_X1 U13976 ( .A(n13935), .B(n13936), .ZN(n13933) );
  XOR2_X1 U13977 ( .A(n13937), .B(n13938), .Z(n13740) );
  XNOR2_X1 U13978 ( .A(n13939), .B(n13940), .ZN(n13938) );
  XOR2_X1 U13979 ( .A(n13941), .B(n13942), .Z(n13744) );
  XOR2_X1 U13980 ( .A(n13943), .B(n13944), .Z(n13941) );
  XOR2_X1 U13981 ( .A(n13945), .B(n13946), .Z(n13675) );
  XOR2_X1 U13982 ( .A(n13947), .B(n13948), .Z(n13945) );
  XNOR2_X1 U13983 ( .A(n13949), .B(n13950), .ZN(n13748) );
  XNOR2_X1 U13984 ( .A(n13951), .B(n13952), .ZN(n13950) );
  XNOR2_X1 U13985 ( .A(n13953), .B(n13954), .ZN(n13752) );
  NAND2_X1 U13986 ( .A1(n13955), .A2(n13956), .ZN(n13953) );
  XOR2_X1 U13987 ( .A(n13957), .B(n13958), .Z(n13756) );
  XOR2_X1 U13988 ( .A(n13959), .B(n13960), .Z(n13957) );
  NOR2_X1 U13989 ( .A1(n10633), .A2(n13725), .ZN(n13960) );
  XOR2_X1 U13990 ( .A(n13961), .B(n13962), .Z(n13760) );
  XNOR2_X1 U13991 ( .A(n13963), .B(n13964), .ZN(n13962) );
  XNOR2_X1 U13992 ( .A(n13965), .B(n13966), .ZN(n13639) );
  XOR2_X1 U13993 ( .A(n13967), .B(n13968), .Z(n13965) );
  XNOR2_X1 U13994 ( .A(n13969), .B(n13970), .ZN(n13631) );
  NAND2_X1 U13995 ( .A1(n13971), .A2(n13972), .ZN(n13969) );
  XOR2_X1 U13996 ( .A(n13973), .B(n13974), .Z(n13767) );
  XNOR2_X1 U13997 ( .A(n13975), .B(n13976), .ZN(n13974) );
  XNOR2_X1 U13998 ( .A(n13977), .B(n13978), .ZN(n13620) );
  NAND2_X1 U13999 ( .A1(n13979), .A2(n13980), .ZN(n13977) );
  XOR2_X1 U14000 ( .A(n13981), .B(n13982), .Z(n13596) );
  XNOR2_X1 U14001 ( .A(n13983), .B(n13984), .ZN(n13981) );
  XNOR2_X1 U14002 ( .A(n13985), .B(n13986), .ZN(n13588) );
  NAND2_X1 U14003 ( .A1(n13987), .A2(n13988), .ZN(n13985) );
  XNOR2_X1 U14004 ( .A(n13989), .B(n13990), .ZN(n13579) );
  XOR2_X1 U14005 ( .A(n13991), .B(n13992), .Z(n13989) );
  XNOR2_X1 U14006 ( .A(n13993), .B(n13994), .ZN(n13571) );
  XNOR2_X1 U14007 ( .A(n13995), .B(n13996), .ZN(n13994) );
  XOR2_X1 U14008 ( .A(n13997), .B(n13998), .Z(n13564) );
  XOR2_X1 U14009 ( .A(n13999), .B(n14000), .Z(n13997) );
  XOR2_X1 U14010 ( .A(n14001), .B(n14002), .Z(n13556) );
  XNOR2_X1 U14011 ( .A(n14003), .B(n14004), .ZN(n14001) );
  XOR2_X1 U14012 ( .A(n14005), .B(n14006), .Z(n13548) );
  XOR2_X1 U14013 ( .A(n14007), .B(n14008), .Z(n14006) );
  XNOR2_X1 U14014 ( .A(n14009), .B(n14010), .ZN(n13539) );
  XOR2_X1 U14015 ( .A(n14011), .B(n14012), .Z(n14010) );
  XOR2_X1 U14016 ( .A(n14013), .B(n14014), .Z(n13532) );
  XOR2_X1 U14017 ( .A(n14015), .B(n14016), .Z(n14013) );
  XOR2_X1 U14018 ( .A(n14017), .B(n14018), .Z(n13771) );
  XOR2_X1 U14019 ( .A(n14019), .B(n14020), .Z(n14017) );
  XNOR2_X1 U14020 ( .A(n14021), .B(n14022), .ZN(n13525) );
  XNOR2_X1 U14021 ( .A(n14023), .B(n14024), .ZN(n14022) );
  XNOR2_X1 U14022 ( .A(n14025), .B(n14026), .ZN(n8605) );
  NAND2_X1 U14023 ( .A1(n8342), .A2(n8343), .ZN(n8341) );
  INV_X1 U14024 ( .A(n14027), .ZN(n8343) );
  NAND2_X1 U14025 ( .A1(n14026), .A2(n14025), .ZN(n14027) );
  NAND2_X1 U14026 ( .A1(n14028), .A2(n14029), .ZN(n14025) );
  NAND2_X1 U14027 ( .A1(n14024), .A2(n14030), .ZN(n14029) );
  INV_X1 U14028 ( .A(n14031), .ZN(n14030) );
  NOR2_X1 U14029 ( .A1(n14021), .A2(n14023), .ZN(n14031) );
  NOR2_X1 U14030 ( .A1(n8690), .A2(n13725), .ZN(n14024) );
  NAND2_X1 U14031 ( .A1(n14021), .A2(n14023), .ZN(n14028) );
  NAND2_X1 U14032 ( .A1(n14032), .A2(n14033), .ZN(n14023) );
  NAND2_X1 U14033 ( .A1(n14020), .A2(n14034), .ZN(n14033) );
  INV_X1 U14034 ( .A(n14035), .ZN(n14034) );
  NOR2_X1 U14035 ( .A1(n14018), .A2(n14019), .ZN(n14035) );
  NOR2_X1 U14036 ( .A1(n8502), .A2(n13725), .ZN(n14020) );
  NAND2_X1 U14037 ( .A1(n14018), .A2(n14019), .ZN(n14032) );
  NAND2_X1 U14038 ( .A1(n14036), .A2(n14037), .ZN(n14019) );
  NAND2_X1 U14039 ( .A1(n14016), .A2(n14038), .ZN(n14037) );
  NAND2_X1 U14040 ( .A1(n14039), .A2(n14040), .ZN(n14038) );
  INV_X1 U14041 ( .A(n14015), .ZN(n14040) );
  INV_X1 U14042 ( .A(n14014), .ZN(n14039) );
  NOR2_X1 U14043 ( .A1(n8497), .A2(n13725), .ZN(n14016) );
  NAND2_X1 U14044 ( .A1(n14014), .A2(n14015), .ZN(n14036) );
  NAND2_X1 U14045 ( .A1(n14041), .A2(n14042), .ZN(n14015) );
  INV_X1 U14046 ( .A(n14043), .ZN(n14042) );
  NOR2_X1 U14047 ( .A1(n14012), .A2(n14044), .ZN(n14043) );
  NOR2_X1 U14048 ( .A1(n14009), .A2(n14011), .ZN(n14044) );
  NAND2_X1 U14049 ( .A1(a_3_), .A2(b_10_), .ZN(n14012) );
  NAND2_X1 U14050 ( .A1(n14009), .A2(n14011), .ZN(n14041) );
  NAND2_X1 U14051 ( .A1(n14045), .A2(n14046), .ZN(n14011) );
  NAND2_X1 U14052 ( .A1(n14008), .A2(n14047), .ZN(n14046) );
  NAND2_X1 U14053 ( .A1(n14005), .A2(n14007), .ZN(n14047) );
  NOR2_X1 U14054 ( .A1(n8712), .A2(n13725), .ZN(n14008) );
  INV_X1 U14055 ( .A(n14048), .ZN(n14045) );
  NOR2_X1 U14056 ( .A1(n14005), .A2(n14007), .ZN(n14048) );
  NOR2_X1 U14057 ( .A1(n14049), .A2(n14050), .ZN(n14007) );
  NOR2_X1 U14058 ( .A1(n14003), .A2(n14051), .ZN(n14050) );
  NOR2_X1 U14059 ( .A1(n14002), .A2(n14004), .ZN(n14051) );
  NAND2_X1 U14060 ( .A1(a_5_), .A2(b_10_), .ZN(n14003) );
  INV_X1 U14061 ( .A(n14052), .ZN(n14049) );
  NAND2_X1 U14062 ( .A1(n14002), .A2(n14004), .ZN(n14052) );
  NAND2_X1 U14063 ( .A1(n14053), .A2(n14054), .ZN(n14004) );
  NAND2_X1 U14064 ( .A1(n14000), .A2(n14055), .ZN(n14054) );
  INV_X1 U14065 ( .A(n14056), .ZN(n14055) );
  NOR2_X1 U14066 ( .A1(n13998), .A2(n13999), .ZN(n14056) );
  NOR2_X1 U14067 ( .A1(n8480), .A2(n13725), .ZN(n14000) );
  NAND2_X1 U14068 ( .A1(n13998), .A2(n13999), .ZN(n14053) );
  NAND2_X1 U14069 ( .A1(n14057), .A2(n14058), .ZN(n13999) );
  NAND2_X1 U14070 ( .A1(n13996), .A2(n14059), .ZN(n14058) );
  NAND2_X1 U14071 ( .A1(n13993), .A2(n13995), .ZN(n14059) );
  NOR2_X1 U14072 ( .A1(n8726), .A2(n13725), .ZN(n13996) );
  INV_X1 U14073 ( .A(n14060), .ZN(n14057) );
  NOR2_X1 U14074 ( .A1(n13995), .A2(n13993), .ZN(n14060) );
  XNOR2_X1 U14075 ( .A(n14061), .B(n14062), .ZN(n13993) );
  XNOR2_X1 U14076 ( .A(n14063), .B(n14064), .ZN(n14062) );
  NAND2_X1 U14077 ( .A1(a_8_), .A2(b_9_), .ZN(n14064) );
  NAND2_X1 U14078 ( .A1(n14065), .A2(n14066), .ZN(n13995) );
  NAND2_X1 U14079 ( .A1(n13990), .A2(n14067), .ZN(n14066) );
  NAND2_X1 U14080 ( .A1(n13992), .A2(n13991), .ZN(n14067) );
  XNOR2_X1 U14081 ( .A(n14068), .B(n14069), .ZN(n13990) );
  XOR2_X1 U14082 ( .A(n14070), .B(n14071), .Z(n14068) );
  INV_X1 U14083 ( .A(n14072), .ZN(n14065) );
  NOR2_X1 U14084 ( .A1(n13991), .A2(n13992), .ZN(n14072) );
  NOR2_X1 U14085 ( .A1(n8731), .A2(n13725), .ZN(n13992) );
  NAND2_X1 U14086 ( .A1(n13987), .A2(n14073), .ZN(n13991) );
  NAND2_X1 U14087 ( .A1(n13986), .A2(n13988), .ZN(n14073) );
  NAND2_X1 U14088 ( .A1(n14074), .A2(n14075), .ZN(n13988) );
  NAND2_X1 U14089 ( .A1(a_9_), .A2(b_10_), .ZN(n14075) );
  XOR2_X1 U14090 ( .A(n14076), .B(n14077), .Z(n13986) );
  XOR2_X1 U14091 ( .A(n14078), .B(n14079), .Z(n14076) );
  NOR2_X1 U14092 ( .A1(n13926), .A2(n8741), .ZN(n14079) );
  INV_X1 U14093 ( .A(n14080), .ZN(n13987) );
  NOR2_X1 U14094 ( .A1(n8736), .A2(n14074), .ZN(n14080) );
  NOR2_X1 U14095 ( .A1(n14081), .A2(n14082), .ZN(n14074) );
  NOR2_X1 U14096 ( .A1(n13984), .A2(n14083), .ZN(n14082) );
  NOR2_X1 U14097 ( .A1(n13982), .A2(n13983), .ZN(n14083) );
  INV_X1 U14098 ( .A(n14084), .ZN(n14081) );
  NAND2_X1 U14099 ( .A1(n13982), .A2(n13983), .ZN(n14084) );
  NAND2_X1 U14100 ( .A1(n13822), .A2(n14085), .ZN(n13983) );
  NAND2_X1 U14101 ( .A1(n13821), .A2(n13823), .ZN(n14085) );
  NAND2_X1 U14102 ( .A1(n14086), .A2(n14087), .ZN(n13823) );
  NAND2_X1 U14103 ( .A1(a_11_), .A2(b_10_), .ZN(n14087) );
  INV_X1 U14104 ( .A(n14088), .ZN(n14086) );
  XOR2_X1 U14105 ( .A(n14089), .B(n14090), .Z(n13821) );
  XOR2_X1 U14106 ( .A(n14091), .B(n14092), .Z(n14089) );
  NOR2_X1 U14107 ( .A1(n13926), .A2(n8750), .ZN(n14092) );
  NAND2_X1 U14108 ( .A1(a_11_), .A2(n14088), .ZN(n13822) );
  NAND2_X1 U14109 ( .A1(n13831), .A2(n14093), .ZN(n14088) );
  NAND2_X1 U14110 ( .A1(n13830), .A2(n13832), .ZN(n14093) );
  NAND2_X1 U14111 ( .A1(n14094), .A2(n14095), .ZN(n13832) );
  NAND2_X1 U14112 ( .A1(a_12_), .A2(b_10_), .ZN(n14095) );
  INV_X1 U14113 ( .A(n14096), .ZN(n14094) );
  XOR2_X1 U14114 ( .A(n14097), .B(n14098), .Z(n13830) );
  XOR2_X1 U14115 ( .A(n14099), .B(n14100), .Z(n14097) );
  NOR2_X1 U14116 ( .A1(n13926), .A2(n8443), .ZN(n14100) );
  NAND2_X1 U14117 ( .A1(a_12_), .A2(n14096), .ZN(n13831) );
  NAND2_X1 U14118 ( .A1(n13979), .A2(n14101), .ZN(n14096) );
  NAND2_X1 U14119 ( .A1(n13978), .A2(n13980), .ZN(n14101) );
  NAND2_X1 U14120 ( .A1(n14102), .A2(n14103), .ZN(n13980) );
  INV_X1 U14121 ( .A(n14104), .ZN(n14103) );
  NAND2_X1 U14122 ( .A1(a_13_), .A2(b_10_), .ZN(n14102) );
  XNOR2_X1 U14123 ( .A(n14105), .B(n14106), .ZN(n13978) );
  NAND2_X1 U14124 ( .A1(n14107), .A2(n14108), .ZN(n14105) );
  NAND2_X1 U14125 ( .A1(n14104), .A2(a_13_), .ZN(n13979) );
  NOR2_X1 U14126 ( .A1(n14109), .A2(n14110), .ZN(n14104) );
  INV_X1 U14127 ( .A(n14111), .ZN(n14110) );
  NAND2_X1 U14128 ( .A1(n13973), .A2(n14112), .ZN(n14111) );
  NAND2_X1 U14129 ( .A1(n13976), .A2(n13975), .ZN(n14112) );
  XNOR2_X1 U14130 ( .A(n14113), .B(n14114), .ZN(n13973) );
  XOR2_X1 U14131 ( .A(n14115), .B(n14116), .Z(n14113) );
  NOR2_X1 U14132 ( .A1(n13926), .A2(n8763), .ZN(n14116) );
  NOR2_X1 U14133 ( .A1(n13975), .A2(n13976), .ZN(n14109) );
  NOR2_X1 U14134 ( .A1(n8438), .A2(n13725), .ZN(n13976) );
  NAND2_X1 U14135 ( .A1(n13971), .A2(n14117), .ZN(n13975) );
  NAND2_X1 U14136 ( .A1(n13970), .A2(n13972), .ZN(n14117) );
  NAND2_X1 U14137 ( .A1(n14118), .A2(n14119), .ZN(n13972) );
  INV_X1 U14138 ( .A(n14120), .ZN(n14119) );
  NAND2_X1 U14139 ( .A1(a_15_), .A2(b_10_), .ZN(n14118) );
  XOR2_X1 U14140 ( .A(n14121), .B(n14122), .Z(n13970) );
  XOR2_X1 U14141 ( .A(n14123), .B(n14124), .Z(n14121) );
  NOR2_X1 U14142 ( .A1(n13926), .A2(n8768), .ZN(n14124) );
  NAND2_X1 U14143 ( .A1(n14120), .A2(a_15_), .ZN(n13971) );
  NOR2_X1 U14144 ( .A1(n14125), .A2(n14126), .ZN(n14120) );
  INV_X1 U14145 ( .A(n14127), .ZN(n14126) );
  NAND2_X1 U14146 ( .A1(n13966), .A2(n14128), .ZN(n14127) );
  NAND2_X1 U14147 ( .A1(n13968), .A2(n13967), .ZN(n14128) );
  XNOR2_X1 U14148 ( .A(n14129), .B(n14130), .ZN(n13966) );
  XOR2_X1 U14149 ( .A(n14131), .B(n14132), .Z(n14129) );
  NOR2_X1 U14150 ( .A1(n13926), .A2(n8772), .ZN(n14132) );
  NOR2_X1 U14151 ( .A1(n13967), .A2(n13968), .ZN(n14125) );
  NOR2_X1 U14152 ( .A1(n8768), .A2(n13725), .ZN(n13968) );
  NAND2_X1 U14153 ( .A1(n13855), .A2(n14133), .ZN(n13967) );
  NAND2_X1 U14154 ( .A1(n13854), .A2(n13856), .ZN(n14133) );
  NAND2_X1 U14155 ( .A1(n14134), .A2(n14135), .ZN(n13856) );
  NAND2_X1 U14156 ( .A1(a_17_), .A2(b_10_), .ZN(n14135) );
  INV_X1 U14157 ( .A(n14136), .ZN(n14134) );
  XOR2_X1 U14158 ( .A(n14137), .B(n14138), .Z(n13854) );
  XOR2_X1 U14159 ( .A(n14139), .B(n14140), .Z(n14137) );
  NOR2_X1 U14160 ( .A1(n13926), .A2(n10616), .ZN(n14140) );
  NAND2_X1 U14161 ( .A1(a_17_), .A2(n14136), .ZN(n13855) );
  NAND2_X1 U14162 ( .A1(n14141), .A2(n14142), .ZN(n14136) );
  NAND2_X1 U14163 ( .A1(n14143), .A2(a_18_), .ZN(n14142) );
  NOR2_X1 U14164 ( .A1(n14144), .A2(n13725), .ZN(n14143) );
  NOR2_X1 U14165 ( .A1(n13863), .A2(n13862), .ZN(n14144) );
  NAND2_X1 U14166 ( .A1(n13863), .A2(n13862), .ZN(n14141) );
  XOR2_X1 U14167 ( .A(n14145), .B(n14146), .Z(n13862) );
  XOR2_X1 U14168 ( .A(n14147), .B(n14148), .Z(n14145) );
  NOR2_X1 U14169 ( .A1(n8881), .A2(n13926), .ZN(n14148) );
  NOR2_X1 U14170 ( .A1(n14149), .A2(n14150), .ZN(n13863) );
  INV_X1 U14171 ( .A(n14151), .ZN(n14150) );
  NAND2_X1 U14172 ( .A1(n13961), .A2(n14152), .ZN(n14151) );
  NAND2_X1 U14173 ( .A1(n13964), .A2(n13963), .ZN(n14152) );
  XNOR2_X1 U14174 ( .A(n14153), .B(n14154), .ZN(n13961) );
  XOR2_X1 U14175 ( .A(n14155), .B(n14156), .Z(n14153) );
  NOR2_X1 U14176 ( .A1(n10633), .A2(n13926), .ZN(n14156) );
  NOR2_X1 U14177 ( .A1(n13963), .A2(n13964), .ZN(n14149) );
  NOR2_X1 U14178 ( .A1(n13725), .A2(n8881), .ZN(n13964) );
  NAND2_X1 U14179 ( .A1(n14157), .A2(n14158), .ZN(n13963) );
  NAND2_X1 U14180 ( .A1(n14159), .A2(b_10_), .ZN(n14158) );
  NOR2_X1 U14181 ( .A1(n14160), .A2(n10633), .ZN(n14159) );
  NOR2_X1 U14182 ( .A1(n13958), .A2(n13959), .ZN(n14160) );
  NAND2_X1 U14183 ( .A1(n13958), .A2(n13959), .ZN(n14157) );
  NAND2_X1 U14184 ( .A1(n13955), .A2(n14161), .ZN(n13959) );
  NAND2_X1 U14185 ( .A1(n13954), .A2(n13956), .ZN(n14161) );
  NAND2_X1 U14186 ( .A1(n14162), .A2(n14163), .ZN(n13956) );
  NAND2_X1 U14187 ( .A1(b_10_), .A2(a_21_), .ZN(n14163) );
  INV_X1 U14188 ( .A(n14164), .ZN(n14162) );
  XNOR2_X1 U14189 ( .A(n14165), .B(n14166), .ZN(n13954) );
  XNOR2_X1 U14190 ( .A(n14167), .B(n14168), .ZN(n14166) );
  NAND2_X1 U14191 ( .A1(a_21_), .A2(n14164), .ZN(n13955) );
  NAND2_X1 U14192 ( .A1(n14169), .A2(n14170), .ZN(n14164) );
  NAND2_X1 U14193 ( .A1(n13952), .A2(n14171), .ZN(n14170) );
  INV_X1 U14194 ( .A(n14172), .ZN(n14171) );
  NOR2_X1 U14195 ( .A1(n13949), .A2(n13951), .ZN(n14172) );
  NOR2_X1 U14196 ( .A1(n13725), .A2(n8803), .ZN(n13952) );
  NAND2_X1 U14197 ( .A1(n13949), .A2(n13951), .ZN(n14169) );
  NAND2_X1 U14198 ( .A1(n14173), .A2(n14174), .ZN(n13951) );
  NAND2_X1 U14199 ( .A1(n13948), .A2(n14175), .ZN(n14174) );
  INV_X1 U14200 ( .A(n14176), .ZN(n14175) );
  NOR2_X1 U14201 ( .A1(n13947), .A2(n13946), .ZN(n14176) );
  NOR2_X1 U14202 ( .A1(n13725), .A2(n8812), .ZN(n13948) );
  NAND2_X1 U14203 ( .A1(n13946), .A2(n13947), .ZN(n14173) );
  NAND2_X1 U14204 ( .A1(n14177), .A2(n14178), .ZN(n13947) );
  NAND2_X1 U14205 ( .A1(n13944), .A2(n14179), .ZN(n14178) );
  INV_X1 U14206 ( .A(n14180), .ZN(n14179) );
  NOR2_X1 U14207 ( .A1(n13942), .A2(n13943), .ZN(n14180) );
  NOR2_X1 U14208 ( .A1(n13725), .A2(n9131), .ZN(n13944) );
  NAND2_X1 U14209 ( .A1(n13942), .A2(n13943), .ZN(n14177) );
  NAND2_X1 U14210 ( .A1(n14181), .A2(n14182), .ZN(n13943) );
  NAND2_X1 U14211 ( .A1(n13940), .A2(n14183), .ZN(n14182) );
  NAND2_X1 U14212 ( .A1(n13937), .A2(n13939), .ZN(n14183) );
  NOR2_X1 U14213 ( .A1(n13725), .A2(n8825), .ZN(n13940) );
  INV_X1 U14214 ( .A(n14184), .ZN(n14181) );
  NOR2_X1 U14215 ( .A1(n13939), .A2(n13937), .ZN(n14184) );
  XNOR2_X1 U14216 ( .A(n14185), .B(n14186), .ZN(n13937) );
  XNOR2_X1 U14217 ( .A(n14187), .B(n14188), .ZN(n14186) );
  NAND2_X1 U14218 ( .A1(n14189), .A2(n14190), .ZN(n13939) );
  NAND2_X1 U14219 ( .A1(n13898), .A2(n14191), .ZN(n14190) );
  NAND2_X1 U14220 ( .A1(n13901), .A2(n13900), .ZN(n14191) );
  XNOR2_X1 U14221 ( .A(n14192), .B(n14193), .ZN(n13898) );
  XOR2_X1 U14222 ( .A(n14194), .B(n14195), .Z(n14193) );
  INV_X1 U14223 ( .A(n14196), .ZN(n14189) );
  NOR2_X1 U14224 ( .A1(n13900), .A2(n13901), .ZN(n14196) );
  NOR2_X1 U14225 ( .A1(n8830), .A2(n13725), .ZN(n13901) );
  NAND2_X1 U14226 ( .A1(n14197), .A2(n14198), .ZN(n13900) );
  NAND2_X1 U14227 ( .A1(n13909), .A2(n14199), .ZN(n14198) );
  NAND2_X1 U14228 ( .A1(n13906), .A2(n13908), .ZN(n14199) );
  NOR2_X1 U14229 ( .A1(n13725), .A2(n8839), .ZN(n13909) );
  INV_X1 U14230 ( .A(n14200), .ZN(n14197) );
  NOR2_X1 U14231 ( .A1(n13906), .A2(n13908), .ZN(n14200) );
  NOR2_X1 U14232 ( .A1(n14201), .A2(n14202), .ZN(n13908) );
  INV_X1 U14233 ( .A(n14203), .ZN(n14202) );
  NAND2_X1 U14234 ( .A1(n13935), .A2(n14204), .ZN(n14203) );
  NAND2_X1 U14235 ( .A1(n13936), .A2(n13934), .ZN(n14204) );
  NOR2_X1 U14236 ( .A1(n13725), .A2(n8844), .ZN(n13935) );
  NOR2_X1 U14237 ( .A1(n13934), .A2(n13936), .ZN(n14201) );
  NOR2_X1 U14238 ( .A1(n14205), .A2(n14206), .ZN(n13936) );
  INV_X1 U14239 ( .A(n14207), .ZN(n14206) );
  NAND2_X1 U14240 ( .A1(n13929), .A2(n14208), .ZN(n14207) );
  NAND2_X1 U14241 ( .A1(n14209), .A2(n13931), .ZN(n14208) );
  NOR2_X1 U14242 ( .A1(n13725), .A2(n9161), .ZN(n13929) );
  NOR2_X1 U14243 ( .A1(n13931), .A2(n14209), .ZN(n14205) );
  INV_X1 U14244 ( .A(n13932), .ZN(n14209) );
  NAND2_X1 U14245 ( .A1(n14210), .A2(n14211), .ZN(n13932) );
  NAND2_X1 U14246 ( .A1(b_8_), .A2(n14212), .ZN(n14211) );
  NAND2_X1 U14247 ( .A1(n8358), .A2(n14213), .ZN(n14212) );
  NAND2_X1 U14248 ( .A1(a_31_), .A2(n13926), .ZN(n14213) );
  NAND2_X1 U14249 ( .A1(b_9_), .A2(n14214), .ZN(n14210) );
  NAND2_X1 U14250 ( .A1(n8362), .A2(n14215), .ZN(n14214) );
  NAND2_X1 U14251 ( .A1(a_30_), .A2(n14216), .ZN(n14215) );
  NAND2_X1 U14252 ( .A1(n14217), .A2(b_9_), .ZN(n13931) );
  NOR2_X1 U14253 ( .A1(n9170), .A2(n13725), .ZN(n14217) );
  XOR2_X1 U14254 ( .A(n14218), .B(n14219), .Z(n13934) );
  XOR2_X1 U14255 ( .A(n14220), .B(n14221), .Z(n14219) );
  XOR2_X1 U14256 ( .A(n14222), .B(n14223), .Z(n13906) );
  XNOR2_X1 U14257 ( .A(n14224), .B(n14225), .ZN(n14222) );
  XNOR2_X1 U14258 ( .A(n14226), .B(n14227), .ZN(n13942) );
  XNOR2_X1 U14259 ( .A(n14228), .B(n14229), .ZN(n14227) );
  XOR2_X1 U14260 ( .A(n14230), .B(n14231), .Z(n13946) );
  XOR2_X1 U14261 ( .A(n14232), .B(n14233), .Z(n14230) );
  XOR2_X1 U14262 ( .A(n14234), .B(n14235), .Z(n13949) );
  XOR2_X1 U14263 ( .A(n14236), .B(n14237), .Z(n14234) );
  XNOR2_X1 U14264 ( .A(n14238), .B(n14239), .ZN(n13958) );
  NAND2_X1 U14265 ( .A1(n14240), .A2(n14241), .ZN(n14238) );
  XOR2_X1 U14266 ( .A(n14242), .B(n14243), .Z(n13982) );
  XOR2_X1 U14267 ( .A(n14244), .B(n14245), .Z(n14242) );
  NOR2_X1 U14268 ( .A1(n13926), .A2(n8452), .ZN(n14245) );
  XOR2_X1 U14269 ( .A(n14246), .B(n14247), .Z(n13998) );
  XNOR2_X1 U14270 ( .A(n14248), .B(n14249), .ZN(n14246) );
  NAND2_X1 U14271 ( .A1(a_7_), .A2(b_9_), .ZN(n14248) );
  XOR2_X1 U14272 ( .A(n14250), .B(n14251), .Z(n14002) );
  XOR2_X1 U14273 ( .A(n14252), .B(n14253), .Z(n14250) );
  NOR2_X1 U14274 ( .A1(n13926), .A2(n8480), .ZN(n14253) );
  XNOR2_X1 U14275 ( .A(n14254), .B(n14255), .ZN(n14005) );
  XOR2_X1 U14276 ( .A(n14256), .B(n14257), .Z(n14254) );
  NOR2_X1 U14277 ( .A1(n13926), .A2(n8717), .ZN(n14257) );
  XOR2_X1 U14278 ( .A(n14258), .B(n14259), .Z(n14009) );
  XOR2_X1 U14279 ( .A(n14260), .B(n14261), .Z(n14258) );
  NOR2_X1 U14280 ( .A1(n13926), .A2(n8712), .ZN(n14261) );
  XNOR2_X1 U14281 ( .A(n14262), .B(n14263), .ZN(n14014) );
  XOR2_X1 U14282 ( .A(n14264), .B(n14265), .Z(n14263) );
  NAND2_X1 U14283 ( .A1(a_3_), .A2(b_9_), .ZN(n14265) );
  XOR2_X1 U14284 ( .A(n14266), .B(n14267), .Z(n14018) );
  XOR2_X1 U14285 ( .A(n14268), .B(n14269), .Z(n14266) );
  NOR2_X1 U14286 ( .A1(n13926), .A2(n8497), .ZN(n14269) );
  XOR2_X1 U14287 ( .A(n14270), .B(n14271), .Z(n14021) );
  XOR2_X1 U14288 ( .A(n14272), .B(n14273), .Z(n14270) );
  NOR2_X1 U14289 ( .A1(n13926), .A2(n8502), .ZN(n14273) );
  XOR2_X1 U14290 ( .A(n14274), .B(n14275), .Z(n14026) );
  XOR2_X1 U14291 ( .A(n14276), .B(n14277), .Z(n14274) );
  NOR2_X1 U14292 ( .A1(n13926), .A2(n8690), .ZN(n14277) );
  NOR2_X1 U14293 ( .A1(n14278), .A2(n8621), .ZN(n8342) );
  INV_X1 U14294 ( .A(n14279), .ZN(n8621) );
  NAND2_X1 U14295 ( .A1(n14280), .A2(n14281), .ZN(n14279) );
  NOR2_X1 U14296 ( .A1(n14281), .A2(n14280), .ZN(n14278) );
  XNOR2_X1 U14297 ( .A(n14282), .B(n14283), .ZN(n14280) );
  XNOR2_X1 U14298 ( .A(n14284), .B(n14285), .ZN(n14282) );
  NAND2_X1 U14299 ( .A1(n14286), .A2(n14287), .ZN(n14281) );
  NAND2_X1 U14300 ( .A1(n14288), .A2(a_0_), .ZN(n14287) );
  NOR2_X1 U14301 ( .A1(n14289), .A2(n13926), .ZN(n14288) );
  NOR2_X1 U14302 ( .A1(n14275), .A2(n14276), .ZN(n14289) );
  NAND2_X1 U14303 ( .A1(n14275), .A2(n14276), .ZN(n14286) );
  NAND2_X1 U14304 ( .A1(n14290), .A2(n14291), .ZN(n14276) );
  NAND2_X1 U14305 ( .A1(n14292), .A2(a_1_), .ZN(n14291) );
  NOR2_X1 U14306 ( .A1(n14293), .A2(n13926), .ZN(n14292) );
  NOR2_X1 U14307 ( .A1(n14271), .A2(n14272), .ZN(n14293) );
  NAND2_X1 U14308 ( .A1(n14271), .A2(n14272), .ZN(n14290) );
  NAND2_X1 U14309 ( .A1(n14294), .A2(n14295), .ZN(n14272) );
  NAND2_X1 U14310 ( .A1(n14296), .A2(a_2_), .ZN(n14295) );
  NOR2_X1 U14311 ( .A1(n14297), .A2(n13926), .ZN(n14296) );
  NOR2_X1 U14312 ( .A1(n14267), .A2(n14268), .ZN(n14297) );
  NAND2_X1 U14313 ( .A1(n14267), .A2(n14268), .ZN(n14294) );
  NAND2_X1 U14314 ( .A1(n14298), .A2(n14299), .ZN(n14268) );
  NAND2_X1 U14315 ( .A1(n14300), .A2(a_3_), .ZN(n14299) );
  NOR2_X1 U14316 ( .A1(n14301), .A2(n13926), .ZN(n14300) );
  NOR2_X1 U14317 ( .A1(n14262), .A2(n14264), .ZN(n14301) );
  NAND2_X1 U14318 ( .A1(n14262), .A2(n14264), .ZN(n14298) );
  NAND2_X1 U14319 ( .A1(n14302), .A2(n14303), .ZN(n14264) );
  NAND2_X1 U14320 ( .A1(n14304), .A2(a_4_), .ZN(n14303) );
  NOR2_X1 U14321 ( .A1(n14305), .A2(n13926), .ZN(n14304) );
  NOR2_X1 U14322 ( .A1(n14259), .A2(n14260), .ZN(n14305) );
  NAND2_X1 U14323 ( .A1(n14259), .A2(n14260), .ZN(n14302) );
  NAND2_X1 U14324 ( .A1(n14306), .A2(n14307), .ZN(n14260) );
  NAND2_X1 U14325 ( .A1(n14308), .A2(a_5_), .ZN(n14307) );
  NOR2_X1 U14326 ( .A1(n14309), .A2(n13926), .ZN(n14308) );
  NOR2_X1 U14327 ( .A1(n14255), .A2(n14256), .ZN(n14309) );
  NAND2_X1 U14328 ( .A1(n14255), .A2(n14256), .ZN(n14306) );
  NAND2_X1 U14329 ( .A1(n14310), .A2(n14311), .ZN(n14256) );
  NAND2_X1 U14330 ( .A1(n14312), .A2(a_6_), .ZN(n14311) );
  NOR2_X1 U14331 ( .A1(n14313), .A2(n13926), .ZN(n14312) );
  NOR2_X1 U14332 ( .A1(n14251), .A2(n14252), .ZN(n14313) );
  NAND2_X1 U14333 ( .A1(n14251), .A2(n14252), .ZN(n14310) );
  NAND2_X1 U14334 ( .A1(n14314), .A2(n14315), .ZN(n14252) );
  NAND2_X1 U14335 ( .A1(n14316), .A2(a_7_), .ZN(n14315) );
  NOR2_X1 U14336 ( .A1(n14317), .A2(n13926), .ZN(n14316) );
  NOR2_X1 U14337 ( .A1(n14247), .A2(n14249), .ZN(n14317) );
  NAND2_X1 U14338 ( .A1(n14247), .A2(n14249), .ZN(n14314) );
  NAND2_X1 U14339 ( .A1(n14318), .A2(n14319), .ZN(n14249) );
  NAND2_X1 U14340 ( .A1(n14320), .A2(a_8_), .ZN(n14319) );
  NOR2_X1 U14341 ( .A1(n14321), .A2(n13926), .ZN(n14320) );
  NOR2_X1 U14342 ( .A1(n14063), .A2(n14061), .ZN(n14321) );
  NAND2_X1 U14343 ( .A1(n14063), .A2(n14061), .ZN(n14318) );
  XNOR2_X1 U14344 ( .A(n14322), .B(n14323), .ZN(n14061) );
  XOR2_X1 U14345 ( .A(n14324), .B(n14325), .Z(n14323) );
  NOR2_X1 U14346 ( .A1(n14326), .A2(n14327), .ZN(n14063) );
  NOR2_X1 U14347 ( .A1(n14069), .A2(n14328), .ZN(n14327) );
  NOR2_X1 U14348 ( .A1(n14329), .A2(n14330), .ZN(n14328) );
  INV_X1 U14349 ( .A(n14070), .ZN(n14330) );
  XNOR2_X1 U14350 ( .A(n14331), .B(n14332), .ZN(n14069) );
  XOR2_X1 U14351 ( .A(n14333), .B(n14334), .Z(n14332) );
  NOR2_X1 U14352 ( .A1(n14070), .A2(n14071), .ZN(n14326) );
  NAND2_X1 U14353 ( .A1(n14335), .A2(n14336), .ZN(n14070) );
  NAND2_X1 U14354 ( .A1(n14337), .A2(a_10_), .ZN(n14336) );
  NOR2_X1 U14355 ( .A1(n14338), .A2(n13926), .ZN(n14337) );
  NOR2_X1 U14356 ( .A1(n14078), .A2(n14077), .ZN(n14338) );
  NAND2_X1 U14357 ( .A1(n14077), .A2(n14078), .ZN(n14335) );
  NAND2_X1 U14358 ( .A1(n14339), .A2(n14340), .ZN(n14078) );
  NAND2_X1 U14359 ( .A1(n14341), .A2(a_11_), .ZN(n14340) );
  NOR2_X1 U14360 ( .A1(n14342), .A2(n13926), .ZN(n14341) );
  NOR2_X1 U14361 ( .A1(n14243), .A2(n14244), .ZN(n14342) );
  NAND2_X1 U14362 ( .A1(n14243), .A2(n14244), .ZN(n14339) );
  NAND2_X1 U14363 ( .A1(n14343), .A2(n14344), .ZN(n14244) );
  NAND2_X1 U14364 ( .A1(n14345), .A2(a_12_), .ZN(n14344) );
  NOR2_X1 U14365 ( .A1(n14346), .A2(n13926), .ZN(n14345) );
  NOR2_X1 U14366 ( .A1(n14090), .A2(n14091), .ZN(n14346) );
  NAND2_X1 U14367 ( .A1(n14090), .A2(n14091), .ZN(n14343) );
  NAND2_X1 U14368 ( .A1(n14347), .A2(n14348), .ZN(n14091) );
  NAND2_X1 U14369 ( .A1(n14349), .A2(a_13_), .ZN(n14348) );
  NOR2_X1 U14370 ( .A1(n14350), .A2(n13926), .ZN(n14349) );
  NOR2_X1 U14371 ( .A1(n14098), .A2(n14099), .ZN(n14350) );
  NAND2_X1 U14372 ( .A1(n14098), .A2(n14099), .ZN(n14347) );
  NAND2_X1 U14373 ( .A1(n14107), .A2(n14351), .ZN(n14099) );
  NAND2_X1 U14374 ( .A1(n14106), .A2(n14108), .ZN(n14351) );
  NAND2_X1 U14375 ( .A1(n14352), .A2(n14353), .ZN(n14108) );
  NAND2_X1 U14376 ( .A1(a_14_), .A2(b_9_), .ZN(n14353) );
  INV_X1 U14377 ( .A(n14354), .ZN(n14352) );
  XNOR2_X1 U14378 ( .A(n14355), .B(n14356), .ZN(n14106) );
  NAND2_X1 U14379 ( .A1(n14357), .A2(n14358), .ZN(n14355) );
  NAND2_X1 U14380 ( .A1(a_14_), .A2(n14354), .ZN(n14107) );
  NAND2_X1 U14381 ( .A1(n14359), .A2(n14360), .ZN(n14354) );
  NAND2_X1 U14382 ( .A1(n14361), .A2(a_15_), .ZN(n14360) );
  NOR2_X1 U14383 ( .A1(n14362), .A2(n13926), .ZN(n14361) );
  NOR2_X1 U14384 ( .A1(n14115), .A2(n14114), .ZN(n14362) );
  NAND2_X1 U14385 ( .A1(n14114), .A2(n14115), .ZN(n14359) );
  NAND2_X1 U14386 ( .A1(n14363), .A2(n14364), .ZN(n14115) );
  NAND2_X1 U14387 ( .A1(n14365), .A2(a_16_), .ZN(n14364) );
  NOR2_X1 U14388 ( .A1(n14366), .A2(n13926), .ZN(n14365) );
  NOR2_X1 U14389 ( .A1(n14122), .A2(n14123), .ZN(n14366) );
  NAND2_X1 U14390 ( .A1(n14122), .A2(n14123), .ZN(n14363) );
  NAND2_X1 U14391 ( .A1(n14367), .A2(n14368), .ZN(n14123) );
  NAND2_X1 U14392 ( .A1(n14369), .A2(a_17_), .ZN(n14368) );
  NOR2_X1 U14393 ( .A1(n14370), .A2(n13926), .ZN(n14369) );
  NOR2_X1 U14394 ( .A1(n14130), .A2(n14131), .ZN(n14370) );
  NAND2_X1 U14395 ( .A1(n14130), .A2(n14131), .ZN(n14367) );
  NAND2_X1 U14396 ( .A1(n14371), .A2(n14372), .ZN(n14131) );
  NAND2_X1 U14397 ( .A1(n14373), .A2(a_18_), .ZN(n14372) );
  NOR2_X1 U14398 ( .A1(n14374), .A2(n13926), .ZN(n14373) );
  NOR2_X1 U14399 ( .A1(n14139), .A2(n14138), .ZN(n14374) );
  NAND2_X1 U14400 ( .A1(n14138), .A2(n14139), .ZN(n14371) );
  NAND2_X1 U14401 ( .A1(n14375), .A2(n14376), .ZN(n14139) );
  NAND2_X1 U14402 ( .A1(n14377), .A2(b_9_), .ZN(n14376) );
  NOR2_X1 U14403 ( .A1(n14378), .A2(n8881), .ZN(n14377) );
  NOR2_X1 U14404 ( .A1(n14146), .A2(n14147), .ZN(n14378) );
  NAND2_X1 U14405 ( .A1(n14146), .A2(n14147), .ZN(n14375) );
  NAND2_X1 U14406 ( .A1(n14379), .A2(n14380), .ZN(n14147) );
  NAND2_X1 U14407 ( .A1(n14381), .A2(b_9_), .ZN(n14380) );
  NOR2_X1 U14408 ( .A1(n14382), .A2(n10633), .ZN(n14381) );
  NOR2_X1 U14409 ( .A1(n14154), .A2(n14155), .ZN(n14382) );
  NAND2_X1 U14410 ( .A1(n14154), .A2(n14155), .ZN(n14379) );
  NAND2_X1 U14411 ( .A1(n14240), .A2(n14383), .ZN(n14155) );
  NAND2_X1 U14412 ( .A1(n14239), .A2(n14241), .ZN(n14383) );
  NAND2_X1 U14413 ( .A1(n14384), .A2(n14385), .ZN(n14241) );
  NAND2_X1 U14414 ( .A1(b_9_), .A2(a_21_), .ZN(n14385) );
  INV_X1 U14415 ( .A(n14386), .ZN(n14384) );
  XNOR2_X1 U14416 ( .A(n14387), .B(n14388), .ZN(n14239) );
  XOR2_X1 U14417 ( .A(n14389), .B(n14390), .Z(n14388) );
  NAND2_X1 U14418 ( .A1(a_21_), .A2(n14386), .ZN(n14240) );
  NAND2_X1 U14419 ( .A1(n14391), .A2(n14392), .ZN(n14386) );
  NAND2_X1 U14420 ( .A1(n14168), .A2(n14393), .ZN(n14392) );
  INV_X1 U14421 ( .A(n14394), .ZN(n14393) );
  NOR2_X1 U14422 ( .A1(n14167), .A2(n14165), .ZN(n14394) );
  NOR2_X1 U14423 ( .A1(n13926), .A2(n8803), .ZN(n14168) );
  NAND2_X1 U14424 ( .A1(n14165), .A2(n14167), .ZN(n14391) );
  NAND2_X1 U14425 ( .A1(n14395), .A2(n14396), .ZN(n14167) );
  NAND2_X1 U14426 ( .A1(n14237), .A2(n14397), .ZN(n14396) );
  INV_X1 U14427 ( .A(n14398), .ZN(n14397) );
  NOR2_X1 U14428 ( .A1(n14236), .A2(n14235), .ZN(n14398) );
  NOR2_X1 U14429 ( .A1(n13926), .A2(n8812), .ZN(n14237) );
  NAND2_X1 U14430 ( .A1(n14235), .A2(n14236), .ZN(n14395) );
  NAND2_X1 U14431 ( .A1(n14399), .A2(n14400), .ZN(n14236) );
  NAND2_X1 U14432 ( .A1(n14233), .A2(n14401), .ZN(n14400) );
  INV_X1 U14433 ( .A(n14402), .ZN(n14401) );
  NOR2_X1 U14434 ( .A1(n14231), .A2(n14232), .ZN(n14402) );
  NOR2_X1 U14435 ( .A1(n13926), .A2(n9131), .ZN(n14233) );
  NAND2_X1 U14436 ( .A1(n14231), .A2(n14232), .ZN(n14399) );
  NAND2_X1 U14437 ( .A1(n14403), .A2(n14404), .ZN(n14232) );
  NAND2_X1 U14438 ( .A1(n14229), .A2(n14405), .ZN(n14404) );
  NAND2_X1 U14439 ( .A1(n14226), .A2(n14228), .ZN(n14405) );
  NOR2_X1 U14440 ( .A1(n13926), .A2(n8825), .ZN(n14229) );
  INV_X1 U14441 ( .A(n14406), .ZN(n14403) );
  NOR2_X1 U14442 ( .A1(n14228), .A2(n14226), .ZN(n14406) );
  XNOR2_X1 U14443 ( .A(n14407), .B(n14408), .ZN(n14226) );
  XNOR2_X1 U14444 ( .A(n14409), .B(n14410), .ZN(n14408) );
  NAND2_X1 U14445 ( .A1(n14411), .A2(n14412), .ZN(n14228) );
  NAND2_X1 U14446 ( .A1(n14185), .A2(n14413), .ZN(n14412) );
  NAND2_X1 U14447 ( .A1(n14188), .A2(n14187), .ZN(n14413) );
  XNOR2_X1 U14448 ( .A(n14414), .B(n14415), .ZN(n14185) );
  XOR2_X1 U14449 ( .A(n14416), .B(n14417), .Z(n14415) );
  INV_X1 U14450 ( .A(n14418), .ZN(n14411) );
  NOR2_X1 U14451 ( .A1(n14187), .A2(n14188), .ZN(n14418) );
  NOR2_X1 U14452 ( .A1(n8830), .A2(n13926), .ZN(n14188) );
  NAND2_X1 U14453 ( .A1(n14419), .A2(n14420), .ZN(n14187) );
  NAND2_X1 U14454 ( .A1(n14195), .A2(n14421), .ZN(n14420) );
  NAND2_X1 U14455 ( .A1(n14192), .A2(n14194), .ZN(n14421) );
  NOR2_X1 U14456 ( .A1(n13926), .A2(n8839), .ZN(n14195) );
  INV_X1 U14457 ( .A(n14422), .ZN(n14419) );
  NOR2_X1 U14458 ( .A1(n14192), .A2(n14194), .ZN(n14422) );
  NOR2_X1 U14459 ( .A1(n14423), .A2(n14424), .ZN(n14194) );
  INV_X1 U14460 ( .A(n14425), .ZN(n14424) );
  NAND2_X1 U14461 ( .A1(n14224), .A2(n14426), .ZN(n14425) );
  NAND2_X1 U14462 ( .A1(n14225), .A2(n14223), .ZN(n14426) );
  NOR2_X1 U14463 ( .A1(n13926), .A2(n8844), .ZN(n14224) );
  NOR2_X1 U14464 ( .A1(n14223), .A2(n14225), .ZN(n14423) );
  NOR2_X1 U14465 ( .A1(n14427), .A2(n14428), .ZN(n14225) );
  INV_X1 U14466 ( .A(n14429), .ZN(n14428) );
  NAND2_X1 U14467 ( .A1(n14218), .A2(n14430), .ZN(n14429) );
  NAND2_X1 U14468 ( .A1(n14431), .A2(n14220), .ZN(n14430) );
  NOR2_X1 U14469 ( .A1(n13926), .A2(n9161), .ZN(n14218) );
  NOR2_X1 U14470 ( .A1(n14220), .A2(n14431), .ZN(n14427) );
  INV_X1 U14471 ( .A(n14221), .ZN(n14431) );
  NAND2_X1 U14472 ( .A1(n14432), .A2(n14433), .ZN(n14221) );
  NAND2_X1 U14473 ( .A1(b_7_), .A2(n14434), .ZN(n14433) );
  NAND2_X1 U14474 ( .A1(n8358), .A2(n14435), .ZN(n14434) );
  NAND2_X1 U14475 ( .A1(a_31_), .A2(n14216), .ZN(n14435) );
  NAND2_X1 U14476 ( .A1(b_8_), .A2(n14436), .ZN(n14432) );
  NAND2_X1 U14477 ( .A1(n8362), .A2(n14437), .ZN(n14436) );
  NAND2_X1 U14478 ( .A1(a_30_), .A2(n14438), .ZN(n14437) );
  NAND2_X1 U14479 ( .A1(n14439), .A2(b_8_), .ZN(n14220) );
  NOR2_X1 U14480 ( .A1(n9170), .A2(n13926), .ZN(n14439) );
  XOR2_X1 U14481 ( .A(n14440), .B(n14441), .Z(n14223) );
  XOR2_X1 U14482 ( .A(n14442), .B(n14443), .Z(n14441) );
  XOR2_X1 U14483 ( .A(n14444), .B(n14445), .Z(n14192) );
  XNOR2_X1 U14484 ( .A(n14446), .B(n14447), .ZN(n14444) );
  XNOR2_X1 U14485 ( .A(n14448), .B(n14449), .ZN(n14231) );
  XNOR2_X1 U14486 ( .A(n14450), .B(n14451), .ZN(n14449) );
  XOR2_X1 U14487 ( .A(n14452), .B(n14453), .Z(n14235) );
  XOR2_X1 U14488 ( .A(n14454), .B(n14455), .Z(n14452) );
  XOR2_X1 U14489 ( .A(n14456), .B(n14457), .Z(n14165) );
  XOR2_X1 U14490 ( .A(n14458), .B(n14459), .Z(n14456) );
  XOR2_X1 U14491 ( .A(n14460), .B(n14461), .Z(n14154) );
  XOR2_X1 U14492 ( .A(n14462), .B(n14463), .Z(n14460) );
  XOR2_X1 U14493 ( .A(n14464), .B(n14465), .Z(n14146) );
  XOR2_X1 U14494 ( .A(n14466), .B(n14467), .Z(n14464) );
  XNOR2_X1 U14495 ( .A(n14468), .B(n14469), .ZN(n14138) );
  NAND2_X1 U14496 ( .A1(n14470), .A2(n14471), .ZN(n14468) );
  XOR2_X1 U14497 ( .A(n14472), .B(n14473), .Z(n14130) );
  XNOR2_X1 U14498 ( .A(n14474), .B(n14475), .ZN(n14473) );
  XNOR2_X1 U14499 ( .A(n14476), .B(n14477), .ZN(n14122) );
  NAND2_X1 U14500 ( .A1(n14478), .A2(n14479), .ZN(n14476) );
  XOR2_X1 U14501 ( .A(n14480), .B(n14481), .Z(n14114) );
  XNOR2_X1 U14502 ( .A(n14482), .B(n14483), .ZN(n14481) );
  XOR2_X1 U14503 ( .A(n14484), .B(n14485), .Z(n14098) );
  XNOR2_X1 U14504 ( .A(n14486), .B(n14487), .ZN(n14485) );
  XOR2_X1 U14505 ( .A(n14488), .B(n14489), .Z(n14090) );
  XOR2_X1 U14506 ( .A(n14490), .B(n14491), .Z(n14489) );
  XNOR2_X1 U14507 ( .A(n14492), .B(n14493), .ZN(n14243) );
  XOR2_X1 U14508 ( .A(n14494), .B(n14495), .Z(n14493) );
  XNOR2_X1 U14509 ( .A(n14496), .B(n14497), .ZN(n14077) );
  XNOR2_X1 U14510 ( .A(n14498), .B(n14499), .ZN(n14497) );
  XNOR2_X1 U14511 ( .A(n14500), .B(n14501), .ZN(n14247) );
  XOR2_X1 U14512 ( .A(n14502), .B(n14503), .Z(n14501) );
  XOR2_X1 U14513 ( .A(n14504), .B(n14505), .Z(n14251) );
  XOR2_X1 U14514 ( .A(n14506), .B(n14507), .Z(n14504) );
  XNOR2_X1 U14515 ( .A(n14508), .B(n14509), .ZN(n14255) );
  XNOR2_X1 U14516 ( .A(n14510), .B(n14511), .ZN(n14509) );
  XOR2_X1 U14517 ( .A(n14512), .B(n14513), .Z(n14259) );
  XOR2_X1 U14518 ( .A(n14514), .B(n14515), .Z(n14512) );
  XOR2_X1 U14519 ( .A(n14516), .B(n14517), .Z(n14262) );
  XOR2_X1 U14520 ( .A(n14518), .B(n14519), .Z(n14516) );
  XNOR2_X1 U14521 ( .A(n14520), .B(n14521), .ZN(n14267) );
  XNOR2_X1 U14522 ( .A(n14522), .B(n14523), .ZN(n14521) );
  XOR2_X1 U14523 ( .A(n14524), .B(n14525), .Z(n14271) );
  XOR2_X1 U14524 ( .A(n14526), .B(n14527), .Z(n14524) );
  XOR2_X1 U14525 ( .A(n14528), .B(n14529), .Z(n14275) );
  XOR2_X1 U14526 ( .A(n14530), .B(n14531), .Z(n14528) );
  XNOR2_X1 U14527 ( .A(n14532), .B(n14533), .ZN(n8345) );
  NAND2_X1 U14528 ( .A1(n8351), .A2(n8352), .ZN(n8350) );
  INV_X1 U14529 ( .A(n14534), .ZN(n8352) );
  NAND2_X1 U14530 ( .A1(n14533), .A2(n14532), .ZN(n14534) );
  NAND2_X1 U14531 ( .A1(n14535), .A2(n14536), .ZN(n14532) );
  NAND2_X1 U14532 ( .A1(n14285), .A2(n14537), .ZN(n14536) );
  INV_X1 U14533 ( .A(n14538), .ZN(n14537) );
  NOR2_X1 U14534 ( .A1(n14283), .A2(n14284), .ZN(n14538) );
  NOR2_X1 U14535 ( .A1(n8690), .A2(n14216), .ZN(n14285) );
  NAND2_X1 U14536 ( .A1(n14283), .A2(n14284), .ZN(n14535) );
  NAND2_X1 U14537 ( .A1(n14539), .A2(n14540), .ZN(n14284) );
  NAND2_X1 U14538 ( .A1(n14531), .A2(n14541), .ZN(n14540) );
  INV_X1 U14539 ( .A(n14542), .ZN(n14541) );
  NOR2_X1 U14540 ( .A1(n14529), .A2(n14530), .ZN(n14542) );
  NOR2_X1 U14541 ( .A1(n8502), .A2(n14216), .ZN(n14531) );
  NAND2_X1 U14542 ( .A1(n14529), .A2(n14530), .ZN(n14539) );
  NAND2_X1 U14543 ( .A1(n14543), .A2(n14544), .ZN(n14530) );
  NAND2_X1 U14544 ( .A1(n14526), .A2(n14545), .ZN(n14544) );
  INV_X1 U14545 ( .A(n14546), .ZN(n14545) );
  NOR2_X1 U14546 ( .A1(n14525), .A2(n14527), .ZN(n14546) );
  NOR2_X1 U14547 ( .A1(n8497), .A2(n14216), .ZN(n14526) );
  NAND2_X1 U14548 ( .A1(n14525), .A2(n14527), .ZN(n14543) );
  NAND2_X1 U14549 ( .A1(n14547), .A2(n14548), .ZN(n14527) );
  NAND2_X1 U14550 ( .A1(n14523), .A2(n14549), .ZN(n14548) );
  INV_X1 U14551 ( .A(n14550), .ZN(n14549) );
  NOR2_X1 U14552 ( .A1(n14520), .A2(n14522), .ZN(n14550) );
  NOR2_X1 U14553 ( .A1(n8707), .A2(n14216), .ZN(n14523) );
  NAND2_X1 U14554 ( .A1(n14520), .A2(n14522), .ZN(n14547) );
  NAND2_X1 U14555 ( .A1(n14551), .A2(n14552), .ZN(n14522) );
  NAND2_X1 U14556 ( .A1(n14519), .A2(n14553), .ZN(n14552) );
  INV_X1 U14557 ( .A(n14554), .ZN(n14553) );
  NOR2_X1 U14558 ( .A1(n14517), .A2(n14518), .ZN(n14554) );
  NOR2_X1 U14559 ( .A1(n8712), .A2(n14216), .ZN(n14519) );
  NAND2_X1 U14560 ( .A1(n14517), .A2(n14518), .ZN(n14551) );
  NAND2_X1 U14561 ( .A1(n14555), .A2(n14556), .ZN(n14518) );
  NAND2_X1 U14562 ( .A1(n14515), .A2(n14557), .ZN(n14556) );
  INV_X1 U14563 ( .A(n14558), .ZN(n14557) );
  NOR2_X1 U14564 ( .A1(n14513), .A2(n14514), .ZN(n14558) );
  NOR2_X1 U14565 ( .A1(n8717), .A2(n14216), .ZN(n14515) );
  NAND2_X1 U14566 ( .A1(n14513), .A2(n14514), .ZN(n14555) );
  NAND2_X1 U14567 ( .A1(n14559), .A2(n14560), .ZN(n14514) );
  NAND2_X1 U14568 ( .A1(n14511), .A2(n14561), .ZN(n14560) );
  INV_X1 U14569 ( .A(n14562), .ZN(n14561) );
  NOR2_X1 U14570 ( .A1(n14508), .A2(n14510), .ZN(n14562) );
  NOR2_X1 U14571 ( .A1(n8480), .A2(n14216), .ZN(n14511) );
  NAND2_X1 U14572 ( .A1(n14508), .A2(n14510), .ZN(n14559) );
  NAND2_X1 U14573 ( .A1(n14563), .A2(n14564), .ZN(n14510) );
  NAND2_X1 U14574 ( .A1(n14507), .A2(n14565), .ZN(n14564) );
  NAND2_X1 U14575 ( .A1(n14505), .A2(n14506), .ZN(n14565) );
  NOR2_X1 U14576 ( .A1(n8726), .A2(n14216), .ZN(n14507) );
  INV_X1 U14577 ( .A(n14566), .ZN(n14563) );
  NOR2_X1 U14578 ( .A1(n14505), .A2(n14506), .ZN(n14566) );
  NAND2_X1 U14579 ( .A1(n14567), .A2(n14568), .ZN(n14506) );
  NAND2_X1 U14580 ( .A1(n14569), .A2(n14503), .ZN(n14568) );
  NAND2_X1 U14581 ( .A1(n14500), .A2(n14502), .ZN(n14569) );
  INV_X1 U14582 ( .A(n14570), .ZN(n14567) );
  NOR2_X1 U14583 ( .A1(n14500), .A2(n14502), .ZN(n14570) );
  NAND2_X1 U14584 ( .A1(n14571), .A2(n14572), .ZN(n14502) );
  NAND2_X1 U14585 ( .A1(n14325), .A2(n14573), .ZN(n14572) );
  NAND2_X1 U14586 ( .A1(n14324), .A2(n14574), .ZN(n14573) );
  INV_X1 U14587 ( .A(n14322), .ZN(n14574) );
  NOR2_X1 U14588 ( .A1(n8736), .A2(n14216), .ZN(n14325) );
  NAND2_X1 U14589 ( .A1(n14322), .A2(n14575), .ZN(n14571) );
  INV_X1 U14590 ( .A(n14324), .ZN(n14575) );
  NOR2_X1 U14591 ( .A1(n14576), .A2(n14577), .ZN(n14324) );
  NOR2_X1 U14592 ( .A1(n14334), .A2(n14578), .ZN(n14577) );
  NOR2_X1 U14593 ( .A1(n14333), .A2(n14331), .ZN(n14578) );
  NAND2_X1 U14594 ( .A1(a_10_), .A2(b_8_), .ZN(n14334) );
  INV_X1 U14595 ( .A(n14579), .ZN(n14576) );
  NAND2_X1 U14596 ( .A1(n14331), .A2(n14333), .ZN(n14579) );
  NAND2_X1 U14597 ( .A1(n14580), .A2(n14581), .ZN(n14333) );
  NAND2_X1 U14598 ( .A1(n14499), .A2(n14582), .ZN(n14581) );
  INV_X1 U14599 ( .A(n14583), .ZN(n14582) );
  NOR2_X1 U14600 ( .A1(n14498), .A2(n14496), .ZN(n14583) );
  NOR2_X1 U14601 ( .A1(n8452), .A2(n14216), .ZN(n14499) );
  NAND2_X1 U14602 ( .A1(n14496), .A2(n14498), .ZN(n14580) );
  NAND2_X1 U14603 ( .A1(n14584), .A2(n14585), .ZN(n14498) );
  INV_X1 U14604 ( .A(n14586), .ZN(n14585) );
  NOR2_X1 U14605 ( .A1(n14495), .A2(n14587), .ZN(n14586) );
  NOR2_X1 U14606 ( .A1(n14492), .A2(n14494), .ZN(n14587) );
  NAND2_X1 U14607 ( .A1(a_12_), .A2(b_8_), .ZN(n14495) );
  NAND2_X1 U14608 ( .A1(n14492), .A2(n14494), .ZN(n14584) );
  NAND2_X1 U14609 ( .A1(n14588), .A2(n14589), .ZN(n14494) );
  NAND2_X1 U14610 ( .A1(n14491), .A2(n14590), .ZN(n14589) );
  INV_X1 U14611 ( .A(n14591), .ZN(n14590) );
  NOR2_X1 U14612 ( .A1(n14488), .A2(n14490), .ZN(n14591) );
  NOR2_X1 U14613 ( .A1(n8443), .A2(n14216), .ZN(n14491) );
  NAND2_X1 U14614 ( .A1(n14488), .A2(n14490), .ZN(n14588) );
  NOR2_X1 U14615 ( .A1(n14592), .A2(n14593), .ZN(n14490) );
  INV_X1 U14616 ( .A(n14594), .ZN(n14593) );
  NAND2_X1 U14617 ( .A1(n14484), .A2(n14595), .ZN(n14594) );
  NAND2_X1 U14618 ( .A1(n14487), .A2(n14486), .ZN(n14595) );
  XNOR2_X1 U14619 ( .A(n14596), .B(n14597), .ZN(n14484) );
  XOR2_X1 U14620 ( .A(n14598), .B(n14599), .Z(n14596) );
  NOR2_X1 U14621 ( .A1(n14438), .A2(n8763), .ZN(n14599) );
  NOR2_X1 U14622 ( .A1(n14486), .A2(n14487), .ZN(n14592) );
  NOR2_X1 U14623 ( .A1(n8438), .A2(n14216), .ZN(n14487) );
  NAND2_X1 U14624 ( .A1(n14357), .A2(n14600), .ZN(n14486) );
  NAND2_X1 U14625 ( .A1(n14356), .A2(n14358), .ZN(n14600) );
  NAND2_X1 U14626 ( .A1(n14601), .A2(n14602), .ZN(n14358) );
  INV_X1 U14627 ( .A(n14603), .ZN(n14602) );
  NAND2_X1 U14628 ( .A1(a_15_), .A2(b_8_), .ZN(n14601) );
  XOR2_X1 U14629 ( .A(n14604), .B(n14605), .Z(n14356) );
  XOR2_X1 U14630 ( .A(n14606), .B(n14607), .Z(n14604) );
  NOR2_X1 U14631 ( .A1(n14438), .A2(n8768), .ZN(n14607) );
  NAND2_X1 U14632 ( .A1(n14603), .A2(a_15_), .ZN(n14357) );
  NOR2_X1 U14633 ( .A1(n14608), .A2(n14609), .ZN(n14603) );
  INV_X1 U14634 ( .A(n14610), .ZN(n14609) );
  NAND2_X1 U14635 ( .A1(n14480), .A2(n14611), .ZN(n14610) );
  NAND2_X1 U14636 ( .A1(n14483), .A2(n14482), .ZN(n14611) );
  XNOR2_X1 U14637 ( .A(n14612), .B(n14613), .ZN(n14480) );
  XOR2_X1 U14638 ( .A(n14614), .B(n14615), .Z(n14612) );
  NOR2_X1 U14639 ( .A1(n14438), .A2(n8772), .ZN(n14615) );
  NOR2_X1 U14640 ( .A1(n14482), .A2(n14483), .ZN(n14608) );
  NOR2_X1 U14641 ( .A1(n8768), .A2(n14216), .ZN(n14483) );
  NAND2_X1 U14642 ( .A1(n14478), .A2(n14616), .ZN(n14482) );
  NAND2_X1 U14643 ( .A1(n14477), .A2(n14479), .ZN(n14616) );
  NAND2_X1 U14644 ( .A1(n14617), .A2(n14618), .ZN(n14479) );
  INV_X1 U14645 ( .A(n14619), .ZN(n14618) );
  NAND2_X1 U14646 ( .A1(a_17_), .A2(b_8_), .ZN(n14617) );
  XOR2_X1 U14647 ( .A(n14620), .B(n14621), .Z(n14477) );
  XOR2_X1 U14648 ( .A(n14622), .B(n14623), .Z(n14620) );
  NOR2_X1 U14649 ( .A1(n14438), .A2(n10616), .ZN(n14623) );
  NAND2_X1 U14650 ( .A1(n14619), .A2(a_17_), .ZN(n14478) );
  NOR2_X1 U14651 ( .A1(n14624), .A2(n14625), .ZN(n14619) );
  INV_X1 U14652 ( .A(n14626), .ZN(n14625) );
  NAND2_X1 U14653 ( .A1(n14472), .A2(n14627), .ZN(n14626) );
  NAND2_X1 U14654 ( .A1(n14475), .A2(n14474), .ZN(n14627) );
  XNOR2_X1 U14655 ( .A(n14628), .B(n14629), .ZN(n14472) );
  XOR2_X1 U14656 ( .A(n14630), .B(n14631), .Z(n14628) );
  NOR2_X1 U14657 ( .A1(n8881), .A2(n14438), .ZN(n14631) );
  NOR2_X1 U14658 ( .A1(n14474), .A2(n14475), .ZN(n14624) );
  NOR2_X1 U14659 ( .A1(n10616), .A2(n14216), .ZN(n14475) );
  NAND2_X1 U14660 ( .A1(n14470), .A2(n14632), .ZN(n14474) );
  NAND2_X1 U14661 ( .A1(n14469), .A2(n14471), .ZN(n14632) );
  NAND2_X1 U14662 ( .A1(n14633), .A2(n14634), .ZN(n14471) );
  NAND2_X1 U14663 ( .A1(b_8_), .A2(a_19_), .ZN(n14634) );
  INV_X1 U14664 ( .A(n14635), .ZN(n14633) );
  XNOR2_X1 U14665 ( .A(n14636), .B(n14637), .ZN(n14469) );
  XOR2_X1 U14666 ( .A(n14638), .B(n14639), .Z(n14637) );
  NAND2_X1 U14667 ( .A1(b_7_), .A2(a_20_), .ZN(n14639) );
  NAND2_X1 U14668 ( .A1(a_19_), .A2(n14635), .ZN(n14470) );
  NAND2_X1 U14669 ( .A1(n14640), .A2(n14641), .ZN(n14635) );
  NAND2_X1 U14670 ( .A1(n14467), .A2(n14642), .ZN(n14641) );
  INV_X1 U14671 ( .A(n14643), .ZN(n14642) );
  NOR2_X1 U14672 ( .A1(n14465), .A2(n14466), .ZN(n14643) );
  NOR2_X1 U14673 ( .A1(n14216), .A2(n10633), .ZN(n14467) );
  NAND2_X1 U14674 ( .A1(n14465), .A2(n14466), .ZN(n14640) );
  NAND2_X1 U14675 ( .A1(n14644), .A2(n14645), .ZN(n14466) );
  NAND2_X1 U14676 ( .A1(n14463), .A2(n14646), .ZN(n14645) );
  NAND2_X1 U14677 ( .A1(n14647), .A2(n14648), .ZN(n14646) );
  INV_X1 U14678 ( .A(n14462), .ZN(n14648) );
  INV_X1 U14679 ( .A(n14461), .ZN(n14647) );
  NOR2_X1 U14680 ( .A1(n14216), .A2(n8798), .ZN(n14463) );
  NAND2_X1 U14681 ( .A1(n14461), .A2(n14462), .ZN(n14644) );
  NAND2_X1 U14682 ( .A1(n14649), .A2(n14650), .ZN(n14462) );
  INV_X1 U14683 ( .A(n14651), .ZN(n14650) );
  NOR2_X1 U14684 ( .A1(n14390), .A2(n14652), .ZN(n14651) );
  NOR2_X1 U14685 ( .A1(n14387), .A2(n14389), .ZN(n14652) );
  NAND2_X1 U14686 ( .A1(b_8_), .A2(a_22_), .ZN(n14390) );
  NAND2_X1 U14687 ( .A1(n14387), .A2(n14389), .ZN(n14649) );
  NAND2_X1 U14688 ( .A1(n14653), .A2(n14654), .ZN(n14389) );
  NAND2_X1 U14689 ( .A1(n14459), .A2(n14655), .ZN(n14654) );
  INV_X1 U14690 ( .A(n14656), .ZN(n14655) );
  NOR2_X1 U14691 ( .A1(n14457), .A2(n14458), .ZN(n14656) );
  NOR2_X1 U14692 ( .A1(n14216), .A2(n8812), .ZN(n14459) );
  NAND2_X1 U14693 ( .A1(n14457), .A2(n14458), .ZN(n14653) );
  NAND2_X1 U14694 ( .A1(n14657), .A2(n14658), .ZN(n14458) );
  NAND2_X1 U14695 ( .A1(n14455), .A2(n14659), .ZN(n14658) );
  INV_X1 U14696 ( .A(n14660), .ZN(n14659) );
  NOR2_X1 U14697 ( .A1(n14453), .A2(n14454), .ZN(n14660) );
  NOR2_X1 U14698 ( .A1(n14216), .A2(n9131), .ZN(n14455) );
  NAND2_X1 U14699 ( .A1(n14453), .A2(n14454), .ZN(n14657) );
  NAND2_X1 U14700 ( .A1(n14661), .A2(n14662), .ZN(n14454) );
  NAND2_X1 U14701 ( .A1(n14451), .A2(n14663), .ZN(n14662) );
  NAND2_X1 U14702 ( .A1(n14448), .A2(n14450), .ZN(n14663) );
  NOR2_X1 U14703 ( .A1(n14216), .A2(n8825), .ZN(n14451) );
  INV_X1 U14704 ( .A(n14664), .ZN(n14661) );
  NOR2_X1 U14705 ( .A1(n14450), .A2(n14448), .ZN(n14664) );
  XNOR2_X1 U14706 ( .A(n14665), .B(n14666), .ZN(n14448) );
  XNOR2_X1 U14707 ( .A(n14667), .B(n14668), .ZN(n14666) );
  NAND2_X1 U14708 ( .A1(n14669), .A2(n14670), .ZN(n14450) );
  NAND2_X1 U14709 ( .A1(n14407), .A2(n14671), .ZN(n14670) );
  NAND2_X1 U14710 ( .A1(n14410), .A2(n14409), .ZN(n14671) );
  XNOR2_X1 U14711 ( .A(n14672), .B(n14673), .ZN(n14407) );
  XOR2_X1 U14712 ( .A(n14674), .B(n14675), .Z(n14673) );
  INV_X1 U14713 ( .A(n14676), .ZN(n14669) );
  NOR2_X1 U14714 ( .A1(n14409), .A2(n14410), .ZN(n14676) );
  NOR2_X1 U14715 ( .A1(n8830), .A2(n14216), .ZN(n14410) );
  NAND2_X1 U14716 ( .A1(n14677), .A2(n14678), .ZN(n14409) );
  NAND2_X1 U14717 ( .A1(n14417), .A2(n14679), .ZN(n14678) );
  NAND2_X1 U14718 ( .A1(n14414), .A2(n14416), .ZN(n14679) );
  NOR2_X1 U14719 ( .A1(n14216), .A2(n8839), .ZN(n14417) );
  INV_X1 U14720 ( .A(n14680), .ZN(n14677) );
  NOR2_X1 U14721 ( .A1(n14414), .A2(n14416), .ZN(n14680) );
  NOR2_X1 U14722 ( .A1(n14681), .A2(n14682), .ZN(n14416) );
  INV_X1 U14723 ( .A(n14683), .ZN(n14682) );
  NAND2_X1 U14724 ( .A1(n14446), .A2(n14684), .ZN(n14683) );
  NAND2_X1 U14725 ( .A1(n14447), .A2(n14445), .ZN(n14684) );
  NOR2_X1 U14726 ( .A1(n14216), .A2(n8844), .ZN(n14446) );
  NOR2_X1 U14727 ( .A1(n14445), .A2(n14447), .ZN(n14681) );
  NOR2_X1 U14728 ( .A1(n14685), .A2(n14686), .ZN(n14447) );
  INV_X1 U14729 ( .A(n14687), .ZN(n14686) );
  NAND2_X1 U14730 ( .A1(n14440), .A2(n14688), .ZN(n14687) );
  NAND2_X1 U14731 ( .A1(n14689), .A2(n14442), .ZN(n14688) );
  NOR2_X1 U14732 ( .A1(n14216), .A2(n9161), .ZN(n14440) );
  NOR2_X1 U14733 ( .A1(n14442), .A2(n14689), .ZN(n14685) );
  INV_X1 U14734 ( .A(n14443), .ZN(n14689) );
  NAND2_X1 U14735 ( .A1(n14690), .A2(n14691), .ZN(n14443) );
  NAND2_X1 U14736 ( .A1(b_6_), .A2(n14692), .ZN(n14691) );
  NAND2_X1 U14737 ( .A1(n8358), .A2(n14693), .ZN(n14692) );
  NAND2_X1 U14738 ( .A1(a_31_), .A2(n14438), .ZN(n14693) );
  NAND2_X1 U14739 ( .A1(b_7_), .A2(n14694), .ZN(n14690) );
  NAND2_X1 U14740 ( .A1(n8362), .A2(n14695), .ZN(n14694) );
  NAND2_X1 U14741 ( .A1(a_30_), .A2(n14696), .ZN(n14695) );
  NAND2_X1 U14742 ( .A1(n14697), .A2(b_7_), .ZN(n14442) );
  NOR2_X1 U14743 ( .A1(n9170), .A2(n14216), .ZN(n14697) );
  XOR2_X1 U14744 ( .A(n14698), .B(n14699), .Z(n14445) );
  XOR2_X1 U14745 ( .A(n14700), .B(n14701), .Z(n14699) );
  XOR2_X1 U14746 ( .A(n14702), .B(n14703), .Z(n14414) );
  XNOR2_X1 U14747 ( .A(n14704), .B(n14705), .ZN(n14702) );
  XNOR2_X1 U14748 ( .A(n14706), .B(n14707), .ZN(n14453) );
  XNOR2_X1 U14749 ( .A(n14708), .B(n14709), .ZN(n14707) );
  XNOR2_X1 U14750 ( .A(n14710), .B(n14711), .ZN(n14457) );
  XNOR2_X1 U14751 ( .A(n14712), .B(n14713), .ZN(n14710) );
  XNOR2_X1 U14752 ( .A(n14714), .B(n14715), .ZN(n14387) );
  XNOR2_X1 U14753 ( .A(n14716), .B(n14717), .ZN(n14714) );
  XNOR2_X1 U14754 ( .A(n14718), .B(n14719), .ZN(n14461) );
  NAND2_X1 U14755 ( .A1(n14720), .A2(n14721), .ZN(n14718) );
  XNOR2_X1 U14756 ( .A(n14722), .B(n14723), .ZN(n14465) );
  NAND2_X1 U14757 ( .A1(n14724), .A2(n14725), .ZN(n14722) );
  XOR2_X1 U14758 ( .A(n14726), .B(n14727), .Z(n14488) );
  XOR2_X1 U14759 ( .A(n14728), .B(n14729), .Z(n14726) );
  NOR2_X1 U14760 ( .A1(n14438), .A2(n8438), .ZN(n14729) );
  XOR2_X1 U14761 ( .A(n14730), .B(n14731), .Z(n14492) );
  XOR2_X1 U14762 ( .A(n14732), .B(n14733), .Z(n14730) );
  NOR2_X1 U14763 ( .A1(n14438), .A2(n8443), .ZN(n14733) );
  XOR2_X1 U14764 ( .A(n14734), .B(n14735), .Z(n14496) );
  XOR2_X1 U14765 ( .A(n14736), .B(n14737), .Z(n14734) );
  NOR2_X1 U14766 ( .A1(n14438), .A2(n8750), .ZN(n14737) );
  XOR2_X1 U14767 ( .A(n14738), .B(n14739), .Z(n14331) );
  XOR2_X1 U14768 ( .A(n14740), .B(n14741), .Z(n14738) );
  NOR2_X1 U14769 ( .A1(n14438), .A2(n8452), .ZN(n14741) );
  XNOR2_X1 U14770 ( .A(n14742), .B(n14743), .ZN(n14322) );
  XOR2_X1 U14771 ( .A(n14744), .B(n14745), .Z(n14743) );
  NAND2_X1 U14772 ( .A1(a_10_), .A2(b_7_), .ZN(n14745) );
  XNOR2_X1 U14773 ( .A(n14746), .B(n14747), .ZN(n14500) );
  XOR2_X1 U14774 ( .A(n14748), .B(n14749), .Z(n14747) );
  NAND2_X1 U14775 ( .A1(a_9_), .A2(b_7_), .ZN(n14749) );
  XOR2_X1 U14776 ( .A(n14750), .B(n14751), .Z(n14505) );
  XOR2_X1 U14777 ( .A(n14752), .B(n14753), .Z(n14751) );
  NAND2_X1 U14778 ( .A1(a_8_), .A2(b_7_), .ZN(n14753) );
  XOR2_X1 U14779 ( .A(n14754), .B(n14755), .Z(n14508) );
  XOR2_X1 U14780 ( .A(n14756), .B(n14757), .Z(n14755) );
  XNOR2_X1 U14781 ( .A(n14758), .B(n14759), .ZN(n14513) );
  XNOR2_X1 U14782 ( .A(n14760), .B(n14761), .ZN(n14759) );
  XNOR2_X1 U14783 ( .A(n14762), .B(n14763), .ZN(n14517) );
  XNOR2_X1 U14784 ( .A(n14764), .B(n14765), .ZN(n14762) );
  XNOR2_X1 U14785 ( .A(n14766), .B(n14767), .ZN(n14520) );
  XNOR2_X1 U14786 ( .A(n14768), .B(n14769), .ZN(n14766) );
  XNOR2_X1 U14787 ( .A(n14770), .B(n14771), .ZN(n14525) );
  XNOR2_X1 U14788 ( .A(n14772), .B(n14773), .ZN(n14770) );
  XNOR2_X1 U14789 ( .A(n14774), .B(n14775), .ZN(n14529) );
  XNOR2_X1 U14790 ( .A(n14776), .B(n14777), .ZN(n14774) );
  XNOR2_X1 U14791 ( .A(n14778), .B(n14779), .ZN(n14283) );
  XNOR2_X1 U14792 ( .A(n14780), .B(n14781), .ZN(n14778) );
  XOR2_X1 U14793 ( .A(n14782), .B(n14783), .Z(n14533) );
  XOR2_X1 U14794 ( .A(n14784), .B(n14785), .Z(n14783) );
  NOR2_X1 U14795 ( .A1(n14786), .A2(n8618), .ZN(n8351) );
  INV_X1 U14796 ( .A(n14787), .ZN(n8618) );
  NAND2_X1 U14797 ( .A1(n14788), .A2(n14789), .ZN(n14787) );
  NOR2_X1 U14798 ( .A1(n14789), .A2(n14788), .ZN(n14786) );
  XNOR2_X1 U14799 ( .A(n14790), .B(n14791), .ZN(n14788) );
  XNOR2_X1 U14800 ( .A(n14792), .B(n14793), .ZN(n14791) );
  NAND2_X1 U14801 ( .A1(n14794), .A2(n14795), .ZN(n14789) );
  NAND2_X1 U14802 ( .A1(n14785), .A2(n14796), .ZN(n14795) );
  NAND2_X1 U14803 ( .A1(n14784), .A2(n14782), .ZN(n14796) );
  INV_X1 U14804 ( .A(n14797), .ZN(n14782) );
  INV_X1 U14805 ( .A(n14798), .ZN(n14784) );
  NOR2_X1 U14806 ( .A1(n8690), .A2(n14438), .ZN(n14785) );
  NAND2_X1 U14807 ( .A1(n14797), .A2(n14798), .ZN(n14794) );
  NAND2_X1 U14808 ( .A1(n14799), .A2(n14800), .ZN(n14798) );
  NAND2_X1 U14809 ( .A1(n14780), .A2(n14801), .ZN(n14800) );
  NAND2_X1 U14810 ( .A1(n14781), .A2(n14779), .ZN(n14801) );
  NOR2_X1 U14811 ( .A1(n8502), .A2(n14438), .ZN(n14780) );
  INV_X1 U14812 ( .A(n14802), .ZN(n14799) );
  NOR2_X1 U14813 ( .A1(n14779), .A2(n14781), .ZN(n14802) );
  NOR2_X1 U14814 ( .A1(n14803), .A2(n14804), .ZN(n14781) );
  INV_X1 U14815 ( .A(n14805), .ZN(n14804) );
  NAND2_X1 U14816 ( .A1(n14776), .A2(n14806), .ZN(n14805) );
  NAND2_X1 U14817 ( .A1(n14777), .A2(n14775), .ZN(n14806) );
  NOR2_X1 U14818 ( .A1(n8497), .A2(n14438), .ZN(n14776) );
  NOR2_X1 U14819 ( .A1(n14775), .A2(n14777), .ZN(n14803) );
  NOR2_X1 U14820 ( .A1(n14807), .A2(n14808), .ZN(n14777) );
  INV_X1 U14821 ( .A(n14809), .ZN(n14808) );
  NAND2_X1 U14822 ( .A1(n14773), .A2(n14810), .ZN(n14809) );
  NAND2_X1 U14823 ( .A1(n14772), .A2(n14771), .ZN(n14810) );
  NOR2_X1 U14824 ( .A1(n8707), .A2(n14438), .ZN(n14773) );
  NOR2_X1 U14825 ( .A1(n14771), .A2(n14772), .ZN(n14807) );
  NOR2_X1 U14826 ( .A1(n14811), .A2(n14812), .ZN(n14772) );
  INV_X1 U14827 ( .A(n14813), .ZN(n14812) );
  NAND2_X1 U14828 ( .A1(n14768), .A2(n14814), .ZN(n14813) );
  NAND2_X1 U14829 ( .A1(n14769), .A2(n14767), .ZN(n14814) );
  NOR2_X1 U14830 ( .A1(n8712), .A2(n14438), .ZN(n14768) );
  NOR2_X1 U14831 ( .A1(n14767), .A2(n14769), .ZN(n14811) );
  NOR2_X1 U14832 ( .A1(n14815), .A2(n14816), .ZN(n14769) );
  INV_X1 U14833 ( .A(n14817), .ZN(n14816) );
  NAND2_X1 U14834 ( .A1(n14765), .A2(n14818), .ZN(n14817) );
  NAND2_X1 U14835 ( .A1(n14764), .A2(n14763), .ZN(n14818) );
  NOR2_X1 U14836 ( .A1(n8717), .A2(n14438), .ZN(n14765) );
  NOR2_X1 U14837 ( .A1(n14763), .A2(n14764), .ZN(n14815) );
  NOR2_X1 U14838 ( .A1(n14819), .A2(n14820), .ZN(n14764) );
  INV_X1 U14839 ( .A(n14821), .ZN(n14820) );
  NAND2_X1 U14840 ( .A1(n14761), .A2(n14822), .ZN(n14821) );
  NAND2_X1 U14841 ( .A1(n14758), .A2(n14760), .ZN(n14822) );
  NOR2_X1 U14842 ( .A1(n8480), .A2(n14438), .ZN(n14761) );
  NOR2_X1 U14843 ( .A1(n14760), .A2(n14758), .ZN(n14819) );
  XOR2_X1 U14844 ( .A(n14823), .B(n14824), .Z(n14758) );
  XOR2_X1 U14845 ( .A(n14825), .B(n14826), .Z(n14824) );
  NAND2_X1 U14846 ( .A1(n14827), .A2(n14828), .ZN(n14760) );
  NAND2_X1 U14847 ( .A1(n14754), .A2(n14829), .ZN(n14828) );
  NAND2_X1 U14848 ( .A1(n14830), .A2(n14756), .ZN(n14829) );
  XNOR2_X1 U14849 ( .A(n14831), .B(n14832), .ZN(n14754) );
  XOR2_X1 U14850 ( .A(n14833), .B(n14834), .Z(n14832) );
  NAND2_X1 U14851 ( .A1(n14835), .A2(n14757), .ZN(n14827) );
  INV_X1 U14852 ( .A(n14756), .ZN(n14835) );
  NAND2_X1 U14853 ( .A1(n14836), .A2(n14837), .ZN(n14756) );
  NAND2_X1 U14854 ( .A1(n14838), .A2(a_8_), .ZN(n14837) );
  NOR2_X1 U14855 ( .A1(n14839), .A2(n14438), .ZN(n14838) );
  NOR2_X1 U14856 ( .A1(n14752), .A2(n14750), .ZN(n14839) );
  NAND2_X1 U14857 ( .A1(n14750), .A2(n14752), .ZN(n14836) );
  NAND2_X1 U14858 ( .A1(n14840), .A2(n14841), .ZN(n14752) );
  NAND2_X1 U14859 ( .A1(n14842), .A2(a_9_), .ZN(n14841) );
  NOR2_X1 U14860 ( .A1(n14843), .A2(n14438), .ZN(n14842) );
  NOR2_X1 U14861 ( .A1(n14746), .A2(n14748), .ZN(n14843) );
  NAND2_X1 U14862 ( .A1(n14746), .A2(n14748), .ZN(n14840) );
  NAND2_X1 U14863 ( .A1(n14844), .A2(n14845), .ZN(n14748) );
  NAND2_X1 U14864 ( .A1(n14846), .A2(a_10_), .ZN(n14845) );
  NOR2_X1 U14865 ( .A1(n14847), .A2(n14438), .ZN(n14846) );
  NOR2_X1 U14866 ( .A1(n14744), .A2(n14742), .ZN(n14847) );
  NAND2_X1 U14867 ( .A1(n14742), .A2(n14744), .ZN(n14844) );
  NAND2_X1 U14868 ( .A1(n14848), .A2(n14849), .ZN(n14744) );
  NAND2_X1 U14869 ( .A1(n14850), .A2(a_11_), .ZN(n14849) );
  NOR2_X1 U14870 ( .A1(n14851), .A2(n14438), .ZN(n14850) );
  NOR2_X1 U14871 ( .A1(n14740), .A2(n14739), .ZN(n14851) );
  NAND2_X1 U14872 ( .A1(n14739), .A2(n14740), .ZN(n14848) );
  NAND2_X1 U14873 ( .A1(n14852), .A2(n14853), .ZN(n14740) );
  NAND2_X1 U14874 ( .A1(n14854), .A2(a_12_), .ZN(n14853) );
  NOR2_X1 U14875 ( .A1(n14855), .A2(n14438), .ZN(n14854) );
  NOR2_X1 U14876 ( .A1(n14736), .A2(n14735), .ZN(n14855) );
  NAND2_X1 U14877 ( .A1(n14735), .A2(n14736), .ZN(n14852) );
  NAND2_X1 U14878 ( .A1(n14856), .A2(n14857), .ZN(n14736) );
  NAND2_X1 U14879 ( .A1(n14858), .A2(a_13_), .ZN(n14857) );
  NOR2_X1 U14880 ( .A1(n14859), .A2(n14438), .ZN(n14858) );
  NOR2_X1 U14881 ( .A1(n14731), .A2(n14732), .ZN(n14859) );
  NAND2_X1 U14882 ( .A1(n14731), .A2(n14732), .ZN(n14856) );
  NAND2_X1 U14883 ( .A1(n14860), .A2(n14861), .ZN(n14732) );
  NAND2_X1 U14884 ( .A1(n14862), .A2(a_14_), .ZN(n14861) );
  NOR2_X1 U14885 ( .A1(n14863), .A2(n14438), .ZN(n14862) );
  NOR2_X1 U14886 ( .A1(n14728), .A2(n14727), .ZN(n14863) );
  NAND2_X1 U14887 ( .A1(n14727), .A2(n14728), .ZN(n14860) );
  NAND2_X1 U14888 ( .A1(n14864), .A2(n14865), .ZN(n14728) );
  NAND2_X1 U14889 ( .A1(n14866), .A2(a_15_), .ZN(n14865) );
  NOR2_X1 U14890 ( .A1(n14867), .A2(n14438), .ZN(n14866) );
  NOR2_X1 U14891 ( .A1(n14597), .A2(n14598), .ZN(n14867) );
  NAND2_X1 U14892 ( .A1(n14597), .A2(n14598), .ZN(n14864) );
  NAND2_X1 U14893 ( .A1(n14868), .A2(n14869), .ZN(n14598) );
  NAND2_X1 U14894 ( .A1(n14870), .A2(a_16_), .ZN(n14869) );
  NOR2_X1 U14895 ( .A1(n14871), .A2(n14438), .ZN(n14870) );
  NOR2_X1 U14896 ( .A1(n14606), .A2(n14605), .ZN(n14871) );
  NAND2_X1 U14897 ( .A1(n14605), .A2(n14606), .ZN(n14868) );
  NAND2_X1 U14898 ( .A1(n14872), .A2(n14873), .ZN(n14606) );
  NAND2_X1 U14899 ( .A1(n14874), .A2(a_17_), .ZN(n14873) );
  NOR2_X1 U14900 ( .A1(n14875), .A2(n14438), .ZN(n14874) );
  NOR2_X1 U14901 ( .A1(n14614), .A2(n14613), .ZN(n14875) );
  NAND2_X1 U14902 ( .A1(n14613), .A2(n14614), .ZN(n14872) );
  NAND2_X1 U14903 ( .A1(n14876), .A2(n14877), .ZN(n14614) );
  NAND2_X1 U14904 ( .A1(n14878), .A2(a_18_), .ZN(n14877) );
  NOR2_X1 U14905 ( .A1(n14879), .A2(n14438), .ZN(n14878) );
  NOR2_X1 U14906 ( .A1(n14622), .A2(n14621), .ZN(n14879) );
  NAND2_X1 U14907 ( .A1(n14621), .A2(n14622), .ZN(n14876) );
  NAND2_X1 U14908 ( .A1(n14880), .A2(n14881), .ZN(n14622) );
  NAND2_X1 U14909 ( .A1(n14882), .A2(b_7_), .ZN(n14881) );
  NOR2_X1 U14910 ( .A1(n14883), .A2(n8881), .ZN(n14882) );
  NOR2_X1 U14911 ( .A1(n14629), .A2(n14630), .ZN(n14883) );
  NAND2_X1 U14912 ( .A1(n14629), .A2(n14630), .ZN(n14880) );
  NAND2_X1 U14913 ( .A1(n14884), .A2(n14885), .ZN(n14630) );
  NAND2_X1 U14914 ( .A1(n14886), .A2(b_7_), .ZN(n14885) );
  NOR2_X1 U14915 ( .A1(n14887), .A2(n10633), .ZN(n14886) );
  NOR2_X1 U14916 ( .A1(n14636), .A2(n14638), .ZN(n14887) );
  NAND2_X1 U14917 ( .A1(n14636), .A2(n14638), .ZN(n14884) );
  NAND2_X1 U14918 ( .A1(n14724), .A2(n14888), .ZN(n14638) );
  NAND2_X1 U14919 ( .A1(n14723), .A2(n14725), .ZN(n14888) );
  NAND2_X1 U14920 ( .A1(n14889), .A2(n14890), .ZN(n14725) );
  NAND2_X1 U14921 ( .A1(b_7_), .A2(a_21_), .ZN(n14890) );
  INV_X1 U14922 ( .A(n14891), .ZN(n14889) );
  XNOR2_X1 U14923 ( .A(n14892), .B(n14893), .ZN(n14723) );
  NAND2_X1 U14924 ( .A1(n14894), .A2(n14895), .ZN(n14892) );
  NAND2_X1 U14925 ( .A1(a_21_), .A2(n14891), .ZN(n14724) );
  NAND2_X1 U14926 ( .A1(n14720), .A2(n14896), .ZN(n14891) );
  NAND2_X1 U14927 ( .A1(n14719), .A2(n14721), .ZN(n14896) );
  NAND2_X1 U14928 ( .A1(n14897), .A2(n14898), .ZN(n14721) );
  NAND2_X1 U14929 ( .A1(b_7_), .A2(a_22_), .ZN(n14898) );
  XNOR2_X1 U14930 ( .A(n14899), .B(n14900), .ZN(n14719) );
  XOR2_X1 U14931 ( .A(n14901), .B(n14902), .Z(n14900) );
  NAND2_X1 U14932 ( .A1(b_6_), .A2(a_23_), .ZN(n14902) );
  INV_X1 U14933 ( .A(n14903), .ZN(n14720) );
  NOR2_X1 U14934 ( .A1(n8803), .A2(n14897), .ZN(n14903) );
  NOR2_X1 U14935 ( .A1(n14904), .A2(n14905), .ZN(n14897) );
  INV_X1 U14936 ( .A(n14906), .ZN(n14905) );
  NAND2_X1 U14937 ( .A1(n14717), .A2(n14907), .ZN(n14906) );
  NAND2_X1 U14938 ( .A1(n14716), .A2(n14715), .ZN(n14907) );
  NOR2_X1 U14939 ( .A1(n14438), .A2(n8812), .ZN(n14717) );
  NOR2_X1 U14940 ( .A1(n14715), .A2(n14716), .ZN(n14904) );
  NOR2_X1 U14941 ( .A1(n14908), .A2(n14909), .ZN(n14716) );
  INV_X1 U14942 ( .A(n14910), .ZN(n14909) );
  NAND2_X1 U14943 ( .A1(n14713), .A2(n14911), .ZN(n14910) );
  NAND2_X1 U14944 ( .A1(n14712), .A2(n14711), .ZN(n14911) );
  NOR2_X1 U14945 ( .A1(n14438), .A2(n9131), .ZN(n14713) );
  NOR2_X1 U14946 ( .A1(n14711), .A2(n14712), .ZN(n14908) );
  NOR2_X1 U14947 ( .A1(n14912), .A2(n14913), .ZN(n14712) );
  INV_X1 U14948 ( .A(n14914), .ZN(n14913) );
  NAND2_X1 U14949 ( .A1(n14709), .A2(n14915), .ZN(n14914) );
  NAND2_X1 U14950 ( .A1(n14706), .A2(n14708), .ZN(n14915) );
  NOR2_X1 U14951 ( .A1(n14438), .A2(n8825), .ZN(n14709) );
  NOR2_X1 U14952 ( .A1(n14708), .A2(n14706), .ZN(n14912) );
  XNOR2_X1 U14953 ( .A(n14916), .B(n14917), .ZN(n14706) );
  XNOR2_X1 U14954 ( .A(n14918), .B(n14919), .ZN(n14917) );
  NAND2_X1 U14955 ( .A1(n14920), .A2(n14921), .ZN(n14708) );
  NAND2_X1 U14956 ( .A1(n14665), .A2(n14922), .ZN(n14921) );
  NAND2_X1 U14957 ( .A1(n14668), .A2(n14667), .ZN(n14922) );
  XNOR2_X1 U14958 ( .A(n14923), .B(n14924), .ZN(n14665) );
  XOR2_X1 U14959 ( .A(n14925), .B(n14926), .Z(n14924) );
  INV_X1 U14960 ( .A(n14927), .ZN(n14920) );
  NOR2_X1 U14961 ( .A1(n14667), .A2(n14668), .ZN(n14927) );
  NOR2_X1 U14962 ( .A1(n8830), .A2(n14438), .ZN(n14668) );
  NAND2_X1 U14963 ( .A1(n14928), .A2(n14929), .ZN(n14667) );
  NAND2_X1 U14964 ( .A1(n14675), .A2(n14930), .ZN(n14929) );
  NAND2_X1 U14965 ( .A1(n14672), .A2(n14674), .ZN(n14930) );
  NOR2_X1 U14966 ( .A1(n14438), .A2(n8839), .ZN(n14675) );
  INV_X1 U14967 ( .A(n14931), .ZN(n14928) );
  NOR2_X1 U14968 ( .A1(n14672), .A2(n14674), .ZN(n14931) );
  NOR2_X1 U14969 ( .A1(n14932), .A2(n14933), .ZN(n14674) );
  INV_X1 U14970 ( .A(n14934), .ZN(n14933) );
  NAND2_X1 U14971 ( .A1(n14704), .A2(n14935), .ZN(n14934) );
  NAND2_X1 U14972 ( .A1(n14705), .A2(n14703), .ZN(n14935) );
  NOR2_X1 U14973 ( .A1(n14438), .A2(n8844), .ZN(n14704) );
  NOR2_X1 U14974 ( .A1(n14703), .A2(n14705), .ZN(n14932) );
  NOR2_X1 U14975 ( .A1(n14936), .A2(n14937), .ZN(n14705) );
  INV_X1 U14976 ( .A(n14938), .ZN(n14937) );
  NAND2_X1 U14977 ( .A1(n14698), .A2(n14939), .ZN(n14938) );
  NAND2_X1 U14978 ( .A1(n14940), .A2(n14700), .ZN(n14939) );
  NOR2_X1 U14979 ( .A1(n14438), .A2(n9161), .ZN(n14698) );
  NOR2_X1 U14980 ( .A1(n14700), .A2(n14940), .ZN(n14936) );
  INV_X1 U14981 ( .A(n14701), .ZN(n14940) );
  NAND2_X1 U14982 ( .A1(n14941), .A2(n14942), .ZN(n14701) );
  NAND2_X1 U14983 ( .A1(b_5_), .A2(n14943), .ZN(n14942) );
  NAND2_X1 U14984 ( .A1(n8358), .A2(n14944), .ZN(n14943) );
  NAND2_X1 U14985 ( .A1(a_31_), .A2(n14696), .ZN(n14944) );
  NAND2_X1 U14986 ( .A1(b_6_), .A2(n14945), .ZN(n14941) );
  NAND2_X1 U14987 ( .A1(n8362), .A2(n14946), .ZN(n14945) );
  NAND2_X1 U14988 ( .A1(a_30_), .A2(n14947), .ZN(n14946) );
  NAND2_X1 U14989 ( .A1(n14948), .A2(b_6_), .ZN(n14700) );
  NOR2_X1 U14990 ( .A1(n9170), .A2(n14438), .ZN(n14948) );
  XOR2_X1 U14991 ( .A(n14949), .B(n14950), .Z(n14703) );
  XOR2_X1 U14992 ( .A(n14951), .B(n14952), .Z(n14950) );
  XOR2_X1 U14993 ( .A(n14953), .B(n14954), .Z(n14672) );
  XNOR2_X1 U14994 ( .A(n14955), .B(n14956), .ZN(n14953) );
  XNOR2_X1 U14995 ( .A(n14957), .B(n14958), .ZN(n14711) );
  XOR2_X1 U14996 ( .A(n14959), .B(n14960), .Z(n14958) );
  XNOR2_X1 U14997 ( .A(n14961), .B(n14962), .ZN(n14715) );
  XOR2_X1 U14998 ( .A(n14963), .B(n14964), .Z(n14961) );
  NOR2_X1 U14999 ( .A1(n9131), .A2(n14696), .ZN(n14964) );
  XNOR2_X1 U15000 ( .A(n14965), .B(n14966), .ZN(n14636) );
  XOR2_X1 U15001 ( .A(n14967), .B(n14968), .Z(n14965) );
  XNOR2_X1 U15002 ( .A(n14969), .B(n14970), .ZN(n14629) );
  NAND2_X1 U15003 ( .A1(n14971), .A2(n14972), .ZN(n14969) );
  XOR2_X1 U15004 ( .A(n14973), .B(n14974), .Z(n14621) );
  XNOR2_X1 U15005 ( .A(n14975), .B(n14976), .ZN(n14974) );
  XNOR2_X1 U15006 ( .A(n14977), .B(n14978), .ZN(n14613) );
  XNOR2_X1 U15007 ( .A(n14979), .B(n14980), .ZN(n14978) );
  XNOR2_X1 U15008 ( .A(n14981), .B(n14982), .ZN(n14605) );
  XNOR2_X1 U15009 ( .A(n14983), .B(n14984), .ZN(n14981) );
  XNOR2_X1 U15010 ( .A(n14985), .B(n14986), .ZN(n14597) );
  XNOR2_X1 U15011 ( .A(n14987), .B(n14988), .ZN(n14986) );
  XNOR2_X1 U15012 ( .A(n14989), .B(n14990), .ZN(n14727) );
  XOR2_X1 U15013 ( .A(n14991), .B(n14992), .Z(n14990) );
  XNOR2_X1 U15014 ( .A(n14993), .B(n14994), .ZN(n14731) );
  XNOR2_X1 U15015 ( .A(n14995), .B(n14996), .ZN(n14994) );
  XNOR2_X1 U15016 ( .A(n14997), .B(n14998), .ZN(n14735) );
  XOR2_X1 U15017 ( .A(n14999), .B(n15000), .Z(n14998) );
  XNOR2_X1 U15018 ( .A(n15001), .B(n15002), .ZN(n14739) );
  XNOR2_X1 U15019 ( .A(n15003), .B(n15004), .ZN(n15002) );
  XNOR2_X1 U15020 ( .A(n15005), .B(n15006), .ZN(n14742) );
  XOR2_X1 U15021 ( .A(n15007), .B(n15008), .Z(n15006) );
  XOR2_X1 U15022 ( .A(n15009), .B(n15010), .Z(n14746) );
  XOR2_X1 U15023 ( .A(n15011), .B(n15012), .Z(n15010) );
  XNOR2_X1 U15024 ( .A(n15013), .B(n15014), .ZN(n14750) );
  XOR2_X1 U15025 ( .A(n15015), .B(n15016), .Z(n15014) );
  XOR2_X1 U15026 ( .A(n15017), .B(n15018), .Z(n14763) );
  XOR2_X1 U15027 ( .A(n15019), .B(n15020), .Z(n15018) );
  XOR2_X1 U15028 ( .A(n15021), .B(n15022), .Z(n14767) );
  XNOR2_X1 U15029 ( .A(n15023), .B(n15024), .ZN(n15022) );
  XOR2_X1 U15030 ( .A(n15025), .B(n15026), .Z(n14771) );
  XNOR2_X1 U15031 ( .A(n15027), .B(n15028), .ZN(n15026) );
  XNOR2_X1 U15032 ( .A(n15029), .B(n15030), .ZN(n14775) );
  XOR2_X1 U15033 ( .A(n15031), .B(n15032), .Z(n15029) );
  XNOR2_X1 U15034 ( .A(n15033), .B(n15034), .ZN(n14779) );
  XOR2_X1 U15035 ( .A(n15035), .B(n15036), .Z(n15033) );
  XOR2_X1 U15036 ( .A(n15037), .B(n15038), .Z(n14797) );
  XOR2_X1 U15037 ( .A(n15039), .B(n15040), .Z(n15037) );
  XNOR2_X1 U15038 ( .A(n15041), .B(n15042), .ZN(n8354) );
  NAND2_X1 U15039 ( .A1(n8378), .A2(n8379), .ZN(n8377) );
  NOR2_X1 U15040 ( .A1(n15041), .A2(n15042), .ZN(n8379) );
  INV_X1 U15041 ( .A(n15043), .ZN(n15042) );
  NAND2_X1 U15042 ( .A1(n15044), .A2(n15045), .ZN(n15043) );
  NAND2_X1 U15043 ( .A1(n14793), .A2(n15046), .ZN(n15045) );
  INV_X1 U15044 ( .A(n15047), .ZN(n15046) );
  NOR2_X1 U15045 ( .A1(n14792), .A2(n14790), .ZN(n15047) );
  NOR2_X1 U15046 ( .A1(n8690), .A2(n14696), .ZN(n14793) );
  NAND2_X1 U15047 ( .A1(n14790), .A2(n14792), .ZN(n15044) );
  NAND2_X1 U15048 ( .A1(n15048), .A2(n15049), .ZN(n14792) );
  NAND2_X1 U15049 ( .A1(n15039), .A2(n15050), .ZN(n15049) );
  INV_X1 U15050 ( .A(n15051), .ZN(n15050) );
  NOR2_X1 U15051 ( .A1(n15038), .A2(n15040), .ZN(n15051) );
  NOR2_X1 U15052 ( .A1(n8502), .A2(n14696), .ZN(n15039) );
  NAND2_X1 U15053 ( .A1(n15038), .A2(n15040), .ZN(n15048) );
  NAND2_X1 U15054 ( .A1(n15052), .A2(n15053), .ZN(n15040) );
  NAND2_X1 U15055 ( .A1(n15036), .A2(n15054), .ZN(n15053) );
  INV_X1 U15056 ( .A(n15055), .ZN(n15054) );
  NOR2_X1 U15057 ( .A1(n15034), .A2(n15035), .ZN(n15055) );
  NOR2_X1 U15058 ( .A1(n8497), .A2(n14696), .ZN(n15036) );
  NAND2_X1 U15059 ( .A1(n15034), .A2(n15035), .ZN(n15052) );
  NAND2_X1 U15060 ( .A1(n15056), .A2(n15057), .ZN(n15035) );
  NAND2_X1 U15061 ( .A1(n15032), .A2(n15058), .ZN(n15057) );
  INV_X1 U15062 ( .A(n15059), .ZN(n15058) );
  NOR2_X1 U15063 ( .A1(n15030), .A2(n15031), .ZN(n15059) );
  NOR2_X1 U15064 ( .A1(n8707), .A2(n14696), .ZN(n15032) );
  NAND2_X1 U15065 ( .A1(n15030), .A2(n15031), .ZN(n15056) );
  NAND2_X1 U15066 ( .A1(n15060), .A2(n15061), .ZN(n15031) );
  NAND2_X1 U15067 ( .A1(n15028), .A2(n15062), .ZN(n15061) );
  INV_X1 U15068 ( .A(n15063), .ZN(n15062) );
  NOR2_X1 U15069 ( .A1(n15025), .A2(n15027), .ZN(n15063) );
  NOR2_X1 U15070 ( .A1(n8712), .A2(n14696), .ZN(n15028) );
  NAND2_X1 U15071 ( .A1(n15025), .A2(n15027), .ZN(n15060) );
  NAND2_X1 U15072 ( .A1(n15064), .A2(n15065), .ZN(n15027) );
  NAND2_X1 U15073 ( .A1(n15024), .A2(n15066), .ZN(n15065) );
  NAND2_X1 U15074 ( .A1(n15021), .A2(n15023), .ZN(n15066) );
  NOR2_X1 U15075 ( .A1(n8717), .A2(n14696), .ZN(n15024) );
  INV_X1 U15076 ( .A(n15067), .ZN(n15064) );
  NOR2_X1 U15077 ( .A1(n15021), .A2(n15023), .ZN(n15067) );
  NAND2_X1 U15078 ( .A1(n15068), .A2(n15069), .ZN(n15023) );
  NAND2_X1 U15079 ( .A1(n15070), .A2(n15020), .ZN(n15069) );
  NAND2_X1 U15080 ( .A1(n15017), .A2(n15019), .ZN(n15070) );
  INV_X1 U15081 ( .A(n15071), .ZN(n15068) );
  NOR2_X1 U15082 ( .A1(n15017), .A2(n15019), .ZN(n15071) );
  NAND2_X1 U15083 ( .A1(n15072), .A2(n15073), .ZN(n15019) );
  INV_X1 U15084 ( .A(n15074), .ZN(n15073) );
  NOR2_X1 U15085 ( .A1(n14826), .A2(n15075), .ZN(n15074) );
  NOR2_X1 U15086 ( .A1(n14825), .A2(n14823), .ZN(n15075) );
  NAND2_X1 U15087 ( .A1(a_7_), .A2(b_6_), .ZN(n14826) );
  NAND2_X1 U15088 ( .A1(n14823), .A2(n14825), .ZN(n15072) );
  NAND2_X1 U15089 ( .A1(n15076), .A2(n15077), .ZN(n14825) );
  NAND2_X1 U15090 ( .A1(n14834), .A2(n15078), .ZN(n15077) );
  NAND2_X1 U15091 ( .A1(n14831), .A2(n14833), .ZN(n15078) );
  NOR2_X1 U15092 ( .A1(n8731), .A2(n14696), .ZN(n14834) );
  NAND2_X1 U15093 ( .A1(n15079), .A2(n15080), .ZN(n15076) );
  INV_X1 U15094 ( .A(n14833), .ZN(n15080) );
  NOR2_X1 U15095 ( .A1(n15081), .A2(n15082), .ZN(n14833) );
  NOR2_X1 U15096 ( .A1(n15016), .A2(n15083), .ZN(n15082) );
  NOR2_X1 U15097 ( .A1(n15015), .A2(n15013), .ZN(n15083) );
  NAND2_X1 U15098 ( .A1(a_9_), .A2(b_6_), .ZN(n15016) );
  INV_X1 U15099 ( .A(n15084), .ZN(n15081) );
  NAND2_X1 U15100 ( .A1(n15013), .A2(n15015), .ZN(n15084) );
  NAND2_X1 U15101 ( .A1(n15085), .A2(n15086), .ZN(n15015) );
  NAND2_X1 U15102 ( .A1(n15012), .A2(n15087), .ZN(n15086) );
  NAND2_X1 U15103 ( .A1(n15009), .A2(n15011), .ZN(n15087) );
  NOR2_X1 U15104 ( .A1(n8741), .A2(n14696), .ZN(n15012) );
  NAND2_X1 U15105 ( .A1(n15088), .A2(n15089), .ZN(n15085) );
  INV_X1 U15106 ( .A(n15011), .ZN(n15089) );
  NOR2_X1 U15107 ( .A1(n15090), .A2(n15091), .ZN(n15011) );
  NOR2_X1 U15108 ( .A1(n15008), .A2(n15092), .ZN(n15091) );
  NOR2_X1 U15109 ( .A1(n15007), .A2(n15005), .ZN(n15092) );
  NAND2_X1 U15110 ( .A1(a_11_), .A2(b_6_), .ZN(n15008) );
  INV_X1 U15111 ( .A(n15093), .ZN(n15090) );
  NAND2_X1 U15112 ( .A1(n15005), .A2(n15007), .ZN(n15093) );
  NAND2_X1 U15113 ( .A1(n15094), .A2(n15095), .ZN(n15007) );
  NAND2_X1 U15114 ( .A1(n15004), .A2(n15096), .ZN(n15095) );
  INV_X1 U15115 ( .A(n15097), .ZN(n15096) );
  NOR2_X1 U15116 ( .A1(n15003), .A2(n15001), .ZN(n15097) );
  NOR2_X1 U15117 ( .A1(n8750), .A2(n14696), .ZN(n15004) );
  NAND2_X1 U15118 ( .A1(n15001), .A2(n15003), .ZN(n15094) );
  NAND2_X1 U15119 ( .A1(n15098), .A2(n15099), .ZN(n15003) );
  INV_X1 U15120 ( .A(n15100), .ZN(n15099) );
  NOR2_X1 U15121 ( .A1(n15000), .A2(n15101), .ZN(n15100) );
  NOR2_X1 U15122 ( .A1(n14999), .A2(n14997), .ZN(n15101) );
  NAND2_X1 U15123 ( .A1(a_13_), .A2(b_6_), .ZN(n15000) );
  NAND2_X1 U15124 ( .A1(n14997), .A2(n14999), .ZN(n15098) );
  NAND2_X1 U15125 ( .A1(n15102), .A2(n15103), .ZN(n14999) );
  NAND2_X1 U15126 ( .A1(n14996), .A2(n15104), .ZN(n15103) );
  INV_X1 U15127 ( .A(n15105), .ZN(n15104) );
  NOR2_X1 U15128 ( .A1(n14993), .A2(n14995), .ZN(n15105) );
  NOR2_X1 U15129 ( .A1(n8438), .A2(n14696), .ZN(n14996) );
  NAND2_X1 U15130 ( .A1(n14993), .A2(n14995), .ZN(n15102) );
  NAND2_X1 U15131 ( .A1(n15106), .A2(n15107), .ZN(n14995) );
  INV_X1 U15132 ( .A(n15108), .ZN(n15107) );
  NOR2_X1 U15133 ( .A1(n14992), .A2(n15109), .ZN(n15108) );
  NOR2_X1 U15134 ( .A1(n14991), .A2(n14989), .ZN(n15109) );
  NAND2_X1 U15135 ( .A1(a_15_), .A2(b_6_), .ZN(n14992) );
  NAND2_X1 U15136 ( .A1(n14989), .A2(n14991), .ZN(n15106) );
  NAND2_X1 U15137 ( .A1(n15110), .A2(n15111), .ZN(n14991) );
  NAND2_X1 U15138 ( .A1(n14988), .A2(n15112), .ZN(n15111) );
  INV_X1 U15139 ( .A(n15113), .ZN(n15112) );
  NOR2_X1 U15140 ( .A1(n14985), .A2(n14987), .ZN(n15113) );
  NOR2_X1 U15141 ( .A1(n8768), .A2(n14696), .ZN(n14988) );
  NAND2_X1 U15142 ( .A1(n14985), .A2(n14987), .ZN(n15110) );
  NAND2_X1 U15143 ( .A1(n15114), .A2(n15115), .ZN(n14987) );
  NAND2_X1 U15144 ( .A1(n14984), .A2(n15116), .ZN(n15115) );
  NAND2_X1 U15145 ( .A1(n14983), .A2(n14982), .ZN(n15116) );
  NOR2_X1 U15146 ( .A1(n8772), .A2(n14696), .ZN(n14984) );
  INV_X1 U15147 ( .A(n15117), .ZN(n15114) );
  NOR2_X1 U15148 ( .A1(n14982), .A2(n14983), .ZN(n15117) );
  NOR2_X1 U15149 ( .A1(n15118), .A2(n15119), .ZN(n14983) );
  INV_X1 U15150 ( .A(n15120), .ZN(n15119) );
  NAND2_X1 U15151 ( .A1(n14980), .A2(n15121), .ZN(n15120) );
  NAND2_X1 U15152 ( .A1(n14977), .A2(n14979), .ZN(n15121) );
  NOR2_X1 U15153 ( .A1(n10616), .A2(n14696), .ZN(n14980) );
  NOR2_X1 U15154 ( .A1(n14979), .A2(n14977), .ZN(n15118) );
  XOR2_X1 U15155 ( .A(n15122), .B(n15123), .Z(n14977) );
  XOR2_X1 U15156 ( .A(n15124), .B(n15125), .Z(n15123) );
  NAND2_X1 U15157 ( .A1(b_5_), .A2(a_19_), .ZN(n15125) );
  NAND2_X1 U15158 ( .A1(n15126), .A2(n15127), .ZN(n14979) );
  NAND2_X1 U15159 ( .A1(n14973), .A2(n15128), .ZN(n15127) );
  NAND2_X1 U15160 ( .A1(n14976), .A2(n14975), .ZN(n15128) );
  XOR2_X1 U15161 ( .A(n15129), .B(n15130), .Z(n14973) );
  XOR2_X1 U15162 ( .A(n15131), .B(n15132), .Z(n15130) );
  NAND2_X1 U15163 ( .A1(b_5_), .A2(a_20_), .ZN(n15132) );
  INV_X1 U15164 ( .A(n15133), .ZN(n15126) );
  NOR2_X1 U15165 ( .A1(n14975), .A2(n14976), .ZN(n15133) );
  NOR2_X1 U15166 ( .A1(n14696), .A2(n8881), .ZN(n14976) );
  NAND2_X1 U15167 ( .A1(n14971), .A2(n15134), .ZN(n14975) );
  NAND2_X1 U15168 ( .A1(n14970), .A2(n14972), .ZN(n15134) );
  NAND2_X1 U15169 ( .A1(n15135), .A2(n15136), .ZN(n14972) );
  INV_X1 U15170 ( .A(n15137), .ZN(n15136) );
  NAND2_X1 U15171 ( .A1(b_6_), .A2(a_20_), .ZN(n15135) );
  XNOR2_X1 U15172 ( .A(n15138), .B(n15139), .ZN(n14970) );
  XOR2_X1 U15173 ( .A(n15140), .B(n15141), .Z(n15139) );
  NAND2_X1 U15174 ( .A1(b_5_), .A2(a_21_), .ZN(n15141) );
  NAND2_X1 U15175 ( .A1(n15137), .A2(a_20_), .ZN(n14971) );
  NOR2_X1 U15176 ( .A1(n15142), .A2(n15143), .ZN(n15137) );
  INV_X1 U15177 ( .A(n15144), .ZN(n15143) );
  NAND2_X1 U15178 ( .A1(n14966), .A2(n15145), .ZN(n15144) );
  NAND2_X1 U15179 ( .A1(n14968), .A2(n14967), .ZN(n15145) );
  XOR2_X1 U15180 ( .A(n15146), .B(n15147), .Z(n14966) );
  XOR2_X1 U15181 ( .A(n15148), .B(n15149), .Z(n15147) );
  NAND2_X1 U15182 ( .A1(b_5_), .A2(a_22_), .ZN(n15149) );
  NOR2_X1 U15183 ( .A1(n14967), .A2(n14968), .ZN(n15142) );
  NOR2_X1 U15184 ( .A1(n14696), .A2(n8798), .ZN(n14968) );
  NAND2_X1 U15185 ( .A1(n14894), .A2(n15150), .ZN(n14967) );
  NAND2_X1 U15186 ( .A1(n14893), .A2(n14895), .ZN(n15150) );
  NAND2_X1 U15187 ( .A1(n15151), .A2(n15152), .ZN(n14895) );
  NAND2_X1 U15188 ( .A1(b_6_), .A2(a_22_), .ZN(n15152) );
  INV_X1 U15189 ( .A(n15153), .ZN(n15151) );
  XNOR2_X1 U15190 ( .A(n15154), .B(n15155), .ZN(n14893) );
  XOR2_X1 U15191 ( .A(n15156), .B(n15157), .Z(n15155) );
  NAND2_X1 U15192 ( .A1(b_5_), .A2(a_23_), .ZN(n15157) );
  NAND2_X1 U15193 ( .A1(a_22_), .A2(n15153), .ZN(n14894) );
  NAND2_X1 U15194 ( .A1(n15158), .A2(n15159), .ZN(n15153) );
  NAND2_X1 U15195 ( .A1(n15160), .A2(b_6_), .ZN(n15159) );
  NOR2_X1 U15196 ( .A1(n15161), .A2(n8812), .ZN(n15160) );
  NOR2_X1 U15197 ( .A1(n14899), .A2(n14901), .ZN(n15161) );
  NAND2_X1 U15198 ( .A1(n14899), .A2(n14901), .ZN(n15158) );
  NAND2_X1 U15199 ( .A1(n15162), .A2(n15163), .ZN(n14901) );
  NAND2_X1 U15200 ( .A1(n15164), .A2(b_6_), .ZN(n15163) );
  NOR2_X1 U15201 ( .A1(n15165), .A2(n9131), .ZN(n15164) );
  NOR2_X1 U15202 ( .A1(n14963), .A2(n14962), .ZN(n15165) );
  NAND2_X1 U15203 ( .A1(n14962), .A2(n14963), .ZN(n15162) );
  NAND2_X1 U15204 ( .A1(n15166), .A2(n15167), .ZN(n14963) );
  NAND2_X1 U15205 ( .A1(n14960), .A2(n15168), .ZN(n15167) );
  INV_X1 U15206 ( .A(n15169), .ZN(n15168) );
  NOR2_X1 U15207 ( .A1(n14957), .A2(n14959), .ZN(n15169) );
  NOR2_X1 U15208 ( .A1(n14696), .A2(n8825), .ZN(n14960) );
  NAND2_X1 U15209 ( .A1(n14957), .A2(n14959), .ZN(n15166) );
  NOR2_X1 U15210 ( .A1(n15170), .A2(n15171), .ZN(n14959) );
  INV_X1 U15211 ( .A(n15172), .ZN(n15171) );
  NAND2_X1 U15212 ( .A1(n14916), .A2(n15173), .ZN(n15172) );
  NAND2_X1 U15213 ( .A1(n14919), .A2(n14918), .ZN(n15173) );
  XNOR2_X1 U15214 ( .A(n15174), .B(n15175), .ZN(n14916) );
  XOR2_X1 U15215 ( .A(n15176), .B(n15177), .Z(n15175) );
  NOR2_X1 U15216 ( .A1(n14918), .A2(n14919), .ZN(n15170) );
  NOR2_X1 U15217 ( .A1(n14696), .A2(n8830), .ZN(n14919) );
  NAND2_X1 U15218 ( .A1(n15178), .A2(n15179), .ZN(n14918) );
  NAND2_X1 U15219 ( .A1(n14926), .A2(n15180), .ZN(n15179) );
  NAND2_X1 U15220 ( .A1(n14923), .A2(n14925), .ZN(n15180) );
  NOR2_X1 U15221 ( .A1(n14696), .A2(n8839), .ZN(n14926) );
  INV_X1 U15222 ( .A(n15181), .ZN(n15178) );
  NOR2_X1 U15223 ( .A1(n14923), .A2(n14925), .ZN(n15181) );
  NOR2_X1 U15224 ( .A1(n15182), .A2(n15183), .ZN(n14925) );
  INV_X1 U15225 ( .A(n15184), .ZN(n15183) );
  NAND2_X1 U15226 ( .A1(n14955), .A2(n15185), .ZN(n15184) );
  NAND2_X1 U15227 ( .A1(n14956), .A2(n14954), .ZN(n15185) );
  NOR2_X1 U15228 ( .A1(n14696), .A2(n8844), .ZN(n14955) );
  NOR2_X1 U15229 ( .A1(n14954), .A2(n14956), .ZN(n15182) );
  NOR2_X1 U15230 ( .A1(n15186), .A2(n15187), .ZN(n14956) );
  INV_X1 U15231 ( .A(n15188), .ZN(n15187) );
  NAND2_X1 U15232 ( .A1(n14949), .A2(n15189), .ZN(n15188) );
  NAND2_X1 U15233 ( .A1(n15190), .A2(n14951), .ZN(n15189) );
  NOR2_X1 U15234 ( .A1(n14696), .A2(n9161), .ZN(n14949) );
  NOR2_X1 U15235 ( .A1(n14951), .A2(n15190), .ZN(n15186) );
  INV_X1 U15236 ( .A(n14952), .ZN(n15190) );
  NAND2_X1 U15237 ( .A1(n15191), .A2(n15192), .ZN(n14952) );
  NAND2_X1 U15238 ( .A1(b_4_), .A2(n15193), .ZN(n15192) );
  NAND2_X1 U15239 ( .A1(n8358), .A2(n15194), .ZN(n15193) );
  NAND2_X1 U15240 ( .A1(a_31_), .A2(n14947), .ZN(n15194) );
  NAND2_X1 U15241 ( .A1(b_5_), .A2(n15195), .ZN(n15191) );
  NAND2_X1 U15242 ( .A1(n8362), .A2(n15196), .ZN(n15195) );
  NAND2_X1 U15243 ( .A1(a_30_), .A2(n15197), .ZN(n15196) );
  NAND2_X1 U15244 ( .A1(n15198), .A2(b_5_), .ZN(n14951) );
  NOR2_X1 U15245 ( .A1(n9170), .A2(n14696), .ZN(n15198) );
  XOR2_X1 U15246 ( .A(n15199), .B(n15200), .Z(n14954) );
  XOR2_X1 U15247 ( .A(n15201), .B(n15202), .Z(n15200) );
  XOR2_X1 U15248 ( .A(n15203), .B(n15204), .Z(n14923) );
  XNOR2_X1 U15249 ( .A(n15205), .B(n15206), .ZN(n15203) );
  XOR2_X1 U15250 ( .A(n15207), .B(n15208), .Z(n14957) );
  XNOR2_X1 U15251 ( .A(n15209), .B(n15210), .ZN(n15208) );
  XNOR2_X1 U15252 ( .A(n15211), .B(n15212), .ZN(n14962) );
  XNOR2_X1 U15253 ( .A(n15213), .B(n15214), .ZN(n15212) );
  XOR2_X1 U15254 ( .A(n15215), .B(n15216), .Z(n14899) );
  XOR2_X1 U15255 ( .A(n15217), .B(n15218), .Z(n15215) );
  NOR2_X1 U15256 ( .A1(n9131), .A2(n14947), .ZN(n15218) );
  XNOR2_X1 U15257 ( .A(n15219), .B(n15220), .ZN(n14982) );
  XOR2_X1 U15258 ( .A(n15221), .B(n15222), .Z(n15219) );
  NOR2_X1 U15259 ( .A1(n14947), .A2(n10616), .ZN(n15222) );
  XOR2_X1 U15260 ( .A(n15223), .B(n15224), .Z(n14985) );
  XOR2_X1 U15261 ( .A(n15225), .B(n15226), .Z(n15223) );
  NOR2_X1 U15262 ( .A1(n14947), .A2(n8772), .ZN(n15226) );
  XOR2_X1 U15263 ( .A(n15227), .B(n15228), .Z(n14989) );
  XOR2_X1 U15264 ( .A(n15229), .B(n15230), .Z(n15227) );
  NOR2_X1 U15265 ( .A1(n14947), .A2(n8768), .ZN(n15230) );
  XOR2_X1 U15266 ( .A(n15231), .B(n15232), .Z(n14993) );
  XOR2_X1 U15267 ( .A(n15233), .B(n15234), .Z(n15231) );
  NOR2_X1 U15268 ( .A1(n14947), .A2(n8763), .ZN(n15234) );
  XOR2_X1 U15269 ( .A(n15235), .B(n15236), .Z(n14997) );
  XOR2_X1 U15270 ( .A(n15237), .B(n15238), .Z(n15235) );
  NOR2_X1 U15271 ( .A1(n14947), .A2(n8438), .ZN(n15238) );
  XOR2_X1 U15272 ( .A(n15239), .B(n15240), .Z(n15001) );
  XOR2_X1 U15273 ( .A(n15241), .B(n15242), .Z(n15239) );
  NOR2_X1 U15274 ( .A1(n14947), .A2(n8443), .ZN(n15242) );
  XOR2_X1 U15275 ( .A(n15243), .B(n15244), .Z(n15005) );
  XOR2_X1 U15276 ( .A(n15245), .B(n15246), .Z(n15243) );
  NOR2_X1 U15277 ( .A1(n14947), .A2(n8750), .ZN(n15246) );
  INV_X1 U15278 ( .A(n15009), .ZN(n15088) );
  XNOR2_X1 U15279 ( .A(n15247), .B(n15248), .ZN(n15009) );
  XOR2_X1 U15280 ( .A(n15249), .B(n15250), .Z(n15247) );
  NOR2_X1 U15281 ( .A1(n14947), .A2(n8452), .ZN(n15250) );
  XOR2_X1 U15282 ( .A(n15251), .B(n15252), .Z(n15013) );
  XOR2_X1 U15283 ( .A(n15253), .B(n15254), .Z(n15251) );
  NOR2_X1 U15284 ( .A1(n14947), .A2(n8741), .ZN(n15254) );
  INV_X1 U15285 ( .A(n14831), .ZN(n15079) );
  XNOR2_X1 U15286 ( .A(n15255), .B(n15256), .ZN(n14831) );
  XOR2_X1 U15287 ( .A(n15257), .B(n15258), .Z(n15255) );
  NOR2_X1 U15288 ( .A1(n14947), .A2(n8736), .ZN(n15258) );
  XOR2_X1 U15289 ( .A(n15259), .B(n15260), .Z(n14823) );
  XOR2_X1 U15290 ( .A(n15261), .B(n15262), .Z(n15259) );
  NOR2_X1 U15291 ( .A1(n14947), .A2(n8731), .ZN(n15262) );
  XOR2_X1 U15292 ( .A(n15263), .B(n15264), .Z(n15017) );
  XOR2_X1 U15293 ( .A(n15265), .B(n15266), .Z(n15263) );
  NOR2_X1 U15294 ( .A1(n14947), .A2(n8726), .ZN(n15266) );
  XNOR2_X1 U15295 ( .A(n15267), .B(n15268), .ZN(n15021) );
  XOR2_X1 U15296 ( .A(n15269), .B(n15270), .Z(n15267) );
  NOR2_X1 U15297 ( .A1(n14947), .A2(n8480), .ZN(n15270) );
  XNOR2_X1 U15298 ( .A(n15271), .B(n15272), .ZN(n15025) );
  XOR2_X1 U15299 ( .A(n15273), .B(n15274), .Z(n15271) );
  XOR2_X1 U15300 ( .A(n15275), .B(n15276), .Z(n15030) );
  XNOR2_X1 U15301 ( .A(n15277), .B(n15278), .ZN(n15276) );
  NAND2_X1 U15302 ( .A1(a_4_), .A2(b_5_), .ZN(n15278) );
  XOR2_X1 U15303 ( .A(n15279), .B(n15280), .Z(n15034) );
  XNOR2_X1 U15304 ( .A(n15281), .B(n15282), .ZN(n15279) );
  NAND2_X1 U15305 ( .A1(a_3_), .A2(b_5_), .ZN(n15281) );
  XOR2_X1 U15306 ( .A(n15283), .B(n15284), .Z(n15038) );
  XOR2_X1 U15307 ( .A(n15285), .B(n15286), .Z(n15283) );
  NOR2_X1 U15308 ( .A1(n14947), .A2(n8497), .ZN(n15286) );
  XOR2_X1 U15309 ( .A(n15287), .B(n15288), .Z(n14790) );
  XOR2_X1 U15310 ( .A(n15289), .B(n15290), .Z(n15287) );
  NOR2_X1 U15311 ( .A1(n14947), .A2(n8502), .ZN(n15290) );
  XNOR2_X1 U15312 ( .A(n15291), .B(n15292), .ZN(n15041) );
  XOR2_X1 U15313 ( .A(n15293), .B(n15294), .Z(n15291) );
  NOR2_X1 U15314 ( .A1(n14947), .A2(n8690), .ZN(n15294) );
  NOR2_X1 U15315 ( .A1(n15295), .A2(n8615), .ZN(n8378) );
  INV_X1 U15316 ( .A(n15296), .ZN(n8615) );
  NAND2_X1 U15317 ( .A1(n15297), .A2(n15298), .ZN(n15296) );
  NOR2_X1 U15318 ( .A1(n15298), .A2(n15297), .ZN(n15295) );
  XNOR2_X1 U15319 ( .A(n15299), .B(n15300), .ZN(n15297) );
  XNOR2_X1 U15320 ( .A(n15301), .B(n15302), .ZN(n15299) );
  NAND2_X1 U15321 ( .A1(n15303), .A2(n15304), .ZN(n15298) );
  NAND2_X1 U15322 ( .A1(n15305), .A2(a_0_), .ZN(n15304) );
  NOR2_X1 U15323 ( .A1(n15306), .A2(n14947), .ZN(n15305) );
  NOR2_X1 U15324 ( .A1(n15292), .A2(n15293), .ZN(n15306) );
  NAND2_X1 U15325 ( .A1(n15292), .A2(n15293), .ZN(n15303) );
  NAND2_X1 U15326 ( .A1(n15307), .A2(n15308), .ZN(n15293) );
  NAND2_X1 U15327 ( .A1(n15309), .A2(a_1_), .ZN(n15308) );
  NOR2_X1 U15328 ( .A1(n15310), .A2(n14947), .ZN(n15309) );
  NOR2_X1 U15329 ( .A1(n15289), .A2(n15288), .ZN(n15310) );
  NAND2_X1 U15330 ( .A1(n15288), .A2(n15289), .ZN(n15307) );
  NAND2_X1 U15331 ( .A1(n15311), .A2(n15312), .ZN(n15289) );
  NAND2_X1 U15332 ( .A1(n15313), .A2(a_2_), .ZN(n15312) );
  NOR2_X1 U15333 ( .A1(n15314), .A2(n14947), .ZN(n15313) );
  NOR2_X1 U15334 ( .A1(n15284), .A2(n15285), .ZN(n15314) );
  NAND2_X1 U15335 ( .A1(n15284), .A2(n15285), .ZN(n15311) );
  NAND2_X1 U15336 ( .A1(n15315), .A2(n15316), .ZN(n15285) );
  NAND2_X1 U15337 ( .A1(n15317), .A2(a_3_), .ZN(n15316) );
  NOR2_X1 U15338 ( .A1(n15318), .A2(n14947), .ZN(n15317) );
  NOR2_X1 U15339 ( .A1(n15280), .A2(n15282), .ZN(n15318) );
  NAND2_X1 U15340 ( .A1(n15280), .A2(n15282), .ZN(n15315) );
  NAND2_X1 U15341 ( .A1(n15319), .A2(n15320), .ZN(n15282) );
  NAND2_X1 U15342 ( .A1(n15321), .A2(a_4_), .ZN(n15320) );
  NOR2_X1 U15343 ( .A1(n15322), .A2(n14947), .ZN(n15321) );
  NOR2_X1 U15344 ( .A1(n15277), .A2(n15275), .ZN(n15322) );
  NAND2_X1 U15345 ( .A1(n15277), .A2(n15275), .ZN(n15319) );
  XOR2_X1 U15346 ( .A(n15323), .B(n15324), .Z(n15275) );
  XOR2_X1 U15347 ( .A(n15325), .B(n15326), .Z(n15323) );
  NOR2_X1 U15348 ( .A1(n15327), .A2(n15328), .ZN(n15277) );
  INV_X1 U15349 ( .A(n15329), .ZN(n15328) );
  NAND2_X1 U15350 ( .A1(n15272), .A2(n15330), .ZN(n15329) );
  NAND2_X1 U15351 ( .A1(n15274), .A2(n15273), .ZN(n15330) );
  XOR2_X1 U15352 ( .A(n15331), .B(n15332), .Z(n15272) );
  XNOR2_X1 U15353 ( .A(n15333), .B(n15334), .ZN(n15332) );
  NOR2_X1 U15354 ( .A1(n15273), .A2(n15274), .ZN(n15327) );
  NAND2_X1 U15355 ( .A1(n15335), .A2(n15336), .ZN(n15273) );
  NAND2_X1 U15356 ( .A1(n15337), .A2(a_6_), .ZN(n15336) );
  NOR2_X1 U15357 ( .A1(n15338), .A2(n14947), .ZN(n15337) );
  NOR2_X1 U15358 ( .A1(n15269), .A2(n15268), .ZN(n15338) );
  NAND2_X1 U15359 ( .A1(n15268), .A2(n15269), .ZN(n15335) );
  NAND2_X1 U15360 ( .A1(n15339), .A2(n15340), .ZN(n15269) );
  NAND2_X1 U15361 ( .A1(n15341), .A2(a_7_), .ZN(n15340) );
  NOR2_X1 U15362 ( .A1(n15342), .A2(n14947), .ZN(n15341) );
  NOR2_X1 U15363 ( .A1(n15264), .A2(n15265), .ZN(n15342) );
  NAND2_X1 U15364 ( .A1(n15264), .A2(n15265), .ZN(n15339) );
  NAND2_X1 U15365 ( .A1(n15343), .A2(n15344), .ZN(n15265) );
  NAND2_X1 U15366 ( .A1(n15345), .A2(a_8_), .ZN(n15344) );
  NOR2_X1 U15367 ( .A1(n15346), .A2(n14947), .ZN(n15345) );
  NOR2_X1 U15368 ( .A1(n15261), .A2(n15260), .ZN(n15346) );
  NAND2_X1 U15369 ( .A1(n15260), .A2(n15261), .ZN(n15343) );
  NAND2_X1 U15370 ( .A1(n15347), .A2(n15348), .ZN(n15261) );
  NAND2_X1 U15371 ( .A1(n15349), .A2(a_9_), .ZN(n15348) );
  NOR2_X1 U15372 ( .A1(n15350), .A2(n14947), .ZN(n15349) );
  NOR2_X1 U15373 ( .A1(n15256), .A2(n15257), .ZN(n15350) );
  NAND2_X1 U15374 ( .A1(n15256), .A2(n15257), .ZN(n15347) );
  NAND2_X1 U15375 ( .A1(n15351), .A2(n15352), .ZN(n15257) );
  NAND2_X1 U15376 ( .A1(n15353), .A2(a_10_), .ZN(n15352) );
  NOR2_X1 U15377 ( .A1(n15354), .A2(n14947), .ZN(n15353) );
  NOR2_X1 U15378 ( .A1(n15253), .A2(n15252), .ZN(n15354) );
  NAND2_X1 U15379 ( .A1(n15252), .A2(n15253), .ZN(n15351) );
  NAND2_X1 U15380 ( .A1(n15355), .A2(n15356), .ZN(n15253) );
  NAND2_X1 U15381 ( .A1(n15357), .A2(a_11_), .ZN(n15356) );
  NOR2_X1 U15382 ( .A1(n15358), .A2(n14947), .ZN(n15357) );
  NOR2_X1 U15383 ( .A1(n15248), .A2(n15249), .ZN(n15358) );
  NAND2_X1 U15384 ( .A1(n15248), .A2(n15249), .ZN(n15355) );
  NAND2_X1 U15385 ( .A1(n15359), .A2(n15360), .ZN(n15249) );
  NAND2_X1 U15386 ( .A1(n15361), .A2(a_12_), .ZN(n15360) );
  NOR2_X1 U15387 ( .A1(n15362), .A2(n14947), .ZN(n15361) );
  NOR2_X1 U15388 ( .A1(n15245), .A2(n15244), .ZN(n15362) );
  NAND2_X1 U15389 ( .A1(n15244), .A2(n15245), .ZN(n15359) );
  NAND2_X1 U15390 ( .A1(n15363), .A2(n15364), .ZN(n15245) );
  NAND2_X1 U15391 ( .A1(n15365), .A2(a_13_), .ZN(n15364) );
  NOR2_X1 U15392 ( .A1(n15366), .A2(n14947), .ZN(n15365) );
  NOR2_X1 U15393 ( .A1(n15241), .A2(n15240), .ZN(n15366) );
  NAND2_X1 U15394 ( .A1(n15240), .A2(n15241), .ZN(n15363) );
  NAND2_X1 U15395 ( .A1(n15367), .A2(n15368), .ZN(n15241) );
  NAND2_X1 U15396 ( .A1(n15369), .A2(a_14_), .ZN(n15368) );
  NOR2_X1 U15397 ( .A1(n15370), .A2(n14947), .ZN(n15369) );
  NOR2_X1 U15398 ( .A1(n15237), .A2(n15236), .ZN(n15370) );
  NAND2_X1 U15399 ( .A1(n15236), .A2(n15237), .ZN(n15367) );
  NAND2_X1 U15400 ( .A1(n15371), .A2(n15372), .ZN(n15237) );
  NAND2_X1 U15401 ( .A1(n15373), .A2(a_15_), .ZN(n15372) );
  NOR2_X1 U15402 ( .A1(n15374), .A2(n14947), .ZN(n15373) );
  NOR2_X1 U15403 ( .A1(n15232), .A2(n15233), .ZN(n15374) );
  NAND2_X1 U15404 ( .A1(n15232), .A2(n15233), .ZN(n15371) );
  NAND2_X1 U15405 ( .A1(n15375), .A2(n15376), .ZN(n15233) );
  NAND2_X1 U15406 ( .A1(n15377), .A2(a_16_), .ZN(n15376) );
  NOR2_X1 U15407 ( .A1(n15378), .A2(n14947), .ZN(n15377) );
  NOR2_X1 U15408 ( .A1(n15229), .A2(n15228), .ZN(n15378) );
  NAND2_X1 U15409 ( .A1(n15228), .A2(n15229), .ZN(n15375) );
  NAND2_X1 U15410 ( .A1(n15379), .A2(n15380), .ZN(n15229) );
  NAND2_X1 U15411 ( .A1(n15381), .A2(a_17_), .ZN(n15380) );
  NOR2_X1 U15412 ( .A1(n15382), .A2(n14947), .ZN(n15381) );
  NOR2_X1 U15413 ( .A1(n15224), .A2(n15225), .ZN(n15382) );
  NAND2_X1 U15414 ( .A1(n15224), .A2(n15225), .ZN(n15379) );
  NAND2_X1 U15415 ( .A1(n15383), .A2(n15384), .ZN(n15225) );
  NAND2_X1 U15416 ( .A1(n15385), .A2(a_18_), .ZN(n15384) );
  NOR2_X1 U15417 ( .A1(n15386), .A2(n14947), .ZN(n15385) );
  NOR2_X1 U15418 ( .A1(n15221), .A2(n15220), .ZN(n15386) );
  NAND2_X1 U15419 ( .A1(n15220), .A2(n15221), .ZN(n15383) );
  NAND2_X1 U15420 ( .A1(n15387), .A2(n15388), .ZN(n15221) );
  NAND2_X1 U15421 ( .A1(n15389), .A2(b_5_), .ZN(n15388) );
  NOR2_X1 U15422 ( .A1(n15390), .A2(n8881), .ZN(n15389) );
  NOR2_X1 U15423 ( .A1(n15122), .A2(n15124), .ZN(n15390) );
  NAND2_X1 U15424 ( .A1(n15122), .A2(n15124), .ZN(n15387) );
  NAND2_X1 U15425 ( .A1(n15391), .A2(n15392), .ZN(n15124) );
  NAND2_X1 U15426 ( .A1(n15393), .A2(b_5_), .ZN(n15392) );
  NOR2_X1 U15427 ( .A1(n15394), .A2(n10633), .ZN(n15393) );
  NOR2_X1 U15428 ( .A1(n15131), .A2(n15129), .ZN(n15394) );
  NAND2_X1 U15429 ( .A1(n15129), .A2(n15131), .ZN(n15391) );
  NAND2_X1 U15430 ( .A1(n15395), .A2(n15396), .ZN(n15131) );
  NAND2_X1 U15431 ( .A1(n15397), .A2(b_5_), .ZN(n15396) );
  NOR2_X1 U15432 ( .A1(n15398), .A2(n8798), .ZN(n15397) );
  NOR2_X1 U15433 ( .A1(n15140), .A2(n15138), .ZN(n15398) );
  NAND2_X1 U15434 ( .A1(n15138), .A2(n15140), .ZN(n15395) );
  NAND2_X1 U15435 ( .A1(n15399), .A2(n15400), .ZN(n15140) );
  NAND2_X1 U15436 ( .A1(n15401), .A2(b_5_), .ZN(n15400) );
  NOR2_X1 U15437 ( .A1(n15402), .A2(n8803), .ZN(n15401) );
  NOR2_X1 U15438 ( .A1(n15146), .A2(n15148), .ZN(n15402) );
  NAND2_X1 U15439 ( .A1(n15146), .A2(n15148), .ZN(n15399) );
  NAND2_X1 U15440 ( .A1(n15403), .A2(n15404), .ZN(n15148) );
  NAND2_X1 U15441 ( .A1(n15405), .A2(b_5_), .ZN(n15404) );
  NOR2_X1 U15442 ( .A1(n15406), .A2(n8812), .ZN(n15405) );
  NOR2_X1 U15443 ( .A1(n15154), .A2(n15156), .ZN(n15406) );
  NAND2_X1 U15444 ( .A1(n15154), .A2(n15156), .ZN(n15403) );
  NAND2_X1 U15445 ( .A1(n15407), .A2(n15408), .ZN(n15156) );
  NAND2_X1 U15446 ( .A1(n15409), .A2(b_5_), .ZN(n15408) );
  NOR2_X1 U15447 ( .A1(n15410), .A2(n9131), .ZN(n15409) );
  NOR2_X1 U15448 ( .A1(n15217), .A2(n15216), .ZN(n15410) );
  NAND2_X1 U15449 ( .A1(n15216), .A2(n15217), .ZN(n15407) );
  NAND2_X1 U15450 ( .A1(n15411), .A2(n15412), .ZN(n15217) );
  NAND2_X1 U15451 ( .A1(n15214), .A2(n15413), .ZN(n15412) );
  NAND2_X1 U15452 ( .A1(n15211), .A2(n15213), .ZN(n15413) );
  NOR2_X1 U15453 ( .A1(n14947), .A2(n8825), .ZN(n15214) );
  INV_X1 U15454 ( .A(n15414), .ZN(n15411) );
  NOR2_X1 U15455 ( .A1(n15213), .A2(n15211), .ZN(n15414) );
  XOR2_X1 U15456 ( .A(n15415), .B(n15416), .Z(n15211) );
  XOR2_X1 U15457 ( .A(n15417), .B(n15418), .Z(n15415) );
  NAND2_X1 U15458 ( .A1(n15419), .A2(n15420), .ZN(n15213) );
  NAND2_X1 U15459 ( .A1(n15207), .A2(n15421), .ZN(n15420) );
  NAND2_X1 U15460 ( .A1(n15210), .A2(n15209), .ZN(n15421) );
  XOR2_X1 U15461 ( .A(n15422), .B(n15423), .Z(n15207) );
  NAND2_X1 U15462 ( .A1(n15424), .A2(n15425), .ZN(n15422) );
  INV_X1 U15463 ( .A(n15426), .ZN(n15419) );
  NOR2_X1 U15464 ( .A1(n15209), .A2(n15210), .ZN(n15426) );
  NOR2_X1 U15465 ( .A1(n14947), .A2(n8830), .ZN(n15210) );
  NAND2_X1 U15466 ( .A1(n15427), .A2(n15428), .ZN(n15209) );
  NAND2_X1 U15467 ( .A1(n15177), .A2(n15429), .ZN(n15428) );
  NAND2_X1 U15468 ( .A1(n15174), .A2(n15176), .ZN(n15429) );
  NOR2_X1 U15469 ( .A1(n14947), .A2(n8839), .ZN(n15177) );
  INV_X1 U15470 ( .A(n15430), .ZN(n15427) );
  NOR2_X1 U15471 ( .A1(n15174), .A2(n15176), .ZN(n15430) );
  NOR2_X1 U15472 ( .A1(n15431), .A2(n15432), .ZN(n15176) );
  INV_X1 U15473 ( .A(n15433), .ZN(n15432) );
  NAND2_X1 U15474 ( .A1(n15205), .A2(n15434), .ZN(n15433) );
  NAND2_X1 U15475 ( .A1(n15206), .A2(n15204), .ZN(n15434) );
  NOR2_X1 U15476 ( .A1(n14947), .A2(n8844), .ZN(n15205) );
  NOR2_X1 U15477 ( .A1(n15204), .A2(n15206), .ZN(n15431) );
  NOR2_X1 U15478 ( .A1(n15435), .A2(n15436), .ZN(n15206) );
  INV_X1 U15479 ( .A(n15437), .ZN(n15436) );
  NAND2_X1 U15480 ( .A1(n15199), .A2(n15438), .ZN(n15437) );
  NAND2_X1 U15481 ( .A1(n15439), .A2(n15201), .ZN(n15438) );
  NOR2_X1 U15482 ( .A1(n14947), .A2(n9161), .ZN(n15199) );
  NOR2_X1 U15483 ( .A1(n15201), .A2(n15439), .ZN(n15435) );
  INV_X1 U15484 ( .A(n15202), .ZN(n15439) );
  NAND2_X1 U15485 ( .A1(n15440), .A2(n15441), .ZN(n15202) );
  NAND2_X1 U15486 ( .A1(b_3_), .A2(n15442), .ZN(n15441) );
  NAND2_X1 U15487 ( .A1(n8358), .A2(n15443), .ZN(n15442) );
  NAND2_X1 U15488 ( .A1(a_31_), .A2(n15197), .ZN(n15443) );
  NAND2_X1 U15489 ( .A1(b_4_), .A2(n15444), .ZN(n15440) );
  NAND2_X1 U15490 ( .A1(n8362), .A2(n15445), .ZN(n15444) );
  NAND2_X1 U15491 ( .A1(a_30_), .A2(n15446), .ZN(n15445) );
  NAND2_X1 U15492 ( .A1(n15447), .A2(b_4_), .ZN(n15201) );
  NOR2_X1 U15493 ( .A1(n9170), .A2(n14947), .ZN(n15447) );
  XOR2_X1 U15494 ( .A(n15448), .B(n15449), .Z(n15204) );
  XOR2_X1 U15495 ( .A(n15450), .B(n15451), .Z(n15449) );
  XOR2_X1 U15496 ( .A(n15452), .B(n15453), .Z(n15174) );
  XNOR2_X1 U15497 ( .A(n15454), .B(n15455), .ZN(n15452) );
  XNOR2_X1 U15498 ( .A(n15456), .B(n15457), .ZN(n15216) );
  XNOR2_X1 U15499 ( .A(n15458), .B(n15459), .ZN(n15457) );
  XNOR2_X1 U15500 ( .A(n15460), .B(n15461), .ZN(n15154) );
  XOR2_X1 U15501 ( .A(n15462), .B(n15463), .Z(n15461) );
  XNOR2_X1 U15502 ( .A(n15464), .B(n15465), .ZN(n15146) );
  XNOR2_X1 U15503 ( .A(n15466), .B(n15467), .ZN(n15464) );
  XNOR2_X1 U15504 ( .A(n15468), .B(n15469), .ZN(n15138) );
  XNOR2_X1 U15505 ( .A(n15470), .B(n15471), .ZN(n15469) );
  XOR2_X1 U15506 ( .A(n15472), .B(n15473), .Z(n15129) );
  XOR2_X1 U15507 ( .A(n15474), .B(n15475), .Z(n15472) );
  XNOR2_X1 U15508 ( .A(n15476), .B(n15477), .ZN(n15122) );
  XNOR2_X1 U15509 ( .A(n15478), .B(n15479), .ZN(n15477) );
  XOR2_X1 U15510 ( .A(n15480), .B(n15481), .Z(n15220) );
  XOR2_X1 U15511 ( .A(n15482), .B(n15483), .Z(n15480) );
  XNOR2_X1 U15512 ( .A(n15484), .B(n15485), .ZN(n15224) );
  XNOR2_X1 U15513 ( .A(n15486), .B(n15487), .ZN(n15485) );
  XOR2_X1 U15514 ( .A(n15488), .B(n15489), .Z(n15228) );
  XOR2_X1 U15515 ( .A(n15490), .B(n15491), .Z(n15488) );
  XNOR2_X1 U15516 ( .A(n15492), .B(n15493), .ZN(n15232) );
  XNOR2_X1 U15517 ( .A(n15494), .B(n15495), .ZN(n15493) );
  XOR2_X1 U15518 ( .A(n15496), .B(n15497), .Z(n15236) );
  XOR2_X1 U15519 ( .A(n15498), .B(n15499), .Z(n15496) );
  XNOR2_X1 U15520 ( .A(n15500), .B(n15501), .ZN(n15240) );
  XNOR2_X1 U15521 ( .A(n15502), .B(n15503), .ZN(n15501) );
  XOR2_X1 U15522 ( .A(n15504), .B(n15505), .Z(n15244) );
  XOR2_X1 U15523 ( .A(n15506), .B(n15507), .Z(n15504) );
  XNOR2_X1 U15524 ( .A(n15508), .B(n15509), .ZN(n15248) );
  XNOR2_X1 U15525 ( .A(n15510), .B(n15511), .ZN(n15509) );
  XOR2_X1 U15526 ( .A(n15512), .B(n15513), .Z(n15252) );
  XOR2_X1 U15527 ( .A(n15514), .B(n15515), .Z(n15512) );
  XNOR2_X1 U15528 ( .A(n15516), .B(n15517), .ZN(n15256) );
  XNOR2_X1 U15529 ( .A(n15518), .B(n15519), .ZN(n15517) );
  XOR2_X1 U15530 ( .A(n15520), .B(n15521), .Z(n15260) );
  XOR2_X1 U15531 ( .A(n15522), .B(n15523), .Z(n15520) );
  XNOR2_X1 U15532 ( .A(n15524), .B(n15525), .ZN(n15264) );
  XNOR2_X1 U15533 ( .A(n15526), .B(n15527), .ZN(n15525) );
  XOR2_X1 U15534 ( .A(n15528), .B(n15529), .Z(n15268) );
  XOR2_X1 U15535 ( .A(n15530), .B(n15531), .Z(n15528) );
  XNOR2_X1 U15536 ( .A(n15532), .B(n15533), .ZN(n15280) );
  XOR2_X1 U15537 ( .A(n15534), .B(n15535), .Z(n15533) );
  XNOR2_X1 U15538 ( .A(n15536), .B(n15537), .ZN(n15284) );
  XNOR2_X1 U15539 ( .A(n15538), .B(n15539), .ZN(n15536) );
  XNOR2_X1 U15540 ( .A(n15540), .B(n15541), .ZN(n15288) );
  XNOR2_X1 U15541 ( .A(n15542), .B(n15543), .ZN(n15541) );
  XNOR2_X1 U15542 ( .A(n15544), .B(n15545), .ZN(n15292) );
  XNOR2_X1 U15543 ( .A(n15546), .B(n15547), .ZN(n15545) );
  XNOR2_X1 U15544 ( .A(n15548), .B(n15549), .ZN(n8421) );
  NAND2_X1 U15545 ( .A1(n8470), .A2(n8471), .ZN(n8469) );
  INV_X1 U15546 ( .A(n15550), .ZN(n8471) );
  NAND2_X1 U15547 ( .A1(n15549), .A2(n15548), .ZN(n15550) );
  NAND2_X1 U15548 ( .A1(n15551), .A2(n15552), .ZN(n15548) );
  NAND2_X1 U15549 ( .A1(n15302), .A2(n15553), .ZN(n15552) );
  INV_X1 U15550 ( .A(n15554), .ZN(n15553) );
  NOR2_X1 U15551 ( .A1(n15300), .A2(n15301), .ZN(n15554) );
  NOR2_X1 U15552 ( .A1(n8690), .A2(n15197), .ZN(n15302) );
  NAND2_X1 U15553 ( .A1(n15300), .A2(n15301), .ZN(n15551) );
  NAND2_X1 U15554 ( .A1(n15555), .A2(n15556), .ZN(n15301) );
  NAND2_X1 U15555 ( .A1(n15547), .A2(n15557), .ZN(n15556) );
  INV_X1 U15556 ( .A(n15558), .ZN(n15557) );
  NOR2_X1 U15557 ( .A1(n15544), .A2(n15546), .ZN(n15558) );
  NOR2_X1 U15558 ( .A1(n8502), .A2(n15197), .ZN(n15547) );
  NAND2_X1 U15559 ( .A1(n15544), .A2(n15546), .ZN(n15555) );
  NAND2_X1 U15560 ( .A1(n15559), .A2(n15560), .ZN(n15546) );
  NAND2_X1 U15561 ( .A1(n15543), .A2(n15561), .ZN(n15560) );
  INV_X1 U15562 ( .A(n15562), .ZN(n15561) );
  NOR2_X1 U15563 ( .A1(n15542), .A2(n15540), .ZN(n15562) );
  NOR2_X1 U15564 ( .A1(n8497), .A2(n15197), .ZN(n15543) );
  NAND2_X1 U15565 ( .A1(n15540), .A2(n15542), .ZN(n15559) );
  NAND2_X1 U15566 ( .A1(n15563), .A2(n15564), .ZN(n15542) );
  NAND2_X1 U15567 ( .A1(n15539), .A2(n15565), .ZN(n15564) );
  INV_X1 U15568 ( .A(n15566), .ZN(n15565) );
  NOR2_X1 U15569 ( .A1(n15537), .A2(n15538), .ZN(n15566) );
  NOR2_X1 U15570 ( .A1(n8707), .A2(n15197), .ZN(n15539) );
  NAND2_X1 U15571 ( .A1(n15537), .A2(n15538), .ZN(n15563) );
  NOR2_X1 U15572 ( .A1(n15567), .A2(n15568), .ZN(n15538) );
  INV_X1 U15573 ( .A(n15569), .ZN(n15568) );
  NAND2_X1 U15574 ( .A1(n15570), .A2(n15535), .ZN(n15569) );
  NAND2_X1 U15575 ( .A1(n15532), .A2(n15534), .ZN(n15570) );
  NOR2_X1 U15576 ( .A1(n15532), .A2(n15534), .ZN(n15567) );
  NAND2_X1 U15577 ( .A1(n15571), .A2(n15572), .ZN(n15534) );
  NAND2_X1 U15578 ( .A1(n15326), .A2(n15573), .ZN(n15572) );
  INV_X1 U15579 ( .A(n15574), .ZN(n15573) );
  NOR2_X1 U15580 ( .A1(n15325), .A2(n15324), .ZN(n15574) );
  NOR2_X1 U15581 ( .A1(n8717), .A2(n15197), .ZN(n15326) );
  NAND2_X1 U15582 ( .A1(n15324), .A2(n15325), .ZN(n15571) );
  NAND2_X1 U15583 ( .A1(n15575), .A2(n15576), .ZN(n15325) );
  NAND2_X1 U15584 ( .A1(n15334), .A2(n15577), .ZN(n15576) );
  INV_X1 U15585 ( .A(n15578), .ZN(n15577) );
  NOR2_X1 U15586 ( .A1(n15331), .A2(n15333), .ZN(n15578) );
  NOR2_X1 U15587 ( .A1(n8480), .A2(n15197), .ZN(n15334) );
  NAND2_X1 U15588 ( .A1(n15331), .A2(n15333), .ZN(n15575) );
  NAND2_X1 U15589 ( .A1(n15579), .A2(n15580), .ZN(n15333) );
  NAND2_X1 U15590 ( .A1(n15531), .A2(n15581), .ZN(n15580) );
  INV_X1 U15591 ( .A(n15582), .ZN(n15581) );
  NOR2_X1 U15592 ( .A1(n15530), .A2(n15529), .ZN(n15582) );
  NOR2_X1 U15593 ( .A1(n8726), .A2(n15197), .ZN(n15531) );
  NAND2_X1 U15594 ( .A1(n15529), .A2(n15530), .ZN(n15579) );
  NAND2_X1 U15595 ( .A1(n15583), .A2(n15584), .ZN(n15530) );
  NAND2_X1 U15596 ( .A1(n15527), .A2(n15585), .ZN(n15584) );
  INV_X1 U15597 ( .A(n15586), .ZN(n15585) );
  NOR2_X1 U15598 ( .A1(n15524), .A2(n15526), .ZN(n15586) );
  NOR2_X1 U15599 ( .A1(n8731), .A2(n15197), .ZN(n15527) );
  NAND2_X1 U15600 ( .A1(n15524), .A2(n15526), .ZN(n15583) );
  NAND2_X1 U15601 ( .A1(n15587), .A2(n15588), .ZN(n15526) );
  NAND2_X1 U15602 ( .A1(n15523), .A2(n15589), .ZN(n15588) );
  INV_X1 U15603 ( .A(n15590), .ZN(n15589) );
  NOR2_X1 U15604 ( .A1(n15522), .A2(n15521), .ZN(n15590) );
  NOR2_X1 U15605 ( .A1(n8736), .A2(n15197), .ZN(n15523) );
  NAND2_X1 U15606 ( .A1(n15521), .A2(n15522), .ZN(n15587) );
  NAND2_X1 U15607 ( .A1(n15591), .A2(n15592), .ZN(n15522) );
  NAND2_X1 U15608 ( .A1(n15519), .A2(n15593), .ZN(n15592) );
  INV_X1 U15609 ( .A(n15594), .ZN(n15593) );
  NOR2_X1 U15610 ( .A1(n15516), .A2(n15518), .ZN(n15594) );
  NOR2_X1 U15611 ( .A1(n8741), .A2(n15197), .ZN(n15519) );
  NAND2_X1 U15612 ( .A1(n15516), .A2(n15518), .ZN(n15591) );
  NAND2_X1 U15613 ( .A1(n15595), .A2(n15596), .ZN(n15518) );
  NAND2_X1 U15614 ( .A1(n15515), .A2(n15597), .ZN(n15596) );
  INV_X1 U15615 ( .A(n15598), .ZN(n15597) );
  NOR2_X1 U15616 ( .A1(n15514), .A2(n15513), .ZN(n15598) );
  NOR2_X1 U15617 ( .A1(n8452), .A2(n15197), .ZN(n15515) );
  NAND2_X1 U15618 ( .A1(n15513), .A2(n15514), .ZN(n15595) );
  NAND2_X1 U15619 ( .A1(n15599), .A2(n15600), .ZN(n15514) );
  NAND2_X1 U15620 ( .A1(n15511), .A2(n15601), .ZN(n15600) );
  INV_X1 U15621 ( .A(n15602), .ZN(n15601) );
  NOR2_X1 U15622 ( .A1(n15508), .A2(n15510), .ZN(n15602) );
  NOR2_X1 U15623 ( .A1(n8750), .A2(n15197), .ZN(n15511) );
  NAND2_X1 U15624 ( .A1(n15508), .A2(n15510), .ZN(n15599) );
  NAND2_X1 U15625 ( .A1(n15603), .A2(n15604), .ZN(n15510) );
  NAND2_X1 U15626 ( .A1(n15506), .A2(n15605), .ZN(n15604) );
  INV_X1 U15627 ( .A(n15606), .ZN(n15605) );
  NOR2_X1 U15628 ( .A1(n15507), .A2(n15505), .ZN(n15606) );
  NOR2_X1 U15629 ( .A1(n8443), .A2(n15197), .ZN(n15506) );
  NAND2_X1 U15630 ( .A1(n15505), .A2(n15507), .ZN(n15603) );
  NAND2_X1 U15631 ( .A1(n15607), .A2(n15608), .ZN(n15507) );
  NAND2_X1 U15632 ( .A1(n15503), .A2(n15609), .ZN(n15608) );
  INV_X1 U15633 ( .A(n15610), .ZN(n15609) );
  NOR2_X1 U15634 ( .A1(n15502), .A2(n15500), .ZN(n15610) );
  NOR2_X1 U15635 ( .A1(n8438), .A2(n15197), .ZN(n15503) );
  NAND2_X1 U15636 ( .A1(n15500), .A2(n15502), .ZN(n15607) );
  NAND2_X1 U15637 ( .A1(n15611), .A2(n15612), .ZN(n15502) );
  NAND2_X1 U15638 ( .A1(n15499), .A2(n15613), .ZN(n15612) );
  INV_X1 U15639 ( .A(n15614), .ZN(n15613) );
  NOR2_X1 U15640 ( .A1(n15498), .A2(n15497), .ZN(n15614) );
  NOR2_X1 U15641 ( .A1(n8763), .A2(n15197), .ZN(n15499) );
  NAND2_X1 U15642 ( .A1(n15497), .A2(n15498), .ZN(n15611) );
  NAND2_X1 U15643 ( .A1(n15615), .A2(n15616), .ZN(n15498) );
  NAND2_X1 U15644 ( .A1(n15495), .A2(n15617), .ZN(n15616) );
  INV_X1 U15645 ( .A(n15618), .ZN(n15617) );
  NOR2_X1 U15646 ( .A1(n15492), .A2(n15494), .ZN(n15618) );
  NOR2_X1 U15647 ( .A1(n8768), .A2(n15197), .ZN(n15495) );
  NAND2_X1 U15648 ( .A1(n15492), .A2(n15494), .ZN(n15615) );
  NAND2_X1 U15649 ( .A1(n15619), .A2(n15620), .ZN(n15494) );
  NAND2_X1 U15650 ( .A1(n15491), .A2(n15621), .ZN(n15620) );
  INV_X1 U15651 ( .A(n15622), .ZN(n15621) );
  NOR2_X1 U15652 ( .A1(n15490), .A2(n15489), .ZN(n15622) );
  NOR2_X1 U15653 ( .A1(n8772), .A2(n15197), .ZN(n15491) );
  NAND2_X1 U15654 ( .A1(n15489), .A2(n15490), .ZN(n15619) );
  NAND2_X1 U15655 ( .A1(n15623), .A2(n15624), .ZN(n15490) );
  NAND2_X1 U15656 ( .A1(n15487), .A2(n15625), .ZN(n15624) );
  INV_X1 U15657 ( .A(n15626), .ZN(n15625) );
  NOR2_X1 U15658 ( .A1(n15484), .A2(n15486), .ZN(n15626) );
  NOR2_X1 U15659 ( .A1(n10616), .A2(n15197), .ZN(n15487) );
  NAND2_X1 U15660 ( .A1(n15484), .A2(n15486), .ZN(n15623) );
  NAND2_X1 U15661 ( .A1(n15627), .A2(n15628), .ZN(n15486) );
  NAND2_X1 U15662 ( .A1(n15483), .A2(n15629), .ZN(n15628) );
  INV_X1 U15663 ( .A(n15630), .ZN(n15629) );
  NOR2_X1 U15664 ( .A1(n15482), .A2(n15481), .ZN(n15630) );
  NOR2_X1 U15665 ( .A1(n15197), .A2(n8881), .ZN(n15483) );
  NAND2_X1 U15666 ( .A1(n15481), .A2(n15482), .ZN(n15627) );
  NAND2_X1 U15667 ( .A1(n15631), .A2(n15632), .ZN(n15482) );
  NAND2_X1 U15668 ( .A1(n15479), .A2(n15633), .ZN(n15632) );
  INV_X1 U15669 ( .A(n15634), .ZN(n15633) );
  NOR2_X1 U15670 ( .A1(n15476), .A2(n15478), .ZN(n15634) );
  NOR2_X1 U15671 ( .A1(n15197), .A2(n10633), .ZN(n15479) );
  NAND2_X1 U15672 ( .A1(n15476), .A2(n15478), .ZN(n15631) );
  NAND2_X1 U15673 ( .A1(n15635), .A2(n15636), .ZN(n15478) );
  NAND2_X1 U15674 ( .A1(n15475), .A2(n15637), .ZN(n15636) );
  INV_X1 U15675 ( .A(n15638), .ZN(n15637) );
  NOR2_X1 U15676 ( .A1(n15474), .A2(n15473), .ZN(n15638) );
  NOR2_X1 U15677 ( .A1(n15197), .A2(n8798), .ZN(n15475) );
  NAND2_X1 U15678 ( .A1(n15473), .A2(n15474), .ZN(n15635) );
  NAND2_X1 U15679 ( .A1(n15639), .A2(n15640), .ZN(n15474) );
  NAND2_X1 U15680 ( .A1(n15471), .A2(n15641), .ZN(n15640) );
  INV_X1 U15681 ( .A(n15642), .ZN(n15641) );
  NOR2_X1 U15682 ( .A1(n15470), .A2(n15468), .ZN(n15642) );
  NOR2_X1 U15683 ( .A1(n15197), .A2(n8803), .ZN(n15471) );
  NAND2_X1 U15684 ( .A1(n15468), .A2(n15470), .ZN(n15639) );
  NAND2_X1 U15685 ( .A1(n15643), .A2(n15644), .ZN(n15470) );
  NAND2_X1 U15686 ( .A1(n15466), .A2(n15645), .ZN(n15644) );
  NAND2_X1 U15687 ( .A1(n15465), .A2(n15467), .ZN(n15645) );
  NOR2_X1 U15688 ( .A1(n15197), .A2(n8812), .ZN(n15466) );
  INV_X1 U15689 ( .A(n15646), .ZN(n15643) );
  NOR2_X1 U15690 ( .A1(n15465), .A2(n15467), .ZN(n15646) );
  NOR2_X1 U15691 ( .A1(n15647), .A2(n15648), .ZN(n15467) );
  NOR2_X1 U15692 ( .A1(n15463), .A2(n15649), .ZN(n15648) );
  NOR2_X1 U15693 ( .A1(n15460), .A2(n15462), .ZN(n15649) );
  NAND2_X1 U15694 ( .A1(b_4_), .A2(a_24_), .ZN(n15463) );
  INV_X1 U15695 ( .A(n15650), .ZN(n15647) );
  NAND2_X1 U15696 ( .A1(n15460), .A2(n15462), .ZN(n15650) );
  NAND2_X1 U15697 ( .A1(n15651), .A2(n15652), .ZN(n15462) );
  NAND2_X1 U15698 ( .A1(n15459), .A2(n15653), .ZN(n15652) );
  NAND2_X1 U15699 ( .A1(n15456), .A2(n15458), .ZN(n15653) );
  NOR2_X1 U15700 ( .A1(n15197), .A2(n8825), .ZN(n15459) );
  INV_X1 U15701 ( .A(n15654), .ZN(n15651) );
  NOR2_X1 U15702 ( .A1(n15458), .A2(n15456), .ZN(n15654) );
  XOR2_X1 U15703 ( .A(n15655), .B(n15656), .Z(n15456) );
  XOR2_X1 U15704 ( .A(n15657), .B(n15658), .Z(n15655) );
  NAND2_X1 U15705 ( .A1(n15659), .A2(n15660), .ZN(n15458) );
  NAND2_X1 U15706 ( .A1(n15416), .A2(n15661), .ZN(n15660) );
  NAND2_X1 U15707 ( .A1(n15418), .A2(n15417), .ZN(n15661) );
  XOR2_X1 U15708 ( .A(n15662), .B(n15663), .Z(n15416) );
  NAND2_X1 U15709 ( .A1(n15664), .A2(n15665), .ZN(n15662) );
  INV_X1 U15710 ( .A(n15666), .ZN(n15659) );
  NOR2_X1 U15711 ( .A1(n15417), .A2(n15418), .ZN(n15666) );
  NOR2_X1 U15712 ( .A1(n15197), .A2(n8830), .ZN(n15418) );
  NAND2_X1 U15713 ( .A1(n15424), .A2(n15667), .ZN(n15417) );
  NAND2_X1 U15714 ( .A1(n15423), .A2(n15425), .ZN(n15667) );
  NAND2_X1 U15715 ( .A1(n15668), .A2(n15669), .ZN(n15425) );
  NAND2_X1 U15716 ( .A1(b_4_), .A2(a_27_), .ZN(n15669) );
  XOR2_X1 U15717 ( .A(n15670), .B(n15671), .Z(n15423) );
  XNOR2_X1 U15718 ( .A(n15672), .B(n15673), .ZN(n15670) );
  NAND2_X1 U15719 ( .A1(b_3_), .A2(a_28_), .ZN(n15672) );
  INV_X1 U15720 ( .A(n15674), .ZN(n15424) );
  NOR2_X1 U15721 ( .A1(n8839), .A2(n15668), .ZN(n15674) );
  NOR2_X1 U15722 ( .A1(n15675), .A2(n15676), .ZN(n15668) );
  INV_X1 U15723 ( .A(n15677), .ZN(n15676) );
  NAND2_X1 U15724 ( .A1(n15454), .A2(n15678), .ZN(n15677) );
  NAND2_X1 U15725 ( .A1(n15455), .A2(n15453), .ZN(n15678) );
  NOR2_X1 U15726 ( .A1(n15197), .A2(n8844), .ZN(n15454) );
  NOR2_X1 U15727 ( .A1(n15453), .A2(n15455), .ZN(n15675) );
  NOR2_X1 U15728 ( .A1(n15679), .A2(n15680), .ZN(n15455) );
  INV_X1 U15729 ( .A(n15681), .ZN(n15680) );
  NAND2_X1 U15730 ( .A1(n15448), .A2(n15682), .ZN(n15681) );
  NAND2_X1 U15731 ( .A1(n15683), .A2(n15450), .ZN(n15682) );
  NOR2_X1 U15732 ( .A1(n15197), .A2(n9161), .ZN(n15448) );
  NOR2_X1 U15733 ( .A1(n15450), .A2(n15683), .ZN(n15679) );
  INV_X1 U15734 ( .A(n15451), .ZN(n15683) );
  NAND2_X1 U15735 ( .A1(n15684), .A2(n15685), .ZN(n15451) );
  NAND2_X1 U15736 ( .A1(b_2_), .A2(n15686), .ZN(n15685) );
  NAND2_X1 U15737 ( .A1(n8358), .A2(n15687), .ZN(n15686) );
  NAND2_X1 U15738 ( .A1(a_31_), .A2(n15446), .ZN(n15687) );
  NAND2_X1 U15739 ( .A1(b_3_), .A2(n15688), .ZN(n15684) );
  NAND2_X1 U15740 ( .A1(n8362), .A2(n15689), .ZN(n15688) );
  NAND2_X1 U15741 ( .A1(a_30_), .A2(n15690), .ZN(n15689) );
  NAND2_X1 U15742 ( .A1(n15691), .A2(b_3_), .ZN(n15450) );
  NOR2_X1 U15743 ( .A1(n9170), .A2(n15197), .ZN(n15691) );
  XOR2_X1 U15744 ( .A(n15692), .B(n15693), .Z(n15453) );
  XNOR2_X1 U15745 ( .A(n15694), .B(n15695), .ZN(n15693) );
  XNOR2_X1 U15746 ( .A(n15696), .B(n15697), .ZN(n15460) );
  XNOR2_X1 U15747 ( .A(n15698), .B(n15699), .ZN(n15697) );
  XOR2_X1 U15748 ( .A(n15700), .B(n15701), .Z(n15465) );
  XNOR2_X1 U15749 ( .A(n15702), .B(n15703), .ZN(n15700) );
  XNOR2_X1 U15750 ( .A(n15704), .B(n15705), .ZN(n15468) );
  NAND2_X1 U15751 ( .A1(n15706), .A2(n15707), .ZN(n15704) );
  XOR2_X1 U15752 ( .A(n15708), .B(n15709), .Z(n15473) );
  XOR2_X1 U15753 ( .A(n15710), .B(n15711), .Z(n15708) );
  NOR2_X1 U15754 ( .A1(n8803), .A2(n15446), .ZN(n15711) );
  XNOR2_X1 U15755 ( .A(n15712), .B(n15713), .ZN(n15476) );
  NAND2_X1 U15756 ( .A1(n15714), .A2(n15715), .ZN(n15712) );
  XOR2_X1 U15757 ( .A(n15716), .B(n15717), .Z(n15481) );
  XOR2_X1 U15758 ( .A(n15718), .B(n15719), .Z(n15716) );
  NOR2_X1 U15759 ( .A1(n10633), .A2(n15446), .ZN(n15719) );
  XNOR2_X1 U15760 ( .A(n15720), .B(n15721), .ZN(n15484) );
  NAND2_X1 U15761 ( .A1(n15722), .A2(n15723), .ZN(n15720) );
  XOR2_X1 U15762 ( .A(n15724), .B(n15725), .Z(n15489) );
  XOR2_X1 U15763 ( .A(n15726), .B(n15727), .Z(n15724) );
  NOR2_X1 U15764 ( .A1(n15446), .A2(n10616), .ZN(n15727) );
  XNOR2_X1 U15765 ( .A(n15728), .B(n15729), .ZN(n15492) );
  NAND2_X1 U15766 ( .A1(n15730), .A2(n15731), .ZN(n15728) );
  XOR2_X1 U15767 ( .A(n15732), .B(n15733), .Z(n15497) );
  XOR2_X1 U15768 ( .A(n15734), .B(n15735), .Z(n15732) );
  NOR2_X1 U15769 ( .A1(n15446), .A2(n8768), .ZN(n15735) );
  XNOR2_X1 U15770 ( .A(n15736), .B(n15737), .ZN(n15500) );
  NAND2_X1 U15771 ( .A1(n15738), .A2(n15739), .ZN(n15736) );
  XOR2_X1 U15772 ( .A(n15740), .B(n15741), .Z(n15505) );
  XOR2_X1 U15773 ( .A(n15742), .B(n15743), .Z(n15740) );
  NOR2_X1 U15774 ( .A1(n15446), .A2(n8438), .ZN(n15743) );
  XNOR2_X1 U15775 ( .A(n15744), .B(n15745), .ZN(n15508) );
  NAND2_X1 U15776 ( .A1(n15746), .A2(n15747), .ZN(n15744) );
  XOR2_X1 U15777 ( .A(n15748), .B(n15749), .Z(n15513) );
  XOR2_X1 U15778 ( .A(n15750), .B(n15751), .Z(n15748) );
  NOR2_X1 U15779 ( .A1(n15446), .A2(n8750), .ZN(n15751) );
  XNOR2_X1 U15780 ( .A(n15752), .B(n15753), .ZN(n15516) );
  NAND2_X1 U15781 ( .A1(n15754), .A2(n15755), .ZN(n15752) );
  XOR2_X1 U15782 ( .A(n15756), .B(n15757), .Z(n15521) );
  XOR2_X1 U15783 ( .A(n15758), .B(n15759), .Z(n15756) );
  NOR2_X1 U15784 ( .A1(n15446), .A2(n8741), .ZN(n15759) );
  XNOR2_X1 U15785 ( .A(n15760), .B(n15761), .ZN(n15524) );
  NAND2_X1 U15786 ( .A1(n15762), .A2(n15763), .ZN(n15760) );
  XOR2_X1 U15787 ( .A(n15764), .B(n15765), .Z(n15529) );
  XOR2_X1 U15788 ( .A(n15766), .B(n15767), .Z(n15764) );
  NOR2_X1 U15789 ( .A1(n15446), .A2(n8731), .ZN(n15767) );
  XNOR2_X1 U15790 ( .A(n15768), .B(n15769), .ZN(n15331) );
  NAND2_X1 U15791 ( .A1(n15770), .A2(n15771), .ZN(n15768) );
  XOR2_X1 U15792 ( .A(n15772), .B(n15773), .Z(n15324) );
  XOR2_X1 U15793 ( .A(n15774), .B(n15775), .Z(n15772) );
  NOR2_X1 U15794 ( .A1(n15446), .A2(n8480), .ZN(n15775) );
  XNOR2_X1 U15795 ( .A(n15776), .B(n15777), .ZN(n15532) );
  NAND2_X1 U15796 ( .A1(n15778), .A2(n15779), .ZN(n15776) );
  XOR2_X1 U15797 ( .A(n15780), .B(n15781), .Z(n15537) );
  XOR2_X1 U15798 ( .A(n15782), .B(n15783), .Z(n15780) );
  NOR2_X1 U15799 ( .A1(n15446), .A2(n8712), .ZN(n15783) );
  XNOR2_X1 U15800 ( .A(n15784), .B(n15785), .ZN(n15540) );
  XOR2_X1 U15801 ( .A(n15786), .B(n15787), .Z(n15784) );
  XOR2_X1 U15802 ( .A(n15788), .B(n15789), .Z(n15544) );
  XNOR2_X1 U15803 ( .A(n15790), .B(n15791), .ZN(n15789) );
  NAND2_X1 U15804 ( .A1(a_2_), .A2(b_3_), .ZN(n15791) );
  XNOR2_X1 U15805 ( .A(n15792), .B(n15793), .ZN(n15300) );
  NAND2_X1 U15806 ( .A1(n15794), .A2(n15795), .ZN(n15792) );
  XOR2_X1 U15807 ( .A(n15796), .B(n15797), .Z(n15549) );
  XOR2_X1 U15808 ( .A(n15798), .B(n15799), .Z(n15796) );
  NOR2_X1 U15809 ( .A1(n15446), .A2(n8690), .ZN(n15799) );
  NOR2_X1 U15810 ( .A1(n15800), .A2(n8612), .ZN(n8470) );
  INV_X1 U15811 ( .A(n15801), .ZN(n8612) );
  NAND2_X1 U15812 ( .A1(n15802), .A2(n15803), .ZN(n15801) );
  NOR2_X1 U15813 ( .A1(n15802), .A2(n15803), .ZN(n15800) );
  NAND2_X1 U15814 ( .A1(n15804), .A2(n15805), .ZN(n15803) );
  NAND2_X1 U15815 ( .A1(n15806), .A2(a_0_), .ZN(n15805) );
  NOR2_X1 U15816 ( .A1(n15807), .A2(n15446), .ZN(n15806) );
  NOR2_X1 U15817 ( .A1(n15797), .A2(n15798), .ZN(n15807) );
  NAND2_X1 U15818 ( .A1(n15797), .A2(n15798), .ZN(n15804) );
  NAND2_X1 U15819 ( .A1(n15794), .A2(n15808), .ZN(n15798) );
  NAND2_X1 U15820 ( .A1(n15793), .A2(n15795), .ZN(n15808) );
  NAND2_X1 U15821 ( .A1(n15809), .A2(n15810), .ZN(n15795) );
  NAND2_X1 U15822 ( .A1(a_1_), .A2(b_3_), .ZN(n15810) );
  INV_X1 U15823 ( .A(n15811), .ZN(n15809) );
  XNOR2_X1 U15824 ( .A(n15812), .B(n15813), .ZN(n15793) );
  XOR2_X1 U15825 ( .A(n15814), .B(n15815), .Z(n15813) );
  NAND2_X1 U15826 ( .A1(a_1_), .A2(n15811), .ZN(n15794) );
  NAND2_X1 U15827 ( .A1(n15816), .A2(n15817), .ZN(n15811) );
  NAND2_X1 U15828 ( .A1(n15818), .A2(a_2_), .ZN(n15817) );
  NOR2_X1 U15829 ( .A1(n15819), .A2(n15446), .ZN(n15818) );
  NOR2_X1 U15830 ( .A1(n15790), .A2(n15788), .ZN(n15819) );
  NAND2_X1 U15831 ( .A1(n15790), .A2(n15788), .ZN(n15816) );
  XNOR2_X1 U15832 ( .A(n15820), .B(n15821), .ZN(n15788) );
  XNOR2_X1 U15833 ( .A(n15822), .B(n15823), .ZN(n15820) );
  NOR2_X1 U15834 ( .A1(n15824), .A2(n15825), .ZN(n15790) );
  INV_X1 U15835 ( .A(n15826), .ZN(n15825) );
  NAND2_X1 U15836 ( .A1(n15785), .A2(n15827), .ZN(n15826) );
  NAND2_X1 U15837 ( .A1(n15787), .A2(n15786), .ZN(n15827) );
  XNOR2_X1 U15838 ( .A(n15828), .B(n15829), .ZN(n15785) );
  XOR2_X1 U15839 ( .A(n15830), .B(n15831), .Z(n15829) );
  NOR2_X1 U15840 ( .A1(n15786), .A2(n15787), .ZN(n15824) );
  NAND2_X1 U15841 ( .A1(n15832), .A2(n15833), .ZN(n15786) );
  NAND2_X1 U15842 ( .A1(n15834), .A2(a_4_), .ZN(n15833) );
  NOR2_X1 U15843 ( .A1(n15835), .A2(n15446), .ZN(n15834) );
  NOR2_X1 U15844 ( .A1(n15782), .A2(n15781), .ZN(n15835) );
  NAND2_X1 U15845 ( .A1(n15781), .A2(n15782), .ZN(n15832) );
  NAND2_X1 U15846 ( .A1(n15778), .A2(n15836), .ZN(n15782) );
  NAND2_X1 U15847 ( .A1(n15777), .A2(n15779), .ZN(n15836) );
  NAND2_X1 U15848 ( .A1(n15837), .A2(n15838), .ZN(n15779) );
  NAND2_X1 U15849 ( .A1(a_5_), .A2(b_3_), .ZN(n15838) );
  INV_X1 U15850 ( .A(n15839), .ZN(n15837) );
  XNOR2_X1 U15851 ( .A(n15840), .B(n15841), .ZN(n15777) );
  XNOR2_X1 U15852 ( .A(n15842), .B(n15843), .ZN(n15841) );
  NAND2_X1 U15853 ( .A1(a_5_), .A2(n15839), .ZN(n15778) );
  NAND2_X1 U15854 ( .A1(n15844), .A2(n15845), .ZN(n15839) );
  NAND2_X1 U15855 ( .A1(n15846), .A2(a_6_), .ZN(n15845) );
  NOR2_X1 U15856 ( .A1(n15847), .A2(n15446), .ZN(n15846) );
  NOR2_X1 U15857 ( .A1(n15774), .A2(n15773), .ZN(n15847) );
  NAND2_X1 U15858 ( .A1(n15773), .A2(n15774), .ZN(n15844) );
  NAND2_X1 U15859 ( .A1(n15770), .A2(n15848), .ZN(n15774) );
  NAND2_X1 U15860 ( .A1(n15769), .A2(n15771), .ZN(n15848) );
  NAND2_X1 U15861 ( .A1(n15849), .A2(n15850), .ZN(n15771) );
  NAND2_X1 U15862 ( .A1(a_7_), .A2(b_3_), .ZN(n15850) );
  INV_X1 U15863 ( .A(n15851), .ZN(n15849) );
  XNOR2_X1 U15864 ( .A(n15852), .B(n15853), .ZN(n15769) );
  XNOR2_X1 U15865 ( .A(n15854), .B(n15855), .ZN(n15853) );
  NAND2_X1 U15866 ( .A1(a_7_), .A2(n15851), .ZN(n15770) );
  NAND2_X1 U15867 ( .A1(n15856), .A2(n15857), .ZN(n15851) );
  NAND2_X1 U15868 ( .A1(n15858), .A2(a_8_), .ZN(n15857) );
  NOR2_X1 U15869 ( .A1(n15859), .A2(n15446), .ZN(n15858) );
  NOR2_X1 U15870 ( .A1(n15766), .A2(n15765), .ZN(n15859) );
  NAND2_X1 U15871 ( .A1(n15765), .A2(n15766), .ZN(n15856) );
  NAND2_X1 U15872 ( .A1(n15762), .A2(n15860), .ZN(n15766) );
  NAND2_X1 U15873 ( .A1(n15761), .A2(n15763), .ZN(n15860) );
  NAND2_X1 U15874 ( .A1(n15861), .A2(n15862), .ZN(n15763) );
  NAND2_X1 U15875 ( .A1(a_9_), .A2(b_3_), .ZN(n15862) );
  INV_X1 U15876 ( .A(n15863), .ZN(n15861) );
  XNOR2_X1 U15877 ( .A(n15864), .B(n15865), .ZN(n15761) );
  XNOR2_X1 U15878 ( .A(n15866), .B(n15867), .ZN(n15865) );
  NAND2_X1 U15879 ( .A1(a_9_), .A2(n15863), .ZN(n15762) );
  NAND2_X1 U15880 ( .A1(n15868), .A2(n15869), .ZN(n15863) );
  NAND2_X1 U15881 ( .A1(n15870), .A2(a_10_), .ZN(n15869) );
  NOR2_X1 U15882 ( .A1(n15871), .A2(n15446), .ZN(n15870) );
  NOR2_X1 U15883 ( .A1(n15758), .A2(n15757), .ZN(n15871) );
  NAND2_X1 U15884 ( .A1(n15757), .A2(n15758), .ZN(n15868) );
  NAND2_X1 U15885 ( .A1(n15754), .A2(n15872), .ZN(n15758) );
  NAND2_X1 U15886 ( .A1(n15753), .A2(n15755), .ZN(n15872) );
  NAND2_X1 U15887 ( .A1(n15873), .A2(n15874), .ZN(n15755) );
  NAND2_X1 U15888 ( .A1(a_11_), .A2(b_3_), .ZN(n15874) );
  INV_X1 U15889 ( .A(n15875), .ZN(n15873) );
  XNOR2_X1 U15890 ( .A(n15876), .B(n15877), .ZN(n15753) );
  XNOR2_X1 U15891 ( .A(n15878), .B(n15879), .ZN(n15877) );
  NAND2_X1 U15892 ( .A1(a_11_), .A2(n15875), .ZN(n15754) );
  NAND2_X1 U15893 ( .A1(n15880), .A2(n15881), .ZN(n15875) );
  NAND2_X1 U15894 ( .A1(n15882), .A2(a_12_), .ZN(n15881) );
  NOR2_X1 U15895 ( .A1(n15883), .A2(n15446), .ZN(n15882) );
  NOR2_X1 U15896 ( .A1(n15750), .A2(n15749), .ZN(n15883) );
  NAND2_X1 U15897 ( .A1(n15749), .A2(n15750), .ZN(n15880) );
  NAND2_X1 U15898 ( .A1(n15746), .A2(n15884), .ZN(n15750) );
  NAND2_X1 U15899 ( .A1(n15745), .A2(n15747), .ZN(n15884) );
  NAND2_X1 U15900 ( .A1(n15885), .A2(n15886), .ZN(n15747) );
  NAND2_X1 U15901 ( .A1(a_13_), .A2(b_3_), .ZN(n15886) );
  INV_X1 U15902 ( .A(n15887), .ZN(n15885) );
  XNOR2_X1 U15903 ( .A(n15888), .B(n15889), .ZN(n15745) );
  XNOR2_X1 U15904 ( .A(n15890), .B(n15891), .ZN(n15889) );
  NAND2_X1 U15905 ( .A1(a_13_), .A2(n15887), .ZN(n15746) );
  NAND2_X1 U15906 ( .A1(n15892), .A2(n15893), .ZN(n15887) );
  NAND2_X1 U15907 ( .A1(n15894), .A2(a_14_), .ZN(n15893) );
  NOR2_X1 U15908 ( .A1(n15895), .A2(n15446), .ZN(n15894) );
  NOR2_X1 U15909 ( .A1(n15742), .A2(n15741), .ZN(n15895) );
  NAND2_X1 U15910 ( .A1(n15741), .A2(n15742), .ZN(n15892) );
  NAND2_X1 U15911 ( .A1(n15738), .A2(n15896), .ZN(n15742) );
  NAND2_X1 U15912 ( .A1(n15737), .A2(n15739), .ZN(n15896) );
  NAND2_X1 U15913 ( .A1(n15897), .A2(n15898), .ZN(n15739) );
  NAND2_X1 U15914 ( .A1(a_15_), .A2(b_3_), .ZN(n15898) );
  INV_X1 U15915 ( .A(n15899), .ZN(n15897) );
  XNOR2_X1 U15916 ( .A(n15900), .B(n15901), .ZN(n15737) );
  XNOR2_X1 U15917 ( .A(n15902), .B(n15903), .ZN(n15900) );
  NAND2_X1 U15918 ( .A1(a_15_), .A2(n15899), .ZN(n15738) );
  NAND2_X1 U15919 ( .A1(n15904), .A2(n15905), .ZN(n15899) );
  NAND2_X1 U15920 ( .A1(n15906), .A2(a_16_), .ZN(n15905) );
  NOR2_X1 U15921 ( .A1(n15907), .A2(n15446), .ZN(n15906) );
  NOR2_X1 U15922 ( .A1(n15734), .A2(n15733), .ZN(n15907) );
  NAND2_X1 U15923 ( .A1(n15733), .A2(n15734), .ZN(n15904) );
  NAND2_X1 U15924 ( .A1(n15730), .A2(n15908), .ZN(n15734) );
  NAND2_X1 U15925 ( .A1(n15729), .A2(n15731), .ZN(n15908) );
  NAND2_X1 U15926 ( .A1(n15909), .A2(n15910), .ZN(n15731) );
  NAND2_X1 U15927 ( .A1(a_17_), .A2(b_3_), .ZN(n15910) );
  INV_X1 U15928 ( .A(n15911), .ZN(n15909) );
  XNOR2_X1 U15929 ( .A(n15912), .B(n15913), .ZN(n15729) );
  XNOR2_X1 U15930 ( .A(n15914), .B(n15915), .ZN(n15912) );
  NAND2_X1 U15931 ( .A1(a_17_), .A2(n15911), .ZN(n15730) );
  NAND2_X1 U15932 ( .A1(n15916), .A2(n15917), .ZN(n15911) );
  NAND2_X1 U15933 ( .A1(n15918), .A2(a_18_), .ZN(n15917) );
  NOR2_X1 U15934 ( .A1(n15919), .A2(n15446), .ZN(n15918) );
  NOR2_X1 U15935 ( .A1(n15726), .A2(n15725), .ZN(n15919) );
  NAND2_X1 U15936 ( .A1(n15725), .A2(n15726), .ZN(n15916) );
  NAND2_X1 U15937 ( .A1(n15722), .A2(n15920), .ZN(n15726) );
  NAND2_X1 U15938 ( .A1(n15721), .A2(n15723), .ZN(n15920) );
  NAND2_X1 U15939 ( .A1(n15921), .A2(n15922), .ZN(n15723) );
  NAND2_X1 U15940 ( .A1(b_3_), .A2(a_19_), .ZN(n15922) );
  INV_X1 U15941 ( .A(n15923), .ZN(n15921) );
  XNOR2_X1 U15942 ( .A(n15924), .B(n15925), .ZN(n15721) );
  XNOR2_X1 U15943 ( .A(n15926), .B(n15927), .ZN(n15924) );
  NAND2_X1 U15944 ( .A1(a_19_), .A2(n15923), .ZN(n15722) );
  NAND2_X1 U15945 ( .A1(n15928), .A2(n15929), .ZN(n15923) );
  NAND2_X1 U15946 ( .A1(n15930), .A2(b_3_), .ZN(n15929) );
  NOR2_X1 U15947 ( .A1(n15931), .A2(n10633), .ZN(n15930) );
  NOR2_X1 U15948 ( .A1(n15718), .A2(n15717), .ZN(n15931) );
  NAND2_X1 U15949 ( .A1(n15717), .A2(n15718), .ZN(n15928) );
  NAND2_X1 U15950 ( .A1(n15714), .A2(n15932), .ZN(n15718) );
  NAND2_X1 U15951 ( .A1(n15713), .A2(n15715), .ZN(n15932) );
  NAND2_X1 U15952 ( .A1(n15933), .A2(n15934), .ZN(n15715) );
  NAND2_X1 U15953 ( .A1(b_3_), .A2(a_21_), .ZN(n15934) );
  INV_X1 U15954 ( .A(n15935), .ZN(n15933) );
  XNOR2_X1 U15955 ( .A(n15936), .B(n15937), .ZN(n15713) );
  XNOR2_X1 U15956 ( .A(n15938), .B(n15939), .ZN(n15936) );
  NAND2_X1 U15957 ( .A1(a_21_), .A2(n15935), .ZN(n15714) );
  NAND2_X1 U15958 ( .A1(n15940), .A2(n15941), .ZN(n15935) );
  NAND2_X1 U15959 ( .A1(n15942), .A2(b_3_), .ZN(n15941) );
  NOR2_X1 U15960 ( .A1(n15943), .A2(n8803), .ZN(n15942) );
  NOR2_X1 U15961 ( .A1(n15710), .A2(n15709), .ZN(n15943) );
  NAND2_X1 U15962 ( .A1(n15709), .A2(n15710), .ZN(n15940) );
  NAND2_X1 U15963 ( .A1(n15706), .A2(n15944), .ZN(n15710) );
  NAND2_X1 U15964 ( .A1(n15705), .A2(n15707), .ZN(n15944) );
  NAND2_X1 U15965 ( .A1(n15945), .A2(n15946), .ZN(n15707) );
  NAND2_X1 U15966 ( .A1(b_3_), .A2(a_23_), .ZN(n15946) );
  XNOR2_X1 U15967 ( .A(n15947), .B(n15948), .ZN(n15705) );
  NAND2_X1 U15968 ( .A1(n15949), .A2(n15950), .ZN(n15947) );
  INV_X1 U15969 ( .A(n15951), .ZN(n15706) );
  NOR2_X1 U15970 ( .A1(n8812), .A2(n15945), .ZN(n15951) );
  NOR2_X1 U15971 ( .A1(n15952), .A2(n15953), .ZN(n15945) );
  INV_X1 U15972 ( .A(n15954), .ZN(n15953) );
  NAND2_X1 U15973 ( .A1(n15703), .A2(n15955), .ZN(n15954) );
  NAND2_X1 U15974 ( .A1(n15702), .A2(n15701), .ZN(n15955) );
  NOR2_X1 U15975 ( .A1(n15446), .A2(n9131), .ZN(n15703) );
  NOR2_X1 U15976 ( .A1(n15701), .A2(n15702), .ZN(n15952) );
  NOR2_X1 U15977 ( .A1(n15956), .A2(n15957), .ZN(n15702) );
  INV_X1 U15978 ( .A(n15958), .ZN(n15957) );
  NAND2_X1 U15979 ( .A1(n15699), .A2(n15959), .ZN(n15958) );
  NAND2_X1 U15980 ( .A1(n15696), .A2(n15698), .ZN(n15959) );
  NOR2_X1 U15981 ( .A1(n15446), .A2(n8825), .ZN(n15699) );
  NOR2_X1 U15982 ( .A1(n15698), .A2(n15696), .ZN(n15956) );
  XOR2_X1 U15983 ( .A(n15960), .B(n15961), .Z(n15696) );
  XOR2_X1 U15984 ( .A(n15962), .B(n15963), .Z(n15961) );
  NAND2_X1 U15985 ( .A1(b_2_), .A2(a_26_), .ZN(n15963) );
  NAND2_X1 U15986 ( .A1(n15964), .A2(n15965), .ZN(n15698) );
  NAND2_X1 U15987 ( .A1(n15656), .A2(n15966), .ZN(n15965) );
  NAND2_X1 U15988 ( .A1(n15658), .A2(n15657), .ZN(n15966) );
  XOR2_X1 U15989 ( .A(n15967), .B(n15968), .Z(n15656) );
  NAND2_X1 U15990 ( .A1(n15969), .A2(n15970), .ZN(n15967) );
  INV_X1 U15991 ( .A(n15971), .ZN(n15964) );
  NOR2_X1 U15992 ( .A1(n15657), .A2(n15658), .ZN(n15971) );
  NOR2_X1 U15993 ( .A1(n15446), .A2(n8830), .ZN(n15658) );
  NAND2_X1 U15994 ( .A1(n15664), .A2(n15972), .ZN(n15657) );
  NAND2_X1 U15995 ( .A1(n15663), .A2(n15665), .ZN(n15972) );
  NAND2_X1 U15996 ( .A1(n15973), .A2(n15974), .ZN(n15665) );
  NAND2_X1 U15997 ( .A1(b_3_), .A2(a_27_), .ZN(n15974) );
  INV_X1 U15998 ( .A(n15975), .ZN(n15973) );
  XOR2_X1 U15999 ( .A(n15976), .B(n15977), .Z(n15663) );
  XNOR2_X1 U16000 ( .A(n15978), .B(n15979), .ZN(n15976) );
  NAND2_X1 U16001 ( .A1(b_2_), .A2(a_28_), .ZN(n15978) );
  NAND2_X1 U16002 ( .A1(a_27_), .A2(n15975), .ZN(n15664) );
  NAND2_X1 U16003 ( .A1(n15980), .A2(n15981), .ZN(n15975) );
  NAND2_X1 U16004 ( .A1(n15982), .A2(b_3_), .ZN(n15981) );
  NOR2_X1 U16005 ( .A1(n15983), .A2(n8844), .ZN(n15982) );
  NOR2_X1 U16006 ( .A1(n15671), .A2(n15673), .ZN(n15983) );
  NAND2_X1 U16007 ( .A1(n15671), .A2(n15673), .ZN(n15980) );
  NAND2_X1 U16008 ( .A1(n15984), .A2(n15985), .ZN(n15673) );
  NAND2_X1 U16009 ( .A1(n15692), .A2(n15986), .ZN(n15985) );
  INV_X1 U16010 ( .A(n15987), .ZN(n15986) );
  NOR2_X1 U16011 ( .A1(n15695), .A2(n15694), .ZN(n15987) );
  NOR2_X1 U16012 ( .A1(n15446), .A2(n9161), .ZN(n15692) );
  NAND2_X1 U16013 ( .A1(n15694), .A2(n15695), .ZN(n15984) );
  NAND2_X1 U16014 ( .A1(n15988), .A2(n15989), .ZN(n15695) );
  NAND2_X1 U16015 ( .A1(b_1_), .A2(n15990), .ZN(n15989) );
  NAND2_X1 U16016 ( .A1(n8358), .A2(n15991), .ZN(n15990) );
  NAND2_X1 U16017 ( .A1(a_31_), .A2(n15690), .ZN(n15991) );
  NAND2_X1 U16018 ( .A1(b_2_), .A2(n15992), .ZN(n15988) );
  NAND2_X1 U16019 ( .A1(n8362), .A2(n15993), .ZN(n15992) );
  NAND2_X1 U16020 ( .A1(a_30_), .A2(n15994), .ZN(n15993) );
  NOR2_X1 U16021 ( .A1(n15995), .A2(n15690), .ZN(n15694) );
  NAND2_X1 U16022 ( .A1(n9926), .A2(b_3_), .ZN(n15995) );
  XNOR2_X1 U16023 ( .A(n15996), .B(n15997), .ZN(n15671) );
  XNOR2_X1 U16024 ( .A(n15998), .B(n15999), .ZN(n15997) );
  XOR2_X1 U16025 ( .A(n16000), .B(n16001), .Z(n15701) );
  NAND2_X1 U16026 ( .A1(n16002), .A2(n16003), .ZN(n16000) );
  XNOR2_X1 U16027 ( .A(n16004), .B(n16005), .ZN(n15709) );
  XOR2_X1 U16028 ( .A(n16006), .B(n16007), .Z(n16005) );
  XNOR2_X1 U16029 ( .A(n16008), .B(n16009), .ZN(n15717) );
  XNOR2_X1 U16030 ( .A(n16010), .B(n16011), .ZN(n16008) );
  XNOR2_X1 U16031 ( .A(n16012), .B(n16013), .ZN(n15725) );
  XNOR2_X1 U16032 ( .A(n16014), .B(n16015), .ZN(n16012) );
  XNOR2_X1 U16033 ( .A(n16016), .B(n16017), .ZN(n15733) );
  XNOR2_X1 U16034 ( .A(n16018), .B(n16019), .ZN(n16016) );
  XNOR2_X1 U16035 ( .A(n16020), .B(n16021), .ZN(n15741) );
  XNOR2_X1 U16036 ( .A(n16022), .B(n16023), .ZN(n16020) );
  XOR2_X1 U16037 ( .A(n16024), .B(n16025), .Z(n15749) );
  XOR2_X1 U16038 ( .A(n16026), .B(n16027), .Z(n16024) );
  XOR2_X1 U16039 ( .A(n16028), .B(n16029), .Z(n15757) );
  XOR2_X1 U16040 ( .A(n16030), .B(n16031), .Z(n16028) );
  XOR2_X1 U16041 ( .A(n16032), .B(n16033), .Z(n15765) );
  XOR2_X1 U16042 ( .A(n16034), .B(n16035), .Z(n16032) );
  XOR2_X1 U16043 ( .A(n16036), .B(n16037), .Z(n15773) );
  XOR2_X1 U16044 ( .A(n16038), .B(n16039), .Z(n16036) );
  XOR2_X1 U16045 ( .A(n16040), .B(n16041), .Z(n15781) );
  XOR2_X1 U16046 ( .A(n16042), .B(n16043), .Z(n16040) );
  XNOR2_X1 U16047 ( .A(n16044), .B(n16045), .ZN(n15797) );
  XNOR2_X1 U16048 ( .A(n16046), .B(n16047), .ZN(n16044) );
  XNOR2_X1 U16049 ( .A(n16048), .B(n16049), .ZN(n15802) );
  XNOR2_X1 U16050 ( .A(n16050), .B(n16051), .ZN(n16048) );
  XNOR2_X1 U16051 ( .A(n16052), .B(n16053), .ZN(n8514) );
  NOR2_X1 U16052 ( .A1(n16054), .A2(n16055), .ZN(n8560) );
  INV_X1 U16053 ( .A(n16056), .ZN(n16055) );
  XOR2_X1 U16054 ( .A(n8608), .B(n16057), .Z(n16054) );
  NOR2_X1 U16055 ( .A1(n16058), .A2(n16056), .ZN(n8561) );
  NAND2_X1 U16056 ( .A1(n16053), .A2(n16052), .ZN(n16056) );
  NAND2_X1 U16057 ( .A1(n16059), .A2(n16060), .ZN(n16052) );
  NAND2_X1 U16058 ( .A1(n16051), .A2(n16061), .ZN(n16060) );
  INV_X1 U16059 ( .A(n16062), .ZN(n16061) );
  NOR2_X1 U16060 ( .A1(n16050), .A2(n16049), .ZN(n16062) );
  NOR2_X1 U16061 ( .A1(n8690), .A2(n15690), .ZN(n16051) );
  NAND2_X1 U16062 ( .A1(n16049), .A2(n16050), .ZN(n16059) );
  NAND2_X1 U16063 ( .A1(n16063), .A2(n16064), .ZN(n16050) );
  NAND2_X1 U16064 ( .A1(n16047), .A2(n16065), .ZN(n16064) );
  INV_X1 U16065 ( .A(n16066), .ZN(n16065) );
  NOR2_X1 U16066 ( .A1(n16045), .A2(n16046), .ZN(n16066) );
  NOR2_X1 U16067 ( .A1(n8502), .A2(n15690), .ZN(n16047) );
  NAND2_X1 U16068 ( .A1(n16045), .A2(n16046), .ZN(n16063) );
  NOR2_X1 U16069 ( .A1(n16067), .A2(n16068), .ZN(n16046) );
  INV_X1 U16070 ( .A(n16069), .ZN(n16068) );
  NAND2_X1 U16071 ( .A1(n16070), .A2(n15815), .ZN(n16069) );
  NAND2_X1 U16072 ( .A1(n15812), .A2(n15814), .ZN(n16070) );
  NOR2_X1 U16073 ( .A1(n15814), .A2(n15812), .ZN(n16067) );
  XOR2_X1 U16074 ( .A(n16071), .B(n16072), .Z(n15812) );
  XOR2_X1 U16075 ( .A(n16073), .B(n16074), .Z(n16071) );
  NAND2_X1 U16076 ( .A1(n16075), .A2(n16076), .ZN(n15814) );
  NAND2_X1 U16077 ( .A1(n15822), .A2(n16077), .ZN(n16076) );
  NAND2_X1 U16078 ( .A1(n15823), .A2(n15821), .ZN(n16077) );
  NOR2_X1 U16079 ( .A1(n8707), .A2(n15690), .ZN(n15822) );
  INV_X1 U16080 ( .A(n16078), .ZN(n16075) );
  NOR2_X1 U16081 ( .A1(n15821), .A2(n15823), .ZN(n16078) );
  NOR2_X1 U16082 ( .A1(n16079), .A2(n16080), .ZN(n15823) );
  INV_X1 U16083 ( .A(n16081), .ZN(n16080) );
  NAND2_X1 U16084 ( .A1(n15831), .A2(n16082), .ZN(n16081) );
  NAND2_X1 U16085 ( .A1(n15830), .A2(n15828), .ZN(n16082) );
  NOR2_X1 U16086 ( .A1(n8712), .A2(n15690), .ZN(n15831) );
  NOR2_X1 U16087 ( .A1(n15828), .A2(n15830), .ZN(n16079) );
  INV_X1 U16088 ( .A(n16083), .ZN(n15830) );
  NAND2_X1 U16089 ( .A1(n16084), .A2(n16085), .ZN(n16083) );
  NAND2_X1 U16090 ( .A1(n16043), .A2(n16086), .ZN(n16085) );
  INV_X1 U16091 ( .A(n16087), .ZN(n16086) );
  NOR2_X1 U16092 ( .A1(n16042), .A2(n16041), .ZN(n16087) );
  NOR2_X1 U16093 ( .A1(n8717), .A2(n15690), .ZN(n16043) );
  NAND2_X1 U16094 ( .A1(n16041), .A2(n16042), .ZN(n16084) );
  NAND2_X1 U16095 ( .A1(n16088), .A2(n16089), .ZN(n16042) );
  NAND2_X1 U16096 ( .A1(n15843), .A2(n16090), .ZN(n16089) );
  INV_X1 U16097 ( .A(n16091), .ZN(n16090) );
  NOR2_X1 U16098 ( .A1(n15842), .A2(n15840), .ZN(n16091) );
  NOR2_X1 U16099 ( .A1(n8480), .A2(n15690), .ZN(n15843) );
  NAND2_X1 U16100 ( .A1(n15840), .A2(n15842), .ZN(n16088) );
  NAND2_X1 U16101 ( .A1(n16092), .A2(n16093), .ZN(n15842) );
  NAND2_X1 U16102 ( .A1(n16038), .A2(n16094), .ZN(n16093) );
  INV_X1 U16103 ( .A(n16095), .ZN(n16094) );
  NOR2_X1 U16104 ( .A1(n16039), .A2(n16037), .ZN(n16095) );
  NOR2_X1 U16105 ( .A1(n8726), .A2(n15690), .ZN(n16038) );
  NAND2_X1 U16106 ( .A1(n16037), .A2(n16039), .ZN(n16092) );
  NAND2_X1 U16107 ( .A1(n16096), .A2(n16097), .ZN(n16039) );
  NAND2_X1 U16108 ( .A1(n15855), .A2(n16098), .ZN(n16097) );
  INV_X1 U16109 ( .A(n16099), .ZN(n16098) );
  NOR2_X1 U16110 ( .A1(n15854), .A2(n15852), .ZN(n16099) );
  NOR2_X1 U16111 ( .A1(n8731), .A2(n15690), .ZN(n15855) );
  NAND2_X1 U16112 ( .A1(n15852), .A2(n15854), .ZN(n16096) );
  NAND2_X1 U16113 ( .A1(n16100), .A2(n16101), .ZN(n15854) );
  NAND2_X1 U16114 ( .A1(n16034), .A2(n16102), .ZN(n16101) );
  INV_X1 U16115 ( .A(n16103), .ZN(n16102) );
  NOR2_X1 U16116 ( .A1(n16035), .A2(n16033), .ZN(n16103) );
  NOR2_X1 U16117 ( .A1(n8736), .A2(n15690), .ZN(n16034) );
  NAND2_X1 U16118 ( .A1(n16033), .A2(n16035), .ZN(n16100) );
  NAND2_X1 U16119 ( .A1(n16104), .A2(n16105), .ZN(n16035) );
  NAND2_X1 U16120 ( .A1(n15867), .A2(n16106), .ZN(n16105) );
  INV_X1 U16121 ( .A(n16107), .ZN(n16106) );
  NOR2_X1 U16122 ( .A1(n15866), .A2(n15864), .ZN(n16107) );
  NOR2_X1 U16123 ( .A1(n8741), .A2(n15690), .ZN(n15867) );
  NAND2_X1 U16124 ( .A1(n15864), .A2(n15866), .ZN(n16104) );
  NAND2_X1 U16125 ( .A1(n16108), .A2(n16109), .ZN(n15866) );
  NAND2_X1 U16126 ( .A1(n16031), .A2(n16110), .ZN(n16109) );
  INV_X1 U16127 ( .A(n16111), .ZN(n16110) );
  NOR2_X1 U16128 ( .A1(n16030), .A2(n16029), .ZN(n16111) );
  NOR2_X1 U16129 ( .A1(n8452), .A2(n15690), .ZN(n16031) );
  NAND2_X1 U16130 ( .A1(n16029), .A2(n16030), .ZN(n16108) );
  NAND2_X1 U16131 ( .A1(n16112), .A2(n16113), .ZN(n16030) );
  NAND2_X1 U16132 ( .A1(n15879), .A2(n16114), .ZN(n16113) );
  INV_X1 U16133 ( .A(n16115), .ZN(n16114) );
  NOR2_X1 U16134 ( .A1(n15878), .A2(n15876), .ZN(n16115) );
  NOR2_X1 U16135 ( .A1(n8750), .A2(n15690), .ZN(n15879) );
  NAND2_X1 U16136 ( .A1(n15876), .A2(n15878), .ZN(n16112) );
  NAND2_X1 U16137 ( .A1(n16116), .A2(n16117), .ZN(n15878) );
  NAND2_X1 U16138 ( .A1(n16026), .A2(n16118), .ZN(n16117) );
  INV_X1 U16139 ( .A(n16119), .ZN(n16118) );
  NOR2_X1 U16140 ( .A1(n16027), .A2(n16025), .ZN(n16119) );
  NOR2_X1 U16141 ( .A1(n8443), .A2(n15690), .ZN(n16026) );
  NAND2_X1 U16142 ( .A1(n16025), .A2(n16027), .ZN(n16116) );
  NAND2_X1 U16143 ( .A1(n16120), .A2(n16121), .ZN(n16027) );
  NAND2_X1 U16144 ( .A1(n15891), .A2(n16122), .ZN(n16121) );
  INV_X1 U16145 ( .A(n16123), .ZN(n16122) );
  NOR2_X1 U16146 ( .A1(n15890), .A2(n15888), .ZN(n16123) );
  NOR2_X1 U16147 ( .A1(n8438), .A2(n15690), .ZN(n15891) );
  NAND2_X1 U16148 ( .A1(n15888), .A2(n15890), .ZN(n16120) );
  NAND2_X1 U16149 ( .A1(n16124), .A2(n16125), .ZN(n15890) );
  NAND2_X1 U16150 ( .A1(n16023), .A2(n16126), .ZN(n16125) );
  NAND2_X1 U16151 ( .A1(n16022), .A2(n16021), .ZN(n16126) );
  NOR2_X1 U16152 ( .A1(n8763), .A2(n15690), .ZN(n16023) );
  INV_X1 U16153 ( .A(n16127), .ZN(n16124) );
  NOR2_X1 U16154 ( .A1(n16021), .A2(n16022), .ZN(n16127) );
  NOR2_X1 U16155 ( .A1(n16128), .A2(n16129), .ZN(n16022) );
  INV_X1 U16156 ( .A(n16130), .ZN(n16129) );
  NAND2_X1 U16157 ( .A1(n15902), .A2(n16131), .ZN(n16130) );
  NAND2_X1 U16158 ( .A1(n15901), .A2(n15903), .ZN(n16131) );
  NOR2_X1 U16159 ( .A1(n8768), .A2(n15690), .ZN(n15902) );
  NOR2_X1 U16160 ( .A1(n15901), .A2(n15903), .ZN(n16128) );
  NOR2_X1 U16161 ( .A1(n16132), .A2(n16133), .ZN(n15903) );
  INV_X1 U16162 ( .A(n16134), .ZN(n16133) );
  NAND2_X1 U16163 ( .A1(n16019), .A2(n16135), .ZN(n16134) );
  NAND2_X1 U16164 ( .A1(n16018), .A2(n16017), .ZN(n16135) );
  NOR2_X1 U16165 ( .A1(n8772), .A2(n15690), .ZN(n16019) );
  NOR2_X1 U16166 ( .A1(n16017), .A2(n16018), .ZN(n16132) );
  NOR2_X1 U16167 ( .A1(n16136), .A2(n16137), .ZN(n16018) );
  INV_X1 U16168 ( .A(n16138), .ZN(n16137) );
  NAND2_X1 U16169 ( .A1(n15914), .A2(n16139), .ZN(n16138) );
  NAND2_X1 U16170 ( .A1(n15915), .A2(n15913), .ZN(n16139) );
  NOR2_X1 U16171 ( .A1(n10616), .A2(n15690), .ZN(n15914) );
  NOR2_X1 U16172 ( .A1(n15913), .A2(n15915), .ZN(n16136) );
  NOR2_X1 U16173 ( .A1(n16140), .A2(n16141), .ZN(n15915) );
  INV_X1 U16174 ( .A(n16142), .ZN(n16141) );
  NAND2_X1 U16175 ( .A1(n16015), .A2(n16143), .ZN(n16142) );
  NAND2_X1 U16176 ( .A1(n16014), .A2(n16013), .ZN(n16143) );
  NOR2_X1 U16177 ( .A1(n15690), .A2(n8881), .ZN(n16015) );
  NOR2_X1 U16178 ( .A1(n16013), .A2(n16014), .ZN(n16140) );
  NOR2_X1 U16179 ( .A1(n16144), .A2(n16145), .ZN(n16014) );
  INV_X1 U16180 ( .A(n16146), .ZN(n16145) );
  NAND2_X1 U16181 ( .A1(n15926), .A2(n16147), .ZN(n16146) );
  NAND2_X1 U16182 ( .A1(n15927), .A2(n15925), .ZN(n16147) );
  NOR2_X1 U16183 ( .A1(n15690), .A2(n10633), .ZN(n15926) );
  NOR2_X1 U16184 ( .A1(n15925), .A2(n15927), .ZN(n16144) );
  NOR2_X1 U16185 ( .A1(n16148), .A2(n16149), .ZN(n15927) );
  INV_X1 U16186 ( .A(n16150), .ZN(n16149) );
  NAND2_X1 U16187 ( .A1(n16011), .A2(n16151), .ZN(n16150) );
  NAND2_X1 U16188 ( .A1(n16010), .A2(n16009), .ZN(n16151) );
  NOR2_X1 U16189 ( .A1(n15690), .A2(n8798), .ZN(n16011) );
  NOR2_X1 U16190 ( .A1(n16009), .A2(n16010), .ZN(n16148) );
  NOR2_X1 U16191 ( .A1(n16152), .A2(n16153), .ZN(n16010) );
  INV_X1 U16192 ( .A(n16154), .ZN(n16153) );
  NAND2_X1 U16193 ( .A1(n15938), .A2(n16155), .ZN(n16154) );
  NAND2_X1 U16194 ( .A1(n15939), .A2(n15937), .ZN(n16155) );
  NOR2_X1 U16195 ( .A1(n15690), .A2(n8803), .ZN(n15938) );
  NOR2_X1 U16196 ( .A1(n15937), .A2(n15939), .ZN(n16152) );
  NOR2_X1 U16197 ( .A1(n16156), .A2(n16157), .ZN(n15939) );
  NOR2_X1 U16198 ( .A1(n16007), .A2(n16158), .ZN(n16157) );
  NOR2_X1 U16199 ( .A1(n16006), .A2(n16004), .ZN(n16158) );
  NAND2_X1 U16200 ( .A1(b_2_), .A2(a_23_), .ZN(n16007) );
  INV_X1 U16201 ( .A(n16159), .ZN(n16156) );
  NAND2_X1 U16202 ( .A1(n16004), .A2(n16006), .ZN(n16159) );
  NAND2_X1 U16203 ( .A1(n15949), .A2(n16160), .ZN(n16006) );
  NAND2_X1 U16204 ( .A1(n15948), .A2(n15950), .ZN(n16160) );
  NAND2_X1 U16205 ( .A1(n16161), .A2(n16162), .ZN(n15950) );
  NAND2_X1 U16206 ( .A1(b_2_), .A2(a_24_), .ZN(n16162) );
  INV_X1 U16207 ( .A(n16163), .ZN(n16161) );
  XOR2_X1 U16208 ( .A(n16164), .B(n16165), .Z(n15948) );
  NOR2_X1 U16209 ( .A1(n8825), .A2(n15994), .ZN(n16165) );
  XOR2_X1 U16210 ( .A(n16166), .B(n16167), .Z(n16164) );
  NAND2_X1 U16211 ( .A1(a_24_), .A2(n16163), .ZN(n15949) );
  NAND2_X1 U16212 ( .A1(n16002), .A2(n16168), .ZN(n16163) );
  NAND2_X1 U16213 ( .A1(n16001), .A2(n16003), .ZN(n16168) );
  NAND2_X1 U16214 ( .A1(n16169), .A2(n16170), .ZN(n16003) );
  NAND2_X1 U16215 ( .A1(b_2_), .A2(a_25_), .ZN(n16170) );
  INV_X1 U16216 ( .A(n16171), .ZN(n16169) );
  XOR2_X1 U16217 ( .A(n16172), .B(n16173), .Z(n16001) );
  NOR2_X1 U16218 ( .A1(n8830), .A2(n15994), .ZN(n16173) );
  XOR2_X1 U16219 ( .A(n16174), .B(n16175), .Z(n16172) );
  NAND2_X1 U16220 ( .A1(a_25_), .A2(n16171), .ZN(n16002) );
  NAND2_X1 U16221 ( .A1(n16176), .A2(n16177), .ZN(n16171) );
  NAND2_X1 U16222 ( .A1(n16178), .A2(b_2_), .ZN(n16177) );
  NOR2_X1 U16223 ( .A1(n16179), .A2(n8830), .ZN(n16178) );
  NOR2_X1 U16224 ( .A1(n15960), .A2(n15962), .ZN(n16179) );
  NAND2_X1 U16225 ( .A1(n15960), .A2(n15962), .ZN(n16176) );
  NAND2_X1 U16226 ( .A1(n15969), .A2(n16180), .ZN(n15962) );
  NAND2_X1 U16227 ( .A1(n15968), .A2(n15970), .ZN(n16180) );
  NAND2_X1 U16228 ( .A1(n16181), .A2(n16182), .ZN(n15970) );
  NAND2_X1 U16229 ( .A1(b_2_), .A2(a_27_), .ZN(n16182) );
  INV_X1 U16230 ( .A(n16183), .ZN(n16181) );
  XOR2_X1 U16231 ( .A(n16184), .B(n16185), .Z(n15968) );
  NOR2_X1 U16232 ( .A1(n16186), .A2(n16187), .ZN(n16185) );
  INV_X1 U16233 ( .A(n16188), .ZN(n16187) );
  NOR2_X1 U16234 ( .A1(n16189), .A2(n16190), .ZN(n16186) );
  NAND2_X1 U16235 ( .A1(a_27_), .A2(n16183), .ZN(n15969) );
  NAND2_X1 U16236 ( .A1(n16191), .A2(n16192), .ZN(n16183) );
  NAND2_X1 U16237 ( .A1(n16193), .A2(b_2_), .ZN(n16192) );
  NOR2_X1 U16238 ( .A1(n16194), .A2(n8844), .ZN(n16193) );
  NOR2_X1 U16239 ( .A1(n15979), .A2(n15977), .ZN(n16194) );
  NAND2_X1 U16240 ( .A1(n15977), .A2(n15979), .ZN(n16191) );
  NAND2_X1 U16241 ( .A1(n16195), .A2(n16196), .ZN(n15979) );
  NAND2_X1 U16242 ( .A1(n15996), .A2(n16197), .ZN(n16196) );
  INV_X1 U16243 ( .A(n16198), .ZN(n16197) );
  NOR2_X1 U16244 ( .A1(n15999), .A2(n15998), .ZN(n16198) );
  NOR2_X1 U16245 ( .A1(n15690), .A2(n9161), .ZN(n15996) );
  NAND2_X1 U16246 ( .A1(n15998), .A2(n15999), .ZN(n16195) );
  NAND2_X1 U16247 ( .A1(n16199), .A2(n16200), .ZN(n15999) );
  NAND2_X1 U16248 ( .A1(b_0_), .A2(n16201), .ZN(n16200) );
  NAND2_X1 U16249 ( .A1(n8358), .A2(n16202), .ZN(n16201) );
  NAND2_X1 U16250 ( .A1(a_31_), .A2(n15994), .ZN(n16202) );
  NAND2_X1 U16251 ( .A1(b_1_), .A2(n16204), .ZN(n16199) );
  NAND2_X1 U16252 ( .A1(n8362), .A2(n16205), .ZN(n16204) );
  NAND2_X1 U16253 ( .A1(a_30_), .A2(n16206), .ZN(n16205) );
  NOR2_X1 U16254 ( .A1(n16203), .A2(a_31_), .ZN(n16207) );
  NOR2_X1 U16255 ( .A1(n16208), .A2(n15994), .ZN(n15998) );
  NAND2_X1 U16256 ( .A1(n9926), .A2(b_2_), .ZN(n16208) );
  INV_X1 U16257 ( .A(n9170), .ZN(n9926) );
  XNOR2_X1 U16258 ( .A(n16209), .B(n16210), .ZN(n15977) );
  XNOR2_X1 U16259 ( .A(n16211), .B(n16212), .ZN(n16210) );
  NAND2_X1 U16260 ( .A1(b_0_), .A2(a_30_), .ZN(n16209) );
  XOR2_X1 U16261 ( .A(n16213), .B(n16214), .Z(n15960) );
  NOR2_X1 U16262 ( .A1(n8839), .A2(n15994), .ZN(n16214) );
  XOR2_X1 U16263 ( .A(n16215), .B(n16216), .Z(n16213) );
  XOR2_X1 U16264 ( .A(n16217), .B(n16218), .Z(n16004) );
  NOR2_X1 U16265 ( .A1(n9131), .A2(n15994), .ZN(n16218) );
  XOR2_X1 U16266 ( .A(n16219), .B(n16220), .Z(n16217) );
  XNOR2_X1 U16267 ( .A(n16221), .B(n16222), .ZN(n15937) );
  NOR2_X1 U16268 ( .A1(n8812), .A2(n15994), .ZN(n16222) );
  XOR2_X1 U16269 ( .A(n16223), .B(n16224), .Z(n16221) );
  XNOR2_X1 U16270 ( .A(n16225), .B(n16226), .ZN(n16009) );
  NOR2_X1 U16271 ( .A1(n8803), .A2(n15994), .ZN(n16226) );
  XOR2_X1 U16272 ( .A(n16227), .B(n16228), .Z(n16225) );
  XNOR2_X1 U16273 ( .A(n16229), .B(n16230), .ZN(n15925) );
  NOR2_X1 U16274 ( .A1(n8798), .A2(n15994), .ZN(n16230) );
  XOR2_X1 U16275 ( .A(n16231), .B(n16232), .Z(n16229) );
  XNOR2_X1 U16276 ( .A(n16233), .B(n16234), .ZN(n16013) );
  NOR2_X1 U16277 ( .A1(n10633), .A2(n15994), .ZN(n16234) );
  XOR2_X1 U16278 ( .A(n16235), .B(n16236), .Z(n16233) );
  XNOR2_X1 U16279 ( .A(n16237), .B(n16238), .ZN(n15913) );
  NOR2_X1 U16280 ( .A1(n8881), .A2(n15994), .ZN(n16238) );
  XOR2_X1 U16281 ( .A(n16239), .B(n16240), .Z(n16237) );
  XNOR2_X1 U16282 ( .A(n16241), .B(n16242), .ZN(n16017) );
  XNOR2_X1 U16283 ( .A(n16243), .B(n16244), .ZN(n16241) );
  XNOR2_X1 U16284 ( .A(n16245), .B(n16246), .ZN(n15901) );
  XOR2_X1 U16285 ( .A(n16247), .B(n16248), .Z(n16246) );
  XNOR2_X1 U16286 ( .A(n16249), .B(n16250), .ZN(n16021) );
  XOR2_X1 U16287 ( .A(n16251), .B(n16252), .Z(n16249) );
  XOR2_X1 U16288 ( .A(n16253), .B(n16254), .Z(n15888) );
  XOR2_X1 U16289 ( .A(n16255), .B(n16256), .Z(n16253) );
  XOR2_X1 U16290 ( .A(n16257), .B(n16258), .Z(n16025) );
  XOR2_X1 U16291 ( .A(n16259), .B(n16260), .Z(n16257) );
  XOR2_X1 U16292 ( .A(n16261), .B(n16262), .Z(n15876) );
  XOR2_X1 U16293 ( .A(n16263), .B(n16264), .Z(n16261) );
  XOR2_X1 U16294 ( .A(n16265), .B(n16266), .Z(n16029) );
  XOR2_X1 U16295 ( .A(n16267), .B(n16268), .Z(n16265) );
  XOR2_X1 U16296 ( .A(n16269), .B(n16270), .Z(n15864) );
  XOR2_X1 U16297 ( .A(n16271), .B(n16272), .Z(n16269) );
  XOR2_X1 U16298 ( .A(n16273), .B(n16274), .Z(n16033) );
  XOR2_X1 U16299 ( .A(n16275), .B(n16276), .Z(n16273) );
  XOR2_X1 U16300 ( .A(n16277), .B(n16278), .Z(n15852) );
  XOR2_X1 U16301 ( .A(n16279), .B(n16280), .Z(n16277) );
  XOR2_X1 U16302 ( .A(n16281), .B(n16282), .Z(n16037) );
  XOR2_X1 U16303 ( .A(n16283), .B(n16284), .Z(n16281) );
  XOR2_X1 U16304 ( .A(n16285), .B(n16286), .Z(n15840) );
  XOR2_X1 U16305 ( .A(n16287), .B(n16288), .Z(n16285) );
  XOR2_X1 U16306 ( .A(n16289), .B(n16290), .Z(n16041) );
  XOR2_X1 U16307 ( .A(n16291), .B(n16292), .Z(n16289) );
  XNOR2_X1 U16308 ( .A(n16293), .B(n16294), .ZN(n15828) );
  XOR2_X1 U16309 ( .A(n16295), .B(n16296), .Z(n16293) );
  XNOR2_X1 U16310 ( .A(n16297), .B(n16298), .ZN(n15821) );
  XOR2_X1 U16311 ( .A(n16299), .B(n16300), .Z(n16297) );
  XOR2_X1 U16312 ( .A(n16301), .B(n16302), .Z(n16045) );
  XOR2_X1 U16313 ( .A(n16303), .B(n16304), .Z(n16301) );
  XOR2_X1 U16314 ( .A(n16305), .B(n16306), .Z(n16049) );
  XOR2_X1 U16315 ( .A(n16307), .B(n16308), .Z(n16305) );
  XOR2_X1 U16316 ( .A(n16309), .B(n16310), .Z(n16053) );
  XOR2_X1 U16317 ( .A(n16311), .B(n16312), .Z(n16309) );
  NAND2_X1 U16318 ( .A1(n16313), .A2(n16057), .ZN(n16058) );
  INV_X1 U16319 ( .A(n8608), .ZN(n16313) );
  NAND2_X1 U16320 ( .A1(n16314), .A2(n16315), .ZN(n8608) );
  NAND2_X1 U16321 ( .A1(n16310), .A2(n16316), .ZN(n16315) );
  INV_X1 U16322 ( .A(n16317), .ZN(n16316) );
  NOR2_X1 U16323 ( .A1(n16311), .A2(n16312), .ZN(n16317) );
  NOR2_X1 U16324 ( .A1(n8502), .A2(n16206), .ZN(n16310) );
  NAND2_X1 U16325 ( .A1(n16312), .A2(n16311), .ZN(n16314) );
  NAND2_X1 U16326 ( .A1(n16318), .A2(n16319), .ZN(n16311) );
  NAND2_X1 U16327 ( .A1(n16306), .A2(n16320), .ZN(n16319) );
  INV_X1 U16328 ( .A(n16321), .ZN(n16320) );
  NOR2_X1 U16329 ( .A1(n16308), .A2(n16307), .ZN(n16321) );
  NOR2_X1 U16330 ( .A1(n8497), .A2(n16206), .ZN(n16306) );
  NAND2_X1 U16331 ( .A1(n16307), .A2(n16308), .ZN(n16318) );
  NAND2_X1 U16332 ( .A1(n16322), .A2(n16323), .ZN(n16308) );
  NAND2_X1 U16333 ( .A1(n16302), .A2(n16324), .ZN(n16323) );
  INV_X1 U16334 ( .A(n16325), .ZN(n16324) );
  NOR2_X1 U16335 ( .A1(n16303), .A2(n16304), .ZN(n16325) );
  NOR2_X1 U16336 ( .A1(n8497), .A2(n15994), .ZN(n16302) );
  NAND2_X1 U16337 ( .A1(n16304), .A2(n16303), .ZN(n16322) );
  NAND2_X1 U16338 ( .A1(n16326), .A2(n16327), .ZN(n16303) );
  NAND2_X1 U16339 ( .A1(n16072), .A2(n16328), .ZN(n16327) );
  INV_X1 U16340 ( .A(n16329), .ZN(n16328) );
  NOR2_X1 U16341 ( .A1(n16074), .A2(n16073), .ZN(n16329) );
  NOR2_X1 U16342 ( .A1(n8707), .A2(n15994), .ZN(n16072) );
  NAND2_X1 U16343 ( .A1(n16073), .A2(n16074), .ZN(n16326) );
  NAND2_X1 U16344 ( .A1(n16330), .A2(n16331), .ZN(n16074) );
  NAND2_X1 U16345 ( .A1(n16298), .A2(n16332), .ZN(n16331) );
  INV_X1 U16346 ( .A(n16333), .ZN(n16332) );
  NOR2_X1 U16347 ( .A1(n16299), .A2(n16300), .ZN(n16333) );
  NOR2_X1 U16348 ( .A1(n8712), .A2(n15994), .ZN(n16298) );
  NAND2_X1 U16349 ( .A1(n16300), .A2(n16299), .ZN(n16330) );
  NAND2_X1 U16350 ( .A1(n16334), .A2(n16335), .ZN(n16299) );
  NAND2_X1 U16351 ( .A1(n16294), .A2(n16336), .ZN(n16335) );
  INV_X1 U16352 ( .A(n16337), .ZN(n16336) );
  NOR2_X1 U16353 ( .A1(n16296), .A2(n16295), .ZN(n16337) );
  NOR2_X1 U16354 ( .A1(n8717), .A2(n15994), .ZN(n16294) );
  NAND2_X1 U16355 ( .A1(n16295), .A2(n16296), .ZN(n16334) );
  NAND2_X1 U16356 ( .A1(n16338), .A2(n16339), .ZN(n16296) );
  NAND2_X1 U16357 ( .A1(n16290), .A2(n16340), .ZN(n16339) );
  INV_X1 U16358 ( .A(n16341), .ZN(n16340) );
  NOR2_X1 U16359 ( .A1(n16291), .A2(n16292), .ZN(n16341) );
  NOR2_X1 U16360 ( .A1(n8480), .A2(n15994), .ZN(n16290) );
  NAND2_X1 U16361 ( .A1(n16292), .A2(n16291), .ZN(n16338) );
  NAND2_X1 U16362 ( .A1(n16342), .A2(n16343), .ZN(n16291) );
  NAND2_X1 U16363 ( .A1(n16286), .A2(n16344), .ZN(n16343) );
  INV_X1 U16364 ( .A(n16345), .ZN(n16344) );
  NOR2_X1 U16365 ( .A1(n16288), .A2(n16287), .ZN(n16345) );
  NOR2_X1 U16366 ( .A1(n8726), .A2(n15994), .ZN(n16286) );
  NAND2_X1 U16367 ( .A1(n16287), .A2(n16288), .ZN(n16342) );
  NAND2_X1 U16368 ( .A1(n16346), .A2(n16347), .ZN(n16288) );
  NAND2_X1 U16369 ( .A1(n16282), .A2(n16348), .ZN(n16347) );
  INV_X1 U16370 ( .A(n16349), .ZN(n16348) );
  NOR2_X1 U16371 ( .A1(n16283), .A2(n16284), .ZN(n16349) );
  NOR2_X1 U16372 ( .A1(n8731), .A2(n15994), .ZN(n16282) );
  NAND2_X1 U16373 ( .A1(n16284), .A2(n16283), .ZN(n16346) );
  NAND2_X1 U16374 ( .A1(n16350), .A2(n16351), .ZN(n16283) );
  NAND2_X1 U16375 ( .A1(n16278), .A2(n16352), .ZN(n16351) );
  INV_X1 U16376 ( .A(n16353), .ZN(n16352) );
  NOR2_X1 U16377 ( .A1(n16280), .A2(n16279), .ZN(n16353) );
  NOR2_X1 U16378 ( .A1(n8736), .A2(n15994), .ZN(n16278) );
  NAND2_X1 U16379 ( .A1(n16279), .A2(n16280), .ZN(n16350) );
  NAND2_X1 U16380 ( .A1(n16354), .A2(n16355), .ZN(n16280) );
  NAND2_X1 U16381 ( .A1(n16274), .A2(n16356), .ZN(n16355) );
  INV_X1 U16382 ( .A(n16357), .ZN(n16356) );
  NOR2_X1 U16383 ( .A1(n16275), .A2(n16276), .ZN(n16357) );
  NOR2_X1 U16384 ( .A1(n8741), .A2(n15994), .ZN(n16274) );
  NAND2_X1 U16385 ( .A1(n16276), .A2(n16275), .ZN(n16354) );
  NAND2_X1 U16386 ( .A1(n16358), .A2(n16359), .ZN(n16275) );
  NAND2_X1 U16387 ( .A1(n16270), .A2(n16360), .ZN(n16359) );
  INV_X1 U16388 ( .A(n16361), .ZN(n16360) );
  NOR2_X1 U16389 ( .A1(n16272), .A2(n16271), .ZN(n16361) );
  NOR2_X1 U16390 ( .A1(n8452), .A2(n15994), .ZN(n16270) );
  NAND2_X1 U16391 ( .A1(n16271), .A2(n16272), .ZN(n16358) );
  NAND2_X1 U16392 ( .A1(n16362), .A2(n16363), .ZN(n16272) );
  NAND2_X1 U16393 ( .A1(n16266), .A2(n16364), .ZN(n16363) );
  INV_X1 U16394 ( .A(n16365), .ZN(n16364) );
  NOR2_X1 U16395 ( .A1(n16267), .A2(n16268), .ZN(n16365) );
  NOR2_X1 U16396 ( .A1(n8750), .A2(n15994), .ZN(n16266) );
  NAND2_X1 U16397 ( .A1(n16268), .A2(n16267), .ZN(n16362) );
  NAND2_X1 U16398 ( .A1(n16366), .A2(n16367), .ZN(n16267) );
  NAND2_X1 U16399 ( .A1(n16262), .A2(n16368), .ZN(n16367) );
  INV_X1 U16400 ( .A(n16369), .ZN(n16368) );
  NOR2_X1 U16401 ( .A1(n16264), .A2(n16263), .ZN(n16369) );
  NOR2_X1 U16402 ( .A1(n8443), .A2(n15994), .ZN(n16262) );
  NAND2_X1 U16403 ( .A1(n16263), .A2(n16264), .ZN(n16366) );
  NAND2_X1 U16404 ( .A1(n16370), .A2(n16371), .ZN(n16264) );
  NAND2_X1 U16405 ( .A1(n16258), .A2(n16372), .ZN(n16371) );
  INV_X1 U16406 ( .A(n16373), .ZN(n16372) );
  NOR2_X1 U16407 ( .A1(n16259), .A2(n16260), .ZN(n16373) );
  NOR2_X1 U16408 ( .A1(n8438), .A2(n15994), .ZN(n16258) );
  NAND2_X1 U16409 ( .A1(n16260), .A2(n16259), .ZN(n16370) );
  NAND2_X1 U16410 ( .A1(n16374), .A2(n16375), .ZN(n16259) );
  NAND2_X1 U16411 ( .A1(n16254), .A2(n16376), .ZN(n16375) );
  INV_X1 U16412 ( .A(n16377), .ZN(n16376) );
  NOR2_X1 U16413 ( .A1(n16256), .A2(n16255), .ZN(n16377) );
  NOR2_X1 U16414 ( .A1(n8763), .A2(n15994), .ZN(n16254) );
  NAND2_X1 U16415 ( .A1(n16255), .A2(n16256), .ZN(n16374) );
  NAND2_X1 U16416 ( .A1(n16378), .A2(n16379), .ZN(n16256) );
  NAND2_X1 U16417 ( .A1(n16250), .A2(n16380), .ZN(n16379) );
  INV_X1 U16418 ( .A(n16381), .ZN(n16380) );
  NOR2_X1 U16419 ( .A1(n16251), .A2(n16252), .ZN(n16381) );
  NOR2_X1 U16420 ( .A1(n8768), .A2(n15994), .ZN(n16250) );
  NAND2_X1 U16421 ( .A1(n16252), .A2(n16251), .ZN(n16378) );
  NAND2_X1 U16422 ( .A1(n16382), .A2(n16383), .ZN(n16251) );
  NAND2_X1 U16423 ( .A1(n16245), .A2(n16384), .ZN(n16383) );
  NAND2_X1 U16424 ( .A1(n16248), .A2(n16247), .ZN(n16384) );
  NOR2_X1 U16425 ( .A1(n8772), .A2(n15994), .ZN(n16245) );
  INV_X1 U16426 ( .A(n16385), .ZN(n16382) );
  NOR2_X1 U16427 ( .A1(n16248), .A2(n16247), .ZN(n16385) );
  NAND2_X1 U16428 ( .A1(a_18_), .A2(b_0_), .ZN(n16247) );
  NAND2_X1 U16429 ( .A1(n16386), .A2(n16387), .ZN(n16248) );
  NAND2_X1 U16430 ( .A1(n16388), .A2(n16244), .ZN(n16387) );
  NAND2_X1 U16431 ( .A1(b_0_), .A2(a_19_), .ZN(n16244) );
  NAND2_X1 U16432 ( .A1(n16242), .A2(n16243), .ZN(n16388) );
  INV_X1 U16433 ( .A(n16389), .ZN(n16386) );
  NOR2_X1 U16434 ( .A1(n16243), .A2(n16242), .ZN(n16389) );
  NOR2_X1 U16435 ( .A1(n10616), .A2(n15994), .ZN(n16242) );
  NAND2_X1 U16436 ( .A1(n16390), .A2(n16391), .ZN(n16243) );
  NAND2_X1 U16437 ( .A1(n16392), .A2(b_1_), .ZN(n16391) );
  NOR2_X1 U16438 ( .A1(n16393), .A2(n8881), .ZN(n16392) );
  NOR2_X1 U16439 ( .A1(n16240), .A2(n16239), .ZN(n16393) );
  NAND2_X1 U16440 ( .A1(n16240), .A2(n16239), .ZN(n16390) );
  NAND2_X1 U16441 ( .A1(n16394), .A2(n16395), .ZN(n16239) );
  NAND2_X1 U16442 ( .A1(n16396), .A2(b_1_), .ZN(n16395) );
  NOR2_X1 U16443 ( .A1(n16397), .A2(n10633), .ZN(n16396) );
  NOR2_X1 U16444 ( .A1(n16236), .A2(n16235), .ZN(n16397) );
  NAND2_X1 U16445 ( .A1(n16236), .A2(n16235), .ZN(n16394) );
  NAND2_X1 U16446 ( .A1(n16398), .A2(n16399), .ZN(n16235) );
  NAND2_X1 U16447 ( .A1(n16400), .A2(b_1_), .ZN(n16399) );
  NOR2_X1 U16448 ( .A1(n16401), .A2(n8798), .ZN(n16400) );
  NOR2_X1 U16449 ( .A1(n16232), .A2(n16231), .ZN(n16401) );
  NAND2_X1 U16450 ( .A1(n16232), .A2(n16231), .ZN(n16398) );
  NAND2_X1 U16451 ( .A1(n16402), .A2(n16403), .ZN(n16231) );
  NAND2_X1 U16452 ( .A1(n16404), .A2(b_1_), .ZN(n16403) );
  NOR2_X1 U16453 ( .A1(n16405), .A2(n8803), .ZN(n16404) );
  NOR2_X1 U16454 ( .A1(n16228), .A2(n16227), .ZN(n16405) );
  NAND2_X1 U16455 ( .A1(n16228), .A2(n16227), .ZN(n16402) );
  NAND2_X1 U16456 ( .A1(n16406), .A2(n16407), .ZN(n16227) );
  NAND2_X1 U16457 ( .A1(n16408), .A2(b_1_), .ZN(n16407) );
  NOR2_X1 U16458 ( .A1(n16409), .A2(n8812), .ZN(n16408) );
  NOR2_X1 U16459 ( .A1(n16224), .A2(n16223), .ZN(n16409) );
  NAND2_X1 U16460 ( .A1(n16224), .A2(n16223), .ZN(n16406) );
  NAND2_X1 U16461 ( .A1(n16410), .A2(n16411), .ZN(n16223) );
  NAND2_X1 U16462 ( .A1(n16412), .A2(b_1_), .ZN(n16411) );
  NOR2_X1 U16463 ( .A1(n16413), .A2(n9131), .ZN(n16412) );
  NOR2_X1 U16464 ( .A1(n16220), .A2(n16219), .ZN(n16413) );
  NAND2_X1 U16465 ( .A1(n16220), .A2(n16219), .ZN(n16410) );
  NAND2_X1 U16466 ( .A1(n16414), .A2(n16415), .ZN(n16219) );
  NAND2_X1 U16467 ( .A1(n16416), .A2(b_1_), .ZN(n16415) );
  NOR2_X1 U16468 ( .A1(n16417), .A2(n8825), .ZN(n16416) );
  NOR2_X1 U16469 ( .A1(n16167), .A2(n16166), .ZN(n16417) );
  NAND2_X1 U16470 ( .A1(n16167), .A2(n16166), .ZN(n16414) );
  NAND2_X1 U16471 ( .A1(n16418), .A2(n16419), .ZN(n16166) );
  NAND2_X1 U16472 ( .A1(n16420), .A2(b_1_), .ZN(n16419) );
  NOR2_X1 U16473 ( .A1(n16421), .A2(n8830), .ZN(n16420) );
  NOR2_X1 U16474 ( .A1(n16175), .A2(n16174), .ZN(n16421) );
  NAND2_X1 U16475 ( .A1(n16175), .A2(n16174), .ZN(n16418) );
  NAND2_X1 U16476 ( .A1(n16422), .A2(n16423), .ZN(n16174) );
  NAND2_X1 U16477 ( .A1(n16424), .A2(b_1_), .ZN(n16423) );
  NOR2_X1 U16478 ( .A1(n16425), .A2(n8839), .ZN(n16424) );
  NOR2_X1 U16479 ( .A1(n16216), .A2(n16215), .ZN(n16425) );
  NAND2_X1 U16480 ( .A1(n16216), .A2(n16215), .ZN(n16422) );
  NAND2_X1 U16481 ( .A1(n16188), .A2(n16426), .ZN(n16215) );
  NAND2_X1 U16482 ( .A1(n16427), .A2(n16184), .ZN(n16426) );
  NAND2_X1 U16483 ( .A1(n16212), .A2(n16428), .ZN(n16184) );
  NAND2_X1 U16484 ( .A1(n16429), .A2(n16211), .ZN(n16428) );
  NOR2_X1 U16485 ( .A1(n15994), .A2(n9161), .ZN(n16211) );
  NOR2_X1 U16486 ( .A1(n16203), .A2(n16206), .ZN(n16429) );
  NAND2_X1 U16487 ( .A1(n16430), .A2(b_0_), .ZN(n16212) );
  NOR2_X1 U16488 ( .A1(n9170), .A2(n15994), .ZN(n16430) );
  NAND2_X1 U16489 ( .A1(a_31_), .A2(a_30_), .ZN(n9170) );
  INV_X1 U16490 ( .A(n16431), .ZN(n16427) );
  NOR2_X1 U16491 ( .A1(n16189), .A2(a_28_), .ZN(n16431) );
  NAND2_X1 U16492 ( .A1(n16190), .A2(n16189), .ZN(n16188) );
  NOR2_X1 U16493 ( .A1(n16206), .A2(n9161), .ZN(n16189) );
  NOR2_X1 U16494 ( .A1(n8844), .A2(n15994), .ZN(n16190) );
  NOR2_X1 U16495 ( .A1(n16206), .A2(n8844), .ZN(n16216) );
  NOR2_X1 U16496 ( .A1(n16206), .A2(n8839), .ZN(n16175) );
  NOR2_X1 U16497 ( .A1(n16206), .A2(n8830), .ZN(n16167) );
  NOR2_X1 U16498 ( .A1(n16206), .A2(n8825), .ZN(n16220) );
  NOR2_X1 U16499 ( .A1(n16206), .A2(n9131), .ZN(n16224) );
  NOR2_X1 U16500 ( .A1(n16206), .A2(n8812), .ZN(n16228) );
  NOR2_X1 U16501 ( .A1(n16206), .A2(n8803), .ZN(n16232) );
  NOR2_X1 U16502 ( .A1(n16206), .A2(n8798), .ZN(n16236) );
  NOR2_X1 U16503 ( .A1(n16206), .A2(n10633), .ZN(n16240) );
  NOR2_X1 U16504 ( .A1(n8772), .A2(n16206), .ZN(n16252) );
  NOR2_X1 U16505 ( .A1(n8768), .A2(n16206), .ZN(n16255) );
  NOR2_X1 U16506 ( .A1(n8763), .A2(n16206), .ZN(n16260) );
  NOR2_X1 U16507 ( .A1(n8438), .A2(n16206), .ZN(n16263) );
  NOR2_X1 U16508 ( .A1(n8443), .A2(n16206), .ZN(n16268) );
  NOR2_X1 U16509 ( .A1(n8750), .A2(n16206), .ZN(n16271) );
  NOR2_X1 U16510 ( .A1(n8452), .A2(n16206), .ZN(n16276) );
  NOR2_X1 U16511 ( .A1(n8741), .A2(n16206), .ZN(n16279) );
  NOR2_X1 U16512 ( .A1(n8736), .A2(n16206), .ZN(n16284) );
  NOR2_X1 U16513 ( .A1(n8731), .A2(n16206), .ZN(n16287) );
  NOR2_X1 U16514 ( .A1(n8726), .A2(n16206), .ZN(n16292) );
  NOR2_X1 U16515 ( .A1(n8480), .A2(n16206), .ZN(n16295) );
  NOR2_X1 U16516 ( .A1(n8717), .A2(n16206), .ZN(n16300) );
  NOR2_X1 U16517 ( .A1(n8712), .A2(n16206), .ZN(n16073) );
  NOR2_X1 U16518 ( .A1(n8707), .A2(n16206), .ZN(n16304) );
  NOR2_X1 U16519 ( .A1(n8690), .A2(n15994), .ZN(n16312) );
  NAND2_X1 U16520 ( .A1(n16432), .A2(n16433), .ZN(Result_add_9_) );
  NAND2_X1 U16521 ( .A1(n14071), .A2(n16434), .ZN(n16433) );
  INV_X1 U16522 ( .A(n14329), .ZN(n14071) );
  NOR2_X1 U16523 ( .A1(n16435), .A2(n16436), .ZN(n16432) );
  NOR2_X1 U16524 ( .A1(b_9_), .A2(n16437), .ZN(n16436) );
  XOR2_X1 U16525 ( .A(n8736), .B(n16434), .Z(n16437) );
  INV_X1 U16526 ( .A(n16438), .ZN(n16435) );
  NAND2_X1 U16527 ( .A1(b_9_), .A2(n16439), .ZN(n16438) );
  NOR2_X1 U16528 ( .A1(n16434), .A2(a_9_), .ZN(n16439) );
  XNOR2_X1 U16529 ( .A(n16440), .B(n16441), .ZN(Result_add_8_) );
  NAND2_X1 U16530 ( .A1(n16442), .A2(n14503), .ZN(n16441) );
  NAND2_X1 U16531 ( .A1(n16443), .A2(n16444), .ZN(Result_add_7_) );
  NAND2_X1 U16532 ( .A1(n14830), .A2(n16445), .ZN(n16444) );
  INV_X1 U16533 ( .A(n14757), .ZN(n14830) );
  NOR2_X1 U16534 ( .A1(n16446), .A2(n16447), .ZN(n16443) );
  NOR2_X1 U16535 ( .A1(b_7_), .A2(n16448), .ZN(n16447) );
  XOR2_X1 U16536 ( .A(n8726), .B(n16445), .Z(n16448) );
  INV_X1 U16537 ( .A(n16449), .ZN(n16446) );
  NAND2_X1 U16538 ( .A1(b_7_), .A2(n16450), .ZN(n16449) );
  NOR2_X1 U16539 ( .A1(n16445), .A2(a_7_), .ZN(n16450) );
  XNOR2_X1 U16540 ( .A(n16451), .B(n16452), .ZN(Result_add_6_) );
  NAND2_X1 U16541 ( .A1(n16453), .A2(n15020), .ZN(n16452) );
  NAND2_X1 U16542 ( .A1(n16454), .A2(n16455), .ZN(Result_add_5_) );
  NAND2_X1 U16543 ( .A1(n15274), .A2(n16456), .ZN(n16455) );
  INV_X1 U16544 ( .A(n16457), .ZN(n15274) );
  NOR2_X1 U16545 ( .A1(n16458), .A2(n16459), .ZN(n16454) );
  NOR2_X1 U16546 ( .A1(b_5_), .A2(n16460), .ZN(n16459) );
  XOR2_X1 U16547 ( .A(n8717), .B(n16456), .Z(n16460) );
  INV_X1 U16548 ( .A(n16461), .ZN(n16458) );
  NAND2_X1 U16549 ( .A1(b_5_), .A2(n16462), .ZN(n16461) );
  NOR2_X1 U16550 ( .A1(n16456), .A2(a_5_), .ZN(n16462) );
  XNOR2_X1 U16551 ( .A(n16463), .B(n16464), .ZN(Result_add_4_) );
  NAND2_X1 U16552 ( .A1(n16465), .A2(n15535), .ZN(n16464) );
  NAND2_X1 U16553 ( .A1(n16466), .A2(n16467), .ZN(Result_add_3_) );
  NAND2_X1 U16554 ( .A1(n15787), .A2(n16468), .ZN(n16467) );
  INV_X1 U16555 ( .A(n16469), .ZN(n15787) );
  NOR2_X1 U16556 ( .A1(n16470), .A2(n16471), .ZN(n16466) );
  NOR2_X1 U16557 ( .A1(b_3_), .A2(n16472), .ZN(n16471) );
  XOR2_X1 U16558 ( .A(n8707), .B(n16468), .Z(n16472) );
  INV_X1 U16559 ( .A(n16473), .ZN(n16470) );
  NAND2_X1 U16560 ( .A1(b_3_), .A2(n16474), .ZN(n16473) );
  NOR2_X1 U16561 ( .A1(n16468), .A2(a_3_), .ZN(n16474) );
  XOR2_X1 U16562 ( .A(b_31_), .B(a_31_), .Z(Result_add_31_) );
  NAND2_X1 U16563 ( .A1(n16475), .A2(n8852), .ZN(Result_add_30_) );
  NAND2_X1 U16564 ( .A1(n16476), .A2(Result_mul_63_), .ZN(n8852) );
  NOR2_X1 U16565 ( .A1(n16203), .A2(n8364), .ZN(n16476) );
  NOR2_X1 U16566 ( .A1(n16477), .A2(n16478), .ZN(n16475) );
  NOR2_X1 U16567 ( .A1(n8364), .A2(n16479), .ZN(n16478) );
  INV_X1 U16568 ( .A(b_30_), .ZN(n8364) );
  NOR2_X1 U16569 ( .A1(b_30_), .A2(n16480), .ZN(n16477) );
  XOR2_X1 U16570 ( .A(n16481), .B(a_30_), .Z(n16480) );
  XNOR2_X1 U16571 ( .A(n16482), .B(n16483), .ZN(Result_add_2_) );
  NAND2_X1 U16572 ( .A1(n16484), .A2(n15815), .ZN(n16483) );
  NAND2_X1 U16573 ( .A1(n16485), .A2(n16486), .ZN(Result_add_29_) );
  NAND2_X1 U16574 ( .A1(n9171), .A2(n16487), .ZN(n16486) );
  NOR2_X1 U16575 ( .A1(n16488), .A2(n16489), .ZN(n16485) );
  NOR2_X1 U16576 ( .A1(b_29_), .A2(n16490), .ZN(n16489) );
  XOR2_X1 U16577 ( .A(n9161), .B(n16487), .Z(n16490) );
  NOR2_X1 U16578 ( .A1(n8860), .A2(n16491), .ZN(n16488) );
  NAND2_X1 U16579 ( .A1(n16492), .A2(n9161), .ZN(n16491) );
  XNOR2_X1 U16580 ( .A(n16493), .B(n16494), .ZN(Result_add_28_) );
  NOR2_X1 U16581 ( .A1(n16495), .A2(n9400), .ZN(n16494) );
  NAND2_X1 U16582 ( .A1(n16496), .A2(n16497), .ZN(Result_add_27_) );
  NAND2_X1 U16583 ( .A1(n9905), .A2(n16498), .ZN(n16497) );
  INV_X1 U16584 ( .A(n9655), .ZN(n9905) );
  NOR2_X1 U16585 ( .A1(n16499), .A2(n16500), .ZN(n16496) );
  NOR2_X1 U16586 ( .A1(b_27_), .A2(n16501), .ZN(n16500) );
  XOR2_X1 U16587 ( .A(n8839), .B(n16498), .Z(n16501) );
  NOR2_X1 U16588 ( .A1(n9421), .A2(n16502), .ZN(n16499) );
  NAND2_X1 U16589 ( .A1(n16503), .A2(n8839), .ZN(n16502) );
  XNOR2_X1 U16590 ( .A(n16504), .B(n16505), .ZN(Result_add_26_) );
  NAND2_X1 U16591 ( .A1(n16506), .A2(n9892), .ZN(n16505) );
  NAND2_X1 U16592 ( .A1(n16507), .A2(n16508), .ZN(Result_add_25_) );
  NAND2_X1 U16593 ( .A1(n10393), .A2(n16509), .ZN(n16508) );
  INV_X1 U16594 ( .A(n10179), .ZN(n10393) );
  NOR2_X1 U16595 ( .A1(n16510), .A2(n16511), .ZN(n16507) );
  NOR2_X1 U16596 ( .A1(b_25_), .A2(n16512), .ZN(n16511) );
  XOR2_X1 U16597 ( .A(n8825), .B(n16509), .Z(n16512) );
  INV_X1 U16598 ( .A(n16513), .ZN(n16510) );
  NAND2_X1 U16599 ( .A1(b_25_), .A2(n16514), .ZN(n16513) );
  NOR2_X1 U16600 ( .A1(n16509), .A2(a_25_), .ZN(n16514) );
  XNOR2_X1 U16601 ( .A(n16515), .B(n16516), .ZN(Result_add_24_) );
  NAND2_X1 U16602 ( .A1(n16517), .A2(n10438), .ZN(n16516) );
  NAND2_X1 U16603 ( .A1(n16518), .A2(n16519), .ZN(Result_add_23_) );
  NAND2_X1 U16604 ( .A1(n10886), .A2(n16520), .ZN(n16519) );
  INV_X1 U16605 ( .A(n10649), .ZN(n10886) );
  NOR2_X1 U16606 ( .A1(n16521), .A2(n16522), .ZN(n16518) );
  NOR2_X1 U16607 ( .A1(b_23_), .A2(n16523), .ZN(n16522) );
  XOR2_X1 U16608 ( .A(n8812), .B(n16520), .Z(n16523) );
  INV_X1 U16609 ( .A(n16524), .ZN(n16521) );
  NAND2_X1 U16610 ( .A1(b_23_), .A2(n16525), .ZN(n16524) );
  NOR2_X1 U16611 ( .A1(n16520), .A2(a_23_), .ZN(n16525) );
  XNOR2_X1 U16612 ( .A(n16526), .B(n16527), .ZN(Result_add_22_) );
  NAND2_X1 U16613 ( .A1(n16528), .A2(n10874), .ZN(n16527) );
  NAND2_X1 U16614 ( .A1(n16529), .A2(n16530), .ZN(Result_add_21_) );
  NAND2_X1 U16615 ( .A1(n11136), .A2(n16531), .ZN(n16530) );
  INV_X1 U16616 ( .A(n16532), .ZN(n11136) );
  NOR2_X1 U16617 ( .A1(n16533), .A2(n16534), .ZN(n16529) );
  NOR2_X1 U16618 ( .A1(b_21_), .A2(n16535), .ZN(n16534) );
  XOR2_X1 U16619 ( .A(n8798), .B(n16531), .Z(n16535) );
  INV_X1 U16620 ( .A(n16536), .ZN(n16533) );
  NAND2_X1 U16621 ( .A1(b_21_), .A2(n16537), .ZN(n16536) );
  NOR2_X1 U16622 ( .A1(n16531), .A2(a_21_), .ZN(n16537) );
  XNOR2_X1 U16623 ( .A(n16538), .B(n16539), .ZN(Result_add_20_) );
  NAND2_X1 U16624 ( .A1(n16540), .A2(n11383), .ZN(n16539) );
  NAND2_X1 U16625 ( .A1(n16541), .A2(n16542), .ZN(Result_add_1_) );
  NAND2_X1 U16626 ( .A1(n16543), .A2(n16544), .ZN(n16542) );
  INV_X1 U16627 ( .A(n16545), .ZN(n16543) );
  NOR2_X1 U16628 ( .A1(n16307), .A2(n16546), .ZN(n16545) );
  NAND2_X1 U16629 ( .A1(n16547), .A2(n16548), .ZN(n16541) );
  INV_X1 U16630 ( .A(n16544), .ZN(n16548) );
  XOR2_X1 U16631 ( .A(b_1_), .B(a_1_), .Z(n16547) );
  NAND2_X1 U16632 ( .A1(n16549), .A2(n16550), .ZN(Result_add_19_) );
  NAND2_X1 U16633 ( .A1(n11740), .A2(n16551), .ZN(n16550) );
  NOR2_X1 U16634 ( .A1(n16552), .A2(n16553), .ZN(n16549) );
  NOR2_X1 U16635 ( .A1(b_19_), .A2(n16554), .ZN(n16553) );
  XOR2_X1 U16636 ( .A(n8881), .B(n16551), .Z(n16554) );
  NOR2_X1 U16637 ( .A1(n11452), .A2(n16555), .ZN(n16552) );
  NAND2_X1 U16638 ( .A1(n16556), .A2(n8881), .ZN(n16555) );
  XNOR2_X1 U16639 ( .A(n16557), .B(n16558), .ZN(Result_add_18_) );
  NOR2_X1 U16640 ( .A1(n16559), .A2(n11871), .ZN(n16558) );
  NAND2_X1 U16641 ( .A1(n16560), .A2(n16561), .ZN(Result_add_17_) );
  NAND2_X1 U16642 ( .A1(n12114), .A2(n16562), .ZN(n16561) );
  NOR2_X1 U16643 ( .A1(n16563), .A2(n16564), .ZN(n16560) );
  NOR2_X1 U16644 ( .A1(b_17_), .A2(n16565), .ZN(n16564) );
  XOR2_X1 U16645 ( .A(n8772), .B(n16562), .Z(n16565) );
  INV_X1 U16646 ( .A(n16566), .ZN(n16562) );
  NOR2_X1 U16647 ( .A1(n11951), .A2(n16567), .ZN(n16563) );
  NAND2_X1 U16648 ( .A1(n16566), .A2(n8772), .ZN(n16567) );
  XNOR2_X1 U16649 ( .A(n16568), .B(n16569), .ZN(Result_add_16_) );
  NOR2_X1 U16650 ( .A1(n16570), .A2(n12361), .ZN(n16569) );
  NAND2_X1 U16651 ( .A1(n16571), .A2(n16572), .ZN(Result_add_15_) );
  NAND2_X1 U16652 ( .A1(n12854), .A2(n16573), .ZN(n16572) );
  INV_X1 U16653 ( .A(n12752), .ZN(n12854) );
  NOR2_X1 U16654 ( .A1(n16574), .A2(n16575), .ZN(n16571) );
  NOR2_X1 U16655 ( .A1(b_15_), .A2(n16576), .ZN(n16575) );
  XOR2_X1 U16656 ( .A(n8763), .B(n16573), .Z(n16576) );
  NOR2_X1 U16657 ( .A1(n12453), .A2(n16577), .ZN(n16574) );
  NAND2_X1 U16658 ( .A1(n16578), .A2(n8763), .ZN(n16577) );
  XNOR2_X1 U16659 ( .A(n16579), .B(n16580), .ZN(Result_add_14_) );
  NAND2_X1 U16660 ( .A1(n16581), .A2(n12840), .ZN(n16580) );
  NAND2_X1 U16661 ( .A1(n16582), .A2(n16583), .ZN(Result_add_13_) );
  NAND2_X1 U16662 ( .A1(n13336), .A2(n16584), .ZN(n16583) );
  INV_X1 U16663 ( .A(n13124), .ZN(n13336) );
  NOR2_X1 U16664 ( .A1(n16585), .A2(n16586), .ZN(n16582) );
  NOR2_X1 U16665 ( .A1(b_13_), .A2(n16587), .ZN(n16586) );
  XOR2_X1 U16666 ( .A(n8443), .B(n16584), .Z(n16587) );
  INV_X1 U16667 ( .A(n16588), .ZN(n16585) );
  NAND2_X1 U16668 ( .A1(b_13_), .A2(n16589), .ZN(n16588) );
  NOR2_X1 U16669 ( .A1(n16584), .A2(a_13_), .ZN(n16589) );
  XNOR2_X1 U16670 ( .A(n16590), .B(n16591), .ZN(Result_add_12_) );
  NAND2_X1 U16671 ( .A1(n16592), .A2(n13479), .ZN(n16591) );
  NAND2_X1 U16672 ( .A1(n16593), .A2(n16594), .ZN(Result_add_11_) );
  NAND2_X1 U16673 ( .A1(n13828), .A2(n16595), .ZN(n16594) );
  INV_X1 U16674 ( .A(n13613), .ZN(n13828) );
  NOR2_X1 U16675 ( .A1(n16596), .A2(n16597), .ZN(n16593) );
  NOR2_X1 U16676 ( .A1(b_11_), .A2(n16598), .ZN(n16597) );
  XOR2_X1 U16677 ( .A(n8452), .B(n16595), .Z(n16598) );
  INV_X1 U16678 ( .A(n16599), .ZN(n16596) );
  NAND2_X1 U16679 ( .A1(b_11_), .A2(n16600), .ZN(n16599) );
  NOR2_X1 U16680 ( .A1(n16595), .A2(a_11_), .ZN(n16600) );
  XNOR2_X1 U16681 ( .A(n16601), .B(n16602), .ZN(Result_add_10_) );
  NAND2_X1 U16682 ( .A1(n16603), .A2(n13984), .ZN(n16602) );
  XOR2_X1 U16683 ( .A(n16604), .B(n16605), .Z(Result_add_0_) );
  NOR2_X1 U16684 ( .A1(n16606), .A2(n16057), .ZN(n16605) );
  NOR2_X1 U16685 ( .A1(n8690), .A2(n16206), .ZN(n16057) );
  NOR2_X1 U16686 ( .A1(b_0_), .A2(a_0_), .ZN(n16606) );
  NOR2_X1 U16687 ( .A1(n16546), .A2(n16607), .ZN(n16604) );
  NOR2_X1 U16688 ( .A1(n16307), .A2(n16544), .ZN(n16607) );
  NAND2_X1 U16689 ( .A1(n15815), .A2(n16608), .ZN(n16544) );
  NAND2_X1 U16690 ( .A1(n16484), .A2(n16482), .ZN(n16608) );
  NAND2_X1 U16691 ( .A1(n16469), .A2(n16609), .ZN(n16482) );
  NAND2_X1 U16692 ( .A1(n16610), .A2(n16468), .ZN(n16609) );
  NAND2_X1 U16693 ( .A1(n15535), .A2(n16611), .ZN(n16468) );
  NAND2_X1 U16694 ( .A1(n16465), .A2(n16463), .ZN(n16611) );
  NAND2_X1 U16695 ( .A1(n16457), .A2(n16612), .ZN(n16463) );
  NAND2_X1 U16696 ( .A1(n16613), .A2(n16456), .ZN(n16612) );
  NAND2_X1 U16697 ( .A1(n15020), .A2(n16614), .ZN(n16456) );
  NAND2_X1 U16698 ( .A1(n16453), .A2(n16451), .ZN(n16614) );
  NAND2_X1 U16699 ( .A1(n14757), .A2(n16615), .ZN(n16451) );
  NAND2_X1 U16700 ( .A1(n16616), .A2(n16445), .ZN(n16615) );
  NAND2_X1 U16701 ( .A1(n14503), .A2(n16617), .ZN(n16445) );
  NAND2_X1 U16702 ( .A1(n16442), .A2(n16440), .ZN(n16617) );
  NAND2_X1 U16703 ( .A1(n14329), .A2(n16618), .ZN(n16440) );
  NAND2_X1 U16704 ( .A1(n16619), .A2(n16434), .ZN(n16618) );
  NAND2_X1 U16705 ( .A1(n13984), .A2(n16620), .ZN(n16434) );
  NAND2_X1 U16706 ( .A1(n16603), .A2(n16601), .ZN(n16620) );
  NAND2_X1 U16707 ( .A1(n13613), .A2(n16621), .ZN(n16601) );
  NAND2_X1 U16708 ( .A1(n16622), .A2(n16595), .ZN(n16621) );
  NAND2_X1 U16709 ( .A1(n13479), .A2(n16623), .ZN(n16595) );
  NAND2_X1 U16710 ( .A1(n16592), .A2(n16590), .ZN(n16623) );
  NAND2_X1 U16711 ( .A1(n13124), .A2(n16624), .ZN(n16590) );
  NAND2_X1 U16712 ( .A1(n16625), .A2(n16584), .ZN(n16624) );
  NAND2_X1 U16713 ( .A1(n12840), .A2(n16626), .ZN(n16584) );
  NAND2_X1 U16714 ( .A1(n16581), .A2(n16579), .ZN(n16626) );
  NAND2_X1 U16715 ( .A1(n12752), .A2(n16627), .ZN(n16579) );
  NAND2_X1 U16716 ( .A1(n16628), .A2(n16573), .ZN(n16627) );
  INV_X1 U16717 ( .A(n16578), .ZN(n16573) );
  NOR2_X1 U16718 ( .A1(n12361), .A2(n16629), .ZN(n16578) );
  NOR2_X1 U16719 ( .A1(n16570), .A2(n16568), .ZN(n16629) );
  NOR2_X1 U16720 ( .A1(n12114), .A2(n16630), .ZN(n16568) );
  NOR2_X1 U16721 ( .A1(n16631), .A2(n16566), .ZN(n16630) );
  NOR2_X1 U16722 ( .A1(n11871), .A2(n16632), .ZN(n16566) );
  NOR2_X1 U16723 ( .A1(n16559), .A2(n16557), .ZN(n16632) );
  NOR2_X1 U16724 ( .A1(n11740), .A2(n16633), .ZN(n16557) );
  NOR2_X1 U16725 ( .A1(n16634), .A2(n16556), .ZN(n16633) );
  INV_X1 U16726 ( .A(n16551), .ZN(n16556) );
  NAND2_X1 U16727 ( .A1(n11383), .A2(n16635), .ZN(n16551) );
  NAND2_X1 U16728 ( .A1(n16540), .A2(n16538), .ZN(n16635) );
  NAND2_X1 U16729 ( .A1(n16532), .A2(n16636), .ZN(n16538) );
  NAND2_X1 U16730 ( .A1(n16637), .A2(n16531), .ZN(n16636) );
  NAND2_X1 U16731 ( .A1(n10874), .A2(n16638), .ZN(n16531) );
  NAND2_X1 U16732 ( .A1(n16528), .A2(n16526), .ZN(n16638) );
  NAND2_X1 U16733 ( .A1(n10649), .A2(n16639), .ZN(n16526) );
  NAND2_X1 U16734 ( .A1(n16640), .A2(n16520), .ZN(n16639) );
  NAND2_X1 U16735 ( .A1(n10438), .A2(n16641), .ZN(n16520) );
  NAND2_X1 U16736 ( .A1(n16517), .A2(n16515), .ZN(n16641) );
  NAND2_X1 U16737 ( .A1(n10179), .A2(n16642), .ZN(n16515) );
  NAND2_X1 U16738 ( .A1(n16643), .A2(n16509), .ZN(n16642) );
  NAND2_X1 U16739 ( .A1(n9892), .A2(n16644), .ZN(n16509) );
  NAND2_X1 U16740 ( .A1(n16506), .A2(n16504), .ZN(n16644) );
  NAND2_X1 U16741 ( .A1(n9655), .A2(n16645), .ZN(n16504) );
  NAND2_X1 U16742 ( .A1(n16646), .A2(n16498), .ZN(n16645) );
  INV_X1 U16743 ( .A(n16503), .ZN(n16498) );
  NOR2_X1 U16744 ( .A1(n9400), .A2(n16647), .ZN(n16503) );
  NOR2_X1 U16745 ( .A1(n16495), .A2(n16493), .ZN(n16647) );
  NOR2_X1 U16746 ( .A1(n9171), .A2(n16648), .ZN(n16493) );
  NOR2_X1 U16747 ( .A1(n16649), .A2(n16492), .ZN(n16648) );
  INV_X1 U16748 ( .A(n16487), .ZN(n16492) );
  NAND2_X1 U16749 ( .A1(n16650), .A2(n16651), .ZN(n16487) );
  NAND2_X1 U16750 ( .A1(b_30_), .A2(n16479), .ZN(n16651) );
  NAND2_X1 U16751 ( .A1(n16481), .A2(n16203), .ZN(n16479) );
  INV_X1 U16752 ( .A(a_30_), .ZN(n16203) );
  NAND2_X1 U16753 ( .A1(Result_mul_63_), .A2(a_30_), .ZN(n16650) );
  INV_X1 U16754 ( .A(n16481), .ZN(Result_mul_63_) );
  NAND2_X1 U16755 ( .A1(b_31_), .A2(a_31_), .ZN(n16481) );
  NOR2_X1 U16756 ( .A1(b_29_), .A2(a_29_), .ZN(n16649) );
  NOR2_X1 U16757 ( .A1(n8860), .A2(n9161), .ZN(n9171) );
  INV_X1 U16758 ( .A(b_29_), .ZN(n8860) );
  NOR2_X1 U16759 ( .A1(b_28_), .A2(a_28_), .ZN(n16495) );
  NOR2_X1 U16760 ( .A1(n9168), .A2(n8844), .ZN(n9400) );
  INV_X1 U16761 ( .A(b_28_), .ZN(n9168) );
  NAND2_X1 U16762 ( .A1(n9421), .A2(n8839), .ZN(n16646) );
  INV_X1 U16763 ( .A(b_27_), .ZN(n9421) );
  NAND2_X1 U16764 ( .A1(b_27_), .A2(a_27_), .ZN(n9655) );
  NAND2_X1 U16765 ( .A1(n9684), .A2(n8830), .ZN(n16506) );
  INV_X1 U16766 ( .A(b_26_), .ZN(n9684) );
  NAND2_X1 U16767 ( .A1(b_26_), .A2(a_26_), .ZN(n9892) );
  NAND2_X1 U16768 ( .A1(n9924), .A2(n8825), .ZN(n16643) );
  INV_X1 U16769 ( .A(b_25_), .ZN(n9924) );
  NAND2_X1 U16770 ( .A1(b_25_), .A2(a_25_), .ZN(n10179) );
  NAND2_X1 U16771 ( .A1(n10170), .A2(n9131), .ZN(n16517) );
  INV_X1 U16772 ( .A(b_24_), .ZN(n10170) );
  NAND2_X1 U16773 ( .A1(b_24_), .A2(a_24_), .ZN(n10438) );
  NAND2_X1 U16774 ( .A1(n10425), .A2(n8812), .ZN(n16640) );
  INV_X1 U16775 ( .A(b_23_), .ZN(n10425) );
  NAND2_X1 U16776 ( .A1(b_23_), .A2(a_23_), .ZN(n10649) );
  NAND2_X1 U16777 ( .A1(n10701), .A2(n8803), .ZN(n16528) );
  INV_X1 U16778 ( .A(a_22_), .ZN(n8803) );
  INV_X1 U16779 ( .A(b_22_), .ZN(n10701) );
  NAND2_X1 U16780 ( .A1(b_22_), .A2(a_22_), .ZN(n10874) );
  NAND2_X1 U16781 ( .A1(n10931), .A2(n8798), .ZN(n16637) );
  INV_X1 U16782 ( .A(a_21_), .ZN(n8798) );
  INV_X1 U16783 ( .A(b_21_), .ZN(n10931) );
  NAND2_X1 U16784 ( .A1(b_21_), .A2(a_21_), .ZN(n16532) );
  NAND2_X1 U16785 ( .A1(n11196), .A2(n10633), .ZN(n16540) );
  INV_X1 U16786 ( .A(b_20_), .ZN(n11196) );
  NAND2_X1 U16787 ( .A1(b_20_), .A2(a_20_), .ZN(n11383) );
  NOR2_X1 U16788 ( .A1(b_19_), .A2(a_19_), .ZN(n16634) );
  NOR2_X1 U16789 ( .A1(n11452), .A2(n8881), .ZN(n11740) );
  INV_X1 U16790 ( .A(b_19_), .ZN(n11452) );
  NOR2_X1 U16791 ( .A1(b_18_), .A2(a_18_), .ZN(n16559) );
  NOR2_X1 U16792 ( .A1(n11711), .A2(n10616), .ZN(n11871) );
  INV_X1 U16793 ( .A(a_18_), .ZN(n10616) );
  INV_X1 U16794 ( .A(b_18_), .ZN(n11711) );
  NOR2_X1 U16795 ( .A1(b_17_), .A2(a_17_), .ZN(n16631) );
  NOR2_X1 U16796 ( .A1(n11951), .A2(n8772), .ZN(n12114) );
  INV_X1 U16797 ( .A(a_17_), .ZN(n8772) );
  INV_X1 U16798 ( .A(b_17_), .ZN(n11951) );
  NOR2_X1 U16799 ( .A1(b_16_), .A2(a_16_), .ZN(n16570) );
  NOR2_X1 U16800 ( .A1(n12199), .A2(n8768), .ZN(n12361) );
  INV_X1 U16801 ( .A(a_16_), .ZN(n8768) );
  INV_X1 U16802 ( .A(b_16_), .ZN(n12199) );
  NAND2_X1 U16803 ( .A1(n12453), .A2(n8763), .ZN(n16628) );
  INV_X1 U16804 ( .A(b_15_), .ZN(n12453) );
  NAND2_X1 U16805 ( .A1(b_15_), .A2(a_15_), .ZN(n12752) );
  NAND2_X1 U16806 ( .A1(n12723), .A2(n8438), .ZN(n16581) );
  INV_X1 U16807 ( .A(a_14_), .ZN(n8438) );
  INV_X1 U16808 ( .A(b_14_), .ZN(n12723) );
  NAND2_X1 U16809 ( .A1(b_14_), .A2(a_14_), .ZN(n12840) );
  NAND2_X1 U16810 ( .A1(n12942), .A2(n8443), .ZN(n16625) );
  INV_X1 U16811 ( .A(a_13_), .ZN(n8443) );
  INV_X1 U16812 ( .A(b_13_), .ZN(n12942) );
  NAND2_X1 U16813 ( .A1(b_13_), .A2(a_13_), .ZN(n13124) );
  NAND2_X1 U16814 ( .A1(n13233), .A2(n8750), .ZN(n16592) );
  INV_X1 U16815 ( .A(b_12_), .ZN(n13233) );
  NAND2_X1 U16816 ( .A1(b_12_), .A2(a_12_), .ZN(n13479) );
  NAND2_X1 U16817 ( .A1(n13436), .A2(n8452), .ZN(n16622) );
  NAND2_X1 U16818 ( .A1(a_11_), .A2(b_11_), .ZN(n13613) );
  NAND2_X1 U16819 ( .A1(n13725), .A2(n8741), .ZN(n16603) );
  INV_X1 U16820 ( .A(a_10_), .ZN(n8741) );
  NAND2_X1 U16821 ( .A1(a_10_), .A2(b_10_), .ZN(n13984) );
  NAND2_X1 U16822 ( .A1(n13926), .A2(n8736), .ZN(n16619) );
  NAND2_X1 U16823 ( .A1(a_9_), .A2(b_9_), .ZN(n14329) );
  NAND2_X1 U16824 ( .A1(n14216), .A2(n8731), .ZN(n16442) );
  INV_X1 U16825 ( .A(a_8_), .ZN(n8731) );
  NAND2_X1 U16826 ( .A1(a_8_), .A2(b_8_), .ZN(n14503) );
  NAND2_X1 U16827 ( .A1(n14438), .A2(n8726), .ZN(n16616) );
  INV_X1 U16828 ( .A(a_7_), .ZN(n8726) );
  NAND2_X1 U16829 ( .A1(a_7_), .A2(b_7_), .ZN(n14757) );
  NAND2_X1 U16830 ( .A1(n14696), .A2(n8480), .ZN(n16453) );
  INV_X1 U16831 ( .A(b_6_), .ZN(n14696) );
  NAND2_X1 U16832 ( .A1(a_6_), .A2(b_6_), .ZN(n15020) );
  NAND2_X1 U16833 ( .A1(n14947), .A2(n8717), .ZN(n16613) );
  NAND2_X1 U16834 ( .A1(a_5_), .A2(b_5_), .ZN(n16457) );
  NAND2_X1 U16835 ( .A1(n15197), .A2(n8712), .ZN(n16465) );
  NAND2_X1 U16836 ( .A1(a_4_), .A2(b_4_), .ZN(n15535) );
  NAND2_X1 U16837 ( .A1(n15446), .A2(n8707), .ZN(n16610) );
  INV_X1 U16838 ( .A(a_3_), .ZN(n8707) );
  NAND2_X1 U16839 ( .A1(a_3_), .A2(b_3_), .ZN(n16469) );
  NAND2_X1 U16840 ( .A1(n15690), .A2(n8497), .ZN(n16484) );
  NAND2_X1 U16841 ( .A1(a_2_), .A2(b_2_), .ZN(n15815) );
  NOR2_X1 U16842 ( .A1(n8502), .A2(n15994), .ZN(n16307) );
  NOR2_X1 U16843 ( .A1(b_1_), .A2(a_1_), .ZN(n16546) );
endmodule

