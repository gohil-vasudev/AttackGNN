module add_mul_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, operation_0_, operation_1_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, Result_17_, 
        Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, Result_23_, 
        Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, Result_29_, 
        Result_30_, Result_31_, Result_32_, Result_33_, Result_34_, Result_35_, 
        Result_36_, Result_37_, Result_38_, Result_39_, Result_40_, Result_41_, 
        Result_42_, Result_43_, Result_44_, Result_45_, Result_46_, Result_47_, 
        Result_48_, Result_49_, Result_50_, Result_51_, Result_52_, Result_53_, 
        Result_54_, Result_55_, Result_56_, Result_57_, Result_58_, Result_59_, 
        Result_60_, Result_61_, Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179;

  AND2_X2 U8018 ( .A1(n8898), .A2(n8899), .ZN(n7987) );
  AND2_X2 U8019 ( .A1(n8898), .A2(operation_0_), .ZN(n7990) );
  AND2_X2 U8020 ( .A1(n8899), .A2(operation_1_), .ZN(n7989) );
  AND2_X2 U8021 ( .A1(operation_0_), .A2(operation_1_), .ZN(n7956) );
  INV_X2 U8022 ( .A(b_18_), .ZN(n8971) );
  INV_X2 U8023 ( .A(b_16_), .ZN(n8963) );
  INV_X2 U8024 ( .A(b_2_), .ZN(n8907) );
  INV_X2 U8025 ( .A(b_17_), .ZN(n8967) );
  INV_X2 U8026 ( .A(b_15_), .ZN(n8959) );
  INV_X2 U8027 ( .A(b_3_), .ZN(n8911) );
  INV_X2 U8028 ( .A(b_4_), .ZN(n8915) );
  INV_X2 U8029 ( .A(b_5_), .ZN(n8919) );
  INV_X2 U8030 ( .A(b_6_), .ZN(n8923) );
  INV_X2 U8031 ( .A(b_7_), .ZN(n8927) );
  INV_X2 U8032 ( .A(b_11_), .ZN(n8943) );
  INV_X2 U8033 ( .A(b_13_), .ZN(n8951) );
  INV_X2 U8034 ( .A(b_8_), .ZN(n8931) );
  INV_X2 U8035 ( .A(b_9_), .ZN(n8935) );
  INV_X2 U8036 ( .A(b_10_), .ZN(n8939) );
  INV_X2 U8037 ( .A(b_12_), .ZN(n8947) );
  INV_X2 U8038 ( .A(b_14_), .ZN(n8955) );
  INV_X2 U8039 ( .A(b_30_), .ZN(n7998) );
  INV_X2 U8040 ( .A(b_20_), .ZN(n8308) );
  INV_X2 U8041 ( .A(b_28_), .ZN(n8075) );
  INV_X2 U8042 ( .A(b_29_), .ZN(n8047) );
  INV_X2 U8043 ( .A(b_22_), .ZN(n8252) );
  INV_X2 U8044 ( .A(b_21_), .ZN(n8280) );
  INV_X2 U8045 ( .A(b_27_), .ZN(n8112) );
  INV_X2 U8046 ( .A(b_23_), .ZN(n8224) );
  INV_X2 U8047 ( .A(b_19_), .ZN(n8336) );
  INV_X2 U8048 ( .A(b_25_), .ZN(n8168) );
  INV_X2 U8049 ( .A(b_26_), .ZN(n8140) );
  INV_X2 U8050 ( .A(b_24_), .ZN(n8196) );
  OR2_X1 U8051 ( .A1(n7954), .A2(n7955), .ZN(Result_9_) );
  AND2_X1 U8052 ( .A1(n7956), .A2(n7957), .ZN(n7954) );
  XOR2_X1 U8053 ( .A(n7958), .B(n7959), .Z(n7957) );
  AND2_X1 U8054 ( .A1(n7960), .A2(n7961), .ZN(n7959) );
  OR2_X1 U8055 ( .A1(n7962), .A2(n7963), .ZN(n7961) );
  INV_X1 U8056 ( .A(n7964), .ZN(n7960) );
  OR2_X1 U8057 ( .A1(n7965), .A2(n7955), .ZN(Result_8_) );
  AND2_X1 U8058 ( .A1(n7966), .A2(n7956), .ZN(n7965) );
  XOR2_X1 U8059 ( .A(n7967), .B(n7968), .Z(n7966) );
  OR2_X1 U8060 ( .A1(n7969), .A2(n7955), .ZN(Result_7_) );
  AND2_X1 U8061 ( .A1(n7956), .A2(n7970), .ZN(n7969) );
  XOR2_X1 U8062 ( .A(n7971), .B(n7972), .Z(n7970) );
  AND2_X1 U8063 ( .A1(n7973), .A2(n7974), .ZN(n7972) );
  OR2_X1 U8064 ( .A1(n7975), .A2(n7976), .ZN(n7974) );
  INV_X1 U8065 ( .A(n7977), .ZN(n7973) );
  OR2_X1 U8066 ( .A1(n7978), .A2(n7955), .ZN(Result_6_) );
  AND2_X1 U8067 ( .A1(n7979), .A2(n7956), .ZN(n7978) );
  XOR2_X1 U8068 ( .A(n7980), .B(n7981), .Z(n7979) );
  OR2_X1 U8069 ( .A1(n7982), .A2(n7983), .ZN(Result_63_) );
  AND2_X1 U8070 ( .A1(n7984), .A2(n7956), .ZN(n7983) );
  AND2_X1 U8071 ( .A1(n7985), .A2(n7986), .ZN(n7982) );
  OR2_X1 U8072 ( .A1(n7987), .A2(n7988), .ZN(n7986) );
  OR2_X1 U8073 ( .A1(n7989), .A2(n7990), .ZN(n7988) );
  OR2_X1 U8074 ( .A1(n7991), .A2(n7992), .ZN(n7985) );
  OR2_X1 U8075 ( .A1(n7993), .A2(n7994), .ZN(Result_62_) );
  OR2_X1 U8076 ( .A1(n7995), .A2(n7996), .ZN(n7994) );
  AND2_X1 U8077 ( .A1(n7997), .A2(n7998), .ZN(n7996) );
  OR2_X1 U8078 ( .A1(n7999), .A2(n8000), .ZN(n7997) );
  AND2_X1 U8079 ( .A1(n8001), .A2(n8002), .ZN(n8000) );
  AND2_X1 U8080 ( .A1(a_30_), .A2(n8003), .ZN(n7999) );
  AND2_X1 U8081 ( .A1(b_30_), .A2(n8004), .ZN(n7995) );
  OR2_X1 U8082 ( .A1(n8005), .A2(n8006), .ZN(n8004) );
  OR2_X1 U8083 ( .A1(n8007), .A2(n8008), .ZN(n8006) );
  AND2_X1 U8084 ( .A1(a_30_), .A2(n8001), .ZN(n8008) );
  OR2_X1 U8085 ( .A1(n8009), .A2(n8010), .ZN(n8001) );
  OR2_X1 U8086 ( .A1(n8011), .A2(n8012), .ZN(n8010) );
  AND2_X1 U8087 ( .A1(n7990), .A2(n7991), .ZN(n8012) );
  AND2_X1 U8088 ( .A1(n7987), .A2(n7984), .ZN(n8011) );
  AND2_X1 U8089 ( .A1(n7989), .A2(n7992), .ZN(n8009) );
  AND2_X1 U8090 ( .A1(n8003), .A2(n8002), .ZN(n8007) );
  OR2_X1 U8091 ( .A1(n8013), .A2(n8014), .ZN(n8003) );
  OR2_X1 U8092 ( .A1(n8015), .A2(n8016), .ZN(n8014) );
  AND2_X1 U8093 ( .A1(n7990), .A2(n8017), .ZN(n8016) );
  INV_X1 U8094 ( .A(n7991), .ZN(n8017) );
  AND2_X1 U8095 ( .A1(n7987), .A2(n8018), .ZN(n8015) );
  AND2_X1 U8096 ( .A1(n7989), .A2(n8019), .ZN(n8013) );
  INV_X1 U8097 ( .A(n7992), .ZN(n8019) );
  AND2_X1 U8098 ( .A1(n7956), .A2(n8020), .ZN(n8005) );
  OR2_X1 U8099 ( .A1(n7991), .A2(n8021), .ZN(n8020) );
  AND2_X1 U8100 ( .A1(n8022), .A2(n7956), .ZN(n7993) );
  AND2_X1 U8101 ( .A1(a_30_), .A2(n8023), .ZN(n8022) );
  OR2_X1 U8102 ( .A1(n8024), .A2(n7992), .ZN(n8023) );
  AND2_X1 U8103 ( .A1(b_31_), .A2(n7998), .ZN(n8024) );
  OR2_X1 U8104 ( .A1(n8025), .A2(n8026), .ZN(Result_61_) );
  OR2_X1 U8105 ( .A1(n8027), .A2(n8028), .ZN(n8026) );
  AND2_X1 U8106 ( .A1(n8029), .A2(n8030), .ZN(n8028) );
  OR2_X1 U8107 ( .A1(n8031), .A2(n8032), .ZN(n8030) );
  OR2_X1 U8108 ( .A1(n8033), .A2(n8034), .ZN(n8032) );
  AND2_X1 U8109 ( .A1(n7990), .A2(n8035), .ZN(n8034) );
  AND2_X1 U8110 ( .A1(n7987), .A2(n8036), .ZN(n8033) );
  INV_X1 U8111 ( .A(n8037), .ZN(n8036) );
  AND2_X1 U8112 ( .A1(n7989), .A2(n8038), .ZN(n8031) );
  INV_X1 U8113 ( .A(n8039), .ZN(n8029) );
  AND2_X1 U8114 ( .A1(n8039), .A2(n8040), .ZN(n8027) );
  OR2_X1 U8115 ( .A1(n8041), .A2(n8042), .ZN(n8040) );
  OR2_X1 U8116 ( .A1(n8043), .A2(n8044), .ZN(n8042) );
  AND2_X1 U8117 ( .A1(n7990), .A2(n8045), .ZN(n8044) );
  INV_X1 U8118 ( .A(n8035), .ZN(n8045) );
  AND2_X1 U8119 ( .A1(n8037), .A2(n7987), .ZN(n8043) );
  AND2_X1 U8120 ( .A1(n7989), .A2(n8046), .ZN(n8041) );
  INV_X1 U8121 ( .A(n8038), .ZN(n8046) );
  XNOR2_X1 U8122 ( .A(a_29_), .B(n8047), .ZN(n8039) );
  AND2_X1 U8123 ( .A1(n8048), .A2(n7956), .ZN(n8025) );
  XNOR2_X1 U8124 ( .A(n8049), .B(n8050), .ZN(n8048) );
  XNOR2_X1 U8125 ( .A(n8051), .B(n8052), .ZN(n8049) );
  OR2_X1 U8126 ( .A1(n8053), .A2(n8054), .ZN(Result_60_) );
  OR2_X1 U8127 ( .A1(n8055), .A2(n8056), .ZN(n8054) );
  AND2_X1 U8128 ( .A1(n8057), .A2(n8058), .ZN(n8056) );
  OR2_X1 U8129 ( .A1(n8059), .A2(n8060), .ZN(n8058) );
  OR2_X1 U8130 ( .A1(n8061), .A2(n8062), .ZN(n8060) );
  AND2_X1 U8131 ( .A1(n7990), .A2(n8063), .ZN(n8062) );
  AND2_X1 U8132 ( .A1(n8064), .A2(n7987), .ZN(n8061) );
  INV_X1 U8133 ( .A(n8065), .ZN(n8064) );
  AND2_X1 U8134 ( .A1(n7989), .A2(n8066), .ZN(n8059) );
  INV_X1 U8135 ( .A(n8067), .ZN(n8057) );
  AND2_X1 U8136 ( .A1(n8067), .A2(n8068), .ZN(n8055) );
  OR2_X1 U8137 ( .A1(n8069), .A2(n8070), .ZN(n8068) );
  OR2_X1 U8138 ( .A1(n8071), .A2(n8072), .ZN(n8070) );
  AND2_X1 U8139 ( .A1(n7990), .A2(n8073), .ZN(n8072) );
  INV_X1 U8140 ( .A(n8063), .ZN(n8073) );
  AND2_X1 U8141 ( .A1(n7987), .A2(n8065), .ZN(n8071) );
  AND2_X1 U8142 ( .A1(n7989), .A2(n8074), .ZN(n8069) );
  INV_X1 U8143 ( .A(n8066), .ZN(n8074) );
  XNOR2_X1 U8144 ( .A(a_28_), .B(n8075), .ZN(n8067) );
  AND2_X1 U8145 ( .A1(n8076), .A2(n7956), .ZN(n8053) );
  XNOR2_X1 U8146 ( .A(n8077), .B(n8078), .ZN(n8076) );
  XOR2_X1 U8147 ( .A(n8079), .B(n8080), .Z(n8078) );
  OR2_X1 U8148 ( .A1(n8081), .A2(n7955), .ZN(Result_5_) );
  AND2_X1 U8149 ( .A1(n7956), .A2(n8082), .ZN(n8081) );
  XOR2_X1 U8150 ( .A(n8083), .B(n8084), .Z(n8082) );
  AND2_X1 U8151 ( .A1(n8085), .A2(n8086), .ZN(n8084) );
  OR2_X1 U8152 ( .A1(n8087), .A2(n8088), .ZN(n8086) );
  INV_X1 U8153 ( .A(n8089), .ZN(n8085) );
  OR2_X1 U8154 ( .A1(n8090), .A2(n8091), .ZN(Result_59_) );
  OR2_X1 U8155 ( .A1(n8092), .A2(n8093), .ZN(n8091) );
  AND2_X1 U8156 ( .A1(n8094), .A2(n8095), .ZN(n8093) );
  OR2_X1 U8157 ( .A1(n8096), .A2(n8097), .ZN(n8095) );
  OR2_X1 U8158 ( .A1(n8098), .A2(n8099), .ZN(n8097) );
  AND2_X1 U8159 ( .A1(n7990), .A2(n8100), .ZN(n8099) );
  AND2_X1 U8160 ( .A1(n8101), .A2(n7987), .ZN(n8098) );
  INV_X1 U8161 ( .A(n8102), .ZN(n8101) );
  AND2_X1 U8162 ( .A1(n7989), .A2(n8103), .ZN(n8096) );
  INV_X1 U8163 ( .A(n8104), .ZN(n8094) );
  AND2_X1 U8164 ( .A1(n8104), .A2(n8105), .ZN(n8092) );
  OR2_X1 U8165 ( .A1(n8106), .A2(n8107), .ZN(n8105) );
  OR2_X1 U8166 ( .A1(n8108), .A2(n8109), .ZN(n8107) );
  AND2_X1 U8167 ( .A1(n7990), .A2(n8110), .ZN(n8109) );
  INV_X1 U8168 ( .A(n8100), .ZN(n8110) );
  AND2_X1 U8169 ( .A1(n7987), .A2(n8102), .ZN(n8108) );
  AND2_X1 U8170 ( .A1(n7989), .A2(n8111), .ZN(n8106) );
  INV_X1 U8171 ( .A(n8103), .ZN(n8111) );
  XNOR2_X1 U8172 ( .A(a_27_), .B(n8112), .ZN(n8104) );
  AND2_X1 U8173 ( .A1(n8113), .A2(n7956), .ZN(n8090) );
  XNOR2_X1 U8174 ( .A(n8114), .B(n8115), .ZN(n8113) );
  XOR2_X1 U8175 ( .A(n8116), .B(n8117), .Z(n8115) );
  OR2_X1 U8176 ( .A1(n8118), .A2(n8119), .ZN(Result_58_) );
  OR2_X1 U8177 ( .A1(n8120), .A2(n8121), .ZN(n8119) );
  AND2_X1 U8178 ( .A1(n8122), .A2(n8123), .ZN(n8121) );
  OR2_X1 U8179 ( .A1(n8124), .A2(n8125), .ZN(n8123) );
  OR2_X1 U8180 ( .A1(n8126), .A2(n8127), .ZN(n8125) );
  AND2_X1 U8181 ( .A1(n7990), .A2(n8128), .ZN(n8127) );
  AND2_X1 U8182 ( .A1(n8129), .A2(n7987), .ZN(n8126) );
  INV_X1 U8183 ( .A(n8130), .ZN(n8129) );
  AND2_X1 U8184 ( .A1(n7989), .A2(n8131), .ZN(n8124) );
  INV_X1 U8185 ( .A(n8132), .ZN(n8122) );
  AND2_X1 U8186 ( .A1(n8132), .A2(n8133), .ZN(n8120) );
  OR2_X1 U8187 ( .A1(n8134), .A2(n8135), .ZN(n8133) );
  OR2_X1 U8188 ( .A1(n8136), .A2(n8137), .ZN(n8135) );
  AND2_X1 U8189 ( .A1(n7990), .A2(n8138), .ZN(n8137) );
  INV_X1 U8190 ( .A(n8128), .ZN(n8138) );
  AND2_X1 U8191 ( .A1(n7987), .A2(n8130), .ZN(n8136) );
  AND2_X1 U8192 ( .A1(n7989), .A2(n8139), .ZN(n8134) );
  INV_X1 U8193 ( .A(n8131), .ZN(n8139) );
  XNOR2_X1 U8194 ( .A(a_26_), .B(n8140), .ZN(n8132) );
  AND2_X1 U8195 ( .A1(n8141), .A2(n7956), .ZN(n8118) );
  XNOR2_X1 U8196 ( .A(n8142), .B(n8143), .ZN(n8141) );
  XOR2_X1 U8197 ( .A(n8144), .B(n8145), .Z(n8143) );
  OR2_X1 U8198 ( .A1(n8146), .A2(n8147), .ZN(Result_57_) );
  OR2_X1 U8199 ( .A1(n8148), .A2(n8149), .ZN(n8147) );
  AND2_X1 U8200 ( .A1(n8150), .A2(n8151), .ZN(n8149) );
  OR2_X1 U8201 ( .A1(n8152), .A2(n8153), .ZN(n8151) );
  OR2_X1 U8202 ( .A1(n8154), .A2(n8155), .ZN(n8153) );
  AND2_X1 U8203 ( .A1(n7990), .A2(n8156), .ZN(n8155) );
  AND2_X1 U8204 ( .A1(n8157), .A2(n7987), .ZN(n8154) );
  INV_X1 U8205 ( .A(n8158), .ZN(n8157) );
  AND2_X1 U8206 ( .A1(n7989), .A2(n8159), .ZN(n8152) );
  INV_X1 U8207 ( .A(n8160), .ZN(n8150) );
  AND2_X1 U8208 ( .A1(n8160), .A2(n8161), .ZN(n8148) );
  OR2_X1 U8209 ( .A1(n8162), .A2(n8163), .ZN(n8161) );
  OR2_X1 U8210 ( .A1(n8164), .A2(n8165), .ZN(n8163) );
  AND2_X1 U8211 ( .A1(n7990), .A2(n8166), .ZN(n8165) );
  INV_X1 U8212 ( .A(n8156), .ZN(n8166) );
  AND2_X1 U8213 ( .A1(n7987), .A2(n8158), .ZN(n8164) );
  AND2_X1 U8214 ( .A1(n7989), .A2(n8167), .ZN(n8162) );
  INV_X1 U8215 ( .A(n8159), .ZN(n8167) );
  XNOR2_X1 U8216 ( .A(a_25_), .B(n8168), .ZN(n8160) );
  AND2_X1 U8217 ( .A1(n8169), .A2(n7956), .ZN(n8146) );
  XNOR2_X1 U8218 ( .A(n8170), .B(n8171), .ZN(n8169) );
  XOR2_X1 U8219 ( .A(n8172), .B(n8173), .Z(n8171) );
  OR2_X1 U8220 ( .A1(n8174), .A2(n8175), .ZN(Result_56_) );
  OR2_X1 U8221 ( .A1(n8176), .A2(n8177), .ZN(n8175) );
  AND2_X1 U8222 ( .A1(n8178), .A2(n8179), .ZN(n8177) );
  OR2_X1 U8223 ( .A1(n8180), .A2(n8181), .ZN(n8179) );
  OR2_X1 U8224 ( .A1(n8182), .A2(n8183), .ZN(n8181) );
  AND2_X1 U8225 ( .A1(n7990), .A2(n8184), .ZN(n8183) );
  AND2_X1 U8226 ( .A1(n8185), .A2(n7987), .ZN(n8182) );
  INV_X1 U8227 ( .A(n8186), .ZN(n8185) );
  AND2_X1 U8228 ( .A1(n7989), .A2(n8187), .ZN(n8180) );
  INV_X1 U8229 ( .A(n8188), .ZN(n8178) );
  AND2_X1 U8230 ( .A1(n8188), .A2(n8189), .ZN(n8176) );
  OR2_X1 U8231 ( .A1(n8190), .A2(n8191), .ZN(n8189) );
  OR2_X1 U8232 ( .A1(n8192), .A2(n8193), .ZN(n8191) );
  AND2_X1 U8233 ( .A1(n7990), .A2(n8194), .ZN(n8193) );
  INV_X1 U8234 ( .A(n8184), .ZN(n8194) );
  AND2_X1 U8235 ( .A1(n7987), .A2(n8186), .ZN(n8192) );
  AND2_X1 U8236 ( .A1(n7989), .A2(n8195), .ZN(n8190) );
  INV_X1 U8237 ( .A(n8187), .ZN(n8195) );
  XNOR2_X1 U8238 ( .A(a_24_), .B(n8196), .ZN(n8188) );
  AND2_X1 U8239 ( .A1(n8197), .A2(n7956), .ZN(n8174) );
  XNOR2_X1 U8240 ( .A(n8198), .B(n8199), .ZN(n8197) );
  XOR2_X1 U8241 ( .A(n8200), .B(n8201), .Z(n8199) );
  OR2_X1 U8242 ( .A1(n8202), .A2(n8203), .ZN(Result_55_) );
  OR2_X1 U8243 ( .A1(n8204), .A2(n8205), .ZN(n8203) );
  AND2_X1 U8244 ( .A1(n8206), .A2(n8207), .ZN(n8205) );
  OR2_X1 U8245 ( .A1(n8208), .A2(n8209), .ZN(n8207) );
  OR2_X1 U8246 ( .A1(n8210), .A2(n8211), .ZN(n8209) );
  AND2_X1 U8247 ( .A1(n7990), .A2(n8212), .ZN(n8211) );
  AND2_X1 U8248 ( .A1(n8213), .A2(n7987), .ZN(n8210) );
  INV_X1 U8249 ( .A(n8214), .ZN(n8213) );
  AND2_X1 U8250 ( .A1(n7989), .A2(n8215), .ZN(n8208) );
  INV_X1 U8251 ( .A(n8216), .ZN(n8206) );
  AND2_X1 U8252 ( .A1(n8216), .A2(n8217), .ZN(n8204) );
  OR2_X1 U8253 ( .A1(n8218), .A2(n8219), .ZN(n8217) );
  OR2_X1 U8254 ( .A1(n8220), .A2(n8221), .ZN(n8219) );
  AND2_X1 U8255 ( .A1(n7990), .A2(n8222), .ZN(n8221) );
  INV_X1 U8256 ( .A(n8212), .ZN(n8222) );
  AND2_X1 U8257 ( .A1(n7987), .A2(n8214), .ZN(n8220) );
  AND2_X1 U8258 ( .A1(n7989), .A2(n8223), .ZN(n8218) );
  INV_X1 U8259 ( .A(n8215), .ZN(n8223) );
  XNOR2_X1 U8260 ( .A(a_23_), .B(n8224), .ZN(n8216) );
  AND2_X1 U8261 ( .A1(n8225), .A2(n7956), .ZN(n8202) );
  XNOR2_X1 U8262 ( .A(n8226), .B(n8227), .ZN(n8225) );
  XOR2_X1 U8263 ( .A(n8228), .B(n8229), .Z(n8227) );
  OR2_X1 U8264 ( .A1(n8230), .A2(n8231), .ZN(Result_54_) );
  OR2_X1 U8265 ( .A1(n8232), .A2(n8233), .ZN(n8231) );
  AND2_X1 U8266 ( .A1(n8234), .A2(n8235), .ZN(n8233) );
  OR2_X1 U8267 ( .A1(n8236), .A2(n8237), .ZN(n8235) );
  OR2_X1 U8268 ( .A1(n8238), .A2(n8239), .ZN(n8237) );
  AND2_X1 U8269 ( .A1(n7990), .A2(n8240), .ZN(n8239) );
  AND2_X1 U8270 ( .A1(n8241), .A2(n7987), .ZN(n8238) );
  INV_X1 U8271 ( .A(n8242), .ZN(n8241) );
  AND2_X1 U8272 ( .A1(n7989), .A2(n8243), .ZN(n8236) );
  INV_X1 U8273 ( .A(n8244), .ZN(n8234) );
  AND2_X1 U8274 ( .A1(n8244), .A2(n8245), .ZN(n8232) );
  OR2_X1 U8275 ( .A1(n8246), .A2(n8247), .ZN(n8245) );
  OR2_X1 U8276 ( .A1(n8248), .A2(n8249), .ZN(n8247) );
  AND2_X1 U8277 ( .A1(n7990), .A2(n8250), .ZN(n8249) );
  INV_X1 U8278 ( .A(n8240), .ZN(n8250) );
  AND2_X1 U8279 ( .A1(n7987), .A2(n8242), .ZN(n8248) );
  AND2_X1 U8280 ( .A1(n7989), .A2(n8251), .ZN(n8246) );
  INV_X1 U8281 ( .A(n8243), .ZN(n8251) );
  XNOR2_X1 U8282 ( .A(a_22_), .B(n8252), .ZN(n8244) );
  AND2_X1 U8283 ( .A1(n8253), .A2(n7956), .ZN(n8230) );
  XNOR2_X1 U8284 ( .A(n8254), .B(n8255), .ZN(n8253) );
  XOR2_X1 U8285 ( .A(n8256), .B(n8257), .Z(n8255) );
  OR2_X1 U8286 ( .A1(n8258), .A2(n8259), .ZN(Result_53_) );
  OR2_X1 U8287 ( .A1(n8260), .A2(n8261), .ZN(n8259) );
  AND2_X1 U8288 ( .A1(n8262), .A2(n8263), .ZN(n8261) );
  OR2_X1 U8289 ( .A1(n8264), .A2(n8265), .ZN(n8263) );
  OR2_X1 U8290 ( .A1(n8266), .A2(n8267), .ZN(n8265) );
  AND2_X1 U8291 ( .A1(n7990), .A2(n8268), .ZN(n8267) );
  AND2_X1 U8292 ( .A1(n8269), .A2(n7987), .ZN(n8266) );
  INV_X1 U8293 ( .A(n8270), .ZN(n8269) );
  AND2_X1 U8294 ( .A1(n7989), .A2(n8271), .ZN(n8264) );
  INV_X1 U8295 ( .A(n8272), .ZN(n8262) );
  AND2_X1 U8296 ( .A1(n8272), .A2(n8273), .ZN(n8260) );
  OR2_X1 U8297 ( .A1(n8274), .A2(n8275), .ZN(n8273) );
  OR2_X1 U8298 ( .A1(n8276), .A2(n8277), .ZN(n8275) );
  AND2_X1 U8299 ( .A1(n7990), .A2(n8278), .ZN(n8277) );
  INV_X1 U8300 ( .A(n8268), .ZN(n8278) );
  AND2_X1 U8301 ( .A1(n7987), .A2(n8270), .ZN(n8276) );
  AND2_X1 U8302 ( .A1(n7989), .A2(n8279), .ZN(n8274) );
  INV_X1 U8303 ( .A(n8271), .ZN(n8279) );
  XNOR2_X1 U8304 ( .A(a_21_), .B(n8280), .ZN(n8272) );
  AND2_X1 U8305 ( .A1(n8281), .A2(n7956), .ZN(n8258) );
  XNOR2_X1 U8306 ( .A(n8282), .B(n8283), .ZN(n8281) );
  XOR2_X1 U8307 ( .A(n8284), .B(n8285), .Z(n8283) );
  OR2_X1 U8308 ( .A1(n8286), .A2(n8287), .ZN(Result_52_) );
  OR2_X1 U8309 ( .A1(n8288), .A2(n8289), .ZN(n8287) );
  AND2_X1 U8310 ( .A1(n8290), .A2(n8291), .ZN(n8289) );
  OR2_X1 U8311 ( .A1(n8292), .A2(n8293), .ZN(n8291) );
  OR2_X1 U8312 ( .A1(n8294), .A2(n8295), .ZN(n8293) );
  AND2_X1 U8313 ( .A1(n7990), .A2(n8296), .ZN(n8295) );
  AND2_X1 U8314 ( .A1(n8297), .A2(n7987), .ZN(n8294) );
  INV_X1 U8315 ( .A(n8298), .ZN(n8297) );
  AND2_X1 U8316 ( .A1(n7989), .A2(n8299), .ZN(n8292) );
  INV_X1 U8317 ( .A(n8300), .ZN(n8290) );
  AND2_X1 U8318 ( .A1(n8300), .A2(n8301), .ZN(n8288) );
  OR2_X1 U8319 ( .A1(n8302), .A2(n8303), .ZN(n8301) );
  OR2_X1 U8320 ( .A1(n8304), .A2(n8305), .ZN(n8303) );
  AND2_X1 U8321 ( .A1(n7990), .A2(n8306), .ZN(n8305) );
  INV_X1 U8322 ( .A(n8296), .ZN(n8306) );
  AND2_X1 U8323 ( .A1(n7987), .A2(n8298), .ZN(n8304) );
  AND2_X1 U8324 ( .A1(n7989), .A2(n8307), .ZN(n8302) );
  INV_X1 U8325 ( .A(n8299), .ZN(n8307) );
  XNOR2_X1 U8326 ( .A(a_20_), .B(n8308), .ZN(n8300) );
  AND2_X1 U8327 ( .A1(n8309), .A2(n7956), .ZN(n8286) );
  XNOR2_X1 U8328 ( .A(n8310), .B(n8311), .ZN(n8309) );
  XOR2_X1 U8329 ( .A(n8312), .B(n8313), .Z(n8311) );
  OR2_X1 U8330 ( .A1(n8314), .A2(n8315), .ZN(Result_51_) );
  OR2_X1 U8331 ( .A1(n8316), .A2(n8317), .ZN(n8315) );
  AND2_X1 U8332 ( .A1(n8318), .A2(n8319), .ZN(n8317) );
  OR2_X1 U8333 ( .A1(n8320), .A2(n8321), .ZN(n8319) );
  OR2_X1 U8334 ( .A1(n8322), .A2(n8323), .ZN(n8321) );
  AND2_X1 U8335 ( .A1(n7990), .A2(n8324), .ZN(n8323) );
  AND2_X1 U8336 ( .A1(n8325), .A2(n7987), .ZN(n8322) );
  INV_X1 U8337 ( .A(n8326), .ZN(n8325) );
  AND2_X1 U8338 ( .A1(n7989), .A2(n8327), .ZN(n8320) );
  INV_X1 U8339 ( .A(n8328), .ZN(n8318) );
  AND2_X1 U8340 ( .A1(n8328), .A2(n8329), .ZN(n8316) );
  OR2_X1 U8341 ( .A1(n8330), .A2(n8331), .ZN(n8329) );
  OR2_X1 U8342 ( .A1(n8332), .A2(n8333), .ZN(n8331) );
  AND2_X1 U8343 ( .A1(n7990), .A2(n8334), .ZN(n8333) );
  INV_X1 U8344 ( .A(n8324), .ZN(n8334) );
  AND2_X1 U8345 ( .A1(n7987), .A2(n8326), .ZN(n8332) );
  AND2_X1 U8346 ( .A1(n7989), .A2(n8335), .ZN(n8330) );
  INV_X1 U8347 ( .A(n8327), .ZN(n8335) );
  XNOR2_X1 U8348 ( .A(a_19_), .B(n8336), .ZN(n8328) );
  AND2_X1 U8349 ( .A1(n8337), .A2(n7956), .ZN(n8314) );
  XNOR2_X1 U8350 ( .A(n8338), .B(n8339), .ZN(n8337) );
  XOR2_X1 U8351 ( .A(n8340), .B(n8341), .Z(n8339) );
  OR2_X1 U8352 ( .A1(n8342), .A2(n8343), .ZN(Result_50_) );
  OR2_X1 U8353 ( .A1(n8344), .A2(n8345), .ZN(n8343) );
  AND2_X1 U8354 ( .A1(n8346), .A2(n8347), .ZN(n8345) );
  OR2_X1 U8355 ( .A1(n8348), .A2(n8349), .ZN(n8347) );
  OR2_X1 U8356 ( .A1(n8350), .A2(n8351), .ZN(n8349) );
  AND2_X1 U8357 ( .A1(n7990), .A2(n8352), .ZN(n8351) );
  INV_X1 U8358 ( .A(n8353), .ZN(n8352) );
  AND2_X1 U8359 ( .A1(n7987), .A2(n8354), .ZN(n8350) );
  AND2_X1 U8360 ( .A1(n7989), .A2(n8355), .ZN(n8348) );
  INV_X1 U8361 ( .A(n8356), .ZN(n8355) );
  AND2_X1 U8362 ( .A1(n8357), .A2(n8358), .ZN(n8344) );
  INV_X1 U8363 ( .A(n8346), .ZN(n8358) );
  AND2_X1 U8364 ( .A1(n8359), .A2(n8360), .ZN(n8346) );
  OR2_X1 U8365 ( .A1(a_18_), .A2(b_18_), .ZN(n8359) );
  OR2_X1 U8366 ( .A1(n8361), .A2(n8362), .ZN(n8357) );
  OR2_X1 U8367 ( .A1(n8363), .A2(n8364), .ZN(n8362) );
  AND2_X1 U8368 ( .A1(n7990), .A2(n8353), .ZN(n8364) );
  AND2_X1 U8369 ( .A1(n8365), .A2(n7987), .ZN(n8363) );
  INV_X1 U8370 ( .A(n8354), .ZN(n8365) );
  AND2_X1 U8371 ( .A1(n7989), .A2(n8356), .ZN(n8361) );
  AND2_X1 U8372 ( .A1(n8366), .A2(n7956), .ZN(n8342) );
  XNOR2_X1 U8373 ( .A(n8367), .B(n8368), .ZN(n8366) );
  XOR2_X1 U8374 ( .A(n8369), .B(n8370), .Z(n8368) );
  OR2_X1 U8375 ( .A1(n8371), .A2(n7955), .ZN(Result_4_) );
  AND2_X1 U8376 ( .A1(n8372), .A2(n7956), .ZN(n8371) );
  XOR2_X1 U8377 ( .A(n8373), .B(n8374), .Z(n8372) );
  OR2_X1 U8378 ( .A1(n8375), .A2(n8376), .ZN(Result_49_) );
  OR2_X1 U8379 ( .A1(n8377), .A2(n8378), .ZN(n8376) );
  AND2_X1 U8380 ( .A1(n8379), .A2(n8380), .ZN(n8378) );
  OR2_X1 U8381 ( .A1(n8381), .A2(n8382), .ZN(n8380) );
  OR2_X1 U8382 ( .A1(n8383), .A2(n8384), .ZN(n8382) );
  AND2_X1 U8383 ( .A1(n7990), .A2(n8385), .ZN(n8384) );
  INV_X1 U8384 ( .A(n8386), .ZN(n8385) );
  AND2_X1 U8385 ( .A1(n7987), .A2(n8387), .ZN(n8383) );
  AND2_X1 U8386 ( .A1(n7989), .A2(n8388), .ZN(n8381) );
  INV_X1 U8387 ( .A(n8389), .ZN(n8388) );
  AND2_X1 U8388 ( .A1(n8390), .A2(n8391), .ZN(n8377) );
  INV_X1 U8389 ( .A(n8379), .ZN(n8391) );
  AND2_X1 U8390 ( .A1(n8392), .A2(n8393), .ZN(n8379) );
  OR2_X1 U8391 ( .A1(a_17_), .A2(b_17_), .ZN(n8392) );
  OR2_X1 U8392 ( .A1(n8394), .A2(n8395), .ZN(n8390) );
  OR2_X1 U8393 ( .A1(n8396), .A2(n8397), .ZN(n8395) );
  AND2_X1 U8394 ( .A1(n7990), .A2(n8386), .ZN(n8397) );
  AND2_X1 U8395 ( .A1(n8398), .A2(n7987), .ZN(n8396) );
  INV_X1 U8396 ( .A(n8387), .ZN(n8398) );
  AND2_X1 U8397 ( .A1(n7989), .A2(n8389), .ZN(n8394) );
  AND2_X1 U8398 ( .A1(n8399), .A2(n7956), .ZN(n8375) );
  XNOR2_X1 U8399 ( .A(n8400), .B(n8401), .ZN(n8399) );
  XOR2_X1 U8400 ( .A(n8402), .B(n8403), .Z(n8401) );
  OR2_X1 U8401 ( .A1(n8404), .A2(n8405), .ZN(Result_48_) );
  OR2_X1 U8402 ( .A1(n8406), .A2(n8407), .ZN(n8405) );
  AND2_X1 U8403 ( .A1(n8408), .A2(n8409), .ZN(n8407) );
  OR2_X1 U8404 ( .A1(n8410), .A2(n8411), .ZN(n8409) );
  OR2_X1 U8405 ( .A1(n8412), .A2(n8413), .ZN(n8411) );
  AND2_X1 U8406 ( .A1(n7990), .A2(n8414), .ZN(n8413) );
  INV_X1 U8407 ( .A(n8415), .ZN(n8414) );
  AND2_X1 U8408 ( .A1(n7987), .A2(n8416), .ZN(n8412) );
  AND2_X1 U8409 ( .A1(n7989), .A2(n8417), .ZN(n8410) );
  INV_X1 U8410 ( .A(n8418), .ZN(n8417) );
  AND2_X1 U8411 ( .A1(n8419), .A2(n8420), .ZN(n8406) );
  INV_X1 U8412 ( .A(n8408), .ZN(n8420) );
  AND2_X1 U8413 ( .A1(n8421), .A2(n8422), .ZN(n8408) );
  OR2_X1 U8414 ( .A1(a_16_), .A2(b_16_), .ZN(n8421) );
  OR2_X1 U8415 ( .A1(n8423), .A2(n8424), .ZN(n8419) );
  OR2_X1 U8416 ( .A1(n8425), .A2(n8426), .ZN(n8424) );
  AND2_X1 U8417 ( .A1(n7990), .A2(n8415), .ZN(n8426) );
  AND2_X1 U8418 ( .A1(n8427), .A2(n7987), .ZN(n8425) );
  INV_X1 U8419 ( .A(n8416), .ZN(n8427) );
  AND2_X1 U8420 ( .A1(n7989), .A2(n8418), .ZN(n8423) );
  AND2_X1 U8421 ( .A1(n8428), .A2(n7956), .ZN(n8404) );
  XNOR2_X1 U8422 ( .A(n8429), .B(n8430), .ZN(n8428) );
  XOR2_X1 U8423 ( .A(n8431), .B(n8432), .Z(n8430) );
  OR2_X1 U8424 ( .A1(n8433), .A2(n8434), .ZN(Result_47_) );
  OR2_X1 U8425 ( .A1(n8435), .A2(n8436), .ZN(n8434) );
  AND2_X1 U8426 ( .A1(n8437), .A2(n8438), .ZN(n8436) );
  OR2_X1 U8427 ( .A1(n8439), .A2(n8440), .ZN(n8438) );
  OR2_X1 U8428 ( .A1(n8441), .A2(n8442), .ZN(n8440) );
  AND2_X1 U8429 ( .A1(n7990), .A2(n8443), .ZN(n8442) );
  INV_X1 U8430 ( .A(n8444), .ZN(n8443) );
  AND2_X1 U8431 ( .A1(n7987), .A2(n8445), .ZN(n8441) );
  AND2_X1 U8432 ( .A1(n7989), .A2(n8446), .ZN(n8439) );
  INV_X1 U8433 ( .A(n8447), .ZN(n8446) );
  AND2_X1 U8434 ( .A1(n8448), .A2(n8449), .ZN(n8435) );
  INV_X1 U8435 ( .A(n8437), .ZN(n8449) );
  AND2_X1 U8436 ( .A1(n8450), .A2(n8451), .ZN(n8437) );
  OR2_X1 U8437 ( .A1(a_15_), .A2(b_15_), .ZN(n8450) );
  OR2_X1 U8438 ( .A1(n8452), .A2(n8453), .ZN(n8448) );
  OR2_X1 U8439 ( .A1(n8454), .A2(n8455), .ZN(n8453) );
  AND2_X1 U8440 ( .A1(n7990), .A2(n8444), .ZN(n8455) );
  AND2_X1 U8441 ( .A1(n8456), .A2(n7987), .ZN(n8454) );
  INV_X1 U8442 ( .A(n8445), .ZN(n8456) );
  AND2_X1 U8443 ( .A1(n7989), .A2(n8447), .ZN(n8452) );
  AND2_X1 U8444 ( .A1(n8457), .A2(n7956), .ZN(n8433) );
  XNOR2_X1 U8445 ( .A(n8458), .B(n8459), .ZN(n8457) );
  XOR2_X1 U8446 ( .A(n8460), .B(n8461), .Z(n8459) );
  OR2_X1 U8447 ( .A1(n8462), .A2(n8463), .ZN(Result_46_) );
  OR2_X1 U8448 ( .A1(n8464), .A2(n8465), .ZN(n8463) );
  AND2_X1 U8449 ( .A1(n8466), .A2(n8467), .ZN(n8465) );
  OR2_X1 U8450 ( .A1(n8468), .A2(n8469), .ZN(n8467) );
  OR2_X1 U8451 ( .A1(n8470), .A2(n8471), .ZN(n8469) );
  AND2_X1 U8452 ( .A1(n7990), .A2(n8472), .ZN(n8471) );
  INV_X1 U8453 ( .A(n8473), .ZN(n8472) );
  AND2_X1 U8454 ( .A1(n7987), .A2(n8474), .ZN(n8470) );
  AND2_X1 U8455 ( .A1(n7989), .A2(n8475), .ZN(n8468) );
  INV_X1 U8456 ( .A(n8476), .ZN(n8475) );
  AND2_X1 U8457 ( .A1(n8477), .A2(n8478), .ZN(n8464) );
  INV_X1 U8458 ( .A(n8466), .ZN(n8478) );
  AND2_X1 U8459 ( .A1(n8479), .A2(n8480), .ZN(n8466) );
  OR2_X1 U8460 ( .A1(a_14_), .A2(b_14_), .ZN(n8479) );
  OR2_X1 U8461 ( .A1(n8481), .A2(n8482), .ZN(n8477) );
  OR2_X1 U8462 ( .A1(n8483), .A2(n8484), .ZN(n8482) );
  AND2_X1 U8463 ( .A1(n7990), .A2(n8473), .ZN(n8484) );
  AND2_X1 U8464 ( .A1(n8485), .A2(n7987), .ZN(n8483) );
  INV_X1 U8465 ( .A(n8474), .ZN(n8485) );
  AND2_X1 U8466 ( .A1(n7989), .A2(n8476), .ZN(n8481) );
  AND2_X1 U8467 ( .A1(n8486), .A2(n7956), .ZN(n8462) );
  XNOR2_X1 U8468 ( .A(n8487), .B(n8488), .ZN(n8486) );
  XOR2_X1 U8469 ( .A(n8489), .B(n8490), .Z(n8488) );
  OR2_X1 U8470 ( .A1(n8491), .A2(n8492), .ZN(Result_45_) );
  OR2_X1 U8471 ( .A1(n8493), .A2(n8494), .ZN(n8492) );
  AND2_X1 U8472 ( .A1(n8495), .A2(n8496), .ZN(n8494) );
  OR2_X1 U8473 ( .A1(n8497), .A2(n8498), .ZN(n8496) );
  OR2_X1 U8474 ( .A1(n8499), .A2(n8500), .ZN(n8498) );
  AND2_X1 U8475 ( .A1(n7990), .A2(n8501), .ZN(n8500) );
  INV_X1 U8476 ( .A(n8502), .ZN(n8501) );
  AND2_X1 U8477 ( .A1(n7987), .A2(n8503), .ZN(n8499) );
  AND2_X1 U8478 ( .A1(n7989), .A2(n8504), .ZN(n8497) );
  INV_X1 U8479 ( .A(n8505), .ZN(n8504) );
  AND2_X1 U8480 ( .A1(n8506), .A2(n8507), .ZN(n8493) );
  INV_X1 U8481 ( .A(n8495), .ZN(n8507) );
  AND2_X1 U8482 ( .A1(n8508), .A2(n8509), .ZN(n8495) );
  OR2_X1 U8483 ( .A1(a_13_), .A2(b_13_), .ZN(n8508) );
  OR2_X1 U8484 ( .A1(n8510), .A2(n8511), .ZN(n8506) );
  OR2_X1 U8485 ( .A1(n8512), .A2(n8513), .ZN(n8511) );
  AND2_X1 U8486 ( .A1(n7990), .A2(n8502), .ZN(n8513) );
  AND2_X1 U8487 ( .A1(n8514), .A2(n7987), .ZN(n8512) );
  INV_X1 U8488 ( .A(n8503), .ZN(n8514) );
  AND2_X1 U8489 ( .A1(n7989), .A2(n8505), .ZN(n8510) );
  AND2_X1 U8490 ( .A1(n8515), .A2(n7956), .ZN(n8491) );
  XNOR2_X1 U8491 ( .A(n8516), .B(n8517), .ZN(n8515) );
  XOR2_X1 U8492 ( .A(n8518), .B(n8519), .Z(n8517) );
  OR2_X1 U8493 ( .A1(n8520), .A2(n8521), .ZN(Result_44_) );
  OR2_X1 U8494 ( .A1(n8522), .A2(n8523), .ZN(n8521) );
  AND2_X1 U8495 ( .A1(n8524), .A2(n8525), .ZN(n8523) );
  OR2_X1 U8496 ( .A1(n8526), .A2(n8527), .ZN(n8525) );
  OR2_X1 U8497 ( .A1(n8528), .A2(n8529), .ZN(n8527) );
  AND2_X1 U8498 ( .A1(n7990), .A2(n8530), .ZN(n8529) );
  INV_X1 U8499 ( .A(n8531), .ZN(n8530) );
  AND2_X1 U8500 ( .A1(n7987), .A2(n8532), .ZN(n8528) );
  AND2_X1 U8501 ( .A1(n7989), .A2(n8533), .ZN(n8526) );
  INV_X1 U8502 ( .A(n8534), .ZN(n8533) );
  AND2_X1 U8503 ( .A1(n8535), .A2(n8536), .ZN(n8522) );
  INV_X1 U8504 ( .A(n8524), .ZN(n8536) );
  AND2_X1 U8505 ( .A1(n8537), .A2(n8538), .ZN(n8524) );
  OR2_X1 U8506 ( .A1(a_12_), .A2(b_12_), .ZN(n8537) );
  OR2_X1 U8507 ( .A1(n8539), .A2(n8540), .ZN(n8535) );
  OR2_X1 U8508 ( .A1(n8541), .A2(n8542), .ZN(n8540) );
  AND2_X1 U8509 ( .A1(n7990), .A2(n8531), .ZN(n8542) );
  AND2_X1 U8510 ( .A1(n8543), .A2(n7987), .ZN(n8541) );
  INV_X1 U8511 ( .A(n8532), .ZN(n8543) );
  AND2_X1 U8512 ( .A1(n7989), .A2(n8534), .ZN(n8539) );
  AND2_X1 U8513 ( .A1(n8544), .A2(n7956), .ZN(n8520) );
  XNOR2_X1 U8514 ( .A(n8545), .B(n8546), .ZN(n8544) );
  XOR2_X1 U8515 ( .A(n8547), .B(n8548), .Z(n8546) );
  OR2_X1 U8516 ( .A1(n8549), .A2(n8550), .ZN(Result_43_) );
  OR2_X1 U8517 ( .A1(n8551), .A2(n8552), .ZN(n8550) );
  AND2_X1 U8518 ( .A1(n8553), .A2(n8554), .ZN(n8552) );
  OR2_X1 U8519 ( .A1(n8555), .A2(n8556), .ZN(n8554) );
  OR2_X1 U8520 ( .A1(n8557), .A2(n8558), .ZN(n8556) );
  AND2_X1 U8521 ( .A1(n7990), .A2(n8559), .ZN(n8558) );
  INV_X1 U8522 ( .A(n8560), .ZN(n8559) );
  AND2_X1 U8523 ( .A1(n7987), .A2(n8561), .ZN(n8557) );
  AND2_X1 U8524 ( .A1(n7989), .A2(n8562), .ZN(n8555) );
  INV_X1 U8525 ( .A(n8563), .ZN(n8562) );
  AND2_X1 U8526 ( .A1(n8564), .A2(n8565), .ZN(n8551) );
  INV_X1 U8527 ( .A(n8553), .ZN(n8565) );
  AND2_X1 U8528 ( .A1(n8566), .A2(n8567), .ZN(n8553) );
  OR2_X1 U8529 ( .A1(a_11_), .A2(b_11_), .ZN(n8566) );
  OR2_X1 U8530 ( .A1(n8568), .A2(n8569), .ZN(n8564) );
  OR2_X1 U8531 ( .A1(n8570), .A2(n8571), .ZN(n8569) );
  AND2_X1 U8532 ( .A1(n7990), .A2(n8560), .ZN(n8571) );
  AND2_X1 U8533 ( .A1(n8572), .A2(n7987), .ZN(n8570) );
  INV_X1 U8534 ( .A(n8561), .ZN(n8572) );
  AND2_X1 U8535 ( .A1(n7989), .A2(n8563), .ZN(n8568) );
  AND2_X1 U8536 ( .A1(n8573), .A2(n7956), .ZN(n8549) );
  XNOR2_X1 U8537 ( .A(n8574), .B(n8575), .ZN(n8573) );
  XOR2_X1 U8538 ( .A(n8576), .B(n8577), .Z(n8575) );
  OR2_X1 U8539 ( .A1(n8578), .A2(n8579), .ZN(Result_42_) );
  OR2_X1 U8540 ( .A1(n8580), .A2(n8581), .ZN(n8579) );
  AND2_X1 U8541 ( .A1(n8582), .A2(n8583), .ZN(n8581) );
  OR2_X1 U8542 ( .A1(n8584), .A2(n8585), .ZN(n8583) );
  OR2_X1 U8543 ( .A1(n8586), .A2(n8587), .ZN(n8585) );
  AND2_X1 U8544 ( .A1(n7990), .A2(n8588), .ZN(n8587) );
  INV_X1 U8545 ( .A(n8589), .ZN(n8588) );
  AND2_X1 U8546 ( .A1(n7987), .A2(n8590), .ZN(n8586) );
  AND2_X1 U8547 ( .A1(n7989), .A2(n8591), .ZN(n8584) );
  INV_X1 U8548 ( .A(n8592), .ZN(n8591) );
  AND2_X1 U8549 ( .A1(n8593), .A2(n8594), .ZN(n8580) );
  INV_X1 U8550 ( .A(n8582), .ZN(n8594) );
  AND2_X1 U8551 ( .A1(n8595), .A2(n8596), .ZN(n8582) );
  OR2_X1 U8552 ( .A1(a_10_), .A2(b_10_), .ZN(n8595) );
  OR2_X1 U8553 ( .A1(n8597), .A2(n8598), .ZN(n8593) );
  OR2_X1 U8554 ( .A1(n8599), .A2(n8600), .ZN(n8598) );
  AND2_X1 U8555 ( .A1(n7990), .A2(n8589), .ZN(n8600) );
  AND2_X1 U8556 ( .A1(n8601), .A2(n7987), .ZN(n8599) );
  INV_X1 U8557 ( .A(n8590), .ZN(n8601) );
  AND2_X1 U8558 ( .A1(n7989), .A2(n8592), .ZN(n8597) );
  AND2_X1 U8559 ( .A1(n8602), .A2(n7956), .ZN(n8578) );
  XNOR2_X1 U8560 ( .A(n8603), .B(n8604), .ZN(n8602) );
  XOR2_X1 U8561 ( .A(n8605), .B(n8606), .Z(n8604) );
  OR2_X1 U8562 ( .A1(n8607), .A2(n8608), .ZN(Result_41_) );
  OR2_X1 U8563 ( .A1(n8609), .A2(n8610), .ZN(n8608) );
  AND2_X1 U8564 ( .A1(n8611), .A2(n8612), .ZN(n8610) );
  OR2_X1 U8565 ( .A1(n8613), .A2(n8614), .ZN(n8612) );
  OR2_X1 U8566 ( .A1(n8615), .A2(n8616), .ZN(n8614) );
  AND2_X1 U8567 ( .A1(n7990), .A2(n8617), .ZN(n8616) );
  INV_X1 U8568 ( .A(n8618), .ZN(n8617) );
  AND2_X1 U8569 ( .A1(n7987), .A2(n8619), .ZN(n8615) );
  AND2_X1 U8570 ( .A1(n7989), .A2(n8620), .ZN(n8613) );
  INV_X1 U8571 ( .A(n8621), .ZN(n8620) );
  AND2_X1 U8572 ( .A1(n8622), .A2(n8623), .ZN(n8609) );
  INV_X1 U8573 ( .A(n8611), .ZN(n8623) );
  AND2_X1 U8574 ( .A1(n8624), .A2(n8625), .ZN(n8611) );
  OR2_X1 U8575 ( .A1(a_9_), .A2(b_9_), .ZN(n8624) );
  OR2_X1 U8576 ( .A1(n8626), .A2(n8627), .ZN(n8622) );
  OR2_X1 U8577 ( .A1(n8628), .A2(n8629), .ZN(n8627) );
  AND2_X1 U8578 ( .A1(n7990), .A2(n8618), .ZN(n8629) );
  AND2_X1 U8579 ( .A1(n8630), .A2(n7987), .ZN(n8628) );
  INV_X1 U8580 ( .A(n8619), .ZN(n8630) );
  AND2_X1 U8581 ( .A1(n7989), .A2(n8621), .ZN(n8626) );
  AND2_X1 U8582 ( .A1(n8631), .A2(n7956), .ZN(n8607) );
  XNOR2_X1 U8583 ( .A(n8632), .B(n8633), .ZN(n8631) );
  XOR2_X1 U8584 ( .A(n8634), .B(n8635), .Z(n8633) );
  OR2_X1 U8585 ( .A1(n8636), .A2(n8637), .ZN(Result_40_) );
  OR2_X1 U8586 ( .A1(n8638), .A2(n8639), .ZN(n8637) );
  AND2_X1 U8587 ( .A1(n8640), .A2(n8641), .ZN(n8639) );
  OR2_X1 U8588 ( .A1(n8642), .A2(n8643), .ZN(n8641) );
  OR2_X1 U8589 ( .A1(n8644), .A2(n8645), .ZN(n8643) );
  AND2_X1 U8590 ( .A1(n7990), .A2(n8646), .ZN(n8645) );
  INV_X1 U8591 ( .A(n8647), .ZN(n8646) );
  AND2_X1 U8592 ( .A1(n7987), .A2(n8648), .ZN(n8644) );
  AND2_X1 U8593 ( .A1(n7989), .A2(n8649), .ZN(n8642) );
  INV_X1 U8594 ( .A(n8650), .ZN(n8649) );
  AND2_X1 U8595 ( .A1(n8651), .A2(n8652), .ZN(n8638) );
  INV_X1 U8596 ( .A(n8640), .ZN(n8652) );
  AND2_X1 U8597 ( .A1(n8653), .A2(n8654), .ZN(n8640) );
  OR2_X1 U8598 ( .A1(a_8_), .A2(b_8_), .ZN(n8653) );
  OR2_X1 U8599 ( .A1(n8655), .A2(n8656), .ZN(n8651) );
  OR2_X1 U8600 ( .A1(n8657), .A2(n8658), .ZN(n8656) );
  AND2_X1 U8601 ( .A1(n7990), .A2(n8647), .ZN(n8658) );
  AND2_X1 U8602 ( .A1(n8659), .A2(n7987), .ZN(n8657) );
  INV_X1 U8603 ( .A(n8648), .ZN(n8659) );
  AND2_X1 U8604 ( .A1(n7989), .A2(n8650), .ZN(n8655) );
  AND2_X1 U8605 ( .A1(n8660), .A2(n7956), .ZN(n8636) );
  XNOR2_X1 U8606 ( .A(n8661), .B(n8662), .ZN(n8660) );
  XOR2_X1 U8607 ( .A(n8663), .B(n8664), .Z(n8662) );
  OR2_X1 U8608 ( .A1(n8665), .A2(n7955), .ZN(Result_3_) );
  AND2_X1 U8609 ( .A1(n7956), .A2(n8666), .ZN(n8665) );
  XOR2_X1 U8610 ( .A(n8667), .B(n8668), .Z(n8666) );
  AND2_X1 U8611 ( .A1(n8669), .A2(n8670), .ZN(n8668) );
  OR2_X1 U8612 ( .A1(n8671), .A2(n8672), .ZN(n8670) );
  INV_X1 U8613 ( .A(n8673), .ZN(n8669) );
  OR2_X1 U8614 ( .A1(n8674), .A2(n8675), .ZN(Result_39_) );
  OR2_X1 U8615 ( .A1(n8676), .A2(n8677), .ZN(n8675) );
  AND2_X1 U8616 ( .A1(n8678), .A2(n8679), .ZN(n8677) );
  OR2_X1 U8617 ( .A1(n8680), .A2(n8681), .ZN(n8679) );
  OR2_X1 U8618 ( .A1(n8682), .A2(n8683), .ZN(n8681) );
  AND2_X1 U8619 ( .A1(n7990), .A2(n8684), .ZN(n8683) );
  INV_X1 U8620 ( .A(n8685), .ZN(n8684) );
  AND2_X1 U8621 ( .A1(n7987), .A2(n8686), .ZN(n8682) );
  AND2_X1 U8622 ( .A1(n7989), .A2(n8687), .ZN(n8680) );
  INV_X1 U8623 ( .A(n8688), .ZN(n8687) );
  AND2_X1 U8624 ( .A1(n8689), .A2(n8690), .ZN(n8676) );
  INV_X1 U8625 ( .A(n8678), .ZN(n8690) );
  AND2_X1 U8626 ( .A1(n8691), .A2(n8692), .ZN(n8678) );
  OR2_X1 U8627 ( .A1(a_7_), .A2(b_7_), .ZN(n8691) );
  OR2_X1 U8628 ( .A1(n8693), .A2(n8694), .ZN(n8689) );
  OR2_X1 U8629 ( .A1(n8695), .A2(n8696), .ZN(n8694) );
  AND2_X1 U8630 ( .A1(n7990), .A2(n8685), .ZN(n8696) );
  AND2_X1 U8631 ( .A1(n8697), .A2(n7987), .ZN(n8695) );
  INV_X1 U8632 ( .A(n8686), .ZN(n8697) );
  AND2_X1 U8633 ( .A1(n7989), .A2(n8688), .ZN(n8693) );
  AND2_X1 U8634 ( .A1(n8698), .A2(n7956), .ZN(n8674) );
  XNOR2_X1 U8635 ( .A(n8699), .B(n8700), .ZN(n8698) );
  XOR2_X1 U8636 ( .A(n8701), .B(n8702), .Z(n8700) );
  OR2_X1 U8637 ( .A1(n8703), .A2(n8704), .ZN(Result_38_) );
  OR2_X1 U8638 ( .A1(n8705), .A2(n8706), .ZN(n8704) );
  AND2_X1 U8639 ( .A1(n8707), .A2(n8708), .ZN(n8706) );
  OR2_X1 U8640 ( .A1(n8709), .A2(n8710), .ZN(n8708) );
  OR2_X1 U8641 ( .A1(n8711), .A2(n8712), .ZN(n8710) );
  AND2_X1 U8642 ( .A1(n7990), .A2(n8713), .ZN(n8712) );
  INV_X1 U8643 ( .A(n8714), .ZN(n8713) );
  AND2_X1 U8644 ( .A1(n7987), .A2(n8715), .ZN(n8711) );
  AND2_X1 U8645 ( .A1(n7989), .A2(n8716), .ZN(n8709) );
  INV_X1 U8646 ( .A(n8717), .ZN(n8716) );
  AND2_X1 U8647 ( .A1(n8718), .A2(n8719), .ZN(n8705) );
  INV_X1 U8648 ( .A(n8707), .ZN(n8719) );
  AND2_X1 U8649 ( .A1(n8720), .A2(n8721), .ZN(n8707) );
  OR2_X1 U8650 ( .A1(a_6_), .A2(b_6_), .ZN(n8720) );
  OR2_X1 U8651 ( .A1(n8722), .A2(n8723), .ZN(n8718) );
  OR2_X1 U8652 ( .A1(n8724), .A2(n8725), .ZN(n8723) );
  AND2_X1 U8653 ( .A1(n7990), .A2(n8714), .ZN(n8725) );
  AND2_X1 U8654 ( .A1(n8726), .A2(n7987), .ZN(n8724) );
  INV_X1 U8655 ( .A(n8715), .ZN(n8726) );
  AND2_X1 U8656 ( .A1(n7989), .A2(n8717), .ZN(n8722) );
  AND2_X1 U8657 ( .A1(n8727), .A2(n7956), .ZN(n8703) );
  XNOR2_X1 U8658 ( .A(n8728), .B(n8729), .ZN(n8727) );
  XOR2_X1 U8659 ( .A(n8730), .B(n8731), .Z(n8729) );
  OR2_X1 U8660 ( .A1(n8732), .A2(n8733), .ZN(Result_37_) );
  OR2_X1 U8661 ( .A1(n8734), .A2(n8735), .ZN(n8733) );
  AND2_X1 U8662 ( .A1(n8736), .A2(n8737), .ZN(n8735) );
  OR2_X1 U8663 ( .A1(n8738), .A2(n8739), .ZN(n8737) );
  OR2_X1 U8664 ( .A1(n8740), .A2(n8741), .ZN(n8739) );
  AND2_X1 U8665 ( .A1(n7990), .A2(n8742), .ZN(n8741) );
  INV_X1 U8666 ( .A(n8743), .ZN(n8742) );
  AND2_X1 U8667 ( .A1(n7987), .A2(n8744), .ZN(n8740) );
  AND2_X1 U8668 ( .A1(n7989), .A2(n8745), .ZN(n8738) );
  INV_X1 U8669 ( .A(n8746), .ZN(n8745) );
  AND2_X1 U8670 ( .A1(n8747), .A2(n8748), .ZN(n8734) );
  INV_X1 U8671 ( .A(n8736), .ZN(n8748) );
  AND2_X1 U8672 ( .A1(n8749), .A2(n8750), .ZN(n8736) );
  OR2_X1 U8673 ( .A1(a_5_), .A2(b_5_), .ZN(n8749) );
  OR2_X1 U8674 ( .A1(n8751), .A2(n8752), .ZN(n8747) );
  OR2_X1 U8675 ( .A1(n8753), .A2(n8754), .ZN(n8752) );
  AND2_X1 U8676 ( .A1(n7990), .A2(n8743), .ZN(n8754) );
  AND2_X1 U8677 ( .A1(n8755), .A2(n7987), .ZN(n8753) );
  INV_X1 U8678 ( .A(n8744), .ZN(n8755) );
  AND2_X1 U8679 ( .A1(n7989), .A2(n8746), .ZN(n8751) );
  AND2_X1 U8680 ( .A1(n8756), .A2(n7956), .ZN(n8732) );
  XNOR2_X1 U8681 ( .A(n8757), .B(n8758), .ZN(n8756) );
  XOR2_X1 U8682 ( .A(n8759), .B(n8760), .Z(n8758) );
  OR2_X1 U8683 ( .A1(n8761), .A2(n8762), .ZN(Result_36_) );
  OR2_X1 U8684 ( .A1(n8763), .A2(n8764), .ZN(n8762) );
  AND2_X1 U8685 ( .A1(n8765), .A2(n8766), .ZN(n8764) );
  OR2_X1 U8686 ( .A1(n8767), .A2(n8768), .ZN(n8766) );
  OR2_X1 U8687 ( .A1(n8769), .A2(n8770), .ZN(n8768) );
  AND2_X1 U8688 ( .A1(n7990), .A2(n8771), .ZN(n8770) );
  INV_X1 U8689 ( .A(n8772), .ZN(n8771) );
  AND2_X1 U8690 ( .A1(n7987), .A2(n8773), .ZN(n8769) );
  AND2_X1 U8691 ( .A1(n7989), .A2(n8774), .ZN(n8767) );
  INV_X1 U8692 ( .A(n8775), .ZN(n8774) );
  AND2_X1 U8693 ( .A1(n8776), .A2(n8777), .ZN(n8763) );
  INV_X1 U8694 ( .A(n8765), .ZN(n8777) );
  AND2_X1 U8695 ( .A1(n8778), .A2(n8779), .ZN(n8765) );
  OR2_X1 U8696 ( .A1(a_4_), .A2(b_4_), .ZN(n8778) );
  OR2_X1 U8697 ( .A1(n8780), .A2(n8781), .ZN(n8776) );
  OR2_X1 U8698 ( .A1(n8782), .A2(n8783), .ZN(n8781) );
  AND2_X1 U8699 ( .A1(n7990), .A2(n8772), .ZN(n8783) );
  AND2_X1 U8700 ( .A1(n8784), .A2(n7987), .ZN(n8782) );
  INV_X1 U8701 ( .A(n8773), .ZN(n8784) );
  AND2_X1 U8702 ( .A1(n7989), .A2(n8775), .ZN(n8780) );
  AND2_X1 U8703 ( .A1(n8785), .A2(n7956), .ZN(n8761) );
  XNOR2_X1 U8704 ( .A(n8786), .B(n8787), .ZN(n8785) );
  XOR2_X1 U8705 ( .A(n8788), .B(n8789), .Z(n8787) );
  OR2_X1 U8706 ( .A1(n8790), .A2(n8791), .ZN(Result_35_) );
  OR2_X1 U8707 ( .A1(n8792), .A2(n8793), .ZN(n8791) );
  AND2_X1 U8708 ( .A1(n8794), .A2(n8795), .ZN(n8793) );
  OR2_X1 U8709 ( .A1(n8796), .A2(n8797), .ZN(n8795) );
  OR2_X1 U8710 ( .A1(n8798), .A2(n8799), .ZN(n8797) );
  AND2_X1 U8711 ( .A1(n7990), .A2(n8800), .ZN(n8799) );
  INV_X1 U8712 ( .A(n8801), .ZN(n8800) );
  AND2_X1 U8713 ( .A1(n7987), .A2(n8802), .ZN(n8798) );
  AND2_X1 U8714 ( .A1(n7989), .A2(n8803), .ZN(n8796) );
  INV_X1 U8715 ( .A(n8804), .ZN(n8803) );
  AND2_X1 U8716 ( .A1(n8805), .A2(n8806), .ZN(n8792) );
  INV_X1 U8717 ( .A(n8794), .ZN(n8806) );
  AND2_X1 U8718 ( .A1(n8807), .A2(n8808), .ZN(n8794) );
  OR2_X1 U8719 ( .A1(a_3_), .A2(b_3_), .ZN(n8807) );
  OR2_X1 U8720 ( .A1(n8809), .A2(n8810), .ZN(n8805) );
  OR2_X1 U8721 ( .A1(n8811), .A2(n8812), .ZN(n8810) );
  AND2_X1 U8722 ( .A1(n7990), .A2(n8801), .ZN(n8812) );
  AND2_X1 U8723 ( .A1(n8813), .A2(n7987), .ZN(n8811) );
  INV_X1 U8724 ( .A(n8802), .ZN(n8813) );
  AND2_X1 U8725 ( .A1(n7989), .A2(n8804), .ZN(n8809) );
  AND2_X1 U8726 ( .A1(n8814), .A2(n7956), .ZN(n8790) );
  XNOR2_X1 U8727 ( .A(n8815), .B(n8816), .ZN(n8814) );
  XOR2_X1 U8728 ( .A(n8817), .B(n8818), .Z(n8816) );
  OR2_X1 U8729 ( .A1(n8819), .A2(n8820), .ZN(Result_34_) );
  OR2_X1 U8730 ( .A1(n8821), .A2(n8822), .ZN(n8820) );
  AND2_X1 U8731 ( .A1(n8823), .A2(n8824), .ZN(n8822) );
  OR2_X1 U8732 ( .A1(n8825), .A2(n8826), .ZN(n8824) );
  OR2_X1 U8733 ( .A1(n8827), .A2(n8828), .ZN(n8826) );
  AND2_X1 U8734 ( .A1(n7990), .A2(n8829), .ZN(n8828) );
  INV_X1 U8735 ( .A(n8830), .ZN(n8829) );
  AND2_X1 U8736 ( .A1(n7987), .A2(n8831), .ZN(n8827) );
  AND2_X1 U8737 ( .A1(n7989), .A2(n8832), .ZN(n8825) );
  INV_X1 U8738 ( .A(n8833), .ZN(n8832) );
  AND2_X1 U8739 ( .A1(n8834), .A2(n8835), .ZN(n8821) );
  INV_X1 U8740 ( .A(n8823), .ZN(n8835) );
  AND2_X1 U8741 ( .A1(n8836), .A2(n8837), .ZN(n8823) );
  OR2_X1 U8742 ( .A1(a_2_), .A2(b_2_), .ZN(n8836) );
  OR2_X1 U8743 ( .A1(n8838), .A2(n8839), .ZN(n8834) );
  OR2_X1 U8744 ( .A1(n8840), .A2(n8841), .ZN(n8839) );
  AND2_X1 U8745 ( .A1(n7990), .A2(n8830), .ZN(n8841) );
  AND2_X1 U8746 ( .A1(n8842), .A2(n7987), .ZN(n8840) );
  INV_X1 U8747 ( .A(n8831), .ZN(n8842) );
  AND2_X1 U8748 ( .A1(n7989), .A2(n8833), .ZN(n8838) );
  AND2_X1 U8749 ( .A1(n8843), .A2(n7956), .ZN(n8819) );
  XNOR2_X1 U8750 ( .A(n8844), .B(n8845), .ZN(n8843) );
  XOR2_X1 U8751 ( .A(n8846), .B(n8847), .Z(n8845) );
  OR2_X1 U8752 ( .A1(n8848), .A2(n8849), .ZN(Result_33_) );
  OR2_X1 U8753 ( .A1(n8850), .A2(n8851), .ZN(n8849) );
  AND2_X1 U8754 ( .A1(n8852), .A2(n8853), .ZN(n8851) );
  OR2_X1 U8755 ( .A1(n8854), .A2(n8855), .ZN(n8853) );
  OR2_X1 U8756 ( .A1(n8856), .A2(n8857), .ZN(n8855) );
  AND2_X1 U8757 ( .A1(n7990), .A2(n8858), .ZN(n8857) );
  INV_X1 U8758 ( .A(n8859), .ZN(n8858) );
  AND2_X1 U8759 ( .A1(n7987), .A2(n8860), .ZN(n8856) );
  AND2_X1 U8760 ( .A1(n7989), .A2(n8861), .ZN(n8854) );
  INV_X1 U8761 ( .A(n8862), .ZN(n8861) );
  AND2_X1 U8762 ( .A1(n8863), .A2(n8864), .ZN(n8850) );
  INV_X1 U8763 ( .A(n8852), .ZN(n8864) );
  AND2_X1 U8764 ( .A1(n8865), .A2(n8866), .ZN(n8852) );
  OR2_X1 U8765 ( .A1(a_1_), .A2(b_1_), .ZN(n8865) );
  OR2_X1 U8766 ( .A1(n8867), .A2(n8868), .ZN(n8863) );
  OR2_X1 U8767 ( .A1(n8869), .A2(n8870), .ZN(n8868) );
  AND2_X1 U8768 ( .A1(n7990), .A2(n8859), .ZN(n8870) );
  AND2_X1 U8769 ( .A1(n8871), .A2(n7987), .ZN(n8869) );
  INV_X1 U8770 ( .A(n8860), .ZN(n8871) );
  AND2_X1 U8771 ( .A1(n7989), .A2(n8862), .ZN(n8867) );
  AND2_X1 U8772 ( .A1(n8872), .A2(n7956), .ZN(n8848) );
  XNOR2_X1 U8773 ( .A(n8873), .B(n8874), .ZN(n8872) );
  XOR2_X1 U8774 ( .A(n8875), .B(n8876), .Z(n8874) );
  OR2_X1 U8775 ( .A1(n8877), .A2(n8878), .ZN(Result_32_) );
  OR2_X1 U8776 ( .A1(n8879), .A2(n8880), .ZN(n8878) );
  AND2_X1 U8777 ( .A1(n8881), .A2(n8882), .ZN(n8880) );
  OR2_X1 U8778 ( .A1(n8883), .A2(n8884), .ZN(n8881) );
  OR2_X1 U8779 ( .A1(n8885), .A2(n8886), .ZN(n8884) );
  AND2_X1 U8780 ( .A1(n7990), .A2(n8887), .ZN(n8886) );
  INV_X1 U8781 ( .A(n8888), .ZN(n8887) );
  AND2_X1 U8782 ( .A1(n7987), .A2(n8889), .ZN(n8885) );
  AND2_X1 U8783 ( .A1(n8890), .A2(n7989), .ZN(n8883) );
  AND2_X1 U8784 ( .A1(n8891), .A2(n8892), .ZN(n8879) );
  OR2_X1 U8785 ( .A1(n8893), .A2(n8894), .ZN(n8892) );
  OR2_X1 U8786 ( .A1(n8895), .A2(n8896), .ZN(n8894) );
  AND2_X1 U8787 ( .A1(n7990), .A2(n8888), .ZN(n8896) );
  AND2_X1 U8788 ( .A1(n8897), .A2(n7987), .ZN(n8895) );
  INV_X1 U8789 ( .A(n8889), .ZN(n8897) );
  OR2_X1 U8790 ( .A1(n8900), .A2(n8901), .ZN(n8889) );
  AND2_X1 U8791 ( .A1(n8902), .A2(n8903), .ZN(n8901) );
  AND2_X1 U8792 ( .A1(n8860), .A2(n8866), .ZN(n8900) );
  OR2_X1 U8793 ( .A1(n8904), .A2(n8905), .ZN(n8860) );
  AND2_X1 U8794 ( .A1(n8906), .A2(n8907), .ZN(n8905) );
  AND2_X1 U8795 ( .A1(n8831), .A2(n8837), .ZN(n8904) );
  OR2_X1 U8796 ( .A1(n8908), .A2(n8909), .ZN(n8831) );
  AND2_X1 U8797 ( .A1(n8910), .A2(n8911), .ZN(n8909) );
  AND2_X1 U8798 ( .A1(n8802), .A2(n8808), .ZN(n8908) );
  OR2_X1 U8799 ( .A1(n8912), .A2(n8913), .ZN(n8802) );
  AND2_X1 U8800 ( .A1(n8914), .A2(n8915), .ZN(n8913) );
  AND2_X1 U8801 ( .A1(n8773), .A2(n8779), .ZN(n8912) );
  OR2_X1 U8802 ( .A1(n8916), .A2(n8917), .ZN(n8773) );
  AND2_X1 U8803 ( .A1(n8918), .A2(n8919), .ZN(n8917) );
  AND2_X1 U8804 ( .A1(n8744), .A2(n8750), .ZN(n8916) );
  OR2_X1 U8805 ( .A1(n8920), .A2(n8921), .ZN(n8744) );
  AND2_X1 U8806 ( .A1(n8922), .A2(n8923), .ZN(n8921) );
  AND2_X1 U8807 ( .A1(n8715), .A2(n8721), .ZN(n8920) );
  OR2_X1 U8808 ( .A1(n8924), .A2(n8925), .ZN(n8715) );
  AND2_X1 U8809 ( .A1(n8926), .A2(n8927), .ZN(n8925) );
  AND2_X1 U8810 ( .A1(n8686), .A2(n8692), .ZN(n8924) );
  OR2_X1 U8811 ( .A1(n8928), .A2(n8929), .ZN(n8686) );
  AND2_X1 U8812 ( .A1(n8930), .A2(n8931), .ZN(n8929) );
  AND2_X1 U8813 ( .A1(n8648), .A2(n8654), .ZN(n8928) );
  OR2_X1 U8814 ( .A1(n8932), .A2(n8933), .ZN(n8648) );
  AND2_X1 U8815 ( .A1(n8934), .A2(n8935), .ZN(n8933) );
  AND2_X1 U8816 ( .A1(n8619), .A2(n8625), .ZN(n8932) );
  OR2_X1 U8817 ( .A1(n8936), .A2(n8937), .ZN(n8619) );
  AND2_X1 U8818 ( .A1(n8938), .A2(n8939), .ZN(n8937) );
  AND2_X1 U8819 ( .A1(n8590), .A2(n8596), .ZN(n8936) );
  OR2_X1 U8820 ( .A1(n8940), .A2(n8941), .ZN(n8590) );
  AND2_X1 U8821 ( .A1(n8942), .A2(n8943), .ZN(n8941) );
  AND2_X1 U8822 ( .A1(n8561), .A2(n8567), .ZN(n8940) );
  OR2_X1 U8823 ( .A1(n8944), .A2(n8945), .ZN(n8561) );
  AND2_X1 U8824 ( .A1(n8946), .A2(n8947), .ZN(n8945) );
  AND2_X1 U8825 ( .A1(n8532), .A2(n8538), .ZN(n8944) );
  OR2_X1 U8826 ( .A1(n8948), .A2(n8949), .ZN(n8532) );
  AND2_X1 U8827 ( .A1(n8950), .A2(n8951), .ZN(n8949) );
  AND2_X1 U8828 ( .A1(n8503), .A2(n8509), .ZN(n8948) );
  OR2_X1 U8829 ( .A1(n8952), .A2(n8953), .ZN(n8503) );
  AND2_X1 U8830 ( .A1(n8954), .A2(n8955), .ZN(n8953) );
  AND2_X1 U8831 ( .A1(n8474), .A2(n8480), .ZN(n8952) );
  OR2_X1 U8832 ( .A1(n8956), .A2(n8957), .ZN(n8474) );
  AND2_X1 U8833 ( .A1(n8958), .A2(n8959), .ZN(n8957) );
  AND2_X1 U8834 ( .A1(n8445), .A2(n8451), .ZN(n8956) );
  OR2_X1 U8835 ( .A1(n8960), .A2(n8961), .ZN(n8445) );
  AND2_X1 U8836 ( .A1(n8962), .A2(n8963), .ZN(n8961) );
  AND2_X1 U8837 ( .A1(n8416), .A2(n8422), .ZN(n8960) );
  OR2_X1 U8838 ( .A1(n8964), .A2(n8965), .ZN(n8416) );
  AND2_X1 U8839 ( .A1(n8966), .A2(n8967), .ZN(n8965) );
  AND2_X1 U8840 ( .A1(n8387), .A2(n8393), .ZN(n8964) );
  OR2_X1 U8841 ( .A1(n8968), .A2(n8969), .ZN(n8387) );
  AND2_X1 U8842 ( .A1(n8970), .A2(n8971), .ZN(n8969) );
  AND2_X1 U8843 ( .A1(n8354), .A2(n8360), .ZN(n8968) );
  OR2_X1 U8844 ( .A1(n8972), .A2(n8973), .ZN(n8354) );
  AND2_X1 U8845 ( .A1(n8974), .A2(n8336), .ZN(n8973) );
  AND2_X1 U8846 ( .A1(n8326), .A2(n8975), .ZN(n8972) );
  OR2_X1 U8847 ( .A1(n8976), .A2(n8977), .ZN(n8326) );
  AND2_X1 U8848 ( .A1(n8978), .A2(n8308), .ZN(n8977) );
  AND2_X1 U8849 ( .A1(n8298), .A2(n8979), .ZN(n8976) );
  OR2_X1 U8850 ( .A1(n8980), .A2(n8981), .ZN(n8298) );
  AND2_X1 U8851 ( .A1(n8982), .A2(n8280), .ZN(n8981) );
  AND2_X1 U8852 ( .A1(n8270), .A2(n8983), .ZN(n8980) );
  OR2_X1 U8853 ( .A1(n8984), .A2(n8985), .ZN(n8270) );
  AND2_X1 U8854 ( .A1(n8986), .A2(n8252), .ZN(n8985) );
  AND2_X1 U8855 ( .A1(n8242), .A2(n8987), .ZN(n8984) );
  OR2_X1 U8856 ( .A1(n8988), .A2(n8989), .ZN(n8242) );
  AND2_X1 U8857 ( .A1(n8990), .A2(n8224), .ZN(n8989) );
  AND2_X1 U8858 ( .A1(n8214), .A2(n8991), .ZN(n8988) );
  OR2_X1 U8859 ( .A1(n8992), .A2(n8993), .ZN(n8214) );
  AND2_X1 U8860 ( .A1(n8994), .A2(n8196), .ZN(n8993) );
  AND2_X1 U8861 ( .A1(n8186), .A2(n8995), .ZN(n8992) );
  OR2_X1 U8862 ( .A1(n8996), .A2(n8997), .ZN(n8186) );
  AND2_X1 U8863 ( .A1(n8998), .A2(n8168), .ZN(n8997) );
  AND2_X1 U8864 ( .A1(n8158), .A2(n8999), .ZN(n8996) );
  OR2_X1 U8865 ( .A1(n9000), .A2(n9001), .ZN(n8158) );
  AND2_X1 U8866 ( .A1(n9002), .A2(n8140), .ZN(n9001) );
  AND2_X1 U8867 ( .A1(n8130), .A2(n9003), .ZN(n9000) );
  OR2_X1 U8868 ( .A1(n9004), .A2(n9005), .ZN(n8130) );
  AND2_X1 U8869 ( .A1(n9006), .A2(n8112), .ZN(n9005) );
  AND2_X1 U8870 ( .A1(n8102), .A2(n9007), .ZN(n9004) );
  OR2_X1 U8871 ( .A1(n9008), .A2(n9009), .ZN(n8102) );
  AND2_X1 U8872 ( .A1(n9010), .A2(n8075), .ZN(n9009) );
  AND2_X1 U8873 ( .A1(n8065), .A2(n9011), .ZN(n9008) );
  OR2_X1 U8874 ( .A1(n9012), .A2(n9013), .ZN(n8065) );
  AND2_X1 U8875 ( .A1(n9014), .A2(n8047), .ZN(n9013) );
  AND2_X1 U8876 ( .A1(n8037), .A2(n9015), .ZN(n9012) );
  AND2_X1 U8877 ( .A1(n9016), .A2(n9017), .ZN(n8037) );
  OR2_X1 U8878 ( .A1(n7998), .A2(n9018), .ZN(n9017) );
  AND2_X1 U8879 ( .A1(n8002), .A2(n8018), .ZN(n9018) );
  INV_X1 U8880 ( .A(n7984), .ZN(n8018) );
  AND2_X1 U8881 ( .A1(a_31_), .A2(b_31_), .ZN(n7984) );
  AND2_X1 U8882 ( .A1(n7989), .A2(n9019), .ZN(n8893) );
  INV_X1 U8883 ( .A(n8882), .ZN(n8891) );
  OR2_X1 U8884 ( .A1(n9020), .A2(n9021), .ZN(n8882) );
  AND2_X1 U8885 ( .A1(n9022), .A2(n7956), .ZN(n8877) );
  XNOR2_X1 U8886 ( .A(n9023), .B(n9024), .ZN(n9022) );
  XOR2_X1 U8887 ( .A(n9025), .B(n9026), .Z(n9024) );
  OR2_X1 U8888 ( .A1(n9027), .A2(n7955), .ZN(Result_31_) );
  AND2_X1 U8889 ( .A1(n7956), .A2(n9028), .ZN(n9027) );
  XNOR2_X1 U8890 ( .A(n9029), .B(n9030), .ZN(n9028) );
  OR2_X1 U8891 ( .A1(n9031), .A2(n7955), .ZN(Result_30_) );
  AND2_X1 U8892 ( .A1(n9032), .A2(n9033), .ZN(n9031) );
  OR2_X1 U8893 ( .A1(n9034), .A2(n9035), .ZN(n9033) );
  AND2_X1 U8894 ( .A1(n9036), .A2(n9030), .ZN(n9034) );
  OR2_X1 U8895 ( .A1(n9037), .A2(n7955), .ZN(Result_2_) );
  AND2_X1 U8896 ( .A1(n9038), .A2(n7956), .ZN(n9037) );
  XOR2_X1 U8897 ( .A(n9039), .B(n9040), .Z(n9038) );
  OR2_X1 U8898 ( .A1(n7955), .A2(n9041), .ZN(Result_29_) );
  OR2_X1 U8899 ( .A1(n9042), .A2(n9043), .ZN(n9041) );
  AND2_X1 U8900 ( .A1(n9044), .A2(n9032), .ZN(n9043) );
  AND2_X1 U8901 ( .A1(n9045), .A2(n7956), .ZN(n9032) );
  INV_X1 U8902 ( .A(n9046), .ZN(n9045) );
  INV_X1 U8903 ( .A(n9047), .ZN(n9044) );
  AND2_X1 U8904 ( .A1(n9048), .A2(n9047), .ZN(n9042) );
  OR2_X1 U8905 ( .A1(n9049), .A2(n9050), .ZN(n9047) );
  AND2_X1 U8906 ( .A1(n7956), .A2(n9046), .ZN(n9048) );
  OR2_X1 U8907 ( .A1(n9051), .A2(n7955), .ZN(Result_28_) );
  AND2_X1 U8908 ( .A1(n9052), .A2(n7956), .ZN(n9051) );
  XOR2_X1 U8909 ( .A(n9053), .B(n9054), .Z(n9052) );
  AND2_X1 U8910 ( .A1(n9055), .A2(n9056), .ZN(n9054) );
  OR2_X1 U8911 ( .A1(n9057), .A2(n7955), .ZN(Result_27_) );
  AND2_X1 U8912 ( .A1(n9058), .A2(n7956), .ZN(n9057) );
  XOR2_X1 U8913 ( .A(n9059), .B(n9060), .Z(n9058) );
  AND2_X1 U8914 ( .A1(n9061), .A2(n9062), .ZN(n9060) );
  INV_X1 U8915 ( .A(n9063), .ZN(n9062) );
  OR2_X1 U8916 ( .A1(n9064), .A2(n7955), .ZN(Result_26_) );
  AND2_X1 U8917 ( .A1(n9065), .A2(n7956), .ZN(n9064) );
  XOR2_X1 U8918 ( .A(n9066), .B(n9067), .Z(n9065) );
  AND2_X1 U8919 ( .A1(n9068), .A2(n9069), .ZN(n9067) );
  INV_X1 U8920 ( .A(n9070), .ZN(n9069) );
  OR2_X1 U8921 ( .A1(n9071), .A2(n7955), .ZN(Result_25_) );
  AND2_X1 U8922 ( .A1(n9072), .A2(n7956), .ZN(n9071) );
  XOR2_X1 U8923 ( .A(n9073), .B(n9074), .Z(n9072) );
  AND2_X1 U8924 ( .A1(n9075), .A2(n9076), .ZN(n9074) );
  OR2_X1 U8925 ( .A1(n9077), .A2(n7955), .ZN(Result_24_) );
  AND2_X1 U8926 ( .A1(n9078), .A2(n7956), .ZN(n9077) );
  XOR2_X1 U8927 ( .A(n9079), .B(n9080), .Z(n9078) );
  AND2_X1 U8928 ( .A1(n9081), .A2(n9082), .ZN(n9080) );
  INV_X1 U8929 ( .A(n9083), .ZN(n9081) );
  OR2_X1 U8930 ( .A1(n9084), .A2(n7955), .ZN(Result_23_) );
  AND2_X1 U8931 ( .A1(n9085), .A2(n7956), .ZN(n9084) );
  XOR2_X1 U8932 ( .A(n9086), .B(n9087), .Z(n9085) );
  AND2_X1 U8933 ( .A1(n9088), .A2(n9089), .ZN(n9087) );
  INV_X1 U8934 ( .A(n9090), .ZN(n9089) );
  OR2_X1 U8935 ( .A1(n9091), .A2(n7955), .ZN(Result_22_) );
  AND2_X1 U8936 ( .A1(n9092), .A2(n7956), .ZN(n9091) );
  XOR2_X1 U8937 ( .A(n9093), .B(n9094), .Z(n9092) );
  AND2_X1 U8938 ( .A1(n9095), .A2(n9096), .ZN(n9094) );
  OR2_X1 U8939 ( .A1(n9097), .A2(n9098), .ZN(n9095) );
  INV_X1 U8940 ( .A(n9099), .ZN(n9097) );
  OR2_X1 U8941 ( .A1(n9100), .A2(n7955), .ZN(Result_21_) );
  AND2_X1 U8942 ( .A1(n9101), .A2(n7956), .ZN(n9100) );
  XOR2_X1 U8943 ( .A(n9102), .B(n9103), .Z(n9101) );
  AND2_X1 U8944 ( .A1(n9104), .A2(n9105), .ZN(n9103) );
  INV_X1 U8945 ( .A(n9106), .ZN(n9105) );
  OR2_X1 U8946 ( .A1(n9107), .A2(n7955), .ZN(Result_20_) );
  AND2_X1 U8947 ( .A1(n9108), .A2(n7956), .ZN(n9107) );
  XOR2_X1 U8948 ( .A(n9109), .B(n9110), .Z(n9108) );
  AND2_X1 U8949 ( .A1(n9111), .A2(n9112), .ZN(n9110) );
  OR2_X1 U8950 ( .A1(n9113), .A2(n7955), .ZN(Result_1_) );
  AND2_X1 U8951 ( .A1(n7956), .A2(n9114), .ZN(n9113) );
  XOR2_X1 U8952 ( .A(n9115), .B(n9116), .Z(n9114) );
  AND2_X1 U8953 ( .A1(n9117), .A2(n9118), .ZN(n9116) );
  OR2_X1 U8954 ( .A1(n9119), .A2(n9120), .ZN(n9118) );
  AND2_X1 U8955 ( .A1(n9121), .A2(n9122), .ZN(n9119) );
  INV_X1 U8956 ( .A(n9123), .ZN(n9117) );
  OR2_X1 U8957 ( .A1(n9124), .A2(n7955), .ZN(Result_19_) );
  AND2_X1 U8958 ( .A1(n9125), .A2(n7956), .ZN(n9124) );
  XOR2_X1 U8959 ( .A(n9126), .B(n9127), .Z(n9125) );
  AND2_X1 U8960 ( .A1(n9128), .A2(n9129), .ZN(n9127) );
  INV_X1 U8961 ( .A(n9130), .ZN(n9129) );
  OR2_X1 U8962 ( .A1(n9131), .A2(n7955), .ZN(Result_18_) );
  AND2_X1 U8963 ( .A1(n9132), .A2(n7956), .ZN(n9131) );
  XOR2_X1 U8964 ( .A(n9133), .B(n9134), .Z(n9132) );
  AND2_X1 U8965 ( .A1(n9135), .A2(n9136), .ZN(n9134) );
  OR2_X1 U8966 ( .A1(n9137), .A2(n9138), .ZN(n9135) );
  INV_X1 U8967 ( .A(n9139), .ZN(n9137) );
  OR2_X1 U8968 ( .A1(n9140), .A2(n7955), .ZN(Result_17_) );
  AND2_X1 U8969 ( .A1(n9141), .A2(n7956), .ZN(n9140) );
  XOR2_X1 U8970 ( .A(n9142), .B(n9143), .Z(n9141) );
  AND2_X1 U8971 ( .A1(n9144), .A2(n9145), .ZN(n9143) );
  INV_X1 U8972 ( .A(n9146), .ZN(n9145) );
  OR2_X1 U8973 ( .A1(n9147), .A2(n7955), .ZN(Result_16_) );
  AND2_X1 U8974 ( .A1(n9148), .A2(n7956), .ZN(n9147) );
  XOR2_X1 U8975 ( .A(n9149), .B(n9150), .Z(n9148) );
  AND2_X1 U8976 ( .A1(n9151), .A2(n9152), .ZN(n9150) );
  INV_X1 U8977 ( .A(n9153), .ZN(n9151) );
  OR2_X1 U8978 ( .A1(n9154), .A2(n7955), .ZN(Result_15_) );
  AND2_X1 U8979 ( .A1(n9155), .A2(n7956), .ZN(n9154) );
  XOR2_X1 U8980 ( .A(n9156), .B(n9157), .Z(n9155) );
  AND2_X1 U8981 ( .A1(n9158), .A2(n9159), .ZN(n9157) );
  OR2_X1 U8982 ( .A1(n9160), .A2(n7955), .ZN(Result_14_) );
  AND2_X1 U8983 ( .A1(n9161), .A2(n7956), .ZN(n9160) );
  XOR2_X1 U8984 ( .A(n9162), .B(n9163), .Z(n9161) );
  AND2_X1 U8985 ( .A1(n9164), .A2(n9165), .ZN(n9163) );
  INV_X1 U8986 ( .A(n9166), .ZN(n9165) );
  OR2_X1 U8987 ( .A1(n9167), .A2(n9168), .ZN(n9164) );
  AND2_X1 U8988 ( .A1(n9169), .A2(n9170), .ZN(n9167) );
  OR2_X1 U8989 ( .A1(n9171), .A2(n7955), .ZN(Result_13_) );
  AND2_X1 U8990 ( .A1(n9172), .A2(n7956), .ZN(n9171) );
  XOR2_X1 U8991 ( .A(n9173), .B(n9174), .Z(n9172) );
  AND2_X1 U8992 ( .A1(n9175), .A2(n9176), .ZN(n9174) );
  OR2_X1 U8993 ( .A1(n9177), .A2(n9178), .ZN(n9176) );
  INV_X1 U8994 ( .A(n9179), .ZN(n9175) );
  OR2_X1 U8995 ( .A1(n9180), .A2(n7955), .ZN(Result_12_) );
  AND2_X1 U8996 ( .A1(n9181), .A2(n7956), .ZN(n9180) );
  XOR2_X1 U8997 ( .A(n9182), .B(n9183), .Z(n9181) );
  OR2_X1 U8998 ( .A1(n9184), .A2(n7955), .ZN(Result_11_) );
  AND2_X1 U8999 ( .A1(n7956), .A2(n9185), .ZN(n9184) );
  XOR2_X1 U9000 ( .A(n9186), .B(n9187), .Z(n9185) );
  AND2_X1 U9001 ( .A1(n9188), .A2(n9189), .ZN(n9187) );
  OR2_X1 U9002 ( .A1(n9190), .A2(n9191), .ZN(n9189) );
  INV_X1 U9003 ( .A(n9192), .ZN(n9188) );
  OR2_X1 U9004 ( .A1(n9193), .A2(n7955), .ZN(Result_10_) );
  AND2_X1 U9005 ( .A1(n9194), .A2(n7956), .ZN(n9193) );
  XOR2_X1 U9006 ( .A(n9195), .B(n9196), .Z(n9194) );
  OR2_X1 U9007 ( .A1(n9197), .A2(n7955), .ZN(Result_0_) );
  OR2_X1 U9008 ( .A1(n9198), .A2(n9199), .ZN(n7955) );
  AND2_X1 U9009 ( .A1(n7989), .A2(n9200), .ZN(n9199) );
  INV_X1 U9010 ( .A(n9201), .ZN(n9200) );
  AND2_X1 U9011 ( .A1(n9202), .A2(n9203), .ZN(n9201) );
  OR2_X1 U9012 ( .A1(n8890), .A2(n9021), .ZN(n9202) );
  INV_X1 U9013 ( .A(n9019), .ZN(n8890) );
  OR2_X1 U9014 ( .A1(n9204), .A2(n9205), .ZN(n9019) );
  AND2_X1 U9015 ( .A1(n8862), .A2(n8902), .ZN(n9205) );
  AND2_X1 U9016 ( .A1(b_1_), .A2(n9206), .ZN(n9204) );
  OR2_X1 U9017 ( .A1(n8902), .A2(n8862), .ZN(n9206) );
  OR2_X1 U9018 ( .A1(n9207), .A2(n9208), .ZN(n8862) );
  AND2_X1 U9019 ( .A1(n8833), .A2(n8906), .ZN(n9208) );
  AND2_X1 U9020 ( .A1(b_2_), .A2(n9209), .ZN(n9207) );
  OR2_X1 U9021 ( .A1(n8906), .A2(n8833), .ZN(n9209) );
  OR2_X1 U9022 ( .A1(n9210), .A2(n9211), .ZN(n8833) );
  AND2_X1 U9023 ( .A1(n8804), .A2(n8910), .ZN(n9211) );
  AND2_X1 U9024 ( .A1(b_3_), .A2(n9212), .ZN(n9210) );
  OR2_X1 U9025 ( .A1(n8910), .A2(n8804), .ZN(n9212) );
  OR2_X1 U9026 ( .A1(n9213), .A2(n9214), .ZN(n8804) );
  AND2_X1 U9027 ( .A1(n8775), .A2(n8914), .ZN(n9214) );
  AND2_X1 U9028 ( .A1(b_4_), .A2(n9215), .ZN(n9213) );
  OR2_X1 U9029 ( .A1(n8914), .A2(n8775), .ZN(n9215) );
  OR2_X1 U9030 ( .A1(n9216), .A2(n9217), .ZN(n8775) );
  AND2_X1 U9031 ( .A1(n8746), .A2(n8918), .ZN(n9217) );
  AND2_X1 U9032 ( .A1(b_5_), .A2(n9218), .ZN(n9216) );
  OR2_X1 U9033 ( .A1(n8918), .A2(n8746), .ZN(n9218) );
  OR2_X1 U9034 ( .A1(n9219), .A2(n9220), .ZN(n8746) );
  AND2_X1 U9035 ( .A1(n8717), .A2(n8922), .ZN(n9220) );
  AND2_X1 U9036 ( .A1(b_6_), .A2(n9221), .ZN(n9219) );
  OR2_X1 U9037 ( .A1(n8922), .A2(n8717), .ZN(n9221) );
  OR2_X1 U9038 ( .A1(n9222), .A2(n9223), .ZN(n8717) );
  AND2_X1 U9039 ( .A1(n8688), .A2(n8926), .ZN(n9223) );
  AND2_X1 U9040 ( .A1(b_7_), .A2(n9224), .ZN(n9222) );
  OR2_X1 U9041 ( .A1(n8926), .A2(n8688), .ZN(n9224) );
  OR2_X1 U9042 ( .A1(n9225), .A2(n9226), .ZN(n8688) );
  AND2_X1 U9043 ( .A1(n8650), .A2(n8930), .ZN(n9226) );
  AND2_X1 U9044 ( .A1(b_8_), .A2(n9227), .ZN(n9225) );
  OR2_X1 U9045 ( .A1(n8930), .A2(n8650), .ZN(n9227) );
  OR2_X1 U9046 ( .A1(n9228), .A2(n9229), .ZN(n8650) );
  AND2_X1 U9047 ( .A1(n8621), .A2(n8934), .ZN(n9229) );
  AND2_X1 U9048 ( .A1(b_9_), .A2(n9230), .ZN(n9228) );
  OR2_X1 U9049 ( .A1(n8934), .A2(n8621), .ZN(n9230) );
  OR2_X1 U9050 ( .A1(n9231), .A2(n9232), .ZN(n8621) );
  AND2_X1 U9051 ( .A1(n8592), .A2(n8938), .ZN(n9232) );
  AND2_X1 U9052 ( .A1(b_10_), .A2(n9233), .ZN(n9231) );
  OR2_X1 U9053 ( .A1(n8938), .A2(n8592), .ZN(n9233) );
  OR2_X1 U9054 ( .A1(n9234), .A2(n9235), .ZN(n8592) );
  AND2_X1 U9055 ( .A1(n8563), .A2(n8942), .ZN(n9235) );
  AND2_X1 U9056 ( .A1(b_11_), .A2(n9236), .ZN(n9234) );
  OR2_X1 U9057 ( .A1(n8942), .A2(n8563), .ZN(n9236) );
  OR2_X1 U9058 ( .A1(n9237), .A2(n9238), .ZN(n8563) );
  AND2_X1 U9059 ( .A1(n8534), .A2(n8946), .ZN(n9238) );
  AND2_X1 U9060 ( .A1(b_12_), .A2(n9239), .ZN(n9237) );
  OR2_X1 U9061 ( .A1(n8946), .A2(n8534), .ZN(n9239) );
  OR2_X1 U9062 ( .A1(n9240), .A2(n9241), .ZN(n8534) );
  AND2_X1 U9063 ( .A1(n8505), .A2(n8950), .ZN(n9241) );
  AND2_X1 U9064 ( .A1(b_13_), .A2(n9242), .ZN(n9240) );
  OR2_X1 U9065 ( .A1(n8950), .A2(n8505), .ZN(n9242) );
  OR2_X1 U9066 ( .A1(n9243), .A2(n9244), .ZN(n8505) );
  AND2_X1 U9067 ( .A1(n8476), .A2(n8954), .ZN(n9244) );
  AND2_X1 U9068 ( .A1(b_14_), .A2(n9245), .ZN(n9243) );
  OR2_X1 U9069 ( .A1(n8954), .A2(n8476), .ZN(n9245) );
  OR2_X1 U9070 ( .A1(n9246), .A2(n9247), .ZN(n8476) );
  AND2_X1 U9071 ( .A1(n8447), .A2(n8958), .ZN(n9247) );
  AND2_X1 U9072 ( .A1(b_15_), .A2(n9248), .ZN(n9246) );
  OR2_X1 U9073 ( .A1(n8958), .A2(n8447), .ZN(n9248) );
  OR2_X1 U9074 ( .A1(n9249), .A2(n9250), .ZN(n8447) );
  AND2_X1 U9075 ( .A1(n8418), .A2(n8962), .ZN(n9250) );
  AND2_X1 U9076 ( .A1(b_16_), .A2(n9251), .ZN(n9249) );
  OR2_X1 U9077 ( .A1(n8962), .A2(n8418), .ZN(n9251) );
  OR2_X1 U9078 ( .A1(n9252), .A2(n9253), .ZN(n8418) );
  AND2_X1 U9079 ( .A1(n8389), .A2(n8966), .ZN(n9253) );
  AND2_X1 U9080 ( .A1(b_17_), .A2(n9254), .ZN(n9252) );
  OR2_X1 U9081 ( .A1(n8966), .A2(n8389), .ZN(n9254) );
  OR2_X1 U9082 ( .A1(n9255), .A2(n9256), .ZN(n8389) );
  AND2_X1 U9083 ( .A1(n8356), .A2(n8970), .ZN(n9256) );
  AND2_X1 U9084 ( .A1(b_18_), .A2(n9257), .ZN(n9255) );
  OR2_X1 U9085 ( .A1(n8970), .A2(n8356), .ZN(n9257) );
  OR2_X1 U9086 ( .A1(n9258), .A2(n9259), .ZN(n8356) );
  AND2_X1 U9087 ( .A1(n8327), .A2(n8974), .ZN(n9259) );
  AND2_X1 U9088 ( .A1(b_19_), .A2(n9260), .ZN(n9258) );
  OR2_X1 U9089 ( .A1(n8974), .A2(n8327), .ZN(n9260) );
  OR2_X1 U9090 ( .A1(n9261), .A2(n9262), .ZN(n8327) );
  AND2_X1 U9091 ( .A1(n8299), .A2(n8978), .ZN(n9262) );
  AND2_X1 U9092 ( .A1(b_20_), .A2(n9263), .ZN(n9261) );
  OR2_X1 U9093 ( .A1(n8978), .A2(n8299), .ZN(n9263) );
  OR2_X1 U9094 ( .A1(n9264), .A2(n9265), .ZN(n8299) );
  AND2_X1 U9095 ( .A1(n8271), .A2(n8982), .ZN(n9265) );
  AND2_X1 U9096 ( .A1(b_21_), .A2(n9266), .ZN(n9264) );
  OR2_X1 U9097 ( .A1(n8982), .A2(n8271), .ZN(n9266) );
  OR2_X1 U9098 ( .A1(n9267), .A2(n9268), .ZN(n8271) );
  AND2_X1 U9099 ( .A1(n8243), .A2(n8986), .ZN(n9268) );
  AND2_X1 U9100 ( .A1(b_22_), .A2(n9269), .ZN(n9267) );
  OR2_X1 U9101 ( .A1(n8986), .A2(n8243), .ZN(n9269) );
  OR2_X1 U9102 ( .A1(n9270), .A2(n9271), .ZN(n8243) );
  AND2_X1 U9103 ( .A1(n8215), .A2(n8990), .ZN(n9271) );
  AND2_X1 U9104 ( .A1(b_23_), .A2(n9272), .ZN(n9270) );
  OR2_X1 U9105 ( .A1(n8990), .A2(n8215), .ZN(n9272) );
  OR2_X1 U9106 ( .A1(n9273), .A2(n9274), .ZN(n8215) );
  AND2_X1 U9107 ( .A1(n8187), .A2(n8994), .ZN(n9274) );
  AND2_X1 U9108 ( .A1(b_24_), .A2(n9275), .ZN(n9273) );
  OR2_X1 U9109 ( .A1(n8994), .A2(n8187), .ZN(n9275) );
  OR2_X1 U9110 ( .A1(n9276), .A2(n9277), .ZN(n8187) );
  AND2_X1 U9111 ( .A1(n8159), .A2(n8998), .ZN(n9277) );
  AND2_X1 U9112 ( .A1(b_25_), .A2(n9278), .ZN(n9276) );
  OR2_X1 U9113 ( .A1(n8998), .A2(n8159), .ZN(n9278) );
  OR2_X1 U9114 ( .A1(n9279), .A2(n9280), .ZN(n8159) );
  AND2_X1 U9115 ( .A1(n8131), .A2(n9002), .ZN(n9280) );
  AND2_X1 U9116 ( .A1(b_26_), .A2(n9281), .ZN(n9279) );
  OR2_X1 U9117 ( .A1(n9002), .A2(n8131), .ZN(n9281) );
  OR2_X1 U9118 ( .A1(n9282), .A2(n9283), .ZN(n8131) );
  AND2_X1 U9119 ( .A1(n8103), .A2(n9006), .ZN(n9283) );
  AND2_X1 U9120 ( .A1(b_27_), .A2(n9284), .ZN(n9282) );
  OR2_X1 U9121 ( .A1(n9006), .A2(n8103), .ZN(n9284) );
  OR2_X1 U9122 ( .A1(n9285), .A2(n9286), .ZN(n8103) );
  AND2_X1 U9123 ( .A1(n8066), .A2(n9010), .ZN(n9286) );
  AND2_X1 U9124 ( .A1(b_28_), .A2(n9287), .ZN(n9285) );
  OR2_X1 U9125 ( .A1(n9010), .A2(n8066), .ZN(n9287) );
  OR2_X1 U9126 ( .A1(n9288), .A2(n9289), .ZN(n8066) );
  AND2_X1 U9127 ( .A1(n8038), .A2(n9014), .ZN(n9289) );
  AND2_X1 U9128 ( .A1(b_29_), .A2(n9290), .ZN(n9288) );
  OR2_X1 U9129 ( .A1(n9014), .A2(n8038), .ZN(n9290) );
  OR2_X1 U9130 ( .A1(n9291), .A2(n9292), .ZN(n8038) );
  AND2_X1 U9131 ( .A1(n7992), .A2(n8002), .ZN(n9292) );
  AND2_X1 U9132 ( .A1(b_30_), .A2(n9293), .ZN(n9291) );
  OR2_X1 U9133 ( .A1(n7992), .A2(n8002), .ZN(n9293) );
  AND2_X1 U9134 ( .A1(n9294), .A2(b_31_), .ZN(n7992) );
  INV_X1 U9135 ( .A(operation_0_), .ZN(n8899) );
  AND2_X1 U9136 ( .A1(n9295), .A2(n7990), .ZN(n9198) );
  INV_X1 U9137 ( .A(operation_1_), .ZN(n8898) );
  AND2_X1 U9138 ( .A1(n9296), .A2(n9203), .ZN(n9295) );
  INV_X1 U9139 ( .A(n9020), .ZN(n9203) );
  AND2_X1 U9140 ( .A1(n9297), .A2(b_0_), .ZN(n9020) );
  OR2_X1 U9141 ( .A1(n9021), .A2(n8888), .ZN(n9296) );
  OR2_X1 U9142 ( .A1(n9298), .A2(n9299), .ZN(n8888) );
  AND2_X1 U9143 ( .A1(a_1_), .A2(n8859), .ZN(n9299) );
  AND2_X1 U9144 ( .A1(n9300), .A2(n8903), .ZN(n9298) );
  OR2_X1 U9145 ( .A1(a_1_), .A2(n8859), .ZN(n9300) );
  OR2_X1 U9146 ( .A1(n9301), .A2(n9302), .ZN(n8859) );
  AND2_X1 U9147 ( .A1(a_2_), .A2(n8830), .ZN(n9302) );
  AND2_X1 U9148 ( .A1(n9303), .A2(n8907), .ZN(n9301) );
  OR2_X1 U9149 ( .A1(a_2_), .A2(n8830), .ZN(n9303) );
  OR2_X1 U9150 ( .A1(n9304), .A2(n9305), .ZN(n8830) );
  AND2_X1 U9151 ( .A1(a_3_), .A2(n8801), .ZN(n9305) );
  AND2_X1 U9152 ( .A1(n9306), .A2(n8911), .ZN(n9304) );
  OR2_X1 U9153 ( .A1(a_3_), .A2(n8801), .ZN(n9306) );
  OR2_X1 U9154 ( .A1(n9307), .A2(n9308), .ZN(n8801) );
  AND2_X1 U9155 ( .A1(a_4_), .A2(n8772), .ZN(n9308) );
  AND2_X1 U9156 ( .A1(n9309), .A2(n8915), .ZN(n9307) );
  OR2_X1 U9157 ( .A1(a_4_), .A2(n8772), .ZN(n9309) );
  OR2_X1 U9158 ( .A1(n9310), .A2(n9311), .ZN(n8772) );
  AND2_X1 U9159 ( .A1(a_5_), .A2(n8743), .ZN(n9311) );
  AND2_X1 U9160 ( .A1(n9312), .A2(n8919), .ZN(n9310) );
  OR2_X1 U9161 ( .A1(a_5_), .A2(n8743), .ZN(n9312) );
  OR2_X1 U9162 ( .A1(n9313), .A2(n9314), .ZN(n8743) );
  AND2_X1 U9163 ( .A1(a_6_), .A2(n8714), .ZN(n9314) );
  AND2_X1 U9164 ( .A1(n9315), .A2(n8923), .ZN(n9313) );
  OR2_X1 U9165 ( .A1(a_6_), .A2(n8714), .ZN(n9315) );
  OR2_X1 U9166 ( .A1(n9316), .A2(n9317), .ZN(n8714) );
  AND2_X1 U9167 ( .A1(a_7_), .A2(n8685), .ZN(n9317) );
  AND2_X1 U9168 ( .A1(n9318), .A2(n8927), .ZN(n9316) );
  OR2_X1 U9169 ( .A1(a_7_), .A2(n8685), .ZN(n9318) );
  OR2_X1 U9170 ( .A1(n9319), .A2(n9320), .ZN(n8685) );
  AND2_X1 U9171 ( .A1(a_8_), .A2(n8647), .ZN(n9320) );
  AND2_X1 U9172 ( .A1(n9321), .A2(n8931), .ZN(n9319) );
  OR2_X1 U9173 ( .A1(a_8_), .A2(n8647), .ZN(n9321) );
  OR2_X1 U9174 ( .A1(n9322), .A2(n9323), .ZN(n8647) );
  AND2_X1 U9175 ( .A1(a_9_), .A2(n8618), .ZN(n9323) );
  AND2_X1 U9176 ( .A1(n9324), .A2(n8935), .ZN(n9322) );
  OR2_X1 U9177 ( .A1(a_9_), .A2(n8618), .ZN(n9324) );
  OR2_X1 U9178 ( .A1(n9325), .A2(n9326), .ZN(n8618) );
  AND2_X1 U9179 ( .A1(a_10_), .A2(n8589), .ZN(n9326) );
  AND2_X1 U9180 ( .A1(n9327), .A2(n8939), .ZN(n9325) );
  OR2_X1 U9181 ( .A1(a_10_), .A2(n8589), .ZN(n9327) );
  OR2_X1 U9182 ( .A1(n9328), .A2(n9329), .ZN(n8589) );
  AND2_X1 U9183 ( .A1(a_11_), .A2(n8560), .ZN(n9329) );
  AND2_X1 U9184 ( .A1(n9330), .A2(n8943), .ZN(n9328) );
  OR2_X1 U9185 ( .A1(a_11_), .A2(n8560), .ZN(n9330) );
  OR2_X1 U9186 ( .A1(n9331), .A2(n9332), .ZN(n8560) );
  AND2_X1 U9187 ( .A1(a_12_), .A2(n8531), .ZN(n9332) );
  AND2_X1 U9188 ( .A1(n9333), .A2(n8947), .ZN(n9331) );
  OR2_X1 U9189 ( .A1(a_12_), .A2(n8531), .ZN(n9333) );
  OR2_X1 U9190 ( .A1(n9334), .A2(n9335), .ZN(n8531) );
  AND2_X1 U9191 ( .A1(a_13_), .A2(n8502), .ZN(n9335) );
  AND2_X1 U9192 ( .A1(n9336), .A2(n8951), .ZN(n9334) );
  OR2_X1 U9193 ( .A1(a_13_), .A2(n8502), .ZN(n9336) );
  OR2_X1 U9194 ( .A1(n9337), .A2(n9338), .ZN(n8502) );
  AND2_X1 U9195 ( .A1(a_14_), .A2(n8473), .ZN(n9338) );
  AND2_X1 U9196 ( .A1(n9339), .A2(n8955), .ZN(n9337) );
  OR2_X1 U9197 ( .A1(a_14_), .A2(n8473), .ZN(n9339) );
  OR2_X1 U9198 ( .A1(n9340), .A2(n9341), .ZN(n8473) );
  AND2_X1 U9199 ( .A1(a_15_), .A2(n8444), .ZN(n9341) );
  AND2_X1 U9200 ( .A1(n9342), .A2(n8959), .ZN(n9340) );
  OR2_X1 U9201 ( .A1(a_15_), .A2(n8444), .ZN(n9342) );
  OR2_X1 U9202 ( .A1(n9343), .A2(n9344), .ZN(n8444) );
  AND2_X1 U9203 ( .A1(a_16_), .A2(n8415), .ZN(n9344) );
  AND2_X1 U9204 ( .A1(n9345), .A2(n8963), .ZN(n9343) );
  OR2_X1 U9205 ( .A1(a_16_), .A2(n8415), .ZN(n9345) );
  OR2_X1 U9206 ( .A1(n9346), .A2(n9347), .ZN(n8415) );
  AND2_X1 U9207 ( .A1(a_17_), .A2(n8386), .ZN(n9347) );
  AND2_X1 U9208 ( .A1(n9348), .A2(n8967), .ZN(n9346) );
  OR2_X1 U9209 ( .A1(a_17_), .A2(n8386), .ZN(n9348) );
  OR2_X1 U9210 ( .A1(n9349), .A2(n9350), .ZN(n8386) );
  AND2_X1 U9211 ( .A1(a_18_), .A2(n8353), .ZN(n9350) );
  AND2_X1 U9212 ( .A1(n9351), .A2(n8971), .ZN(n9349) );
  OR2_X1 U9213 ( .A1(a_18_), .A2(n8353), .ZN(n9351) );
  OR2_X1 U9214 ( .A1(n9352), .A2(n9353), .ZN(n8353) );
  AND2_X1 U9215 ( .A1(a_19_), .A2(n8324), .ZN(n9353) );
  AND2_X1 U9216 ( .A1(n9354), .A2(n8336), .ZN(n9352) );
  OR2_X1 U9217 ( .A1(a_19_), .A2(n8324), .ZN(n9354) );
  OR2_X1 U9218 ( .A1(n9355), .A2(n9356), .ZN(n8324) );
  AND2_X1 U9219 ( .A1(a_20_), .A2(n8296), .ZN(n9356) );
  AND2_X1 U9220 ( .A1(n9357), .A2(n8308), .ZN(n9355) );
  OR2_X1 U9221 ( .A1(a_20_), .A2(n8296), .ZN(n9357) );
  OR2_X1 U9222 ( .A1(n9358), .A2(n9359), .ZN(n8296) );
  AND2_X1 U9223 ( .A1(a_21_), .A2(n8268), .ZN(n9359) );
  AND2_X1 U9224 ( .A1(n9360), .A2(n8280), .ZN(n9358) );
  OR2_X1 U9225 ( .A1(a_21_), .A2(n8268), .ZN(n9360) );
  OR2_X1 U9226 ( .A1(n9361), .A2(n9362), .ZN(n8268) );
  AND2_X1 U9227 ( .A1(a_22_), .A2(n8240), .ZN(n9362) );
  AND2_X1 U9228 ( .A1(n9363), .A2(n8252), .ZN(n9361) );
  OR2_X1 U9229 ( .A1(a_22_), .A2(n8240), .ZN(n9363) );
  OR2_X1 U9230 ( .A1(n9364), .A2(n9365), .ZN(n8240) );
  AND2_X1 U9231 ( .A1(a_23_), .A2(n8212), .ZN(n9365) );
  AND2_X1 U9232 ( .A1(n9366), .A2(n8224), .ZN(n9364) );
  OR2_X1 U9233 ( .A1(a_23_), .A2(n8212), .ZN(n9366) );
  OR2_X1 U9234 ( .A1(n9367), .A2(n9368), .ZN(n8212) );
  AND2_X1 U9235 ( .A1(a_24_), .A2(n8184), .ZN(n9368) );
  AND2_X1 U9236 ( .A1(n9369), .A2(n8196), .ZN(n9367) );
  OR2_X1 U9237 ( .A1(a_24_), .A2(n8184), .ZN(n9369) );
  OR2_X1 U9238 ( .A1(n9370), .A2(n9371), .ZN(n8184) );
  AND2_X1 U9239 ( .A1(a_25_), .A2(n8156), .ZN(n9371) );
  AND2_X1 U9240 ( .A1(n9372), .A2(n8168), .ZN(n9370) );
  OR2_X1 U9241 ( .A1(a_25_), .A2(n8156), .ZN(n9372) );
  OR2_X1 U9242 ( .A1(n9373), .A2(n9374), .ZN(n8156) );
  AND2_X1 U9243 ( .A1(a_26_), .A2(n8128), .ZN(n9374) );
  AND2_X1 U9244 ( .A1(n9375), .A2(n8140), .ZN(n9373) );
  OR2_X1 U9245 ( .A1(a_26_), .A2(n8128), .ZN(n9375) );
  OR2_X1 U9246 ( .A1(n9376), .A2(n9377), .ZN(n8128) );
  AND2_X1 U9247 ( .A1(a_27_), .A2(n8100), .ZN(n9377) );
  AND2_X1 U9248 ( .A1(n9378), .A2(n8112), .ZN(n9376) );
  OR2_X1 U9249 ( .A1(a_27_), .A2(n8100), .ZN(n9378) );
  OR2_X1 U9250 ( .A1(n9379), .A2(n9380), .ZN(n8100) );
  AND2_X1 U9251 ( .A1(a_28_), .A2(n8063), .ZN(n9380) );
  AND2_X1 U9252 ( .A1(n9381), .A2(n8075), .ZN(n9379) );
  OR2_X1 U9253 ( .A1(a_28_), .A2(n8063), .ZN(n9381) );
  OR2_X1 U9254 ( .A1(n9382), .A2(n9383), .ZN(n8063) );
  AND2_X1 U9255 ( .A1(a_29_), .A2(n8035), .ZN(n9383) );
  AND2_X1 U9256 ( .A1(n9384), .A2(n8047), .ZN(n9382) );
  OR2_X1 U9257 ( .A1(a_29_), .A2(n8035), .ZN(n9384) );
  OR2_X1 U9258 ( .A1(n9385), .A2(n9386), .ZN(n8035) );
  AND2_X1 U9259 ( .A1(a_30_), .A2(n7991), .ZN(n9386) );
  AND2_X1 U9260 ( .A1(n9387), .A2(n7998), .ZN(n9385) );
  OR2_X1 U9261 ( .A1(n7991), .A2(a_30_), .ZN(n9387) );
  AND2_X1 U9262 ( .A1(n9388), .A2(a_31_), .ZN(n7991) );
  AND2_X1 U9263 ( .A1(n9389), .A2(a_0_), .ZN(n9021) );
  AND2_X1 U9264 ( .A1(n7956), .A2(n9390), .ZN(n9197) );
  OR2_X1 U9265 ( .A1(n9391), .A2(n9392), .ZN(n9390) );
  OR2_X1 U9266 ( .A1(n9123), .A2(n9393), .ZN(n9392) );
  AND2_X1 U9267 ( .A1(n9115), .A2(n9120), .ZN(n9393) );
  AND2_X1 U9268 ( .A1(n9039), .A2(n9040), .ZN(n9115) );
  XNOR2_X1 U9269 ( .A(n9122), .B(n9394), .ZN(n9040) );
  OR2_X1 U9270 ( .A1(n9395), .A2(n9396), .ZN(n9039) );
  OR2_X1 U9271 ( .A1(n9397), .A2(n8673), .ZN(n9395) );
  AND2_X1 U9272 ( .A1(n8671), .A2(n8672), .ZN(n8673) );
  AND2_X1 U9273 ( .A1(n9398), .A2(n9399), .ZN(n8672) );
  INV_X1 U9274 ( .A(n9400), .ZN(n9398) );
  AND2_X1 U9275 ( .A1(n8667), .A2(n8671), .ZN(n9397) );
  INV_X1 U9276 ( .A(n9401), .ZN(n8671) );
  OR2_X1 U9277 ( .A1(n9402), .A2(n9396), .ZN(n9401) );
  INV_X1 U9278 ( .A(n9403), .ZN(n9396) );
  OR2_X1 U9279 ( .A1(n9404), .A2(n9405), .ZN(n9403) );
  AND2_X1 U9280 ( .A1(n9404), .A2(n9405), .ZN(n9402) );
  OR2_X1 U9281 ( .A1(n9406), .A2(n9407), .ZN(n9405) );
  AND2_X1 U9282 ( .A1(n9408), .A2(n9409), .ZN(n9407) );
  AND2_X1 U9283 ( .A1(n9410), .A2(n9411), .ZN(n9406) );
  OR2_X1 U9284 ( .A1(n9409), .A2(n9408), .ZN(n9411) );
  XOR2_X1 U9285 ( .A(n9412), .B(n9413), .Z(n9404) );
  XOR2_X1 U9286 ( .A(n9414), .B(n9415), .Z(n9413) );
  AND2_X1 U9287 ( .A1(n8373), .A2(n8374), .ZN(n8667) );
  XNOR2_X1 U9288 ( .A(n9399), .B(n9400), .ZN(n8374) );
  OR2_X1 U9289 ( .A1(n9416), .A2(n9417), .ZN(n9400) );
  AND2_X1 U9290 ( .A1(n9418), .A2(n9419), .ZN(n9417) );
  AND2_X1 U9291 ( .A1(n9420), .A2(n9421), .ZN(n9416) );
  OR2_X1 U9292 ( .A1(n9419), .A2(n9418), .ZN(n9421) );
  XNOR2_X1 U9293 ( .A(n9410), .B(n9422), .ZN(n9399) );
  XOR2_X1 U9294 ( .A(n9409), .B(n9408), .Z(n9422) );
  OR2_X1 U9295 ( .A1(n9297), .A2(n8911), .ZN(n9408) );
  OR2_X1 U9296 ( .A1(n9423), .A2(n9424), .ZN(n9409) );
  AND2_X1 U9297 ( .A1(n9425), .A2(n9426), .ZN(n9424) );
  AND2_X1 U9298 ( .A1(n9427), .A2(n9428), .ZN(n9423) );
  OR2_X1 U9299 ( .A1(n9426), .A2(n9425), .ZN(n9428) );
  XOR2_X1 U9300 ( .A(n9429), .B(n9430), .Z(n9410) );
  XOR2_X1 U9301 ( .A(n9431), .B(n9432), .Z(n9430) );
  OR2_X1 U9302 ( .A1(n9433), .A2(n9434), .ZN(n8373) );
  OR2_X1 U9303 ( .A1(n9435), .A2(n8089), .ZN(n9433) );
  AND2_X1 U9304 ( .A1(n8087), .A2(n8088), .ZN(n8089) );
  AND2_X1 U9305 ( .A1(n9436), .A2(n9437), .ZN(n8088) );
  INV_X1 U9306 ( .A(n9438), .ZN(n9436) );
  AND2_X1 U9307 ( .A1(n8083), .A2(n8087), .ZN(n9435) );
  INV_X1 U9308 ( .A(n9439), .ZN(n8087) );
  OR2_X1 U9309 ( .A1(n9440), .A2(n9434), .ZN(n9439) );
  INV_X1 U9310 ( .A(n9441), .ZN(n9434) );
  OR2_X1 U9311 ( .A1(n9442), .A2(n9443), .ZN(n9441) );
  AND2_X1 U9312 ( .A1(n9442), .A2(n9443), .ZN(n9440) );
  OR2_X1 U9313 ( .A1(n9444), .A2(n9445), .ZN(n9443) );
  AND2_X1 U9314 ( .A1(n9446), .A2(n9447), .ZN(n9445) );
  AND2_X1 U9315 ( .A1(n9448), .A2(n9449), .ZN(n9444) );
  OR2_X1 U9316 ( .A1(n9447), .A2(n9446), .ZN(n9449) );
  XOR2_X1 U9317 ( .A(n9420), .B(n9450), .Z(n9442) );
  XOR2_X1 U9318 ( .A(n9419), .B(n9418), .Z(n9450) );
  OR2_X1 U9319 ( .A1(n9297), .A2(n8915), .ZN(n9418) );
  OR2_X1 U9320 ( .A1(n9451), .A2(n9452), .ZN(n9419) );
  AND2_X1 U9321 ( .A1(n9453), .A2(n9454), .ZN(n9452) );
  AND2_X1 U9322 ( .A1(n9455), .A2(n9456), .ZN(n9451) );
  OR2_X1 U9323 ( .A1(n9454), .A2(n9453), .ZN(n9456) );
  XOR2_X1 U9324 ( .A(n9427), .B(n9457), .Z(n9420) );
  XOR2_X1 U9325 ( .A(n9426), .B(n9425), .Z(n9457) );
  OR2_X1 U9326 ( .A1(n8902), .A2(n8911), .ZN(n9425) );
  OR2_X1 U9327 ( .A1(n9458), .A2(n9459), .ZN(n9426) );
  AND2_X1 U9328 ( .A1(n9460), .A2(n9461), .ZN(n9459) );
  AND2_X1 U9329 ( .A1(n9462), .A2(n9463), .ZN(n9458) );
  OR2_X1 U9330 ( .A1(n9461), .A2(n9460), .ZN(n9463) );
  XOR2_X1 U9331 ( .A(n9464), .B(n9465), .Z(n9427) );
  XOR2_X1 U9332 ( .A(n9466), .B(n8837), .Z(n9465) );
  AND2_X1 U9333 ( .A1(n7980), .A2(n7981), .ZN(n8083) );
  XNOR2_X1 U9334 ( .A(n9437), .B(n9438), .ZN(n7981) );
  OR2_X1 U9335 ( .A1(n9467), .A2(n9468), .ZN(n9438) );
  AND2_X1 U9336 ( .A1(n9469), .A2(n9470), .ZN(n9468) );
  AND2_X1 U9337 ( .A1(n9471), .A2(n9472), .ZN(n9467) );
  OR2_X1 U9338 ( .A1(n9470), .A2(n9469), .ZN(n9472) );
  XNOR2_X1 U9339 ( .A(n9448), .B(n9473), .ZN(n9437) );
  XOR2_X1 U9340 ( .A(n9447), .B(n9446), .Z(n9473) );
  OR2_X1 U9341 ( .A1(n9297), .A2(n8919), .ZN(n9446) );
  OR2_X1 U9342 ( .A1(n9474), .A2(n9475), .ZN(n9447) );
  AND2_X1 U9343 ( .A1(n9476), .A2(n9477), .ZN(n9475) );
  AND2_X1 U9344 ( .A1(n9478), .A2(n9479), .ZN(n9474) );
  OR2_X1 U9345 ( .A1(n9477), .A2(n9476), .ZN(n9479) );
  XOR2_X1 U9346 ( .A(n9455), .B(n9480), .Z(n9448) );
  XOR2_X1 U9347 ( .A(n9454), .B(n9453), .Z(n9480) );
  OR2_X1 U9348 ( .A1(n8902), .A2(n8915), .ZN(n9453) );
  OR2_X1 U9349 ( .A1(n9481), .A2(n9482), .ZN(n9454) );
  AND2_X1 U9350 ( .A1(n9483), .A2(n9484), .ZN(n9482) );
  AND2_X1 U9351 ( .A1(n9485), .A2(n9486), .ZN(n9481) );
  OR2_X1 U9352 ( .A1(n9484), .A2(n9483), .ZN(n9486) );
  XOR2_X1 U9353 ( .A(n9462), .B(n9487), .Z(n9455) );
  XOR2_X1 U9354 ( .A(n9461), .B(n9460), .Z(n9487) );
  OR2_X1 U9355 ( .A1(n8906), .A2(n8911), .ZN(n9460) );
  OR2_X1 U9356 ( .A1(n9488), .A2(n9489), .ZN(n9461) );
  AND2_X1 U9357 ( .A1(n8808), .A2(n9490), .ZN(n9489) );
  AND2_X1 U9358 ( .A1(n9491), .A2(n9492), .ZN(n9488) );
  OR2_X1 U9359 ( .A1(n9490), .A2(n8808), .ZN(n9492) );
  XOR2_X1 U9360 ( .A(n9493), .B(n9494), .Z(n9462) );
  XOR2_X1 U9361 ( .A(n9495), .B(n9496), .Z(n9494) );
  OR2_X1 U9362 ( .A1(n9497), .A2(n9498), .ZN(n7980) );
  OR2_X1 U9363 ( .A1(n9499), .A2(n7977), .ZN(n9497) );
  AND2_X1 U9364 ( .A1(n7975), .A2(n7976), .ZN(n7977) );
  AND2_X1 U9365 ( .A1(n9500), .A2(n9501), .ZN(n7976) );
  INV_X1 U9366 ( .A(n9502), .ZN(n9500) );
  AND2_X1 U9367 ( .A1(n7971), .A2(n7975), .ZN(n9499) );
  INV_X1 U9368 ( .A(n9503), .ZN(n7975) );
  OR2_X1 U9369 ( .A1(n9504), .A2(n9498), .ZN(n9503) );
  INV_X1 U9370 ( .A(n9505), .ZN(n9498) );
  OR2_X1 U9371 ( .A1(n9506), .A2(n9507), .ZN(n9505) );
  AND2_X1 U9372 ( .A1(n9506), .A2(n9507), .ZN(n9504) );
  OR2_X1 U9373 ( .A1(n9508), .A2(n9509), .ZN(n9507) );
  AND2_X1 U9374 ( .A1(n9510), .A2(n9511), .ZN(n9509) );
  AND2_X1 U9375 ( .A1(n9512), .A2(n9513), .ZN(n9508) );
  OR2_X1 U9376 ( .A1(n9511), .A2(n9510), .ZN(n9513) );
  XOR2_X1 U9377 ( .A(n9471), .B(n9514), .Z(n9506) );
  XOR2_X1 U9378 ( .A(n9470), .B(n9469), .Z(n9514) );
  OR2_X1 U9379 ( .A1(n9297), .A2(n8923), .ZN(n9469) );
  OR2_X1 U9380 ( .A1(n9515), .A2(n9516), .ZN(n9470) );
  AND2_X1 U9381 ( .A1(n9517), .A2(n9518), .ZN(n9516) );
  AND2_X1 U9382 ( .A1(n9519), .A2(n9520), .ZN(n9515) );
  OR2_X1 U9383 ( .A1(n9518), .A2(n9517), .ZN(n9520) );
  XOR2_X1 U9384 ( .A(n9478), .B(n9521), .Z(n9471) );
  XOR2_X1 U9385 ( .A(n9477), .B(n9476), .Z(n9521) );
  OR2_X1 U9386 ( .A1(n8902), .A2(n8919), .ZN(n9476) );
  OR2_X1 U9387 ( .A1(n9522), .A2(n9523), .ZN(n9477) );
  AND2_X1 U9388 ( .A1(n9524), .A2(n9525), .ZN(n9523) );
  AND2_X1 U9389 ( .A1(n9526), .A2(n9527), .ZN(n9522) );
  OR2_X1 U9390 ( .A1(n9525), .A2(n9524), .ZN(n9527) );
  XOR2_X1 U9391 ( .A(n9485), .B(n9528), .Z(n9478) );
  XOR2_X1 U9392 ( .A(n9484), .B(n9483), .Z(n9528) );
  OR2_X1 U9393 ( .A1(n8906), .A2(n8915), .ZN(n9483) );
  OR2_X1 U9394 ( .A1(n9529), .A2(n9530), .ZN(n9484) );
  AND2_X1 U9395 ( .A1(n9531), .A2(n9532), .ZN(n9530) );
  AND2_X1 U9396 ( .A1(n9533), .A2(n9534), .ZN(n9529) );
  OR2_X1 U9397 ( .A1(n9532), .A2(n9531), .ZN(n9534) );
  XOR2_X1 U9398 ( .A(n9491), .B(n9535), .Z(n9485) );
  XOR2_X1 U9399 ( .A(n9490), .B(n8808), .Z(n9535) );
  OR2_X1 U9400 ( .A1(n8910), .A2(n8911), .ZN(n8808) );
  OR2_X1 U9401 ( .A1(n9536), .A2(n9537), .ZN(n9490) );
  AND2_X1 U9402 ( .A1(n9538), .A2(n9539), .ZN(n9537) );
  AND2_X1 U9403 ( .A1(n9540), .A2(n9541), .ZN(n9536) );
  OR2_X1 U9404 ( .A1(n9539), .A2(n9538), .ZN(n9541) );
  XOR2_X1 U9405 ( .A(n9542), .B(n9543), .Z(n9491) );
  XOR2_X1 U9406 ( .A(n9544), .B(n9545), .Z(n9543) );
  AND2_X1 U9407 ( .A1(n7967), .A2(n7968), .ZN(n7971) );
  XNOR2_X1 U9408 ( .A(n9501), .B(n9502), .ZN(n7968) );
  OR2_X1 U9409 ( .A1(n9546), .A2(n9547), .ZN(n9502) );
  AND2_X1 U9410 ( .A1(n9548), .A2(n9549), .ZN(n9547) );
  AND2_X1 U9411 ( .A1(n9550), .A2(n9551), .ZN(n9546) );
  OR2_X1 U9412 ( .A1(n9549), .A2(n9548), .ZN(n9551) );
  XNOR2_X1 U9413 ( .A(n9512), .B(n9552), .ZN(n9501) );
  XOR2_X1 U9414 ( .A(n9511), .B(n9510), .Z(n9552) );
  OR2_X1 U9415 ( .A1(n9297), .A2(n8927), .ZN(n9510) );
  OR2_X1 U9416 ( .A1(n9553), .A2(n9554), .ZN(n9511) );
  AND2_X1 U9417 ( .A1(n9555), .A2(n9556), .ZN(n9554) );
  AND2_X1 U9418 ( .A1(n9557), .A2(n9558), .ZN(n9553) );
  OR2_X1 U9419 ( .A1(n9556), .A2(n9555), .ZN(n9558) );
  XOR2_X1 U9420 ( .A(n9519), .B(n9559), .Z(n9512) );
  XOR2_X1 U9421 ( .A(n9518), .B(n9517), .Z(n9559) );
  OR2_X1 U9422 ( .A1(n8902), .A2(n8923), .ZN(n9517) );
  OR2_X1 U9423 ( .A1(n9560), .A2(n9561), .ZN(n9518) );
  AND2_X1 U9424 ( .A1(n9562), .A2(n9563), .ZN(n9561) );
  AND2_X1 U9425 ( .A1(n9564), .A2(n9565), .ZN(n9560) );
  OR2_X1 U9426 ( .A1(n9563), .A2(n9562), .ZN(n9565) );
  XOR2_X1 U9427 ( .A(n9526), .B(n9566), .Z(n9519) );
  XOR2_X1 U9428 ( .A(n9525), .B(n9524), .Z(n9566) );
  OR2_X1 U9429 ( .A1(n8906), .A2(n8919), .ZN(n9524) );
  OR2_X1 U9430 ( .A1(n9567), .A2(n9568), .ZN(n9525) );
  AND2_X1 U9431 ( .A1(n9569), .A2(n9570), .ZN(n9568) );
  AND2_X1 U9432 ( .A1(n9571), .A2(n9572), .ZN(n9567) );
  OR2_X1 U9433 ( .A1(n9570), .A2(n9569), .ZN(n9572) );
  XOR2_X1 U9434 ( .A(n9533), .B(n9573), .Z(n9526) );
  XOR2_X1 U9435 ( .A(n9532), .B(n9531), .Z(n9573) );
  OR2_X1 U9436 ( .A1(n8910), .A2(n8915), .ZN(n9531) );
  OR2_X1 U9437 ( .A1(n9574), .A2(n9575), .ZN(n9532) );
  AND2_X1 U9438 ( .A1(n8779), .A2(n9576), .ZN(n9575) );
  AND2_X1 U9439 ( .A1(n9577), .A2(n9578), .ZN(n9574) );
  OR2_X1 U9440 ( .A1(n9576), .A2(n8779), .ZN(n9578) );
  XOR2_X1 U9441 ( .A(n9540), .B(n9579), .Z(n9533) );
  XOR2_X1 U9442 ( .A(n9539), .B(n9538), .Z(n9579) );
  OR2_X1 U9443 ( .A1(n8914), .A2(n8911), .ZN(n9538) );
  OR2_X1 U9444 ( .A1(n9580), .A2(n9581), .ZN(n9539) );
  AND2_X1 U9445 ( .A1(n9582), .A2(n9583), .ZN(n9581) );
  AND2_X1 U9446 ( .A1(n9584), .A2(n9585), .ZN(n9580) );
  OR2_X1 U9447 ( .A1(n9583), .A2(n9582), .ZN(n9585) );
  XOR2_X1 U9448 ( .A(n9586), .B(n9587), .Z(n9540) );
  XOR2_X1 U9449 ( .A(n9588), .B(n9589), .Z(n9587) );
  OR2_X1 U9450 ( .A1(n9590), .A2(n9591), .ZN(n7967) );
  OR2_X1 U9451 ( .A1(n9592), .A2(n7964), .ZN(n9590) );
  AND2_X1 U9452 ( .A1(n7962), .A2(n7963), .ZN(n7964) );
  AND2_X1 U9453 ( .A1(n9593), .A2(n9594), .ZN(n7963) );
  INV_X1 U9454 ( .A(n9595), .ZN(n9593) );
  AND2_X1 U9455 ( .A1(n7958), .A2(n7962), .ZN(n9592) );
  INV_X1 U9456 ( .A(n9596), .ZN(n7962) );
  OR2_X1 U9457 ( .A1(n9597), .A2(n9591), .ZN(n9596) );
  INV_X1 U9458 ( .A(n9598), .ZN(n9591) );
  OR2_X1 U9459 ( .A1(n9599), .A2(n9600), .ZN(n9598) );
  AND2_X1 U9460 ( .A1(n9599), .A2(n9600), .ZN(n9597) );
  OR2_X1 U9461 ( .A1(n9601), .A2(n9602), .ZN(n9600) );
  AND2_X1 U9462 ( .A1(n9603), .A2(n9604), .ZN(n9602) );
  AND2_X1 U9463 ( .A1(n9605), .A2(n9606), .ZN(n9601) );
  OR2_X1 U9464 ( .A1(n9604), .A2(n9603), .ZN(n9606) );
  XOR2_X1 U9465 ( .A(n9550), .B(n9607), .Z(n9599) );
  XOR2_X1 U9466 ( .A(n9549), .B(n9548), .Z(n9607) );
  OR2_X1 U9467 ( .A1(n9297), .A2(n8931), .ZN(n9548) );
  OR2_X1 U9468 ( .A1(n9608), .A2(n9609), .ZN(n9549) );
  AND2_X1 U9469 ( .A1(n9610), .A2(n9611), .ZN(n9609) );
  AND2_X1 U9470 ( .A1(n9612), .A2(n9613), .ZN(n9608) );
  OR2_X1 U9471 ( .A1(n9611), .A2(n9610), .ZN(n9613) );
  XOR2_X1 U9472 ( .A(n9557), .B(n9614), .Z(n9550) );
  XOR2_X1 U9473 ( .A(n9556), .B(n9555), .Z(n9614) );
  OR2_X1 U9474 ( .A1(n8902), .A2(n8927), .ZN(n9555) );
  OR2_X1 U9475 ( .A1(n9615), .A2(n9616), .ZN(n9556) );
  AND2_X1 U9476 ( .A1(n9617), .A2(n9618), .ZN(n9616) );
  AND2_X1 U9477 ( .A1(n9619), .A2(n9620), .ZN(n9615) );
  OR2_X1 U9478 ( .A1(n9618), .A2(n9617), .ZN(n9620) );
  XOR2_X1 U9479 ( .A(n9564), .B(n9621), .Z(n9557) );
  XOR2_X1 U9480 ( .A(n9563), .B(n9562), .Z(n9621) );
  OR2_X1 U9481 ( .A1(n8906), .A2(n8923), .ZN(n9562) );
  OR2_X1 U9482 ( .A1(n9622), .A2(n9623), .ZN(n9563) );
  AND2_X1 U9483 ( .A1(n9624), .A2(n9625), .ZN(n9623) );
  AND2_X1 U9484 ( .A1(n9626), .A2(n9627), .ZN(n9622) );
  OR2_X1 U9485 ( .A1(n9625), .A2(n9624), .ZN(n9627) );
  XOR2_X1 U9486 ( .A(n9571), .B(n9628), .Z(n9564) );
  XOR2_X1 U9487 ( .A(n9570), .B(n9569), .Z(n9628) );
  OR2_X1 U9488 ( .A1(n8910), .A2(n8919), .ZN(n9569) );
  OR2_X1 U9489 ( .A1(n9629), .A2(n9630), .ZN(n9570) );
  AND2_X1 U9490 ( .A1(n9631), .A2(n9632), .ZN(n9630) );
  AND2_X1 U9491 ( .A1(n9633), .A2(n9634), .ZN(n9629) );
  OR2_X1 U9492 ( .A1(n9632), .A2(n9631), .ZN(n9634) );
  XOR2_X1 U9493 ( .A(n9577), .B(n9635), .Z(n9571) );
  XOR2_X1 U9494 ( .A(n9576), .B(n8779), .Z(n9635) );
  OR2_X1 U9495 ( .A1(n8914), .A2(n8915), .ZN(n8779) );
  OR2_X1 U9496 ( .A1(n9636), .A2(n9637), .ZN(n9576) );
  AND2_X1 U9497 ( .A1(n9638), .A2(n9639), .ZN(n9637) );
  AND2_X1 U9498 ( .A1(n9640), .A2(n9641), .ZN(n9636) );
  OR2_X1 U9499 ( .A1(n9639), .A2(n9638), .ZN(n9641) );
  XOR2_X1 U9500 ( .A(n9584), .B(n9642), .Z(n9577) );
  XOR2_X1 U9501 ( .A(n9583), .B(n9582), .Z(n9642) );
  OR2_X1 U9502 ( .A1(n8918), .A2(n8911), .ZN(n9582) );
  OR2_X1 U9503 ( .A1(n9643), .A2(n9644), .ZN(n9583) );
  AND2_X1 U9504 ( .A1(n9645), .A2(n9646), .ZN(n9644) );
  AND2_X1 U9505 ( .A1(n9647), .A2(n9648), .ZN(n9643) );
  OR2_X1 U9506 ( .A1(n9646), .A2(n9645), .ZN(n9648) );
  XOR2_X1 U9507 ( .A(n9649), .B(n9650), .Z(n9584) );
  XOR2_X1 U9508 ( .A(n9651), .B(n9652), .Z(n9650) );
  AND2_X1 U9509 ( .A1(n9195), .A2(n9196), .ZN(n7958) );
  XNOR2_X1 U9510 ( .A(n9594), .B(n9595), .ZN(n9196) );
  OR2_X1 U9511 ( .A1(n9653), .A2(n9654), .ZN(n9595) );
  AND2_X1 U9512 ( .A1(n9655), .A2(n9656), .ZN(n9654) );
  AND2_X1 U9513 ( .A1(n9657), .A2(n9658), .ZN(n9653) );
  OR2_X1 U9514 ( .A1(n9656), .A2(n9655), .ZN(n9658) );
  XNOR2_X1 U9515 ( .A(n9605), .B(n9659), .ZN(n9594) );
  XOR2_X1 U9516 ( .A(n9604), .B(n9603), .Z(n9659) );
  OR2_X1 U9517 ( .A1(n9297), .A2(n8935), .ZN(n9603) );
  OR2_X1 U9518 ( .A1(n9660), .A2(n9661), .ZN(n9604) );
  AND2_X1 U9519 ( .A1(n9662), .A2(n9663), .ZN(n9661) );
  AND2_X1 U9520 ( .A1(n9664), .A2(n9665), .ZN(n9660) );
  OR2_X1 U9521 ( .A1(n9663), .A2(n9662), .ZN(n9665) );
  XOR2_X1 U9522 ( .A(n9612), .B(n9666), .Z(n9605) );
  XOR2_X1 U9523 ( .A(n9611), .B(n9610), .Z(n9666) );
  OR2_X1 U9524 ( .A1(n8902), .A2(n8931), .ZN(n9610) );
  OR2_X1 U9525 ( .A1(n9667), .A2(n9668), .ZN(n9611) );
  AND2_X1 U9526 ( .A1(n9669), .A2(n9670), .ZN(n9668) );
  AND2_X1 U9527 ( .A1(n9671), .A2(n9672), .ZN(n9667) );
  OR2_X1 U9528 ( .A1(n9670), .A2(n9669), .ZN(n9672) );
  XOR2_X1 U9529 ( .A(n9619), .B(n9673), .Z(n9612) );
  XOR2_X1 U9530 ( .A(n9618), .B(n9617), .Z(n9673) );
  OR2_X1 U9531 ( .A1(n8906), .A2(n8927), .ZN(n9617) );
  OR2_X1 U9532 ( .A1(n9674), .A2(n9675), .ZN(n9618) );
  AND2_X1 U9533 ( .A1(n9676), .A2(n9677), .ZN(n9675) );
  AND2_X1 U9534 ( .A1(n9678), .A2(n9679), .ZN(n9674) );
  OR2_X1 U9535 ( .A1(n9677), .A2(n9676), .ZN(n9679) );
  XOR2_X1 U9536 ( .A(n9626), .B(n9680), .Z(n9619) );
  XOR2_X1 U9537 ( .A(n9625), .B(n9624), .Z(n9680) );
  OR2_X1 U9538 ( .A1(n8910), .A2(n8923), .ZN(n9624) );
  OR2_X1 U9539 ( .A1(n9681), .A2(n9682), .ZN(n9625) );
  AND2_X1 U9540 ( .A1(n9683), .A2(n9684), .ZN(n9682) );
  AND2_X1 U9541 ( .A1(n9685), .A2(n9686), .ZN(n9681) );
  OR2_X1 U9542 ( .A1(n9684), .A2(n9683), .ZN(n9686) );
  XOR2_X1 U9543 ( .A(n9633), .B(n9687), .Z(n9626) );
  XOR2_X1 U9544 ( .A(n9632), .B(n9631), .Z(n9687) );
  OR2_X1 U9545 ( .A1(n8914), .A2(n8919), .ZN(n9631) );
  OR2_X1 U9546 ( .A1(n9688), .A2(n9689), .ZN(n9632) );
  AND2_X1 U9547 ( .A1(n8750), .A2(n9690), .ZN(n9689) );
  AND2_X1 U9548 ( .A1(n9691), .A2(n9692), .ZN(n9688) );
  OR2_X1 U9549 ( .A1(n9690), .A2(n8750), .ZN(n9692) );
  XOR2_X1 U9550 ( .A(n9640), .B(n9693), .Z(n9633) );
  XOR2_X1 U9551 ( .A(n9639), .B(n9638), .Z(n9693) );
  OR2_X1 U9552 ( .A1(n8918), .A2(n8915), .ZN(n9638) );
  OR2_X1 U9553 ( .A1(n9694), .A2(n9695), .ZN(n9639) );
  AND2_X1 U9554 ( .A1(n9696), .A2(n9697), .ZN(n9695) );
  AND2_X1 U9555 ( .A1(n9698), .A2(n9699), .ZN(n9694) );
  OR2_X1 U9556 ( .A1(n9697), .A2(n9696), .ZN(n9699) );
  XOR2_X1 U9557 ( .A(n9647), .B(n9700), .Z(n9640) );
  XOR2_X1 U9558 ( .A(n9646), .B(n9645), .Z(n9700) );
  OR2_X1 U9559 ( .A1(n8922), .A2(n8911), .ZN(n9645) );
  OR2_X1 U9560 ( .A1(n9701), .A2(n9702), .ZN(n9646) );
  AND2_X1 U9561 ( .A1(n9703), .A2(n9704), .ZN(n9702) );
  AND2_X1 U9562 ( .A1(n9705), .A2(n9706), .ZN(n9701) );
  OR2_X1 U9563 ( .A1(n9704), .A2(n9703), .ZN(n9706) );
  XOR2_X1 U9564 ( .A(n9707), .B(n9708), .Z(n9647) );
  XOR2_X1 U9565 ( .A(n9709), .B(n9710), .Z(n9708) );
  OR2_X1 U9566 ( .A1(n9711), .A2(n9712), .ZN(n9195) );
  OR2_X1 U9567 ( .A1(n9713), .A2(n9192), .ZN(n9712) );
  AND2_X1 U9568 ( .A1(n9190), .A2(n9191), .ZN(n9192) );
  AND2_X1 U9569 ( .A1(n9714), .A2(n9715), .ZN(n9191) );
  INV_X1 U9570 ( .A(n9716), .ZN(n9714) );
  AND2_X1 U9571 ( .A1(n9186), .A2(n9190), .ZN(n9713) );
  INV_X1 U9572 ( .A(n9717), .ZN(n9190) );
  OR2_X1 U9573 ( .A1(n9718), .A2(n9711), .ZN(n9717) );
  AND2_X1 U9574 ( .A1(n9719), .A2(n9720), .ZN(n9718) );
  AND2_X1 U9575 ( .A1(n9182), .A2(n9183), .ZN(n9186) );
  XNOR2_X1 U9576 ( .A(n9715), .B(n9716), .ZN(n9183) );
  OR2_X1 U9577 ( .A1(n9721), .A2(n9722), .ZN(n9716) );
  AND2_X1 U9578 ( .A1(n9723), .A2(n9724), .ZN(n9722) );
  AND2_X1 U9579 ( .A1(n9725), .A2(n9726), .ZN(n9721) );
  OR2_X1 U9580 ( .A1(n9724), .A2(n9723), .ZN(n9726) );
  XNOR2_X1 U9581 ( .A(n9727), .B(n9728), .ZN(n9715) );
  XOR2_X1 U9582 ( .A(n9729), .B(n9730), .Z(n9728) );
  OR2_X1 U9583 ( .A1(n9731), .A2(n9732), .ZN(n9182) );
  OR2_X1 U9584 ( .A1(n9733), .A2(n9179), .ZN(n9732) );
  AND2_X1 U9585 ( .A1(n9177), .A2(n9178), .ZN(n9179) );
  AND2_X1 U9586 ( .A1(n9734), .A2(n9735), .ZN(n9178) );
  INV_X1 U9587 ( .A(n9736), .ZN(n9734) );
  AND2_X1 U9588 ( .A1(n9177), .A2(n9173), .ZN(n9733) );
  OR2_X1 U9589 ( .A1(n9737), .A2(n9166), .ZN(n9173) );
  AND2_X1 U9590 ( .A1(n9169), .A2(n9738), .ZN(n9166) );
  AND2_X1 U9591 ( .A1(n9170), .A2(n9168), .ZN(n9738) );
  AND2_X1 U9592 ( .A1(n9168), .A2(n9162), .ZN(n9737) );
  OR2_X1 U9593 ( .A1(n9739), .A2(n9740), .ZN(n9162) );
  INV_X1 U9594 ( .A(n9159), .ZN(n9740) );
  OR2_X1 U9595 ( .A1(n9741), .A2(n9742), .ZN(n9159) );
  OR2_X1 U9596 ( .A1(n9743), .A2(n9744), .ZN(n9742) );
  AND2_X1 U9597 ( .A1(n9156), .A2(n9158), .ZN(n9739) );
  INV_X1 U9598 ( .A(n9745), .ZN(n9158) );
  AND2_X1 U9599 ( .A1(n9746), .A2(n9744), .ZN(n9745) );
  XNOR2_X1 U9600 ( .A(n9170), .B(n9169), .ZN(n9744) );
  INV_X1 U9601 ( .A(n9747), .ZN(n9169) );
  OR2_X1 U9602 ( .A1(n9748), .A2(n9749), .ZN(n9747) );
  AND2_X1 U9603 ( .A1(n9750), .A2(n9751), .ZN(n9749) );
  AND2_X1 U9604 ( .A1(n9752), .A2(n9753), .ZN(n9748) );
  OR2_X1 U9605 ( .A1(n9751), .A2(n9750), .ZN(n9753) );
  XNOR2_X1 U9606 ( .A(n9754), .B(n9755), .ZN(n9170) );
  XOR2_X1 U9607 ( .A(n9756), .B(n9757), .Z(n9755) );
  OR2_X1 U9608 ( .A1(n9741), .A2(n9743), .ZN(n9746) );
  OR2_X1 U9609 ( .A1(n9758), .A2(n9153), .ZN(n9156) );
  AND2_X1 U9610 ( .A1(n9759), .A2(n9760), .ZN(n9153) );
  AND2_X1 U9611 ( .A1(n9149), .A2(n9152), .ZN(n9758) );
  OR2_X1 U9612 ( .A1(n9760), .A2(n9759), .ZN(n9152) );
  XOR2_X1 U9613 ( .A(n9743), .B(n9741), .Z(n9759) );
  OR2_X1 U9614 ( .A1(n9761), .A2(n9762), .ZN(n9741) );
  AND2_X1 U9615 ( .A1(n9763), .A2(n9764), .ZN(n9762) );
  AND2_X1 U9616 ( .A1(n9765), .A2(n9766), .ZN(n9761) );
  OR2_X1 U9617 ( .A1(n9763), .A2(n9764), .ZN(n9766) );
  XOR2_X1 U9618 ( .A(n9752), .B(n9767), .Z(n9743) );
  XOR2_X1 U9619 ( .A(n9751), .B(n9750), .Z(n9767) );
  OR2_X1 U9620 ( .A1(n9297), .A2(n8959), .ZN(n9750) );
  OR2_X1 U9621 ( .A1(n9768), .A2(n9769), .ZN(n9751) );
  AND2_X1 U9622 ( .A1(n9770), .A2(n9771), .ZN(n9769) );
  AND2_X1 U9623 ( .A1(n9772), .A2(n9773), .ZN(n9768) );
  OR2_X1 U9624 ( .A1(n9771), .A2(n9770), .ZN(n9773) );
  XOR2_X1 U9625 ( .A(n9774), .B(n9775), .Z(n9752) );
  XOR2_X1 U9626 ( .A(n9776), .B(n9777), .Z(n9775) );
  INV_X1 U9627 ( .A(n9778), .ZN(n9760) );
  OR2_X1 U9628 ( .A1(n9779), .A2(n9146), .ZN(n9149) );
  AND2_X1 U9629 ( .A1(n9780), .A2(n9781), .ZN(n9146) );
  AND2_X1 U9630 ( .A1(n9778), .A2(n9782), .ZN(n9780) );
  INV_X1 U9631 ( .A(n9783), .ZN(n9782) );
  AND2_X1 U9632 ( .A1(n9784), .A2(n9785), .ZN(n9783) );
  OR2_X1 U9633 ( .A1(n9784), .A2(n9785), .ZN(n9778) );
  AND2_X1 U9634 ( .A1(n9144), .A2(n9142), .ZN(n9779) );
  OR2_X1 U9635 ( .A1(n9786), .A2(n9787), .ZN(n9142) );
  AND2_X1 U9636 ( .A1(n9133), .A2(n9136), .ZN(n9787) );
  OR2_X1 U9637 ( .A1(n9788), .A2(n9139), .ZN(n9136) );
  OR2_X1 U9638 ( .A1(n9789), .A2(n9130), .ZN(n9133) );
  AND2_X1 U9639 ( .A1(n9790), .A2(n9791), .ZN(n9130) );
  AND2_X1 U9640 ( .A1(n9126), .A2(n9128), .ZN(n9789) );
  OR2_X1 U9641 ( .A1(n9791), .A2(n9790), .ZN(n9128) );
  XOR2_X1 U9642 ( .A(n9792), .B(n9793), .Z(n9790) );
  OR2_X1 U9643 ( .A1(n9794), .A2(n9795), .ZN(n9126) );
  INV_X1 U9644 ( .A(n9112), .ZN(n9795) );
  OR2_X1 U9645 ( .A1(n9796), .A2(n9797), .ZN(n9112) );
  AND2_X1 U9646 ( .A1(n9109), .A2(n9111), .ZN(n9794) );
  INV_X1 U9647 ( .A(n9798), .ZN(n9111) );
  AND2_X1 U9648 ( .A1(n9797), .A2(n9796), .ZN(n9798) );
  OR2_X1 U9649 ( .A1(n9799), .A2(n9791), .ZN(n9797) );
  INV_X1 U9650 ( .A(n9800), .ZN(n9791) );
  OR2_X1 U9651 ( .A1(n9801), .A2(n9802), .ZN(n9800) );
  AND2_X1 U9652 ( .A1(n9801), .A2(n9802), .ZN(n9799) );
  OR2_X1 U9653 ( .A1(n9803), .A2(n9804), .ZN(n9802) );
  AND2_X1 U9654 ( .A1(n9805), .A2(n9806), .ZN(n9804) );
  AND2_X1 U9655 ( .A1(n9807), .A2(n9808), .ZN(n9803) );
  OR2_X1 U9656 ( .A1(n9805), .A2(n9806), .ZN(n9807) );
  XOR2_X1 U9657 ( .A(n9809), .B(n9810), .Z(n9801) );
  XOR2_X1 U9658 ( .A(n9811), .B(n9812), .Z(n9810) );
  OR2_X1 U9659 ( .A1(n9813), .A2(n9106), .ZN(n9109) );
  AND2_X1 U9660 ( .A1(n9814), .A2(n9815), .ZN(n9106) );
  AND2_X1 U9661 ( .A1(n9104), .A2(n9102), .ZN(n9813) );
  OR2_X1 U9662 ( .A1(n9816), .A2(n9817), .ZN(n9102) );
  AND2_X1 U9663 ( .A1(n9096), .A2(n9093), .ZN(n9817) );
  OR2_X1 U9664 ( .A1(n9818), .A2(n9090), .ZN(n9093) );
  AND2_X1 U9665 ( .A1(n9819), .A2(n9820), .ZN(n9090) );
  AND2_X1 U9666 ( .A1(n9088), .A2(n9086), .ZN(n9818) );
  OR2_X1 U9667 ( .A1(n9821), .A2(n9083), .ZN(n9086) );
  AND2_X1 U9668 ( .A1(n9822), .A2(n9823), .ZN(n9083) );
  AND2_X1 U9669 ( .A1(n9079), .A2(n9082), .ZN(n9821) );
  OR2_X1 U9670 ( .A1(n9823), .A2(n9822), .ZN(n9082) );
  XNOR2_X1 U9671 ( .A(n9824), .B(n9825), .ZN(n9822) );
  OR2_X1 U9672 ( .A1(n9826), .A2(n9827), .ZN(n9079) );
  INV_X1 U9673 ( .A(n9075), .ZN(n9827) );
  OR2_X1 U9674 ( .A1(n9828), .A2(n9829), .ZN(n9075) );
  AND2_X1 U9675 ( .A1(n9073), .A2(n9076), .ZN(n9826) );
  INV_X1 U9676 ( .A(n9830), .ZN(n9076) );
  AND2_X1 U9677 ( .A1(n9829), .A2(n9828), .ZN(n9830) );
  OR2_X1 U9678 ( .A1(n9831), .A2(n9823), .ZN(n9828) );
  INV_X1 U9679 ( .A(n9832), .ZN(n9823) );
  OR2_X1 U9680 ( .A1(n9833), .A2(n9834), .ZN(n9832) );
  AND2_X1 U9681 ( .A1(n9833), .A2(n9834), .ZN(n9831) );
  OR2_X1 U9682 ( .A1(n9835), .A2(n9836), .ZN(n9834) );
  AND2_X1 U9683 ( .A1(n9837), .A2(n9838), .ZN(n9836) );
  AND2_X1 U9684 ( .A1(n9839), .A2(n9840), .ZN(n9835) );
  OR2_X1 U9685 ( .A1(n9837), .A2(n9838), .ZN(n9840) );
  XOR2_X1 U9686 ( .A(n9841), .B(n9842), .Z(n9833) );
  XOR2_X1 U9687 ( .A(n9843), .B(n9844), .Z(n9842) );
  OR2_X1 U9688 ( .A1(n9845), .A2(n9846), .ZN(n9829) );
  OR2_X1 U9689 ( .A1(n9847), .A2(n9070), .ZN(n9073) );
  AND2_X1 U9690 ( .A1(n9848), .A2(n9849), .ZN(n9070) );
  AND2_X1 U9691 ( .A1(n9068), .A2(n9066), .ZN(n9847) );
  OR2_X1 U9692 ( .A1(n9850), .A2(n9063), .ZN(n9066) );
  AND2_X1 U9693 ( .A1(n9851), .A2(n9852), .ZN(n9063) );
  AND2_X1 U9694 ( .A1(n9061), .A2(n9059), .ZN(n9850) );
  OR2_X1 U9695 ( .A1(n9853), .A2(n9854), .ZN(n9059) );
  INV_X1 U9696 ( .A(n9056), .ZN(n9854) );
  OR2_X1 U9697 ( .A1(n9855), .A2(n9856), .ZN(n9056) );
  OR2_X1 U9698 ( .A1(n9857), .A2(n9858), .ZN(n9856) );
  XNOR2_X1 U9699 ( .A(n9859), .B(n9860), .ZN(n9858) );
  INV_X1 U9700 ( .A(n9861), .ZN(n9857) );
  AND2_X1 U9701 ( .A1(n9055), .A2(n9053), .ZN(n9853) );
  OR2_X1 U9702 ( .A1(n9862), .A2(n9049), .ZN(n9053) );
  INV_X1 U9703 ( .A(n9863), .ZN(n9049) );
  OR2_X1 U9704 ( .A1(n9864), .A2(n9865), .ZN(n9863) );
  OR2_X1 U9705 ( .A1(n9866), .A2(n9867), .ZN(n9865) );
  AND2_X1 U9706 ( .A1(n9046), .A2(n9868), .ZN(n9862) );
  INV_X1 U9707 ( .A(n9050), .ZN(n9868) );
  AND2_X1 U9708 ( .A1(n9869), .A2(n9866), .ZN(n9050) );
  XNOR2_X1 U9709 ( .A(n9861), .B(n9870), .ZN(n9866) );
  OR2_X1 U9710 ( .A1(n9864), .A2(n9867), .ZN(n9869) );
  AND2_X1 U9711 ( .A1(n9036), .A2(n9871), .ZN(n9046) );
  AND2_X1 U9712 ( .A1(n9030), .A2(n9035), .ZN(n9871) );
  XOR2_X1 U9713 ( .A(n9867), .B(n9864), .Z(n9035) );
  OR2_X1 U9714 ( .A1(n9872), .A2(n9873), .ZN(n9864) );
  AND2_X1 U9715 ( .A1(n9874), .A2(n9875), .ZN(n9873) );
  AND2_X1 U9716 ( .A1(n9876), .A2(n9877), .ZN(n9872) );
  OR2_X1 U9717 ( .A1(n9874), .A2(n9875), .ZN(n9877) );
  XOR2_X1 U9718 ( .A(n9878), .B(n9879), .Z(n9867) );
  XOR2_X1 U9719 ( .A(n9880), .B(n9881), .Z(n9879) );
  XNOR2_X1 U9720 ( .A(n9876), .B(n9882), .ZN(n9030) );
  XOR2_X1 U9721 ( .A(n9875), .B(n9874), .Z(n9882) );
  OR2_X1 U9722 ( .A1(n9297), .A2(n7998), .ZN(n9874) );
  OR2_X1 U9723 ( .A1(n9883), .A2(n9884), .ZN(n9875) );
  AND2_X1 U9724 ( .A1(n9885), .A2(n9886), .ZN(n9884) );
  AND2_X1 U9725 ( .A1(n9887), .A2(n9888), .ZN(n9883) );
  OR2_X1 U9726 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  XOR2_X1 U9727 ( .A(n9889), .B(n9890), .Z(n9876) );
  XOR2_X1 U9728 ( .A(n9891), .B(n9892), .Z(n9890) );
  INV_X1 U9729 ( .A(n9029), .ZN(n9036) );
  OR2_X1 U9730 ( .A1(n9893), .A2(n9894), .ZN(n9029) );
  AND2_X1 U9731 ( .A1(n9026), .A2(n9025), .ZN(n9894) );
  AND2_X1 U9732 ( .A1(n9023), .A2(n9895), .ZN(n9893) );
  OR2_X1 U9733 ( .A1(n9026), .A2(n9025), .ZN(n9895) );
  OR2_X1 U9734 ( .A1(n9896), .A2(n9897), .ZN(n9025) );
  AND2_X1 U9735 ( .A1(n8876), .A2(n8875), .ZN(n9897) );
  AND2_X1 U9736 ( .A1(n8873), .A2(n9898), .ZN(n9896) );
  OR2_X1 U9737 ( .A1(n8876), .A2(n8875), .ZN(n9898) );
  OR2_X1 U9738 ( .A1(n9899), .A2(n9900), .ZN(n8875) );
  AND2_X1 U9739 ( .A1(n8847), .A2(n8846), .ZN(n9900) );
  AND2_X1 U9740 ( .A1(n8844), .A2(n9901), .ZN(n9899) );
  OR2_X1 U9741 ( .A1(n8847), .A2(n8846), .ZN(n9901) );
  OR2_X1 U9742 ( .A1(n9902), .A2(n9903), .ZN(n8846) );
  AND2_X1 U9743 ( .A1(n8818), .A2(n8817), .ZN(n9903) );
  AND2_X1 U9744 ( .A1(n8815), .A2(n9904), .ZN(n9902) );
  OR2_X1 U9745 ( .A1(n8818), .A2(n8817), .ZN(n9904) );
  OR2_X1 U9746 ( .A1(n9905), .A2(n9906), .ZN(n8817) );
  AND2_X1 U9747 ( .A1(n8789), .A2(n8788), .ZN(n9906) );
  AND2_X1 U9748 ( .A1(n8786), .A2(n9907), .ZN(n9905) );
  OR2_X1 U9749 ( .A1(n8789), .A2(n8788), .ZN(n9907) );
  OR2_X1 U9750 ( .A1(n9908), .A2(n9909), .ZN(n8788) );
  AND2_X1 U9751 ( .A1(n8760), .A2(n8759), .ZN(n9909) );
  AND2_X1 U9752 ( .A1(n8757), .A2(n9910), .ZN(n9908) );
  OR2_X1 U9753 ( .A1(n8760), .A2(n8759), .ZN(n9910) );
  OR2_X1 U9754 ( .A1(n9911), .A2(n9912), .ZN(n8759) );
  AND2_X1 U9755 ( .A1(n8731), .A2(n8730), .ZN(n9912) );
  AND2_X1 U9756 ( .A1(n8728), .A2(n9913), .ZN(n9911) );
  OR2_X1 U9757 ( .A1(n8731), .A2(n8730), .ZN(n9913) );
  OR2_X1 U9758 ( .A1(n9914), .A2(n9915), .ZN(n8730) );
  AND2_X1 U9759 ( .A1(n8702), .A2(n8701), .ZN(n9915) );
  AND2_X1 U9760 ( .A1(n8699), .A2(n9916), .ZN(n9914) );
  OR2_X1 U9761 ( .A1(n8702), .A2(n8701), .ZN(n9916) );
  OR2_X1 U9762 ( .A1(n9917), .A2(n9918), .ZN(n8701) );
  AND2_X1 U9763 ( .A1(n8664), .A2(n8663), .ZN(n9918) );
  AND2_X1 U9764 ( .A1(n8661), .A2(n9919), .ZN(n9917) );
  OR2_X1 U9765 ( .A1(n8664), .A2(n8663), .ZN(n9919) );
  OR2_X1 U9766 ( .A1(n9920), .A2(n9921), .ZN(n8663) );
  AND2_X1 U9767 ( .A1(n8635), .A2(n8634), .ZN(n9921) );
  AND2_X1 U9768 ( .A1(n8632), .A2(n9922), .ZN(n9920) );
  OR2_X1 U9769 ( .A1(n8635), .A2(n8634), .ZN(n9922) );
  OR2_X1 U9770 ( .A1(n9923), .A2(n9924), .ZN(n8634) );
  AND2_X1 U9771 ( .A1(n8606), .A2(n8605), .ZN(n9924) );
  AND2_X1 U9772 ( .A1(n8603), .A2(n9925), .ZN(n9923) );
  OR2_X1 U9773 ( .A1(n8606), .A2(n8605), .ZN(n9925) );
  OR2_X1 U9774 ( .A1(n9926), .A2(n9927), .ZN(n8605) );
  AND2_X1 U9775 ( .A1(n8577), .A2(n8576), .ZN(n9927) );
  AND2_X1 U9776 ( .A1(n8574), .A2(n9928), .ZN(n9926) );
  OR2_X1 U9777 ( .A1(n8577), .A2(n8576), .ZN(n9928) );
  OR2_X1 U9778 ( .A1(n9929), .A2(n9930), .ZN(n8576) );
  AND2_X1 U9779 ( .A1(n8548), .A2(n8547), .ZN(n9930) );
  AND2_X1 U9780 ( .A1(n8545), .A2(n9931), .ZN(n9929) );
  OR2_X1 U9781 ( .A1(n8548), .A2(n8547), .ZN(n9931) );
  OR2_X1 U9782 ( .A1(n9932), .A2(n9933), .ZN(n8547) );
  AND2_X1 U9783 ( .A1(n8519), .A2(n8518), .ZN(n9933) );
  AND2_X1 U9784 ( .A1(n8516), .A2(n9934), .ZN(n9932) );
  OR2_X1 U9785 ( .A1(n8519), .A2(n8518), .ZN(n9934) );
  OR2_X1 U9786 ( .A1(n9935), .A2(n9936), .ZN(n8518) );
  AND2_X1 U9787 ( .A1(n8490), .A2(n8489), .ZN(n9936) );
  AND2_X1 U9788 ( .A1(n8487), .A2(n9937), .ZN(n9935) );
  OR2_X1 U9789 ( .A1(n8490), .A2(n8489), .ZN(n9937) );
  OR2_X1 U9790 ( .A1(n9938), .A2(n9939), .ZN(n8489) );
  AND2_X1 U9791 ( .A1(n8461), .A2(n8460), .ZN(n9939) );
  AND2_X1 U9792 ( .A1(n8458), .A2(n9940), .ZN(n9938) );
  OR2_X1 U9793 ( .A1(n8461), .A2(n8460), .ZN(n9940) );
  OR2_X1 U9794 ( .A1(n9941), .A2(n9942), .ZN(n8460) );
  AND2_X1 U9795 ( .A1(n8432), .A2(n8431), .ZN(n9942) );
  AND2_X1 U9796 ( .A1(n8429), .A2(n9943), .ZN(n9941) );
  OR2_X1 U9797 ( .A1(n8432), .A2(n8431), .ZN(n9943) );
  OR2_X1 U9798 ( .A1(n9944), .A2(n9945), .ZN(n8431) );
  AND2_X1 U9799 ( .A1(n8403), .A2(n8402), .ZN(n9945) );
  AND2_X1 U9800 ( .A1(n8400), .A2(n9946), .ZN(n9944) );
  OR2_X1 U9801 ( .A1(n8403), .A2(n8402), .ZN(n9946) );
  OR2_X1 U9802 ( .A1(n9947), .A2(n9948), .ZN(n8402) );
  AND2_X1 U9803 ( .A1(n8370), .A2(n8369), .ZN(n9948) );
  AND2_X1 U9804 ( .A1(n8367), .A2(n9949), .ZN(n9947) );
  OR2_X1 U9805 ( .A1(n8370), .A2(n8369), .ZN(n9949) );
  OR2_X1 U9806 ( .A1(n9950), .A2(n9951), .ZN(n8369) );
  AND2_X1 U9807 ( .A1(n8341), .A2(n8340), .ZN(n9951) );
  AND2_X1 U9808 ( .A1(n8338), .A2(n9952), .ZN(n9950) );
  OR2_X1 U9809 ( .A1(n8341), .A2(n8340), .ZN(n9952) );
  OR2_X1 U9810 ( .A1(n9953), .A2(n9954), .ZN(n8340) );
  AND2_X1 U9811 ( .A1(n8313), .A2(n8312), .ZN(n9954) );
  AND2_X1 U9812 ( .A1(n8310), .A2(n9955), .ZN(n9953) );
  OR2_X1 U9813 ( .A1(n8313), .A2(n8312), .ZN(n9955) );
  OR2_X1 U9814 ( .A1(n9956), .A2(n9957), .ZN(n8312) );
  AND2_X1 U9815 ( .A1(n8285), .A2(n8284), .ZN(n9957) );
  AND2_X1 U9816 ( .A1(n8282), .A2(n9958), .ZN(n9956) );
  OR2_X1 U9817 ( .A1(n8285), .A2(n8284), .ZN(n9958) );
  OR2_X1 U9818 ( .A1(n9959), .A2(n9960), .ZN(n8284) );
  AND2_X1 U9819 ( .A1(n8257), .A2(n8256), .ZN(n9960) );
  AND2_X1 U9820 ( .A1(n8254), .A2(n9961), .ZN(n9959) );
  OR2_X1 U9821 ( .A1(n8257), .A2(n8256), .ZN(n9961) );
  OR2_X1 U9822 ( .A1(n9962), .A2(n9963), .ZN(n8256) );
  AND2_X1 U9823 ( .A1(n8229), .A2(n8228), .ZN(n9963) );
  AND2_X1 U9824 ( .A1(n8226), .A2(n9964), .ZN(n9962) );
  OR2_X1 U9825 ( .A1(n8229), .A2(n8228), .ZN(n9964) );
  OR2_X1 U9826 ( .A1(n9965), .A2(n9966), .ZN(n8228) );
  AND2_X1 U9827 ( .A1(n8201), .A2(n8200), .ZN(n9966) );
  AND2_X1 U9828 ( .A1(n8198), .A2(n9967), .ZN(n9965) );
  OR2_X1 U9829 ( .A1(n8201), .A2(n8200), .ZN(n9967) );
  OR2_X1 U9830 ( .A1(n9968), .A2(n9969), .ZN(n8200) );
  AND2_X1 U9831 ( .A1(n8173), .A2(n8172), .ZN(n9969) );
  AND2_X1 U9832 ( .A1(n8170), .A2(n9970), .ZN(n9968) );
  OR2_X1 U9833 ( .A1(n8173), .A2(n8172), .ZN(n9970) );
  OR2_X1 U9834 ( .A1(n9971), .A2(n9972), .ZN(n8172) );
  AND2_X1 U9835 ( .A1(n8145), .A2(n8144), .ZN(n9972) );
  AND2_X1 U9836 ( .A1(n8142), .A2(n9973), .ZN(n9971) );
  OR2_X1 U9837 ( .A1(n8145), .A2(n8144), .ZN(n9973) );
  OR2_X1 U9838 ( .A1(n9974), .A2(n9975), .ZN(n8144) );
  AND2_X1 U9839 ( .A1(n8117), .A2(n8116), .ZN(n9975) );
  AND2_X1 U9840 ( .A1(n8114), .A2(n9976), .ZN(n9974) );
  OR2_X1 U9841 ( .A1(n8117), .A2(n8116), .ZN(n9976) );
  OR2_X1 U9842 ( .A1(n9977), .A2(n9978), .ZN(n8116) );
  AND2_X1 U9843 ( .A1(n8080), .A2(n8079), .ZN(n9978) );
  AND2_X1 U9844 ( .A1(n8077), .A2(n9979), .ZN(n9977) );
  OR2_X1 U9845 ( .A1(n8080), .A2(n8079), .ZN(n9979) );
  OR2_X1 U9846 ( .A1(n9980), .A2(n9981), .ZN(n8079) );
  AND2_X1 U9847 ( .A1(n8050), .A2(n8051), .ZN(n9981) );
  AND2_X1 U9848 ( .A1(n9982), .A2(n9983), .ZN(n9980) );
  OR2_X1 U9849 ( .A1(n8050), .A2(n8051), .ZN(n9983) );
  OR2_X1 U9850 ( .A1(n9014), .A2(n9388), .ZN(n8051) );
  OR2_X1 U9851 ( .A1(n7998), .A2(n9016), .ZN(n8050) );
  OR2_X1 U9852 ( .A1(n9388), .A2(n9984), .ZN(n9016) );
  INV_X1 U9853 ( .A(n8052), .ZN(n9982) );
  OR2_X1 U9854 ( .A1(n9985), .A2(n9986), .ZN(n8052) );
  AND2_X1 U9855 ( .A1(b_30_), .A2(n9987), .ZN(n9986) );
  OR2_X1 U9856 ( .A1(n9988), .A2(n9989), .ZN(n9987) );
  AND2_X1 U9857 ( .A1(a_30_), .A2(n8047), .ZN(n9988) );
  AND2_X1 U9858 ( .A1(b_29_), .A2(n9990), .ZN(n9985) );
  OR2_X1 U9859 ( .A1(n9991), .A2(n8021), .ZN(n9990) );
  AND2_X1 U9860 ( .A1(a_31_), .A2(n7998), .ZN(n9991) );
  OR2_X1 U9861 ( .A1(n9010), .A2(n9388), .ZN(n8080) );
  XOR2_X1 U9862 ( .A(n9992), .B(n9993), .Z(n8077) );
  XNOR2_X1 U9863 ( .A(n9994), .B(n9995), .ZN(n9992) );
  OR2_X1 U9864 ( .A1(n9006), .A2(n9388), .ZN(n8117) );
  XOR2_X1 U9865 ( .A(n9996), .B(n9997), .Z(n8114) );
  XOR2_X1 U9866 ( .A(n9998), .B(n9999), .Z(n9997) );
  OR2_X1 U9867 ( .A1(n9002), .A2(n9388), .ZN(n8145) );
  XNOR2_X1 U9868 ( .A(n10000), .B(n10001), .ZN(n8142) );
  XNOR2_X1 U9869 ( .A(n10002), .B(n10003), .ZN(n10000) );
  OR2_X1 U9870 ( .A1(n8998), .A2(n9388), .ZN(n8173) );
  XOR2_X1 U9871 ( .A(n10004), .B(n10005), .Z(n8170) );
  XOR2_X1 U9872 ( .A(n10006), .B(n10007), .Z(n10005) );
  OR2_X1 U9873 ( .A1(n8994), .A2(n9388), .ZN(n8201) );
  XOR2_X1 U9874 ( .A(n10008), .B(n10009), .Z(n8198) );
  XOR2_X1 U9875 ( .A(n10010), .B(n10011), .Z(n10009) );
  OR2_X1 U9876 ( .A1(n8990), .A2(n9388), .ZN(n8229) );
  XOR2_X1 U9877 ( .A(n10012), .B(n10013), .Z(n8226) );
  XOR2_X1 U9878 ( .A(n10014), .B(n10015), .Z(n10013) );
  OR2_X1 U9879 ( .A1(n8986), .A2(n9388), .ZN(n8257) );
  XOR2_X1 U9880 ( .A(n10016), .B(n10017), .Z(n8254) );
  XOR2_X1 U9881 ( .A(n10018), .B(n10019), .Z(n10017) );
  OR2_X1 U9882 ( .A1(n8982), .A2(n9388), .ZN(n8285) );
  XOR2_X1 U9883 ( .A(n10020), .B(n10021), .Z(n8282) );
  XOR2_X1 U9884 ( .A(n10022), .B(n10023), .Z(n10021) );
  OR2_X1 U9885 ( .A1(n8978), .A2(n9388), .ZN(n8313) );
  XOR2_X1 U9886 ( .A(n10024), .B(n10025), .Z(n8310) );
  XOR2_X1 U9887 ( .A(n10026), .B(n10027), .Z(n10025) );
  OR2_X1 U9888 ( .A1(n8974), .A2(n9388), .ZN(n8341) );
  XOR2_X1 U9889 ( .A(n10028), .B(n10029), .Z(n8338) );
  XOR2_X1 U9890 ( .A(n10030), .B(n10031), .Z(n10029) );
  OR2_X1 U9891 ( .A1(n8970), .A2(n9388), .ZN(n8370) );
  XOR2_X1 U9892 ( .A(n10032), .B(n10033), .Z(n8367) );
  XOR2_X1 U9893 ( .A(n10034), .B(n10035), .Z(n10033) );
  OR2_X1 U9894 ( .A1(n8966), .A2(n9388), .ZN(n8403) );
  XOR2_X1 U9895 ( .A(n10036), .B(n10037), .Z(n8400) );
  XOR2_X1 U9896 ( .A(n10038), .B(n10039), .Z(n10037) );
  OR2_X1 U9897 ( .A1(n8962), .A2(n9388), .ZN(n8432) );
  XOR2_X1 U9898 ( .A(n10040), .B(n10041), .Z(n8429) );
  XOR2_X1 U9899 ( .A(n10042), .B(n10043), .Z(n10041) );
  OR2_X1 U9900 ( .A1(n8958), .A2(n9388), .ZN(n8461) );
  XOR2_X1 U9901 ( .A(n10044), .B(n10045), .Z(n8458) );
  XOR2_X1 U9902 ( .A(n10046), .B(n10047), .Z(n10045) );
  OR2_X1 U9903 ( .A1(n8954), .A2(n9388), .ZN(n8490) );
  XOR2_X1 U9904 ( .A(n10048), .B(n10049), .Z(n8487) );
  XOR2_X1 U9905 ( .A(n10050), .B(n10051), .Z(n10049) );
  OR2_X1 U9906 ( .A1(n8950), .A2(n9388), .ZN(n8519) );
  XOR2_X1 U9907 ( .A(n10052), .B(n10053), .Z(n8516) );
  XOR2_X1 U9908 ( .A(n10054), .B(n10055), .Z(n10053) );
  OR2_X1 U9909 ( .A1(n8946), .A2(n9388), .ZN(n8548) );
  XOR2_X1 U9910 ( .A(n10056), .B(n10057), .Z(n8545) );
  XOR2_X1 U9911 ( .A(n10058), .B(n10059), .Z(n10057) );
  OR2_X1 U9912 ( .A1(n8942), .A2(n9388), .ZN(n8577) );
  XOR2_X1 U9913 ( .A(n10060), .B(n10061), .Z(n8574) );
  XOR2_X1 U9914 ( .A(n10062), .B(n10063), .Z(n10061) );
  OR2_X1 U9915 ( .A1(n8938), .A2(n9388), .ZN(n8606) );
  XOR2_X1 U9916 ( .A(n10064), .B(n10065), .Z(n8603) );
  XOR2_X1 U9917 ( .A(n10066), .B(n10067), .Z(n10065) );
  OR2_X1 U9918 ( .A1(n8934), .A2(n9388), .ZN(n8635) );
  XOR2_X1 U9919 ( .A(n10068), .B(n10069), .Z(n8632) );
  XOR2_X1 U9920 ( .A(n10070), .B(n10071), .Z(n10069) );
  OR2_X1 U9921 ( .A1(n8930), .A2(n9388), .ZN(n8664) );
  XOR2_X1 U9922 ( .A(n10072), .B(n10073), .Z(n8661) );
  XOR2_X1 U9923 ( .A(n10074), .B(n10075), .Z(n10073) );
  OR2_X1 U9924 ( .A1(n8926), .A2(n9388), .ZN(n8702) );
  XOR2_X1 U9925 ( .A(n10076), .B(n10077), .Z(n8699) );
  XOR2_X1 U9926 ( .A(n10078), .B(n10079), .Z(n10077) );
  OR2_X1 U9927 ( .A1(n8922), .A2(n9388), .ZN(n8731) );
  XOR2_X1 U9928 ( .A(n10080), .B(n10081), .Z(n8728) );
  XOR2_X1 U9929 ( .A(n10082), .B(n10083), .Z(n10081) );
  OR2_X1 U9930 ( .A1(n8918), .A2(n9388), .ZN(n8760) );
  XOR2_X1 U9931 ( .A(n10084), .B(n10085), .Z(n8757) );
  XOR2_X1 U9932 ( .A(n10086), .B(n10087), .Z(n10085) );
  OR2_X1 U9933 ( .A1(n8914), .A2(n9388), .ZN(n8789) );
  XOR2_X1 U9934 ( .A(n10088), .B(n10089), .Z(n8786) );
  XOR2_X1 U9935 ( .A(n10090), .B(n10091), .Z(n10089) );
  OR2_X1 U9936 ( .A1(n8910), .A2(n9388), .ZN(n8818) );
  XOR2_X1 U9937 ( .A(n10092), .B(n10093), .Z(n8815) );
  XOR2_X1 U9938 ( .A(n10094), .B(n10095), .Z(n10093) );
  OR2_X1 U9939 ( .A1(n8906), .A2(n9388), .ZN(n8847) );
  XOR2_X1 U9940 ( .A(n10096), .B(n10097), .Z(n8844) );
  XOR2_X1 U9941 ( .A(n10098), .B(n10099), .Z(n10097) );
  OR2_X1 U9942 ( .A1(n8902), .A2(n9388), .ZN(n8876) );
  XOR2_X1 U9943 ( .A(n10100), .B(n10101), .Z(n8873) );
  XOR2_X1 U9944 ( .A(n10102), .B(n10103), .Z(n10101) );
  OR2_X1 U9945 ( .A1(n9297), .A2(n9388), .ZN(n9026) );
  INV_X1 U9946 ( .A(b_31_), .ZN(n9388) );
  XOR2_X1 U9947 ( .A(n9885), .B(n10104), .Z(n9023) );
  XOR2_X1 U9948 ( .A(n9888), .B(n9886), .Z(n10104) );
  OR2_X1 U9949 ( .A1(n8902), .A2(n7998), .ZN(n9886) );
  OR2_X1 U9950 ( .A1(n10105), .A2(n10106), .ZN(n9888) );
  AND2_X1 U9951 ( .A1(n10100), .A2(n10103), .ZN(n10106) );
  AND2_X1 U9952 ( .A1(n10107), .A2(n10102), .ZN(n10105) );
  OR2_X1 U9953 ( .A1(n10108), .A2(n10109), .ZN(n10102) );
  AND2_X1 U9954 ( .A1(n10096), .A2(n10099), .ZN(n10109) );
  AND2_X1 U9955 ( .A1(n10110), .A2(n10098), .ZN(n10108) );
  OR2_X1 U9956 ( .A1(n10111), .A2(n10112), .ZN(n10098) );
  AND2_X1 U9957 ( .A1(n10092), .A2(n10095), .ZN(n10112) );
  AND2_X1 U9958 ( .A1(n10113), .A2(n10094), .ZN(n10111) );
  OR2_X1 U9959 ( .A1(n10114), .A2(n10115), .ZN(n10094) );
  AND2_X1 U9960 ( .A1(n10088), .A2(n10091), .ZN(n10115) );
  AND2_X1 U9961 ( .A1(n10116), .A2(n10090), .ZN(n10114) );
  OR2_X1 U9962 ( .A1(n10117), .A2(n10118), .ZN(n10090) );
  AND2_X1 U9963 ( .A1(n10084), .A2(n10087), .ZN(n10118) );
  AND2_X1 U9964 ( .A1(n10119), .A2(n10086), .ZN(n10117) );
  OR2_X1 U9965 ( .A1(n10120), .A2(n10121), .ZN(n10086) );
  AND2_X1 U9966 ( .A1(n10080), .A2(n10083), .ZN(n10121) );
  AND2_X1 U9967 ( .A1(n10122), .A2(n10082), .ZN(n10120) );
  OR2_X1 U9968 ( .A1(n10123), .A2(n10124), .ZN(n10082) );
  AND2_X1 U9969 ( .A1(n10076), .A2(n10079), .ZN(n10124) );
  AND2_X1 U9970 ( .A1(n10125), .A2(n10078), .ZN(n10123) );
  OR2_X1 U9971 ( .A1(n10126), .A2(n10127), .ZN(n10078) );
  AND2_X1 U9972 ( .A1(n10072), .A2(n10075), .ZN(n10127) );
  AND2_X1 U9973 ( .A1(n10128), .A2(n10074), .ZN(n10126) );
  OR2_X1 U9974 ( .A1(n10129), .A2(n10130), .ZN(n10074) );
  AND2_X1 U9975 ( .A1(n10068), .A2(n10071), .ZN(n10130) );
  AND2_X1 U9976 ( .A1(n10131), .A2(n10070), .ZN(n10129) );
  OR2_X1 U9977 ( .A1(n10132), .A2(n10133), .ZN(n10070) );
  AND2_X1 U9978 ( .A1(n10064), .A2(n10067), .ZN(n10133) );
  AND2_X1 U9979 ( .A1(n10134), .A2(n10066), .ZN(n10132) );
  OR2_X1 U9980 ( .A1(n10135), .A2(n10136), .ZN(n10066) );
  AND2_X1 U9981 ( .A1(n10060), .A2(n10063), .ZN(n10136) );
  AND2_X1 U9982 ( .A1(n10137), .A2(n10062), .ZN(n10135) );
  OR2_X1 U9983 ( .A1(n10138), .A2(n10139), .ZN(n10062) );
  AND2_X1 U9984 ( .A1(n10056), .A2(n10059), .ZN(n10139) );
  AND2_X1 U9985 ( .A1(n10140), .A2(n10058), .ZN(n10138) );
  OR2_X1 U9986 ( .A1(n10141), .A2(n10142), .ZN(n10058) );
  AND2_X1 U9987 ( .A1(n10052), .A2(n10055), .ZN(n10142) );
  AND2_X1 U9988 ( .A1(n10143), .A2(n10054), .ZN(n10141) );
  OR2_X1 U9989 ( .A1(n10144), .A2(n10145), .ZN(n10054) );
  AND2_X1 U9990 ( .A1(n10048), .A2(n10051), .ZN(n10145) );
  AND2_X1 U9991 ( .A1(n10146), .A2(n10050), .ZN(n10144) );
  OR2_X1 U9992 ( .A1(n10147), .A2(n10148), .ZN(n10050) );
  AND2_X1 U9993 ( .A1(n10044), .A2(n10047), .ZN(n10148) );
  AND2_X1 U9994 ( .A1(n10149), .A2(n10046), .ZN(n10147) );
  OR2_X1 U9995 ( .A1(n10150), .A2(n10151), .ZN(n10046) );
  AND2_X1 U9996 ( .A1(n10040), .A2(n10043), .ZN(n10151) );
  AND2_X1 U9997 ( .A1(n10152), .A2(n10042), .ZN(n10150) );
  OR2_X1 U9998 ( .A1(n10153), .A2(n10154), .ZN(n10042) );
  AND2_X1 U9999 ( .A1(n10036), .A2(n10039), .ZN(n10154) );
  AND2_X1 U10000 ( .A1(n10155), .A2(n10038), .ZN(n10153) );
  OR2_X1 U10001 ( .A1(n10156), .A2(n10157), .ZN(n10038) );
  AND2_X1 U10002 ( .A1(n10032), .A2(n10035), .ZN(n10157) );
  AND2_X1 U10003 ( .A1(n10158), .A2(n10034), .ZN(n10156) );
  OR2_X1 U10004 ( .A1(n10159), .A2(n10160), .ZN(n10034) );
  AND2_X1 U10005 ( .A1(n10028), .A2(n10031), .ZN(n10160) );
  AND2_X1 U10006 ( .A1(n10161), .A2(n10030), .ZN(n10159) );
  OR2_X1 U10007 ( .A1(n10162), .A2(n10163), .ZN(n10030) );
  AND2_X1 U10008 ( .A1(n10024), .A2(n10027), .ZN(n10163) );
  AND2_X1 U10009 ( .A1(n10164), .A2(n10026), .ZN(n10162) );
  OR2_X1 U10010 ( .A1(n10165), .A2(n10166), .ZN(n10026) );
  AND2_X1 U10011 ( .A1(n10020), .A2(n10023), .ZN(n10166) );
  AND2_X1 U10012 ( .A1(n10167), .A2(n10022), .ZN(n10165) );
  OR2_X1 U10013 ( .A1(n10168), .A2(n10169), .ZN(n10022) );
  AND2_X1 U10014 ( .A1(n10016), .A2(n10019), .ZN(n10169) );
  AND2_X1 U10015 ( .A1(n10170), .A2(n10018), .ZN(n10168) );
  OR2_X1 U10016 ( .A1(n10171), .A2(n10172), .ZN(n10018) );
  AND2_X1 U10017 ( .A1(n10012), .A2(n10015), .ZN(n10172) );
  AND2_X1 U10018 ( .A1(n10173), .A2(n10014), .ZN(n10171) );
  OR2_X1 U10019 ( .A1(n10174), .A2(n10175), .ZN(n10014) );
  AND2_X1 U10020 ( .A1(n10008), .A2(n10011), .ZN(n10175) );
  AND2_X1 U10021 ( .A1(n10176), .A2(n10010), .ZN(n10174) );
  OR2_X1 U10022 ( .A1(n10177), .A2(n10178), .ZN(n10010) );
  AND2_X1 U10023 ( .A1(n10004), .A2(n10007), .ZN(n10178) );
  AND2_X1 U10024 ( .A1(n10179), .A2(n10006), .ZN(n10177) );
  OR2_X1 U10025 ( .A1(n10180), .A2(n10181), .ZN(n10006) );
  AND2_X1 U10026 ( .A1(n10001), .A2(n10002), .ZN(n10181) );
  AND2_X1 U10027 ( .A1(n10182), .A2(n10003), .ZN(n10180) );
  OR2_X1 U10028 ( .A1(n10183), .A2(n10184), .ZN(n10003) );
  AND2_X1 U10029 ( .A1(n9996), .A2(n9999), .ZN(n10184) );
  AND2_X1 U10030 ( .A1(n10185), .A2(n9998), .ZN(n10183) );
  OR2_X1 U10031 ( .A1(n10186), .A2(n10187), .ZN(n9998) );
  AND2_X1 U10032 ( .A1(n9993), .A2(n9994), .ZN(n10187) );
  AND2_X1 U10033 ( .A1(n10188), .A2(n10189), .ZN(n10186) );
  OR2_X1 U10034 ( .A1(n9994), .A2(n9993), .ZN(n10189) );
  OR2_X1 U10035 ( .A1(n9014), .A2(n7998), .ZN(n9993) );
  OR2_X1 U10036 ( .A1(n9984), .A2(n10190), .ZN(n9994) );
  OR2_X1 U10037 ( .A1(n7998), .A2(n8047), .ZN(n10190) );
  INV_X1 U10038 ( .A(n9995), .ZN(n10188) );
  OR2_X1 U10039 ( .A1(n10191), .A2(n10192), .ZN(n9995) );
  AND2_X1 U10040 ( .A1(b_29_), .A2(n10193), .ZN(n10192) );
  OR2_X1 U10041 ( .A1(n10194), .A2(n9989), .ZN(n10193) );
  AND2_X1 U10042 ( .A1(a_30_), .A2(n8075), .ZN(n10194) );
  AND2_X1 U10043 ( .A1(b_28_), .A2(n10195), .ZN(n10191) );
  OR2_X1 U10044 ( .A1(n10196), .A2(n8021), .ZN(n10195) );
  AND2_X1 U10045 ( .A1(a_31_), .A2(n8047), .ZN(n10196) );
  OR2_X1 U10046 ( .A1(n9999), .A2(n9996), .ZN(n10185) );
  XOR2_X1 U10047 ( .A(n10197), .B(n9015), .Z(n9996) );
  XNOR2_X1 U10048 ( .A(n10198), .B(n10199), .ZN(n10197) );
  OR2_X1 U10049 ( .A1(n9010), .A2(n7998), .ZN(n9999) );
  OR2_X1 U10050 ( .A1(n10002), .A2(n10001), .ZN(n10182) );
  XOR2_X1 U10051 ( .A(n10200), .B(n10201), .Z(n10001) );
  XOR2_X1 U10052 ( .A(n10202), .B(n10203), .Z(n10201) );
  OR2_X1 U10053 ( .A1(n9006), .A2(n7998), .ZN(n10002) );
  OR2_X1 U10054 ( .A1(n10007), .A2(n10004), .ZN(n10179) );
  XOR2_X1 U10055 ( .A(n10204), .B(n10205), .Z(n10004) );
  XOR2_X1 U10056 ( .A(n10206), .B(n10207), .Z(n10205) );
  OR2_X1 U10057 ( .A1(n9002), .A2(n7998), .ZN(n10007) );
  OR2_X1 U10058 ( .A1(n10011), .A2(n10008), .ZN(n10176) );
  XOR2_X1 U10059 ( .A(n10208), .B(n10209), .Z(n10008) );
  XOR2_X1 U10060 ( .A(n10210), .B(n10211), .Z(n10209) );
  OR2_X1 U10061 ( .A1(n8998), .A2(n7998), .ZN(n10011) );
  OR2_X1 U10062 ( .A1(n10015), .A2(n10012), .ZN(n10173) );
  XOR2_X1 U10063 ( .A(n10212), .B(n10213), .Z(n10012) );
  XOR2_X1 U10064 ( .A(n10214), .B(n10215), .Z(n10213) );
  OR2_X1 U10065 ( .A1(n8994), .A2(n7998), .ZN(n10015) );
  OR2_X1 U10066 ( .A1(n10019), .A2(n10016), .ZN(n10170) );
  XOR2_X1 U10067 ( .A(n10216), .B(n10217), .Z(n10016) );
  XOR2_X1 U10068 ( .A(n10218), .B(n10219), .Z(n10217) );
  OR2_X1 U10069 ( .A1(n8990), .A2(n7998), .ZN(n10019) );
  OR2_X1 U10070 ( .A1(n10023), .A2(n10020), .ZN(n10167) );
  XOR2_X1 U10071 ( .A(n10220), .B(n10221), .Z(n10020) );
  XOR2_X1 U10072 ( .A(n10222), .B(n10223), .Z(n10221) );
  OR2_X1 U10073 ( .A1(n8986), .A2(n7998), .ZN(n10023) );
  OR2_X1 U10074 ( .A1(n10027), .A2(n10024), .ZN(n10164) );
  XOR2_X1 U10075 ( .A(n10224), .B(n10225), .Z(n10024) );
  XOR2_X1 U10076 ( .A(n10226), .B(n10227), .Z(n10225) );
  OR2_X1 U10077 ( .A1(n8982), .A2(n7998), .ZN(n10027) );
  OR2_X1 U10078 ( .A1(n10031), .A2(n10028), .ZN(n10161) );
  XOR2_X1 U10079 ( .A(n10228), .B(n10229), .Z(n10028) );
  XOR2_X1 U10080 ( .A(n10230), .B(n10231), .Z(n10229) );
  OR2_X1 U10081 ( .A1(n8978), .A2(n7998), .ZN(n10031) );
  OR2_X1 U10082 ( .A1(n10035), .A2(n10032), .ZN(n10158) );
  XOR2_X1 U10083 ( .A(n10232), .B(n10233), .Z(n10032) );
  XOR2_X1 U10084 ( .A(n10234), .B(n10235), .Z(n10233) );
  OR2_X1 U10085 ( .A1(n8974), .A2(n7998), .ZN(n10035) );
  OR2_X1 U10086 ( .A1(n10039), .A2(n10036), .ZN(n10155) );
  XOR2_X1 U10087 ( .A(n10236), .B(n10237), .Z(n10036) );
  XOR2_X1 U10088 ( .A(n10238), .B(n10239), .Z(n10237) );
  OR2_X1 U10089 ( .A1(n8970), .A2(n7998), .ZN(n10039) );
  OR2_X1 U10090 ( .A1(n10043), .A2(n10040), .ZN(n10152) );
  XOR2_X1 U10091 ( .A(n10240), .B(n10241), .Z(n10040) );
  XOR2_X1 U10092 ( .A(n10242), .B(n10243), .Z(n10241) );
  OR2_X1 U10093 ( .A1(n8966), .A2(n7998), .ZN(n10043) );
  OR2_X1 U10094 ( .A1(n10047), .A2(n10044), .ZN(n10149) );
  XOR2_X1 U10095 ( .A(n10244), .B(n10245), .Z(n10044) );
  XOR2_X1 U10096 ( .A(n10246), .B(n10247), .Z(n10245) );
  OR2_X1 U10097 ( .A1(n8962), .A2(n7998), .ZN(n10047) );
  OR2_X1 U10098 ( .A1(n10051), .A2(n10048), .ZN(n10146) );
  XOR2_X1 U10099 ( .A(n10248), .B(n10249), .Z(n10048) );
  XOR2_X1 U10100 ( .A(n10250), .B(n10251), .Z(n10249) );
  OR2_X1 U10101 ( .A1(n8958), .A2(n7998), .ZN(n10051) );
  OR2_X1 U10102 ( .A1(n10055), .A2(n10052), .ZN(n10143) );
  XOR2_X1 U10103 ( .A(n10252), .B(n10253), .Z(n10052) );
  XOR2_X1 U10104 ( .A(n10254), .B(n10255), .Z(n10253) );
  OR2_X1 U10105 ( .A1(n8954), .A2(n7998), .ZN(n10055) );
  OR2_X1 U10106 ( .A1(n10059), .A2(n10056), .ZN(n10140) );
  XOR2_X1 U10107 ( .A(n10256), .B(n10257), .Z(n10056) );
  XOR2_X1 U10108 ( .A(n10258), .B(n10259), .Z(n10257) );
  OR2_X1 U10109 ( .A1(n8950), .A2(n7998), .ZN(n10059) );
  OR2_X1 U10110 ( .A1(n10063), .A2(n10060), .ZN(n10137) );
  XOR2_X1 U10111 ( .A(n10260), .B(n10261), .Z(n10060) );
  XOR2_X1 U10112 ( .A(n10262), .B(n10263), .Z(n10261) );
  OR2_X1 U10113 ( .A1(n8946), .A2(n7998), .ZN(n10063) );
  OR2_X1 U10114 ( .A1(n10067), .A2(n10064), .ZN(n10134) );
  XOR2_X1 U10115 ( .A(n10264), .B(n10265), .Z(n10064) );
  XOR2_X1 U10116 ( .A(n10266), .B(n10267), .Z(n10265) );
  OR2_X1 U10117 ( .A1(n8942), .A2(n7998), .ZN(n10067) );
  OR2_X1 U10118 ( .A1(n10071), .A2(n10068), .ZN(n10131) );
  XOR2_X1 U10119 ( .A(n10268), .B(n10269), .Z(n10068) );
  XOR2_X1 U10120 ( .A(n10270), .B(n10271), .Z(n10269) );
  OR2_X1 U10121 ( .A1(n8938), .A2(n7998), .ZN(n10071) );
  OR2_X1 U10122 ( .A1(n10075), .A2(n10072), .ZN(n10128) );
  XOR2_X1 U10123 ( .A(n10272), .B(n10273), .Z(n10072) );
  XOR2_X1 U10124 ( .A(n10274), .B(n10275), .Z(n10273) );
  OR2_X1 U10125 ( .A1(n8934), .A2(n7998), .ZN(n10075) );
  OR2_X1 U10126 ( .A1(n10079), .A2(n10076), .ZN(n10125) );
  XOR2_X1 U10127 ( .A(n10276), .B(n10277), .Z(n10076) );
  XOR2_X1 U10128 ( .A(n10278), .B(n10279), .Z(n10277) );
  OR2_X1 U10129 ( .A1(n8930), .A2(n7998), .ZN(n10079) );
  OR2_X1 U10130 ( .A1(n10083), .A2(n10080), .ZN(n10122) );
  XOR2_X1 U10131 ( .A(n10280), .B(n10281), .Z(n10080) );
  XOR2_X1 U10132 ( .A(n10282), .B(n10283), .Z(n10281) );
  OR2_X1 U10133 ( .A1(n8926), .A2(n7998), .ZN(n10083) );
  OR2_X1 U10134 ( .A1(n10087), .A2(n10084), .ZN(n10119) );
  XOR2_X1 U10135 ( .A(n10284), .B(n10285), .Z(n10084) );
  XOR2_X1 U10136 ( .A(n10286), .B(n10287), .Z(n10285) );
  OR2_X1 U10137 ( .A1(n8922), .A2(n7998), .ZN(n10087) );
  OR2_X1 U10138 ( .A1(n10091), .A2(n10088), .ZN(n10116) );
  XOR2_X1 U10139 ( .A(n10288), .B(n10289), .Z(n10088) );
  XOR2_X1 U10140 ( .A(n10290), .B(n10291), .Z(n10289) );
  OR2_X1 U10141 ( .A1(n8918), .A2(n7998), .ZN(n10091) );
  OR2_X1 U10142 ( .A1(n10095), .A2(n10092), .ZN(n10113) );
  XOR2_X1 U10143 ( .A(n10292), .B(n10293), .Z(n10092) );
  XOR2_X1 U10144 ( .A(n10294), .B(n10295), .Z(n10293) );
  OR2_X1 U10145 ( .A1(n8914), .A2(n7998), .ZN(n10095) );
  OR2_X1 U10146 ( .A1(n10099), .A2(n10096), .ZN(n10110) );
  XOR2_X1 U10147 ( .A(n10296), .B(n10297), .Z(n10096) );
  XOR2_X1 U10148 ( .A(n10298), .B(n10299), .Z(n10297) );
  OR2_X1 U10149 ( .A1(n8910), .A2(n7998), .ZN(n10099) );
  OR2_X1 U10150 ( .A1(n10103), .A2(n10100), .ZN(n10107) );
  XOR2_X1 U10151 ( .A(n10300), .B(n10301), .Z(n10100) );
  XOR2_X1 U10152 ( .A(n10302), .B(n10303), .Z(n10301) );
  OR2_X1 U10153 ( .A1(n8906), .A2(n7998), .ZN(n10103) );
  XNOR2_X1 U10154 ( .A(n10304), .B(n10305), .ZN(n9885) );
  XNOR2_X1 U10155 ( .A(n10306), .B(n10307), .ZN(n10304) );
  OR2_X1 U10156 ( .A1(n10308), .A2(n10309), .ZN(n9055) );
  XNOR2_X1 U10157 ( .A(n10310), .B(n9859), .ZN(n10309) );
  AND2_X1 U10158 ( .A1(n9870), .A2(n9861), .ZN(n10308) );
  XNOR2_X1 U10159 ( .A(n10311), .B(n10312), .ZN(n9861) );
  XOR2_X1 U10160 ( .A(n10313), .B(n10314), .Z(n10312) );
  INV_X1 U10161 ( .A(n9855), .ZN(n9870) );
  OR2_X1 U10162 ( .A1(n10315), .A2(n10316), .ZN(n9855) );
  AND2_X1 U10163 ( .A1(n9881), .A2(n9880), .ZN(n10316) );
  AND2_X1 U10164 ( .A1(n9878), .A2(n10317), .ZN(n10315) );
  OR2_X1 U10165 ( .A1(n9880), .A2(n9881), .ZN(n10317) );
  OR2_X1 U10166 ( .A1(n9297), .A2(n8047), .ZN(n9881) );
  OR2_X1 U10167 ( .A1(n10318), .A2(n10319), .ZN(n9880) );
  AND2_X1 U10168 ( .A1(n9892), .A2(n9891), .ZN(n10319) );
  AND2_X1 U10169 ( .A1(n9889), .A2(n10320), .ZN(n10318) );
  OR2_X1 U10170 ( .A1(n9891), .A2(n9892), .ZN(n10320) );
  OR2_X1 U10171 ( .A1(n8902), .A2(n8047), .ZN(n9892) );
  OR2_X1 U10172 ( .A1(n10321), .A2(n10322), .ZN(n9891) );
  AND2_X1 U10173 ( .A1(n10307), .A2(n10306), .ZN(n10322) );
  AND2_X1 U10174 ( .A1(n10305), .A2(n10323), .ZN(n10321) );
  OR2_X1 U10175 ( .A1(n10306), .A2(n10307), .ZN(n10323) );
  OR2_X1 U10176 ( .A1(n10324), .A2(n10325), .ZN(n10307) );
  AND2_X1 U10177 ( .A1(n10303), .A2(n10302), .ZN(n10325) );
  AND2_X1 U10178 ( .A1(n10300), .A2(n10326), .ZN(n10324) );
  OR2_X1 U10179 ( .A1(n10302), .A2(n10303), .ZN(n10326) );
  OR2_X1 U10180 ( .A1(n8910), .A2(n8047), .ZN(n10303) );
  OR2_X1 U10181 ( .A1(n10327), .A2(n10328), .ZN(n10302) );
  AND2_X1 U10182 ( .A1(n10299), .A2(n10298), .ZN(n10328) );
  AND2_X1 U10183 ( .A1(n10296), .A2(n10329), .ZN(n10327) );
  OR2_X1 U10184 ( .A1(n10298), .A2(n10299), .ZN(n10329) );
  OR2_X1 U10185 ( .A1(n8914), .A2(n8047), .ZN(n10299) );
  OR2_X1 U10186 ( .A1(n10330), .A2(n10331), .ZN(n10298) );
  AND2_X1 U10187 ( .A1(n10295), .A2(n10294), .ZN(n10331) );
  AND2_X1 U10188 ( .A1(n10292), .A2(n10332), .ZN(n10330) );
  OR2_X1 U10189 ( .A1(n10294), .A2(n10295), .ZN(n10332) );
  OR2_X1 U10190 ( .A1(n8918), .A2(n8047), .ZN(n10295) );
  OR2_X1 U10191 ( .A1(n10333), .A2(n10334), .ZN(n10294) );
  AND2_X1 U10192 ( .A1(n10291), .A2(n10290), .ZN(n10334) );
  AND2_X1 U10193 ( .A1(n10288), .A2(n10335), .ZN(n10333) );
  OR2_X1 U10194 ( .A1(n10290), .A2(n10291), .ZN(n10335) );
  OR2_X1 U10195 ( .A1(n8922), .A2(n8047), .ZN(n10291) );
  OR2_X1 U10196 ( .A1(n10336), .A2(n10337), .ZN(n10290) );
  AND2_X1 U10197 ( .A1(n10287), .A2(n10286), .ZN(n10337) );
  AND2_X1 U10198 ( .A1(n10284), .A2(n10338), .ZN(n10336) );
  OR2_X1 U10199 ( .A1(n10286), .A2(n10287), .ZN(n10338) );
  OR2_X1 U10200 ( .A1(n8926), .A2(n8047), .ZN(n10287) );
  OR2_X1 U10201 ( .A1(n10339), .A2(n10340), .ZN(n10286) );
  AND2_X1 U10202 ( .A1(n10283), .A2(n10282), .ZN(n10340) );
  AND2_X1 U10203 ( .A1(n10280), .A2(n10341), .ZN(n10339) );
  OR2_X1 U10204 ( .A1(n10282), .A2(n10283), .ZN(n10341) );
  OR2_X1 U10205 ( .A1(n8930), .A2(n8047), .ZN(n10283) );
  OR2_X1 U10206 ( .A1(n10342), .A2(n10343), .ZN(n10282) );
  AND2_X1 U10207 ( .A1(n10279), .A2(n10278), .ZN(n10343) );
  AND2_X1 U10208 ( .A1(n10276), .A2(n10344), .ZN(n10342) );
  OR2_X1 U10209 ( .A1(n10278), .A2(n10279), .ZN(n10344) );
  OR2_X1 U10210 ( .A1(n8934), .A2(n8047), .ZN(n10279) );
  OR2_X1 U10211 ( .A1(n10345), .A2(n10346), .ZN(n10278) );
  AND2_X1 U10212 ( .A1(n10275), .A2(n10274), .ZN(n10346) );
  AND2_X1 U10213 ( .A1(n10272), .A2(n10347), .ZN(n10345) );
  OR2_X1 U10214 ( .A1(n10274), .A2(n10275), .ZN(n10347) );
  OR2_X1 U10215 ( .A1(n8938), .A2(n8047), .ZN(n10275) );
  OR2_X1 U10216 ( .A1(n10348), .A2(n10349), .ZN(n10274) );
  AND2_X1 U10217 ( .A1(n10271), .A2(n10270), .ZN(n10349) );
  AND2_X1 U10218 ( .A1(n10268), .A2(n10350), .ZN(n10348) );
  OR2_X1 U10219 ( .A1(n10270), .A2(n10271), .ZN(n10350) );
  OR2_X1 U10220 ( .A1(n8942), .A2(n8047), .ZN(n10271) );
  OR2_X1 U10221 ( .A1(n10351), .A2(n10352), .ZN(n10270) );
  AND2_X1 U10222 ( .A1(n10267), .A2(n10266), .ZN(n10352) );
  AND2_X1 U10223 ( .A1(n10264), .A2(n10353), .ZN(n10351) );
  OR2_X1 U10224 ( .A1(n10266), .A2(n10267), .ZN(n10353) );
  OR2_X1 U10225 ( .A1(n8946), .A2(n8047), .ZN(n10267) );
  OR2_X1 U10226 ( .A1(n10354), .A2(n10355), .ZN(n10266) );
  AND2_X1 U10227 ( .A1(n10263), .A2(n10262), .ZN(n10355) );
  AND2_X1 U10228 ( .A1(n10260), .A2(n10356), .ZN(n10354) );
  OR2_X1 U10229 ( .A1(n10262), .A2(n10263), .ZN(n10356) );
  OR2_X1 U10230 ( .A1(n8950), .A2(n8047), .ZN(n10263) );
  OR2_X1 U10231 ( .A1(n10357), .A2(n10358), .ZN(n10262) );
  AND2_X1 U10232 ( .A1(n10259), .A2(n10258), .ZN(n10358) );
  AND2_X1 U10233 ( .A1(n10256), .A2(n10359), .ZN(n10357) );
  OR2_X1 U10234 ( .A1(n10258), .A2(n10259), .ZN(n10359) );
  OR2_X1 U10235 ( .A1(n8954), .A2(n8047), .ZN(n10259) );
  OR2_X1 U10236 ( .A1(n10360), .A2(n10361), .ZN(n10258) );
  AND2_X1 U10237 ( .A1(n10255), .A2(n10254), .ZN(n10361) );
  AND2_X1 U10238 ( .A1(n10252), .A2(n10362), .ZN(n10360) );
  OR2_X1 U10239 ( .A1(n10254), .A2(n10255), .ZN(n10362) );
  OR2_X1 U10240 ( .A1(n8958), .A2(n8047), .ZN(n10255) );
  OR2_X1 U10241 ( .A1(n10363), .A2(n10364), .ZN(n10254) );
  AND2_X1 U10242 ( .A1(n10251), .A2(n10250), .ZN(n10364) );
  AND2_X1 U10243 ( .A1(n10248), .A2(n10365), .ZN(n10363) );
  OR2_X1 U10244 ( .A1(n10250), .A2(n10251), .ZN(n10365) );
  OR2_X1 U10245 ( .A1(n8962), .A2(n8047), .ZN(n10251) );
  OR2_X1 U10246 ( .A1(n10366), .A2(n10367), .ZN(n10250) );
  AND2_X1 U10247 ( .A1(n10247), .A2(n10246), .ZN(n10367) );
  AND2_X1 U10248 ( .A1(n10244), .A2(n10368), .ZN(n10366) );
  OR2_X1 U10249 ( .A1(n10246), .A2(n10247), .ZN(n10368) );
  OR2_X1 U10250 ( .A1(n8966), .A2(n8047), .ZN(n10247) );
  OR2_X1 U10251 ( .A1(n10369), .A2(n10370), .ZN(n10246) );
  AND2_X1 U10252 ( .A1(n10243), .A2(n10242), .ZN(n10370) );
  AND2_X1 U10253 ( .A1(n10240), .A2(n10371), .ZN(n10369) );
  OR2_X1 U10254 ( .A1(n10242), .A2(n10243), .ZN(n10371) );
  OR2_X1 U10255 ( .A1(n8970), .A2(n8047), .ZN(n10243) );
  OR2_X1 U10256 ( .A1(n10372), .A2(n10373), .ZN(n10242) );
  AND2_X1 U10257 ( .A1(n10239), .A2(n10238), .ZN(n10373) );
  AND2_X1 U10258 ( .A1(n10236), .A2(n10374), .ZN(n10372) );
  OR2_X1 U10259 ( .A1(n10238), .A2(n10239), .ZN(n10374) );
  OR2_X1 U10260 ( .A1(n8974), .A2(n8047), .ZN(n10239) );
  OR2_X1 U10261 ( .A1(n10375), .A2(n10376), .ZN(n10238) );
  AND2_X1 U10262 ( .A1(n10235), .A2(n10234), .ZN(n10376) );
  AND2_X1 U10263 ( .A1(n10232), .A2(n10377), .ZN(n10375) );
  OR2_X1 U10264 ( .A1(n10234), .A2(n10235), .ZN(n10377) );
  OR2_X1 U10265 ( .A1(n8978), .A2(n8047), .ZN(n10235) );
  OR2_X1 U10266 ( .A1(n10378), .A2(n10379), .ZN(n10234) );
  AND2_X1 U10267 ( .A1(n10231), .A2(n10230), .ZN(n10379) );
  AND2_X1 U10268 ( .A1(n10228), .A2(n10380), .ZN(n10378) );
  OR2_X1 U10269 ( .A1(n10230), .A2(n10231), .ZN(n10380) );
  OR2_X1 U10270 ( .A1(n8982), .A2(n8047), .ZN(n10231) );
  OR2_X1 U10271 ( .A1(n10381), .A2(n10382), .ZN(n10230) );
  AND2_X1 U10272 ( .A1(n10227), .A2(n10226), .ZN(n10382) );
  AND2_X1 U10273 ( .A1(n10224), .A2(n10383), .ZN(n10381) );
  OR2_X1 U10274 ( .A1(n10226), .A2(n10227), .ZN(n10383) );
  OR2_X1 U10275 ( .A1(n8986), .A2(n8047), .ZN(n10227) );
  OR2_X1 U10276 ( .A1(n10384), .A2(n10385), .ZN(n10226) );
  AND2_X1 U10277 ( .A1(n10223), .A2(n10222), .ZN(n10385) );
  AND2_X1 U10278 ( .A1(n10220), .A2(n10386), .ZN(n10384) );
  OR2_X1 U10279 ( .A1(n10222), .A2(n10223), .ZN(n10386) );
  OR2_X1 U10280 ( .A1(n8990), .A2(n8047), .ZN(n10223) );
  OR2_X1 U10281 ( .A1(n10387), .A2(n10388), .ZN(n10222) );
  AND2_X1 U10282 ( .A1(n10219), .A2(n10218), .ZN(n10388) );
  AND2_X1 U10283 ( .A1(n10216), .A2(n10389), .ZN(n10387) );
  OR2_X1 U10284 ( .A1(n10218), .A2(n10219), .ZN(n10389) );
  OR2_X1 U10285 ( .A1(n8994), .A2(n8047), .ZN(n10219) );
  OR2_X1 U10286 ( .A1(n10390), .A2(n10391), .ZN(n10218) );
  AND2_X1 U10287 ( .A1(n10215), .A2(n10214), .ZN(n10391) );
  AND2_X1 U10288 ( .A1(n10212), .A2(n10392), .ZN(n10390) );
  OR2_X1 U10289 ( .A1(n10214), .A2(n10215), .ZN(n10392) );
  OR2_X1 U10290 ( .A1(n8998), .A2(n8047), .ZN(n10215) );
  OR2_X1 U10291 ( .A1(n10393), .A2(n10394), .ZN(n10214) );
  AND2_X1 U10292 ( .A1(n10211), .A2(n10210), .ZN(n10394) );
  AND2_X1 U10293 ( .A1(n10208), .A2(n10395), .ZN(n10393) );
  OR2_X1 U10294 ( .A1(n10210), .A2(n10211), .ZN(n10395) );
  OR2_X1 U10295 ( .A1(n9002), .A2(n8047), .ZN(n10211) );
  OR2_X1 U10296 ( .A1(n10396), .A2(n10397), .ZN(n10210) );
  AND2_X1 U10297 ( .A1(n10207), .A2(n10206), .ZN(n10397) );
  AND2_X1 U10298 ( .A1(n10204), .A2(n10398), .ZN(n10396) );
  OR2_X1 U10299 ( .A1(n10206), .A2(n10207), .ZN(n10398) );
  OR2_X1 U10300 ( .A1(n9006), .A2(n8047), .ZN(n10207) );
  OR2_X1 U10301 ( .A1(n10399), .A2(n10400), .ZN(n10206) );
  AND2_X1 U10302 ( .A1(n10203), .A2(n10202), .ZN(n10400) );
  AND2_X1 U10303 ( .A1(n10200), .A2(n10401), .ZN(n10399) );
  OR2_X1 U10304 ( .A1(n10202), .A2(n10203), .ZN(n10401) );
  OR2_X1 U10305 ( .A1(n9010), .A2(n8047), .ZN(n10203) );
  OR2_X1 U10306 ( .A1(n10402), .A2(n10403), .ZN(n10202) );
  AND2_X1 U10307 ( .A1(n9015), .A2(n10198), .ZN(n10403) );
  AND2_X1 U10308 ( .A1(n10404), .A2(n10405), .ZN(n10402) );
  OR2_X1 U10309 ( .A1(n10198), .A2(n9015), .ZN(n10405) );
  OR2_X1 U10310 ( .A1(n9014), .A2(n8047), .ZN(n9015) );
  OR2_X1 U10311 ( .A1(n9984), .A2(n10406), .ZN(n10198) );
  OR2_X1 U10312 ( .A1(n8047), .A2(n8075), .ZN(n10406) );
  INV_X1 U10313 ( .A(n10199), .ZN(n10404) );
  OR2_X1 U10314 ( .A1(n10407), .A2(n10408), .ZN(n10199) );
  AND2_X1 U10315 ( .A1(b_28_), .A2(n10409), .ZN(n10408) );
  OR2_X1 U10316 ( .A1(n10410), .A2(n9989), .ZN(n10409) );
  AND2_X1 U10317 ( .A1(a_30_), .A2(n8112), .ZN(n10410) );
  AND2_X1 U10318 ( .A1(b_27_), .A2(n10411), .ZN(n10407) );
  OR2_X1 U10319 ( .A1(n10412), .A2(n8021), .ZN(n10411) );
  AND2_X1 U10320 ( .A1(a_31_), .A2(n8075), .ZN(n10412) );
  XOR2_X1 U10321 ( .A(n10413), .B(n10414), .Z(n10200) );
  XNOR2_X1 U10322 ( .A(n10415), .B(n10416), .ZN(n10413) );
  XOR2_X1 U10323 ( .A(n10417), .B(n10418), .Z(n10204) );
  XOR2_X1 U10324 ( .A(n10419), .B(n9011), .Z(n10418) );
  XOR2_X1 U10325 ( .A(n10420), .B(n10421), .Z(n10208) );
  XOR2_X1 U10326 ( .A(n10422), .B(n10423), .Z(n10421) );
  XOR2_X1 U10327 ( .A(n10424), .B(n10425), .Z(n10212) );
  XOR2_X1 U10328 ( .A(n10426), .B(n10427), .Z(n10425) );
  XOR2_X1 U10329 ( .A(n10428), .B(n10429), .Z(n10216) );
  XOR2_X1 U10330 ( .A(n10430), .B(n10431), .Z(n10429) );
  XOR2_X1 U10331 ( .A(n10432), .B(n10433), .Z(n10220) );
  XOR2_X1 U10332 ( .A(n10434), .B(n10435), .Z(n10433) );
  XOR2_X1 U10333 ( .A(n10436), .B(n10437), .Z(n10224) );
  XOR2_X1 U10334 ( .A(n10438), .B(n10439), .Z(n10437) );
  XOR2_X1 U10335 ( .A(n10440), .B(n10441), .Z(n10228) );
  XOR2_X1 U10336 ( .A(n10442), .B(n10443), .Z(n10441) );
  XOR2_X1 U10337 ( .A(n10444), .B(n10445), .Z(n10232) );
  XOR2_X1 U10338 ( .A(n10446), .B(n10447), .Z(n10445) );
  XOR2_X1 U10339 ( .A(n10448), .B(n10449), .Z(n10236) );
  XOR2_X1 U10340 ( .A(n10450), .B(n10451), .Z(n10449) );
  XOR2_X1 U10341 ( .A(n10452), .B(n10453), .Z(n10240) );
  XOR2_X1 U10342 ( .A(n10454), .B(n10455), .Z(n10453) );
  XOR2_X1 U10343 ( .A(n10456), .B(n10457), .Z(n10244) );
  XOR2_X1 U10344 ( .A(n10458), .B(n10459), .Z(n10457) );
  XOR2_X1 U10345 ( .A(n10460), .B(n10461), .Z(n10248) );
  XOR2_X1 U10346 ( .A(n10462), .B(n10463), .Z(n10461) );
  XOR2_X1 U10347 ( .A(n10464), .B(n10465), .Z(n10252) );
  XOR2_X1 U10348 ( .A(n10466), .B(n10467), .Z(n10465) );
  XOR2_X1 U10349 ( .A(n10468), .B(n10469), .Z(n10256) );
  XOR2_X1 U10350 ( .A(n10470), .B(n10471), .Z(n10469) );
  XOR2_X1 U10351 ( .A(n10472), .B(n10473), .Z(n10260) );
  XOR2_X1 U10352 ( .A(n10474), .B(n10475), .Z(n10473) );
  XOR2_X1 U10353 ( .A(n10476), .B(n10477), .Z(n10264) );
  XOR2_X1 U10354 ( .A(n10478), .B(n10479), .Z(n10477) );
  XOR2_X1 U10355 ( .A(n10480), .B(n10481), .Z(n10268) );
  XOR2_X1 U10356 ( .A(n10482), .B(n10483), .Z(n10481) );
  XOR2_X1 U10357 ( .A(n10484), .B(n10485), .Z(n10272) );
  XOR2_X1 U10358 ( .A(n10486), .B(n10487), .Z(n10485) );
  XOR2_X1 U10359 ( .A(n10488), .B(n10489), .Z(n10276) );
  XOR2_X1 U10360 ( .A(n10490), .B(n10491), .Z(n10489) );
  XOR2_X1 U10361 ( .A(n10492), .B(n10493), .Z(n10280) );
  XOR2_X1 U10362 ( .A(n10494), .B(n10495), .Z(n10493) );
  XOR2_X1 U10363 ( .A(n10496), .B(n10497), .Z(n10284) );
  XOR2_X1 U10364 ( .A(n10498), .B(n10499), .Z(n10497) );
  XOR2_X1 U10365 ( .A(n10500), .B(n10501), .Z(n10288) );
  XOR2_X1 U10366 ( .A(n10502), .B(n10503), .Z(n10501) );
  XOR2_X1 U10367 ( .A(n10504), .B(n10505), .Z(n10292) );
  XOR2_X1 U10368 ( .A(n10506), .B(n10507), .Z(n10505) );
  XOR2_X1 U10369 ( .A(n10508), .B(n10509), .Z(n10296) );
  XOR2_X1 U10370 ( .A(n10510), .B(n10511), .Z(n10509) );
  XOR2_X1 U10371 ( .A(n10512), .B(n10513), .Z(n10300) );
  XOR2_X1 U10372 ( .A(n10514), .B(n10515), .Z(n10513) );
  OR2_X1 U10373 ( .A1(n8906), .A2(n8047), .ZN(n10306) );
  XOR2_X1 U10374 ( .A(n10516), .B(n10517), .Z(n10305) );
  XOR2_X1 U10375 ( .A(n10518), .B(n10519), .Z(n10517) );
  XNOR2_X1 U10376 ( .A(n10520), .B(n10521), .ZN(n9889) );
  XNOR2_X1 U10377 ( .A(n10522), .B(n10523), .ZN(n10520) );
  XOR2_X1 U10378 ( .A(n10524), .B(n10525), .Z(n9878) );
  XOR2_X1 U10379 ( .A(n10526), .B(n10527), .Z(n10525) );
  OR2_X1 U10380 ( .A1(n9852), .A2(n9851), .ZN(n9061) );
  INV_X1 U10381 ( .A(n10528), .ZN(n9851) );
  OR2_X1 U10382 ( .A1(n10529), .A2(n9849), .ZN(n10528) );
  AND2_X1 U10383 ( .A1(n10530), .A2(n10531), .ZN(n10529) );
  AND2_X1 U10384 ( .A1(n9859), .A2(n9860), .ZN(n9852) );
  INV_X1 U10385 ( .A(n10310), .ZN(n9860) );
  OR2_X1 U10386 ( .A1(n10532), .A2(n10533), .ZN(n10310) );
  AND2_X1 U10387 ( .A1(n10314), .A2(n10313), .ZN(n10533) );
  AND2_X1 U10388 ( .A1(n10311), .A2(n10534), .ZN(n10532) );
  OR2_X1 U10389 ( .A1(n10313), .A2(n10314), .ZN(n10534) );
  OR2_X1 U10390 ( .A1(n9297), .A2(n8075), .ZN(n10314) );
  OR2_X1 U10391 ( .A1(n10535), .A2(n10536), .ZN(n10313) );
  AND2_X1 U10392 ( .A1(n10527), .A2(n10526), .ZN(n10536) );
  AND2_X1 U10393 ( .A1(n10524), .A2(n10537), .ZN(n10535) );
  OR2_X1 U10394 ( .A1(n10526), .A2(n10527), .ZN(n10537) );
  OR2_X1 U10395 ( .A1(n8902), .A2(n8075), .ZN(n10527) );
  OR2_X1 U10396 ( .A1(n10538), .A2(n10539), .ZN(n10526) );
  AND2_X1 U10397 ( .A1(n10523), .A2(n10522), .ZN(n10539) );
  AND2_X1 U10398 ( .A1(n10521), .A2(n10540), .ZN(n10538) );
  OR2_X1 U10399 ( .A1(n10522), .A2(n10523), .ZN(n10540) );
  OR2_X1 U10400 ( .A1(n10541), .A2(n10542), .ZN(n10523) );
  AND2_X1 U10401 ( .A1(n10519), .A2(n10518), .ZN(n10542) );
  AND2_X1 U10402 ( .A1(n10516), .A2(n10543), .ZN(n10541) );
  OR2_X1 U10403 ( .A1(n10518), .A2(n10519), .ZN(n10543) );
  OR2_X1 U10404 ( .A1(n8910), .A2(n8075), .ZN(n10519) );
  OR2_X1 U10405 ( .A1(n10544), .A2(n10545), .ZN(n10518) );
  AND2_X1 U10406 ( .A1(n10515), .A2(n10514), .ZN(n10545) );
  AND2_X1 U10407 ( .A1(n10512), .A2(n10546), .ZN(n10544) );
  OR2_X1 U10408 ( .A1(n10514), .A2(n10515), .ZN(n10546) );
  OR2_X1 U10409 ( .A1(n8914), .A2(n8075), .ZN(n10515) );
  OR2_X1 U10410 ( .A1(n10547), .A2(n10548), .ZN(n10514) );
  AND2_X1 U10411 ( .A1(n10511), .A2(n10510), .ZN(n10548) );
  AND2_X1 U10412 ( .A1(n10508), .A2(n10549), .ZN(n10547) );
  OR2_X1 U10413 ( .A1(n10510), .A2(n10511), .ZN(n10549) );
  OR2_X1 U10414 ( .A1(n8918), .A2(n8075), .ZN(n10511) );
  OR2_X1 U10415 ( .A1(n10550), .A2(n10551), .ZN(n10510) );
  AND2_X1 U10416 ( .A1(n10507), .A2(n10506), .ZN(n10551) );
  AND2_X1 U10417 ( .A1(n10504), .A2(n10552), .ZN(n10550) );
  OR2_X1 U10418 ( .A1(n10506), .A2(n10507), .ZN(n10552) );
  OR2_X1 U10419 ( .A1(n8922), .A2(n8075), .ZN(n10507) );
  OR2_X1 U10420 ( .A1(n10553), .A2(n10554), .ZN(n10506) );
  AND2_X1 U10421 ( .A1(n10503), .A2(n10502), .ZN(n10554) );
  AND2_X1 U10422 ( .A1(n10500), .A2(n10555), .ZN(n10553) );
  OR2_X1 U10423 ( .A1(n10502), .A2(n10503), .ZN(n10555) );
  OR2_X1 U10424 ( .A1(n8926), .A2(n8075), .ZN(n10503) );
  OR2_X1 U10425 ( .A1(n10556), .A2(n10557), .ZN(n10502) );
  AND2_X1 U10426 ( .A1(n10499), .A2(n10498), .ZN(n10557) );
  AND2_X1 U10427 ( .A1(n10496), .A2(n10558), .ZN(n10556) );
  OR2_X1 U10428 ( .A1(n10498), .A2(n10499), .ZN(n10558) );
  OR2_X1 U10429 ( .A1(n8930), .A2(n8075), .ZN(n10499) );
  OR2_X1 U10430 ( .A1(n10559), .A2(n10560), .ZN(n10498) );
  AND2_X1 U10431 ( .A1(n10495), .A2(n10494), .ZN(n10560) );
  AND2_X1 U10432 ( .A1(n10492), .A2(n10561), .ZN(n10559) );
  OR2_X1 U10433 ( .A1(n10494), .A2(n10495), .ZN(n10561) );
  OR2_X1 U10434 ( .A1(n8934), .A2(n8075), .ZN(n10495) );
  OR2_X1 U10435 ( .A1(n10562), .A2(n10563), .ZN(n10494) );
  AND2_X1 U10436 ( .A1(n10491), .A2(n10490), .ZN(n10563) );
  AND2_X1 U10437 ( .A1(n10488), .A2(n10564), .ZN(n10562) );
  OR2_X1 U10438 ( .A1(n10490), .A2(n10491), .ZN(n10564) );
  OR2_X1 U10439 ( .A1(n8938), .A2(n8075), .ZN(n10491) );
  OR2_X1 U10440 ( .A1(n10565), .A2(n10566), .ZN(n10490) );
  AND2_X1 U10441 ( .A1(n10487), .A2(n10486), .ZN(n10566) );
  AND2_X1 U10442 ( .A1(n10484), .A2(n10567), .ZN(n10565) );
  OR2_X1 U10443 ( .A1(n10486), .A2(n10487), .ZN(n10567) );
  OR2_X1 U10444 ( .A1(n8942), .A2(n8075), .ZN(n10487) );
  OR2_X1 U10445 ( .A1(n10568), .A2(n10569), .ZN(n10486) );
  AND2_X1 U10446 ( .A1(n10483), .A2(n10482), .ZN(n10569) );
  AND2_X1 U10447 ( .A1(n10480), .A2(n10570), .ZN(n10568) );
  OR2_X1 U10448 ( .A1(n10482), .A2(n10483), .ZN(n10570) );
  OR2_X1 U10449 ( .A1(n8946), .A2(n8075), .ZN(n10483) );
  OR2_X1 U10450 ( .A1(n10571), .A2(n10572), .ZN(n10482) );
  AND2_X1 U10451 ( .A1(n10479), .A2(n10478), .ZN(n10572) );
  AND2_X1 U10452 ( .A1(n10476), .A2(n10573), .ZN(n10571) );
  OR2_X1 U10453 ( .A1(n10478), .A2(n10479), .ZN(n10573) );
  OR2_X1 U10454 ( .A1(n8950), .A2(n8075), .ZN(n10479) );
  OR2_X1 U10455 ( .A1(n10574), .A2(n10575), .ZN(n10478) );
  AND2_X1 U10456 ( .A1(n10475), .A2(n10474), .ZN(n10575) );
  AND2_X1 U10457 ( .A1(n10472), .A2(n10576), .ZN(n10574) );
  OR2_X1 U10458 ( .A1(n10474), .A2(n10475), .ZN(n10576) );
  OR2_X1 U10459 ( .A1(n8954), .A2(n8075), .ZN(n10475) );
  OR2_X1 U10460 ( .A1(n10577), .A2(n10578), .ZN(n10474) );
  AND2_X1 U10461 ( .A1(n10471), .A2(n10470), .ZN(n10578) );
  AND2_X1 U10462 ( .A1(n10468), .A2(n10579), .ZN(n10577) );
  OR2_X1 U10463 ( .A1(n10470), .A2(n10471), .ZN(n10579) );
  OR2_X1 U10464 ( .A1(n8958), .A2(n8075), .ZN(n10471) );
  OR2_X1 U10465 ( .A1(n10580), .A2(n10581), .ZN(n10470) );
  AND2_X1 U10466 ( .A1(n10467), .A2(n10466), .ZN(n10581) );
  AND2_X1 U10467 ( .A1(n10464), .A2(n10582), .ZN(n10580) );
  OR2_X1 U10468 ( .A1(n10466), .A2(n10467), .ZN(n10582) );
  OR2_X1 U10469 ( .A1(n8962), .A2(n8075), .ZN(n10467) );
  OR2_X1 U10470 ( .A1(n10583), .A2(n10584), .ZN(n10466) );
  AND2_X1 U10471 ( .A1(n10463), .A2(n10462), .ZN(n10584) );
  AND2_X1 U10472 ( .A1(n10460), .A2(n10585), .ZN(n10583) );
  OR2_X1 U10473 ( .A1(n10462), .A2(n10463), .ZN(n10585) );
  OR2_X1 U10474 ( .A1(n8966), .A2(n8075), .ZN(n10463) );
  OR2_X1 U10475 ( .A1(n10586), .A2(n10587), .ZN(n10462) );
  AND2_X1 U10476 ( .A1(n10459), .A2(n10458), .ZN(n10587) );
  AND2_X1 U10477 ( .A1(n10456), .A2(n10588), .ZN(n10586) );
  OR2_X1 U10478 ( .A1(n10458), .A2(n10459), .ZN(n10588) );
  OR2_X1 U10479 ( .A1(n8970), .A2(n8075), .ZN(n10459) );
  OR2_X1 U10480 ( .A1(n10589), .A2(n10590), .ZN(n10458) );
  AND2_X1 U10481 ( .A1(n10455), .A2(n10454), .ZN(n10590) );
  AND2_X1 U10482 ( .A1(n10452), .A2(n10591), .ZN(n10589) );
  OR2_X1 U10483 ( .A1(n10454), .A2(n10455), .ZN(n10591) );
  OR2_X1 U10484 ( .A1(n8974), .A2(n8075), .ZN(n10455) );
  OR2_X1 U10485 ( .A1(n10592), .A2(n10593), .ZN(n10454) );
  AND2_X1 U10486 ( .A1(n10451), .A2(n10450), .ZN(n10593) );
  AND2_X1 U10487 ( .A1(n10448), .A2(n10594), .ZN(n10592) );
  OR2_X1 U10488 ( .A1(n10450), .A2(n10451), .ZN(n10594) );
  OR2_X1 U10489 ( .A1(n8978), .A2(n8075), .ZN(n10451) );
  OR2_X1 U10490 ( .A1(n10595), .A2(n10596), .ZN(n10450) );
  AND2_X1 U10491 ( .A1(n10447), .A2(n10446), .ZN(n10596) );
  AND2_X1 U10492 ( .A1(n10444), .A2(n10597), .ZN(n10595) );
  OR2_X1 U10493 ( .A1(n10446), .A2(n10447), .ZN(n10597) );
  OR2_X1 U10494 ( .A1(n8982), .A2(n8075), .ZN(n10447) );
  OR2_X1 U10495 ( .A1(n10598), .A2(n10599), .ZN(n10446) );
  AND2_X1 U10496 ( .A1(n10443), .A2(n10442), .ZN(n10599) );
  AND2_X1 U10497 ( .A1(n10440), .A2(n10600), .ZN(n10598) );
  OR2_X1 U10498 ( .A1(n10442), .A2(n10443), .ZN(n10600) );
  OR2_X1 U10499 ( .A1(n8986), .A2(n8075), .ZN(n10443) );
  OR2_X1 U10500 ( .A1(n10601), .A2(n10602), .ZN(n10442) );
  AND2_X1 U10501 ( .A1(n10439), .A2(n10438), .ZN(n10602) );
  AND2_X1 U10502 ( .A1(n10436), .A2(n10603), .ZN(n10601) );
  OR2_X1 U10503 ( .A1(n10438), .A2(n10439), .ZN(n10603) );
  OR2_X1 U10504 ( .A1(n8990), .A2(n8075), .ZN(n10439) );
  OR2_X1 U10505 ( .A1(n10604), .A2(n10605), .ZN(n10438) );
  AND2_X1 U10506 ( .A1(n10435), .A2(n10434), .ZN(n10605) );
  AND2_X1 U10507 ( .A1(n10432), .A2(n10606), .ZN(n10604) );
  OR2_X1 U10508 ( .A1(n10434), .A2(n10435), .ZN(n10606) );
  OR2_X1 U10509 ( .A1(n8994), .A2(n8075), .ZN(n10435) );
  OR2_X1 U10510 ( .A1(n10607), .A2(n10608), .ZN(n10434) );
  AND2_X1 U10511 ( .A1(n10431), .A2(n10430), .ZN(n10608) );
  AND2_X1 U10512 ( .A1(n10428), .A2(n10609), .ZN(n10607) );
  OR2_X1 U10513 ( .A1(n10430), .A2(n10431), .ZN(n10609) );
  OR2_X1 U10514 ( .A1(n8998), .A2(n8075), .ZN(n10431) );
  OR2_X1 U10515 ( .A1(n10610), .A2(n10611), .ZN(n10430) );
  AND2_X1 U10516 ( .A1(n10427), .A2(n10426), .ZN(n10611) );
  AND2_X1 U10517 ( .A1(n10424), .A2(n10612), .ZN(n10610) );
  OR2_X1 U10518 ( .A1(n10426), .A2(n10427), .ZN(n10612) );
  OR2_X1 U10519 ( .A1(n9002), .A2(n8075), .ZN(n10427) );
  OR2_X1 U10520 ( .A1(n10613), .A2(n10614), .ZN(n10426) );
  AND2_X1 U10521 ( .A1(n10423), .A2(n10422), .ZN(n10614) );
  AND2_X1 U10522 ( .A1(n10420), .A2(n10615), .ZN(n10613) );
  OR2_X1 U10523 ( .A1(n10422), .A2(n10423), .ZN(n10615) );
  OR2_X1 U10524 ( .A1(n9006), .A2(n8075), .ZN(n10423) );
  OR2_X1 U10525 ( .A1(n10616), .A2(n10617), .ZN(n10422) );
  AND2_X1 U10526 ( .A1(n9011), .A2(n10419), .ZN(n10617) );
  AND2_X1 U10527 ( .A1(n10417), .A2(n10618), .ZN(n10616) );
  OR2_X1 U10528 ( .A1(n10419), .A2(n9011), .ZN(n10618) );
  OR2_X1 U10529 ( .A1(n9010), .A2(n8075), .ZN(n9011) );
  OR2_X1 U10530 ( .A1(n10619), .A2(n10620), .ZN(n10419) );
  AND2_X1 U10531 ( .A1(n10414), .A2(n10415), .ZN(n10620) );
  AND2_X1 U10532 ( .A1(n10621), .A2(n10622), .ZN(n10619) );
  OR2_X1 U10533 ( .A1(n10415), .A2(n10414), .ZN(n10622) );
  OR2_X1 U10534 ( .A1(n9014), .A2(n8075), .ZN(n10414) );
  OR2_X1 U10535 ( .A1(n9984), .A2(n10623), .ZN(n10415) );
  OR2_X1 U10536 ( .A1(n8075), .A2(n8112), .ZN(n10623) );
  INV_X1 U10537 ( .A(n10416), .ZN(n10621) );
  OR2_X1 U10538 ( .A1(n10624), .A2(n10625), .ZN(n10416) );
  AND2_X1 U10539 ( .A1(b_27_), .A2(n10626), .ZN(n10625) );
  OR2_X1 U10540 ( .A1(n10627), .A2(n9989), .ZN(n10626) );
  AND2_X1 U10541 ( .A1(a_30_), .A2(n8140), .ZN(n10627) );
  AND2_X1 U10542 ( .A1(b_26_), .A2(n10628), .ZN(n10624) );
  OR2_X1 U10543 ( .A1(n10629), .A2(n8021), .ZN(n10628) );
  AND2_X1 U10544 ( .A1(a_31_), .A2(n8112), .ZN(n10629) );
  XOR2_X1 U10545 ( .A(n10630), .B(n10631), .Z(n10417) );
  XNOR2_X1 U10546 ( .A(n10632), .B(n10633), .ZN(n10630) );
  XOR2_X1 U10547 ( .A(n10634), .B(n10635), .Z(n10420) );
  XOR2_X1 U10548 ( .A(n10636), .B(n10637), .Z(n10635) );
  XOR2_X1 U10549 ( .A(n10638), .B(n10639), .Z(n10424) );
  XOR2_X1 U10550 ( .A(n10640), .B(n9007), .Z(n10639) );
  XOR2_X1 U10551 ( .A(n10641), .B(n10642), .Z(n10428) );
  XOR2_X1 U10552 ( .A(n10643), .B(n10644), .Z(n10642) );
  XOR2_X1 U10553 ( .A(n10645), .B(n10646), .Z(n10432) );
  XOR2_X1 U10554 ( .A(n10647), .B(n10648), .Z(n10646) );
  XOR2_X1 U10555 ( .A(n10649), .B(n10650), .Z(n10436) );
  XOR2_X1 U10556 ( .A(n10651), .B(n10652), .Z(n10650) );
  XOR2_X1 U10557 ( .A(n10653), .B(n10654), .Z(n10440) );
  XOR2_X1 U10558 ( .A(n10655), .B(n10656), .Z(n10654) );
  XOR2_X1 U10559 ( .A(n10657), .B(n10658), .Z(n10444) );
  XOR2_X1 U10560 ( .A(n10659), .B(n10660), .Z(n10658) );
  XOR2_X1 U10561 ( .A(n10661), .B(n10662), .Z(n10448) );
  XOR2_X1 U10562 ( .A(n10663), .B(n10664), .Z(n10662) );
  XOR2_X1 U10563 ( .A(n10665), .B(n10666), .Z(n10452) );
  XOR2_X1 U10564 ( .A(n10667), .B(n10668), .Z(n10666) );
  XOR2_X1 U10565 ( .A(n10669), .B(n10670), .Z(n10456) );
  XOR2_X1 U10566 ( .A(n10671), .B(n10672), .Z(n10670) );
  XOR2_X1 U10567 ( .A(n10673), .B(n10674), .Z(n10460) );
  XOR2_X1 U10568 ( .A(n10675), .B(n10676), .Z(n10674) );
  XOR2_X1 U10569 ( .A(n10677), .B(n10678), .Z(n10464) );
  XOR2_X1 U10570 ( .A(n10679), .B(n10680), .Z(n10678) );
  XOR2_X1 U10571 ( .A(n10681), .B(n10682), .Z(n10468) );
  XOR2_X1 U10572 ( .A(n10683), .B(n10684), .Z(n10682) );
  XOR2_X1 U10573 ( .A(n10685), .B(n10686), .Z(n10472) );
  XOR2_X1 U10574 ( .A(n10687), .B(n10688), .Z(n10686) );
  XOR2_X1 U10575 ( .A(n10689), .B(n10690), .Z(n10476) );
  XOR2_X1 U10576 ( .A(n10691), .B(n10692), .Z(n10690) );
  XOR2_X1 U10577 ( .A(n10693), .B(n10694), .Z(n10480) );
  XOR2_X1 U10578 ( .A(n10695), .B(n10696), .Z(n10694) );
  XOR2_X1 U10579 ( .A(n10697), .B(n10698), .Z(n10484) );
  XOR2_X1 U10580 ( .A(n10699), .B(n10700), .Z(n10698) );
  XOR2_X1 U10581 ( .A(n10701), .B(n10702), .Z(n10488) );
  XOR2_X1 U10582 ( .A(n10703), .B(n10704), .Z(n10702) );
  XOR2_X1 U10583 ( .A(n10705), .B(n10706), .Z(n10492) );
  XOR2_X1 U10584 ( .A(n10707), .B(n10708), .Z(n10706) );
  XOR2_X1 U10585 ( .A(n10709), .B(n10710), .Z(n10496) );
  XOR2_X1 U10586 ( .A(n10711), .B(n10712), .Z(n10710) );
  XOR2_X1 U10587 ( .A(n10713), .B(n10714), .Z(n10500) );
  XOR2_X1 U10588 ( .A(n10715), .B(n10716), .Z(n10714) );
  XOR2_X1 U10589 ( .A(n10717), .B(n10718), .Z(n10504) );
  XOR2_X1 U10590 ( .A(n10719), .B(n10720), .Z(n10718) );
  XNOR2_X1 U10591 ( .A(n10721), .B(n10722), .ZN(n10508) );
  XNOR2_X1 U10592 ( .A(n10723), .B(n10724), .ZN(n10721) );
  XOR2_X1 U10593 ( .A(n10725), .B(n10726), .Z(n10512) );
  XOR2_X1 U10594 ( .A(n10727), .B(n10728), .Z(n10726) );
  XOR2_X1 U10595 ( .A(n10729), .B(n10730), .Z(n10516) );
  XOR2_X1 U10596 ( .A(n10731), .B(n10732), .Z(n10730) );
  OR2_X1 U10597 ( .A1(n8906), .A2(n8075), .ZN(n10522) );
  XOR2_X1 U10598 ( .A(n10733), .B(n10734), .Z(n10521) );
  XOR2_X1 U10599 ( .A(n10735), .B(n10736), .Z(n10734) );
  XNOR2_X1 U10600 ( .A(n10737), .B(n10738), .ZN(n10524) );
  XNOR2_X1 U10601 ( .A(n10739), .B(n10740), .ZN(n10737) );
  XOR2_X1 U10602 ( .A(n10741), .B(n10742), .Z(n10311) );
  XOR2_X1 U10603 ( .A(n10743), .B(n10744), .Z(n10742) );
  XNOR2_X1 U10604 ( .A(n10745), .B(n10746), .ZN(n9859) );
  XOR2_X1 U10605 ( .A(n10747), .B(n10748), .Z(n10746) );
  OR2_X1 U10606 ( .A1(n9849), .A2(n9848), .ZN(n9068) );
  XOR2_X1 U10607 ( .A(n9845), .B(n9846), .Z(n9848) );
  OR2_X1 U10608 ( .A1(n10749), .A2(n10750), .ZN(n9846) );
  AND2_X1 U10609 ( .A1(n10751), .A2(n10752), .ZN(n10750) );
  AND2_X1 U10610 ( .A1(n10753), .A2(n10754), .ZN(n10749) );
  OR2_X1 U10611 ( .A1(n10751), .A2(n10752), .ZN(n10754) );
  XOR2_X1 U10612 ( .A(n9839), .B(n10755), .Z(n9845) );
  XOR2_X1 U10613 ( .A(n9838), .B(n9837), .Z(n10755) );
  OR2_X1 U10614 ( .A1(n9297), .A2(n8168), .ZN(n9837) );
  OR2_X1 U10615 ( .A1(n10756), .A2(n10757), .ZN(n9838) );
  AND2_X1 U10616 ( .A1(n10758), .A2(n10759), .ZN(n10757) );
  AND2_X1 U10617 ( .A1(n10760), .A2(n10761), .ZN(n10756) );
  OR2_X1 U10618 ( .A1(n10758), .A2(n10759), .ZN(n10761) );
  XNOR2_X1 U10619 ( .A(n10762), .B(n10763), .ZN(n9839) );
  XNOR2_X1 U10620 ( .A(n10764), .B(n10765), .ZN(n10762) );
  INV_X1 U10621 ( .A(n10766), .ZN(n9849) );
  OR2_X1 U10622 ( .A1(n10530), .A2(n10531), .ZN(n10766) );
  OR2_X1 U10623 ( .A1(n10767), .A2(n10768), .ZN(n10531) );
  AND2_X1 U10624 ( .A1(n10745), .A2(n10748), .ZN(n10768) );
  AND2_X1 U10625 ( .A1(n10769), .A2(n10747), .ZN(n10767) );
  OR2_X1 U10626 ( .A1(n10770), .A2(n10771), .ZN(n10747) );
  AND2_X1 U10627 ( .A1(n10744), .A2(n10743), .ZN(n10771) );
  AND2_X1 U10628 ( .A1(n10741), .A2(n10772), .ZN(n10770) );
  OR2_X1 U10629 ( .A1(n10743), .A2(n10744), .ZN(n10772) );
  OR2_X1 U10630 ( .A1(n8902), .A2(n8112), .ZN(n10744) );
  OR2_X1 U10631 ( .A1(n10773), .A2(n10774), .ZN(n10743) );
  AND2_X1 U10632 ( .A1(n10740), .A2(n10739), .ZN(n10774) );
  AND2_X1 U10633 ( .A1(n10738), .A2(n10775), .ZN(n10773) );
  OR2_X1 U10634 ( .A1(n10739), .A2(n10740), .ZN(n10775) );
  OR2_X1 U10635 ( .A1(n10776), .A2(n10777), .ZN(n10740) );
  AND2_X1 U10636 ( .A1(n10736), .A2(n10735), .ZN(n10777) );
  AND2_X1 U10637 ( .A1(n10733), .A2(n10778), .ZN(n10776) );
  OR2_X1 U10638 ( .A1(n10735), .A2(n10736), .ZN(n10778) );
  OR2_X1 U10639 ( .A1(n8910), .A2(n8112), .ZN(n10736) );
  OR2_X1 U10640 ( .A1(n10779), .A2(n10780), .ZN(n10735) );
  AND2_X1 U10641 ( .A1(n10732), .A2(n10731), .ZN(n10780) );
  AND2_X1 U10642 ( .A1(n10729), .A2(n10781), .ZN(n10779) );
  OR2_X1 U10643 ( .A1(n10731), .A2(n10732), .ZN(n10781) );
  OR2_X1 U10644 ( .A1(n8914), .A2(n8112), .ZN(n10732) );
  OR2_X1 U10645 ( .A1(n10782), .A2(n10783), .ZN(n10731) );
  AND2_X1 U10646 ( .A1(n10728), .A2(n10727), .ZN(n10783) );
  AND2_X1 U10647 ( .A1(n10725), .A2(n10784), .ZN(n10782) );
  OR2_X1 U10648 ( .A1(n10727), .A2(n10728), .ZN(n10784) );
  OR2_X1 U10649 ( .A1(n8918), .A2(n8112), .ZN(n10728) );
  OR2_X1 U10650 ( .A1(n10785), .A2(n10786), .ZN(n10727) );
  AND2_X1 U10651 ( .A1(n10724), .A2(n10723), .ZN(n10786) );
  AND2_X1 U10652 ( .A1(n10722), .A2(n10787), .ZN(n10785) );
  OR2_X1 U10653 ( .A1(n10723), .A2(n10724), .ZN(n10787) );
  OR2_X1 U10654 ( .A1(n10788), .A2(n10789), .ZN(n10724) );
  AND2_X1 U10655 ( .A1(n10720), .A2(n10719), .ZN(n10789) );
  AND2_X1 U10656 ( .A1(n10717), .A2(n10790), .ZN(n10788) );
  OR2_X1 U10657 ( .A1(n10719), .A2(n10720), .ZN(n10790) );
  OR2_X1 U10658 ( .A1(n8926), .A2(n8112), .ZN(n10720) );
  OR2_X1 U10659 ( .A1(n10791), .A2(n10792), .ZN(n10719) );
  AND2_X1 U10660 ( .A1(n10716), .A2(n10715), .ZN(n10792) );
  AND2_X1 U10661 ( .A1(n10713), .A2(n10793), .ZN(n10791) );
  OR2_X1 U10662 ( .A1(n10715), .A2(n10716), .ZN(n10793) );
  OR2_X1 U10663 ( .A1(n8930), .A2(n8112), .ZN(n10716) );
  OR2_X1 U10664 ( .A1(n10794), .A2(n10795), .ZN(n10715) );
  AND2_X1 U10665 ( .A1(n10712), .A2(n10711), .ZN(n10795) );
  AND2_X1 U10666 ( .A1(n10709), .A2(n10796), .ZN(n10794) );
  OR2_X1 U10667 ( .A1(n10711), .A2(n10712), .ZN(n10796) );
  OR2_X1 U10668 ( .A1(n8934), .A2(n8112), .ZN(n10712) );
  OR2_X1 U10669 ( .A1(n10797), .A2(n10798), .ZN(n10711) );
  AND2_X1 U10670 ( .A1(n10708), .A2(n10707), .ZN(n10798) );
  AND2_X1 U10671 ( .A1(n10705), .A2(n10799), .ZN(n10797) );
  OR2_X1 U10672 ( .A1(n10707), .A2(n10708), .ZN(n10799) );
  OR2_X1 U10673 ( .A1(n8938), .A2(n8112), .ZN(n10708) );
  OR2_X1 U10674 ( .A1(n10800), .A2(n10801), .ZN(n10707) );
  AND2_X1 U10675 ( .A1(n10704), .A2(n10703), .ZN(n10801) );
  AND2_X1 U10676 ( .A1(n10701), .A2(n10802), .ZN(n10800) );
  OR2_X1 U10677 ( .A1(n10703), .A2(n10704), .ZN(n10802) );
  OR2_X1 U10678 ( .A1(n8942), .A2(n8112), .ZN(n10704) );
  OR2_X1 U10679 ( .A1(n10803), .A2(n10804), .ZN(n10703) );
  AND2_X1 U10680 ( .A1(n10700), .A2(n10699), .ZN(n10804) );
  AND2_X1 U10681 ( .A1(n10697), .A2(n10805), .ZN(n10803) );
  OR2_X1 U10682 ( .A1(n10699), .A2(n10700), .ZN(n10805) );
  OR2_X1 U10683 ( .A1(n8946), .A2(n8112), .ZN(n10700) );
  OR2_X1 U10684 ( .A1(n10806), .A2(n10807), .ZN(n10699) );
  AND2_X1 U10685 ( .A1(n10696), .A2(n10695), .ZN(n10807) );
  AND2_X1 U10686 ( .A1(n10693), .A2(n10808), .ZN(n10806) );
  OR2_X1 U10687 ( .A1(n10695), .A2(n10696), .ZN(n10808) );
  OR2_X1 U10688 ( .A1(n8950), .A2(n8112), .ZN(n10696) );
  OR2_X1 U10689 ( .A1(n10809), .A2(n10810), .ZN(n10695) );
  AND2_X1 U10690 ( .A1(n10692), .A2(n10691), .ZN(n10810) );
  AND2_X1 U10691 ( .A1(n10689), .A2(n10811), .ZN(n10809) );
  OR2_X1 U10692 ( .A1(n10691), .A2(n10692), .ZN(n10811) );
  OR2_X1 U10693 ( .A1(n8954), .A2(n8112), .ZN(n10692) );
  OR2_X1 U10694 ( .A1(n10812), .A2(n10813), .ZN(n10691) );
  AND2_X1 U10695 ( .A1(n10688), .A2(n10687), .ZN(n10813) );
  AND2_X1 U10696 ( .A1(n10685), .A2(n10814), .ZN(n10812) );
  OR2_X1 U10697 ( .A1(n10687), .A2(n10688), .ZN(n10814) );
  OR2_X1 U10698 ( .A1(n8958), .A2(n8112), .ZN(n10688) );
  OR2_X1 U10699 ( .A1(n10815), .A2(n10816), .ZN(n10687) );
  AND2_X1 U10700 ( .A1(n10684), .A2(n10683), .ZN(n10816) );
  AND2_X1 U10701 ( .A1(n10681), .A2(n10817), .ZN(n10815) );
  OR2_X1 U10702 ( .A1(n10683), .A2(n10684), .ZN(n10817) );
  OR2_X1 U10703 ( .A1(n8962), .A2(n8112), .ZN(n10684) );
  OR2_X1 U10704 ( .A1(n10818), .A2(n10819), .ZN(n10683) );
  AND2_X1 U10705 ( .A1(n10680), .A2(n10679), .ZN(n10819) );
  AND2_X1 U10706 ( .A1(n10677), .A2(n10820), .ZN(n10818) );
  OR2_X1 U10707 ( .A1(n10679), .A2(n10680), .ZN(n10820) );
  OR2_X1 U10708 ( .A1(n8966), .A2(n8112), .ZN(n10680) );
  OR2_X1 U10709 ( .A1(n10821), .A2(n10822), .ZN(n10679) );
  AND2_X1 U10710 ( .A1(n10676), .A2(n10675), .ZN(n10822) );
  AND2_X1 U10711 ( .A1(n10673), .A2(n10823), .ZN(n10821) );
  OR2_X1 U10712 ( .A1(n10675), .A2(n10676), .ZN(n10823) );
  OR2_X1 U10713 ( .A1(n8970), .A2(n8112), .ZN(n10676) );
  OR2_X1 U10714 ( .A1(n10824), .A2(n10825), .ZN(n10675) );
  AND2_X1 U10715 ( .A1(n10672), .A2(n10671), .ZN(n10825) );
  AND2_X1 U10716 ( .A1(n10669), .A2(n10826), .ZN(n10824) );
  OR2_X1 U10717 ( .A1(n10671), .A2(n10672), .ZN(n10826) );
  OR2_X1 U10718 ( .A1(n8974), .A2(n8112), .ZN(n10672) );
  OR2_X1 U10719 ( .A1(n10827), .A2(n10828), .ZN(n10671) );
  AND2_X1 U10720 ( .A1(n10668), .A2(n10667), .ZN(n10828) );
  AND2_X1 U10721 ( .A1(n10665), .A2(n10829), .ZN(n10827) );
  OR2_X1 U10722 ( .A1(n10667), .A2(n10668), .ZN(n10829) );
  OR2_X1 U10723 ( .A1(n8978), .A2(n8112), .ZN(n10668) );
  OR2_X1 U10724 ( .A1(n10830), .A2(n10831), .ZN(n10667) );
  AND2_X1 U10725 ( .A1(n10664), .A2(n10663), .ZN(n10831) );
  AND2_X1 U10726 ( .A1(n10661), .A2(n10832), .ZN(n10830) );
  OR2_X1 U10727 ( .A1(n10663), .A2(n10664), .ZN(n10832) );
  OR2_X1 U10728 ( .A1(n8982), .A2(n8112), .ZN(n10664) );
  OR2_X1 U10729 ( .A1(n10833), .A2(n10834), .ZN(n10663) );
  AND2_X1 U10730 ( .A1(n10660), .A2(n10659), .ZN(n10834) );
  AND2_X1 U10731 ( .A1(n10657), .A2(n10835), .ZN(n10833) );
  OR2_X1 U10732 ( .A1(n10659), .A2(n10660), .ZN(n10835) );
  OR2_X1 U10733 ( .A1(n8986), .A2(n8112), .ZN(n10660) );
  OR2_X1 U10734 ( .A1(n10836), .A2(n10837), .ZN(n10659) );
  AND2_X1 U10735 ( .A1(n10656), .A2(n10655), .ZN(n10837) );
  AND2_X1 U10736 ( .A1(n10653), .A2(n10838), .ZN(n10836) );
  OR2_X1 U10737 ( .A1(n10655), .A2(n10656), .ZN(n10838) );
  OR2_X1 U10738 ( .A1(n8990), .A2(n8112), .ZN(n10656) );
  OR2_X1 U10739 ( .A1(n10839), .A2(n10840), .ZN(n10655) );
  AND2_X1 U10740 ( .A1(n10652), .A2(n10651), .ZN(n10840) );
  AND2_X1 U10741 ( .A1(n10649), .A2(n10841), .ZN(n10839) );
  OR2_X1 U10742 ( .A1(n10651), .A2(n10652), .ZN(n10841) );
  OR2_X1 U10743 ( .A1(n8994), .A2(n8112), .ZN(n10652) );
  OR2_X1 U10744 ( .A1(n10842), .A2(n10843), .ZN(n10651) );
  AND2_X1 U10745 ( .A1(n10648), .A2(n10647), .ZN(n10843) );
  AND2_X1 U10746 ( .A1(n10645), .A2(n10844), .ZN(n10842) );
  OR2_X1 U10747 ( .A1(n10647), .A2(n10648), .ZN(n10844) );
  OR2_X1 U10748 ( .A1(n8998), .A2(n8112), .ZN(n10648) );
  OR2_X1 U10749 ( .A1(n10845), .A2(n10846), .ZN(n10647) );
  AND2_X1 U10750 ( .A1(n10644), .A2(n10643), .ZN(n10846) );
  AND2_X1 U10751 ( .A1(n10641), .A2(n10847), .ZN(n10845) );
  OR2_X1 U10752 ( .A1(n10643), .A2(n10644), .ZN(n10847) );
  OR2_X1 U10753 ( .A1(n9002), .A2(n8112), .ZN(n10644) );
  OR2_X1 U10754 ( .A1(n10848), .A2(n10849), .ZN(n10643) );
  AND2_X1 U10755 ( .A1(n9007), .A2(n10640), .ZN(n10849) );
  AND2_X1 U10756 ( .A1(n10638), .A2(n10850), .ZN(n10848) );
  OR2_X1 U10757 ( .A1(n10640), .A2(n9007), .ZN(n10850) );
  OR2_X1 U10758 ( .A1(n9006), .A2(n8112), .ZN(n9007) );
  OR2_X1 U10759 ( .A1(n10851), .A2(n10852), .ZN(n10640) );
  AND2_X1 U10760 ( .A1(n10637), .A2(n10636), .ZN(n10852) );
  AND2_X1 U10761 ( .A1(n10634), .A2(n10853), .ZN(n10851) );
  OR2_X1 U10762 ( .A1(n10636), .A2(n10637), .ZN(n10853) );
  OR2_X1 U10763 ( .A1(n9010), .A2(n8112), .ZN(n10637) );
  OR2_X1 U10764 ( .A1(n10854), .A2(n10855), .ZN(n10636) );
  AND2_X1 U10765 ( .A1(n10631), .A2(n10632), .ZN(n10855) );
  AND2_X1 U10766 ( .A1(n10856), .A2(n10857), .ZN(n10854) );
  OR2_X1 U10767 ( .A1(n10632), .A2(n10631), .ZN(n10857) );
  OR2_X1 U10768 ( .A1(n9014), .A2(n8112), .ZN(n10631) );
  OR2_X1 U10769 ( .A1(n9984), .A2(n10858), .ZN(n10632) );
  OR2_X1 U10770 ( .A1(n8112), .A2(n8140), .ZN(n10858) );
  INV_X1 U10771 ( .A(n10633), .ZN(n10856) );
  OR2_X1 U10772 ( .A1(n10859), .A2(n10860), .ZN(n10633) );
  AND2_X1 U10773 ( .A1(b_26_), .A2(n10861), .ZN(n10860) );
  OR2_X1 U10774 ( .A1(n10862), .A2(n9989), .ZN(n10861) );
  AND2_X1 U10775 ( .A1(a_30_), .A2(n8168), .ZN(n10862) );
  AND2_X1 U10776 ( .A1(b_25_), .A2(n10863), .ZN(n10859) );
  OR2_X1 U10777 ( .A1(n10864), .A2(n8021), .ZN(n10863) );
  AND2_X1 U10778 ( .A1(a_31_), .A2(n8140), .ZN(n10864) );
  XOR2_X1 U10779 ( .A(n10865), .B(n10866), .Z(n10634) );
  XNOR2_X1 U10780 ( .A(n10867), .B(n10868), .ZN(n10865) );
  XOR2_X1 U10781 ( .A(n10869), .B(n10870), .Z(n10638) );
  XOR2_X1 U10782 ( .A(n10871), .B(n10872), .Z(n10870) );
  XOR2_X1 U10783 ( .A(n10873), .B(n10874), .Z(n10641) );
  XOR2_X1 U10784 ( .A(n10875), .B(n10876), .Z(n10874) );
  XOR2_X1 U10785 ( .A(n10877), .B(n10878), .Z(n10645) );
  XOR2_X1 U10786 ( .A(n10879), .B(n9003), .Z(n10878) );
  XOR2_X1 U10787 ( .A(n10880), .B(n10881), .Z(n10649) );
  XOR2_X1 U10788 ( .A(n10882), .B(n10883), .Z(n10881) );
  XOR2_X1 U10789 ( .A(n10884), .B(n10885), .Z(n10653) );
  XOR2_X1 U10790 ( .A(n10886), .B(n10887), .Z(n10885) );
  XOR2_X1 U10791 ( .A(n10888), .B(n10889), .Z(n10657) );
  XOR2_X1 U10792 ( .A(n10890), .B(n10891), .Z(n10889) );
  XOR2_X1 U10793 ( .A(n10892), .B(n10893), .Z(n10661) );
  XOR2_X1 U10794 ( .A(n10894), .B(n10895), .Z(n10893) );
  XOR2_X1 U10795 ( .A(n10896), .B(n10897), .Z(n10665) );
  XOR2_X1 U10796 ( .A(n10898), .B(n10899), .Z(n10897) );
  XOR2_X1 U10797 ( .A(n10900), .B(n10901), .Z(n10669) );
  XOR2_X1 U10798 ( .A(n10902), .B(n10903), .Z(n10901) );
  XOR2_X1 U10799 ( .A(n10904), .B(n10905), .Z(n10673) );
  XOR2_X1 U10800 ( .A(n10906), .B(n10907), .Z(n10905) );
  XOR2_X1 U10801 ( .A(n10908), .B(n10909), .Z(n10677) );
  XOR2_X1 U10802 ( .A(n10910), .B(n10911), .Z(n10909) );
  XOR2_X1 U10803 ( .A(n10912), .B(n10913), .Z(n10681) );
  XOR2_X1 U10804 ( .A(n10914), .B(n10915), .Z(n10913) );
  XOR2_X1 U10805 ( .A(n10916), .B(n10917), .Z(n10685) );
  XOR2_X1 U10806 ( .A(n10918), .B(n10919), .Z(n10917) );
  XOR2_X1 U10807 ( .A(n10920), .B(n10921), .Z(n10689) );
  XOR2_X1 U10808 ( .A(n10922), .B(n10923), .Z(n10921) );
  XOR2_X1 U10809 ( .A(n10924), .B(n10925), .Z(n10693) );
  XOR2_X1 U10810 ( .A(n10926), .B(n10927), .Z(n10925) );
  XOR2_X1 U10811 ( .A(n10928), .B(n10929), .Z(n10697) );
  XOR2_X1 U10812 ( .A(n10930), .B(n10931), .Z(n10929) );
  XOR2_X1 U10813 ( .A(n10932), .B(n10933), .Z(n10701) );
  XOR2_X1 U10814 ( .A(n10934), .B(n10935), .Z(n10933) );
  XOR2_X1 U10815 ( .A(n10936), .B(n10937), .Z(n10705) );
  XOR2_X1 U10816 ( .A(n10938), .B(n10939), .Z(n10937) );
  XOR2_X1 U10817 ( .A(n10940), .B(n10941), .Z(n10709) );
  XOR2_X1 U10818 ( .A(n10942), .B(n10943), .Z(n10941) );
  XOR2_X1 U10819 ( .A(n10944), .B(n10945), .Z(n10713) );
  XOR2_X1 U10820 ( .A(n10946), .B(n10947), .Z(n10945) );
  XOR2_X1 U10821 ( .A(n10948), .B(n10949), .Z(n10717) );
  XOR2_X1 U10822 ( .A(n10950), .B(n10951), .Z(n10949) );
  OR2_X1 U10823 ( .A1(n8922), .A2(n8112), .ZN(n10723) );
  XOR2_X1 U10824 ( .A(n10952), .B(n10953), .Z(n10722) );
  XOR2_X1 U10825 ( .A(n10954), .B(n10955), .Z(n10953) );
  XNOR2_X1 U10826 ( .A(n10956), .B(n10957), .ZN(n10725) );
  XNOR2_X1 U10827 ( .A(n10958), .B(n10959), .ZN(n10956) );
  XOR2_X1 U10828 ( .A(n10960), .B(n10961), .Z(n10729) );
  XOR2_X1 U10829 ( .A(n10962), .B(n10963), .Z(n10961) );
  XOR2_X1 U10830 ( .A(n10964), .B(n10965), .Z(n10733) );
  XOR2_X1 U10831 ( .A(n10966), .B(n10967), .Z(n10965) );
  OR2_X1 U10832 ( .A1(n8906), .A2(n8112), .ZN(n10739) );
  XOR2_X1 U10833 ( .A(n10968), .B(n10969), .Z(n10738) );
  XOR2_X1 U10834 ( .A(n10970), .B(n10971), .Z(n10969) );
  XOR2_X1 U10835 ( .A(n10972), .B(n10973), .Z(n10741) );
  XOR2_X1 U10836 ( .A(n10974), .B(n10975), .Z(n10973) );
  OR2_X1 U10837 ( .A1(n10745), .A2(n10748), .ZN(n10769) );
  OR2_X1 U10838 ( .A1(n9297), .A2(n8112), .ZN(n10748) );
  XOR2_X1 U10839 ( .A(n10976), .B(n10977), .Z(n10745) );
  XOR2_X1 U10840 ( .A(n10978), .B(n10979), .Z(n10977) );
  XOR2_X1 U10841 ( .A(n10753), .B(n10980), .Z(n10530) );
  XOR2_X1 U10842 ( .A(n10752), .B(n10751), .Z(n10980) );
  OR2_X1 U10843 ( .A1(n9297), .A2(n8140), .ZN(n10751) );
  OR2_X1 U10844 ( .A1(n10981), .A2(n10982), .ZN(n10752) );
  AND2_X1 U10845 ( .A1(n10979), .A2(n10978), .ZN(n10982) );
  AND2_X1 U10846 ( .A1(n10976), .A2(n10983), .ZN(n10981) );
  OR2_X1 U10847 ( .A1(n10979), .A2(n10978), .ZN(n10983) );
  OR2_X1 U10848 ( .A1(n10984), .A2(n10985), .ZN(n10978) );
  AND2_X1 U10849 ( .A1(n10975), .A2(n10974), .ZN(n10985) );
  AND2_X1 U10850 ( .A1(n10972), .A2(n10986), .ZN(n10984) );
  OR2_X1 U10851 ( .A1(n10975), .A2(n10974), .ZN(n10986) );
  OR2_X1 U10852 ( .A1(n10987), .A2(n10988), .ZN(n10974) );
  AND2_X1 U10853 ( .A1(n10971), .A2(n10970), .ZN(n10988) );
  AND2_X1 U10854 ( .A1(n10968), .A2(n10989), .ZN(n10987) );
  OR2_X1 U10855 ( .A1(n10971), .A2(n10970), .ZN(n10989) );
  OR2_X1 U10856 ( .A1(n10990), .A2(n10991), .ZN(n10970) );
  AND2_X1 U10857 ( .A1(n10967), .A2(n10966), .ZN(n10991) );
  AND2_X1 U10858 ( .A1(n10964), .A2(n10992), .ZN(n10990) );
  OR2_X1 U10859 ( .A1(n10967), .A2(n10966), .ZN(n10992) );
  OR2_X1 U10860 ( .A1(n10993), .A2(n10994), .ZN(n10966) );
  AND2_X1 U10861 ( .A1(n10963), .A2(n10962), .ZN(n10994) );
  AND2_X1 U10862 ( .A1(n10960), .A2(n10995), .ZN(n10993) );
  OR2_X1 U10863 ( .A1(n10963), .A2(n10962), .ZN(n10995) );
  OR2_X1 U10864 ( .A1(n10996), .A2(n10997), .ZN(n10962) );
  AND2_X1 U10865 ( .A1(n10959), .A2(n10958), .ZN(n10997) );
  AND2_X1 U10866 ( .A1(n10957), .A2(n10998), .ZN(n10996) );
  OR2_X1 U10867 ( .A1(n10959), .A2(n10958), .ZN(n10998) );
  OR2_X1 U10868 ( .A1(n8922), .A2(n8140), .ZN(n10958) );
  OR2_X1 U10869 ( .A1(n10999), .A2(n11000), .ZN(n10959) );
  AND2_X1 U10870 ( .A1(n10955), .A2(n10954), .ZN(n11000) );
  AND2_X1 U10871 ( .A1(n10952), .A2(n11001), .ZN(n10999) );
  OR2_X1 U10872 ( .A1(n10955), .A2(n10954), .ZN(n11001) );
  OR2_X1 U10873 ( .A1(n11002), .A2(n11003), .ZN(n10954) );
  AND2_X1 U10874 ( .A1(n10951), .A2(n10950), .ZN(n11003) );
  AND2_X1 U10875 ( .A1(n10948), .A2(n11004), .ZN(n11002) );
  OR2_X1 U10876 ( .A1(n10951), .A2(n10950), .ZN(n11004) );
  OR2_X1 U10877 ( .A1(n11005), .A2(n11006), .ZN(n10950) );
  AND2_X1 U10878 ( .A1(n10947), .A2(n10946), .ZN(n11006) );
  AND2_X1 U10879 ( .A1(n10944), .A2(n11007), .ZN(n11005) );
  OR2_X1 U10880 ( .A1(n10947), .A2(n10946), .ZN(n11007) );
  OR2_X1 U10881 ( .A1(n11008), .A2(n11009), .ZN(n10946) );
  AND2_X1 U10882 ( .A1(n10943), .A2(n10942), .ZN(n11009) );
  AND2_X1 U10883 ( .A1(n10940), .A2(n11010), .ZN(n11008) );
  OR2_X1 U10884 ( .A1(n10943), .A2(n10942), .ZN(n11010) );
  OR2_X1 U10885 ( .A1(n11011), .A2(n11012), .ZN(n10942) );
  AND2_X1 U10886 ( .A1(n10939), .A2(n10938), .ZN(n11012) );
  AND2_X1 U10887 ( .A1(n10936), .A2(n11013), .ZN(n11011) );
  OR2_X1 U10888 ( .A1(n10939), .A2(n10938), .ZN(n11013) );
  OR2_X1 U10889 ( .A1(n11014), .A2(n11015), .ZN(n10938) );
  AND2_X1 U10890 ( .A1(n10935), .A2(n10934), .ZN(n11015) );
  AND2_X1 U10891 ( .A1(n10932), .A2(n11016), .ZN(n11014) );
  OR2_X1 U10892 ( .A1(n10935), .A2(n10934), .ZN(n11016) );
  OR2_X1 U10893 ( .A1(n11017), .A2(n11018), .ZN(n10934) );
  AND2_X1 U10894 ( .A1(n10931), .A2(n10930), .ZN(n11018) );
  AND2_X1 U10895 ( .A1(n10928), .A2(n11019), .ZN(n11017) );
  OR2_X1 U10896 ( .A1(n10931), .A2(n10930), .ZN(n11019) );
  OR2_X1 U10897 ( .A1(n11020), .A2(n11021), .ZN(n10930) );
  AND2_X1 U10898 ( .A1(n10927), .A2(n10926), .ZN(n11021) );
  AND2_X1 U10899 ( .A1(n10924), .A2(n11022), .ZN(n11020) );
  OR2_X1 U10900 ( .A1(n10927), .A2(n10926), .ZN(n11022) );
  OR2_X1 U10901 ( .A1(n11023), .A2(n11024), .ZN(n10926) );
  AND2_X1 U10902 ( .A1(n10923), .A2(n10922), .ZN(n11024) );
  AND2_X1 U10903 ( .A1(n10920), .A2(n11025), .ZN(n11023) );
  OR2_X1 U10904 ( .A1(n10923), .A2(n10922), .ZN(n11025) );
  OR2_X1 U10905 ( .A1(n11026), .A2(n11027), .ZN(n10922) );
  AND2_X1 U10906 ( .A1(n10919), .A2(n10918), .ZN(n11027) );
  AND2_X1 U10907 ( .A1(n10916), .A2(n11028), .ZN(n11026) );
  OR2_X1 U10908 ( .A1(n10919), .A2(n10918), .ZN(n11028) );
  OR2_X1 U10909 ( .A1(n11029), .A2(n11030), .ZN(n10918) );
  AND2_X1 U10910 ( .A1(n10915), .A2(n10914), .ZN(n11030) );
  AND2_X1 U10911 ( .A1(n10912), .A2(n11031), .ZN(n11029) );
  OR2_X1 U10912 ( .A1(n10915), .A2(n10914), .ZN(n11031) );
  OR2_X1 U10913 ( .A1(n11032), .A2(n11033), .ZN(n10914) );
  AND2_X1 U10914 ( .A1(n10911), .A2(n10910), .ZN(n11033) );
  AND2_X1 U10915 ( .A1(n10908), .A2(n11034), .ZN(n11032) );
  OR2_X1 U10916 ( .A1(n10911), .A2(n10910), .ZN(n11034) );
  OR2_X1 U10917 ( .A1(n11035), .A2(n11036), .ZN(n10910) );
  AND2_X1 U10918 ( .A1(n10907), .A2(n10906), .ZN(n11036) );
  AND2_X1 U10919 ( .A1(n10904), .A2(n11037), .ZN(n11035) );
  OR2_X1 U10920 ( .A1(n10907), .A2(n10906), .ZN(n11037) );
  OR2_X1 U10921 ( .A1(n11038), .A2(n11039), .ZN(n10906) );
  AND2_X1 U10922 ( .A1(n10903), .A2(n10902), .ZN(n11039) );
  AND2_X1 U10923 ( .A1(n10900), .A2(n11040), .ZN(n11038) );
  OR2_X1 U10924 ( .A1(n10903), .A2(n10902), .ZN(n11040) );
  OR2_X1 U10925 ( .A1(n11041), .A2(n11042), .ZN(n10902) );
  AND2_X1 U10926 ( .A1(n10899), .A2(n10898), .ZN(n11042) );
  AND2_X1 U10927 ( .A1(n10896), .A2(n11043), .ZN(n11041) );
  OR2_X1 U10928 ( .A1(n10899), .A2(n10898), .ZN(n11043) );
  OR2_X1 U10929 ( .A1(n11044), .A2(n11045), .ZN(n10898) );
  AND2_X1 U10930 ( .A1(n10895), .A2(n10894), .ZN(n11045) );
  AND2_X1 U10931 ( .A1(n10892), .A2(n11046), .ZN(n11044) );
  OR2_X1 U10932 ( .A1(n10895), .A2(n10894), .ZN(n11046) );
  OR2_X1 U10933 ( .A1(n11047), .A2(n11048), .ZN(n10894) );
  AND2_X1 U10934 ( .A1(n10891), .A2(n10890), .ZN(n11048) );
  AND2_X1 U10935 ( .A1(n10888), .A2(n11049), .ZN(n11047) );
  OR2_X1 U10936 ( .A1(n10891), .A2(n10890), .ZN(n11049) );
  OR2_X1 U10937 ( .A1(n11050), .A2(n11051), .ZN(n10890) );
  AND2_X1 U10938 ( .A1(n10887), .A2(n10886), .ZN(n11051) );
  AND2_X1 U10939 ( .A1(n10884), .A2(n11052), .ZN(n11050) );
  OR2_X1 U10940 ( .A1(n10887), .A2(n10886), .ZN(n11052) );
  OR2_X1 U10941 ( .A1(n11053), .A2(n11054), .ZN(n10886) );
  AND2_X1 U10942 ( .A1(n10883), .A2(n10882), .ZN(n11054) );
  AND2_X1 U10943 ( .A1(n10880), .A2(n11055), .ZN(n11053) );
  OR2_X1 U10944 ( .A1(n10883), .A2(n10882), .ZN(n11055) );
  OR2_X1 U10945 ( .A1(n11056), .A2(n11057), .ZN(n10882) );
  AND2_X1 U10946 ( .A1(n9003), .A2(n10879), .ZN(n11057) );
  AND2_X1 U10947 ( .A1(n10877), .A2(n11058), .ZN(n11056) );
  OR2_X1 U10948 ( .A1(n9003), .A2(n10879), .ZN(n11058) );
  OR2_X1 U10949 ( .A1(n11059), .A2(n11060), .ZN(n10879) );
  AND2_X1 U10950 ( .A1(n10876), .A2(n10875), .ZN(n11060) );
  AND2_X1 U10951 ( .A1(n10873), .A2(n11061), .ZN(n11059) );
  OR2_X1 U10952 ( .A1(n10876), .A2(n10875), .ZN(n11061) );
  OR2_X1 U10953 ( .A1(n11062), .A2(n11063), .ZN(n10875) );
  AND2_X1 U10954 ( .A1(n10872), .A2(n10871), .ZN(n11063) );
  AND2_X1 U10955 ( .A1(n10869), .A2(n11064), .ZN(n11062) );
  OR2_X1 U10956 ( .A1(n10872), .A2(n10871), .ZN(n11064) );
  OR2_X1 U10957 ( .A1(n11065), .A2(n11066), .ZN(n10871) );
  AND2_X1 U10958 ( .A1(n10866), .A2(n10867), .ZN(n11066) );
  AND2_X1 U10959 ( .A1(n11067), .A2(n11068), .ZN(n11065) );
  OR2_X1 U10960 ( .A1(n10866), .A2(n10867), .ZN(n11068) );
  OR2_X1 U10961 ( .A1(n9984), .A2(n11069), .ZN(n10867) );
  OR2_X1 U10962 ( .A1(n8140), .A2(n8168), .ZN(n11069) );
  OR2_X1 U10963 ( .A1(n9014), .A2(n8140), .ZN(n10866) );
  INV_X1 U10964 ( .A(n10868), .ZN(n11067) );
  OR2_X1 U10965 ( .A1(n11070), .A2(n11071), .ZN(n10868) );
  AND2_X1 U10966 ( .A1(b_25_), .A2(n11072), .ZN(n11071) );
  OR2_X1 U10967 ( .A1(n11073), .A2(n9989), .ZN(n11072) );
  AND2_X1 U10968 ( .A1(a_30_), .A2(n8196), .ZN(n11073) );
  AND2_X1 U10969 ( .A1(b_24_), .A2(n11074), .ZN(n11070) );
  OR2_X1 U10970 ( .A1(n11075), .A2(n8021), .ZN(n11074) );
  AND2_X1 U10971 ( .A1(a_31_), .A2(n8168), .ZN(n11075) );
  OR2_X1 U10972 ( .A1(n9010), .A2(n8140), .ZN(n10872) );
  XOR2_X1 U10973 ( .A(n11076), .B(n11077), .Z(n10869) );
  XNOR2_X1 U10974 ( .A(n11078), .B(n11079), .ZN(n11076) );
  OR2_X1 U10975 ( .A1(n9006), .A2(n8140), .ZN(n10876) );
  XOR2_X1 U10976 ( .A(n11080), .B(n11081), .Z(n10873) );
  XOR2_X1 U10977 ( .A(n11082), .B(n11083), .Z(n11081) );
  OR2_X1 U10978 ( .A1(n9002), .A2(n8140), .ZN(n9003) );
  XOR2_X1 U10979 ( .A(n11084), .B(n11085), .Z(n10877) );
  XOR2_X1 U10980 ( .A(n11086), .B(n11087), .Z(n11085) );
  OR2_X1 U10981 ( .A1(n8998), .A2(n8140), .ZN(n10883) );
  XOR2_X1 U10982 ( .A(n11088), .B(n11089), .Z(n10880) );
  XOR2_X1 U10983 ( .A(n11090), .B(n11091), .Z(n11089) );
  OR2_X1 U10984 ( .A1(n8994), .A2(n8140), .ZN(n10887) );
  XOR2_X1 U10985 ( .A(n11092), .B(n11093), .Z(n10884) );
  XOR2_X1 U10986 ( .A(n11094), .B(n8999), .Z(n11093) );
  OR2_X1 U10987 ( .A1(n8990), .A2(n8140), .ZN(n10891) );
  XOR2_X1 U10988 ( .A(n11095), .B(n11096), .Z(n10888) );
  XOR2_X1 U10989 ( .A(n11097), .B(n11098), .Z(n11096) );
  OR2_X1 U10990 ( .A1(n8986), .A2(n8140), .ZN(n10895) );
  XOR2_X1 U10991 ( .A(n11099), .B(n11100), .Z(n10892) );
  XOR2_X1 U10992 ( .A(n11101), .B(n11102), .Z(n11100) );
  OR2_X1 U10993 ( .A1(n8982), .A2(n8140), .ZN(n10899) );
  XOR2_X1 U10994 ( .A(n11103), .B(n11104), .Z(n10896) );
  XOR2_X1 U10995 ( .A(n11105), .B(n11106), .Z(n11104) );
  OR2_X1 U10996 ( .A1(n8978), .A2(n8140), .ZN(n10903) );
  XOR2_X1 U10997 ( .A(n11107), .B(n11108), .Z(n10900) );
  XOR2_X1 U10998 ( .A(n11109), .B(n11110), .Z(n11108) );
  OR2_X1 U10999 ( .A1(n8974), .A2(n8140), .ZN(n10907) );
  XOR2_X1 U11000 ( .A(n11111), .B(n11112), .Z(n10904) );
  XOR2_X1 U11001 ( .A(n11113), .B(n11114), .Z(n11112) );
  OR2_X1 U11002 ( .A1(n8970), .A2(n8140), .ZN(n10911) );
  XOR2_X1 U11003 ( .A(n11115), .B(n11116), .Z(n10908) );
  XOR2_X1 U11004 ( .A(n11117), .B(n11118), .Z(n11116) );
  OR2_X1 U11005 ( .A1(n8966), .A2(n8140), .ZN(n10915) );
  XOR2_X1 U11006 ( .A(n11119), .B(n11120), .Z(n10912) );
  XOR2_X1 U11007 ( .A(n11121), .B(n11122), .Z(n11120) );
  OR2_X1 U11008 ( .A1(n8962), .A2(n8140), .ZN(n10919) );
  XOR2_X1 U11009 ( .A(n11123), .B(n11124), .Z(n10916) );
  XOR2_X1 U11010 ( .A(n11125), .B(n11126), .Z(n11124) );
  OR2_X1 U11011 ( .A1(n8958), .A2(n8140), .ZN(n10923) );
  XOR2_X1 U11012 ( .A(n11127), .B(n11128), .Z(n10920) );
  XOR2_X1 U11013 ( .A(n11129), .B(n11130), .Z(n11128) );
  OR2_X1 U11014 ( .A1(n8954), .A2(n8140), .ZN(n10927) );
  XOR2_X1 U11015 ( .A(n11131), .B(n11132), .Z(n10924) );
  XOR2_X1 U11016 ( .A(n11133), .B(n11134), .Z(n11132) );
  OR2_X1 U11017 ( .A1(n8950), .A2(n8140), .ZN(n10931) );
  XOR2_X1 U11018 ( .A(n11135), .B(n11136), .Z(n10928) );
  XOR2_X1 U11019 ( .A(n11137), .B(n11138), .Z(n11136) );
  OR2_X1 U11020 ( .A1(n8946), .A2(n8140), .ZN(n10935) );
  XOR2_X1 U11021 ( .A(n11139), .B(n11140), .Z(n10932) );
  XOR2_X1 U11022 ( .A(n11141), .B(n11142), .Z(n11140) );
  OR2_X1 U11023 ( .A1(n8942), .A2(n8140), .ZN(n10939) );
  XOR2_X1 U11024 ( .A(n11143), .B(n11144), .Z(n10936) );
  XOR2_X1 U11025 ( .A(n11145), .B(n11146), .Z(n11144) );
  OR2_X1 U11026 ( .A1(n8938), .A2(n8140), .ZN(n10943) );
  XOR2_X1 U11027 ( .A(n11147), .B(n11148), .Z(n10940) );
  XOR2_X1 U11028 ( .A(n11149), .B(n11150), .Z(n11148) );
  OR2_X1 U11029 ( .A1(n8934), .A2(n8140), .ZN(n10947) );
  XNOR2_X1 U11030 ( .A(n11151), .B(n11152), .ZN(n10944) );
  XNOR2_X1 U11031 ( .A(n11153), .B(n11154), .ZN(n11151) );
  OR2_X1 U11032 ( .A1(n8930), .A2(n8140), .ZN(n10951) );
  XOR2_X1 U11033 ( .A(n11155), .B(n11156), .Z(n10948) );
  XOR2_X1 U11034 ( .A(n11157), .B(n11158), .Z(n11156) );
  OR2_X1 U11035 ( .A1(n8926), .A2(n8140), .ZN(n10955) );
  XOR2_X1 U11036 ( .A(n11159), .B(n11160), .Z(n10952) );
  XOR2_X1 U11037 ( .A(n11161), .B(n11162), .Z(n11160) );
  XOR2_X1 U11038 ( .A(n11163), .B(n11164), .Z(n10957) );
  XOR2_X1 U11039 ( .A(n11165), .B(n11166), .Z(n11164) );
  OR2_X1 U11040 ( .A1(n8918), .A2(n8140), .ZN(n10963) );
  XNOR2_X1 U11041 ( .A(n11167), .B(n11168), .ZN(n10960) );
  XNOR2_X1 U11042 ( .A(n11169), .B(n11170), .ZN(n11167) );
  OR2_X1 U11043 ( .A1(n8914), .A2(n8140), .ZN(n10967) );
  XOR2_X1 U11044 ( .A(n11171), .B(n11172), .Z(n10964) );
  XOR2_X1 U11045 ( .A(n11173), .B(n11174), .Z(n11172) );
  OR2_X1 U11046 ( .A1(n8910), .A2(n8140), .ZN(n10971) );
  XOR2_X1 U11047 ( .A(n11175), .B(n11176), .Z(n10968) );
  XOR2_X1 U11048 ( .A(n11177), .B(n11178), .Z(n11176) );
  OR2_X1 U11049 ( .A1(n8906), .A2(n8140), .ZN(n10975) );
  XOR2_X1 U11050 ( .A(n11179), .B(n11180), .Z(n10972) );
  XOR2_X1 U11051 ( .A(n11181), .B(n11182), .Z(n11180) );
  OR2_X1 U11052 ( .A1(n8902), .A2(n8140), .ZN(n10979) );
  XOR2_X1 U11053 ( .A(n11183), .B(n11184), .Z(n10976) );
  XOR2_X1 U11054 ( .A(n11185), .B(n11186), .Z(n11184) );
  XOR2_X1 U11055 ( .A(n10760), .B(n11187), .Z(n10753) );
  XOR2_X1 U11056 ( .A(n10759), .B(n10758), .Z(n11187) );
  OR2_X1 U11057 ( .A1(n8902), .A2(n8168), .ZN(n10758) );
  OR2_X1 U11058 ( .A1(n11188), .A2(n11189), .ZN(n10759) );
  AND2_X1 U11059 ( .A1(n11186), .A2(n11185), .ZN(n11189) );
  AND2_X1 U11060 ( .A1(n11183), .A2(n11190), .ZN(n11188) );
  OR2_X1 U11061 ( .A1(n11186), .A2(n11185), .ZN(n11190) );
  OR2_X1 U11062 ( .A1(n11191), .A2(n11192), .ZN(n11185) );
  AND2_X1 U11063 ( .A1(n11182), .A2(n11181), .ZN(n11192) );
  AND2_X1 U11064 ( .A1(n11179), .A2(n11193), .ZN(n11191) );
  OR2_X1 U11065 ( .A1(n11182), .A2(n11181), .ZN(n11193) );
  OR2_X1 U11066 ( .A1(n11194), .A2(n11195), .ZN(n11181) );
  AND2_X1 U11067 ( .A1(n11178), .A2(n11177), .ZN(n11195) );
  AND2_X1 U11068 ( .A1(n11175), .A2(n11196), .ZN(n11194) );
  OR2_X1 U11069 ( .A1(n11178), .A2(n11177), .ZN(n11196) );
  OR2_X1 U11070 ( .A1(n11197), .A2(n11198), .ZN(n11177) );
  AND2_X1 U11071 ( .A1(n11174), .A2(n11173), .ZN(n11198) );
  AND2_X1 U11072 ( .A1(n11171), .A2(n11199), .ZN(n11197) );
  OR2_X1 U11073 ( .A1(n11174), .A2(n11173), .ZN(n11199) );
  OR2_X1 U11074 ( .A1(n11200), .A2(n11201), .ZN(n11173) );
  AND2_X1 U11075 ( .A1(n11170), .A2(n11169), .ZN(n11201) );
  AND2_X1 U11076 ( .A1(n11168), .A2(n11202), .ZN(n11200) );
  OR2_X1 U11077 ( .A1(n11170), .A2(n11169), .ZN(n11202) );
  OR2_X1 U11078 ( .A1(n8922), .A2(n8168), .ZN(n11169) );
  OR2_X1 U11079 ( .A1(n11203), .A2(n11204), .ZN(n11170) );
  AND2_X1 U11080 ( .A1(n11166), .A2(n11165), .ZN(n11204) );
  AND2_X1 U11081 ( .A1(n11163), .A2(n11205), .ZN(n11203) );
  OR2_X1 U11082 ( .A1(n11166), .A2(n11165), .ZN(n11205) );
  OR2_X1 U11083 ( .A1(n11206), .A2(n11207), .ZN(n11165) );
  AND2_X1 U11084 ( .A1(n11162), .A2(n11161), .ZN(n11207) );
  AND2_X1 U11085 ( .A1(n11159), .A2(n11208), .ZN(n11206) );
  OR2_X1 U11086 ( .A1(n11162), .A2(n11161), .ZN(n11208) );
  OR2_X1 U11087 ( .A1(n11209), .A2(n11210), .ZN(n11161) );
  AND2_X1 U11088 ( .A1(n11158), .A2(n11157), .ZN(n11210) );
  AND2_X1 U11089 ( .A1(n11155), .A2(n11211), .ZN(n11209) );
  OR2_X1 U11090 ( .A1(n11158), .A2(n11157), .ZN(n11211) );
  OR2_X1 U11091 ( .A1(n11212), .A2(n11213), .ZN(n11157) );
  AND2_X1 U11092 ( .A1(n11154), .A2(n11153), .ZN(n11213) );
  AND2_X1 U11093 ( .A1(n11152), .A2(n11214), .ZN(n11212) );
  OR2_X1 U11094 ( .A1(n11154), .A2(n11153), .ZN(n11214) );
  OR2_X1 U11095 ( .A1(n8938), .A2(n8168), .ZN(n11153) );
  OR2_X1 U11096 ( .A1(n11215), .A2(n11216), .ZN(n11154) );
  AND2_X1 U11097 ( .A1(n11150), .A2(n11149), .ZN(n11216) );
  AND2_X1 U11098 ( .A1(n11147), .A2(n11217), .ZN(n11215) );
  OR2_X1 U11099 ( .A1(n11150), .A2(n11149), .ZN(n11217) );
  OR2_X1 U11100 ( .A1(n11218), .A2(n11219), .ZN(n11149) );
  AND2_X1 U11101 ( .A1(n11146), .A2(n11145), .ZN(n11219) );
  AND2_X1 U11102 ( .A1(n11143), .A2(n11220), .ZN(n11218) );
  OR2_X1 U11103 ( .A1(n11146), .A2(n11145), .ZN(n11220) );
  OR2_X1 U11104 ( .A1(n11221), .A2(n11222), .ZN(n11145) );
  AND2_X1 U11105 ( .A1(n11142), .A2(n11141), .ZN(n11222) );
  AND2_X1 U11106 ( .A1(n11139), .A2(n11223), .ZN(n11221) );
  OR2_X1 U11107 ( .A1(n11142), .A2(n11141), .ZN(n11223) );
  OR2_X1 U11108 ( .A1(n11224), .A2(n11225), .ZN(n11141) );
  AND2_X1 U11109 ( .A1(n11138), .A2(n11137), .ZN(n11225) );
  AND2_X1 U11110 ( .A1(n11135), .A2(n11226), .ZN(n11224) );
  OR2_X1 U11111 ( .A1(n11138), .A2(n11137), .ZN(n11226) );
  OR2_X1 U11112 ( .A1(n11227), .A2(n11228), .ZN(n11137) );
  AND2_X1 U11113 ( .A1(n11134), .A2(n11133), .ZN(n11228) );
  AND2_X1 U11114 ( .A1(n11131), .A2(n11229), .ZN(n11227) );
  OR2_X1 U11115 ( .A1(n11134), .A2(n11133), .ZN(n11229) );
  OR2_X1 U11116 ( .A1(n11230), .A2(n11231), .ZN(n11133) );
  AND2_X1 U11117 ( .A1(n11130), .A2(n11129), .ZN(n11231) );
  AND2_X1 U11118 ( .A1(n11127), .A2(n11232), .ZN(n11230) );
  OR2_X1 U11119 ( .A1(n11130), .A2(n11129), .ZN(n11232) );
  OR2_X1 U11120 ( .A1(n11233), .A2(n11234), .ZN(n11129) );
  AND2_X1 U11121 ( .A1(n11126), .A2(n11125), .ZN(n11234) );
  AND2_X1 U11122 ( .A1(n11123), .A2(n11235), .ZN(n11233) );
  OR2_X1 U11123 ( .A1(n11126), .A2(n11125), .ZN(n11235) );
  OR2_X1 U11124 ( .A1(n11236), .A2(n11237), .ZN(n11125) );
  AND2_X1 U11125 ( .A1(n11122), .A2(n11121), .ZN(n11237) );
  AND2_X1 U11126 ( .A1(n11119), .A2(n11238), .ZN(n11236) );
  OR2_X1 U11127 ( .A1(n11122), .A2(n11121), .ZN(n11238) );
  OR2_X1 U11128 ( .A1(n11239), .A2(n11240), .ZN(n11121) );
  AND2_X1 U11129 ( .A1(n11118), .A2(n11117), .ZN(n11240) );
  AND2_X1 U11130 ( .A1(n11115), .A2(n11241), .ZN(n11239) );
  OR2_X1 U11131 ( .A1(n11118), .A2(n11117), .ZN(n11241) );
  OR2_X1 U11132 ( .A1(n11242), .A2(n11243), .ZN(n11117) );
  AND2_X1 U11133 ( .A1(n11114), .A2(n11113), .ZN(n11243) );
  AND2_X1 U11134 ( .A1(n11111), .A2(n11244), .ZN(n11242) );
  OR2_X1 U11135 ( .A1(n11114), .A2(n11113), .ZN(n11244) );
  OR2_X1 U11136 ( .A1(n11245), .A2(n11246), .ZN(n11113) );
  AND2_X1 U11137 ( .A1(n11110), .A2(n11109), .ZN(n11246) );
  AND2_X1 U11138 ( .A1(n11107), .A2(n11247), .ZN(n11245) );
  OR2_X1 U11139 ( .A1(n11110), .A2(n11109), .ZN(n11247) );
  OR2_X1 U11140 ( .A1(n11248), .A2(n11249), .ZN(n11109) );
  AND2_X1 U11141 ( .A1(n11106), .A2(n11105), .ZN(n11249) );
  AND2_X1 U11142 ( .A1(n11103), .A2(n11250), .ZN(n11248) );
  OR2_X1 U11143 ( .A1(n11106), .A2(n11105), .ZN(n11250) );
  OR2_X1 U11144 ( .A1(n11251), .A2(n11252), .ZN(n11105) );
  AND2_X1 U11145 ( .A1(n11102), .A2(n11101), .ZN(n11252) );
  AND2_X1 U11146 ( .A1(n11099), .A2(n11253), .ZN(n11251) );
  OR2_X1 U11147 ( .A1(n11102), .A2(n11101), .ZN(n11253) );
  OR2_X1 U11148 ( .A1(n11254), .A2(n11255), .ZN(n11101) );
  AND2_X1 U11149 ( .A1(n11098), .A2(n11097), .ZN(n11255) );
  AND2_X1 U11150 ( .A1(n11095), .A2(n11256), .ZN(n11254) );
  OR2_X1 U11151 ( .A1(n11098), .A2(n11097), .ZN(n11256) );
  OR2_X1 U11152 ( .A1(n11257), .A2(n11258), .ZN(n11097) );
  AND2_X1 U11153 ( .A1(n8999), .A2(n11094), .ZN(n11258) );
  AND2_X1 U11154 ( .A1(n11092), .A2(n11259), .ZN(n11257) );
  OR2_X1 U11155 ( .A1(n8999), .A2(n11094), .ZN(n11259) );
  OR2_X1 U11156 ( .A1(n11260), .A2(n11261), .ZN(n11094) );
  AND2_X1 U11157 ( .A1(n11091), .A2(n11090), .ZN(n11261) );
  AND2_X1 U11158 ( .A1(n11088), .A2(n11262), .ZN(n11260) );
  OR2_X1 U11159 ( .A1(n11091), .A2(n11090), .ZN(n11262) );
  OR2_X1 U11160 ( .A1(n11263), .A2(n11264), .ZN(n11090) );
  AND2_X1 U11161 ( .A1(n11087), .A2(n11086), .ZN(n11264) );
  AND2_X1 U11162 ( .A1(n11084), .A2(n11265), .ZN(n11263) );
  OR2_X1 U11163 ( .A1(n11087), .A2(n11086), .ZN(n11265) );
  OR2_X1 U11164 ( .A1(n11266), .A2(n11267), .ZN(n11086) );
  AND2_X1 U11165 ( .A1(n11083), .A2(n11082), .ZN(n11267) );
  AND2_X1 U11166 ( .A1(n11080), .A2(n11268), .ZN(n11266) );
  OR2_X1 U11167 ( .A1(n11083), .A2(n11082), .ZN(n11268) );
  OR2_X1 U11168 ( .A1(n11269), .A2(n11270), .ZN(n11082) );
  AND2_X1 U11169 ( .A1(n11077), .A2(n11078), .ZN(n11270) );
  AND2_X1 U11170 ( .A1(n11271), .A2(n11272), .ZN(n11269) );
  OR2_X1 U11171 ( .A1(n11077), .A2(n11078), .ZN(n11272) );
  OR2_X1 U11172 ( .A1(n9984), .A2(n11273), .ZN(n11078) );
  OR2_X1 U11173 ( .A1(n8168), .A2(n8196), .ZN(n11273) );
  OR2_X1 U11174 ( .A1(n9014), .A2(n8168), .ZN(n11077) );
  INV_X1 U11175 ( .A(n11079), .ZN(n11271) );
  OR2_X1 U11176 ( .A1(n11274), .A2(n11275), .ZN(n11079) );
  AND2_X1 U11177 ( .A1(b_24_), .A2(n11276), .ZN(n11275) );
  OR2_X1 U11178 ( .A1(n11277), .A2(n9989), .ZN(n11276) );
  AND2_X1 U11179 ( .A1(a_30_), .A2(n8224), .ZN(n11277) );
  AND2_X1 U11180 ( .A1(b_23_), .A2(n11278), .ZN(n11274) );
  OR2_X1 U11181 ( .A1(n11279), .A2(n8021), .ZN(n11278) );
  AND2_X1 U11182 ( .A1(a_31_), .A2(n8196), .ZN(n11279) );
  OR2_X1 U11183 ( .A1(n9010), .A2(n8168), .ZN(n11083) );
  XOR2_X1 U11184 ( .A(n11280), .B(n11281), .Z(n11080) );
  XNOR2_X1 U11185 ( .A(n11282), .B(n11283), .ZN(n11280) );
  OR2_X1 U11186 ( .A1(n9006), .A2(n8168), .ZN(n11087) );
  XOR2_X1 U11187 ( .A(n11284), .B(n11285), .Z(n11084) );
  XOR2_X1 U11188 ( .A(n11286), .B(n11287), .Z(n11285) );
  OR2_X1 U11189 ( .A1(n9002), .A2(n8168), .ZN(n11091) );
  XOR2_X1 U11190 ( .A(n11288), .B(n11289), .Z(n11088) );
  XOR2_X1 U11191 ( .A(n11290), .B(n11291), .Z(n11289) );
  OR2_X1 U11192 ( .A1(n8998), .A2(n8168), .ZN(n8999) );
  XOR2_X1 U11193 ( .A(n11292), .B(n11293), .Z(n11092) );
  XOR2_X1 U11194 ( .A(n11294), .B(n11295), .Z(n11293) );
  OR2_X1 U11195 ( .A1(n8994), .A2(n8168), .ZN(n11098) );
  XOR2_X1 U11196 ( .A(n11296), .B(n11297), .Z(n11095) );
  XOR2_X1 U11197 ( .A(n11298), .B(n11299), .Z(n11297) );
  OR2_X1 U11198 ( .A1(n8990), .A2(n8168), .ZN(n11102) );
  XOR2_X1 U11199 ( .A(n11300), .B(n11301), .Z(n11099) );
  XOR2_X1 U11200 ( .A(n11302), .B(n8995), .Z(n11301) );
  OR2_X1 U11201 ( .A1(n8986), .A2(n8168), .ZN(n11106) );
  XOR2_X1 U11202 ( .A(n11303), .B(n11304), .Z(n11103) );
  XOR2_X1 U11203 ( .A(n11305), .B(n11306), .Z(n11304) );
  OR2_X1 U11204 ( .A1(n8982), .A2(n8168), .ZN(n11110) );
  XOR2_X1 U11205 ( .A(n11307), .B(n11308), .Z(n11107) );
  XOR2_X1 U11206 ( .A(n11309), .B(n11310), .Z(n11308) );
  OR2_X1 U11207 ( .A1(n8978), .A2(n8168), .ZN(n11114) );
  XOR2_X1 U11208 ( .A(n11311), .B(n11312), .Z(n11111) );
  XOR2_X1 U11209 ( .A(n11313), .B(n11314), .Z(n11312) );
  OR2_X1 U11210 ( .A1(n8974), .A2(n8168), .ZN(n11118) );
  XOR2_X1 U11211 ( .A(n11315), .B(n11316), .Z(n11115) );
  XOR2_X1 U11212 ( .A(n11317), .B(n11318), .Z(n11316) );
  OR2_X1 U11213 ( .A1(n8970), .A2(n8168), .ZN(n11122) );
  XOR2_X1 U11214 ( .A(n11319), .B(n11320), .Z(n11119) );
  XOR2_X1 U11215 ( .A(n11321), .B(n11322), .Z(n11320) );
  OR2_X1 U11216 ( .A1(n8966), .A2(n8168), .ZN(n11126) );
  XOR2_X1 U11217 ( .A(n11323), .B(n11324), .Z(n11123) );
  XOR2_X1 U11218 ( .A(n11325), .B(n11326), .Z(n11324) );
  OR2_X1 U11219 ( .A1(n8962), .A2(n8168), .ZN(n11130) );
  XOR2_X1 U11220 ( .A(n11327), .B(n11328), .Z(n11127) );
  XOR2_X1 U11221 ( .A(n11329), .B(n11330), .Z(n11328) );
  OR2_X1 U11222 ( .A1(n8958), .A2(n8168), .ZN(n11134) );
  XOR2_X1 U11223 ( .A(n11331), .B(n11332), .Z(n11131) );
  XOR2_X1 U11224 ( .A(n11333), .B(n11334), .Z(n11332) );
  OR2_X1 U11225 ( .A1(n8954), .A2(n8168), .ZN(n11138) );
  XOR2_X1 U11226 ( .A(n11335), .B(n11336), .Z(n11135) );
  XOR2_X1 U11227 ( .A(n11337), .B(n11338), .Z(n11336) );
  OR2_X1 U11228 ( .A1(n8950), .A2(n8168), .ZN(n11142) );
  XOR2_X1 U11229 ( .A(n11339), .B(n11340), .Z(n11139) );
  XOR2_X1 U11230 ( .A(n11341), .B(n11342), .Z(n11340) );
  OR2_X1 U11231 ( .A1(n8946), .A2(n8168), .ZN(n11146) );
  XOR2_X1 U11232 ( .A(n11343), .B(n11344), .Z(n11143) );
  XOR2_X1 U11233 ( .A(n11345), .B(n11346), .Z(n11344) );
  OR2_X1 U11234 ( .A1(n8942), .A2(n8168), .ZN(n11150) );
  XOR2_X1 U11235 ( .A(n11347), .B(n11348), .Z(n11147) );
  XOR2_X1 U11236 ( .A(n11349), .B(n11350), .Z(n11348) );
  XOR2_X1 U11237 ( .A(n11351), .B(n11352), .Z(n11152) );
  XOR2_X1 U11238 ( .A(n11353), .B(n11354), .Z(n11352) );
  OR2_X1 U11239 ( .A1(n8934), .A2(n8168), .ZN(n11158) );
  XNOR2_X1 U11240 ( .A(n11355), .B(n11356), .ZN(n11155) );
  XNOR2_X1 U11241 ( .A(n11357), .B(n11358), .ZN(n11355) );
  OR2_X1 U11242 ( .A1(n8930), .A2(n8168), .ZN(n11162) );
  XOR2_X1 U11243 ( .A(n11359), .B(n11360), .Z(n11159) );
  XOR2_X1 U11244 ( .A(n11361), .B(n11362), .Z(n11360) );
  OR2_X1 U11245 ( .A1(n8926), .A2(n8168), .ZN(n11166) );
  XOR2_X1 U11246 ( .A(n11363), .B(n11364), .Z(n11163) );
  XOR2_X1 U11247 ( .A(n11365), .B(n11366), .Z(n11364) );
  XOR2_X1 U11248 ( .A(n11367), .B(n11368), .Z(n11168) );
  XOR2_X1 U11249 ( .A(n11369), .B(n11370), .Z(n11368) );
  OR2_X1 U11250 ( .A1(n8918), .A2(n8168), .ZN(n11174) );
  XNOR2_X1 U11251 ( .A(n11371), .B(n11372), .ZN(n11171) );
  XNOR2_X1 U11252 ( .A(n11373), .B(n11374), .ZN(n11371) );
  OR2_X1 U11253 ( .A1(n8914), .A2(n8168), .ZN(n11178) );
  XOR2_X1 U11254 ( .A(n11375), .B(n11376), .Z(n11175) );
  XOR2_X1 U11255 ( .A(n11377), .B(n11378), .Z(n11376) );
  OR2_X1 U11256 ( .A1(n8910), .A2(n8168), .ZN(n11182) );
  XOR2_X1 U11257 ( .A(n11379), .B(n11380), .Z(n11179) );
  XOR2_X1 U11258 ( .A(n11381), .B(n11382), .Z(n11380) );
  OR2_X1 U11259 ( .A1(n8906), .A2(n8168), .ZN(n11186) );
  XNOR2_X1 U11260 ( .A(n11383), .B(n11384), .ZN(n11183) );
  XNOR2_X1 U11261 ( .A(n11385), .B(n11386), .ZN(n11383) );
  XOR2_X1 U11262 ( .A(n11387), .B(n11388), .Z(n10760) );
  XOR2_X1 U11263 ( .A(n11389), .B(n11390), .Z(n11388) );
  OR2_X1 U11264 ( .A1(n9820), .A2(n9819), .ZN(n9088) );
  INV_X1 U11265 ( .A(n11391), .ZN(n9819) );
  OR2_X1 U11266 ( .A1(n11392), .A2(n11393), .ZN(n11391) );
  AND2_X1 U11267 ( .A1(n11394), .A2(n11395), .ZN(n11392) );
  AND2_X1 U11268 ( .A1(n9824), .A2(n11396), .ZN(n9820) );
  INV_X1 U11269 ( .A(n9825), .ZN(n11396) );
  OR2_X1 U11270 ( .A1(n11397), .A2(n11398), .ZN(n9825) );
  AND2_X1 U11271 ( .A1(n9844), .A2(n9843), .ZN(n11398) );
  AND2_X1 U11272 ( .A1(n9841), .A2(n11399), .ZN(n11397) );
  OR2_X1 U11273 ( .A1(n9843), .A2(n9844), .ZN(n11399) );
  OR2_X1 U11274 ( .A1(n9297), .A2(n8196), .ZN(n9844) );
  OR2_X1 U11275 ( .A1(n11400), .A2(n11401), .ZN(n9843) );
  AND2_X1 U11276 ( .A1(n10765), .A2(n10764), .ZN(n11401) );
  AND2_X1 U11277 ( .A1(n10763), .A2(n11402), .ZN(n11400) );
  OR2_X1 U11278 ( .A1(n10764), .A2(n10765), .ZN(n11402) );
  OR2_X1 U11279 ( .A1(n11403), .A2(n11404), .ZN(n10765) );
  AND2_X1 U11280 ( .A1(n11390), .A2(n11389), .ZN(n11404) );
  AND2_X1 U11281 ( .A1(n11387), .A2(n11405), .ZN(n11403) );
  OR2_X1 U11282 ( .A1(n11389), .A2(n11390), .ZN(n11405) );
  OR2_X1 U11283 ( .A1(n8906), .A2(n8196), .ZN(n11390) );
  OR2_X1 U11284 ( .A1(n11406), .A2(n11407), .ZN(n11389) );
  AND2_X1 U11285 ( .A1(n11386), .A2(n11385), .ZN(n11407) );
  AND2_X1 U11286 ( .A1(n11384), .A2(n11408), .ZN(n11406) );
  OR2_X1 U11287 ( .A1(n11385), .A2(n11386), .ZN(n11408) );
  OR2_X1 U11288 ( .A1(n11409), .A2(n11410), .ZN(n11386) );
  AND2_X1 U11289 ( .A1(n11382), .A2(n11381), .ZN(n11410) );
  AND2_X1 U11290 ( .A1(n11379), .A2(n11411), .ZN(n11409) );
  OR2_X1 U11291 ( .A1(n11381), .A2(n11382), .ZN(n11411) );
  OR2_X1 U11292 ( .A1(n8914), .A2(n8196), .ZN(n11382) );
  OR2_X1 U11293 ( .A1(n11412), .A2(n11413), .ZN(n11381) );
  AND2_X1 U11294 ( .A1(n11378), .A2(n11377), .ZN(n11413) );
  AND2_X1 U11295 ( .A1(n11375), .A2(n11414), .ZN(n11412) );
  OR2_X1 U11296 ( .A1(n11377), .A2(n11378), .ZN(n11414) );
  OR2_X1 U11297 ( .A1(n8918), .A2(n8196), .ZN(n11378) );
  OR2_X1 U11298 ( .A1(n11415), .A2(n11416), .ZN(n11377) );
  AND2_X1 U11299 ( .A1(n11374), .A2(n11373), .ZN(n11416) );
  AND2_X1 U11300 ( .A1(n11372), .A2(n11417), .ZN(n11415) );
  OR2_X1 U11301 ( .A1(n11373), .A2(n11374), .ZN(n11417) );
  OR2_X1 U11302 ( .A1(n11418), .A2(n11419), .ZN(n11374) );
  AND2_X1 U11303 ( .A1(n11370), .A2(n11369), .ZN(n11419) );
  AND2_X1 U11304 ( .A1(n11367), .A2(n11420), .ZN(n11418) );
  OR2_X1 U11305 ( .A1(n11369), .A2(n11370), .ZN(n11420) );
  OR2_X1 U11306 ( .A1(n8926), .A2(n8196), .ZN(n11370) );
  OR2_X1 U11307 ( .A1(n11421), .A2(n11422), .ZN(n11369) );
  AND2_X1 U11308 ( .A1(n11366), .A2(n11365), .ZN(n11422) );
  AND2_X1 U11309 ( .A1(n11363), .A2(n11423), .ZN(n11421) );
  OR2_X1 U11310 ( .A1(n11365), .A2(n11366), .ZN(n11423) );
  OR2_X1 U11311 ( .A1(n8930), .A2(n8196), .ZN(n11366) );
  OR2_X1 U11312 ( .A1(n11424), .A2(n11425), .ZN(n11365) );
  AND2_X1 U11313 ( .A1(n11362), .A2(n11361), .ZN(n11425) );
  AND2_X1 U11314 ( .A1(n11359), .A2(n11426), .ZN(n11424) );
  OR2_X1 U11315 ( .A1(n11361), .A2(n11362), .ZN(n11426) );
  OR2_X1 U11316 ( .A1(n8934), .A2(n8196), .ZN(n11362) );
  OR2_X1 U11317 ( .A1(n11427), .A2(n11428), .ZN(n11361) );
  AND2_X1 U11318 ( .A1(n11358), .A2(n11357), .ZN(n11428) );
  AND2_X1 U11319 ( .A1(n11356), .A2(n11429), .ZN(n11427) );
  OR2_X1 U11320 ( .A1(n11357), .A2(n11358), .ZN(n11429) );
  OR2_X1 U11321 ( .A1(n11430), .A2(n11431), .ZN(n11358) );
  AND2_X1 U11322 ( .A1(n11354), .A2(n11353), .ZN(n11431) );
  AND2_X1 U11323 ( .A1(n11351), .A2(n11432), .ZN(n11430) );
  OR2_X1 U11324 ( .A1(n11353), .A2(n11354), .ZN(n11432) );
  OR2_X1 U11325 ( .A1(n8942), .A2(n8196), .ZN(n11354) );
  OR2_X1 U11326 ( .A1(n11433), .A2(n11434), .ZN(n11353) );
  AND2_X1 U11327 ( .A1(n11350), .A2(n11349), .ZN(n11434) );
  AND2_X1 U11328 ( .A1(n11347), .A2(n11435), .ZN(n11433) );
  OR2_X1 U11329 ( .A1(n11349), .A2(n11350), .ZN(n11435) );
  OR2_X1 U11330 ( .A1(n8946), .A2(n8196), .ZN(n11350) );
  OR2_X1 U11331 ( .A1(n11436), .A2(n11437), .ZN(n11349) );
  AND2_X1 U11332 ( .A1(n11346), .A2(n11345), .ZN(n11437) );
  AND2_X1 U11333 ( .A1(n11343), .A2(n11438), .ZN(n11436) );
  OR2_X1 U11334 ( .A1(n11345), .A2(n11346), .ZN(n11438) );
  OR2_X1 U11335 ( .A1(n8950), .A2(n8196), .ZN(n11346) );
  OR2_X1 U11336 ( .A1(n11439), .A2(n11440), .ZN(n11345) );
  AND2_X1 U11337 ( .A1(n11342), .A2(n11341), .ZN(n11440) );
  AND2_X1 U11338 ( .A1(n11339), .A2(n11441), .ZN(n11439) );
  OR2_X1 U11339 ( .A1(n11341), .A2(n11342), .ZN(n11441) );
  OR2_X1 U11340 ( .A1(n8954), .A2(n8196), .ZN(n11342) );
  OR2_X1 U11341 ( .A1(n11442), .A2(n11443), .ZN(n11341) );
  AND2_X1 U11342 ( .A1(n11338), .A2(n11337), .ZN(n11443) );
  AND2_X1 U11343 ( .A1(n11335), .A2(n11444), .ZN(n11442) );
  OR2_X1 U11344 ( .A1(n11337), .A2(n11338), .ZN(n11444) );
  OR2_X1 U11345 ( .A1(n8958), .A2(n8196), .ZN(n11338) );
  OR2_X1 U11346 ( .A1(n11445), .A2(n11446), .ZN(n11337) );
  AND2_X1 U11347 ( .A1(n11334), .A2(n11333), .ZN(n11446) );
  AND2_X1 U11348 ( .A1(n11331), .A2(n11447), .ZN(n11445) );
  OR2_X1 U11349 ( .A1(n11333), .A2(n11334), .ZN(n11447) );
  OR2_X1 U11350 ( .A1(n8962), .A2(n8196), .ZN(n11334) );
  OR2_X1 U11351 ( .A1(n11448), .A2(n11449), .ZN(n11333) );
  AND2_X1 U11352 ( .A1(n11330), .A2(n11329), .ZN(n11449) );
  AND2_X1 U11353 ( .A1(n11327), .A2(n11450), .ZN(n11448) );
  OR2_X1 U11354 ( .A1(n11329), .A2(n11330), .ZN(n11450) );
  OR2_X1 U11355 ( .A1(n8966), .A2(n8196), .ZN(n11330) );
  OR2_X1 U11356 ( .A1(n11451), .A2(n11452), .ZN(n11329) );
  AND2_X1 U11357 ( .A1(n11326), .A2(n11325), .ZN(n11452) );
  AND2_X1 U11358 ( .A1(n11323), .A2(n11453), .ZN(n11451) );
  OR2_X1 U11359 ( .A1(n11325), .A2(n11326), .ZN(n11453) );
  OR2_X1 U11360 ( .A1(n8970), .A2(n8196), .ZN(n11326) );
  OR2_X1 U11361 ( .A1(n11454), .A2(n11455), .ZN(n11325) );
  AND2_X1 U11362 ( .A1(n11322), .A2(n11321), .ZN(n11455) );
  AND2_X1 U11363 ( .A1(n11319), .A2(n11456), .ZN(n11454) );
  OR2_X1 U11364 ( .A1(n11321), .A2(n11322), .ZN(n11456) );
  OR2_X1 U11365 ( .A1(n8974), .A2(n8196), .ZN(n11322) );
  OR2_X1 U11366 ( .A1(n11457), .A2(n11458), .ZN(n11321) );
  AND2_X1 U11367 ( .A1(n11318), .A2(n11317), .ZN(n11458) );
  AND2_X1 U11368 ( .A1(n11315), .A2(n11459), .ZN(n11457) );
  OR2_X1 U11369 ( .A1(n11317), .A2(n11318), .ZN(n11459) );
  OR2_X1 U11370 ( .A1(n8978), .A2(n8196), .ZN(n11318) );
  OR2_X1 U11371 ( .A1(n11460), .A2(n11461), .ZN(n11317) );
  AND2_X1 U11372 ( .A1(n11314), .A2(n11313), .ZN(n11461) );
  AND2_X1 U11373 ( .A1(n11311), .A2(n11462), .ZN(n11460) );
  OR2_X1 U11374 ( .A1(n11313), .A2(n11314), .ZN(n11462) );
  OR2_X1 U11375 ( .A1(n8982), .A2(n8196), .ZN(n11314) );
  OR2_X1 U11376 ( .A1(n11463), .A2(n11464), .ZN(n11313) );
  AND2_X1 U11377 ( .A1(n11310), .A2(n11309), .ZN(n11464) );
  AND2_X1 U11378 ( .A1(n11307), .A2(n11465), .ZN(n11463) );
  OR2_X1 U11379 ( .A1(n11309), .A2(n11310), .ZN(n11465) );
  OR2_X1 U11380 ( .A1(n8986), .A2(n8196), .ZN(n11310) );
  OR2_X1 U11381 ( .A1(n11466), .A2(n11467), .ZN(n11309) );
  AND2_X1 U11382 ( .A1(n11306), .A2(n11305), .ZN(n11467) );
  AND2_X1 U11383 ( .A1(n11303), .A2(n11468), .ZN(n11466) );
  OR2_X1 U11384 ( .A1(n11305), .A2(n11306), .ZN(n11468) );
  OR2_X1 U11385 ( .A1(n8990), .A2(n8196), .ZN(n11306) );
  OR2_X1 U11386 ( .A1(n11469), .A2(n11470), .ZN(n11305) );
  AND2_X1 U11387 ( .A1(n8995), .A2(n11302), .ZN(n11470) );
  AND2_X1 U11388 ( .A1(n11300), .A2(n11471), .ZN(n11469) );
  OR2_X1 U11389 ( .A1(n11302), .A2(n8995), .ZN(n11471) );
  OR2_X1 U11390 ( .A1(n8994), .A2(n8196), .ZN(n8995) );
  OR2_X1 U11391 ( .A1(n11472), .A2(n11473), .ZN(n11302) );
  AND2_X1 U11392 ( .A1(n11299), .A2(n11298), .ZN(n11473) );
  AND2_X1 U11393 ( .A1(n11296), .A2(n11474), .ZN(n11472) );
  OR2_X1 U11394 ( .A1(n11298), .A2(n11299), .ZN(n11474) );
  OR2_X1 U11395 ( .A1(n8998), .A2(n8196), .ZN(n11299) );
  OR2_X1 U11396 ( .A1(n11475), .A2(n11476), .ZN(n11298) );
  AND2_X1 U11397 ( .A1(n11295), .A2(n11294), .ZN(n11476) );
  AND2_X1 U11398 ( .A1(n11292), .A2(n11477), .ZN(n11475) );
  OR2_X1 U11399 ( .A1(n11294), .A2(n11295), .ZN(n11477) );
  OR2_X1 U11400 ( .A1(n9002), .A2(n8196), .ZN(n11295) );
  OR2_X1 U11401 ( .A1(n11478), .A2(n11479), .ZN(n11294) );
  AND2_X1 U11402 ( .A1(n11291), .A2(n11290), .ZN(n11479) );
  AND2_X1 U11403 ( .A1(n11288), .A2(n11480), .ZN(n11478) );
  OR2_X1 U11404 ( .A1(n11290), .A2(n11291), .ZN(n11480) );
  OR2_X1 U11405 ( .A1(n9006), .A2(n8196), .ZN(n11291) );
  OR2_X1 U11406 ( .A1(n11481), .A2(n11482), .ZN(n11290) );
  AND2_X1 U11407 ( .A1(n11287), .A2(n11286), .ZN(n11482) );
  AND2_X1 U11408 ( .A1(n11284), .A2(n11483), .ZN(n11481) );
  OR2_X1 U11409 ( .A1(n11286), .A2(n11287), .ZN(n11483) );
  OR2_X1 U11410 ( .A1(n9010), .A2(n8196), .ZN(n11287) );
  OR2_X1 U11411 ( .A1(n11484), .A2(n11485), .ZN(n11286) );
  AND2_X1 U11412 ( .A1(n11281), .A2(n11282), .ZN(n11485) );
  AND2_X1 U11413 ( .A1(n11486), .A2(n11487), .ZN(n11484) );
  OR2_X1 U11414 ( .A1(n11282), .A2(n11281), .ZN(n11487) );
  OR2_X1 U11415 ( .A1(n9014), .A2(n8196), .ZN(n11281) );
  OR2_X1 U11416 ( .A1(n9984), .A2(n11488), .ZN(n11282) );
  OR2_X1 U11417 ( .A1(n8196), .A2(n8224), .ZN(n11488) );
  INV_X1 U11418 ( .A(n11283), .ZN(n11486) );
  OR2_X1 U11419 ( .A1(n11489), .A2(n11490), .ZN(n11283) );
  AND2_X1 U11420 ( .A1(b_23_), .A2(n11491), .ZN(n11490) );
  OR2_X1 U11421 ( .A1(n11492), .A2(n9989), .ZN(n11491) );
  AND2_X1 U11422 ( .A1(a_30_), .A2(n8252), .ZN(n11492) );
  AND2_X1 U11423 ( .A1(b_22_), .A2(n11493), .ZN(n11489) );
  OR2_X1 U11424 ( .A1(n11494), .A2(n8021), .ZN(n11493) );
  AND2_X1 U11425 ( .A1(a_31_), .A2(n8224), .ZN(n11494) );
  XOR2_X1 U11426 ( .A(n11495), .B(n11496), .Z(n11284) );
  XNOR2_X1 U11427 ( .A(n11497), .B(n11498), .ZN(n11495) );
  XOR2_X1 U11428 ( .A(n11499), .B(n11500), .Z(n11288) );
  XOR2_X1 U11429 ( .A(n11501), .B(n11502), .Z(n11500) );
  XOR2_X1 U11430 ( .A(n11503), .B(n11504), .Z(n11292) );
  XOR2_X1 U11431 ( .A(n11505), .B(n11506), .Z(n11504) );
  XOR2_X1 U11432 ( .A(n11507), .B(n11508), .Z(n11296) );
  XOR2_X1 U11433 ( .A(n11509), .B(n11510), .Z(n11508) );
  XOR2_X1 U11434 ( .A(n11511), .B(n11512), .Z(n11300) );
  XOR2_X1 U11435 ( .A(n11513), .B(n11514), .Z(n11512) );
  XOR2_X1 U11436 ( .A(n11515), .B(n11516), .Z(n11303) );
  XOR2_X1 U11437 ( .A(n11517), .B(n11518), .Z(n11516) );
  XOR2_X1 U11438 ( .A(n11519), .B(n11520), .Z(n11307) );
  XOR2_X1 U11439 ( .A(n11521), .B(n8991), .Z(n11520) );
  XOR2_X1 U11440 ( .A(n11522), .B(n11523), .Z(n11311) );
  XOR2_X1 U11441 ( .A(n11524), .B(n11525), .Z(n11523) );
  XOR2_X1 U11442 ( .A(n11526), .B(n11527), .Z(n11315) );
  XOR2_X1 U11443 ( .A(n11528), .B(n11529), .Z(n11527) );
  XOR2_X1 U11444 ( .A(n11530), .B(n11531), .Z(n11319) );
  XOR2_X1 U11445 ( .A(n11532), .B(n11533), .Z(n11531) );
  XOR2_X1 U11446 ( .A(n11534), .B(n11535), .Z(n11323) );
  XOR2_X1 U11447 ( .A(n11536), .B(n11537), .Z(n11535) );
  XOR2_X1 U11448 ( .A(n11538), .B(n11539), .Z(n11327) );
  XOR2_X1 U11449 ( .A(n11540), .B(n11541), .Z(n11539) );
  XOR2_X1 U11450 ( .A(n11542), .B(n11543), .Z(n11331) );
  XOR2_X1 U11451 ( .A(n11544), .B(n11545), .Z(n11543) );
  XOR2_X1 U11452 ( .A(n11546), .B(n11547), .Z(n11335) );
  XOR2_X1 U11453 ( .A(n11548), .B(n11549), .Z(n11547) );
  XOR2_X1 U11454 ( .A(n11550), .B(n11551), .Z(n11339) );
  XOR2_X1 U11455 ( .A(n11552), .B(n11553), .Z(n11551) );
  XNOR2_X1 U11456 ( .A(n11554), .B(n11555), .ZN(n11343) );
  XNOR2_X1 U11457 ( .A(n11556), .B(n11557), .ZN(n11554) );
  XOR2_X1 U11458 ( .A(n11558), .B(n11559), .Z(n11347) );
  XOR2_X1 U11459 ( .A(n11560), .B(n11561), .Z(n11559) );
  XOR2_X1 U11460 ( .A(n11562), .B(n11563), .Z(n11351) );
  XOR2_X1 U11461 ( .A(n11564), .B(n11565), .Z(n11563) );
  OR2_X1 U11462 ( .A1(n8938), .A2(n8196), .ZN(n11357) );
  XOR2_X1 U11463 ( .A(n11566), .B(n11567), .Z(n11356) );
  XOR2_X1 U11464 ( .A(n11568), .B(n11569), .Z(n11567) );
  XNOR2_X1 U11465 ( .A(n11570), .B(n11571), .ZN(n11359) );
  XNOR2_X1 U11466 ( .A(n11572), .B(n11573), .ZN(n11570) );
  XOR2_X1 U11467 ( .A(n11574), .B(n11575), .Z(n11363) );
  XOR2_X1 U11468 ( .A(n11576), .B(n11577), .Z(n11575) );
  XOR2_X1 U11469 ( .A(n11578), .B(n11579), .Z(n11367) );
  XOR2_X1 U11470 ( .A(n11580), .B(n11581), .Z(n11579) );
  OR2_X1 U11471 ( .A1(n8922), .A2(n8196), .ZN(n11373) );
  XOR2_X1 U11472 ( .A(n11582), .B(n11583), .Z(n11372) );
  XOR2_X1 U11473 ( .A(n11584), .B(n11585), .Z(n11583) );
  XNOR2_X1 U11474 ( .A(n11586), .B(n11587), .ZN(n11375) );
  XNOR2_X1 U11475 ( .A(n11588), .B(n11589), .ZN(n11586) );
  XOR2_X1 U11476 ( .A(n11590), .B(n11591), .Z(n11379) );
  XOR2_X1 U11477 ( .A(n11592), .B(n11593), .Z(n11591) );
  OR2_X1 U11478 ( .A1(n8910), .A2(n8196), .ZN(n11385) );
  XOR2_X1 U11479 ( .A(n11594), .B(n11595), .Z(n11384) );
  XOR2_X1 U11480 ( .A(n11596), .B(n11597), .Z(n11595) );
  XOR2_X1 U11481 ( .A(n11598), .B(n11599), .Z(n11387) );
  XOR2_X1 U11482 ( .A(n11600), .B(n11601), .Z(n11599) );
  OR2_X1 U11483 ( .A1(n8902), .A2(n8196), .ZN(n10764) );
  XOR2_X1 U11484 ( .A(n11602), .B(n11603), .Z(n10763) );
  XOR2_X1 U11485 ( .A(n11604), .B(n11605), .Z(n11603) );
  XOR2_X1 U11486 ( .A(n11606), .B(n11607), .Z(n9841) );
  XOR2_X1 U11487 ( .A(n11608), .B(n11609), .Z(n11607) );
  XNOR2_X1 U11488 ( .A(n11610), .B(n11611), .ZN(n9824) );
  XOR2_X1 U11489 ( .A(n11612), .B(n11613), .Z(n11611) );
  OR2_X1 U11490 ( .A1(n11393), .A2(n9099), .ZN(n9096) );
  AND2_X1 U11491 ( .A1(n11393), .A2(n9099), .ZN(n9816) );
  XNOR2_X1 U11492 ( .A(n11614), .B(n11615), .ZN(n9099) );
  INV_X1 U11493 ( .A(n9098), .ZN(n11393) );
  OR2_X1 U11494 ( .A1(n11394), .A2(n11395), .ZN(n9098) );
  OR2_X1 U11495 ( .A1(n11616), .A2(n11617), .ZN(n11395) );
  AND2_X1 U11496 ( .A1(n11610), .A2(n11613), .ZN(n11617) );
  AND2_X1 U11497 ( .A1(n11618), .A2(n11612), .ZN(n11616) );
  OR2_X1 U11498 ( .A1(n11619), .A2(n11620), .ZN(n11612) );
  AND2_X1 U11499 ( .A1(n11609), .A2(n11608), .ZN(n11620) );
  AND2_X1 U11500 ( .A1(n11606), .A2(n11621), .ZN(n11619) );
  OR2_X1 U11501 ( .A1(n11609), .A2(n11608), .ZN(n11621) );
  OR2_X1 U11502 ( .A1(n11622), .A2(n11623), .ZN(n11608) );
  AND2_X1 U11503 ( .A1(n11605), .A2(n11604), .ZN(n11623) );
  AND2_X1 U11504 ( .A1(n11602), .A2(n11624), .ZN(n11622) );
  OR2_X1 U11505 ( .A1(n11605), .A2(n11604), .ZN(n11624) );
  OR2_X1 U11506 ( .A1(n11625), .A2(n11626), .ZN(n11604) );
  AND2_X1 U11507 ( .A1(n11601), .A2(n11600), .ZN(n11626) );
  AND2_X1 U11508 ( .A1(n11598), .A2(n11627), .ZN(n11625) );
  OR2_X1 U11509 ( .A1(n11601), .A2(n11600), .ZN(n11627) );
  OR2_X1 U11510 ( .A1(n11628), .A2(n11629), .ZN(n11600) );
  AND2_X1 U11511 ( .A1(n11597), .A2(n11596), .ZN(n11629) );
  AND2_X1 U11512 ( .A1(n11594), .A2(n11630), .ZN(n11628) );
  OR2_X1 U11513 ( .A1(n11597), .A2(n11596), .ZN(n11630) );
  OR2_X1 U11514 ( .A1(n11631), .A2(n11632), .ZN(n11596) );
  AND2_X1 U11515 ( .A1(n11593), .A2(n11592), .ZN(n11632) );
  AND2_X1 U11516 ( .A1(n11590), .A2(n11633), .ZN(n11631) );
  OR2_X1 U11517 ( .A1(n11593), .A2(n11592), .ZN(n11633) );
  OR2_X1 U11518 ( .A1(n11634), .A2(n11635), .ZN(n11592) );
  AND2_X1 U11519 ( .A1(n11589), .A2(n11588), .ZN(n11635) );
  AND2_X1 U11520 ( .A1(n11587), .A2(n11636), .ZN(n11634) );
  OR2_X1 U11521 ( .A1(n11589), .A2(n11588), .ZN(n11636) );
  OR2_X1 U11522 ( .A1(n8922), .A2(n8224), .ZN(n11588) );
  OR2_X1 U11523 ( .A1(n11637), .A2(n11638), .ZN(n11589) );
  AND2_X1 U11524 ( .A1(n11585), .A2(n11584), .ZN(n11638) );
  AND2_X1 U11525 ( .A1(n11582), .A2(n11639), .ZN(n11637) );
  OR2_X1 U11526 ( .A1(n11585), .A2(n11584), .ZN(n11639) );
  OR2_X1 U11527 ( .A1(n11640), .A2(n11641), .ZN(n11584) );
  AND2_X1 U11528 ( .A1(n11581), .A2(n11580), .ZN(n11641) );
  AND2_X1 U11529 ( .A1(n11578), .A2(n11642), .ZN(n11640) );
  OR2_X1 U11530 ( .A1(n11581), .A2(n11580), .ZN(n11642) );
  OR2_X1 U11531 ( .A1(n11643), .A2(n11644), .ZN(n11580) );
  AND2_X1 U11532 ( .A1(n11577), .A2(n11576), .ZN(n11644) );
  AND2_X1 U11533 ( .A1(n11574), .A2(n11645), .ZN(n11643) );
  OR2_X1 U11534 ( .A1(n11577), .A2(n11576), .ZN(n11645) );
  OR2_X1 U11535 ( .A1(n11646), .A2(n11647), .ZN(n11576) );
  AND2_X1 U11536 ( .A1(n11573), .A2(n11572), .ZN(n11647) );
  AND2_X1 U11537 ( .A1(n11571), .A2(n11648), .ZN(n11646) );
  OR2_X1 U11538 ( .A1(n11573), .A2(n11572), .ZN(n11648) );
  OR2_X1 U11539 ( .A1(n8938), .A2(n8224), .ZN(n11572) );
  OR2_X1 U11540 ( .A1(n11649), .A2(n11650), .ZN(n11573) );
  AND2_X1 U11541 ( .A1(n11569), .A2(n11568), .ZN(n11650) );
  AND2_X1 U11542 ( .A1(n11566), .A2(n11651), .ZN(n11649) );
  OR2_X1 U11543 ( .A1(n11569), .A2(n11568), .ZN(n11651) );
  OR2_X1 U11544 ( .A1(n11652), .A2(n11653), .ZN(n11568) );
  AND2_X1 U11545 ( .A1(n11565), .A2(n11564), .ZN(n11653) );
  AND2_X1 U11546 ( .A1(n11562), .A2(n11654), .ZN(n11652) );
  OR2_X1 U11547 ( .A1(n11565), .A2(n11564), .ZN(n11654) );
  OR2_X1 U11548 ( .A1(n11655), .A2(n11656), .ZN(n11564) );
  AND2_X1 U11549 ( .A1(n11561), .A2(n11560), .ZN(n11656) );
  AND2_X1 U11550 ( .A1(n11558), .A2(n11657), .ZN(n11655) );
  OR2_X1 U11551 ( .A1(n11561), .A2(n11560), .ZN(n11657) );
  OR2_X1 U11552 ( .A1(n11658), .A2(n11659), .ZN(n11560) );
  AND2_X1 U11553 ( .A1(n11557), .A2(n11556), .ZN(n11659) );
  AND2_X1 U11554 ( .A1(n11555), .A2(n11660), .ZN(n11658) );
  OR2_X1 U11555 ( .A1(n11557), .A2(n11556), .ZN(n11660) );
  OR2_X1 U11556 ( .A1(n8954), .A2(n8224), .ZN(n11556) );
  OR2_X1 U11557 ( .A1(n11661), .A2(n11662), .ZN(n11557) );
  AND2_X1 U11558 ( .A1(n11553), .A2(n11552), .ZN(n11662) );
  AND2_X1 U11559 ( .A1(n11550), .A2(n11663), .ZN(n11661) );
  OR2_X1 U11560 ( .A1(n11553), .A2(n11552), .ZN(n11663) );
  OR2_X1 U11561 ( .A1(n11664), .A2(n11665), .ZN(n11552) );
  AND2_X1 U11562 ( .A1(n11549), .A2(n11548), .ZN(n11665) );
  AND2_X1 U11563 ( .A1(n11546), .A2(n11666), .ZN(n11664) );
  OR2_X1 U11564 ( .A1(n11549), .A2(n11548), .ZN(n11666) );
  OR2_X1 U11565 ( .A1(n11667), .A2(n11668), .ZN(n11548) );
  AND2_X1 U11566 ( .A1(n11545), .A2(n11544), .ZN(n11668) );
  AND2_X1 U11567 ( .A1(n11542), .A2(n11669), .ZN(n11667) );
  OR2_X1 U11568 ( .A1(n11545), .A2(n11544), .ZN(n11669) );
  OR2_X1 U11569 ( .A1(n11670), .A2(n11671), .ZN(n11544) );
  AND2_X1 U11570 ( .A1(n11541), .A2(n11540), .ZN(n11671) );
  AND2_X1 U11571 ( .A1(n11538), .A2(n11672), .ZN(n11670) );
  OR2_X1 U11572 ( .A1(n11541), .A2(n11540), .ZN(n11672) );
  OR2_X1 U11573 ( .A1(n11673), .A2(n11674), .ZN(n11540) );
  AND2_X1 U11574 ( .A1(n11537), .A2(n11536), .ZN(n11674) );
  AND2_X1 U11575 ( .A1(n11534), .A2(n11675), .ZN(n11673) );
  OR2_X1 U11576 ( .A1(n11537), .A2(n11536), .ZN(n11675) );
  OR2_X1 U11577 ( .A1(n11676), .A2(n11677), .ZN(n11536) );
  AND2_X1 U11578 ( .A1(n11533), .A2(n11532), .ZN(n11677) );
  AND2_X1 U11579 ( .A1(n11530), .A2(n11678), .ZN(n11676) );
  OR2_X1 U11580 ( .A1(n11533), .A2(n11532), .ZN(n11678) );
  OR2_X1 U11581 ( .A1(n11679), .A2(n11680), .ZN(n11532) );
  AND2_X1 U11582 ( .A1(n11529), .A2(n11528), .ZN(n11680) );
  AND2_X1 U11583 ( .A1(n11526), .A2(n11681), .ZN(n11679) );
  OR2_X1 U11584 ( .A1(n11529), .A2(n11528), .ZN(n11681) );
  OR2_X1 U11585 ( .A1(n11682), .A2(n11683), .ZN(n11528) );
  AND2_X1 U11586 ( .A1(n11525), .A2(n11524), .ZN(n11683) );
  AND2_X1 U11587 ( .A1(n11522), .A2(n11684), .ZN(n11682) );
  OR2_X1 U11588 ( .A1(n11525), .A2(n11524), .ZN(n11684) );
  OR2_X1 U11589 ( .A1(n11685), .A2(n11686), .ZN(n11524) );
  AND2_X1 U11590 ( .A1(n8991), .A2(n11521), .ZN(n11686) );
  AND2_X1 U11591 ( .A1(n11519), .A2(n11687), .ZN(n11685) );
  OR2_X1 U11592 ( .A1(n8991), .A2(n11521), .ZN(n11687) );
  OR2_X1 U11593 ( .A1(n11688), .A2(n11689), .ZN(n11521) );
  AND2_X1 U11594 ( .A1(n11518), .A2(n11517), .ZN(n11689) );
  AND2_X1 U11595 ( .A1(n11515), .A2(n11690), .ZN(n11688) );
  OR2_X1 U11596 ( .A1(n11518), .A2(n11517), .ZN(n11690) );
  OR2_X1 U11597 ( .A1(n11691), .A2(n11692), .ZN(n11517) );
  AND2_X1 U11598 ( .A1(n11514), .A2(n11513), .ZN(n11692) );
  AND2_X1 U11599 ( .A1(n11511), .A2(n11693), .ZN(n11691) );
  OR2_X1 U11600 ( .A1(n11514), .A2(n11513), .ZN(n11693) );
  OR2_X1 U11601 ( .A1(n11694), .A2(n11695), .ZN(n11513) );
  AND2_X1 U11602 ( .A1(n11510), .A2(n11509), .ZN(n11695) );
  AND2_X1 U11603 ( .A1(n11507), .A2(n11696), .ZN(n11694) );
  OR2_X1 U11604 ( .A1(n11510), .A2(n11509), .ZN(n11696) );
  OR2_X1 U11605 ( .A1(n11697), .A2(n11698), .ZN(n11509) );
  AND2_X1 U11606 ( .A1(n11506), .A2(n11505), .ZN(n11698) );
  AND2_X1 U11607 ( .A1(n11503), .A2(n11699), .ZN(n11697) );
  OR2_X1 U11608 ( .A1(n11506), .A2(n11505), .ZN(n11699) );
  OR2_X1 U11609 ( .A1(n11700), .A2(n11701), .ZN(n11505) );
  AND2_X1 U11610 ( .A1(n11502), .A2(n11501), .ZN(n11701) );
  AND2_X1 U11611 ( .A1(n11499), .A2(n11702), .ZN(n11700) );
  OR2_X1 U11612 ( .A1(n11502), .A2(n11501), .ZN(n11702) );
  OR2_X1 U11613 ( .A1(n11703), .A2(n11704), .ZN(n11501) );
  AND2_X1 U11614 ( .A1(n11496), .A2(n11497), .ZN(n11704) );
  AND2_X1 U11615 ( .A1(n11705), .A2(n11706), .ZN(n11703) );
  OR2_X1 U11616 ( .A1(n11496), .A2(n11497), .ZN(n11706) );
  OR2_X1 U11617 ( .A1(n9984), .A2(n11707), .ZN(n11497) );
  OR2_X1 U11618 ( .A1(n8224), .A2(n8252), .ZN(n11707) );
  OR2_X1 U11619 ( .A1(n9014), .A2(n8224), .ZN(n11496) );
  INV_X1 U11620 ( .A(n11498), .ZN(n11705) );
  OR2_X1 U11621 ( .A1(n11708), .A2(n11709), .ZN(n11498) );
  AND2_X1 U11622 ( .A1(b_22_), .A2(n11710), .ZN(n11709) );
  OR2_X1 U11623 ( .A1(n11711), .A2(n9989), .ZN(n11710) );
  AND2_X1 U11624 ( .A1(a_30_), .A2(n8280), .ZN(n11711) );
  AND2_X1 U11625 ( .A1(b_21_), .A2(n11712), .ZN(n11708) );
  OR2_X1 U11626 ( .A1(n11713), .A2(n8021), .ZN(n11712) );
  AND2_X1 U11627 ( .A1(a_31_), .A2(n8252), .ZN(n11713) );
  OR2_X1 U11628 ( .A1(n9010), .A2(n8224), .ZN(n11502) );
  XOR2_X1 U11629 ( .A(n11714), .B(n11715), .Z(n11499) );
  XNOR2_X1 U11630 ( .A(n11716), .B(n11717), .ZN(n11714) );
  OR2_X1 U11631 ( .A1(n9006), .A2(n8224), .ZN(n11506) );
  XOR2_X1 U11632 ( .A(n11718), .B(n11719), .Z(n11503) );
  XOR2_X1 U11633 ( .A(n11720), .B(n11721), .Z(n11719) );
  OR2_X1 U11634 ( .A1(n9002), .A2(n8224), .ZN(n11510) );
  XOR2_X1 U11635 ( .A(n11722), .B(n11723), .Z(n11507) );
  XOR2_X1 U11636 ( .A(n11724), .B(n11725), .Z(n11723) );
  OR2_X1 U11637 ( .A1(n8998), .A2(n8224), .ZN(n11514) );
  XOR2_X1 U11638 ( .A(n11726), .B(n11727), .Z(n11511) );
  XOR2_X1 U11639 ( .A(n11728), .B(n11729), .Z(n11727) );
  OR2_X1 U11640 ( .A1(n8994), .A2(n8224), .ZN(n11518) );
  XOR2_X1 U11641 ( .A(n11730), .B(n11731), .Z(n11515) );
  XOR2_X1 U11642 ( .A(n11732), .B(n11733), .Z(n11731) );
  OR2_X1 U11643 ( .A1(n8990), .A2(n8224), .ZN(n8991) );
  XOR2_X1 U11644 ( .A(n11734), .B(n11735), .Z(n11519) );
  XOR2_X1 U11645 ( .A(n11736), .B(n11737), .Z(n11735) );
  OR2_X1 U11646 ( .A1(n8986), .A2(n8224), .ZN(n11525) );
  XOR2_X1 U11647 ( .A(n11738), .B(n11739), .Z(n11522) );
  XOR2_X1 U11648 ( .A(n11740), .B(n11741), .Z(n11739) );
  OR2_X1 U11649 ( .A1(n8982), .A2(n8224), .ZN(n11529) );
  XOR2_X1 U11650 ( .A(n11742), .B(n11743), .Z(n11526) );
  XOR2_X1 U11651 ( .A(n11744), .B(n8987), .Z(n11743) );
  OR2_X1 U11652 ( .A1(n8978), .A2(n8224), .ZN(n11533) );
  XOR2_X1 U11653 ( .A(n11745), .B(n11746), .Z(n11530) );
  XOR2_X1 U11654 ( .A(n11747), .B(n11748), .Z(n11746) );
  OR2_X1 U11655 ( .A1(n8974), .A2(n8224), .ZN(n11537) );
  XOR2_X1 U11656 ( .A(n11749), .B(n11750), .Z(n11534) );
  XOR2_X1 U11657 ( .A(n11751), .B(n11752), .Z(n11750) );
  OR2_X1 U11658 ( .A1(n8970), .A2(n8224), .ZN(n11541) );
  XOR2_X1 U11659 ( .A(n11753), .B(n11754), .Z(n11538) );
  XOR2_X1 U11660 ( .A(n11755), .B(n11756), .Z(n11754) );
  OR2_X1 U11661 ( .A1(n8966), .A2(n8224), .ZN(n11545) );
  XOR2_X1 U11662 ( .A(n11757), .B(n11758), .Z(n11542) );
  XOR2_X1 U11663 ( .A(n11759), .B(n11760), .Z(n11758) );
  OR2_X1 U11664 ( .A1(n8962), .A2(n8224), .ZN(n11549) );
  XOR2_X1 U11665 ( .A(n11761), .B(n11762), .Z(n11546) );
  XOR2_X1 U11666 ( .A(n11763), .B(n11764), .Z(n11762) );
  OR2_X1 U11667 ( .A1(n8958), .A2(n8224), .ZN(n11553) );
  XOR2_X1 U11668 ( .A(n11765), .B(n11766), .Z(n11550) );
  XOR2_X1 U11669 ( .A(n11767), .B(n11768), .Z(n11766) );
  XOR2_X1 U11670 ( .A(n11769), .B(n11770), .Z(n11555) );
  XOR2_X1 U11671 ( .A(n11771), .B(n11772), .Z(n11770) );
  OR2_X1 U11672 ( .A1(n8950), .A2(n8224), .ZN(n11561) );
  XOR2_X1 U11673 ( .A(n11773), .B(n11774), .Z(n11558) );
  XOR2_X1 U11674 ( .A(n11775), .B(n11776), .Z(n11774) );
  OR2_X1 U11675 ( .A1(n8946), .A2(n8224), .ZN(n11565) );
  XOR2_X1 U11676 ( .A(n11777), .B(n11778), .Z(n11562) );
  XOR2_X1 U11677 ( .A(n11779), .B(n11780), .Z(n11778) );
  OR2_X1 U11678 ( .A1(n8942), .A2(n8224), .ZN(n11569) );
  XOR2_X1 U11679 ( .A(n11781), .B(n11782), .Z(n11566) );
  XOR2_X1 U11680 ( .A(n11783), .B(n11784), .Z(n11782) );
  XOR2_X1 U11681 ( .A(n11785), .B(n11786), .Z(n11571) );
  XOR2_X1 U11682 ( .A(n11787), .B(n11788), .Z(n11786) );
  OR2_X1 U11683 ( .A1(n8934), .A2(n8224), .ZN(n11577) );
  XOR2_X1 U11684 ( .A(n11789), .B(n11790), .Z(n11574) );
  XOR2_X1 U11685 ( .A(n11791), .B(n11792), .Z(n11790) );
  OR2_X1 U11686 ( .A1(n8930), .A2(n8224), .ZN(n11581) );
  XOR2_X1 U11687 ( .A(n11793), .B(n11794), .Z(n11578) );
  XOR2_X1 U11688 ( .A(n11795), .B(n11796), .Z(n11794) );
  OR2_X1 U11689 ( .A1(n8926), .A2(n8224), .ZN(n11585) );
  XOR2_X1 U11690 ( .A(n11797), .B(n11798), .Z(n11582) );
  XOR2_X1 U11691 ( .A(n11799), .B(n11800), .Z(n11798) );
  XOR2_X1 U11692 ( .A(n11801), .B(n11802), .Z(n11587) );
  XOR2_X1 U11693 ( .A(n11803), .B(n11804), .Z(n11802) );
  OR2_X1 U11694 ( .A1(n8918), .A2(n8224), .ZN(n11593) );
  XOR2_X1 U11695 ( .A(n11805), .B(n11806), .Z(n11590) );
  XOR2_X1 U11696 ( .A(n11807), .B(n11808), .Z(n11806) );
  OR2_X1 U11697 ( .A1(n8914), .A2(n8224), .ZN(n11597) );
  XOR2_X1 U11698 ( .A(n11809), .B(n11810), .Z(n11594) );
  XOR2_X1 U11699 ( .A(n11811), .B(n11812), .Z(n11810) );
  OR2_X1 U11700 ( .A1(n8910), .A2(n8224), .ZN(n11601) );
  XOR2_X1 U11701 ( .A(n11813), .B(n11814), .Z(n11598) );
  XOR2_X1 U11702 ( .A(n11815), .B(n11816), .Z(n11814) );
  OR2_X1 U11703 ( .A1(n8906), .A2(n8224), .ZN(n11605) );
  XOR2_X1 U11704 ( .A(n11817), .B(n11818), .Z(n11602) );
  XOR2_X1 U11705 ( .A(n11819), .B(n11820), .Z(n11818) );
  OR2_X1 U11706 ( .A1(n8902), .A2(n8224), .ZN(n11609) );
  XOR2_X1 U11707 ( .A(n11821), .B(n11822), .Z(n11606) );
  XOR2_X1 U11708 ( .A(n11823), .B(n11824), .Z(n11822) );
  OR2_X1 U11709 ( .A1(n11610), .A2(n11613), .ZN(n11618) );
  OR2_X1 U11710 ( .A1(n9297), .A2(n8224), .ZN(n11613) );
  XOR2_X1 U11711 ( .A(n11825), .B(n11826), .Z(n11610) );
  XOR2_X1 U11712 ( .A(n11827), .B(n11828), .Z(n11826) );
  XOR2_X1 U11713 ( .A(n11829), .B(n11830), .Z(n11394) );
  XOR2_X1 U11714 ( .A(n11831), .B(n11832), .Z(n11830) );
  OR2_X1 U11715 ( .A1(n9815), .A2(n9814), .ZN(n9104) );
  AND2_X1 U11716 ( .A1(n11833), .A2(n9796), .ZN(n9814) );
  OR2_X1 U11717 ( .A1(n11834), .A2(n11835), .ZN(n9796) );
  INV_X1 U11718 ( .A(n11836), .ZN(n11833) );
  AND2_X1 U11719 ( .A1(n11834), .A2(n11835), .ZN(n11836) );
  OR2_X1 U11720 ( .A1(n11837), .A2(n11838), .ZN(n11835) );
  AND2_X1 U11721 ( .A1(n11839), .A2(n11840), .ZN(n11838) );
  AND2_X1 U11722 ( .A1(n11841), .A2(n11842), .ZN(n11837) );
  OR2_X1 U11723 ( .A1(n11839), .A2(n11840), .ZN(n11841) );
  XOR2_X1 U11724 ( .A(n9805), .B(n11843), .Z(n11834) );
  XOR2_X1 U11725 ( .A(n9808), .B(n9806), .Z(n11843) );
  OR2_X1 U11726 ( .A1(n9297), .A2(n8308), .ZN(n9806) );
  OR2_X1 U11727 ( .A1(n11844), .A2(n11845), .ZN(n9808) );
  AND2_X1 U11728 ( .A1(n11846), .A2(n11847), .ZN(n11845) );
  AND2_X1 U11729 ( .A1(n11848), .A2(n11849), .ZN(n11844) );
  OR2_X1 U11730 ( .A1(n11846), .A2(n11847), .ZN(n11848) );
  XOR2_X1 U11731 ( .A(n11850), .B(n11851), .Z(n9805) );
  XOR2_X1 U11732 ( .A(n11852), .B(n11853), .Z(n11851) );
  AND2_X1 U11733 ( .A1(n11614), .A2(n11854), .ZN(n9815) );
  INV_X1 U11734 ( .A(n11615), .ZN(n11854) );
  OR2_X1 U11735 ( .A1(n11855), .A2(n11856), .ZN(n11615) );
  AND2_X1 U11736 ( .A1(n11829), .A2(n11832), .ZN(n11856) );
  AND2_X1 U11737 ( .A1(n11857), .A2(n11831), .ZN(n11855) );
  OR2_X1 U11738 ( .A1(n11858), .A2(n11859), .ZN(n11831) );
  AND2_X1 U11739 ( .A1(n11825), .A2(n11828), .ZN(n11859) );
  AND2_X1 U11740 ( .A1(n11860), .A2(n11827), .ZN(n11858) );
  OR2_X1 U11741 ( .A1(n11861), .A2(n11862), .ZN(n11827) );
  AND2_X1 U11742 ( .A1(n11821), .A2(n11824), .ZN(n11862) );
  AND2_X1 U11743 ( .A1(n11863), .A2(n11823), .ZN(n11861) );
  OR2_X1 U11744 ( .A1(n11864), .A2(n11865), .ZN(n11823) );
  AND2_X1 U11745 ( .A1(n11820), .A2(n11819), .ZN(n11865) );
  AND2_X1 U11746 ( .A1(n11817), .A2(n11866), .ZN(n11864) );
  OR2_X1 U11747 ( .A1(n11819), .A2(n11820), .ZN(n11866) );
  OR2_X1 U11748 ( .A1(n8910), .A2(n8252), .ZN(n11820) );
  OR2_X1 U11749 ( .A1(n11867), .A2(n11868), .ZN(n11819) );
  AND2_X1 U11750 ( .A1(n11816), .A2(n11815), .ZN(n11868) );
  AND2_X1 U11751 ( .A1(n11813), .A2(n11869), .ZN(n11867) );
  OR2_X1 U11752 ( .A1(n11815), .A2(n11816), .ZN(n11869) );
  OR2_X1 U11753 ( .A1(n8914), .A2(n8252), .ZN(n11816) );
  OR2_X1 U11754 ( .A1(n11870), .A2(n11871), .ZN(n11815) );
  AND2_X1 U11755 ( .A1(n11812), .A2(n11811), .ZN(n11871) );
  AND2_X1 U11756 ( .A1(n11809), .A2(n11872), .ZN(n11870) );
  OR2_X1 U11757 ( .A1(n11811), .A2(n11812), .ZN(n11872) );
  OR2_X1 U11758 ( .A1(n8918), .A2(n8252), .ZN(n11812) );
  OR2_X1 U11759 ( .A1(n11873), .A2(n11874), .ZN(n11811) );
  AND2_X1 U11760 ( .A1(n11808), .A2(n11807), .ZN(n11874) );
  AND2_X1 U11761 ( .A1(n11805), .A2(n11875), .ZN(n11873) );
  OR2_X1 U11762 ( .A1(n11807), .A2(n11808), .ZN(n11875) );
  OR2_X1 U11763 ( .A1(n8922), .A2(n8252), .ZN(n11808) );
  OR2_X1 U11764 ( .A1(n11876), .A2(n11877), .ZN(n11807) );
  AND2_X1 U11765 ( .A1(n11804), .A2(n11803), .ZN(n11877) );
  AND2_X1 U11766 ( .A1(n11801), .A2(n11878), .ZN(n11876) );
  OR2_X1 U11767 ( .A1(n11803), .A2(n11804), .ZN(n11878) );
  OR2_X1 U11768 ( .A1(n8926), .A2(n8252), .ZN(n11804) );
  OR2_X1 U11769 ( .A1(n11879), .A2(n11880), .ZN(n11803) );
  AND2_X1 U11770 ( .A1(n11800), .A2(n11799), .ZN(n11880) );
  AND2_X1 U11771 ( .A1(n11797), .A2(n11881), .ZN(n11879) );
  OR2_X1 U11772 ( .A1(n11799), .A2(n11800), .ZN(n11881) );
  OR2_X1 U11773 ( .A1(n8930), .A2(n8252), .ZN(n11800) );
  OR2_X1 U11774 ( .A1(n11882), .A2(n11883), .ZN(n11799) );
  AND2_X1 U11775 ( .A1(n11796), .A2(n11795), .ZN(n11883) );
  AND2_X1 U11776 ( .A1(n11793), .A2(n11884), .ZN(n11882) );
  OR2_X1 U11777 ( .A1(n11795), .A2(n11796), .ZN(n11884) );
  OR2_X1 U11778 ( .A1(n8934), .A2(n8252), .ZN(n11796) );
  OR2_X1 U11779 ( .A1(n11885), .A2(n11886), .ZN(n11795) );
  AND2_X1 U11780 ( .A1(n11792), .A2(n11791), .ZN(n11886) );
  AND2_X1 U11781 ( .A1(n11789), .A2(n11887), .ZN(n11885) );
  OR2_X1 U11782 ( .A1(n11791), .A2(n11792), .ZN(n11887) );
  OR2_X1 U11783 ( .A1(n8938), .A2(n8252), .ZN(n11792) );
  OR2_X1 U11784 ( .A1(n11888), .A2(n11889), .ZN(n11791) );
  AND2_X1 U11785 ( .A1(n11788), .A2(n11787), .ZN(n11889) );
  AND2_X1 U11786 ( .A1(n11785), .A2(n11890), .ZN(n11888) );
  OR2_X1 U11787 ( .A1(n11787), .A2(n11788), .ZN(n11890) );
  OR2_X1 U11788 ( .A1(n8942), .A2(n8252), .ZN(n11788) );
  OR2_X1 U11789 ( .A1(n11891), .A2(n11892), .ZN(n11787) );
  AND2_X1 U11790 ( .A1(n11784), .A2(n11783), .ZN(n11892) );
  AND2_X1 U11791 ( .A1(n11781), .A2(n11893), .ZN(n11891) );
  OR2_X1 U11792 ( .A1(n11783), .A2(n11784), .ZN(n11893) );
  OR2_X1 U11793 ( .A1(n8946), .A2(n8252), .ZN(n11784) );
  OR2_X1 U11794 ( .A1(n11894), .A2(n11895), .ZN(n11783) );
  AND2_X1 U11795 ( .A1(n11780), .A2(n11779), .ZN(n11895) );
  AND2_X1 U11796 ( .A1(n11777), .A2(n11896), .ZN(n11894) );
  OR2_X1 U11797 ( .A1(n11779), .A2(n11780), .ZN(n11896) );
  OR2_X1 U11798 ( .A1(n8950), .A2(n8252), .ZN(n11780) );
  OR2_X1 U11799 ( .A1(n11897), .A2(n11898), .ZN(n11779) );
  AND2_X1 U11800 ( .A1(n11776), .A2(n11775), .ZN(n11898) );
  AND2_X1 U11801 ( .A1(n11773), .A2(n11899), .ZN(n11897) );
  OR2_X1 U11802 ( .A1(n11775), .A2(n11776), .ZN(n11899) );
  OR2_X1 U11803 ( .A1(n8954), .A2(n8252), .ZN(n11776) );
  OR2_X1 U11804 ( .A1(n11900), .A2(n11901), .ZN(n11775) );
  AND2_X1 U11805 ( .A1(n11772), .A2(n11771), .ZN(n11901) );
  AND2_X1 U11806 ( .A1(n11769), .A2(n11902), .ZN(n11900) );
  OR2_X1 U11807 ( .A1(n11771), .A2(n11772), .ZN(n11902) );
  OR2_X1 U11808 ( .A1(n8958), .A2(n8252), .ZN(n11772) );
  OR2_X1 U11809 ( .A1(n11903), .A2(n11904), .ZN(n11771) );
  AND2_X1 U11810 ( .A1(n11768), .A2(n11767), .ZN(n11904) );
  AND2_X1 U11811 ( .A1(n11765), .A2(n11905), .ZN(n11903) );
  OR2_X1 U11812 ( .A1(n11767), .A2(n11768), .ZN(n11905) );
  OR2_X1 U11813 ( .A1(n8962), .A2(n8252), .ZN(n11768) );
  OR2_X1 U11814 ( .A1(n11906), .A2(n11907), .ZN(n11767) );
  AND2_X1 U11815 ( .A1(n11764), .A2(n11763), .ZN(n11907) );
  AND2_X1 U11816 ( .A1(n11761), .A2(n11908), .ZN(n11906) );
  OR2_X1 U11817 ( .A1(n11763), .A2(n11764), .ZN(n11908) );
  OR2_X1 U11818 ( .A1(n8966), .A2(n8252), .ZN(n11764) );
  OR2_X1 U11819 ( .A1(n11909), .A2(n11910), .ZN(n11763) );
  AND2_X1 U11820 ( .A1(n11760), .A2(n11759), .ZN(n11910) );
  AND2_X1 U11821 ( .A1(n11757), .A2(n11911), .ZN(n11909) );
  OR2_X1 U11822 ( .A1(n11759), .A2(n11760), .ZN(n11911) );
  OR2_X1 U11823 ( .A1(n8970), .A2(n8252), .ZN(n11760) );
  OR2_X1 U11824 ( .A1(n11912), .A2(n11913), .ZN(n11759) );
  AND2_X1 U11825 ( .A1(n11756), .A2(n11755), .ZN(n11913) );
  AND2_X1 U11826 ( .A1(n11753), .A2(n11914), .ZN(n11912) );
  OR2_X1 U11827 ( .A1(n11755), .A2(n11756), .ZN(n11914) );
  OR2_X1 U11828 ( .A1(n8974), .A2(n8252), .ZN(n11756) );
  OR2_X1 U11829 ( .A1(n11915), .A2(n11916), .ZN(n11755) );
  AND2_X1 U11830 ( .A1(n11752), .A2(n11751), .ZN(n11916) );
  AND2_X1 U11831 ( .A1(n11749), .A2(n11917), .ZN(n11915) );
  OR2_X1 U11832 ( .A1(n11751), .A2(n11752), .ZN(n11917) );
  OR2_X1 U11833 ( .A1(n8978), .A2(n8252), .ZN(n11752) );
  OR2_X1 U11834 ( .A1(n11918), .A2(n11919), .ZN(n11751) );
  AND2_X1 U11835 ( .A1(n11748), .A2(n11747), .ZN(n11919) );
  AND2_X1 U11836 ( .A1(n11745), .A2(n11920), .ZN(n11918) );
  OR2_X1 U11837 ( .A1(n11747), .A2(n11748), .ZN(n11920) );
  OR2_X1 U11838 ( .A1(n8982), .A2(n8252), .ZN(n11748) );
  OR2_X1 U11839 ( .A1(n11921), .A2(n11922), .ZN(n11747) );
  AND2_X1 U11840 ( .A1(n8987), .A2(n11744), .ZN(n11922) );
  AND2_X1 U11841 ( .A1(n11742), .A2(n11923), .ZN(n11921) );
  OR2_X1 U11842 ( .A1(n11744), .A2(n8987), .ZN(n11923) );
  OR2_X1 U11843 ( .A1(n8986), .A2(n8252), .ZN(n8987) );
  OR2_X1 U11844 ( .A1(n11924), .A2(n11925), .ZN(n11744) );
  AND2_X1 U11845 ( .A1(n11741), .A2(n11740), .ZN(n11925) );
  AND2_X1 U11846 ( .A1(n11738), .A2(n11926), .ZN(n11924) );
  OR2_X1 U11847 ( .A1(n11740), .A2(n11741), .ZN(n11926) );
  OR2_X1 U11848 ( .A1(n8990), .A2(n8252), .ZN(n11741) );
  OR2_X1 U11849 ( .A1(n11927), .A2(n11928), .ZN(n11740) );
  AND2_X1 U11850 ( .A1(n11737), .A2(n11736), .ZN(n11928) );
  AND2_X1 U11851 ( .A1(n11734), .A2(n11929), .ZN(n11927) );
  OR2_X1 U11852 ( .A1(n11736), .A2(n11737), .ZN(n11929) );
  OR2_X1 U11853 ( .A1(n8994), .A2(n8252), .ZN(n11737) );
  OR2_X1 U11854 ( .A1(n11930), .A2(n11931), .ZN(n11736) );
  AND2_X1 U11855 ( .A1(n11733), .A2(n11732), .ZN(n11931) );
  AND2_X1 U11856 ( .A1(n11730), .A2(n11932), .ZN(n11930) );
  OR2_X1 U11857 ( .A1(n11732), .A2(n11733), .ZN(n11932) );
  OR2_X1 U11858 ( .A1(n8998), .A2(n8252), .ZN(n11733) );
  OR2_X1 U11859 ( .A1(n11933), .A2(n11934), .ZN(n11732) );
  AND2_X1 U11860 ( .A1(n11729), .A2(n11728), .ZN(n11934) );
  AND2_X1 U11861 ( .A1(n11726), .A2(n11935), .ZN(n11933) );
  OR2_X1 U11862 ( .A1(n11728), .A2(n11729), .ZN(n11935) );
  OR2_X1 U11863 ( .A1(n9002), .A2(n8252), .ZN(n11729) );
  OR2_X1 U11864 ( .A1(n11936), .A2(n11937), .ZN(n11728) );
  AND2_X1 U11865 ( .A1(n11725), .A2(n11724), .ZN(n11937) );
  AND2_X1 U11866 ( .A1(n11722), .A2(n11938), .ZN(n11936) );
  OR2_X1 U11867 ( .A1(n11724), .A2(n11725), .ZN(n11938) );
  OR2_X1 U11868 ( .A1(n9006), .A2(n8252), .ZN(n11725) );
  OR2_X1 U11869 ( .A1(n11939), .A2(n11940), .ZN(n11724) );
  AND2_X1 U11870 ( .A1(n11721), .A2(n11720), .ZN(n11940) );
  AND2_X1 U11871 ( .A1(n11718), .A2(n11941), .ZN(n11939) );
  OR2_X1 U11872 ( .A1(n11720), .A2(n11721), .ZN(n11941) );
  OR2_X1 U11873 ( .A1(n9010), .A2(n8252), .ZN(n11721) );
  OR2_X1 U11874 ( .A1(n11942), .A2(n11943), .ZN(n11720) );
  AND2_X1 U11875 ( .A1(n11715), .A2(n11716), .ZN(n11943) );
  AND2_X1 U11876 ( .A1(n11944), .A2(n11945), .ZN(n11942) );
  OR2_X1 U11877 ( .A1(n11716), .A2(n11715), .ZN(n11945) );
  OR2_X1 U11878 ( .A1(n9014), .A2(n8252), .ZN(n11715) );
  OR2_X1 U11879 ( .A1(n9984), .A2(n11946), .ZN(n11716) );
  OR2_X1 U11880 ( .A1(n8252), .A2(n8280), .ZN(n11946) );
  INV_X1 U11881 ( .A(n11717), .ZN(n11944) );
  OR2_X1 U11882 ( .A1(n11947), .A2(n11948), .ZN(n11717) );
  AND2_X1 U11883 ( .A1(b_21_), .A2(n11949), .ZN(n11948) );
  OR2_X1 U11884 ( .A1(n11950), .A2(n9989), .ZN(n11949) );
  AND2_X1 U11885 ( .A1(a_30_), .A2(n8308), .ZN(n11950) );
  AND2_X1 U11886 ( .A1(b_20_), .A2(n11951), .ZN(n11947) );
  OR2_X1 U11887 ( .A1(n11952), .A2(n8021), .ZN(n11951) );
  AND2_X1 U11888 ( .A1(a_31_), .A2(n8280), .ZN(n11952) );
  XOR2_X1 U11889 ( .A(n11953), .B(n11954), .Z(n11718) );
  XNOR2_X1 U11890 ( .A(n11955), .B(n11956), .ZN(n11953) );
  XOR2_X1 U11891 ( .A(n11957), .B(n11958), .Z(n11722) );
  XOR2_X1 U11892 ( .A(n11959), .B(n11960), .Z(n11958) );
  XOR2_X1 U11893 ( .A(n11961), .B(n11962), .Z(n11726) );
  XOR2_X1 U11894 ( .A(n11963), .B(n11964), .Z(n11962) );
  XOR2_X1 U11895 ( .A(n11965), .B(n11966), .Z(n11730) );
  XOR2_X1 U11896 ( .A(n11967), .B(n11968), .Z(n11966) );
  XOR2_X1 U11897 ( .A(n11969), .B(n11970), .Z(n11734) );
  XOR2_X1 U11898 ( .A(n11971), .B(n11972), .Z(n11970) );
  XOR2_X1 U11899 ( .A(n11973), .B(n11974), .Z(n11738) );
  XOR2_X1 U11900 ( .A(n11975), .B(n11976), .Z(n11974) );
  XOR2_X1 U11901 ( .A(n11977), .B(n11978), .Z(n11742) );
  XOR2_X1 U11902 ( .A(n11979), .B(n11980), .Z(n11978) );
  XOR2_X1 U11903 ( .A(n11981), .B(n11982), .Z(n11745) );
  XOR2_X1 U11904 ( .A(n11983), .B(n11984), .Z(n11982) );
  XOR2_X1 U11905 ( .A(n11985), .B(n11986), .Z(n11749) );
  XOR2_X1 U11906 ( .A(n11987), .B(n8983), .Z(n11986) );
  XOR2_X1 U11907 ( .A(n11988), .B(n11989), .Z(n11753) );
  XOR2_X1 U11908 ( .A(n11990), .B(n11991), .Z(n11989) );
  XOR2_X1 U11909 ( .A(n11992), .B(n11993), .Z(n11757) );
  XOR2_X1 U11910 ( .A(n11994), .B(n11995), .Z(n11993) );
  XOR2_X1 U11911 ( .A(n11996), .B(n11997), .Z(n11761) );
  XOR2_X1 U11912 ( .A(n11998), .B(n11999), .Z(n11997) );
  XOR2_X1 U11913 ( .A(n12000), .B(n12001), .Z(n11765) );
  XOR2_X1 U11914 ( .A(n12002), .B(n12003), .Z(n12001) );
  XOR2_X1 U11915 ( .A(n12004), .B(n12005), .Z(n11769) );
  XOR2_X1 U11916 ( .A(n12006), .B(n12007), .Z(n12005) );
  XOR2_X1 U11917 ( .A(n12008), .B(n12009), .Z(n11773) );
  XOR2_X1 U11918 ( .A(n12010), .B(n12011), .Z(n12009) );
  XOR2_X1 U11919 ( .A(n12012), .B(n12013), .Z(n11777) );
  XOR2_X1 U11920 ( .A(n12014), .B(n12015), .Z(n12013) );
  XOR2_X1 U11921 ( .A(n12016), .B(n12017), .Z(n11781) );
  XOR2_X1 U11922 ( .A(n12018), .B(n12019), .Z(n12017) );
  XOR2_X1 U11923 ( .A(n12020), .B(n12021), .Z(n11785) );
  XOR2_X1 U11924 ( .A(n12022), .B(n12023), .Z(n12021) );
  XOR2_X1 U11925 ( .A(n12024), .B(n12025), .Z(n11789) );
  XOR2_X1 U11926 ( .A(n12026), .B(n12027), .Z(n12025) );
  XOR2_X1 U11927 ( .A(n12028), .B(n12029), .Z(n11793) );
  XOR2_X1 U11928 ( .A(n12030), .B(n12031), .Z(n12029) );
  XOR2_X1 U11929 ( .A(n12032), .B(n12033), .Z(n11797) );
  XOR2_X1 U11930 ( .A(n12034), .B(n12035), .Z(n12033) );
  XOR2_X1 U11931 ( .A(n12036), .B(n12037), .Z(n11801) );
  XOR2_X1 U11932 ( .A(n12038), .B(n12039), .Z(n12037) );
  XOR2_X1 U11933 ( .A(n12040), .B(n12041), .Z(n11805) );
  XOR2_X1 U11934 ( .A(n12042), .B(n12043), .Z(n12041) );
  XOR2_X1 U11935 ( .A(n12044), .B(n12045), .Z(n11809) );
  XOR2_X1 U11936 ( .A(n12046), .B(n12047), .Z(n12045) );
  XOR2_X1 U11937 ( .A(n12048), .B(n12049), .Z(n11813) );
  XOR2_X1 U11938 ( .A(n12050), .B(n12051), .Z(n12049) );
  XOR2_X1 U11939 ( .A(n12052), .B(n12053), .Z(n11817) );
  XOR2_X1 U11940 ( .A(n12054), .B(n12055), .Z(n12053) );
  OR2_X1 U11941 ( .A1(n11821), .A2(n11824), .ZN(n11863) );
  OR2_X1 U11942 ( .A1(n8906), .A2(n8252), .ZN(n11824) );
  XOR2_X1 U11943 ( .A(n12056), .B(n12057), .Z(n11821) );
  XOR2_X1 U11944 ( .A(n12058), .B(n12059), .Z(n12057) );
  OR2_X1 U11945 ( .A1(n11825), .A2(n11828), .ZN(n11860) );
  OR2_X1 U11946 ( .A1(n8902), .A2(n8252), .ZN(n11828) );
  XOR2_X1 U11947 ( .A(n12060), .B(n12061), .Z(n11825) );
  XOR2_X1 U11948 ( .A(n12062), .B(n12063), .Z(n12061) );
  OR2_X1 U11949 ( .A1(n11829), .A2(n11832), .ZN(n11857) );
  OR2_X1 U11950 ( .A1(n9297), .A2(n8252), .ZN(n11832) );
  XOR2_X1 U11951 ( .A(n12064), .B(n12065), .Z(n11829) );
  XOR2_X1 U11952 ( .A(n12066), .B(n12067), .Z(n12065) );
  XNOR2_X1 U11953 ( .A(n11839), .B(n12068), .ZN(n11614) );
  XOR2_X1 U11954 ( .A(n11842), .B(n11840), .Z(n12068) );
  OR2_X1 U11955 ( .A1(n9297), .A2(n8280), .ZN(n11840) );
  OR2_X1 U11956 ( .A1(n12069), .A2(n12070), .ZN(n11842) );
  AND2_X1 U11957 ( .A1(n12064), .A2(n12067), .ZN(n12070) );
  AND2_X1 U11958 ( .A1(n12071), .A2(n12066), .ZN(n12069) );
  OR2_X1 U11959 ( .A1(n12072), .A2(n12073), .ZN(n12066) );
  AND2_X1 U11960 ( .A1(n12060), .A2(n12063), .ZN(n12073) );
  AND2_X1 U11961 ( .A1(n12074), .A2(n12062), .ZN(n12072) );
  OR2_X1 U11962 ( .A1(n12075), .A2(n12076), .ZN(n12062) );
  AND2_X1 U11963 ( .A1(n12056), .A2(n12059), .ZN(n12076) );
  AND2_X1 U11964 ( .A1(n12077), .A2(n12058), .ZN(n12075) );
  OR2_X1 U11965 ( .A1(n12078), .A2(n12079), .ZN(n12058) );
  AND2_X1 U11966 ( .A1(n12052), .A2(n12055), .ZN(n12079) );
  AND2_X1 U11967 ( .A1(n12080), .A2(n12054), .ZN(n12078) );
  OR2_X1 U11968 ( .A1(n12081), .A2(n12082), .ZN(n12054) );
  AND2_X1 U11969 ( .A1(n12051), .A2(n12050), .ZN(n12082) );
  AND2_X1 U11970 ( .A1(n12048), .A2(n12083), .ZN(n12081) );
  OR2_X1 U11971 ( .A1(n12051), .A2(n12050), .ZN(n12083) );
  OR2_X1 U11972 ( .A1(n12084), .A2(n12085), .ZN(n12050) );
  AND2_X1 U11973 ( .A1(n12047), .A2(n12046), .ZN(n12085) );
  AND2_X1 U11974 ( .A1(n12044), .A2(n12086), .ZN(n12084) );
  OR2_X1 U11975 ( .A1(n12047), .A2(n12046), .ZN(n12086) );
  OR2_X1 U11976 ( .A1(n12087), .A2(n12088), .ZN(n12046) );
  AND2_X1 U11977 ( .A1(n12043), .A2(n12042), .ZN(n12088) );
  AND2_X1 U11978 ( .A1(n12040), .A2(n12089), .ZN(n12087) );
  OR2_X1 U11979 ( .A1(n12043), .A2(n12042), .ZN(n12089) );
  OR2_X1 U11980 ( .A1(n12090), .A2(n12091), .ZN(n12042) );
  AND2_X1 U11981 ( .A1(n12039), .A2(n12038), .ZN(n12091) );
  AND2_X1 U11982 ( .A1(n12036), .A2(n12092), .ZN(n12090) );
  OR2_X1 U11983 ( .A1(n12039), .A2(n12038), .ZN(n12092) );
  OR2_X1 U11984 ( .A1(n12093), .A2(n12094), .ZN(n12038) );
  AND2_X1 U11985 ( .A1(n12035), .A2(n12034), .ZN(n12094) );
  AND2_X1 U11986 ( .A1(n12032), .A2(n12095), .ZN(n12093) );
  OR2_X1 U11987 ( .A1(n12035), .A2(n12034), .ZN(n12095) );
  OR2_X1 U11988 ( .A1(n12096), .A2(n12097), .ZN(n12034) );
  AND2_X1 U11989 ( .A1(n12031), .A2(n12030), .ZN(n12097) );
  AND2_X1 U11990 ( .A1(n12028), .A2(n12098), .ZN(n12096) );
  OR2_X1 U11991 ( .A1(n12031), .A2(n12030), .ZN(n12098) );
  OR2_X1 U11992 ( .A1(n12099), .A2(n12100), .ZN(n12030) );
  AND2_X1 U11993 ( .A1(n12027), .A2(n12026), .ZN(n12100) );
  AND2_X1 U11994 ( .A1(n12024), .A2(n12101), .ZN(n12099) );
  OR2_X1 U11995 ( .A1(n12027), .A2(n12026), .ZN(n12101) );
  OR2_X1 U11996 ( .A1(n12102), .A2(n12103), .ZN(n12026) );
  AND2_X1 U11997 ( .A1(n12023), .A2(n12022), .ZN(n12103) );
  AND2_X1 U11998 ( .A1(n12020), .A2(n12104), .ZN(n12102) );
  OR2_X1 U11999 ( .A1(n12023), .A2(n12022), .ZN(n12104) );
  OR2_X1 U12000 ( .A1(n12105), .A2(n12106), .ZN(n12022) );
  AND2_X1 U12001 ( .A1(n12019), .A2(n12018), .ZN(n12106) );
  AND2_X1 U12002 ( .A1(n12016), .A2(n12107), .ZN(n12105) );
  OR2_X1 U12003 ( .A1(n12019), .A2(n12018), .ZN(n12107) );
  OR2_X1 U12004 ( .A1(n12108), .A2(n12109), .ZN(n12018) );
  AND2_X1 U12005 ( .A1(n12015), .A2(n12014), .ZN(n12109) );
  AND2_X1 U12006 ( .A1(n12012), .A2(n12110), .ZN(n12108) );
  OR2_X1 U12007 ( .A1(n12015), .A2(n12014), .ZN(n12110) );
  OR2_X1 U12008 ( .A1(n12111), .A2(n12112), .ZN(n12014) );
  AND2_X1 U12009 ( .A1(n12011), .A2(n12010), .ZN(n12112) );
  AND2_X1 U12010 ( .A1(n12008), .A2(n12113), .ZN(n12111) );
  OR2_X1 U12011 ( .A1(n12011), .A2(n12010), .ZN(n12113) );
  OR2_X1 U12012 ( .A1(n12114), .A2(n12115), .ZN(n12010) );
  AND2_X1 U12013 ( .A1(n12007), .A2(n12006), .ZN(n12115) );
  AND2_X1 U12014 ( .A1(n12004), .A2(n12116), .ZN(n12114) );
  OR2_X1 U12015 ( .A1(n12007), .A2(n12006), .ZN(n12116) );
  OR2_X1 U12016 ( .A1(n12117), .A2(n12118), .ZN(n12006) );
  AND2_X1 U12017 ( .A1(n12003), .A2(n12002), .ZN(n12118) );
  AND2_X1 U12018 ( .A1(n12000), .A2(n12119), .ZN(n12117) );
  OR2_X1 U12019 ( .A1(n12003), .A2(n12002), .ZN(n12119) );
  OR2_X1 U12020 ( .A1(n12120), .A2(n12121), .ZN(n12002) );
  AND2_X1 U12021 ( .A1(n11999), .A2(n11998), .ZN(n12121) );
  AND2_X1 U12022 ( .A1(n11996), .A2(n12122), .ZN(n12120) );
  OR2_X1 U12023 ( .A1(n11999), .A2(n11998), .ZN(n12122) );
  OR2_X1 U12024 ( .A1(n12123), .A2(n12124), .ZN(n11998) );
  AND2_X1 U12025 ( .A1(n11995), .A2(n11994), .ZN(n12124) );
  AND2_X1 U12026 ( .A1(n11992), .A2(n12125), .ZN(n12123) );
  OR2_X1 U12027 ( .A1(n11995), .A2(n11994), .ZN(n12125) );
  OR2_X1 U12028 ( .A1(n12126), .A2(n12127), .ZN(n11994) );
  AND2_X1 U12029 ( .A1(n11991), .A2(n11990), .ZN(n12127) );
  AND2_X1 U12030 ( .A1(n11988), .A2(n12128), .ZN(n12126) );
  OR2_X1 U12031 ( .A1(n11991), .A2(n11990), .ZN(n12128) );
  OR2_X1 U12032 ( .A1(n12129), .A2(n12130), .ZN(n11990) );
  AND2_X1 U12033 ( .A1(n8983), .A2(n11987), .ZN(n12130) );
  AND2_X1 U12034 ( .A1(n11985), .A2(n12131), .ZN(n12129) );
  OR2_X1 U12035 ( .A1(n8983), .A2(n11987), .ZN(n12131) );
  OR2_X1 U12036 ( .A1(n12132), .A2(n12133), .ZN(n11987) );
  AND2_X1 U12037 ( .A1(n11984), .A2(n11983), .ZN(n12133) );
  AND2_X1 U12038 ( .A1(n11981), .A2(n12134), .ZN(n12132) );
  OR2_X1 U12039 ( .A1(n11984), .A2(n11983), .ZN(n12134) );
  OR2_X1 U12040 ( .A1(n12135), .A2(n12136), .ZN(n11983) );
  AND2_X1 U12041 ( .A1(n11980), .A2(n11979), .ZN(n12136) );
  AND2_X1 U12042 ( .A1(n11977), .A2(n12137), .ZN(n12135) );
  OR2_X1 U12043 ( .A1(n11980), .A2(n11979), .ZN(n12137) );
  OR2_X1 U12044 ( .A1(n12138), .A2(n12139), .ZN(n11979) );
  AND2_X1 U12045 ( .A1(n11976), .A2(n11975), .ZN(n12139) );
  AND2_X1 U12046 ( .A1(n11973), .A2(n12140), .ZN(n12138) );
  OR2_X1 U12047 ( .A1(n11976), .A2(n11975), .ZN(n12140) );
  OR2_X1 U12048 ( .A1(n12141), .A2(n12142), .ZN(n11975) );
  AND2_X1 U12049 ( .A1(n11972), .A2(n11971), .ZN(n12142) );
  AND2_X1 U12050 ( .A1(n11969), .A2(n12143), .ZN(n12141) );
  OR2_X1 U12051 ( .A1(n11972), .A2(n11971), .ZN(n12143) );
  OR2_X1 U12052 ( .A1(n12144), .A2(n12145), .ZN(n11971) );
  AND2_X1 U12053 ( .A1(n11968), .A2(n11967), .ZN(n12145) );
  AND2_X1 U12054 ( .A1(n11965), .A2(n12146), .ZN(n12144) );
  OR2_X1 U12055 ( .A1(n11968), .A2(n11967), .ZN(n12146) );
  OR2_X1 U12056 ( .A1(n12147), .A2(n12148), .ZN(n11967) );
  AND2_X1 U12057 ( .A1(n11964), .A2(n11963), .ZN(n12148) );
  AND2_X1 U12058 ( .A1(n11961), .A2(n12149), .ZN(n12147) );
  OR2_X1 U12059 ( .A1(n11964), .A2(n11963), .ZN(n12149) );
  OR2_X1 U12060 ( .A1(n12150), .A2(n12151), .ZN(n11963) );
  AND2_X1 U12061 ( .A1(n11960), .A2(n11959), .ZN(n12151) );
  AND2_X1 U12062 ( .A1(n11957), .A2(n12152), .ZN(n12150) );
  OR2_X1 U12063 ( .A1(n11960), .A2(n11959), .ZN(n12152) );
  OR2_X1 U12064 ( .A1(n12153), .A2(n12154), .ZN(n11959) );
  AND2_X1 U12065 ( .A1(n11954), .A2(n11955), .ZN(n12154) );
  AND2_X1 U12066 ( .A1(n12155), .A2(n12156), .ZN(n12153) );
  OR2_X1 U12067 ( .A1(n11954), .A2(n11955), .ZN(n12156) );
  OR2_X1 U12068 ( .A1(n9984), .A2(n12157), .ZN(n11955) );
  OR2_X1 U12069 ( .A1(n8280), .A2(n8308), .ZN(n12157) );
  OR2_X1 U12070 ( .A1(n9014), .A2(n8280), .ZN(n11954) );
  INV_X1 U12071 ( .A(n11956), .ZN(n12155) );
  OR2_X1 U12072 ( .A1(n12158), .A2(n12159), .ZN(n11956) );
  AND2_X1 U12073 ( .A1(b_20_), .A2(n12160), .ZN(n12159) );
  OR2_X1 U12074 ( .A1(n12161), .A2(n9989), .ZN(n12160) );
  AND2_X1 U12075 ( .A1(a_30_), .A2(n8336), .ZN(n12161) );
  AND2_X1 U12076 ( .A1(b_19_), .A2(n12162), .ZN(n12158) );
  OR2_X1 U12077 ( .A1(n12163), .A2(n8021), .ZN(n12162) );
  AND2_X1 U12078 ( .A1(a_31_), .A2(n8308), .ZN(n12163) );
  OR2_X1 U12079 ( .A1(n9010), .A2(n8280), .ZN(n11960) );
  XOR2_X1 U12080 ( .A(n12164), .B(n12165), .Z(n11957) );
  XNOR2_X1 U12081 ( .A(n12166), .B(n12167), .ZN(n12164) );
  OR2_X1 U12082 ( .A1(n9006), .A2(n8280), .ZN(n11964) );
  XOR2_X1 U12083 ( .A(n12168), .B(n12169), .Z(n11961) );
  XOR2_X1 U12084 ( .A(n12170), .B(n12171), .Z(n12169) );
  OR2_X1 U12085 ( .A1(n9002), .A2(n8280), .ZN(n11968) );
  XOR2_X1 U12086 ( .A(n12172), .B(n12173), .Z(n11965) );
  XOR2_X1 U12087 ( .A(n12174), .B(n12175), .Z(n12173) );
  OR2_X1 U12088 ( .A1(n8998), .A2(n8280), .ZN(n11972) );
  XOR2_X1 U12089 ( .A(n12176), .B(n12177), .Z(n11969) );
  XOR2_X1 U12090 ( .A(n12178), .B(n12179), .Z(n12177) );
  OR2_X1 U12091 ( .A1(n8994), .A2(n8280), .ZN(n11976) );
  XOR2_X1 U12092 ( .A(n12180), .B(n12181), .Z(n11973) );
  XOR2_X1 U12093 ( .A(n12182), .B(n12183), .Z(n12181) );
  OR2_X1 U12094 ( .A1(n8990), .A2(n8280), .ZN(n11980) );
  XOR2_X1 U12095 ( .A(n12184), .B(n12185), .Z(n11977) );
  XOR2_X1 U12096 ( .A(n12186), .B(n12187), .Z(n12185) );
  OR2_X1 U12097 ( .A1(n8986), .A2(n8280), .ZN(n11984) );
  XOR2_X1 U12098 ( .A(n12188), .B(n12189), .Z(n11981) );
  XOR2_X1 U12099 ( .A(n12190), .B(n12191), .Z(n12189) );
  OR2_X1 U12100 ( .A1(n8982), .A2(n8280), .ZN(n8983) );
  XOR2_X1 U12101 ( .A(n12192), .B(n12193), .Z(n11985) );
  XOR2_X1 U12102 ( .A(n12194), .B(n12195), .Z(n12193) );
  OR2_X1 U12103 ( .A1(n8978), .A2(n8280), .ZN(n11991) );
  XOR2_X1 U12104 ( .A(n12196), .B(n12197), .Z(n11988) );
  XOR2_X1 U12105 ( .A(n12198), .B(n12199), .Z(n12197) );
  OR2_X1 U12106 ( .A1(n8974), .A2(n8280), .ZN(n11995) );
  XOR2_X1 U12107 ( .A(n12200), .B(n12201), .Z(n11992) );
  XOR2_X1 U12108 ( .A(n12202), .B(n8979), .Z(n12201) );
  OR2_X1 U12109 ( .A1(n8970), .A2(n8280), .ZN(n11999) );
  XOR2_X1 U12110 ( .A(n12203), .B(n12204), .Z(n11996) );
  XOR2_X1 U12111 ( .A(n12205), .B(n12206), .Z(n12204) );
  OR2_X1 U12112 ( .A1(n8966), .A2(n8280), .ZN(n12003) );
  XOR2_X1 U12113 ( .A(n12207), .B(n12208), .Z(n12000) );
  XOR2_X1 U12114 ( .A(n12209), .B(n12210), .Z(n12208) );
  OR2_X1 U12115 ( .A1(n8962), .A2(n8280), .ZN(n12007) );
  XOR2_X1 U12116 ( .A(n12211), .B(n12212), .Z(n12004) );
  XOR2_X1 U12117 ( .A(n12213), .B(n12214), .Z(n12212) );
  OR2_X1 U12118 ( .A1(n8958), .A2(n8280), .ZN(n12011) );
  XOR2_X1 U12119 ( .A(n12215), .B(n12216), .Z(n12008) );
  XOR2_X1 U12120 ( .A(n12217), .B(n12218), .Z(n12216) );
  OR2_X1 U12121 ( .A1(n8954), .A2(n8280), .ZN(n12015) );
  XOR2_X1 U12122 ( .A(n12219), .B(n12220), .Z(n12012) );
  XOR2_X1 U12123 ( .A(n12221), .B(n12222), .Z(n12220) );
  OR2_X1 U12124 ( .A1(n8950), .A2(n8280), .ZN(n12019) );
  XOR2_X1 U12125 ( .A(n12223), .B(n12224), .Z(n12016) );
  XOR2_X1 U12126 ( .A(n12225), .B(n12226), .Z(n12224) );
  OR2_X1 U12127 ( .A1(n8946), .A2(n8280), .ZN(n12023) );
  XOR2_X1 U12128 ( .A(n12227), .B(n12228), .Z(n12020) );
  XOR2_X1 U12129 ( .A(n12229), .B(n12230), .Z(n12228) );
  OR2_X1 U12130 ( .A1(n8942), .A2(n8280), .ZN(n12027) );
  XOR2_X1 U12131 ( .A(n12231), .B(n12232), .Z(n12024) );
  XOR2_X1 U12132 ( .A(n12233), .B(n12234), .Z(n12232) );
  OR2_X1 U12133 ( .A1(n8938), .A2(n8280), .ZN(n12031) );
  XOR2_X1 U12134 ( .A(n12235), .B(n12236), .Z(n12028) );
  XOR2_X1 U12135 ( .A(n12237), .B(n12238), .Z(n12236) );
  OR2_X1 U12136 ( .A1(n8934), .A2(n8280), .ZN(n12035) );
  XOR2_X1 U12137 ( .A(n12239), .B(n12240), .Z(n12032) );
  XOR2_X1 U12138 ( .A(n12241), .B(n12242), .Z(n12240) );
  OR2_X1 U12139 ( .A1(n8930), .A2(n8280), .ZN(n12039) );
  XOR2_X1 U12140 ( .A(n12243), .B(n12244), .Z(n12036) );
  XOR2_X1 U12141 ( .A(n12245), .B(n12246), .Z(n12244) );
  OR2_X1 U12142 ( .A1(n8926), .A2(n8280), .ZN(n12043) );
  XOR2_X1 U12143 ( .A(n12247), .B(n12248), .Z(n12040) );
  XOR2_X1 U12144 ( .A(n12249), .B(n12250), .Z(n12248) );
  OR2_X1 U12145 ( .A1(n8922), .A2(n8280), .ZN(n12047) );
  XOR2_X1 U12146 ( .A(n12251), .B(n12252), .Z(n12044) );
  XOR2_X1 U12147 ( .A(n12253), .B(n12254), .Z(n12252) );
  OR2_X1 U12148 ( .A1(n8918), .A2(n8280), .ZN(n12051) );
  XOR2_X1 U12149 ( .A(n12255), .B(n12256), .Z(n12048) );
  XOR2_X1 U12150 ( .A(n12257), .B(n12258), .Z(n12256) );
  OR2_X1 U12151 ( .A1(n12052), .A2(n12055), .ZN(n12080) );
  OR2_X1 U12152 ( .A1(n8914), .A2(n8280), .ZN(n12055) );
  XOR2_X1 U12153 ( .A(n12259), .B(n12260), .Z(n12052) );
  XOR2_X1 U12154 ( .A(n12261), .B(n12262), .Z(n12260) );
  OR2_X1 U12155 ( .A1(n12056), .A2(n12059), .ZN(n12077) );
  OR2_X1 U12156 ( .A1(n8910), .A2(n8280), .ZN(n12059) );
  XOR2_X1 U12157 ( .A(n12263), .B(n12264), .Z(n12056) );
  XOR2_X1 U12158 ( .A(n12265), .B(n12266), .Z(n12264) );
  OR2_X1 U12159 ( .A1(n12060), .A2(n12063), .ZN(n12074) );
  OR2_X1 U12160 ( .A1(n8906), .A2(n8280), .ZN(n12063) );
  XOR2_X1 U12161 ( .A(n12267), .B(n12268), .Z(n12060) );
  XOR2_X1 U12162 ( .A(n12269), .B(n12270), .Z(n12268) );
  OR2_X1 U12163 ( .A1(n12064), .A2(n12067), .ZN(n12071) );
  OR2_X1 U12164 ( .A1(n8902), .A2(n8280), .ZN(n12067) );
  XOR2_X1 U12165 ( .A(n12271), .B(n12272), .Z(n12064) );
  XOR2_X1 U12166 ( .A(n12273), .B(n12274), .Z(n12272) );
  XOR2_X1 U12167 ( .A(n11846), .B(n12275), .Z(n11839) );
  XOR2_X1 U12168 ( .A(n11849), .B(n11847), .Z(n12275) );
  OR2_X1 U12169 ( .A1(n8902), .A2(n8308), .ZN(n11847) );
  OR2_X1 U12170 ( .A1(n12276), .A2(n12277), .ZN(n11849) );
  AND2_X1 U12171 ( .A1(n12271), .A2(n12274), .ZN(n12277) );
  AND2_X1 U12172 ( .A1(n12278), .A2(n12273), .ZN(n12276) );
  OR2_X1 U12173 ( .A1(n12279), .A2(n12280), .ZN(n12273) );
  AND2_X1 U12174 ( .A1(n12267), .A2(n12270), .ZN(n12280) );
  AND2_X1 U12175 ( .A1(n12281), .A2(n12269), .ZN(n12279) );
  OR2_X1 U12176 ( .A1(n12282), .A2(n12283), .ZN(n12269) );
  AND2_X1 U12177 ( .A1(n12263), .A2(n12266), .ZN(n12283) );
  AND2_X1 U12178 ( .A1(n12284), .A2(n12265), .ZN(n12282) );
  OR2_X1 U12179 ( .A1(n12285), .A2(n12286), .ZN(n12265) );
  AND2_X1 U12180 ( .A1(n12259), .A2(n12262), .ZN(n12286) );
  AND2_X1 U12181 ( .A1(n12287), .A2(n12261), .ZN(n12285) );
  OR2_X1 U12182 ( .A1(n12288), .A2(n12289), .ZN(n12261) );
  AND2_X1 U12183 ( .A1(n12255), .A2(n12258), .ZN(n12289) );
  AND2_X1 U12184 ( .A1(n12290), .A2(n12257), .ZN(n12288) );
  OR2_X1 U12185 ( .A1(n12291), .A2(n12292), .ZN(n12257) );
  AND2_X1 U12186 ( .A1(n12254), .A2(n12253), .ZN(n12292) );
  AND2_X1 U12187 ( .A1(n12251), .A2(n12293), .ZN(n12291) );
  OR2_X1 U12188 ( .A1(n12254), .A2(n12253), .ZN(n12293) );
  OR2_X1 U12189 ( .A1(n12294), .A2(n12295), .ZN(n12253) );
  AND2_X1 U12190 ( .A1(n12250), .A2(n12249), .ZN(n12295) );
  AND2_X1 U12191 ( .A1(n12247), .A2(n12296), .ZN(n12294) );
  OR2_X1 U12192 ( .A1(n12250), .A2(n12249), .ZN(n12296) );
  OR2_X1 U12193 ( .A1(n12297), .A2(n12298), .ZN(n12249) );
  AND2_X1 U12194 ( .A1(n12246), .A2(n12245), .ZN(n12298) );
  AND2_X1 U12195 ( .A1(n12243), .A2(n12299), .ZN(n12297) );
  OR2_X1 U12196 ( .A1(n12246), .A2(n12245), .ZN(n12299) );
  OR2_X1 U12197 ( .A1(n12300), .A2(n12301), .ZN(n12245) );
  AND2_X1 U12198 ( .A1(n12242), .A2(n12241), .ZN(n12301) );
  AND2_X1 U12199 ( .A1(n12239), .A2(n12302), .ZN(n12300) );
  OR2_X1 U12200 ( .A1(n12242), .A2(n12241), .ZN(n12302) );
  OR2_X1 U12201 ( .A1(n12303), .A2(n12304), .ZN(n12241) );
  AND2_X1 U12202 ( .A1(n12238), .A2(n12237), .ZN(n12304) );
  AND2_X1 U12203 ( .A1(n12235), .A2(n12305), .ZN(n12303) );
  OR2_X1 U12204 ( .A1(n12238), .A2(n12237), .ZN(n12305) );
  OR2_X1 U12205 ( .A1(n12306), .A2(n12307), .ZN(n12237) );
  AND2_X1 U12206 ( .A1(n12234), .A2(n12233), .ZN(n12307) );
  AND2_X1 U12207 ( .A1(n12231), .A2(n12308), .ZN(n12306) );
  OR2_X1 U12208 ( .A1(n12234), .A2(n12233), .ZN(n12308) );
  OR2_X1 U12209 ( .A1(n12309), .A2(n12310), .ZN(n12233) );
  AND2_X1 U12210 ( .A1(n12230), .A2(n12229), .ZN(n12310) );
  AND2_X1 U12211 ( .A1(n12227), .A2(n12311), .ZN(n12309) );
  OR2_X1 U12212 ( .A1(n12230), .A2(n12229), .ZN(n12311) );
  OR2_X1 U12213 ( .A1(n12312), .A2(n12313), .ZN(n12229) );
  AND2_X1 U12214 ( .A1(n12226), .A2(n12225), .ZN(n12313) );
  AND2_X1 U12215 ( .A1(n12223), .A2(n12314), .ZN(n12312) );
  OR2_X1 U12216 ( .A1(n12226), .A2(n12225), .ZN(n12314) );
  OR2_X1 U12217 ( .A1(n12315), .A2(n12316), .ZN(n12225) );
  AND2_X1 U12218 ( .A1(n12222), .A2(n12221), .ZN(n12316) );
  AND2_X1 U12219 ( .A1(n12219), .A2(n12317), .ZN(n12315) );
  OR2_X1 U12220 ( .A1(n12222), .A2(n12221), .ZN(n12317) );
  OR2_X1 U12221 ( .A1(n12318), .A2(n12319), .ZN(n12221) );
  AND2_X1 U12222 ( .A1(n12218), .A2(n12217), .ZN(n12319) );
  AND2_X1 U12223 ( .A1(n12215), .A2(n12320), .ZN(n12318) );
  OR2_X1 U12224 ( .A1(n12218), .A2(n12217), .ZN(n12320) );
  OR2_X1 U12225 ( .A1(n12321), .A2(n12322), .ZN(n12217) );
  AND2_X1 U12226 ( .A1(n12214), .A2(n12213), .ZN(n12322) );
  AND2_X1 U12227 ( .A1(n12211), .A2(n12323), .ZN(n12321) );
  OR2_X1 U12228 ( .A1(n12214), .A2(n12213), .ZN(n12323) );
  OR2_X1 U12229 ( .A1(n12324), .A2(n12325), .ZN(n12213) );
  AND2_X1 U12230 ( .A1(n12210), .A2(n12209), .ZN(n12325) );
  AND2_X1 U12231 ( .A1(n12207), .A2(n12326), .ZN(n12324) );
  OR2_X1 U12232 ( .A1(n12210), .A2(n12209), .ZN(n12326) );
  OR2_X1 U12233 ( .A1(n12327), .A2(n12328), .ZN(n12209) );
  AND2_X1 U12234 ( .A1(n12206), .A2(n12205), .ZN(n12328) );
  AND2_X1 U12235 ( .A1(n12203), .A2(n12329), .ZN(n12327) );
  OR2_X1 U12236 ( .A1(n12206), .A2(n12205), .ZN(n12329) );
  OR2_X1 U12237 ( .A1(n12330), .A2(n12331), .ZN(n12205) );
  AND2_X1 U12238 ( .A1(n8979), .A2(n12202), .ZN(n12331) );
  AND2_X1 U12239 ( .A1(n12200), .A2(n12332), .ZN(n12330) );
  OR2_X1 U12240 ( .A1(n8979), .A2(n12202), .ZN(n12332) );
  OR2_X1 U12241 ( .A1(n12333), .A2(n12334), .ZN(n12202) );
  AND2_X1 U12242 ( .A1(n12199), .A2(n12198), .ZN(n12334) );
  AND2_X1 U12243 ( .A1(n12196), .A2(n12335), .ZN(n12333) );
  OR2_X1 U12244 ( .A1(n12199), .A2(n12198), .ZN(n12335) );
  OR2_X1 U12245 ( .A1(n12336), .A2(n12337), .ZN(n12198) );
  AND2_X1 U12246 ( .A1(n12195), .A2(n12194), .ZN(n12337) );
  AND2_X1 U12247 ( .A1(n12192), .A2(n12338), .ZN(n12336) );
  OR2_X1 U12248 ( .A1(n12195), .A2(n12194), .ZN(n12338) );
  OR2_X1 U12249 ( .A1(n12339), .A2(n12340), .ZN(n12194) );
  AND2_X1 U12250 ( .A1(n12191), .A2(n12190), .ZN(n12340) );
  AND2_X1 U12251 ( .A1(n12188), .A2(n12341), .ZN(n12339) );
  OR2_X1 U12252 ( .A1(n12191), .A2(n12190), .ZN(n12341) );
  OR2_X1 U12253 ( .A1(n12342), .A2(n12343), .ZN(n12190) );
  AND2_X1 U12254 ( .A1(n12187), .A2(n12186), .ZN(n12343) );
  AND2_X1 U12255 ( .A1(n12184), .A2(n12344), .ZN(n12342) );
  OR2_X1 U12256 ( .A1(n12187), .A2(n12186), .ZN(n12344) );
  OR2_X1 U12257 ( .A1(n12345), .A2(n12346), .ZN(n12186) );
  AND2_X1 U12258 ( .A1(n12183), .A2(n12182), .ZN(n12346) );
  AND2_X1 U12259 ( .A1(n12180), .A2(n12347), .ZN(n12345) );
  OR2_X1 U12260 ( .A1(n12183), .A2(n12182), .ZN(n12347) );
  OR2_X1 U12261 ( .A1(n12348), .A2(n12349), .ZN(n12182) );
  AND2_X1 U12262 ( .A1(n12179), .A2(n12178), .ZN(n12349) );
  AND2_X1 U12263 ( .A1(n12176), .A2(n12350), .ZN(n12348) );
  OR2_X1 U12264 ( .A1(n12179), .A2(n12178), .ZN(n12350) );
  OR2_X1 U12265 ( .A1(n12351), .A2(n12352), .ZN(n12178) );
  AND2_X1 U12266 ( .A1(n12175), .A2(n12174), .ZN(n12352) );
  AND2_X1 U12267 ( .A1(n12172), .A2(n12353), .ZN(n12351) );
  OR2_X1 U12268 ( .A1(n12175), .A2(n12174), .ZN(n12353) );
  OR2_X1 U12269 ( .A1(n12354), .A2(n12355), .ZN(n12174) );
  AND2_X1 U12270 ( .A1(n12171), .A2(n12170), .ZN(n12355) );
  AND2_X1 U12271 ( .A1(n12168), .A2(n12356), .ZN(n12354) );
  OR2_X1 U12272 ( .A1(n12171), .A2(n12170), .ZN(n12356) );
  OR2_X1 U12273 ( .A1(n12357), .A2(n12358), .ZN(n12170) );
  AND2_X1 U12274 ( .A1(n12165), .A2(n12166), .ZN(n12358) );
  AND2_X1 U12275 ( .A1(n12359), .A2(n12360), .ZN(n12357) );
  OR2_X1 U12276 ( .A1(n12165), .A2(n12166), .ZN(n12360) );
  OR2_X1 U12277 ( .A1(n9984), .A2(n12361), .ZN(n12166) );
  OR2_X1 U12278 ( .A1(n8308), .A2(n8336), .ZN(n12361) );
  OR2_X1 U12279 ( .A1(n9014), .A2(n8308), .ZN(n12165) );
  INV_X1 U12280 ( .A(n12167), .ZN(n12359) );
  OR2_X1 U12281 ( .A1(n12362), .A2(n12363), .ZN(n12167) );
  AND2_X1 U12282 ( .A1(b_19_), .A2(n12364), .ZN(n12363) );
  OR2_X1 U12283 ( .A1(n12365), .A2(n9989), .ZN(n12364) );
  AND2_X1 U12284 ( .A1(a_30_), .A2(n8971), .ZN(n12365) );
  AND2_X1 U12285 ( .A1(b_18_), .A2(n12366), .ZN(n12362) );
  OR2_X1 U12286 ( .A1(n12367), .A2(n8021), .ZN(n12366) );
  AND2_X1 U12287 ( .A1(a_31_), .A2(n8336), .ZN(n12367) );
  OR2_X1 U12288 ( .A1(n9010), .A2(n8308), .ZN(n12171) );
  XOR2_X1 U12289 ( .A(n12368), .B(n12369), .Z(n12168) );
  XNOR2_X1 U12290 ( .A(n12370), .B(n12371), .ZN(n12368) );
  OR2_X1 U12291 ( .A1(n9006), .A2(n8308), .ZN(n12175) );
  XOR2_X1 U12292 ( .A(n12372), .B(n12373), .Z(n12172) );
  XOR2_X1 U12293 ( .A(n12374), .B(n12375), .Z(n12373) );
  OR2_X1 U12294 ( .A1(n9002), .A2(n8308), .ZN(n12179) );
  XOR2_X1 U12295 ( .A(n12376), .B(n12377), .Z(n12176) );
  XOR2_X1 U12296 ( .A(n12378), .B(n12379), .Z(n12377) );
  OR2_X1 U12297 ( .A1(n8998), .A2(n8308), .ZN(n12183) );
  XOR2_X1 U12298 ( .A(n12380), .B(n12381), .Z(n12180) );
  XOR2_X1 U12299 ( .A(n12382), .B(n12383), .Z(n12381) );
  OR2_X1 U12300 ( .A1(n8994), .A2(n8308), .ZN(n12187) );
  XOR2_X1 U12301 ( .A(n12384), .B(n12385), .Z(n12184) );
  XOR2_X1 U12302 ( .A(n12386), .B(n12387), .Z(n12385) );
  OR2_X1 U12303 ( .A1(n8990), .A2(n8308), .ZN(n12191) );
  XOR2_X1 U12304 ( .A(n12388), .B(n12389), .Z(n12188) );
  XOR2_X1 U12305 ( .A(n12390), .B(n12391), .Z(n12389) );
  OR2_X1 U12306 ( .A1(n8986), .A2(n8308), .ZN(n12195) );
  XOR2_X1 U12307 ( .A(n12392), .B(n12393), .Z(n12192) );
  XOR2_X1 U12308 ( .A(n12394), .B(n12395), .Z(n12393) );
  OR2_X1 U12309 ( .A1(n8982), .A2(n8308), .ZN(n12199) );
  XOR2_X1 U12310 ( .A(n12396), .B(n12397), .Z(n12196) );
  XOR2_X1 U12311 ( .A(n12398), .B(n12399), .Z(n12397) );
  OR2_X1 U12312 ( .A1(n8978), .A2(n8308), .ZN(n8979) );
  XOR2_X1 U12313 ( .A(n12400), .B(n12401), .Z(n12200) );
  XOR2_X1 U12314 ( .A(n12402), .B(n12403), .Z(n12401) );
  OR2_X1 U12315 ( .A1(n8974), .A2(n8308), .ZN(n12206) );
  XOR2_X1 U12316 ( .A(n12404), .B(n12405), .Z(n12203) );
  XOR2_X1 U12317 ( .A(n12406), .B(n12407), .Z(n12405) );
  OR2_X1 U12318 ( .A1(n8970), .A2(n8308), .ZN(n12210) );
  XOR2_X1 U12319 ( .A(n12408), .B(n12409), .Z(n12207) );
  XOR2_X1 U12320 ( .A(n12410), .B(n8975), .Z(n12409) );
  OR2_X1 U12321 ( .A1(n8966), .A2(n8308), .ZN(n12214) );
  XOR2_X1 U12322 ( .A(n12411), .B(n12412), .Z(n12211) );
  XOR2_X1 U12323 ( .A(n12413), .B(n12414), .Z(n12412) );
  OR2_X1 U12324 ( .A1(n8962), .A2(n8308), .ZN(n12218) );
  XOR2_X1 U12325 ( .A(n12415), .B(n12416), .Z(n12215) );
  XOR2_X1 U12326 ( .A(n12417), .B(n12418), .Z(n12416) );
  OR2_X1 U12327 ( .A1(n8958), .A2(n8308), .ZN(n12222) );
  XOR2_X1 U12328 ( .A(n12419), .B(n12420), .Z(n12219) );
  XOR2_X1 U12329 ( .A(n12421), .B(n12422), .Z(n12420) );
  OR2_X1 U12330 ( .A1(n8954), .A2(n8308), .ZN(n12226) );
  XOR2_X1 U12331 ( .A(n12423), .B(n12424), .Z(n12223) );
  XOR2_X1 U12332 ( .A(n12425), .B(n12426), .Z(n12424) );
  OR2_X1 U12333 ( .A1(n8950), .A2(n8308), .ZN(n12230) );
  XOR2_X1 U12334 ( .A(n12427), .B(n12428), .Z(n12227) );
  XOR2_X1 U12335 ( .A(n12429), .B(n12430), .Z(n12428) );
  OR2_X1 U12336 ( .A1(n8946), .A2(n8308), .ZN(n12234) );
  XOR2_X1 U12337 ( .A(n12431), .B(n12432), .Z(n12231) );
  XOR2_X1 U12338 ( .A(n12433), .B(n12434), .Z(n12432) );
  OR2_X1 U12339 ( .A1(n8942), .A2(n8308), .ZN(n12238) );
  XOR2_X1 U12340 ( .A(n12435), .B(n12436), .Z(n12235) );
  XOR2_X1 U12341 ( .A(n12437), .B(n12438), .Z(n12436) );
  OR2_X1 U12342 ( .A1(n8938), .A2(n8308), .ZN(n12242) );
  XOR2_X1 U12343 ( .A(n12439), .B(n12440), .Z(n12239) );
  XOR2_X1 U12344 ( .A(n12441), .B(n12442), .Z(n12440) );
  OR2_X1 U12345 ( .A1(n8934), .A2(n8308), .ZN(n12246) );
  XOR2_X1 U12346 ( .A(n12443), .B(n12444), .Z(n12243) );
  XOR2_X1 U12347 ( .A(n12445), .B(n12446), .Z(n12444) );
  OR2_X1 U12348 ( .A1(n8930), .A2(n8308), .ZN(n12250) );
  XOR2_X1 U12349 ( .A(n12447), .B(n12448), .Z(n12247) );
  XOR2_X1 U12350 ( .A(n12449), .B(n12450), .Z(n12448) );
  OR2_X1 U12351 ( .A1(n8926), .A2(n8308), .ZN(n12254) );
  XOR2_X1 U12352 ( .A(n12451), .B(n12452), .Z(n12251) );
  XOR2_X1 U12353 ( .A(n12453), .B(n12454), .Z(n12452) );
  OR2_X1 U12354 ( .A1(n12255), .A2(n12258), .ZN(n12290) );
  OR2_X1 U12355 ( .A1(n8922), .A2(n8308), .ZN(n12258) );
  XOR2_X1 U12356 ( .A(n12455), .B(n12456), .Z(n12255) );
  XOR2_X1 U12357 ( .A(n12457), .B(n12458), .Z(n12456) );
  OR2_X1 U12358 ( .A1(n12259), .A2(n12262), .ZN(n12287) );
  OR2_X1 U12359 ( .A1(n8918), .A2(n8308), .ZN(n12262) );
  XOR2_X1 U12360 ( .A(n12459), .B(n12460), .Z(n12259) );
  XOR2_X1 U12361 ( .A(n12461), .B(n12462), .Z(n12460) );
  OR2_X1 U12362 ( .A1(n12263), .A2(n12266), .ZN(n12284) );
  OR2_X1 U12363 ( .A1(n8914), .A2(n8308), .ZN(n12266) );
  XOR2_X1 U12364 ( .A(n12463), .B(n12464), .Z(n12263) );
  XOR2_X1 U12365 ( .A(n12465), .B(n12466), .Z(n12464) );
  OR2_X1 U12366 ( .A1(n12267), .A2(n12270), .ZN(n12281) );
  OR2_X1 U12367 ( .A1(n8910), .A2(n8308), .ZN(n12270) );
  XOR2_X1 U12368 ( .A(n12467), .B(n12468), .Z(n12267) );
  XOR2_X1 U12369 ( .A(n12469), .B(n12470), .Z(n12468) );
  OR2_X1 U12370 ( .A1(n12271), .A2(n12274), .ZN(n12278) );
  OR2_X1 U12371 ( .A1(n8906), .A2(n8308), .ZN(n12274) );
  XOR2_X1 U12372 ( .A(n12471), .B(n12472), .Z(n12271) );
  XOR2_X1 U12373 ( .A(n12473), .B(n12474), .Z(n12472) );
  XOR2_X1 U12374 ( .A(n12475), .B(n12476), .Z(n11846) );
  XOR2_X1 U12375 ( .A(n12477), .B(n12478), .Z(n12476) );
  AND2_X1 U12376 ( .A1(n9788), .A2(n9139), .ZN(n9786) );
  XOR2_X1 U12377 ( .A(n12479), .B(n12480), .Z(n9139) );
  INV_X1 U12378 ( .A(n9138), .ZN(n9788) );
  OR2_X1 U12379 ( .A1(n9792), .A2(n9793), .ZN(n9138) );
  OR2_X1 U12380 ( .A1(n12481), .A2(n12482), .ZN(n9793) );
  AND2_X1 U12381 ( .A1(n9809), .A2(n9812), .ZN(n12482) );
  AND2_X1 U12382 ( .A1(n12483), .A2(n9811), .ZN(n12481) );
  OR2_X1 U12383 ( .A1(n12484), .A2(n12485), .ZN(n9811) );
  AND2_X1 U12384 ( .A1(n11850), .A2(n11853), .ZN(n12485) );
  AND2_X1 U12385 ( .A1(n12486), .A2(n11852), .ZN(n12484) );
  OR2_X1 U12386 ( .A1(n12487), .A2(n12488), .ZN(n11852) );
  AND2_X1 U12387 ( .A1(n12475), .A2(n12478), .ZN(n12488) );
  AND2_X1 U12388 ( .A1(n12489), .A2(n12477), .ZN(n12487) );
  OR2_X1 U12389 ( .A1(n12490), .A2(n12491), .ZN(n12477) );
  AND2_X1 U12390 ( .A1(n12471), .A2(n12474), .ZN(n12491) );
  AND2_X1 U12391 ( .A1(n12492), .A2(n12473), .ZN(n12490) );
  OR2_X1 U12392 ( .A1(n12493), .A2(n12494), .ZN(n12473) );
  AND2_X1 U12393 ( .A1(n12467), .A2(n12470), .ZN(n12494) );
  AND2_X1 U12394 ( .A1(n12495), .A2(n12469), .ZN(n12493) );
  OR2_X1 U12395 ( .A1(n12496), .A2(n12497), .ZN(n12469) );
  AND2_X1 U12396 ( .A1(n12463), .A2(n12466), .ZN(n12497) );
  AND2_X1 U12397 ( .A1(n12498), .A2(n12465), .ZN(n12496) );
  OR2_X1 U12398 ( .A1(n12499), .A2(n12500), .ZN(n12465) );
  AND2_X1 U12399 ( .A1(n12459), .A2(n12462), .ZN(n12500) );
  AND2_X1 U12400 ( .A1(n12501), .A2(n12461), .ZN(n12499) );
  OR2_X1 U12401 ( .A1(n12502), .A2(n12503), .ZN(n12461) );
  AND2_X1 U12402 ( .A1(n12455), .A2(n12458), .ZN(n12503) );
  AND2_X1 U12403 ( .A1(n12504), .A2(n12457), .ZN(n12502) );
  OR2_X1 U12404 ( .A1(n12505), .A2(n12506), .ZN(n12457) );
  AND2_X1 U12405 ( .A1(n12451), .A2(n12454), .ZN(n12506) );
  AND2_X1 U12406 ( .A1(n12507), .A2(n12453), .ZN(n12505) );
  OR2_X1 U12407 ( .A1(n12508), .A2(n12509), .ZN(n12453) );
  AND2_X1 U12408 ( .A1(n12450), .A2(n12449), .ZN(n12509) );
  AND2_X1 U12409 ( .A1(n12447), .A2(n12510), .ZN(n12508) );
  OR2_X1 U12410 ( .A1(n12450), .A2(n12449), .ZN(n12510) );
  OR2_X1 U12411 ( .A1(n12511), .A2(n12512), .ZN(n12449) );
  AND2_X1 U12412 ( .A1(n12446), .A2(n12445), .ZN(n12512) );
  AND2_X1 U12413 ( .A1(n12443), .A2(n12513), .ZN(n12511) );
  OR2_X1 U12414 ( .A1(n12446), .A2(n12445), .ZN(n12513) );
  OR2_X1 U12415 ( .A1(n12514), .A2(n12515), .ZN(n12445) );
  AND2_X1 U12416 ( .A1(n12442), .A2(n12441), .ZN(n12515) );
  AND2_X1 U12417 ( .A1(n12439), .A2(n12516), .ZN(n12514) );
  OR2_X1 U12418 ( .A1(n12442), .A2(n12441), .ZN(n12516) );
  OR2_X1 U12419 ( .A1(n12517), .A2(n12518), .ZN(n12441) );
  AND2_X1 U12420 ( .A1(n12438), .A2(n12437), .ZN(n12518) );
  AND2_X1 U12421 ( .A1(n12435), .A2(n12519), .ZN(n12517) );
  OR2_X1 U12422 ( .A1(n12438), .A2(n12437), .ZN(n12519) );
  OR2_X1 U12423 ( .A1(n12520), .A2(n12521), .ZN(n12437) );
  AND2_X1 U12424 ( .A1(n12434), .A2(n12433), .ZN(n12521) );
  AND2_X1 U12425 ( .A1(n12431), .A2(n12522), .ZN(n12520) );
  OR2_X1 U12426 ( .A1(n12434), .A2(n12433), .ZN(n12522) );
  OR2_X1 U12427 ( .A1(n12523), .A2(n12524), .ZN(n12433) );
  AND2_X1 U12428 ( .A1(n12430), .A2(n12429), .ZN(n12524) );
  AND2_X1 U12429 ( .A1(n12427), .A2(n12525), .ZN(n12523) );
  OR2_X1 U12430 ( .A1(n12430), .A2(n12429), .ZN(n12525) );
  OR2_X1 U12431 ( .A1(n12526), .A2(n12527), .ZN(n12429) );
  AND2_X1 U12432 ( .A1(n12426), .A2(n12425), .ZN(n12527) );
  AND2_X1 U12433 ( .A1(n12423), .A2(n12528), .ZN(n12526) );
  OR2_X1 U12434 ( .A1(n12426), .A2(n12425), .ZN(n12528) );
  OR2_X1 U12435 ( .A1(n12529), .A2(n12530), .ZN(n12425) );
  AND2_X1 U12436 ( .A1(n12422), .A2(n12421), .ZN(n12530) );
  AND2_X1 U12437 ( .A1(n12419), .A2(n12531), .ZN(n12529) );
  OR2_X1 U12438 ( .A1(n12422), .A2(n12421), .ZN(n12531) );
  OR2_X1 U12439 ( .A1(n12532), .A2(n12533), .ZN(n12421) );
  AND2_X1 U12440 ( .A1(n12418), .A2(n12417), .ZN(n12533) );
  AND2_X1 U12441 ( .A1(n12415), .A2(n12534), .ZN(n12532) );
  OR2_X1 U12442 ( .A1(n12418), .A2(n12417), .ZN(n12534) );
  OR2_X1 U12443 ( .A1(n12535), .A2(n12536), .ZN(n12417) );
  AND2_X1 U12444 ( .A1(n12414), .A2(n12413), .ZN(n12536) );
  AND2_X1 U12445 ( .A1(n12411), .A2(n12537), .ZN(n12535) );
  OR2_X1 U12446 ( .A1(n12414), .A2(n12413), .ZN(n12537) );
  OR2_X1 U12447 ( .A1(n12538), .A2(n12539), .ZN(n12413) );
  AND2_X1 U12448 ( .A1(n8975), .A2(n12410), .ZN(n12539) );
  AND2_X1 U12449 ( .A1(n12408), .A2(n12540), .ZN(n12538) );
  OR2_X1 U12450 ( .A1(n8975), .A2(n12410), .ZN(n12540) );
  OR2_X1 U12451 ( .A1(n12541), .A2(n12542), .ZN(n12410) );
  AND2_X1 U12452 ( .A1(n12407), .A2(n12406), .ZN(n12542) );
  AND2_X1 U12453 ( .A1(n12404), .A2(n12543), .ZN(n12541) );
  OR2_X1 U12454 ( .A1(n12407), .A2(n12406), .ZN(n12543) );
  OR2_X1 U12455 ( .A1(n12544), .A2(n12545), .ZN(n12406) );
  AND2_X1 U12456 ( .A1(n12403), .A2(n12402), .ZN(n12545) );
  AND2_X1 U12457 ( .A1(n12400), .A2(n12546), .ZN(n12544) );
  OR2_X1 U12458 ( .A1(n12403), .A2(n12402), .ZN(n12546) );
  OR2_X1 U12459 ( .A1(n12547), .A2(n12548), .ZN(n12402) );
  AND2_X1 U12460 ( .A1(n12399), .A2(n12398), .ZN(n12548) );
  AND2_X1 U12461 ( .A1(n12396), .A2(n12549), .ZN(n12547) );
  OR2_X1 U12462 ( .A1(n12399), .A2(n12398), .ZN(n12549) );
  OR2_X1 U12463 ( .A1(n12550), .A2(n12551), .ZN(n12398) );
  AND2_X1 U12464 ( .A1(n12395), .A2(n12394), .ZN(n12551) );
  AND2_X1 U12465 ( .A1(n12392), .A2(n12552), .ZN(n12550) );
  OR2_X1 U12466 ( .A1(n12395), .A2(n12394), .ZN(n12552) );
  OR2_X1 U12467 ( .A1(n12553), .A2(n12554), .ZN(n12394) );
  AND2_X1 U12468 ( .A1(n12391), .A2(n12390), .ZN(n12554) );
  AND2_X1 U12469 ( .A1(n12388), .A2(n12555), .ZN(n12553) );
  OR2_X1 U12470 ( .A1(n12391), .A2(n12390), .ZN(n12555) );
  OR2_X1 U12471 ( .A1(n12556), .A2(n12557), .ZN(n12390) );
  AND2_X1 U12472 ( .A1(n12387), .A2(n12386), .ZN(n12557) );
  AND2_X1 U12473 ( .A1(n12384), .A2(n12558), .ZN(n12556) );
  OR2_X1 U12474 ( .A1(n12387), .A2(n12386), .ZN(n12558) );
  OR2_X1 U12475 ( .A1(n12559), .A2(n12560), .ZN(n12386) );
  AND2_X1 U12476 ( .A1(n12383), .A2(n12382), .ZN(n12560) );
  AND2_X1 U12477 ( .A1(n12380), .A2(n12561), .ZN(n12559) );
  OR2_X1 U12478 ( .A1(n12383), .A2(n12382), .ZN(n12561) );
  OR2_X1 U12479 ( .A1(n12562), .A2(n12563), .ZN(n12382) );
  AND2_X1 U12480 ( .A1(n12379), .A2(n12378), .ZN(n12563) );
  AND2_X1 U12481 ( .A1(n12376), .A2(n12564), .ZN(n12562) );
  OR2_X1 U12482 ( .A1(n12379), .A2(n12378), .ZN(n12564) );
  OR2_X1 U12483 ( .A1(n12565), .A2(n12566), .ZN(n12378) );
  AND2_X1 U12484 ( .A1(n12375), .A2(n12374), .ZN(n12566) );
  AND2_X1 U12485 ( .A1(n12372), .A2(n12567), .ZN(n12565) );
  OR2_X1 U12486 ( .A1(n12375), .A2(n12374), .ZN(n12567) );
  OR2_X1 U12487 ( .A1(n12568), .A2(n12569), .ZN(n12374) );
  AND2_X1 U12488 ( .A1(n12369), .A2(n12370), .ZN(n12569) );
  AND2_X1 U12489 ( .A1(n12570), .A2(n12571), .ZN(n12568) );
  OR2_X1 U12490 ( .A1(n12369), .A2(n12370), .ZN(n12571) );
  OR2_X1 U12491 ( .A1(n9984), .A2(n12572), .ZN(n12370) );
  OR2_X1 U12492 ( .A1(n8336), .A2(n8971), .ZN(n12572) );
  OR2_X1 U12493 ( .A1(n9014), .A2(n8336), .ZN(n12369) );
  INV_X1 U12494 ( .A(n12371), .ZN(n12570) );
  OR2_X1 U12495 ( .A1(n12573), .A2(n12574), .ZN(n12371) );
  AND2_X1 U12496 ( .A1(b_18_), .A2(n12575), .ZN(n12574) );
  OR2_X1 U12497 ( .A1(n12576), .A2(n9989), .ZN(n12575) );
  AND2_X1 U12498 ( .A1(a_30_), .A2(n8967), .ZN(n12576) );
  AND2_X1 U12499 ( .A1(b_17_), .A2(n12577), .ZN(n12573) );
  OR2_X1 U12500 ( .A1(n12578), .A2(n8021), .ZN(n12577) );
  AND2_X1 U12501 ( .A1(a_31_), .A2(n8971), .ZN(n12578) );
  OR2_X1 U12502 ( .A1(n9010), .A2(n8336), .ZN(n12375) );
  XOR2_X1 U12503 ( .A(n12579), .B(n12580), .Z(n12372) );
  XNOR2_X1 U12504 ( .A(n12581), .B(n12582), .ZN(n12579) );
  OR2_X1 U12505 ( .A1(n9006), .A2(n8336), .ZN(n12379) );
  XOR2_X1 U12506 ( .A(n12583), .B(n12584), .Z(n12376) );
  XOR2_X1 U12507 ( .A(n12585), .B(n12586), .Z(n12584) );
  OR2_X1 U12508 ( .A1(n9002), .A2(n8336), .ZN(n12383) );
  XOR2_X1 U12509 ( .A(n12587), .B(n12588), .Z(n12380) );
  XOR2_X1 U12510 ( .A(n12589), .B(n12590), .Z(n12588) );
  OR2_X1 U12511 ( .A1(n8998), .A2(n8336), .ZN(n12387) );
  XOR2_X1 U12512 ( .A(n12591), .B(n12592), .Z(n12384) );
  XOR2_X1 U12513 ( .A(n12593), .B(n12594), .Z(n12592) );
  OR2_X1 U12514 ( .A1(n8994), .A2(n8336), .ZN(n12391) );
  XOR2_X1 U12515 ( .A(n12595), .B(n12596), .Z(n12388) );
  XOR2_X1 U12516 ( .A(n12597), .B(n12598), .Z(n12596) );
  OR2_X1 U12517 ( .A1(n8990), .A2(n8336), .ZN(n12395) );
  XOR2_X1 U12518 ( .A(n12599), .B(n12600), .Z(n12392) );
  XOR2_X1 U12519 ( .A(n12601), .B(n12602), .Z(n12600) );
  OR2_X1 U12520 ( .A1(n8986), .A2(n8336), .ZN(n12399) );
  XOR2_X1 U12521 ( .A(n12603), .B(n12604), .Z(n12396) );
  XOR2_X1 U12522 ( .A(n12605), .B(n12606), .Z(n12604) );
  OR2_X1 U12523 ( .A1(n8982), .A2(n8336), .ZN(n12403) );
  XOR2_X1 U12524 ( .A(n12607), .B(n12608), .Z(n12400) );
  XOR2_X1 U12525 ( .A(n12609), .B(n12610), .Z(n12608) );
  OR2_X1 U12526 ( .A1(n8978), .A2(n8336), .ZN(n12407) );
  XOR2_X1 U12527 ( .A(n12611), .B(n12612), .Z(n12404) );
  XOR2_X1 U12528 ( .A(n12613), .B(n12614), .Z(n12612) );
  OR2_X1 U12529 ( .A1(n8974), .A2(n8336), .ZN(n8975) );
  XOR2_X1 U12530 ( .A(n12615), .B(n12616), .Z(n12408) );
  XOR2_X1 U12531 ( .A(n12617), .B(n12618), .Z(n12616) );
  OR2_X1 U12532 ( .A1(n8970), .A2(n8336), .ZN(n12414) );
  XOR2_X1 U12533 ( .A(n12619), .B(n12620), .Z(n12411) );
  XOR2_X1 U12534 ( .A(n12621), .B(n12622), .Z(n12620) );
  OR2_X1 U12535 ( .A1(n8966), .A2(n8336), .ZN(n12418) );
  XOR2_X1 U12536 ( .A(n12623), .B(n12624), .Z(n12415) );
  XOR2_X1 U12537 ( .A(n12625), .B(n8360), .Z(n12624) );
  OR2_X1 U12538 ( .A1(n8962), .A2(n8336), .ZN(n12422) );
  XOR2_X1 U12539 ( .A(n12626), .B(n12627), .Z(n12419) );
  XOR2_X1 U12540 ( .A(n12628), .B(n12629), .Z(n12627) );
  OR2_X1 U12541 ( .A1(n8958), .A2(n8336), .ZN(n12426) );
  XOR2_X1 U12542 ( .A(n12630), .B(n12631), .Z(n12423) );
  XOR2_X1 U12543 ( .A(n12632), .B(n12633), .Z(n12631) );
  OR2_X1 U12544 ( .A1(n8954), .A2(n8336), .ZN(n12430) );
  XOR2_X1 U12545 ( .A(n12634), .B(n12635), .Z(n12427) );
  XOR2_X1 U12546 ( .A(n12636), .B(n12637), .Z(n12635) );
  OR2_X1 U12547 ( .A1(n8950), .A2(n8336), .ZN(n12434) );
  XOR2_X1 U12548 ( .A(n12638), .B(n12639), .Z(n12431) );
  XOR2_X1 U12549 ( .A(n12640), .B(n12641), .Z(n12639) );
  OR2_X1 U12550 ( .A1(n8946), .A2(n8336), .ZN(n12438) );
  XOR2_X1 U12551 ( .A(n12642), .B(n12643), .Z(n12435) );
  XOR2_X1 U12552 ( .A(n12644), .B(n12645), .Z(n12643) );
  OR2_X1 U12553 ( .A1(n8942), .A2(n8336), .ZN(n12442) );
  XOR2_X1 U12554 ( .A(n12646), .B(n12647), .Z(n12439) );
  XOR2_X1 U12555 ( .A(n12648), .B(n12649), .Z(n12647) );
  OR2_X1 U12556 ( .A1(n8938), .A2(n8336), .ZN(n12446) );
  XOR2_X1 U12557 ( .A(n12650), .B(n12651), .Z(n12443) );
  XOR2_X1 U12558 ( .A(n12652), .B(n12653), .Z(n12651) );
  OR2_X1 U12559 ( .A1(n8934), .A2(n8336), .ZN(n12450) );
  XOR2_X1 U12560 ( .A(n12654), .B(n12655), .Z(n12447) );
  XOR2_X1 U12561 ( .A(n12656), .B(n12657), .Z(n12655) );
  OR2_X1 U12562 ( .A1(n12451), .A2(n12454), .ZN(n12507) );
  OR2_X1 U12563 ( .A1(n8930), .A2(n8336), .ZN(n12454) );
  XOR2_X1 U12564 ( .A(n12658), .B(n12659), .Z(n12451) );
  XOR2_X1 U12565 ( .A(n12660), .B(n12661), .Z(n12659) );
  OR2_X1 U12566 ( .A1(n12455), .A2(n12458), .ZN(n12504) );
  OR2_X1 U12567 ( .A1(n8926), .A2(n8336), .ZN(n12458) );
  XOR2_X1 U12568 ( .A(n12662), .B(n12663), .Z(n12455) );
  XOR2_X1 U12569 ( .A(n12664), .B(n12665), .Z(n12663) );
  OR2_X1 U12570 ( .A1(n12459), .A2(n12462), .ZN(n12501) );
  OR2_X1 U12571 ( .A1(n8922), .A2(n8336), .ZN(n12462) );
  XOR2_X1 U12572 ( .A(n12666), .B(n12667), .Z(n12459) );
  XOR2_X1 U12573 ( .A(n12668), .B(n12669), .Z(n12667) );
  OR2_X1 U12574 ( .A1(n12463), .A2(n12466), .ZN(n12498) );
  OR2_X1 U12575 ( .A1(n8918), .A2(n8336), .ZN(n12466) );
  XOR2_X1 U12576 ( .A(n12670), .B(n12671), .Z(n12463) );
  XOR2_X1 U12577 ( .A(n12672), .B(n12673), .Z(n12671) );
  OR2_X1 U12578 ( .A1(n12467), .A2(n12470), .ZN(n12495) );
  OR2_X1 U12579 ( .A1(n8914), .A2(n8336), .ZN(n12470) );
  XOR2_X1 U12580 ( .A(n12674), .B(n12675), .Z(n12467) );
  XOR2_X1 U12581 ( .A(n12676), .B(n12677), .Z(n12675) );
  OR2_X1 U12582 ( .A1(n12471), .A2(n12474), .ZN(n12492) );
  OR2_X1 U12583 ( .A1(n8910), .A2(n8336), .ZN(n12474) );
  XOR2_X1 U12584 ( .A(n12678), .B(n12679), .Z(n12471) );
  XOR2_X1 U12585 ( .A(n12680), .B(n12681), .Z(n12679) );
  OR2_X1 U12586 ( .A1(n12475), .A2(n12478), .ZN(n12489) );
  OR2_X1 U12587 ( .A1(n8906), .A2(n8336), .ZN(n12478) );
  XOR2_X1 U12588 ( .A(n12682), .B(n12683), .Z(n12475) );
  XOR2_X1 U12589 ( .A(n12684), .B(n12685), .Z(n12683) );
  OR2_X1 U12590 ( .A1(n11850), .A2(n11853), .ZN(n12486) );
  OR2_X1 U12591 ( .A1(n8902), .A2(n8336), .ZN(n11853) );
  XOR2_X1 U12592 ( .A(n12686), .B(n12687), .Z(n11850) );
  XOR2_X1 U12593 ( .A(n12688), .B(n12689), .Z(n12687) );
  OR2_X1 U12594 ( .A1(n9809), .A2(n9812), .ZN(n12483) );
  OR2_X1 U12595 ( .A1(n9297), .A2(n8336), .ZN(n9812) );
  XOR2_X1 U12596 ( .A(n12690), .B(n12691), .Z(n9809) );
  XOR2_X1 U12597 ( .A(n12692), .B(n12693), .Z(n12691) );
  XOR2_X1 U12598 ( .A(n12694), .B(n12695), .Z(n9792) );
  XOR2_X1 U12599 ( .A(n12696), .B(n12697), .Z(n12695) );
  OR2_X1 U12600 ( .A1(n9781), .A2(n12698), .ZN(n9144) );
  XOR2_X1 U12601 ( .A(n9785), .B(n9784), .Z(n12698) );
  XOR2_X1 U12602 ( .A(n9765), .B(n12699), .Z(n9784) );
  XOR2_X1 U12603 ( .A(n9764), .B(n9763), .Z(n12699) );
  OR2_X1 U12604 ( .A1(n9297), .A2(n8963), .ZN(n9763) );
  OR2_X1 U12605 ( .A1(n12700), .A2(n12701), .ZN(n9764) );
  AND2_X1 U12606 ( .A1(n12702), .A2(n12703), .ZN(n12701) );
  AND2_X1 U12607 ( .A1(n12704), .A2(n12705), .ZN(n12700) );
  OR2_X1 U12608 ( .A1(n12702), .A2(n12703), .ZN(n12705) );
  XOR2_X1 U12609 ( .A(n9772), .B(n12706), .Z(n9765) );
  XOR2_X1 U12610 ( .A(n9771), .B(n9770), .Z(n12706) );
  OR2_X1 U12611 ( .A1(n8902), .A2(n8959), .ZN(n9770) );
  OR2_X1 U12612 ( .A1(n12707), .A2(n12708), .ZN(n9771) );
  AND2_X1 U12613 ( .A1(n12709), .A2(n12710), .ZN(n12708) );
  AND2_X1 U12614 ( .A1(n12711), .A2(n12712), .ZN(n12707) );
  OR2_X1 U12615 ( .A1(n12710), .A2(n12709), .ZN(n12712) );
  XOR2_X1 U12616 ( .A(n12713), .B(n12714), .Z(n9772) );
  XOR2_X1 U12617 ( .A(n12715), .B(n12716), .Z(n12714) );
  OR2_X1 U12618 ( .A1(n12717), .A2(n12718), .ZN(n9785) );
  AND2_X1 U12619 ( .A1(n12719), .A2(n12720), .ZN(n12718) );
  AND2_X1 U12620 ( .A1(n12721), .A2(n12722), .ZN(n12717) );
  OR2_X1 U12621 ( .A1(n12719), .A2(n12720), .ZN(n12722) );
  AND2_X1 U12622 ( .A1(n12479), .A2(n12480), .ZN(n9781) );
  INV_X1 U12623 ( .A(n12723), .ZN(n12480) );
  OR2_X1 U12624 ( .A1(n12724), .A2(n12725), .ZN(n12723) );
  AND2_X1 U12625 ( .A1(n12697), .A2(n12696), .ZN(n12725) );
  AND2_X1 U12626 ( .A1(n12694), .A2(n12726), .ZN(n12724) );
  OR2_X1 U12627 ( .A1(n12696), .A2(n12697), .ZN(n12726) );
  OR2_X1 U12628 ( .A1(n9297), .A2(n8971), .ZN(n12697) );
  OR2_X1 U12629 ( .A1(n12727), .A2(n12728), .ZN(n12696) );
  AND2_X1 U12630 ( .A1(n12693), .A2(n12692), .ZN(n12728) );
  AND2_X1 U12631 ( .A1(n12690), .A2(n12729), .ZN(n12727) );
  OR2_X1 U12632 ( .A1(n12692), .A2(n12693), .ZN(n12729) );
  OR2_X1 U12633 ( .A1(n8902), .A2(n8971), .ZN(n12693) );
  OR2_X1 U12634 ( .A1(n12730), .A2(n12731), .ZN(n12692) );
  AND2_X1 U12635 ( .A1(n12689), .A2(n12688), .ZN(n12731) );
  AND2_X1 U12636 ( .A1(n12686), .A2(n12732), .ZN(n12730) );
  OR2_X1 U12637 ( .A1(n12688), .A2(n12689), .ZN(n12732) );
  OR2_X1 U12638 ( .A1(n8906), .A2(n8971), .ZN(n12689) );
  OR2_X1 U12639 ( .A1(n12733), .A2(n12734), .ZN(n12688) );
  AND2_X1 U12640 ( .A1(n12685), .A2(n12684), .ZN(n12734) );
  AND2_X1 U12641 ( .A1(n12682), .A2(n12735), .ZN(n12733) );
  OR2_X1 U12642 ( .A1(n12684), .A2(n12685), .ZN(n12735) );
  OR2_X1 U12643 ( .A1(n8910), .A2(n8971), .ZN(n12685) );
  OR2_X1 U12644 ( .A1(n12736), .A2(n12737), .ZN(n12684) );
  AND2_X1 U12645 ( .A1(n12681), .A2(n12680), .ZN(n12737) );
  AND2_X1 U12646 ( .A1(n12678), .A2(n12738), .ZN(n12736) );
  OR2_X1 U12647 ( .A1(n12680), .A2(n12681), .ZN(n12738) );
  OR2_X1 U12648 ( .A1(n8914), .A2(n8971), .ZN(n12681) );
  OR2_X1 U12649 ( .A1(n12739), .A2(n12740), .ZN(n12680) );
  AND2_X1 U12650 ( .A1(n12677), .A2(n12676), .ZN(n12740) );
  AND2_X1 U12651 ( .A1(n12674), .A2(n12741), .ZN(n12739) );
  OR2_X1 U12652 ( .A1(n12676), .A2(n12677), .ZN(n12741) );
  OR2_X1 U12653 ( .A1(n8918), .A2(n8971), .ZN(n12677) );
  OR2_X1 U12654 ( .A1(n12742), .A2(n12743), .ZN(n12676) );
  AND2_X1 U12655 ( .A1(n12673), .A2(n12672), .ZN(n12743) );
  AND2_X1 U12656 ( .A1(n12670), .A2(n12744), .ZN(n12742) );
  OR2_X1 U12657 ( .A1(n12672), .A2(n12673), .ZN(n12744) );
  OR2_X1 U12658 ( .A1(n8922), .A2(n8971), .ZN(n12673) );
  OR2_X1 U12659 ( .A1(n12745), .A2(n12746), .ZN(n12672) );
  AND2_X1 U12660 ( .A1(n12669), .A2(n12668), .ZN(n12746) );
  AND2_X1 U12661 ( .A1(n12666), .A2(n12747), .ZN(n12745) );
  OR2_X1 U12662 ( .A1(n12668), .A2(n12669), .ZN(n12747) );
  OR2_X1 U12663 ( .A1(n8926), .A2(n8971), .ZN(n12669) );
  OR2_X1 U12664 ( .A1(n12748), .A2(n12749), .ZN(n12668) );
  AND2_X1 U12665 ( .A1(n12665), .A2(n12664), .ZN(n12749) );
  AND2_X1 U12666 ( .A1(n12662), .A2(n12750), .ZN(n12748) );
  OR2_X1 U12667 ( .A1(n12664), .A2(n12665), .ZN(n12750) );
  OR2_X1 U12668 ( .A1(n8930), .A2(n8971), .ZN(n12665) );
  OR2_X1 U12669 ( .A1(n12751), .A2(n12752), .ZN(n12664) );
  AND2_X1 U12670 ( .A1(n12661), .A2(n12660), .ZN(n12752) );
  AND2_X1 U12671 ( .A1(n12658), .A2(n12753), .ZN(n12751) );
  OR2_X1 U12672 ( .A1(n12660), .A2(n12661), .ZN(n12753) );
  OR2_X1 U12673 ( .A1(n8934), .A2(n8971), .ZN(n12661) );
  OR2_X1 U12674 ( .A1(n12754), .A2(n12755), .ZN(n12660) );
  AND2_X1 U12675 ( .A1(n12657), .A2(n12656), .ZN(n12755) );
  AND2_X1 U12676 ( .A1(n12654), .A2(n12756), .ZN(n12754) );
  OR2_X1 U12677 ( .A1(n12656), .A2(n12657), .ZN(n12756) );
  OR2_X1 U12678 ( .A1(n8938), .A2(n8971), .ZN(n12657) );
  OR2_X1 U12679 ( .A1(n12757), .A2(n12758), .ZN(n12656) );
  AND2_X1 U12680 ( .A1(n12653), .A2(n12652), .ZN(n12758) );
  AND2_X1 U12681 ( .A1(n12650), .A2(n12759), .ZN(n12757) );
  OR2_X1 U12682 ( .A1(n12652), .A2(n12653), .ZN(n12759) );
  OR2_X1 U12683 ( .A1(n8942), .A2(n8971), .ZN(n12653) );
  OR2_X1 U12684 ( .A1(n12760), .A2(n12761), .ZN(n12652) );
  AND2_X1 U12685 ( .A1(n12649), .A2(n12648), .ZN(n12761) );
  AND2_X1 U12686 ( .A1(n12646), .A2(n12762), .ZN(n12760) );
  OR2_X1 U12687 ( .A1(n12648), .A2(n12649), .ZN(n12762) );
  OR2_X1 U12688 ( .A1(n8946), .A2(n8971), .ZN(n12649) );
  OR2_X1 U12689 ( .A1(n12763), .A2(n12764), .ZN(n12648) );
  AND2_X1 U12690 ( .A1(n12645), .A2(n12644), .ZN(n12764) );
  AND2_X1 U12691 ( .A1(n12642), .A2(n12765), .ZN(n12763) );
  OR2_X1 U12692 ( .A1(n12644), .A2(n12645), .ZN(n12765) );
  OR2_X1 U12693 ( .A1(n8950), .A2(n8971), .ZN(n12645) );
  OR2_X1 U12694 ( .A1(n12766), .A2(n12767), .ZN(n12644) );
  AND2_X1 U12695 ( .A1(n12641), .A2(n12640), .ZN(n12767) );
  AND2_X1 U12696 ( .A1(n12638), .A2(n12768), .ZN(n12766) );
  OR2_X1 U12697 ( .A1(n12640), .A2(n12641), .ZN(n12768) );
  OR2_X1 U12698 ( .A1(n8954), .A2(n8971), .ZN(n12641) );
  OR2_X1 U12699 ( .A1(n12769), .A2(n12770), .ZN(n12640) );
  AND2_X1 U12700 ( .A1(n12637), .A2(n12636), .ZN(n12770) );
  AND2_X1 U12701 ( .A1(n12634), .A2(n12771), .ZN(n12769) );
  OR2_X1 U12702 ( .A1(n12636), .A2(n12637), .ZN(n12771) );
  OR2_X1 U12703 ( .A1(n8958), .A2(n8971), .ZN(n12637) );
  OR2_X1 U12704 ( .A1(n12772), .A2(n12773), .ZN(n12636) );
  AND2_X1 U12705 ( .A1(n12633), .A2(n12632), .ZN(n12773) );
  AND2_X1 U12706 ( .A1(n12630), .A2(n12774), .ZN(n12772) );
  OR2_X1 U12707 ( .A1(n12632), .A2(n12633), .ZN(n12774) );
  OR2_X1 U12708 ( .A1(n8962), .A2(n8971), .ZN(n12633) );
  OR2_X1 U12709 ( .A1(n12775), .A2(n12776), .ZN(n12632) );
  AND2_X1 U12710 ( .A1(n12629), .A2(n12628), .ZN(n12776) );
  AND2_X1 U12711 ( .A1(n12626), .A2(n12777), .ZN(n12775) );
  OR2_X1 U12712 ( .A1(n12628), .A2(n12629), .ZN(n12777) );
  OR2_X1 U12713 ( .A1(n8966), .A2(n8971), .ZN(n12629) );
  OR2_X1 U12714 ( .A1(n12778), .A2(n12779), .ZN(n12628) );
  AND2_X1 U12715 ( .A1(n8360), .A2(n12625), .ZN(n12779) );
  AND2_X1 U12716 ( .A1(n12623), .A2(n12780), .ZN(n12778) );
  OR2_X1 U12717 ( .A1(n12625), .A2(n8360), .ZN(n12780) );
  OR2_X1 U12718 ( .A1(n8970), .A2(n8971), .ZN(n8360) );
  OR2_X1 U12719 ( .A1(n12781), .A2(n12782), .ZN(n12625) );
  AND2_X1 U12720 ( .A1(n12622), .A2(n12621), .ZN(n12782) );
  AND2_X1 U12721 ( .A1(n12619), .A2(n12783), .ZN(n12781) );
  OR2_X1 U12722 ( .A1(n12621), .A2(n12622), .ZN(n12783) );
  OR2_X1 U12723 ( .A1(n8974), .A2(n8971), .ZN(n12622) );
  OR2_X1 U12724 ( .A1(n12784), .A2(n12785), .ZN(n12621) );
  AND2_X1 U12725 ( .A1(n12618), .A2(n12617), .ZN(n12785) );
  AND2_X1 U12726 ( .A1(n12615), .A2(n12786), .ZN(n12784) );
  OR2_X1 U12727 ( .A1(n12617), .A2(n12618), .ZN(n12786) );
  OR2_X1 U12728 ( .A1(n8978), .A2(n8971), .ZN(n12618) );
  OR2_X1 U12729 ( .A1(n12787), .A2(n12788), .ZN(n12617) );
  AND2_X1 U12730 ( .A1(n12614), .A2(n12613), .ZN(n12788) );
  AND2_X1 U12731 ( .A1(n12611), .A2(n12789), .ZN(n12787) );
  OR2_X1 U12732 ( .A1(n12613), .A2(n12614), .ZN(n12789) );
  OR2_X1 U12733 ( .A1(n8982), .A2(n8971), .ZN(n12614) );
  OR2_X1 U12734 ( .A1(n12790), .A2(n12791), .ZN(n12613) );
  AND2_X1 U12735 ( .A1(n12610), .A2(n12609), .ZN(n12791) );
  AND2_X1 U12736 ( .A1(n12607), .A2(n12792), .ZN(n12790) );
  OR2_X1 U12737 ( .A1(n12609), .A2(n12610), .ZN(n12792) );
  OR2_X1 U12738 ( .A1(n8986), .A2(n8971), .ZN(n12610) );
  OR2_X1 U12739 ( .A1(n12793), .A2(n12794), .ZN(n12609) );
  AND2_X1 U12740 ( .A1(n12606), .A2(n12605), .ZN(n12794) );
  AND2_X1 U12741 ( .A1(n12603), .A2(n12795), .ZN(n12793) );
  OR2_X1 U12742 ( .A1(n12605), .A2(n12606), .ZN(n12795) );
  OR2_X1 U12743 ( .A1(n8990), .A2(n8971), .ZN(n12606) );
  OR2_X1 U12744 ( .A1(n12796), .A2(n12797), .ZN(n12605) );
  AND2_X1 U12745 ( .A1(n12602), .A2(n12601), .ZN(n12797) );
  AND2_X1 U12746 ( .A1(n12599), .A2(n12798), .ZN(n12796) );
  OR2_X1 U12747 ( .A1(n12601), .A2(n12602), .ZN(n12798) );
  OR2_X1 U12748 ( .A1(n8994), .A2(n8971), .ZN(n12602) );
  OR2_X1 U12749 ( .A1(n12799), .A2(n12800), .ZN(n12601) );
  AND2_X1 U12750 ( .A1(n12598), .A2(n12597), .ZN(n12800) );
  AND2_X1 U12751 ( .A1(n12595), .A2(n12801), .ZN(n12799) );
  OR2_X1 U12752 ( .A1(n12597), .A2(n12598), .ZN(n12801) );
  OR2_X1 U12753 ( .A1(n8998), .A2(n8971), .ZN(n12598) );
  OR2_X1 U12754 ( .A1(n12802), .A2(n12803), .ZN(n12597) );
  AND2_X1 U12755 ( .A1(n12594), .A2(n12593), .ZN(n12803) );
  AND2_X1 U12756 ( .A1(n12591), .A2(n12804), .ZN(n12802) );
  OR2_X1 U12757 ( .A1(n12593), .A2(n12594), .ZN(n12804) );
  OR2_X1 U12758 ( .A1(n9002), .A2(n8971), .ZN(n12594) );
  OR2_X1 U12759 ( .A1(n12805), .A2(n12806), .ZN(n12593) );
  AND2_X1 U12760 ( .A1(n12590), .A2(n12589), .ZN(n12806) );
  AND2_X1 U12761 ( .A1(n12587), .A2(n12807), .ZN(n12805) );
  OR2_X1 U12762 ( .A1(n12589), .A2(n12590), .ZN(n12807) );
  OR2_X1 U12763 ( .A1(n9006), .A2(n8971), .ZN(n12590) );
  OR2_X1 U12764 ( .A1(n12808), .A2(n12809), .ZN(n12589) );
  AND2_X1 U12765 ( .A1(n12586), .A2(n12585), .ZN(n12809) );
  AND2_X1 U12766 ( .A1(n12583), .A2(n12810), .ZN(n12808) );
  OR2_X1 U12767 ( .A1(n12585), .A2(n12586), .ZN(n12810) );
  OR2_X1 U12768 ( .A1(n9010), .A2(n8971), .ZN(n12586) );
  OR2_X1 U12769 ( .A1(n12811), .A2(n12812), .ZN(n12585) );
  AND2_X1 U12770 ( .A1(n12580), .A2(n12581), .ZN(n12812) );
  AND2_X1 U12771 ( .A1(n12813), .A2(n12814), .ZN(n12811) );
  OR2_X1 U12772 ( .A1(n12581), .A2(n12580), .ZN(n12814) );
  OR2_X1 U12773 ( .A1(n9014), .A2(n8971), .ZN(n12580) );
  OR2_X1 U12774 ( .A1(n9984), .A2(n12815), .ZN(n12581) );
  OR2_X1 U12775 ( .A1(n8971), .A2(n8967), .ZN(n12815) );
  INV_X1 U12776 ( .A(n12582), .ZN(n12813) );
  OR2_X1 U12777 ( .A1(n12816), .A2(n12817), .ZN(n12582) );
  AND2_X1 U12778 ( .A1(b_17_), .A2(n12818), .ZN(n12817) );
  OR2_X1 U12779 ( .A1(n12819), .A2(n9989), .ZN(n12818) );
  AND2_X1 U12780 ( .A1(a_30_), .A2(n8963), .ZN(n12819) );
  AND2_X1 U12781 ( .A1(b_16_), .A2(n12820), .ZN(n12816) );
  OR2_X1 U12782 ( .A1(n12821), .A2(n8021), .ZN(n12820) );
  AND2_X1 U12783 ( .A1(a_31_), .A2(n8967), .ZN(n12821) );
  XOR2_X1 U12784 ( .A(n12822), .B(n12823), .Z(n12583) );
  XNOR2_X1 U12785 ( .A(n12824), .B(n12825), .ZN(n12822) );
  XOR2_X1 U12786 ( .A(n12826), .B(n12827), .Z(n12587) );
  XOR2_X1 U12787 ( .A(n12828), .B(n12829), .Z(n12827) );
  XOR2_X1 U12788 ( .A(n12830), .B(n12831), .Z(n12591) );
  XOR2_X1 U12789 ( .A(n12832), .B(n12833), .Z(n12831) );
  XOR2_X1 U12790 ( .A(n12834), .B(n12835), .Z(n12595) );
  XOR2_X1 U12791 ( .A(n12836), .B(n12837), .Z(n12835) );
  XOR2_X1 U12792 ( .A(n12838), .B(n12839), .Z(n12599) );
  XOR2_X1 U12793 ( .A(n12840), .B(n12841), .Z(n12839) );
  XOR2_X1 U12794 ( .A(n12842), .B(n12843), .Z(n12603) );
  XOR2_X1 U12795 ( .A(n12844), .B(n12845), .Z(n12843) );
  XOR2_X1 U12796 ( .A(n12846), .B(n12847), .Z(n12607) );
  XOR2_X1 U12797 ( .A(n12848), .B(n12849), .Z(n12847) );
  XOR2_X1 U12798 ( .A(n12850), .B(n12851), .Z(n12611) );
  XOR2_X1 U12799 ( .A(n12852), .B(n12853), .Z(n12851) );
  XOR2_X1 U12800 ( .A(n12854), .B(n12855), .Z(n12615) );
  XOR2_X1 U12801 ( .A(n12856), .B(n12857), .Z(n12855) );
  XOR2_X1 U12802 ( .A(n12858), .B(n12859), .Z(n12619) );
  XOR2_X1 U12803 ( .A(n12860), .B(n12861), .Z(n12859) );
  XOR2_X1 U12804 ( .A(n12862), .B(n12863), .Z(n12623) );
  XOR2_X1 U12805 ( .A(n12864), .B(n12865), .Z(n12863) );
  XOR2_X1 U12806 ( .A(n12866), .B(n12867), .Z(n12626) );
  XOR2_X1 U12807 ( .A(n12868), .B(n12869), .Z(n12867) );
  XOR2_X1 U12808 ( .A(n12870), .B(n12871), .Z(n12630) );
  XOR2_X1 U12809 ( .A(n12872), .B(n8393), .Z(n12871) );
  XOR2_X1 U12810 ( .A(n12873), .B(n12874), .Z(n12634) );
  XOR2_X1 U12811 ( .A(n12875), .B(n12876), .Z(n12874) );
  XOR2_X1 U12812 ( .A(n12877), .B(n12878), .Z(n12638) );
  XOR2_X1 U12813 ( .A(n12879), .B(n12880), .Z(n12878) );
  XOR2_X1 U12814 ( .A(n12881), .B(n12882), .Z(n12642) );
  XOR2_X1 U12815 ( .A(n12883), .B(n12884), .Z(n12882) );
  XOR2_X1 U12816 ( .A(n12885), .B(n12886), .Z(n12646) );
  XOR2_X1 U12817 ( .A(n12887), .B(n12888), .Z(n12886) );
  XOR2_X1 U12818 ( .A(n12889), .B(n12890), .Z(n12650) );
  XOR2_X1 U12819 ( .A(n12891), .B(n12892), .Z(n12890) );
  XOR2_X1 U12820 ( .A(n12893), .B(n12894), .Z(n12654) );
  XOR2_X1 U12821 ( .A(n12895), .B(n12896), .Z(n12894) );
  XOR2_X1 U12822 ( .A(n12897), .B(n12898), .Z(n12658) );
  XOR2_X1 U12823 ( .A(n12899), .B(n12900), .Z(n12898) );
  XOR2_X1 U12824 ( .A(n12901), .B(n12902), .Z(n12662) );
  XOR2_X1 U12825 ( .A(n12903), .B(n12904), .Z(n12902) );
  XOR2_X1 U12826 ( .A(n12905), .B(n12906), .Z(n12666) );
  XOR2_X1 U12827 ( .A(n12907), .B(n12908), .Z(n12906) );
  XOR2_X1 U12828 ( .A(n12909), .B(n12910), .Z(n12670) );
  XOR2_X1 U12829 ( .A(n12911), .B(n12912), .Z(n12910) );
  XOR2_X1 U12830 ( .A(n12913), .B(n12914), .Z(n12674) );
  XOR2_X1 U12831 ( .A(n12915), .B(n12916), .Z(n12914) );
  XOR2_X1 U12832 ( .A(n12917), .B(n12918), .Z(n12678) );
  XOR2_X1 U12833 ( .A(n12919), .B(n12920), .Z(n12918) );
  XOR2_X1 U12834 ( .A(n12921), .B(n12922), .Z(n12682) );
  XOR2_X1 U12835 ( .A(n12923), .B(n12924), .Z(n12922) );
  XOR2_X1 U12836 ( .A(n12925), .B(n12926), .Z(n12686) );
  XOR2_X1 U12837 ( .A(n12927), .B(n12928), .Z(n12926) );
  XOR2_X1 U12838 ( .A(n12929), .B(n12930), .Z(n12690) );
  XOR2_X1 U12839 ( .A(n12931), .B(n12932), .Z(n12930) );
  XOR2_X1 U12840 ( .A(n12933), .B(n12934), .Z(n12694) );
  XOR2_X1 U12841 ( .A(n12935), .B(n12936), .Z(n12934) );
  XNOR2_X1 U12842 ( .A(n12721), .B(n12937), .ZN(n12479) );
  XOR2_X1 U12843 ( .A(n12720), .B(n12719), .Z(n12937) );
  OR2_X1 U12844 ( .A1(n9297), .A2(n8967), .ZN(n12719) );
  OR2_X1 U12845 ( .A1(n12938), .A2(n12939), .ZN(n12720) );
  AND2_X1 U12846 ( .A1(n12936), .A2(n12935), .ZN(n12939) );
  AND2_X1 U12847 ( .A1(n12933), .A2(n12940), .ZN(n12938) );
  OR2_X1 U12848 ( .A1(n12936), .A2(n12935), .ZN(n12940) );
  OR2_X1 U12849 ( .A1(n12941), .A2(n12942), .ZN(n12935) );
  AND2_X1 U12850 ( .A1(n12932), .A2(n12931), .ZN(n12942) );
  AND2_X1 U12851 ( .A1(n12929), .A2(n12943), .ZN(n12941) );
  OR2_X1 U12852 ( .A1(n12932), .A2(n12931), .ZN(n12943) );
  OR2_X1 U12853 ( .A1(n12944), .A2(n12945), .ZN(n12931) );
  AND2_X1 U12854 ( .A1(n12928), .A2(n12927), .ZN(n12945) );
  AND2_X1 U12855 ( .A1(n12925), .A2(n12946), .ZN(n12944) );
  OR2_X1 U12856 ( .A1(n12928), .A2(n12927), .ZN(n12946) );
  OR2_X1 U12857 ( .A1(n12947), .A2(n12948), .ZN(n12927) );
  AND2_X1 U12858 ( .A1(n12924), .A2(n12923), .ZN(n12948) );
  AND2_X1 U12859 ( .A1(n12921), .A2(n12949), .ZN(n12947) );
  OR2_X1 U12860 ( .A1(n12924), .A2(n12923), .ZN(n12949) );
  OR2_X1 U12861 ( .A1(n12950), .A2(n12951), .ZN(n12923) );
  AND2_X1 U12862 ( .A1(n12920), .A2(n12919), .ZN(n12951) );
  AND2_X1 U12863 ( .A1(n12917), .A2(n12952), .ZN(n12950) );
  OR2_X1 U12864 ( .A1(n12920), .A2(n12919), .ZN(n12952) );
  OR2_X1 U12865 ( .A1(n12953), .A2(n12954), .ZN(n12919) );
  AND2_X1 U12866 ( .A1(n12916), .A2(n12915), .ZN(n12954) );
  AND2_X1 U12867 ( .A1(n12913), .A2(n12955), .ZN(n12953) );
  OR2_X1 U12868 ( .A1(n12916), .A2(n12915), .ZN(n12955) );
  OR2_X1 U12869 ( .A1(n12956), .A2(n12957), .ZN(n12915) );
  AND2_X1 U12870 ( .A1(n12912), .A2(n12911), .ZN(n12957) );
  AND2_X1 U12871 ( .A1(n12909), .A2(n12958), .ZN(n12956) );
  OR2_X1 U12872 ( .A1(n12912), .A2(n12911), .ZN(n12958) );
  OR2_X1 U12873 ( .A1(n12959), .A2(n12960), .ZN(n12911) );
  AND2_X1 U12874 ( .A1(n12908), .A2(n12907), .ZN(n12960) );
  AND2_X1 U12875 ( .A1(n12905), .A2(n12961), .ZN(n12959) );
  OR2_X1 U12876 ( .A1(n12908), .A2(n12907), .ZN(n12961) );
  OR2_X1 U12877 ( .A1(n12962), .A2(n12963), .ZN(n12907) );
  AND2_X1 U12878 ( .A1(n12904), .A2(n12903), .ZN(n12963) );
  AND2_X1 U12879 ( .A1(n12901), .A2(n12964), .ZN(n12962) );
  OR2_X1 U12880 ( .A1(n12904), .A2(n12903), .ZN(n12964) );
  OR2_X1 U12881 ( .A1(n12965), .A2(n12966), .ZN(n12903) );
  AND2_X1 U12882 ( .A1(n12900), .A2(n12899), .ZN(n12966) );
  AND2_X1 U12883 ( .A1(n12897), .A2(n12967), .ZN(n12965) );
  OR2_X1 U12884 ( .A1(n12900), .A2(n12899), .ZN(n12967) );
  OR2_X1 U12885 ( .A1(n12968), .A2(n12969), .ZN(n12899) );
  AND2_X1 U12886 ( .A1(n12896), .A2(n12895), .ZN(n12969) );
  AND2_X1 U12887 ( .A1(n12893), .A2(n12970), .ZN(n12968) );
  OR2_X1 U12888 ( .A1(n12896), .A2(n12895), .ZN(n12970) );
  OR2_X1 U12889 ( .A1(n12971), .A2(n12972), .ZN(n12895) );
  AND2_X1 U12890 ( .A1(n12892), .A2(n12891), .ZN(n12972) );
  AND2_X1 U12891 ( .A1(n12889), .A2(n12973), .ZN(n12971) );
  OR2_X1 U12892 ( .A1(n12892), .A2(n12891), .ZN(n12973) );
  OR2_X1 U12893 ( .A1(n12974), .A2(n12975), .ZN(n12891) );
  AND2_X1 U12894 ( .A1(n12888), .A2(n12887), .ZN(n12975) );
  AND2_X1 U12895 ( .A1(n12885), .A2(n12976), .ZN(n12974) );
  OR2_X1 U12896 ( .A1(n12888), .A2(n12887), .ZN(n12976) );
  OR2_X1 U12897 ( .A1(n12977), .A2(n12978), .ZN(n12887) );
  AND2_X1 U12898 ( .A1(n12884), .A2(n12883), .ZN(n12978) );
  AND2_X1 U12899 ( .A1(n12881), .A2(n12979), .ZN(n12977) );
  OR2_X1 U12900 ( .A1(n12884), .A2(n12883), .ZN(n12979) );
  OR2_X1 U12901 ( .A1(n12980), .A2(n12981), .ZN(n12883) );
  AND2_X1 U12902 ( .A1(n12880), .A2(n12879), .ZN(n12981) );
  AND2_X1 U12903 ( .A1(n12877), .A2(n12982), .ZN(n12980) );
  OR2_X1 U12904 ( .A1(n12880), .A2(n12879), .ZN(n12982) );
  OR2_X1 U12905 ( .A1(n12983), .A2(n12984), .ZN(n12879) );
  AND2_X1 U12906 ( .A1(n12876), .A2(n12875), .ZN(n12984) );
  AND2_X1 U12907 ( .A1(n12873), .A2(n12985), .ZN(n12983) );
  OR2_X1 U12908 ( .A1(n12876), .A2(n12875), .ZN(n12985) );
  OR2_X1 U12909 ( .A1(n12986), .A2(n12987), .ZN(n12875) );
  AND2_X1 U12910 ( .A1(n8393), .A2(n12872), .ZN(n12987) );
  AND2_X1 U12911 ( .A1(n12870), .A2(n12988), .ZN(n12986) );
  OR2_X1 U12912 ( .A1(n8393), .A2(n12872), .ZN(n12988) );
  OR2_X1 U12913 ( .A1(n12989), .A2(n12990), .ZN(n12872) );
  AND2_X1 U12914 ( .A1(n12869), .A2(n12868), .ZN(n12990) );
  AND2_X1 U12915 ( .A1(n12866), .A2(n12991), .ZN(n12989) );
  OR2_X1 U12916 ( .A1(n12869), .A2(n12868), .ZN(n12991) );
  OR2_X1 U12917 ( .A1(n12992), .A2(n12993), .ZN(n12868) );
  AND2_X1 U12918 ( .A1(n12865), .A2(n12864), .ZN(n12993) );
  AND2_X1 U12919 ( .A1(n12862), .A2(n12994), .ZN(n12992) );
  OR2_X1 U12920 ( .A1(n12865), .A2(n12864), .ZN(n12994) );
  OR2_X1 U12921 ( .A1(n12995), .A2(n12996), .ZN(n12864) );
  AND2_X1 U12922 ( .A1(n12861), .A2(n12860), .ZN(n12996) );
  AND2_X1 U12923 ( .A1(n12858), .A2(n12997), .ZN(n12995) );
  OR2_X1 U12924 ( .A1(n12861), .A2(n12860), .ZN(n12997) );
  OR2_X1 U12925 ( .A1(n12998), .A2(n12999), .ZN(n12860) );
  AND2_X1 U12926 ( .A1(n12857), .A2(n12856), .ZN(n12999) );
  AND2_X1 U12927 ( .A1(n12854), .A2(n13000), .ZN(n12998) );
  OR2_X1 U12928 ( .A1(n12857), .A2(n12856), .ZN(n13000) );
  OR2_X1 U12929 ( .A1(n13001), .A2(n13002), .ZN(n12856) );
  AND2_X1 U12930 ( .A1(n12853), .A2(n12852), .ZN(n13002) );
  AND2_X1 U12931 ( .A1(n12850), .A2(n13003), .ZN(n13001) );
  OR2_X1 U12932 ( .A1(n12853), .A2(n12852), .ZN(n13003) );
  OR2_X1 U12933 ( .A1(n13004), .A2(n13005), .ZN(n12852) );
  AND2_X1 U12934 ( .A1(n12849), .A2(n12848), .ZN(n13005) );
  AND2_X1 U12935 ( .A1(n12846), .A2(n13006), .ZN(n13004) );
  OR2_X1 U12936 ( .A1(n12849), .A2(n12848), .ZN(n13006) );
  OR2_X1 U12937 ( .A1(n13007), .A2(n13008), .ZN(n12848) );
  AND2_X1 U12938 ( .A1(n12845), .A2(n12844), .ZN(n13008) );
  AND2_X1 U12939 ( .A1(n12842), .A2(n13009), .ZN(n13007) );
  OR2_X1 U12940 ( .A1(n12845), .A2(n12844), .ZN(n13009) );
  OR2_X1 U12941 ( .A1(n13010), .A2(n13011), .ZN(n12844) );
  AND2_X1 U12942 ( .A1(n12841), .A2(n12840), .ZN(n13011) );
  AND2_X1 U12943 ( .A1(n12838), .A2(n13012), .ZN(n13010) );
  OR2_X1 U12944 ( .A1(n12841), .A2(n12840), .ZN(n13012) );
  OR2_X1 U12945 ( .A1(n13013), .A2(n13014), .ZN(n12840) );
  AND2_X1 U12946 ( .A1(n12837), .A2(n12836), .ZN(n13014) );
  AND2_X1 U12947 ( .A1(n12834), .A2(n13015), .ZN(n13013) );
  OR2_X1 U12948 ( .A1(n12837), .A2(n12836), .ZN(n13015) );
  OR2_X1 U12949 ( .A1(n13016), .A2(n13017), .ZN(n12836) );
  AND2_X1 U12950 ( .A1(n12833), .A2(n12832), .ZN(n13017) );
  AND2_X1 U12951 ( .A1(n12830), .A2(n13018), .ZN(n13016) );
  OR2_X1 U12952 ( .A1(n12833), .A2(n12832), .ZN(n13018) );
  OR2_X1 U12953 ( .A1(n13019), .A2(n13020), .ZN(n12832) );
  AND2_X1 U12954 ( .A1(n12829), .A2(n12828), .ZN(n13020) );
  AND2_X1 U12955 ( .A1(n12826), .A2(n13021), .ZN(n13019) );
  OR2_X1 U12956 ( .A1(n12829), .A2(n12828), .ZN(n13021) );
  OR2_X1 U12957 ( .A1(n13022), .A2(n13023), .ZN(n12828) );
  AND2_X1 U12958 ( .A1(n12823), .A2(n12824), .ZN(n13023) );
  AND2_X1 U12959 ( .A1(n13024), .A2(n13025), .ZN(n13022) );
  OR2_X1 U12960 ( .A1(n12823), .A2(n12824), .ZN(n13025) );
  OR2_X1 U12961 ( .A1(n9984), .A2(n13026), .ZN(n12824) );
  OR2_X1 U12962 ( .A1(n8967), .A2(n8963), .ZN(n13026) );
  OR2_X1 U12963 ( .A1(n9014), .A2(n8967), .ZN(n12823) );
  INV_X1 U12964 ( .A(n12825), .ZN(n13024) );
  OR2_X1 U12965 ( .A1(n13027), .A2(n13028), .ZN(n12825) );
  AND2_X1 U12966 ( .A1(b_16_), .A2(n13029), .ZN(n13028) );
  OR2_X1 U12967 ( .A1(n13030), .A2(n9989), .ZN(n13029) );
  AND2_X1 U12968 ( .A1(a_30_), .A2(n8959), .ZN(n13030) );
  AND2_X1 U12969 ( .A1(b_15_), .A2(n13031), .ZN(n13027) );
  OR2_X1 U12970 ( .A1(n13032), .A2(n8021), .ZN(n13031) );
  AND2_X1 U12971 ( .A1(a_31_), .A2(n8963), .ZN(n13032) );
  OR2_X1 U12972 ( .A1(n9010), .A2(n8967), .ZN(n12829) );
  XOR2_X1 U12973 ( .A(n13033), .B(n13034), .Z(n12826) );
  XNOR2_X1 U12974 ( .A(n13035), .B(n13036), .ZN(n13033) );
  OR2_X1 U12975 ( .A1(n9006), .A2(n8967), .ZN(n12833) );
  XOR2_X1 U12976 ( .A(n13037), .B(n13038), .Z(n12830) );
  XOR2_X1 U12977 ( .A(n13039), .B(n13040), .Z(n13038) );
  OR2_X1 U12978 ( .A1(n9002), .A2(n8967), .ZN(n12837) );
  XOR2_X1 U12979 ( .A(n13041), .B(n13042), .Z(n12834) );
  XOR2_X1 U12980 ( .A(n13043), .B(n13044), .Z(n13042) );
  OR2_X1 U12981 ( .A1(n8998), .A2(n8967), .ZN(n12841) );
  XOR2_X1 U12982 ( .A(n13045), .B(n13046), .Z(n12838) );
  XOR2_X1 U12983 ( .A(n13047), .B(n13048), .Z(n13046) );
  OR2_X1 U12984 ( .A1(n8994), .A2(n8967), .ZN(n12845) );
  XOR2_X1 U12985 ( .A(n13049), .B(n13050), .Z(n12842) );
  XOR2_X1 U12986 ( .A(n13051), .B(n13052), .Z(n13050) );
  OR2_X1 U12987 ( .A1(n8990), .A2(n8967), .ZN(n12849) );
  XOR2_X1 U12988 ( .A(n13053), .B(n13054), .Z(n12846) );
  XOR2_X1 U12989 ( .A(n13055), .B(n13056), .Z(n13054) );
  OR2_X1 U12990 ( .A1(n8986), .A2(n8967), .ZN(n12853) );
  XOR2_X1 U12991 ( .A(n13057), .B(n13058), .Z(n12850) );
  XOR2_X1 U12992 ( .A(n13059), .B(n13060), .Z(n13058) );
  OR2_X1 U12993 ( .A1(n8982), .A2(n8967), .ZN(n12857) );
  XOR2_X1 U12994 ( .A(n13061), .B(n13062), .Z(n12854) );
  XOR2_X1 U12995 ( .A(n13063), .B(n13064), .Z(n13062) );
  OR2_X1 U12996 ( .A1(n8978), .A2(n8967), .ZN(n12861) );
  XOR2_X1 U12997 ( .A(n13065), .B(n13066), .Z(n12858) );
  XOR2_X1 U12998 ( .A(n13067), .B(n13068), .Z(n13066) );
  OR2_X1 U12999 ( .A1(n8974), .A2(n8967), .ZN(n12865) );
  XOR2_X1 U13000 ( .A(n13069), .B(n13070), .Z(n12862) );
  XOR2_X1 U13001 ( .A(n13071), .B(n13072), .Z(n13070) );
  OR2_X1 U13002 ( .A1(n8970), .A2(n8967), .ZN(n12869) );
  XOR2_X1 U13003 ( .A(n13073), .B(n13074), .Z(n12866) );
  XOR2_X1 U13004 ( .A(n13075), .B(n13076), .Z(n13074) );
  OR2_X1 U13005 ( .A1(n8966), .A2(n8967), .ZN(n8393) );
  XOR2_X1 U13006 ( .A(n13077), .B(n13078), .Z(n12870) );
  XOR2_X1 U13007 ( .A(n13079), .B(n13080), .Z(n13078) );
  OR2_X1 U13008 ( .A1(n8962), .A2(n8967), .ZN(n12876) );
  XOR2_X1 U13009 ( .A(n13081), .B(n13082), .Z(n12873) );
  XOR2_X1 U13010 ( .A(n13083), .B(n13084), .Z(n13082) );
  OR2_X1 U13011 ( .A1(n8958), .A2(n8967), .ZN(n12880) );
  XOR2_X1 U13012 ( .A(n13085), .B(n13086), .Z(n12877) );
  XOR2_X1 U13013 ( .A(n13087), .B(n8422), .Z(n13086) );
  OR2_X1 U13014 ( .A1(n8954), .A2(n8967), .ZN(n12884) );
  XOR2_X1 U13015 ( .A(n13088), .B(n13089), .Z(n12881) );
  XOR2_X1 U13016 ( .A(n13090), .B(n13091), .Z(n13089) );
  OR2_X1 U13017 ( .A1(n8950), .A2(n8967), .ZN(n12888) );
  XOR2_X1 U13018 ( .A(n13092), .B(n13093), .Z(n12885) );
  XOR2_X1 U13019 ( .A(n13094), .B(n13095), .Z(n13093) );
  OR2_X1 U13020 ( .A1(n8946), .A2(n8967), .ZN(n12892) );
  XOR2_X1 U13021 ( .A(n13096), .B(n13097), .Z(n12889) );
  XOR2_X1 U13022 ( .A(n13098), .B(n13099), .Z(n13097) );
  OR2_X1 U13023 ( .A1(n8942), .A2(n8967), .ZN(n12896) );
  XOR2_X1 U13024 ( .A(n13100), .B(n13101), .Z(n12893) );
  XOR2_X1 U13025 ( .A(n13102), .B(n13103), .Z(n13101) );
  OR2_X1 U13026 ( .A1(n8938), .A2(n8967), .ZN(n12900) );
  XOR2_X1 U13027 ( .A(n13104), .B(n13105), .Z(n12897) );
  XOR2_X1 U13028 ( .A(n13106), .B(n13107), .Z(n13105) );
  OR2_X1 U13029 ( .A1(n8934), .A2(n8967), .ZN(n12904) );
  XOR2_X1 U13030 ( .A(n13108), .B(n13109), .Z(n12901) );
  XOR2_X1 U13031 ( .A(n13110), .B(n13111), .Z(n13109) );
  OR2_X1 U13032 ( .A1(n8930), .A2(n8967), .ZN(n12908) );
  XOR2_X1 U13033 ( .A(n13112), .B(n13113), .Z(n12905) );
  XOR2_X1 U13034 ( .A(n13114), .B(n13115), .Z(n13113) );
  OR2_X1 U13035 ( .A1(n8926), .A2(n8967), .ZN(n12912) );
  XOR2_X1 U13036 ( .A(n13116), .B(n13117), .Z(n12909) );
  XOR2_X1 U13037 ( .A(n13118), .B(n13119), .Z(n13117) );
  OR2_X1 U13038 ( .A1(n8922), .A2(n8967), .ZN(n12916) );
  XOR2_X1 U13039 ( .A(n13120), .B(n13121), .Z(n12913) );
  XOR2_X1 U13040 ( .A(n13122), .B(n13123), .Z(n13121) );
  OR2_X1 U13041 ( .A1(n8918), .A2(n8967), .ZN(n12920) );
  XOR2_X1 U13042 ( .A(n13124), .B(n13125), .Z(n12917) );
  XOR2_X1 U13043 ( .A(n13126), .B(n13127), .Z(n13125) );
  OR2_X1 U13044 ( .A1(n8914), .A2(n8967), .ZN(n12924) );
  XOR2_X1 U13045 ( .A(n13128), .B(n13129), .Z(n12921) );
  XOR2_X1 U13046 ( .A(n13130), .B(n13131), .Z(n13129) );
  OR2_X1 U13047 ( .A1(n8910), .A2(n8967), .ZN(n12928) );
  XOR2_X1 U13048 ( .A(n13132), .B(n13133), .Z(n12925) );
  XOR2_X1 U13049 ( .A(n13134), .B(n13135), .Z(n13133) );
  OR2_X1 U13050 ( .A1(n8906), .A2(n8967), .ZN(n12932) );
  XOR2_X1 U13051 ( .A(n13136), .B(n13137), .Z(n12929) );
  XOR2_X1 U13052 ( .A(n13138), .B(n13139), .Z(n13137) );
  OR2_X1 U13053 ( .A1(n8902), .A2(n8967), .ZN(n12936) );
  XOR2_X1 U13054 ( .A(n13140), .B(n13141), .Z(n12933) );
  XOR2_X1 U13055 ( .A(n13142), .B(n13143), .Z(n13141) );
  XOR2_X1 U13056 ( .A(n12704), .B(n13144), .Z(n12721) );
  XOR2_X1 U13057 ( .A(n12703), .B(n12702), .Z(n13144) );
  OR2_X1 U13058 ( .A1(n8902), .A2(n8963), .ZN(n12702) );
  OR2_X1 U13059 ( .A1(n13145), .A2(n13146), .ZN(n12703) );
  AND2_X1 U13060 ( .A1(n13143), .A2(n13142), .ZN(n13146) );
  AND2_X1 U13061 ( .A1(n13140), .A2(n13147), .ZN(n13145) );
  OR2_X1 U13062 ( .A1(n13143), .A2(n13142), .ZN(n13147) );
  OR2_X1 U13063 ( .A1(n13148), .A2(n13149), .ZN(n13142) );
  AND2_X1 U13064 ( .A1(n13139), .A2(n13138), .ZN(n13149) );
  AND2_X1 U13065 ( .A1(n13136), .A2(n13150), .ZN(n13148) );
  OR2_X1 U13066 ( .A1(n13139), .A2(n13138), .ZN(n13150) );
  OR2_X1 U13067 ( .A1(n13151), .A2(n13152), .ZN(n13138) );
  AND2_X1 U13068 ( .A1(n13135), .A2(n13134), .ZN(n13152) );
  AND2_X1 U13069 ( .A1(n13132), .A2(n13153), .ZN(n13151) );
  OR2_X1 U13070 ( .A1(n13135), .A2(n13134), .ZN(n13153) );
  OR2_X1 U13071 ( .A1(n13154), .A2(n13155), .ZN(n13134) );
  AND2_X1 U13072 ( .A1(n13131), .A2(n13130), .ZN(n13155) );
  AND2_X1 U13073 ( .A1(n13128), .A2(n13156), .ZN(n13154) );
  OR2_X1 U13074 ( .A1(n13131), .A2(n13130), .ZN(n13156) );
  OR2_X1 U13075 ( .A1(n13157), .A2(n13158), .ZN(n13130) );
  AND2_X1 U13076 ( .A1(n13127), .A2(n13126), .ZN(n13158) );
  AND2_X1 U13077 ( .A1(n13124), .A2(n13159), .ZN(n13157) );
  OR2_X1 U13078 ( .A1(n13127), .A2(n13126), .ZN(n13159) );
  OR2_X1 U13079 ( .A1(n13160), .A2(n13161), .ZN(n13126) );
  AND2_X1 U13080 ( .A1(n13123), .A2(n13122), .ZN(n13161) );
  AND2_X1 U13081 ( .A1(n13120), .A2(n13162), .ZN(n13160) );
  OR2_X1 U13082 ( .A1(n13123), .A2(n13122), .ZN(n13162) );
  OR2_X1 U13083 ( .A1(n13163), .A2(n13164), .ZN(n13122) );
  AND2_X1 U13084 ( .A1(n13119), .A2(n13118), .ZN(n13164) );
  AND2_X1 U13085 ( .A1(n13116), .A2(n13165), .ZN(n13163) );
  OR2_X1 U13086 ( .A1(n13119), .A2(n13118), .ZN(n13165) );
  OR2_X1 U13087 ( .A1(n13166), .A2(n13167), .ZN(n13118) );
  AND2_X1 U13088 ( .A1(n13115), .A2(n13114), .ZN(n13167) );
  AND2_X1 U13089 ( .A1(n13112), .A2(n13168), .ZN(n13166) );
  OR2_X1 U13090 ( .A1(n13115), .A2(n13114), .ZN(n13168) );
  OR2_X1 U13091 ( .A1(n13169), .A2(n13170), .ZN(n13114) );
  AND2_X1 U13092 ( .A1(n13111), .A2(n13110), .ZN(n13170) );
  AND2_X1 U13093 ( .A1(n13108), .A2(n13171), .ZN(n13169) );
  OR2_X1 U13094 ( .A1(n13111), .A2(n13110), .ZN(n13171) );
  OR2_X1 U13095 ( .A1(n13172), .A2(n13173), .ZN(n13110) );
  AND2_X1 U13096 ( .A1(n13107), .A2(n13106), .ZN(n13173) );
  AND2_X1 U13097 ( .A1(n13104), .A2(n13174), .ZN(n13172) );
  OR2_X1 U13098 ( .A1(n13107), .A2(n13106), .ZN(n13174) );
  OR2_X1 U13099 ( .A1(n13175), .A2(n13176), .ZN(n13106) );
  AND2_X1 U13100 ( .A1(n13103), .A2(n13102), .ZN(n13176) );
  AND2_X1 U13101 ( .A1(n13100), .A2(n13177), .ZN(n13175) );
  OR2_X1 U13102 ( .A1(n13103), .A2(n13102), .ZN(n13177) );
  OR2_X1 U13103 ( .A1(n13178), .A2(n13179), .ZN(n13102) );
  AND2_X1 U13104 ( .A1(n13096), .A2(n13099), .ZN(n13179) );
  AND2_X1 U13105 ( .A1(n13180), .A2(n13098), .ZN(n13178) );
  OR2_X1 U13106 ( .A1(n13181), .A2(n13182), .ZN(n13098) );
  AND2_X1 U13107 ( .A1(n13095), .A2(n13094), .ZN(n13182) );
  AND2_X1 U13108 ( .A1(n13092), .A2(n13183), .ZN(n13181) );
  OR2_X1 U13109 ( .A1(n13095), .A2(n13094), .ZN(n13183) );
  OR2_X1 U13110 ( .A1(n13184), .A2(n13185), .ZN(n13094) );
  AND2_X1 U13111 ( .A1(n13088), .A2(n13091), .ZN(n13185) );
  AND2_X1 U13112 ( .A1(n13186), .A2(n13090), .ZN(n13184) );
  OR2_X1 U13113 ( .A1(n13187), .A2(n13188), .ZN(n13090) );
  AND2_X1 U13114 ( .A1(n13085), .A2(n8422), .ZN(n13188) );
  AND2_X1 U13115 ( .A1(n13189), .A2(n13087), .ZN(n13187) );
  OR2_X1 U13116 ( .A1(n13190), .A2(n13191), .ZN(n13087) );
  AND2_X1 U13117 ( .A1(n13081), .A2(n13084), .ZN(n13191) );
  AND2_X1 U13118 ( .A1(n13192), .A2(n13083), .ZN(n13190) );
  OR2_X1 U13119 ( .A1(n13193), .A2(n13194), .ZN(n13083) );
  AND2_X1 U13120 ( .A1(n13077), .A2(n13080), .ZN(n13194) );
  AND2_X1 U13121 ( .A1(n13195), .A2(n13079), .ZN(n13193) );
  OR2_X1 U13122 ( .A1(n13196), .A2(n13197), .ZN(n13079) );
  AND2_X1 U13123 ( .A1(n13073), .A2(n13076), .ZN(n13197) );
  AND2_X1 U13124 ( .A1(n13198), .A2(n13075), .ZN(n13196) );
  OR2_X1 U13125 ( .A1(n13199), .A2(n13200), .ZN(n13075) );
  AND2_X1 U13126 ( .A1(n13069), .A2(n13072), .ZN(n13200) );
  AND2_X1 U13127 ( .A1(n13201), .A2(n13071), .ZN(n13199) );
  OR2_X1 U13128 ( .A1(n13202), .A2(n13203), .ZN(n13071) );
  AND2_X1 U13129 ( .A1(n13065), .A2(n13068), .ZN(n13203) );
  AND2_X1 U13130 ( .A1(n13204), .A2(n13067), .ZN(n13202) );
  OR2_X1 U13131 ( .A1(n13205), .A2(n13206), .ZN(n13067) );
  AND2_X1 U13132 ( .A1(n13061), .A2(n13064), .ZN(n13206) );
  AND2_X1 U13133 ( .A1(n13207), .A2(n13063), .ZN(n13205) );
  OR2_X1 U13134 ( .A1(n13208), .A2(n13209), .ZN(n13063) );
  AND2_X1 U13135 ( .A1(n13057), .A2(n13060), .ZN(n13209) );
  AND2_X1 U13136 ( .A1(n13210), .A2(n13059), .ZN(n13208) );
  OR2_X1 U13137 ( .A1(n13211), .A2(n13212), .ZN(n13059) );
  AND2_X1 U13138 ( .A1(n13053), .A2(n13056), .ZN(n13212) );
  AND2_X1 U13139 ( .A1(n13213), .A2(n13055), .ZN(n13211) );
  OR2_X1 U13140 ( .A1(n13214), .A2(n13215), .ZN(n13055) );
  AND2_X1 U13141 ( .A1(n13049), .A2(n13052), .ZN(n13215) );
  AND2_X1 U13142 ( .A1(n13216), .A2(n13051), .ZN(n13214) );
  OR2_X1 U13143 ( .A1(n13217), .A2(n13218), .ZN(n13051) );
  AND2_X1 U13144 ( .A1(n13045), .A2(n13048), .ZN(n13218) );
  AND2_X1 U13145 ( .A1(n13219), .A2(n13047), .ZN(n13217) );
  OR2_X1 U13146 ( .A1(n13220), .A2(n13221), .ZN(n13047) );
  AND2_X1 U13147 ( .A1(n13041), .A2(n13044), .ZN(n13221) );
  AND2_X1 U13148 ( .A1(n13222), .A2(n13043), .ZN(n13220) );
  OR2_X1 U13149 ( .A1(n13223), .A2(n13224), .ZN(n13043) );
  AND2_X1 U13150 ( .A1(n13037), .A2(n13040), .ZN(n13224) );
  AND2_X1 U13151 ( .A1(n13225), .A2(n13039), .ZN(n13223) );
  OR2_X1 U13152 ( .A1(n13226), .A2(n13227), .ZN(n13039) );
  AND2_X1 U13153 ( .A1(n13034), .A2(n13035), .ZN(n13227) );
  AND2_X1 U13154 ( .A1(n13228), .A2(n13229), .ZN(n13226) );
  OR2_X1 U13155 ( .A1(n13034), .A2(n13035), .ZN(n13229) );
  OR2_X1 U13156 ( .A1(n9984), .A2(n13230), .ZN(n13035) );
  OR2_X1 U13157 ( .A1(n8963), .A2(n8959), .ZN(n13230) );
  OR2_X1 U13158 ( .A1(n9014), .A2(n8963), .ZN(n13034) );
  INV_X1 U13159 ( .A(n13036), .ZN(n13228) );
  OR2_X1 U13160 ( .A1(n13231), .A2(n13232), .ZN(n13036) );
  AND2_X1 U13161 ( .A1(b_15_), .A2(n13233), .ZN(n13232) );
  OR2_X1 U13162 ( .A1(n13234), .A2(n9989), .ZN(n13233) );
  AND2_X1 U13163 ( .A1(a_30_), .A2(n8955), .ZN(n13234) );
  AND2_X1 U13164 ( .A1(b_14_), .A2(n13235), .ZN(n13231) );
  OR2_X1 U13165 ( .A1(n13236), .A2(n8021), .ZN(n13235) );
  AND2_X1 U13166 ( .A1(a_31_), .A2(n8959), .ZN(n13236) );
  OR2_X1 U13167 ( .A1(n13037), .A2(n13040), .ZN(n13225) );
  OR2_X1 U13168 ( .A1(n9010), .A2(n8963), .ZN(n13040) );
  XOR2_X1 U13169 ( .A(n13237), .B(n13238), .Z(n13037) );
  XNOR2_X1 U13170 ( .A(n13239), .B(n13240), .ZN(n13237) );
  OR2_X1 U13171 ( .A1(n13041), .A2(n13044), .ZN(n13222) );
  OR2_X1 U13172 ( .A1(n9006), .A2(n8963), .ZN(n13044) );
  XOR2_X1 U13173 ( .A(n13241), .B(n13242), .Z(n13041) );
  XOR2_X1 U13174 ( .A(n13243), .B(n13244), .Z(n13242) );
  OR2_X1 U13175 ( .A1(n13045), .A2(n13048), .ZN(n13219) );
  OR2_X1 U13176 ( .A1(n9002), .A2(n8963), .ZN(n13048) );
  XOR2_X1 U13177 ( .A(n13245), .B(n13246), .Z(n13045) );
  XOR2_X1 U13178 ( .A(n13247), .B(n13248), .Z(n13246) );
  OR2_X1 U13179 ( .A1(n13049), .A2(n13052), .ZN(n13216) );
  OR2_X1 U13180 ( .A1(n8998), .A2(n8963), .ZN(n13052) );
  XOR2_X1 U13181 ( .A(n13249), .B(n13250), .Z(n13049) );
  XOR2_X1 U13182 ( .A(n13251), .B(n13252), .Z(n13250) );
  OR2_X1 U13183 ( .A1(n13053), .A2(n13056), .ZN(n13213) );
  OR2_X1 U13184 ( .A1(n8994), .A2(n8963), .ZN(n13056) );
  XOR2_X1 U13185 ( .A(n13253), .B(n13254), .Z(n13053) );
  XOR2_X1 U13186 ( .A(n13255), .B(n13256), .Z(n13254) );
  OR2_X1 U13187 ( .A1(n13057), .A2(n13060), .ZN(n13210) );
  OR2_X1 U13188 ( .A1(n8990), .A2(n8963), .ZN(n13060) );
  XOR2_X1 U13189 ( .A(n13257), .B(n13258), .Z(n13057) );
  XOR2_X1 U13190 ( .A(n13259), .B(n13260), .Z(n13258) );
  OR2_X1 U13191 ( .A1(n13061), .A2(n13064), .ZN(n13207) );
  OR2_X1 U13192 ( .A1(n8986), .A2(n8963), .ZN(n13064) );
  XOR2_X1 U13193 ( .A(n13261), .B(n13262), .Z(n13061) );
  XOR2_X1 U13194 ( .A(n13263), .B(n13264), .Z(n13262) );
  OR2_X1 U13195 ( .A1(n13065), .A2(n13068), .ZN(n13204) );
  OR2_X1 U13196 ( .A1(n8982), .A2(n8963), .ZN(n13068) );
  XOR2_X1 U13197 ( .A(n13265), .B(n13266), .Z(n13065) );
  XOR2_X1 U13198 ( .A(n13267), .B(n13268), .Z(n13266) );
  OR2_X1 U13199 ( .A1(n13069), .A2(n13072), .ZN(n13201) );
  OR2_X1 U13200 ( .A1(n8978), .A2(n8963), .ZN(n13072) );
  XOR2_X1 U13201 ( .A(n13269), .B(n13270), .Z(n13069) );
  XOR2_X1 U13202 ( .A(n13271), .B(n13272), .Z(n13270) );
  OR2_X1 U13203 ( .A1(n13073), .A2(n13076), .ZN(n13198) );
  OR2_X1 U13204 ( .A1(n8974), .A2(n8963), .ZN(n13076) );
  XOR2_X1 U13205 ( .A(n13273), .B(n13274), .Z(n13073) );
  XOR2_X1 U13206 ( .A(n13275), .B(n13276), .Z(n13274) );
  OR2_X1 U13207 ( .A1(n13077), .A2(n13080), .ZN(n13195) );
  OR2_X1 U13208 ( .A1(n8970), .A2(n8963), .ZN(n13080) );
  XOR2_X1 U13209 ( .A(n13277), .B(n13278), .Z(n13077) );
  XOR2_X1 U13210 ( .A(n13279), .B(n13280), .Z(n13278) );
  OR2_X1 U13211 ( .A1(n13081), .A2(n13084), .ZN(n13192) );
  OR2_X1 U13212 ( .A1(n8966), .A2(n8963), .ZN(n13084) );
  XOR2_X1 U13213 ( .A(n13281), .B(n13282), .Z(n13081) );
  XOR2_X1 U13214 ( .A(n13283), .B(n13284), .Z(n13282) );
  OR2_X1 U13215 ( .A1(n13085), .A2(n8422), .ZN(n13189) );
  OR2_X1 U13216 ( .A1(n8962), .A2(n8963), .ZN(n8422) );
  XOR2_X1 U13217 ( .A(n13285), .B(n13286), .Z(n13085) );
  XOR2_X1 U13218 ( .A(n13287), .B(n13288), .Z(n13286) );
  OR2_X1 U13219 ( .A1(n13088), .A2(n13091), .ZN(n13186) );
  OR2_X1 U13220 ( .A1(n8958), .A2(n8963), .ZN(n13091) );
  XOR2_X1 U13221 ( .A(n13289), .B(n13290), .Z(n13088) );
  XOR2_X1 U13222 ( .A(n13291), .B(n13292), .Z(n13290) );
  OR2_X1 U13223 ( .A1(n8954), .A2(n8963), .ZN(n13095) );
  XOR2_X1 U13224 ( .A(n13293), .B(n13294), .Z(n13092) );
  XOR2_X1 U13225 ( .A(n13295), .B(n8451), .Z(n13294) );
  OR2_X1 U13226 ( .A1(n13096), .A2(n13099), .ZN(n13180) );
  OR2_X1 U13227 ( .A1(n8950), .A2(n8963), .ZN(n13099) );
  XOR2_X1 U13228 ( .A(n13296), .B(n13297), .Z(n13096) );
  XOR2_X1 U13229 ( .A(n13298), .B(n13299), .Z(n13297) );
  OR2_X1 U13230 ( .A1(n8946), .A2(n8963), .ZN(n13103) );
  XOR2_X1 U13231 ( .A(n13300), .B(n13301), .Z(n13100) );
  XOR2_X1 U13232 ( .A(n13302), .B(n13303), .Z(n13301) );
  OR2_X1 U13233 ( .A1(n8942), .A2(n8963), .ZN(n13107) );
  XOR2_X1 U13234 ( .A(n13304), .B(n13305), .Z(n13104) );
  XOR2_X1 U13235 ( .A(n13306), .B(n13307), .Z(n13305) );
  OR2_X1 U13236 ( .A1(n8938), .A2(n8963), .ZN(n13111) );
  XOR2_X1 U13237 ( .A(n13308), .B(n13309), .Z(n13108) );
  XOR2_X1 U13238 ( .A(n13310), .B(n13311), .Z(n13309) );
  OR2_X1 U13239 ( .A1(n8934), .A2(n8963), .ZN(n13115) );
  XOR2_X1 U13240 ( .A(n13312), .B(n13313), .Z(n13112) );
  XOR2_X1 U13241 ( .A(n13314), .B(n13315), .Z(n13313) );
  OR2_X1 U13242 ( .A1(n8930), .A2(n8963), .ZN(n13119) );
  XOR2_X1 U13243 ( .A(n13316), .B(n13317), .Z(n13116) );
  XOR2_X1 U13244 ( .A(n13318), .B(n13319), .Z(n13317) );
  OR2_X1 U13245 ( .A1(n8926), .A2(n8963), .ZN(n13123) );
  XOR2_X1 U13246 ( .A(n13320), .B(n13321), .Z(n13120) );
  XOR2_X1 U13247 ( .A(n13322), .B(n13323), .Z(n13321) );
  OR2_X1 U13248 ( .A1(n8922), .A2(n8963), .ZN(n13127) );
  XOR2_X1 U13249 ( .A(n13324), .B(n13325), .Z(n13124) );
  XOR2_X1 U13250 ( .A(n13326), .B(n13327), .Z(n13325) );
  OR2_X1 U13251 ( .A1(n8918), .A2(n8963), .ZN(n13131) );
  XOR2_X1 U13252 ( .A(n13328), .B(n13329), .Z(n13128) );
  XOR2_X1 U13253 ( .A(n13330), .B(n13331), .Z(n13329) );
  OR2_X1 U13254 ( .A1(n8914), .A2(n8963), .ZN(n13135) );
  XOR2_X1 U13255 ( .A(n13332), .B(n13333), .Z(n13132) );
  XOR2_X1 U13256 ( .A(n13334), .B(n13335), .Z(n13333) );
  OR2_X1 U13257 ( .A1(n8910), .A2(n8963), .ZN(n13139) );
  XOR2_X1 U13258 ( .A(n13336), .B(n13337), .Z(n13136) );
  XOR2_X1 U13259 ( .A(n13338), .B(n13339), .Z(n13337) );
  OR2_X1 U13260 ( .A1(n8906), .A2(n8963), .ZN(n13143) );
  XOR2_X1 U13261 ( .A(n13340), .B(n13341), .Z(n13140) );
  XOR2_X1 U13262 ( .A(n13342), .B(n13343), .Z(n13341) );
  XOR2_X1 U13263 ( .A(n12711), .B(n13344), .Z(n12704) );
  XOR2_X1 U13264 ( .A(n12710), .B(n12709), .Z(n13344) );
  OR2_X1 U13265 ( .A1(n8906), .A2(n8959), .ZN(n12709) );
  OR2_X1 U13266 ( .A1(n13345), .A2(n13346), .ZN(n12710) );
  AND2_X1 U13267 ( .A1(n13343), .A2(n13342), .ZN(n13346) );
  AND2_X1 U13268 ( .A1(n13340), .A2(n13347), .ZN(n13345) );
  OR2_X1 U13269 ( .A1(n13342), .A2(n13343), .ZN(n13347) );
  OR2_X1 U13270 ( .A1(n8910), .A2(n8959), .ZN(n13343) );
  OR2_X1 U13271 ( .A1(n13348), .A2(n13349), .ZN(n13342) );
  AND2_X1 U13272 ( .A1(n13339), .A2(n13338), .ZN(n13349) );
  AND2_X1 U13273 ( .A1(n13336), .A2(n13350), .ZN(n13348) );
  OR2_X1 U13274 ( .A1(n13338), .A2(n13339), .ZN(n13350) );
  OR2_X1 U13275 ( .A1(n8914), .A2(n8959), .ZN(n13339) );
  OR2_X1 U13276 ( .A1(n13351), .A2(n13352), .ZN(n13338) );
  AND2_X1 U13277 ( .A1(n13335), .A2(n13334), .ZN(n13352) );
  AND2_X1 U13278 ( .A1(n13332), .A2(n13353), .ZN(n13351) );
  OR2_X1 U13279 ( .A1(n13334), .A2(n13335), .ZN(n13353) );
  OR2_X1 U13280 ( .A1(n8918), .A2(n8959), .ZN(n13335) );
  OR2_X1 U13281 ( .A1(n13354), .A2(n13355), .ZN(n13334) );
  AND2_X1 U13282 ( .A1(n13331), .A2(n13330), .ZN(n13355) );
  AND2_X1 U13283 ( .A1(n13328), .A2(n13356), .ZN(n13354) );
  OR2_X1 U13284 ( .A1(n13330), .A2(n13331), .ZN(n13356) );
  OR2_X1 U13285 ( .A1(n8922), .A2(n8959), .ZN(n13331) );
  OR2_X1 U13286 ( .A1(n13357), .A2(n13358), .ZN(n13330) );
  AND2_X1 U13287 ( .A1(n13327), .A2(n13326), .ZN(n13358) );
  AND2_X1 U13288 ( .A1(n13324), .A2(n13359), .ZN(n13357) );
  OR2_X1 U13289 ( .A1(n13326), .A2(n13327), .ZN(n13359) );
  OR2_X1 U13290 ( .A1(n8926), .A2(n8959), .ZN(n13327) );
  OR2_X1 U13291 ( .A1(n13360), .A2(n13361), .ZN(n13326) );
  AND2_X1 U13292 ( .A1(n13323), .A2(n13322), .ZN(n13361) );
  AND2_X1 U13293 ( .A1(n13320), .A2(n13362), .ZN(n13360) );
  OR2_X1 U13294 ( .A1(n13322), .A2(n13323), .ZN(n13362) );
  OR2_X1 U13295 ( .A1(n8930), .A2(n8959), .ZN(n13323) );
  OR2_X1 U13296 ( .A1(n13363), .A2(n13364), .ZN(n13322) );
  AND2_X1 U13297 ( .A1(n13319), .A2(n13318), .ZN(n13364) );
  AND2_X1 U13298 ( .A1(n13316), .A2(n13365), .ZN(n13363) );
  OR2_X1 U13299 ( .A1(n13318), .A2(n13319), .ZN(n13365) );
  OR2_X1 U13300 ( .A1(n8934), .A2(n8959), .ZN(n13319) );
  OR2_X1 U13301 ( .A1(n13366), .A2(n13367), .ZN(n13318) );
  AND2_X1 U13302 ( .A1(n13315), .A2(n13314), .ZN(n13367) );
  AND2_X1 U13303 ( .A1(n13312), .A2(n13368), .ZN(n13366) );
  OR2_X1 U13304 ( .A1(n13314), .A2(n13315), .ZN(n13368) );
  OR2_X1 U13305 ( .A1(n8938), .A2(n8959), .ZN(n13315) );
  OR2_X1 U13306 ( .A1(n13369), .A2(n13370), .ZN(n13314) );
  AND2_X1 U13307 ( .A1(n13311), .A2(n13310), .ZN(n13370) );
  AND2_X1 U13308 ( .A1(n13308), .A2(n13371), .ZN(n13369) );
  OR2_X1 U13309 ( .A1(n13310), .A2(n13311), .ZN(n13371) );
  OR2_X1 U13310 ( .A1(n8942), .A2(n8959), .ZN(n13311) );
  OR2_X1 U13311 ( .A1(n13372), .A2(n13373), .ZN(n13310) );
  AND2_X1 U13312 ( .A1(n13307), .A2(n13306), .ZN(n13373) );
  AND2_X1 U13313 ( .A1(n13304), .A2(n13374), .ZN(n13372) );
  OR2_X1 U13314 ( .A1(n13306), .A2(n13307), .ZN(n13374) );
  OR2_X1 U13315 ( .A1(n8946), .A2(n8959), .ZN(n13307) );
  OR2_X1 U13316 ( .A1(n13375), .A2(n13376), .ZN(n13306) );
  AND2_X1 U13317 ( .A1(n13303), .A2(n13302), .ZN(n13376) );
  AND2_X1 U13318 ( .A1(n13300), .A2(n13377), .ZN(n13375) );
  OR2_X1 U13319 ( .A1(n13302), .A2(n13303), .ZN(n13377) );
  OR2_X1 U13320 ( .A1(n8950), .A2(n8959), .ZN(n13303) );
  OR2_X1 U13321 ( .A1(n13378), .A2(n13379), .ZN(n13302) );
  AND2_X1 U13322 ( .A1(n13299), .A2(n13298), .ZN(n13379) );
  AND2_X1 U13323 ( .A1(n13296), .A2(n13380), .ZN(n13378) );
  OR2_X1 U13324 ( .A1(n13298), .A2(n13299), .ZN(n13380) );
  OR2_X1 U13325 ( .A1(n8954), .A2(n8959), .ZN(n13299) );
  OR2_X1 U13326 ( .A1(n13381), .A2(n13382), .ZN(n13298) );
  AND2_X1 U13327 ( .A1(n8451), .A2(n13295), .ZN(n13382) );
  AND2_X1 U13328 ( .A1(n13293), .A2(n13383), .ZN(n13381) );
  OR2_X1 U13329 ( .A1(n13295), .A2(n8451), .ZN(n13383) );
  OR2_X1 U13330 ( .A1(n8958), .A2(n8959), .ZN(n8451) );
  OR2_X1 U13331 ( .A1(n13384), .A2(n13385), .ZN(n13295) );
  AND2_X1 U13332 ( .A1(n13292), .A2(n13291), .ZN(n13385) );
  AND2_X1 U13333 ( .A1(n13289), .A2(n13386), .ZN(n13384) );
  OR2_X1 U13334 ( .A1(n13291), .A2(n13292), .ZN(n13386) );
  OR2_X1 U13335 ( .A1(n8962), .A2(n8959), .ZN(n13292) );
  OR2_X1 U13336 ( .A1(n13387), .A2(n13388), .ZN(n13291) );
  AND2_X1 U13337 ( .A1(n13288), .A2(n13287), .ZN(n13388) );
  AND2_X1 U13338 ( .A1(n13285), .A2(n13389), .ZN(n13387) );
  OR2_X1 U13339 ( .A1(n13287), .A2(n13288), .ZN(n13389) );
  OR2_X1 U13340 ( .A1(n8966), .A2(n8959), .ZN(n13288) );
  OR2_X1 U13341 ( .A1(n13390), .A2(n13391), .ZN(n13287) );
  AND2_X1 U13342 ( .A1(n13284), .A2(n13283), .ZN(n13391) );
  AND2_X1 U13343 ( .A1(n13281), .A2(n13392), .ZN(n13390) );
  OR2_X1 U13344 ( .A1(n13283), .A2(n13284), .ZN(n13392) );
  OR2_X1 U13345 ( .A1(n8970), .A2(n8959), .ZN(n13284) );
  OR2_X1 U13346 ( .A1(n13393), .A2(n13394), .ZN(n13283) );
  AND2_X1 U13347 ( .A1(n13280), .A2(n13279), .ZN(n13394) );
  AND2_X1 U13348 ( .A1(n13277), .A2(n13395), .ZN(n13393) );
  OR2_X1 U13349 ( .A1(n13279), .A2(n13280), .ZN(n13395) );
  OR2_X1 U13350 ( .A1(n8974), .A2(n8959), .ZN(n13280) );
  OR2_X1 U13351 ( .A1(n13396), .A2(n13397), .ZN(n13279) );
  AND2_X1 U13352 ( .A1(n13276), .A2(n13275), .ZN(n13397) );
  AND2_X1 U13353 ( .A1(n13273), .A2(n13398), .ZN(n13396) );
  OR2_X1 U13354 ( .A1(n13275), .A2(n13276), .ZN(n13398) );
  OR2_X1 U13355 ( .A1(n8978), .A2(n8959), .ZN(n13276) );
  OR2_X1 U13356 ( .A1(n13399), .A2(n13400), .ZN(n13275) );
  AND2_X1 U13357 ( .A1(n13272), .A2(n13271), .ZN(n13400) );
  AND2_X1 U13358 ( .A1(n13269), .A2(n13401), .ZN(n13399) );
  OR2_X1 U13359 ( .A1(n13271), .A2(n13272), .ZN(n13401) );
  OR2_X1 U13360 ( .A1(n8982), .A2(n8959), .ZN(n13272) );
  OR2_X1 U13361 ( .A1(n13402), .A2(n13403), .ZN(n13271) );
  AND2_X1 U13362 ( .A1(n13268), .A2(n13267), .ZN(n13403) );
  AND2_X1 U13363 ( .A1(n13265), .A2(n13404), .ZN(n13402) );
  OR2_X1 U13364 ( .A1(n13267), .A2(n13268), .ZN(n13404) );
  OR2_X1 U13365 ( .A1(n8986), .A2(n8959), .ZN(n13268) );
  OR2_X1 U13366 ( .A1(n13405), .A2(n13406), .ZN(n13267) );
  AND2_X1 U13367 ( .A1(n13264), .A2(n13263), .ZN(n13406) );
  AND2_X1 U13368 ( .A1(n13261), .A2(n13407), .ZN(n13405) );
  OR2_X1 U13369 ( .A1(n13263), .A2(n13264), .ZN(n13407) );
  OR2_X1 U13370 ( .A1(n8990), .A2(n8959), .ZN(n13264) );
  OR2_X1 U13371 ( .A1(n13408), .A2(n13409), .ZN(n13263) );
  AND2_X1 U13372 ( .A1(n13260), .A2(n13259), .ZN(n13409) );
  AND2_X1 U13373 ( .A1(n13257), .A2(n13410), .ZN(n13408) );
  OR2_X1 U13374 ( .A1(n13259), .A2(n13260), .ZN(n13410) );
  OR2_X1 U13375 ( .A1(n8994), .A2(n8959), .ZN(n13260) );
  OR2_X1 U13376 ( .A1(n13411), .A2(n13412), .ZN(n13259) );
  AND2_X1 U13377 ( .A1(n13256), .A2(n13255), .ZN(n13412) );
  AND2_X1 U13378 ( .A1(n13253), .A2(n13413), .ZN(n13411) );
  OR2_X1 U13379 ( .A1(n13255), .A2(n13256), .ZN(n13413) );
  OR2_X1 U13380 ( .A1(n8998), .A2(n8959), .ZN(n13256) );
  OR2_X1 U13381 ( .A1(n13414), .A2(n13415), .ZN(n13255) );
  AND2_X1 U13382 ( .A1(n13252), .A2(n13251), .ZN(n13415) );
  AND2_X1 U13383 ( .A1(n13249), .A2(n13416), .ZN(n13414) );
  OR2_X1 U13384 ( .A1(n13251), .A2(n13252), .ZN(n13416) );
  OR2_X1 U13385 ( .A1(n9002), .A2(n8959), .ZN(n13252) );
  OR2_X1 U13386 ( .A1(n13417), .A2(n13418), .ZN(n13251) );
  AND2_X1 U13387 ( .A1(n13248), .A2(n13247), .ZN(n13418) );
  AND2_X1 U13388 ( .A1(n13245), .A2(n13419), .ZN(n13417) );
  OR2_X1 U13389 ( .A1(n13247), .A2(n13248), .ZN(n13419) );
  OR2_X1 U13390 ( .A1(n9006), .A2(n8959), .ZN(n13248) );
  OR2_X1 U13391 ( .A1(n13420), .A2(n13421), .ZN(n13247) );
  AND2_X1 U13392 ( .A1(n13244), .A2(n13243), .ZN(n13421) );
  AND2_X1 U13393 ( .A1(n13241), .A2(n13422), .ZN(n13420) );
  OR2_X1 U13394 ( .A1(n13243), .A2(n13244), .ZN(n13422) );
  OR2_X1 U13395 ( .A1(n9010), .A2(n8959), .ZN(n13244) );
  OR2_X1 U13396 ( .A1(n13423), .A2(n13424), .ZN(n13243) );
  AND2_X1 U13397 ( .A1(n13238), .A2(n13239), .ZN(n13424) );
  AND2_X1 U13398 ( .A1(n13425), .A2(n13426), .ZN(n13423) );
  OR2_X1 U13399 ( .A1(n13239), .A2(n13238), .ZN(n13426) );
  OR2_X1 U13400 ( .A1(n9014), .A2(n8959), .ZN(n13238) );
  OR2_X1 U13401 ( .A1(n9984), .A2(n13427), .ZN(n13239) );
  OR2_X1 U13402 ( .A1(n8959), .A2(n8955), .ZN(n13427) );
  INV_X1 U13403 ( .A(n13240), .ZN(n13425) );
  OR2_X1 U13404 ( .A1(n13428), .A2(n13429), .ZN(n13240) );
  AND2_X1 U13405 ( .A1(b_14_), .A2(n13430), .ZN(n13429) );
  OR2_X1 U13406 ( .A1(n13431), .A2(n9989), .ZN(n13430) );
  AND2_X1 U13407 ( .A1(a_30_), .A2(n8951), .ZN(n13431) );
  AND2_X1 U13408 ( .A1(b_13_), .A2(n13432), .ZN(n13428) );
  OR2_X1 U13409 ( .A1(n13433), .A2(n8021), .ZN(n13432) );
  AND2_X1 U13410 ( .A1(a_31_), .A2(n8955), .ZN(n13433) );
  XOR2_X1 U13411 ( .A(n13434), .B(n13435), .Z(n13241) );
  XNOR2_X1 U13412 ( .A(n13436), .B(n13437), .ZN(n13434) );
  XOR2_X1 U13413 ( .A(n13438), .B(n13439), .Z(n13245) );
  XOR2_X1 U13414 ( .A(n13440), .B(n13441), .Z(n13439) );
  XOR2_X1 U13415 ( .A(n13442), .B(n13443), .Z(n13249) );
  XOR2_X1 U13416 ( .A(n13444), .B(n13445), .Z(n13443) );
  XOR2_X1 U13417 ( .A(n13446), .B(n13447), .Z(n13253) );
  XOR2_X1 U13418 ( .A(n13448), .B(n13449), .Z(n13447) );
  XOR2_X1 U13419 ( .A(n13450), .B(n13451), .Z(n13257) );
  XOR2_X1 U13420 ( .A(n13452), .B(n13453), .Z(n13451) );
  XOR2_X1 U13421 ( .A(n13454), .B(n13455), .Z(n13261) );
  XOR2_X1 U13422 ( .A(n13456), .B(n13457), .Z(n13455) );
  XOR2_X1 U13423 ( .A(n13458), .B(n13459), .Z(n13265) );
  XOR2_X1 U13424 ( .A(n13460), .B(n13461), .Z(n13459) );
  XOR2_X1 U13425 ( .A(n13462), .B(n13463), .Z(n13269) );
  XOR2_X1 U13426 ( .A(n13464), .B(n13465), .Z(n13463) );
  XOR2_X1 U13427 ( .A(n13466), .B(n13467), .Z(n13273) );
  XOR2_X1 U13428 ( .A(n13468), .B(n13469), .Z(n13467) );
  XOR2_X1 U13429 ( .A(n13470), .B(n13471), .Z(n13277) );
  XOR2_X1 U13430 ( .A(n13472), .B(n13473), .Z(n13471) );
  XOR2_X1 U13431 ( .A(n13474), .B(n13475), .Z(n13281) );
  XOR2_X1 U13432 ( .A(n13476), .B(n13477), .Z(n13475) );
  XOR2_X1 U13433 ( .A(n13478), .B(n13479), .Z(n13285) );
  XOR2_X1 U13434 ( .A(n13480), .B(n13481), .Z(n13479) );
  XOR2_X1 U13435 ( .A(n13482), .B(n13483), .Z(n13289) );
  XOR2_X1 U13436 ( .A(n13484), .B(n13485), .Z(n13483) );
  XOR2_X1 U13437 ( .A(n13486), .B(n13487), .Z(n13293) );
  XOR2_X1 U13438 ( .A(n13488), .B(n13489), .Z(n13487) );
  XOR2_X1 U13439 ( .A(n13490), .B(n13491), .Z(n13296) );
  XOR2_X1 U13440 ( .A(n13492), .B(n13493), .Z(n13491) );
  XOR2_X1 U13441 ( .A(n13494), .B(n13495), .Z(n13300) );
  XOR2_X1 U13442 ( .A(n13496), .B(n8480), .Z(n13495) );
  XOR2_X1 U13443 ( .A(n13497), .B(n13498), .Z(n13304) );
  XOR2_X1 U13444 ( .A(n13499), .B(n13500), .Z(n13498) );
  XOR2_X1 U13445 ( .A(n13501), .B(n13502), .Z(n13308) );
  XOR2_X1 U13446 ( .A(n13503), .B(n13504), .Z(n13502) );
  XOR2_X1 U13447 ( .A(n13505), .B(n13506), .Z(n13312) );
  XOR2_X1 U13448 ( .A(n13507), .B(n13508), .Z(n13506) );
  XOR2_X1 U13449 ( .A(n13509), .B(n13510), .Z(n13316) );
  XOR2_X1 U13450 ( .A(n13511), .B(n13512), .Z(n13510) );
  XOR2_X1 U13451 ( .A(n13513), .B(n13514), .Z(n13320) );
  XOR2_X1 U13452 ( .A(n13515), .B(n13516), .Z(n13514) );
  XOR2_X1 U13453 ( .A(n13517), .B(n13518), .Z(n13324) );
  XOR2_X1 U13454 ( .A(n13519), .B(n13520), .Z(n13518) );
  XOR2_X1 U13455 ( .A(n13521), .B(n13522), .Z(n13328) );
  XOR2_X1 U13456 ( .A(n13523), .B(n13524), .Z(n13522) );
  XOR2_X1 U13457 ( .A(n13525), .B(n13526), .Z(n13332) );
  XOR2_X1 U13458 ( .A(n13527), .B(n13528), .Z(n13526) );
  XOR2_X1 U13459 ( .A(n13529), .B(n13530), .Z(n13336) );
  XOR2_X1 U13460 ( .A(n13531), .B(n13532), .Z(n13530) );
  XOR2_X1 U13461 ( .A(n13533), .B(n13534), .Z(n13340) );
  XOR2_X1 U13462 ( .A(n13535), .B(n13536), .Z(n13534) );
  XOR2_X1 U13463 ( .A(n13537), .B(n13538), .Z(n12711) );
  XOR2_X1 U13464 ( .A(n13539), .B(n13540), .Z(n13538) );
  XNOR2_X1 U13465 ( .A(n9735), .B(n9736), .ZN(n9168) );
  OR2_X1 U13466 ( .A1(n13541), .A2(n13542), .ZN(n9736) );
  AND2_X1 U13467 ( .A1(n9757), .A2(n9756), .ZN(n13542) );
  AND2_X1 U13468 ( .A1(n9754), .A2(n13543), .ZN(n13541) );
  OR2_X1 U13469 ( .A1(n9756), .A2(n9757), .ZN(n13543) );
  OR2_X1 U13470 ( .A1(n9297), .A2(n8955), .ZN(n9757) );
  OR2_X1 U13471 ( .A1(n13544), .A2(n13545), .ZN(n9756) );
  AND2_X1 U13472 ( .A1(n9777), .A2(n9776), .ZN(n13545) );
  AND2_X1 U13473 ( .A1(n9774), .A2(n13546), .ZN(n13544) );
  OR2_X1 U13474 ( .A1(n9776), .A2(n9777), .ZN(n13546) );
  OR2_X1 U13475 ( .A1(n8902), .A2(n8955), .ZN(n9777) );
  OR2_X1 U13476 ( .A1(n13547), .A2(n13548), .ZN(n9776) );
  AND2_X1 U13477 ( .A1(n12716), .A2(n12715), .ZN(n13548) );
  AND2_X1 U13478 ( .A1(n12713), .A2(n13549), .ZN(n13547) );
  OR2_X1 U13479 ( .A1(n12715), .A2(n12716), .ZN(n13549) );
  OR2_X1 U13480 ( .A1(n8906), .A2(n8955), .ZN(n12716) );
  OR2_X1 U13481 ( .A1(n13550), .A2(n13551), .ZN(n12715) );
  AND2_X1 U13482 ( .A1(n13540), .A2(n13539), .ZN(n13551) );
  AND2_X1 U13483 ( .A1(n13537), .A2(n13552), .ZN(n13550) );
  OR2_X1 U13484 ( .A1(n13539), .A2(n13540), .ZN(n13552) );
  OR2_X1 U13485 ( .A1(n8910), .A2(n8955), .ZN(n13540) );
  OR2_X1 U13486 ( .A1(n13553), .A2(n13554), .ZN(n13539) );
  AND2_X1 U13487 ( .A1(n13536), .A2(n13535), .ZN(n13554) );
  AND2_X1 U13488 ( .A1(n13533), .A2(n13555), .ZN(n13553) );
  OR2_X1 U13489 ( .A1(n13535), .A2(n13536), .ZN(n13555) );
  OR2_X1 U13490 ( .A1(n8914), .A2(n8955), .ZN(n13536) );
  OR2_X1 U13491 ( .A1(n13556), .A2(n13557), .ZN(n13535) );
  AND2_X1 U13492 ( .A1(n13532), .A2(n13531), .ZN(n13557) );
  AND2_X1 U13493 ( .A1(n13529), .A2(n13558), .ZN(n13556) );
  OR2_X1 U13494 ( .A1(n13531), .A2(n13532), .ZN(n13558) );
  OR2_X1 U13495 ( .A1(n8918), .A2(n8955), .ZN(n13532) );
  OR2_X1 U13496 ( .A1(n13559), .A2(n13560), .ZN(n13531) );
  AND2_X1 U13497 ( .A1(n13528), .A2(n13527), .ZN(n13560) );
  AND2_X1 U13498 ( .A1(n13525), .A2(n13561), .ZN(n13559) );
  OR2_X1 U13499 ( .A1(n13527), .A2(n13528), .ZN(n13561) );
  OR2_X1 U13500 ( .A1(n8922), .A2(n8955), .ZN(n13528) );
  OR2_X1 U13501 ( .A1(n13562), .A2(n13563), .ZN(n13527) );
  AND2_X1 U13502 ( .A1(n13524), .A2(n13523), .ZN(n13563) );
  AND2_X1 U13503 ( .A1(n13521), .A2(n13564), .ZN(n13562) );
  OR2_X1 U13504 ( .A1(n13523), .A2(n13524), .ZN(n13564) );
  OR2_X1 U13505 ( .A1(n8926), .A2(n8955), .ZN(n13524) );
  OR2_X1 U13506 ( .A1(n13565), .A2(n13566), .ZN(n13523) );
  AND2_X1 U13507 ( .A1(n13520), .A2(n13519), .ZN(n13566) );
  AND2_X1 U13508 ( .A1(n13517), .A2(n13567), .ZN(n13565) );
  OR2_X1 U13509 ( .A1(n13519), .A2(n13520), .ZN(n13567) );
  OR2_X1 U13510 ( .A1(n8930), .A2(n8955), .ZN(n13520) );
  OR2_X1 U13511 ( .A1(n13568), .A2(n13569), .ZN(n13519) );
  AND2_X1 U13512 ( .A1(n13516), .A2(n13515), .ZN(n13569) );
  AND2_X1 U13513 ( .A1(n13513), .A2(n13570), .ZN(n13568) );
  OR2_X1 U13514 ( .A1(n13515), .A2(n13516), .ZN(n13570) );
  OR2_X1 U13515 ( .A1(n8934), .A2(n8955), .ZN(n13516) );
  OR2_X1 U13516 ( .A1(n13571), .A2(n13572), .ZN(n13515) );
  AND2_X1 U13517 ( .A1(n13512), .A2(n13511), .ZN(n13572) );
  AND2_X1 U13518 ( .A1(n13509), .A2(n13573), .ZN(n13571) );
  OR2_X1 U13519 ( .A1(n13511), .A2(n13512), .ZN(n13573) );
  OR2_X1 U13520 ( .A1(n8938), .A2(n8955), .ZN(n13512) );
  OR2_X1 U13521 ( .A1(n13574), .A2(n13575), .ZN(n13511) );
  AND2_X1 U13522 ( .A1(n13508), .A2(n13507), .ZN(n13575) );
  AND2_X1 U13523 ( .A1(n13505), .A2(n13576), .ZN(n13574) );
  OR2_X1 U13524 ( .A1(n13507), .A2(n13508), .ZN(n13576) );
  OR2_X1 U13525 ( .A1(n8942), .A2(n8955), .ZN(n13508) );
  OR2_X1 U13526 ( .A1(n13577), .A2(n13578), .ZN(n13507) );
  AND2_X1 U13527 ( .A1(n13504), .A2(n13503), .ZN(n13578) );
  AND2_X1 U13528 ( .A1(n13501), .A2(n13579), .ZN(n13577) );
  OR2_X1 U13529 ( .A1(n13503), .A2(n13504), .ZN(n13579) );
  OR2_X1 U13530 ( .A1(n8946), .A2(n8955), .ZN(n13504) );
  OR2_X1 U13531 ( .A1(n13580), .A2(n13581), .ZN(n13503) );
  AND2_X1 U13532 ( .A1(n13500), .A2(n13499), .ZN(n13581) );
  AND2_X1 U13533 ( .A1(n13497), .A2(n13582), .ZN(n13580) );
  OR2_X1 U13534 ( .A1(n13499), .A2(n13500), .ZN(n13582) );
  OR2_X1 U13535 ( .A1(n8950), .A2(n8955), .ZN(n13500) );
  OR2_X1 U13536 ( .A1(n13583), .A2(n13584), .ZN(n13499) );
  AND2_X1 U13537 ( .A1(n8480), .A2(n13496), .ZN(n13584) );
  AND2_X1 U13538 ( .A1(n13494), .A2(n13585), .ZN(n13583) );
  OR2_X1 U13539 ( .A1(n13496), .A2(n8480), .ZN(n13585) );
  OR2_X1 U13540 ( .A1(n8954), .A2(n8955), .ZN(n8480) );
  OR2_X1 U13541 ( .A1(n13586), .A2(n13587), .ZN(n13496) );
  AND2_X1 U13542 ( .A1(n13493), .A2(n13492), .ZN(n13587) );
  AND2_X1 U13543 ( .A1(n13490), .A2(n13588), .ZN(n13586) );
  OR2_X1 U13544 ( .A1(n13492), .A2(n13493), .ZN(n13588) );
  OR2_X1 U13545 ( .A1(n8958), .A2(n8955), .ZN(n13493) );
  OR2_X1 U13546 ( .A1(n13589), .A2(n13590), .ZN(n13492) );
  AND2_X1 U13547 ( .A1(n13489), .A2(n13488), .ZN(n13590) );
  AND2_X1 U13548 ( .A1(n13486), .A2(n13591), .ZN(n13589) );
  OR2_X1 U13549 ( .A1(n13488), .A2(n13489), .ZN(n13591) );
  OR2_X1 U13550 ( .A1(n8962), .A2(n8955), .ZN(n13489) );
  OR2_X1 U13551 ( .A1(n13592), .A2(n13593), .ZN(n13488) );
  AND2_X1 U13552 ( .A1(n13485), .A2(n13484), .ZN(n13593) );
  AND2_X1 U13553 ( .A1(n13482), .A2(n13594), .ZN(n13592) );
  OR2_X1 U13554 ( .A1(n13484), .A2(n13485), .ZN(n13594) );
  OR2_X1 U13555 ( .A1(n8966), .A2(n8955), .ZN(n13485) );
  OR2_X1 U13556 ( .A1(n13595), .A2(n13596), .ZN(n13484) );
  AND2_X1 U13557 ( .A1(n13481), .A2(n13480), .ZN(n13596) );
  AND2_X1 U13558 ( .A1(n13478), .A2(n13597), .ZN(n13595) );
  OR2_X1 U13559 ( .A1(n13480), .A2(n13481), .ZN(n13597) );
  OR2_X1 U13560 ( .A1(n8970), .A2(n8955), .ZN(n13481) );
  OR2_X1 U13561 ( .A1(n13598), .A2(n13599), .ZN(n13480) );
  AND2_X1 U13562 ( .A1(n13477), .A2(n13476), .ZN(n13599) );
  AND2_X1 U13563 ( .A1(n13474), .A2(n13600), .ZN(n13598) );
  OR2_X1 U13564 ( .A1(n13476), .A2(n13477), .ZN(n13600) );
  OR2_X1 U13565 ( .A1(n8974), .A2(n8955), .ZN(n13477) );
  OR2_X1 U13566 ( .A1(n13601), .A2(n13602), .ZN(n13476) );
  AND2_X1 U13567 ( .A1(n13473), .A2(n13472), .ZN(n13602) );
  AND2_X1 U13568 ( .A1(n13470), .A2(n13603), .ZN(n13601) );
  OR2_X1 U13569 ( .A1(n13472), .A2(n13473), .ZN(n13603) );
  OR2_X1 U13570 ( .A1(n8978), .A2(n8955), .ZN(n13473) );
  OR2_X1 U13571 ( .A1(n13604), .A2(n13605), .ZN(n13472) );
  AND2_X1 U13572 ( .A1(n13469), .A2(n13468), .ZN(n13605) );
  AND2_X1 U13573 ( .A1(n13466), .A2(n13606), .ZN(n13604) );
  OR2_X1 U13574 ( .A1(n13468), .A2(n13469), .ZN(n13606) );
  OR2_X1 U13575 ( .A1(n8982), .A2(n8955), .ZN(n13469) );
  OR2_X1 U13576 ( .A1(n13607), .A2(n13608), .ZN(n13468) );
  AND2_X1 U13577 ( .A1(n13465), .A2(n13464), .ZN(n13608) );
  AND2_X1 U13578 ( .A1(n13462), .A2(n13609), .ZN(n13607) );
  OR2_X1 U13579 ( .A1(n13464), .A2(n13465), .ZN(n13609) );
  OR2_X1 U13580 ( .A1(n8986), .A2(n8955), .ZN(n13465) );
  OR2_X1 U13581 ( .A1(n13610), .A2(n13611), .ZN(n13464) );
  AND2_X1 U13582 ( .A1(n13461), .A2(n13460), .ZN(n13611) );
  AND2_X1 U13583 ( .A1(n13458), .A2(n13612), .ZN(n13610) );
  OR2_X1 U13584 ( .A1(n13460), .A2(n13461), .ZN(n13612) );
  OR2_X1 U13585 ( .A1(n8990), .A2(n8955), .ZN(n13461) );
  OR2_X1 U13586 ( .A1(n13613), .A2(n13614), .ZN(n13460) );
  AND2_X1 U13587 ( .A1(n13457), .A2(n13456), .ZN(n13614) );
  AND2_X1 U13588 ( .A1(n13454), .A2(n13615), .ZN(n13613) );
  OR2_X1 U13589 ( .A1(n13456), .A2(n13457), .ZN(n13615) );
  OR2_X1 U13590 ( .A1(n8994), .A2(n8955), .ZN(n13457) );
  OR2_X1 U13591 ( .A1(n13616), .A2(n13617), .ZN(n13456) );
  AND2_X1 U13592 ( .A1(n13453), .A2(n13452), .ZN(n13617) );
  AND2_X1 U13593 ( .A1(n13450), .A2(n13618), .ZN(n13616) );
  OR2_X1 U13594 ( .A1(n13452), .A2(n13453), .ZN(n13618) );
  OR2_X1 U13595 ( .A1(n8998), .A2(n8955), .ZN(n13453) );
  OR2_X1 U13596 ( .A1(n13619), .A2(n13620), .ZN(n13452) );
  AND2_X1 U13597 ( .A1(n13449), .A2(n13448), .ZN(n13620) );
  AND2_X1 U13598 ( .A1(n13446), .A2(n13621), .ZN(n13619) );
  OR2_X1 U13599 ( .A1(n13448), .A2(n13449), .ZN(n13621) );
  OR2_X1 U13600 ( .A1(n9002), .A2(n8955), .ZN(n13449) );
  OR2_X1 U13601 ( .A1(n13622), .A2(n13623), .ZN(n13448) );
  AND2_X1 U13602 ( .A1(n13445), .A2(n13444), .ZN(n13623) );
  AND2_X1 U13603 ( .A1(n13442), .A2(n13624), .ZN(n13622) );
  OR2_X1 U13604 ( .A1(n13444), .A2(n13445), .ZN(n13624) );
  OR2_X1 U13605 ( .A1(n9006), .A2(n8955), .ZN(n13445) );
  OR2_X1 U13606 ( .A1(n13625), .A2(n13626), .ZN(n13444) );
  AND2_X1 U13607 ( .A1(n13441), .A2(n13440), .ZN(n13626) );
  AND2_X1 U13608 ( .A1(n13438), .A2(n13627), .ZN(n13625) );
  OR2_X1 U13609 ( .A1(n13440), .A2(n13441), .ZN(n13627) );
  OR2_X1 U13610 ( .A1(n9010), .A2(n8955), .ZN(n13441) );
  OR2_X1 U13611 ( .A1(n13628), .A2(n13629), .ZN(n13440) );
  AND2_X1 U13612 ( .A1(n13435), .A2(n13436), .ZN(n13629) );
  AND2_X1 U13613 ( .A1(n13630), .A2(n13631), .ZN(n13628) );
  OR2_X1 U13614 ( .A1(n13436), .A2(n13435), .ZN(n13631) );
  OR2_X1 U13615 ( .A1(n9014), .A2(n8955), .ZN(n13435) );
  OR2_X1 U13616 ( .A1(n9984), .A2(n13632), .ZN(n13436) );
  OR2_X1 U13617 ( .A1(n8955), .A2(n8951), .ZN(n13632) );
  INV_X1 U13618 ( .A(n13437), .ZN(n13630) );
  OR2_X1 U13619 ( .A1(n13633), .A2(n13634), .ZN(n13437) );
  AND2_X1 U13620 ( .A1(b_13_), .A2(n13635), .ZN(n13634) );
  OR2_X1 U13621 ( .A1(n13636), .A2(n9989), .ZN(n13635) );
  AND2_X1 U13622 ( .A1(a_30_), .A2(n8947), .ZN(n13636) );
  AND2_X1 U13623 ( .A1(b_12_), .A2(n13637), .ZN(n13633) );
  OR2_X1 U13624 ( .A1(n13638), .A2(n8021), .ZN(n13637) );
  AND2_X1 U13625 ( .A1(a_31_), .A2(n8951), .ZN(n13638) );
  XOR2_X1 U13626 ( .A(n13639), .B(n13640), .Z(n13438) );
  XNOR2_X1 U13627 ( .A(n13641), .B(n13642), .ZN(n13639) );
  XOR2_X1 U13628 ( .A(n13643), .B(n13644), .Z(n13442) );
  XOR2_X1 U13629 ( .A(n13645), .B(n13646), .Z(n13644) );
  XOR2_X1 U13630 ( .A(n13647), .B(n13648), .Z(n13446) );
  XOR2_X1 U13631 ( .A(n13649), .B(n13650), .Z(n13648) );
  XOR2_X1 U13632 ( .A(n13651), .B(n13652), .Z(n13450) );
  XOR2_X1 U13633 ( .A(n13653), .B(n13654), .Z(n13652) );
  XOR2_X1 U13634 ( .A(n13655), .B(n13656), .Z(n13454) );
  XOR2_X1 U13635 ( .A(n13657), .B(n13658), .Z(n13656) );
  XOR2_X1 U13636 ( .A(n13659), .B(n13660), .Z(n13458) );
  XOR2_X1 U13637 ( .A(n13661), .B(n13662), .Z(n13660) );
  XOR2_X1 U13638 ( .A(n13663), .B(n13664), .Z(n13462) );
  XOR2_X1 U13639 ( .A(n13665), .B(n13666), .Z(n13664) );
  XOR2_X1 U13640 ( .A(n13667), .B(n13668), .Z(n13466) );
  XOR2_X1 U13641 ( .A(n13669), .B(n13670), .Z(n13668) );
  XOR2_X1 U13642 ( .A(n13671), .B(n13672), .Z(n13470) );
  XOR2_X1 U13643 ( .A(n13673), .B(n13674), .Z(n13672) );
  XOR2_X1 U13644 ( .A(n13675), .B(n13676), .Z(n13474) );
  XOR2_X1 U13645 ( .A(n13677), .B(n13678), .Z(n13676) );
  XOR2_X1 U13646 ( .A(n13679), .B(n13680), .Z(n13478) );
  XOR2_X1 U13647 ( .A(n13681), .B(n13682), .Z(n13680) );
  XOR2_X1 U13648 ( .A(n13683), .B(n13684), .Z(n13482) );
  XOR2_X1 U13649 ( .A(n13685), .B(n13686), .Z(n13684) );
  XOR2_X1 U13650 ( .A(n13687), .B(n13688), .Z(n13486) );
  XOR2_X1 U13651 ( .A(n13689), .B(n13690), .Z(n13688) );
  XOR2_X1 U13652 ( .A(n13691), .B(n13692), .Z(n13490) );
  XOR2_X1 U13653 ( .A(n13693), .B(n13694), .Z(n13692) );
  XOR2_X1 U13654 ( .A(n13695), .B(n13696), .Z(n13494) );
  XOR2_X1 U13655 ( .A(n13697), .B(n13698), .Z(n13696) );
  XOR2_X1 U13656 ( .A(n13699), .B(n13700), .Z(n13497) );
  XOR2_X1 U13657 ( .A(n13701), .B(n13702), .Z(n13700) );
  XOR2_X1 U13658 ( .A(n13703), .B(n13704), .Z(n13501) );
  XOR2_X1 U13659 ( .A(n13705), .B(n8509), .Z(n13704) );
  XOR2_X1 U13660 ( .A(n13706), .B(n13707), .Z(n13505) );
  XOR2_X1 U13661 ( .A(n13708), .B(n13709), .Z(n13707) );
  XOR2_X1 U13662 ( .A(n13710), .B(n13711), .Z(n13509) );
  XOR2_X1 U13663 ( .A(n13712), .B(n13713), .Z(n13711) );
  XOR2_X1 U13664 ( .A(n13714), .B(n13715), .Z(n13513) );
  XOR2_X1 U13665 ( .A(n13716), .B(n13717), .Z(n13715) );
  XOR2_X1 U13666 ( .A(n13718), .B(n13719), .Z(n13517) );
  XOR2_X1 U13667 ( .A(n13720), .B(n13721), .Z(n13719) );
  XOR2_X1 U13668 ( .A(n13722), .B(n13723), .Z(n13521) );
  XOR2_X1 U13669 ( .A(n13724), .B(n13725), .Z(n13723) );
  XOR2_X1 U13670 ( .A(n13726), .B(n13727), .Z(n13525) );
  XOR2_X1 U13671 ( .A(n13728), .B(n13729), .Z(n13727) );
  XOR2_X1 U13672 ( .A(n13730), .B(n13731), .Z(n13529) );
  XOR2_X1 U13673 ( .A(n13732), .B(n13733), .Z(n13731) );
  XOR2_X1 U13674 ( .A(n13734), .B(n13735), .Z(n13533) );
  XOR2_X1 U13675 ( .A(n13736), .B(n13737), .Z(n13735) );
  XOR2_X1 U13676 ( .A(n13738), .B(n13739), .Z(n13537) );
  XOR2_X1 U13677 ( .A(n13740), .B(n13741), .Z(n13739) );
  XOR2_X1 U13678 ( .A(n13742), .B(n13743), .Z(n12713) );
  XOR2_X1 U13679 ( .A(n13744), .B(n13745), .Z(n13743) );
  XOR2_X1 U13680 ( .A(n13746), .B(n13747), .Z(n9774) );
  XOR2_X1 U13681 ( .A(n13748), .B(n13749), .Z(n13747) );
  XOR2_X1 U13682 ( .A(n13750), .B(n13751), .Z(n9754) );
  XOR2_X1 U13683 ( .A(n13752), .B(n13753), .Z(n13751) );
  XNOR2_X1 U13684 ( .A(n13754), .B(n13755), .ZN(n9735) );
  XOR2_X1 U13685 ( .A(n13756), .B(n13757), .Z(n13755) );
  INV_X1 U13686 ( .A(n13758), .ZN(n9177) );
  OR2_X1 U13687 ( .A1(n13759), .A2(n9731), .ZN(n13758) );
  AND2_X1 U13688 ( .A1(n13760), .A2(n13761), .ZN(n13759) );
  INV_X1 U13689 ( .A(n13762), .ZN(n9731) );
  OR2_X1 U13690 ( .A1(n13760), .A2(n13761), .ZN(n13762) );
  OR2_X1 U13691 ( .A1(n13763), .A2(n13764), .ZN(n13761) );
  AND2_X1 U13692 ( .A1(n13757), .A2(n13756), .ZN(n13764) );
  AND2_X1 U13693 ( .A1(n13754), .A2(n13765), .ZN(n13763) );
  OR2_X1 U13694 ( .A1(n13757), .A2(n13756), .ZN(n13765) );
  OR2_X1 U13695 ( .A1(n13766), .A2(n13767), .ZN(n13756) );
  AND2_X1 U13696 ( .A1(n13753), .A2(n13752), .ZN(n13767) );
  AND2_X1 U13697 ( .A1(n13750), .A2(n13768), .ZN(n13766) );
  OR2_X1 U13698 ( .A1(n13753), .A2(n13752), .ZN(n13768) );
  OR2_X1 U13699 ( .A1(n13769), .A2(n13770), .ZN(n13752) );
  AND2_X1 U13700 ( .A1(n13749), .A2(n13748), .ZN(n13770) );
  AND2_X1 U13701 ( .A1(n13746), .A2(n13771), .ZN(n13769) );
  OR2_X1 U13702 ( .A1(n13749), .A2(n13748), .ZN(n13771) );
  OR2_X1 U13703 ( .A1(n13772), .A2(n13773), .ZN(n13748) );
  AND2_X1 U13704 ( .A1(n13745), .A2(n13744), .ZN(n13773) );
  AND2_X1 U13705 ( .A1(n13742), .A2(n13774), .ZN(n13772) );
  OR2_X1 U13706 ( .A1(n13745), .A2(n13744), .ZN(n13774) );
  OR2_X1 U13707 ( .A1(n13775), .A2(n13776), .ZN(n13744) );
  AND2_X1 U13708 ( .A1(n13741), .A2(n13740), .ZN(n13776) );
  AND2_X1 U13709 ( .A1(n13738), .A2(n13777), .ZN(n13775) );
  OR2_X1 U13710 ( .A1(n13741), .A2(n13740), .ZN(n13777) );
  OR2_X1 U13711 ( .A1(n13778), .A2(n13779), .ZN(n13740) );
  AND2_X1 U13712 ( .A1(n13737), .A2(n13736), .ZN(n13779) );
  AND2_X1 U13713 ( .A1(n13734), .A2(n13780), .ZN(n13778) );
  OR2_X1 U13714 ( .A1(n13737), .A2(n13736), .ZN(n13780) );
  OR2_X1 U13715 ( .A1(n13781), .A2(n13782), .ZN(n13736) );
  AND2_X1 U13716 ( .A1(n13733), .A2(n13732), .ZN(n13782) );
  AND2_X1 U13717 ( .A1(n13730), .A2(n13783), .ZN(n13781) );
  OR2_X1 U13718 ( .A1(n13733), .A2(n13732), .ZN(n13783) );
  OR2_X1 U13719 ( .A1(n13784), .A2(n13785), .ZN(n13732) );
  AND2_X1 U13720 ( .A1(n13729), .A2(n13728), .ZN(n13785) );
  AND2_X1 U13721 ( .A1(n13726), .A2(n13786), .ZN(n13784) );
  OR2_X1 U13722 ( .A1(n13729), .A2(n13728), .ZN(n13786) );
  OR2_X1 U13723 ( .A1(n13787), .A2(n13788), .ZN(n13728) );
  AND2_X1 U13724 ( .A1(n13725), .A2(n13724), .ZN(n13788) );
  AND2_X1 U13725 ( .A1(n13722), .A2(n13789), .ZN(n13787) );
  OR2_X1 U13726 ( .A1(n13725), .A2(n13724), .ZN(n13789) );
  OR2_X1 U13727 ( .A1(n13790), .A2(n13791), .ZN(n13724) );
  AND2_X1 U13728 ( .A1(n13721), .A2(n13720), .ZN(n13791) );
  AND2_X1 U13729 ( .A1(n13718), .A2(n13792), .ZN(n13790) );
  OR2_X1 U13730 ( .A1(n13721), .A2(n13720), .ZN(n13792) );
  OR2_X1 U13731 ( .A1(n13793), .A2(n13794), .ZN(n13720) );
  AND2_X1 U13732 ( .A1(n13717), .A2(n13716), .ZN(n13794) );
  AND2_X1 U13733 ( .A1(n13714), .A2(n13795), .ZN(n13793) );
  OR2_X1 U13734 ( .A1(n13717), .A2(n13716), .ZN(n13795) );
  OR2_X1 U13735 ( .A1(n13796), .A2(n13797), .ZN(n13716) );
  AND2_X1 U13736 ( .A1(n13713), .A2(n13712), .ZN(n13797) );
  AND2_X1 U13737 ( .A1(n13710), .A2(n13798), .ZN(n13796) );
  OR2_X1 U13738 ( .A1(n13713), .A2(n13712), .ZN(n13798) );
  OR2_X1 U13739 ( .A1(n13799), .A2(n13800), .ZN(n13712) );
  AND2_X1 U13740 ( .A1(n13709), .A2(n13708), .ZN(n13800) );
  AND2_X1 U13741 ( .A1(n13706), .A2(n13801), .ZN(n13799) );
  OR2_X1 U13742 ( .A1(n13709), .A2(n13708), .ZN(n13801) );
  OR2_X1 U13743 ( .A1(n13802), .A2(n13803), .ZN(n13708) );
  AND2_X1 U13744 ( .A1(n8509), .A2(n13705), .ZN(n13803) );
  AND2_X1 U13745 ( .A1(n13703), .A2(n13804), .ZN(n13802) );
  OR2_X1 U13746 ( .A1(n8509), .A2(n13705), .ZN(n13804) );
  OR2_X1 U13747 ( .A1(n13805), .A2(n13806), .ZN(n13705) );
  AND2_X1 U13748 ( .A1(n13702), .A2(n13701), .ZN(n13806) );
  AND2_X1 U13749 ( .A1(n13699), .A2(n13807), .ZN(n13805) );
  OR2_X1 U13750 ( .A1(n13702), .A2(n13701), .ZN(n13807) );
  OR2_X1 U13751 ( .A1(n13808), .A2(n13809), .ZN(n13701) );
  AND2_X1 U13752 ( .A1(n13698), .A2(n13697), .ZN(n13809) );
  AND2_X1 U13753 ( .A1(n13695), .A2(n13810), .ZN(n13808) );
  OR2_X1 U13754 ( .A1(n13698), .A2(n13697), .ZN(n13810) );
  OR2_X1 U13755 ( .A1(n13811), .A2(n13812), .ZN(n13697) );
  AND2_X1 U13756 ( .A1(n13694), .A2(n13693), .ZN(n13812) );
  AND2_X1 U13757 ( .A1(n13691), .A2(n13813), .ZN(n13811) );
  OR2_X1 U13758 ( .A1(n13694), .A2(n13693), .ZN(n13813) );
  OR2_X1 U13759 ( .A1(n13814), .A2(n13815), .ZN(n13693) );
  AND2_X1 U13760 ( .A1(n13690), .A2(n13689), .ZN(n13815) );
  AND2_X1 U13761 ( .A1(n13687), .A2(n13816), .ZN(n13814) );
  OR2_X1 U13762 ( .A1(n13690), .A2(n13689), .ZN(n13816) );
  OR2_X1 U13763 ( .A1(n13817), .A2(n13818), .ZN(n13689) );
  AND2_X1 U13764 ( .A1(n13686), .A2(n13685), .ZN(n13818) );
  AND2_X1 U13765 ( .A1(n13683), .A2(n13819), .ZN(n13817) );
  OR2_X1 U13766 ( .A1(n13686), .A2(n13685), .ZN(n13819) );
  OR2_X1 U13767 ( .A1(n13820), .A2(n13821), .ZN(n13685) );
  AND2_X1 U13768 ( .A1(n13682), .A2(n13681), .ZN(n13821) );
  AND2_X1 U13769 ( .A1(n13679), .A2(n13822), .ZN(n13820) );
  OR2_X1 U13770 ( .A1(n13682), .A2(n13681), .ZN(n13822) );
  OR2_X1 U13771 ( .A1(n13823), .A2(n13824), .ZN(n13681) );
  AND2_X1 U13772 ( .A1(n13678), .A2(n13677), .ZN(n13824) );
  AND2_X1 U13773 ( .A1(n13675), .A2(n13825), .ZN(n13823) );
  OR2_X1 U13774 ( .A1(n13678), .A2(n13677), .ZN(n13825) );
  OR2_X1 U13775 ( .A1(n13826), .A2(n13827), .ZN(n13677) );
  AND2_X1 U13776 ( .A1(n13674), .A2(n13673), .ZN(n13827) );
  AND2_X1 U13777 ( .A1(n13671), .A2(n13828), .ZN(n13826) );
  OR2_X1 U13778 ( .A1(n13674), .A2(n13673), .ZN(n13828) );
  OR2_X1 U13779 ( .A1(n13829), .A2(n13830), .ZN(n13673) );
  AND2_X1 U13780 ( .A1(n13670), .A2(n13669), .ZN(n13830) );
  AND2_X1 U13781 ( .A1(n13667), .A2(n13831), .ZN(n13829) );
  OR2_X1 U13782 ( .A1(n13670), .A2(n13669), .ZN(n13831) );
  OR2_X1 U13783 ( .A1(n13832), .A2(n13833), .ZN(n13669) );
  AND2_X1 U13784 ( .A1(n13666), .A2(n13665), .ZN(n13833) );
  AND2_X1 U13785 ( .A1(n13663), .A2(n13834), .ZN(n13832) );
  OR2_X1 U13786 ( .A1(n13666), .A2(n13665), .ZN(n13834) );
  OR2_X1 U13787 ( .A1(n13835), .A2(n13836), .ZN(n13665) );
  AND2_X1 U13788 ( .A1(n13662), .A2(n13661), .ZN(n13836) );
  AND2_X1 U13789 ( .A1(n13659), .A2(n13837), .ZN(n13835) );
  OR2_X1 U13790 ( .A1(n13662), .A2(n13661), .ZN(n13837) );
  OR2_X1 U13791 ( .A1(n13838), .A2(n13839), .ZN(n13661) );
  AND2_X1 U13792 ( .A1(n13658), .A2(n13657), .ZN(n13839) );
  AND2_X1 U13793 ( .A1(n13655), .A2(n13840), .ZN(n13838) );
  OR2_X1 U13794 ( .A1(n13658), .A2(n13657), .ZN(n13840) );
  OR2_X1 U13795 ( .A1(n13841), .A2(n13842), .ZN(n13657) );
  AND2_X1 U13796 ( .A1(n13654), .A2(n13653), .ZN(n13842) );
  AND2_X1 U13797 ( .A1(n13651), .A2(n13843), .ZN(n13841) );
  OR2_X1 U13798 ( .A1(n13654), .A2(n13653), .ZN(n13843) );
  OR2_X1 U13799 ( .A1(n13844), .A2(n13845), .ZN(n13653) );
  AND2_X1 U13800 ( .A1(n13650), .A2(n13649), .ZN(n13845) );
  AND2_X1 U13801 ( .A1(n13647), .A2(n13846), .ZN(n13844) );
  OR2_X1 U13802 ( .A1(n13650), .A2(n13649), .ZN(n13846) );
  OR2_X1 U13803 ( .A1(n13847), .A2(n13848), .ZN(n13649) );
  AND2_X1 U13804 ( .A1(n13646), .A2(n13645), .ZN(n13848) );
  AND2_X1 U13805 ( .A1(n13643), .A2(n13849), .ZN(n13847) );
  OR2_X1 U13806 ( .A1(n13646), .A2(n13645), .ZN(n13849) );
  OR2_X1 U13807 ( .A1(n13850), .A2(n13851), .ZN(n13645) );
  AND2_X1 U13808 ( .A1(n13640), .A2(n13641), .ZN(n13851) );
  AND2_X1 U13809 ( .A1(n13852), .A2(n13853), .ZN(n13850) );
  OR2_X1 U13810 ( .A1(n13640), .A2(n13641), .ZN(n13853) );
  OR2_X1 U13811 ( .A1(n9984), .A2(n13854), .ZN(n13641) );
  OR2_X1 U13812 ( .A1(n8951), .A2(n8947), .ZN(n13854) );
  OR2_X1 U13813 ( .A1(n9014), .A2(n8951), .ZN(n13640) );
  INV_X1 U13814 ( .A(n13642), .ZN(n13852) );
  OR2_X1 U13815 ( .A1(n13855), .A2(n13856), .ZN(n13642) );
  AND2_X1 U13816 ( .A1(b_12_), .A2(n13857), .ZN(n13856) );
  OR2_X1 U13817 ( .A1(n13858), .A2(n9989), .ZN(n13857) );
  AND2_X1 U13818 ( .A1(a_30_), .A2(n8943), .ZN(n13858) );
  AND2_X1 U13819 ( .A1(b_11_), .A2(n13859), .ZN(n13855) );
  OR2_X1 U13820 ( .A1(n13860), .A2(n8021), .ZN(n13859) );
  AND2_X1 U13821 ( .A1(a_31_), .A2(n8947), .ZN(n13860) );
  OR2_X1 U13822 ( .A1(n9010), .A2(n8951), .ZN(n13646) );
  XOR2_X1 U13823 ( .A(n13861), .B(n13862), .Z(n13643) );
  XNOR2_X1 U13824 ( .A(n13863), .B(n13864), .ZN(n13861) );
  OR2_X1 U13825 ( .A1(n9006), .A2(n8951), .ZN(n13650) );
  XOR2_X1 U13826 ( .A(n13865), .B(n13866), .Z(n13647) );
  XOR2_X1 U13827 ( .A(n13867), .B(n13868), .Z(n13866) );
  OR2_X1 U13828 ( .A1(n9002), .A2(n8951), .ZN(n13654) );
  XOR2_X1 U13829 ( .A(n13869), .B(n13870), .Z(n13651) );
  XOR2_X1 U13830 ( .A(n13871), .B(n13872), .Z(n13870) );
  OR2_X1 U13831 ( .A1(n8998), .A2(n8951), .ZN(n13658) );
  XOR2_X1 U13832 ( .A(n13873), .B(n13874), .Z(n13655) );
  XOR2_X1 U13833 ( .A(n13875), .B(n13876), .Z(n13874) );
  OR2_X1 U13834 ( .A1(n8994), .A2(n8951), .ZN(n13662) );
  XOR2_X1 U13835 ( .A(n13877), .B(n13878), .Z(n13659) );
  XOR2_X1 U13836 ( .A(n13879), .B(n13880), .Z(n13878) );
  OR2_X1 U13837 ( .A1(n8990), .A2(n8951), .ZN(n13666) );
  XOR2_X1 U13838 ( .A(n13881), .B(n13882), .Z(n13663) );
  XOR2_X1 U13839 ( .A(n13883), .B(n13884), .Z(n13882) );
  OR2_X1 U13840 ( .A1(n8986), .A2(n8951), .ZN(n13670) );
  XOR2_X1 U13841 ( .A(n13885), .B(n13886), .Z(n13667) );
  XOR2_X1 U13842 ( .A(n13887), .B(n13888), .Z(n13886) );
  OR2_X1 U13843 ( .A1(n8982), .A2(n8951), .ZN(n13674) );
  XOR2_X1 U13844 ( .A(n13889), .B(n13890), .Z(n13671) );
  XOR2_X1 U13845 ( .A(n13891), .B(n13892), .Z(n13890) );
  OR2_X1 U13846 ( .A1(n8978), .A2(n8951), .ZN(n13678) );
  XOR2_X1 U13847 ( .A(n13893), .B(n13894), .Z(n13675) );
  XOR2_X1 U13848 ( .A(n13895), .B(n13896), .Z(n13894) );
  OR2_X1 U13849 ( .A1(n8974), .A2(n8951), .ZN(n13682) );
  XOR2_X1 U13850 ( .A(n13897), .B(n13898), .Z(n13679) );
  XOR2_X1 U13851 ( .A(n13899), .B(n13900), .Z(n13898) );
  OR2_X1 U13852 ( .A1(n8970), .A2(n8951), .ZN(n13686) );
  XOR2_X1 U13853 ( .A(n13901), .B(n13902), .Z(n13683) );
  XOR2_X1 U13854 ( .A(n13903), .B(n13904), .Z(n13902) );
  OR2_X1 U13855 ( .A1(n8966), .A2(n8951), .ZN(n13690) );
  XOR2_X1 U13856 ( .A(n13905), .B(n13906), .Z(n13687) );
  XOR2_X1 U13857 ( .A(n13907), .B(n13908), .Z(n13906) );
  OR2_X1 U13858 ( .A1(n8962), .A2(n8951), .ZN(n13694) );
  XOR2_X1 U13859 ( .A(n13909), .B(n13910), .Z(n13691) );
  XOR2_X1 U13860 ( .A(n13911), .B(n13912), .Z(n13910) );
  OR2_X1 U13861 ( .A1(n8958), .A2(n8951), .ZN(n13698) );
  XOR2_X1 U13862 ( .A(n13913), .B(n13914), .Z(n13695) );
  XOR2_X1 U13863 ( .A(n13915), .B(n13916), .Z(n13914) );
  OR2_X1 U13864 ( .A1(n8954), .A2(n8951), .ZN(n13702) );
  XOR2_X1 U13865 ( .A(n13917), .B(n13918), .Z(n13699) );
  XOR2_X1 U13866 ( .A(n13919), .B(n13920), .Z(n13918) );
  OR2_X1 U13867 ( .A1(n8950), .A2(n8951), .ZN(n8509) );
  XOR2_X1 U13868 ( .A(n13921), .B(n13922), .Z(n13703) );
  XOR2_X1 U13869 ( .A(n13923), .B(n13924), .Z(n13922) );
  OR2_X1 U13870 ( .A1(n8946), .A2(n8951), .ZN(n13709) );
  XOR2_X1 U13871 ( .A(n13925), .B(n13926), .Z(n13706) );
  XOR2_X1 U13872 ( .A(n13927), .B(n13928), .Z(n13926) );
  OR2_X1 U13873 ( .A1(n8942), .A2(n8951), .ZN(n13713) );
  XOR2_X1 U13874 ( .A(n13929), .B(n13930), .Z(n13710) );
  XOR2_X1 U13875 ( .A(n13931), .B(n8538), .Z(n13930) );
  OR2_X1 U13876 ( .A1(n8938), .A2(n8951), .ZN(n13717) );
  XOR2_X1 U13877 ( .A(n13932), .B(n13933), .Z(n13714) );
  XOR2_X1 U13878 ( .A(n13934), .B(n13935), .Z(n13933) );
  OR2_X1 U13879 ( .A1(n8934), .A2(n8951), .ZN(n13721) );
  XOR2_X1 U13880 ( .A(n13936), .B(n13937), .Z(n13718) );
  XOR2_X1 U13881 ( .A(n13938), .B(n13939), .Z(n13937) );
  OR2_X1 U13882 ( .A1(n8930), .A2(n8951), .ZN(n13725) );
  XOR2_X1 U13883 ( .A(n13940), .B(n13941), .Z(n13722) );
  XOR2_X1 U13884 ( .A(n13942), .B(n13943), .Z(n13941) );
  OR2_X1 U13885 ( .A1(n8926), .A2(n8951), .ZN(n13729) );
  XOR2_X1 U13886 ( .A(n13944), .B(n13945), .Z(n13726) );
  XOR2_X1 U13887 ( .A(n13946), .B(n13947), .Z(n13945) );
  OR2_X1 U13888 ( .A1(n8922), .A2(n8951), .ZN(n13733) );
  XOR2_X1 U13889 ( .A(n13948), .B(n13949), .Z(n13730) );
  XOR2_X1 U13890 ( .A(n13950), .B(n13951), .Z(n13949) );
  OR2_X1 U13891 ( .A1(n8918), .A2(n8951), .ZN(n13737) );
  XOR2_X1 U13892 ( .A(n13952), .B(n13953), .Z(n13734) );
  XOR2_X1 U13893 ( .A(n13954), .B(n13955), .Z(n13953) );
  OR2_X1 U13894 ( .A1(n8914), .A2(n8951), .ZN(n13741) );
  XOR2_X1 U13895 ( .A(n13956), .B(n13957), .Z(n13738) );
  XOR2_X1 U13896 ( .A(n13958), .B(n13959), .Z(n13957) );
  OR2_X1 U13897 ( .A1(n8910), .A2(n8951), .ZN(n13745) );
  XOR2_X1 U13898 ( .A(n13960), .B(n13961), .Z(n13742) );
  XOR2_X1 U13899 ( .A(n13962), .B(n13963), .Z(n13961) );
  OR2_X1 U13900 ( .A1(n8906), .A2(n8951), .ZN(n13749) );
  XOR2_X1 U13901 ( .A(n13964), .B(n13965), .Z(n13746) );
  XOR2_X1 U13902 ( .A(n13966), .B(n13967), .Z(n13965) );
  OR2_X1 U13903 ( .A1(n8902), .A2(n8951), .ZN(n13753) );
  XOR2_X1 U13904 ( .A(n13968), .B(n13969), .Z(n13750) );
  XOR2_X1 U13905 ( .A(n13970), .B(n13971), .Z(n13969) );
  OR2_X1 U13906 ( .A1(n9297), .A2(n8951), .ZN(n13757) );
  XOR2_X1 U13907 ( .A(n13972), .B(n13973), .Z(n13754) );
  XOR2_X1 U13908 ( .A(n13974), .B(n13975), .Z(n13973) );
  XOR2_X1 U13909 ( .A(n9725), .B(n13976), .Z(n13760) );
  XOR2_X1 U13910 ( .A(n9724), .B(n9723), .Z(n13976) );
  OR2_X1 U13911 ( .A1(n9297), .A2(n8947), .ZN(n9723) );
  OR2_X1 U13912 ( .A1(n13977), .A2(n13978), .ZN(n9724) );
  AND2_X1 U13913 ( .A1(n13975), .A2(n13974), .ZN(n13978) );
  AND2_X1 U13914 ( .A1(n13972), .A2(n13979), .ZN(n13977) );
  OR2_X1 U13915 ( .A1(n13974), .A2(n13975), .ZN(n13979) );
  OR2_X1 U13916 ( .A1(n8902), .A2(n8947), .ZN(n13975) );
  OR2_X1 U13917 ( .A1(n13980), .A2(n13981), .ZN(n13974) );
  AND2_X1 U13918 ( .A1(n13971), .A2(n13970), .ZN(n13981) );
  AND2_X1 U13919 ( .A1(n13968), .A2(n13982), .ZN(n13980) );
  OR2_X1 U13920 ( .A1(n13970), .A2(n13971), .ZN(n13982) );
  OR2_X1 U13921 ( .A1(n8906), .A2(n8947), .ZN(n13971) );
  OR2_X1 U13922 ( .A1(n13983), .A2(n13984), .ZN(n13970) );
  AND2_X1 U13923 ( .A1(n13967), .A2(n13966), .ZN(n13984) );
  AND2_X1 U13924 ( .A1(n13964), .A2(n13985), .ZN(n13983) );
  OR2_X1 U13925 ( .A1(n13966), .A2(n13967), .ZN(n13985) );
  OR2_X1 U13926 ( .A1(n8910), .A2(n8947), .ZN(n13967) );
  OR2_X1 U13927 ( .A1(n13986), .A2(n13987), .ZN(n13966) );
  AND2_X1 U13928 ( .A1(n13963), .A2(n13962), .ZN(n13987) );
  AND2_X1 U13929 ( .A1(n13960), .A2(n13988), .ZN(n13986) );
  OR2_X1 U13930 ( .A1(n13962), .A2(n13963), .ZN(n13988) );
  OR2_X1 U13931 ( .A1(n8914), .A2(n8947), .ZN(n13963) );
  OR2_X1 U13932 ( .A1(n13989), .A2(n13990), .ZN(n13962) );
  AND2_X1 U13933 ( .A1(n13959), .A2(n13958), .ZN(n13990) );
  AND2_X1 U13934 ( .A1(n13956), .A2(n13991), .ZN(n13989) );
  OR2_X1 U13935 ( .A1(n13958), .A2(n13959), .ZN(n13991) );
  OR2_X1 U13936 ( .A1(n8918), .A2(n8947), .ZN(n13959) );
  OR2_X1 U13937 ( .A1(n13992), .A2(n13993), .ZN(n13958) );
  AND2_X1 U13938 ( .A1(n13955), .A2(n13954), .ZN(n13993) );
  AND2_X1 U13939 ( .A1(n13952), .A2(n13994), .ZN(n13992) );
  OR2_X1 U13940 ( .A1(n13954), .A2(n13955), .ZN(n13994) );
  OR2_X1 U13941 ( .A1(n8922), .A2(n8947), .ZN(n13955) );
  OR2_X1 U13942 ( .A1(n13995), .A2(n13996), .ZN(n13954) );
  AND2_X1 U13943 ( .A1(n13951), .A2(n13950), .ZN(n13996) );
  AND2_X1 U13944 ( .A1(n13948), .A2(n13997), .ZN(n13995) );
  OR2_X1 U13945 ( .A1(n13950), .A2(n13951), .ZN(n13997) );
  OR2_X1 U13946 ( .A1(n8926), .A2(n8947), .ZN(n13951) );
  OR2_X1 U13947 ( .A1(n13998), .A2(n13999), .ZN(n13950) );
  AND2_X1 U13948 ( .A1(n13947), .A2(n13946), .ZN(n13999) );
  AND2_X1 U13949 ( .A1(n13944), .A2(n14000), .ZN(n13998) );
  OR2_X1 U13950 ( .A1(n13946), .A2(n13947), .ZN(n14000) );
  OR2_X1 U13951 ( .A1(n8930), .A2(n8947), .ZN(n13947) );
  OR2_X1 U13952 ( .A1(n14001), .A2(n14002), .ZN(n13946) );
  AND2_X1 U13953 ( .A1(n13943), .A2(n13942), .ZN(n14002) );
  AND2_X1 U13954 ( .A1(n13940), .A2(n14003), .ZN(n14001) );
  OR2_X1 U13955 ( .A1(n13942), .A2(n13943), .ZN(n14003) );
  OR2_X1 U13956 ( .A1(n8934), .A2(n8947), .ZN(n13943) );
  OR2_X1 U13957 ( .A1(n14004), .A2(n14005), .ZN(n13942) );
  AND2_X1 U13958 ( .A1(n13939), .A2(n13938), .ZN(n14005) );
  AND2_X1 U13959 ( .A1(n13936), .A2(n14006), .ZN(n14004) );
  OR2_X1 U13960 ( .A1(n13938), .A2(n13939), .ZN(n14006) );
  OR2_X1 U13961 ( .A1(n8938), .A2(n8947), .ZN(n13939) );
  OR2_X1 U13962 ( .A1(n14007), .A2(n14008), .ZN(n13938) );
  AND2_X1 U13963 ( .A1(n13935), .A2(n13934), .ZN(n14008) );
  AND2_X1 U13964 ( .A1(n13932), .A2(n14009), .ZN(n14007) );
  OR2_X1 U13965 ( .A1(n13934), .A2(n13935), .ZN(n14009) );
  OR2_X1 U13966 ( .A1(n8942), .A2(n8947), .ZN(n13935) );
  OR2_X1 U13967 ( .A1(n14010), .A2(n14011), .ZN(n13934) );
  AND2_X1 U13968 ( .A1(n8538), .A2(n13931), .ZN(n14011) );
  AND2_X1 U13969 ( .A1(n13929), .A2(n14012), .ZN(n14010) );
  OR2_X1 U13970 ( .A1(n13931), .A2(n8538), .ZN(n14012) );
  OR2_X1 U13971 ( .A1(n8946), .A2(n8947), .ZN(n8538) );
  OR2_X1 U13972 ( .A1(n14013), .A2(n14014), .ZN(n13931) );
  AND2_X1 U13973 ( .A1(n13928), .A2(n13927), .ZN(n14014) );
  AND2_X1 U13974 ( .A1(n13925), .A2(n14015), .ZN(n14013) );
  OR2_X1 U13975 ( .A1(n13927), .A2(n13928), .ZN(n14015) );
  OR2_X1 U13976 ( .A1(n8950), .A2(n8947), .ZN(n13928) );
  OR2_X1 U13977 ( .A1(n14016), .A2(n14017), .ZN(n13927) );
  AND2_X1 U13978 ( .A1(n13924), .A2(n13923), .ZN(n14017) );
  AND2_X1 U13979 ( .A1(n13921), .A2(n14018), .ZN(n14016) );
  OR2_X1 U13980 ( .A1(n13923), .A2(n13924), .ZN(n14018) );
  OR2_X1 U13981 ( .A1(n8954), .A2(n8947), .ZN(n13924) );
  OR2_X1 U13982 ( .A1(n14019), .A2(n14020), .ZN(n13923) );
  AND2_X1 U13983 ( .A1(n13920), .A2(n13919), .ZN(n14020) );
  AND2_X1 U13984 ( .A1(n13917), .A2(n14021), .ZN(n14019) );
  OR2_X1 U13985 ( .A1(n13919), .A2(n13920), .ZN(n14021) );
  OR2_X1 U13986 ( .A1(n8958), .A2(n8947), .ZN(n13920) );
  OR2_X1 U13987 ( .A1(n14022), .A2(n14023), .ZN(n13919) );
  AND2_X1 U13988 ( .A1(n13916), .A2(n13915), .ZN(n14023) );
  AND2_X1 U13989 ( .A1(n13913), .A2(n14024), .ZN(n14022) );
  OR2_X1 U13990 ( .A1(n13915), .A2(n13916), .ZN(n14024) );
  OR2_X1 U13991 ( .A1(n8962), .A2(n8947), .ZN(n13916) );
  OR2_X1 U13992 ( .A1(n14025), .A2(n14026), .ZN(n13915) );
  AND2_X1 U13993 ( .A1(n13912), .A2(n13911), .ZN(n14026) );
  AND2_X1 U13994 ( .A1(n13909), .A2(n14027), .ZN(n14025) );
  OR2_X1 U13995 ( .A1(n13911), .A2(n13912), .ZN(n14027) );
  OR2_X1 U13996 ( .A1(n8966), .A2(n8947), .ZN(n13912) );
  OR2_X1 U13997 ( .A1(n14028), .A2(n14029), .ZN(n13911) );
  AND2_X1 U13998 ( .A1(n13908), .A2(n13907), .ZN(n14029) );
  AND2_X1 U13999 ( .A1(n13905), .A2(n14030), .ZN(n14028) );
  OR2_X1 U14000 ( .A1(n13907), .A2(n13908), .ZN(n14030) );
  OR2_X1 U14001 ( .A1(n8970), .A2(n8947), .ZN(n13908) );
  OR2_X1 U14002 ( .A1(n14031), .A2(n14032), .ZN(n13907) );
  AND2_X1 U14003 ( .A1(n13904), .A2(n13903), .ZN(n14032) );
  AND2_X1 U14004 ( .A1(n13901), .A2(n14033), .ZN(n14031) );
  OR2_X1 U14005 ( .A1(n13903), .A2(n13904), .ZN(n14033) );
  OR2_X1 U14006 ( .A1(n8974), .A2(n8947), .ZN(n13904) );
  OR2_X1 U14007 ( .A1(n14034), .A2(n14035), .ZN(n13903) );
  AND2_X1 U14008 ( .A1(n13900), .A2(n13899), .ZN(n14035) );
  AND2_X1 U14009 ( .A1(n13897), .A2(n14036), .ZN(n14034) );
  OR2_X1 U14010 ( .A1(n13899), .A2(n13900), .ZN(n14036) );
  OR2_X1 U14011 ( .A1(n8978), .A2(n8947), .ZN(n13900) );
  OR2_X1 U14012 ( .A1(n14037), .A2(n14038), .ZN(n13899) );
  AND2_X1 U14013 ( .A1(n13896), .A2(n13895), .ZN(n14038) );
  AND2_X1 U14014 ( .A1(n13893), .A2(n14039), .ZN(n14037) );
  OR2_X1 U14015 ( .A1(n13895), .A2(n13896), .ZN(n14039) );
  OR2_X1 U14016 ( .A1(n8982), .A2(n8947), .ZN(n13896) );
  OR2_X1 U14017 ( .A1(n14040), .A2(n14041), .ZN(n13895) );
  AND2_X1 U14018 ( .A1(n13892), .A2(n13891), .ZN(n14041) );
  AND2_X1 U14019 ( .A1(n13889), .A2(n14042), .ZN(n14040) );
  OR2_X1 U14020 ( .A1(n13891), .A2(n13892), .ZN(n14042) );
  OR2_X1 U14021 ( .A1(n8986), .A2(n8947), .ZN(n13892) );
  OR2_X1 U14022 ( .A1(n14043), .A2(n14044), .ZN(n13891) );
  AND2_X1 U14023 ( .A1(n13888), .A2(n13887), .ZN(n14044) );
  AND2_X1 U14024 ( .A1(n13885), .A2(n14045), .ZN(n14043) );
  OR2_X1 U14025 ( .A1(n13887), .A2(n13888), .ZN(n14045) );
  OR2_X1 U14026 ( .A1(n8990), .A2(n8947), .ZN(n13888) );
  OR2_X1 U14027 ( .A1(n14046), .A2(n14047), .ZN(n13887) );
  AND2_X1 U14028 ( .A1(n13884), .A2(n13883), .ZN(n14047) );
  AND2_X1 U14029 ( .A1(n13881), .A2(n14048), .ZN(n14046) );
  OR2_X1 U14030 ( .A1(n13883), .A2(n13884), .ZN(n14048) );
  OR2_X1 U14031 ( .A1(n8994), .A2(n8947), .ZN(n13884) );
  OR2_X1 U14032 ( .A1(n14049), .A2(n14050), .ZN(n13883) );
  AND2_X1 U14033 ( .A1(n13880), .A2(n13879), .ZN(n14050) );
  AND2_X1 U14034 ( .A1(n13877), .A2(n14051), .ZN(n14049) );
  OR2_X1 U14035 ( .A1(n13879), .A2(n13880), .ZN(n14051) );
  OR2_X1 U14036 ( .A1(n8998), .A2(n8947), .ZN(n13880) );
  OR2_X1 U14037 ( .A1(n14052), .A2(n14053), .ZN(n13879) );
  AND2_X1 U14038 ( .A1(n13876), .A2(n13875), .ZN(n14053) );
  AND2_X1 U14039 ( .A1(n13873), .A2(n14054), .ZN(n14052) );
  OR2_X1 U14040 ( .A1(n13875), .A2(n13876), .ZN(n14054) );
  OR2_X1 U14041 ( .A1(n9002), .A2(n8947), .ZN(n13876) );
  OR2_X1 U14042 ( .A1(n14055), .A2(n14056), .ZN(n13875) );
  AND2_X1 U14043 ( .A1(n13872), .A2(n13871), .ZN(n14056) );
  AND2_X1 U14044 ( .A1(n13869), .A2(n14057), .ZN(n14055) );
  OR2_X1 U14045 ( .A1(n13871), .A2(n13872), .ZN(n14057) );
  OR2_X1 U14046 ( .A1(n9006), .A2(n8947), .ZN(n13872) );
  OR2_X1 U14047 ( .A1(n14058), .A2(n14059), .ZN(n13871) );
  AND2_X1 U14048 ( .A1(n13868), .A2(n13867), .ZN(n14059) );
  AND2_X1 U14049 ( .A1(n13865), .A2(n14060), .ZN(n14058) );
  OR2_X1 U14050 ( .A1(n13867), .A2(n13868), .ZN(n14060) );
  OR2_X1 U14051 ( .A1(n9010), .A2(n8947), .ZN(n13868) );
  OR2_X1 U14052 ( .A1(n14061), .A2(n14062), .ZN(n13867) );
  AND2_X1 U14053 ( .A1(n13862), .A2(n13863), .ZN(n14062) );
  AND2_X1 U14054 ( .A1(n14063), .A2(n14064), .ZN(n14061) );
  OR2_X1 U14055 ( .A1(n13863), .A2(n13862), .ZN(n14064) );
  OR2_X1 U14056 ( .A1(n9014), .A2(n8947), .ZN(n13862) );
  OR2_X1 U14057 ( .A1(n9984), .A2(n14065), .ZN(n13863) );
  OR2_X1 U14058 ( .A1(n8947), .A2(n8943), .ZN(n14065) );
  INV_X1 U14059 ( .A(n13864), .ZN(n14063) );
  OR2_X1 U14060 ( .A1(n14066), .A2(n14067), .ZN(n13864) );
  AND2_X1 U14061 ( .A1(b_11_), .A2(n14068), .ZN(n14067) );
  OR2_X1 U14062 ( .A1(n14069), .A2(n9989), .ZN(n14068) );
  AND2_X1 U14063 ( .A1(a_30_), .A2(n8939), .ZN(n14069) );
  AND2_X1 U14064 ( .A1(b_10_), .A2(n14070), .ZN(n14066) );
  OR2_X1 U14065 ( .A1(n14071), .A2(n8021), .ZN(n14070) );
  AND2_X1 U14066 ( .A1(a_31_), .A2(n8943), .ZN(n14071) );
  XOR2_X1 U14067 ( .A(n14072), .B(n14073), .Z(n13865) );
  XNOR2_X1 U14068 ( .A(n14074), .B(n14075), .ZN(n14072) );
  XOR2_X1 U14069 ( .A(n14076), .B(n14077), .Z(n13869) );
  XOR2_X1 U14070 ( .A(n14078), .B(n14079), .Z(n14077) );
  XOR2_X1 U14071 ( .A(n14080), .B(n14081), .Z(n13873) );
  XOR2_X1 U14072 ( .A(n14082), .B(n14083), .Z(n14081) );
  XOR2_X1 U14073 ( .A(n14084), .B(n14085), .Z(n13877) );
  XOR2_X1 U14074 ( .A(n14086), .B(n14087), .Z(n14085) );
  XOR2_X1 U14075 ( .A(n14088), .B(n14089), .Z(n13881) );
  XOR2_X1 U14076 ( .A(n14090), .B(n14091), .Z(n14089) );
  XOR2_X1 U14077 ( .A(n14092), .B(n14093), .Z(n13885) );
  XOR2_X1 U14078 ( .A(n14094), .B(n14095), .Z(n14093) );
  XOR2_X1 U14079 ( .A(n14096), .B(n14097), .Z(n13889) );
  XOR2_X1 U14080 ( .A(n14098), .B(n14099), .Z(n14097) );
  XOR2_X1 U14081 ( .A(n14100), .B(n14101), .Z(n13893) );
  XOR2_X1 U14082 ( .A(n14102), .B(n14103), .Z(n14101) );
  XOR2_X1 U14083 ( .A(n14104), .B(n14105), .Z(n13897) );
  XOR2_X1 U14084 ( .A(n14106), .B(n14107), .Z(n14105) );
  XOR2_X1 U14085 ( .A(n14108), .B(n14109), .Z(n13901) );
  XOR2_X1 U14086 ( .A(n14110), .B(n14111), .Z(n14109) );
  XOR2_X1 U14087 ( .A(n14112), .B(n14113), .Z(n13905) );
  XOR2_X1 U14088 ( .A(n14114), .B(n14115), .Z(n14113) );
  XOR2_X1 U14089 ( .A(n14116), .B(n14117), .Z(n13909) );
  XOR2_X1 U14090 ( .A(n14118), .B(n14119), .Z(n14117) );
  XOR2_X1 U14091 ( .A(n14120), .B(n14121), .Z(n13913) );
  XOR2_X1 U14092 ( .A(n14122), .B(n14123), .Z(n14121) );
  XOR2_X1 U14093 ( .A(n14124), .B(n14125), .Z(n13917) );
  XOR2_X1 U14094 ( .A(n14126), .B(n14127), .Z(n14125) );
  XOR2_X1 U14095 ( .A(n14128), .B(n14129), .Z(n13921) );
  XOR2_X1 U14096 ( .A(n14130), .B(n14131), .Z(n14129) );
  XOR2_X1 U14097 ( .A(n14132), .B(n14133), .Z(n13925) );
  XOR2_X1 U14098 ( .A(n14134), .B(n14135), .Z(n14133) );
  XOR2_X1 U14099 ( .A(n14136), .B(n14137), .Z(n13929) );
  XOR2_X1 U14100 ( .A(n14138), .B(n14139), .Z(n14137) );
  XOR2_X1 U14101 ( .A(n14140), .B(n14141), .Z(n13932) );
  XOR2_X1 U14102 ( .A(n14142), .B(n14143), .Z(n14141) );
  XOR2_X1 U14103 ( .A(n14144), .B(n14145), .Z(n13936) );
  XOR2_X1 U14104 ( .A(n14146), .B(n8567), .Z(n14145) );
  XOR2_X1 U14105 ( .A(n14147), .B(n14148), .Z(n13940) );
  XOR2_X1 U14106 ( .A(n14149), .B(n14150), .Z(n14148) );
  XOR2_X1 U14107 ( .A(n14151), .B(n14152), .Z(n13944) );
  XOR2_X1 U14108 ( .A(n14153), .B(n14154), .Z(n14152) );
  XOR2_X1 U14109 ( .A(n14155), .B(n14156), .Z(n13948) );
  XOR2_X1 U14110 ( .A(n14157), .B(n14158), .Z(n14156) );
  XOR2_X1 U14111 ( .A(n14159), .B(n14160), .Z(n13952) );
  XOR2_X1 U14112 ( .A(n14161), .B(n14162), .Z(n14160) );
  XOR2_X1 U14113 ( .A(n14163), .B(n14164), .Z(n13956) );
  XOR2_X1 U14114 ( .A(n14165), .B(n14166), .Z(n14164) );
  XOR2_X1 U14115 ( .A(n14167), .B(n14168), .Z(n13960) );
  XOR2_X1 U14116 ( .A(n14169), .B(n14170), .Z(n14168) );
  XOR2_X1 U14117 ( .A(n14171), .B(n14172), .Z(n13964) );
  XOR2_X1 U14118 ( .A(n14173), .B(n14174), .Z(n14172) );
  XOR2_X1 U14119 ( .A(n14175), .B(n14176), .Z(n13968) );
  XOR2_X1 U14120 ( .A(n14177), .B(n14178), .Z(n14176) );
  XOR2_X1 U14121 ( .A(n14179), .B(n14180), .Z(n13972) );
  XOR2_X1 U14122 ( .A(n14181), .B(n14182), .Z(n14180) );
  XOR2_X1 U14123 ( .A(n14183), .B(n14184), .Z(n9725) );
  XOR2_X1 U14124 ( .A(n14185), .B(n14186), .Z(n14184) );
  INV_X1 U14125 ( .A(n14187), .ZN(n9711) );
  OR2_X1 U14126 ( .A1(n9719), .A2(n9720), .ZN(n14187) );
  OR2_X1 U14127 ( .A1(n14188), .A2(n14189), .ZN(n9720) );
  AND2_X1 U14128 ( .A1(n9730), .A2(n9729), .ZN(n14189) );
  AND2_X1 U14129 ( .A1(n9727), .A2(n14190), .ZN(n14188) );
  OR2_X1 U14130 ( .A1(n9730), .A2(n9729), .ZN(n14190) );
  OR2_X1 U14131 ( .A1(n14191), .A2(n14192), .ZN(n9729) );
  AND2_X1 U14132 ( .A1(n14186), .A2(n14185), .ZN(n14192) );
  AND2_X1 U14133 ( .A1(n14183), .A2(n14193), .ZN(n14191) );
  OR2_X1 U14134 ( .A1(n14186), .A2(n14185), .ZN(n14193) );
  OR2_X1 U14135 ( .A1(n14194), .A2(n14195), .ZN(n14185) );
  AND2_X1 U14136 ( .A1(n14182), .A2(n14181), .ZN(n14195) );
  AND2_X1 U14137 ( .A1(n14179), .A2(n14196), .ZN(n14194) );
  OR2_X1 U14138 ( .A1(n14182), .A2(n14181), .ZN(n14196) );
  OR2_X1 U14139 ( .A1(n14197), .A2(n14198), .ZN(n14181) );
  AND2_X1 U14140 ( .A1(n14178), .A2(n14177), .ZN(n14198) );
  AND2_X1 U14141 ( .A1(n14175), .A2(n14199), .ZN(n14197) );
  OR2_X1 U14142 ( .A1(n14178), .A2(n14177), .ZN(n14199) );
  OR2_X1 U14143 ( .A1(n14200), .A2(n14201), .ZN(n14177) );
  AND2_X1 U14144 ( .A1(n14174), .A2(n14173), .ZN(n14201) );
  AND2_X1 U14145 ( .A1(n14171), .A2(n14202), .ZN(n14200) );
  OR2_X1 U14146 ( .A1(n14174), .A2(n14173), .ZN(n14202) );
  OR2_X1 U14147 ( .A1(n14203), .A2(n14204), .ZN(n14173) );
  AND2_X1 U14148 ( .A1(n14170), .A2(n14169), .ZN(n14204) );
  AND2_X1 U14149 ( .A1(n14167), .A2(n14205), .ZN(n14203) );
  OR2_X1 U14150 ( .A1(n14170), .A2(n14169), .ZN(n14205) );
  OR2_X1 U14151 ( .A1(n14206), .A2(n14207), .ZN(n14169) );
  AND2_X1 U14152 ( .A1(n14166), .A2(n14165), .ZN(n14207) );
  AND2_X1 U14153 ( .A1(n14163), .A2(n14208), .ZN(n14206) );
  OR2_X1 U14154 ( .A1(n14166), .A2(n14165), .ZN(n14208) );
  OR2_X1 U14155 ( .A1(n14209), .A2(n14210), .ZN(n14165) );
  AND2_X1 U14156 ( .A1(n14162), .A2(n14161), .ZN(n14210) );
  AND2_X1 U14157 ( .A1(n14159), .A2(n14211), .ZN(n14209) );
  OR2_X1 U14158 ( .A1(n14162), .A2(n14161), .ZN(n14211) );
  OR2_X1 U14159 ( .A1(n14212), .A2(n14213), .ZN(n14161) );
  AND2_X1 U14160 ( .A1(n14158), .A2(n14157), .ZN(n14213) );
  AND2_X1 U14161 ( .A1(n14155), .A2(n14214), .ZN(n14212) );
  OR2_X1 U14162 ( .A1(n14158), .A2(n14157), .ZN(n14214) );
  OR2_X1 U14163 ( .A1(n14215), .A2(n14216), .ZN(n14157) );
  AND2_X1 U14164 ( .A1(n14154), .A2(n14153), .ZN(n14216) );
  AND2_X1 U14165 ( .A1(n14151), .A2(n14217), .ZN(n14215) );
  OR2_X1 U14166 ( .A1(n14154), .A2(n14153), .ZN(n14217) );
  OR2_X1 U14167 ( .A1(n14218), .A2(n14219), .ZN(n14153) );
  AND2_X1 U14168 ( .A1(n14150), .A2(n14149), .ZN(n14219) );
  AND2_X1 U14169 ( .A1(n14147), .A2(n14220), .ZN(n14218) );
  OR2_X1 U14170 ( .A1(n14150), .A2(n14149), .ZN(n14220) );
  OR2_X1 U14171 ( .A1(n14221), .A2(n14222), .ZN(n14149) );
  AND2_X1 U14172 ( .A1(n8567), .A2(n14146), .ZN(n14222) );
  AND2_X1 U14173 ( .A1(n14144), .A2(n14223), .ZN(n14221) );
  OR2_X1 U14174 ( .A1(n8567), .A2(n14146), .ZN(n14223) );
  OR2_X1 U14175 ( .A1(n14224), .A2(n14225), .ZN(n14146) );
  AND2_X1 U14176 ( .A1(n14143), .A2(n14142), .ZN(n14225) );
  AND2_X1 U14177 ( .A1(n14140), .A2(n14226), .ZN(n14224) );
  OR2_X1 U14178 ( .A1(n14143), .A2(n14142), .ZN(n14226) );
  OR2_X1 U14179 ( .A1(n14227), .A2(n14228), .ZN(n14142) );
  AND2_X1 U14180 ( .A1(n14139), .A2(n14138), .ZN(n14228) );
  AND2_X1 U14181 ( .A1(n14136), .A2(n14229), .ZN(n14227) );
  OR2_X1 U14182 ( .A1(n14139), .A2(n14138), .ZN(n14229) );
  OR2_X1 U14183 ( .A1(n14230), .A2(n14231), .ZN(n14138) );
  AND2_X1 U14184 ( .A1(n14135), .A2(n14134), .ZN(n14231) );
  AND2_X1 U14185 ( .A1(n14132), .A2(n14232), .ZN(n14230) );
  OR2_X1 U14186 ( .A1(n14135), .A2(n14134), .ZN(n14232) );
  OR2_X1 U14187 ( .A1(n14233), .A2(n14234), .ZN(n14134) );
  AND2_X1 U14188 ( .A1(n14131), .A2(n14130), .ZN(n14234) );
  AND2_X1 U14189 ( .A1(n14128), .A2(n14235), .ZN(n14233) );
  OR2_X1 U14190 ( .A1(n14131), .A2(n14130), .ZN(n14235) );
  OR2_X1 U14191 ( .A1(n14236), .A2(n14237), .ZN(n14130) );
  AND2_X1 U14192 ( .A1(n14127), .A2(n14126), .ZN(n14237) );
  AND2_X1 U14193 ( .A1(n14124), .A2(n14238), .ZN(n14236) );
  OR2_X1 U14194 ( .A1(n14127), .A2(n14126), .ZN(n14238) );
  OR2_X1 U14195 ( .A1(n14239), .A2(n14240), .ZN(n14126) );
  AND2_X1 U14196 ( .A1(n14123), .A2(n14122), .ZN(n14240) );
  AND2_X1 U14197 ( .A1(n14120), .A2(n14241), .ZN(n14239) );
  OR2_X1 U14198 ( .A1(n14123), .A2(n14122), .ZN(n14241) );
  OR2_X1 U14199 ( .A1(n14242), .A2(n14243), .ZN(n14122) );
  AND2_X1 U14200 ( .A1(n14119), .A2(n14118), .ZN(n14243) );
  AND2_X1 U14201 ( .A1(n14116), .A2(n14244), .ZN(n14242) );
  OR2_X1 U14202 ( .A1(n14119), .A2(n14118), .ZN(n14244) );
  OR2_X1 U14203 ( .A1(n14245), .A2(n14246), .ZN(n14118) );
  AND2_X1 U14204 ( .A1(n14115), .A2(n14114), .ZN(n14246) );
  AND2_X1 U14205 ( .A1(n14112), .A2(n14247), .ZN(n14245) );
  OR2_X1 U14206 ( .A1(n14115), .A2(n14114), .ZN(n14247) );
  OR2_X1 U14207 ( .A1(n14248), .A2(n14249), .ZN(n14114) );
  AND2_X1 U14208 ( .A1(n14111), .A2(n14110), .ZN(n14249) );
  AND2_X1 U14209 ( .A1(n14108), .A2(n14250), .ZN(n14248) );
  OR2_X1 U14210 ( .A1(n14111), .A2(n14110), .ZN(n14250) );
  OR2_X1 U14211 ( .A1(n14251), .A2(n14252), .ZN(n14110) );
  AND2_X1 U14212 ( .A1(n14107), .A2(n14106), .ZN(n14252) );
  AND2_X1 U14213 ( .A1(n14104), .A2(n14253), .ZN(n14251) );
  OR2_X1 U14214 ( .A1(n14107), .A2(n14106), .ZN(n14253) );
  OR2_X1 U14215 ( .A1(n14254), .A2(n14255), .ZN(n14106) );
  AND2_X1 U14216 ( .A1(n14103), .A2(n14102), .ZN(n14255) );
  AND2_X1 U14217 ( .A1(n14100), .A2(n14256), .ZN(n14254) );
  OR2_X1 U14218 ( .A1(n14103), .A2(n14102), .ZN(n14256) );
  OR2_X1 U14219 ( .A1(n14257), .A2(n14258), .ZN(n14102) );
  AND2_X1 U14220 ( .A1(n14099), .A2(n14098), .ZN(n14258) );
  AND2_X1 U14221 ( .A1(n14096), .A2(n14259), .ZN(n14257) );
  OR2_X1 U14222 ( .A1(n14099), .A2(n14098), .ZN(n14259) );
  OR2_X1 U14223 ( .A1(n14260), .A2(n14261), .ZN(n14098) );
  AND2_X1 U14224 ( .A1(n14095), .A2(n14094), .ZN(n14261) );
  AND2_X1 U14225 ( .A1(n14092), .A2(n14262), .ZN(n14260) );
  OR2_X1 U14226 ( .A1(n14095), .A2(n14094), .ZN(n14262) );
  OR2_X1 U14227 ( .A1(n14263), .A2(n14264), .ZN(n14094) );
  AND2_X1 U14228 ( .A1(n14091), .A2(n14090), .ZN(n14264) );
  AND2_X1 U14229 ( .A1(n14088), .A2(n14265), .ZN(n14263) );
  OR2_X1 U14230 ( .A1(n14091), .A2(n14090), .ZN(n14265) );
  OR2_X1 U14231 ( .A1(n14266), .A2(n14267), .ZN(n14090) );
  AND2_X1 U14232 ( .A1(n14087), .A2(n14086), .ZN(n14267) );
  AND2_X1 U14233 ( .A1(n14084), .A2(n14268), .ZN(n14266) );
  OR2_X1 U14234 ( .A1(n14087), .A2(n14086), .ZN(n14268) );
  OR2_X1 U14235 ( .A1(n14269), .A2(n14270), .ZN(n14086) );
  AND2_X1 U14236 ( .A1(n14083), .A2(n14082), .ZN(n14270) );
  AND2_X1 U14237 ( .A1(n14080), .A2(n14271), .ZN(n14269) );
  OR2_X1 U14238 ( .A1(n14083), .A2(n14082), .ZN(n14271) );
  OR2_X1 U14239 ( .A1(n14272), .A2(n14273), .ZN(n14082) );
  AND2_X1 U14240 ( .A1(n14079), .A2(n14078), .ZN(n14273) );
  AND2_X1 U14241 ( .A1(n14076), .A2(n14274), .ZN(n14272) );
  OR2_X1 U14242 ( .A1(n14079), .A2(n14078), .ZN(n14274) );
  OR2_X1 U14243 ( .A1(n14275), .A2(n14276), .ZN(n14078) );
  AND2_X1 U14244 ( .A1(n14073), .A2(n14074), .ZN(n14276) );
  AND2_X1 U14245 ( .A1(n14277), .A2(n14278), .ZN(n14275) );
  OR2_X1 U14246 ( .A1(n14073), .A2(n14074), .ZN(n14278) );
  OR2_X1 U14247 ( .A1(n9984), .A2(n14279), .ZN(n14074) );
  OR2_X1 U14248 ( .A1(n8943), .A2(n8939), .ZN(n14279) );
  OR2_X1 U14249 ( .A1(n9014), .A2(n8943), .ZN(n14073) );
  INV_X1 U14250 ( .A(n14075), .ZN(n14277) );
  OR2_X1 U14251 ( .A1(n14280), .A2(n14281), .ZN(n14075) );
  AND2_X1 U14252 ( .A1(b_9_), .A2(n14282), .ZN(n14281) );
  OR2_X1 U14253 ( .A1(n14283), .A2(n8021), .ZN(n14282) );
  AND2_X1 U14254 ( .A1(a_31_), .A2(n8939), .ZN(n14283) );
  AND2_X1 U14255 ( .A1(b_10_), .A2(n14284), .ZN(n14280) );
  OR2_X1 U14256 ( .A1(n14285), .A2(n9989), .ZN(n14284) );
  AND2_X1 U14257 ( .A1(a_30_), .A2(n8935), .ZN(n14285) );
  OR2_X1 U14258 ( .A1(n9010), .A2(n8943), .ZN(n14079) );
  XOR2_X1 U14259 ( .A(n14286), .B(n14287), .Z(n14076) );
  XNOR2_X1 U14260 ( .A(n14288), .B(n14289), .ZN(n14286) );
  OR2_X1 U14261 ( .A1(n9006), .A2(n8943), .ZN(n14083) );
  XOR2_X1 U14262 ( .A(n14290), .B(n14291), .Z(n14080) );
  XOR2_X1 U14263 ( .A(n14292), .B(n14293), .Z(n14291) );
  OR2_X1 U14264 ( .A1(n9002), .A2(n8943), .ZN(n14087) );
  XNOR2_X1 U14265 ( .A(n14294), .B(n14295), .ZN(n14084) );
  XNOR2_X1 U14266 ( .A(n14296), .B(n14297), .ZN(n14294) );
  OR2_X1 U14267 ( .A1(n8998), .A2(n8943), .ZN(n14091) );
  XOR2_X1 U14268 ( .A(n14298), .B(n14299), .Z(n14088) );
  XOR2_X1 U14269 ( .A(n14300), .B(n14301), .Z(n14299) );
  OR2_X1 U14270 ( .A1(n8994), .A2(n8943), .ZN(n14095) );
  XOR2_X1 U14271 ( .A(n14302), .B(n14303), .Z(n14092) );
  XOR2_X1 U14272 ( .A(n14304), .B(n14305), .Z(n14303) );
  OR2_X1 U14273 ( .A1(n8990), .A2(n8943), .ZN(n14099) );
  XOR2_X1 U14274 ( .A(n14306), .B(n14307), .Z(n14096) );
  XOR2_X1 U14275 ( .A(n14308), .B(n14309), .Z(n14307) );
  OR2_X1 U14276 ( .A1(n8986), .A2(n8943), .ZN(n14103) );
  XOR2_X1 U14277 ( .A(n14310), .B(n14311), .Z(n14100) );
  XOR2_X1 U14278 ( .A(n14312), .B(n14313), .Z(n14311) );
  OR2_X1 U14279 ( .A1(n8982), .A2(n8943), .ZN(n14107) );
  XOR2_X1 U14280 ( .A(n14314), .B(n14315), .Z(n14104) );
  XOR2_X1 U14281 ( .A(n14316), .B(n14317), .Z(n14315) );
  OR2_X1 U14282 ( .A1(n8978), .A2(n8943), .ZN(n14111) );
  XOR2_X1 U14283 ( .A(n14318), .B(n14319), .Z(n14108) );
  XOR2_X1 U14284 ( .A(n14320), .B(n14321), .Z(n14319) );
  OR2_X1 U14285 ( .A1(n8974), .A2(n8943), .ZN(n14115) );
  XOR2_X1 U14286 ( .A(n14322), .B(n14323), .Z(n14112) );
  XOR2_X1 U14287 ( .A(n14324), .B(n14325), .Z(n14323) );
  OR2_X1 U14288 ( .A1(n8970), .A2(n8943), .ZN(n14119) );
  XOR2_X1 U14289 ( .A(n14326), .B(n14327), .Z(n14116) );
  XOR2_X1 U14290 ( .A(n14328), .B(n14329), .Z(n14327) );
  OR2_X1 U14291 ( .A1(n8966), .A2(n8943), .ZN(n14123) );
  XOR2_X1 U14292 ( .A(n14330), .B(n14331), .Z(n14120) );
  XOR2_X1 U14293 ( .A(n14332), .B(n14333), .Z(n14331) );
  OR2_X1 U14294 ( .A1(n8962), .A2(n8943), .ZN(n14127) );
  XOR2_X1 U14295 ( .A(n14334), .B(n14335), .Z(n14124) );
  XOR2_X1 U14296 ( .A(n14336), .B(n14337), .Z(n14335) );
  OR2_X1 U14297 ( .A1(n8958), .A2(n8943), .ZN(n14131) );
  XOR2_X1 U14298 ( .A(n14338), .B(n14339), .Z(n14128) );
  XOR2_X1 U14299 ( .A(n14340), .B(n14341), .Z(n14339) );
  OR2_X1 U14300 ( .A1(n8954), .A2(n8943), .ZN(n14135) );
  XOR2_X1 U14301 ( .A(n14342), .B(n14343), .Z(n14132) );
  XOR2_X1 U14302 ( .A(n14344), .B(n14345), .Z(n14343) );
  OR2_X1 U14303 ( .A1(n8950), .A2(n8943), .ZN(n14139) );
  XOR2_X1 U14304 ( .A(n14346), .B(n14347), .Z(n14136) );
  XOR2_X1 U14305 ( .A(n14348), .B(n14349), .Z(n14347) );
  OR2_X1 U14306 ( .A1(n8946), .A2(n8943), .ZN(n14143) );
  XOR2_X1 U14307 ( .A(n14350), .B(n14351), .Z(n14140) );
  XOR2_X1 U14308 ( .A(n14352), .B(n14353), .Z(n14351) );
  OR2_X1 U14309 ( .A1(n8942), .A2(n8943), .ZN(n8567) );
  XOR2_X1 U14310 ( .A(n14354), .B(n14355), .Z(n14144) );
  XOR2_X1 U14311 ( .A(n14356), .B(n14357), .Z(n14355) );
  OR2_X1 U14312 ( .A1(n8938), .A2(n8943), .ZN(n14150) );
  XOR2_X1 U14313 ( .A(n14358), .B(n14359), .Z(n14147) );
  XOR2_X1 U14314 ( .A(n14360), .B(n14361), .Z(n14359) );
  OR2_X1 U14315 ( .A1(n8934), .A2(n8943), .ZN(n14154) );
  XOR2_X1 U14316 ( .A(n14362), .B(n14363), .Z(n14151) );
  XOR2_X1 U14317 ( .A(n14364), .B(n8596), .Z(n14363) );
  OR2_X1 U14318 ( .A1(n8930), .A2(n8943), .ZN(n14158) );
  XOR2_X1 U14319 ( .A(n14365), .B(n14366), .Z(n14155) );
  XOR2_X1 U14320 ( .A(n14367), .B(n14368), .Z(n14366) );
  OR2_X1 U14321 ( .A1(n8926), .A2(n8943), .ZN(n14162) );
  XOR2_X1 U14322 ( .A(n14369), .B(n14370), .Z(n14159) );
  XOR2_X1 U14323 ( .A(n14371), .B(n14372), .Z(n14370) );
  OR2_X1 U14324 ( .A1(n8922), .A2(n8943), .ZN(n14166) );
  XOR2_X1 U14325 ( .A(n14373), .B(n14374), .Z(n14163) );
  XOR2_X1 U14326 ( .A(n14375), .B(n14376), .Z(n14374) );
  OR2_X1 U14327 ( .A1(n8918), .A2(n8943), .ZN(n14170) );
  XOR2_X1 U14328 ( .A(n14377), .B(n14378), .Z(n14167) );
  XOR2_X1 U14329 ( .A(n14379), .B(n14380), .Z(n14378) );
  OR2_X1 U14330 ( .A1(n8914), .A2(n8943), .ZN(n14174) );
  XOR2_X1 U14331 ( .A(n14381), .B(n14382), .Z(n14171) );
  XOR2_X1 U14332 ( .A(n14383), .B(n14384), .Z(n14382) );
  OR2_X1 U14333 ( .A1(n8910), .A2(n8943), .ZN(n14178) );
  XOR2_X1 U14334 ( .A(n14385), .B(n14386), .Z(n14175) );
  XOR2_X1 U14335 ( .A(n14387), .B(n14388), .Z(n14386) );
  OR2_X1 U14336 ( .A1(n8906), .A2(n8943), .ZN(n14182) );
  XOR2_X1 U14337 ( .A(n14389), .B(n14390), .Z(n14179) );
  XOR2_X1 U14338 ( .A(n14391), .B(n14392), .Z(n14390) );
  OR2_X1 U14339 ( .A1(n8902), .A2(n8943), .ZN(n14186) );
  XOR2_X1 U14340 ( .A(n14393), .B(n14394), .Z(n14183) );
  XOR2_X1 U14341 ( .A(n14395), .B(n14396), .Z(n14394) );
  OR2_X1 U14342 ( .A1(n9297), .A2(n8943), .ZN(n9730) );
  XOR2_X1 U14343 ( .A(n14397), .B(n14398), .Z(n9727) );
  XOR2_X1 U14344 ( .A(n14399), .B(n14400), .Z(n14398) );
  XOR2_X1 U14345 ( .A(n9657), .B(n14401), .Z(n9719) );
  XOR2_X1 U14346 ( .A(n9656), .B(n9655), .Z(n14401) );
  OR2_X1 U14347 ( .A1(n9297), .A2(n8939), .ZN(n9655) );
  OR2_X1 U14348 ( .A1(n14402), .A2(n14403), .ZN(n9656) );
  AND2_X1 U14349 ( .A1(n14400), .A2(n14399), .ZN(n14403) );
  AND2_X1 U14350 ( .A1(n14397), .A2(n14404), .ZN(n14402) );
  OR2_X1 U14351 ( .A1(n14399), .A2(n14400), .ZN(n14404) );
  OR2_X1 U14352 ( .A1(n8902), .A2(n8939), .ZN(n14400) );
  OR2_X1 U14353 ( .A1(n14405), .A2(n14406), .ZN(n14399) );
  AND2_X1 U14354 ( .A1(n14396), .A2(n14395), .ZN(n14406) );
  AND2_X1 U14355 ( .A1(n14393), .A2(n14407), .ZN(n14405) );
  OR2_X1 U14356 ( .A1(n14395), .A2(n14396), .ZN(n14407) );
  OR2_X1 U14357 ( .A1(n8906), .A2(n8939), .ZN(n14396) );
  OR2_X1 U14358 ( .A1(n14408), .A2(n14409), .ZN(n14395) );
  AND2_X1 U14359 ( .A1(n14392), .A2(n14391), .ZN(n14409) );
  AND2_X1 U14360 ( .A1(n14389), .A2(n14410), .ZN(n14408) );
  OR2_X1 U14361 ( .A1(n14391), .A2(n14392), .ZN(n14410) );
  OR2_X1 U14362 ( .A1(n8910), .A2(n8939), .ZN(n14392) );
  OR2_X1 U14363 ( .A1(n14411), .A2(n14412), .ZN(n14391) );
  AND2_X1 U14364 ( .A1(n14388), .A2(n14387), .ZN(n14412) );
  AND2_X1 U14365 ( .A1(n14385), .A2(n14413), .ZN(n14411) );
  OR2_X1 U14366 ( .A1(n14387), .A2(n14388), .ZN(n14413) );
  OR2_X1 U14367 ( .A1(n8914), .A2(n8939), .ZN(n14388) );
  OR2_X1 U14368 ( .A1(n14414), .A2(n14415), .ZN(n14387) );
  AND2_X1 U14369 ( .A1(n14384), .A2(n14383), .ZN(n14415) );
  AND2_X1 U14370 ( .A1(n14381), .A2(n14416), .ZN(n14414) );
  OR2_X1 U14371 ( .A1(n14383), .A2(n14384), .ZN(n14416) );
  OR2_X1 U14372 ( .A1(n8918), .A2(n8939), .ZN(n14384) );
  OR2_X1 U14373 ( .A1(n14417), .A2(n14418), .ZN(n14383) );
  AND2_X1 U14374 ( .A1(n14380), .A2(n14379), .ZN(n14418) );
  AND2_X1 U14375 ( .A1(n14377), .A2(n14419), .ZN(n14417) );
  OR2_X1 U14376 ( .A1(n14379), .A2(n14380), .ZN(n14419) );
  OR2_X1 U14377 ( .A1(n8922), .A2(n8939), .ZN(n14380) );
  OR2_X1 U14378 ( .A1(n14420), .A2(n14421), .ZN(n14379) );
  AND2_X1 U14379 ( .A1(n14376), .A2(n14375), .ZN(n14421) );
  AND2_X1 U14380 ( .A1(n14373), .A2(n14422), .ZN(n14420) );
  OR2_X1 U14381 ( .A1(n14375), .A2(n14376), .ZN(n14422) );
  OR2_X1 U14382 ( .A1(n8926), .A2(n8939), .ZN(n14376) );
  OR2_X1 U14383 ( .A1(n14423), .A2(n14424), .ZN(n14375) );
  AND2_X1 U14384 ( .A1(n14372), .A2(n14371), .ZN(n14424) );
  AND2_X1 U14385 ( .A1(n14369), .A2(n14425), .ZN(n14423) );
  OR2_X1 U14386 ( .A1(n14371), .A2(n14372), .ZN(n14425) );
  OR2_X1 U14387 ( .A1(n8930), .A2(n8939), .ZN(n14372) );
  OR2_X1 U14388 ( .A1(n14426), .A2(n14427), .ZN(n14371) );
  AND2_X1 U14389 ( .A1(n14368), .A2(n14367), .ZN(n14427) );
  AND2_X1 U14390 ( .A1(n14365), .A2(n14428), .ZN(n14426) );
  OR2_X1 U14391 ( .A1(n14367), .A2(n14368), .ZN(n14428) );
  OR2_X1 U14392 ( .A1(n8934), .A2(n8939), .ZN(n14368) );
  OR2_X1 U14393 ( .A1(n14429), .A2(n14430), .ZN(n14367) );
  AND2_X1 U14394 ( .A1(n8596), .A2(n14364), .ZN(n14430) );
  AND2_X1 U14395 ( .A1(n14362), .A2(n14431), .ZN(n14429) );
  OR2_X1 U14396 ( .A1(n14364), .A2(n8596), .ZN(n14431) );
  OR2_X1 U14397 ( .A1(n8938), .A2(n8939), .ZN(n8596) );
  OR2_X1 U14398 ( .A1(n14432), .A2(n14433), .ZN(n14364) );
  AND2_X1 U14399 ( .A1(n14361), .A2(n14360), .ZN(n14433) );
  AND2_X1 U14400 ( .A1(n14358), .A2(n14434), .ZN(n14432) );
  OR2_X1 U14401 ( .A1(n14360), .A2(n14361), .ZN(n14434) );
  OR2_X1 U14402 ( .A1(n8942), .A2(n8939), .ZN(n14361) );
  OR2_X1 U14403 ( .A1(n14435), .A2(n14436), .ZN(n14360) );
  AND2_X1 U14404 ( .A1(n14357), .A2(n14356), .ZN(n14436) );
  AND2_X1 U14405 ( .A1(n14354), .A2(n14437), .ZN(n14435) );
  OR2_X1 U14406 ( .A1(n14356), .A2(n14357), .ZN(n14437) );
  OR2_X1 U14407 ( .A1(n8946), .A2(n8939), .ZN(n14357) );
  OR2_X1 U14408 ( .A1(n14438), .A2(n14439), .ZN(n14356) );
  AND2_X1 U14409 ( .A1(n14353), .A2(n14352), .ZN(n14439) );
  AND2_X1 U14410 ( .A1(n14350), .A2(n14440), .ZN(n14438) );
  OR2_X1 U14411 ( .A1(n14352), .A2(n14353), .ZN(n14440) );
  OR2_X1 U14412 ( .A1(n8950), .A2(n8939), .ZN(n14353) );
  OR2_X1 U14413 ( .A1(n14441), .A2(n14442), .ZN(n14352) );
  AND2_X1 U14414 ( .A1(n14349), .A2(n14348), .ZN(n14442) );
  AND2_X1 U14415 ( .A1(n14346), .A2(n14443), .ZN(n14441) );
  OR2_X1 U14416 ( .A1(n14348), .A2(n14349), .ZN(n14443) );
  OR2_X1 U14417 ( .A1(n8954), .A2(n8939), .ZN(n14349) );
  OR2_X1 U14418 ( .A1(n14444), .A2(n14445), .ZN(n14348) );
  AND2_X1 U14419 ( .A1(n14345), .A2(n14344), .ZN(n14445) );
  AND2_X1 U14420 ( .A1(n14342), .A2(n14446), .ZN(n14444) );
  OR2_X1 U14421 ( .A1(n14344), .A2(n14345), .ZN(n14446) );
  OR2_X1 U14422 ( .A1(n8958), .A2(n8939), .ZN(n14345) );
  OR2_X1 U14423 ( .A1(n14447), .A2(n14448), .ZN(n14344) );
  AND2_X1 U14424 ( .A1(n14341), .A2(n14340), .ZN(n14448) );
  AND2_X1 U14425 ( .A1(n14338), .A2(n14449), .ZN(n14447) );
  OR2_X1 U14426 ( .A1(n14340), .A2(n14341), .ZN(n14449) );
  OR2_X1 U14427 ( .A1(n8962), .A2(n8939), .ZN(n14341) );
  OR2_X1 U14428 ( .A1(n14450), .A2(n14451), .ZN(n14340) );
  AND2_X1 U14429 ( .A1(n14337), .A2(n14336), .ZN(n14451) );
  AND2_X1 U14430 ( .A1(n14334), .A2(n14452), .ZN(n14450) );
  OR2_X1 U14431 ( .A1(n14336), .A2(n14337), .ZN(n14452) );
  OR2_X1 U14432 ( .A1(n8966), .A2(n8939), .ZN(n14337) );
  OR2_X1 U14433 ( .A1(n14453), .A2(n14454), .ZN(n14336) );
  AND2_X1 U14434 ( .A1(n14333), .A2(n14332), .ZN(n14454) );
  AND2_X1 U14435 ( .A1(n14330), .A2(n14455), .ZN(n14453) );
  OR2_X1 U14436 ( .A1(n14332), .A2(n14333), .ZN(n14455) );
  OR2_X1 U14437 ( .A1(n8970), .A2(n8939), .ZN(n14333) );
  OR2_X1 U14438 ( .A1(n14456), .A2(n14457), .ZN(n14332) );
  AND2_X1 U14439 ( .A1(n14326), .A2(n14329), .ZN(n14457) );
  AND2_X1 U14440 ( .A1(n14458), .A2(n14328), .ZN(n14456) );
  OR2_X1 U14441 ( .A1(n14459), .A2(n14460), .ZN(n14328) );
  AND2_X1 U14442 ( .A1(n14325), .A2(n14324), .ZN(n14460) );
  AND2_X1 U14443 ( .A1(n14322), .A2(n14461), .ZN(n14459) );
  OR2_X1 U14444 ( .A1(n14324), .A2(n14325), .ZN(n14461) );
  OR2_X1 U14445 ( .A1(n8978), .A2(n8939), .ZN(n14325) );
  OR2_X1 U14446 ( .A1(n14462), .A2(n14463), .ZN(n14324) );
  AND2_X1 U14447 ( .A1(n14318), .A2(n14321), .ZN(n14463) );
  AND2_X1 U14448 ( .A1(n14464), .A2(n14320), .ZN(n14462) );
  OR2_X1 U14449 ( .A1(n14465), .A2(n14466), .ZN(n14320) );
  AND2_X1 U14450 ( .A1(n14314), .A2(n14317), .ZN(n14466) );
  AND2_X1 U14451 ( .A1(n14467), .A2(n14316), .ZN(n14465) );
  OR2_X1 U14452 ( .A1(n14468), .A2(n14469), .ZN(n14316) );
  AND2_X1 U14453 ( .A1(n14310), .A2(n14313), .ZN(n14469) );
  AND2_X1 U14454 ( .A1(n14470), .A2(n14312), .ZN(n14468) );
  OR2_X1 U14455 ( .A1(n14471), .A2(n14472), .ZN(n14312) );
  AND2_X1 U14456 ( .A1(n14306), .A2(n14309), .ZN(n14472) );
  AND2_X1 U14457 ( .A1(n14473), .A2(n14308), .ZN(n14471) );
  OR2_X1 U14458 ( .A1(n14474), .A2(n14475), .ZN(n14308) );
  AND2_X1 U14459 ( .A1(n14302), .A2(n14305), .ZN(n14475) );
  AND2_X1 U14460 ( .A1(n14476), .A2(n14304), .ZN(n14474) );
  OR2_X1 U14461 ( .A1(n14477), .A2(n14478), .ZN(n14304) );
  AND2_X1 U14462 ( .A1(n14298), .A2(n14301), .ZN(n14478) );
  AND2_X1 U14463 ( .A1(n14479), .A2(n14300), .ZN(n14477) );
  OR2_X1 U14464 ( .A1(n14480), .A2(n14481), .ZN(n14300) );
  AND2_X1 U14465 ( .A1(n14295), .A2(n14296), .ZN(n14481) );
  AND2_X1 U14466 ( .A1(n14482), .A2(n14297), .ZN(n14480) );
  OR2_X1 U14467 ( .A1(n14483), .A2(n14484), .ZN(n14297) );
  AND2_X1 U14468 ( .A1(n14290), .A2(n14293), .ZN(n14484) );
  AND2_X1 U14469 ( .A1(n14485), .A2(n14292), .ZN(n14483) );
  OR2_X1 U14470 ( .A1(n14486), .A2(n14487), .ZN(n14292) );
  AND2_X1 U14471 ( .A1(n14287), .A2(n14288), .ZN(n14487) );
  AND2_X1 U14472 ( .A1(n14488), .A2(n14489), .ZN(n14486) );
  OR2_X1 U14473 ( .A1(n14288), .A2(n14287), .ZN(n14489) );
  OR2_X1 U14474 ( .A1(n9014), .A2(n8939), .ZN(n14287) );
  OR2_X1 U14475 ( .A1(n9984), .A2(n14490), .ZN(n14288) );
  OR2_X1 U14476 ( .A1(n8939), .A2(n8935), .ZN(n14490) );
  INV_X1 U14477 ( .A(n14289), .ZN(n14488) );
  OR2_X1 U14478 ( .A1(n14491), .A2(n14492), .ZN(n14289) );
  AND2_X1 U14479 ( .A1(b_9_), .A2(n14493), .ZN(n14492) );
  OR2_X1 U14480 ( .A1(n14494), .A2(n9989), .ZN(n14493) );
  AND2_X1 U14481 ( .A1(a_30_), .A2(n8931), .ZN(n14494) );
  AND2_X1 U14482 ( .A1(b_8_), .A2(n14495), .ZN(n14491) );
  OR2_X1 U14483 ( .A1(n14496), .A2(n8021), .ZN(n14495) );
  AND2_X1 U14484 ( .A1(a_31_), .A2(n8935), .ZN(n14496) );
  OR2_X1 U14485 ( .A1(n14293), .A2(n14290), .ZN(n14485) );
  XOR2_X1 U14486 ( .A(n14497), .B(n14498), .Z(n14290) );
  XNOR2_X1 U14487 ( .A(n14499), .B(n14500), .ZN(n14497) );
  OR2_X1 U14488 ( .A1(n9010), .A2(n8939), .ZN(n14293) );
  OR2_X1 U14489 ( .A1(n14296), .A2(n14295), .ZN(n14482) );
  XOR2_X1 U14490 ( .A(n14501), .B(n14502), .Z(n14295) );
  XOR2_X1 U14491 ( .A(n14503), .B(n14504), .Z(n14502) );
  OR2_X1 U14492 ( .A1(n9006), .A2(n8939), .ZN(n14296) );
  OR2_X1 U14493 ( .A1(n14301), .A2(n14298), .ZN(n14479) );
  XNOR2_X1 U14494 ( .A(n14505), .B(n14506), .ZN(n14298) );
  XNOR2_X1 U14495 ( .A(n14507), .B(n14508), .ZN(n14505) );
  OR2_X1 U14496 ( .A1(n9002), .A2(n8939), .ZN(n14301) );
  OR2_X1 U14497 ( .A1(n14305), .A2(n14302), .ZN(n14476) );
  XOR2_X1 U14498 ( .A(n14509), .B(n14510), .Z(n14302) );
  XOR2_X1 U14499 ( .A(n14511), .B(n14512), .Z(n14510) );
  OR2_X1 U14500 ( .A1(n8998), .A2(n8939), .ZN(n14305) );
  OR2_X1 U14501 ( .A1(n14309), .A2(n14306), .ZN(n14473) );
  XOR2_X1 U14502 ( .A(n14513), .B(n14514), .Z(n14306) );
  XOR2_X1 U14503 ( .A(n14515), .B(n14516), .Z(n14514) );
  OR2_X1 U14504 ( .A1(n8994), .A2(n8939), .ZN(n14309) );
  OR2_X1 U14505 ( .A1(n14313), .A2(n14310), .ZN(n14470) );
  XOR2_X1 U14506 ( .A(n14517), .B(n14518), .Z(n14310) );
  XOR2_X1 U14507 ( .A(n14519), .B(n14520), .Z(n14518) );
  OR2_X1 U14508 ( .A1(n8990), .A2(n8939), .ZN(n14313) );
  OR2_X1 U14509 ( .A1(n14317), .A2(n14314), .ZN(n14467) );
  XOR2_X1 U14510 ( .A(n14521), .B(n14522), .Z(n14314) );
  XOR2_X1 U14511 ( .A(n14523), .B(n14524), .Z(n14522) );
  OR2_X1 U14512 ( .A1(n8986), .A2(n8939), .ZN(n14317) );
  OR2_X1 U14513 ( .A1(n14321), .A2(n14318), .ZN(n14464) );
  XOR2_X1 U14514 ( .A(n14525), .B(n14526), .Z(n14318) );
  XOR2_X1 U14515 ( .A(n14527), .B(n14528), .Z(n14526) );
  OR2_X1 U14516 ( .A1(n8982), .A2(n8939), .ZN(n14321) );
  XOR2_X1 U14517 ( .A(n14529), .B(n14530), .Z(n14322) );
  XOR2_X1 U14518 ( .A(n14531), .B(n14532), .Z(n14530) );
  OR2_X1 U14519 ( .A1(n14329), .A2(n14326), .ZN(n14458) );
  XOR2_X1 U14520 ( .A(n14533), .B(n14534), .Z(n14326) );
  XOR2_X1 U14521 ( .A(n14535), .B(n14536), .Z(n14534) );
  OR2_X1 U14522 ( .A1(n8974), .A2(n8939), .ZN(n14329) );
  XOR2_X1 U14523 ( .A(n14537), .B(n14538), .Z(n14330) );
  XOR2_X1 U14524 ( .A(n14539), .B(n14540), .Z(n14538) );
  XOR2_X1 U14525 ( .A(n14541), .B(n14542), .Z(n14334) );
  XOR2_X1 U14526 ( .A(n14543), .B(n14544), .Z(n14542) );
  XOR2_X1 U14527 ( .A(n14545), .B(n14546), .Z(n14338) );
  XOR2_X1 U14528 ( .A(n14547), .B(n14548), .Z(n14546) );
  XOR2_X1 U14529 ( .A(n14549), .B(n14550), .Z(n14342) );
  XOR2_X1 U14530 ( .A(n14551), .B(n14552), .Z(n14550) );
  XOR2_X1 U14531 ( .A(n14553), .B(n14554), .Z(n14346) );
  XOR2_X1 U14532 ( .A(n14555), .B(n14556), .Z(n14554) );
  XOR2_X1 U14533 ( .A(n14557), .B(n14558), .Z(n14350) );
  XOR2_X1 U14534 ( .A(n14559), .B(n14560), .Z(n14558) );
  XOR2_X1 U14535 ( .A(n14561), .B(n14562), .Z(n14354) );
  XOR2_X1 U14536 ( .A(n14563), .B(n14564), .Z(n14562) );
  XOR2_X1 U14537 ( .A(n14565), .B(n14566), .Z(n14358) );
  XOR2_X1 U14538 ( .A(n14567), .B(n14568), .Z(n14566) );
  XOR2_X1 U14539 ( .A(n14569), .B(n14570), .Z(n14362) );
  XOR2_X1 U14540 ( .A(n14571), .B(n14572), .Z(n14570) );
  XOR2_X1 U14541 ( .A(n14573), .B(n14574), .Z(n14365) );
  XOR2_X1 U14542 ( .A(n14575), .B(n14576), .Z(n14574) );
  XOR2_X1 U14543 ( .A(n14577), .B(n14578), .Z(n14369) );
  XOR2_X1 U14544 ( .A(n14579), .B(n8625), .Z(n14578) );
  XOR2_X1 U14545 ( .A(n14580), .B(n14581), .Z(n14373) );
  XOR2_X1 U14546 ( .A(n14582), .B(n14583), .Z(n14581) );
  XOR2_X1 U14547 ( .A(n14584), .B(n14585), .Z(n14377) );
  XOR2_X1 U14548 ( .A(n14586), .B(n14587), .Z(n14585) );
  XOR2_X1 U14549 ( .A(n14588), .B(n14589), .Z(n14381) );
  XOR2_X1 U14550 ( .A(n14590), .B(n14591), .Z(n14589) );
  XOR2_X1 U14551 ( .A(n14592), .B(n14593), .Z(n14385) );
  XOR2_X1 U14552 ( .A(n14594), .B(n14595), .Z(n14593) );
  XOR2_X1 U14553 ( .A(n14596), .B(n14597), .Z(n14389) );
  XOR2_X1 U14554 ( .A(n14598), .B(n14599), .Z(n14597) );
  XOR2_X1 U14555 ( .A(n14600), .B(n14601), .Z(n14393) );
  XOR2_X1 U14556 ( .A(n14602), .B(n14603), .Z(n14601) );
  XOR2_X1 U14557 ( .A(n14604), .B(n14605), .Z(n14397) );
  XOR2_X1 U14558 ( .A(n14606), .B(n14607), .Z(n14605) );
  XOR2_X1 U14559 ( .A(n9664), .B(n14608), .Z(n9657) );
  XOR2_X1 U14560 ( .A(n9663), .B(n9662), .Z(n14608) );
  OR2_X1 U14561 ( .A1(n8902), .A2(n8935), .ZN(n9662) );
  OR2_X1 U14562 ( .A1(n14609), .A2(n14610), .ZN(n9663) );
  AND2_X1 U14563 ( .A1(n14607), .A2(n14606), .ZN(n14610) );
  AND2_X1 U14564 ( .A1(n14604), .A2(n14611), .ZN(n14609) );
  OR2_X1 U14565 ( .A1(n14606), .A2(n14607), .ZN(n14611) );
  OR2_X1 U14566 ( .A1(n8906), .A2(n8935), .ZN(n14607) );
  OR2_X1 U14567 ( .A1(n14612), .A2(n14613), .ZN(n14606) );
  AND2_X1 U14568 ( .A1(n14603), .A2(n14602), .ZN(n14613) );
  AND2_X1 U14569 ( .A1(n14600), .A2(n14614), .ZN(n14612) );
  OR2_X1 U14570 ( .A1(n14602), .A2(n14603), .ZN(n14614) );
  OR2_X1 U14571 ( .A1(n8910), .A2(n8935), .ZN(n14603) );
  OR2_X1 U14572 ( .A1(n14615), .A2(n14616), .ZN(n14602) );
  AND2_X1 U14573 ( .A1(n14599), .A2(n14598), .ZN(n14616) );
  AND2_X1 U14574 ( .A1(n14596), .A2(n14617), .ZN(n14615) );
  OR2_X1 U14575 ( .A1(n14598), .A2(n14599), .ZN(n14617) );
  OR2_X1 U14576 ( .A1(n8914), .A2(n8935), .ZN(n14599) );
  OR2_X1 U14577 ( .A1(n14618), .A2(n14619), .ZN(n14598) );
  AND2_X1 U14578 ( .A1(n14595), .A2(n14594), .ZN(n14619) );
  AND2_X1 U14579 ( .A1(n14592), .A2(n14620), .ZN(n14618) );
  OR2_X1 U14580 ( .A1(n14594), .A2(n14595), .ZN(n14620) );
  OR2_X1 U14581 ( .A1(n8918), .A2(n8935), .ZN(n14595) );
  OR2_X1 U14582 ( .A1(n14621), .A2(n14622), .ZN(n14594) );
  AND2_X1 U14583 ( .A1(n14591), .A2(n14590), .ZN(n14622) );
  AND2_X1 U14584 ( .A1(n14588), .A2(n14623), .ZN(n14621) );
  OR2_X1 U14585 ( .A1(n14590), .A2(n14591), .ZN(n14623) );
  OR2_X1 U14586 ( .A1(n8922), .A2(n8935), .ZN(n14591) );
  OR2_X1 U14587 ( .A1(n14624), .A2(n14625), .ZN(n14590) );
  AND2_X1 U14588 ( .A1(n14587), .A2(n14586), .ZN(n14625) );
  AND2_X1 U14589 ( .A1(n14584), .A2(n14626), .ZN(n14624) );
  OR2_X1 U14590 ( .A1(n14586), .A2(n14587), .ZN(n14626) );
  OR2_X1 U14591 ( .A1(n8926), .A2(n8935), .ZN(n14587) );
  OR2_X1 U14592 ( .A1(n14627), .A2(n14628), .ZN(n14586) );
  AND2_X1 U14593 ( .A1(n14583), .A2(n14582), .ZN(n14628) );
  AND2_X1 U14594 ( .A1(n14580), .A2(n14629), .ZN(n14627) );
  OR2_X1 U14595 ( .A1(n14582), .A2(n14583), .ZN(n14629) );
  OR2_X1 U14596 ( .A1(n8930), .A2(n8935), .ZN(n14583) );
  OR2_X1 U14597 ( .A1(n14630), .A2(n14631), .ZN(n14582) );
  AND2_X1 U14598 ( .A1(n8625), .A2(n14579), .ZN(n14631) );
  AND2_X1 U14599 ( .A1(n14577), .A2(n14632), .ZN(n14630) );
  OR2_X1 U14600 ( .A1(n14579), .A2(n8625), .ZN(n14632) );
  OR2_X1 U14601 ( .A1(n8934), .A2(n8935), .ZN(n8625) );
  OR2_X1 U14602 ( .A1(n14633), .A2(n14634), .ZN(n14579) );
  AND2_X1 U14603 ( .A1(n14576), .A2(n14575), .ZN(n14634) );
  AND2_X1 U14604 ( .A1(n14573), .A2(n14635), .ZN(n14633) );
  OR2_X1 U14605 ( .A1(n14575), .A2(n14576), .ZN(n14635) );
  OR2_X1 U14606 ( .A1(n8938), .A2(n8935), .ZN(n14576) );
  OR2_X1 U14607 ( .A1(n14636), .A2(n14637), .ZN(n14575) );
  AND2_X1 U14608 ( .A1(n14572), .A2(n14571), .ZN(n14637) );
  AND2_X1 U14609 ( .A1(n14569), .A2(n14638), .ZN(n14636) );
  OR2_X1 U14610 ( .A1(n14571), .A2(n14572), .ZN(n14638) );
  OR2_X1 U14611 ( .A1(n8942), .A2(n8935), .ZN(n14572) );
  OR2_X1 U14612 ( .A1(n14639), .A2(n14640), .ZN(n14571) );
  AND2_X1 U14613 ( .A1(n14568), .A2(n14567), .ZN(n14640) );
  AND2_X1 U14614 ( .A1(n14565), .A2(n14641), .ZN(n14639) );
  OR2_X1 U14615 ( .A1(n14567), .A2(n14568), .ZN(n14641) );
  OR2_X1 U14616 ( .A1(n8946), .A2(n8935), .ZN(n14568) );
  OR2_X1 U14617 ( .A1(n14642), .A2(n14643), .ZN(n14567) );
  AND2_X1 U14618 ( .A1(n14564), .A2(n14563), .ZN(n14643) );
  AND2_X1 U14619 ( .A1(n14561), .A2(n14644), .ZN(n14642) );
  OR2_X1 U14620 ( .A1(n14563), .A2(n14564), .ZN(n14644) );
  OR2_X1 U14621 ( .A1(n8950), .A2(n8935), .ZN(n14564) );
  OR2_X1 U14622 ( .A1(n14645), .A2(n14646), .ZN(n14563) );
  AND2_X1 U14623 ( .A1(n14560), .A2(n14559), .ZN(n14646) );
  AND2_X1 U14624 ( .A1(n14557), .A2(n14647), .ZN(n14645) );
  OR2_X1 U14625 ( .A1(n14559), .A2(n14560), .ZN(n14647) );
  OR2_X1 U14626 ( .A1(n8954), .A2(n8935), .ZN(n14560) );
  OR2_X1 U14627 ( .A1(n14648), .A2(n14649), .ZN(n14559) );
  AND2_X1 U14628 ( .A1(n14556), .A2(n14555), .ZN(n14649) );
  AND2_X1 U14629 ( .A1(n14553), .A2(n14650), .ZN(n14648) );
  OR2_X1 U14630 ( .A1(n14555), .A2(n14556), .ZN(n14650) );
  OR2_X1 U14631 ( .A1(n8958), .A2(n8935), .ZN(n14556) );
  OR2_X1 U14632 ( .A1(n14651), .A2(n14652), .ZN(n14555) );
  AND2_X1 U14633 ( .A1(n14552), .A2(n14551), .ZN(n14652) );
  AND2_X1 U14634 ( .A1(n14549), .A2(n14653), .ZN(n14651) );
  OR2_X1 U14635 ( .A1(n14551), .A2(n14552), .ZN(n14653) );
  OR2_X1 U14636 ( .A1(n8962), .A2(n8935), .ZN(n14552) );
  OR2_X1 U14637 ( .A1(n14654), .A2(n14655), .ZN(n14551) );
  AND2_X1 U14638 ( .A1(n14548), .A2(n14547), .ZN(n14655) );
  AND2_X1 U14639 ( .A1(n14545), .A2(n14656), .ZN(n14654) );
  OR2_X1 U14640 ( .A1(n14547), .A2(n14548), .ZN(n14656) );
  OR2_X1 U14641 ( .A1(n8966), .A2(n8935), .ZN(n14548) );
  OR2_X1 U14642 ( .A1(n14657), .A2(n14658), .ZN(n14547) );
  AND2_X1 U14643 ( .A1(n14544), .A2(n14543), .ZN(n14658) );
  AND2_X1 U14644 ( .A1(n14541), .A2(n14659), .ZN(n14657) );
  OR2_X1 U14645 ( .A1(n14543), .A2(n14544), .ZN(n14659) );
  OR2_X1 U14646 ( .A1(n8970), .A2(n8935), .ZN(n14544) );
  OR2_X1 U14647 ( .A1(n14660), .A2(n14661), .ZN(n14543) );
  AND2_X1 U14648 ( .A1(n14540), .A2(n14539), .ZN(n14661) );
  AND2_X1 U14649 ( .A1(n14537), .A2(n14662), .ZN(n14660) );
  OR2_X1 U14650 ( .A1(n14539), .A2(n14540), .ZN(n14662) );
  OR2_X1 U14651 ( .A1(n8974), .A2(n8935), .ZN(n14540) );
  OR2_X1 U14652 ( .A1(n14663), .A2(n14664), .ZN(n14539) );
  AND2_X1 U14653 ( .A1(n14533), .A2(n14536), .ZN(n14664) );
  AND2_X1 U14654 ( .A1(n14665), .A2(n14535), .ZN(n14663) );
  OR2_X1 U14655 ( .A1(n14666), .A2(n14667), .ZN(n14535) );
  AND2_X1 U14656 ( .A1(n14532), .A2(n14531), .ZN(n14667) );
  AND2_X1 U14657 ( .A1(n14529), .A2(n14668), .ZN(n14666) );
  OR2_X1 U14658 ( .A1(n14531), .A2(n14532), .ZN(n14668) );
  OR2_X1 U14659 ( .A1(n8982), .A2(n8935), .ZN(n14532) );
  OR2_X1 U14660 ( .A1(n14669), .A2(n14670), .ZN(n14531) );
  AND2_X1 U14661 ( .A1(n14525), .A2(n14528), .ZN(n14670) );
  AND2_X1 U14662 ( .A1(n14671), .A2(n14527), .ZN(n14669) );
  OR2_X1 U14663 ( .A1(n14672), .A2(n14673), .ZN(n14527) );
  AND2_X1 U14664 ( .A1(n14521), .A2(n14524), .ZN(n14673) );
  AND2_X1 U14665 ( .A1(n14674), .A2(n14523), .ZN(n14672) );
  OR2_X1 U14666 ( .A1(n14675), .A2(n14676), .ZN(n14523) );
  AND2_X1 U14667 ( .A1(n14517), .A2(n14520), .ZN(n14676) );
  AND2_X1 U14668 ( .A1(n14677), .A2(n14519), .ZN(n14675) );
  OR2_X1 U14669 ( .A1(n14678), .A2(n14679), .ZN(n14519) );
  AND2_X1 U14670 ( .A1(n14513), .A2(n14516), .ZN(n14679) );
  AND2_X1 U14671 ( .A1(n14680), .A2(n14515), .ZN(n14678) );
  OR2_X1 U14672 ( .A1(n14681), .A2(n14682), .ZN(n14515) );
  AND2_X1 U14673 ( .A1(n14509), .A2(n14512), .ZN(n14682) );
  AND2_X1 U14674 ( .A1(n14683), .A2(n14511), .ZN(n14681) );
  OR2_X1 U14675 ( .A1(n14684), .A2(n14685), .ZN(n14511) );
  AND2_X1 U14676 ( .A1(n14506), .A2(n14507), .ZN(n14685) );
  AND2_X1 U14677 ( .A1(n14686), .A2(n14508), .ZN(n14684) );
  OR2_X1 U14678 ( .A1(n14687), .A2(n14688), .ZN(n14508) );
  AND2_X1 U14679 ( .A1(n14501), .A2(n14504), .ZN(n14688) );
  AND2_X1 U14680 ( .A1(n14689), .A2(n14503), .ZN(n14687) );
  OR2_X1 U14681 ( .A1(n14690), .A2(n14691), .ZN(n14503) );
  AND2_X1 U14682 ( .A1(n14498), .A2(n14499), .ZN(n14691) );
  AND2_X1 U14683 ( .A1(n14692), .A2(n14693), .ZN(n14690) );
  OR2_X1 U14684 ( .A1(n14499), .A2(n14498), .ZN(n14693) );
  OR2_X1 U14685 ( .A1(n9014), .A2(n8935), .ZN(n14498) );
  OR2_X1 U14686 ( .A1(n9984), .A2(n14694), .ZN(n14499) );
  OR2_X1 U14687 ( .A1(n8935), .A2(n8931), .ZN(n14694) );
  INV_X1 U14688 ( .A(n14500), .ZN(n14692) );
  OR2_X1 U14689 ( .A1(n14695), .A2(n14696), .ZN(n14500) );
  AND2_X1 U14690 ( .A1(b_8_), .A2(n14697), .ZN(n14696) );
  OR2_X1 U14691 ( .A1(n14698), .A2(n9989), .ZN(n14697) );
  AND2_X1 U14692 ( .A1(a_30_), .A2(n8927), .ZN(n14698) );
  AND2_X1 U14693 ( .A1(b_7_), .A2(n14699), .ZN(n14695) );
  OR2_X1 U14694 ( .A1(n14700), .A2(n8021), .ZN(n14699) );
  AND2_X1 U14695 ( .A1(a_31_), .A2(n8931), .ZN(n14700) );
  OR2_X1 U14696 ( .A1(n14504), .A2(n14501), .ZN(n14689) );
  XOR2_X1 U14697 ( .A(n14701), .B(n14702), .Z(n14501) );
  XNOR2_X1 U14698 ( .A(n14703), .B(n14704), .ZN(n14701) );
  OR2_X1 U14699 ( .A1(n9010), .A2(n8935), .ZN(n14504) );
  OR2_X1 U14700 ( .A1(n14507), .A2(n14506), .ZN(n14686) );
  XOR2_X1 U14701 ( .A(n14705), .B(n14706), .Z(n14506) );
  XOR2_X1 U14702 ( .A(n14707), .B(n14708), .Z(n14706) );
  OR2_X1 U14703 ( .A1(n9006), .A2(n8935), .ZN(n14507) );
  OR2_X1 U14704 ( .A1(n14512), .A2(n14509), .ZN(n14683) );
  XNOR2_X1 U14705 ( .A(n14709), .B(n14710), .ZN(n14509) );
  XNOR2_X1 U14706 ( .A(n14711), .B(n14712), .ZN(n14709) );
  OR2_X1 U14707 ( .A1(n9002), .A2(n8935), .ZN(n14512) );
  OR2_X1 U14708 ( .A1(n14516), .A2(n14513), .ZN(n14680) );
  XOR2_X1 U14709 ( .A(n14713), .B(n14714), .Z(n14513) );
  XOR2_X1 U14710 ( .A(n14715), .B(n14716), .Z(n14714) );
  OR2_X1 U14711 ( .A1(n8998), .A2(n8935), .ZN(n14516) );
  OR2_X1 U14712 ( .A1(n14520), .A2(n14517), .ZN(n14677) );
  XOR2_X1 U14713 ( .A(n14717), .B(n14718), .Z(n14517) );
  XOR2_X1 U14714 ( .A(n14719), .B(n14720), .Z(n14718) );
  OR2_X1 U14715 ( .A1(n8994), .A2(n8935), .ZN(n14520) );
  OR2_X1 U14716 ( .A1(n14524), .A2(n14521), .ZN(n14674) );
  XOR2_X1 U14717 ( .A(n14721), .B(n14722), .Z(n14521) );
  XOR2_X1 U14718 ( .A(n14723), .B(n14724), .Z(n14722) );
  OR2_X1 U14719 ( .A1(n8990), .A2(n8935), .ZN(n14524) );
  OR2_X1 U14720 ( .A1(n14528), .A2(n14525), .ZN(n14671) );
  XOR2_X1 U14721 ( .A(n14725), .B(n14726), .Z(n14525) );
  XOR2_X1 U14722 ( .A(n14727), .B(n14728), .Z(n14726) );
  OR2_X1 U14723 ( .A1(n8986), .A2(n8935), .ZN(n14528) );
  XOR2_X1 U14724 ( .A(n14729), .B(n14730), .Z(n14529) );
  XOR2_X1 U14725 ( .A(n14731), .B(n14732), .Z(n14730) );
  OR2_X1 U14726 ( .A1(n14536), .A2(n14533), .ZN(n14665) );
  XOR2_X1 U14727 ( .A(n14733), .B(n14734), .Z(n14533) );
  XOR2_X1 U14728 ( .A(n14735), .B(n14736), .Z(n14734) );
  OR2_X1 U14729 ( .A1(n8978), .A2(n8935), .ZN(n14536) );
  XOR2_X1 U14730 ( .A(n14737), .B(n14738), .Z(n14537) );
  XOR2_X1 U14731 ( .A(n14739), .B(n14740), .Z(n14738) );
  XOR2_X1 U14732 ( .A(n14741), .B(n14742), .Z(n14541) );
  XOR2_X1 U14733 ( .A(n14743), .B(n14744), .Z(n14742) );
  XOR2_X1 U14734 ( .A(n14745), .B(n14746), .Z(n14545) );
  XOR2_X1 U14735 ( .A(n14747), .B(n14748), .Z(n14746) );
  XOR2_X1 U14736 ( .A(n14749), .B(n14750), .Z(n14549) );
  XOR2_X1 U14737 ( .A(n14751), .B(n14752), .Z(n14750) );
  XOR2_X1 U14738 ( .A(n14753), .B(n14754), .Z(n14553) );
  XOR2_X1 U14739 ( .A(n14755), .B(n14756), .Z(n14754) );
  XOR2_X1 U14740 ( .A(n14757), .B(n14758), .Z(n14557) );
  XOR2_X1 U14741 ( .A(n14759), .B(n14760), .Z(n14758) );
  XOR2_X1 U14742 ( .A(n14761), .B(n14762), .Z(n14561) );
  XOR2_X1 U14743 ( .A(n14763), .B(n14764), .Z(n14762) );
  XOR2_X1 U14744 ( .A(n14765), .B(n14766), .Z(n14565) );
  XOR2_X1 U14745 ( .A(n14767), .B(n14768), .Z(n14766) );
  XOR2_X1 U14746 ( .A(n14769), .B(n14770), .Z(n14569) );
  XOR2_X1 U14747 ( .A(n14771), .B(n14772), .Z(n14770) );
  XOR2_X1 U14748 ( .A(n14773), .B(n14774), .Z(n14573) );
  XOR2_X1 U14749 ( .A(n14775), .B(n14776), .Z(n14774) );
  XOR2_X1 U14750 ( .A(n14777), .B(n14778), .Z(n14577) );
  XOR2_X1 U14751 ( .A(n14779), .B(n14780), .Z(n14778) );
  XOR2_X1 U14752 ( .A(n14781), .B(n14782), .Z(n14580) );
  XOR2_X1 U14753 ( .A(n14783), .B(n14784), .Z(n14782) );
  XOR2_X1 U14754 ( .A(n14785), .B(n14786), .Z(n14584) );
  XOR2_X1 U14755 ( .A(n14787), .B(n8654), .Z(n14786) );
  XOR2_X1 U14756 ( .A(n14788), .B(n14789), .Z(n14588) );
  XOR2_X1 U14757 ( .A(n14790), .B(n14791), .Z(n14789) );
  XOR2_X1 U14758 ( .A(n14792), .B(n14793), .Z(n14592) );
  XOR2_X1 U14759 ( .A(n14794), .B(n14795), .Z(n14793) );
  XOR2_X1 U14760 ( .A(n14796), .B(n14797), .Z(n14596) );
  XOR2_X1 U14761 ( .A(n14798), .B(n14799), .Z(n14797) );
  XOR2_X1 U14762 ( .A(n14800), .B(n14801), .Z(n14600) );
  XOR2_X1 U14763 ( .A(n14802), .B(n14803), .Z(n14801) );
  XOR2_X1 U14764 ( .A(n14804), .B(n14805), .Z(n14604) );
  XOR2_X1 U14765 ( .A(n14806), .B(n14807), .Z(n14805) );
  XOR2_X1 U14766 ( .A(n9671), .B(n14808), .Z(n9664) );
  XOR2_X1 U14767 ( .A(n9670), .B(n9669), .Z(n14808) );
  OR2_X1 U14768 ( .A1(n8906), .A2(n8931), .ZN(n9669) );
  OR2_X1 U14769 ( .A1(n14809), .A2(n14810), .ZN(n9670) );
  AND2_X1 U14770 ( .A1(n14807), .A2(n14806), .ZN(n14810) );
  AND2_X1 U14771 ( .A1(n14804), .A2(n14811), .ZN(n14809) );
  OR2_X1 U14772 ( .A1(n14806), .A2(n14807), .ZN(n14811) );
  OR2_X1 U14773 ( .A1(n8910), .A2(n8931), .ZN(n14807) );
  OR2_X1 U14774 ( .A1(n14812), .A2(n14813), .ZN(n14806) );
  AND2_X1 U14775 ( .A1(n14803), .A2(n14802), .ZN(n14813) );
  AND2_X1 U14776 ( .A1(n14800), .A2(n14814), .ZN(n14812) );
  OR2_X1 U14777 ( .A1(n14802), .A2(n14803), .ZN(n14814) );
  OR2_X1 U14778 ( .A1(n8914), .A2(n8931), .ZN(n14803) );
  OR2_X1 U14779 ( .A1(n14815), .A2(n14816), .ZN(n14802) );
  AND2_X1 U14780 ( .A1(n14799), .A2(n14798), .ZN(n14816) );
  AND2_X1 U14781 ( .A1(n14796), .A2(n14817), .ZN(n14815) );
  OR2_X1 U14782 ( .A1(n14798), .A2(n14799), .ZN(n14817) );
  OR2_X1 U14783 ( .A1(n8918), .A2(n8931), .ZN(n14799) );
  OR2_X1 U14784 ( .A1(n14818), .A2(n14819), .ZN(n14798) );
  AND2_X1 U14785 ( .A1(n14795), .A2(n14794), .ZN(n14819) );
  AND2_X1 U14786 ( .A1(n14792), .A2(n14820), .ZN(n14818) );
  OR2_X1 U14787 ( .A1(n14794), .A2(n14795), .ZN(n14820) );
  OR2_X1 U14788 ( .A1(n8922), .A2(n8931), .ZN(n14795) );
  OR2_X1 U14789 ( .A1(n14821), .A2(n14822), .ZN(n14794) );
  AND2_X1 U14790 ( .A1(n14791), .A2(n14790), .ZN(n14822) );
  AND2_X1 U14791 ( .A1(n14788), .A2(n14823), .ZN(n14821) );
  OR2_X1 U14792 ( .A1(n14790), .A2(n14791), .ZN(n14823) );
  OR2_X1 U14793 ( .A1(n8926), .A2(n8931), .ZN(n14791) );
  OR2_X1 U14794 ( .A1(n14824), .A2(n14825), .ZN(n14790) );
  AND2_X1 U14795 ( .A1(n8654), .A2(n14787), .ZN(n14825) );
  AND2_X1 U14796 ( .A1(n14785), .A2(n14826), .ZN(n14824) );
  OR2_X1 U14797 ( .A1(n14787), .A2(n8654), .ZN(n14826) );
  OR2_X1 U14798 ( .A1(n8930), .A2(n8931), .ZN(n8654) );
  OR2_X1 U14799 ( .A1(n14827), .A2(n14828), .ZN(n14787) );
  AND2_X1 U14800 ( .A1(n14784), .A2(n14783), .ZN(n14828) );
  AND2_X1 U14801 ( .A1(n14781), .A2(n14829), .ZN(n14827) );
  OR2_X1 U14802 ( .A1(n14783), .A2(n14784), .ZN(n14829) );
  OR2_X1 U14803 ( .A1(n8934), .A2(n8931), .ZN(n14784) );
  OR2_X1 U14804 ( .A1(n14830), .A2(n14831), .ZN(n14783) );
  AND2_X1 U14805 ( .A1(n14780), .A2(n14779), .ZN(n14831) );
  AND2_X1 U14806 ( .A1(n14777), .A2(n14832), .ZN(n14830) );
  OR2_X1 U14807 ( .A1(n14779), .A2(n14780), .ZN(n14832) );
  OR2_X1 U14808 ( .A1(n8938), .A2(n8931), .ZN(n14780) );
  OR2_X1 U14809 ( .A1(n14833), .A2(n14834), .ZN(n14779) );
  AND2_X1 U14810 ( .A1(n14776), .A2(n14775), .ZN(n14834) );
  AND2_X1 U14811 ( .A1(n14773), .A2(n14835), .ZN(n14833) );
  OR2_X1 U14812 ( .A1(n14775), .A2(n14776), .ZN(n14835) );
  OR2_X1 U14813 ( .A1(n8942), .A2(n8931), .ZN(n14776) );
  OR2_X1 U14814 ( .A1(n14836), .A2(n14837), .ZN(n14775) );
  AND2_X1 U14815 ( .A1(n14772), .A2(n14771), .ZN(n14837) );
  AND2_X1 U14816 ( .A1(n14769), .A2(n14838), .ZN(n14836) );
  OR2_X1 U14817 ( .A1(n14771), .A2(n14772), .ZN(n14838) );
  OR2_X1 U14818 ( .A1(n8946), .A2(n8931), .ZN(n14772) );
  OR2_X1 U14819 ( .A1(n14839), .A2(n14840), .ZN(n14771) );
  AND2_X1 U14820 ( .A1(n14768), .A2(n14767), .ZN(n14840) );
  AND2_X1 U14821 ( .A1(n14765), .A2(n14841), .ZN(n14839) );
  OR2_X1 U14822 ( .A1(n14767), .A2(n14768), .ZN(n14841) );
  OR2_X1 U14823 ( .A1(n8950), .A2(n8931), .ZN(n14768) );
  OR2_X1 U14824 ( .A1(n14842), .A2(n14843), .ZN(n14767) );
  AND2_X1 U14825 ( .A1(n14764), .A2(n14763), .ZN(n14843) );
  AND2_X1 U14826 ( .A1(n14761), .A2(n14844), .ZN(n14842) );
  OR2_X1 U14827 ( .A1(n14763), .A2(n14764), .ZN(n14844) );
  OR2_X1 U14828 ( .A1(n8954), .A2(n8931), .ZN(n14764) );
  OR2_X1 U14829 ( .A1(n14845), .A2(n14846), .ZN(n14763) );
  AND2_X1 U14830 ( .A1(n14760), .A2(n14759), .ZN(n14846) );
  AND2_X1 U14831 ( .A1(n14757), .A2(n14847), .ZN(n14845) );
  OR2_X1 U14832 ( .A1(n14759), .A2(n14760), .ZN(n14847) );
  OR2_X1 U14833 ( .A1(n8958), .A2(n8931), .ZN(n14760) );
  OR2_X1 U14834 ( .A1(n14848), .A2(n14849), .ZN(n14759) );
  AND2_X1 U14835 ( .A1(n14756), .A2(n14755), .ZN(n14849) );
  AND2_X1 U14836 ( .A1(n14753), .A2(n14850), .ZN(n14848) );
  OR2_X1 U14837 ( .A1(n14755), .A2(n14756), .ZN(n14850) );
  OR2_X1 U14838 ( .A1(n8962), .A2(n8931), .ZN(n14756) );
  OR2_X1 U14839 ( .A1(n14851), .A2(n14852), .ZN(n14755) );
  AND2_X1 U14840 ( .A1(n14752), .A2(n14751), .ZN(n14852) );
  AND2_X1 U14841 ( .A1(n14749), .A2(n14853), .ZN(n14851) );
  OR2_X1 U14842 ( .A1(n14751), .A2(n14752), .ZN(n14853) );
  OR2_X1 U14843 ( .A1(n8966), .A2(n8931), .ZN(n14752) );
  OR2_X1 U14844 ( .A1(n14854), .A2(n14855), .ZN(n14751) );
  AND2_X1 U14845 ( .A1(n14748), .A2(n14747), .ZN(n14855) );
  AND2_X1 U14846 ( .A1(n14745), .A2(n14856), .ZN(n14854) );
  OR2_X1 U14847 ( .A1(n14747), .A2(n14748), .ZN(n14856) );
  OR2_X1 U14848 ( .A1(n8970), .A2(n8931), .ZN(n14748) );
  OR2_X1 U14849 ( .A1(n14857), .A2(n14858), .ZN(n14747) );
  AND2_X1 U14850 ( .A1(n14744), .A2(n14743), .ZN(n14858) );
  AND2_X1 U14851 ( .A1(n14741), .A2(n14859), .ZN(n14857) );
  OR2_X1 U14852 ( .A1(n14743), .A2(n14744), .ZN(n14859) );
  OR2_X1 U14853 ( .A1(n8974), .A2(n8931), .ZN(n14744) );
  OR2_X1 U14854 ( .A1(n14860), .A2(n14861), .ZN(n14743) );
  AND2_X1 U14855 ( .A1(n14740), .A2(n14739), .ZN(n14861) );
  AND2_X1 U14856 ( .A1(n14737), .A2(n14862), .ZN(n14860) );
  OR2_X1 U14857 ( .A1(n14739), .A2(n14740), .ZN(n14862) );
  OR2_X1 U14858 ( .A1(n8978), .A2(n8931), .ZN(n14740) );
  OR2_X1 U14859 ( .A1(n14863), .A2(n14864), .ZN(n14739) );
  AND2_X1 U14860 ( .A1(n14733), .A2(n14736), .ZN(n14864) );
  AND2_X1 U14861 ( .A1(n14865), .A2(n14735), .ZN(n14863) );
  OR2_X1 U14862 ( .A1(n14866), .A2(n14867), .ZN(n14735) );
  AND2_X1 U14863 ( .A1(n14732), .A2(n14731), .ZN(n14867) );
  AND2_X1 U14864 ( .A1(n14729), .A2(n14868), .ZN(n14866) );
  OR2_X1 U14865 ( .A1(n14731), .A2(n14732), .ZN(n14868) );
  OR2_X1 U14866 ( .A1(n8986), .A2(n8931), .ZN(n14732) );
  OR2_X1 U14867 ( .A1(n14869), .A2(n14870), .ZN(n14731) );
  AND2_X1 U14868 ( .A1(n14725), .A2(n14728), .ZN(n14870) );
  AND2_X1 U14869 ( .A1(n14871), .A2(n14727), .ZN(n14869) );
  OR2_X1 U14870 ( .A1(n14872), .A2(n14873), .ZN(n14727) );
  AND2_X1 U14871 ( .A1(n14721), .A2(n14724), .ZN(n14873) );
  AND2_X1 U14872 ( .A1(n14874), .A2(n14723), .ZN(n14872) );
  OR2_X1 U14873 ( .A1(n14875), .A2(n14876), .ZN(n14723) );
  AND2_X1 U14874 ( .A1(n14717), .A2(n14720), .ZN(n14876) );
  AND2_X1 U14875 ( .A1(n14877), .A2(n14719), .ZN(n14875) );
  OR2_X1 U14876 ( .A1(n14878), .A2(n14879), .ZN(n14719) );
  AND2_X1 U14877 ( .A1(n14713), .A2(n14716), .ZN(n14879) );
  AND2_X1 U14878 ( .A1(n14880), .A2(n14715), .ZN(n14878) );
  OR2_X1 U14879 ( .A1(n14881), .A2(n14882), .ZN(n14715) );
  AND2_X1 U14880 ( .A1(n14710), .A2(n14711), .ZN(n14882) );
  AND2_X1 U14881 ( .A1(n14883), .A2(n14712), .ZN(n14881) );
  OR2_X1 U14882 ( .A1(n14884), .A2(n14885), .ZN(n14712) );
  AND2_X1 U14883 ( .A1(n14705), .A2(n14708), .ZN(n14885) );
  AND2_X1 U14884 ( .A1(n14886), .A2(n14707), .ZN(n14884) );
  OR2_X1 U14885 ( .A1(n14887), .A2(n14888), .ZN(n14707) );
  AND2_X1 U14886 ( .A1(n14702), .A2(n14703), .ZN(n14888) );
  AND2_X1 U14887 ( .A1(n14889), .A2(n14890), .ZN(n14887) );
  OR2_X1 U14888 ( .A1(n14703), .A2(n14702), .ZN(n14890) );
  OR2_X1 U14889 ( .A1(n9014), .A2(n8931), .ZN(n14702) );
  OR2_X1 U14890 ( .A1(n9984), .A2(n14891), .ZN(n14703) );
  OR2_X1 U14891 ( .A1(n8931), .A2(n8927), .ZN(n14891) );
  INV_X1 U14892 ( .A(n14704), .ZN(n14889) );
  OR2_X1 U14893 ( .A1(n14892), .A2(n14893), .ZN(n14704) );
  AND2_X1 U14894 ( .A1(b_7_), .A2(n14894), .ZN(n14893) );
  OR2_X1 U14895 ( .A1(n14895), .A2(n9989), .ZN(n14894) );
  AND2_X1 U14896 ( .A1(a_30_), .A2(n8923), .ZN(n14895) );
  AND2_X1 U14897 ( .A1(b_6_), .A2(n14896), .ZN(n14892) );
  OR2_X1 U14898 ( .A1(n14897), .A2(n8021), .ZN(n14896) );
  AND2_X1 U14899 ( .A1(a_31_), .A2(n8927), .ZN(n14897) );
  OR2_X1 U14900 ( .A1(n14708), .A2(n14705), .ZN(n14886) );
  XOR2_X1 U14901 ( .A(n14898), .B(n14899), .Z(n14705) );
  XNOR2_X1 U14902 ( .A(n14900), .B(n14901), .ZN(n14898) );
  OR2_X1 U14903 ( .A1(n9010), .A2(n8931), .ZN(n14708) );
  OR2_X1 U14904 ( .A1(n14711), .A2(n14710), .ZN(n14883) );
  XOR2_X1 U14905 ( .A(n14902), .B(n14903), .Z(n14710) );
  XOR2_X1 U14906 ( .A(n14904), .B(n14905), .Z(n14903) );
  OR2_X1 U14907 ( .A1(n9006), .A2(n8931), .ZN(n14711) );
  OR2_X1 U14908 ( .A1(n14716), .A2(n14713), .ZN(n14880) );
  XNOR2_X1 U14909 ( .A(n14906), .B(n14907), .ZN(n14713) );
  XNOR2_X1 U14910 ( .A(n14908), .B(n14909), .ZN(n14906) );
  OR2_X1 U14911 ( .A1(n9002), .A2(n8931), .ZN(n14716) );
  OR2_X1 U14912 ( .A1(n14720), .A2(n14717), .ZN(n14877) );
  XOR2_X1 U14913 ( .A(n14910), .B(n14911), .Z(n14717) );
  XOR2_X1 U14914 ( .A(n14912), .B(n14913), .Z(n14911) );
  OR2_X1 U14915 ( .A1(n8998), .A2(n8931), .ZN(n14720) );
  OR2_X1 U14916 ( .A1(n14724), .A2(n14721), .ZN(n14874) );
  XOR2_X1 U14917 ( .A(n14914), .B(n14915), .Z(n14721) );
  XOR2_X1 U14918 ( .A(n14916), .B(n14917), .Z(n14915) );
  OR2_X1 U14919 ( .A1(n8994), .A2(n8931), .ZN(n14724) );
  OR2_X1 U14920 ( .A1(n14728), .A2(n14725), .ZN(n14871) );
  XOR2_X1 U14921 ( .A(n14918), .B(n14919), .Z(n14725) );
  XOR2_X1 U14922 ( .A(n14920), .B(n14921), .Z(n14919) );
  OR2_X1 U14923 ( .A1(n8990), .A2(n8931), .ZN(n14728) );
  XOR2_X1 U14924 ( .A(n14922), .B(n14923), .Z(n14729) );
  XOR2_X1 U14925 ( .A(n14924), .B(n14925), .Z(n14923) );
  OR2_X1 U14926 ( .A1(n14736), .A2(n14733), .ZN(n14865) );
  XOR2_X1 U14927 ( .A(n14926), .B(n14927), .Z(n14733) );
  XOR2_X1 U14928 ( .A(n14928), .B(n14929), .Z(n14927) );
  OR2_X1 U14929 ( .A1(n8982), .A2(n8931), .ZN(n14736) );
  XOR2_X1 U14930 ( .A(n14930), .B(n14931), .Z(n14737) );
  XOR2_X1 U14931 ( .A(n14932), .B(n14933), .Z(n14931) );
  XOR2_X1 U14932 ( .A(n14934), .B(n14935), .Z(n14741) );
  XOR2_X1 U14933 ( .A(n14936), .B(n14937), .Z(n14935) );
  XOR2_X1 U14934 ( .A(n14938), .B(n14939), .Z(n14745) );
  XOR2_X1 U14935 ( .A(n14940), .B(n14941), .Z(n14939) );
  XOR2_X1 U14936 ( .A(n14942), .B(n14943), .Z(n14749) );
  XOR2_X1 U14937 ( .A(n14944), .B(n14945), .Z(n14943) );
  XOR2_X1 U14938 ( .A(n14946), .B(n14947), .Z(n14753) );
  XOR2_X1 U14939 ( .A(n14948), .B(n14949), .Z(n14947) );
  XOR2_X1 U14940 ( .A(n14950), .B(n14951), .Z(n14757) );
  XOR2_X1 U14941 ( .A(n14952), .B(n14953), .Z(n14951) );
  XOR2_X1 U14942 ( .A(n14954), .B(n14955), .Z(n14761) );
  XOR2_X1 U14943 ( .A(n14956), .B(n14957), .Z(n14955) );
  XOR2_X1 U14944 ( .A(n14958), .B(n14959), .Z(n14765) );
  XOR2_X1 U14945 ( .A(n14960), .B(n14961), .Z(n14959) );
  XOR2_X1 U14946 ( .A(n14962), .B(n14963), .Z(n14769) );
  XOR2_X1 U14947 ( .A(n14964), .B(n14965), .Z(n14963) );
  XOR2_X1 U14948 ( .A(n14966), .B(n14967), .Z(n14773) );
  XOR2_X1 U14949 ( .A(n14968), .B(n14969), .Z(n14967) );
  XOR2_X1 U14950 ( .A(n14970), .B(n14971), .Z(n14777) );
  XOR2_X1 U14951 ( .A(n14972), .B(n14973), .Z(n14971) );
  XOR2_X1 U14952 ( .A(n14974), .B(n14975), .Z(n14781) );
  XOR2_X1 U14953 ( .A(n14976), .B(n14977), .Z(n14975) );
  XOR2_X1 U14954 ( .A(n14978), .B(n14979), .Z(n14785) );
  XOR2_X1 U14955 ( .A(n14980), .B(n14981), .Z(n14979) );
  XOR2_X1 U14956 ( .A(n14982), .B(n14983), .Z(n14788) );
  XOR2_X1 U14957 ( .A(n14984), .B(n14985), .Z(n14983) );
  XOR2_X1 U14958 ( .A(n14986), .B(n14987), .Z(n14792) );
  XOR2_X1 U14959 ( .A(n14988), .B(n8692), .Z(n14987) );
  XOR2_X1 U14960 ( .A(n14989), .B(n14990), .Z(n14796) );
  XOR2_X1 U14961 ( .A(n14991), .B(n14992), .Z(n14990) );
  XOR2_X1 U14962 ( .A(n14993), .B(n14994), .Z(n14800) );
  XOR2_X1 U14963 ( .A(n14995), .B(n14996), .Z(n14994) );
  XOR2_X1 U14964 ( .A(n14997), .B(n14998), .Z(n14804) );
  XOR2_X1 U14965 ( .A(n14999), .B(n15000), .Z(n14998) );
  XOR2_X1 U14966 ( .A(n9678), .B(n15001), .Z(n9671) );
  XOR2_X1 U14967 ( .A(n9677), .B(n9676), .Z(n15001) );
  OR2_X1 U14968 ( .A1(n8910), .A2(n8927), .ZN(n9676) );
  OR2_X1 U14969 ( .A1(n15002), .A2(n15003), .ZN(n9677) );
  AND2_X1 U14970 ( .A1(n15000), .A2(n14999), .ZN(n15003) );
  AND2_X1 U14971 ( .A1(n14997), .A2(n15004), .ZN(n15002) );
  OR2_X1 U14972 ( .A1(n14999), .A2(n15000), .ZN(n15004) );
  OR2_X1 U14973 ( .A1(n8914), .A2(n8927), .ZN(n15000) );
  OR2_X1 U14974 ( .A1(n15005), .A2(n15006), .ZN(n14999) );
  AND2_X1 U14975 ( .A1(n14996), .A2(n14995), .ZN(n15006) );
  AND2_X1 U14976 ( .A1(n14993), .A2(n15007), .ZN(n15005) );
  OR2_X1 U14977 ( .A1(n14995), .A2(n14996), .ZN(n15007) );
  OR2_X1 U14978 ( .A1(n8918), .A2(n8927), .ZN(n14996) );
  OR2_X1 U14979 ( .A1(n15008), .A2(n15009), .ZN(n14995) );
  AND2_X1 U14980 ( .A1(n14992), .A2(n14991), .ZN(n15009) );
  AND2_X1 U14981 ( .A1(n14989), .A2(n15010), .ZN(n15008) );
  OR2_X1 U14982 ( .A1(n14991), .A2(n14992), .ZN(n15010) );
  OR2_X1 U14983 ( .A1(n8922), .A2(n8927), .ZN(n14992) );
  OR2_X1 U14984 ( .A1(n15011), .A2(n15012), .ZN(n14991) );
  AND2_X1 U14985 ( .A1(n8692), .A2(n14988), .ZN(n15012) );
  AND2_X1 U14986 ( .A1(n14986), .A2(n15013), .ZN(n15011) );
  OR2_X1 U14987 ( .A1(n14988), .A2(n8692), .ZN(n15013) );
  OR2_X1 U14988 ( .A1(n8926), .A2(n8927), .ZN(n8692) );
  OR2_X1 U14989 ( .A1(n15014), .A2(n15015), .ZN(n14988) );
  AND2_X1 U14990 ( .A1(n14985), .A2(n14984), .ZN(n15015) );
  AND2_X1 U14991 ( .A1(n14982), .A2(n15016), .ZN(n15014) );
  OR2_X1 U14992 ( .A1(n14984), .A2(n14985), .ZN(n15016) );
  OR2_X1 U14993 ( .A1(n8930), .A2(n8927), .ZN(n14985) );
  OR2_X1 U14994 ( .A1(n15017), .A2(n15018), .ZN(n14984) );
  AND2_X1 U14995 ( .A1(n14981), .A2(n14980), .ZN(n15018) );
  AND2_X1 U14996 ( .A1(n14978), .A2(n15019), .ZN(n15017) );
  OR2_X1 U14997 ( .A1(n14980), .A2(n14981), .ZN(n15019) );
  OR2_X1 U14998 ( .A1(n8934), .A2(n8927), .ZN(n14981) );
  OR2_X1 U14999 ( .A1(n15020), .A2(n15021), .ZN(n14980) );
  AND2_X1 U15000 ( .A1(n14977), .A2(n14976), .ZN(n15021) );
  AND2_X1 U15001 ( .A1(n14974), .A2(n15022), .ZN(n15020) );
  OR2_X1 U15002 ( .A1(n14976), .A2(n14977), .ZN(n15022) );
  OR2_X1 U15003 ( .A1(n8938), .A2(n8927), .ZN(n14977) );
  OR2_X1 U15004 ( .A1(n15023), .A2(n15024), .ZN(n14976) );
  AND2_X1 U15005 ( .A1(n14973), .A2(n14972), .ZN(n15024) );
  AND2_X1 U15006 ( .A1(n14970), .A2(n15025), .ZN(n15023) );
  OR2_X1 U15007 ( .A1(n14972), .A2(n14973), .ZN(n15025) );
  OR2_X1 U15008 ( .A1(n8942), .A2(n8927), .ZN(n14973) );
  OR2_X1 U15009 ( .A1(n15026), .A2(n15027), .ZN(n14972) );
  AND2_X1 U15010 ( .A1(n14969), .A2(n14968), .ZN(n15027) );
  AND2_X1 U15011 ( .A1(n14966), .A2(n15028), .ZN(n15026) );
  OR2_X1 U15012 ( .A1(n14968), .A2(n14969), .ZN(n15028) );
  OR2_X1 U15013 ( .A1(n8946), .A2(n8927), .ZN(n14969) );
  OR2_X1 U15014 ( .A1(n15029), .A2(n15030), .ZN(n14968) );
  AND2_X1 U15015 ( .A1(n14965), .A2(n14964), .ZN(n15030) );
  AND2_X1 U15016 ( .A1(n14962), .A2(n15031), .ZN(n15029) );
  OR2_X1 U15017 ( .A1(n14964), .A2(n14965), .ZN(n15031) );
  OR2_X1 U15018 ( .A1(n8950), .A2(n8927), .ZN(n14965) );
  OR2_X1 U15019 ( .A1(n15032), .A2(n15033), .ZN(n14964) );
  AND2_X1 U15020 ( .A1(n14961), .A2(n14960), .ZN(n15033) );
  AND2_X1 U15021 ( .A1(n14958), .A2(n15034), .ZN(n15032) );
  OR2_X1 U15022 ( .A1(n14960), .A2(n14961), .ZN(n15034) );
  OR2_X1 U15023 ( .A1(n8954), .A2(n8927), .ZN(n14961) );
  OR2_X1 U15024 ( .A1(n15035), .A2(n15036), .ZN(n14960) );
  AND2_X1 U15025 ( .A1(n14957), .A2(n14956), .ZN(n15036) );
  AND2_X1 U15026 ( .A1(n14954), .A2(n15037), .ZN(n15035) );
  OR2_X1 U15027 ( .A1(n14956), .A2(n14957), .ZN(n15037) );
  OR2_X1 U15028 ( .A1(n8958), .A2(n8927), .ZN(n14957) );
  OR2_X1 U15029 ( .A1(n15038), .A2(n15039), .ZN(n14956) );
  AND2_X1 U15030 ( .A1(n14953), .A2(n14952), .ZN(n15039) );
  AND2_X1 U15031 ( .A1(n14950), .A2(n15040), .ZN(n15038) );
  OR2_X1 U15032 ( .A1(n14952), .A2(n14953), .ZN(n15040) );
  OR2_X1 U15033 ( .A1(n8962), .A2(n8927), .ZN(n14953) );
  OR2_X1 U15034 ( .A1(n15041), .A2(n15042), .ZN(n14952) );
  AND2_X1 U15035 ( .A1(n14949), .A2(n14948), .ZN(n15042) );
  AND2_X1 U15036 ( .A1(n14946), .A2(n15043), .ZN(n15041) );
  OR2_X1 U15037 ( .A1(n14948), .A2(n14949), .ZN(n15043) );
  OR2_X1 U15038 ( .A1(n8966), .A2(n8927), .ZN(n14949) );
  OR2_X1 U15039 ( .A1(n15044), .A2(n15045), .ZN(n14948) );
  AND2_X1 U15040 ( .A1(n14945), .A2(n14944), .ZN(n15045) );
  AND2_X1 U15041 ( .A1(n14942), .A2(n15046), .ZN(n15044) );
  OR2_X1 U15042 ( .A1(n14944), .A2(n14945), .ZN(n15046) );
  OR2_X1 U15043 ( .A1(n8970), .A2(n8927), .ZN(n14945) );
  OR2_X1 U15044 ( .A1(n15047), .A2(n15048), .ZN(n14944) );
  AND2_X1 U15045 ( .A1(n14941), .A2(n14940), .ZN(n15048) );
  AND2_X1 U15046 ( .A1(n14938), .A2(n15049), .ZN(n15047) );
  OR2_X1 U15047 ( .A1(n14940), .A2(n14941), .ZN(n15049) );
  OR2_X1 U15048 ( .A1(n8974), .A2(n8927), .ZN(n14941) );
  OR2_X1 U15049 ( .A1(n15050), .A2(n15051), .ZN(n14940) );
  AND2_X1 U15050 ( .A1(n14937), .A2(n14936), .ZN(n15051) );
  AND2_X1 U15051 ( .A1(n14934), .A2(n15052), .ZN(n15050) );
  OR2_X1 U15052 ( .A1(n14936), .A2(n14937), .ZN(n15052) );
  OR2_X1 U15053 ( .A1(n8978), .A2(n8927), .ZN(n14937) );
  OR2_X1 U15054 ( .A1(n15053), .A2(n15054), .ZN(n14936) );
  AND2_X1 U15055 ( .A1(n14933), .A2(n14932), .ZN(n15054) );
  AND2_X1 U15056 ( .A1(n14930), .A2(n15055), .ZN(n15053) );
  OR2_X1 U15057 ( .A1(n14932), .A2(n14933), .ZN(n15055) );
  OR2_X1 U15058 ( .A1(n8982), .A2(n8927), .ZN(n14933) );
  OR2_X1 U15059 ( .A1(n15056), .A2(n15057), .ZN(n14932) );
  AND2_X1 U15060 ( .A1(n14926), .A2(n14929), .ZN(n15057) );
  AND2_X1 U15061 ( .A1(n15058), .A2(n14928), .ZN(n15056) );
  OR2_X1 U15062 ( .A1(n15059), .A2(n15060), .ZN(n14928) );
  AND2_X1 U15063 ( .A1(n14925), .A2(n14924), .ZN(n15060) );
  AND2_X1 U15064 ( .A1(n14922), .A2(n15061), .ZN(n15059) );
  OR2_X1 U15065 ( .A1(n14924), .A2(n14925), .ZN(n15061) );
  OR2_X1 U15066 ( .A1(n8990), .A2(n8927), .ZN(n14925) );
  OR2_X1 U15067 ( .A1(n15062), .A2(n15063), .ZN(n14924) );
  AND2_X1 U15068 ( .A1(n14918), .A2(n14921), .ZN(n15063) );
  AND2_X1 U15069 ( .A1(n15064), .A2(n14920), .ZN(n15062) );
  OR2_X1 U15070 ( .A1(n15065), .A2(n15066), .ZN(n14920) );
  AND2_X1 U15071 ( .A1(n14914), .A2(n14917), .ZN(n15066) );
  AND2_X1 U15072 ( .A1(n15067), .A2(n14916), .ZN(n15065) );
  OR2_X1 U15073 ( .A1(n15068), .A2(n15069), .ZN(n14916) );
  AND2_X1 U15074 ( .A1(n14910), .A2(n14913), .ZN(n15069) );
  AND2_X1 U15075 ( .A1(n15070), .A2(n14912), .ZN(n15068) );
  OR2_X1 U15076 ( .A1(n15071), .A2(n15072), .ZN(n14912) );
  AND2_X1 U15077 ( .A1(n14907), .A2(n14908), .ZN(n15072) );
  AND2_X1 U15078 ( .A1(n15073), .A2(n14909), .ZN(n15071) );
  OR2_X1 U15079 ( .A1(n15074), .A2(n15075), .ZN(n14909) );
  AND2_X1 U15080 ( .A1(n14902), .A2(n14905), .ZN(n15075) );
  AND2_X1 U15081 ( .A1(n15076), .A2(n14904), .ZN(n15074) );
  OR2_X1 U15082 ( .A1(n15077), .A2(n15078), .ZN(n14904) );
  AND2_X1 U15083 ( .A1(n14899), .A2(n14900), .ZN(n15078) );
  AND2_X1 U15084 ( .A1(n15079), .A2(n15080), .ZN(n15077) );
  OR2_X1 U15085 ( .A1(n14900), .A2(n14899), .ZN(n15080) );
  OR2_X1 U15086 ( .A1(n9014), .A2(n8927), .ZN(n14899) );
  OR2_X1 U15087 ( .A1(n9984), .A2(n15081), .ZN(n14900) );
  OR2_X1 U15088 ( .A1(n8927), .A2(n8923), .ZN(n15081) );
  INV_X1 U15089 ( .A(n14901), .ZN(n15079) );
  OR2_X1 U15090 ( .A1(n15082), .A2(n15083), .ZN(n14901) );
  AND2_X1 U15091 ( .A1(b_6_), .A2(n15084), .ZN(n15083) );
  OR2_X1 U15092 ( .A1(n15085), .A2(n9989), .ZN(n15084) );
  AND2_X1 U15093 ( .A1(a_30_), .A2(n8919), .ZN(n15085) );
  AND2_X1 U15094 ( .A1(b_5_), .A2(n15086), .ZN(n15082) );
  OR2_X1 U15095 ( .A1(n15087), .A2(n8021), .ZN(n15086) );
  AND2_X1 U15096 ( .A1(a_31_), .A2(n8923), .ZN(n15087) );
  OR2_X1 U15097 ( .A1(n14905), .A2(n14902), .ZN(n15076) );
  XOR2_X1 U15098 ( .A(n15088), .B(n15089), .Z(n14902) );
  XNOR2_X1 U15099 ( .A(n15090), .B(n15091), .ZN(n15088) );
  OR2_X1 U15100 ( .A1(n9010), .A2(n8927), .ZN(n14905) );
  OR2_X1 U15101 ( .A1(n14908), .A2(n14907), .ZN(n15073) );
  XOR2_X1 U15102 ( .A(n15092), .B(n15093), .Z(n14907) );
  XOR2_X1 U15103 ( .A(n15094), .B(n15095), .Z(n15093) );
  OR2_X1 U15104 ( .A1(n9006), .A2(n8927), .ZN(n14908) );
  OR2_X1 U15105 ( .A1(n14913), .A2(n14910), .ZN(n15070) );
  XNOR2_X1 U15106 ( .A(n15096), .B(n15097), .ZN(n14910) );
  XNOR2_X1 U15107 ( .A(n15098), .B(n15099), .ZN(n15096) );
  OR2_X1 U15108 ( .A1(n9002), .A2(n8927), .ZN(n14913) );
  OR2_X1 U15109 ( .A1(n14917), .A2(n14914), .ZN(n15067) );
  XOR2_X1 U15110 ( .A(n15100), .B(n15101), .Z(n14914) );
  XOR2_X1 U15111 ( .A(n15102), .B(n15103), .Z(n15101) );
  OR2_X1 U15112 ( .A1(n8998), .A2(n8927), .ZN(n14917) );
  OR2_X1 U15113 ( .A1(n14921), .A2(n14918), .ZN(n15064) );
  XOR2_X1 U15114 ( .A(n15104), .B(n15105), .Z(n14918) );
  XOR2_X1 U15115 ( .A(n15106), .B(n15107), .Z(n15105) );
  OR2_X1 U15116 ( .A1(n8994), .A2(n8927), .ZN(n14921) );
  XOR2_X1 U15117 ( .A(n15108), .B(n15109), .Z(n14922) );
  XOR2_X1 U15118 ( .A(n15110), .B(n15111), .Z(n15109) );
  OR2_X1 U15119 ( .A1(n14929), .A2(n14926), .ZN(n15058) );
  XOR2_X1 U15120 ( .A(n15112), .B(n15113), .Z(n14926) );
  XOR2_X1 U15121 ( .A(n15114), .B(n15115), .Z(n15113) );
  OR2_X1 U15122 ( .A1(n8986), .A2(n8927), .ZN(n14929) );
  XOR2_X1 U15123 ( .A(n15116), .B(n15117), .Z(n14930) );
  XOR2_X1 U15124 ( .A(n15118), .B(n15119), .Z(n15117) );
  XOR2_X1 U15125 ( .A(n15120), .B(n15121), .Z(n14934) );
  XOR2_X1 U15126 ( .A(n15122), .B(n15123), .Z(n15121) );
  XOR2_X1 U15127 ( .A(n15124), .B(n15125), .Z(n14938) );
  XOR2_X1 U15128 ( .A(n15126), .B(n15127), .Z(n15125) );
  XOR2_X1 U15129 ( .A(n15128), .B(n15129), .Z(n14942) );
  XOR2_X1 U15130 ( .A(n15130), .B(n15131), .Z(n15129) );
  XOR2_X1 U15131 ( .A(n15132), .B(n15133), .Z(n14946) );
  XOR2_X1 U15132 ( .A(n15134), .B(n15135), .Z(n15133) );
  XOR2_X1 U15133 ( .A(n15136), .B(n15137), .Z(n14950) );
  XOR2_X1 U15134 ( .A(n15138), .B(n15139), .Z(n15137) );
  XOR2_X1 U15135 ( .A(n15140), .B(n15141), .Z(n14954) );
  XOR2_X1 U15136 ( .A(n15142), .B(n15143), .Z(n15141) );
  XOR2_X1 U15137 ( .A(n15144), .B(n15145), .Z(n14958) );
  XOR2_X1 U15138 ( .A(n15146), .B(n15147), .Z(n15145) );
  XOR2_X1 U15139 ( .A(n15148), .B(n15149), .Z(n14962) );
  XOR2_X1 U15140 ( .A(n15150), .B(n15151), .Z(n15149) );
  XOR2_X1 U15141 ( .A(n15152), .B(n15153), .Z(n14966) );
  XOR2_X1 U15142 ( .A(n15154), .B(n15155), .Z(n15153) );
  XOR2_X1 U15143 ( .A(n15156), .B(n15157), .Z(n14970) );
  XOR2_X1 U15144 ( .A(n15158), .B(n15159), .Z(n15157) );
  XOR2_X1 U15145 ( .A(n15160), .B(n15161), .Z(n14974) );
  XOR2_X1 U15146 ( .A(n15162), .B(n15163), .Z(n15161) );
  XOR2_X1 U15147 ( .A(n15164), .B(n15165), .Z(n14978) );
  XOR2_X1 U15148 ( .A(n15166), .B(n15167), .Z(n15165) );
  XOR2_X1 U15149 ( .A(n15168), .B(n15169), .Z(n14982) );
  XOR2_X1 U15150 ( .A(n15170), .B(n15171), .Z(n15169) );
  XOR2_X1 U15151 ( .A(n15172), .B(n15173), .Z(n14986) );
  XOR2_X1 U15152 ( .A(n15174), .B(n15175), .Z(n15173) );
  XOR2_X1 U15153 ( .A(n15176), .B(n15177), .Z(n14989) );
  XOR2_X1 U15154 ( .A(n15178), .B(n15179), .Z(n15177) );
  XOR2_X1 U15155 ( .A(n15180), .B(n15181), .Z(n14993) );
  XOR2_X1 U15156 ( .A(n15182), .B(n8721), .Z(n15181) );
  XOR2_X1 U15157 ( .A(n15183), .B(n15184), .Z(n14997) );
  XOR2_X1 U15158 ( .A(n15185), .B(n15186), .Z(n15184) );
  XOR2_X1 U15159 ( .A(n9685), .B(n15187), .Z(n9678) );
  XOR2_X1 U15160 ( .A(n9684), .B(n9683), .Z(n15187) );
  OR2_X1 U15161 ( .A1(n8914), .A2(n8923), .ZN(n9683) );
  OR2_X1 U15162 ( .A1(n15188), .A2(n15189), .ZN(n9684) );
  AND2_X1 U15163 ( .A1(n15186), .A2(n15185), .ZN(n15189) );
  AND2_X1 U15164 ( .A1(n15183), .A2(n15190), .ZN(n15188) );
  OR2_X1 U15165 ( .A1(n15185), .A2(n15186), .ZN(n15190) );
  OR2_X1 U15166 ( .A1(n8918), .A2(n8923), .ZN(n15186) );
  OR2_X1 U15167 ( .A1(n15191), .A2(n15192), .ZN(n15185) );
  AND2_X1 U15168 ( .A1(n8721), .A2(n15182), .ZN(n15192) );
  AND2_X1 U15169 ( .A1(n15180), .A2(n15193), .ZN(n15191) );
  OR2_X1 U15170 ( .A1(n15182), .A2(n8721), .ZN(n15193) );
  OR2_X1 U15171 ( .A1(n8922), .A2(n8923), .ZN(n8721) );
  OR2_X1 U15172 ( .A1(n15194), .A2(n15195), .ZN(n15182) );
  AND2_X1 U15173 ( .A1(n15179), .A2(n15178), .ZN(n15195) );
  AND2_X1 U15174 ( .A1(n15176), .A2(n15196), .ZN(n15194) );
  OR2_X1 U15175 ( .A1(n15178), .A2(n15179), .ZN(n15196) );
  OR2_X1 U15176 ( .A1(n8926), .A2(n8923), .ZN(n15179) );
  OR2_X1 U15177 ( .A1(n15197), .A2(n15198), .ZN(n15178) );
  AND2_X1 U15178 ( .A1(n15175), .A2(n15174), .ZN(n15198) );
  AND2_X1 U15179 ( .A1(n15172), .A2(n15199), .ZN(n15197) );
  OR2_X1 U15180 ( .A1(n15174), .A2(n15175), .ZN(n15199) );
  OR2_X1 U15181 ( .A1(n8930), .A2(n8923), .ZN(n15175) );
  OR2_X1 U15182 ( .A1(n15200), .A2(n15201), .ZN(n15174) );
  AND2_X1 U15183 ( .A1(n15171), .A2(n15170), .ZN(n15201) );
  AND2_X1 U15184 ( .A1(n15168), .A2(n15202), .ZN(n15200) );
  OR2_X1 U15185 ( .A1(n15170), .A2(n15171), .ZN(n15202) );
  OR2_X1 U15186 ( .A1(n8934), .A2(n8923), .ZN(n15171) );
  OR2_X1 U15187 ( .A1(n15203), .A2(n15204), .ZN(n15170) );
  AND2_X1 U15188 ( .A1(n15167), .A2(n15166), .ZN(n15204) );
  AND2_X1 U15189 ( .A1(n15164), .A2(n15205), .ZN(n15203) );
  OR2_X1 U15190 ( .A1(n15166), .A2(n15167), .ZN(n15205) );
  OR2_X1 U15191 ( .A1(n8938), .A2(n8923), .ZN(n15167) );
  OR2_X1 U15192 ( .A1(n15206), .A2(n15207), .ZN(n15166) );
  AND2_X1 U15193 ( .A1(n15163), .A2(n15162), .ZN(n15207) );
  AND2_X1 U15194 ( .A1(n15160), .A2(n15208), .ZN(n15206) );
  OR2_X1 U15195 ( .A1(n15162), .A2(n15163), .ZN(n15208) );
  OR2_X1 U15196 ( .A1(n8942), .A2(n8923), .ZN(n15163) );
  OR2_X1 U15197 ( .A1(n15209), .A2(n15210), .ZN(n15162) );
  AND2_X1 U15198 ( .A1(n15159), .A2(n15158), .ZN(n15210) );
  AND2_X1 U15199 ( .A1(n15156), .A2(n15211), .ZN(n15209) );
  OR2_X1 U15200 ( .A1(n15158), .A2(n15159), .ZN(n15211) );
  OR2_X1 U15201 ( .A1(n8946), .A2(n8923), .ZN(n15159) );
  OR2_X1 U15202 ( .A1(n15212), .A2(n15213), .ZN(n15158) );
  AND2_X1 U15203 ( .A1(n15155), .A2(n15154), .ZN(n15213) );
  AND2_X1 U15204 ( .A1(n15152), .A2(n15214), .ZN(n15212) );
  OR2_X1 U15205 ( .A1(n15154), .A2(n15155), .ZN(n15214) );
  OR2_X1 U15206 ( .A1(n8950), .A2(n8923), .ZN(n15155) );
  OR2_X1 U15207 ( .A1(n15215), .A2(n15216), .ZN(n15154) );
  AND2_X1 U15208 ( .A1(n15151), .A2(n15150), .ZN(n15216) );
  AND2_X1 U15209 ( .A1(n15148), .A2(n15217), .ZN(n15215) );
  OR2_X1 U15210 ( .A1(n15150), .A2(n15151), .ZN(n15217) );
  OR2_X1 U15211 ( .A1(n8954), .A2(n8923), .ZN(n15151) );
  OR2_X1 U15212 ( .A1(n15218), .A2(n15219), .ZN(n15150) );
  AND2_X1 U15213 ( .A1(n15147), .A2(n15146), .ZN(n15219) );
  AND2_X1 U15214 ( .A1(n15144), .A2(n15220), .ZN(n15218) );
  OR2_X1 U15215 ( .A1(n15146), .A2(n15147), .ZN(n15220) );
  OR2_X1 U15216 ( .A1(n8958), .A2(n8923), .ZN(n15147) );
  OR2_X1 U15217 ( .A1(n15221), .A2(n15222), .ZN(n15146) );
  AND2_X1 U15218 ( .A1(n15143), .A2(n15142), .ZN(n15222) );
  AND2_X1 U15219 ( .A1(n15140), .A2(n15223), .ZN(n15221) );
  OR2_X1 U15220 ( .A1(n15142), .A2(n15143), .ZN(n15223) );
  OR2_X1 U15221 ( .A1(n8962), .A2(n8923), .ZN(n15143) );
  OR2_X1 U15222 ( .A1(n15224), .A2(n15225), .ZN(n15142) );
  AND2_X1 U15223 ( .A1(n15139), .A2(n15138), .ZN(n15225) );
  AND2_X1 U15224 ( .A1(n15136), .A2(n15226), .ZN(n15224) );
  OR2_X1 U15225 ( .A1(n15138), .A2(n15139), .ZN(n15226) );
  OR2_X1 U15226 ( .A1(n8966), .A2(n8923), .ZN(n15139) );
  OR2_X1 U15227 ( .A1(n15227), .A2(n15228), .ZN(n15138) );
  AND2_X1 U15228 ( .A1(n15135), .A2(n15134), .ZN(n15228) );
  AND2_X1 U15229 ( .A1(n15132), .A2(n15229), .ZN(n15227) );
  OR2_X1 U15230 ( .A1(n15134), .A2(n15135), .ZN(n15229) );
  OR2_X1 U15231 ( .A1(n8970), .A2(n8923), .ZN(n15135) );
  OR2_X1 U15232 ( .A1(n15230), .A2(n15231), .ZN(n15134) );
  AND2_X1 U15233 ( .A1(n15131), .A2(n15130), .ZN(n15231) );
  AND2_X1 U15234 ( .A1(n15128), .A2(n15232), .ZN(n15230) );
  OR2_X1 U15235 ( .A1(n15130), .A2(n15131), .ZN(n15232) );
  OR2_X1 U15236 ( .A1(n8974), .A2(n8923), .ZN(n15131) );
  OR2_X1 U15237 ( .A1(n15233), .A2(n15234), .ZN(n15130) );
  AND2_X1 U15238 ( .A1(n15127), .A2(n15126), .ZN(n15234) );
  AND2_X1 U15239 ( .A1(n15124), .A2(n15235), .ZN(n15233) );
  OR2_X1 U15240 ( .A1(n15126), .A2(n15127), .ZN(n15235) );
  OR2_X1 U15241 ( .A1(n8978), .A2(n8923), .ZN(n15127) );
  OR2_X1 U15242 ( .A1(n15236), .A2(n15237), .ZN(n15126) );
  AND2_X1 U15243 ( .A1(n15123), .A2(n15122), .ZN(n15237) );
  AND2_X1 U15244 ( .A1(n15120), .A2(n15238), .ZN(n15236) );
  OR2_X1 U15245 ( .A1(n15122), .A2(n15123), .ZN(n15238) );
  OR2_X1 U15246 ( .A1(n8982), .A2(n8923), .ZN(n15123) );
  OR2_X1 U15247 ( .A1(n15239), .A2(n15240), .ZN(n15122) );
  AND2_X1 U15248 ( .A1(n15119), .A2(n15118), .ZN(n15240) );
  AND2_X1 U15249 ( .A1(n15116), .A2(n15241), .ZN(n15239) );
  OR2_X1 U15250 ( .A1(n15118), .A2(n15119), .ZN(n15241) );
  OR2_X1 U15251 ( .A1(n8986), .A2(n8923), .ZN(n15119) );
  OR2_X1 U15252 ( .A1(n15242), .A2(n15243), .ZN(n15118) );
  AND2_X1 U15253 ( .A1(n15112), .A2(n15115), .ZN(n15243) );
  AND2_X1 U15254 ( .A1(n15244), .A2(n15114), .ZN(n15242) );
  OR2_X1 U15255 ( .A1(n15245), .A2(n15246), .ZN(n15114) );
  AND2_X1 U15256 ( .A1(n15111), .A2(n15110), .ZN(n15246) );
  AND2_X1 U15257 ( .A1(n15108), .A2(n15247), .ZN(n15245) );
  OR2_X1 U15258 ( .A1(n15110), .A2(n15111), .ZN(n15247) );
  OR2_X1 U15259 ( .A1(n8994), .A2(n8923), .ZN(n15111) );
  OR2_X1 U15260 ( .A1(n15248), .A2(n15249), .ZN(n15110) );
  AND2_X1 U15261 ( .A1(n15104), .A2(n15107), .ZN(n15249) );
  AND2_X1 U15262 ( .A1(n15250), .A2(n15106), .ZN(n15248) );
  OR2_X1 U15263 ( .A1(n15251), .A2(n15252), .ZN(n15106) );
  AND2_X1 U15264 ( .A1(n15100), .A2(n15103), .ZN(n15252) );
  AND2_X1 U15265 ( .A1(n15253), .A2(n15102), .ZN(n15251) );
  OR2_X1 U15266 ( .A1(n15254), .A2(n15255), .ZN(n15102) );
  AND2_X1 U15267 ( .A1(n15097), .A2(n15098), .ZN(n15255) );
  AND2_X1 U15268 ( .A1(n15256), .A2(n15099), .ZN(n15254) );
  OR2_X1 U15269 ( .A1(n15257), .A2(n15258), .ZN(n15099) );
  AND2_X1 U15270 ( .A1(n15092), .A2(n15095), .ZN(n15258) );
  AND2_X1 U15271 ( .A1(n15259), .A2(n15094), .ZN(n15257) );
  OR2_X1 U15272 ( .A1(n15260), .A2(n15261), .ZN(n15094) );
  AND2_X1 U15273 ( .A1(n15089), .A2(n15090), .ZN(n15261) );
  AND2_X1 U15274 ( .A1(n15262), .A2(n15263), .ZN(n15260) );
  OR2_X1 U15275 ( .A1(n15090), .A2(n15089), .ZN(n15263) );
  OR2_X1 U15276 ( .A1(n9014), .A2(n8923), .ZN(n15089) );
  OR2_X1 U15277 ( .A1(n9984), .A2(n15264), .ZN(n15090) );
  OR2_X1 U15278 ( .A1(n8923), .A2(n8919), .ZN(n15264) );
  INV_X1 U15279 ( .A(n15091), .ZN(n15262) );
  OR2_X1 U15280 ( .A1(n15265), .A2(n15266), .ZN(n15091) );
  AND2_X1 U15281 ( .A1(b_5_), .A2(n15267), .ZN(n15266) );
  OR2_X1 U15282 ( .A1(n15268), .A2(n9989), .ZN(n15267) );
  AND2_X1 U15283 ( .A1(a_30_), .A2(n8915), .ZN(n15268) );
  AND2_X1 U15284 ( .A1(b_4_), .A2(n15269), .ZN(n15265) );
  OR2_X1 U15285 ( .A1(n15270), .A2(n8021), .ZN(n15269) );
  AND2_X1 U15286 ( .A1(a_31_), .A2(n8919), .ZN(n15270) );
  OR2_X1 U15287 ( .A1(n15095), .A2(n15092), .ZN(n15259) );
  XOR2_X1 U15288 ( .A(n15271), .B(n15272), .Z(n15092) );
  XNOR2_X1 U15289 ( .A(n15273), .B(n15274), .ZN(n15271) );
  OR2_X1 U15290 ( .A1(n9010), .A2(n8923), .ZN(n15095) );
  OR2_X1 U15291 ( .A1(n15098), .A2(n15097), .ZN(n15256) );
  XOR2_X1 U15292 ( .A(n15275), .B(n15276), .Z(n15097) );
  XOR2_X1 U15293 ( .A(n15277), .B(n15278), .Z(n15276) );
  OR2_X1 U15294 ( .A1(n9006), .A2(n8923), .ZN(n15098) );
  OR2_X1 U15295 ( .A1(n15103), .A2(n15100), .ZN(n15253) );
  XNOR2_X1 U15296 ( .A(n15279), .B(n15280), .ZN(n15100) );
  XNOR2_X1 U15297 ( .A(n15281), .B(n15282), .ZN(n15279) );
  OR2_X1 U15298 ( .A1(n9002), .A2(n8923), .ZN(n15103) );
  OR2_X1 U15299 ( .A1(n15107), .A2(n15104), .ZN(n15250) );
  XOR2_X1 U15300 ( .A(n15283), .B(n15284), .Z(n15104) );
  XOR2_X1 U15301 ( .A(n15285), .B(n15286), .Z(n15284) );
  OR2_X1 U15302 ( .A1(n8998), .A2(n8923), .ZN(n15107) );
  XOR2_X1 U15303 ( .A(n15287), .B(n15288), .Z(n15108) );
  XOR2_X1 U15304 ( .A(n15289), .B(n15290), .Z(n15288) );
  OR2_X1 U15305 ( .A1(n15115), .A2(n15112), .ZN(n15244) );
  XOR2_X1 U15306 ( .A(n15291), .B(n15292), .Z(n15112) );
  XOR2_X1 U15307 ( .A(n15293), .B(n15294), .Z(n15292) );
  OR2_X1 U15308 ( .A1(n8990), .A2(n8923), .ZN(n15115) );
  XOR2_X1 U15309 ( .A(n15295), .B(n15296), .Z(n15116) );
  XOR2_X1 U15310 ( .A(n15297), .B(n15298), .Z(n15296) );
  XOR2_X1 U15311 ( .A(n15299), .B(n15300), .Z(n15120) );
  XOR2_X1 U15312 ( .A(n15301), .B(n15302), .Z(n15300) );
  XOR2_X1 U15313 ( .A(n15303), .B(n15304), .Z(n15124) );
  XOR2_X1 U15314 ( .A(n15305), .B(n15306), .Z(n15304) );
  XOR2_X1 U15315 ( .A(n15307), .B(n15308), .Z(n15128) );
  XOR2_X1 U15316 ( .A(n15309), .B(n15310), .Z(n15308) );
  XOR2_X1 U15317 ( .A(n15311), .B(n15312), .Z(n15132) );
  XOR2_X1 U15318 ( .A(n15313), .B(n15314), .Z(n15312) );
  XOR2_X1 U15319 ( .A(n15315), .B(n15316), .Z(n15136) );
  XOR2_X1 U15320 ( .A(n15317), .B(n15318), .Z(n15316) );
  XOR2_X1 U15321 ( .A(n15319), .B(n15320), .Z(n15140) );
  XOR2_X1 U15322 ( .A(n15321), .B(n15322), .Z(n15320) );
  XOR2_X1 U15323 ( .A(n15323), .B(n15324), .Z(n15144) );
  XOR2_X1 U15324 ( .A(n15325), .B(n15326), .Z(n15324) );
  XOR2_X1 U15325 ( .A(n15327), .B(n15328), .Z(n15148) );
  XOR2_X1 U15326 ( .A(n15329), .B(n15330), .Z(n15328) );
  XOR2_X1 U15327 ( .A(n15331), .B(n15332), .Z(n15152) );
  XOR2_X1 U15328 ( .A(n15333), .B(n15334), .Z(n15332) );
  XOR2_X1 U15329 ( .A(n15335), .B(n15336), .Z(n15156) );
  XOR2_X1 U15330 ( .A(n15337), .B(n15338), .Z(n15336) );
  XOR2_X1 U15331 ( .A(n15339), .B(n15340), .Z(n15160) );
  XOR2_X1 U15332 ( .A(n15341), .B(n15342), .Z(n15340) );
  XOR2_X1 U15333 ( .A(n15343), .B(n15344), .Z(n15164) );
  XOR2_X1 U15334 ( .A(n15345), .B(n15346), .Z(n15344) );
  XOR2_X1 U15335 ( .A(n15347), .B(n15348), .Z(n15168) );
  XOR2_X1 U15336 ( .A(n15349), .B(n15350), .Z(n15348) );
  XOR2_X1 U15337 ( .A(n15351), .B(n15352), .Z(n15172) );
  XOR2_X1 U15338 ( .A(n15353), .B(n15354), .Z(n15352) );
  XOR2_X1 U15339 ( .A(n15355), .B(n15356), .Z(n15176) );
  XOR2_X1 U15340 ( .A(n15357), .B(n15358), .Z(n15356) );
  XOR2_X1 U15341 ( .A(n15359), .B(n15360), .Z(n15180) );
  XOR2_X1 U15342 ( .A(n15361), .B(n15362), .Z(n15360) );
  XOR2_X1 U15343 ( .A(n15363), .B(n15364), .Z(n15183) );
  XOR2_X1 U15344 ( .A(n15365), .B(n15366), .Z(n15364) );
  XOR2_X1 U15345 ( .A(n9691), .B(n15367), .Z(n9685) );
  XOR2_X1 U15346 ( .A(n9690), .B(n8750), .Z(n15367) );
  OR2_X1 U15347 ( .A1(n8918), .A2(n8919), .ZN(n8750) );
  OR2_X1 U15348 ( .A1(n15368), .A2(n15369), .ZN(n9690) );
  AND2_X1 U15349 ( .A1(n15366), .A2(n15365), .ZN(n15369) );
  AND2_X1 U15350 ( .A1(n15363), .A2(n15370), .ZN(n15368) );
  OR2_X1 U15351 ( .A1(n15365), .A2(n15366), .ZN(n15370) );
  OR2_X1 U15352 ( .A1(n8922), .A2(n8919), .ZN(n15366) );
  OR2_X1 U15353 ( .A1(n15371), .A2(n15372), .ZN(n15365) );
  AND2_X1 U15354 ( .A1(n15362), .A2(n15361), .ZN(n15372) );
  AND2_X1 U15355 ( .A1(n15359), .A2(n15373), .ZN(n15371) );
  OR2_X1 U15356 ( .A1(n15361), .A2(n15362), .ZN(n15373) );
  OR2_X1 U15357 ( .A1(n8926), .A2(n8919), .ZN(n15362) );
  OR2_X1 U15358 ( .A1(n15374), .A2(n15375), .ZN(n15361) );
  AND2_X1 U15359 ( .A1(n15358), .A2(n15357), .ZN(n15375) );
  AND2_X1 U15360 ( .A1(n15355), .A2(n15376), .ZN(n15374) );
  OR2_X1 U15361 ( .A1(n15357), .A2(n15358), .ZN(n15376) );
  OR2_X1 U15362 ( .A1(n8930), .A2(n8919), .ZN(n15358) );
  OR2_X1 U15363 ( .A1(n15377), .A2(n15378), .ZN(n15357) );
  AND2_X1 U15364 ( .A1(n15354), .A2(n15353), .ZN(n15378) );
  AND2_X1 U15365 ( .A1(n15351), .A2(n15379), .ZN(n15377) );
  OR2_X1 U15366 ( .A1(n15353), .A2(n15354), .ZN(n15379) );
  OR2_X1 U15367 ( .A1(n8934), .A2(n8919), .ZN(n15354) );
  OR2_X1 U15368 ( .A1(n15380), .A2(n15381), .ZN(n15353) );
  AND2_X1 U15369 ( .A1(n15350), .A2(n15349), .ZN(n15381) );
  AND2_X1 U15370 ( .A1(n15347), .A2(n15382), .ZN(n15380) );
  OR2_X1 U15371 ( .A1(n15349), .A2(n15350), .ZN(n15382) );
  OR2_X1 U15372 ( .A1(n8938), .A2(n8919), .ZN(n15350) );
  OR2_X1 U15373 ( .A1(n15383), .A2(n15384), .ZN(n15349) );
  AND2_X1 U15374 ( .A1(n15346), .A2(n15345), .ZN(n15384) );
  AND2_X1 U15375 ( .A1(n15343), .A2(n15385), .ZN(n15383) );
  OR2_X1 U15376 ( .A1(n15345), .A2(n15346), .ZN(n15385) );
  OR2_X1 U15377 ( .A1(n8942), .A2(n8919), .ZN(n15346) );
  OR2_X1 U15378 ( .A1(n15386), .A2(n15387), .ZN(n15345) );
  AND2_X1 U15379 ( .A1(n15342), .A2(n15341), .ZN(n15387) );
  AND2_X1 U15380 ( .A1(n15339), .A2(n15388), .ZN(n15386) );
  OR2_X1 U15381 ( .A1(n15341), .A2(n15342), .ZN(n15388) );
  OR2_X1 U15382 ( .A1(n8946), .A2(n8919), .ZN(n15342) );
  OR2_X1 U15383 ( .A1(n15389), .A2(n15390), .ZN(n15341) );
  AND2_X1 U15384 ( .A1(n15338), .A2(n15337), .ZN(n15390) );
  AND2_X1 U15385 ( .A1(n15335), .A2(n15391), .ZN(n15389) );
  OR2_X1 U15386 ( .A1(n15337), .A2(n15338), .ZN(n15391) );
  OR2_X1 U15387 ( .A1(n8950), .A2(n8919), .ZN(n15338) );
  OR2_X1 U15388 ( .A1(n15392), .A2(n15393), .ZN(n15337) );
  AND2_X1 U15389 ( .A1(n15334), .A2(n15333), .ZN(n15393) );
  AND2_X1 U15390 ( .A1(n15331), .A2(n15394), .ZN(n15392) );
  OR2_X1 U15391 ( .A1(n15333), .A2(n15334), .ZN(n15394) );
  OR2_X1 U15392 ( .A1(n8954), .A2(n8919), .ZN(n15334) );
  OR2_X1 U15393 ( .A1(n15395), .A2(n15396), .ZN(n15333) );
  AND2_X1 U15394 ( .A1(n15330), .A2(n15329), .ZN(n15396) );
  AND2_X1 U15395 ( .A1(n15327), .A2(n15397), .ZN(n15395) );
  OR2_X1 U15396 ( .A1(n15329), .A2(n15330), .ZN(n15397) );
  OR2_X1 U15397 ( .A1(n8958), .A2(n8919), .ZN(n15330) );
  OR2_X1 U15398 ( .A1(n15398), .A2(n15399), .ZN(n15329) );
  AND2_X1 U15399 ( .A1(n15326), .A2(n15325), .ZN(n15399) );
  AND2_X1 U15400 ( .A1(n15323), .A2(n15400), .ZN(n15398) );
  OR2_X1 U15401 ( .A1(n15325), .A2(n15326), .ZN(n15400) );
  OR2_X1 U15402 ( .A1(n8962), .A2(n8919), .ZN(n15326) );
  OR2_X1 U15403 ( .A1(n15401), .A2(n15402), .ZN(n15325) );
  AND2_X1 U15404 ( .A1(n15322), .A2(n15321), .ZN(n15402) );
  AND2_X1 U15405 ( .A1(n15319), .A2(n15403), .ZN(n15401) );
  OR2_X1 U15406 ( .A1(n15321), .A2(n15322), .ZN(n15403) );
  OR2_X1 U15407 ( .A1(n8966), .A2(n8919), .ZN(n15322) );
  OR2_X1 U15408 ( .A1(n15404), .A2(n15405), .ZN(n15321) );
  AND2_X1 U15409 ( .A1(n15318), .A2(n15317), .ZN(n15405) );
  AND2_X1 U15410 ( .A1(n15315), .A2(n15406), .ZN(n15404) );
  OR2_X1 U15411 ( .A1(n15317), .A2(n15318), .ZN(n15406) );
  OR2_X1 U15412 ( .A1(n8970), .A2(n8919), .ZN(n15318) );
  OR2_X1 U15413 ( .A1(n15407), .A2(n15408), .ZN(n15317) );
  AND2_X1 U15414 ( .A1(n15314), .A2(n15313), .ZN(n15408) );
  AND2_X1 U15415 ( .A1(n15311), .A2(n15409), .ZN(n15407) );
  OR2_X1 U15416 ( .A1(n15313), .A2(n15314), .ZN(n15409) );
  OR2_X1 U15417 ( .A1(n8974), .A2(n8919), .ZN(n15314) );
  OR2_X1 U15418 ( .A1(n15410), .A2(n15411), .ZN(n15313) );
  AND2_X1 U15419 ( .A1(n15310), .A2(n15309), .ZN(n15411) );
  AND2_X1 U15420 ( .A1(n15307), .A2(n15412), .ZN(n15410) );
  OR2_X1 U15421 ( .A1(n15309), .A2(n15310), .ZN(n15412) );
  OR2_X1 U15422 ( .A1(n8978), .A2(n8919), .ZN(n15310) );
  OR2_X1 U15423 ( .A1(n15413), .A2(n15414), .ZN(n15309) );
  AND2_X1 U15424 ( .A1(n15306), .A2(n15305), .ZN(n15414) );
  AND2_X1 U15425 ( .A1(n15303), .A2(n15415), .ZN(n15413) );
  OR2_X1 U15426 ( .A1(n15305), .A2(n15306), .ZN(n15415) );
  OR2_X1 U15427 ( .A1(n8982), .A2(n8919), .ZN(n15306) );
  OR2_X1 U15428 ( .A1(n15416), .A2(n15417), .ZN(n15305) );
  AND2_X1 U15429 ( .A1(n15302), .A2(n15301), .ZN(n15417) );
  AND2_X1 U15430 ( .A1(n15299), .A2(n15418), .ZN(n15416) );
  OR2_X1 U15431 ( .A1(n15301), .A2(n15302), .ZN(n15418) );
  OR2_X1 U15432 ( .A1(n8986), .A2(n8919), .ZN(n15302) );
  OR2_X1 U15433 ( .A1(n15419), .A2(n15420), .ZN(n15301) );
  AND2_X1 U15434 ( .A1(n15298), .A2(n15297), .ZN(n15420) );
  AND2_X1 U15435 ( .A1(n15295), .A2(n15421), .ZN(n15419) );
  OR2_X1 U15436 ( .A1(n15297), .A2(n15298), .ZN(n15421) );
  OR2_X1 U15437 ( .A1(n8990), .A2(n8919), .ZN(n15298) );
  OR2_X1 U15438 ( .A1(n15422), .A2(n15423), .ZN(n15297) );
  AND2_X1 U15439 ( .A1(n15291), .A2(n15294), .ZN(n15423) );
  AND2_X1 U15440 ( .A1(n15424), .A2(n15293), .ZN(n15422) );
  OR2_X1 U15441 ( .A1(n15425), .A2(n15426), .ZN(n15293) );
  AND2_X1 U15442 ( .A1(n15290), .A2(n15289), .ZN(n15426) );
  AND2_X1 U15443 ( .A1(n15287), .A2(n15427), .ZN(n15425) );
  OR2_X1 U15444 ( .A1(n15289), .A2(n15290), .ZN(n15427) );
  OR2_X1 U15445 ( .A1(n8998), .A2(n8919), .ZN(n15290) );
  OR2_X1 U15446 ( .A1(n15428), .A2(n15429), .ZN(n15289) );
  AND2_X1 U15447 ( .A1(n15283), .A2(n15286), .ZN(n15429) );
  AND2_X1 U15448 ( .A1(n15430), .A2(n15285), .ZN(n15428) );
  OR2_X1 U15449 ( .A1(n15431), .A2(n15432), .ZN(n15285) );
  AND2_X1 U15450 ( .A1(n15280), .A2(n15281), .ZN(n15432) );
  AND2_X1 U15451 ( .A1(n15433), .A2(n15282), .ZN(n15431) );
  OR2_X1 U15452 ( .A1(n15434), .A2(n15435), .ZN(n15282) );
  AND2_X1 U15453 ( .A1(n15275), .A2(n15278), .ZN(n15435) );
  AND2_X1 U15454 ( .A1(n15436), .A2(n15277), .ZN(n15434) );
  OR2_X1 U15455 ( .A1(n15437), .A2(n15438), .ZN(n15277) );
  AND2_X1 U15456 ( .A1(n15272), .A2(n15273), .ZN(n15438) );
  AND2_X1 U15457 ( .A1(n15439), .A2(n15440), .ZN(n15437) );
  OR2_X1 U15458 ( .A1(n15273), .A2(n15272), .ZN(n15440) );
  OR2_X1 U15459 ( .A1(n9014), .A2(n8919), .ZN(n15272) );
  OR2_X1 U15460 ( .A1(n9984), .A2(n15441), .ZN(n15273) );
  OR2_X1 U15461 ( .A1(n8919), .A2(n8915), .ZN(n15441) );
  INV_X1 U15462 ( .A(n15274), .ZN(n15439) );
  OR2_X1 U15463 ( .A1(n15442), .A2(n15443), .ZN(n15274) );
  AND2_X1 U15464 ( .A1(b_4_), .A2(n15444), .ZN(n15443) );
  OR2_X1 U15465 ( .A1(n15445), .A2(n9989), .ZN(n15444) );
  AND2_X1 U15466 ( .A1(a_30_), .A2(n8911), .ZN(n15445) );
  AND2_X1 U15467 ( .A1(b_3_), .A2(n15446), .ZN(n15442) );
  OR2_X1 U15468 ( .A1(n15447), .A2(n8021), .ZN(n15446) );
  AND2_X1 U15469 ( .A1(a_31_), .A2(n8915), .ZN(n15447) );
  OR2_X1 U15470 ( .A1(n15278), .A2(n15275), .ZN(n15436) );
  XOR2_X1 U15471 ( .A(n15448), .B(n15449), .Z(n15275) );
  XNOR2_X1 U15472 ( .A(n15450), .B(n15451), .ZN(n15448) );
  OR2_X1 U15473 ( .A1(n9010), .A2(n8919), .ZN(n15278) );
  OR2_X1 U15474 ( .A1(n15281), .A2(n15280), .ZN(n15433) );
  XOR2_X1 U15475 ( .A(n15452), .B(n15453), .Z(n15280) );
  XOR2_X1 U15476 ( .A(n15454), .B(n15455), .Z(n15453) );
  OR2_X1 U15477 ( .A1(n9006), .A2(n8919), .ZN(n15281) );
  OR2_X1 U15478 ( .A1(n15286), .A2(n15283), .ZN(n15430) );
  XNOR2_X1 U15479 ( .A(n15456), .B(n15457), .ZN(n15283) );
  XNOR2_X1 U15480 ( .A(n15458), .B(n15459), .ZN(n15456) );
  OR2_X1 U15481 ( .A1(n9002), .A2(n8919), .ZN(n15286) );
  XOR2_X1 U15482 ( .A(n15460), .B(n15461), .Z(n15287) );
  XOR2_X1 U15483 ( .A(n15462), .B(n15463), .Z(n15461) );
  OR2_X1 U15484 ( .A1(n15294), .A2(n15291), .ZN(n15424) );
  XOR2_X1 U15485 ( .A(n15464), .B(n15465), .Z(n15291) );
  XOR2_X1 U15486 ( .A(n15466), .B(n15467), .Z(n15465) );
  OR2_X1 U15487 ( .A1(n8994), .A2(n8919), .ZN(n15294) );
  XOR2_X1 U15488 ( .A(n15468), .B(n15469), .Z(n15295) );
  XOR2_X1 U15489 ( .A(n15470), .B(n15471), .Z(n15469) );
  XOR2_X1 U15490 ( .A(n15472), .B(n15473), .Z(n15299) );
  XOR2_X1 U15491 ( .A(n15474), .B(n15475), .Z(n15473) );
  XOR2_X1 U15492 ( .A(n15476), .B(n15477), .Z(n15303) );
  XOR2_X1 U15493 ( .A(n15478), .B(n15479), .Z(n15477) );
  XOR2_X1 U15494 ( .A(n15480), .B(n15481), .Z(n15307) );
  XOR2_X1 U15495 ( .A(n15482), .B(n15483), .Z(n15481) );
  XOR2_X1 U15496 ( .A(n15484), .B(n15485), .Z(n15311) );
  XOR2_X1 U15497 ( .A(n15486), .B(n15487), .Z(n15485) );
  XOR2_X1 U15498 ( .A(n15488), .B(n15489), .Z(n15315) );
  XOR2_X1 U15499 ( .A(n15490), .B(n15491), .Z(n15489) );
  XOR2_X1 U15500 ( .A(n15492), .B(n15493), .Z(n15319) );
  XOR2_X1 U15501 ( .A(n15494), .B(n15495), .Z(n15493) );
  XOR2_X1 U15502 ( .A(n15496), .B(n15497), .Z(n15323) );
  XOR2_X1 U15503 ( .A(n15498), .B(n15499), .Z(n15497) );
  XOR2_X1 U15504 ( .A(n15500), .B(n15501), .Z(n15327) );
  XOR2_X1 U15505 ( .A(n15502), .B(n15503), .Z(n15501) );
  XOR2_X1 U15506 ( .A(n15504), .B(n15505), .Z(n15331) );
  XOR2_X1 U15507 ( .A(n15506), .B(n15507), .Z(n15505) );
  XOR2_X1 U15508 ( .A(n15508), .B(n15509), .Z(n15335) );
  XOR2_X1 U15509 ( .A(n15510), .B(n15511), .Z(n15509) );
  XOR2_X1 U15510 ( .A(n15512), .B(n15513), .Z(n15339) );
  XOR2_X1 U15511 ( .A(n15514), .B(n15515), .Z(n15513) );
  XOR2_X1 U15512 ( .A(n15516), .B(n15517), .Z(n15343) );
  XOR2_X1 U15513 ( .A(n15518), .B(n15519), .Z(n15517) );
  XOR2_X1 U15514 ( .A(n15520), .B(n15521), .Z(n15347) );
  XOR2_X1 U15515 ( .A(n15522), .B(n15523), .Z(n15521) );
  XOR2_X1 U15516 ( .A(n15524), .B(n15525), .Z(n15351) );
  XOR2_X1 U15517 ( .A(n15526), .B(n15527), .Z(n15525) );
  XOR2_X1 U15518 ( .A(n15528), .B(n15529), .Z(n15355) );
  XOR2_X1 U15519 ( .A(n15530), .B(n15531), .Z(n15529) );
  XOR2_X1 U15520 ( .A(n15532), .B(n15533), .Z(n15359) );
  XOR2_X1 U15521 ( .A(n15534), .B(n15535), .Z(n15533) );
  XOR2_X1 U15522 ( .A(n15536), .B(n15537), .Z(n15363) );
  XOR2_X1 U15523 ( .A(n15538), .B(n15539), .Z(n15537) );
  XOR2_X1 U15524 ( .A(n9698), .B(n15540), .Z(n9691) );
  XOR2_X1 U15525 ( .A(n9697), .B(n9696), .Z(n15540) );
  OR2_X1 U15526 ( .A1(n8922), .A2(n8915), .ZN(n9696) );
  OR2_X1 U15527 ( .A1(n15541), .A2(n15542), .ZN(n9697) );
  AND2_X1 U15528 ( .A1(n15539), .A2(n15538), .ZN(n15542) );
  AND2_X1 U15529 ( .A1(n15536), .A2(n15543), .ZN(n15541) );
  OR2_X1 U15530 ( .A1(n15538), .A2(n15539), .ZN(n15543) );
  OR2_X1 U15531 ( .A1(n8926), .A2(n8915), .ZN(n15539) );
  OR2_X1 U15532 ( .A1(n15544), .A2(n15545), .ZN(n15538) );
  AND2_X1 U15533 ( .A1(n15535), .A2(n15534), .ZN(n15545) );
  AND2_X1 U15534 ( .A1(n15532), .A2(n15546), .ZN(n15544) );
  OR2_X1 U15535 ( .A1(n15534), .A2(n15535), .ZN(n15546) );
  OR2_X1 U15536 ( .A1(n8930), .A2(n8915), .ZN(n15535) );
  OR2_X1 U15537 ( .A1(n15547), .A2(n15548), .ZN(n15534) );
  AND2_X1 U15538 ( .A1(n15531), .A2(n15530), .ZN(n15548) );
  AND2_X1 U15539 ( .A1(n15528), .A2(n15549), .ZN(n15547) );
  OR2_X1 U15540 ( .A1(n15530), .A2(n15531), .ZN(n15549) );
  OR2_X1 U15541 ( .A1(n8934), .A2(n8915), .ZN(n15531) );
  OR2_X1 U15542 ( .A1(n15550), .A2(n15551), .ZN(n15530) );
  AND2_X1 U15543 ( .A1(n15527), .A2(n15526), .ZN(n15551) );
  AND2_X1 U15544 ( .A1(n15524), .A2(n15552), .ZN(n15550) );
  OR2_X1 U15545 ( .A1(n15526), .A2(n15527), .ZN(n15552) );
  OR2_X1 U15546 ( .A1(n8938), .A2(n8915), .ZN(n15527) );
  OR2_X1 U15547 ( .A1(n15553), .A2(n15554), .ZN(n15526) );
  AND2_X1 U15548 ( .A1(n15523), .A2(n15522), .ZN(n15554) );
  AND2_X1 U15549 ( .A1(n15520), .A2(n15555), .ZN(n15553) );
  OR2_X1 U15550 ( .A1(n15522), .A2(n15523), .ZN(n15555) );
  OR2_X1 U15551 ( .A1(n8942), .A2(n8915), .ZN(n15523) );
  OR2_X1 U15552 ( .A1(n15556), .A2(n15557), .ZN(n15522) );
  AND2_X1 U15553 ( .A1(n15519), .A2(n15518), .ZN(n15557) );
  AND2_X1 U15554 ( .A1(n15516), .A2(n15558), .ZN(n15556) );
  OR2_X1 U15555 ( .A1(n15518), .A2(n15519), .ZN(n15558) );
  OR2_X1 U15556 ( .A1(n8946), .A2(n8915), .ZN(n15519) );
  OR2_X1 U15557 ( .A1(n15559), .A2(n15560), .ZN(n15518) );
  AND2_X1 U15558 ( .A1(n15515), .A2(n15514), .ZN(n15560) );
  AND2_X1 U15559 ( .A1(n15512), .A2(n15561), .ZN(n15559) );
  OR2_X1 U15560 ( .A1(n15514), .A2(n15515), .ZN(n15561) );
  OR2_X1 U15561 ( .A1(n8950), .A2(n8915), .ZN(n15515) );
  OR2_X1 U15562 ( .A1(n15562), .A2(n15563), .ZN(n15514) );
  AND2_X1 U15563 ( .A1(n15511), .A2(n15510), .ZN(n15563) );
  AND2_X1 U15564 ( .A1(n15508), .A2(n15564), .ZN(n15562) );
  OR2_X1 U15565 ( .A1(n15510), .A2(n15511), .ZN(n15564) );
  OR2_X1 U15566 ( .A1(n8954), .A2(n8915), .ZN(n15511) );
  OR2_X1 U15567 ( .A1(n15565), .A2(n15566), .ZN(n15510) );
  AND2_X1 U15568 ( .A1(n15507), .A2(n15506), .ZN(n15566) );
  AND2_X1 U15569 ( .A1(n15504), .A2(n15567), .ZN(n15565) );
  OR2_X1 U15570 ( .A1(n15506), .A2(n15507), .ZN(n15567) );
  OR2_X1 U15571 ( .A1(n8958), .A2(n8915), .ZN(n15507) );
  OR2_X1 U15572 ( .A1(n15568), .A2(n15569), .ZN(n15506) );
  AND2_X1 U15573 ( .A1(n15503), .A2(n15502), .ZN(n15569) );
  AND2_X1 U15574 ( .A1(n15500), .A2(n15570), .ZN(n15568) );
  OR2_X1 U15575 ( .A1(n15502), .A2(n15503), .ZN(n15570) );
  OR2_X1 U15576 ( .A1(n8962), .A2(n8915), .ZN(n15503) );
  OR2_X1 U15577 ( .A1(n15571), .A2(n15572), .ZN(n15502) );
  AND2_X1 U15578 ( .A1(n15499), .A2(n15498), .ZN(n15572) );
  AND2_X1 U15579 ( .A1(n15496), .A2(n15573), .ZN(n15571) );
  OR2_X1 U15580 ( .A1(n15498), .A2(n15499), .ZN(n15573) );
  OR2_X1 U15581 ( .A1(n8966), .A2(n8915), .ZN(n15499) );
  OR2_X1 U15582 ( .A1(n15574), .A2(n15575), .ZN(n15498) );
  AND2_X1 U15583 ( .A1(n15495), .A2(n15494), .ZN(n15575) );
  AND2_X1 U15584 ( .A1(n15492), .A2(n15576), .ZN(n15574) );
  OR2_X1 U15585 ( .A1(n15494), .A2(n15495), .ZN(n15576) );
  OR2_X1 U15586 ( .A1(n8970), .A2(n8915), .ZN(n15495) );
  OR2_X1 U15587 ( .A1(n15577), .A2(n15578), .ZN(n15494) );
  AND2_X1 U15588 ( .A1(n15491), .A2(n15490), .ZN(n15578) );
  AND2_X1 U15589 ( .A1(n15488), .A2(n15579), .ZN(n15577) );
  OR2_X1 U15590 ( .A1(n15490), .A2(n15491), .ZN(n15579) );
  OR2_X1 U15591 ( .A1(n8974), .A2(n8915), .ZN(n15491) );
  OR2_X1 U15592 ( .A1(n15580), .A2(n15581), .ZN(n15490) );
  AND2_X1 U15593 ( .A1(n15487), .A2(n15486), .ZN(n15581) );
  AND2_X1 U15594 ( .A1(n15484), .A2(n15582), .ZN(n15580) );
  OR2_X1 U15595 ( .A1(n15486), .A2(n15487), .ZN(n15582) );
  OR2_X1 U15596 ( .A1(n8978), .A2(n8915), .ZN(n15487) );
  OR2_X1 U15597 ( .A1(n15583), .A2(n15584), .ZN(n15486) );
  AND2_X1 U15598 ( .A1(n15483), .A2(n15482), .ZN(n15584) );
  AND2_X1 U15599 ( .A1(n15480), .A2(n15585), .ZN(n15583) );
  OR2_X1 U15600 ( .A1(n15482), .A2(n15483), .ZN(n15585) );
  OR2_X1 U15601 ( .A1(n8982), .A2(n8915), .ZN(n15483) );
  OR2_X1 U15602 ( .A1(n15586), .A2(n15587), .ZN(n15482) );
  AND2_X1 U15603 ( .A1(n15479), .A2(n15478), .ZN(n15587) );
  AND2_X1 U15604 ( .A1(n15476), .A2(n15588), .ZN(n15586) );
  OR2_X1 U15605 ( .A1(n15478), .A2(n15479), .ZN(n15588) );
  OR2_X1 U15606 ( .A1(n8986), .A2(n8915), .ZN(n15479) );
  OR2_X1 U15607 ( .A1(n15589), .A2(n15590), .ZN(n15478) );
  AND2_X1 U15608 ( .A1(n15475), .A2(n15474), .ZN(n15590) );
  AND2_X1 U15609 ( .A1(n15472), .A2(n15591), .ZN(n15589) );
  OR2_X1 U15610 ( .A1(n15474), .A2(n15475), .ZN(n15591) );
  OR2_X1 U15611 ( .A1(n8990), .A2(n8915), .ZN(n15475) );
  OR2_X1 U15612 ( .A1(n15592), .A2(n15593), .ZN(n15474) );
  AND2_X1 U15613 ( .A1(n15471), .A2(n15470), .ZN(n15593) );
  AND2_X1 U15614 ( .A1(n15468), .A2(n15594), .ZN(n15592) );
  OR2_X1 U15615 ( .A1(n15470), .A2(n15471), .ZN(n15594) );
  OR2_X1 U15616 ( .A1(n8994), .A2(n8915), .ZN(n15471) );
  OR2_X1 U15617 ( .A1(n15595), .A2(n15596), .ZN(n15470) );
  AND2_X1 U15618 ( .A1(n15464), .A2(n15467), .ZN(n15596) );
  AND2_X1 U15619 ( .A1(n15597), .A2(n15466), .ZN(n15595) );
  OR2_X1 U15620 ( .A1(n15598), .A2(n15599), .ZN(n15466) );
  AND2_X1 U15621 ( .A1(n15463), .A2(n15462), .ZN(n15599) );
  AND2_X1 U15622 ( .A1(n15460), .A2(n15600), .ZN(n15598) );
  OR2_X1 U15623 ( .A1(n15462), .A2(n15463), .ZN(n15600) );
  OR2_X1 U15624 ( .A1(n9002), .A2(n8915), .ZN(n15463) );
  OR2_X1 U15625 ( .A1(n15601), .A2(n15602), .ZN(n15462) );
  AND2_X1 U15626 ( .A1(n15457), .A2(n15458), .ZN(n15602) );
  AND2_X1 U15627 ( .A1(n15603), .A2(n15459), .ZN(n15601) );
  OR2_X1 U15628 ( .A1(n15604), .A2(n15605), .ZN(n15459) );
  AND2_X1 U15629 ( .A1(n15452), .A2(n15455), .ZN(n15605) );
  AND2_X1 U15630 ( .A1(n15606), .A2(n15454), .ZN(n15604) );
  OR2_X1 U15631 ( .A1(n15607), .A2(n15608), .ZN(n15454) );
  AND2_X1 U15632 ( .A1(n15449), .A2(n15450), .ZN(n15608) );
  AND2_X1 U15633 ( .A1(n15609), .A2(n15610), .ZN(n15607) );
  OR2_X1 U15634 ( .A1(n15450), .A2(n15449), .ZN(n15610) );
  OR2_X1 U15635 ( .A1(n9014), .A2(n8915), .ZN(n15449) );
  OR2_X1 U15636 ( .A1(n9984), .A2(n15611), .ZN(n15450) );
  OR2_X1 U15637 ( .A1(n8915), .A2(n8911), .ZN(n15611) );
  INV_X1 U15638 ( .A(n15451), .ZN(n15609) );
  OR2_X1 U15639 ( .A1(n15612), .A2(n15613), .ZN(n15451) );
  AND2_X1 U15640 ( .A1(b_3_), .A2(n15614), .ZN(n15613) );
  OR2_X1 U15641 ( .A1(n15615), .A2(n9989), .ZN(n15614) );
  AND2_X1 U15642 ( .A1(a_30_), .A2(n8907), .ZN(n15615) );
  AND2_X1 U15643 ( .A1(b_2_), .A2(n15616), .ZN(n15612) );
  OR2_X1 U15644 ( .A1(n15617), .A2(n8021), .ZN(n15616) );
  AND2_X1 U15645 ( .A1(a_31_), .A2(n8911), .ZN(n15617) );
  OR2_X1 U15646 ( .A1(n15455), .A2(n15452), .ZN(n15606) );
  XOR2_X1 U15647 ( .A(n15618), .B(n15619), .Z(n15452) );
  XNOR2_X1 U15648 ( .A(n15620), .B(n15621), .ZN(n15618) );
  OR2_X1 U15649 ( .A1(n9010), .A2(n8915), .ZN(n15455) );
  OR2_X1 U15650 ( .A1(n15458), .A2(n15457), .ZN(n15603) );
  XOR2_X1 U15651 ( .A(n15622), .B(n15623), .Z(n15457) );
  XOR2_X1 U15652 ( .A(n15624), .B(n15625), .Z(n15623) );
  OR2_X1 U15653 ( .A1(n9006), .A2(n8915), .ZN(n15458) );
  XNOR2_X1 U15654 ( .A(n15626), .B(n15627), .ZN(n15460) );
  XNOR2_X1 U15655 ( .A(n15628), .B(n15629), .ZN(n15626) );
  OR2_X1 U15656 ( .A1(n15467), .A2(n15464), .ZN(n15597) );
  XOR2_X1 U15657 ( .A(n15630), .B(n15631), .Z(n15464) );
  XOR2_X1 U15658 ( .A(n15632), .B(n15633), .Z(n15631) );
  OR2_X1 U15659 ( .A1(n8998), .A2(n8915), .ZN(n15467) );
  XOR2_X1 U15660 ( .A(n15634), .B(n15635), .Z(n15468) );
  XOR2_X1 U15661 ( .A(n15636), .B(n15637), .Z(n15635) );
  XOR2_X1 U15662 ( .A(n15638), .B(n15639), .Z(n15472) );
  XOR2_X1 U15663 ( .A(n15640), .B(n15641), .Z(n15639) );
  XOR2_X1 U15664 ( .A(n15642), .B(n15643), .Z(n15476) );
  XOR2_X1 U15665 ( .A(n15644), .B(n15645), .Z(n15643) );
  XOR2_X1 U15666 ( .A(n15646), .B(n15647), .Z(n15480) );
  XOR2_X1 U15667 ( .A(n15648), .B(n15649), .Z(n15647) );
  XOR2_X1 U15668 ( .A(n15650), .B(n15651), .Z(n15484) );
  XOR2_X1 U15669 ( .A(n15652), .B(n15653), .Z(n15651) );
  XOR2_X1 U15670 ( .A(n15654), .B(n15655), .Z(n15488) );
  XOR2_X1 U15671 ( .A(n15656), .B(n15657), .Z(n15655) );
  XOR2_X1 U15672 ( .A(n15658), .B(n15659), .Z(n15492) );
  XOR2_X1 U15673 ( .A(n15660), .B(n15661), .Z(n15659) );
  XOR2_X1 U15674 ( .A(n15662), .B(n15663), .Z(n15496) );
  XOR2_X1 U15675 ( .A(n15664), .B(n15665), .Z(n15663) );
  XOR2_X1 U15676 ( .A(n15666), .B(n15667), .Z(n15500) );
  XOR2_X1 U15677 ( .A(n15668), .B(n15669), .Z(n15667) );
  XOR2_X1 U15678 ( .A(n15670), .B(n15671), .Z(n15504) );
  XOR2_X1 U15679 ( .A(n15672), .B(n15673), .Z(n15671) );
  XOR2_X1 U15680 ( .A(n15674), .B(n15675), .Z(n15508) );
  XOR2_X1 U15681 ( .A(n15676), .B(n15677), .Z(n15675) );
  XOR2_X1 U15682 ( .A(n15678), .B(n15679), .Z(n15512) );
  XOR2_X1 U15683 ( .A(n15680), .B(n15681), .Z(n15679) );
  XOR2_X1 U15684 ( .A(n15682), .B(n15683), .Z(n15516) );
  XOR2_X1 U15685 ( .A(n15684), .B(n15685), .Z(n15683) );
  XOR2_X1 U15686 ( .A(n15686), .B(n15687), .Z(n15520) );
  XOR2_X1 U15687 ( .A(n15688), .B(n15689), .Z(n15687) );
  XOR2_X1 U15688 ( .A(n15690), .B(n15691), .Z(n15524) );
  XOR2_X1 U15689 ( .A(n15692), .B(n15693), .Z(n15691) );
  XOR2_X1 U15690 ( .A(n15694), .B(n15695), .Z(n15528) );
  XOR2_X1 U15691 ( .A(n15696), .B(n15697), .Z(n15695) );
  XOR2_X1 U15692 ( .A(n15698), .B(n15699), .Z(n15532) );
  XOR2_X1 U15693 ( .A(n15700), .B(n15701), .Z(n15699) );
  XOR2_X1 U15694 ( .A(n15702), .B(n15703), .Z(n15536) );
  XOR2_X1 U15695 ( .A(n15704), .B(n15705), .Z(n15703) );
  XOR2_X1 U15696 ( .A(n9705), .B(n15706), .Z(n9698) );
  XOR2_X1 U15697 ( .A(n9704), .B(n9703), .Z(n15706) );
  OR2_X1 U15698 ( .A1(n8926), .A2(n8911), .ZN(n9703) );
  OR2_X1 U15699 ( .A1(n15707), .A2(n15708), .ZN(n9704) );
  AND2_X1 U15700 ( .A1(n15705), .A2(n15704), .ZN(n15708) );
  AND2_X1 U15701 ( .A1(n15702), .A2(n15709), .ZN(n15707) );
  OR2_X1 U15702 ( .A1(n15704), .A2(n15705), .ZN(n15709) );
  OR2_X1 U15703 ( .A1(n8930), .A2(n8911), .ZN(n15705) );
  OR2_X1 U15704 ( .A1(n15710), .A2(n15711), .ZN(n15704) );
  AND2_X1 U15705 ( .A1(n15701), .A2(n15700), .ZN(n15711) );
  AND2_X1 U15706 ( .A1(n15698), .A2(n15712), .ZN(n15710) );
  OR2_X1 U15707 ( .A1(n15700), .A2(n15701), .ZN(n15712) );
  OR2_X1 U15708 ( .A1(n8934), .A2(n8911), .ZN(n15701) );
  OR2_X1 U15709 ( .A1(n15713), .A2(n15714), .ZN(n15700) );
  AND2_X1 U15710 ( .A1(n15697), .A2(n15696), .ZN(n15714) );
  AND2_X1 U15711 ( .A1(n15694), .A2(n15715), .ZN(n15713) );
  OR2_X1 U15712 ( .A1(n15696), .A2(n15697), .ZN(n15715) );
  OR2_X1 U15713 ( .A1(n8938), .A2(n8911), .ZN(n15697) );
  OR2_X1 U15714 ( .A1(n15716), .A2(n15717), .ZN(n15696) );
  AND2_X1 U15715 ( .A1(n15693), .A2(n15692), .ZN(n15717) );
  AND2_X1 U15716 ( .A1(n15690), .A2(n15718), .ZN(n15716) );
  OR2_X1 U15717 ( .A1(n15692), .A2(n15693), .ZN(n15718) );
  OR2_X1 U15718 ( .A1(n8942), .A2(n8911), .ZN(n15693) );
  OR2_X1 U15719 ( .A1(n15719), .A2(n15720), .ZN(n15692) );
  AND2_X1 U15720 ( .A1(n15689), .A2(n15688), .ZN(n15720) );
  AND2_X1 U15721 ( .A1(n15686), .A2(n15721), .ZN(n15719) );
  OR2_X1 U15722 ( .A1(n15688), .A2(n15689), .ZN(n15721) );
  OR2_X1 U15723 ( .A1(n8946), .A2(n8911), .ZN(n15689) );
  OR2_X1 U15724 ( .A1(n15722), .A2(n15723), .ZN(n15688) );
  AND2_X1 U15725 ( .A1(n15685), .A2(n15684), .ZN(n15723) );
  AND2_X1 U15726 ( .A1(n15682), .A2(n15724), .ZN(n15722) );
  OR2_X1 U15727 ( .A1(n15684), .A2(n15685), .ZN(n15724) );
  OR2_X1 U15728 ( .A1(n8950), .A2(n8911), .ZN(n15685) );
  OR2_X1 U15729 ( .A1(n15725), .A2(n15726), .ZN(n15684) );
  AND2_X1 U15730 ( .A1(n15681), .A2(n15680), .ZN(n15726) );
  AND2_X1 U15731 ( .A1(n15678), .A2(n15727), .ZN(n15725) );
  OR2_X1 U15732 ( .A1(n15680), .A2(n15681), .ZN(n15727) );
  OR2_X1 U15733 ( .A1(n8954), .A2(n8911), .ZN(n15681) );
  OR2_X1 U15734 ( .A1(n15728), .A2(n15729), .ZN(n15680) );
  AND2_X1 U15735 ( .A1(n15677), .A2(n15676), .ZN(n15729) );
  AND2_X1 U15736 ( .A1(n15674), .A2(n15730), .ZN(n15728) );
  OR2_X1 U15737 ( .A1(n15676), .A2(n15677), .ZN(n15730) );
  OR2_X1 U15738 ( .A1(n8958), .A2(n8911), .ZN(n15677) );
  OR2_X1 U15739 ( .A1(n15731), .A2(n15732), .ZN(n15676) );
  AND2_X1 U15740 ( .A1(n15673), .A2(n15672), .ZN(n15732) );
  AND2_X1 U15741 ( .A1(n15670), .A2(n15733), .ZN(n15731) );
  OR2_X1 U15742 ( .A1(n15672), .A2(n15673), .ZN(n15733) );
  OR2_X1 U15743 ( .A1(n8962), .A2(n8911), .ZN(n15673) );
  OR2_X1 U15744 ( .A1(n15734), .A2(n15735), .ZN(n15672) );
  AND2_X1 U15745 ( .A1(n15669), .A2(n15668), .ZN(n15735) );
  AND2_X1 U15746 ( .A1(n15666), .A2(n15736), .ZN(n15734) );
  OR2_X1 U15747 ( .A1(n15668), .A2(n15669), .ZN(n15736) );
  OR2_X1 U15748 ( .A1(n8966), .A2(n8911), .ZN(n15669) );
  OR2_X1 U15749 ( .A1(n15737), .A2(n15738), .ZN(n15668) );
  AND2_X1 U15750 ( .A1(n15665), .A2(n15664), .ZN(n15738) );
  AND2_X1 U15751 ( .A1(n15662), .A2(n15739), .ZN(n15737) );
  OR2_X1 U15752 ( .A1(n15664), .A2(n15665), .ZN(n15739) );
  OR2_X1 U15753 ( .A1(n8970), .A2(n8911), .ZN(n15665) );
  OR2_X1 U15754 ( .A1(n15740), .A2(n15741), .ZN(n15664) );
  AND2_X1 U15755 ( .A1(n15661), .A2(n15660), .ZN(n15741) );
  AND2_X1 U15756 ( .A1(n15658), .A2(n15742), .ZN(n15740) );
  OR2_X1 U15757 ( .A1(n15660), .A2(n15661), .ZN(n15742) );
  OR2_X1 U15758 ( .A1(n8974), .A2(n8911), .ZN(n15661) );
  OR2_X1 U15759 ( .A1(n15743), .A2(n15744), .ZN(n15660) );
  AND2_X1 U15760 ( .A1(n15657), .A2(n15656), .ZN(n15744) );
  AND2_X1 U15761 ( .A1(n15654), .A2(n15745), .ZN(n15743) );
  OR2_X1 U15762 ( .A1(n15656), .A2(n15657), .ZN(n15745) );
  OR2_X1 U15763 ( .A1(n8978), .A2(n8911), .ZN(n15657) );
  OR2_X1 U15764 ( .A1(n15746), .A2(n15747), .ZN(n15656) );
  AND2_X1 U15765 ( .A1(n15653), .A2(n15652), .ZN(n15747) );
  AND2_X1 U15766 ( .A1(n15650), .A2(n15748), .ZN(n15746) );
  OR2_X1 U15767 ( .A1(n15652), .A2(n15653), .ZN(n15748) );
  OR2_X1 U15768 ( .A1(n8982), .A2(n8911), .ZN(n15653) );
  OR2_X1 U15769 ( .A1(n15749), .A2(n15750), .ZN(n15652) );
  AND2_X1 U15770 ( .A1(n15649), .A2(n15648), .ZN(n15750) );
  AND2_X1 U15771 ( .A1(n15646), .A2(n15751), .ZN(n15749) );
  OR2_X1 U15772 ( .A1(n15648), .A2(n15649), .ZN(n15751) );
  OR2_X1 U15773 ( .A1(n8986), .A2(n8911), .ZN(n15649) );
  OR2_X1 U15774 ( .A1(n15752), .A2(n15753), .ZN(n15648) );
  AND2_X1 U15775 ( .A1(n15645), .A2(n15644), .ZN(n15753) );
  AND2_X1 U15776 ( .A1(n15642), .A2(n15754), .ZN(n15752) );
  OR2_X1 U15777 ( .A1(n15644), .A2(n15645), .ZN(n15754) );
  OR2_X1 U15778 ( .A1(n8990), .A2(n8911), .ZN(n15645) );
  OR2_X1 U15779 ( .A1(n15755), .A2(n15756), .ZN(n15644) );
  AND2_X1 U15780 ( .A1(n15641), .A2(n15640), .ZN(n15756) );
  AND2_X1 U15781 ( .A1(n15638), .A2(n15757), .ZN(n15755) );
  OR2_X1 U15782 ( .A1(n15640), .A2(n15641), .ZN(n15757) );
  OR2_X1 U15783 ( .A1(n8994), .A2(n8911), .ZN(n15641) );
  OR2_X1 U15784 ( .A1(n15758), .A2(n15759), .ZN(n15640) );
  AND2_X1 U15785 ( .A1(n15637), .A2(n15636), .ZN(n15759) );
  AND2_X1 U15786 ( .A1(n15634), .A2(n15760), .ZN(n15758) );
  OR2_X1 U15787 ( .A1(n15636), .A2(n15637), .ZN(n15760) );
  OR2_X1 U15788 ( .A1(n8998), .A2(n8911), .ZN(n15637) );
  OR2_X1 U15789 ( .A1(n15761), .A2(n15762), .ZN(n15636) );
  AND2_X1 U15790 ( .A1(n15630), .A2(n15633), .ZN(n15762) );
  AND2_X1 U15791 ( .A1(n15763), .A2(n15632), .ZN(n15761) );
  OR2_X1 U15792 ( .A1(n15764), .A2(n15765), .ZN(n15632) );
  AND2_X1 U15793 ( .A1(n15628), .A2(n15629), .ZN(n15765) );
  AND2_X1 U15794 ( .A1(n15627), .A2(n15766), .ZN(n15764) );
  OR2_X1 U15795 ( .A1(n15629), .A2(n15628), .ZN(n15766) );
  OR2_X1 U15796 ( .A1(n9006), .A2(n8911), .ZN(n15628) );
  OR2_X1 U15797 ( .A1(n15767), .A2(n15768), .ZN(n15629) );
  AND2_X1 U15798 ( .A1(n15622), .A2(n15625), .ZN(n15768) );
  AND2_X1 U15799 ( .A1(n15769), .A2(n15624), .ZN(n15767) );
  OR2_X1 U15800 ( .A1(n15770), .A2(n15771), .ZN(n15624) );
  AND2_X1 U15801 ( .A1(n15619), .A2(n15620), .ZN(n15771) );
  AND2_X1 U15802 ( .A1(n15772), .A2(n15773), .ZN(n15770) );
  OR2_X1 U15803 ( .A1(n15620), .A2(n15619), .ZN(n15773) );
  OR2_X1 U15804 ( .A1(n9014), .A2(n8911), .ZN(n15619) );
  OR2_X1 U15805 ( .A1(n9984), .A2(n15774), .ZN(n15620) );
  OR2_X1 U15806 ( .A1(n8911), .A2(n8907), .ZN(n15774) );
  INV_X1 U15807 ( .A(n15621), .ZN(n15772) );
  OR2_X1 U15808 ( .A1(n15775), .A2(n15776), .ZN(n15621) );
  AND2_X1 U15809 ( .A1(b_2_), .A2(n15777), .ZN(n15776) );
  OR2_X1 U15810 ( .A1(n15778), .A2(n9989), .ZN(n15777) );
  AND2_X1 U15811 ( .A1(a_30_), .A2(n8903), .ZN(n15778) );
  AND2_X1 U15812 ( .A1(b_1_), .A2(n15779), .ZN(n15775) );
  OR2_X1 U15813 ( .A1(n15780), .A2(n8021), .ZN(n15779) );
  AND2_X1 U15814 ( .A1(a_31_), .A2(n8907), .ZN(n15780) );
  OR2_X1 U15815 ( .A1(n15625), .A2(n15622), .ZN(n15769) );
  XOR2_X1 U15816 ( .A(n15781), .B(n15782), .Z(n15622) );
  XNOR2_X1 U15817 ( .A(n15783), .B(n15784), .ZN(n15781) );
  OR2_X1 U15818 ( .A1(n9010), .A2(n8911), .ZN(n15625) );
  XOR2_X1 U15819 ( .A(n15785), .B(n15786), .Z(n15627) );
  XOR2_X1 U15820 ( .A(n15787), .B(n15788), .Z(n15786) );
  OR2_X1 U15821 ( .A1(n15633), .A2(n15630), .ZN(n15763) );
  XOR2_X1 U15822 ( .A(n15789), .B(n15790), .Z(n15630) );
  XOR2_X1 U15823 ( .A(n15791), .B(n15792), .Z(n15790) );
  OR2_X1 U15824 ( .A1(n9002), .A2(n8911), .ZN(n15633) );
  XOR2_X1 U15825 ( .A(n15793), .B(n15794), .Z(n15634) );
  XOR2_X1 U15826 ( .A(n15795), .B(n15796), .Z(n15794) );
  XOR2_X1 U15827 ( .A(n15797), .B(n15798), .Z(n15638) );
  XOR2_X1 U15828 ( .A(n15799), .B(n15800), .Z(n15798) );
  XOR2_X1 U15829 ( .A(n15801), .B(n15802), .Z(n15642) );
  XOR2_X1 U15830 ( .A(n15803), .B(n15804), .Z(n15802) );
  XOR2_X1 U15831 ( .A(n15805), .B(n15806), .Z(n15646) );
  XOR2_X1 U15832 ( .A(n15807), .B(n15808), .Z(n15806) );
  XOR2_X1 U15833 ( .A(n15809), .B(n15810), .Z(n15650) );
  XOR2_X1 U15834 ( .A(n15811), .B(n15812), .Z(n15810) );
  XOR2_X1 U15835 ( .A(n15813), .B(n15814), .Z(n15654) );
  XOR2_X1 U15836 ( .A(n15815), .B(n15816), .Z(n15814) );
  XOR2_X1 U15837 ( .A(n15817), .B(n15818), .Z(n15658) );
  XOR2_X1 U15838 ( .A(n15819), .B(n15820), .Z(n15818) );
  XOR2_X1 U15839 ( .A(n15821), .B(n15822), .Z(n15662) );
  XOR2_X1 U15840 ( .A(n15823), .B(n15824), .Z(n15822) );
  XOR2_X1 U15841 ( .A(n15825), .B(n15826), .Z(n15666) );
  XOR2_X1 U15842 ( .A(n15827), .B(n15828), .Z(n15826) );
  XOR2_X1 U15843 ( .A(n15829), .B(n15830), .Z(n15670) );
  XOR2_X1 U15844 ( .A(n15831), .B(n15832), .Z(n15830) );
  XOR2_X1 U15845 ( .A(n15833), .B(n15834), .Z(n15674) );
  XOR2_X1 U15846 ( .A(n15835), .B(n15836), .Z(n15834) );
  XOR2_X1 U15847 ( .A(n15837), .B(n15838), .Z(n15678) );
  XOR2_X1 U15848 ( .A(n15839), .B(n15840), .Z(n15838) );
  XOR2_X1 U15849 ( .A(n15841), .B(n15842), .Z(n15682) );
  XOR2_X1 U15850 ( .A(n15843), .B(n15844), .Z(n15842) );
  XOR2_X1 U15851 ( .A(n15845), .B(n15846), .Z(n15686) );
  XOR2_X1 U15852 ( .A(n15847), .B(n15848), .Z(n15846) );
  XOR2_X1 U15853 ( .A(n15849), .B(n15850), .Z(n15690) );
  XOR2_X1 U15854 ( .A(n15851), .B(n15852), .Z(n15850) );
  XOR2_X1 U15855 ( .A(n15853), .B(n15854), .Z(n15694) );
  XOR2_X1 U15856 ( .A(n15855), .B(n15856), .Z(n15854) );
  XOR2_X1 U15857 ( .A(n15857), .B(n15858), .Z(n15698) );
  XOR2_X1 U15858 ( .A(n15859), .B(n15860), .Z(n15858) );
  XOR2_X1 U15859 ( .A(n15861), .B(n15862), .Z(n15702) );
  XOR2_X1 U15860 ( .A(n15863), .B(n15864), .Z(n15862) );
  XOR2_X1 U15861 ( .A(n15865), .B(n15866), .Z(n9705) );
  XOR2_X1 U15862 ( .A(n15867), .B(n15868), .Z(n15866) );
  AND2_X1 U15863 ( .A1(n9121), .A2(n15869), .ZN(n9123) );
  AND2_X1 U15864 ( .A1(n9122), .A2(n9120), .ZN(n15869) );
  XOR2_X1 U15865 ( .A(n15870), .B(n15871), .Z(n9120) );
  OR2_X1 U15866 ( .A1(n9389), .A2(n9297), .ZN(n15870) );
  XNOR2_X1 U15867 ( .A(n15872), .B(n15873), .ZN(n9122) );
  XOR2_X1 U15868 ( .A(n15874), .B(n15875), .Z(n15873) );
  INV_X1 U15869 ( .A(n9394), .ZN(n9121) );
  OR2_X1 U15870 ( .A1(n15876), .A2(n15877), .ZN(n9394) );
  AND2_X1 U15871 ( .A1(n9415), .A2(n9414), .ZN(n15877) );
  AND2_X1 U15872 ( .A1(n9412), .A2(n15878), .ZN(n15876) );
  OR2_X1 U15873 ( .A1(n9414), .A2(n9415), .ZN(n15878) );
  OR2_X1 U15874 ( .A1(n9297), .A2(n8907), .ZN(n9415) );
  OR2_X1 U15875 ( .A1(n15879), .A2(n15880), .ZN(n9414) );
  AND2_X1 U15876 ( .A1(n9432), .A2(n9431), .ZN(n15880) );
  AND2_X1 U15877 ( .A1(n9429), .A2(n15881), .ZN(n15879) );
  OR2_X1 U15878 ( .A1(n9431), .A2(n9432), .ZN(n15881) );
  OR2_X1 U15879 ( .A1(n8902), .A2(n8907), .ZN(n9432) );
  OR2_X1 U15880 ( .A1(n15882), .A2(n15883), .ZN(n9431) );
  AND2_X1 U15881 ( .A1(n8837), .A2(n9466), .ZN(n15883) );
  AND2_X1 U15882 ( .A1(n9464), .A2(n15884), .ZN(n15882) );
  OR2_X1 U15883 ( .A1(n9466), .A2(n8837), .ZN(n15884) );
  OR2_X1 U15884 ( .A1(n8906), .A2(n8907), .ZN(n8837) );
  OR2_X1 U15885 ( .A1(n15885), .A2(n15886), .ZN(n9466) );
  AND2_X1 U15886 ( .A1(n9496), .A2(n9495), .ZN(n15886) );
  AND2_X1 U15887 ( .A1(n9493), .A2(n15887), .ZN(n15885) );
  OR2_X1 U15888 ( .A1(n9495), .A2(n9496), .ZN(n15887) );
  OR2_X1 U15889 ( .A1(n8910), .A2(n8907), .ZN(n9496) );
  OR2_X1 U15890 ( .A1(n15888), .A2(n15889), .ZN(n9495) );
  AND2_X1 U15891 ( .A1(n9545), .A2(n9544), .ZN(n15889) );
  AND2_X1 U15892 ( .A1(n9542), .A2(n15890), .ZN(n15888) );
  OR2_X1 U15893 ( .A1(n9544), .A2(n9545), .ZN(n15890) );
  OR2_X1 U15894 ( .A1(n8914), .A2(n8907), .ZN(n9545) );
  OR2_X1 U15895 ( .A1(n15891), .A2(n15892), .ZN(n9544) );
  AND2_X1 U15896 ( .A1(n9589), .A2(n9588), .ZN(n15892) );
  AND2_X1 U15897 ( .A1(n9586), .A2(n15893), .ZN(n15891) );
  OR2_X1 U15898 ( .A1(n9588), .A2(n9589), .ZN(n15893) );
  OR2_X1 U15899 ( .A1(n8918), .A2(n8907), .ZN(n9589) );
  OR2_X1 U15900 ( .A1(n15894), .A2(n15895), .ZN(n9588) );
  AND2_X1 U15901 ( .A1(n9652), .A2(n9651), .ZN(n15895) );
  AND2_X1 U15902 ( .A1(n9649), .A2(n15896), .ZN(n15894) );
  OR2_X1 U15903 ( .A1(n9651), .A2(n9652), .ZN(n15896) );
  OR2_X1 U15904 ( .A1(n8922), .A2(n8907), .ZN(n9652) );
  OR2_X1 U15905 ( .A1(n15897), .A2(n15898), .ZN(n9651) );
  AND2_X1 U15906 ( .A1(n9710), .A2(n9709), .ZN(n15898) );
  AND2_X1 U15907 ( .A1(n9707), .A2(n15899), .ZN(n15897) );
  OR2_X1 U15908 ( .A1(n9709), .A2(n9710), .ZN(n15899) );
  OR2_X1 U15909 ( .A1(n8926), .A2(n8907), .ZN(n9710) );
  OR2_X1 U15910 ( .A1(n15900), .A2(n15901), .ZN(n9709) );
  AND2_X1 U15911 ( .A1(n15868), .A2(n15867), .ZN(n15901) );
  AND2_X1 U15912 ( .A1(n15865), .A2(n15902), .ZN(n15900) );
  OR2_X1 U15913 ( .A1(n15867), .A2(n15868), .ZN(n15902) );
  OR2_X1 U15914 ( .A1(n8930), .A2(n8907), .ZN(n15868) );
  OR2_X1 U15915 ( .A1(n15903), .A2(n15904), .ZN(n15867) );
  AND2_X1 U15916 ( .A1(n15864), .A2(n15863), .ZN(n15904) );
  AND2_X1 U15917 ( .A1(n15861), .A2(n15905), .ZN(n15903) );
  OR2_X1 U15918 ( .A1(n15863), .A2(n15864), .ZN(n15905) );
  OR2_X1 U15919 ( .A1(n8934), .A2(n8907), .ZN(n15864) );
  OR2_X1 U15920 ( .A1(n15906), .A2(n15907), .ZN(n15863) );
  AND2_X1 U15921 ( .A1(n15860), .A2(n15859), .ZN(n15907) );
  AND2_X1 U15922 ( .A1(n15857), .A2(n15908), .ZN(n15906) );
  OR2_X1 U15923 ( .A1(n15859), .A2(n15860), .ZN(n15908) );
  OR2_X1 U15924 ( .A1(n8938), .A2(n8907), .ZN(n15860) );
  OR2_X1 U15925 ( .A1(n15909), .A2(n15910), .ZN(n15859) );
  AND2_X1 U15926 ( .A1(n15856), .A2(n15855), .ZN(n15910) );
  AND2_X1 U15927 ( .A1(n15853), .A2(n15911), .ZN(n15909) );
  OR2_X1 U15928 ( .A1(n15855), .A2(n15856), .ZN(n15911) );
  OR2_X1 U15929 ( .A1(n8942), .A2(n8907), .ZN(n15856) );
  OR2_X1 U15930 ( .A1(n15912), .A2(n15913), .ZN(n15855) );
  AND2_X1 U15931 ( .A1(n15852), .A2(n15851), .ZN(n15913) );
  AND2_X1 U15932 ( .A1(n15849), .A2(n15914), .ZN(n15912) );
  OR2_X1 U15933 ( .A1(n15851), .A2(n15852), .ZN(n15914) );
  OR2_X1 U15934 ( .A1(n8946), .A2(n8907), .ZN(n15852) );
  OR2_X1 U15935 ( .A1(n15915), .A2(n15916), .ZN(n15851) );
  AND2_X1 U15936 ( .A1(n15848), .A2(n15847), .ZN(n15916) );
  AND2_X1 U15937 ( .A1(n15845), .A2(n15917), .ZN(n15915) );
  OR2_X1 U15938 ( .A1(n15847), .A2(n15848), .ZN(n15917) );
  OR2_X1 U15939 ( .A1(n8950), .A2(n8907), .ZN(n15848) );
  OR2_X1 U15940 ( .A1(n15918), .A2(n15919), .ZN(n15847) );
  AND2_X1 U15941 ( .A1(n15844), .A2(n15843), .ZN(n15919) );
  AND2_X1 U15942 ( .A1(n15841), .A2(n15920), .ZN(n15918) );
  OR2_X1 U15943 ( .A1(n15843), .A2(n15844), .ZN(n15920) );
  OR2_X1 U15944 ( .A1(n8954), .A2(n8907), .ZN(n15844) );
  OR2_X1 U15945 ( .A1(n15921), .A2(n15922), .ZN(n15843) );
  AND2_X1 U15946 ( .A1(n15840), .A2(n15839), .ZN(n15922) );
  AND2_X1 U15947 ( .A1(n15837), .A2(n15923), .ZN(n15921) );
  OR2_X1 U15948 ( .A1(n15839), .A2(n15840), .ZN(n15923) );
  OR2_X1 U15949 ( .A1(n8958), .A2(n8907), .ZN(n15840) );
  OR2_X1 U15950 ( .A1(n15924), .A2(n15925), .ZN(n15839) );
  AND2_X1 U15951 ( .A1(n15836), .A2(n15835), .ZN(n15925) );
  AND2_X1 U15952 ( .A1(n15833), .A2(n15926), .ZN(n15924) );
  OR2_X1 U15953 ( .A1(n15835), .A2(n15836), .ZN(n15926) );
  OR2_X1 U15954 ( .A1(n8962), .A2(n8907), .ZN(n15836) );
  OR2_X1 U15955 ( .A1(n15927), .A2(n15928), .ZN(n15835) );
  AND2_X1 U15956 ( .A1(n15832), .A2(n15831), .ZN(n15928) );
  AND2_X1 U15957 ( .A1(n15829), .A2(n15929), .ZN(n15927) );
  OR2_X1 U15958 ( .A1(n15831), .A2(n15832), .ZN(n15929) );
  OR2_X1 U15959 ( .A1(n8966), .A2(n8907), .ZN(n15832) );
  OR2_X1 U15960 ( .A1(n15930), .A2(n15931), .ZN(n15831) );
  AND2_X1 U15961 ( .A1(n15828), .A2(n15827), .ZN(n15931) );
  AND2_X1 U15962 ( .A1(n15825), .A2(n15932), .ZN(n15930) );
  OR2_X1 U15963 ( .A1(n15827), .A2(n15828), .ZN(n15932) );
  OR2_X1 U15964 ( .A1(n8970), .A2(n8907), .ZN(n15828) );
  OR2_X1 U15965 ( .A1(n15933), .A2(n15934), .ZN(n15827) );
  AND2_X1 U15966 ( .A1(n15824), .A2(n15823), .ZN(n15934) );
  AND2_X1 U15967 ( .A1(n15821), .A2(n15935), .ZN(n15933) );
  OR2_X1 U15968 ( .A1(n15823), .A2(n15824), .ZN(n15935) );
  OR2_X1 U15969 ( .A1(n8974), .A2(n8907), .ZN(n15824) );
  OR2_X1 U15970 ( .A1(n15936), .A2(n15937), .ZN(n15823) );
  AND2_X1 U15971 ( .A1(n15820), .A2(n15819), .ZN(n15937) );
  AND2_X1 U15972 ( .A1(n15817), .A2(n15938), .ZN(n15936) );
  OR2_X1 U15973 ( .A1(n15819), .A2(n15820), .ZN(n15938) );
  OR2_X1 U15974 ( .A1(n8978), .A2(n8907), .ZN(n15820) );
  OR2_X1 U15975 ( .A1(n15939), .A2(n15940), .ZN(n15819) );
  AND2_X1 U15976 ( .A1(n15816), .A2(n15815), .ZN(n15940) );
  AND2_X1 U15977 ( .A1(n15813), .A2(n15941), .ZN(n15939) );
  OR2_X1 U15978 ( .A1(n15815), .A2(n15816), .ZN(n15941) );
  OR2_X1 U15979 ( .A1(n8982), .A2(n8907), .ZN(n15816) );
  OR2_X1 U15980 ( .A1(n15942), .A2(n15943), .ZN(n15815) );
  AND2_X1 U15981 ( .A1(n15812), .A2(n15811), .ZN(n15943) );
  AND2_X1 U15982 ( .A1(n15809), .A2(n15944), .ZN(n15942) );
  OR2_X1 U15983 ( .A1(n15811), .A2(n15812), .ZN(n15944) );
  OR2_X1 U15984 ( .A1(n8986), .A2(n8907), .ZN(n15812) );
  OR2_X1 U15985 ( .A1(n15945), .A2(n15946), .ZN(n15811) );
  AND2_X1 U15986 ( .A1(n15808), .A2(n15807), .ZN(n15946) );
  AND2_X1 U15987 ( .A1(n15805), .A2(n15947), .ZN(n15945) );
  OR2_X1 U15988 ( .A1(n15807), .A2(n15808), .ZN(n15947) );
  OR2_X1 U15989 ( .A1(n8990), .A2(n8907), .ZN(n15808) );
  OR2_X1 U15990 ( .A1(n15948), .A2(n15949), .ZN(n15807) );
  AND2_X1 U15991 ( .A1(n15804), .A2(n15803), .ZN(n15949) );
  AND2_X1 U15992 ( .A1(n15801), .A2(n15950), .ZN(n15948) );
  OR2_X1 U15993 ( .A1(n15803), .A2(n15804), .ZN(n15950) );
  OR2_X1 U15994 ( .A1(n8994), .A2(n8907), .ZN(n15804) );
  OR2_X1 U15995 ( .A1(n15951), .A2(n15952), .ZN(n15803) );
  AND2_X1 U15996 ( .A1(n15800), .A2(n15799), .ZN(n15952) );
  AND2_X1 U15997 ( .A1(n15797), .A2(n15953), .ZN(n15951) );
  OR2_X1 U15998 ( .A1(n15799), .A2(n15800), .ZN(n15953) );
  OR2_X1 U15999 ( .A1(n8998), .A2(n8907), .ZN(n15800) );
  OR2_X1 U16000 ( .A1(n15954), .A2(n15955), .ZN(n15799) );
  AND2_X1 U16001 ( .A1(n15796), .A2(n15795), .ZN(n15955) );
  AND2_X1 U16002 ( .A1(n15793), .A2(n15956), .ZN(n15954) );
  OR2_X1 U16003 ( .A1(n15795), .A2(n15796), .ZN(n15956) );
  OR2_X1 U16004 ( .A1(n9002), .A2(n8907), .ZN(n15796) );
  OR2_X1 U16005 ( .A1(n15957), .A2(n15958), .ZN(n15795) );
  AND2_X1 U16006 ( .A1(n15789), .A2(n15792), .ZN(n15958) );
  AND2_X1 U16007 ( .A1(n15959), .A2(n15791), .ZN(n15957) );
  OR2_X1 U16008 ( .A1(n15960), .A2(n15961), .ZN(n15791) );
  AND2_X1 U16009 ( .A1(n15788), .A2(n15787), .ZN(n15961) );
  AND2_X1 U16010 ( .A1(n15785), .A2(n15962), .ZN(n15960) );
  OR2_X1 U16011 ( .A1(n15787), .A2(n15788), .ZN(n15962) );
  OR2_X1 U16012 ( .A1(n9010), .A2(n8907), .ZN(n15788) );
  OR2_X1 U16013 ( .A1(n15963), .A2(n15964), .ZN(n15787) );
  AND2_X1 U16014 ( .A1(n15782), .A2(n15783), .ZN(n15964) );
  AND2_X1 U16015 ( .A1(n15965), .A2(n15966), .ZN(n15963) );
  OR2_X1 U16016 ( .A1(n15783), .A2(n15782), .ZN(n15966) );
  OR2_X1 U16017 ( .A1(n9014), .A2(n8907), .ZN(n15782) );
  OR2_X1 U16018 ( .A1(n9984), .A2(n15967), .ZN(n15783) );
  OR2_X1 U16019 ( .A1(n8907), .A2(n8903), .ZN(n15967) );
  INV_X1 U16020 ( .A(n15784), .ZN(n15965) );
  OR2_X1 U16021 ( .A1(n15968), .A2(n15969), .ZN(n15784) );
  AND2_X1 U16022 ( .A1(b_1_), .A2(n15970), .ZN(n15969) );
  OR2_X1 U16023 ( .A1(n15971), .A2(n9989), .ZN(n15970) );
  AND2_X1 U16024 ( .A1(n9294), .A2(a_30_), .ZN(n9989) );
  AND2_X1 U16025 ( .A1(a_30_), .A2(n9389), .ZN(n15971) );
  AND2_X1 U16026 ( .A1(b_0_), .A2(n15972), .ZN(n15968) );
  OR2_X1 U16027 ( .A1(n15973), .A2(n8021), .ZN(n15972) );
  AND2_X1 U16028 ( .A1(n8002), .A2(a_31_), .ZN(n8021) );
  AND2_X1 U16029 ( .A1(a_31_), .A2(n8903), .ZN(n15973) );
  XOR2_X1 U16030 ( .A(n15974), .B(n15975), .Z(n15785) );
  XOR2_X1 U16031 ( .A(n15976), .B(n15977), .Z(n15974) );
  OR2_X1 U16032 ( .A1(n15792), .A2(n15789), .ZN(n15959) );
  XNOR2_X1 U16033 ( .A(n15978), .B(n15979), .ZN(n15789) );
  XNOR2_X1 U16034 ( .A(n15980), .B(n15981), .ZN(n15979) );
  OR2_X1 U16035 ( .A1(n9006), .A2(n8907), .ZN(n15792) );
  XNOR2_X1 U16036 ( .A(n15982), .B(n15983), .ZN(n15793) );
  XNOR2_X1 U16037 ( .A(n15984), .B(n15985), .ZN(n15982) );
  XNOR2_X1 U16038 ( .A(n15986), .B(n15987), .ZN(n15797) );
  XNOR2_X1 U16039 ( .A(n15988), .B(n15989), .ZN(n15986) );
  XNOR2_X1 U16040 ( .A(n15990), .B(n15991), .ZN(n15801) );
  XNOR2_X1 U16041 ( .A(n15992), .B(n15993), .ZN(n15990) );
  XNOR2_X1 U16042 ( .A(n15994), .B(n15995), .ZN(n15805) );
  XNOR2_X1 U16043 ( .A(n15996), .B(n15997), .ZN(n15994) );
  XNOR2_X1 U16044 ( .A(n15998), .B(n15999), .ZN(n15809) );
  XNOR2_X1 U16045 ( .A(n16000), .B(n16001), .ZN(n15998) );
  XNOR2_X1 U16046 ( .A(n16002), .B(n16003), .ZN(n15813) );
  XNOR2_X1 U16047 ( .A(n16004), .B(n16005), .ZN(n16002) );
  XNOR2_X1 U16048 ( .A(n16006), .B(n16007), .ZN(n15817) );
  XNOR2_X1 U16049 ( .A(n16008), .B(n16009), .ZN(n16006) );
  XNOR2_X1 U16050 ( .A(n16010), .B(n16011), .ZN(n15821) );
  XNOR2_X1 U16051 ( .A(n16012), .B(n16013), .ZN(n16010) );
  XNOR2_X1 U16052 ( .A(n16014), .B(n16015), .ZN(n15825) );
  XNOR2_X1 U16053 ( .A(n16016), .B(n16017), .ZN(n16014) );
  XNOR2_X1 U16054 ( .A(n16018), .B(n16019), .ZN(n15829) );
  XNOR2_X1 U16055 ( .A(n16020), .B(n16021), .ZN(n16018) );
  XNOR2_X1 U16056 ( .A(n16022), .B(n16023), .ZN(n15833) );
  XNOR2_X1 U16057 ( .A(n16024), .B(n16025), .ZN(n16022) );
  XNOR2_X1 U16058 ( .A(n16026), .B(n16027), .ZN(n15837) );
  XNOR2_X1 U16059 ( .A(n16028), .B(n16029), .ZN(n16026) );
  XNOR2_X1 U16060 ( .A(n16030), .B(n16031), .ZN(n15841) );
  XNOR2_X1 U16061 ( .A(n16032), .B(n16033), .ZN(n16030) );
  XNOR2_X1 U16062 ( .A(n16034), .B(n16035), .ZN(n15845) );
  XNOR2_X1 U16063 ( .A(n16036), .B(n16037), .ZN(n16034) );
  XNOR2_X1 U16064 ( .A(n16038), .B(n16039), .ZN(n15849) );
  XNOR2_X1 U16065 ( .A(n16040), .B(n16041), .ZN(n16038) );
  XNOR2_X1 U16066 ( .A(n16042), .B(n16043), .ZN(n15853) );
  XNOR2_X1 U16067 ( .A(n16044), .B(n16045), .ZN(n16042) );
  XNOR2_X1 U16068 ( .A(n16046), .B(n16047), .ZN(n15857) );
  XNOR2_X1 U16069 ( .A(n16048), .B(n16049), .ZN(n16046) );
  XNOR2_X1 U16070 ( .A(n16050), .B(n16051), .ZN(n15861) );
  XNOR2_X1 U16071 ( .A(n16052), .B(n16053), .ZN(n16050) );
  XNOR2_X1 U16072 ( .A(n16054), .B(n16055), .ZN(n15865) );
  XNOR2_X1 U16073 ( .A(n16056), .B(n16057), .ZN(n16054) );
  XOR2_X1 U16074 ( .A(n16058), .B(n16059), .Z(n9707) );
  XOR2_X1 U16075 ( .A(n16060), .B(n16061), .Z(n16059) );
  XOR2_X1 U16076 ( .A(n16062), .B(n16063), .Z(n9649) );
  XOR2_X1 U16077 ( .A(n16064), .B(n16065), .Z(n16063) );
  XOR2_X1 U16078 ( .A(n16066), .B(n16067), .Z(n9586) );
  XOR2_X1 U16079 ( .A(n16068), .B(n16069), .Z(n16067) );
  XOR2_X1 U16080 ( .A(n16070), .B(n16071), .Z(n9542) );
  XOR2_X1 U16081 ( .A(n16072), .B(n16073), .Z(n16071) );
  XOR2_X1 U16082 ( .A(n16074), .B(n16075), .Z(n9493) );
  XOR2_X1 U16083 ( .A(n16076), .B(n16077), .Z(n16075) );
  XOR2_X1 U16084 ( .A(n16078), .B(n16079), .Z(n9464) );
  XOR2_X1 U16085 ( .A(n16080), .B(n16081), .Z(n16079) );
  XOR2_X1 U16086 ( .A(n16082), .B(n16083), .Z(n9429) );
  XOR2_X1 U16087 ( .A(n16084), .B(n16085), .Z(n16083) );
  XOR2_X1 U16088 ( .A(n16086), .B(n16087), .Z(n9412) );
  XOR2_X1 U16089 ( .A(n16088), .B(n8866), .Z(n16087) );
  INV_X1 U16090 ( .A(n16089), .ZN(n9391) );
  OR2_X1 U16091 ( .A1(n15871), .A2(n9297), .ZN(n16089) );
  OR2_X1 U16092 ( .A1(n16090), .A2(n16091), .ZN(n15871) );
  AND2_X1 U16093 ( .A1(n15872), .A2(n15874), .ZN(n16091) );
  AND2_X1 U16094 ( .A1(n16092), .A2(n15875), .ZN(n16090) );
  OR2_X1 U16095 ( .A1(n9297), .A2(n8903), .ZN(n15875) );
  INV_X1 U16096 ( .A(a_0_), .ZN(n9297) );
  OR2_X1 U16097 ( .A1(n15874), .A2(n15872), .ZN(n16092) );
  OR2_X1 U16098 ( .A1(n9389), .A2(n8902), .ZN(n15872) );
  OR2_X1 U16099 ( .A1(n16093), .A2(n16094), .ZN(n15874) );
  AND2_X1 U16100 ( .A1(n16086), .A2(n16088), .ZN(n16094) );
  AND2_X1 U16101 ( .A1(n16095), .A2(n8866), .ZN(n16093) );
  OR2_X1 U16102 ( .A1(n8902), .A2(n8903), .ZN(n8866) );
  INV_X1 U16103 ( .A(a_1_), .ZN(n8902) );
  OR2_X1 U16104 ( .A1(n16088), .A2(n16086), .ZN(n16095) );
  OR2_X1 U16105 ( .A1(n9389), .A2(n8906), .ZN(n16086) );
  OR2_X1 U16106 ( .A1(n16096), .A2(n16097), .ZN(n16088) );
  AND2_X1 U16107 ( .A1(n16082), .A2(n16084), .ZN(n16097) );
  AND2_X1 U16108 ( .A1(n16098), .A2(n16085), .ZN(n16096) );
  OR2_X1 U16109 ( .A1(n9389), .A2(n8910), .ZN(n16085) );
  OR2_X1 U16110 ( .A1(n16084), .A2(n16082), .ZN(n16098) );
  OR2_X1 U16111 ( .A1(n8906), .A2(n8903), .ZN(n16082) );
  INV_X1 U16112 ( .A(a_2_), .ZN(n8906) );
  OR2_X1 U16113 ( .A1(n16099), .A2(n16100), .ZN(n16084) );
  AND2_X1 U16114 ( .A1(n16078), .A2(n16080), .ZN(n16100) );
  AND2_X1 U16115 ( .A1(n16101), .A2(n16081), .ZN(n16099) );
  OR2_X1 U16116 ( .A1(n9389), .A2(n8914), .ZN(n16081) );
  OR2_X1 U16117 ( .A1(n16080), .A2(n16078), .ZN(n16101) );
  OR2_X1 U16118 ( .A1(n8910), .A2(n8903), .ZN(n16078) );
  INV_X1 U16119 ( .A(a_3_), .ZN(n8910) );
  OR2_X1 U16120 ( .A1(n16102), .A2(n16103), .ZN(n16080) );
  AND2_X1 U16121 ( .A1(n16074), .A2(n16076), .ZN(n16103) );
  AND2_X1 U16122 ( .A1(n16104), .A2(n16077), .ZN(n16102) );
  OR2_X1 U16123 ( .A1(n9389), .A2(n8918), .ZN(n16077) );
  OR2_X1 U16124 ( .A1(n16076), .A2(n16074), .ZN(n16104) );
  OR2_X1 U16125 ( .A1(n8914), .A2(n8903), .ZN(n16074) );
  INV_X1 U16126 ( .A(a_4_), .ZN(n8914) );
  OR2_X1 U16127 ( .A1(n16105), .A2(n16106), .ZN(n16076) );
  AND2_X1 U16128 ( .A1(n16070), .A2(n16072), .ZN(n16106) );
  AND2_X1 U16129 ( .A1(n16107), .A2(n16073), .ZN(n16105) );
  OR2_X1 U16130 ( .A1(n9389), .A2(n8922), .ZN(n16073) );
  OR2_X1 U16131 ( .A1(n16072), .A2(n16070), .ZN(n16107) );
  OR2_X1 U16132 ( .A1(n8918), .A2(n8903), .ZN(n16070) );
  INV_X1 U16133 ( .A(a_5_), .ZN(n8918) );
  OR2_X1 U16134 ( .A1(n16108), .A2(n16109), .ZN(n16072) );
  AND2_X1 U16135 ( .A1(n16066), .A2(n16068), .ZN(n16109) );
  AND2_X1 U16136 ( .A1(n16110), .A2(n16069), .ZN(n16108) );
  OR2_X1 U16137 ( .A1(n9389), .A2(n8926), .ZN(n16069) );
  OR2_X1 U16138 ( .A1(n16068), .A2(n16066), .ZN(n16110) );
  OR2_X1 U16139 ( .A1(n8922), .A2(n8903), .ZN(n16066) );
  INV_X1 U16140 ( .A(a_6_), .ZN(n8922) );
  OR2_X1 U16141 ( .A1(n16111), .A2(n16112), .ZN(n16068) );
  AND2_X1 U16142 ( .A1(n16062), .A2(n16064), .ZN(n16112) );
  AND2_X1 U16143 ( .A1(n16113), .A2(n16065), .ZN(n16111) );
  OR2_X1 U16144 ( .A1(n9389), .A2(n8930), .ZN(n16065) );
  OR2_X1 U16145 ( .A1(n16064), .A2(n16062), .ZN(n16113) );
  OR2_X1 U16146 ( .A1(n8926), .A2(n8903), .ZN(n16062) );
  INV_X1 U16147 ( .A(a_7_), .ZN(n8926) );
  OR2_X1 U16148 ( .A1(n16114), .A2(n16115), .ZN(n16064) );
  AND2_X1 U16149 ( .A1(n16058), .A2(n16060), .ZN(n16115) );
  AND2_X1 U16150 ( .A1(n16116), .A2(n16061), .ZN(n16114) );
  OR2_X1 U16151 ( .A1(n9389), .A2(n8934), .ZN(n16061) );
  OR2_X1 U16152 ( .A1(n16060), .A2(n16058), .ZN(n16116) );
  OR2_X1 U16153 ( .A1(n8930), .A2(n8903), .ZN(n16058) );
  INV_X1 U16154 ( .A(a_8_), .ZN(n8930) );
  OR2_X1 U16155 ( .A1(n16117), .A2(n16118), .ZN(n16060) );
  AND2_X1 U16156 ( .A1(n16055), .A2(n16057), .ZN(n16118) );
  AND2_X1 U16157 ( .A1(n16119), .A2(n16056), .ZN(n16117) );
  OR2_X1 U16158 ( .A1(n9389), .A2(n8938), .ZN(n16056) );
  OR2_X1 U16159 ( .A1(n16057), .A2(n16055), .ZN(n16119) );
  OR2_X1 U16160 ( .A1(n8934), .A2(n8903), .ZN(n16055) );
  INV_X1 U16161 ( .A(a_9_), .ZN(n8934) );
  OR2_X1 U16162 ( .A1(n16120), .A2(n16121), .ZN(n16057) );
  AND2_X1 U16163 ( .A1(n16051), .A2(n16053), .ZN(n16121) );
  AND2_X1 U16164 ( .A1(n16122), .A2(n16052), .ZN(n16120) );
  OR2_X1 U16165 ( .A1(n9389), .A2(n8942), .ZN(n16052) );
  OR2_X1 U16166 ( .A1(n16053), .A2(n16051), .ZN(n16122) );
  OR2_X1 U16167 ( .A1(n8938), .A2(n8903), .ZN(n16051) );
  INV_X1 U16168 ( .A(a_10_), .ZN(n8938) );
  OR2_X1 U16169 ( .A1(n16123), .A2(n16124), .ZN(n16053) );
  AND2_X1 U16170 ( .A1(n16047), .A2(n16049), .ZN(n16124) );
  AND2_X1 U16171 ( .A1(n16125), .A2(n16048), .ZN(n16123) );
  OR2_X1 U16172 ( .A1(n9389), .A2(n8946), .ZN(n16048) );
  OR2_X1 U16173 ( .A1(n16049), .A2(n16047), .ZN(n16125) );
  OR2_X1 U16174 ( .A1(n8942), .A2(n8903), .ZN(n16047) );
  INV_X1 U16175 ( .A(a_11_), .ZN(n8942) );
  OR2_X1 U16176 ( .A1(n16126), .A2(n16127), .ZN(n16049) );
  AND2_X1 U16177 ( .A1(n16043), .A2(n16045), .ZN(n16127) );
  AND2_X1 U16178 ( .A1(n16128), .A2(n16044), .ZN(n16126) );
  OR2_X1 U16179 ( .A1(n9389), .A2(n8950), .ZN(n16044) );
  OR2_X1 U16180 ( .A1(n16045), .A2(n16043), .ZN(n16128) );
  OR2_X1 U16181 ( .A1(n8946), .A2(n8903), .ZN(n16043) );
  INV_X1 U16182 ( .A(a_12_), .ZN(n8946) );
  OR2_X1 U16183 ( .A1(n16129), .A2(n16130), .ZN(n16045) );
  AND2_X1 U16184 ( .A1(n16039), .A2(n16041), .ZN(n16130) );
  AND2_X1 U16185 ( .A1(n16131), .A2(n16040), .ZN(n16129) );
  OR2_X1 U16186 ( .A1(n9389), .A2(n8954), .ZN(n16040) );
  OR2_X1 U16187 ( .A1(n16041), .A2(n16039), .ZN(n16131) );
  OR2_X1 U16188 ( .A1(n8950), .A2(n8903), .ZN(n16039) );
  INV_X1 U16189 ( .A(a_13_), .ZN(n8950) );
  OR2_X1 U16190 ( .A1(n16132), .A2(n16133), .ZN(n16041) );
  AND2_X1 U16191 ( .A1(n16035), .A2(n16037), .ZN(n16133) );
  AND2_X1 U16192 ( .A1(n16134), .A2(n16036), .ZN(n16132) );
  OR2_X1 U16193 ( .A1(n9389), .A2(n8958), .ZN(n16036) );
  OR2_X1 U16194 ( .A1(n16037), .A2(n16035), .ZN(n16134) );
  OR2_X1 U16195 ( .A1(n8954), .A2(n8903), .ZN(n16035) );
  INV_X1 U16196 ( .A(a_14_), .ZN(n8954) );
  OR2_X1 U16197 ( .A1(n16135), .A2(n16136), .ZN(n16037) );
  AND2_X1 U16198 ( .A1(n16031), .A2(n16033), .ZN(n16136) );
  AND2_X1 U16199 ( .A1(n16137), .A2(n16032), .ZN(n16135) );
  OR2_X1 U16200 ( .A1(n9389), .A2(n8962), .ZN(n16032) );
  OR2_X1 U16201 ( .A1(n16033), .A2(n16031), .ZN(n16137) );
  OR2_X1 U16202 ( .A1(n8958), .A2(n8903), .ZN(n16031) );
  INV_X1 U16203 ( .A(a_15_), .ZN(n8958) );
  OR2_X1 U16204 ( .A1(n16138), .A2(n16139), .ZN(n16033) );
  AND2_X1 U16205 ( .A1(n16027), .A2(n16029), .ZN(n16139) );
  AND2_X1 U16206 ( .A1(n16140), .A2(n16028), .ZN(n16138) );
  OR2_X1 U16207 ( .A1(n9389), .A2(n8966), .ZN(n16028) );
  OR2_X1 U16208 ( .A1(n16029), .A2(n16027), .ZN(n16140) );
  OR2_X1 U16209 ( .A1(n8962), .A2(n8903), .ZN(n16027) );
  INV_X1 U16210 ( .A(a_16_), .ZN(n8962) );
  OR2_X1 U16211 ( .A1(n16141), .A2(n16142), .ZN(n16029) );
  AND2_X1 U16212 ( .A1(n16023), .A2(n16025), .ZN(n16142) );
  AND2_X1 U16213 ( .A1(n16143), .A2(n16024), .ZN(n16141) );
  OR2_X1 U16214 ( .A1(n9389), .A2(n8970), .ZN(n16024) );
  OR2_X1 U16215 ( .A1(n16025), .A2(n16023), .ZN(n16143) );
  OR2_X1 U16216 ( .A1(n8966), .A2(n8903), .ZN(n16023) );
  INV_X1 U16217 ( .A(a_17_), .ZN(n8966) );
  OR2_X1 U16218 ( .A1(n16144), .A2(n16145), .ZN(n16025) );
  AND2_X1 U16219 ( .A1(n16019), .A2(n16021), .ZN(n16145) );
  AND2_X1 U16220 ( .A1(n16146), .A2(n16020), .ZN(n16144) );
  OR2_X1 U16221 ( .A1(n9389), .A2(n8974), .ZN(n16020) );
  OR2_X1 U16222 ( .A1(n16021), .A2(n16019), .ZN(n16146) );
  OR2_X1 U16223 ( .A1(n8970), .A2(n8903), .ZN(n16019) );
  INV_X1 U16224 ( .A(a_18_), .ZN(n8970) );
  OR2_X1 U16225 ( .A1(n16147), .A2(n16148), .ZN(n16021) );
  AND2_X1 U16226 ( .A1(n16015), .A2(n16017), .ZN(n16148) );
  AND2_X1 U16227 ( .A1(n16149), .A2(n16016), .ZN(n16147) );
  OR2_X1 U16228 ( .A1(n9389), .A2(n8978), .ZN(n16016) );
  OR2_X1 U16229 ( .A1(n16017), .A2(n16015), .ZN(n16149) );
  OR2_X1 U16230 ( .A1(n8974), .A2(n8903), .ZN(n16015) );
  INV_X1 U16231 ( .A(a_19_), .ZN(n8974) );
  OR2_X1 U16232 ( .A1(n16150), .A2(n16151), .ZN(n16017) );
  AND2_X1 U16233 ( .A1(n16011), .A2(n16013), .ZN(n16151) );
  AND2_X1 U16234 ( .A1(n16152), .A2(n16012), .ZN(n16150) );
  OR2_X1 U16235 ( .A1(n9389), .A2(n8982), .ZN(n16012) );
  OR2_X1 U16236 ( .A1(n16013), .A2(n16011), .ZN(n16152) );
  OR2_X1 U16237 ( .A1(n8978), .A2(n8903), .ZN(n16011) );
  INV_X1 U16238 ( .A(a_20_), .ZN(n8978) );
  OR2_X1 U16239 ( .A1(n16153), .A2(n16154), .ZN(n16013) );
  AND2_X1 U16240 ( .A1(n16007), .A2(n16009), .ZN(n16154) );
  AND2_X1 U16241 ( .A1(n16155), .A2(n16008), .ZN(n16153) );
  OR2_X1 U16242 ( .A1(n9389), .A2(n8986), .ZN(n16008) );
  OR2_X1 U16243 ( .A1(n16009), .A2(n16007), .ZN(n16155) );
  OR2_X1 U16244 ( .A1(n8982), .A2(n8903), .ZN(n16007) );
  INV_X1 U16245 ( .A(a_21_), .ZN(n8982) );
  OR2_X1 U16246 ( .A1(n16156), .A2(n16157), .ZN(n16009) );
  AND2_X1 U16247 ( .A1(n16003), .A2(n16005), .ZN(n16157) );
  AND2_X1 U16248 ( .A1(n16158), .A2(n16004), .ZN(n16156) );
  OR2_X1 U16249 ( .A1(n9389), .A2(n8990), .ZN(n16004) );
  OR2_X1 U16250 ( .A1(n16005), .A2(n16003), .ZN(n16158) );
  OR2_X1 U16251 ( .A1(n8986), .A2(n8903), .ZN(n16003) );
  INV_X1 U16252 ( .A(a_22_), .ZN(n8986) );
  OR2_X1 U16253 ( .A1(n16159), .A2(n16160), .ZN(n16005) );
  AND2_X1 U16254 ( .A1(n15999), .A2(n16001), .ZN(n16160) );
  AND2_X1 U16255 ( .A1(n16161), .A2(n16000), .ZN(n16159) );
  OR2_X1 U16256 ( .A1(n9389), .A2(n8994), .ZN(n16000) );
  OR2_X1 U16257 ( .A1(n16001), .A2(n15999), .ZN(n16161) );
  OR2_X1 U16258 ( .A1(n8990), .A2(n8903), .ZN(n15999) );
  INV_X1 U16259 ( .A(a_23_), .ZN(n8990) );
  OR2_X1 U16260 ( .A1(n16162), .A2(n16163), .ZN(n16001) );
  AND2_X1 U16261 ( .A1(n15995), .A2(n15997), .ZN(n16163) );
  AND2_X1 U16262 ( .A1(n16164), .A2(n15996), .ZN(n16162) );
  OR2_X1 U16263 ( .A1(n9389), .A2(n8998), .ZN(n15996) );
  OR2_X1 U16264 ( .A1(n15997), .A2(n15995), .ZN(n16164) );
  OR2_X1 U16265 ( .A1(n8994), .A2(n8903), .ZN(n15995) );
  INV_X1 U16266 ( .A(a_24_), .ZN(n8994) );
  OR2_X1 U16267 ( .A1(n16165), .A2(n16166), .ZN(n15997) );
  AND2_X1 U16268 ( .A1(n15991), .A2(n15993), .ZN(n16166) );
  AND2_X1 U16269 ( .A1(n16167), .A2(n15992), .ZN(n16165) );
  OR2_X1 U16270 ( .A1(n9389), .A2(n9002), .ZN(n15992) );
  OR2_X1 U16271 ( .A1(n15993), .A2(n15991), .ZN(n16167) );
  OR2_X1 U16272 ( .A1(n8998), .A2(n8903), .ZN(n15991) );
  INV_X1 U16273 ( .A(a_25_), .ZN(n8998) );
  OR2_X1 U16274 ( .A1(n16168), .A2(n16169), .ZN(n15993) );
  AND2_X1 U16275 ( .A1(n15987), .A2(n15989), .ZN(n16169) );
  AND2_X1 U16276 ( .A1(n16170), .A2(n15988), .ZN(n16168) );
  OR2_X1 U16277 ( .A1(n9389), .A2(n9006), .ZN(n15988) );
  OR2_X1 U16278 ( .A1(n15989), .A2(n15987), .ZN(n16170) );
  OR2_X1 U16279 ( .A1(n9002), .A2(n8903), .ZN(n15987) );
  INV_X1 U16280 ( .A(a_26_), .ZN(n9002) );
  OR2_X1 U16281 ( .A1(n16171), .A2(n16172), .ZN(n15989) );
  AND2_X1 U16282 ( .A1(n15983), .A2(n15985), .ZN(n16172) );
  AND2_X1 U16283 ( .A1(n16173), .A2(n15984), .ZN(n16171) );
  OR2_X1 U16284 ( .A1(n9389), .A2(n9010), .ZN(n15984) );
  OR2_X1 U16285 ( .A1(n15985), .A2(n15983), .ZN(n16173) );
  OR2_X1 U16286 ( .A1(n9006), .A2(n8903), .ZN(n15983) );
  INV_X1 U16287 ( .A(a_27_), .ZN(n9006) );
  OR2_X1 U16288 ( .A1(n16174), .A2(n16175), .ZN(n15985) );
  AND2_X1 U16289 ( .A1(n15978), .A2(n15981), .ZN(n16175) );
  AND2_X1 U16290 ( .A1(n15980), .A2(n16176), .ZN(n16174) );
  OR2_X1 U16291 ( .A1(n15981), .A2(n15978), .ZN(n16176) );
  OR2_X1 U16292 ( .A1(n9010), .A2(n8903), .ZN(n15978) );
  INV_X1 U16293 ( .A(a_28_), .ZN(n9010) );
  OR2_X1 U16294 ( .A1(n9389), .A2(n9014), .ZN(n15981) );
  INV_X1 U16295 ( .A(a_29_), .ZN(n9014) );
  AND2_X1 U16296 ( .A1(n16177), .A2(n15977), .ZN(n15980) );
  OR2_X1 U16297 ( .A1(n9984), .A2(n16178), .ZN(n15977) );
  OR2_X1 U16298 ( .A1(n9389), .A2(n8903), .ZN(n16178) );
  INV_X1 U16299 ( .A(b_1_), .ZN(n8903) );
  INV_X1 U16300 ( .A(b_0_), .ZN(n9389) );
  OR2_X1 U16301 ( .A1(n9294), .A2(n8002), .ZN(n9984) );
  INV_X1 U16302 ( .A(a_30_), .ZN(n8002) );
  INV_X1 U16303 ( .A(a_31_), .ZN(n9294) );
  INV_X1 U16304 ( .A(n16179), .ZN(n16177) );
  AND2_X1 U16305 ( .A1(n15975), .A2(n15976), .ZN(n16179) );
  AND2_X1 U16306 ( .A1(a_29_), .A2(b_1_), .ZN(n15976) );
  AND2_X1 U16307 ( .A1(a_30_), .A2(b_0_), .ZN(n15975) );
endmodule

