module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, n3515, WX660, WX661, n3513, WX662, WX663,
         n3511, WX664, WX665, n3509, WX666, WX667, n3507, WX668, WX669, n3505,
         WX670, WX671, n3503, WX672, WX673, n3501, WX674, WX675, n3499, WX676,
         WX677, n3497, WX678, WX679, n3495, WX680, WX681, n3493, WX682, WX683,
         n3491, WX684, WX685, n3489, WX686, WX688, WX689, n3485, WX690, WX691,
         n3483, WX692, WX693, n3481, WX694, WX695, n3479, WX696, WX697, n3477,
         WX698, WX699, n3475, WX700, WX701, n3473, WX702, WX703, n3471, WX704,
         WX705, n3469, WX706, WX707, n3467, WX708, WX709, WX710, WX711, WX712,
         WX713, WX714, WX715, WX716, WX717, WX718, WX719, WX720, WX721, WX722,
         WX724, WX725, WX726, WX727, WX728, WX729, WX730, WX731, WX732, WX733,
         WX734, WX735, WX736, WX737, WX738, WX739, WX740, WX741, WX742, WX743,
         WX744, WX745, WX746, WX747, WX748, WX749, WX750, WX751, WX752, WX753,
         WX754, WX755, WX756, WX757, WX758, WX760, WX761, WX762, WX763, WX764,
         WX765, WX766, WX767, WX768, WX769, WX770, WX771, WX772, WX773, WX774,
         WX775, WX776, WX777, WX778, WX779, WX780, WX781, WX782, WX783, WX784,
         WX785, WX786, WX787, WX788, WX789, WX790, WX791, WX792, WX793, WX794,
         WX796, WX797, WX798, WX799, WX800, WX801, WX802, WX803, WX804, WX805,
         WX806, WX807, WX808, WX809, WX810, WX811, WX812, WX813, WX814, WX815,
         WX816, WX817, WX818, WX819, WX820, WX821, WX822, WX823, WX824, WX825,
         WX826, WX827, WX828, WX829, WX830, WX832, WX833, WX834, WX835, WX836,
         WX837, WX838, WX839, WX840, WX841, WX842, WX843, WX844, WX845, WX846,
         WX847, WX848, WX849, WX850, WX851, WX852, WX853, WX854, WX855, WX856,
         WX857, WX858, WX859, WX860, WX861, WX862, WX863, WX864, WX865, WX866,
         WX868, WX869, WX870, WX871, WX872, WX873, WX874, WX875, WX876, WX877,
         WX878, WX879, WX880, WX881, WX882, WX883, WX884, WX885, WX886, WX887,
         WX888, WX889, WX890, WX891, WX892, WX893, WX894, WX895, WX896, WX897,
         WX898, WX899, WX1264, DFF_160_n1, WX1266, WX1268, DFF_162_n1, WX1270,
         WX1272, DFF_164_n1, WX1274, DFF_165_n1, WX1276, DFF_166_n1, WX1278,
         DFF_167_n1, WX1280, DFF_168_n1, WX1282, DFF_169_n1, WX1284, WX1286,
         DFF_171_n1, WX1288, DFF_172_n1, WX1290, DFF_173_n1, WX1292,
         DFF_174_n1, WX1294, WX1296, DFF_176_n1, WX1298, DFF_177_n1, WX1300,
         DFF_178_n1, WX1302, WX1304, DFF_180_n1, WX1306, DFF_181_n1, WX1308,
         DFF_182_n1, WX1310, DFF_183_n1, WX1312, DFF_184_n1, WX1314,
         DFF_185_n1, WX1316, DFF_186_n1, WX1318, DFF_187_n1, WX1320,
         DFF_188_n1, WX1322, DFF_189_n1, WX1324, DFF_190_n1, WX1326,
         DFF_191_n1, WX1778, n8702, n8701, n8700, n8699, n8696, n8695, n8694,
         n8693, n8692, n8691, n8690, n8689, n8688, n8687, n8686, n8685, n8684,
         n8683, n8682, n8681, n8680, n8677, n8676, n8675, n8674, n8673, n8672,
         n8671, WX1839, n8670, WX1937, n8669, WX1939, n8668, WX1941, n8667,
         WX1943, n8666, WX1945, n8665, WX1947, n8664, WX1949, n8663, WX1951,
         n8662, WX1953, n8661, WX1955, WX1957, n8658, WX1959, n8657, WX1961,
         n8656, WX1963, n8655, WX1965, n8654, WX1967, n8653, WX1969, WX1970,
         WX1971, WX1972, WX1973, WX1974, WX1975, WX1976, WX1977, WX1978,
         WX1979, WX1980, WX1981, WX1982, WX1983, WX1984, WX1985, WX1986,
         WX1987, WX1988, WX1989, WX1990, WX1991, WX1993, WX1994, WX1995,
         WX1996, WX1997, WX1998, WX1999, WX2000, WX2001, WX2002, WX2003,
         WX2004, WX2005, WX2006, WX2007, WX2008, WX2009, WX2010, WX2011,
         WX2012, WX2013, WX2014, WX2015, WX2016, WX2017, WX2018, WX2019,
         WX2020, WX2021, WX2022, WX2023, WX2024, WX2025, WX2026, WX2027,
         WX2029, WX2030, WX2031, WX2032, WX2033, WX2034, WX2035, WX2036, n3783,
         WX2037, WX2038, WX2039, WX2040, WX2041, WX2042, WX2043, WX2044, n3775,
         WX2045, WX2046, WX2047, WX2048, WX2049, WX2050, WX2051, WX2052,
         WX2053, WX2054, WX2055, WX2056, n3763, WX2057, WX2058, WX2059, WX2060,
         WX2061, WX2062, WX2063, WX2065, WX2066, WX2067, WX2068, WX2069,
         WX2070, WX2071, WX2072, WX2073, WX2074, WX2075, WX2076, WX2077,
         WX2078, WX2079, WX2080, WX2081, WX2082, WX2083, WX2084, WX2085,
         WX2086, WX2087, WX2088, WX2089, WX2090, WX2091, WX2092, WX2093,
         WX2094, WX2095, WX2096, WX2097, WX2098, WX2099, WX2101, WX2102,
         WX2103, WX2104, WX2105, WX2106, WX2107, WX2108, WX2109, WX2110,
         WX2111, WX2112, WX2113, WX2114, WX2115, WX2116, WX2117, WX2118,
         WX2119, WX2120, WX2121, WX2122, WX2123, WX2124, WX2125, WX2126,
         WX2127, WX2128, WX2129, WX2130, WX2131, WX2132, WX2133, WX2134,
         WX2135, WX2137, WX2138, WX2139, WX2140, WX2141, WX2142, WX2143,
         WX2144, WX2145, WX2146, WX2147, WX2148, WX2149, WX2150, WX2151,
         WX2152, WX2153, WX2154, WX2155, WX2156, WX2157, WX2158, WX2159,
         WX2160, WX2161, WX2162, WX2163, WX2164, WX2165, WX2166, WX2167,
         WX2168, WX2169, WX2170, WX2171, WX2173, WX2174, WX2175, WX2176,
         WX2177, WX2178, WX2179, WX2180, WX2181, WX2182, WX2183, WX2184,
         WX2185, WX2186, WX2187, WX2188, WX2189, WX2190, WX2191, WX2192,
         WX2557, DFF_352_n1, WX2559, DFF_353_n1, WX2561, DFF_354_n1, WX2563,
         WX2565, DFF_356_n1, WX2567, DFF_357_n1, WX2569, DFF_358_n1, WX2571,
         WX2573, DFF_360_n1, WX2575, DFF_361_n1, WX2577, WX2579, DFF_363_n1,
         WX2581, DFF_364_n1, WX2583, DFF_365_n1, WX2585, DFF_366_n1, WX2587,
         WX2589, DFF_368_n1, WX2591, DFF_369_n1, WX2593, DFF_370_n1, WX2595,
         DFF_371_n1, WX2597, DFF_372_n1, WX2599, DFF_373_n1, WX2601,
         DFF_374_n1, WX2603, DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609,
         DFF_378_n1, WX2611, DFF_379_n1, WX2613, DFF_380_n1, WX2615,
         DFF_381_n1, WX2617, DFF_382_n1, WX2619, DFF_383_n1, WX3071, n8644,
         n8643, n8642, n8641, n8640, n8639, n8638, n8637, n8636, n8635, n8632,
         n8631, n8630, n8629, n8628, n8627, n8626, n8625, n8624, n8623, n8622,
         n8621, n8620, n8619, n8618, n8617, n8616, n8613, WX3132, n8612,
         WX3230, n8611, WX3232, n8610, WX3234, n8609, WX3236, n8608, WX3238,
         n8607, WX3240, n8606, WX3242, n8605, WX3244, n8604, WX3246, n8603,
         WX3248, n8602, WX3250, n8601, WX3252, n8600, WX3254, n8599, WX3256,
         n8598, WX3258, n8597, WX3260, WX3262, WX3263, WX3264, WX3265, WX3266,
         WX3267, WX3268, WX3269, WX3270, WX3271, WX3272, WX3273, WX3274,
         WX3275, WX3276, WX3277, WX3278, WX3279, WX3280, WX3281, WX3282,
         WX3283, WX3284, WX3285, WX3286, WX3287, WX3288, WX3289, WX3290,
         WX3291, WX3292, WX3293, WX3294, WX3295, WX3296, WX3298, WX3299,
         WX3300, WX3301, WX3302, WX3303, WX3304, WX3305, WX3306, WX3307,
         WX3308, WX3309, WX3310, WX3311, WX3312, WX3313, WX3314, WX3315,
         WX3316, WX3317, WX3318, WX3319, WX3320, WX3321, WX3322, WX3323,
         WX3324, WX3325, WX3326, WX3327, WX3328, WX3329, WX3330, WX3331,
         WX3332, WX3334, WX3335, WX3336, WX3337, WX3338, WX3339, WX3340,
         WX3341, n3739, WX3342, WX3343, WX3344, WX3345, n3735, WX3346, WX3347,
         WX3348, WX3349, WX3350, WX3351, WX3352, WX3353, WX3354, WX3355,
         WX3356, WX3357, WX3358, WX3359, WX3360, WX3361, WX3362, WX3363,
         WX3364, WX3365, WX3366, WX3367, WX3368, WX3370, WX3371, WX3372,
         WX3373, WX3374, WX3375, WX3376, WX3377, WX3378, WX3379, WX3380,
         WX3381, WX3382, WX3383, WX3384, WX3385, WX3386, WX3387, WX3388,
         WX3389, WX3390, WX3391, WX3392, WX3393, WX3394, WX3395, WX3396,
         WX3397, WX3398, WX3399, WX3400, WX3401, WX3402, WX3403, WX3404,
         WX3406, WX3407, WX3408, WX3409, WX3410, WX3411, WX3412, WX3413,
         WX3414, WX3415, WX3416, WX3417, WX3418, WX3419, WX3420, WX3421,
         WX3422, WX3423, WX3424, WX3425, WX3426, WX3427, WX3428, WX3429,
         WX3430, WX3431, WX3432, WX3433, WX3434, WX3435, WX3436, WX3437,
         WX3438, WX3440, WX3441, WX3442, WX3443, WX3444, WX3445, WX3446,
         WX3447, WX3448, WX3449, WX3450, WX3451, WX3452, WX3453, WX3454,
         WX3455, WX3456, WX3457, WX3458, WX3459, WX3460, WX3461, WX3462,
         WX3463, WX3464, WX3465, WX3466, WX3467, WX3468, WX3469, WX3470,
         WX3471, WX3472, WX3474, WX3475, WX3476, WX3477, WX3478, WX3479,
         WX3480, WX3481, WX3482, WX3483, WX3484, WX3485, WX3850, DFF_544_n1,
         WX3852, DFF_545_n1, WX3854, DFF_546_n1, WX3856, WX3858, DFF_548_n1,
         WX3860, DFF_549_n1, WX3862, DFF_550_n1, WX3864, DFF_551_n1, WX3866,
         DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872, DFF_555_n1, WX3874,
         DFF_556_n1, WX3876, DFF_557_n1, WX3878, DFF_558_n1, WX3880, WX3882,
         DFF_560_n1, WX3884, DFF_561_n1, WX3886, DFF_562_n1, WX3888,
         DFF_563_n1, WX3890, DFF_564_n1, WX3892, DFF_565_n1, WX3894,
         DFF_566_n1, WX3896, DFF_567_n1, WX3898, DFF_568_n1, WX3900,
         DFF_569_n1, WX3902, DFF_570_n1, WX3904, WX3906, DFF_572_n1, WX3908,
         DFF_573_n1, WX3910, DFF_574_n1, WX3912, DFF_575_n1, WX4364, n8586,
         n8585, n8584, n8583, n8582, n8581, n8580, n8579, n8578, n8577, n8576,
         n8573, n8572, n8571, n8570, n8569, n8568, n8567, n8566, n8565, n8564,
         n8563, n8562, n8561, n8560, n8559, n8558, n8555, WX4425, n8554,
         WX4523, n8553, WX4525, n8552, WX4527, n8551, WX4529, n8550, WX4531,
         n8549, WX4533, n8548, WX4535, n8547, WX4537, n8546, WX4539, n8545,
         WX4541, n8544, WX4543, n8543, WX4545, n8542, WX4547, n8541, WX4549,
         n8540, WX4551, WX4553, n8537, WX4555, WX4556, WX4557, WX4558, WX4559,
         WX4560, WX4561, WX4562, WX4563, WX4564, WX4565, WX4566, WX4567,
         WX4568, WX4569, WX4570, WX4571, WX4572, WX4573, WX4574, WX4575,
         WX4576, WX4577, WX4578, WX4579, WX4580, WX4581, WX4582, WX4583,
         WX4584, WX4585, WX4587, WX4588, WX4589, WX4590, WX4591, WX4592,
         WX4593, WX4594, WX4595, WX4596, WX4597, WX4598, WX4599, WX4600,
         WX4601, WX4602, WX4603, WX4604, WX4605, WX4606, WX4607, WX4608,
         WX4609, WX4610, WX4611, WX4612, WX4613, WX4614, WX4615, WX4616,
         WX4617, WX4618, WX4619, WX4621, WX4622, WX4623, WX4624, n3717, WX4625,
         WX4626, WX4627, WX4628, n3713, WX4629, WX4630, WX4631, WX4632, WX4633,
         WX4634, WX4635, WX4636, WX4637, WX4638, WX4639, WX4640, WX4641,
         WX4642, WX4643, WX4644, WX4645, WX4646, WX4647, WX4648, WX4649,
         WX4650, n3691, WX4651, WX4652, WX4653, WX4655, WX4656, WX4657, WX4658,
         WX4659, WX4660, WX4661, WX4662, WX4663, WX4664, WX4665, WX4666,
         WX4667, WX4668, WX4669, WX4670, WX4671, WX4672, WX4673, WX4674,
         WX4675, WX4676, WX4677, WX4678, WX4679, WX4680, WX4681, WX4682,
         WX4683, WX4684, WX4685, WX4686, WX4687, WX4689, WX4690, WX4691,
         WX4692, WX4693, WX4694, WX4695, WX4696, WX4697, WX4698, WX4699,
         WX4700, WX4701, WX4702, WX4703, WX4704, WX4705, WX4706, WX4707,
         WX4708, WX4709, WX4710, WX4711, WX4712, WX4713, WX4714, WX4715,
         WX4716, WX4717, WX4718, WX4719, WX4720, WX4721, WX4723, WX4724,
         WX4725, WX4726, WX4727, WX4728, WX4729, WX4730, WX4731, WX4732,
         WX4733, WX4734, WX4735, WX4736, WX4737, WX4738, WX4739, WX4740,
         WX4741, WX4742, WX4743, WX4744, WX4745, WX4746, WX4747, WX4748,
         WX4749, WX4750, WX4751, WX4752, WX4753, WX4754, WX4755, WX4757,
         WX4758, WX4759, WX4760, WX4761, WX4762, WX4763, WX4764, WX4765,
         WX4766, WX4767, WX4768, WX4769, WX4770, WX4771, WX4772, WX4773,
         WX4774, WX4775, WX4776, WX4777, WX4778, WX5143, DFF_736_n1, WX5145,
         DFF_737_n1, WX5147, DFF_738_n1, WX5149, WX5151, DFF_740_n1, WX5153,
         WX5155, DFF_742_n1, WX5157, DFF_743_n1, WX5159, DFF_744_n1, WX5161,
         DFF_745_n1, WX5163, WX5165, DFF_747_n1, WX5167, DFF_748_n1, WX5169,
         DFF_749_n1, WX5171, DFF_750_n1, WX5173, WX5175, DFF_752_n1, WX5177,
         DFF_753_n1, WX5179, DFF_754_n1, WX5181, DFF_755_n1, WX5183,
         DFF_756_n1, WX5185, DFF_757_n1, WX5187, WX5189, DFF_759_n1, WX5191,
         DFF_760_n1, WX5193, DFF_761_n1, WX5195, DFF_762_n1, WX5197,
         DFF_763_n1, WX5199, DFF_764_n1, WX5201, DFF_765_n1, WX5203,
         DFF_766_n1, WX5205, DFF_767_n1, WX5657, n8528, n8527, n8526, n8525,
         n8524, n8523, n8520, n8519, n8518, n8517, n8516, n8515, n8514, n8513,
         n8512, n8511, n8510, n8509, n8508, n8507, n8506, n8505, n8502, n8501,
         n8500, n8499, n8498, n8497, WX5718, n8496, WX5816, n8495, WX5818,
         n8494, WX5820, n8493, WX5822, n8492, WX5824, n8491, WX5826, n8490,
         WX5828, n8489, WX5830, n8488, WX5832, n8487, WX5834, WX5836, n8484,
         WX5838, n8483, WX5840, n8482, WX5842, n8481, WX5844, n8480, WX5846,
         n8479, WX5848, WX5849, WX5850, WX5851, WX5852, WX5853, WX5854, WX5855,
         WX5856, WX5857, WX5858, WX5859, WX5860, WX5861, WX5862, WX5863,
         WX5864, WX5865, WX5866, WX5867, WX5868, WX5870, WX5871, WX5872,
         WX5873, WX5874, WX5875, WX5876, WX5877, WX5878, WX5879, WX5880,
         WX5881, WX5882, WX5883, WX5884, WX5885, WX5886, WX5887, WX5888,
         WX5889, WX5890, WX5891, WX5892, WX5893, WX5894, WX5895, WX5896,
         WX5897, WX5898, WX5899, WX5900, WX5901, WX5902, WX5904, WX5905,
         WX5906, WX5907, WX5908, WX5909, WX5910, WX5911, WX5912, WX5913,
         WX5914, WX5915, WX5916, WX5917, WX5918, WX5919, WX5920, WX5921,
         WX5922, WX5923, WX5924, WX5925, WX5926, WX5927, WX5928, WX5929,
         WX5930, WX5931, WX5932, WX5933, n3669, WX5934, WX5935, WX5936, WX5938,
         WX5939, WX5940, WX5941, n3661, WX5942, WX5943, WX5944, WX5945, WX5946,
         WX5947, WX5948, WX5949, WX5950, WX5951, WX5952, WX5953, WX5954,
         WX5955, WX5956, WX5957, WX5958, WX5959, WX5960, WX5961, WX5962,
         WX5963, WX5964, WX5965, WX5966, WX5967, WX5968, WX5969, WX5970,
         WX5972, WX5973, WX5974, WX5975, WX5976, WX5977, WX5978, WX5979,
         WX5980, WX5981, WX5982, WX5983, WX5984, WX5985, WX5986, WX5987,
         WX5988, WX5989, WX5990, WX5991, WX5992, WX5993, WX5994, WX5995,
         WX5996, WX5997, WX5998, WX5999, WX6000, WX6001, WX6002, WX6003,
         WX6004, WX6006, WX6007, WX6008, WX6009, WX6010, WX6011, WX6012,
         WX6013, WX6014, WX6015, WX6016, WX6017, WX6018, WX6019, WX6020,
         WX6021, WX6022, WX6023, WX6024, WX6025, WX6026, WX6027, WX6028,
         WX6029, WX6030, WX6031, WX6032, WX6033, WX6034, WX6035, WX6036,
         WX6037, WX6038, WX6040, WX6041, WX6042, WX6043, WX6044, WX6045,
         WX6046, WX6047, WX6048, WX6049, WX6050, WX6051, WX6052, WX6053,
         WX6054, WX6055, WX6056, WX6057, WX6058, WX6059, WX6060, WX6061,
         WX6062, WX6063, WX6064, WX6065, WX6066, WX6067, WX6068, WX6069,
         WX6070, WX6071, WX6436, WX6438, DFF_929_n1, WX6440, DFF_930_n1,
         WX6442, WX6444, DFF_932_n1, WX6446, DFF_933_n1, WX6448, DFF_934_n1,
         WX6450, DFF_935_n1, WX6452, DFF_936_n1, WX6454, DFF_937_n1, WX6456,
         WX6458, DFF_939_n1, WX6460, DFF_940_n1, WX6462, DFF_941_n1, WX6464,
         DFF_942_n1, WX6466, WX6468, DFF_944_n1, WX6470, WX6472, DFF_946_n1,
         WX6474, DFF_947_n1, WX6476, DFF_948_n1, WX6478, DFF_949_n1, WX6480,
         DFF_950_n1, WX6482, DFF_951_n1, WX6484, DFF_952_n1, WX6486,
         DFF_953_n1, WX6488, DFF_954_n1, WX6490, DFF_955_n1, WX6492,
         DFF_956_n1, WX6494, DFF_957_n1, WX6496, DFF_958_n1, WX6498,
         DFF_959_n1, WX6950, n8470, n8467, n8466, n8465, n8464, n8463, n8462,
         n8461, n8460, n8459, n8458, n8457, n8456, n8455, n8454, n8453, n8452,
         n8449, n8448, n8447, n8446, n8445, n8444, n8443, n8442, n8441, n8440,
         n8439, WX7011, n8438, WX7109, n8437, WX7111, n8436, WX7113, n8435,
         WX7115, n8434, WX7117, WX7119, n8431, WX7121, n8430, WX7123, n8429,
         WX7125, n8428, WX7127, n8427, WX7129, n8426, WX7131, n8425, WX7133,
         n8424, WX7135, n8423, WX7137, n8422, WX7139, n8421, WX7141, WX7142,
         WX7143, WX7144, WX7145, WX7146, WX7147, WX7148, WX7149, WX7150,
         WX7151, WX7153, WX7154, WX7155, WX7156, WX7157, WX7158, WX7159,
         WX7160, WX7161, WX7162, WX7163, WX7164, WX7165, WX7166, WX7167,
         WX7168, WX7169, WX7170, WX7171, WX7172, WX7173, WX7174, WX7175,
         WX7176, WX7177, WX7178, WX7179, WX7180, WX7181, WX7182, WX7183,
         WX7184, WX7185, WX7187, WX7188, WX7189, WX7190, WX7191, WX7192,
         WX7193, WX7194, WX7195, WX7196, WX7197, WX7198, WX7199, WX7200,
         WX7201, WX7202, WX7203, WX7204, WX7205, WX7206, WX7207, WX7208,
         WX7209, WX7210, WX7211, WX7212, WX7213, WX7214, WX7215, WX7216, n3647,
         WX7217, WX7218, WX7219, WX7221, WX7222, WX7223, WX7224, n3639, WX7225,
         WX7226, WX7227, WX7228, n3635, WX7229, WX7230, WX7231, WX7232, WX7233,
         WX7234, WX7235, WX7236, WX7237, WX7238, WX7239, WX7240, WX7241,
         WX7242, WX7243, WX7244, WX7245, WX7246, WX7247, WX7248, WX7249,
         WX7250, WX7251, WX7252, WX7253, WX7255, WX7256, WX7257, WX7258,
         WX7259, WX7260, WX7261, WX7262, WX7263, WX7264, WX7265, WX7266,
         WX7267, WX7268, WX7269, WX7270, WX7271, WX7272, WX7273, WX7274,
         WX7275, WX7276, WX7277, WX7278, WX7279, WX7280, WX7281, WX7282,
         WX7283, WX7284, WX7285, WX7286, WX7287, WX7289, WX7290, WX7291,
         WX7292, WX7293, WX7294, WX7295, WX7296, WX7297, WX7298, WX7299,
         WX7300, WX7301, WX7302, WX7303, WX7304, WX7305, WX7306, WX7307,
         WX7308, WX7309, WX7310, WX7311, WX7312, WX7313, WX7314, WX7315,
         WX7316, WX7317, WX7318, WX7319, WX7320, WX7321, WX7323, WX7324,
         WX7325, WX7326, WX7327, WX7328, WX7329, WX7330, WX7331, WX7332,
         WX7333, WX7334, WX7335, WX7336, WX7337, WX7338, WX7339, WX7340,
         WX7341, WX7342, WX7343, WX7344, WX7345, WX7346, WX7347, WX7348,
         WX7349, WX7350, WX7351, WX7352, WX7353, WX7354, WX7355, WX7357,
         WX7358, WX7359, WX7360, WX7361, WX7362, WX7363, WX7364, WX7729,
         DFF_1120_n1, WX7731, DFF_1121_n1, WX7733, DFF_1122_n1, WX7735, WX7737,
         DFF_1124_n1, WX7739, DFF_1125_n1, WX7741, DFF_1126_n1, WX7743,
         DFF_1127_n1, WX7745, DFF_1128_n1, WX7747, DFF_1129_n1, WX7749, WX7751,
         DFF_1131_n1, WX7753, WX7755, DFF_1133_n1, WX7757, DFF_1134_n1, WX7759,
         WX7761, DFF_1136_n1, WX7763, DFF_1137_n1, WX7765, DFF_1138_n1, WX7767,
         DFF_1139_n1, WX7769, DFF_1140_n1, WX7771, DFF_1141_n1, WX7773,
         DFF_1142_n1, WX7775, DFF_1143_n1, WX7777, DFF_1144_n1, WX7779,
         DFF_1145_n1, WX7781, DFF_1146_n1, WX7783, DFF_1147_n1, WX7785,
         DFF_1148_n1, WX7787, WX7789, DFF_1150_n1, WX7791, DFF_1151_n1, WX8243,
         n8411, n8410, n8409, n8408, n8407, n8406, n8405, n8404, n8403, n8402,
         n8401, n8400, n8399, n8396, n8395, n8394, n8393, n8392, n8391, n8390,
         n8389, n8388, n8387, n8386, n8385, n8384, n8383, n8382, n8381, WX8304,
         WX8402, n8378, WX8404, n8377, WX8406, n8376, WX8408, n8375, WX8410,
         n8374, WX8412, n8373, WX8414, n8372, WX8416, n8371, WX8418, n8370,
         WX8420, n8369, WX8422, n8368, WX8424, n8367, WX8426, n8366, WX8428,
         n8365, WX8430, n8364, WX8432, n8363, WX8434, WX8436, WX8437, WX8438,
         WX8439, WX8440, WX8441, WX8442, WX8443, WX8444, WX8445, WX8446,
         WX8447, WX8448, WX8449, WX8450, WX8451, WX8452, WX8453, WX8454,
         WX8455, WX8456, WX8457, WX8458, WX8459, WX8460, WX8461, WX8462,
         WX8463, WX8464, WX8465, WX8466, WX8467, WX8468, WX8470, WX8471,
         WX8472, WX8473, WX8474, WX8475, WX8476, WX8477, WX8478, WX8479,
         WX8480, WX8481, WX8482, WX8483, WX8484, WX8485, WX8486, WX8487,
         WX8488, WX8489, WX8490, WX8491, WX8492, WX8493, WX8494, WX8495,
         WX8496, WX8497, WX8498, WX8499, n3625, WX8500, WX8501, WX8502, WX8504,
         WX8505, WX8506, WX8507, n3617, WX8508, WX8509, WX8510, WX8511, n3613,
         WX8512, WX8513, WX8514, WX8515, WX8516, WX8517, WX8518, WX8519,
         WX8520, WX8521, WX8522, WX8523, WX8524, WX8525, WX8526, WX8527,
         WX8528, WX8529, WX8530, WX8531, WX8532, WX8533, WX8534, WX8535,
         WX8536, WX8538, WX8539, WX8540, WX8541, WX8542, WX8543, WX8544,
         WX8545, WX8546, WX8547, WX8548, WX8549, WX8550, WX8551, WX8552,
         WX8553, WX8554, WX8555, WX8556, WX8557, WX8558, WX8559, WX8560,
         WX8561, WX8562, WX8563, WX8564, WX8565, WX8566, WX8567, WX8568,
         WX8569, WX8570, WX8572, WX8573, WX8574, WX8575, WX8576, WX8577,
         WX8578, WX8579, WX8580, WX8581, WX8582, WX8583, WX8584, WX8585,
         WX8586, WX8587, WX8588, WX8589, WX8590, WX8591, WX8592, WX8593,
         WX8594, WX8595, WX8596, WX8597, WX8598, WX8599, WX8600, WX8601,
         WX8602, WX8603, WX8604, WX8606, WX8607, WX8608, WX8609, WX8610,
         WX8611, WX8612, WX8613, WX8614, WX8615, WX8616, WX8617, WX8618,
         WX8619, WX8620, WX8621, WX8622, WX8623, WX8624, WX8625, WX8626,
         WX8627, WX8628, WX8629, WX8630, WX8631, WX8632, WX8633, WX8634,
         WX8635, WX8636, WX8637, WX8638, WX8640, WX8641, WX8642, WX8643,
         WX8644, WX8645, WX8646, WX8647, WX8648, WX8649, WX8650, WX8651,
         WX8652, WX8653, WX8654, WX8655, WX8656, WX8657, WX9022, DFF_1312_n1,
         WX9024, DFF_1313_n1, WX9026, DFF_1314_n1, WX9028, WX9030, DFF_1316_n1,
         WX9032, DFF_1317_n1, WX9034, DFF_1318_n1, WX9036, WX9038, DFF_1320_n1,
         WX9040, DFF_1321_n1, WX9042, WX9044, DFF_1323_n1, WX9046, DFF_1324_n1,
         WX9048, DFF_1325_n1, WX9050, DFF_1326_n1, WX9052, WX9054, DFF_1328_n1,
         WX9056, DFF_1329_n1, WX9058, DFF_1330_n1, WX9060, DFF_1331_n1, WX9062,
         DFF_1332_n1, WX9064, DFF_1333_n1, WX9066, DFF_1334_n1, WX9068,
         DFF_1335_n1, WX9070, WX9072, DFF_1337_n1, WX9074, DFF_1338_n1, WX9076,
         DFF_1339_n1, WX9078, DFF_1340_n1, WX9080, DFF_1341_n1, WX9082,
         DFF_1342_n1, WX9084, DFF_1343_n1, WX9536, n8353, n8352, n8351, n8350,
         n8349, n8348, n8347, n8346, n8343, n8342, n8341, n8340, n8339, n8338,
         n8337, n8336, n8335, n8334, n8333, n8332, n8331, n8330, n8329, n8328,
         n8325, n8324, n8323, n8322, WX9597, n8321, WX9695, n8320, WX9697,
         n8319, WX9699, n8318, WX9701, n8317, WX9703, n8316, WX9705, n8315,
         WX9707, n8314, WX9709, n8313, WX9711, n8312, WX9713, n8311, WX9715,
         n8310, WX9717, WX9719, n8307, WX9721, n8306, WX9723, n8305, WX9725,
         n8304, WX9727, WX9728, WX9729, WX9730, WX9731, WX9732, WX9733, WX9734,
         WX9735, WX9736, WX9737, WX9738, WX9739, WX9740, WX9741, WX9742,
         WX9743, WX9744, WX9745, WX9746, WX9747, WX9748, WX9749, WX9750,
         WX9751, WX9753, WX9754, WX9755, WX9756, WX9757, WX9758, WX9759,
         WX9760, WX9761, WX9762, WX9763, WX9764, WX9765, WX9766, WX9767,
         WX9768, WX9769, WX9770, WX9771, WX9772, WX9773, WX9774, WX9775,
         WX9776, WX9777, WX9778, WX9779, WX9780, WX9781, WX9782, WX9783,
         WX9784, WX9785, WX9787, WX9788, WX9789, WX9790, WX9791, WX9792,
         WX9793, WX9794, n3591, WX9795, WX9796, WX9797, WX9798, WX9799, WX9800,
         WX9801, WX9802, WX9803, WX9804, WX9805, WX9806, WX9807, WX9808,
         WX9809, WX9810, WX9811, WX9812, WX9813, WX9814, WX9815, WX9816, n3569,
         WX9817, WX9818, WX9819, WX9821, WX9822, WX9823, WX9824, WX9825,
         WX9826, WX9827, WX9828, WX9829, WX9830, WX9831, WX9832, WX9833,
         WX9834, WX9835, WX9836, WX9837, WX9838, WX9839, WX9840, WX9841,
         WX9842, WX9843, WX9844, WX9845, WX9846, WX9847, WX9848, WX9849,
         WX9850, WX9851, WX9852, WX9853, WX9855, WX9856, WX9857, WX9858,
         WX9859, WX9860, WX9861, WX9862, WX9863, WX9864, WX9865, WX9866,
         WX9867, WX9868, WX9869, WX9870, WX9871, WX9872, WX9873, WX9874,
         WX9875, WX9876, WX9877, WX9878, WX9879, WX9880, WX9881, WX9882,
         WX9883, WX9884, WX9885, WX9886, WX9887, WX9889, WX9890, WX9891,
         WX9892, WX9893, WX9894, WX9895, WX9896, WX9897, WX9898, WX9899,
         WX9900, WX9901, WX9902, WX9903, WX9904, WX9905, WX9906, WX9907,
         WX9908, WX9909, WX9910, WX9911, WX9912, WX9913, WX9914, WX9915,
         WX9916, WX9917, WX9918, WX9919, WX9920, WX9921, WX9923, WX9924,
         WX9925, WX9926, WX9927, WX9928, WX9929, WX9930, WX9931, WX9932,
         WX9933, WX9934, WX9935, WX9936, WX9937, WX9938, WX9939, WX9940,
         WX9941, WX9942, WX9943, WX9944, WX9945, WX9946, WX9947, WX9948,
         WX9949, WX9950, WX10315, DFF_1504_n1, WX10317, DFF_1505_n1, WX10319,
         WX10321, WX10323, DFF_1508_n1, WX10325, DFF_1509_n1, WX10327,
         DFF_1510_n1, WX10329, DFF_1511_n1, WX10331, DFF_1512_n1, WX10333,
         DFF_1513_n1, WX10335, WX10337, DFF_1515_n1, WX10339, DFF_1516_n1,
         WX10341, DFF_1517_n1, WX10343, DFF_1518_n1, WX10345, DFF_1519_n1,
         WX10347, DFF_1520_n1, WX10349, DFF_1521_n1, WX10351, DFF_1522_n1,
         WX10353, WX10355, DFF_1524_n1, WX10357, DFF_1525_n1, WX10359,
         DFF_1526_n1, WX10361, DFF_1527_n1, WX10363, DFF_1528_n1, WX10365,
         DFF_1529_n1, WX10367, DFF_1530_n1, WX10369, DFF_1531_n1, WX10371,
         DFF_1532_n1, WX10373, DFF_1533_n1, WX10375, DFF_1534_n1, WX10377,
         DFF_1535_n1, WX10829, n8295, n8294, n8293, n8290, n8289, n8288, n8287,
         n8286, n8285, n8284, n8283, n8282, n8281, n8280, n8279, n8278, n8277,
         n8276, n8275, n8272, n8271, n8270, n8269, n8268, n8267, n8266, n8265,
         n8264, WX10890, n8263, WX10988, n8262, WX10990, n8261, WX10992, n8260,
         WX10994, n8259, WX10996, n8258, WX10998, n8257, WX11000, WX11002,
         n8254, WX11004, n8253, WX11006, n8252, WX11008, n8251, WX11010, n8250,
         WX11012, n8249, WX11014, n8248, WX11016, n8247, WX11018, n8246,
         WX11020, WX11021, WX11022, WX11023, WX11024, WX11025, WX11026,
         WX11027, WX11028, WX11029, WX11030, WX11031, WX11032, WX11033,
         WX11034, WX11036, WX11037, WX11038, WX11039, WX11040, WX11041,
         WX11042, WX11043, WX11044, WX11045, WX11046, WX11047, WX11048,
         WX11049, WX11050, WX11051, WX11052, WX11053, WX11054, WX11055,
         WX11056, WX11057, WX11058, WX11059, WX11060, WX11061, WX11062,
         WX11063, WX11064, WX11065, WX11066, WX11067, WX11068, WX11070,
         WX11071, WX11072, WX11073, WX11074, WX11075, WX11076, WX11077,
         WX11078, WX11079, WX11080, WX11081, WX11082, WX11083, WX11084,
         WX11085, WX11086, WX11087, WX11088, WX11089, WX11090, WX11091,
         WX11092, WX11093, WX11094, WX11095, WX11096, WX11097, WX11098,
         WX11099, n3547, WX11100, WX11101, WX11102, WX11104, WX11105, WX11106,
         WX11107, n3539, WX11108, WX11109, WX11110, WX11111, n3535, WX11112,
         WX11113, WX11114, WX11115, WX11116, WX11117, WX11118, WX11119,
         WX11120, WX11121, WX11122, WX11123, WX11124, WX11125, WX11126,
         WX11127, WX11128, WX11129, WX11130, WX11131, WX11132, WX11133,
         WX11134, WX11135, WX11136, WX11138, WX11139, WX11140, WX11141,
         WX11142, WX11143, WX11144, WX11145, WX11146, WX11147, WX11148,
         WX11149, WX11150, WX11151, WX11152, WX11153, WX11154, WX11155,
         WX11156, WX11157, WX11158, WX11159, WX11160, WX11161, WX11162,
         WX11163, WX11164, WX11165, WX11166, WX11167, WX11168, WX11169,
         WX11170, WX11172, WX11173, WX11174, WX11175, WX11176, WX11177,
         WX11178, WX11179, WX11180, WX11181, WX11182, WX11183, WX11184,
         WX11185, WX11186, WX11187, WX11188, WX11189, WX11190, WX11191,
         WX11192, WX11193, WX11194, WX11195, WX11196, WX11197, WX11198,
         WX11199, WX11200, WX11201, WX11202, WX11203, WX11204, WX11206,
         WX11207, WX11208, WX11209, WX11210, WX11211, WX11212, WX11213,
         WX11214, WX11215, WX11216, WX11217, WX11218, WX11219, WX11220,
         WX11221, WX11222, WX11223, WX11224, WX11225, WX11226, WX11227,
         WX11228, WX11229, WX11230, WX11231, WX11232, WX11233, WX11234,
         WX11235, WX11236, WX11237, WX11238, WX11240, WX11241, WX11242,
         WX11243, WX11608, DFF_1696_n1, WX11610, DFF_1697_n1, WX11612,
         DFF_1698_n1, WX11614, WX11616, DFF_1700_n1, WX11618, DFF_1701_n1,
         WX11620, DFF_1702_n1, WX11622, DFF_1703_n1, WX11624, DFF_1704_n1,
         WX11626, DFF_1705_n1, WX11628, WX11630, DFF_1707_n1, WX11632,
         DFF_1708_n1, WX11634, DFF_1709_n1, WX11636, WX11638, WX11640,
         DFF_1712_n1, WX11642, DFF_1713_n1, WX11644, DFF_1714_n1, WX11646,
         DFF_1715_n1, WX11648, DFF_1716_n1, WX11650, DFF_1717_n1, WX11652,
         DFF_1718_n1, WX11654, DFF_1719_n1, WX11656, DFF_1720_n1, WX11658,
         DFF_1721_n1, WX11660, DFF_1722_n1, WX11662, DFF_1723_n1, WX11664,
         DFF_1724_n1, WX11666, DFF_1725_n1, WX11668, DFF_1726_n1, WX11670,
         n2245, n2153, n3278, n2152, n2148, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4,
         Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         Tj_Trigger, Stage4, Stage1_1, Stage1_2, Stage1_3, Stage1_4, Stage1,
         Stage2_i, Stage2_7, Stage2_8, Stage2_9, Stage2_10, Stage2, Stage3_i,
         Stage3_12, Stage3_13, Stage3_14, Stage3_15, Stage4_i, Stage4_17,
         Stage4_18, Stage4_19, Stage4_20, Stage4_21, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n2181, n2182, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7862, n7863, n7865, n7866, n7867,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7886, n7887, n7888, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7937, n7938, n7940, n7941, n7942,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7957, n7958, n7960, n7961, n7962, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7977,
         n7978, n7980, n7981, n7982, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8030, n8031,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8051, n8052, n8053,
         n8054, n8055, n8056, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8093, n8094, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8255, n8256, n8273, n8274, n8291, n8292, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8308, n8309, n8326,
         n8327, n8344, n8345, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8362, n8379, n8380, n8397, n8398, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8433, n8450, n8451, n8468, n8469, n8471,
         n8472, n8474, n8475, n8476, n8477, n8478, n8485, n8486, n8503, n8504,
         n8521, n8522, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8538, n8539, n8556, n8557, n8574, n8575, n8587, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8614, n8615, n8633, n8634, n8645,
         n8646, n8648, n8649, n8650, n8651, n8652, n8659, n8660, n8678, n8679,
         n8697, n8698, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, U3558_n1, U3871_n1, U3991_n1, U5716_n1, U5717_n1, U5718_n1,
         U5719_n1, U5720_n1, U5721_n1, U5722_n1, U5723_n1, U5724_n1, U5725_n1,
         U5726_n1, U5727_n1, U5728_n1, U5729_n1, U5730_n1, U5731_n1, U5732_n1,
         U5733_n1, U5734_n1, U5735_n1, U5736_n1, U5737_n1, U5738_n1, U5739_n1,
         U5740_n1, U5741_n1, U5742_n1, U5743_n1, U5744_n1, U5745_n1, U5746_n1,
         U5747_n1, U5748_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1, U5753_n1,
         U5754_n1, U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1, U5760_n1,
         U5761_n1, U5762_n1, U5763_n1, U5764_n1, U5765_n1, U5766_n1, U5767_n1,
         U5768_n1, U5769_n1, U5770_n1, U5771_n1, U5772_n1, U5773_n1, U5774_n1,
         U5775_n1, U5776_n1, U5777_n1, U5778_n1, U5779_n1, U5780_n1, U5781_n1,
         U5782_n1, U5783_n1, U5784_n1, U5785_n1, U5786_n1, U5787_n1, U5788_n1,
         U5789_n1, U5790_n1, U5791_n1, U5792_n1, U5793_n1, U5794_n1, U5795_n1,
         U5796_n1, U5797_n1, U5798_n1, U5799_n1, U5800_n1, U5801_n1, U5802_n1,
         U5803_n1, U5804_n1, U5805_n1, U5806_n1, U5807_n1, U5808_n1, U5809_n1,
         U5810_n1, U5811_n1, U5812_n1, U5813_n1, U5814_n1, U5815_n1, U5816_n1,
         U5817_n1, U5818_n1, U5819_n1, U5820_n1, U5821_n1, U5822_n1, U5823_n1,
         U5824_n1, U5825_n1, U5826_n1, U5827_n1, U5828_n1, U5829_n1, U5830_n1,
         U5831_n1, U5832_n1, U5833_n1, U5834_n1, U5835_n1, U5836_n1, U5837_n1,
         U5838_n1, U5839_n1, U5840_n1, U5841_n1, U5842_n1, U5843_n1, U5844_n1,
         U5845_n1, U5846_n1, U5847_n1, U5848_n1, U5849_n1, U5850_n1, U5851_n1,
         U5852_n1, U5853_n1, U5854_n1, U5855_n1, U5856_n1, U5857_n1, U5858_n1,
         U5859_n1, U5860_n1, U5861_n1, U5862_n1, U5863_n1, U5864_n1, U5865_n1,
         U5866_n1, U5867_n1, U5868_n1, U5869_n1, U5870_n1, U5871_n1, U5872_n1,
         U5873_n1, U5874_n1, U5875_n1, U5876_n1, U5877_n1, U5878_n1, U5879_n1,
         U5880_n1, U5881_n1, U5882_n1, U5883_n1, U5884_n1, U5885_n1, U5886_n1,
         U5887_n1, U5888_n1, U5889_n1, U5890_n1, U5891_n1, U5892_n1, U5893_n1,
         U5894_n1, U5895_n1, U5896_n1, U5897_n1, U5898_n1, U5899_n1, U5900_n1,
         U5901_n1, U5902_n1, U5903_n1, U5904_n1, U5905_n1, U5906_n1, U5907_n1,
         U5908_n1, U5909_n1, U5910_n1, U5911_n1, U5912_n1, U5913_n1, U5914_n1,
         U5915_n1, U5916_n1, U5917_n1, U5918_n1, U5919_n1, U5920_n1, U5921_n1,
         U5922_n1, U5923_n1, U5924_n1, U5925_n1, U5926_n1, U5927_n1, U5928_n1,
         U5929_n1, U5930_n1, U5931_n1, U5932_n1, U5933_n1, U5934_n1, U5935_n1,
         U5936_n1, U5937_n1, U5938_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1,
         U5943_n1, U5944_n1, U5945_n1, U5946_n1, U5947_n1, U5948_n1, U5949_n1,
         U5950_n1, U5951_n1, U5952_n1, U5953_n1, U5954_n1, U5955_n1, U5956_n1,
         U5957_n1, U5958_n1, U5959_n1, U5960_n1, U5961_n1, U5962_n1, U5963_n1,
         U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1, U5969_n1, U5970_n1,
         U5971_n1, U5972_n1, U5973_n1, U5974_n1, U5975_n1, U5976_n1, U5977_n1,
         U5978_n1, U5979_n1, U5980_n1, U5981_n1, U5982_n1, U5983_n1, U5984_n1,
         U5985_n1, U5986_n1, U5987_n1, U5988_n1, U5989_n1, U5990_n1, U5991_n1,
         U5992_n1, U5993_n1, U5994_n1, U5995_n1, U5996_n1, U5997_n1, U5998_n1,
         U5999_n1, U6000_n1, U6001_n1, U6002_n1, U6003_n1, U6004_n1, U6005_n1,
         U6006_n1, U6007_n1, U6008_n1, U6009_n1, U6010_n1, U6011_n1, U6012_n1,
         U6013_n1, U6014_n1, U6015_n1, U6016_n1, U6017_n1, U6018_n1, U6019_n1,
         U6020_n1, U6021_n1, U6022_n1, U6023_n1, U6024_n1, U6025_n1, U6026_n1,
         U6027_n1, U6028_n1, U6029_n1, U6030_n1, U6031_n1, U6032_n1, U6033_n1,
         U6034_n1, U6035_n1, U6036_n1, U6037_n1, U6038_n1, U6039_n1, U6040_n1,
         U6041_n1, U6042_n1, U6043_n1, U6044_n1, U6045_n1, U6046_n1, U6047_n1,
         U6048_n1, U6049_n1, U6050_n1, U6051_n1, U6052_n1, U6053_n1, U6054_n1,
         U6055_n1, U6056_n1, U6057_n1, U6058_n1, U6059_n1, U6060_n1, U6061_n1,
         U6062_n1, U6063_n1, U6064_n1, U6065_n1, U6066_n1, U6067_n1, U6068_n1,
         U6069_n1, U6070_n1, U6071_n1, U6072_n1, U6073_n1, U6074_n1, U6075_n1,
         U6076_n1, U6077_n1, U6078_n1, U6079_n1, U6080_n1, U6081_n1, U6082_n1,
         U6083_n1, U6084_n1, U6085_n1, U6086_n1, U6087_n1, U6088_n1, U6089_n1,
         U6090_n1, U6091_n1, U6092_n1, U6093_n1, U6094_n1, U6095_n1, U6096_n1,
         U6097_n1, U6098_n1, U6099_n1, U6100_n1, U6101_n1, U6102_n1, U6103_n1,
         U6104_n1, U6105_n1, U6106_n1, U6107_n1, U6108_n1, U6109_n1, U6110_n1,
         U6111_n1, U6112_n1, U6113_n1, U6114_n1, U6115_n1, U6116_n1, U6117_n1,
         U6118_n1, U6119_n1, U6120_n1, U6121_n1, U6122_n1, U6123_n1, U6124_n1,
         U6125_n1, U6126_n1, U6127_n1, U6128_n1, U6129_n1, U6130_n1, U6131_n1,
         U6132_n1, U6133_n1, U6134_n1, U6135_n1, U6136_n1, U6137_n1, U6138_n1,
         U6139_n1, U6140_n1, U6141_n1, U6142_n1, U6143_n1, U6144_n1, U6145_n1,
         U6146_n1, U6147_n1, U6148_n1, U6149_n1, U6150_n1, U6151_n1, U6152_n1,
         U6153_n1, U6154_n1, U6155_n1, U6156_n1, U6157_n1, U6158_n1, U6159_n1,
         U6160_n1, U6161_n1, U6162_n1, U6163_n1, U6164_n1, U6165_n1, U6166_n1,
         U6167_n1, U6168_n1, U6169_n1, U6170_n1, U6171_n1, U6172_n1, U6173_n1,
         U6174_n1, U6175_n1, U6176_n1, U6177_n1, U6178_n1, U6179_n1, U6180_n1,
         U6181_n1, U6182_n1, U6183_n1, U6184_n1, U6185_n1, U6186_n1, U6187_n1,
         U6188_n1, U6189_n1, U6190_n1, U6191_n1, U6192_n1, U6193_n1, U6194_n1,
         U6195_n1, U6196_n1, U6197_n1, U6198_n1, U6199_n1, U6200_n1, U6201_n1,
         U6202_n1, U6203_n1, U6204_n1, U6205_n1, U6206_n1, U6207_n1, U6208_n1,
         U6209_n1, U6210_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1,
         U6216_n1, U6217_n1, U6218_n1, U6219_n1, U6220_n1, U6221_n1, U6222_n1,
         U6223_n1, U6224_n1, U6225_n1, U6226_n1, U6227_n1, U6228_n1, U6229_n1,
         U6230_n1, U6231_n1, U6232_n1, U6233_n1, U6234_n1, U6235_n1, U6236_n1,
         U6237_n1, U6238_n1, U6239_n1, U6240_n1, U6241_n1, U6242_n1, U6243_n1,
         U6244_n1, U6245_n1, U6246_n1, U6247_n1, U6248_n1, U6249_n1, U6250_n1,
         U6251_n1, U6252_n1, U6253_n1, U6254_n1, U6255_n1, U6256_n1, U6257_n1,
         U6258_n1, U6259_n1, U6260_n1, U6261_n1, U6262_n1, U6263_n1, U6264_n1,
         U6265_n1, U6266_n1, U6267_n1, U6268_n1, U6269_n1, U6270_n1, U6271_n1,
         U6272_n1, U6273_n1, U6274_n1, U6275_n1, U6276_n1, U6277_n1, U6278_n1,
         U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1,
         U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1,
         U6293_n1, U6294_n1, U6295_n1, U6296_n1, U6297_n1, U6298_n1, U6299_n1,
         U6300_n1, U6301_n1, U6302_n1, U6303_n1, U6304_n1, U6305_n1, U6306_n1,
         U6307_n1, U6308_n1, U6309_n1, U6310_n1, U6311_n1, U6312_n1, U6313_n1,
         U6314_n1, U6315_n1, U6316_n1, U6317_n1, U6318_n1, U6319_n1, U6320_n1,
         U6321_n1, U6322_n1, U6323_n1, U6324_n1, U6325_n1, U6326_n1, U6327_n1,
         U6328_n1, U6329_n1, U6330_n1, U6331_n1, U6332_n1, U6333_n1, U6334_n1,
         U6335_n1, U6336_n1, U6337_n1, U6338_n1, U6339_n1, U6340_n1, U6341_n1,
         U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1,
         U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1,
         U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1,
         U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1,
         U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6376_n1,
         U6377_n1, U6378_n1, U6379_n1, U6380_n1, U6381_n1, U6382_n1, U6383_n1,
         U6384_n1, U6385_n1, U6386_n1, U6387_n1, U6388_n1, U6389_n1, U6390_n1,
         U6391_n1, U6392_n1, U6393_n1, U6394_n1, U6395_n1, U6396_n1, U6397_n1,
         U6398_n1, U6399_n1, U6400_n1, U6401_n1, U6402_n1, U6403_n1, U6404_n1,
         U6405_n1, U6406_n1, U6407_n1, U6408_n1, U6409_n1, U6410_n1, U6411_n1,
         U6412_n1, U6413_n1, U6414_n1, U6415_n1, U6416_n1, U6417_n1, U6418_n1,
         U6419_n1, U6420_n1, U6421_n1, U6422_n1, U6423_n1, U6424_n1, U6425_n1,
         U6426_n1, U6427_n1, U6428_n1, U6429_n1, U6430_n1, U6431_n1, U6432_n1,
         U6433_n1, U6434_n1, U6435_n1, U6436_n1, U6437_n1, U6438_n1, U6439_n1,
         U6440_n1, U6441_n1, U6442_n1, U6443_n1, U6444_n1, U6445_n1, U6446_n1,
         U6447_n1, U6448_n1, U6449_n1, U6450_n1, U6451_n1, U6452_n1, U6453_n1,
         U6454_n1, U6455_n1, U6456_n1, U6457_n1, U6458_n1, U6459_n1, U6460_n1,
         U6461_n1, U6462_n1, U6463_n1, U6464_n1, U6465_n1, U6466_n1, U6467_n1,
         U6468_n1, U6469_n1, U6470_n1, U6471_n1, U6472_n1, U6473_n1, U6474_n1,
         U6475_n1, U6476_n1, U6477_n1, U6478_n1, U6479_n1, U6480_n1, U6481_n1,
         U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n9341), .CLK(n9493), .Q(
        WX485) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n9482), .CLK(n9495), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n9482), .CLK(n9495), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n9482), .CLK(n9495), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n9482), .CLK(n9495), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n9482), .CLK(n9495), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n9482), .CLK(n9495), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n9482), .CLK(n9495), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n9482), .CLK(n9495), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n9340), .CLK(n9494), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n9337), .CLK(n9494), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n9338), .CLK(n9494), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n9341), .CLK(n9494), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n9342), .CLK(n9494), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(test_se), .CLK(n9494), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n9343), .CLK(n9494), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n9339), .CLK(n9494), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n9340), .CLK(n9494), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n9337), .CLK(n9494), .Q(
        WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n9338), .CLK(n9494), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n9341), .CLK(n9494), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(test_se), .CLK(n9493), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n9343), .CLK(n9493), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n9339), .CLK(n9493), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n9340), .CLK(n9493), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n9337), .CLK(n9493), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n9338), .CLK(n9493), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n9341), .CLK(n9493), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n9339), .CLK(n9493), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n9340), .CLK(n9493), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n9337), .CLK(n9493), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n9338), .CLK(n9493), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n9482), .CLK(n9495), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n9482), .CLK(n9495), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n9482), .CLK(n9495), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n9482), .CLK(n9495), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n9481), .CLK(n9496), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n9481), .CLK(n9496), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n9481), .CLK(n9496), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n9481), .CLK(n9496), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n9481), .CLK(n9496), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n9481), .CLK(n9496), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n9480), .CLK(n9497), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n9480), .CLK(n9497), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n9480), .CLK(n9497), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n9480), .CLK(n9497), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n9480), .CLK(n9497), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n9479), .CLK(n9498), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n9479), .CLK(n9498), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n9479), .CLK(n9498), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n9478), .CLK(n9499), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n9478), .CLK(n9499), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n9478), .CLK(n9499), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n9477), .CLK(n9500), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n9477), .CLK(n9500), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n9477), .CLK(n9500), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n9476), .CLK(n9501), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n9476), .CLK(n9501), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n9476), .CLK(n9501), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n9475), .CLK(n9502), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n9475), .CLK(n9502), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n9475), .CLK(n9502), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n9474), .CLK(n9503), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n9474), .CLK(n9503), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n9474), .CLK(n9503), .Q(
        WX709), .QN(n8772) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n9473), .CLK(n9504), .Q(
        WX711), .QN(n8660) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n9473), .CLK(n9504), .Q(
        WX713), .QN(n8709) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n9481), .CLK(n9496), .Q(
        WX715), .QN(n8718) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n9481), .CLK(n9496), .Q(
        WX717), .QN(n8724) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n9481), .CLK(n9496), .Q(
        WX719), .QN(n8727) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n9481), .CLK(n9496), .Q(
        WX721), .QN(n8736) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n9481), .CLK(n9496), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n9481), .CLK(n9496), .Q(
        WX725), .QN(n8747) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n9480), .CLK(n9497), .Q(
        WX727), .QN(n8759) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n9480), .CLK(n9497), .Q(
        WX729), .QN(n8765) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n9480), .CLK(n9497), .Q(
        WX731) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n9480), .CLK(n9497), .Q(
        WX733), .QN(n8706) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n9480), .CLK(n9497), .Q(
        WX735), .QN(n8721) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n9479), .CLK(n9498), .Q(
        WX737), .QN(n8733) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n9479), .CLK(n9498), .Q(
        WX739), .QN(n8748) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n9479), .CLK(n9498), .Q(
        WX741), .QN(n8762) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n9479), .CLK(n9498), .Q(
        WX743), .QN(n8777) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n9478), .CLK(n9499), .Q(
        WX745), .QN(n8712) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n9478), .CLK(n9499), .Q(
        WX747), .QN(n8739) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n9478), .CLK(n9499), .Q(
        WX749), .QN(n8785) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n9477), .CLK(n9500), .Q(
        WX751), .QN(n8730) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n9477), .CLK(n9500), .Q(
        WX753), .QN(n8740) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n9477), .CLK(n9500), .Q(
        WX755), .QN(n8752) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n9476), .CLK(n9501), .Q(
        WX757), .QN(n8780) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n9476), .CLK(n9501), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n9476), .CLK(n9501), .Q(
        WX761), .QN(n8755) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n9475), .CLK(n9502), .Q(
        WX763), .QN(n8758) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n9475), .CLK(n9502), .Q(
        WX765), .QN(n8703) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n9475), .CLK(n9502), .Q(
        WX767), .QN(n8778) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n9474), .CLK(n9503), .Q(
        WX769), .QN(n8714) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n9474), .CLK(n9503), .Q(
        WX771), .QN(n8786) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n9474), .CLK(n9503), .Q(
        WX773), .QN(n8773) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n9473), .CLK(n9504), .Q(
        WX775), .QN(n8678) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n9473), .CLK(n9504), .Q(
        WX777), .QN(n8707) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n9473), .CLK(n9504), .Q(
        WX779), .QN(n8716) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n9473), .CLK(n9504), .Q(
        WX781), .QN(n8722) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n9473), .CLK(n9504), .Q(
        WX783), .QN(n8725) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n9472), .CLK(n9505), .Q(
        WX785), .QN(n8734) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n9472), .CLK(n9505), .Q(
        WX787), .QN(n8743) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n9472), .CLK(n9505), .Q(
        WX789), .QN(n8745) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n9472), .CLK(n9505), .Q(
        WX791), .QN(n8760) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n9472), .CLK(n9505), .Q(
        WX793), .QN(n8766) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n9472), .CLK(n9505), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n9480), .CLK(n9497), 
        .Q(WX797), .QN(n8704) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n9480), .CLK(n9497), .Q(
        WX799), .QN(n8719) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n9479), .CLK(n9498), .Q(
        WX801), .QN(n8731) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n9479), .CLK(n9498), .Q(
        WX803), .QN(n8749) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n9479), .CLK(n9498), .Q(
        WX805), .QN(n8763) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n9479), .CLK(n9498), .Q(
        WX807), .QN(n8775) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n9478), .CLK(n9499), .Q(
        WX809), .QN(n8710) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n9478), .CLK(n9499), .Q(
        WX811), .QN(n8737) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n9478), .CLK(n9499), .Q(
        WX813), .QN(n8783) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n9477), .CLK(n9500), .Q(
        WX815), .QN(n8728) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n9477), .CLK(n9500), .Q(
        WX817), .QN(n8741) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n9477), .CLK(n9500), .Q(
        WX819), .QN(n8750) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n9476), .CLK(n9501), .Q(
        WX821), .QN(n8781) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n9476), .CLK(n9501), .Q(
        WX823), .QN(n8768) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n9476), .CLK(n9501), .Q(
        WX825), .QN(n8753) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n9475), .CLK(n9502), .Q(
        WX827), .QN(n8756) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n9475), .CLK(n9502), .Q(
        WX829), .QN(n8697) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n9475), .CLK(n9502), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n9474), .CLK(n9503), 
        .Q(WX833) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n9474), .CLK(n9503), .Q(
        WX835), .QN(n8787) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n9474), .CLK(n9503), .Q(
        WX837), .QN(n8774) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n9473), .CLK(n9504), .Q(
        WX839), .QN(n8679) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n9473), .CLK(n9504), .Q(
        WX841), .QN(n8708) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n9473), .CLK(n9504), .Q(
        WX843), .QN(n8717) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n9473), .CLK(n9504), .Q(
        WX845), .QN(n8723) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n9473), .CLK(n9504), .Q(
        WX847), .QN(n8726) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n9472), .CLK(n9505), .Q(
        WX849), .QN(n8735) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n9472), .CLK(n9505), .Q(
        WX851), .QN(n8744) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n9472), .CLK(n9505), .Q(
        WX853), .QN(n8746) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n9472), .CLK(n9505), .Q(
        WX855), .QN(n8761) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n9472), .CLK(n9505), .Q(
        WX857), .QN(n8767) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n9472), .CLK(n9505), .Q(
        WX859), .QN(n8770) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n9471), .CLK(n9506), .Q(
        WX861), .QN(n8705) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n9471), .CLK(n9506), .Q(
        WX863), .QN(n8720) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n9471), .CLK(n9506), .Q(
        WX865), .QN(n8732) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n9471), .CLK(n9506), .Q(
        test_so8), .QN(n8797) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n9479), .CLK(n9498), 
        .Q(WX869), .QN(n8764) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n9478), .CLK(n9499), .Q(
        WX871), .QN(n8776) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n9478), .CLK(n9499), .Q(
        WX873), .QN(n8711) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n9478), .CLK(n9499), .Q(
        WX875), .QN(n8738) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n9477), .CLK(n9500), .Q(
        WX877), .QN(n8784) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n9477), .CLK(n9500), .Q(
        WX879), .QN(n8729) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n9477), .CLK(n9500), .Q(
        WX881), .QN(n8742) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n9476), .CLK(n9501), .Q(
        WX883), .QN(n8751) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n9476), .CLK(n9501), .Q(
        WX885), .QN(n8782) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n9476), .CLK(n9501), .Q(
        WX887), .QN(n8769) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n9475), .CLK(n9502), .Q(
        WX889), .QN(n8754) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n9475), .CLK(n9502), .Q(
        WX891), .QN(n8757) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n9475), .CLK(n9502), .Q(
        WX893), .QN(n8698) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n9474), .CLK(n9503), .Q(
        WX895) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n9474), .CLK(n9503), .Q(
        WX897), .QN(n8713) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n9474), .CLK(n9503), .Q(
        WX899), .QN(n8788) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n9345), .CLK(n9635), .Q(
        CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n9345), .CLK(n9635), 
        .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n9345), .CLK(n9635), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n9345), .CLK(n9635), 
        .Q(CRC_OUT_9_3) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n9345), .CLK(n9635), 
        .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n9345), .CLK(n9635), 
        .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n9345), .CLK(n9635), 
        .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n9345), .CLK(n9635), 
        .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n9344), .CLK(n9636), 
        .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n9344), .CLK(n9636), 
        .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n9344), .CLK(n9636), 
        .Q(CRC_OUT_9_10) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n9344), .CLK(n9636), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n9344), .CLK(n9636), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n9344), .CLK(n9636), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n9344), .CLK(n9636), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n9344), .CLK(n9636), .Q(CRC_OUT_9_15) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n9344), .CLK(n9636), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n9344), .CLK(n9636), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n9344), .CLK(n9636), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n9344), .CLK(n9636), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n9471), .CLK(n9506), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n9471), .CLK(n9506), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n9471), .CLK(n9506), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n9471), .CLK(n9506), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n9471), .CLK(n9506), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n9471), .CLK(n9506), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n9471), .CLK(n9506), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n9471), .CLK(n9506), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n9339), .CLK(n9507), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n9343), .CLK(n9507), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(test_se), .CLK(
        n9507), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n9342), .CLK(n9507), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n250), .SI(CRC_OUT_9_31), .SE(n9341), .CLK(n9507), 
        .Q(WX1778) );
  SDFFX1 DFF_193_Q_reg ( .D(n251), .SI(WX1778), .SE(n9469), .CLK(n9509), .Q(
        n8702), .QN(n9030) );
  SDFFX1 DFF_194_Q_reg ( .D(n252), .SI(n8702), .SE(n9469), .CLK(n9509), .Q(
        n8701), .QN(n9029) );
  SDFFX1 DFF_195_Q_reg ( .D(n253), .SI(n8701), .SE(n9469), .CLK(n9509), .Q(
        n8700), .QN(n9028) );
  SDFFX1 DFF_196_Q_reg ( .D(n254), .SI(n8700), .SE(n9469), .CLK(n9509), .Q(
        n8699), .QN(n9027) );
  SDFFX1 DFF_197_Q_reg ( .D(n255), .SI(n8699), .SE(n9469), .CLK(n9509), .Q(
        test_so11), .QN(n9073) );
  SDFFX1 DFF_198_Q_reg ( .D(n256), .SI(test_si12), .SE(n9469), .CLK(n9509), 
        .Q(n8696), .QN(n9026) );
  SDFFX1 DFF_199_Q_reg ( .D(n257), .SI(n8696), .SE(n9469), .CLK(n9509), .Q(
        n8695), .QN(n9025) );
  SDFFX1 DFF_200_Q_reg ( .D(n258), .SI(n8695), .SE(n9469), .CLK(n9509), .Q(
        n8694), .QN(n9024) );
  SDFFX1 DFF_201_Q_reg ( .D(n259), .SI(n8694), .SE(n9469), .CLK(n9509), .Q(
        n8693), .QN(n9023) );
  SDFFX1 DFF_202_Q_reg ( .D(n260), .SI(n8693), .SE(n9469), .CLK(n9509), .Q(
        n8692), .QN(n9022) );
  SDFFX1 DFF_203_Q_reg ( .D(n261), .SI(n8692), .SE(n9469), .CLK(n9509), .Q(
        n8691), .QN(n9021) );
  SDFFX1 DFF_204_Q_reg ( .D(n262), .SI(n8691), .SE(n9469), .CLK(n9509), .Q(
        n8690), .QN(n9020) );
  SDFFX1 DFF_205_Q_reg ( .D(n263), .SI(n8690), .SE(n9470), .CLK(n9508), .Q(
        n8689), .QN(n9019) );
  SDFFX1 DFF_206_Q_reg ( .D(n264), .SI(n8689), .SE(n9470), .CLK(n9508), .Q(
        n8688), .QN(n9018) );
  SDFFX1 DFF_207_Q_reg ( .D(n265), .SI(n8688), .SE(n9470), .CLK(n9508), .Q(
        n8687), .QN(n9017) );
  SDFFX1 DFF_208_Q_reg ( .D(n266), .SI(n8687), .SE(n9470), .CLK(n9508), .Q(
        n8686), .QN(n9016) );
  SDFFX1 DFF_209_Q_reg ( .D(n267), .SI(n8686), .SE(n9470), .CLK(n9508), .Q(
        n8685), .QN(n9015) );
  SDFFX1 DFF_210_Q_reg ( .D(n268), .SI(n8685), .SE(n9470), .CLK(n9508), .Q(
        n8684), .QN(n9014) );
  SDFFX1 DFF_211_Q_reg ( .D(n269), .SI(n8684), .SE(n9470), .CLK(n9508), .Q(
        n8683), .QN(n9013) );
  SDFFX1 DFF_212_Q_reg ( .D(n270), .SI(n8683), .SE(n9470), .CLK(n9508), .Q(
        n8682), .QN(n9012) );
  SDFFX1 DFF_213_Q_reg ( .D(n271), .SI(n8682), .SE(n9470), .CLK(n9508), .Q(
        n8681), .QN(n9011) );
  SDFFX1 DFF_214_Q_reg ( .D(n272), .SI(n8681), .SE(n9470), .CLK(n9508), .Q(
        n8680), .QN(n9010) );
  SDFFX1 DFF_215_Q_reg ( .D(n273), .SI(n8680), .SE(n9470), .CLK(n9508), .Q(
        test_so12), .QN(n9072) );
  SDFFX1 DFF_216_Q_reg ( .D(n274), .SI(test_si13), .SE(n9470), .CLK(n9508), 
        .Q(n8677), .QN(n9009) );
  SDFFX1 DFF_217_Q_reg ( .D(n275), .SI(n8677), .SE(n9342), .CLK(n9507), .Q(
        n8676), .QN(n9008) );
  SDFFX1 DFF_218_Q_reg ( .D(n276), .SI(n8676), .SE(test_se), .CLK(n9507), .Q(
        n8675), .QN(n9007) );
  SDFFX1 DFF_219_Q_reg ( .D(n277), .SI(n8675), .SE(n9343), .CLK(n9507), .Q(
        n8674), .QN(n9006) );
  SDFFX1 DFF_220_Q_reg ( .D(n278), .SI(n8674), .SE(n9339), .CLK(n9507), .Q(
        n8673), .QN(n9005) );
  SDFFX1 DFF_221_Q_reg ( .D(n279), .SI(n8673), .SE(n9340), .CLK(n9507), .Q(
        n8672), .QN(n9004) );
  SDFFX1 DFF_222_Q_reg ( .D(n280), .SI(n8672), .SE(n9337), .CLK(n9507), .Q(
        n8671), .QN(n9003) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n9338), .CLK(n9507), .Q(
        n8670), .QN(n9002) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n9468), .CLK(n9510), .Q(
        n8669), .QN(n16027) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n9468), .CLK(n9510), .Q(
        n8668), .QN(n16028) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n9468), .CLK(n9510), .Q(
        n8667), .QN(n16029) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n9468), .CLK(n9510), .Q(
        n8666), .QN(n16030) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n9467), .CLK(n9511), .Q(
        n8665), .QN(n16031) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n9467), .CLK(n9511), .Q(
        n8664), .QN(n16032) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n9467), .CLK(n9511), .Q(
        n8663), .QN(n16033) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n9466), .CLK(n9512), .Q(
        n8662), .QN(n16034) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n9466), .CLK(n9512), .Q(
        n8661), .QN(n16035) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n9345), .CLK(n9635), .Q(
        test_so13), .QN(n8824) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n9465), .CLK(n9513), 
        .Q(n8658), .QN(n16036) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n9465), .CLK(n9513), .Q(
        n8657), .QN(n16037) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n9465), .CLK(n9513), .Q(
        n8656), .QN(n16038) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n9465), .CLK(n9513), .Q(
        n8655), .QN(n16039) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n9464), .CLK(n9514), .Q(
        n8654), .QN(n16040) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n9464), .CLK(n9514), .Q(
        n8653), .QN(n16041) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n9464), .CLK(n9514), .Q(
        WX1970), .QN(n8093) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n9463), .CLK(n9515), .Q(
        WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n9463), .CLK(n9515), .Q(
        WX1974), .QN(n8090) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n9463), .CLK(n9515), .Q(
        WX1976), .QN(n8088) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n9462), .CLK(n9516), .Q(
        WX1978), .QN(n8086) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n9462), .CLK(n9516), .Q(
        WX1980), .QN(n8084) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n9462), .CLK(n9516), .Q(
        WX1982), .QN(n8082) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n9461), .CLK(n9517), .Q(
        WX1984), .QN(n8080) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n9461), .CLK(n9517), .Q(
        WX1986), .QN(n8078) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n9461), .CLK(n9517), .Q(
        WX1988), .QN(n8076) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n9340), .CLK(n9518), .Q(
        WX1990), .QN(n8074) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n9342), .CLK(n9518), .Q(
        test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n9460), .CLK(n9519), 
        .Q(WX1994), .QN(n8071) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n9460), .CLK(n9519), .Q(
        WX1996), .QN(n8069) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n9460), .CLK(n9519), .Q(
        WX1998), .QN(n8067) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n9460), .CLK(n9519), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n9468), .CLK(n9510), .Q(
        WX2002), .QN(n7625) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n9468), .CLK(n9510), .Q(
        WX2004), .QN(n7851) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n9468), .CLK(n9510), .Q(
        WX2006), .QN(n7849) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n9468), .CLK(n9510), .Q(
        WX2008), .QN(n7847) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n9467), .CLK(n9511), .Q(
        WX2010), .QN(n7845) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n9467), .CLK(n9511), .Q(
        WX2012), .QN(n7843) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n9467), .CLK(n9511), .Q(
        WX2014), .QN(n7841) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n9466), .CLK(n9512), .Q(
        WX2016), .QN(n7839) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n9466), .CLK(n9512), .Q(
        WX2018), .QN(n7837) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n9466), .CLK(n9512), .Q(
        WX2020), .QN(n7835) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n9466), .CLK(n9512), .Q(
        WX2022), .QN(n7833) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n9465), .CLK(n9513), .Q(
        WX2024), .QN(n7831) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n9465), .CLK(n9513), .Q(
        WX2026), .QN(n7829) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n9464), .CLK(n9514), .Q(
        test_so15), .QN(n8814) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n9464), .CLK(n9514), 
        .Q(WX2030), .QN(n7826) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n9464), .CLK(n9514), .Q(
        WX2032), .QN(n7824) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n9463), .CLK(n9515), .Q(
        WX2034) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n9463), .CLK(n9515), .Q(
        WX2036), .QN(n3783) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n9463), .CLK(n9515), .Q(
        WX2038) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n9462), .CLK(n9516), .Q(
        WX2040) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n9462), .CLK(n9516), .Q(
        WX2042) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n9462), .CLK(n9516), .Q(
        WX2044), .QN(n3775) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n9461), .CLK(n9517), .Q(
        WX2046) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n9461), .CLK(n9517), .Q(
        WX2048) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n9461), .CLK(n9517), .Q(
        WX2050) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n9341), .CLK(n9518), .Q(
        WX2052) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n9339), .CLK(n9518), .Q(
        WX2054) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n9341), .CLK(n9518), .Q(
        WX2056), .QN(n3763) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n9340), .CLK(n9518), .Q(
        WX2058) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n9460), .CLK(n9519), .Q(
        WX2060) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n9460), .CLK(n9519), .Q(
        WX2062) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n9459), .CLK(n9520), .Q(
        test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n9468), .CLK(n9510), 
        .Q(WX2066), .QN(n7626) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n9468), .CLK(n9510), .Q(
        WX2068), .QN(n7852) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n9468), .CLK(n9510), .Q(
        WX2070), .QN(n7850) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n9468), .CLK(n9510), .Q(
        WX2072), .QN(n7848) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n9467), .CLK(n9511), .Q(
        WX2074), .QN(n7846) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n9467), .CLK(n9511), .Q(
        WX2076), .QN(n7844) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n9467), .CLK(n9511), .Q(
        WX2078), .QN(n7842) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n9466), .CLK(n9512), .Q(
        WX2080), .QN(n7840) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n9466), .CLK(n9512), .Q(
        WX2082), .QN(n7838) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n9466), .CLK(n9512), .Q(
        WX2084), .QN(n7836) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n9465), .CLK(n9513), .Q(
        WX2086), .QN(n7834) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n9465), .CLK(n9513), .Q(
        WX2088), .QN(n7832) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n9465), .CLK(n9513), .Q(
        WX2090), .QN(n7830) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n9464), .CLK(n9514), .Q(
        WX2092), .QN(n7828) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n9464), .CLK(n9514), .Q(
        WX2094), .QN(n7827) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n9464), .CLK(n9514), .Q(
        WX2096), .QN(n7825) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n9463), .CLK(n9515), .Q(
        WX2098), .QN(n8094) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n9463), .CLK(n9515), .Q(
        test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n9463), .CLK(n9515), 
        .Q(WX2102), .QN(n8091) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n9462), .CLK(n9516), .Q(
        WX2104), .QN(n8089) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n9462), .CLK(n9516), .Q(
        WX2106), .QN(n8087) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n9462), .CLK(n9516), .Q(
        WX2108), .QN(n8085) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n9461), .CLK(n9517), .Q(
        WX2110), .QN(n8083) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n9461), .CLK(n9517), .Q(
        WX2112), .QN(n8081) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n9461), .CLK(n9517), .Q(
        WX2114), .QN(n8079) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n9338), .CLK(n9518), .Q(
        WX2116), .QN(n8077) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n9343), .CLK(n9518), .Q(
        WX2118), .QN(n8075) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n9338), .CLK(n9518), .Q(
        WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n9460), .CLK(n9519), .Q(
        WX2122), .QN(n8072) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n9460), .CLK(n9519), .Q(
        WX2124), .QN(n8070) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n9460), .CLK(n9519), .Q(
        WX2126), .QN(n8068) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n9459), .CLK(n9520), .Q(
        WX2128), .QN(n8066) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n9459), .CLK(n9520), .Q(
        WX2130), .QN(n8557) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n9459), .CLK(n9520), .Q(
        WX2132), .QN(n8574) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n9459), .CLK(n9520), .Q(
        WX2134), .QN(n8575) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n9459), .CLK(n9520), .Q(
        test_so18), .QN(n8802) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n9467), .CLK(n9511), 
        .Q(WX2138), .QN(n8587) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n9467), .CLK(n9511), .Q(
        WX2140) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n9467), .CLK(n9511), .Q(
        WX2142), .QN(n8589) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n9466), .CLK(n9512), .Q(
        WX2144), .QN(n8590) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n9466), .CLK(n9512), .Q(
        WX2146), .QN(n8591) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n9466), .CLK(n9512), .Q(
        WX2148), .QN(n8592) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n9465), .CLK(n9513), .Q(
        WX2150), .QN(n8593) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n9465), .CLK(n9513), .Q(
        WX2152), .QN(n8594) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n9465), .CLK(n9513), .Q(
        WX2154), .QN(n8595) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n9464), .CLK(n9514), .Q(
        WX2156), .QN(n8596) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n9464), .CLK(n9514), .Q(
        WX2158), .QN(n8614) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n9464), .CLK(n9514), .Q(
        WX2160), .QN(n8122) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n9463), .CLK(n9515), .Q(
        WX2162), .QN(n8615) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n9463), .CLK(n9515), .Q(
        WX2164), .QN(n8633) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n9463), .CLK(n9515), .Q(
        WX2166), .QN(n8634) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n9462), .CLK(n9516), .Q(
        WX2168), .QN(n8645) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n9462), .CLK(n9516), .Q(
        WX2170), .QN(n8123) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n9462), .CLK(n9516), .Q(
        test_so19), .QN(n8792) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n9461), .CLK(n9517), 
        .Q(WX2174), .QN(n8646) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n9461), .CLK(n9517), .Q(
        WX2176) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n9461), .CLK(n9517), .Q(
        WX2178), .QN(n8648) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n9337), .CLK(n9518), .Q(
        WX2180), .QN(n8649) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(test_se), .CLK(n9518), 
        .Q(WX2182), .QN(n8650) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n9337), .CLK(n9518), .Q(
        WX2184), .QN(n8124) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n9460), .CLK(n9519), .Q(
        WX2186), .QN(n8651) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n9460), .CLK(n9519), .Q(
        WX2188), .QN(n8652) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n9460), .CLK(n9519), .Q(
        WX2190), .QN(n8659) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n9459), .CLK(n9520), .Q(
        WX2192), .QN(n8132) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n9348), .CLK(n9632), .Q(
        CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n9348), .CLK(n9632), 
        .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n9348), .CLK(n9632), 
        .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n9348), .CLK(n9632), 
        .Q(CRC_OUT_8_3) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n9347), .CLK(n9633), 
        .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n9347), .CLK(n9633), 
        .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n9347), .CLK(n9633), 
        .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n9347), .CLK(n9633), 
        .Q(test_so20) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n9347), .CLK(n9633), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n9347), .CLK(n9633), 
        .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n9347), .CLK(n9633), 
        .Q(CRC_OUT_8_10) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n9347), .CLK(n9633), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n9347), .CLK(n9633), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n9347), .CLK(n9633), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n9347), .CLK(n9633), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n9347), .CLK(n9633), .Q(CRC_OUT_8_15) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n9346), .CLK(n9634), .Q(test_so21) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n9346), .CLK(n9634), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n9346), .CLK(n9634), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n9345), .CLK(n9635), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n9345), .CLK(n9635), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n9345), .CLK(n9635), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n9459), .CLK(n9520), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n491), .SI(CRC_OUT_8_31), .SE(n9459), .CLK(n9520), 
        .Q(WX3071) );
  SDFFX1 DFF_385_Q_reg ( .D(n492), .SI(WX3071), .SE(n9456), .CLK(n9523), .Q(
        n8644), .QN(n9001) );
  SDFFX1 DFF_386_Q_reg ( .D(n493), .SI(n8644), .SE(n9456), .CLK(n9523), .Q(
        n8643), .QN(n9000) );
  SDFFX1 DFF_387_Q_reg ( .D(n494), .SI(n8643), .SE(n9456), .CLK(n9523), .Q(
        n8642), .QN(n8999) );
  SDFFX1 DFF_388_Q_reg ( .D(n495), .SI(n8642), .SE(n9456), .CLK(n9523), .Q(
        n8641), .QN(n8998) );
  SDFFX1 DFF_389_Q_reg ( .D(n496), .SI(n8641), .SE(n9457), .CLK(n9522), .Q(
        n8640), .QN(n8997) );
  SDFFX1 DFF_390_Q_reg ( .D(n497), .SI(n8640), .SE(n9457), .CLK(n9522), .Q(
        n8639), .QN(n8996) );
  SDFFX1 DFF_391_Q_reg ( .D(n498), .SI(n8639), .SE(n9457), .CLK(n9522), .Q(
        n8638), .QN(n8995) );
  SDFFX1 DFF_392_Q_reg ( .D(n499), .SI(n8638), .SE(n9457), .CLK(n9522), .Q(
        n8637), .QN(n8994) );
  SDFFX1 DFF_393_Q_reg ( .D(n500), .SI(n8637), .SE(n9457), .CLK(n9522), .Q(
        n8636), .QN(n8993) );
  SDFFX1 DFF_394_Q_reg ( .D(n501), .SI(n8636), .SE(n9457), .CLK(n9522), .Q(
        n8635), .QN(n8992) );
  SDFFX1 DFF_395_Q_reg ( .D(n502), .SI(n8635), .SE(n9457), .CLK(n9522), .Q(
        test_so22), .QN(n9071) );
  SDFFX1 DFF_396_Q_reg ( .D(n503), .SI(test_si23), .SE(n9457), .CLK(n9522), 
        .Q(n8632), .QN(n8991) );
  SDFFX1 DFF_397_Q_reg ( .D(n504), .SI(n8632), .SE(n9457), .CLK(n9522), .Q(
        n8631), .QN(n8990) );
  SDFFX1 DFF_398_Q_reg ( .D(n505), .SI(n8631), .SE(n9457), .CLK(n9522), .Q(
        n8630), .QN(n8989) );
  SDFFX1 DFF_399_Q_reg ( .D(n506), .SI(n8630), .SE(n9457), .CLK(n9522), .Q(
        n8629), .QN(n8988) );
  SDFFX1 DFF_400_Q_reg ( .D(n507), .SI(n8629), .SE(n9457), .CLK(n9522), .Q(
        n8628), .QN(n8987) );
  SDFFX1 DFF_401_Q_reg ( .D(n508), .SI(n8628), .SE(n9458), .CLK(n9521), .Q(
        n8627), .QN(n8986) );
  SDFFX1 DFF_402_Q_reg ( .D(n509), .SI(n8627), .SE(n9458), .CLK(n9521), .Q(
        n8626), .QN(n8985) );
  SDFFX1 DFF_403_Q_reg ( .D(n510), .SI(n8626), .SE(n9458), .CLK(n9521), .Q(
        n8625), .QN(n8984) );
  SDFFX1 DFF_404_Q_reg ( .D(n511), .SI(n8625), .SE(n9458), .CLK(n9521), .Q(
        n8624), .QN(n8983) );
  SDFFX1 DFF_405_Q_reg ( .D(n512), .SI(n8624), .SE(n9458), .CLK(n9521), .Q(
        n8623), .QN(n8982) );
  SDFFX1 DFF_406_Q_reg ( .D(n513), .SI(n8623), .SE(n9458), .CLK(n9521), .Q(
        n8622), .QN(n8981) );
  SDFFX1 DFF_407_Q_reg ( .D(n514), .SI(n8622), .SE(n9458), .CLK(n9521), .Q(
        n8621), .QN(n8980) );
  SDFFX1 DFF_408_Q_reg ( .D(n515), .SI(n8621), .SE(n9458), .CLK(n9521), .Q(
        n8620), .QN(n8979) );
  SDFFX1 DFF_409_Q_reg ( .D(n516), .SI(n8620), .SE(n9458), .CLK(n9521), .Q(
        n8619), .QN(n8978) );
  SDFFX1 DFF_410_Q_reg ( .D(n517), .SI(n8619), .SE(n9458), .CLK(n9521), .Q(
        n8618), .QN(n8977) );
  SDFFX1 DFF_411_Q_reg ( .D(n518), .SI(n8618), .SE(n9458), .CLK(n9521), .Q(
        n8617), .QN(n8976) );
  SDFFX1 DFF_412_Q_reg ( .D(n519), .SI(n8617), .SE(n9458), .CLK(n9521), .Q(
        n8616), .QN(n8975) );
  SDFFX1 DFF_413_Q_reg ( .D(n520), .SI(n8616), .SE(n9459), .CLK(n9520), .Q(
        test_so23), .QN(n9070) );
  SDFFX1 DFF_414_Q_reg ( .D(n521), .SI(test_si24), .SE(n9459), .CLK(n9520), 
        .Q(n8613), .QN(n8974) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n9459), .CLK(n9520), .Q(
        n8612), .QN(n8973) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n9456), .CLK(n9523), .Q(
        n8611), .QN(n16042) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n9456), .CLK(n9523), .Q(
        n8610), .QN(n16043) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n9456), .CLK(n9523), .Q(
        n8609), .QN(n16044) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n9456), .CLK(n9523), .Q(
        n8608), .QN(n16045) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n9455), .CLK(n9524), .Q(
        n8607), .QN(n16046) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n9455), .CLK(n9524), .Q(
        n8606), .QN(n16047) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n9455), .CLK(n9524), .Q(
        n8605), .QN(n16048) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n9455), .CLK(n9524), .Q(
        n8604), .QN(n16049) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n9455), .CLK(n9524), .Q(
        n8603), .QN(n16050) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n9454), .CLK(n9525), .Q(
        n8602), .QN(n16051) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n9454), .CLK(n9525), .Q(
        n8601), .QN(n16052) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n9453), .CLK(n9526), .Q(
        n8600), .QN(n16053) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n9453), .CLK(n9526), .Q(
        n8599), .QN(n16054) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n9453), .CLK(n9526), .Q(
        n8598), .QN(n16055) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n9453), .CLK(n9526), .Q(
        n8597), .QN(n16056) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n9348), .CLK(n9632), .Q(
        test_so24), .QN(n8823) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n9340), .CLK(n9527), 
        .Q(WX3263), .QN(n8063) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n9339), .CLK(n9527), .Q(
        WX3265), .QN(n8061) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n9452), .CLK(n9528), .Q(
        WX3267), .QN(n8059) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n9452), .CLK(n9528), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n9452), .CLK(n9528), .Q(
        WX3271), .QN(n8055) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n9451), .CLK(n9529), .Q(
        WX3273), .QN(n8053) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n9451), .CLK(n9529), .Q(
        WX3275), .QN(n8051) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n9451), .CLK(n9529), .Q(
        WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n9450), .CLK(n9530), .Q(
        WX3279), .QN(n8048) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n9450), .CLK(n9530), .Q(
        WX3281), .QN(n8046) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n9450), .CLK(n9530), .Q(
        WX3283), .QN(n8044) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n9449), .CLK(n9531), .Q(
        WX3285), .QN(n8042) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n9449), .CLK(n9531), .Q(
        WX3287), .QN(n8040) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n9449), .CLK(n9531), .Q(
        WX3289), .QN(n8038) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n9448), .CLK(n9532), .Q(
        WX3291), .QN(n8036) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n9448), .CLK(n9532), .Q(
        WX3293), .QN(n8034) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n9456), .CLK(n9523), .Q(
        WX3295), .QN(n7623) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n9456), .CLK(n9523), .Q(
        test_so25), .QN(n8816) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n9456), .CLK(n9523), 
        .Q(WX3299), .QN(n7821) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n9456), .CLK(n9523), .Q(
        WX3301), .QN(n7819) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n9455), .CLK(n9524), .Q(
        WX3303), .QN(n7817) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n9455), .CLK(n9524), .Q(
        WX3305), .QN(n7816) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n9455), .CLK(n9524), .Q(
        WX3307), .QN(n7814) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n9455), .CLK(n9524), .Q(
        WX3309), .QN(n7812) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n9455), .CLK(n9524), .Q(
        WX3311), .QN(n7810) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n9454), .CLK(n9525), .Q(
        WX3313), .QN(n7808) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n9454), .CLK(n9525), .Q(
        WX3315), .QN(n7806) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n9454), .CLK(n9525), .Q(
        WX3317), .QN(n7804) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n9453), .CLK(n9526), .Q(
        WX3319), .QN(n7802) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n9453), .CLK(n9526), .Q(
        WX3321), .QN(n7800) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n9453), .CLK(n9526), .Q(
        WX3323), .QN(n7798) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n9343), .CLK(n9527), .Q(
        WX3325), .QN(n7796) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n9341), .CLK(n9527), .Q(
        WX3327) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n9343), .CLK(n9527), .Q(
        WX3329) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n9452), .CLK(n9528), .Q(
        WX3331) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n9452), .CLK(n9528), .Q(
        test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n9452), .CLK(n9528), 
        .Q(WX3335) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n9451), .CLK(n9529), .Q(
        WX3337) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n9451), .CLK(n9529), .Q(
        WX3339) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n9451), .CLK(n9529), .Q(
        WX3341), .QN(n3739) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n9450), .CLK(n9530), .Q(
        WX3343) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n9450), .CLK(n9530), .Q(
        WX3345), .QN(n3735) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n9450), .CLK(n9530), .Q(
        WX3347) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n9449), .CLK(n9531), .Q(
        WX3349) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n9449), .CLK(n9531), .Q(
        WX3351) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n9449), .CLK(n9531), .Q(
        WX3353) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n9448), .CLK(n9532), .Q(
        WX3355) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n9448), .CLK(n9532), .Q(
        WX3357) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n9448), .CLK(n9532), .Q(
        WX3359), .QN(n7624) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n9448), .CLK(n9532), .Q(
        WX3361), .QN(n7823) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n9447), .CLK(n9533), .Q(
        WX3363), .QN(n7822) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n9447), .CLK(n9533), .Q(
        WX3365), .QN(n7820) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n9447), .CLK(n9533), .Q(
        WX3367), .QN(n7818) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n9447), .CLK(n9533), .Q(
        test_so27), .QN(n8815) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n9455), .CLK(n9524), 
        .Q(WX3371), .QN(n7815) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n9455), .CLK(n9524), .Q(
        WX3373), .QN(n7813) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n9454), .CLK(n9525), .Q(
        WX3375), .QN(n7811) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n9454), .CLK(n9525), .Q(
        WX3377), .QN(n7809) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n9454), .CLK(n9525), .Q(
        WX3379), .QN(n7807) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n9454), .CLK(n9525), .Q(
        WX3381), .QN(n7805) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n9453), .CLK(n9526), .Q(
        WX3383), .QN(n7803) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n9453), .CLK(n9526), .Q(
        WX3385), .QN(n7801) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n9453), .CLK(n9526), .Q(
        WX3387), .QN(n7799) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(test_se), .CLK(n9527), 
        .Q(WX3389), .QN(n7797) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n9338), .CLK(n9527), .Q(
        WX3391), .QN(n8064) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(test_se), .CLK(n9527), 
        .Q(WX3393), .QN(n8062) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n9452), .CLK(n9528), .Q(
        WX3395), .QN(n8060) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n9452), .CLK(n9528), .Q(
        WX3397), .QN(n8058) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n9452), .CLK(n9528), .Q(
        WX3399), .QN(n8056) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n9451), .CLK(n9529), .Q(
        WX3401), .QN(n8054) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n9451), .CLK(n9529), .Q(
        WX3403), .QN(n8052) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n9451), .CLK(n9529), .Q(
        test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n9450), .CLK(n9530), 
        .Q(WX3407), .QN(n8049) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n9450), .CLK(n9530), .Q(
        WX3409), .QN(n8047) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n9450), .CLK(n9530), .Q(
        WX3411), .QN(n8045) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n9449), .CLK(n9531), .Q(
        WX3413), .QN(n8043) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n9449), .CLK(n9531), .Q(
        WX3415), .QN(n8041) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n9449), .CLK(n9531), .Q(
        WX3417), .QN(n8039) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n9448), .CLK(n9532), .Q(
        WX3419), .QN(n8037) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n9448), .CLK(n9532), .Q(
        WX3421), .QN(n8035) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n9448), .CLK(n9532), .Q(
        WX3423), .QN(n8469) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n9448), .CLK(n9532), .Q(
        WX3425), .QN(n8471) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n9447), .CLK(n9533), .Q(
        WX3427), .QN(n8472) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n9447), .CLK(n9533), .Q(
        WX3429) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n9447), .CLK(n9533), .Q(
        WX3431), .QN(n8474) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n9447), .CLK(n9533), .Q(
        WX3433), .QN(n8475) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n9447), .CLK(n9533), .Q(
        WX3435), .QN(n8476) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n9447), .CLK(n9533), .Q(
        WX3437), .QN(n8477) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n9447), .CLK(n9533), .Q(
        test_so29), .QN(n8801) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n9454), .CLK(n9525), 
        .Q(WX3441), .QN(n8478) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n9454), .CLK(n9525), .Q(
        WX3443), .QN(n8485) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n9454), .CLK(n9525), .Q(
        WX3445), .QN(n8486) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n9453), .CLK(n9526), .Q(
        WX3447), .QN(n8503) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n9453), .CLK(n9526), .Q(
        WX3449), .QN(n8504) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n9339), .CLK(n9527), .Q(
        WX3451), .QN(n8521) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n9342), .CLK(n9527), .Q(
        WX3453), .QN(n8119) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n9337), .CLK(n9527), .Q(
        WX3455), .QN(n8522) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n9342), .CLK(n9527), .Q(
        WX3457), .QN(n8529) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n9452), .CLK(n9528), .Q(
        WX3459), .QN(n8530) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n9452), .CLK(n9528), .Q(
        WX3461), .QN(n8531) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n9452), .CLK(n9528), .Q(
        WX3463) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n9451), .CLK(n9529), .Q(
        WX3465), .QN(n8532) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n9451), .CLK(n9529), .Q(
        WX3467), .QN(n8533) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n9451), .CLK(n9529), .Q(
        WX3469), .QN(n8534) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n9450), .CLK(n9530), .Q(
        WX3471), .QN(n8535) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n9450), .CLK(n9530), .Q(
        test_so30), .QN(n8791) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n9450), .CLK(n9530), 
        .Q(WX3475), .QN(n8536) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n9449), .CLK(n9531), .Q(
        WX3477), .QN(n8121) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n9449), .CLK(n9531), .Q(
        WX3479), .QN(n8538) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n9449), .CLK(n9531), .Q(
        WX3481), .QN(n8539) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n9448), .CLK(n9532), .Q(
        WX3483), .QN(n8556) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n9448), .CLK(n9532), .Q(
        WX3485), .QN(n8131) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n9350), .CLK(n9630), .Q(
        CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n9350), .CLK(n9630), 
        .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n9350), .CLK(n9630), 
        .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n9350), .CLK(n9630), 
        .Q(CRC_OUT_7_3) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n9350), .CLK(n9630), 
        .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n9350), .CLK(n9630), 
        .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n9350), .CLK(n9630), 
        .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n9349), .CLK(n9631), 
        .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n9349), .CLK(n9631), 
        .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n9349), .CLK(n9631), 
        .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n9349), .CLK(n9631), 
        .Q(test_so31) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n9349), .CLK(n9631), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n9349), .CLK(n9631), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n9349), .CLK(n9631), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n9349), .CLK(n9631), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n9349), .CLK(n9631), .Q(CRC_OUT_7_15) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n9349), .CLK(n9631), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n9349), .CLK(n9631), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n9349), .CLK(n9631), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n9348), .CLK(n9632), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n9348), .CLK(n9632), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n9348), .CLK(n9632), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n9348), .CLK(n9632), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n9348), .CLK(n9632), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n9348), .CLK(n9632), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n9348), .CLK(n9632), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n9447), .CLK(n9533), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n9446), .CLK(n9534), .Q(test_so32) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n9446), .CLK(n9534), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n9446), .CLK(n9534), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n9446), .CLK(n9534), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n9446), .CLK(n9534), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n732), .SI(CRC_OUT_7_31), .SE(n9446), .CLK(n9534), 
        .Q(WX4364) );
  SDFFX1 DFF_577_Q_reg ( .D(n733), .SI(WX4364), .SE(n9443), .CLK(n9537), .Q(
        n8586), .QN(n8972) );
  SDFFX1 DFF_578_Q_reg ( .D(n734), .SI(n8586), .SE(n9444), .CLK(n9536), .Q(
        n8585), .QN(n8971) );
  SDFFX1 DFF_579_Q_reg ( .D(n735), .SI(n8585), .SE(n9444), .CLK(n9536), .Q(
        n8584), .QN(n8970) );
  SDFFX1 DFF_580_Q_reg ( .D(n736), .SI(n8584), .SE(n9444), .CLK(n9536), .Q(
        n8583), .QN(n8969) );
  SDFFX1 DFF_581_Q_reg ( .D(n737), .SI(n8583), .SE(n9444), .CLK(n9536), .Q(
        n8582), .QN(n8968) );
  SDFFX1 DFF_582_Q_reg ( .D(n738), .SI(n8582), .SE(n9444), .CLK(n9536), .Q(
        n8581), .QN(n8967) );
  SDFFX1 DFF_583_Q_reg ( .D(n739), .SI(n8581), .SE(n9444), .CLK(n9536), .Q(
        n8580), .QN(n8966) );
  SDFFX1 DFF_584_Q_reg ( .D(n740), .SI(n8580), .SE(n9444), .CLK(n9536), .Q(
        n8579), .QN(n8965) );
  SDFFX1 DFF_585_Q_reg ( .D(n741), .SI(n8579), .SE(n9444), .CLK(n9536), .Q(
        n8578), .QN(n8964) );
  SDFFX1 DFF_586_Q_reg ( .D(n742), .SI(n8578), .SE(n9444), .CLK(n9536), .Q(
        n8577), .QN(n8963) );
  SDFFX1 DFF_587_Q_reg ( .D(n743), .SI(n8577), .SE(n9444), .CLK(n9536), .Q(
        n8576), .QN(n8962) );
  SDFFX1 DFF_588_Q_reg ( .D(n744), .SI(n8576), .SE(n9444), .CLK(n9536), .Q(
        test_so33), .QN(n9069) );
  SDFFX1 DFF_589_Q_reg ( .D(n745), .SI(test_si34), .SE(n9444), .CLK(n9536), 
        .Q(n8573), .QN(n8961) );
  SDFFX1 DFF_590_Q_reg ( .D(n746), .SI(n8573), .SE(n9445), .CLK(n9535), .Q(
        n8572), .QN(n8960) );
  SDFFX1 DFF_591_Q_reg ( .D(n747), .SI(n8572), .SE(n9445), .CLK(n9535), .Q(
        n8571), .QN(n8959) );
  SDFFX1 DFF_592_Q_reg ( .D(n748), .SI(n8571), .SE(n9445), .CLK(n9535), .Q(
        n8570), .QN(n8958) );
  SDFFX1 DFF_593_Q_reg ( .D(n749), .SI(n8570), .SE(n9445), .CLK(n9535), .Q(
        n8569), .QN(n8957) );
  SDFFX1 DFF_594_Q_reg ( .D(n750), .SI(n8569), .SE(n9445), .CLK(n9535), .Q(
        n8568), .QN(n8956) );
  SDFFX1 DFF_595_Q_reg ( .D(n751), .SI(n8568), .SE(n9445), .CLK(n9535), .Q(
        n8567), .QN(n8955) );
  SDFFX1 DFF_596_Q_reg ( .D(n752), .SI(n8567), .SE(n9445), .CLK(n9535), .Q(
        n8566), .QN(n8954) );
  SDFFX1 DFF_597_Q_reg ( .D(n753), .SI(n8566), .SE(n9445), .CLK(n9535), .Q(
        n8565), .QN(n8953) );
  SDFFX1 DFF_598_Q_reg ( .D(n754), .SI(n8565), .SE(n9445), .CLK(n9535), .Q(
        n8564), .QN(n8952) );
  SDFFX1 DFF_599_Q_reg ( .D(n755), .SI(n8564), .SE(n9445), .CLK(n9535), .Q(
        n8563), .QN(n8951) );
  SDFFX1 DFF_600_Q_reg ( .D(n756), .SI(n8563), .SE(n9445), .CLK(n9535), .Q(
        n8562), .QN(n8950) );
  SDFFX1 DFF_601_Q_reg ( .D(n757), .SI(n8562), .SE(n9445), .CLK(n9535), .Q(
        n8561), .QN(n8949) );
  SDFFX1 DFF_602_Q_reg ( .D(n758), .SI(n8561), .SE(n9446), .CLK(n9534), .Q(
        n8560), .QN(n8948) );
  SDFFX1 DFF_603_Q_reg ( .D(n759), .SI(n8560), .SE(n9446), .CLK(n9534), .Q(
        n8559), .QN(n8947) );
  SDFFX1 DFF_604_Q_reg ( .D(n760), .SI(n8559), .SE(n9446), .CLK(n9534), .Q(
        n8558), .QN(n8946) );
  SDFFX1 DFF_605_Q_reg ( .D(n761), .SI(n8558), .SE(n9446), .CLK(n9534), .Q(
        test_so34), .QN(n9068) );
  SDFFX1 DFF_606_Q_reg ( .D(n762), .SI(test_si35), .SE(n9446), .CLK(n9534), 
        .Q(n8555), .QN(n8945) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n9446), .CLK(n9534), .Q(
        n8554), .QN(n8944) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n9443), .CLK(n9537), .Q(
        n8553), .QN(n16057) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n9443), .CLK(n9537), .Q(
        n8552), .QN(n16058) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n9443), .CLK(n9537), .Q(
        n8551), .QN(n16059) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n9443), .CLK(n9537), .Q(
        n8550), .QN(n16060) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n9443), .CLK(n9537), .Q(
        n8549), .QN(n16061) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n9442), .CLK(n9538), .Q(
        n8548), .QN(n16062) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n9442), .CLK(n9538), .Q(
        n8547), .QN(n16063) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n9441), .CLK(n9539), .Q(
        n8546), .QN(n16064) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n9441), .CLK(n9539), .Q(
        n8545), .QN(n16065) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n9441), .CLK(n9539), .Q(
        n8544), .QN(n16066) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n9441), .CLK(n9539), .Q(
        n8543), .QN(n16067) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n9440), .CLK(n9540), .Q(
        n8542), .QN(n16068) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n9440), .CLK(n9540), .Q(
        n8541), .QN(n16069) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n9439), .CLK(n9541), .Q(
        n8540), .QN(n16070) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n9439), .CLK(n9541), .Q(
        test_so35), .QN(n8822) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n9439), .CLK(n9541), 
        .Q(n8537), .QN(n16071) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n9439), .CLK(n9541), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n9438), .CLK(n9542), .Q(
        WX4558), .QN(n8030) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n9438), .CLK(n9542), .Q(
        WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n9438), .CLK(n9542), .Q(
        WX4562), .QN(n8027) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n9437), .CLK(n9543), .Q(
        WX4564), .QN(n8025) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n9437), .CLK(n9543), .Q(
        WX4566), .QN(n8023) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n9437), .CLK(n9543), .Q(
        WX4568), .QN(n8021) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n9436), .CLK(n9544), .Q(
        WX4570), .QN(n8019) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n9436), .CLK(n9544), .Q(
        WX4572), .QN(n8017) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n9436), .CLK(n9544), .Q(
        WX4574), .QN(n8015) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n9435), .CLK(n9545), .Q(
        WX4576), .QN(n8013) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n9435), .CLK(n9545), .Q(
        WX4578), .QN(n8011) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n9435), .CLK(n9545), .Q(
        WX4580), .QN(n8009) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n9434), .CLK(n9546), .Q(
        WX4582), .QN(n8007) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n9434), .CLK(n9546), .Q(
        WX4584), .QN(n8005) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n9434), .CLK(n9546), .Q(
        test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n9443), .CLK(n9537), 
        .Q(WX4588), .QN(n7621) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n9443), .CLK(n9537), .Q(
        WX4590), .QN(n7795) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n9443), .CLK(n9537), .Q(
        WX4592), .QN(n7793) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n9443), .CLK(n9537), .Q(
        WX4594), .QN(n7791) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n9442), .CLK(n9538), .Q(
        WX4596), .QN(n7789) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n9442), .CLK(n9538), .Q(
        WX4598), .QN(n7787) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n9442), .CLK(n9538), .Q(
        WX4600), .QN(n7785) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n9442), .CLK(n9538), .Q(
        WX4602), .QN(n7783) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n9441), .CLK(n9539), .Q(
        WX4604), .QN(n7781) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n9441), .CLK(n9539), .Q(
        WX4606), .QN(n7779) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n9440), .CLK(n9540), .Q(
        WX4608), .QN(n7777) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n9440), .CLK(n9540), .Q(
        WX4610), .QN(n7775) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n9440), .CLK(n9540), .Q(
        WX4612), .QN(n7773) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n9440), .CLK(n9540), .Q(
        WX4614), .QN(n7771) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n9439), .CLK(n9541), .Q(
        WX4616), .QN(n7769) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n9439), .CLK(n9541), .Q(
        WX4618), .QN(n7767) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n9438), .CLK(n9542), .Q(
        test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n9438), .CLK(n9542), 
        .Q(WX4622) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n9438), .CLK(n9542), .Q(
        WX4624), .QN(n3717) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n9437), .CLK(n9543), .Q(
        WX4626) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n9437), .CLK(n9543), .Q(
        WX4628), .QN(n3713) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n9437), .CLK(n9543), .Q(
        WX4630) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n9436), .CLK(n9544), .Q(
        WX4632) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n9436), .CLK(n9544), .Q(
        WX4634) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n9436), .CLK(n9544), .Q(
        WX4636) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n9435), .CLK(n9545), .Q(
        WX4638) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n9435), .CLK(n9545), .Q(
        WX4640) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n9435), .CLK(n9545), .Q(
        WX4642) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n9434), .CLK(n9546), .Q(
        WX4644) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n9434), .CLK(n9546), .Q(
        WX4646) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n9434), .CLK(n9546), .Q(
        WX4648) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n9433), .CLK(n9547), .Q(
        WX4650), .QN(n3691) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n9433), .CLK(n9547), .Q(
        WX4652), .QN(n7622) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n9433), .CLK(n9547), .Q(
        test_so38), .QN(n8813) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n9443), .CLK(n9537), 
        .Q(WX4656), .QN(n7794) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n9443), .CLK(n9537), .Q(
        WX4658), .QN(n7792) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n9442), .CLK(n9538), .Q(
        WX4660), .QN(n7790) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n9442), .CLK(n9538), .Q(
        WX4662), .QN(n7788) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n9442), .CLK(n9538), .Q(
        WX4664), .QN(n7786) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n9441), .CLK(n9539), .Q(
        WX4666), .QN(n7784) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n9441), .CLK(n9539), .Q(
        WX4668), .QN(n7782) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n9441), .CLK(n9539), .Q(
        WX4670), .QN(n7780) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n9440), .CLK(n9540), .Q(
        WX4672), .QN(n7778) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n9440), .CLK(n9540), .Q(
        WX4674), .QN(n7776) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n9440), .CLK(n9540), .Q(
        WX4676), .QN(n7774) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n9439), .CLK(n9541), .Q(
        WX4678), .QN(n7772) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n9439), .CLK(n9541), .Q(
        WX4680), .QN(n7770) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n9439), .CLK(n9541), .Q(
        WX4682), .QN(n7768) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n9438), .CLK(n9542), .Q(
        WX4684), .QN(n8033) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n9438), .CLK(n9542), .Q(
        WX4686), .QN(n8031) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n9438), .CLK(n9542), .Q(
        test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n9437), .CLK(n9543), 
        .Q(WX4690), .QN(n8028) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n9437), .CLK(n9543), .Q(
        WX4692), .QN(n8026) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n9437), .CLK(n9543), .Q(
        WX4694), .QN(n8024) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n9436), .CLK(n9544), .Q(
        WX4696), .QN(n8022) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n9436), .CLK(n9544), .Q(
        WX4698), .QN(n8020) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n9436), .CLK(n9544), .Q(
        WX4700), .QN(n8018) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n9435), .CLK(n9545), .Q(
        WX4702), .QN(n8016) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n9435), .CLK(n9545), .Q(
        WX4704), .QN(n8014) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n9435), .CLK(n9545), .Q(
        WX4706), .QN(n8012) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n9434), .CLK(n9546), .Q(
        WX4708), .QN(n8010) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n9434), .CLK(n9546), .Q(
        WX4710), .QN(n8008) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n9434), .CLK(n9546), .Q(
        WX4712), .QN(n8006) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n9433), .CLK(n9547), .Q(
        WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n9433), .CLK(n9547), .Q(
        WX4716), .QN(n8354) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n9433), .CLK(n9547), .Q(
        WX4718), .QN(n8355) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n9433), .CLK(n9547), .Q(
        WX4720), .QN(n8356) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n9433), .CLK(n9547), .Q(
        test_so40), .QN(n8800) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n9442), .CLK(n9538), 
        .Q(WX4724), .QN(n8357) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n9442), .CLK(n9538), .Q(
        WX4726), .QN(n8358) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n9442), .CLK(n9538), .Q(
        WX4728), .QN(n8359) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n9441), .CLK(n9539), .Q(
        WX4730), .QN(n8360) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n9441), .CLK(n9539), .Q(
        WX4732) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n9441), .CLK(n9539), .Q(
        WX4734), .QN(n8362) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n9440), .CLK(n9540), .Q(
        WX4736), .QN(n8379) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n9440), .CLK(n9540), .Q(
        WX4738), .QN(n8380) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n9440), .CLK(n9540), .Q(
        WX4740), .QN(n8397) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n9439), .CLK(n9541), .Q(
        WX4742), .QN(n8398) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n9439), .CLK(n9541), .Q(
        WX4744), .QN(n8412) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n9439), .CLK(n9541), .Q(
        WX4746), .QN(n8117) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n9438), .CLK(n9542), .Q(
        WX4748), .QN(n8413) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n9438), .CLK(n9542), .Q(
        WX4750), .QN(n8414) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n9438), .CLK(n9542), .Q(
        WX4752), .QN(n8415) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n9437), .CLK(n9543), .Q(
        WX4754), .QN(n8416) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n9437), .CLK(n9543), .Q(
        test_so41), .QN(n8796) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n9437), .CLK(n9543), 
        .Q(WX4758), .QN(n8417) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n9436), .CLK(n9544), .Q(
        WX4760), .QN(n8418) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n9436), .CLK(n9544), .Q(
        WX4762), .QN(n8419) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n9436), .CLK(n9544), .Q(
        WX4764), .QN(n8420) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n9435), .CLK(n9545), .Q(
        WX4766) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n9435), .CLK(n9545), .Q(
        WX4768), .QN(n8433) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n9435), .CLK(n9545), .Q(
        WX4770), .QN(n8118) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n9434), .CLK(n9546), .Q(
        WX4772), .QN(n8450) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n9434), .CLK(n9546), .Q(
        WX4774), .QN(n8451) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n9434), .CLK(n9546), .Q(
        WX4776), .QN(n8468) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n9433), .CLK(n9547), .Q(
        WX4778), .QN(n8130) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n9353), .CLK(n9627), .Q(
        CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_3) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n9352), .CLK(n9628), 
        .Q(test_so42) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n9352), .CLK(n9628), 
        .Q(CRC_OUT_6_10) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n9352), .CLK(n9628), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n9352), .CLK(n9628), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_15) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n9351), .CLK(n9629), .Q(test_so43) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n9351), .CLK(n9629), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n9351), .CLK(n9629), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n9350), .CLK(n9630), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n9350), .CLK(n9630), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n9350), .CLK(n9630), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n9350), .CLK(n9630), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n9350), .CLK(n9630), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n9433), .CLK(n9547), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n9433), .CLK(n9547), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n973), .SI(CRC_OUT_6_31), .SE(n9433), .CLK(n9547), 
        .Q(WX5657) );
  SDFFX1 DFF_769_Q_reg ( .D(n974), .SI(WX5657), .SE(n9430), .CLK(n9550), .Q(
        n8528), .QN(n8943) );
  SDFFX1 DFF_770_Q_reg ( .D(n975), .SI(n8528), .SE(n9430), .CLK(n9550), .Q(
        n8527), .QN(n8942) );
  SDFFX1 DFF_771_Q_reg ( .D(n976), .SI(n8527), .SE(n9430), .CLK(n9550), .Q(
        n8526), .QN(n8941) );
  SDFFX1 DFF_772_Q_reg ( .D(n977), .SI(n8526), .SE(n9430), .CLK(n9550), .Q(
        n8525), .QN(n8940) );
  SDFFX1 DFF_773_Q_reg ( .D(n978), .SI(n8525), .SE(n9430), .CLK(n9550), .Q(
        n8524), .QN(n8939) );
  SDFFX1 DFF_774_Q_reg ( .D(n979), .SI(n8524), .SE(n9430), .CLK(n9550), .Q(
        n8523), .QN(n8938) );
  SDFFX1 DFF_775_Q_reg ( .D(n980), .SI(n8523), .SE(n9430), .CLK(n9550), .Q(
        test_so44), .QN(n9067) );
  SDFFX1 DFF_776_Q_reg ( .D(n981), .SI(test_si45), .SE(n9431), .CLK(n9549), 
        .Q(n8520), .QN(n8937) );
  SDFFX1 DFF_777_Q_reg ( .D(n982), .SI(n8520), .SE(n9431), .CLK(n9549), .Q(
        n8519), .QN(n8936) );
  SDFFX1 DFF_778_Q_reg ( .D(n983), .SI(n8519), .SE(n9431), .CLK(n9549), .Q(
        n8518), .QN(n8935) );
  SDFFX1 DFF_779_Q_reg ( .D(n984), .SI(n8518), .SE(n9431), .CLK(n9549), .Q(
        n8517), .QN(n8934) );
  SDFFX1 DFF_780_Q_reg ( .D(n985), .SI(n8517), .SE(n9431), .CLK(n9549), .Q(
        n8516), .QN(n8933) );
  SDFFX1 DFF_781_Q_reg ( .D(n986), .SI(n8516), .SE(n9431), .CLK(n9549), .Q(
        n8515), .QN(n8932) );
  SDFFX1 DFF_782_Q_reg ( .D(n987), .SI(n8515), .SE(n9431), .CLK(n9549), .Q(
        n8514), .QN(n8931) );
  SDFFX1 DFF_783_Q_reg ( .D(n988), .SI(n8514), .SE(n9431), .CLK(n9549), .Q(
        n8513), .QN(n8930) );
  SDFFX1 DFF_784_Q_reg ( .D(n989), .SI(n8513), .SE(n9431), .CLK(n9549), .Q(
        n8512), .QN(n8929) );
  SDFFX1 DFF_785_Q_reg ( .D(n990), .SI(n8512), .SE(n9431), .CLK(n9549), .Q(
        n8511), .QN(n8928) );
  SDFFX1 DFF_786_Q_reg ( .D(n991), .SI(n8511), .SE(n9431), .CLK(n9549), .Q(
        n8510), .QN(n8927) );
  SDFFX1 DFF_787_Q_reg ( .D(n992), .SI(n8510), .SE(n9431), .CLK(n9549), .Q(
        n8509), .QN(n8926) );
  SDFFX1 DFF_788_Q_reg ( .D(n993), .SI(n8509), .SE(n9432), .CLK(n9548), .Q(
        n8508), .QN(n8925) );
  SDFFX1 DFF_789_Q_reg ( .D(n994), .SI(n8508), .SE(n9432), .CLK(n9548), .Q(
        n8507), .QN(n8924) );
  SDFFX1 DFF_790_Q_reg ( .D(n995), .SI(n8507), .SE(n9432), .CLK(n9548), .Q(
        n8506), .QN(n8923) );
  SDFFX1 DFF_791_Q_reg ( .D(n996), .SI(n8506), .SE(n9432), .CLK(n9548), .Q(
        n8505), .QN(n8922) );
  SDFFX1 DFF_792_Q_reg ( .D(n997), .SI(n8505), .SE(n9432), .CLK(n9548), .Q(
        test_so45), .QN(n9066) );
  SDFFX1 DFF_793_Q_reg ( .D(n998), .SI(test_si46), .SE(n9432), .CLK(n9548), 
        .Q(n8502), .QN(n8921) );
  SDFFX1 DFF_794_Q_reg ( .D(n999), .SI(n8502), .SE(n9432), .CLK(n9548), .Q(
        n8501), .QN(n8920) );
  SDFFX1 DFF_795_Q_reg ( .D(n1000), .SI(n8501), .SE(n9432), .CLK(n9548), .Q(
        n8500), .QN(n8919) );
  SDFFX1 DFF_796_Q_reg ( .D(n1001), .SI(n8500), .SE(n9432), .CLK(n9548), .Q(
        n8499), .QN(n8918) );
  SDFFX1 DFF_797_Q_reg ( .D(n1002), .SI(n8499), .SE(n9432), .CLK(n9548), .Q(
        n8498), .QN(n8917) );
  SDFFX1 DFF_798_Q_reg ( .D(n1003), .SI(n8498), .SE(n9432), .CLK(n9548), .Q(
        n8497), .QN(n8916) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n9432), .CLK(n9548), .Q(
        n8496), .QN(n8915) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n9430), .CLK(n9550), .Q(
        n8495), .QN(n16072) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n9430), .CLK(n9550), .Q(
        n8494), .QN(n16073) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n9430), .CLK(n9550), .Q(
        n8493), .QN(n16074) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n9429), .CLK(n9551), .Q(
        n8492), .QN(n16075) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n9429), .CLK(n9551), .Q(
        n8491), .QN(n16076) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n9429), .CLK(n9551), .Q(
        n8490), .QN(n16077) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n9429), .CLK(n9551), .Q(
        n8489), .QN(n16078) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n9429), .CLK(n9551), .Q(
        n8488), .QN(n16079) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n9429), .CLK(n9551), .Q(
        n8487), .QN(n16080) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n9353), .CLK(n9627), .Q(
        test_so46), .QN(n8821) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n9428), .CLK(n9552), 
        .Q(n8484), .QN(n16081) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n9428), .CLK(n9552), .Q(
        n8483), .QN(n16082) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n9428), .CLK(n9552), .Q(
        n8482), .QN(n16083) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n9427), .CLK(n9553), .Q(
        n8481), .QN(n16084) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n9427), .CLK(n9553), .Q(
        n8480), .QN(n16085) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n9427), .CLK(n9553), .Q(
        n8479), .QN(n16086) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n9427), .CLK(n9553), .Q(
        WX5849), .QN(n8002) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n9427), .CLK(n9553), .Q(
        WX5851), .QN(n8000) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n9426), .CLK(n9554), .Q(
        WX5853), .QN(n7998) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n9426), .CLK(n9554), .Q(
        WX5855), .QN(n7996) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n9426), .CLK(n9554), .Q(
        WX5857), .QN(n7994) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n9425), .CLK(n9555), .Q(
        WX5859), .QN(n7992) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n9425), .CLK(n9555), .Q(
        WX5861), .QN(n7990) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n9425), .CLK(n9555), .Q(
        WX5863), .QN(n7988) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n9424), .CLK(n9556), .Q(
        WX5865), .QN(n7986) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n9424), .CLK(n9556), .Q(
        WX5867), .QN(n7984) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n9424), .CLK(n9556), .Q(
        test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n9423), .CLK(n9557), 
        .Q(WX5871), .QN(n7981) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n9423), .CLK(n9557), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n9423), .CLK(n9557), .Q(
        WX5875), .QN(n7977) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n9422), .CLK(n9558), .Q(
        WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n9422), .CLK(n9558), .Q(
        WX5879), .QN(n7974) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n9430), .CLK(n9550), .Q(
        WX5881), .QN(n7619) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n9430), .CLK(n9550), .Q(
        WX5883), .QN(n7765) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n9429), .CLK(n9551), .Q(
        WX5885), .QN(n7763) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n9429), .CLK(n9551), .Q(
        WX5887), .QN(n7761) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n9429), .CLK(n9551), .Q(
        WX5889), .QN(n7759) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n9429), .CLK(n9551), .Q(
        WX5891), .QN(n7757) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n9429), .CLK(n9551), .Q(
        WX5893), .QN(n7755) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n9429), .CLK(n9551), .Q(
        WX5895), .QN(n7753) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n9428), .CLK(n9552), .Q(
        WX5897), .QN(n7751) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n9428), .CLK(n9552), .Q(
        WX5899), .QN(n7749) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n9428), .CLK(n9552), .Q(
        WX5901), .QN(n7747) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n9428), .CLK(n9552), .Q(
        test_so48), .QN(n8812) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n9428), .CLK(n9552), 
        .Q(WX5905), .QN(n7744) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n9428), .CLK(n9552), .Q(
        WX5907), .QN(n7743) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n9427), .CLK(n9553), .Q(
        WX5909), .QN(n7741) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n9427), .CLK(n9553), .Q(
        WX5911), .QN(n7739) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n9427), .CLK(n9553), .Q(
        WX5913) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n9426), .CLK(n9554), .Q(
        WX5915) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n9426), .CLK(n9554), .Q(
        WX5917) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n9426), .CLK(n9554), .Q(
        WX5919) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n9425), .CLK(n9555), .Q(
        WX5921) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n9425), .CLK(n9555), .Q(
        WX5923) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n9425), .CLK(n9555), .Q(
        WX5925) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n9424), .CLK(n9556), .Q(
        WX5927) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n9424), .CLK(n9556), .Q(
        WX5929) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n9424), .CLK(n9556), .Q(
        WX5931) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n9423), .CLK(n9557), .Q(
        WX5933), .QN(n3669) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n9423), .CLK(n9557), .Q(
        WX5935) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n9423), .CLK(n9557), .Q(
        test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n9422), .CLK(n9558), 
        .Q(WX5939) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n9422), .CLK(n9558), .Q(
        WX5941), .QN(n3661) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n9422), .CLK(n9558), .Q(
        WX5943) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n9422), .CLK(n9558), .Q(
        WX5945), .QN(n7620) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n9421), .CLK(n9559), .Q(
        WX5947), .QN(n7766) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n9421), .CLK(n9559), .Q(
        WX5949), .QN(n7764) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n9421), .CLK(n9559), .Q(
        WX5951), .QN(n7762) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n9421), .CLK(n9559), .Q(
        WX5953), .QN(n7760) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n9421), .CLK(n9559), .Q(
        WX5955), .QN(n7758) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n9421), .CLK(n9559), .Q(
        WX5957), .QN(n7756) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n9420), .CLK(n9560), .Q(
        WX5959), .QN(n7754) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n9420), .CLK(n9560), .Q(
        WX5961), .QN(n7752) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n9420), .CLK(n9560), .Q(
        WX5963), .QN(n7750) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n9420), .CLK(n9560), .Q(
        WX5965), .QN(n7748) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n9428), .CLK(n9552), .Q(
        WX5967), .QN(n7746) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n9428), .CLK(n9552), .Q(
        WX5969), .QN(n7745) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n9428), .CLK(n9552), .Q(
        test_so50), .QN(n8811) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n9427), .CLK(n9553), 
        .Q(WX5973), .QN(n7742) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n9427), .CLK(n9553), .Q(
        WX5975), .QN(n7740) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n9427), .CLK(n9553), .Q(
        WX5977), .QN(n8003) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n9426), .CLK(n9554), .Q(
        WX5979), .QN(n8001) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n9426), .CLK(n9554), .Q(
        WX5981), .QN(n7999) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n9426), .CLK(n9554), .Q(
        WX5983), .QN(n7997) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n9425), .CLK(n9555), .Q(
        WX5985), .QN(n7995) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n9425), .CLK(n9555), .Q(
        WX5987), .QN(n7993) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n9425), .CLK(n9555), .Q(
        WX5989), .QN(n7991) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n9424), .CLK(n9556), .Q(
        WX5991), .QN(n7989) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n9424), .CLK(n9556), .Q(
        WX5993), .QN(n7987) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n9424), .CLK(n9556), .Q(
        WX5995), .QN(n7985) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n9423), .CLK(n9557), .Q(
        WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n9423), .CLK(n9557), .Q(
        WX5999), .QN(n7982) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n9423), .CLK(n9557), .Q(
        WX6001), .QN(n7980) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n9422), .CLK(n9558), .Q(
        WX6003), .QN(n7978) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n9422), .CLK(n9558), .Q(
        test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n9422), .CLK(n9558), 
        .Q(WX6007), .QN(n7975) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n9421), .CLK(n9559), .Q(
        WX6009), .QN(n8238) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n9421), .CLK(n9559), .Q(
        WX6011), .QN(n8239) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n9421), .CLK(n9559), .Q(
        WX6013), .QN(n8240) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n9421), .CLK(n9559), .Q(
        WX6015), .QN(n8241) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n9421), .CLK(n9559), .Q(
        WX6017), .QN(n8242) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n9421), .CLK(n9559), .Q(
        WX6019), .QN(n8243) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n9420), .CLK(n9560), .Q(
        WX6021), .QN(n8244) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n9420), .CLK(n9560), .Q(
        WX6023), .QN(n8245) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n9420), .CLK(n9560), .Q(
        WX6025), .QN(n8255) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n9420), .CLK(n9560), .Q(
        WX6027), .QN(n8256) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n9420), .CLK(n9560), .Q(
        WX6029), .QN(n8273) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n9420), .CLK(n9560), .Q(
        WX6031), .QN(n8274) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n9420), .CLK(n9560), .Q(
        WX6033), .QN(n8291) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n9420), .CLK(n9560), .Q(
        WX6035), .QN(n8292) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n9419), .CLK(n9561), .Q(
        WX6037), .QN(n8296) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n9419), .CLK(n9561), .Q(
        test_so52), .QN(n8826) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n9427), .CLK(n9553), 
        .Q(WX6041), .QN(n8297) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n9426), .CLK(n9554), .Q(
        WX6043), .QN(n8298) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n9426), .CLK(n9554), .Q(
        WX6045), .QN(n8299) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n9426), .CLK(n9554), .Q(
        WX6047), .QN(n8300) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n9425), .CLK(n9555), .Q(
        WX6049), .QN(n8115) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n9425), .CLK(n9555), .Q(
        WX6051), .QN(n8301) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n9425), .CLK(n9555), .Q(
        WX6053), .QN(n8302) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n9424), .CLK(n9556), .Q(
        WX6055), .QN(n8303) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n9424), .CLK(n9556), .Q(
        WX6057), .QN(n8308) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n9424), .CLK(n9556), .Q(
        WX6059), .QN(n8309) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n9423), .CLK(n9557), .Q(
        WX6061), .QN(n8326) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n9423), .CLK(n9557), .Q(
        WX6063), .QN(n8116) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n9423), .CLK(n9557), .Q(
        WX6065), .QN(n8327) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n9422), .CLK(n9558), .Q(
        WX6067), .QN(n8344) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n9422), .CLK(n9558), .Q(
        WX6069), .QN(n8345) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n9422), .CLK(n9558), .Q(
        WX6071), .QN(n8129) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n9354), .CLK(n9626), .Q(
        test_so53) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_3) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n9354), .CLK(n9626), 
        .Q(CRC_OUT_5_10) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n9353), .CLK(n9627), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n9353), .CLK(n9627), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n9353), .CLK(n9627), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n9353), .CLK(n9627), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n9353), .CLK(n9627), .Q(CRC_OUT_5_15) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n9353), .CLK(n9627), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n9353), .CLK(n9627), .Q(test_so54), .QN(n8827) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n9353), .CLK(n9627), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n9353), .CLK(n9627), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n9353), .CLK(n9627), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n9419), .CLK(n9561), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n9418), .CLK(n9562), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n1214), .SI(CRC_OUT_5_31), .SE(n9418), .CLK(n9562), 
        .Q(WX6950) );
  SDFFX1 DFF_961_Q_reg ( .D(n1215), .SI(WX6950), .SE(n9416), .CLK(n9564), .Q(
        n8470), .QN(n8914) );
  SDFFX1 DFF_962_Q_reg ( .D(n1216), .SI(n8470), .SE(n9416), .CLK(n9564), .Q(
        test_so55), .QN(n9065) );
  SDFFX1 DFF_963_Q_reg ( .D(n1217), .SI(test_si56), .SE(n9416), .CLK(n9564), 
        .Q(n8467), .QN(n8913) );
  SDFFX1 DFF_964_Q_reg ( .D(n1218), .SI(n8467), .SE(n9416), .CLK(n9564), .Q(
        n8466), .QN(n8912) );
  SDFFX1 DFF_965_Q_reg ( .D(n1219), .SI(n8466), .SE(n9416), .CLK(n9564), .Q(
        n8465), .QN(n8911) );
  SDFFX1 DFF_966_Q_reg ( .D(n1220), .SI(n8465), .SE(n9416), .CLK(n9564), .Q(
        n8464), .QN(n8910) );
  SDFFX1 DFF_967_Q_reg ( .D(n1221), .SI(n8464), .SE(n9416), .CLK(n9564), .Q(
        n8463), .QN(n8909) );
  SDFFX1 DFF_968_Q_reg ( .D(n1222), .SI(n8463), .SE(n9416), .CLK(n9564), .Q(
        n8462), .QN(n8908) );
  SDFFX1 DFF_969_Q_reg ( .D(n1223), .SI(n8462), .SE(n9416), .CLK(n9564), .Q(
        n8461), .QN(n8907) );
  SDFFX1 DFF_970_Q_reg ( .D(n1224), .SI(n8461), .SE(n9417), .CLK(n9563), .Q(
        n8460), .QN(n8906) );
  SDFFX1 DFF_971_Q_reg ( .D(n1225), .SI(n8460), .SE(n9417), .CLK(n9563), .Q(
        n8459), .QN(n8905) );
  SDFFX1 DFF_972_Q_reg ( .D(n1226), .SI(n8459), .SE(n9417), .CLK(n9563), .Q(
        n8458), .QN(n8904) );
  SDFFX1 DFF_973_Q_reg ( .D(n1227), .SI(n8458), .SE(n9417), .CLK(n9563), .Q(
        n8457), .QN(n8903) );
  SDFFX1 DFF_974_Q_reg ( .D(n1228), .SI(n8457), .SE(n9417), .CLK(n9563), .Q(
        n8456), .QN(n8902) );
  SDFFX1 DFF_975_Q_reg ( .D(n1229), .SI(n8456), .SE(n9417), .CLK(n9563), .Q(
        n8455), .QN(n8901) );
  SDFFX1 DFF_976_Q_reg ( .D(n1230), .SI(n8455), .SE(n9417), .CLK(n9563), .Q(
        n8454), .QN(n8900) );
  SDFFX1 DFF_977_Q_reg ( .D(n1231), .SI(n8454), .SE(n9417), .CLK(n9563), .Q(
        n8453), .QN(n8899) );
  SDFFX1 DFF_978_Q_reg ( .D(n1232), .SI(n8453), .SE(n9417), .CLK(n9563), .Q(
        n8452), .QN(n8898) );
  SDFFX1 DFF_979_Q_reg ( .D(n1233), .SI(n8452), .SE(n9417), .CLK(n9563), .Q(
        test_so56), .QN(n9064) );
  SDFFX1 DFF_980_Q_reg ( .D(n1234), .SI(test_si57), .SE(n9417), .CLK(n9563), 
        .Q(n8449), .QN(n8897) );
  SDFFX1 DFF_981_Q_reg ( .D(n1235), .SI(n8449), .SE(n9417), .CLK(n9563), .Q(
        n8448), .QN(n8896) );
  SDFFX1 DFF_982_Q_reg ( .D(n1236), .SI(n8448), .SE(n9418), .CLK(n9562), .Q(
        n8447), .QN(n8895) );
  SDFFX1 DFF_983_Q_reg ( .D(n1237), .SI(n8447), .SE(n9418), .CLK(n9562), .Q(
        n8446), .QN(n8894) );
  SDFFX1 DFF_984_Q_reg ( .D(n1238), .SI(n8446), .SE(n9418), .CLK(n9562), .Q(
        n8445), .QN(n8893) );
  SDFFX1 DFF_985_Q_reg ( .D(n1239), .SI(n8445), .SE(n9418), .CLK(n9562), .Q(
        n8444), .QN(n8892) );
  SDFFX1 DFF_986_Q_reg ( .D(n1240), .SI(n8444), .SE(n9418), .CLK(n9562), .Q(
        n8443), .QN(n8891) );
  SDFFX1 DFF_987_Q_reg ( .D(n1241), .SI(n8443), .SE(n9418), .CLK(n9562), .Q(
        n8442), .QN(n8890) );
  SDFFX1 DFF_988_Q_reg ( .D(n1242), .SI(n8442), .SE(n9418), .CLK(n9562), .Q(
        n8441), .QN(n8889) );
  SDFFX1 DFF_989_Q_reg ( .D(n1243), .SI(n8441), .SE(n9418), .CLK(n9562), .Q(
        n8440), .QN(n8888) );
  SDFFX1 DFF_990_Q_reg ( .D(n1244), .SI(n8440), .SE(n9418), .CLK(n9562), .Q(
        n8439), .QN(n8887) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n9418), .CLK(n9562), .Q(
        n8438), .QN(n8886) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n9416), .CLK(n9564), .Q(
        n8437), .QN(n16087) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n9415), .CLK(n9565), .Q(
        n8436), .QN(n16088) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n9415), .CLK(n9565), .Q(
        n8435), .QN(n16089) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n9415), .CLK(n9565), .Q(
        n8434), .QN(n16090) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n9415), .CLK(n9565), .Q(
        test_so57), .QN(n8820) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n9415), .CLK(n9565), 
        .Q(n8431), .QN(n16091) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n9415), .CLK(n9565), .Q(
        n8430), .QN(n16092) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n9414), .CLK(n9566), .Q(
        n8429), .QN(n16093) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n9414), .CLK(n9566), .Q(
        n8428), .QN(n16094) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n9414), .CLK(n9566), .Q(
        n8427), .QN(n16095) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n9414), .CLK(n9566), .Q(
        n8426), .QN(n16096) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n9413), .CLK(n9567), .Q(
        n8425), .QN(n16097) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n9413), .CLK(n9567), .Q(
        n8424), .QN(n16098) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n9413), .CLK(n9567), .Q(
        n8423), .QN(n16099) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n9412), .CLK(n9568), .Q(
        n8422), .QN(n16100) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n9412), .CLK(n9568), .Q(
        n8421), .QN(n16101) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n9412), .CLK(n9568), .Q(
        WX7142), .QN(n7972) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n9411), .CLK(n9569), 
        .Q(WX7144), .QN(n7970) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n9411), .CLK(n9569), 
        .Q(WX7146), .QN(n7968) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n9411), .CLK(n9569), 
        .Q(WX7148), .QN(n7966) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n9410), .CLK(n9570), 
        .Q(WX7150), .QN(n7964) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n9410), .CLK(n9570), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n9410), .CLK(n9570), 
        .Q(WX7154), .QN(n7961) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n9409), .CLK(n9571), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n9409), .CLK(n9571), 
        .Q(WX7158), .QN(n7957) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n9409), .CLK(n9571), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n9408), .CLK(n9572), 
        .Q(WX7162), .QN(n7954) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n9408), .CLK(n9572), 
        .Q(WX7164), .QN(n7952) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n9408), .CLK(n9572), 
        .Q(WX7166), .QN(n7950) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n9407), .CLK(n9573), 
        .Q(WX7168), .QN(n7948) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n9407), .CLK(n9573), 
        .Q(WX7170), .QN(n7946) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n9407), .CLK(n9573), 
        .Q(WX7172), .QN(n7944) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n9416), .CLK(n9564), 
        .Q(WX7174), .QN(n7617) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n9416), .CLK(n9564), 
        .Q(WX7176), .QN(n7737) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n9415), .CLK(n9565), 
        .Q(WX7178), .QN(n7735) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n9415), .CLK(n9565), 
        .Q(WX7180), .QN(n7733) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n9415), .CLK(n9565), 
        .Q(WX7182), .QN(n7731) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n9415), .CLK(n9565), 
        .Q(WX7184), .QN(n7729) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n9415), .CLK(n9565), 
        .Q(test_so59), .QN(n8810) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n9414), .CLK(n9566), 
        .Q(WX7188), .QN(n7726) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n9414), .CLK(n9566), 
        .Q(WX7190), .QN(n7725) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n9414), .CLK(n9566), 
        .Q(WX7192), .QN(n7723) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n9414), .CLK(n9566), 
        .Q(WX7194), .QN(n7721) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n9413), .CLK(n9567), 
        .Q(WX7196), .QN(n7719) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n9413), .CLK(n9567), 
        .Q(WX7198), .QN(n7717) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n9413), .CLK(n9567), 
        .Q(WX7200), .QN(n7715) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n9412), .CLK(n9568), 
        .Q(WX7202), .QN(n7713) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n9412), .CLK(n9568), 
        .Q(WX7204), .QN(n7711) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n9412), .CLK(n9568), 
        .Q(WX7206) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n9411), .CLK(n9569), 
        .Q(WX7208) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n9411), .CLK(n9569), 
        .Q(WX7210) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n9411), .CLK(n9569), 
        .Q(WX7212) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n9410), .CLK(n9570), 
        .Q(WX7214) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n9410), .CLK(n9570), 
        .Q(WX7216), .QN(n3647) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n9410), .CLK(n9570), 
        .Q(WX7218) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n9409), .CLK(n9571), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n9409), .CLK(n9571), 
        .Q(WX7222) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n9409), .CLK(n9571), 
        .Q(WX7224), .QN(n3639) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n9408), .CLK(n9572), 
        .Q(WX7226) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n9408), .CLK(n9572), 
        .Q(WX7228), .QN(n3635) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n9408), .CLK(n9572), 
        .Q(WX7230) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n9407), .CLK(n9573), 
        .Q(WX7232) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n9407), .CLK(n9573), 
        .Q(WX7234) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n9407), .CLK(n9573), 
        .Q(WX7236) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n9406), .CLK(n9574), 
        .Q(WX7238), .QN(n7618) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n9406), .CLK(n9574), 
        .Q(WX7240), .QN(n7738) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n9406), .CLK(n9574), 
        .Q(WX7242), .QN(n7736) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n9406), .CLK(n9574), 
        .Q(WX7244), .QN(n7734) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n9406), .CLK(n9574), 
        .Q(WX7246), .QN(n7732) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n9406), .CLK(n9574), 
        .Q(WX7248), .QN(n7730) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n9415), .CLK(n9565), 
        .Q(WX7250), .QN(n7728) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n9414), .CLK(n9566), 
        .Q(WX7252), .QN(n7727) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n9414), .CLK(n9566), 
        .Q(test_so61), .QN(n8809) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n9414), .CLK(n9566), 
        .Q(WX7256), .QN(n7724) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n9414), .CLK(n9566), 
        .Q(WX7258), .QN(n7722) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n9413), .CLK(n9567), 
        .Q(WX7260), .QN(n7720) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n9413), .CLK(n9567), 
        .Q(WX7262), .QN(n7718) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n9413), .CLK(n9567), 
        .Q(WX7264), .QN(n7716) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n9412), .CLK(n9568), 
        .Q(WX7266), .QN(n7714) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n9412), .CLK(n9568), 
        .Q(WX7268), .QN(n7712) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n9412), .CLK(n9568), 
        .Q(WX7270), .QN(n7973) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n9411), .CLK(n9569), 
        .Q(WX7272), .QN(n7971) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n9411), .CLK(n9569), 
        .Q(WX7274), .QN(n7969) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n9411), .CLK(n9569), 
        .Q(WX7276), .QN(n7967) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n9410), .CLK(n9570), 
        .Q(WX7278), .QN(n7965) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n9410), .CLK(n9570), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n9410), .CLK(n9570), 
        .Q(WX7282), .QN(n7962) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n9409), .CLK(n9571), 
        .Q(WX7284), .QN(n7960) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n9409), .CLK(n9571), 
        .Q(WX7286), .QN(n7958) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n9409), .CLK(n9571), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n9408), .CLK(n9572), 
        .Q(WX7290), .QN(n7955) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n9408), .CLK(n9572), 
        .Q(WX7292), .QN(n7953) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n9408), .CLK(n9572), 
        .Q(WX7294), .QN(n7951) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n9407), .CLK(n9573), 
        .Q(WX7296), .QN(n7949) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n9407), .CLK(n9573), 
        .Q(WX7298), .QN(n7947) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n9407), .CLK(n9573), 
        .Q(WX7300), .QN(n7945) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n9406), .CLK(n9574), 
        .Q(WX7302), .QN(n8211) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n9406), .CLK(n9574), 
        .Q(WX7304) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n9406), .CLK(n9574), 
        .Q(WX7306), .QN(n8213) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n9406), .CLK(n9574), 
        .Q(WX7308), .QN(n8214) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n9406), .CLK(n9574), 
        .Q(WX7310), .QN(n8215) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n9406), .CLK(n9574), 
        .Q(WX7312), .QN(n8216) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n9405), .CLK(n9575), 
        .Q(WX7314), .QN(n8217) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n9405), .CLK(n9575), 
        .Q(WX7316), .QN(n8218) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n9405), .CLK(n9575), 
        .Q(WX7318), .QN(n8219) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n9405), .CLK(n9575), 
        .Q(WX7320), .QN(n8220) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n9405), .CLK(n9575), 
        .Q(test_so63), .QN(n8799) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n9413), .CLK(n9567), 
        .Q(WX7324), .QN(n8221) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n9413), .CLK(n9567), 
        .Q(WX7326), .QN(n8222) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n9413), .CLK(n9567), 
        .Q(WX7328), .QN(n8223) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n9412), .CLK(n9568), 
        .Q(WX7330), .QN(n8224) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n9412), .CLK(n9568), 
        .Q(WX7332), .QN(n8113) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n9412), .CLK(n9568), 
        .Q(WX7334), .QN(n8225) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n9411), .CLK(n9569), 
        .Q(WX7336), .QN(n8226) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n9411), .CLK(n9569), 
        .Q(WX7338) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n9411), .CLK(n9569), 
        .Q(WX7340), .QN(n8228) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n9410), .CLK(n9570), 
        .Q(WX7342), .QN(n8114) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n9410), .CLK(n9570), 
        .Q(WX7344), .QN(n8229) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n9410), .CLK(n9570), 
        .Q(WX7346), .QN(n8230) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n9409), .CLK(n9571), 
        .Q(WX7348), .QN(n8231) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n9409), .CLK(n9571), 
        .Q(WX7350), .QN(n8232) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n9409), .CLK(n9571), 
        .Q(WX7352), .QN(n8233) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n9408), .CLK(n9572), 
        .Q(WX7354), .QN(n8234) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n9408), .CLK(n9572), 
        .Q(test_so64), .QN(n8795) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n9408), .CLK(n9572), 
        .Q(WX7358), .QN(n8235) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n9407), .CLK(n9573), 
        .Q(WX7360), .QN(n8236) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n9407), .CLK(n9573), 
        .Q(WX7362), .QN(n8237) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n9407), .CLK(n9573), 
        .Q(WX7364), .QN(n8128) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n9357), .CLK(n9623), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_3) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n9356), .CLK(n9624), .Q(CRC_OUT_4_10) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n9356), .CLK(
        n9624), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n9356), .CLK(
        n9624), .Q(test_so65) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n9355), .CLK(n9625), 
        .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_15) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n9355), .CLK(
        n9625), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n9354), .CLK(
        n9626), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n9405), .CLK(
        n9575), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n9405), .CLK(
        n9575), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n9405), .CLK(
        n9575), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n9405), .CLK(
        n9575), .Q(test_so66) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n9405), .CLK(n9575), 
        .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n9405), .CLK(
        n9575), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n1455), .SI(CRC_OUT_4_31), .SE(n9405), .CLK(n9575), .Q(WX8243) );
  SDFFX1 DFF_1153_Q_reg ( .D(n1456), .SI(WX8243), .SE(n9402), .CLK(n9578), .Q(
        n8411), .QN(n8885) );
  SDFFX1 DFF_1154_Q_reg ( .D(n1457), .SI(n8411), .SE(n9402), .CLK(n9578), .Q(
        n8410), .QN(n8884) );
  SDFFX1 DFF_1155_Q_reg ( .D(n1458), .SI(n8410), .SE(n9402), .CLK(n9578), .Q(
        n8409), .QN(n8883) );
  SDFFX1 DFF_1156_Q_reg ( .D(n1459), .SI(n8409), .SE(n9402), .CLK(n9578), .Q(
        n8408), .QN(n8882) );
  SDFFX1 DFF_1157_Q_reg ( .D(n1460), .SI(n8408), .SE(n9402), .CLK(n9578), .Q(
        n8407), .QN(n8881) );
  SDFFX1 DFF_1158_Q_reg ( .D(n1461), .SI(n8407), .SE(n9402), .CLK(n9578), .Q(
        n8406), .QN(n8880) );
  SDFFX1 DFF_1159_Q_reg ( .D(n1462), .SI(n8406), .SE(n9402), .CLK(n9578), .Q(
        n8405), .QN(n8879) );
  SDFFX1 DFF_1160_Q_reg ( .D(n1463), .SI(n8405), .SE(n9403), .CLK(n9577), .Q(
        n8404), .QN(n8878) );
  SDFFX1 DFF_1161_Q_reg ( .D(n1464), .SI(n8404), .SE(n9403), .CLK(n9577), .Q(
        n8403), .QN(n8877) );
  SDFFX1 DFF_1162_Q_reg ( .D(n1465), .SI(n8403), .SE(n9403), .CLK(n9577), .Q(
        n8402), .QN(n8876) );
  SDFFX1 DFF_1163_Q_reg ( .D(n1466), .SI(n8402), .SE(n9403), .CLK(n9577), .Q(
        n8401), .QN(n8875) );
  SDFFX1 DFF_1164_Q_reg ( .D(n1467), .SI(n8401), .SE(n9403), .CLK(n9577), .Q(
        n8400), .QN(n8874) );
  SDFFX1 DFF_1165_Q_reg ( .D(n1468), .SI(n8400), .SE(n9403), .CLK(n9577), .Q(
        n8399), .QN(n8873) );
  SDFFX1 DFF_1166_Q_reg ( .D(n1469), .SI(n8399), .SE(n9403), .CLK(n9577), .Q(
        test_so67), .QN(n9063) );
  SDFFX1 DFF_1167_Q_reg ( .D(n1470), .SI(test_si68), .SE(n9403), .CLK(n9577), 
        .Q(n8396), .QN(n8872) );
  SDFFX1 DFF_1168_Q_reg ( .D(n1471), .SI(n8396), .SE(n9403), .CLK(n9577), .Q(
        n8395), .QN(n8871) );
  SDFFX1 DFF_1169_Q_reg ( .D(n1472), .SI(n8395), .SE(n9403), .CLK(n9577), .Q(
        n8394), .QN(n8870) );
  SDFFX1 DFF_1170_Q_reg ( .D(n1473), .SI(n8394), .SE(n9403), .CLK(n9577), .Q(
        n8393), .QN(n8869) );
  SDFFX1 DFF_1171_Q_reg ( .D(n1474), .SI(n8393), .SE(n9403), .CLK(n9577), .Q(
        n8392), .QN(n8868) );
  SDFFX1 DFF_1172_Q_reg ( .D(n1475), .SI(n8392), .SE(n9404), .CLK(n9576), .Q(
        n8391), .QN(n8867) );
  SDFFX1 DFF_1173_Q_reg ( .D(n1476), .SI(n8391), .SE(n9404), .CLK(n9576), .Q(
        n8390), .QN(n8866) );
  SDFFX1 DFF_1174_Q_reg ( .D(n1477), .SI(n8390), .SE(n9404), .CLK(n9576), .Q(
        n8389), .QN(n8865) );
  SDFFX1 DFF_1175_Q_reg ( .D(n1478), .SI(n8389), .SE(n9404), .CLK(n9576), .Q(
        n8388), .QN(n8864) );
  SDFFX1 DFF_1176_Q_reg ( .D(n1479), .SI(n8388), .SE(n9404), .CLK(n9576), .Q(
        n8387), .QN(n8863) );
  SDFFX1 DFF_1177_Q_reg ( .D(n1480), .SI(n8387), .SE(n9404), .CLK(n9576), .Q(
        n8386), .QN(n8862) );
  SDFFX1 DFF_1178_Q_reg ( .D(n1481), .SI(n8386), .SE(n9404), .CLK(n9576), .Q(
        n8385), .QN(n8861) );
  SDFFX1 DFF_1179_Q_reg ( .D(n1482), .SI(n8385), .SE(n9404), .CLK(n9576), .Q(
        n8384), .QN(n8860) );
  SDFFX1 DFF_1180_Q_reg ( .D(n1483), .SI(n8384), .SE(n9404), .CLK(n9576), .Q(
        n8383), .QN(n8859) );
  SDFFX1 DFF_1181_Q_reg ( .D(n1484), .SI(n8383), .SE(n9404), .CLK(n9576), .Q(
        n8382), .QN(n8858) );
  SDFFX1 DFF_1182_Q_reg ( .D(n1485), .SI(n8382), .SE(n9404), .CLK(n9576), .Q(
        n8381), .QN(n8857) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n9404), .CLK(n9576), .Q(
        test_so68), .QN(n9062) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n9402), .CLK(n9578), 
        .Q(n8378), .QN(n16102) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n9402), .CLK(n9578), .Q(
        n8377), .QN(n16103) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n9402), .CLK(n9578), .Q(
        n8376), .QN(n16104) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n9401), .CLK(n9579), .Q(
        n8375), .QN(n16105) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n9401), .CLK(n9579), .Q(
        n8374), .QN(n16106) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n9401), .CLK(n9579), .Q(
        n8373), .QN(n16107) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n9401), .CLK(n9579), .Q(
        n8372), .QN(n16108) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n9400), .CLK(n9580), .Q(
        n8371), .QN(n16109) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n9400), .CLK(n9580), .Q(
        n8370), .QN(n16110) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n9399), .CLK(n9581), .Q(
        n8369), .QN(n16111) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n9399), .CLK(n9581), .Q(
        n8368), .QN(n16112) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n9399), .CLK(n9581), .Q(
        n8367), .QN(n16113) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n9399), .CLK(n9581), .Q(
        n8366), .QN(n16114) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n9398), .CLK(n9582), .Q(
        n8365), .QN(n16115) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n9398), .CLK(n9582), .Q(
        n8364), .QN(n16116) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n9397), .CLK(n9583), .Q(
        n8363), .QN(n16117) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n9397), .CLK(n9583), .Q(
        test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n9397), .CLK(n9583), 
        .Q(WX8437), .QN(n7941) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n9397), .CLK(n9583), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n9396), .CLK(n9584), 
        .Q(WX8441), .QN(n7937) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n9396), .CLK(n9584), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n9396), .CLK(n9584), 
        .Q(WX8445), .QN(n7934) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n9395), .CLK(n9585), 
        .Q(WX8447), .QN(n7932) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n9395), .CLK(n9585), 
        .Q(WX8449), .QN(n7930) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n9395), .CLK(n9585), 
        .Q(WX8451), .QN(n7928) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n9394), .CLK(n9586), 
        .Q(WX8453), .QN(n7926) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n9394), .CLK(n9586), 
        .Q(WX8455), .QN(n7924) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n9394), .CLK(n9586), 
        .Q(WX8457), .QN(n7922) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n9393), .CLK(n9587), 
        .Q(WX8459), .QN(n7920) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n9393), .CLK(n9587), 
        .Q(WX8461), .QN(n7918) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n9393), .CLK(n9587), 
        .Q(WX8463), .QN(n7916) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n9392), .CLK(n9588), 
        .Q(WX8465), .QN(n7914) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n9402), .CLK(n9578), 
        .Q(WX8467), .QN(n7615) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n9402), .CLK(n9578), 
        .Q(test_so70), .QN(n8808) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n9401), .CLK(n9579), 
        .Q(WX8471), .QN(n7708) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n9401), .CLK(n9579), 
        .Q(WX8473), .QN(n7707) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n9401), .CLK(n9579), 
        .Q(WX8475), .QN(n7705) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n9401), .CLK(n9579), 
        .Q(WX8477), .QN(n7703) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n9401), .CLK(n9579), 
        .Q(WX8479), .QN(n7701) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n9400), .CLK(n9580), 
        .Q(WX8481), .QN(n7699) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n9400), .CLK(n9580), 
        .Q(WX8483), .QN(n7697) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n9400), .CLK(n9580), 
        .Q(WX8485), .QN(n7695) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n9399), .CLK(n9581), 
        .Q(WX8487), .QN(n7693) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n9399), .CLK(n9581), 
        .Q(WX8489), .QN(n7691) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n9399), .CLK(n9581), 
        .Q(WX8491), .QN(n7689) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n9398), .CLK(n9582), 
        .Q(WX8493), .QN(n7687) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n9398), .CLK(n9582), 
        .Q(WX8495), .QN(n7685) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n9398), .CLK(n9582), 
        .Q(WX8497), .QN(n7683) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n9397), .CLK(n9583), 
        .Q(WX8499), .QN(n3625) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n9397), .CLK(n9583), 
        .Q(WX8501) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n9397), .CLK(n9583), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n9396), .CLK(n9584), 
        .Q(WX8505) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n9396), .CLK(n9584), 
        .Q(WX8507), .QN(n3617) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n9396), .CLK(n9584), 
        .Q(WX8509) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n9395), .CLK(n9585), 
        .Q(WX8511), .QN(n3613) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n9395), .CLK(n9585), 
        .Q(WX8513) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n9395), .CLK(n9585), 
        .Q(WX8515) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n9394), .CLK(n9586), 
        .Q(WX8517) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n9394), .CLK(n9586), 
        .Q(WX8519) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n9394), .CLK(n9586), 
        .Q(WX8521) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n9393), .CLK(n9587), 
        .Q(WX8523) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n9393), .CLK(n9587), 
        .Q(WX8525) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n9393), .CLK(n9587), 
        .Q(WX8527) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n9392), .CLK(n9588), 
        .Q(WX8529) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n9392), .CLK(n9588), 
        .Q(WX8531), .QN(n7616) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n9392), .CLK(n9588), 
        .Q(WX8533), .QN(n7710) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n9392), .CLK(n9588), 
        .Q(WX8535), .QN(n7709) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n9392), .CLK(n9588), 
        .Q(test_so72), .QN(n8807) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n9401), .CLK(n9579), 
        .Q(WX8539), .QN(n7706) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n9401), .CLK(n9579), 
        .Q(WX8541), .QN(n7704) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n9401), .CLK(n9579), 
        .Q(WX8543), .QN(n7702) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n9400), .CLK(n9580), 
        .Q(WX8545), .QN(n7700) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n9400), .CLK(n9580), 
        .Q(WX8547), .QN(n7698) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n9400), .CLK(n9580), 
        .Q(WX8549), .QN(n7696) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n9399), .CLK(n9581), 
        .Q(WX8551), .QN(n7694) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n9399), .CLK(n9581), 
        .Q(WX8553), .QN(n7692) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n9399), .CLK(n9581), 
        .Q(WX8555), .QN(n7690) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n9398), .CLK(n9582), 
        .Q(WX8557), .QN(n7688) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n9398), .CLK(n9582), 
        .Q(WX8559), .QN(n7686) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n9398), .CLK(n9582), 
        .Q(WX8561), .QN(n7684) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n9397), .CLK(n9583), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n9397), .CLK(n9583), 
        .Q(WX8565), .QN(n7942) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n9397), .CLK(n9583), 
        .Q(WX8567), .QN(n7940) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n9396), .CLK(n9584), 
        .Q(WX8569), .QN(n7938) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n9396), .CLK(n9584), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n9396), .CLK(n9584), 
        .Q(WX8573), .QN(n7935) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n9395), .CLK(n9585), 
        .Q(WX8575), .QN(n7933) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n9395), .CLK(n9585), 
        .Q(WX8577), .QN(n7931) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n9395), .CLK(n9585), 
        .Q(WX8579), .QN(n7929) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n9394), .CLK(n9586), 
        .Q(WX8581), .QN(n7927) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n9394), .CLK(n9586), 
        .Q(WX8583), .QN(n7925) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n9394), .CLK(n9586), 
        .Q(WX8585), .QN(n7923) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n9393), .CLK(n9587), 
        .Q(WX8587), .QN(n7921) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n9393), .CLK(n9587), 
        .Q(WX8589), .QN(n7919) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n9393), .CLK(n9587), 
        .Q(WX8591), .QN(n7917) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n9392), .CLK(n9588), 
        .Q(WX8593), .QN(n7915) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n9392), .CLK(n9588), 
        .Q(WX8595), .QN(n8185) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n9392), .CLK(n9588), 
        .Q(WX8597), .QN(n8186) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n9392), .CLK(n9588), 
        .Q(WX8599), .QN(n8187) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n9391), .CLK(n9589), 
        .Q(WX8601), .QN(n8188) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n9391), .CLK(n9589), 
        .Q(WX8603), .QN(n8189) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n9391), .CLK(n9589), 
        .Q(test_so74), .QN(n8798) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n9400), .CLK(n9580), 
        .Q(WX8607) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n9400), .CLK(n9580), 
        .Q(WX8609), .QN(n8191) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n9400), .CLK(n9580), 
        .Q(WX8611), .QN(n8192) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n9400), .CLK(n9580), 
        .Q(WX8613), .QN(n8193) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n9399), .CLK(n9581), 
        .Q(WX8615), .QN(n8194) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n9399), .CLK(n9581), 
        .Q(WX8617), .QN(n8195) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n9398), .CLK(n9582), 
        .Q(WX8619), .QN(n8196) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n9398), .CLK(n9582), 
        .Q(WX8621), .QN(n8197) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n9398), .CLK(n9582), 
        .Q(WX8623), .QN(n8198) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n9398), .CLK(n9582), 
        .Q(WX8625), .QN(n8110) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n9397), .CLK(n9583), 
        .Q(WX8627), .QN(n8199) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n9397), .CLK(n9583), 
        .Q(WX8629), .QN(n8200) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n9396), .CLK(n9584), 
        .Q(WX8631), .QN(n8201) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n9396), .CLK(n9584), 
        .Q(WX8633), .QN(n8202) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n9396), .CLK(n9584), 
        .Q(WX8635), .QN(n8111) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n9395), .CLK(n9585), 
        .Q(WX8637), .QN(n8203) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n9395), .CLK(n9585), 
        .Q(test_so75), .QN(n8790) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n9395), .CLK(n9585), 
        .Q(WX8641) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n9394), .CLK(n9586), 
        .Q(WX8643), .QN(n8205) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n9394), .CLK(n9586), 
        .Q(WX8645), .QN(n8206) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n9394), .CLK(n9586), 
        .Q(WX8647), .QN(n8207) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n9393), .CLK(n9587), 
        .Q(WX8649), .QN(n8112) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n9393), .CLK(n9587), 
        .Q(WX8651), .QN(n8208) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n9393), .CLK(n9587), 
        .Q(WX8653), .QN(n8209) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n9392), .CLK(n9588), 
        .Q(WX8655), .QN(n8210) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n9392), .CLK(n9588), 
        .Q(WX8657), .QN(n8127) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n9359), .CLK(n9621), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n9359), .CLK(n9621), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n9359), .CLK(n9621), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n9359), .CLK(n9621), .Q(CRC_OUT_3_3) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n9359), .CLK(n9621), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n9358), .CLK(n9622), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n9358), .CLK(n9622), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n9358), .CLK(n9622), .Q(test_so76) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n9358), .CLK(n9622), 
        .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n9358), .CLK(n9622), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n9358), .CLK(n9622), .Q(CRC_OUT_3_10) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n9358), .CLK(
        n9622), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n9358), .CLK(
        n9622), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n9358), .CLK(
        n9622), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n9358), .CLK(
        n9622), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n9358), .CLK(
        n9622), .Q(CRC_OUT_3_15) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n9358), .CLK(
        n9622), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n9357), .CLK(
        n9623), .Q(test_so77) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n9357), .CLK(n9623), 
        .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n9357), .CLK(
        n9623), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n9391), .CLK(
        n9589), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n9391), .CLK(
        n9589), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n9391), .CLK(
        n9589), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n9391), .CLK(
        n9589), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n1697), .SI(CRC_OUT_3_31), .SE(n9391), .CLK(n9589), .Q(WX9536) );
  SDFFX1 DFF_1345_Q_reg ( .D(n1698), .SI(WX9536), .SE(n9388), .CLK(n9592), .Q(
        n8353), .QN(n8856) );
  SDFFX1 DFF_1346_Q_reg ( .D(n1699), .SI(n8353), .SE(n9388), .CLK(n9592), .Q(
        n8352), .QN(n8855) );
  SDFFX1 DFF_1347_Q_reg ( .D(n1700), .SI(n8352), .SE(n9388), .CLK(n9592), .Q(
        n8351), .QN(n8854) );
  SDFFX1 DFF_1348_Q_reg ( .D(n1701), .SI(n8351), .SE(n9389), .CLK(n9591), .Q(
        n8350), .QN(n8853) );
  SDFFX1 DFF_1349_Q_reg ( .D(n1702), .SI(n8350), .SE(n9389), .CLK(n9591), .Q(
        n8349), .QN(n8852) );
  SDFFX1 DFF_1350_Q_reg ( .D(n1703), .SI(n8349), .SE(n9389), .CLK(n9591), .Q(
        n8348), .QN(n8851) );
  SDFFX1 DFF_1351_Q_reg ( .D(n1704), .SI(n8348), .SE(n9389), .CLK(n9591), .Q(
        n8347), .QN(n8850) );
  SDFFX1 DFF_1352_Q_reg ( .D(n1705), .SI(n8347), .SE(n9389), .CLK(n9591), .Q(
        n8346), .QN(n8849) );
  SDFFX1 DFF_1353_Q_reg ( .D(n1706), .SI(n8346), .SE(n9389), .CLK(n9591), .Q(
        test_so78), .QN(n9061) );
  SDFFX1 DFF_1354_Q_reg ( .D(n1707), .SI(test_si79), .SE(n9389), .CLK(n9591), 
        .Q(n8343), .QN(n8848) );
  SDFFX1 DFF_1355_Q_reg ( .D(n1708), .SI(n8343), .SE(n9389), .CLK(n9591), .Q(
        n8342), .QN(n8847) );
  SDFFX1 DFF_1356_Q_reg ( .D(n1709), .SI(n8342), .SE(n9389), .CLK(n9591), .Q(
        n8341), .QN(n8846) );
  SDFFX1 DFF_1357_Q_reg ( .D(n1710), .SI(n8341), .SE(n9389), .CLK(n9591), .Q(
        n8340), .QN(n8845) );
  SDFFX1 DFF_1358_Q_reg ( .D(n1711), .SI(n8340), .SE(n9389), .CLK(n9591), .Q(
        n8339), .QN(n8844) );
  SDFFX1 DFF_1359_Q_reg ( .D(n1712), .SI(n8339), .SE(n9389), .CLK(n9591), .Q(
        n8338), .QN(n8843) );
  SDFFX1 DFF_1360_Q_reg ( .D(n1713), .SI(n8338), .SE(n9390), .CLK(n9590), .Q(
        n8337), .QN(n8842) );
  SDFFX1 DFF_1361_Q_reg ( .D(n1714), .SI(n8337), .SE(n9390), .CLK(n9590), .Q(
        n8336), .QN(n8841) );
  SDFFX1 DFF_1362_Q_reg ( .D(n1715), .SI(n8336), .SE(n9390), .CLK(n9590), .Q(
        n8335), .QN(n8840) );
  SDFFX1 DFF_1363_Q_reg ( .D(n1716), .SI(n8335), .SE(n9390), .CLK(n9590), .Q(
        n8334), .QN(n8839) );
  SDFFX1 DFF_1364_Q_reg ( .D(n1717), .SI(n8334), .SE(n9390), .CLK(n9590), .Q(
        n8333), .QN(n8838) );
  SDFFX1 DFF_1365_Q_reg ( .D(n1718), .SI(n8333), .SE(n9390), .CLK(n9590), .Q(
        n8332), .QN(n8837) );
  SDFFX1 DFF_1366_Q_reg ( .D(n1719), .SI(n8332), .SE(n9390), .CLK(n9590), .Q(
        n8331), .QN(n8836) );
  SDFFX1 DFF_1367_Q_reg ( .D(n1720), .SI(n8331), .SE(n9390), .CLK(n9590), .Q(
        n8330), .QN(n8835) );
  SDFFX1 DFF_1368_Q_reg ( .D(n1721), .SI(n8330), .SE(n9390), .CLK(n9590), .Q(
        n8329), .QN(n8834) );
  SDFFX1 DFF_1369_Q_reg ( .D(n1722), .SI(n8329), .SE(n9390), .CLK(n9590), .Q(
        n8328), .QN(n8833) );
  SDFFX1 DFF_1370_Q_reg ( .D(n1723), .SI(n8328), .SE(n9390), .CLK(n9590), .Q(
        test_so79), .QN(n9060) );
  SDFFX1 DFF_1371_Q_reg ( .D(n1724), .SI(test_si80), .SE(n9390), .CLK(n9590), 
        .Q(n8325), .QN(n8832) );
  SDFFX1 DFF_1372_Q_reg ( .D(n1725), .SI(n8325), .SE(n9391), .CLK(n9589), .Q(
        n8324), .QN(n8831) );
  SDFFX1 DFF_1373_Q_reg ( .D(n1726), .SI(n8324), .SE(n9391), .CLK(n9589), .Q(
        n8323), .QN(n8830) );
  SDFFX1 DFF_1374_Q_reg ( .D(n1727), .SI(n8323), .SE(n9391), .CLK(n9589), .Q(
        n8322), .QN(n8829) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n9391), .CLK(n9589), .Q(
        n8321), .QN(n8828) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n9388), .CLK(n9592), .Q(
        n8320), .QN(n16118) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n9388), .CLK(n9592), .Q(
        n8319), .QN(n16119) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n9388), .CLK(n9592), .Q(
        n8318), .QN(n16120) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n9388), .CLK(n9592), .Q(
        n8317), .QN(n16121) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n9388), .CLK(n9592), .Q(
        n8316), .QN(n16122) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n9387), .CLK(n9593), .Q(
        n8315), .QN(n16123) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n9387), .CLK(n9593), .Q(
        n8314), .QN(n16124) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n9387), .CLK(n9593), .Q(
        n8313), .QN(n16125) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n9387), .CLK(n9593), .Q(
        n8312), .QN(n16126) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n9387), .CLK(n9593), .Q(
        n8311), .QN(n16127) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n9387), .CLK(n9593), .Q(
        n8310), .QN(n16128) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n9359), .CLK(n9621), .Q(
        test_so80), .QN(n8819) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n9386), .CLK(n9594), 
        .Q(n8307), .QN(n16129) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n9386), .CLK(n9594), .Q(
        n8306), .QN(n16130) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n9386), .CLK(n9594), .Q(
        n8305), .QN(n16131) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n9385), .CLK(n9595), .Q(
        n8304), .QN(n16132) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n9385), .CLK(n9595), .Q(
        WX9728), .QN(n7912) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n9385), .CLK(n9595), 
        .Q(WX9730), .QN(n7910) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n9385), .CLK(n9595), 
        .Q(WX9732), .QN(n7908) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n9385), .CLK(n9595), 
        .Q(WX9734), .QN(n7906) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n9384), .CLK(n9596), 
        .Q(WX9736), .QN(n7904) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n9384), .CLK(n9596), 
        .Q(WX9738), .QN(n7902) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n9384), .CLK(n9596), 
        .Q(WX9740), .QN(n7900) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n9383), .CLK(n9597), 
        .Q(WX9742), .QN(n7898) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n9383), .CLK(n9597), 
        .Q(WX9744), .QN(n7896) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n9383), .CLK(n9597), 
        .Q(WX9746), .QN(n7894) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n9382), .CLK(n9598), 
        .Q(WX9748), .QN(n7892) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n9382), .CLK(n9598), 
        .Q(WX9750), .QN(n7890) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n9382), .CLK(n9598), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n9381), .CLK(n9599), 
        .Q(WX9754), .QN(n7887) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n9381), .CLK(n9599), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n9381), .CLK(n9599), 
        .Q(WX9758), .QN(n7883) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n9388), .CLK(n9592), 
        .Q(WX9760), .QN(n7613) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n9388), .CLK(n9592), 
        .Q(WX9762), .QN(n7681) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n9388), .CLK(n9592), 
        .Q(WX9764), .QN(n7679) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n9388), .CLK(n9592), 
        .Q(WX9766), .QN(n7677) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n9387), .CLK(n9593), 
        .Q(WX9768), .QN(n7675) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n9387), .CLK(n9593), 
        .Q(WX9770), .QN(n7673) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n9387), .CLK(n9593), 
        .Q(WX9772), .QN(n7671) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n9387), .CLK(n9593), 
        .Q(WX9774), .QN(n7669) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n9387), .CLK(n9593), 
        .Q(WX9776), .QN(n7667) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n9387), .CLK(n9593), 
        .Q(WX9778), .QN(n7665) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n9386), .CLK(n9594), 
        .Q(WX9780), .QN(n7663) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n9386), .CLK(n9594), 
        .Q(WX9782), .QN(n7661) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n9386), .CLK(n9594), 
        .Q(WX9784), .QN(n7659) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n9386), .CLK(n9594), 
        .Q(test_so82), .QN(n8806) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n9386), .CLK(n9594), 
        .Q(WX9788), .QN(n7656) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n9386), .CLK(n9594), 
        .Q(WX9790), .QN(n7655) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n9385), .CLK(n9595), 
        .Q(WX9792) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n9385), .CLK(n9595), 
        .Q(WX9794), .QN(n3591) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n9385), .CLK(n9595), 
        .Q(WX9796) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n9384), .CLK(n9596), 
        .Q(WX9798) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n9384), .CLK(n9596), 
        .Q(WX9800) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n9384), .CLK(n9596), 
        .Q(WX9802) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n9383), .CLK(n9597), 
        .Q(WX9804) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n9383), .CLK(n9597), 
        .Q(WX9806) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n9383), .CLK(n9597), 
        .Q(WX9808) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n9382), .CLK(n9598), 
        .Q(WX9810) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n9382), .CLK(n9598), 
        .Q(WX9812) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n9382), .CLK(n9598), 
        .Q(WX9814) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n9381), .CLK(n9599), 
        .Q(WX9816), .QN(n3569) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n9381), .CLK(n9599), 
        .Q(WX9818) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n9381), .CLK(n9599), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n9380), .CLK(n9600), 
        .Q(WX9822) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n9380), .CLK(n9600), 
        .Q(WX9824), .QN(n7614) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n9380), .CLK(n9600), 
        .Q(WX9826), .QN(n7682) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n9380), .CLK(n9600), 
        .Q(WX9828), .QN(n7680) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n9380), .CLK(n9600), 
        .Q(WX9830), .QN(n7678) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n9380), .CLK(n9600), 
        .Q(WX9832), .QN(n7676) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n9379), .CLK(n9601), 
        .Q(WX9834), .QN(n7674) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n9379), .CLK(n9601), 
        .Q(WX9836), .QN(n7672) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n9379), .CLK(n9601), 
        .Q(WX9838), .QN(n7670) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n9379), .CLK(n9601), 
        .Q(WX9840), .QN(n7668) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n9379), .CLK(n9601), 
        .Q(WX9842), .QN(n7666) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n9379), .CLK(n9601), 
        .Q(WX9844), .QN(n7664) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n9378), .CLK(n9602), 
        .Q(WX9846), .QN(n7662) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n9378), .CLK(n9602), 
        .Q(WX9848), .QN(n7660) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n9386), .CLK(n9594), 
        .Q(WX9850), .QN(n7658) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n9386), .CLK(n9594), 
        .Q(WX9852), .QN(n7657) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n9386), .CLK(n9594), 
        .Q(test_so84), .QN(n8805) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n9385), .CLK(n9595), 
        .Q(WX9856), .QN(n7913) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n9385), .CLK(n9595), 
        .Q(WX9858), .QN(n7911) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n9385), .CLK(n9595), 
        .Q(WX9860), .QN(n7909) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n9384), .CLK(n9596), 
        .Q(WX9862), .QN(n7907) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n9384), .CLK(n9596), 
        .Q(WX9864), .QN(n7905) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n9384), .CLK(n9596), 
        .Q(WX9866), .QN(n7903) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n9383), .CLK(n9597), 
        .Q(WX9868), .QN(n7901) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n9383), .CLK(n9597), 
        .Q(WX9870), .QN(n7899) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n9383), .CLK(n9597), 
        .Q(WX9872), .QN(n7897) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n9382), .CLK(n9598), 
        .Q(WX9874), .QN(n7895) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n9382), .CLK(n9598), 
        .Q(WX9876), .QN(n7893) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n9382), .CLK(n9598), 
        .Q(WX9878), .QN(n7891) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n9381), .CLK(n9599), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n9381), .CLK(n9599), 
        .Q(WX9882), .QN(n7888) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n9381), .CLK(n9599), 
        .Q(WX9884), .QN(n7886) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n9380), .CLK(n9600), 
        .Q(WX9886), .QN(n7884) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n9380), .CLK(n9600), 
        .Q(test_so85), .QN(n8804) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n9380), .CLK(n9600), 
        .Q(WX9890), .QN(n8159) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n9380), .CLK(n9600), 
        .Q(WX9892), .QN(n8160) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n9380), .CLK(n9600), 
        .Q(WX9894), .QN(n8161) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n9379), .CLK(n9601), 
        .Q(WX9896), .QN(n8162) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n9379), .CLK(n9601), 
        .Q(WX9898), .QN(n8163) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n9379), .CLK(n9601), 
        .Q(WX9900), .QN(n8164) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n9379), .CLK(n9601), 
        .Q(WX9902), .QN(n8165) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n9379), .CLK(n9601), 
        .Q(WX9904), .QN(n8166) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n9379), .CLK(n9601), 
        .Q(WX9906), .QN(n8167) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n9378), .CLK(n9602), 
        .Q(WX9908), .QN(n8168) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n9378), .CLK(n9602), 
        .Q(WX9910), .QN(n8169) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n9378), .CLK(n9602), 
        .Q(WX9912), .QN(n8170) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n9378), .CLK(n9602), 
        .Q(WX9914), .QN(n8171) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n9378), .CLK(n9602), 
        .Q(WX9916), .QN(n8172) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n9378), .CLK(n9602), 
        .Q(WX9918), .QN(n8107) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n9378), .CLK(n9602), 
        .Q(WX9920), .QN(n8173) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n9378), .CLK(n9602), 
        .Q(test_so86), .QN(n8794) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n9385), .CLK(n9595), 
        .Q(WX9924), .QN(n8174) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n9384), .CLK(n9596), 
        .Q(WX9926), .QN(n8175) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n9384), .CLK(n9596), 
        .Q(WX9928), .QN(n8108) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n9384), .CLK(n9596), 
        .Q(WX9930), .QN(n8176) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n9383), .CLK(n9597), 
        .Q(WX9932), .QN(n8177) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n9383), .CLK(n9597), 
        .Q(WX9934), .QN(n8178) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n9383), .CLK(n9597), 
        .Q(WX9936), .QN(n8179) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n9382), .CLK(n9598), 
        .Q(WX9938), .QN(n8180) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n9382), .CLK(n9598), 
        .Q(WX9940), .QN(n8181) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n9382), .CLK(n9598), 
        .Q(WX9942), .QN(n8109) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n9381), .CLK(n9599), 
        .Q(WX9944), .QN(n8182) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n9381), .CLK(n9599), 
        .Q(WX9946), .QN(n8183) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n9381), .CLK(n9599), 
        .Q(WX9948), .QN(n8184) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n9380), .CLK(n9600), 
        .Q(WX9950), .QN(n8126) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n9361), .CLK(n9619), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n9360), .CLK(
        n9620), .Q(test_so87) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n9360), .CLK(n9620), 
        .Q(CRC_OUT_2_3) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_10) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n9360), .CLK(
        n9620), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n9359), .CLK(
        n9621), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n9359), .CLK(
        n9621), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n9359), .CLK(
        n9621), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n9359), .CLK(
        n9621), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n9359), .CLK(
        n9621), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n9359), .CLK(
        n9621), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n9378), .CLK(
        n9602), .Q(test_so88) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n9378), .CLK(n9602), 
        .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n9377), .CLK(
        n9603), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n1938), .SI(CRC_OUT_2_31), .SE(n9377), .CLK(n9603), .Q(WX10829) );
  SDFFX1 DFF_1537_Q_reg ( .D(n1939), .SI(WX10829), .SE(n9374), .CLK(n9606), 
        .Q(n8295), .QN(n9059) );
  SDFFX1 DFF_1538_Q_reg ( .D(n1940), .SI(n8295), .SE(n9374), .CLK(n9606), .Q(
        n8294), .QN(n9058) );
  SDFFX1 DFF_1539_Q_reg ( .D(n1941), .SI(n8294), .SE(n9374), .CLK(n9606), .Q(
        n8293), .QN(n9057) );
  SDFFX1 DFF_1540_Q_reg ( .D(n1942), .SI(n8293), .SE(n9374), .CLK(n9606), .Q(
        test_so89), .QN(n9075) );
  SDFFX1 DFF_1541_Q_reg ( .D(n1943), .SI(test_si90), .SE(n9374), .CLK(n9606), 
        .Q(n8290), .QN(n9056) );
  SDFFX1 DFF_1542_Q_reg ( .D(n1944), .SI(n8290), .SE(n9374), .CLK(n9606), .Q(
        n8289), .QN(n9055) );
  SDFFX1 DFF_1543_Q_reg ( .D(n1945), .SI(n8289), .SE(n9374), .CLK(n9606), .Q(
        n8288), .QN(n9054) );
  SDFFX1 DFF_1544_Q_reg ( .D(n1946), .SI(n8288), .SE(n9375), .CLK(n9605), .Q(
        n8287), .QN(n9053) );
  SDFFX1 DFF_1545_Q_reg ( .D(n1947), .SI(n8287), .SE(n9375), .CLK(n9605), .Q(
        n8286), .QN(n9052) );
  SDFFX1 DFF_1546_Q_reg ( .D(n1948), .SI(n8286), .SE(n9375), .CLK(n9605), .Q(
        n8285), .QN(n9051) );
  SDFFX1 DFF_1547_Q_reg ( .D(n1949), .SI(n8285), .SE(n9375), .CLK(n9605), .Q(
        n8284), .QN(n9050) );
  SDFFX1 DFF_1548_Q_reg ( .D(n1950), .SI(n8284), .SE(n9375), .CLK(n9605), .Q(
        n8283), .QN(n9049) );
  SDFFX1 DFF_1549_Q_reg ( .D(n1951), .SI(n8283), .SE(n9375), .CLK(n9605), .Q(
        n8282), .QN(n9048) );
  SDFFX1 DFF_1550_Q_reg ( .D(n1952), .SI(n8282), .SE(n9375), .CLK(n9605), .Q(
        n8281), .QN(n9047) );
  SDFFX1 DFF_1551_Q_reg ( .D(n1953), .SI(n8281), .SE(n9375), .CLK(n9605), .Q(
        n8280), .QN(n9046) );
  SDFFX1 DFF_1552_Q_reg ( .D(n1954), .SI(n8280), .SE(n9375), .CLK(n9605), .Q(
        n8279), .QN(n9045) );
  SDFFX1 DFF_1553_Q_reg ( .D(n1955), .SI(n8279), .SE(n9375), .CLK(n9605), .Q(
        n8278), .QN(n9044) );
  SDFFX1 DFF_1554_Q_reg ( .D(n1956), .SI(n8278), .SE(n9375), .CLK(n9605), .Q(
        n8277), .QN(n9043) );
  SDFFX1 DFF_1555_Q_reg ( .D(n1957), .SI(n8277), .SE(n9375), .CLK(n9605), .Q(
        n8276), .QN(n9042) );
  SDFFX1 DFF_1556_Q_reg ( .D(n1958), .SI(n8276), .SE(n9376), .CLK(n9604), .Q(
        n8275), .QN(n9041) );
  SDFFX1 DFF_1557_Q_reg ( .D(n1959), .SI(n8275), .SE(n9376), .CLK(n9604), .Q(
        test_so90), .QN(n9074) );
  SDFFX1 DFF_1558_Q_reg ( .D(n1960), .SI(test_si91), .SE(n9376), .CLK(n9604), 
        .Q(n8272), .QN(n9040) );
  SDFFX1 DFF_1559_Q_reg ( .D(n1961), .SI(n8272), .SE(n9376), .CLK(n9604), .Q(
        n8271), .QN(n9039) );
  SDFFX1 DFF_1560_Q_reg ( .D(n1962), .SI(n8271), .SE(n9376), .CLK(n9604), .Q(
        n8270), .QN(n9038) );
  SDFFX1 DFF_1561_Q_reg ( .D(n1963), .SI(n8270), .SE(n9376), .CLK(n9604), .Q(
        n8269), .QN(n9037) );
  SDFFX1 DFF_1562_Q_reg ( .D(n1964), .SI(n8269), .SE(n9376), .CLK(n9604), .Q(
        n8268), .QN(n9036) );
  SDFFX1 DFF_1563_Q_reg ( .D(n1965), .SI(n8268), .SE(n9376), .CLK(n9604), .Q(
        n8267), .QN(n9035) );
  SDFFX1 DFF_1564_Q_reg ( .D(n1966), .SI(n8267), .SE(n9376), .CLK(n9604), .Q(
        n8266), .QN(n9034) );
  SDFFX1 DFF_1565_Q_reg ( .D(n1967), .SI(n8266), .SE(n9376), .CLK(n9604), .Q(
        n8265), .QN(n9033) );
  SDFFX1 DFF_1566_Q_reg ( .D(n1968), .SI(n8265), .SE(n9376), .CLK(n9604), .Q(
        n8264), .QN(n9032) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n9376), .CLK(n9604), 
        .Q(n8263), .QN(n9031) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n9374), .CLK(n9606), 
        .Q(n8262), .QN(n16133) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n9374), .CLK(n9606), 
        .Q(n8261), .QN(n16134) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n9374), .CLK(n9606), 
        .Q(n8260), .QN(n16135) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n9373), .CLK(n9607), 
        .Q(n8259), .QN(n16136) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n9373), .CLK(n9607), 
        .Q(n8258), .QN(n16137) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n9373), .CLK(n9607), 
        .Q(n8257), .QN(n16138) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n9373), .CLK(n9607), 
        .Q(test_so91), .QN(n8825) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n9373), .CLK(n9607), 
        .Q(n8254), .QN(n16139) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n9373), .CLK(n9607), 
        .Q(n8253), .QN(n16140) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n9372), .CLK(n9608), 
        .Q(n8252), .QN(n16141) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n9372), .CLK(n9608), 
        .Q(n8251), .QN(n16142) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n9372), .CLK(n9608), 
        .Q(n8250), .QN(n16143) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n9371), .CLK(n9609), 
        .Q(n8249), .QN(n16144) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n9371), .CLK(n9609), 
        .Q(n8248), .QN(n16145) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n9371), .CLK(n9609), 
        .Q(n8247), .QN(n16146) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n9371), .CLK(n9609), 
        .Q(n8246), .QN(n16147) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n9370), .CLK(n9610), 
        .Q(WX11021), .QN(n7881) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n9370), .CLK(n9610), 
        .Q(WX11023), .QN(n7879) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n9370), .CLK(n9610), 
        .Q(WX11025), .QN(n7877) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n9369), .CLK(n9611), 
        .Q(WX11027), .QN(n7875) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n9369), .CLK(n9611), 
        .Q(WX11029), .QN(n7873) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n9369), .CLK(n9611), 
        .Q(WX11031), .QN(n7871) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n9368), .CLK(n9612), 
        .Q(WX11033), .QN(n7869) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n9368), .CLK(n9612), 
        .Q(test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n9367), .CLK(n9613), 
        .Q(WX11037), .QN(n7866) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n9367), .CLK(n9613), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n9367), .CLK(n9613), 
        .Q(WX11041), .QN(n7862) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n9367), .CLK(n9613), 
        .Q(WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n9366), .CLK(n9614), 
        .Q(WX11045), .QN(n7859) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n9366), .CLK(n9614), 
        .Q(WX11047), .QN(n7857) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n9366), .CLK(n9614), 
        .Q(WX11049), .QN(n7855) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n9365), .CLK(n9615), 
        .Q(WX11051), .QN(n7853) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n9374), .CLK(n9606), 
        .Q(WX11053), .QN(n7611) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n9374), .CLK(n9606), 
        .Q(WX11055), .QN(n7653) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n9373), .CLK(n9607), 
        .Q(WX11057), .QN(n7651) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n9373), .CLK(n9607), 
        .Q(WX11059), .QN(n7649) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n9373), .CLK(n9607), 
        .Q(WX11061), .QN(n7647) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n9373), .CLK(n9607), 
        .Q(WX11063), .QN(n7645) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n9373), .CLK(n9607), 
        .Q(WX11065), .QN(n7643) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n9373), .CLK(n9607), 
        .Q(WX11067), .QN(n7641) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n9372), .CLK(n9608), 
        .Q(test_so93), .QN(n8818) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n9372), .CLK(n9608), 
        .Q(WX11071), .QN(n7638) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n9372), .CLK(n9608), 
        .Q(WX11073), .QN(n7637) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n9372), .CLK(n9608), 
        .Q(WX11075), .QN(n7635) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n9372), .CLK(n9608), 
        .Q(WX11077), .QN(n7633) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n9371), .CLK(n9609), 
        .Q(WX11079), .QN(n7631) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n9371), .CLK(n9609), 
        .Q(WX11081), .QN(n7629) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n9371), .CLK(n9609), 
        .Q(WX11083), .QN(n7627) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n9370), .CLK(n9610), 
        .Q(WX11085) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n9370), .CLK(n9610), 
        .Q(WX11087) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n9370), .CLK(n9610), 
        .Q(WX11089) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n9369), .CLK(n9611), 
        .Q(WX11091) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n9369), .CLK(n9611), 
        .Q(WX11093) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n9369), .CLK(n9611), 
        .Q(WX11095) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n9368), .CLK(n9612), 
        .Q(WX11097) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n9368), .CLK(n9612), 
        .Q(WX11099), .QN(n3547) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n9368), .CLK(n9612), 
        .Q(WX11101) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n9367), .CLK(n9613), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n9367), .CLK(n9613), 
        .Q(WX11105) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n9367), .CLK(n9613), 
        .Q(WX11107), .QN(n3539) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n9366), .CLK(n9614), 
        .Q(WX11109) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n9366), .CLK(n9614), 
        .Q(WX11111), .QN(n3535) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n9366), .CLK(n9614), 
        .Q(WX11113) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n9365), .CLK(n9615), 
        .Q(WX11115) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n9365), .CLK(n9615), 
        .Q(WX11117), .QN(n7612) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n9365), .CLK(n9615), 
        .Q(WX11119), .QN(n7654) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n9365), .CLK(n9615), 
        .Q(WX11121), .QN(n7652) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n9364), .CLK(n9616), 
        .Q(WX11123), .QN(n7650) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n9364), .CLK(n9616), 
        .Q(WX11125), .QN(n7648) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n9364), .CLK(n9616), 
        .Q(WX11127), .QN(n7646) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n9364), .CLK(n9616), 
        .Q(WX11129), .QN(n7644) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n9364), .CLK(n9616), 
        .Q(WX11131), .QN(n7642) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n9372), .CLK(n9608), 
        .Q(WX11133), .QN(n7640) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n9372), .CLK(n9608), 
        .Q(WX11135), .QN(n7639) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n9372), .CLK(n9608), 
        .Q(test_so95), .QN(n8817) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n9372), .CLK(n9608), 
        .Q(WX11139), .QN(n7636) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n9371), .CLK(n9609), 
        .Q(WX11141), .QN(n7634) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n9371), .CLK(n9609), 
        .Q(WX11143), .QN(n7632) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n9371), .CLK(n9609), 
        .Q(WX11145), .QN(n7630) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n9370), .CLK(n9610), 
        .Q(WX11147), .QN(n7628) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n9370), .CLK(n9610), 
        .Q(WX11149), .QN(n7882) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n9370), .CLK(n9610), 
        .Q(WX11151), .QN(n7880) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n9369), .CLK(n9611), 
        .Q(WX11153), .QN(n7878) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n9369), .CLK(n9611), 
        .Q(WX11155), .QN(n7876) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155), .SE(n9369), .CLK(n9611), 
        .Q(WX11157), .QN(n7874) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(n9368), .CLK(n9612), 
        .Q(WX11159), .QN(n7872) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(n9368), .CLK(n9612), 
        .Q(WX11161), .QN(n7870) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(n9368), .CLK(n9612), 
        .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(n9368), .CLK(n9612), 
        .Q(WX11165), .QN(n7867) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(n9367), .CLK(n9613), 
        .Q(WX11167), .QN(n7865) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(n9367), .CLK(n9613), 
        .Q(WX11169), .QN(n7863) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(n9366), .CLK(n9614), 
        .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n9366), .CLK(n9614), 
        .Q(WX11173), .QN(n7860) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n9366), .CLK(n9614), 
        .Q(WX11175), .QN(n7858) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n9365), .CLK(n9615), 
        .Q(WX11177), .QN(n7856) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n9365), .CLK(n9615), 
        .Q(WX11179), .QN(n7854) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n9365), .CLK(n9615), 
        .Q(WX11181), .QN(n8133) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n9365), .CLK(n9615), 
        .Q(WX11183), .QN(n8134) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n9365), .CLK(n9615), 
        .Q(WX11185), .QN(n8135) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n9364), .CLK(n9616), 
        .Q(WX11187), .QN(n8136) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n9364), .CLK(n9616), 
        .Q(WX11189), .QN(n8137) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n9364), .CLK(n9616), 
        .Q(WX11191), .QN(n8138) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n9364), .CLK(n9616), 
        .Q(WX11193), .QN(n8139) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n9364), .CLK(n9616), 
        .Q(WX11195), .QN(n8140) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n9364), .CLK(n9616), 
        .Q(WX11197), .QN(n8141) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n9364), .CLK(n9616), 
        .Q(WX11199), .QN(n8142) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n9363), .CLK(n9617), 
        .Q(WX11201), .QN(n8143) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n9363), .CLK(n9617), 
        .Q(WX11203), .QN(n8144) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n9363), .CLK(n9617), 
        .Q(test_so97), .QN(n8803) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n9371), .CLK(n9609), 
        .Q(WX11207), .QN(n8145) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n9371), .CLK(n9609), 
        .Q(WX11209), .QN(n8146) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n9370), .CLK(n9610), 
        .Q(WX11211), .QN(n8104) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n9370), .CLK(n9610), 
        .Q(WX11213) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n9370), .CLK(n9610), 
        .Q(WX11215), .QN(n8148) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n9369), .CLK(n9611), 
        .Q(WX11217), .QN(n8149) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n9369), .CLK(n9611), 
        .Q(WX11219), .QN(n8150) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n9369), .CLK(n9611), 
        .Q(WX11221), .QN(n8105) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n9368), .CLK(n9612), 
        .Q(WX11223), .QN(n8151) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n9368), .CLK(n9612), 
        .Q(WX11225), .QN(n8152) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n9368), .CLK(n9612), 
        .Q(WX11227), .QN(n8153) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n9367), .CLK(n9613), 
        .Q(WX11229), .QN(n8154) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n9367), .CLK(n9613), 
        .Q(WX11231), .QN(n8155) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n9367), .CLK(n9613), 
        .Q(WX11233), .QN(n8156) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n9366), .CLK(n9614), 
        .Q(WX11235), .QN(n8106) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n9366), .CLK(n9614), 
        .Q(WX11237), .QN(n8157) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n9366), .CLK(n9614), 
        .Q(test_so98), .QN(n8793) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n9365), .CLK(n9615), 
        .Q(WX11241), .QN(n8158) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n9365), .CLK(n9615), 
        .Q(WX11243), .QN(n8125) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n9363), .CLK(n9617), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_3) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_10) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n9362), .CLK(
        n9618), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n9361), .CLK(
        n9619), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n9361), .CLK(n9619), .Q(CRC_OUT_1_15) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n9361), .CLK(
        n9619), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n9363), .CLK(
        n9617), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n9363), .CLK(
        n9617), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n9363), .CLK(
        n9617), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n9363), .CLK(
        n9617), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n9363), .CLK(
        n9617), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n9363), .CLK(
        n9617), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n9363), .CLK(
        n9617), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n9363), .CLK(
        n9617), .Q(test_so100), .QN(n8789) );
  NOR2X0 Trojan1 ( .IN1(WX3442), .IN2(WX5974), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(WX806), .IN2(WX782), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(WX11632), .IN2(n507), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(WX5964), .IN2(WX3324), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(WX8634), .IN2(WX3330), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n519), .IN2(n511), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(WX862), .IN2(WX7227), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(WX11616), .IN2(n1955), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(n9490), .Q(
        Tj_Trigger) );
  NAND3X4 TrojanPayload1 ( .IN1(WX547), .IN2(Tj_Trigger), .IN3(Stage4), .QN(
        Stage1_1) );
  INVX8 TrojanPayload2 ( .INP(Stage1_1), .ZN(Stage1_2) );
  INVX8 TrojanPayload3 ( .INP(Stage1_2), .ZN(Stage1_3) );
  INVX8 TrojanPayload4 ( .INP(Stage1_3), .ZN(Stage1_4) );
  INVX8 TrojanPayload5 ( .INP(Stage1_4), .ZN(Stage1) );
  MUX21X2 TrojanPayload6 ( .IN1(WX544), .IN2(Stage1), .S(1'b0), .Q(Stage2_i)
         );
  INVX8 TrojanPayload7 ( .INP(Stage2_i), .ZN(Stage2_7) );
  INVX8 TrojanPayload8 ( .INP(Stage2_7), .ZN(Stage2_8) );
  INVX8 TrojanPayload9 ( .INP(Stage2_8), .ZN(Stage2_9) );
  INVX8 TrojanPayload10 ( .INP(Stage2_9), .ZN(Stage2_10) );
  INVX8 TrojanPayload11 ( .INP(Stage2_10), .ZN(Stage2) );
  MUX21X2 TrojanPayload12 ( .IN1(WX706), .IN2(Stage2), .S(1'b0), .Q(Stage3_i)
         );
  INVX8 TrojanPayload13 ( .INP(Stage3_i), .ZN(Stage3_12) );
  INVX8 TrojanPayload14 ( .INP(Stage3_12), .ZN(Stage3_13) );
  INVX8 TrojanPayload15 ( .INP(Stage3_13), .ZN(Stage3_14) );
  INVX8 TrojanPayload16 ( .INP(Stage3_14), .ZN(Stage3_15) );
  INVX8 TrojanPayload17 ( .INP(Stage3_15) );
  MUX21X2 TrojanPayload18 ( .IN1(n3467), .IN2(1'b0), .S(1'b0), .Q(Stage4_i) );
  INVX8 TrojanPayload19 ( .INP(Stage4_i), .ZN(Stage4_17) );
  INVX8 TrojanPayload20 ( .INP(Stage4_17), .ZN(Stage4_18) );
  INVX8 TrojanPayload21 ( .INP(Stage4_18), .ZN(Stage4_19) );
  INVX8 TrojanPayload22 ( .INP(Stage4_19), .ZN(Stage4_20) );
  INVX8 TrojanPayload23 ( .INP(Stage4_20), .ZN(Stage4_21) );
  INVX8 TrojanPayload24 ( .INP(Stage4_21), .ZN(Stage4) );
  INVX0 U8973 ( .INP(n9791), .ZN(n9076) );
  INVX0 U8974 ( .INP(n9076), .ZN(n9077) );
  INVX0 U8975 ( .INP(n9076), .ZN(n9078) );
  INVX0 U8976 ( .INP(n9076), .ZN(n9079) );
  INVX0 U8977 ( .INP(n9790), .ZN(n9080) );
  INVX0 U8978 ( .INP(n9080), .ZN(n9081) );
  INVX0 U8979 ( .INP(n9080), .ZN(n9082) );
  INVX0 U8980 ( .INP(n9080), .ZN(n9083) );
  NBUFFX2 U8981 ( .INP(n9244), .Z(n9227) );
  NBUFFX2 U8982 ( .INP(n9244), .Z(n9228) );
  NBUFFX2 U8983 ( .INP(n9244), .Z(n9230) );
  NBUFFX2 U8984 ( .INP(n9244), .Z(n9229) );
  NBUFFX2 U8985 ( .INP(n9245), .Z(n9223) );
  NBUFFX2 U8986 ( .INP(n9244), .Z(n9231) );
  NBUFFX2 U8987 ( .INP(n9243), .Z(n9232) );
  NBUFFX2 U8988 ( .INP(n9243), .Z(n9233) );
  NBUFFX2 U8989 ( .INP(n9243), .Z(n9234) );
  NBUFFX2 U8990 ( .INP(n9243), .Z(n9236) );
  NBUFFX2 U8991 ( .INP(n9242), .Z(n9237) );
  NBUFFX2 U8992 ( .INP(n9242), .Z(n9238) );
  NBUFFX2 U8993 ( .INP(n9242), .Z(n9239) );
  NBUFFX2 U8994 ( .INP(n9242), .Z(n9240) );
  NBUFFX2 U8995 ( .INP(n9245), .Z(n9226) );
  NBUFFX2 U8996 ( .INP(n9245), .Z(n9225) );
  NBUFFX2 U8997 ( .INP(n9245), .Z(n9224) );
  NBUFFX2 U8998 ( .INP(n9243), .Z(n9235) );
  NBUFFX2 U8999 ( .INP(n9260), .Z(n9147) );
  NBUFFX2 U9000 ( .INP(n9261), .Z(n9146) );
  NBUFFX2 U9001 ( .INP(n9261), .Z(n9145) );
  NBUFFX2 U9002 ( .INP(n9261), .Z(n9144) );
  NBUFFX2 U9003 ( .INP(n9261), .Z(n9143) );
  NBUFFX2 U9004 ( .INP(n9261), .Z(n9142) );
  NBUFFX2 U9005 ( .INP(n9262), .Z(n9141) );
  NBUFFX2 U9006 ( .INP(n9262), .Z(n9139) );
  NBUFFX2 U9007 ( .INP(n9262), .Z(n9138) );
  NBUFFX2 U9008 ( .INP(n9262), .Z(n9137) );
  NBUFFX2 U9009 ( .INP(n9262), .Z(n9140) );
  NBUFFX2 U9010 ( .INP(n9259), .Z(n9152) );
  NBUFFX2 U9011 ( .INP(n9259), .Z(n9154) );
  NBUFFX2 U9012 ( .INP(n9259), .Z(n9153) );
  NBUFFX2 U9013 ( .INP(n9260), .Z(n9151) );
  NBUFFX2 U9014 ( .INP(n9260), .Z(n9150) );
  NBUFFX2 U9015 ( .INP(n9260), .Z(n9149) );
  NBUFFX2 U9016 ( .INP(n9260), .Z(n9148) );
  NBUFFX2 U9017 ( .INP(n9259), .Z(n9155) );
  NBUFFX2 U9018 ( .INP(n9258), .Z(n9157) );
  NBUFFX2 U9019 ( .INP(n9259), .Z(n9156) );
  NBUFFX2 U9020 ( .INP(n9257), .Z(n9163) );
  NBUFFX2 U9021 ( .INP(n9258), .Z(n9158) );
  NBUFFX2 U9022 ( .INP(n9258), .Z(n9159) );
  NBUFFX2 U9023 ( .INP(n9258), .Z(n9160) );
  NBUFFX2 U9024 ( .INP(n9258), .Z(n9161) );
  NBUFFX2 U9025 ( .INP(n9257), .Z(n9162) );
  NBUFFX2 U9026 ( .INP(n9251), .Z(n9195) );
  NBUFFX2 U9027 ( .INP(n9251), .Z(n9196) );
  NBUFFX2 U9028 ( .INP(n9250), .Z(n9198) );
  NBUFFX2 U9029 ( .INP(n9250), .Z(n9199) );
  NBUFFX2 U9030 ( .INP(n9250), .Z(n9200) );
  NBUFFX2 U9031 ( .INP(n9250), .Z(n9201) );
  NBUFFX2 U9032 ( .INP(n9249), .Z(n9202) );
  NBUFFX2 U9033 ( .INP(n9254), .Z(n9180) );
  NBUFFX2 U9034 ( .INP(n9254), .Z(n9181) );
  NBUFFX2 U9035 ( .INP(n9253), .Z(n9182) );
  NBUFFX2 U9036 ( .INP(n9253), .Z(n9183) );
  NBUFFX2 U9037 ( .INP(n9253), .Z(n9184) );
  NBUFFX2 U9038 ( .INP(n9253), .Z(n9185) );
  NBUFFX2 U9039 ( .INP(n9253), .Z(n9186) );
  NBUFFX2 U9040 ( .INP(n9252), .Z(n9187) );
  NBUFFX2 U9041 ( .INP(n9252), .Z(n9188) );
  NBUFFX2 U9042 ( .INP(n9252), .Z(n9189) );
  NBUFFX2 U9043 ( .INP(n9252), .Z(n9190) );
  NBUFFX2 U9044 ( .INP(n9246), .Z(n9221) );
  NBUFFX2 U9045 ( .INP(n9245), .Z(n9222) );
  NBUFFX2 U9046 ( .INP(n9246), .Z(n9220) );
  NBUFFX2 U9047 ( .INP(n9248), .Z(n9210) );
  NBUFFX2 U9048 ( .INP(n9248), .Z(n9209) );
  NBUFFX2 U9049 ( .INP(n9249), .Z(n9206) );
  NBUFFX2 U9050 ( .INP(n9249), .Z(n9205) );
  NBUFFX2 U9051 ( .INP(n9249), .Z(n9204) );
  NBUFFX2 U9052 ( .INP(n9248), .Z(n9207) );
  NBUFFX2 U9053 ( .INP(n9246), .Z(n9219) );
  NBUFFX2 U9054 ( .INP(n9246), .Z(n9218) );
  NBUFFX2 U9055 ( .INP(n9246), .Z(n9217) );
  NBUFFX2 U9056 ( .INP(n9247), .Z(n9216) );
  NBUFFX2 U9057 ( .INP(n9247), .Z(n9214) );
  NBUFFX2 U9058 ( .INP(n9247), .Z(n9213) );
  NBUFFX2 U9059 ( .INP(n9247), .Z(n9212) );
  NBUFFX2 U9060 ( .INP(n9248), .Z(n9211) );
  NBUFFX2 U9061 ( .INP(n9247), .Z(n9215) );
  NBUFFX2 U9062 ( .INP(n9248), .Z(n9208) );
  NBUFFX2 U9063 ( .INP(n9251), .Z(n9194) );
  NBUFFX2 U9064 ( .INP(n9256), .Z(n9170) );
  NBUFFX2 U9065 ( .INP(n9256), .Z(n9169) );
  NBUFFX2 U9066 ( .INP(n9256), .Z(n9167) );
  NBUFFX2 U9067 ( .INP(n9257), .Z(n9166) );
  NBUFFX2 U9068 ( .INP(n9257), .Z(n9165) );
  NBUFFX2 U9069 ( .INP(n9242), .Z(n9241) );
  NBUFFX2 U9070 ( .INP(n9256), .Z(n9168) );
  NBUFFX2 U9071 ( .INP(n9256), .Z(n9171) );
  NBUFFX2 U9072 ( .INP(n9255), .Z(n9172) );
  NBUFFX2 U9073 ( .INP(n9255), .Z(n9173) );
  NBUFFX2 U9074 ( .INP(n9255), .Z(n9174) );
  NBUFFX2 U9075 ( .INP(n9255), .Z(n9175) );
  NBUFFX2 U9076 ( .INP(n9255), .Z(n9176) );
  NBUFFX2 U9077 ( .INP(n9254), .Z(n9177) );
  NBUFFX2 U9078 ( .INP(n9254), .Z(n9178) );
  NBUFFX2 U9079 ( .INP(n9254), .Z(n9179) );
  NBUFFX2 U9080 ( .INP(n9249), .Z(n9203) );
  NBUFFX2 U9081 ( .INP(n9250), .Z(n9197) );
  NBUFFX2 U9082 ( .INP(n9252), .Z(n9191) );
  NBUFFX2 U9083 ( .INP(n9251), .Z(n9192) );
  NBUFFX2 U9084 ( .INP(n9251), .Z(n9193) );
  NBUFFX2 U9085 ( .INP(n9257), .Z(n9164) );
  NBUFFX2 U9086 ( .INP(n9264), .Z(n9272) );
  NBUFFX2 U9087 ( .INP(n9269), .Z(n9287) );
  NBUFFX2 U9088 ( .INP(n9264), .Z(n9273) );
  NBUFFX2 U9089 ( .INP(n9264), .Z(n9274) );
  NBUFFX2 U9090 ( .INP(n9265), .Z(n9275) );
  NBUFFX2 U9091 ( .INP(n9265), .Z(n9276) );
  NBUFFX2 U9092 ( .INP(n9266), .Z(n9280) );
  NBUFFX2 U9093 ( .INP(n9267), .Z(n9281) );
  NBUFFX2 U9094 ( .INP(n9267), .Z(n9282) );
  NBUFFX2 U9095 ( .INP(n9267), .Z(n9283) );
  NBUFFX2 U9096 ( .INP(n9268), .Z(n9284) );
  NBUFFX2 U9097 ( .INP(n9268), .Z(n9285) );
  NBUFFX2 U9098 ( .INP(n9268), .Z(n9286) );
  NBUFFX2 U9099 ( .INP(n9265), .Z(n9277) );
  NBUFFX2 U9100 ( .INP(n9266), .Z(n9278) );
  NBUFFX2 U9101 ( .INP(n9266), .Z(n9279) );
  NBUFFX2 U9102 ( .INP(n9315), .Z(n9313) );
  NBUFFX2 U9103 ( .INP(n9319), .Z(n9291) );
  NBUFFX2 U9104 ( .INP(n9319), .Z(n9292) );
  NBUFFX2 U9105 ( .INP(n9319), .Z(n9293) );
  NBUFFX2 U9106 ( .INP(n9319), .Z(n9294) );
  NBUFFX2 U9107 ( .INP(n9317), .Z(n9301) );
  NBUFFX2 U9108 ( .INP(n9317), .Z(n9303) );
  NBUFFX2 U9109 ( .INP(n9317), .Z(n9304) );
  NBUFFX2 U9110 ( .INP(n9316), .Z(n9305) );
  NBUFFX2 U9111 ( .INP(n9316), .Z(n9306) );
  NBUFFX2 U9112 ( .INP(n9316), .Z(n9307) );
  NBUFFX2 U9113 ( .INP(n9318), .Z(n9295) );
  NBUFFX2 U9114 ( .INP(n9318), .Z(n9296) );
  NBUFFX2 U9115 ( .INP(n9317), .Z(n9302) );
  NBUFFX2 U9116 ( .INP(n9318), .Z(n9297) );
  NBUFFX2 U9117 ( .INP(n9318), .Z(n9298) );
  NBUFFX2 U9118 ( .INP(n9318), .Z(n9299) );
  NBUFFX2 U9119 ( .INP(n9317), .Z(n9300) );
  NBUFFX2 U9120 ( .INP(n9316), .Z(n9309) );
  NBUFFX2 U9121 ( .INP(n9316), .Z(n9308) );
  NBUFFX2 U9122 ( .INP(n9315), .Z(n9310) );
  NBUFFX2 U9123 ( .INP(n9315), .Z(n9311) );
  NBUFFX2 U9124 ( .INP(n9315), .Z(n9312) );
  NBUFFX2 U9125 ( .INP(n9315), .Z(n9314) );
  NBUFFX2 U9126 ( .INP(n9665), .Z(n9496) );
  NBUFFX2 U9127 ( .INP(n9665), .Z(n9494) );
  NBUFFX2 U9128 ( .INP(n9665), .Z(n9495) );
  NBUFFX2 U9129 ( .INP(n9665), .Z(n9493) );
  NBUFFX2 U9130 ( .INP(n9640), .Z(n9618) );
  NBUFFX2 U9131 ( .INP(n9640), .Z(n9617) );
  NBUFFX2 U9132 ( .INP(n9641), .Z(n9616) );
  NBUFFX2 U9133 ( .INP(n9641), .Z(n9615) );
  NBUFFX2 U9134 ( .INP(n9641), .Z(n9614) );
  NBUFFX2 U9135 ( .INP(n9641), .Z(n9613) );
  NBUFFX2 U9136 ( .INP(n9641), .Z(n9612) );
  NBUFFX2 U9137 ( .INP(n9642), .Z(n9611) );
  NBUFFX2 U9138 ( .INP(n9642), .Z(n9610) );
  NBUFFX2 U9139 ( .INP(n9642), .Z(n9609) );
  NBUFFX2 U9140 ( .INP(n9642), .Z(n9608) );
  NBUFFX2 U9141 ( .INP(n9642), .Z(n9607) );
  NBUFFX2 U9142 ( .INP(n9643), .Z(n9604) );
  NBUFFX2 U9143 ( .INP(n9643), .Z(n9605) );
  NBUFFX2 U9144 ( .INP(n9643), .Z(n9606) );
  NBUFFX2 U9145 ( .INP(n9643), .Z(n9603) );
  NBUFFX2 U9146 ( .INP(n9640), .Z(n9620) );
  NBUFFX2 U9147 ( .INP(n9640), .Z(n9619) );
  NBUFFX2 U9148 ( .INP(n9643), .Z(n9602) );
  NBUFFX2 U9149 ( .INP(n9644), .Z(n9601) );
  NBUFFX2 U9150 ( .INP(n9644), .Z(n9600) );
  NBUFFX2 U9151 ( .INP(n9644), .Z(n9599) );
  NBUFFX2 U9152 ( .INP(n9644), .Z(n9598) );
  NBUFFX2 U9153 ( .INP(n9644), .Z(n9597) );
  NBUFFX2 U9154 ( .INP(n9645), .Z(n9596) );
  NBUFFX2 U9155 ( .INP(n9645), .Z(n9595) );
  NBUFFX2 U9156 ( .INP(n9645), .Z(n9594) );
  NBUFFX2 U9157 ( .INP(n9645), .Z(n9593) );
  NBUFFX2 U9158 ( .INP(n9646), .Z(n9590) );
  NBUFFX2 U9159 ( .INP(n9646), .Z(n9591) );
  NBUFFX2 U9160 ( .INP(n9645), .Z(n9592) );
  NBUFFX2 U9161 ( .INP(n9639), .Z(n9622) );
  NBUFFX2 U9162 ( .INP(n9640), .Z(n9621) );
  NBUFFX2 U9163 ( .INP(n9646), .Z(n9589) );
  NBUFFX2 U9164 ( .INP(n9646), .Z(n9588) );
  NBUFFX2 U9165 ( .INP(n9646), .Z(n9587) );
  NBUFFX2 U9166 ( .INP(n9647), .Z(n9586) );
  NBUFFX2 U9167 ( .INP(n9647), .Z(n9585) );
  NBUFFX2 U9168 ( .INP(n9647), .Z(n9584) );
  NBUFFX2 U9169 ( .INP(n9647), .Z(n9583) );
  NBUFFX2 U9170 ( .INP(n9647), .Z(n9582) );
  NBUFFX2 U9171 ( .INP(n9648), .Z(n9581) );
  NBUFFX2 U9172 ( .INP(n9648), .Z(n9580) );
  NBUFFX2 U9173 ( .INP(n9648), .Z(n9579) );
  NBUFFX2 U9174 ( .INP(n9649), .Z(n9576) );
  NBUFFX2 U9175 ( .INP(n9648), .Z(n9577) );
  NBUFFX2 U9176 ( .INP(n9648), .Z(n9578) );
  NBUFFX2 U9177 ( .INP(n9639), .Z(n9625) );
  NBUFFX2 U9178 ( .INP(n9639), .Z(n9624) );
  NBUFFX2 U9179 ( .INP(n9639), .Z(n9623) );
  NBUFFX2 U9180 ( .INP(n9649), .Z(n9575) );
  NBUFFX2 U9181 ( .INP(n9649), .Z(n9574) );
  NBUFFX2 U9182 ( .INP(n9649), .Z(n9573) );
  NBUFFX2 U9183 ( .INP(n9649), .Z(n9572) );
  NBUFFX2 U9184 ( .INP(n9650), .Z(n9571) );
  NBUFFX2 U9185 ( .INP(n9650), .Z(n9570) );
  NBUFFX2 U9186 ( .INP(n9650), .Z(n9569) );
  NBUFFX2 U9187 ( .INP(n9650), .Z(n9568) );
  NBUFFX2 U9188 ( .INP(n9650), .Z(n9567) );
  NBUFFX2 U9189 ( .INP(n9651), .Z(n9566) );
  NBUFFX2 U9190 ( .INP(n9651), .Z(n9565) );
  NBUFFX2 U9191 ( .INP(n9651), .Z(n9563) );
  NBUFFX2 U9192 ( .INP(n9651), .Z(n9564) );
  NBUFFX2 U9193 ( .INP(n9651), .Z(n9562) );
  NBUFFX2 U9194 ( .INP(n9639), .Z(n9626) );
  NBUFFX2 U9195 ( .INP(n9652), .Z(n9561) );
  NBUFFX2 U9196 ( .INP(n9652), .Z(n9560) );
  NBUFFX2 U9197 ( .INP(n9652), .Z(n9559) );
  NBUFFX2 U9198 ( .INP(n9652), .Z(n9558) );
  NBUFFX2 U9199 ( .INP(n9652), .Z(n9557) );
  NBUFFX2 U9200 ( .INP(n9653), .Z(n9556) );
  NBUFFX2 U9201 ( .INP(n9653), .Z(n9555) );
  NBUFFX2 U9202 ( .INP(n9653), .Z(n9554) );
  NBUFFX2 U9203 ( .INP(n9653), .Z(n9553) );
  NBUFFX2 U9204 ( .INP(n9653), .Z(n9552) );
  NBUFFX2 U9205 ( .INP(n9654), .Z(n9551) );
  NBUFFX2 U9206 ( .INP(n9654), .Z(n9548) );
  NBUFFX2 U9207 ( .INP(n9654), .Z(n9549) );
  NBUFFX2 U9208 ( .INP(n9654), .Z(n9550) );
  NBUFFX2 U9209 ( .INP(n9638), .Z(n9629) );
  NBUFFX2 U9210 ( .INP(n9638), .Z(n9628) );
  NBUFFX2 U9211 ( .INP(n9638), .Z(n9627) );
  NBUFFX2 U9212 ( .INP(n9654), .Z(n9547) );
  NBUFFX2 U9213 ( .INP(n9655), .Z(n9546) );
  NBUFFX2 U9214 ( .INP(n9655), .Z(n9545) );
  NBUFFX2 U9215 ( .INP(n9655), .Z(n9544) );
  NBUFFX2 U9216 ( .INP(n9655), .Z(n9543) );
  NBUFFX2 U9217 ( .INP(n9655), .Z(n9542) );
  NBUFFX2 U9218 ( .INP(n9656), .Z(n9541) );
  NBUFFX2 U9219 ( .INP(n9656), .Z(n9540) );
  NBUFFX2 U9220 ( .INP(n9656), .Z(n9539) );
  NBUFFX2 U9221 ( .INP(n9656), .Z(n9538) );
  NBUFFX2 U9222 ( .INP(n9657), .Z(n9535) );
  NBUFFX2 U9223 ( .INP(n9657), .Z(n9536) );
  NBUFFX2 U9224 ( .INP(n9656), .Z(n9537) );
  NBUFFX2 U9225 ( .INP(n9657), .Z(n9534) );
  NBUFFX2 U9226 ( .INP(n9638), .Z(n9631) );
  NBUFFX2 U9227 ( .INP(n9638), .Z(n9630) );
  NBUFFX2 U9228 ( .INP(n9657), .Z(n9533) );
  NBUFFX2 U9229 ( .INP(n9657), .Z(n9532) );
  NBUFFX2 U9230 ( .INP(n9658), .Z(n9531) );
  NBUFFX2 U9231 ( .INP(n9658), .Z(n9530) );
  NBUFFX2 U9232 ( .INP(n9658), .Z(n9529) );
  NBUFFX2 U9233 ( .INP(n9658), .Z(n9528) );
  NBUFFX2 U9234 ( .INP(n9658), .Z(n9527) );
  NBUFFX2 U9235 ( .INP(n9659), .Z(n9526) );
  NBUFFX2 U9236 ( .INP(n9659), .Z(n9525) );
  NBUFFX2 U9237 ( .INP(n9659), .Z(n9524) );
  NBUFFX2 U9238 ( .INP(n9660), .Z(n9521) );
  NBUFFX2 U9239 ( .INP(n9659), .Z(n9522) );
  NBUFFX2 U9240 ( .INP(n9659), .Z(n9523) );
  NBUFFX2 U9241 ( .INP(n9637), .Z(n9634) );
  NBUFFX2 U9242 ( .INP(n9637), .Z(n9633) );
  NBUFFX2 U9243 ( .INP(n9637), .Z(n9632) );
  NBUFFX2 U9244 ( .INP(n9660), .Z(n9520) );
  NBUFFX2 U9245 ( .INP(n9660), .Z(n9519) );
  NBUFFX2 U9246 ( .INP(n9660), .Z(n9518) );
  NBUFFX2 U9247 ( .INP(n9660), .Z(n9517) );
  NBUFFX2 U9248 ( .INP(n9661), .Z(n9516) );
  NBUFFX2 U9249 ( .INP(n9661), .Z(n9515) );
  NBUFFX2 U9250 ( .INP(n9661), .Z(n9514) );
  NBUFFX2 U9251 ( .INP(n9661), .Z(n9513) );
  NBUFFX2 U9252 ( .INP(n9661), .Z(n9512) );
  NBUFFX2 U9253 ( .INP(n9662), .Z(n9511) );
  NBUFFX2 U9254 ( .INP(n9662), .Z(n9510) );
  NBUFFX2 U9255 ( .INP(n9662), .Z(n9508) );
  NBUFFX2 U9256 ( .INP(n9662), .Z(n9509) );
  NBUFFX2 U9257 ( .INP(n9662), .Z(n9507) );
  NBUFFX2 U9258 ( .INP(n9637), .Z(n9636) );
  NBUFFX2 U9259 ( .INP(n9637), .Z(n9635) );
  NBUFFX2 U9260 ( .INP(n9663), .Z(n9506) );
  NBUFFX2 U9261 ( .INP(n9663), .Z(n9505) );
  NBUFFX2 U9262 ( .INP(n9663), .Z(n9504) );
  NBUFFX2 U9263 ( .INP(n9663), .Z(n9503) );
  NBUFFX2 U9264 ( .INP(n9663), .Z(n9502) );
  NBUFFX2 U9265 ( .INP(n9664), .Z(n9501) );
  NBUFFX2 U9266 ( .INP(n9664), .Z(n9500) );
  NBUFFX2 U9267 ( .INP(n9664), .Z(n9499) );
  NBUFFX2 U9268 ( .INP(n9664), .Z(n9498) );
  NBUFFX2 U9269 ( .INP(n9664), .Z(n9497) );
  NBUFFX2 U9270 ( .INP(n9269), .Z(n9288) );
  NBUFFX2 U9271 ( .INP(n9263), .Z(n9136) );
  NBUFFX2 U9272 ( .INP(n9263), .Z(n9135) );
  NBUFFX2 U9273 ( .INP(n9271), .Z(n9264) );
  NBUFFX2 U9274 ( .INP(n9270), .Z(n9267) );
  NBUFFX2 U9275 ( .INP(n9270), .Z(n9268) );
  NBUFFX2 U9276 ( .INP(n9271), .Z(n9265) );
  NBUFFX2 U9277 ( .INP(n9271), .Z(n9266) );
  NBUFFX2 U9278 ( .INP(n9270), .Z(n9269) );
  NBUFFX2 U9279 ( .INP(n9112), .Z(n9116) );
  NBUFFX2 U9280 ( .INP(n9112), .Z(n9115) );
  NBUFFX2 U9281 ( .INP(n9112), .Z(n9117) );
  NBUFFX2 U9282 ( .INP(n9113), .Z(n9119) );
  NBUFFX2 U9283 ( .INP(n9113), .Z(n9118) );
  NBUFFX2 U9284 ( .INP(n9114), .Z(n9121) );
  NBUFFX2 U9285 ( .INP(n9114), .Z(n9122) );
  NBUFFX2 U9286 ( .INP(n9113), .Z(n9120) );
  NBUFFX2 U9287 ( .INP(n9084), .Z(n9091) );
  NBUFFX2 U9288 ( .INP(n9088), .Z(n9110) );
  NBUFFX2 U9289 ( .INP(n9088), .Z(n9109) );
  NBUFFX2 U9290 ( .INP(n9084), .Z(n9089) );
  NBUFFX2 U9291 ( .INP(n9084), .Z(n9090) );
  NBUFFX2 U9292 ( .INP(n9087), .Z(n9107) );
  NBUFFX2 U9293 ( .INP(n9087), .Z(n9105) );
  NBUFFX2 U9294 ( .INP(n9086), .Z(n9103) );
  NBUFFX2 U9295 ( .INP(n9086), .Z(n9102) );
  NBUFFX2 U9296 ( .INP(n9086), .Z(n9101) );
  NBUFFX2 U9297 ( .INP(n9086), .Z(n9100) );
  NBUFFX2 U9298 ( .INP(n9086), .Z(n9099) );
  NBUFFX2 U9299 ( .INP(n9085), .Z(n9098) );
  NBUFFX2 U9300 ( .INP(n9085), .Z(n9097) );
  NBUFFX2 U9301 ( .INP(n9085), .Z(n9096) );
  NBUFFX2 U9302 ( .INP(n9085), .Z(n9095) );
  NBUFFX2 U9303 ( .INP(n9087), .Z(n9106) );
  NBUFFX2 U9304 ( .INP(n9087), .Z(n9108) );
  NBUFFX2 U9305 ( .INP(n9087), .Z(n9104) );
  NBUFFX2 U9306 ( .INP(n9084), .Z(n9092) );
  NBUFFX2 U9307 ( .INP(n9084), .Z(n9093) );
  NBUFFX2 U9308 ( .INP(n9085), .Z(n9094) );
  NBUFFX2 U9309 ( .INP(n9114), .Z(n9123) );
  NBUFFX2 U9310 ( .INP(n9088), .Z(n9111) );
  NBUFFX2 U9311 ( .INP(n2148), .Z(n9270) );
  NBUFFX2 U9312 ( .INP(n2148), .Z(n9271) );
  INVX0 U9313 ( .INP(n9341), .ZN(n9491) );
  INVX0 U9314 ( .INP(n9340), .ZN(n9490) );
  INVX0 U9315 ( .INP(n9340), .ZN(n9489) );
  INVX0 U9316 ( .INP(n9339), .ZN(n9488) );
  INVX0 U9317 ( .INP(n9339), .ZN(n9487) );
  INVX0 U9318 ( .INP(n9338), .ZN(n9486) );
  INVX0 U9319 ( .INP(n9338), .ZN(n9485) );
  INVX0 U9320 ( .INP(n9341), .ZN(n9492) );
  INVX0 U9321 ( .INP(n9337), .ZN(n9484) );
  INVX0 U9322 ( .INP(n9337), .ZN(n9483) );
  NBUFFX2 U9323 ( .INP(n10355), .Z(n9114) );
  NBUFFX2 U9324 ( .INP(n10355), .Z(n9112) );
  NBUFFX2 U9325 ( .INP(n10355), .Z(n9113) );
  NBUFFX2 U9326 ( .INP(n9342), .Z(n9340) );
  NBUFFX2 U9327 ( .INP(n9342), .Z(n9339) );
  NBUFFX2 U9328 ( .INP(n9343), .Z(n9338) );
  NBUFFX2 U9329 ( .INP(n9342), .Z(n9341) );
  NBUFFX2 U9330 ( .INP(n9343), .Z(n9337) );
  INVX0 U9331 ( .INP(n2153), .ZN(n9336) );
  NBUFFX2 U9332 ( .INP(n9680), .Z(n9084) );
  NBUFFX2 U9333 ( .INP(n9680), .Z(n9085) );
  NBUFFX2 U9334 ( .INP(n9680), .Z(n9086) );
  NBUFFX2 U9335 ( .INP(n9680), .Z(n9087) );
  NBUFFX2 U9336 ( .INP(n9680), .Z(n9088) );
  NBUFFX2 U9337 ( .INP(n9134), .Z(n9124) );
  NBUFFX2 U9338 ( .INP(n9134), .Z(n9125) );
  NBUFFX2 U9339 ( .INP(n9133), .Z(n9126) );
  NBUFFX2 U9340 ( .INP(n9133), .Z(n9127) );
  NBUFFX2 U9341 ( .INP(n9133), .Z(n9128) );
  NBUFFX2 U9342 ( .INP(n9132), .Z(n9129) );
  NBUFFX2 U9343 ( .INP(n9132), .Z(n9130) );
  NBUFFX2 U9344 ( .INP(n9132), .Z(n9131) );
  NBUFFX2 U9345 ( .INP(n2181), .Z(n9132) );
  NBUFFX2 U9346 ( .INP(n2181), .Z(n9133) );
  NBUFFX2 U9347 ( .INP(n2181), .Z(n9134) );
  NBUFFX2 U9348 ( .INP(n9124), .Z(n9242) );
  NBUFFX2 U9349 ( .INP(n9124), .Z(n9243) );
  NBUFFX2 U9350 ( .INP(n9124), .Z(n9244) );
  NBUFFX2 U9351 ( .INP(n9125), .Z(n9245) );
  NBUFFX2 U9352 ( .INP(n9125), .Z(n9246) );
  NBUFFX2 U9353 ( .INP(n9125), .Z(n9247) );
  NBUFFX2 U9354 ( .INP(n9126), .Z(n9248) );
  NBUFFX2 U9355 ( .INP(n9126), .Z(n9249) );
  NBUFFX2 U9356 ( .INP(n9126), .Z(n9250) );
  NBUFFX2 U9357 ( .INP(n9127), .Z(n9251) );
  NBUFFX2 U9358 ( .INP(n9127), .Z(n9252) );
  NBUFFX2 U9359 ( .INP(n9127), .Z(n9253) );
  NBUFFX2 U9360 ( .INP(n9128), .Z(n9254) );
  NBUFFX2 U9361 ( .INP(n9128), .Z(n9255) );
  NBUFFX2 U9362 ( .INP(n9128), .Z(n9256) );
  NBUFFX2 U9363 ( .INP(n9129), .Z(n9257) );
  NBUFFX2 U9364 ( .INP(n9129), .Z(n9258) );
  NBUFFX2 U9365 ( .INP(n9129), .Z(n9259) );
  NBUFFX2 U9366 ( .INP(n9130), .Z(n9260) );
  NBUFFX2 U9367 ( .INP(n9130), .Z(n9261) );
  NBUFFX2 U9368 ( .INP(n9130), .Z(n9262) );
  NBUFFX2 U9369 ( .INP(n9131), .Z(n9263) );
  NBUFFX2 U9370 ( .INP(n2152), .Z(n9289) );
  NBUFFX2 U9371 ( .INP(n2152), .Z(n9290) );
  NBUFFX2 U9372 ( .INP(n9289), .Z(n9315) );
  NBUFFX2 U9373 ( .INP(n9289), .Z(n9316) );
  NBUFFX2 U9374 ( .INP(n9289), .Z(n9317) );
  NBUFFX2 U9375 ( .INP(n9290), .Z(n9318) );
  NBUFFX2 U9376 ( .INP(n9290), .Z(n9319) );
  INVX0 U9377 ( .INP(n9336), .ZN(n9320) );
  INVX0 U9378 ( .INP(n9336), .ZN(n9321) );
  INVX0 U9379 ( .INP(n9336), .ZN(n9322) );
  INVX0 U9380 ( .INP(n9336), .ZN(n9323) );
  INVX0 U9381 ( .INP(n9336), .ZN(n9324) );
  INVX0 U9382 ( .INP(n9336), .ZN(n9325) );
  INVX0 U9383 ( .INP(n9336), .ZN(n9326) );
  INVX0 U9384 ( .INP(n9336), .ZN(n9327) );
  INVX0 U9385 ( .INP(n9336), .ZN(n9328) );
  INVX0 U9386 ( .INP(n9336), .ZN(n9329) );
  INVX0 U9387 ( .INP(n9336), .ZN(n9330) );
  INVX0 U9388 ( .INP(n9336), .ZN(n9331) );
  INVX0 U9389 ( .INP(n9336), .ZN(n9332) );
  INVX0 U9390 ( .INP(n9336), .ZN(n9333) );
  INVX0 U9391 ( .INP(n9336), .ZN(n9334) );
  INVX0 U9392 ( .INP(n9336), .ZN(n9335) );
  NBUFFX2 U9393 ( .INP(test_se), .Z(n9342) );
  NBUFFX2 U9394 ( .INP(test_se), .Z(n9343) );
  INVX0 U9395 ( .INP(n9491), .ZN(n9344) );
  INVX0 U9396 ( .INP(n9491), .ZN(n9345) );
  INVX0 U9397 ( .INP(n9486), .ZN(n9346) );
  INVX0 U9398 ( .INP(n9488), .ZN(n9347) );
  INVX0 U9399 ( .INP(n9489), .ZN(n9348) );
  INVX0 U9400 ( .INP(n9490), .ZN(n9349) );
  INVX0 U9401 ( .INP(n9489), .ZN(n9350) );
  INVX0 U9402 ( .INP(n9488), .ZN(n9351) );
  INVX0 U9403 ( .INP(n9487), .ZN(n9352) );
  INVX0 U9404 ( .INP(n9491), .ZN(n9353) );
  INVX0 U9405 ( .INP(n9492), .ZN(n9354) );
  INVX0 U9406 ( .INP(n9488), .ZN(n9355) );
  INVX0 U9407 ( .INP(n9492), .ZN(n9356) );
  INVX0 U9408 ( .INP(n9492), .ZN(n9357) );
  INVX0 U9409 ( .INP(n9492), .ZN(n9358) );
  INVX0 U9410 ( .INP(n9492), .ZN(n9359) );
  INVX0 U9411 ( .INP(n9492), .ZN(n9360) );
  INVX0 U9412 ( .INP(n9492), .ZN(n9361) );
  INVX0 U9413 ( .INP(n9491), .ZN(n9362) );
  INVX0 U9414 ( .INP(n9491), .ZN(n9363) );
  INVX0 U9415 ( .INP(n9491), .ZN(n9364) );
  INVX0 U9416 ( .INP(n9491), .ZN(n9365) );
  INVX0 U9417 ( .INP(n9491), .ZN(n9366) );
  INVX0 U9418 ( .INP(n9491), .ZN(n9367) );
  INVX0 U9419 ( .INP(n9490), .ZN(n9368) );
  INVX0 U9420 ( .INP(n9490), .ZN(n9369) );
  INVX0 U9421 ( .INP(n9490), .ZN(n9370) );
  INVX0 U9422 ( .INP(n9490), .ZN(n9371) );
  INVX0 U9423 ( .INP(n9490), .ZN(n9372) );
  INVX0 U9424 ( .INP(n9490), .ZN(n9373) );
  INVX0 U9425 ( .INP(n9489), .ZN(n9374) );
  INVX0 U9426 ( .INP(n9489), .ZN(n9375) );
  INVX0 U9427 ( .INP(n9489), .ZN(n9376) );
  INVX0 U9428 ( .INP(n9489), .ZN(n9377) );
  INVX0 U9429 ( .INP(n9489), .ZN(n9378) );
  INVX0 U9430 ( .INP(n9489), .ZN(n9379) );
  INVX0 U9431 ( .INP(n9488), .ZN(n9380) );
  INVX0 U9432 ( .INP(n9488), .ZN(n9381) );
  INVX0 U9433 ( .INP(n9488), .ZN(n9382) );
  INVX0 U9434 ( .INP(n9488), .ZN(n9383) );
  INVX0 U9435 ( .INP(n9488), .ZN(n9384) );
  INVX0 U9436 ( .INP(n9488), .ZN(n9385) );
  INVX0 U9437 ( .INP(n9487), .ZN(n9386) );
  INVX0 U9438 ( .INP(n9487), .ZN(n9387) );
  INVX0 U9439 ( .INP(n9487), .ZN(n9388) );
  INVX0 U9440 ( .INP(n9487), .ZN(n9389) );
  INVX0 U9441 ( .INP(n9487), .ZN(n9390) );
  INVX0 U9442 ( .INP(n9487), .ZN(n9391) );
  INVX0 U9443 ( .INP(n9486), .ZN(n9392) );
  INVX0 U9444 ( .INP(n9486), .ZN(n9393) );
  INVX0 U9445 ( .INP(n9486), .ZN(n9394) );
  INVX0 U9446 ( .INP(n9486), .ZN(n9395) );
  INVX0 U9447 ( .INP(n9486), .ZN(n9396) );
  INVX0 U9448 ( .INP(n9486), .ZN(n9397) );
  INVX0 U9449 ( .INP(n9485), .ZN(n9398) );
  INVX0 U9450 ( .INP(n9485), .ZN(n9399) );
  INVX0 U9451 ( .INP(n9485), .ZN(n9400) );
  INVX0 U9452 ( .INP(n9485), .ZN(n9401) );
  INVX0 U9453 ( .INP(n9485), .ZN(n9402) );
  INVX0 U9454 ( .INP(n9485), .ZN(n9403) );
  INVX0 U9455 ( .INP(n9484), .ZN(n9404) );
  INVX0 U9456 ( .INP(n9484), .ZN(n9405) );
  INVX0 U9457 ( .INP(n9484), .ZN(n9406) );
  INVX0 U9458 ( .INP(n9484), .ZN(n9407) );
  INVX0 U9459 ( .INP(n9484), .ZN(n9408) );
  INVX0 U9460 ( .INP(n9484), .ZN(n9409) );
  INVX0 U9461 ( .INP(n9483), .ZN(n9410) );
  INVX0 U9462 ( .INP(n9483), .ZN(n9411) );
  INVX0 U9463 ( .INP(n9483), .ZN(n9412) );
  INVX0 U9464 ( .INP(n9483), .ZN(n9413) );
  INVX0 U9465 ( .INP(n9483), .ZN(n9414) );
  INVX0 U9466 ( .INP(n9483), .ZN(n9415) );
  INVX0 U9467 ( .INP(n9486), .ZN(n9416) );
  INVX0 U9468 ( .INP(n9485), .ZN(n9417) );
  INVX0 U9469 ( .INP(n9484), .ZN(n9418) );
  INVX0 U9470 ( .INP(n9483), .ZN(n9419) );
  INVX0 U9471 ( .INP(n9486), .ZN(n9420) );
  INVX0 U9472 ( .INP(n9490), .ZN(n9421) );
  INVX0 U9473 ( .INP(n9486), .ZN(n9422) );
  INVX0 U9474 ( .INP(n9485), .ZN(n9423) );
  INVX0 U9475 ( .INP(n9484), .ZN(n9424) );
  INVX0 U9476 ( .INP(n9483), .ZN(n9425) );
  INVX0 U9477 ( .INP(n9490), .ZN(n9426) );
  INVX0 U9478 ( .INP(n9485), .ZN(n9427) );
  INVX0 U9479 ( .INP(n9484), .ZN(n9428) );
  INVX0 U9480 ( .INP(n9483), .ZN(n9429) );
  INVX0 U9481 ( .INP(n9489), .ZN(n9430) );
  INVX0 U9482 ( .INP(n9489), .ZN(n9431) );
  INVX0 U9483 ( .INP(n9484), .ZN(n9432) );
  INVX0 U9484 ( .INP(n9490), .ZN(n9433) );
  INVX0 U9485 ( .INP(n9491), .ZN(n9434) );
  INVX0 U9486 ( .INP(n9483), .ZN(n9435) );
  INVX0 U9487 ( .INP(n9490), .ZN(n9436) );
  INVX0 U9488 ( .INP(n9489), .ZN(n9437) );
  INVX0 U9489 ( .INP(n9488), .ZN(n9438) );
  INVX0 U9490 ( .INP(n9487), .ZN(n9439) );
  INVX0 U9491 ( .INP(n9487), .ZN(n9440) );
  INVX0 U9492 ( .INP(n9491), .ZN(n9441) );
  INVX0 U9493 ( .INP(n9492), .ZN(n9442) );
  INVX0 U9494 ( .INP(n9486), .ZN(n9443) );
  INVX0 U9495 ( .INP(n9485), .ZN(n9444) );
  INVX0 U9496 ( .INP(n9484), .ZN(n9445) );
  INVX0 U9497 ( .INP(n9488), .ZN(n9446) );
  INVX0 U9498 ( .INP(n9487), .ZN(n9447) );
  INVX0 U9499 ( .INP(n9491), .ZN(n9448) );
  INVX0 U9500 ( .INP(n9492), .ZN(n9449) );
  INVX0 U9501 ( .INP(n9490), .ZN(n9450) );
  INVX0 U9502 ( .INP(n9489), .ZN(n9451) );
  INVX0 U9503 ( .INP(n9491), .ZN(n9452) );
  INVX0 U9504 ( .INP(n9486), .ZN(n9453) );
  INVX0 U9505 ( .INP(n9485), .ZN(n9454) );
  INVX0 U9506 ( .INP(n9484), .ZN(n9455) );
  INVX0 U9507 ( .INP(n9483), .ZN(n9456) );
  INVX0 U9508 ( .INP(n9484), .ZN(n9457) );
  INVX0 U9509 ( .INP(n9483), .ZN(n9458) );
  INVX0 U9510 ( .INP(n9487), .ZN(n9459) );
  INVX0 U9511 ( .INP(n9487), .ZN(n9460) );
  INVX0 U9512 ( .INP(n9483), .ZN(n9461) );
  INVX0 U9513 ( .INP(n9485), .ZN(n9462) );
  INVX0 U9514 ( .INP(n9487), .ZN(n9463) );
  INVX0 U9515 ( .INP(n9486), .ZN(n9464) );
  INVX0 U9516 ( .INP(n9485), .ZN(n9465) );
  INVX0 U9517 ( .INP(n9484), .ZN(n9466) );
  INVX0 U9518 ( .INP(n9483), .ZN(n9467) );
  INVX0 U9519 ( .INP(n9488), .ZN(n9468) );
  INVX0 U9520 ( .INP(n9487), .ZN(n9469) );
  INVX0 U9521 ( .INP(n9491), .ZN(n9470) );
  INVX0 U9522 ( .INP(n9490), .ZN(n9471) );
  INVX0 U9523 ( .INP(n9486), .ZN(n9472) );
  INVX0 U9524 ( .INP(n9485), .ZN(n9473) );
  INVX0 U9525 ( .INP(n9488), .ZN(n9474) );
  INVX0 U9526 ( .INP(n9488), .ZN(n9475) );
  INVX0 U9527 ( .INP(n9489), .ZN(n9476) );
  INVX0 U9528 ( .INP(n9490), .ZN(n9477) );
  INVX0 U9529 ( .INP(n9489), .ZN(n9478) );
  INVX0 U9530 ( .INP(n9486), .ZN(n9479) );
  INVX0 U9531 ( .INP(n9485), .ZN(n9480) );
  INVX0 U9532 ( .INP(n9484), .ZN(n9481) );
  INVX0 U9533 ( .INP(n9483), .ZN(n9482) );
  NBUFFX2 U9534 ( .INP(n9675), .Z(n9637) );
  NBUFFX2 U9535 ( .INP(n9675), .Z(n9638) );
  NBUFFX2 U9536 ( .INP(n9674), .Z(n9639) );
  NBUFFX2 U9537 ( .INP(n9674), .Z(n9640) );
  NBUFFX2 U9538 ( .INP(n9674), .Z(n9641) );
  NBUFFX2 U9539 ( .INP(n9673), .Z(n9642) );
  NBUFFX2 U9540 ( .INP(n9673), .Z(n9643) );
  NBUFFX2 U9541 ( .INP(n9673), .Z(n9644) );
  NBUFFX2 U9542 ( .INP(n9672), .Z(n9645) );
  NBUFFX2 U9543 ( .INP(n9672), .Z(n9646) );
  NBUFFX2 U9544 ( .INP(n9672), .Z(n9647) );
  NBUFFX2 U9545 ( .INP(n9671), .Z(n9648) );
  NBUFFX2 U9546 ( .INP(n9671), .Z(n9649) );
  NBUFFX2 U9547 ( .INP(n9671), .Z(n9650) );
  NBUFFX2 U9548 ( .INP(n9670), .Z(n9651) );
  NBUFFX2 U9549 ( .INP(n9670), .Z(n9652) );
  NBUFFX2 U9550 ( .INP(n9670), .Z(n9653) );
  NBUFFX2 U9551 ( .INP(n9669), .Z(n9654) );
  NBUFFX2 U9552 ( .INP(n9669), .Z(n9655) );
  NBUFFX2 U9553 ( .INP(n9669), .Z(n9656) );
  NBUFFX2 U9554 ( .INP(n9668), .Z(n9657) );
  NBUFFX2 U9555 ( .INP(n9668), .Z(n9658) );
  NBUFFX2 U9556 ( .INP(n9668), .Z(n9659) );
  NBUFFX2 U9557 ( .INP(n9667), .Z(n9660) );
  NBUFFX2 U9558 ( .INP(n9667), .Z(n9661) );
  NBUFFX2 U9559 ( .INP(n9667), .Z(n9662) );
  NBUFFX2 U9560 ( .INP(n9666), .Z(n9663) );
  NBUFFX2 U9561 ( .INP(n9666), .Z(n9664) );
  NBUFFX2 U9562 ( .INP(n9666), .Z(n9665) );
  NBUFFX2 U9563 ( .INP(CK), .Z(n9666) );
  NBUFFX2 U9564 ( .INP(CK), .Z(n9667) );
  NBUFFX2 U9565 ( .INP(n9675), .Z(n9668) );
  NBUFFX2 U9566 ( .INP(CK), .Z(n9669) );
  NBUFFX2 U9567 ( .INP(n9671), .Z(n9670) );
  NBUFFX2 U9568 ( .INP(CK), .Z(n9671) );
  NBUFFX2 U9569 ( .INP(n9666), .Z(n9672) );
  NBUFFX2 U9570 ( .INP(n9667), .Z(n9673) );
  NBUFFX2 U9571 ( .INP(n9669), .Z(n9674) );
  NBUFFX2 U9572 ( .INP(n9506), .Z(n9675) );
  NOR2X0 U9573 ( .IN1(TM1), .IN2(n9158), .QN(n3278) );
  NOR2X0 U9574 ( .IN1(n16132), .IN2(n9158), .QN(WX9789) );
  NOR2X0 U9575 ( .IN1(n16131), .IN2(n9158), .QN(WX9787) );
  NOR2X0 U9576 ( .IN1(n16130), .IN2(n9158), .QN(WX9785) );
  NOR2X0 U9577 ( .IN1(n16129), .IN2(n9158), .QN(WX9783) );
  NOR2X0 U9578 ( .IN1(n9236), .IN2(n8819), .QN(WX9781) );
  NOR2X0 U9579 ( .IN1(n16128), .IN2(n9158), .QN(WX9779) );
  NOR2X0 U9580 ( .IN1(n16127), .IN2(n9157), .QN(WX9777) );
  NOR2X0 U9581 ( .IN1(n16126), .IN2(n9157), .QN(WX9775) );
  NOR2X0 U9582 ( .IN1(n16125), .IN2(n9157), .QN(WX9773) );
  NOR2X0 U9583 ( .IN1(n16124), .IN2(n9157), .QN(WX9771) );
  NOR2X0 U9584 ( .IN1(n16123), .IN2(n9157), .QN(WX9769) );
  NOR2X0 U9585 ( .IN1(n16122), .IN2(n9157), .QN(WX9767) );
  NOR2X0 U9586 ( .IN1(n16121), .IN2(n9157), .QN(WX9765) );
  NOR2X0 U9587 ( .IN1(n16120), .IN2(n9156), .QN(WX9763) );
  NOR2X0 U9588 ( .IN1(n16119), .IN2(n9156), .QN(WX9761) );
  NOR2X0 U9589 ( .IN1(n16118), .IN2(n9156), .QN(WX9759) );
  NAND4X0 U9590 ( .IN1(n9676), .IN2(n9677), .IN3(n9678), .IN4(n9679), .QN(
        WX9757) );
  NAND2X0 U9591 ( .IN1(n9100), .IN2(n9681), .QN(n9679) );
  NAND2X0 U9592 ( .IN1(n9322), .IN2(n9682), .QN(n9678) );
  NAND2X0 U9593 ( .IN1(n9272), .IN2(n1727), .QN(n9677) );
  NOR2X0 U9594 ( .IN1(n9231), .IN2(n8828), .QN(n1727) );
  NAND2X0 U9595 ( .IN1(n9291), .IN2(CRC_OUT_2_0), .QN(n9676) );
  NAND4X0 U9596 ( .IN1(n9683), .IN2(n9684), .IN3(n9685), .IN4(n9686), .QN(
        WX9755) );
  NAND3X0 U9597 ( .IN1(n9687), .IN2(n9688), .IN3(n9089), .QN(n9686) );
  NAND2X0 U9598 ( .IN1(n9331), .IN2(n9689), .QN(n9685) );
  NAND2X0 U9599 ( .IN1(n1726), .IN2(n9272), .QN(n9684) );
  NOR2X0 U9600 ( .IN1(n9233), .IN2(n8829), .QN(n1726) );
  NAND2X0 U9601 ( .IN1(n9308), .IN2(CRC_OUT_2_1), .QN(n9683) );
  NAND4X0 U9602 ( .IN1(n9690), .IN2(n9691), .IN3(n9692), .IN4(n9693), .QN(
        WX9753) );
  NAND3X0 U9603 ( .IN1(n9694), .IN2(n9695), .IN3(n9320), .QN(n9693) );
  NAND2X0 U9604 ( .IN1(n9100), .IN2(n9696), .QN(n9692) );
  NAND2X0 U9605 ( .IN1(n1725), .IN2(n9272), .QN(n9691) );
  NOR2X0 U9606 ( .IN1(n9233), .IN2(n8830), .QN(n1725) );
  NAND2X0 U9607 ( .IN1(test_so87), .IN2(n9314), .QN(n9690) );
  NAND4X0 U9608 ( .IN1(n9697), .IN2(n9698), .IN3(n9699), .IN4(n9700), .QN(
        WX9751) );
  NAND3X0 U9609 ( .IN1(n9701), .IN2(n9702), .IN3(n9089), .QN(n9700) );
  NAND2X0 U9610 ( .IN1(n9328), .IN2(n9703), .QN(n9699) );
  NAND2X0 U9611 ( .IN1(n1724), .IN2(n9272), .QN(n9698) );
  NOR2X0 U9612 ( .IN1(n9233), .IN2(n8831), .QN(n1724) );
  NAND2X0 U9613 ( .IN1(n9302), .IN2(CRC_OUT_2_3), .QN(n9697) );
  NAND4X0 U9614 ( .IN1(n9704), .IN2(n9705), .IN3(n9706), .IN4(n9707), .QN(
        WX9749) );
  NAND3X0 U9615 ( .IN1(n9708), .IN2(n9709), .IN3(n9320), .QN(n9707) );
  NAND2X0 U9616 ( .IN1(n9100), .IN2(n9710), .QN(n9706) );
  NAND2X0 U9617 ( .IN1(n1723), .IN2(n9272), .QN(n9705) );
  NOR2X0 U9618 ( .IN1(n9233), .IN2(n8832), .QN(n1723) );
  NAND2X0 U9619 ( .IN1(n9302), .IN2(CRC_OUT_2_4), .QN(n9704) );
  NAND4X0 U9620 ( .IN1(n9711), .IN2(n9712), .IN3(n9713), .IN4(n9714), .QN(
        WX9747) );
  NAND2X0 U9621 ( .IN1(n9100), .IN2(n9715), .QN(n9714) );
  NAND2X0 U9622 ( .IN1(n9328), .IN2(n9716), .QN(n9713) );
  NAND2X0 U9623 ( .IN1(n1722), .IN2(n9272), .QN(n9712) );
  NOR2X0 U9624 ( .IN1(n9060), .IN2(n9155), .QN(n1722) );
  NAND2X0 U9625 ( .IN1(n9302), .IN2(CRC_OUT_2_5), .QN(n9711) );
  NAND4X0 U9626 ( .IN1(n9717), .IN2(n9718), .IN3(n9719), .IN4(n9720), .QN(
        WX9745) );
  NAND3X0 U9627 ( .IN1(n9721), .IN2(n9722), .IN3(n9320), .QN(n9720) );
  NAND2X0 U9628 ( .IN1(n9100), .IN2(n9723), .QN(n9719) );
  NAND2X0 U9629 ( .IN1(n1721), .IN2(n9272), .QN(n9718) );
  NOR2X0 U9630 ( .IN1(n9234), .IN2(n8833), .QN(n1721) );
  NAND2X0 U9631 ( .IN1(n9302), .IN2(CRC_OUT_2_6), .QN(n9717) );
  NAND4X0 U9632 ( .IN1(n9724), .IN2(n9725), .IN3(n9726), .IN4(n9727), .QN(
        WX9743) );
  NAND2X0 U9633 ( .IN1(n9100), .IN2(n9728), .QN(n9727) );
  NAND2X0 U9634 ( .IN1(n9328), .IN2(n9729), .QN(n9726) );
  NAND2X0 U9635 ( .IN1(n1720), .IN2(n9272), .QN(n9725) );
  NOR2X0 U9636 ( .IN1(n9234), .IN2(n8834), .QN(n1720) );
  NAND2X0 U9637 ( .IN1(n9303), .IN2(CRC_OUT_2_7), .QN(n9724) );
  NAND4X0 U9638 ( .IN1(n9730), .IN2(n9731), .IN3(n9732), .IN4(n9733), .QN(
        WX9741) );
  NAND3X0 U9639 ( .IN1(n9734), .IN2(n9735), .IN3(n9320), .QN(n9733) );
  NAND2X0 U9640 ( .IN1(n9100), .IN2(n9736), .QN(n9732) );
  NAND2X0 U9641 ( .IN1(n1719), .IN2(n9272), .QN(n9731) );
  NOR2X0 U9642 ( .IN1(n9234), .IN2(n8835), .QN(n1719) );
  NAND2X0 U9643 ( .IN1(n9303), .IN2(CRC_OUT_2_8), .QN(n9730) );
  NAND4X0 U9644 ( .IN1(n9737), .IN2(n9738), .IN3(n9739), .IN4(n9740), .QN(
        WX9739) );
  NAND2X0 U9645 ( .IN1(n9100), .IN2(n9741), .QN(n9740) );
  NAND2X0 U9646 ( .IN1(n9328), .IN2(n9742), .QN(n9739) );
  NAND2X0 U9647 ( .IN1(n1718), .IN2(n9272), .QN(n9738) );
  NOR2X0 U9648 ( .IN1(n9234), .IN2(n8836), .QN(n1718) );
  NAND2X0 U9649 ( .IN1(n9303), .IN2(CRC_OUT_2_9), .QN(n9737) );
  NAND4X0 U9650 ( .IN1(n9743), .IN2(n9744), .IN3(n9745), .IN4(n9746), .QN(
        WX9737) );
  NAND2X0 U9651 ( .IN1(n9100), .IN2(n9747), .QN(n9746) );
  NAND2X0 U9652 ( .IN1(n9328), .IN2(n9748), .QN(n9745) );
  NAND2X0 U9653 ( .IN1(n1717), .IN2(n9272), .QN(n9744) );
  NOR2X0 U9654 ( .IN1(n9234), .IN2(n8837), .QN(n1717) );
  NAND2X0 U9655 ( .IN1(n9303), .IN2(CRC_OUT_2_10), .QN(n9743) );
  NAND4X0 U9656 ( .IN1(n9749), .IN2(n9750), .IN3(n9751), .IN4(n9752), .QN(
        WX9735) );
  NAND2X0 U9657 ( .IN1(n9100), .IN2(n9753), .QN(n9752) );
  NAND2X0 U9658 ( .IN1(n9328), .IN2(n9754), .QN(n9751) );
  NAND2X0 U9659 ( .IN1(n1716), .IN2(n9272), .QN(n9750) );
  NOR2X0 U9660 ( .IN1(n9234), .IN2(n8838), .QN(n1716) );
  NAND2X0 U9661 ( .IN1(n9303), .IN2(CRC_OUT_2_11), .QN(n9749) );
  NAND4X0 U9662 ( .IN1(n9755), .IN2(n9756), .IN3(n9757), .IN4(n9758), .QN(
        WX9733) );
  NAND2X0 U9663 ( .IN1(n9099), .IN2(n9759), .QN(n9758) );
  NAND2X0 U9664 ( .IN1(n9328), .IN2(n9760), .QN(n9757) );
  NAND2X0 U9665 ( .IN1(n1715), .IN2(n9272), .QN(n9756) );
  NOR2X0 U9666 ( .IN1(n9234), .IN2(n8839), .QN(n1715) );
  NAND2X0 U9667 ( .IN1(n9303), .IN2(CRC_OUT_2_12), .QN(n9755) );
  NAND4X0 U9668 ( .IN1(n9761), .IN2(n9762), .IN3(n9763), .IN4(n9764), .QN(
        WX9731) );
  NAND2X0 U9669 ( .IN1(n9099), .IN2(n9765), .QN(n9764) );
  NAND2X0 U9670 ( .IN1(n9328), .IN2(n9766), .QN(n9763) );
  NAND2X0 U9671 ( .IN1(n1714), .IN2(n9272), .QN(n9762) );
  NOR2X0 U9672 ( .IN1(n9234), .IN2(n8840), .QN(n1714) );
  NAND2X0 U9673 ( .IN1(n9303), .IN2(CRC_OUT_2_13), .QN(n9761) );
  NAND4X0 U9674 ( .IN1(n9767), .IN2(n9768), .IN3(n9769), .IN4(n9770), .QN(
        WX9729) );
  NAND3X0 U9675 ( .IN1(n9771), .IN2(n9772), .IN3(n9089), .QN(n9770) );
  NAND2X0 U9676 ( .IN1(n9328), .IN2(n9773), .QN(n9769) );
  NAND2X0 U9677 ( .IN1(n1713), .IN2(n9272), .QN(n9768) );
  NOR2X0 U9678 ( .IN1(n9234), .IN2(n8841), .QN(n1713) );
  NAND2X0 U9679 ( .IN1(n9303), .IN2(CRC_OUT_2_14), .QN(n9767) );
  NAND4X0 U9680 ( .IN1(n9774), .IN2(n9775), .IN3(n9776), .IN4(n9777), .QN(
        WX9727) );
  NAND2X0 U9681 ( .IN1(n9099), .IN2(n9778), .QN(n9777) );
  NAND2X0 U9682 ( .IN1(n9328), .IN2(n9779), .QN(n9776) );
  NAND2X0 U9683 ( .IN1(n1712), .IN2(n9272), .QN(n9775) );
  NOR2X0 U9684 ( .IN1(n9234), .IN2(n8842), .QN(n1712) );
  NAND2X0 U9685 ( .IN1(n9303), .IN2(CRC_OUT_2_15), .QN(n9774) );
  NAND4X0 U9686 ( .IN1(n9780), .IN2(n9781), .IN3(n9782), .IN4(n9783), .QN(
        WX9725) );
  NAND2X0 U9687 ( .IN1(n9784), .IN2(n9785), .QN(n9783) );
  NAND3X0 U9688 ( .IN1(n9786), .IN2(n9787), .IN3(n9788), .QN(n9784) );
  NAND2X0 U9689 ( .IN1(n9328), .IN2(n9789), .QN(n9788) );
  NAND2X0 U9690 ( .IN1(n9083), .IN2(n8246), .QN(n9787) );
  NAND2X0 U9691 ( .IN1(n9077), .IN2(n16147), .QN(n9786) );
  NAND2X0 U9692 ( .IN1(n9792), .IN2(n9110), .QN(n9782) );
  NAND2X0 U9693 ( .IN1(n1711), .IN2(n9273), .QN(n9781) );
  NOR2X0 U9694 ( .IN1(n9235), .IN2(n8843), .QN(n1711) );
  NAND2X0 U9695 ( .IN1(n9303), .IN2(CRC_OUT_2_16), .QN(n9780) );
  NAND4X0 U9696 ( .IN1(n9793), .IN2(n9794), .IN3(n9795), .IN4(n9796), .QN(
        WX9723) );
  NAND2X0 U9697 ( .IN1(n9797), .IN2(n9798), .QN(n9796) );
  NAND2X0 U9698 ( .IN1(n9799), .IN2(n9800), .QN(n9797) );
  NAND2X0 U9699 ( .IN1(n9099), .IN2(n9801), .QN(n9800) );
  NAND2X0 U9700 ( .IN1(n9099), .IN2(n8305), .QN(n9799) );
  NAND2X0 U9701 ( .IN1(n9802), .IN2(n9803), .QN(n9795) );
  NAND3X0 U9702 ( .IN1(n9804), .IN2(n9805), .IN3(n9806), .QN(n9802) );
  NAND2X0 U9703 ( .IN1(n9328), .IN2(n9807), .QN(n9806) );
  NAND2X0 U9704 ( .IN1(n9082), .IN2(n8247), .QN(n9805) );
  NAND2X0 U9705 ( .IN1(n16146), .IN2(n9079), .QN(n9804) );
  NAND2X0 U9706 ( .IN1(n1710), .IN2(n9273), .QN(n9794) );
  NOR2X0 U9707 ( .IN1(n9235), .IN2(n8844), .QN(n1710) );
  NAND2X0 U9708 ( .IN1(n9303), .IN2(CRC_OUT_2_17), .QN(n9793) );
  NAND4X0 U9709 ( .IN1(n9808), .IN2(n9809), .IN3(n9810), .IN4(n9811), .QN(
        WX9721) );
  NAND2X0 U9710 ( .IN1(n9812), .IN2(n9813), .QN(n9811) );
  NAND3X0 U9711 ( .IN1(n9814), .IN2(n9815), .IN3(n9816), .QN(n9812) );
  NAND2X0 U9712 ( .IN1(n9328), .IN2(n9817), .QN(n9816) );
  NAND2X0 U9713 ( .IN1(n9081), .IN2(n8248), .QN(n9815) );
  NAND2X0 U9714 ( .IN1(n16145), .IN2(n9078), .QN(n9814) );
  NAND2X0 U9715 ( .IN1(n9818), .IN2(n9110), .QN(n9810) );
  NAND2X0 U9716 ( .IN1(n1709), .IN2(n9273), .QN(n9809) );
  NOR2X0 U9717 ( .IN1(n9235), .IN2(n8845), .QN(n1709) );
  NAND2X0 U9718 ( .IN1(n9303), .IN2(CRC_OUT_2_18), .QN(n9808) );
  NAND4X0 U9719 ( .IN1(n9819), .IN2(n9820), .IN3(n9821), .IN4(n9822), .QN(
        WX9719) );
  NAND2X0 U9720 ( .IN1(n9823), .IN2(n9824), .QN(n9822) );
  NAND2X0 U9721 ( .IN1(n9825), .IN2(n9826), .QN(n9823) );
  NAND2X0 U9722 ( .IN1(n9099), .IN2(n9827), .QN(n9826) );
  NAND2X0 U9723 ( .IN1(n9099), .IN2(n8307), .QN(n9825) );
  NAND2X0 U9724 ( .IN1(n9828), .IN2(n9335), .QN(n9821) );
  NAND2X0 U9725 ( .IN1(n1708), .IN2(n9273), .QN(n9820) );
  NOR2X0 U9726 ( .IN1(n9235), .IN2(n8846), .QN(n1708) );
  NAND2X0 U9727 ( .IN1(test_so88), .IN2(n9313), .QN(n9819) );
  NAND4X0 U9728 ( .IN1(n9829), .IN2(n9830), .IN3(n9831), .IN4(n9832), .QN(
        WX9717) );
  NAND2X0 U9729 ( .IN1(n9833), .IN2(n9834), .QN(n9832) );
  NAND2X0 U9730 ( .IN1(n9835), .IN2(n9836), .QN(n9833) );
  NAND2X0 U9731 ( .IN1(n9099), .IN2(n9837), .QN(n9836) );
  NAND2X0 U9732 ( .IN1(n8169), .IN2(n9110), .QN(n9835) );
  NAND2X0 U9733 ( .IN1(n9838), .IN2(n9839), .QN(n9831) );
  NAND3X0 U9734 ( .IN1(n9840), .IN2(n9841), .IN3(n9842), .QN(n9838) );
  NAND2X0 U9735 ( .IN1(n9328), .IN2(n9843), .QN(n9842) );
  NAND2X0 U9736 ( .IN1(n9081), .IN2(n8250), .QN(n9841) );
  NAND2X0 U9737 ( .IN1(n16143), .IN2(n9077), .QN(n9840) );
  NAND2X0 U9738 ( .IN1(n1707), .IN2(n9273), .QN(n9830) );
  NOR2X0 U9739 ( .IN1(n9238), .IN2(n8847), .QN(n1707) );
  NAND2X0 U9740 ( .IN1(n9304), .IN2(CRC_OUT_2_20), .QN(n9829) );
  NAND4X0 U9741 ( .IN1(n9844), .IN2(n9845), .IN3(n9846), .IN4(n9847), .QN(
        WX9715) );
  NAND2X0 U9742 ( .IN1(n9848), .IN2(n9849), .QN(n9847) );
  NAND2X0 U9743 ( .IN1(n9850), .IN2(n9851), .QN(n9848) );
  NAND2X0 U9744 ( .IN1(n9099), .IN2(n9852), .QN(n9851) );
  NAND2X0 U9745 ( .IN1(n9099), .IN2(n8310), .QN(n9850) );
  NAND2X0 U9746 ( .IN1(n9853), .IN2(n9335), .QN(n9846) );
  NAND2X0 U9747 ( .IN1(n1706), .IN2(n9273), .QN(n9845) );
  NOR2X0 U9748 ( .IN1(n9239), .IN2(n8848), .QN(n1706) );
  NAND2X0 U9749 ( .IN1(n9304), .IN2(CRC_OUT_2_21), .QN(n9844) );
  NAND4X0 U9750 ( .IN1(n9854), .IN2(n9855), .IN3(n9856), .IN4(n9857), .QN(
        WX9713) );
  NAND2X0 U9751 ( .IN1(n9858), .IN2(n9859), .QN(n9857) );
  NAND2X0 U9752 ( .IN1(n9860), .IN2(n9861), .QN(n9858) );
  NAND2X0 U9753 ( .IN1(n9099), .IN2(n9862), .QN(n9861) );
  NAND2X0 U9754 ( .IN1(n9099), .IN2(n8311), .QN(n9860) );
  NAND2X0 U9755 ( .IN1(n9863), .IN2(n9864), .QN(n9856) );
  NAND3X0 U9756 ( .IN1(n9865), .IN2(n9866), .IN3(n9867), .QN(n9863) );
  NAND2X0 U9757 ( .IN1(n9328), .IN2(n9868), .QN(n9867) );
  NAND2X0 U9758 ( .IN1(n9083), .IN2(n8252), .QN(n9866) );
  NAND2X0 U9759 ( .IN1(n16141), .IN2(n9077), .QN(n9865) );
  NAND2X0 U9760 ( .IN1(n1705), .IN2(n9273), .QN(n9855) );
  NOR2X0 U9761 ( .IN1(n9061), .IN2(n9155), .QN(n1705) );
  NAND2X0 U9762 ( .IN1(n9304), .IN2(CRC_OUT_2_22), .QN(n9854) );
  NAND4X0 U9763 ( .IN1(n9869), .IN2(n9870), .IN3(n9871), .IN4(n9872), .QN(
        WX9711) );
  NAND2X0 U9764 ( .IN1(n9873), .IN2(n9874), .QN(n9872) );
  NAND2X0 U9765 ( .IN1(n9875), .IN2(n9876), .QN(n9873) );
  NAND2X0 U9766 ( .IN1(n9099), .IN2(n9877), .QN(n9876) );
  NAND2X0 U9767 ( .IN1(n9099), .IN2(n8312), .QN(n9875) );
  NAND2X0 U9768 ( .IN1(n9878), .IN2(n9335), .QN(n9871) );
  NAND2X0 U9769 ( .IN1(n1704), .IN2(n9273), .QN(n9870) );
  NOR2X0 U9770 ( .IN1(n9239), .IN2(n8849), .QN(n1704) );
  NAND2X0 U9771 ( .IN1(n9304), .IN2(CRC_OUT_2_23), .QN(n9869) );
  NAND4X0 U9772 ( .IN1(n9879), .IN2(n9880), .IN3(n9881), .IN4(n9882), .QN(
        WX9709) );
  NAND2X0 U9773 ( .IN1(n9883), .IN2(n9884), .QN(n9882) );
  NAND2X0 U9774 ( .IN1(n9885), .IN2(n9886), .QN(n9883) );
  NAND2X0 U9775 ( .IN1(n9099), .IN2(n9887), .QN(n9886) );
  NAND2X0 U9776 ( .IN1(n9099), .IN2(n8313), .QN(n9885) );
  NAND2X0 U9777 ( .IN1(n9888), .IN2(n9889), .QN(n9881) );
  NAND3X0 U9778 ( .IN1(n9890), .IN2(n9891), .IN3(n9892), .QN(n9888) );
  NAND2X0 U9779 ( .IN1(n9328), .IN2(n9893), .QN(n9892) );
  NAND2X0 U9780 ( .IN1(n9082), .IN2(n8254), .QN(n9891) );
  NAND2X0 U9781 ( .IN1(n16139), .IN2(n9079), .QN(n9890) );
  NAND2X0 U9782 ( .IN1(n1703), .IN2(n9273), .QN(n9880) );
  NOR2X0 U9783 ( .IN1(n9239), .IN2(n8850), .QN(n1703) );
  NAND2X0 U9784 ( .IN1(n9304), .IN2(CRC_OUT_2_24), .QN(n9879) );
  NAND4X0 U9785 ( .IN1(n9894), .IN2(n9895), .IN3(n9896), .IN4(n9897), .QN(
        WX9707) );
  NAND2X0 U9786 ( .IN1(n9898), .IN2(n9899), .QN(n9897) );
  NAND2X0 U9787 ( .IN1(n9900), .IN2(n9901), .QN(n9898) );
  NAND2X0 U9788 ( .IN1(n9099), .IN2(n9902), .QN(n9901) );
  NAND2X0 U9789 ( .IN1(n9099), .IN2(n8314), .QN(n9900) );
  NAND2X0 U9790 ( .IN1(n9903), .IN2(n9904), .QN(n9896) );
  NAND3X0 U9791 ( .IN1(n9905), .IN2(n9906), .IN3(n9907), .QN(n9903) );
  NAND2X0 U9792 ( .IN1(n9328), .IN2(n9908), .QN(n9907) );
  NAND2X0 U9793 ( .IN1(n9791), .IN2(WX11193), .QN(n9906) );
  NAND2X0 U9794 ( .IN1(n9081), .IN2(n8139), .QN(n9905) );
  NAND2X0 U9795 ( .IN1(n1702), .IN2(n9273), .QN(n9895) );
  NOR2X0 U9796 ( .IN1(n9239), .IN2(n8851), .QN(n1702) );
  NAND2X0 U9797 ( .IN1(n9304), .IN2(CRC_OUT_2_25), .QN(n9894) );
  NAND4X0 U9798 ( .IN1(n9909), .IN2(n9910), .IN3(n9911), .IN4(n9912), .QN(
        WX9705) );
  NAND2X0 U9799 ( .IN1(n9913), .IN2(n9914), .QN(n9912) );
  NAND2X0 U9800 ( .IN1(n9915), .IN2(n9916), .QN(n9913) );
  NAND2X0 U9801 ( .IN1(n9098), .IN2(n9917), .QN(n9916) );
  NAND2X0 U9802 ( .IN1(n9098), .IN2(n8315), .QN(n9915) );
  NAND2X0 U9803 ( .IN1(n9918), .IN2(n9919), .QN(n9911) );
  NAND3X0 U9804 ( .IN1(n9920), .IN2(n9921), .IN3(n9922), .QN(n9918) );
  NAND2X0 U9805 ( .IN1(n9329), .IN2(n9923), .QN(n9922) );
  NAND2X0 U9806 ( .IN1(n9790), .IN2(n8257), .QN(n9921) );
  NAND2X0 U9807 ( .IN1(n16138), .IN2(n9078), .QN(n9920) );
  NAND2X0 U9808 ( .IN1(n1701), .IN2(n9273), .QN(n9910) );
  NOR2X0 U9809 ( .IN1(n9239), .IN2(n8852), .QN(n1701) );
  NAND2X0 U9810 ( .IN1(n9304), .IN2(CRC_OUT_2_26), .QN(n9909) );
  NAND4X0 U9811 ( .IN1(n9924), .IN2(n9925), .IN3(n9926), .IN4(n9927), .QN(
        WX9703) );
  NAND2X0 U9812 ( .IN1(n9928), .IN2(n9929), .QN(n9927) );
  NAND2X0 U9813 ( .IN1(n9930), .IN2(n9931), .QN(n9928) );
  NAND2X0 U9814 ( .IN1(n9098), .IN2(n9932), .QN(n9931) );
  NAND2X0 U9815 ( .IN1(n9098), .IN2(n8316), .QN(n9930) );
  NAND2X0 U9816 ( .IN1(n9933), .IN2(n9934), .QN(n9926) );
  NAND3X0 U9817 ( .IN1(n9935), .IN2(n9936), .IN3(n9937), .QN(n9933) );
  NAND2X0 U9818 ( .IN1(n9329), .IN2(n9938), .QN(n9937) );
  NAND2X0 U9819 ( .IN1(n9083), .IN2(n8258), .QN(n9936) );
  NAND2X0 U9820 ( .IN1(n16137), .IN2(n9077), .QN(n9935) );
  NAND2X0 U9821 ( .IN1(n1700), .IN2(n9273), .QN(n9925) );
  NOR2X0 U9822 ( .IN1(n9239), .IN2(n8853), .QN(n1700) );
  NAND2X0 U9823 ( .IN1(n9304), .IN2(CRC_OUT_2_27), .QN(n9924) );
  NAND4X0 U9824 ( .IN1(n9939), .IN2(n9940), .IN3(n9941), .IN4(n9942), .QN(
        WX9701) );
  NAND2X0 U9825 ( .IN1(n9943), .IN2(n9944), .QN(n9942) );
  NAND2X0 U9826 ( .IN1(n9945), .IN2(n9946), .QN(n9943) );
  NAND2X0 U9827 ( .IN1(n9098), .IN2(n9947), .QN(n9946) );
  NAND2X0 U9828 ( .IN1(n9098), .IN2(n8317), .QN(n9945) );
  NAND2X0 U9829 ( .IN1(n9948), .IN2(n9949), .QN(n9941) );
  NAND3X0 U9830 ( .IN1(n9950), .IN2(n9951), .IN3(n9952), .QN(n9948) );
  NAND2X0 U9831 ( .IN1(n9329), .IN2(n9953), .QN(n9952) );
  NAND2X0 U9832 ( .IN1(n9082), .IN2(n8259), .QN(n9951) );
  NAND2X0 U9833 ( .IN1(n16136), .IN2(n9791), .QN(n9950) );
  NAND2X0 U9834 ( .IN1(n1699), .IN2(n9273), .QN(n9940) );
  NOR2X0 U9835 ( .IN1(n9239), .IN2(n8854), .QN(n1699) );
  NAND2X0 U9836 ( .IN1(n9304), .IN2(CRC_OUT_2_28), .QN(n9939) );
  NAND4X0 U9837 ( .IN1(n9954), .IN2(n9955), .IN3(n9956), .IN4(n9957), .QN(
        WX9699) );
  NAND2X0 U9838 ( .IN1(n9958), .IN2(n9959), .QN(n9957) );
  NAND2X0 U9839 ( .IN1(n9960), .IN2(n9961), .QN(n9958) );
  NAND2X0 U9840 ( .IN1(n9098), .IN2(n9962), .QN(n9961) );
  NAND2X0 U9841 ( .IN1(n9098), .IN2(n8318), .QN(n9960) );
  NAND2X0 U9842 ( .IN1(n9963), .IN2(n9964), .QN(n9956) );
  NAND3X0 U9843 ( .IN1(n9965), .IN2(n9966), .IN3(n9967), .QN(n9963) );
  NAND2X0 U9844 ( .IN1(n9329), .IN2(n9968), .QN(n9967) );
  NAND2X0 U9845 ( .IN1(n9081), .IN2(n8260), .QN(n9966) );
  NAND2X0 U9846 ( .IN1(n16135), .IN2(n9079), .QN(n9965) );
  NAND2X0 U9847 ( .IN1(n1698), .IN2(n9273), .QN(n9955) );
  NOR2X0 U9848 ( .IN1(n9240), .IN2(n8855), .QN(n1698) );
  NAND2X0 U9849 ( .IN1(n9304), .IN2(CRC_OUT_2_29), .QN(n9954) );
  NAND4X0 U9850 ( .IN1(n9969), .IN2(n9970), .IN3(n9971), .IN4(n9972), .QN(
        WX9697) );
  NAND2X0 U9851 ( .IN1(n9973), .IN2(n9974), .QN(n9972) );
  NAND2X0 U9852 ( .IN1(n9975), .IN2(n9976), .QN(n9973) );
  NAND2X0 U9853 ( .IN1(n9098), .IN2(n9977), .QN(n9976) );
  NAND2X0 U9854 ( .IN1(n9098), .IN2(n8319), .QN(n9975) );
  NAND2X0 U9855 ( .IN1(n9978), .IN2(n9979), .QN(n9971) );
  NAND3X0 U9856 ( .IN1(n9980), .IN2(n9981), .IN3(n9982), .QN(n9978) );
  NAND2X0 U9857 ( .IN1(n9329), .IN2(n9983), .QN(n9982) );
  NAND2X0 U9858 ( .IN1(n9790), .IN2(n8261), .QN(n9981) );
  NAND2X0 U9859 ( .IN1(n16134), .IN2(n9078), .QN(n9980) );
  NAND2X0 U9860 ( .IN1(n1697), .IN2(n9273), .QN(n9970) );
  NOR2X0 U9861 ( .IN1(n9240), .IN2(n8856), .QN(n1697) );
  NAND2X0 U9862 ( .IN1(n9304), .IN2(CRC_OUT_2_30), .QN(n9969) );
  NAND4X0 U9863 ( .IN1(n9984), .IN2(n9985), .IN3(n9986), .IN4(n9987), .QN(
        WX9695) );
  NAND2X0 U9864 ( .IN1(n9988), .IN2(n9989), .QN(n9987) );
  NAND3X0 U9865 ( .IN1(n9990), .IN2(n9991), .IN3(n9992), .QN(n9988) );
  NAND2X0 U9866 ( .IN1(n9329), .IN2(n9993), .QN(n9992) );
  NAND2X0 U9867 ( .IN1(n9083), .IN2(n8262), .QN(n9991) );
  NAND2X0 U9868 ( .IN1(n16133), .IN2(n9077), .QN(n9990) );
  NAND2X0 U9869 ( .IN1(n9994), .IN2(n9110), .QN(n9986) );
  NAND2X0 U9870 ( .IN1(n9304), .IN2(CRC_OUT_2_31), .QN(n9985) );
  NAND2X0 U9871 ( .IN1(n2245), .IN2(WX9536), .QN(n9984) );
  NOR2X0 U9872 ( .IN1(n9240), .IN2(WX9536), .QN(WX9597) );
  NOR3X0 U9873 ( .IN1(n9146), .IN2(n9995), .IN3(n9996), .QN(WX9084) );
  NOR2X0 U9874 ( .IN1(n8185), .IN2(CRC_OUT_3_30), .QN(n9996) );
  NOR2X0 U9875 ( .IN1(DFF_1342_n1), .IN2(WX8595), .QN(n9995) );
  NOR3X0 U9876 ( .IN1(n9146), .IN2(n9997), .IN3(n9998), .QN(WX9082) );
  NOR2X0 U9877 ( .IN1(n8186), .IN2(CRC_OUT_3_29), .QN(n9998) );
  NOR2X0 U9878 ( .IN1(DFF_1341_n1), .IN2(WX8597), .QN(n9997) );
  NOR3X0 U9879 ( .IN1(n9146), .IN2(n9999), .IN3(n10000), .QN(WX9080) );
  NOR2X0 U9880 ( .IN1(n8187), .IN2(CRC_OUT_3_28), .QN(n10000) );
  NOR2X0 U9881 ( .IN1(DFF_1340_n1), .IN2(WX8599), .QN(n9999) );
  NOR3X0 U9882 ( .IN1(n9146), .IN2(n10001), .IN3(n10002), .QN(WX9078) );
  NOR2X0 U9883 ( .IN1(n8188), .IN2(CRC_OUT_3_27), .QN(n10002) );
  NOR2X0 U9884 ( .IN1(DFF_1339_n1), .IN2(WX8601), .QN(n10001) );
  NOR3X0 U9885 ( .IN1(n9146), .IN2(n10003), .IN3(n10004), .QN(WX9076) );
  NOR2X0 U9886 ( .IN1(n8189), .IN2(CRC_OUT_3_26), .QN(n10004) );
  NOR2X0 U9887 ( .IN1(DFF_1338_n1), .IN2(WX8603), .QN(n10003) );
  NOR2X0 U9888 ( .IN1(n9240), .IN2(n10005), .QN(WX9074) );
  NOR2X0 U9889 ( .IN1(n10006), .IN2(n10007), .QN(n10005) );
  NOR2X0 U9890 ( .IN1(test_so74), .IN2(CRC_OUT_3_25), .QN(n10007) );
  NOR2X0 U9891 ( .IN1(DFF_1337_n1), .IN2(n8798), .QN(n10006) );
  NOR2X0 U9892 ( .IN1(n9240), .IN2(n10008), .QN(WX9072) );
  NOR2X0 U9893 ( .IN1(n10009), .IN2(n10010), .QN(n10008) );
  NOR2X0 U9894 ( .IN1(test_so77), .IN2(WX8607), .QN(n10010) );
  INVX0 U9895 ( .INP(n10011), .ZN(n10009) );
  NAND2X0 U9896 ( .IN1(WX8607), .IN2(test_so77), .QN(n10011) );
  NOR3X0 U9897 ( .IN1(n9146), .IN2(n10012), .IN3(n10013), .QN(WX9070) );
  NOR2X0 U9898 ( .IN1(n8191), .IN2(CRC_OUT_3_23), .QN(n10013) );
  NOR2X0 U9899 ( .IN1(DFF_1335_n1), .IN2(WX8609), .QN(n10012) );
  NOR3X0 U9900 ( .IN1(n9145), .IN2(n10014), .IN3(n10015), .QN(WX9068) );
  NOR2X0 U9901 ( .IN1(n8192), .IN2(CRC_OUT_3_22), .QN(n10015) );
  NOR2X0 U9902 ( .IN1(DFF_1334_n1), .IN2(WX8611), .QN(n10014) );
  NOR3X0 U9903 ( .IN1(n9145), .IN2(n10016), .IN3(n10017), .QN(WX9066) );
  NOR2X0 U9904 ( .IN1(n8193), .IN2(CRC_OUT_3_21), .QN(n10017) );
  NOR2X0 U9905 ( .IN1(DFF_1333_n1), .IN2(WX8613), .QN(n10016) );
  NOR3X0 U9906 ( .IN1(n9145), .IN2(n10018), .IN3(n10019), .QN(WX9064) );
  NOR2X0 U9907 ( .IN1(n8194), .IN2(CRC_OUT_3_20), .QN(n10019) );
  NOR2X0 U9908 ( .IN1(DFF_1332_n1), .IN2(WX8615), .QN(n10018) );
  NOR3X0 U9909 ( .IN1(n9145), .IN2(n10020), .IN3(n10021), .QN(WX9062) );
  NOR2X0 U9910 ( .IN1(n8195), .IN2(CRC_OUT_3_19), .QN(n10021) );
  NOR2X0 U9911 ( .IN1(DFF_1331_n1), .IN2(WX8617), .QN(n10020) );
  NOR3X0 U9912 ( .IN1(n9145), .IN2(n10022), .IN3(n10023), .QN(WX9060) );
  NOR2X0 U9913 ( .IN1(n8196), .IN2(CRC_OUT_3_18), .QN(n10023) );
  NOR2X0 U9914 ( .IN1(DFF_1330_n1), .IN2(WX8619), .QN(n10022) );
  NOR3X0 U9915 ( .IN1(n9145), .IN2(n10024), .IN3(n10025), .QN(WX9058) );
  NOR2X0 U9916 ( .IN1(n8197), .IN2(CRC_OUT_3_17), .QN(n10025) );
  NOR2X0 U9917 ( .IN1(DFF_1329_n1), .IN2(WX8621), .QN(n10024) );
  NOR3X0 U9918 ( .IN1(n9145), .IN2(n10026), .IN3(n10027), .QN(WX9056) );
  NOR2X0 U9919 ( .IN1(n8198), .IN2(CRC_OUT_3_16), .QN(n10027) );
  NOR2X0 U9920 ( .IN1(DFF_1328_n1), .IN2(WX8623), .QN(n10026) );
  NOR2X0 U9921 ( .IN1(n9240), .IN2(n10028), .QN(WX9054) );
  NOR2X0 U9922 ( .IN1(n10029), .IN2(n10030), .QN(n10028) );
  INVX0 U9923 ( .INP(n10031), .ZN(n10030) );
  NAND2X0 U9924 ( .IN1(CRC_OUT_3_15), .IN2(n10032), .QN(n10031) );
  NOR2X0 U9925 ( .IN1(n10032), .IN2(CRC_OUT_3_15), .QN(n10029) );
  NAND2X0 U9926 ( .IN1(n10033), .IN2(n10034), .QN(n10032) );
  NAND2X0 U9927 ( .IN1(n8110), .IN2(CRC_OUT_3_31), .QN(n10034) );
  NAND2X0 U9928 ( .IN1(DFF_1343_n1), .IN2(WX8625), .QN(n10033) );
  NOR3X0 U9929 ( .IN1(n9145), .IN2(n10035), .IN3(n10036), .QN(WX9052) );
  NOR2X0 U9930 ( .IN1(n8199), .IN2(CRC_OUT_3_14), .QN(n10036) );
  NOR2X0 U9931 ( .IN1(DFF_1326_n1), .IN2(WX8627), .QN(n10035) );
  NOR3X0 U9932 ( .IN1(n9145), .IN2(n10037), .IN3(n10038), .QN(WX9050) );
  NOR2X0 U9933 ( .IN1(n8200), .IN2(CRC_OUT_3_13), .QN(n10038) );
  NOR2X0 U9934 ( .IN1(DFF_1325_n1), .IN2(WX8629), .QN(n10037) );
  NOR3X0 U9935 ( .IN1(n9145), .IN2(n10039), .IN3(n10040), .QN(WX9048) );
  NOR2X0 U9936 ( .IN1(n8201), .IN2(CRC_OUT_3_12), .QN(n10040) );
  NOR2X0 U9937 ( .IN1(DFF_1324_n1), .IN2(WX8631), .QN(n10039) );
  NOR3X0 U9938 ( .IN1(n9145), .IN2(n10041), .IN3(n10042), .QN(WX9046) );
  NOR2X0 U9939 ( .IN1(n8202), .IN2(CRC_OUT_3_11), .QN(n10042) );
  NOR2X0 U9940 ( .IN1(DFF_1323_n1), .IN2(WX8633), .QN(n10041) );
  NOR2X0 U9941 ( .IN1(n9225), .IN2(n10043), .QN(WX9044) );
  NOR2X0 U9942 ( .IN1(n10044), .IN2(n10045), .QN(n10043) );
  INVX0 U9943 ( .INP(n10046), .ZN(n10045) );
  NAND2X0 U9944 ( .IN1(CRC_OUT_3_10), .IN2(n10047), .QN(n10046) );
  NOR2X0 U9945 ( .IN1(n10047), .IN2(CRC_OUT_3_10), .QN(n10044) );
  NAND2X0 U9946 ( .IN1(n10048), .IN2(n10049), .QN(n10047) );
  NAND2X0 U9947 ( .IN1(n8111), .IN2(CRC_OUT_3_31), .QN(n10049) );
  NAND2X0 U9948 ( .IN1(DFF_1343_n1), .IN2(WX8635), .QN(n10048) );
  NOR3X0 U9949 ( .IN1(n9145), .IN2(n10050), .IN3(n10051), .QN(WX9042) );
  NOR2X0 U9950 ( .IN1(n8203), .IN2(CRC_OUT_3_9), .QN(n10051) );
  NOR2X0 U9951 ( .IN1(DFF_1321_n1), .IN2(WX8637), .QN(n10050) );
  NOR2X0 U9952 ( .IN1(n9225), .IN2(n10052), .QN(WX9040) );
  NOR2X0 U9953 ( .IN1(n10053), .IN2(n10054), .QN(n10052) );
  NOR2X0 U9954 ( .IN1(test_so75), .IN2(CRC_OUT_3_8), .QN(n10054) );
  NOR2X0 U9955 ( .IN1(DFF_1320_n1), .IN2(n8790), .QN(n10053) );
  NOR2X0 U9956 ( .IN1(n9225), .IN2(n10055), .QN(WX9038) );
  NOR2X0 U9957 ( .IN1(n10056), .IN2(n10057), .QN(n10055) );
  NOR2X0 U9958 ( .IN1(test_so76), .IN2(WX8641), .QN(n10057) );
  INVX0 U9959 ( .INP(n10058), .ZN(n10056) );
  NAND2X0 U9960 ( .IN1(WX8641), .IN2(test_so76), .QN(n10058) );
  NOR3X0 U9961 ( .IN1(n9144), .IN2(n10059), .IN3(n10060), .QN(WX9036) );
  NOR2X0 U9962 ( .IN1(n8205), .IN2(CRC_OUT_3_6), .QN(n10060) );
  NOR2X0 U9963 ( .IN1(DFF_1318_n1), .IN2(WX8643), .QN(n10059) );
  NOR3X0 U9964 ( .IN1(n9144), .IN2(n10061), .IN3(n10062), .QN(WX9034) );
  NOR2X0 U9965 ( .IN1(n8206), .IN2(CRC_OUT_3_5), .QN(n10062) );
  NOR2X0 U9966 ( .IN1(DFF_1317_n1), .IN2(WX8645), .QN(n10061) );
  NOR3X0 U9967 ( .IN1(n9144), .IN2(n10063), .IN3(n10064), .QN(WX9032) );
  NOR2X0 U9968 ( .IN1(n8207), .IN2(CRC_OUT_3_4), .QN(n10064) );
  NOR2X0 U9969 ( .IN1(DFF_1316_n1), .IN2(WX8647), .QN(n10063) );
  NOR2X0 U9970 ( .IN1(n9225), .IN2(n10065), .QN(WX9030) );
  NOR2X0 U9971 ( .IN1(n10066), .IN2(n10067), .QN(n10065) );
  INVX0 U9972 ( .INP(n10068), .ZN(n10067) );
  NAND2X0 U9973 ( .IN1(CRC_OUT_3_3), .IN2(n10069), .QN(n10068) );
  NOR2X0 U9974 ( .IN1(n10069), .IN2(CRC_OUT_3_3), .QN(n10066) );
  NAND2X0 U9975 ( .IN1(n10070), .IN2(n10071), .QN(n10069) );
  NAND2X0 U9976 ( .IN1(n8112), .IN2(CRC_OUT_3_31), .QN(n10071) );
  NAND2X0 U9977 ( .IN1(DFF_1343_n1), .IN2(WX8649), .QN(n10070) );
  NOR3X0 U9978 ( .IN1(n9144), .IN2(n10072), .IN3(n10073), .QN(WX9028) );
  NOR2X0 U9979 ( .IN1(n8208), .IN2(CRC_OUT_3_2), .QN(n10073) );
  NOR2X0 U9980 ( .IN1(DFF_1314_n1), .IN2(WX8651), .QN(n10072) );
  NOR3X0 U9981 ( .IN1(n9144), .IN2(n10074), .IN3(n10075), .QN(WX9026) );
  NOR2X0 U9982 ( .IN1(n8209), .IN2(CRC_OUT_3_1), .QN(n10075) );
  NOR2X0 U9983 ( .IN1(DFF_1313_n1), .IN2(WX8653), .QN(n10074) );
  NOR3X0 U9984 ( .IN1(n9144), .IN2(n10076), .IN3(n10077), .QN(WX9024) );
  NOR2X0 U9985 ( .IN1(n8210), .IN2(CRC_OUT_3_0), .QN(n10077) );
  NOR2X0 U9986 ( .IN1(DFF_1312_n1), .IN2(WX8655), .QN(n10076) );
  NOR3X0 U9987 ( .IN1(n9144), .IN2(n10078), .IN3(n10079), .QN(WX9022) );
  NOR2X0 U9988 ( .IN1(n8127), .IN2(CRC_OUT_3_31), .QN(n10079) );
  NOR2X0 U9989 ( .IN1(DFF_1343_n1), .IN2(WX8657), .QN(n10078) );
  NOR2X0 U9990 ( .IN1(n16117), .IN2(n9155), .QN(WX8496) );
  NOR2X0 U9991 ( .IN1(n16116), .IN2(n9155), .QN(WX8494) );
  NOR2X0 U9992 ( .IN1(n16115), .IN2(n9156), .QN(WX8492) );
  NOR2X0 U9993 ( .IN1(n16114), .IN2(n9158), .QN(WX8490) );
  NOR2X0 U9994 ( .IN1(n16113), .IN2(n9155), .QN(WX8488) );
  NOR2X0 U9995 ( .IN1(n16112), .IN2(n9156), .QN(WX8486) );
  NOR2X0 U9996 ( .IN1(n16111), .IN2(n9155), .QN(WX8484) );
  NOR2X0 U9997 ( .IN1(n16110), .IN2(n9156), .QN(WX8482) );
  NOR2X0 U9998 ( .IN1(n16109), .IN2(n9156), .QN(WX8480) );
  NOR2X0 U9999 ( .IN1(n16108), .IN2(n9155), .QN(WX8478) );
  NOR2X0 U10000 ( .IN1(n16107), .IN2(n9155), .QN(WX8476) );
  NOR2X0 U10001 ( .IN1(n16106), .IN2(n9156), .QN(WX8474) );
  NOR2X0 U10002 ( .IN1(n16105), .IN2(n9155), .QN(WX8472) );
  NOR2X0 U10003 ( .IN1(n16104), .IN2(n9155), .QN(WX8470) );
  NOR2X0 U10004 ( .IN1(n16103), .IN2(n9156), .QN(WX8468) );
  NOR2X0 U10005 ( .IN1(n16102), .IN2(n9156), .QN(WX8466) );
  NAND4X0 U10006 ( .IN1(n10080), .IN2(n10081), .IN3(n10082), .IN4(n10083), 
        .QN(WX8464) );
  NAND2X0 U10007 ( .IN1(n9329), .IN2(n9681), .QN(n10083) );
  NAND2X0 U10008 ( .IN1(n10084), .IN2(n10085), .QN(n9681) );
  INVX0 U10009 ( .INP(n10086), .ZN(n10085) );
  NOR2X0 U10010 ( .IN1(n10087), .IN2(n10088), .QN(n10086) );
  NAND2X0 U10011 ( .IN1(n10088), .IN2(n10087), .QN(n10084) );
  NOR2X0 U10012 ( .IN1(n10089), .IN2(n10090), .QN(n10087) );
  NOR2X0 U10013 ( .IN1(WX9950), .IN2(n7884), .QN(n10090) );
  INVX0 U10014 ( .INP(n10091), .ZN(n10089) );
  NAND2X0 U10015 ( .IN1(n7884), .IN2(WX9950), .QN(n10091) );
  NAND2X0 U10016 ( .IN1(n10092), .IN2(n10093), .QN(n10088) );
  NAND2X0 U10017 ( .IN1(n7883), .IN2(WX9822), .QN(n10093) );
  INVX0 U10018 ( .INP(n10094), .ZN(n10092) );
  NOR2X0 U10019 ( .IN1(WX9822), .IN2(n7883), .QN(n10094) );
  NAND2X0 U10020 ( .IN1(n9098), .IN2(n10095), .QN(n10082) );
  NAND2X0 U10021 ( .IN1(n1485), .IN2(n9273), .QN(n10081) );
  NOR2X0 U10022 ( .IN1(n9062), .IN2(n9155), .QN(n1485) );
  NAND2X0 U10023 ( .IN1(n9305), .IN2(CRC_OUT_3_0), .QN(n10080) );
  NAND4X0 U10024 ( .IN1(n10096), .IN2(n10097), .IN3(n10098), .IN4(n10099), 
        .QN(WX8462) );
  NAND3X0 U10025 ( .IN1(n9687), .IN2(n9688), .IN3(n9321), .QN(n10099) );
  NAND3X0 U10026 ( .IN1(n10100), .IN2(n10101), .IN3(n10102), .QN(n9688) );
  INVX0 U10027 ( .INP(n10103), .ZN(n10102) );
  NAND2X0 U10028 ( .IN1(n10103), .IN2(n10104), .QN(n9687) );
  NAND2X0 U10029 ( .IN1(n10100), .IN2(n10101), .QN(n10104) );
  NAND2X0 U10030 ( .IN1(n8184), .IN2(WX9884), .QN(n10101) );
  NAND2X0 U10031 ( .IN1(n7886), .IN2(WX9948), .QN(n10100) );
  NOR2X0 U10032 ( .IN1(n10105), .IN2(n10106), .QN(n10103) );
  INVX0 U10033 ( .INP(n10107), .ZN(n10106) );
  NAND2X0 U10034 ( .IN1(test_so83), .IN2(WX9756), .QN(n10107) );
  NOR2X0 U10035 ( .IN1(WX9756), .IN2(test_so83), .QN(n10105) );
  NAND2X0 U10036 ( .IN1(n9098), .IN2(n10108), .QN(n10098) );
  NAND2X0 U10037 ( .IN1(n1484), .IN2(n9273), .QN(n10097) );
  NOR2X0 U10038 ( .IN1(n9227), .IN2(n8857), .QN(n1484) );
  NAND2X0 U10039 ( .IN1(n9305), .IN2(CRC_OUT_3_1), .QN(n10096) );
  NAND4X0 U10040 ( .IN1(n10109), .IN2(n10110), .IN3(n10111), .IN4(n10112), 
        .QN(WX8460) );
  NAND2X0 U10041 ( .IN1(n9329), .IN2(n9696), .QN(n10112) );
  NAND2X0 U10042 ( .IN1(n10113), .IN2(n10114), .QN(n9696) );
  INVX0 U10043 ( .INP(n10115), .ZN(n10114) );
  NOR2X0 U10044 ( .IN1(n10116), .IN2(n10117), .QN(n10115) );
  NAND2X0 U10045 ( .IN1(n10117), .IN2(n10116), .QN(n10113) );
  NOR2X0 U10046 ( .IN1(n10118), .IN2(n10119), .QN(n10116) );
  NOR2X0 U10047 ( .IN1(WX9946), .IN2(n7888), .QN(n10119) );
  INVX0 U10048 ( .INP(n10120), .ZN(n10118) );
  NAND2X0 U10049 ( .IN1(n7888), .IN2(WX9946), .QN(n10120) );
  NAND2X0 U10050 ( .IN1(n10121), .IN2(n10122), .QN(n10117) );
  NAND2X0 U10051 ( .IN1(n7887), .IN2(WX9818), .QN(n10122) );
  INVX0 U10052 ( .INP(n10123), .ZN(n10121) );
  NOR2X0 U10053 ( .IN1(WX9818), .IN2(n7887), .QN(n10123) );
  NAND2X0 U10054 ( .IN1(n9098), .IN2(n10124), .QN(n10111) );
  NAND2X0 U10055 ( .IN1(n1483), .IN2(n9274), .QN(n10110) );
  NOR2X0 U10056 ( .IN1(n9227), .IN2(n8858), .QN(n1483) );
  NAND2X0 U10057 ( .IN1(n9305), .IN2(CRC_OUT_3_2), .QN(n10109) );
  NAND4X0 U10058 ( .IN1(n10125), .IN2(n10126), .IN3(n10127), .IN4(n10128), 
        .QN(WX8458) );
  NAND3X0 U10059 ( .IN1(n9701), .IN2(n9702), .IN3(n9320), .QN(n10128) );
  NAND3X0 U10060 ( .IN1(n10129), .IN2(n10130), .IN3(n10131), .QN(n9702) );
  INVX0 U10061 ( .INP(n10132), .ZN(n10131) );
  NAND2X0 U10062 ( .IN1(n10132), .IN2(n10133), .QN(n9701) );
  NAND2X0 U10063 ( .IN1(n10129), .IN2(n10130), .QN(n10133) );
  NAND2X0 U10064 ( .IN1(n8182), .IN2(WX9816), .QN(n10130) );
  NAND2X0 U10065 ( .IN1(n3569), .IN2(WX9944), .QN(n10129) );
  NOR2X0 U10066 ( .IN1(n10134), .IN2(n10135), .QN(n10132) );
  INVX0 U10067 ( .INP(n10136), .ZN(n10135) );
  NAND2X0 U10068 ( .IN1(test_so81), .IN2(WX9880), .QN(n10136) );
  NOR2X0 U10069 ( .IN1(WX9880), .IN2(test_so81), .QN(n10134) );
  NAND2X0 U10070 ( .IN1(n9098), .IN2(n10137), .QN(n10127) );
  NAND2X0 U10071 ( .IN1(n1482), .IN2(n9274), .QN(n10126) );
  NOR2X0 U10072 ( .IN1(n9227), .IN2(n8859), .QN(n1482) );
  NAND2X0 U10073 ( .IN1(n9305), .IN2(CRC_OUT_3_3), .QN(n10125) );
  NAND4X0 U10074 ( .IN1(n10138), .IN2(n10139), .IN3(n10140), .IN4(n10141), 
        .QN(WX8456) );
  NAND2X0 U10075 ( .IN1(n9329), .IN2(n9710), .QN(n10141) );
  NAND2X0 U10076 ( .IN1(n10142), .IN2(n10143), .QN(n9710) );
  INVX0 U10077 ( .INP(n10144), .ZN(n10143) );
  NOR2X0 U10078 ( .IN1(n10145), .IN2(n10146), .QN(n10144) );
  NAND2X0 U10079 ( .IN1(n10146), .IN2(n10145), .QN(n10142) );
  NOR2X0 U10080 ( .IN1(n10147), .IN2(n10148), .QN(n10145) );
  NOR2X0 U10081 ( .IN1(WX9942), .IN2(n7891), .QN(n10148) );
  INVX0 U10082 ( .INP(n10149), .ZN(n10147) );
  NAND2X0 U10083 ( .IN1(n7891), .IN2(WX9942), .QN(n10149) );
  NAND2X0 U10084 ( .IN1(n10150), .IN2(n10151), .QN(n10146) );
  NAND2X0 U10085 ( .IN1(n7890), .IN2(WX9814), .QN(n10151) );
  INVX0 U10086 ( .INP(n10152), .ZN(n10150) );
  NOR2X0 U10087 ( .IN1(WX9814), .IN2(n7890), .QN(n10152) );
  NAND2X0 U10088 ( .IN1(n9098), .IN2(n10153), .QN(n10140) );
  NAND2X0 U10089 ( .IN1(n1481), .IN2(n9274), .QN(n10139) );
  NOR2X0 U10090 ( .IN1(n9227), .IN2(n8860), .QN(n1481) );
  NAND2X0 U10091 ( .IN1(n9305), .IN2(CRC_OUT_3_4), .QN(n10138) );
  NAND4X0 U10092 ( .IN1(n10154), .IN2(n10155), .IN3(n10156), .IN4(n10157), 
        .QN(WX8454) );
  NAND2X0 U10093 ( .IN1(n9329), .IN2(n9715), .QN(n10157) );
  NAND2X0 U10094 ( .IN1(n10158), .IN2(n10159), .QN(n9715) );
  INVX0 U10095 ( .INP(n10160), .ZN(n10159) );
  NOR2X0 U10096 ( .IN1(n10161), .IN2(n10162), .QN(n10160) );
  NAND2X0 U10097 ( .IN1(n10162), .IN2(n10161), .QN(n10158) );
  NOR2X0 U10098 ( .IN1(n10163), .IN2(n10164), .QN(n10161) );
  NOR2X0 U10099 ( .IN1(WX9940), .IN2(n7893), .QN(n10164) );
  INVX0 U10100 ( .INP(n10165), .ZN(n10163) );
  NAND2X0 U10101 ( .IN1(n7893), .IN2(WX9940), .QN(n10165) );
  NAND2X0 U10102 ( .IN1(n10166), .IN2(n10167), .QN(n10162) );
  NAND2X0 U10103 ( .IN1(n7892), .IN2(WX9812), .QN(n10167) );
  INVX0 U10104 ( .INP(n10168), .ZN(n10166) );
  NOR2X0 U10105 ( .IN1(WX9812), .IN2(n7892), .QN(n10168) );
  NAND2X0 U10106 ( .IN1(n9098), .IN2(n10169), .QN(n10156) );
  NAND2X0 U10107 ( .IN1(n1480), .IN2(n9274), .QN(n10155) );
  NOR2X0 U10108 ( .IN1(n9227), .IN2(n8861), .QN(n1480) );
  NAND2X0 U10109 ( .IN1(n9305), .IN2(CRC_OUT_3_5), .QN(n10154) );
  NAND4X0 U10110 ( .IN1(n10170), .IN2(n10171), .IN3(n10172), .IN4(n10173), 
        .QN(WX8452) );
  NAND2X0 U10111 ( .IN1(n9329), .IN2(n9723), .QN(n10173) );
  NAND2X0 U10112 ( .IN1(n10174), .IN2(n10175), .QN(n9723) );
  INVX0 U10113 ( .INP(n10176), .ZN(n10175) );
  NOR2X0 U10114 ( .IN1(n10177), .IN2(n10178), .QN(n10176) );
  NAND2X0 U10115 ( .IN1(n10178), .IN2(n10177), .QN(n10174) );
  NOR2X0 U10116 ( .IN1(n10179), .IN2(n10180), .QN(n10177) );
  NOR2X0 U10117 ( .IN1(WX9938), .IN2(n7895), .QN(n10180) );
  INVX0 U10118 ( .INP(n10181), .ZN(n10179) );
  NAND2X0 U10119 ( .IN1(n7895), .IN2(WX9938), .QN(n10181) );
  NAND2X0 U10120 ( .IN1(n10182), .IN2(n10183), .QN(n10178) );
  NAND2X0 U10121 ( .IN1(n7894), .IN2(WX9810), .QN(n10183) );
  INVX0 U10122 ( .INP(n10184), .ZN(n10182) );
  NOR2X0 U10123 ( .IN1(WX9810), .IN2(n7894), .QN(n10184) );
  NAND2X0 U10124 ( .IN1(n9098), .IN2(n10185), .QN(n10172) );
  NAND2X0 U10125 ( .IN1(n1479), .IN2(n9274), .QN(n10171) );
  NOR2X0 U10126 ( .IN1(n9227), .IN2(n8862), .QN(n1479) );
  NAND2X0 U10127 ( .IN1(n9305), .IN2(CRC_OUT_3_6), .QN(n10170) );
  NAND4X0 U10128 ( .IN1(n10186), .IN2(n10187), .IN3(n10188), .IN4(n10189), 
        .QN(WX8450) );
  NAND2X0 U10129 ( .IN1(n9329), .IN2(n9728), .QN(n10189) );
  NAND2X0 U10130 ( .IN1(n10190), .IN2(n10191), .QN(n9728) );
  INVX0 U10131 ( .INP(n10192), .ZN(n10191) );
  NOR2X0 U10132 ( .IN1(n10193), .IN2(n10194), .QN(n10192) );
  NAND2X0 U10133 ( .IN1(n10194), .IN2(n10193), .QN(n10190) );
  NOR2X0 U10134 ( .IN1(n10195), .IN2(n10196), .QN(n10193) );
  NOR2X0 U10135 ( .IN1(WX9936), .IN2(n7897), .QN(n10196) );
  INVX0 U10136 ( .INP(n10197), .ZN(n10195) );
  NAND2X0 U10137 ( .IN1(n7897), .IN2(WX9936), .QN(n10197) );
  NAND2X0 U10138 ( .IN1(n10198), .IN2(n10199), .QN(n10194) );
  NAND2X0 U10139 ( .IN1(n7896), .IN2(WX9808), .QN(n10199) );
  INVX0 U10140 ( .INP(n10200), .ZN(n10198) );
  NOR2X0 U10141 ( .IN1(WX9808), .IN2(n7896), .QN(n10200) );
  NAND2X0 U10142 ( .IN1(n9098), .IN2(n10201), .QN(n10188) );
  NAND2X0 U10143 ( .IN1(n1478), .IN2(n9274), .QN(n10187) );
  NOR2X0 U10144 ( .IN1(n9227), .IN2(n8863), .QN(n1478) );
  NAND2X0 U10145 ( .IN1(test_so76), .IN2(n9314), .QN(n10186) );
  NAND4X0 U10146 ( .IN1(n10202), .IN2(n10203), .IN3(n10204), .IN4(n10205), 
        .QN(WX8448) );
  NAND2X0 U10147 ( .IN1(n9329), .IN2(n9736), .QN(n10205) );
  NAND2X0 U10148 ( .IN1(n10206), .IN2(n10207), .QN(n9736) );
  INVX0 U10149 ( .INP(n10208), .ZN(n10207) );
  NOR2X0 U10150 ( .IN1(n10209), .IN2(n10210), .QN(n10208) );
  NAND2X0 U10151 ( .IN1(n10210), .IN2(n10209), .QN(n10206) );
  NOR2X0 U10152 ( .IN1(n10211), .IN2(n10212), .QN(n10209) );
  NOR2X0 U10153 ( .IN1(WX9934), .IN2(n7899), .QN(n10212) );
  INVX0 U10154 ( .INP(n10213), .ZN(n10211) );
  NAND2X0 U10155 ( .IN1(n7899), .IN2(WX9934), .QN(n10213) );
  NAND2X0 U10156 ( .IN1(n10214), .IN2(n10215), .QN(n10210) );
  NAND2X0 U10157 ( .IN1(n7898), .IN2(WX9806), .QN(n10215) );
  INVX0 U10158 ( .INP(n10216), .ZN(n10214) );
  NOR2X0 U10159 ( .IN1(WX9806), .IN2(n7898), .QN(n10216) );
  NAND2X0 U10160 ( .IN1(n9097), .IN2(n10217), .QN(n10204) );
  NAND2X0 U10161 ( .IN1(n1477), .IN2(n9274), .QN(n10203) );
  NOR2X0 U10162 ( .IN1(n9227), .IN2(n8864), .QN(n1477) );
  NAND2X0 U10163 ( .IN1(n9305), .IN2(CRC_OUT_3_8), .QN(n10202) );
  NAND4X0 U10164 ( .IN1(n10218), .IN2(n10219), .IN3(n10220), .IN4(n10221), 
        .QN(WX8446) );
  NAND3X0 U10165 ( .IN1(n10222), .IN2(n10223), .IN3(n9091), .QN(n10221) );
  NAND2X0 U10166 ( .IN1(n9329), .IN2(n9741), .QN(n10220) );
  NAND2X0 U10167 ( .IN1(n10224), .IN2(n10225), .QN(n9741) );
  INVX0 U10168 ( .INP(n10226), .ZN(n10225) );
  NOR2X0 U10169 ( .IN1(n10227), .IN2(n10228), .QN(n10226) );
  NAND2X0 U10170 ( .IN1(n10228), .IN2(n10227), .QN(n10224) );
  NOR2X0 U10171 ( .IN1(n10229), .IN2(n10230), .QN(n10227) );
  NOR2X0 U10172 ( .IN1(WX9932), .IN2(n7901), .QN(n10230) );
  INVX0 U10173 ( .INP(n10231), .ZN(n10229) );
  NAND2X0 U10174 ( .IN1(n7901), .IN2(WX9932), .QN(n10231) );
  NAND2X0 U10175 ( .IN1(n10232), .IN2(n10233), .QN(n10228) );
  NAND2X0 U10176 ( .IN1(n7900), .IN2(WX9804), .QN(n10233) );
  INVX0 U10177 ( .INP(n10234), .ZN(n10232) );
  NOR2X0 U10178 ( .IN1(WX9804), .IN2(n7900), .QN(n10234) );
  NAND2X0 U10179 ( .IN1(n1476), .IN2(n9274), .QN(n10219) );
  NOR2X0 U10180 ( .IN1(n9228), .IN2(n8865), .QN(n1476) );
  NAND2X0 U10181 ( .IN1(n9305), .IN2(CRC_OUT_3_9), .QN(n10218) );
  NAND4X0 U10182 ( .IN1(n10235), .IN2(n10236), .IN3(n10237), .IN4(n10238), 
        .QN(WX8444) );
  NAND2X0 U10183 ( .IN1(n9329), .IN2(n9747), .QN(n10238) );
  NAND2X0 U10184 ( .IN1(n10239), .IN2(n10240), .QN(n9747) );
  INVX0 U10185 ( .INP(n10241), .ZN(n10240) );
  NOR2X0 U10186 ( .IN1(n10242), .IN2(n10243), .QN(n10241) );
  NAND2X0 U10187 ( .IN1(n10243), .IN2(n10242), .QN(n10239) );
  NOR2X0 U10188 ( .IN1(n10244), .IN2(n10245), .QN(n10242) );
  NOR2X0 U10189 ( .IN1(WX9930), .IN2(n7903), .QN(n10245) );
  INVX0 U10190 ( .INP(n10246), .ZN(n10244) );
  NAND2X0 U10191 ( .IN1(n7903), .IN2(WX9930), .QN(n10246) );
  NAND2X0 U10192 ( .IN1(n10247), .IN2(n10248), .QN(n10243) );
  NAND2X0 U10193 ( .IN1(n7902), .IN2(WX9802), .QN(n10248) );
  INVX0 U10194 ( .INP(n10249), .ZN(n10247) );
  NOR2X0 U10195 ( .IN1(WX9802), .IN2(n7902), .QN(n10249) );
  NAND2X0 U10196 ( .IN1(n9097), .IN2(n10250), .QN(n10237) );
  NAND2X0 U10197 ( .IN1(n1475), .IN2(n9274), .QN(n10236) );
  NOR2X0 U10198 ( .IN1(n9229), .IN2(n8866), .QN(n1475) );
  NAND2X0 U10199 ( .IN1(n9305), .IN2(CRC_OUT_3_10), .QN(n10235) );
  NAND4X0 U10200 ( .IN1(n10251), .IN2(n10252), .IN3(n10253), .IN4(n10254), 
        .QN(WX8442) );
  NAND3X0 U10201 ( .IN1(n10255), .IN2(n10256), .IN3(n9090), .QN(n10254) );
  NAND2X0 U10202 ( .IN1(n9329), .IN2(n9753), .QN(n10253) );
  NAND2X0 U10203 ( .IN1(n10257), .IN2(n10258), .QN(n9753) );
  INVX0 U10204 ( .INP(n10259), .ZN(n10258) );
  NOR2X0 U10205 ( .IN1(n10260), .IN2(n10261), .QN(n10259) );
  NAND2X0 U10206 ( .IN1(n10261), .IN2(n10260), .QN(n10257) );
  NOR2X0 U10207 ( .IN1(n10262), .IN2(n10263), .QN(n10260) );
  NOR2X0 U10208 ( .IN1(WX9928), .IN2(n7905), .QN(n10263) );
  INVX0 U10209 ( .INP(n10264), .ZN(n10262) );
  NAND2X0 U10210 ( .IN1(n7905), .IN2(WX9928), .QN(n10264) );
  NAND2X0 U10211 ( .IN1(n10265), .IN2(n10266), .QN(n10261) );
  NAND2X0 U10212 ( .IN1(n7904), .IN2(WX9800), .QN(n10266) );
  INVX0 U10213 ( .INP(n10267), .ZN(n10265) );
  NOR2X0 U10214 ( .IN1(WX9800), .IN2(n7904), .QN(n10267) );
  NAND2X0 U10215 ( .IN1(n1474), .IN2(n9274), .QN(n10252) );
  NOR2X0 U10216 ( .IN1(n9229), .IN2(n8867), .QN(n1474) );
  NAND2X0 U10217 ( .IN1(n9305), .IN2(CRC_OUT_3_11), .QN(n10251) );
  NAND4X0 U10218 ( .IN1(n10268), .IN2(n10269), .IN3(n10270), .IN4(n10271), 
        .QN(WX8440) );
  NAND2X0 U10219 ( .IN1(n9329), .IN2(n9759), .QN(n10271) );
  NAND2X0 U10220 ( .IN1(n10272), .IN2(n10273), .QN(n9759) );
  INVX0 U10221 ( .INP(n10274), .ZN(n10273) );
  NOR2X0 U10222 ( .IN1(n10275), .IN2(n10276), .QN(n10274) );
  NAND2X0 U10223 ( .IN1(n10276), .IN2(n10275), .QN(n10272) );
  NOR2X0 U10224 ( .IN1(n10277), .IN2(n10278), .QN(n10275) );
  NOR2X0 U10225 ( .IN1(WX9926), .IN2(n7907), .QN(n10278) );
  INVX0 U10226 ( .INP(n10279), .ZN(n10277) );
  NAND2X0 U10227 ( .IN1(n7907), .IN2(WX9926), .QN(n10279) );
  NAND2X0 U10228 ( .IN1(n10280), .IN2(n10281), .QN(n10276) );
  NAND2X0 U10229 ( .IN1(n7906), .IN2(WX9798), .QN(n10281) );
  INVX0 U10230 ( .INP(n10282), .ZN(n10280) );
  NOR2X0 U10231 ( .IN1(WX9798), .IN2(n7906), .QN(n10282) );
  NAND2X0 U10232 ( .IN1(n9097), .IN2(n10283), .QN(n10270) );
  NAND2X0 U10233 ( .IN1(n1473), .IN2(n9274), .QN(n10269) );
  NOR2X0 U10234 ( .IN1(n9229), .IN2(n8868), .QN(n1473) );
  NAND2X0 U10235 ( .IN1(n9305), .IN2(CRC_OUT_3_12), .QN(n10268) );
  NAND4X0 U10236 ( .IN1(n10284), .IN2(n10285), .IN3(n10286), .IN4(n10287), 
        .QN(WX8438) );
  NAND3X0 U10237 ( .IN1(n10288), .IN2(n10289), .IN3(n9091), .QN(n10287) );
  NAND2X0 U10238 ( .IN1(n9329), .IN2(n9765), .QN(n10286) );
  NAND2X0 U10239 ( .IN1(n10290), .IN2(n10291), .QN(n9765) );
  INVX0 U10240 ( .INP(n10292), .ZN(n10291) );
  NOR2X0 U10241 ( .IN1(n10293), .IN2(n10294), .QN(n10292) );
  NAND2X0 U10242 ( .IN1(n10294), .IN2(n10293), .QN(n10290) );
  NOR2X0 U10243 ( .IN1(n10295), .IN2(n10296), .QN(n10293) );
  NOR2X0 U10244 ( .IN1(WX9924), .IN2(n7909), .QN(n10296) );
  INVX0 U10245 ( .INP(n10297), .ZN(n10295) );
  NAND2X0 U10246 ( .IN1(n7909), .IN2(WX9924), .QN(n10297) );
  NAND2X0 U10247 ( .IN1(n10298), .IN2(n10299), .QN(n10294) );
  NAND2X0 U10248 ( .IN1(n7908), .IN2(WX9796), .QN(n10299) );
  INVX0 U10249 ( .INP(n10300), .ZN(n10298) );
  NOR2X0 U10250 ( .IN1(WX9796), .IN2(n7908), .QN(n10300) );
  NAND2X0 U10251 ( .IN1(n1472), .IN2(n9274), .QN(n10285) );
  NOR2X0 U10252 ( .IN1(n9230), .IN2(n8869), .QN(n1472) );
  NAND2X0 U10253 ( .IN1(n9306), .IN2(CRC_OUT_3_13), .QN(n10284) );
  NAND4X0 U10254 ( .IN1(n10301), .IN2(n10302), .IN3(n10303), .IN4(n10304), 
        .QN(WX8436) );
  NAND3X0 U10255 ( .IN1(n9771), .IN2(n9772), .IN3(n9321), .QN(n10304) );
  NAND3X0 U10256 ( .IN1(n10305), .IN2(n10306), .IN3(n10307), .QN(n9772) );
  INVX0 U10257 ( .INP(n10308), .ZN(n10307) );
  NAND2X0 U10258 ( .IN1(n10308), .IN2(n10309), .QN(n9771) );
  NAND2X0 U10259 ( .IN1(n10305), .IN2(n10306), .QN(n10309) );
  NAND2X0 U10260 ( .IN1(n7911), .IN2(WX9794), .QN(n10306) );
  NAND2X0 U10261 ( .IN1(n3591), .IN2(WX9858), .QN(n10305) );
  NOR2X0 U10262 ( .IN1(n10310), .IN2(n10311), .QN(n10308) );
  NOR2X0 U10263 ( .IN1(n8794), .IN2(n7910), .QN(n10311) );
  INVX0 U10264 ( .INP(n10312), .ZN(n10310) );
  NAND2X0 U10265 ( .IN1(n7910), .IN2(n8794), .QN(n10312) );
  NAND2X0 U10266 ( .IN1(n9097), .IN2(n10313), .QN(n10303) );
  NAND2X0 U10267 ( .IN1(n1471), .IN2(n9274), .QN(n10302) );
  NOR2X0 U10268 ( .IN1(n9230), .IN2(n8870), .QN(n1471) );
  NAND2X0 U10269 ( .IN1(n9306), .IN2(CRC_OUT_3_14), .QN(n10301) );
  NAND4X0 U10270 ( .IN1(n10314), .IN2(n10315), .IN3(n10316), .IN4(n10317), 
        .QN(WX8434) );
  NAND3X0 U10271 ( .IN1(n10318), .IN2(n10319), .IN3(n9091), .QN(n10317) );
  NAND2X0 U10272 ( .IN1(n9330), .IN2(n9778), .QN(n10316) );
  NAND2X0 U10273 ( .IN1(n10320), .IN2(n10321), .QN(n9778) );
  INVX0 U10274 ( .INP(n10322), .ZN(n10321) );
  NOR2X0 U10275 ( .IN1(n10323), .IN2(n10324), .QN(n10322) );
  NAND2X0 U10276 ( .IN1(n10324), .IN2(n10323), .QN(n10320) );
  NOR2X0 U10277 ( .IN1(n10325), .IN2(n10326), .QN(n10323) );
  NOR2X0 U10278 ( .IN1(WX9920), .IN2(n7913), .QN(n10326) );
  INVX0 U10279 ( .INP(n10327), .ZN(n10325) );
  NAND2X0 U10280 ( .IN1(n7913), .IN2(WX9920), .QN(n10327) );
  NAND2X0 U10281 ( .IN1(n10328), .IN2(n10329), .QN(n10324) );
  NAND2X0 U10282 ( .IN1(n7912), .IN2(WX9792), .QN(n10329) );
  INVX0 U10283 ( .INP(n10330), .ZN(n10328) );
  NOR2X0 U10284 ( .IN1(WX9792), .IN2(n7912), .QN(n10330) );
  NAND2X0 U10285 ( .IN1(n1470), .IN2(n9274), .QN(n10315) );
  NOR2X0 U10286 ( .IN1(n9230), .IN2(n8871), .QN(n1470) );
  NAND2X0 U10287 ( .IN1(n9306), .IN2(CRC_OUT_3_15), .QN(n10314) );
  NAND4X0 U10288 ( .IN1(n10331), .IN2(n10332), .IN3(n10333), .IN4(n10334), 
        .QN(WX8432) );
  NAND2X0 U10289 ( .IN1(n10335), .IN2(n10336), .QN(n10334) );
  NAND2X0 U10290 ( .IN1(n10337), .IN2(n10338), .QN(n10335) );
  NAND2X0 U10291 ( .IN1(n9097), .IN2(n10339), .QN(n10338) );
  NAND2X0 U10292 ( .IN1(n9097), .IN2(n8363), .QN(n10337) );
  NAND2X0 U10293 ( .IN1(n9792), .IN2(n2153), .QN(n10333) );
  NOR2X0 U10294 ( .IN1(n10340), .IN2(n10341), .QN(n9792) );
  INVX0 U10295 ( .INP(n10342), .ZN(n10341) );
  NAND2X0 U10296 ( .IN1(n10343), .IN2(n10344), .QN(n10342) );
  NOR2X0 U10297 ( .IN1(n10344), .IN2(n10343), .QN(n10340) );
  NAND2X0 U10298 ( .IN1(n10345), .IN2(n10346), .QN(n10343) );
  NAND2X0 U10299 ( .IN1(n8107), .IN2(n10347), .QN(n10346) );
  INVX0 U10300 ( .INP(n10348), .ZN(n10347) );
  NAND2X0 U10301 ( .IN1(n10348), .IN2(WX9918), .QN(n10345) );
  NAND2X0 U10302 ( .IN1(n10349), .IN2(n10350), .QN(n10348) );
  INVX0 U10303 ( .INP(n10351), .ZN(n10350) );
  NOR2X0 U10304 ( .IN1(n8805), .IN2(n16132), .QN(n10351) );
  NAND2X0 U10305 ( .IN1(n16132), .IN2(n8805), .QN(n10349) );
  NOR2X0 U10306 ( .IN1(n10352), .IN2(n10353), .QN(n10344) );
  INVX0 U10307 ( .INP(n10354), .ZN(n10353) );
  NAND2X0 U10308 ( .IN1(n7655), .IN2(n9120), .QN(n10354) );
  NOR2X0 U10309 ( .IN1(n9115), .IN2(n7655), .QN(n10352) );
  NAND2X0 U10310 ( .IN1(n1469), .IN2(n9274), .QN(n10332) );
  NOR2X0 U10311 ( .IN1(n9230), .IN2(n8872), .QN(n1469) );
  NAND2X0 U10312 ( .IN1(n9306), .IN2(CRC_OUT_3_16), .QN(n10331) );
  NAND4X0 U10313 ( .IN1(n10356), .IN2(n10357), .IN3(n10358), .IN4(n10359), 
        .QN(WX8430) );
  NAND2X0 U10314 ( .IN1(n10360), .IN2(n9798), .QN(n10359) );
  NAND2X0 U10315 ( .IN1(n10361), .IN2(n9801), .QN(n9798) );
  NAND2X0 U10316 ( .IN1(n10362), .IN2(n10363), .QN(n10361) );
  NAND2X0 U10317 ( .IN1(n16131), .IN2(n9120), .QN(n10363) );
  NAND2X0 U10318 ( .IN1(TM1), .IN2(n8305), .QN(n10362) );
  NAND3X0 U10319 ( .IN1(n10364), .IN2(n10365), .IN3(n10366), .QN(n10360) );
  NAND2X0 U10320 ( .IN1(n9330), .IN2(n9801), .QN(n10366) );
  NAND2X0 U10321 ( .IN1(n10367), .IN2(n10368), .QN(n9801) );
  NAND2X0 U10322 ( .IN1(n7656), .IN2(n10369), .QN(n10368) );
  INVX0 U10323 ( .INP(n10370), .ZN(n10367) );
  NOR2X0 U10324 ( .IN1(n10369), .IN2(n7656), .QN(n10370) );
  NOR2X0 U10325 ( .IN1(n10371), .IN2(n10372), .QN(n10369) );
  NOR2X0 U10326 ( .IN1(WX9916), .IN2(n7657), .QN(n10372) );
  INVX0 U10327 ( .INP(n10373), .ZN(n10371) );
  NAND2X0 U10328 ( .IN1(n7657), .IN2(WX9916), .QN(n10373) );
  NAND2X0 U10329 ( .IN1(n9082), .IN2(n8305), .QN(n10365) );
  NAND2X0 U10330 ( .IN1(n16131), .IN2(n9791), .QN(n10364) );
  NAND2X0 U10331 ( .IN1(n10374), .IN2(n10375), .QN(n10358) );
  NAND2X0 U10332 ( .IN1(n10376), .IN2(n10377), .QN(n10374) );
  NAND2X0 U10333 ( .IN1(n9097), .IN2(n10378), .QN(n10377) );
  NAND2X0 U10334 ( .IN1(n9097), .IN2(n8364), .QN(n10376) );
  NAND2X0 U10335 ( .IN1(n1468), .IN2(n9274), .QN(n10357) );
  NOR2X0 U10336 ( .IN1(n9063), .IN2(n9156), .QN(n1468) );
  NAND2X0 U10337 ( .IN1(n9306), .IN2(CRC_OUT_3_17), .QN(n10356) );
  NAND4X0 U10338 ( .IN1(n10379), .IN2(n10380), .IN3(n10381), .IN4(n10382), 
        .QN(WX8428) );
  NAND2X0 U10339 ( .IN1(n10383), .IN2(n10384), .QN(n10382) );
  NAND2X0 U10340 ( .IN1(n10385), .IN2(n10386), .QN(n10383) );
  NAND2X0 U10341 ( .IN1(n9097), .IN2(n10387), .QN(n10386) );
  NAND2X0 U10342 ( .IN1(n9097), .IN2(n8365), .QN(n10385) );
  NAND2X0 U10343 ( .IN1(n9818), .IN2(n2153), .QN(n10381) );
  NOR2X0 U10344 ( .IN1(n10388), .IN2(n10389), .QN(n9818) );
  INVX0 U10345 ( .INP(n10390), .ZN(n10389) );
  NAND2X0 U10346 ( .IN1(n10391), .IN2(n10392), .QN(n10390) );
  NOR2X0 U10347 ( .IN1(n10392), .IN2(n10391), .QN(n10388) );
  NAND2X0 U10348 ( .IN1(n10393), .IN2(n10394), .QN(n10391) );
  NAND2X0 U10349 ( .IN1(n8171), .IN2(n10395), .QN(n10394) );
  INVX0 U10350 ( .INP(n10396), .ZN(n10395) );
  NAND2X0 U10351 ( .IN1(n10396), .IN2(WX9914), .QN(n10393) );
  NAND2X0 U10352 ( .IN1(n10397), .IN2(n10398), .QN(n10396) );
  INVX0 U10353 ( .INP(n10399), .ZN(n10398) );
  NOR2X0 U10354 ( .IN1(n8806), .IN2(n16130), .QN(n10399) );
  NAND2X0 U10355 ( .IN1(n16130), .IN2(n8806), .QN(n10397) );
  NOR2X0 U10356 ( .IN1(n10400), .IN2(n10401), .QN(n10392) );
  INVX0 U10357 ( .INP(n10402), .ZN(n10401) );
  NAND2X0 U10358 ( .IN1(n7658), .IN2(n9120), .QN(n10402) );
  NOR2X0 U10359 ( .IN1(n9115), .IN2(n7658), .QN(n10400) );
  NAND2X0 U10360 ( .IN1(n1467), .IN2(n9274), .QN(n10380) );
  NOR2X0 U10361 ( .IN1(n9230), .IN2(n8873), .QN(n1467) );
  NAND2X0 U10362 ( .IN1(n9306), .IN2(CRC_OUT_3_18), .QN(n10379) );
  NAND4X0 U10363 ( .IN1(n10403), .IN2(n10404), .IN3(n10405), .IN4(n10406), 
        .QN(WX8426) );
  NAND2X0 U10364 ( .IN1(n10407), .IN2(n9824), .QN(n10406) );
  NAND2X0 U10365 ( .IN1(n10408), .IN2(n9827), .QN(n9824) );
  NAND2X0 U10366 ( .IN1(n10409), .IN2(n10410), .QN(n10408) );
  NAND2X0 U10367 ( .IN1(n16129), .IN2(n9120), .QN(n10410) );
  NAND2X0 U10368 ( .IN1(TM1), .IN2(n8307), .QN(n10409) );
  NAND3X0 U10369 ( .IN1(n10411), .IN2(n10412), .IN3(n10413), .QN(n10407) );
  NAND2X0 U10370 ( .IN1(n9330), .IN2(n9827), .QN(n10413) );
  NAND2X0 U10371 ( .IN1(n10414), .IN2(n10415), .QN(n9827) );
  NAND2X0 U10372 ( .IN1(n7659), .IN2(n10416), .QN(n10415) );
  INVX0 U10373 ( .INP(n10417), .ZN(n10414) );
  NOR2X0 U10374 ( .IN1(n10416), .IN2(n7659), .QN(n10417) );
  NOR2X0 U10375 ( .IN1(n10418), .IN2(n10419), .QN(n10416) );
  NOR2X0 U10376 ( .IN1(WX9912), .IN2(n7660), .QN(n10419) );
  INVX0 U10377 ( .INP(n10420), .ZN(n10418) );
  NAND2X0 U10378 ( .IN1(n7660), .IN2(WX9912), .QN(n10420) );
  NAND2X0 U10379 ( .IN1(n9081), .IN2(n8307), .QN(n10412) );
  NAND2X0 U10380 ( .IN1(n16129), .IN2(n9079), .QN(n10411) );
  NAND2X0 U10381 ( .IN1(n10421), .IN2(n10422), .QN(n10405) );
  NAND2X0 U10382 ( .IN1(n10423), .IN2(n10424), .QN(n10421) );
  NAND2X0 U10383 ( .IN1(n9097), .IN2(n10425), .QN(n10424) );
  NAND2X0 U10384 ( .IN1(n9097), .IN2(n8366), .QN(n10423) );
  NAND2X0 U10385 ( .IN1(n1466), .IN2(n9275), .QN(n10404) );
  NOR2X0 U10386 ( .IN1(n9230), .IN2(n8874), .QN(n1466) );
  NAND2X0 U10387 ( .IN1(n9306), .IN2(CRC_OUT_3_19), .QN(n10403) );
  NAND4X0 U10388 ( .IN1(n10426), .IN2(n10427), .IN3(n10428), .IN4(n10429), 
        .QN(WX8424) );
  NAND2X0 U10389 ( .IN1(n10430), .IN2(n9834), .QN(n10429) );
  NAND3X0 U10390 ( .IN1(n10431), .IN2(n10432), .IN3(n9837), .QN(n9834) );
  NAND2X0 U10391 ( .IN1(n8169), .IN2(n9120), .QN(n10432) );
  NAND2X0 U10392 ( .IN1(TM1), .IN2(WX9910), .QN(n10431) );
  NAND3X0 U10393 ( .IN1(n10433), .IN2(n10434), .IN3(n10435), .QN(n10430) );
  NAND2X0 U10394 ( .IN1(n9330), .IN2(n9837), .QN(n10435) );
  NAND2X0 U10395 ( .IN1(n10436), .IN2(n10437), .QN(n9837) );
  NAND2X0 U10396 ( .IN1(n10438), .IN2(WX9846), .QN(n10437) );
  NAND2X0 U10397 ( .IN1(n10439), .IN2(n10440), .QN(n10438) );
  NAND3X0 U10398 ( .IN1(n10439), .IN2(n10440), .IN3(n7662), .QN(n10436) );
  NAND2X0 U10399 ( .IN1(test_so80), .IN2(WX9782), .QN(n10440) );
  NAND2X0 U10400 ( .IN1(n7661), .IN2(n8819), .QN(n10439) );
  NAND2X0 U10401 ( .IN1(n9079), .IN2(WX9910), .QN(n10434) );
  NAND2X0 U10402 ( .IN1(n9790), .IN2(n8169), .QN(n10433) );
  NAND2X0 U10403 ( .IN1(n10441), .IN2(n10442), .QN(n10428) );
  NAND2X0 U10404 ( .IN1(n10443), .IN2(n10444), .QN(n10441) );
  NAND2X0 U10405 ( .IN1(n9097), .IN2(n10445), .QN(n10444) );
  NAND2X0 U10406 ( .IN1(n9097), .IN2(n8367), .QN(n10443) );
  NAND2X0 U10407 ( .IN1(n1465), .IN2(n9275), .QN(n10427) );
  NOR2X0 U10408 ( .IN1(n9230), .IN2(n8875), .QN(n1465) );
  NAND2X0 U10409 ( .IN1(n9306), .IN2(CRC_OUT_3_20), .QN(n10426) );
  NAND4X0 U10410 ( .IN1(n10446), .IN2(n10447), .IN3(n10448), .IN4(n10449), 
        .QN(WX8422) );
  NAND2X0 U10411 ( .IN1(n10450), .IN2(n9849), .QN(n10449) );
  NAND2X0 U10412 ( .IN1(n10451), .IN2(n9852), .QN(n9849) );
  NAND2X0 U10413 ( .IN1(n10452), .IN2(n10453), .QN(n10451) );
  NAND2X0 U10414 ( .IN1(n16128), .IN2(n9120), .QN(n10453) );
  NAND2X0 U10415 ( .IN1(TM1), .IN2(n8310), .QN(n10452) );
  NAND3X0 U10416 ( .IN1(n10454), .IN2(n10455), .IN3(n10456), .QN(n10450) );
  NAND2X0 U10417 ( .IN1(n9330), .IN2(n9852), .QN(n10456) );
  NAND2X0 U10418 ( .IN1(n10457), .IN2(n10458), .QN(n9852) );
  NAND2X0 U10419 ( .IN1(n7663), .IN2(n10459), .QN(n10458) );
  INVX0 U10420 ( .INP(n10460), .ZN(n10457) );
  NOR2X0 U10421 ( .IN1(n10459), .IN2(n7663), .QN(n10460) );
  NOR2X0 U10422 ( .IN1(n10461), .IN2(n10462), .QN(n10459) );
  NOR2X0 U10423 ( .IN1(WX9908), .IN2(n7664), .QN(n10462) );
  INVX0 U10424 ( .INP(n10463), .ZN(n10461) );
  NAND2X0 U10425 ( .IN1(n7664), .IN2(WX9908), .QN(n10463) );
  NAND2X0 U10426 ( .IN1(n9083), .IN2(n8310), .QN(n10455) );
  NAND2X0 U10427 ( .IN1(n16128), .IN2(n9078), .QN(n10454) );
  NAND2X0 U10428 ( .IN1(n10464), .IN2(n10465), .QN(n10448) );
  NAND2X0 U10429 ( .IN1(n10466), .IN2(n10467), .QN(n10464) );
  NAND2X0 U10430 ( .IN1(n9097), .IN2(n10468), .QN(n10467) );
  NAND2X0 U10431 ( .IN1(n9097), .IN2(n8368), .QN(n10466) );
  NAND2X0 U10432 ( .IN1(n1464), .IN2(n9275), .QN(n10447) );
  NOR2X0 U10433 ( .IN1(n9230), .IN2(n8876), .QN(n1464) );
  NAND2X0 U10434 ( .IN1(n9306), .IN2(CRC_OUT_3_21), .QN(n10446) );
  NAND4X0 U10435 ( .IN1(n10469), .IN2(n10470), .IN3(n10471), .IN4(n10472), 
        .QN(WX8420) );
  NAND2X0 U10436 ( .IN1(n10473), .IN2(n9859), .QN(n10472) );
  NAND2X0 U10437 ( .IN1(n10474), .IN2(n9862), .QN(n9859) );
  NAND2X0 U10438 ( .IN1(n10475), .IN2(n10476), .QN(n10474) );
  NAND2X0 U10439 ( .IN1(n16127), .IN2(n9120), .QN(n10476) );
  NAND2X0 U10440 ( .IN1(TM1), .IN2(n8311), .QN(n10475) );
  NAND3X0 U10441 ( .IN1(n10477), .IN2(n10478), .IN3(n10479), .QN(n10473) );
  NAND2X0 U10442 ( .IN1(n9330), .IN2(n9862), .QN(n10479) );
  NAND2X0 U10443 ( .IN1(n10480), .IN2(n10481), .QN(n9862) );
  NAND2X0 U10444 ( .IN1(n7665), .IN2(n10482), .QN(n10481) );
  INVX0 U10445 ( .INP(n10483), .ZN(n10480) );
  NOR2X0 U10446 ( .IN1(n10482), .IN2(n7665), .QN(n10483) );
  NOR2X0 U10447 ( .IN1(n10484), .IN2(n10485), .QN(n10482) );
  NOR2X0 U10448 ( .IN1(WX9906), .IN2(n7666), .QN(n10485) );
  INVX0 U10449 ( .INP(n10486), .ZN(n10484) );
  NAND2X0 U10450 ( .IN1(n7666), .IN2(WX9906), .QN(n10486) );
  NAND2X0 U10451 ( .IN1(n9082), .IN2(n8311), .QN(n10478) );
  NAND2X0 U10452 ( .IN1(n16127), .IN2(n9077), .QN(n10477) );
  NAND2X0 U10453 ( .IN1(n10487), .IN2(n10488), .QN(n10471) );
  NAND2X0 U10454 ( .IN1(n10489), .IN2(n10490), .QN(n10487) );
  NAND2X0 U10455 ( .IN1(n9097), .IN2(n10491), .QN(n10490) );
  NAND2X0 U10456 ( .IN1(n9097), .IN2(n8369), .QN(n10489) );
  NAND2X0 U10457 ( .IN1(n1463), .IN2(n9275), .QN(n10470) );
  NOR2X0 U10458 ( .IN1(n9230), .IN2(n8877), .QN(n1463) );
  NAND2X0 U10459 ( .IN1(n9306), .IN2(CRC_OUT_3_22), .QN(n10469) );
  NAND4X0 U10460 ( .IN1(n10492), .IN2(n10493), .IN3(n10494), .IN4(n10495), 
        .QN(WX8418) );
  NAND2X0 U10461 ( .IN1(n10496), .IN2(n9874), .QN(n10495) );
  NAND2X0 U10462 ( .IN1(n10497), .IN2(n9877), .QN(n9874) );
  NAND2X0 U10463 ( .IN1(n10498), .IN2(n10499), .QN(n10497) );
  NAND2X0 U10464 ( .IN1(n16126), .IN2(n9119), .QN(n10499) );
  NAND2X0 U10465 ( .IN1(TM1), .IN2(n8312), .QN(n10498) );
  NAND3X0 U10466 ( .IN1(n10500), .IN2(n10501), .IN3(n10502), .QN(n10496) );
  NAND2X0 U10467 ( .IN1(n9330), .IN2(n9877), .QN(n10502) );
  NAND2X0 U10468 ( .IN1(n10503), .IN2(n10504), .QN(n9877) );
  NAND2X0 U10469 ( .IN1(n7667), .IN2(n10505), .QN(n10504) );
  INVX0 U10470 ( .INP(n10506), .ZN(n10503) );
  NOR2X0 U10471 ( .IN1(n10505), .IN2(n7667), .QN(n10506) );
  NOR2X0 U10472 ( .IN1(n10507), .IN2(n10508), .QN(n10505) );
  NOR2X0 U10473 ( .IN1(WX9904), .IN2(n7668), .QN(n10508) );
  INVX0 U10474 ( .INP(n10509), .ZN(n10507) );
  NAND2X0 U10475 ( .IN1(n7668), .IN2(WX9904), .QN(n10509) );
  NAND2X0 U10476 ( .IN1(n9081), .IN2(n8312), .QN(n10501) );
  NAND2X0 U10477 ( .IN1(n16126), .IN2(n9791), .QN(n10500) );
  NAND2X0 U10478 ( .IN1(n10510), .IN2(n10511), .QN(n10494) );
  NAND2X0 U10479 ( .IN1(n10512), .IN2(n10513), .QN(n10510) );
  NAND2X0 U10480 ( .IN1(n9096), .IN2(n10514), .QN(n10513) );
  NAND2X0 U10481 ( .IN1(n9096), .IN2(n8370), .QN(n10512) );
  NAND2X0 U10482 ( .IN1(n1462), .IN2(n9275), .QN(n10493) );
  NOR2X0 U10483 ( .IN1(n9230), .IN2(n8878), .QN(n1462) );
  NAND2X0 U10484 ( .IN1(n9306), .IN2(CRC_OUT_3_23), .QN(n10492) );
  NAND4X0 U10485 ( .IN1(n10515), .IN2(n10516), .IN3(n10517), .IN4(n10518), 
        .QN(WX8416) );
  NAND2X0 U10486 ( .IN1(n10519), .IN2(n9884), .QN(n10518) );
  NAND2X0 U10487 ( .IN1(n10520), .IN2(n9887), .QN(n9884) );
  NAND2X0 U10488 ( .IN1(n10521), .IN2(n10522), .QN(n10520) );
  NAND2X0 U10489 ( .IN1(n16125), .IN2(n9119), .QN(n10522) );
  NAND2X0 U10490 ( .IN1(TM1), .IN2(n8313), .QN(n10521) );
  NAND3X0 U10491 ( .IN1(n10523), .IN2(n10524), .IN3(n10525), .QN(n10519) );
  NAND2X0 U10492 ( .IN1(n9330), .IN2(n9887), .QN(n10525) );
  NAND2X0 U10493 ( .IN1(n10526), .IN2(n10527), .QN(n9887) );
  NAND2X0 U10494 ( .IN1(n7669), .IN2(n10528), .QN(n10527) );
  INVX0 U10495 ( .INP(n10529), .ZN(n10526) );
  NOR2X0 U10496 ( .IN1(n10528), .IN2(n7669), .QN(n10529) );
  NOR2X0 U10497 ( .IN1(n10530), .IN2(n10531), .QN(n10528) );
  NOR2X0 U10498 ( .IN1(WX9902), .IN2(n7670), .QN(n10531) );
  INVX0 U10499 ( .INP(n10532), .ZN(n10530) );
  NAND2X0 U10500 ( .IN1(n7670), .IN2(WX9902), .QN(n10532) );
  NAND2X0 U10501 ( .IN1(n9790), .IN2(n8313), .QN(n10524) );
  NAND2X0 U10502 ( .IN1(n16125), .IN2(n9079), .QN(n10523) );
  NAND2X0 U10503 ( .IN1(n10533), .IN2(n10534), .QN(n10517) );
  NAND2X0 U10504 ( .IN1(n10535), .IN2(n10536), .QN(n10533) );
  NAND2X0 U10505 ( .IN1(n9096), .IN2(n10537), .QN(n10536) );
  NAND2X0 U10506 ( .IN1(n9096), .IN2(n8371), .QN(n10535) );
  NAND2X0 U10507 ( .IN1(n1461), .IN2(n9275), .QN(n10516) );
  NOR2X0 U10508 ( .IN1(n9231), .IN2(n8879), .QN(n1461) );
  NAND2X0 U10509 ( .IN1(test_so77), .IN2(n9313), .QN(n10515) );
  NAND4X0 U10510 ( .IN1(n10538), .IN2(n10539), .IN3(n10540), .IN4(n10541), 
        .QN(WX8414) );
  NAND2X0 U10511 ( .IN1(n10542), .IN2(n9899), .QN(n10541) );
  NAND2X0 U10512 ( .IN1(n10543), .IN2(n9902), .QN(n9899) );
  NAND2X0 U10513 ( .IN1(n10544), .IN2(n10545), .QN(n10543) );
  NAND2X0 U10514 ( .IN1(n16124), .IN2(n9119), .QN(n10545) );
  NAND2X0 U10515 ( .IN1(TM1), .IN2(n8314), .QN(n10544) );
  NAND3X0 U10516 ( .IN1(n10546), .IN2(n10547), .IN3(n10548), .QN(n10542) );
  NAND2X0 U10517 ( .IN1(n9330), .IN2(n9902), .QN(n10548) );
  NAND2X0 U10518 ( .IN1(n10549), .IN2(n10550), .QN(n9902) );
  NAND2X0 U10519 ( .IN1(n7671), .IN2(n10551), .QN(n10550) );
  INVX0 U10520 ( .INP(n10552), .ZN(n10549) );
  NOR2X0 U10521 ( .IN1(n10551), .IN2(n7671), .QN(n10552) );
  NOR2X0 U10522 ( .IN1(n10553), .IN2(n10554), .QN(n10551) );
  NOR2X0 U10523 ( .IN1(WX9900), .IN2(n7672), .QN(n10554) );
  INVX0 U10524 ( .INP(n10555), .ZN(n10553) );
  NAND2X0 U10525 ( .IN1(n7672), .IN2(WX9900), .QN(n10555) );
  NAND2X0 U10526 ( .IN1(n9083), .IN2(n8314), .QN(n10547) );
  NAND2X0 U10527 ( .IN1(n16124), .IN2(n9078), .QN(n10546) );
  NAND2X0 U10528 ( .IN1(n10556), .IN2(n10557), .QN(n10540) );
  NAND2X0 U10529 ( .IN1(n10558), .IN2(n10559), .QN(n10556) );
  NAND2X0 U10530 ( .IN1(n9096), .IN2(n10560), .QN(n10559) );
  NAND2X0 U10531 ( .IN1(n9096), .IN2(n8372), .QN(n10558) );
  NAND2X0 U10532 ( .IN1(n1460), .IN2(n9275), .QN(n10539) );
  NOR2X0 U10533 ( .IN1(n9231), .IN2(n8880), .QN(n1460) );
  NAND2X0 U10534 ( .IN1(n9306), .IN2(CRC_OUT_3_25), .QN(n10538) );
  NAND4X0 U10535 ( .IN1(n10561), .IN2(n10562), .IN3(n10563), .IN4(n10564), 
        .QN(WX8412) );
  NAND2X0 U10536 ( .IN1(n10565), .IN2(n9914), .QN(n10564) );
  NAND2X0 U10537 ( .IN1(n10566), .IN2(n9917), .QN(n9914) );
  NAND2X0 U10538 ( .IN1(n10567), .IN2(n10568), .QN(n10566) );
  NAND2X0 U10539 ( .IN1(n16123), .IN2(n9119), .QN(n10568) );
  NAND2X0 U10540 ( .IN1(TM1), .IN2(n8315), .QN(n10567) );
  NAND3X0 U10541 ( .IN1(n10569), .IN2(n10570), .IN3(n10571), .QN(n10565) );
  NAND2X0 U10542 ( .IN1(n9330), .IN2(n9917), .QN(n10571) );
  NAND2X0 U10543 ( .IN1(n10572), .IN2(n10573), .QN(n9917) );
  NAND2X0 U10544 ( .IN1(n7673), .IN2(n10574), .QN(n10573) );
  INVX0 U10545 ( .INP(n10575), .ZN(n10572) );
  NOR2X0 U10546 ( .IN1(n10574), .IN2(n7673), .QN(n10575) );
  NOR2X0 U10547 ( .IN1(n10576), .IN2(n10577), .QN(n10574) );
  NOR2X0 U10548 ( .IN1(WX9898), .IN2(n7674), .QN(n10577) );
  INVX0 U10549 ( .INP(n10578), .ZN(n10576) );
  NAND2X0 U10550 ( .IN1(n7674), .IN2(WX9898), .QN(n10578) );
  NAND2X0 U10551 ( .IN1(n9082), .IN2(n8315), .QN(n10570) );
  NAND2X0 U10552 ( .IN1(n16123), .IN2(n9077), .QN(n10569) );
  NAND2X0 U10553 ( .IN1(n10579), .IN2(n9109), .QN(n10563) );
  NAND2X0 U10554 ( .IN1(n1459), .IN2(n9275), .QN(n10562) );
  NOR2X0 U10555 ( .IN1(n9231), .IN2(n8881), .QN(n1459) );
  NAND2X0 U10556 ( .IN1(n9307), .IN2(CRC_OUT_3_26), .QN(n10561) );
  NAND4X0 U10557 ( .IN1(n10580), .IN2(n10581), .IN3(n10582), .IN4(n10583), 
        .QN(WX8410) );
  NAND2X0 U10558 ( .IN1(n10584), .IN2(n9929), .QN(n10583) );
  NAND2X0 U10559 ( .IN1(n10585), .IN2(n9932), .QN(n9929) );
  NAND2X0 U10560 ( .IN1(n10586), .IN2(n10587), .QN(n10585) );
  NAND2X0 U10561 ( .IN1(n16122), .IN2(n9119), .QN(n10587) );
  NAND2X0 U10562 ( .IN1(TM1), .IN2(n8316), .QN(n10586) );
  NAND3X0 U10563 ( .IN1(n10588), .IN2(n10589), .IN3(n10590), .QN(n10584) );
  NAND2X0 U10564 ( .IN1(n9330), .IN2(n9932), .QN(n10590) );
  NAND2X0 U10565 ( .IN1(n10591), .IN2(n10592), .QN(n9932) );
  NAND2X0 U10566 ( .IN1(n7675), .IN2(n10593), .QN(n10592) );
  INVX0 U10567 ( .INP(n10594), .ZN(n10591) );
  NOR2X0 U10568 ( .IN1(n10593), .IN2(n7675), .QN(n10594) );
  NOR2X0 U10569 ( .IN1(n10595), .IN2(n10596), .QN(n10593) );
  NOR2X0 U10570 ( .IN1(WX9896), .IN2(n7676), .QN(n10596) );
  INVX0 U10571 ( .INP(n10597), .ZN(n10595) );
  NAND2X0 U10572 ( .IN1(n7676), .IN2(WX9896), .QN(n10597) );
  NAND2X0 U10573 ( .IN1(n9081), .IN2(n8316), .QN(n10589) );
  NAND2X0 U10574 ( .IN1(n16122), .IN2(n9791), .QN(n10588) );
  NAND2X0 U10575 ( .IN1(n10598), .IN2(n10599), .QN(n10582) );
  NAND2X0 U10576 ( .IN1(n10600), .IN2(n10601), .QN(n10598) );
  NAND2X0 U10577 ( .IN1(n9096), .IN2(n10602), .QN(n10601) );
  NAND2X0 U10578 ( .IN1(n9096), .IN2(n8374), .QN(n10600) );
  NAND2X0 U10579 ( .IN1(n1458), .IN2(n9275), .QN(n10581) );
  NOR2X0 U10580 ( .IN1(n9231), .IN2(n8882), .QN(n1458) );
  NAND2X0 U10581 ( .IN1(n9307), .IN2(CRC_OUT_3_27), .QN(n10580) );
  NAND4X0 U10582 ( .IN1(n10603), .IN2(n10604), .IN3(n10605), .IN4(n10606), 
        .QN(WX8408) );
  NAND2X0 U10583 ( .IN1(n10607), .IN2(n9944), .QN(n10606) );
  NAND2X0 U10584 ( .IN1(n10608), .IN2(n9947), .QN(n9944) );
  NAND2X0 U10585 ( .IN1(n10609), .IN2(n10610), .QN(n10608) );
  NAND2X0 U10586 ( .IN1(n16121), .IN2(n9119), .QN(n10610) );
  NAND2X0 U10587 ( .IN1(TM1), .IN2(n8317), .QN(n10609) );
  NAND3X0 U10588 ( .IN1(n10611), .IN2(n10612), .IN3(n10613), .QN(n10607) );
  NAND2X0 U10589 ( .IN1(n9330), .IN2(n9947), .QN(n10613) );
  NAND2X0 U10590 ( .IN1(n10614), .IN2(n10615), .QN(n9947) );
  NAND2X0 U10591 ( .IN1(n7677), .IN2(n10616), .QN(n10615) );
  INVX0 U10592 ( .INP(n10617), .ZN(n10614) );
  NOR2X0 U10593 ( .IN1(n10616), .IN2(n7677), .QN(n10617) );
  NOR2X0 U10594 ( .IN1(n10618), .IN2(n10619), .QN(n10616) );
  NOR2X0 U10595 ( .IN1(WX9894), .IN2(n7678), .QN(n10619) );
  INVX0 U10596 ( .INP(n10620), .ZN(n10618) );
  NAND2X0 U10597 ( .IN1(n7678), .IN2(WX9894), .QN(n10620) );
  NAND2X0 U10598 ( .IN1(n9790), .IN2(n8317), .QN(n10612) );
  NAND2X0 U10599 ( .IN1(n16121), .IN2(n9079), .QN(n10611) );
  NAND2X0 U10600 ( .IN1(n10621), .IN2(n9110), .QN(n10605) );
  NAND2X0 U10601 ( .IN1(n1457), .IN2(n9275), .QN(n10604) );
  NOR2X0 U10602 ( .IN1(n9231), .IN2(n8883), .QN(n1457) );
  NAND2X0 U10603 ( .IN1(n9307), .IN2(CRC_OUT_3_28), .QN(n10603) );
  NAND4X0 U10604 ( .IN1(n10622), .IN2(n10623), .IN3(n10624), .IN4(n10625), 
        .QN(WX8406) );
  NAND2X0 U10605 ( .IN1(n10626), .IN2(n9959), .QN(n10625) );
  NAND2X0 U10606 ( .IN1(n10627), .IN2(n9962), .QN(n9959) );
  NAND2X0 U10607 ( .IN1(n10628), .IN2(n10629), .QN(n10627) );
  NAND2X0 U10608 ( .IN1(n16120), .IN2(n9119), .QN(n10629) );
  NAND2X0 U10609 ( .IN1(TM1), .IN2(n8318), .QN(n10628) );
  NAND3X0 U10610 ( .IN1(n10630), .IN2(n10631), .IN3(n10632), .QN(n10626) );
  NAND2X0 U10611 ( .IN1(n9330), .IN2(n9962), .QN(n10632) );
  NAND2X0 U10612 ( .IN1(n10633), .IN2(n10634), .QN(n9962) );
  NAND2X0 U10613 ( .IN1(n7679), .IN2(n10635), .QN(n10634) );
  INVX0 U10614 ( .INP(n10636), .ZN(n10633) );
  NOR2X0 U10615 ( .IN1(n10635), .IN2(n7679), .QN(n10636) );
  NOR2X0 U10616 ( .IN1(n10637), .IN2(n10638), .QN(n10635) );
  NOR2X0 U10617 ( .IN1(WX9892), .IN2(n7680), .QN(n10638) );
  INVX0 U10618 ( .INP(n10639), .ZN(n10637) );
  NAND2X0 U10619 ( .IN1(n7680), .IN2(WX9892), .QN(n10639) );
  NAND2X0 U10620 ( .IN1(n9083), .IN2(n8318), .QN(n10631) );
  NAND2X0 U10621 ( .IN1(n16120), .IN2(n9078), .QN(n10630) );
  NAND2X0 U10622 ( .IN1(n10640), .IN2(n10641), .QN(n10624) );
  NAND2X0 U10623 ( .IN1(n10642), .IN2(n10643), .QN(n10640) );
  NAND2X0 U10624 ( .IN1(n9096), .IN2(n10644), .QN(n10643) );
  NAND2X0 U10625 ( .IN1(n9096), .IN2(n8376), .QN(n10642) );
  NAND2X0 U10626 ( .IN1(n1456), .IN2(n9275), .QN(n10623) );
  NOR2X0 U10627 ( .IN1(n9231), .IN2(n8884), .QN(n1456) );
  NAND2X0 U10628 ( .IN1(n9307), .IN2(CRC_OUT_3_29), .QN(n10622) );
  NAND4X0 U10629 ( .IN1(n10645), .IN2(n10646), .IN3(n10647), .IN4(n10648), 
        .QN(WX8404) );
  NAND2X0 U10630 ( .IN1(n10649), .IN2(n9974), .QN(n10648) );
  NAND2X0 U10631 ( .IN1(n10650), .IN2(n9977), .QN(n9974) );
  NAND2X0 U10632 ( .IN1(n10651), .IN2(n10652), .QN(n10650) );
  NAND2X0 U10633 ( .IN1(n16119), .IN2(n9119), .QN(n10652) );
  NAND2X0 U10634 ( .IN1(TM1), .IN2(n8319), .QN(n10651) );
  NAND3X0 U10635 ( .IN1(n10653), .IN2(n10654), .IN3(n10655), .QN(n10649) );
  NAND2X0 U10636 ( .IN1(n9330), .IN2(n9977), .QN(n10655) );
  NAND2X0 U10637 ( .IN1(n10656), .IN2(n10657), .QN(n9977) );
  NAND2X0 U10638 ( .IN1(n7681), .IN2(n10658), .QN(n10657) );
  INVX0 U10639 ( .INP(n10659), .ZN(n10656) );
  NOR2X0 U10640 ( .IN1(n10658), .IN2(n7681), .QN(n10659) );
  NOR2X0 U10641 ( .IN1(n10660), .IN2(n10661), .QN(n10658) );
  NOR2X0 U10642 ( .IN1(WX9890), .IN2(n7682), .QN(n10661) );
  INVX0 U10643 ( .INP(n10662), .ZN(n10660) );
  NAND2X0 U10644 ( .IN1(n7682), .IN2(WX9890), .QN(n10662) );
  NAND2X0 U10645 ( .IN1(n9082), .IN2(n8319), .QN(n10654) );
  NAND2X0 U10646 ( .IN1(n16119), .IN2(n9077), .QN(n10653) );
  NAND2X0 U10647 ( .IN1(n10663), .IN2(n9110), .QN(n10647) );
  NAND2X0 U10648 ( .IN1(n1455), .IN2(n9275), .QN(n10646) );
  NOR2X0 U10649 ( .IN1(n9231), .IN2(n8885), .QN(n1455) );
  NAND2X0 U10650 ( .IN1(n9307), .IN2(CRC_OUT_3_30), .QN(n10645) );
  NAND4X0 U10651 ( .IN1(n10664), .IN2(n10665), .IN3(n10666), .IN4(n10667), 
        .QN(WX8402) );
  NAND2X0 U10652 ( .IN1(n10668), .IN2(n10669), .QN(n10667) );
  NAND2X0 U10653 ( .IN1(n10670), .IN2(n10671), .QN(n10668) );
  NAND2X0 U10654 ( .IN1(n9096), .IN2(n10672), .QN(n10671) );
  NAND2X0 U10655 ( .IN1(n9096), .IN2(n8378), .QN(n10670) );
  NAND2X0 U10656 ( .IN1(n9994), .IN2(n9334), .QN(n10666) );
  NOR2X0 U10657 ( .IN1(n10673), .IN2(n10674), .QN(n9994) );
  INVX0 U10658 ( .INP(n10675), .ZN(n10674) );
  NAND2X0 U10659 ( .IN1(n10676), .IN2(n10677), .QN(n10675) );
  NOR2X0 U10660 ( .IN1(n10677), .IN2(n10676), .QN(n10673) );
  NAND2X0 U10661 ( .IN1(n10678), .IN2(n10679), .QN(n10676) );
  NAND2X0 U10662 ( .IN1(n10680), .IN2(WX9824), .QN(n10679) );
  NAND2X0 U10663 ( .IN1(n10681), .IN2(n10682), .QN(n10680) );
  NAND3X0 U10664 ( .IN1(n10681), .IN2(n10682), .IN3(n7614), .QN(n10678) );
  NAND2X0 U10665 ( .IN1(test_so85), .IN2(WX9760), .QN(n10682) );
  NAND2X0 U10666 ( .IN1(n7613), .IN2(n8804), .QN(n10681) );
  NOR2X0 U10667 ( .IN1(n10683), .IN2(n10684), .QN(n10677) );
  INVX0 U10668 ( .INP(n10685), .ZN(n10684) );
  NAND2X0 U10669 ( .IN1(n16118), .IN2(n9119), .QN(n10685) );
  NOR2X0 U10670 ( .IN1(n9116), .IN2(n16118), .QN(n10683) );
  NAND2X0 U10671 ( .IN1(n9307), .IN2(CRC_OUT_3_31), .QN(n10665) );
  NAND2X0 U10672 ( .IN1(n2245), .IN2(WX8243), .QN(n10664) );
  NOR2X0 U10673 ( .IN1(n9231), .IN2(WX8243), .QN(WX8304) );
  NOR3X0 U10674 ( .IN1(n9144), .IN2(n10686), .IN3(n10687), .QN(WX7791) );
  NOR2X0 U10675 ( .IN1(n8211), .IN2(CRC_OUT_4_30), .QN(n10687) );
  NOR2X0 U10676 ( .IN1(DFF_1150_n1), .IN2(WX7302), .QN(n10686) );
  NOR2X0 U10677 ( .IN1(n9231), .IN2(n10688), .QN(WX7789) );
  NOR2X0 U10678 ( .IN1(n10689), .IN2(n10690), .QN(n10688) );
  NOR2X0 U10679 ( .IN1(test_so66), .IN2(WX7304), .QN(n10690) );
  INVX0 U10680 ( .INP(n10691), .ZN(n10689) );
  NAND2X0 U10681 ( .IN1(WX7304), .IN2(test_so66), .QN(n10691) );
  NOR3X0 U10682 ( .IN1(n9144), .IN2(n10692), .IN3(n10693), .QN(WX7787) );
  NOR2X0 U10683 ( .IN1(n8213), .IN2(CRC_OUT_4_28), .QN(n10693) );
  NOR2X0 U10684 ( .IN1(DFF_1148_n1), .IN2(WX7306), .QN(n10692) );
  NOR3X0 U10685 ( .IN1(n9144), .IN2(n10694), .IN3(n10695), .QN(WX7785) );
  NOR2X0 U10686 ( .IN1(n8214), .IN2(CRC_OUT_4_27), .QN(n10695) );
  NOR2X0 U10687 ( .IN1(DFF_1147_n1), .IN2(WX7308), .QN(n10694) );
  NOR3X0 U10688 ( .IN1(n9144), .IN2(n10696), .IN3(n10697), .QN(WX7783) );
  NOR2X0 U10689 ( .IN1(n8215), .IN2(CRC_OUT_4_26), .QN(n10697) );
  NOR2X0 U10690 ( .IN1(DFF_1146_n1), .IN2(WX7310), .QN(n10696) );
  NOR3X0 U10691 ( .IN1(n9144), .IN2(n10698), .IN3(n10699), .QN(WX7781) );
  NOR2X0 U10692 ( .IN1(n8216), .IN2(CRC_OUT_4_25), .QN(n10699) );
  NOR2X0 U10693 ( .IN1(DFF_1145_n1), .IN2(WX7312), .QN(n10698) );
  NOR3X0 U10694 ( .IN1(n9143), .IN2(n10700), .IN3(n10701), .QN(WX7779) );
  NOR2X0 U10695 ( .IN1(n8217), .IN2(CRC_OUT_4_24), .QN(n10701) );
  NOR2X0 U10696 ( .IN1(DFF_1144_n1), .IN2(WX7314), .QN(n10700) );
  NOR3X0 U10697 ( .IN1(n9143), .IN2(n10702), .IN3(n10703), .QN(WX7777) );
  NOR2X0 U10698 ( .IN1(n8218), .IN2(CRC_OUT_4_23), .QN(n10703) );
  NOR2X0 U10699 ( .IN1(DFF_1143_n1), .IN2(WX7316), .QN(n10702) );
  NOR3X0 U10700 ( .IN1(n9143), .IN2(n10704), .IN3(n10705), .QN(WX7775) );
  NOR2X0 U10701 ( .IN1(n8219), .IN2(CRC_OUT_4_22), .QN(n10705) );
  NOR2X0 U10702 ( .IN1(DFF_1142_n1), .IN2(WX7318), .QN(n10704) );
  NOR3X0 U10703 ( .IN1(n9143), .IN2(n10706), .IN3(n10707), .QN(WX7773) );
  NOR2X0 U10704 ( .IN1(n8220), .IN2(CRC_OUT_4_21), .QN(n10707) );
  NOR2X0 U10705 ( .IN1(DFF_1141_n1), .IN2(WX7320), .QN(n10706) );
  NOR2X0 U10706 ( .IN1(n9230), .IN2(n10708), .QN(WX7771) );
  NOR2X0 U10707 ( .IN1(n10709), .IN2(n10710), .QN(n10708) );
  NOR2X0 U10708 ( .IN1(test_so63), .IN2(CRC_OUT_4_20), .QN(n10710) );
  NOR2X0 U10709 ( .IN1(DFF_1140_n1), .IN2(n8799), .QN(n10709) );
  NOR3X0 U10710 ( .IN1(n9143), .IN2(n10711), .IN3(n10712), .QN(WX7769) );
  NOR2X0 U10711 ( .IN1(n8221), .IN2(CRC_OUT_4_19), .QN(n10712) );
  NOR2X0 U10712 ( .IN1(DFF_1139_n1), .IN2(WX7324), .QN(n10711) );
  NOR3X0 U10713 ( .IN1(n9143), .IN2(n10713), .IN3(n10714), .QN(WX7767) );
  NOR2X0 U10714 ( .IN1(n8222), .IN2(CRC_OUT_4_18), .QN(n10714) );
  NOR2X0 U10715 ( .IN1(DFF_1138_n1), .IN2(WX7326), .QN(n10713) );
  NOR3X0 U10716 ( .IN1(n9143), .IN2(n10715), .IN3(n10716), .QN(WX7765) );
  NOR2X0 U10717 ( .IN1(n8223), .IN2(CRC_OUT_4_17), .QN(n10716) );
  NOR2X0 U10718 ( .IN1(DFF_1137_n1), .IN2(WX7328), .QN(n10715) );
  NOR3X0 U10719 ( .IN1(n9143), .IN2(n10717), .IN3(n10718), .QN(WX7763) );
  NOR2X0 U10720 ( .IN1(n8224), .IN2(CRC_OUT_4_16), .QN(n10718) );
  NOR2X0 U10721 ( .IN1(DFF_1136_n1), .IN2(WX7330), .QN(n10717) );
  NOR2X0 U10722 ( .IN1(n9230), .IN2(n10719), .QN(WX7761) );
  NOR2X0 U10723 ( .IN1(n10720), .IN2(n10721), .QN(n10719) );
  INVX0 U10724 ( .INP(n10722), .ZN(n10721) );
  NAND2X0 U10725 ( .IN1(CRC_OUT_4_15), .IN2(n10723), .QN(n10722) );
  NOR2X0 U10726 ( .IN1(n10723), .IN2(CRC_OUT_4_15), .QN(n10720) );
  NAND2X0 U10727 ( .IN1(n10724), .IN2(n10725), .QN(n10723) );
  NAND2X0 U10728 ( .IN1(n8113), .IN2(CRC_OUT_4_31), .QN(n10725) );
  NAND2X0 U10729 ( .IN1(DFF_1151_n1), .IN2(WX7332), .QN(n10724) );
  NOR3X0 U10730 ( .IN1(n9143), .IN2(n10726), .IN3(n10727), .QN(WX7759) );
  NOR2X0 U10731 ( .IN1(n8225), .IN2(CRC_OUT_4_14), .QN(n10727) );
  NOR2X0 U10732 ( .IN1(DFF_1134_n1), .IN2(WX7334), .QN(n10726) );
  NOR3X0 U10733 ( .IN1(n9143), .IN2(n10728), .IN3(n10729), .QN(WX7757) );
  NOR2X0 U10734 ( .IN1(n8226), .IN2(CRC_OUT_4_13), .QN(n10729) );
  NOR2X0 U10735 ( .IN1(DFF_1133_n1), .IN2(WX7336), .QN(n10728) );
  NOR2X0 U10736 ( .IN1(n9229), .IN2(n10730), .QN(WX7755) );
  NOR2X0 U10737 ( .IN1(n10731), .IN2(n10732), .QN(n10730) );
  NOR2X0 U10738 ( .IN1(test_so65), .IN2(WX7338), .QN(n10732) );
  INVX0 U10739 ( .INP(n10733), .ZN(n10731) );
  NAND2X0 U10740 ( .IN1(WX7338), .IN2(test_so65), .QN(n10733) );
  NOR3X0 U10741 ( .IN1(n9143), .IN2(n10734), .IN3(n10735), .QN(WX7753) );
  NOR2X0 U10742 ( .IN1(n8228), .IN2(CRC_OUT_4_11), .QN(n10735) );
  NOR2X0 U10743 ( .IN1(DFF_1131_n1), .IN2(WX7340), .QN(n10734) );
  NOR2X0 U10744 ( .IN1(n9229), .IN2(n10736), .QN(WX7751) );
  NOR2X0 U10745 ( .IN1(n10737), .IN2(n10738), .QN(n10736) );
  INVX0 U10746 ( .INP(n10739), .ZN(n10738) );
  NAND2X0 U10747 ( .IN1(CRC_OUT_4_10), .IN2(n10740), .QN(n10739) );
  NOR2X0 U10748 ( .IN1(n10740), .IN2(CRC_OUT_4_10), .QN(n10737) );
  NAND2X0 U10749 ( .IN1(n10741), .IN2(n10742), .QN(n10740) );
  NAND2X0 U10750 ( .IN1(n8114), .IN2(CRC_OUT_4_31), .QN(n10742) );
  NAND2X0 U10751 ( .IN1(DFF_1151_n1), .IN2(WX7342), .QN(n10741) );
  NOR3X0 U10752 ( .IN1(n9143), .IN2(n10743), .IN3(n10744), .QN(WX7749) );
  NOR2X0 U10753 ( .IN1(n8229), .IN2(CRC_OUT_4_9), .QN(n10744) );
  NOR2X0 U10754 ( .IN1(DFF_1129_n1), .IN2(WX7344), .QN(n10743) );
  NOR3X0 U10755 ( .IN1(n9142), .IN2(n10745), .IN3(n10746), .QN(WX7747) );
  NOR2X0 U10756 ( .IN1(n8230), .IN2(CRC_OUT_4_8), .QN(n10746) );
  NOR2X0 U10757 ( .IN1(DFF_1128_n1), .IN2(WX7346), .QN(n10745) );
  NOR3X0 U10758 ( .IN1(n9142), .IN2(n10747), .IN3(n10748), .QN(WX7745) );
  NOR2X0 U10759 ( .IN1(n8231), .IN2(CRC_OUT_4_7), .QN(n10748) );
  NOR2X0 U10760 ( .IN1(DFF_1127_n1), .IN2(WX7348), .QN(n10747) );
  NOR3X0 U10761 ( .IN1(n9142), .IN2(n10749), .IN3(n10750), .QN(WX7743) );
  NOR2X0 U10762 ( .IN1(n8232), .IN2(CRC_OUT_4_6), .QN(n10750) );
  NOR2X0 U10763 ( .IN1(DFF_1126_n1), .IN2(WX7350), .QN(n10749) );
  NOR3X0 U10764 ( .IN1(n9142), .IN2(n10751), .IN3(n10752), .QN(WX7741) );
  NOR2X0 U10765 ( .IN1(n8233), .IN2(CRC_OUT_4_5), .QN(n10752) );
  NOR2X0 U10766 ( .IN1(DFF_1125_n1), .IN2(WX7352), .QN(n10751) );
  NOR3X0 U10767 ( .IN1(n9142), .IN2(n10753), .IN3(n10754), .QN(WX7739) );
  NOR2X0 U10768 ( .IN1(n8234), .IN2(CRC_OUT_4_4), .QN(n10754) );
  NOR2X0 U10769 ( .IN1(DFF_1124_n1), .IN2(WX7354), .QN(n10753) );
  NOR3X0 U10770 ( .IN1(n9142), .IN2(n10755), .IN3(n10756), .QN(WX7737) );
  INVX0 U10771 ( .INP(n10757), .ZN(n10756) );
  NAND2X0 U10772 ( .IN1(CRC_OUT_4_3), .IN2(n10758), .QN(n10757) );
  NOR2X0 U10773 ( .IN1(n10758), .IN2(CRC_OUT_4_3), .QN(n10755) );
  NAND2X0 U10774 ( .IN1(n10759), .IN2(n10760), .QN(n10758) );
  NAND2X0 U10775 ( .IN1(test_so64), .IN2(CRC_OUT_4_31), .QN(n10760) );
  NAND2X0 U10776 ( .IN1(DFF_1151_n1), .IN2(n8795), .QN(n10759) );
  NOR3X0 U10777 ( .IN1(n9142), .IN2(n10761), .IN3(n10762), .QN(WX7735) );
  NOR2X0 U10778 ( .IN1(n8235), .IN2(CRC_OUT_4_2), .QN(n10762) );
  NOR2X0 U10779 ( .IN1(DFF_1122_n1), .IN2(WX7358), .QN(n10761) );
  NOR3X0 U10780 ( .IN1(n9142), .IN2(n10763), .IN3(n10764), .QN(WX7733) );
  NOR2X0 U10781 ( .IN1(n8236), .IN2(CRC_OUT_4_1), .QN(n10764) );
  NOR2X0 U10782 ( .IN1(DFF_1121_n1), .IN2(WX7360), .QN(n10763) );
  NOR3X0 U10783 ( .IN1(n9142), .IN2(n10765), .IN3(n10766), .QN(WX7731) );
  NOR2X0 U10784 ( .IN1(n8237), .IN2(CRC_OUT_4_0), .QN(n10766) );
  NOR2X0 U10785 ( .IN1(DFF_1120_n1), .IN2(WX7362), .QN(n10765) );
  NOR3X0 U10786 ( .IN1(n9142), .IN2(n10767), .IN3(n10768), .QN(WX7729) );
  NOR2X0 U10787 ( .IN1(n8128), .IN2(CRC_OUT_4_31), .QN(n10768) );
  NOR2X0 U10788 ( .IN1(DFF_1151_n1), .IN2(WX7364), .QN(n10767) );
  NOR2X0 U10789 ( .IN1(n16101), .IN2(n9164), .QN(WX7203) );
  NOR2X0 U10790 ( .IN1(n16100), .IN2(n9164), .QN(WX7201) );
  NOR2X0 U10791 ( .IN1(n16099), .IN2(n9163), .QN(WX7199) );
  NOR2X0 U10792 ( .IN1(n16098), .IN2(n9164), .QN(WX7197) );
  NOR2X0 U10793 ( .IN1(n16097), .IN2(n9164), .QN(WX7195) );
  NOR2X0 U10794 ( .IN1(n16096), .IN2(n9163), .QN(WX7193) );
  NOR2X0 U10795 ( .IN1(n16095), .IN2(n9163), .QN(WX7191) );
  NOR2X0 U10796 ( .IN1(n16094), .IN2(n9163), .QN(WX7189) );
  NOR2X0 U10797 ( .IN1(n16093), .IN2(n9163), .QN(WX7187) );
  NOR2X0 U10798 ( .IN1(n16092), .IN2(n9163), .QN(WX7185) );
  NOR2X0 U10799 ( .IN1(n16091), .IN2(n9163), .QN(WX7183) );
  NOR2X0 U10800 ( .IN1(n9226), .IN2(n8820), .QN(WX7181) );
  NOR2X0 U10801 ( .IN1(n16090), .IN2(n9163), .QN(WX7179) );
  NOR2X0 U10802 ( .IN1(n16089), .IN2(n9163), .QN(WX7177) );
  NOR2X0 U10803 ( .IN1(n16088), .IN2(n9163), .QN(WX7175) );
  NOR2X0 U10804 ( .IN1(n16087), .IN2(n9163), .QN(WX7173) );
  NAND4X0 U10805 ( .IN1(n10769), .IN2(n10770), .IN3(n10771), .IN4(n10772), 
        .QN(WX7171) );
  NAND2X0 U10806 ( .IN1(n9330), .IN2(n10095), .QN(n10772) );
  NAND2X0 U10807 ( .IN1(n10773), .IN2(n10774), .QN(n10095) );
  INVX0 U10808 ( .INP(n10775), .ZN(n10774) );
  NOR2X0 U10809 ( .IN1(n10776), .IN2(n10777), .QN(n10775) );
  NAND2X0 U10810 ( .IN1(n10777), .IN2(n10776), .QN(n10773) );
  NOR2X0 U10811 ( .IN1(n10778), .IN2(n10779), .QN(n10776) );
  NOR2X0 U10812 ( .IN1(WX8657), .IN2(n7915), .QN(n10779) );
  INVX0 U10813 ( .INP(n10780), .ZN(n10778) );
  NAND2X0 U10814 ( .IN1(n7915), .IN2(WX8657), .QN(n10780) );
  NAND2X0 U10815 ( .IN1(n10781), .IN2(n10782), .QN(n10777) );
  NAND2X0 U10816 ( .IN1(n7914), .IN2(WX8529), .QN(n10782) );
  INVX0 U10817 ( .INP(n10783), .ZN(n10781) );
  NOR2X0 U10818 ( .IN1(WX8529), .IN2(n7914), .QN(n10783) );
  NAND2X0 U10819 ( .IN1(n9096), .IN2(n10784), .QN(n10771) );
  NAND2X0 U10820 ( .IN1(n1244), .IN2(n9275), .QN(n10770) );
  NOR2X0 U10821 ( .IN1(n9226), .IN2(n8886), .QN(n1244) );
  NAND2X0 U10822 ( .IN1(n9307), .IN2(CRC_OUT_4_0), .QN(n10769) );
  NAND4X0 U10823 ( .IN1(n10785), .IN2(n10786), .IN3(n10787), .IN4(n10788), 
        .QN(WX7169) );
  NAND2X0 U10824 ( .IN1(n9330), .IN2(n10108), .QN(n10788) );
  NAND2X0 U10825 ( .IN1(n10789), .IN2(n10790), .QN(n10108) );
  INVX0 U10826 ( .INP(n10791), .ZN(n10790) );
  NOR2X0 U10827 ( .IN1(n10792), .IN2(n10793), .QN(n10791) );
  NAND2X0 U10828 ( .IN1(n10793), .IN2(n10792), .QN(n10789) );
  NOR2X0 U10829 ( .IN1(n10794), .IN2(n10795), .QN(n10792) );
  NOR2X0 U10830 ( .IN1(WX8655), .IN2(n7917), .QN(n10795) );
  INVX0 U10831 ( .INP(n10796), .ZN(n10794) );
  NAND2X0 U10832 ( .IN1(n7917), .IN2(WX8655), .QN(n10796) );
  NAND2X0 U10833 ( .IN1(n10797), .IN2(n10798), .QN(n10793) );
  NAND2X0 U10834 ( .IN1(n7916), .IN2(WX8527), .QN(n10798) );
  INVX0 U10835 ( .INP(n10799), .ZN(n10797) );
  NOR2X0 U10836 ( .IN1(WX8527), .IN2(n7916), .QN(n10799) );
  NAND2X0 U10837 ( .IN1(n9096), .IN2(n10800), .QN(n10787) );
  NAND2X0 U10838 ( .IN1(n1243), .IN2(n9275), .QN(n10786) );
  NOR2X0 U10839 ( .IN1(n9226), .IN2(n8887), .QN(n1243) );
  NAND2X0 U10840 ( .IN1(n9307), .IN2(CRC_OUT_4_1), .QN(n10785) );
  NAND4X0 U10841 ( .IN1(n10801), .IN2(n10802), .IN3(n10803), .IN4(n10804), 
        .QN(WX7167) );
  NAND2X0 U10842 ( .IN1(n9330), .IN2(n10124), .QN(n10804) );
  NAND2X0 U10843 ( .IN1(n10805), .IN2(n10806), .QN(n10124) );
  INVX0 U10844 ( .INP(n10807), .ZN(n10806) );
  NOR2X0 U10845 ( .IN1(n10808), .IN2(n10809), .QN(n10807) );
  NAND2X0 U10846 ( .IN1(n10809), .IN2(n10808), .QN(n10805) );
  NOR2X0 U10847 ( .IN1(n10810), .IN2(n10811), .QN(n10808) );
  NOR2X0 U10848 ( .IN1(WX8653), .IN2(n7919), .QN(n10811) );
  INVX0 U10849 ( .INP(n10812), .ZN(n10810) );
  NAND2X0 U10850 ( .IN1(n7919), .IN2(WX8653), .QN(n10812) );
  NAND2X0 U10851 ( .IN1(n10813), .IN2(n10814), .QN(n10809) );
  NAND2X0 U10852 ( .IN1(n7918), .IN2(WX8525), .QN(n10814) );
  INVX0 U10853 ( .INP(n10815), .ZN(n10813) );
  NOR2X0 U10854 ( .IN1(WX8525), .IN2(n7918), .QN(n10815) );
  NAND2X0 U10855 ( .IN1(n9096), .IN2(n10816), .QN(n10803) );
  NAND2X0 U10856 ( .IN1(n1242), .IN2(n9275), .QN(n10802) );
  NOR2X0 U10857 ( .IN1(n9226), .IN2(n8888), .QN(n1242) );
  NAND2X0 U10858 ( .IN1(n9307), .IN2(CRC_OUT_4_2), .QN(n10801) );
  NAND4X0 U10859 ( .IN1(n10817), .IN2(n10818), .IN3(n10819), .IN4(n10820), 
        .QN(WX7165) );
  NAND2X0 U10860 ( .IN1(n9330), .IN2(n10137), .QN(n10820) );
  NAND2X0 U10861 ( .IN1(n10821), .IN2(n10822), .QN(n10137) );
  INVX0 U10862 ( .INP(n10823), .ZN(n10822) );
  NOR2X0 U10863 ( .IN1(n10824), .IN2(n10825), .QN(n10823) );
  NAND2X0 U10864 ( .IN1(n10825), .IN2(n10824), .QN(n10821) );
  NOR2X0 U10865 ( .IN1(n10826), .IN2(n10827), .QN(n10824) );
  NOR2X0 U10866 ( .IN1(WX8651), .IN2(n7921), .QN(n10827) );
  INVX0 U10867 ( .INP(n10828), .ZN(n10826) );
  NAND2X0 U10868 ( .IN1(n7921), .IN2(WX8651), .QN(n10828) );
  NAND2X0 U10869 ( .IN1(n10829), .IN2(n10830), .QN(n10825) );
  NAND2X0 U10870 ( .IN1(n7920), .IN2(WX8523), .QN(n10830) );
  INVX0 U10871 ( .INP(n10831), .ZN(n10829) );
  NOR2X0 U10872 ( .IN1(WX8523), .IN2(n7920), .QN(n10831) );
  NAND2X0 U10873 ( .IN1(n9096), .IN2(n10832), .QN(n10819) );
  NAND2X0 U10874 ( .IN1(n1241), .IN2(n9275), .QN(n10818) );
  NOR2X0 U10875 ( .IN1(n9226), .IN2(n8889), .QN(n1241) );
  NAND2X0 U10876 ( .IN1(n9307), .IN2(CRC_OUT_4_3), .QN(n10817) );
  NAND4X0 U10877 ( .IN1(n10833), .IN2(n10834), .IN3(n10835), .IN4(n10836), 
        .QN(WX7163) );
  NAND3X0 U10878 ( .IN1(n10837), .IN2(n10838), .IN3(n9089), .QN(n10836) );
  NAND2X0 U10879 ( .IN1(n9331), .IN2(n10153), .QN(n10835) );
  NAND2X0 U10880 ( .IN1(n10839), .IN2(n10840), .QN(n10153) );
  INVX0 U10881 ( .INP(n10841), .ZN(n10840) );
  NOR2X0 U10882 ( .IN1(n10842), .IN2(n10843), .QN(n10841) );
  NAND2X0 U10883 ( .IN1(n10843), .IN2(n10842), .QN(n10839) );
  NOR2X0 U10884 ( .IN1(n10844), .IN2(n10845), .QN(n10842) );
  NOR2X0 U10885 ( .IN1(WX8649), .IN2(n7923), .QN(n10845) );
  INVX0 U10886 ( .INP(n10846), .ZN(n10844) );
  NAND2X0 U10887 ( .IN1(n7923), .IN2(WX8649), .QN(n10846) );
  NAND2X0 U10888 ( .IN1(n10847), .IN2(n10848), .QN(n10843) );
  NAND2X0 U10889 ( .IN1(n7922), .IN2(WX8521), .QN(n10848) );
  INVX0 U10890 ( .INP(n10849), .ZN(n10847) );
  NOR2X0 U10891 ( .IN1(WX8521), .IN2(n7922), .QN(n10849) );
  NAND2X0 U10892 ( .IN1(n1240), .IN2(n9275), .QN(n10834) );
  NOR2X0 U10893 ( .IN1(n9224), .IN2(n8890), .QN(n1240) );
  NAND2X0 U10894 ( .IN1(n9307), .IN2(CRC_OUT_4_4), .QN(n10833) );
  NAND4X0 U10895 ( .IN1(n10850), .IN2(n10851), .IN3(n10852), .IN4(n10853), 
        .QN(WX7161) );
  NAND2X0 U10896 ( .IN1(n9331), .IN2(n10169), .QN(n10853) );
  NAND2X0 U10897 ( .IN1(n10854), .IN2(n10855), .QN(n10169) );
  INVX0 U10898 ( .INP(n10856), .ZN(n10855) );
  NOR2X0 U10899 ( .IN1(n10857), .IN2(n10858), .QN(n10856) );
  NAND2X0 U10900 ( .IN1(n10858), .IN2(n10857), .QN(n10854) );
  NOR2X0 U10901 ( .IN1(n10859), .IN2(n10860), .QN(n10857) );
  NOR2X0 U10902 ( .IN1(WX8647), .IN2(n7925), .QN(n10860) );
  INVX0 U10903 ( .INP(n10861), .ZN(n10859) );
  NAND2X0 U10904 ( .IN1(n7925), .IN2(WX8647), .QN(n10861) );
  NAND2X0 U10905 ( .IN1(n10862), .IN2(n10863), .QN(n10858) );
  NAND2X0 U10906 ( .IN1(n7924), .IN2(WX8519), .QN(n10863) );
  INVX0 U10907 ( .INP(n10864), .ZN(n10862) );
  NOR2X0 U10908 ( .IN1(WX8519), .IN2(n7924), .QN(n10864) );
  NAND2X0 U10909 ( .IN1(n9096), .IN2(n10865), .QN(n10852) );
  NAND2X0 U10910 ( .IN1(n1239), .IN2(n9276), .QN(n10851) );
  NOR2X0 U10911 ( .IN1(n9223), .IN2(n8891), .QN(n1239) );
  NAND2X0 U10912 ( .IN1(n9307), .IN2(CRC_OUT_4_5), .QN(n10850) );
  NAND4X0 U10913 ( .IN1(n10866), .IN2(n10867), .IN3(n10868), .IN4(n10869), 
        .QN(WX7159) );
  NAND3X0 U10914 ( .IN1(n10870), .IN2(n10871), .IN3(n9089), .QN(n10869) );
  NAND2X0 U10915 ( .IN1(n9331), .IN2(n10185), .QN(n10868) );
  NAND2X0 U10916 ( .IN1(n10872), .IN2(n10873), .QN(n10185) );
  INVX0 U10917 ( .INP(n10874), .ZN(n10873) );
  NOR2X0 U10918 ( .IN1(n10875), .IN2(n10876), .QN(n10874) );
  NAND2X0 U10919 ( .IN1(n10876), .IN2(n10875), .QN(n10872) );
  NOR2X0 U10920 ( .IN1(n10877), .IN2(n10878), .QN(n10875) );
  NOR2X0 U10921 ( .IN1(WX8645), .IN2(n7927), .QN(n10878) );
  INVX0 U10922 ( .INP(n10879), .ZN(n10877) );
  NAND2X0 U10923 ( .IN1(n7927), .IN2(WX8645), .QN(n10879) );
  NAND2X0 U10924 ( .IN1(n10880), .IN2(n10881), .QN(n10876) );
  NAND2X0 U10925 ( .IN1(n7926), .IN2(WX8517), .QN(n10881) );
  INVX0 U10926 ( .INP(n10882), .ZN(n10880) );
  NOR2X0 U10927 ( .IN1(WX8517), .IN2(n7926), .QN(n10882) );
  NAND2X0 U10928 ( .IN1(n1238), .IN2(n9276), .QN(n10867) );
  NOR2X0 U10929 ( .IN1(n9223), .IN2(n8892), .QN(n1238) );
  NAND2X0 U10930 ( .IN1(n9308), .IN2(CRC_OUT_4_6), .QN(n10866) );
  NAND4X0 U10931 ( .IN1(n10883), .IN2(n10884), .IN3(n10885), .IN4(n10886), 
        .QN(WX7157) );
  NAND2X0 U10932 ( .IN1(n9331), .IN2(n10201), .QN(n10886) );
  NAND2X0 U10933 ( .IN1(n10887), .IN2(n10888), .QN(n10201) );
  INVX0 U10934 ( .INP(n10889), .ZN(n10888) );
  NOR2X0 U10935 ( .IN1(n10890), .IN2(n10891), .QN(n10889) );
  NAND2X0 U10936 ( .IN1(n10891), .IN2(n10890), .QN(n10887) );
  NOR2X0 U10937 ( .IN1(n10892), .IN2(n10893), .QN(n10890) );
  NOR2X0 U10938 ( .IN1(WX8643), .IN2(n7929), .QN(n10893) );
  INVX0 U10939 ( .INP(n10894), .ZN(n10892) );
  NAND2X0 U10940 ( .IN1(n7929), .IN2(WX8643), .QN(n10894) );
  NAND2X0 U10941 ( .IN1(n10895), .IN2(n10896), .QN(n10891) );
  NAND2X0 U10942 ( .IN1(n7928), .IN2(WX8515), .QN(n10896) );
  INVX0 U10943 ( .INP(n10897), .ZN(n10895) );
  NOR2X0 U10944 ( .IN1(WX8515), .IN2(n7928), .QN(n10897) );
  NAND2X0 U10945 ( .IN1(n9096), .IN2(n10898), .QN(n10885) );
  NAND2X0 U10946 ( .IN1(n1237), .IN2(n9276), .QN(n10884) );
  NOR2X0 U10947 ( .IN1(n9223), .IN2(n8893), .QN(n1237) );
  NAND2X0 U10948 ( .IN1(n9308), .IN2(CRC_OUT_4_7), .QN(n10883) );
  NAND4X0 U10949 ( .IN1(n10899), .IN2(n10900), .IN3(n10901), .IN4(n10902), 
        .QN(WX7155) );
  NAND3X0 U10950 ( .IN1(n10903), .IN2(n10904), .IN3(n9089), .QN(n10902) );
  NAND2X0 U10951 ( .IN1(n9331), .IN2(n10217), .QN(n10901) );
  NAND2X0 U10952 ( .IN1(n10905), .IN2(n10906), .QN(n10217) );
  INVX0 U10953 ( .INP(n10907), .ZN(n10906) );
  NOR2X0 U10954 ( .IN1(n10908), .IN2(n10909), .QN(n10907) );
  NAND2X0 U10955 ( .IN1(n10909), .IN2(n10908), .QN(n10905) );
  NOR2X0 U10956 ( .IN1(n10910), .IN2(n10911), .QN(n10908) );
  NOR2X0 U10957 ( .IN1(WX8641), .IN2(n7931), .QN(n10911) );
  INVX0 U10958 ( .INP(n10912), .ZN(n10910) );
  NAND2X0 U10959 ( .IN1(n7931), .IN2(WX8641), .QN(n10912) );
  NAND2X0 U10960 ( .IN1(n10913), .IN2(n10914), .QN(n10909) );
  NAND2X0 U10961 ( .IN1(n7930), .IN2(WX8513), .QN(n10914) );
  INVX0 U10962 ( .INP(n10915), .ZN(n10913) );
  NOR2X0 U10963 ( .IN1(WX8513), .IN2(n7930), .QN(n10915) );
  NAND2X0 U10964 ( .IN1(n1236), .IN2(n9276), .QN(n10900) );
  NOR2X0 U10965 ( .IN1(n9223), .IN2(n8894), .QN(n1236) );
  NAND2X0 U10966 ( .IN1(n9308), .IN2(CRC_OUT_4_8), .QN(n10899) );
  NAND4X0 U10967 ( .IN1(n10916), .IN2(n10917), .IN3(n10918), .IN4(n10919), 
        .QN(WX7153) );
  NAND3X0 U10968 ( .IN1(n10222), .IN2(n10223), .IN3(n9322), .QN(n10919) );
  NAND3X0 U10969 ( .IN1(n10920), .IN2(n10921), .IN3(n10922), .QN(n10223) );
  INVX0 U10970 ( .INP(n10923), .ZN(n10922) );
  NAND2X0 U10971 ( .IN1(n10923), .IN2(n10924), .QN(n10222) );
  NAND2X0 U10972 ( .IN1(n10920), .IN2(n10921), .QN(n10924) );
  NAND2X0 U10973 ( .IN1(n7933), .IN2(WX8511), .QN(n10921) );
  NAND2X0 U10974 ( .IN1(n3613), .IN2(WX8575), .QN(n10920) );
  NOR2X0 U10975 ( .IN1(n10925), .IN2(n10926), .QN(n10923) );
  NOR2X0 U10976 ( .IN1(n8790), .IN2(n7932), .QN(n10926) );
  INVX0 U10977 ( .INP(n10927), .ZN(n10925) );
  NAND2X0 U10978 ( .IN1(n7932), .IN2(n8790), .QN(n10927) );
  NAND2X0 U10979 ( .IN1(n9095), .IN2(n10928), .QN(n10918) );
  NAND2X0 U10980 ( .IN1(n1235), .IN2(n9276), .QN(n10917) );
  NOR2X0 U10981 ( .IN1(n9223), .IN2(n8895), .QN(n1235) );
  NAND2X0 U10982 ( .IN1(n9308), .IN2(CRC_OUT_4_9), .QN(n10916) );
  NAND4X0 U10983 ( .IN1(n10929), .IN2(n10930), .IN3(n10931), .IN4(n10932), 
        .QN(WX7151) );
  NAND3X0 U10984 ( .IN1(n10933), .IN2(n10934), .IN3(n9089), .QN(n10932) );
  NAND2X0 U10985 ( .IN1(n9331), .IN2(n10250), .QN(n10931) );
  NAND2X0 U10986 ( .IN1(n10935), .IN2(n10936), .QN(n10250) );
  INVX0 U10987 ( .INP(n10937), .ZN(n10936) );
  NOR2X0 U10988 ( .IN1(n10938), .IN2(n10939), .QN(n10937) );
  NAND2X0 U10989 ( .IN1(n10939), .IN2(n10938), .QN(n10935) );
  NOR2X0 U10990 ( .IN1(n10940), .IN2(n10941), .QN(n10938) );
  NOR2X0 U10991 ( .IN1(WX8637), .IN2(n7935), .QN(n10941) );
  INVX0 U10992 ( .INP(n10942), .ZN(n10940) );
  NAND2X0 U10993 ( .IN1(n7935), .IN2(WX8637), .QN(n10942) );
  NAND2X0 U10994 ( .IN1(n10943), .IN2(n10944), .QN(n10939) );
  NAND2X0 U10995 ( .IN1(n7934), .IN2(WX8509), .QN(n10944) );
  INVX0 U10996 ( .INP(n10945), .ZN(n10943) );
  NOR2X0 U10997 ( .IN1(WX8509), .IN2(n7934), .QN(n10945) );
  NAND2X0 U10998 ( .IN1(n1234), .IN2(n9276), .QN(n10930) );
  NOR2X0 U10999 ( .IN1(n9223), .IN2(n8896), .QN(n1234) );
  NAND2X0 U11000 ( .IN1(n9308), .IN2(CRC_OUT_4_10), .QN(n10929) );
  NAND4X0 U11001 ( .IN1(n10946), .IN2(n10947), .IN3(n10948), .IN4(n10949), 
        .QN(WX7149) );
  NAND3X0 U11002 ( .IN1(n10255), .IN2(n10256), .IN3(n9322), .QN(n10949) );
  NAND3X0 U11003 ( .IN1(n10950), .IN2(n10951), .IN3(n10952), .QN(n10256) );
  INVX0 U11004 ( .INP(n10953), .ZN(n10952) );
  NAND2X0 U11005 ( .IN1(n10953), .IN2(n10954), .QN(n10255) );
  NAND2X0 U11006 ( .IN1(n10950), .IN2(n10951), .QN(n10954) );
  NAND2X0 U11007 ( .IN1(n8111), .IN2(WX8507), .QN(n10951) );
  NAND2X0 U11008 ( .IN1(n3617), .IN2(WX8635), .QN(n10950) );
  NOR2X0 U11009 ( .IN1(n10955), .IN2(n10956), .QN(n10953) );
  INVX0 U11010 ( .INP(n10957), .ZN(n10956) );
  NAND2X0 U11011 ( .IN1(test_so73), .IN2(WX8443), .QN(n10957) );
  NOR2X0 U11012 ( .IN1(WX8443), .IN2(test_so73), .QN(n10955) );
  NAND2X0 U11013 ( .IN1(n9095), .IN2(n10958), .QN(n10948) );
  NAND2X0 U11014 ( .IN1(n1233), .IN2(n9276), .QN(n10947) );
  NOR2X0 U11015 ( .IN1(n9223), .IN2(n8897), .QN(n1233) );
  NAND2X0 U11016 ( .IN1(n9308), .IN2(CRC_OUT_4_11), .QN(n10946) );
  NAND4X0 U11017 ( .IN1(n10959), .IN2(n10960), .IN3(n10961), .IN4(n10962), 
        .QN(WX7147) );
  NAND2X0 U11018 ( .IN1(n9331), .IN2(n10283), .QN(n10962) );
  NAND2X0 U11019 ( .IN1(n10963), .IN2(n10964), .QN(n10283) );
  INVX0 U11020 ( .INP(n10965), .ZN(n10964) );
  NOR2X0 U11021 ( .IN1(n10966), .IN2(n10967), .QN(n10965) );
  NAND2X0 U11022 ( .IN1(n10967), .IN2(n10966), .QN(n10963) );
  NOR2X0 U11023 ( .IN1(n10968), .IN2(n10969), .QN(n10966) );
  NOR2X0 U11024 ( .IN1(WX8633), .IN2(n7938), .QN(n10969) );
  INVX0 U11025 ( .INP(n10970), .ZN(n10968) );
  NAND2X0 U11026 ( .IN1(n7938), .IN2(WX8633), .QN(n10970) );
  NAND2X0 U11027 ( .IN1(n10971), .IN2(n10972), .QN(n10967) );
  NAND2X0 U11028 ( .IN1(n7937), .IN2(WX8505), .QN(n10972) );
  INVX0 U11029 ( .INP(n10973), .ZN(n10971) );
  NOR2X0 U11030 ( .IN1(WX8505), .IN2(n7937), .QN(n10973) );
  NAND2X0 U11031 ( .IN1(n9095), .IN2(n10974), .QN(n10961) );
  NAND2X0 U11032 ( .IN1(n1232), .IN2(n9276), .QN(n10960) );
  NOR2X0 U11033 ( .IN1(n9064), .IN2(n9163), .QN(n1232) );
  NAND2X0 U11034 ( .IN1(test_so65), .IN2(n9313), .QN(n10959) );
  NAND4X0 U11035 ( .IN1(n10975), .IN2(n10976), .IN3(n10977), .IN4(n10978), 
        .QN(WX7145) );
  NAND3X0 U11036 ( .IN1(n10288), .IN2(n10289), .IN3(n9322), .QN(n10978) );
  NAND3X0 U11037 ( .IN1(n10979), .IN2(n10980), .IN3(n10981), .QN(n10289) );
  INVX0 U11038 ( .INP(n10982), .ZN(n10981) );
  NAND2X0 U11039 ( .IN1(n10982), .IN2(n10983), .QN(n10288) );
  NAND2X0 U11040 ( .IN1(n10979), .IN2(n10980), .QN(n10983) );
  NAND2X0 U11041 ( .IN1(n8201), .IN2(WX8567), .QN(n10980) );
  NAND2X0 U11042 ( .IN1(n7940), .IN2(WX8631), .QN(n10979) );
  NOR2X0 U11043 ( .IN1(n10984), .IN2(n10985), .QN(n10982) );
  INVX0 U11044 ( .INP(n10986), .ZN(n10985) );
  NAND2X0 U11045 ( .IN1(test_so71), .IN2(WX8439), .QN(n10986) );
  NOR2X0 U11046 ( .IN1(WX8439), .IN2(test_so71), .QN(n10984) );
  NAND2X0 U11047 ( .IN1(n9095), .IN2(n10987), .QN(n10977) );
  NAND2X0 U11048 ( .IN1(n1231), .IN2(n9276), .QN(n10976) );
  NOR2X0 U11049 ( .IN1(n9223), .IN2(n8898), .QN(n1231) );
  NAND2X0 U11050 ( .IN1(n9308), .IN2(CRC_OUT_4_13), .QN(n10975) );
  NAND4X0 U11051 ( .IN1(n10988), .IN2(n10989), .IN3(n10990), .IN4(n10991), 
        .QN(WX7143) );
  NAND2X0 U11052 ( .IN1(n9331), .IN2(n10313), .QN(n10991) );
  NAND2X0 U11053 ( .IN1(n10992), .IN2(n10993), .QN(n10313) );
  INVX0 U11054 ( .INP(n10994), .ZN(n10993) );
  NOR2X0 U11055 ( .IN1(n10995), .IN2(n10996), .QN(n10994) );
  NAND2X0 U11056 ( .IN1(n10996), .IN2(n10995), .QN(n10992) );
  NOR2X0 U11057 ( .IN1(n10997), .IN2(n10998), .QN(n10995) );
  NOR2X0 U11058 ( .IN1(WX8629), .IN2(n7942), .QN(n10998) );
  INVX0 U11059 ( .INP(n10999), .ZN(n10997) );
  NAND2X0 U11060 ( .IN1(n7942), .IN2(WX8629), .QN(n10999) );
  NAND2X0 U11061 ( .IN1(n11000), .IN2(n11001), .QN(n10996) );
  NAND2X0 U11062 ( .IN1(n7941), .IN2(WX8501), .QN(n11001) );
  INVX0 U11063 ( .INP(n11002), .ZN(n11000) );
  NOR2X0 U11064 ( .IN1(WX8501), .IN2(n7941), .QN(n11002) );
  NAND2X0 U11065 ( .IN1(n9095), .IN2(n11003), .QN(n10990) );
  NAND2X0 U11066 ( .IN1(n1230), .IN2(n9276), .QN(n10989) );
  NOR2X0 U11067 ( .IN1(n9223), .IN2(n8899), .QN(n1230) );
  NAND2X0 U11068 ( .IN1(n9308), .IN2(CRC_OUT_4_14), .QN(n10988) );
  NAND4X0 U11069 ( .IN1(n11004), .IN2(n11005), .IN3(n11006), .IN4(n11007), 
        .QN(WX7141) );
  NAND3X0 U11070 ( .IN1(n10318), .IN2(n10319), .IN3(n9321), .QN(n11007) );
  NAND3X0 U11071 ( .IN1(n11008), .IN2(n11009), .IN3(n11010), .QN(n10319) );
  INVX0 U11072 ( .INP(n11011), .ZN(n11010) );
  NAND2X0 U11073 ( .IN1(n11011), .IN2(n11012), .QN(n10318) );
  NAND2X0 U11074 ( .IN1(n11008), .IN2(n11009), .QN(n11012) );
  NAND2X0 U11075 ( .IN1(n8199), .IN2(WX8499), .QN(n11009) );
  NAND2X0 U11076 ( .IN1(n3625), .IN2(WX8627), .QN(n11008) );
  NOR2X0 U11077 ( .IN1(n11013), .IN2(n11014), .QN(n11011) );
  INVX0 U11078 ( .INP(n11015), .ZN(n11014) );
  NAND2X0 U11079 ( .IN1(test_so69), .IN2(WX8563), .QN(n11015) );
  NOR2X0 U11080 ( .IN1(WX8563), .IN2(test_so69), .QN(n11013) );
  NAND2X0 U11081 ( .IN1(n9093), .IN2(n11016), .QN(n11006) );
  NAND2X0 U11082 ( .IN1(n1229), .IN2(n9276), .QN(n11005) );
  NOR2X0 U11083 ( .IN1(n9224), .IN2(n8900), .QN(n1229) );
  NAND2X0 U11084 ( .IN1(n9308), .IN2(CRC_OUT_4_15), .QN(n11004) );
  NAND4X0 U11085 ( .IN1(n11017), .IN2(n11018), .IN3(n11019), .IN4(n11020), 
        .QN(WX7139) );
  NAND2X0 U11086 ( .IN1(n11021), .IN2(n10336), .QN(n11020) );
  NAND2X0 U11087 ( .IN1(n11022), .IN2(n10339), .QN(n10336) );
  NAND2X0 U11088 ( .IN1(n11023), .IN2(n11024), .QN(n11022) );
  NAND2X0 U11089 ( .IN1(n16117), .IN2(n9119), .QN(n11024) );
  NAND2X0 U11090 ( .IN1(TM1), .IN2(n8363), .QN(n11023) );
  NAND3X0 U11091 ( .IN1(n11025), .IN2(n11026), .IN3(n11027), .QN(n11021) );
  NAND2X0 U11092 ( .IN1(n9331), .IN2(n10339), .QN(n11027) );
  NAND2X0 U11093 ( .IN1(n11028), .IN2(n11029), .QN(n10339) );
  NAND2X0 U11094 ( .IN1(n7683), .IN2(n11030), .QN(n11029) );
  INVX0 U11095 ( .INP(n11031), .ZN(n11028) );
  NOR2X0 U11096 ( .IN1(n11030), .IN2(n7683), .QN(n11031) );
  NOR2X0 U11097 ( .IN1(n11032), .IN2(n11033), .QN(n11030) );
  NOR2X0 U11098 ( .IN1(WX8625), .IN2(n7684), .QN(n11033) );
  INVX0 U11099 ( .INP(n11034), .ZN(n11032) );
  NAND2X0 U11100 ( .IN1(n7684), .IN2(WX8625), .QN(n11034) );
  NAND2X0 U11101 ( .IN1(n9081), .IN2(n8363), .QN(n11026) );
  NAND2X0 U11102 ( .IN1(n16117), .IN2(n9791), .QN(n11025) );
  NAND2X0 U11103 ( .IN1(n11035), .IN2(n11036), .QN(n11019) );
  NAND2X0 U11104 ( .IN1(n11037), .IN2(n11038), .QN(n11035) );
  NAND2X0 U11105 ( .IN1(n9091), .IN2(n11039), .QN(n11038) );
  NAND2X0 U11106 ( .IN1(n9091), .IN2(n8421), .QN(n11037) );
  NAND2X0 U11107 ( .IN1(n1228), .IN2(n9276), .QN(n11018) );
  NOR2X0 U11108 ( .IN1(n9224), .IN2(n8901), .QN(n1228) );
  NAND2X0 U11109 ( .IN1(n9309), .IN2(CRC_OUT_4_16), .QN(n11017) );
  NAND4X0 U11110 ( .IN1(n11040), .IN2(n11041), .IN3(n11042), .IN4(n11043), 
        .QN(WX7137) );
  NAND2X0 U11111 ( .IN1(n11044), .IN2(n10375), .QN(n11043) );
  NAND2X0 U11112 ( .IN1(n11045), .IN2(n10378), .QN(n10375) );
  NAND2X0 U11113 ( .IN1(n11046), .IN2(n11047), .QN(n11045) );
  NAND2X0 U11114 ( .IN1(n16116), .IN2(n9119), .QN(n11047) );
  NAND2X0 U11115 ( .IN1(TM1), .IN2(n8364), .QN(n11046) );
  NAND3X0 U11116 ( .IN1(n11048), .IN2(n11049), .IN3(n11050), .QN(n11044) );
  NAND2X0 U11117 ( .IN1(n9331), .IN2(n10378), .QN(n11050) );
  NAND2X0 U11118 ( .IN1(n11051), .IN2(n11052), .QN(n10378) );
  NAND2X0 U11119 ( .IN1(n7685), .IN2(n11053), .QN(n11052) );
  INVX0 U11120 ( .INP(n11054), .ZN(n11051) );
  NOR2X0 U11121 ( .IN1(n11053), .IN2(n7685), .QN(n11054) );
  NOR2X0 U11122 ( .IN1(n11055), .IN2(n11056), .QN(n11053) );
  NOR2X0 U11123 ( .IN1(WX8623), .IN2(n7686), .QN(n11056) );
  INVX0 U11124 ( .INP(n11057), .ZN(n11055) );
  NAND2X0 U11125 ( .IN1(n7686), .IN2(WX8623), .QN(n11057) );
  NAND2X0 U11126 ( .IN1(n9790), .IN2(n8364), .QN(n11049) );
  NAND2X0 U11127 ( .IN1(n16116), .IN2(n9079), .QN(n11048) );
  NAND2X0 U11128 ( .IN1(n11058), .IN2(n11059), .QN(n11042) );
  NAND2X0 U11129 ( .IN1(n11060), .IN2(n11061), .QN(n11058) );
  NAND2X0 U11130 ( .IN1(n9091), .IN2(n11062), .QN(n11061) );
  NAND2X0 U11131 ( .IN1(n9092), .IN2(n8422), .QN(n11060) );
  NAND2X0 U11132 ( .IN1(n1227), .IN2(n9276), .QN(n11041) );
  NOR2X0 U11133 ( .IN1(n9224), .IN2(n8902), .QN(n1227) );
  NAND2X0 U11134 ( .IN1(n9309), .IN2(CRC_OUT_4_17), .QN(n11040) );
  NAND4X0 U11135 ( .IN1(n11063), .IN2(n11064), .IN3(n11065), .IN4(n11066), 
        .QN(WX7135) );
  NAND2X0 U11136 ( .IN1(n11067), .IN2(n10384), .QN(n11066) );
  NAND2X0 U11137 ( .IN1(n11068), .IN2(n10387), .QN(n10384) );
  NAND2X0 U11138 ( .IN1(n11069), .IN2(n11070), .QN(n11068) );
  NAND2X0 U11139 ( .IN1(n16115), .IN2(n9119), .QN(n11070) );
  NAND2X0 U11140 ( .IN1(TM1), .IN2(n8365), .QN(n11069) );
  NAND3X0 U11141 ( .IN1(n11071), .IN2(n11072), .IN3(n11073), .QN(n11067) );
  NAND2X0 U11142 ( .IN1(n9331), .IN2(n10387), .QN(n11073) );
  NAND2X0 U11143 ( .IN1(n11074), .IN2(n11075), .QN(n10387) );
  NAND2X0 U11144 ( .IN1(n7687), .IN2(n11076), .QN(n11075) );
  INVX0 U11145 ( .INP(n11077), .ZN(n11074) );
  NOR2X0 U11146 ( .IN1(n11076), .IN2(n7687), .QN(n11077) );
  NOR2X0 U11147 ( .IN1(n11078), .IN2(n11079), .QN(n11076) );
  NOR2X0 U11148 ( .IN1(WX8621), .IN2(n7688), .QN(n11079) );
  INVX0 U11149 ( .INP(n11080), .ZN(n11078) );
  NAND2X0 U11150 ( .IN1(n7688), .IN2(WX8621), .QN(n11080) );
  NAND2X0 U11151 ( .IN1(n9083), .IN2(n8365), .QN(n11072) );
  NAND2X0 U11152 ( .IN1(n16115), .IN2(n9078), .QN(n11071) );
  NAND2X0 U11153 ( .IN1(n11081), .IN2(n11082), .QN(n11065) );
  NAND2X0 U11154 ( .IN1(n11083), .IN2(n11084), .QN(n11081) );
  NAND2X0 U11155 ( .IN1(n9091), .IN2(n11085), .QN(n11084) );
  NAND2X0 U11156 ( .IN1(n9092), .IN2(n8423), .QN(n11083) );
  NAND2X0 U11157 ( .IN1(n1226), .IN2(n9276), .QN(n11064) );
  NOR2X0 U11158 ( .IN1(n9224), .IN2(n8903), .QN(n1226) );
  NAND2X0 U11159 ( .IN1(n9309), .IN2(CRC_OUT_4_18), .QN(n11063) );
  NAND4X0 U11160 ( .IN1(n11086), .IN2(n11087), .IN3(n11088), .IN4(n11089), 
        .QN(WX7133) );
  NAND2X0 U11161 ( .IN1(n11090), .IN2(n10422), .QN(n11089) );
  NAND2X0 U11162 ( .IN1(n11091), .IN2(n10425), .QN(n10422) );
  NAND2X0 U11163 ( .IN1(n11092), .IN2(n11093), .QN(n11091) );
  NAND2X0 U11164 ( .IN1(n16114), .IN2(n9119), .QN(n11093) );
  NAND2X0 U11165 ( .IN1(TM1), .IN2(n8366), .QN(n11092) );
  NAND3X0 U11166 ( .IN1(n11094), .IN2(n11095), .IN3(n11096), .QN(n11090) );
  NAND2X0 U11167 ( .IN1(n9331), .IN2(n10425), .QN(n11096) );
  NAND2X0 U11168 ( .IN1(n11097), .IN2(n11098), .QN(n10425) );
  NAND2X0 U11169 ( .IN1(n7689), .IN2(n11099), .QN(n11098) );
  INVX0 U11170 ( .INP(n11100), .ZN(n11097) );
  NOR2X0 U11171 ( .IN1(n11099), .IN2(n7689), .QN(n11100) );
  NOR2X0 U11172 ( .IN1(n11101), .IN2(n11102), .QN(n11099) );
  NOR2X0 U11173 ( .IN1(WX8619), .IN2(n7690), .QN(n11102) );
  INVX0 U11174 ( .INP(n11103), .ZN(n11101) );
  NAND2X0 U11175 ( .IN1(n7690), .IN2(WX8619), .QN(n11103) );
  NAND2X0 U11176 ( .IN1(n9082), .IN2(n8366), .QN(n11095) );
  NAND2X0 U11177 ( .IN1(n16114), .IN2(n9077), .QN(n11094) );
  NAND2X0 U11178 ( .IN1(n11104), .IN2(n11105), .QN(n11088) );
  NAND2X0 U11179 ( .IN1(n11106), .IN2(n11107), .QN(n11104) );
  NAND2X0 U11180 ( .IN1(n9091), .IN2(n11108), .QN(n11107) );
  NAND2X0 U11181 ( .IN1(n9092), .IN2(n8424), .QN(n11106) );
  NAND2X0 U11182 ( .IN1(n1225), .IN2(n9276), .QN(n11087) );
  NOR2X0 U11183 ( .IN1(n9224), .IN2(n8904), .QN(n1225) );
  NAND2X0 U11184 ( .IN1(n9308), .IN2(CRC_OUT_4_19), .QN(n11086) );
  NAND4X0 U11185 ( .IN1(n11109), .IN2(n11110), .IN3(n11111), .IN4(n11112), 
        .QN(WX7131) );
  NAND2X0 U11186 ( .IN1(n11113), .IN2(n10442), .QN(n11112) );
  NAND2X0 U11187 ( .IN1(n11114), .IN2(n10445), .QN(n10442) );
  NAND2X0 U11188 ( .IN1(n11115), .IN2(n11116), .QN(n11114) );
  NAND2X0 U11189 ( .IN1(n16113), .IN2(n9119), .QN(n11116) );
  NAND2X0 U11190 ( .IN1(TM1), .IN2(n8367), .QN(n11115) );
  NAND3X0 U11191 ( .IN1(n11117), .IN2(n11118), .IN3(n11119), .QN(n11113) );
  NAND2X0 U11192 ( .IN1(n9331), .IN2(n10445), .QN(n11119) );
  NAND2X0 U11193 ( .IN1(n11120), .IN2(n11121), .QN(n10445) );
  NAND2X0 U11194 ( .IN1(n7691), .IN2(n11122), .QN(n11121) );
  INVX0 U11195 ( .INP(n11123), .ZN(n11120) );
  NOR2X0 U11196 ( .IN1(n11122), .IN2(n7691), .QN(n11123) );
  NOR2X0 U11197 ( .IN1(n11124), .IN2(n11125), .QN(n11122) );
  NOR2X0 U11198 ( .IN1(WX8617), .IN2(n7692), .QN(n11125) );
  INVX0 U11199 ( .INP(n11126), .ZN(n11124) );
  NAND2X0 U11200 ( .IN1(n7692), .IN2(WX8617), .QN(n11126) );
  NAND2X0 U11201 ( .IN1(n9081), .IN2(n8367), .QN(n11118) );
  NAND2X0 U11202 ( .IN1(n16113), .IN2(n9791), .QN(n11117) );
  NAND2X0 U11203 ( .IN1(n11127), .IN2(n11128), .QN(n11111) );
  NAND2X0 U11204 ( .IN1(n11129), .IN2(n11130), .QN(n11127) );
  NAND2X0 U11205 ( .IN1(n9092), .IN2(n11131), .QN(n11130) );
  NAND2X0 U11206 ( .IN1(n9091), .IN2(n8425), .QN(n11129) );
  NAND2X0 U11207 ( .IN1(n1224), .IN2(n9276), .QN(n11110) );
  NOR2X0 U11208 ( .IN1(n9224), .IN2(n8905), .QN(n1224) );
  NAND2X0 U11209 ( .IN1(n9309), .IN2(CRC_OUT_4_20), .QN(n11109) );
  NAND4X0 U11210 ( .IN1(n11132), .IN2(n11133), .IN3(n11134), .IN4(n11135), 
        .QN(WX7129) );
  NAND2X0 U11211 ( .IN1(n11136), .IN2(n10465), .QN(n11135) );
  NAND2X0 U11212 ( .IN1(n11137), .IN2(n10468), .QN(n10465) );
  NAND2X0 U11213 ( .IN1(n11138), .IN2(n11139), .QN(n11137) );
  NAND2X0 U11214 ( .IN1(n16112), .IN2(n9119), .QN(n11139) );
  NAND2X0 U11215 ( .IN1(TM1), .IN2(n8368), .QN(n11138) );
  NAND3X0 U11216 ( .IN1(n11140), .IN2(n11141), .IN3(n11142), .QN(n11136) );
  NAND2X0 U11217 ( .IN1(n9331), .IN2(n10468), .QN(n11142) );
  NAND2X0 U11218 ( .IN1(n11143), .IN2(n11144), .QN(n10468) );
  NAND2X0 U11219 ( .IN1(n7693), .IN2(n11145), .QN(n11144) );
  INVX0 U11220 ( .INP(n11146), .ZN(n11143) );
  NOR2X0 U11221 ( .IN1(n11145), .IN2(n7693), .QN(n11146) );
  NOR2X0 U11222 ( .IN1(n11147), .IN2(n11148), .QN(n11145) );
  NOR2X0 U11223 ( .IN1(WX8615), .IN2(n7694), .QN(n11148) );
  INVX0 U11224 ( .INP(n11149), .ZN(n11147) );
  NAND2X0 U11225 ( .IN1(n7694), .IN2(WX8615), .QN(n11149) );
  NAND2X0 U11226 ( .IN1(n9790), .IN2(n8368), .QN(n11141) );
  NAND2X0 U11227 ( .IN1(n16112), .IN2(n9079), .QN(n11140) );
  NAND2X0 U11228 ( .IN1(n11150), .IN2(n9111), .QN(n11134) );
  NAND2X0 U11229 ( .IN1(n1223), .IN2(n9276), .QN(n11133) );
  NOR2X0 U11230 ( .IN1(n9224), .IN2(n8906), .QN(n1223) );
  NAND2X0 U11231 ( .IN1(n9309), .IN2(CRC_OUT_4_21), .QN(n11132) );
  NAND4X0 U11232 ( .IN1(n11151), .IN2(n11152), .IN3(n11153), .IN4(n11154), 
        .QN(WX7127) );
  NAND2X0 U11233 ( .IN1(n11155), .IN2(n10488), .QN(n11154) );
  NAND2X0 U11234 ( .IN1(n11156), .IN2(n10491), .QN(n10488) );
  NAND2X0 U11235 ( .IN1(n11157), .IN2(n11158), .QN(n11156) );
  NAND2X0 U11236 ( .IN1(n16111), .IN2(n9119), .QN(n11158) );
  NAND2X0 U11237 ( .IN1(TM1), .IN2(n8369), .QN(n11157) );
  NAND3X0 U11238 ( .IN1(n11159), .IN2(n11160), .IN3(n11161), .QN(n11155) );
  NAND2X0 U11239 ( .IN1(n9331), .IN2(n10491), .QN(n11161) );
  NAND2X0 U11240 ( .IN1(n11162), .IN2(n11163), .QN(n10491) );
  NAND2X0 U11241 ( .IN1(n7695), .IN2(n11164), .QN(n11163) );
  INVX0 U11242 ( .INP(n11165), .ZN(n11162) );
  NOR2X0 U11243 ( .IN1(n11164), .IN2(n7695), .QN(n11165) );
  NOR2X0 U11244 ( .IN1(n11166), .IN2(n11167), .QN(n11164) );
  NOR2X0 U11245 ( .IN1(WX8613), .IN2(n7696), .QN(n11167) );
  INVX0 U11246 ( .INP(n11168), .ZN(n11166) );
  NAND2X0 U11247 ( .IN1(n7696), .IN2(WX8613), .QN(n11168) );
  NAND2X0 U11248 ( .IN1(n9083), .IN2(n8369), .QN(n11160) );
  NAND2X0 U11249 ( .IN1(n16111), .IN2(n9078), .QN(n11159) );
  NAND2X0 U11250 ( .IN1(n11169), .IN2(n11170), .QN(n11153) );
  NAND2X0 U11251 ( .IN1(n11171), .IN2(n11172), .QN(n11169) );
  NAND2X0 U11252 ( .IN1(n9091), .IN2(n11173), .QN(n11172) );
  NAND2X0 U11253 ( .IN1(n9092), .IN2(n8427), .QN(n11171) );
  NAND2X0 U11254 ( .IN1(n1222), .IN2(n9277), .QN(n11152) );
  NOR2X0 U11255 ( .IN1(n9224), .IN2(n8907), .QN(n1222) );
  NAND2X0 U11256 ( .IN1(n9309), .IN2(CRC_OUT_4_22), .QN(n11151) );
  NAND4X0 U11257 ( .IN1(n11174), .IN2(n11175), .IN3(n11176), .IN4(n11177), 
        .QN(WX7125) );
  NAND2X0 U11258 ( .IN1(n11178), .IN2(n10511), .QN(n11177) );
  NAND2X0 U11259 ( .IN1(n11179), .IN2(n10514), .QN(n10511) );
  NAND2X0 U11260 ( .IN1(n11180), .IN2(n11181), .QN(n11179) );
  NAND2X0 U11261 ( .IN1(n16110), .IN2(n9119), .QN(n11181) );
  NAND2X0 U11262 ( .IN1(TM1), .IN2(n8370), .QN(n11180) );
  NAND3X0 U11263 ( .IN1(n11182), .IN2(n11183), .IN3(n11184), .QN(n11178) );
  NAND2X0 U11264 ( .IN1(n9331), .IN2(n10514), .QN(n11184) );
  NAND2X0 U11265 ( .IN1(n11185), .IN2(n11186), .QN(n10514) );
  NAND2X0 U11266 ( .IN1(n7697), .IN2(n11187), .QN(n11186) );
  INVX0 U11267 ( .INP(n11188), .ZN(n11185) );
  NOR2X0 U11268 ( .IN1(n11187), .IN2(n7697), .QN(n11188) );
  NOR2X0 U11269 ( .IN1(n11189), .IN2(n11190), .QN(n11187) );
  NOR2X0 U11270 ( .IN1(WX8611), .IN2(n7698), .QN(n11190) );
  INVX0 U11271 ( .INP(n11191), .ZN(n11189) );
  NAND2X0 U11272 ( .IN1(n7698), .IN2(WX8611), .QN(n11191) );
  NAND2X0 U11273 ( .IN1(n9082), .IN2(n8370), .QN(n11183) );
  NAND2X0 U11274 ( .IN1(n16110), .IN2(n9077), .QN(n11182) );
  NAND2X0 U11275 ( .IN1(n11192), .IN2(n9110), .QN(n11176) );
  NAND2X0 U11276 ( .IN1(n1221), .IN2(n9277), .QN(n11175) );
  NOR2X0 U11277 ( .IN1(n9224), .IN2(n8908), .QN(n1221) );
  NAND2X0 U11278 ( .IN1(n9309), .IN2(CRC_OUT_4_23), .QN(n11174) );
  NAND4X0 U11279 ( .IN1(n11193), .IN2(n11194), .IN3(n11195), .IN4(n11196), 
        .QN(WX7123) );
  NAND2X0 U11280 ( .IN1(n11197), .IN2(n10534), .QN(n11196) );
  NAND2X0 U11281 ( .IN1(n11198), .IN2(n10537), .QN(n10534) );
  NAND2X0 U11282 ( .IN1(n11199), .IN2(n11200), .QN(n11198) );
  NAND2X0 U11283 ( .IN1(n16109), .IN2(n9119), .QN(n11200) );
  NAND2X0 U11284 ( .IN1(TM1), .IN2(n8371), .QN(n11199) );
  NAND3X0 U11285 ( .IN1(n11201), .IN2(n11202), .IN3(n11203), .QN(n11197) );
  NAND2X0 U11286 ( .IN1(n9332), .IN2(n10537), .QN(n11203) );
  NAND2X0 U11287 ( .IN1(n11204), .IN2(n11205), .QN(n10537) );
  NAND2X0 U11288 ( .IN1(n7699), .IN2(n11206), .QN(n11205) );
  INVX0 U11289 ( .INP(n11207), .ZN(n11204) );
  NOR2X0 U11290 ( .IN1(n11206), .IN2(n7699), .QN(n11207) );
  NOR2X0 U11291 ( .IN1(n11208), .IN2(n11209), .QN(n11206) );
  NOR2X0 U11292 ( .IN1(WX8609), .IN2(n7700), .QN(n11209) );
  INVX0 U11293 ( .INP(n11210), .ZN(n11208) );
  NAND2X0 U11294 ( .IN1(n7700), .IN2(WX8609), .QN(n11210) );
  NAND2X0 U11295 ( .IN1(n9081), .IN2(n8371), .QN(n11202) );
  NAND2X0 U11296 ( .IN1(n16109), .IN2(n9791), .QN(n11201) );
  NAND2X0 U11297 ( .IN1(n11211), .IN2(n11212), .QN(n11195) );
  NAND2X0 U11298 ( .IN1(n11213), .IN2(n11214), .QN(n11211) );
  NAND2X0 U11299 ( .IN1(n9091), .IN2(n11215), .QN(n11214) );
  NAND2X0 U11300 ( .IN1(n9091), .IN2(n8429), .QN(n11213) );
  NAND2X0 U11301 ( .IN1(n1220), .IN2(n9277), .QN(n11194) );
  NOR2X0 U11302 ( .IN1(n9224), .IN2(n8909), .QN(n1220) );
  NAND2X0 U11303 ( .IN1(n9309), .IN2(CRC_OUT_4_24), .QN(n11193) );
  NAND4X0 U11304 ( .IN1(n11216), .IN2(n11217), .IN3(n11218), .IN4(n11219), 
        .QN(WX7121) );
  NAND2X0 U11305 ( .IN1(n11220), .IN2(n10557), .QN(n11219) );
  NAND2X0 U11306 ( .IN1(n11221), .IN2(n10560), .QN(n10557) );
  NAND2X0 U11307 ( .IN1(n11222), .IN2(n11223), .QN(n11221) );
  NAND2X0 U11308 ( .IN1(n16108), .IN2(n9119), .QN(n11223) );
  NAND2X0 U11309 ( .IN1(TM1), .IN2(n8372), .QN(n11222) );
  NAND3X0 U11310 ( .IN1(n11224), .IN2(n11225), .IN3(n11226), .QN(n11220) );
  NAND2X0 U11311 ( .IN1(n9332), .IN2(n10560), .QN(n11226) );
  NAND2X0 U11312 ( .IN1(n11227), .IN2(n11228), .QN(n10560) );
  NAND2X0 U11313 ( .IN1(n7701), .IN2(n11229), .QN(n11228) );
  INVX0 U11314 ( .INP(n11230), .ZN(n11227) );
  NOR2X0 U11315 ( .IN1(n11229), .IN2(n7701), .QN(n11230) );
  NOR2X0 U11316 ( .IN1(n11231), .IN2(n11232), .QN(n11229) );
  NOR2X0 U11317 ( .IN1(WX8607), .IN2(n7702), .QN(n11232) );
  INVX0 U11318 ( .INP(n11233), .ZN(n11231) );
  NAND2X0 U11319 ( .IN1(n7702), .IN2(WX8607), .QN(n11233) );
  NAND2X0 U11320 ( .IN1(n9790), .IN2(n8372), .QN(n11225) );
  NAND2X0 U11321 ( .IN1(n16108), .IN2(n9079), .QN(n11224) );
  NAND2X0 U11322 ( .IN1(n11234), .IN2(n9110), .QN(n11218) );
  NAND2X0 U11323 ( .IN1(n1219), .IN2(n9277), .QN(n11217) );
  NOR2X0 U11324 ( .IN1(n9224), .IN2(n8910), .QN(n1219) );
  NAND2X0 U11325 ( .IN1(n9309), .IN2(CRC_OUT_4_25), .QN(n11216) );
  NAND4X0 U11326 ( .IN1(n11235), .IN2(n11236), .IN3(n11237), .IN4(n11238), 
        .QN(WX7119) );
  NAND2X0 U11327 ( .IN1(n11239), .IN2(n11240), .QN(n11238) );
  NAND2X0 U11328 ( .IN1(n11241), .IN2(n11242), .QN(n11239) );
  NAND2X0 U11329 ( .IN1(n9092), .IN2(n11243), .QN(n11242) );
  NAND2X0 U11330 ( .IN1(n9091), .IN2(n8431), .QN(n11241) );
  NAND2X0 U11331 ( .IN1(n10579), .IN2(n2153), .QN(n11237) );
  NOR2X0 U11332 ( .IN1(n11244), .IN2(n11245), .QN(n10579) );
  INVX0 U11333 ( .INP(n11246), .ZN(n11245) );
  NAND2X0 U11334 ( .IN1(n11247), .IN2(n11248), .QN(n11246) );
  NOR2X0 U11335 ( .IN1(n11248), .IN2(n11247), .QN(n11244) );
  NAND2X0 U11336 ( .IN1(n11249), .IN2(n11250), .QN(n11247) );
  NAND2X0 U11337 ( .IN1(n11251), .IN2(WX8541), .QN(n11250) );
  NAND2X0 U11338 ( .IN1(n11252), .IN2(n11253), .QN(n11251) );
  NAND3X0 U11339 ( .IN1(n11252), .IN2(n11253), .IN3(n7704), .QN(n11249) );
  NAND2X0 U11340 ( .IN1(test_so74), .IN2(WX8477), .QN(n11253) );
  NAND2X0 U11341 ( .IN1(n7703), .IN2(n8798), .QN(n11252) );
  NOR2X0 U11342 ( .IN1(n11254), .IN2(n11255), .QN(n11248) );
  INVX0 U11343 ( .INP(n11256), .ZN(n11255) );
  NAND2X0 U11344 ( .IN1(n16107), .IN2(n9119), .QN(n11256) );
  NOR2X0 U11345 ( .IN1(n9117), .IN2(n16107), .QN(n11254) );
  NAND2X0 U11346 ( .IN1(n1218), .IN2(n9277), .QN(n11236) );
  NOR2X0 U11347 ( .IN1(n9224), .IN2(n8911), .QN(n1218) );
  NAND2X0 U11348 ( .IN1(n9310), .IN2(CRC_OUT_4_26), .QN(n11235) );
  NAND4X0 U11349 ( .IN1(n11257), .IN2(n11258), .IN3(n11259), .IN4(n11260), 
        .QN(WX7117) );
  NAND2X0 U11350 ( .IN1(n11261), .IN2(n10599), .QN(n11260) );
  NAND2X0 U11351 ( .IN1(n11262), .IN2(n10602), .QN(n10599) );
  NAND2X0 U11352 ( .IN1(n11263), .IN2(n11264), .QN(n11262) );
  NAND2X0 U11353 ( .IN1(n16106), .IN2(n9119), .QN(n11264) );
  NAND2X0 U11354 ( .IN1(TM1), .IN2(n8374), .QN(n11263) );
  NAND3X0 U11355 ( .IN1(n11265), .IN2(n11266), .IN3(n11267), .QN(n11261) );
  NAND2X0 U11356 ( .IN1(n9332), .IN2(n10602), .QN(n11267) );
  NAND2X0 U11357 ( .IN1(n11268), .IN2(n11269), .QN(n10602) );
  NAND2X0 U11358 ( .IN1(n7705), .IN2(n11270), .QN(n11269) );
  INVX0 U11359 ( .INP(n11271), .ZN(n11268) );
  NOR2X0 U11360 ( .IN1(n11270), .IN2(n7705), .QN(n11271) );
  NOR2X0 U11361 ( .IN1(n11272), .IN2(n11273), .QN(n11270) );
  NOR2X0 U11362 ( .IN1(WX8603), .IN2(n7706), .QN(n11273) );
  INVX0 U11363 ( .INP(n11274), .ZN(n11272) );
  NAND2X0 U11364 ( .IN1(n7706), .IN2(WX8603), .QN(n11274) );
  NAND2X0 U11365 ( .IN1(n9083), .IN2(n8374), .QN(n11266) );
  NAND2X0 U11366 ( .IN1(n16106), .IN2(n9078), .QN(n11265) );
  NAND2X0 U11367 ( .IN1(n11275), .IN2(n11276), .QN(n11259) );
  NAND2X0 U11368 ( .IN1(n11277), .IN2(n11278), .QN(n11275) );
  NAND2X0 U11369 ( .IN1(n9092), .IN2(n11279), .QN(n11278) );
  NAND2X0 U11370 ( .IN1(n8215), .IN2(n9110), .QN(n11277) );
  NAND2X0 U11371 ( .IN1(n1217), .IN2(n9277), .QN(n11258) );
  NOR2X0 U11372 ( .IN1(n9224), .IN2(n8912), .QN(n1217) );
  NAND2X0 U11373 ( .IN1(n9310), .IN2(CRC_OUT_4_27), .QN(n11257) );
  NAND4X0 U11374 ( .IN1(n11280), .IN2(n11281), .IN3(n11282), .IN4(n11283), 
        .QN(WX7115) );
  NAND2X0 U11375 ( .IN1(n11284), .IN2(n11285), .QN(n11283) );
  NAND2X0 U11376 ( .IN1(n11286), .IN2(n11287), .QN(n11284) );
  NAND2X0 U11377 ( .IN1(n9092), .IN2(n11288), .QN(n11287) );
  NAND2X0 U11378 ( .IN1(n9092), .IN2(n8434), .QN(n11286) );
  NAND2X0 U11379 ( .IN1(n10621), .IN2(n2153), .QN(n11282) );
  NOR2X0 U11380 ( .IN1(n11289), .IN2(n11290), .QN(n10621) );
  INVX0 U11381 ( .INP(n11291), .ZN(n11290) );
  NAND2X0 U11382 ( .IN1(n11292), .IN2(n11293), .QN(n11291) );
  NOR2X0 U11383 ( .IN1(n11293), .IN2(n11292), .QN(n11289) );
  NAND2X0 U11384 ( .IN1(n11294), .IN2(n11295), .QN(n11292) );
  NAND2X0 U11385 ( .IN1(n8188), .IN2(n11296), .QN(n11295) );
  INVX0 U11386 ( .INP(n11297), .ZN(n11296) );
  NAND2X0 U11387 ( .IN1(n11297), .IN2(WX8601), .QN(n11294) );
  NAND2X0 U11388 ( .IN1(n11298), .IN2(n11299), .QN(n11297) );
  INVX0 U11389 ( .INP(n11300), .ZN(n11299) );
  NOR2X0 U11390 ( .IN1(n8807), .IN2(n16105), .QN(n11300) );
  NAND2X0 U11391 ( .IN1(n16105), .IN2(n8807), .QN(n11298) );
  NOR2X0 U11392 ( .IN1(n11301), .IN2(n11302), .QN(n11293) );
  INVX0 U11393 ( .INP(n11303), .ZN(n11302) );
  NAND2X0 U11394 ( .IN1(n7707), .IN2(n9119), .QN(n11303) );
  NOR2X0 U11395 ( .IN1(n9116), .IN2(n7707), .QN(n11301) );
  NAND2X0 U11396 ( .IN1(n1216), .IN2(n9277), .QN(n11281) );
  NOR2X0 U11397 ( .IN1(n9225), .IN2(n8913), .QN(n1216) );
  NAND2X0 U11398 ( .IN1(n9310), .IN2(CRC_OUT_4_28), .QN(n11280) );
  NAND4X0 U11399 ( .IN1(n11304), .IN2(n11305), .IN3(n11306), .IN4(n11307), 
        .QN(WX7113) );
  NAND2X0 U11400 ( .IN1(n11308), .IN2(n10641), .QN(n11307) );
  NAND2X0 U11401 ( .IN1(n11309), .IN2(n10644), .QN(n10641) );
  NAND2X0 U11402 ( .IN1(n11310), .IN2(n11311), .QN(n11309) );
  NAND2X0 U11403 ( .IN1(n16104), .IN2(n9119), .QN(n11311) );
  NAND2X0 U11404 ( .IN1(TM1), .IN2(n8376), .QN(n11310) );
  NAND3X0 U11405 ( .IN1(n11312), .IN2(n11313), .IN3(n11314), .QN(n11308) );
  NAND2X0 U11406 ( .IN1(n9332), .IN2(n10644), .QN(n11314) );
  NAND2X0 U11407 ( .IN1(n11315), .IN2(n11316), .QN(n10644) );
  NAND2X0 U11408 ( .IN1(n7708), .IN2(n11317), .QN(n11316) );
  INVX0 U11409 ( .INP(n11318), .ZN(n11315) );
  NOR2X0 U11410 ( .IN1(n11317), .IN2(n7708), .QN(n11318) );
  NOR2X0 U11411 ( .IN1(n11319), .IN2(n11320), .QN(n11317) );
  NOR2X0 U11412 ( .IN1(WX8599), .IN2(n7709), .QN(n11320) );
  INVX0 U11413 ( .INP(n11321), .ZN(n11319) );
  NAND2X0 U11414 ( .IN1(n7709), .IN2(WX8599), .QN(n11321) );
  NAND2X0 U11415 ( .IN1(n9082), .IN2(n8376), .QN(n11313) );
  NAND2X0 U11416 ( .IN1(n16104), .IN2(n9077), .QN(n11312) );
  NAND2X0 U11417 ( .IN1(n11322), .IN2(n11323), .QN(n11306) );
  NAND2X0 U11418 ( .IN1(n11324), .IN2(n11325), .QN(n11322) );
  NAND2X0 U11419 ( .IN1(n9092), .IN2(n11326), .QN(n11325) );
  NAND2X0 U11420 ( .IN1(n9092), .IN2(n8435), .QN(n11324) );
  NAND2X0 U11421 ( .IN1(n1215), .IN2(n9277), .QN(n11305) );
  NOR2X0 U11422 ( .IN1(n9065), .IN2(n9163), .QN(n1215) );
  NAND2X0 U11423 ( .IN1(test_so66), .IN2(n9314), .QN(n11304) );
  NAND4X0 U11424 ( .IN1(n11327), .IN2(n11328), .IN3(n11329), .IN4(n11330), 
        .QN(WX7111) );
  NAND2X0 U11425 ( .IN1(n11331), .IN2(n11332), .QN(n11330) );
  NAND2X0 U11426 ( .IN1(n11333), .IN2(n11334), .QN(n11331) );
  NAND2X0 U11427 ( .IN1(n9092), .IN2(n11335), .QN(n11334) );
  NAND2X0 U11428 ( .IN1(n9092), .IN2(n8436), .QN(n11333) );
  NAND2X0 U11429 ( .IN1(n10663), .IN2(n2153), .QN(n11329) );
  NOR2X0 U11430 ( .IN1(n11336), .IN2(n11337), .QN(n10663) );
  INVX0 U11431 ( .INP(n11338), .ZN(n11337) );
  NAND2X0 U11432 ( .IN1(n11339), .IN2(n11340), .QN(n11338) );
  NOR2X0 U11433 ( .IN1(n11340), .IN2(n11339), .QN(n11336) );
  NAND2X0 U11434 ( .IN1(n11341), .IN2(n11342), .QN(n11339) );
  NAND2X0 U11435 ( .IN1(n8186), .IN2(n11343), .QN(n11342) );
  INVX0 U11436 ( .INP(n11344), .ZN(n11343) );
  NAND2X0 U11437 ( .IN1(n11344), .IN2(WX8597), .QN(n11341) );
  NAND2X0 U11438 ( .IN1(n11345), .IN2(n11346), .QN(n11344) );
  INVX0 U11439 ( .INP(n11347), .ZN(n11346) );
  NOR2X0 U11440 ( .IN1(n8808), .IN2(n16103), .QN(n11347) );
  NAND2X0 U11441 ( .IN1(n16103), .IN2(n8808), .QN(n11345) );
  NOR2X0 U11442 ( .IN1(n11348), .IN2(n11349), .QN(n11340) );
  INVX0 U11443 ( .INP(n11350), .ZN(n11349) );
  NAND2X0 U11444 ( .IN1(n7710), .IN2(n9118), .QN(n11350) );
  NOR2X0 U11445 ( .IN1(n9117), .IN2(n7710), .QN(n11348) );
  NAND2X0 U11446 ( .IN1(n1214), .IN2(n9277), .QN(n11328) );
  NOR2X0 U11447 ( .IN1(n9225), .IN2(n8914), .QN(n1214) );
  NAND2X0 U11448 ( .IN1(n9310), .IN2(CRC_OUT_4_30), .QN(n11327) );
  NAND4X0 U11449 ( .IN1(n11351), .IN2(n11352), .IN3(n11353), .IN4(n11354), 
        .QN(WX7109) );
  NAND2X0 U11450 ( .IN1(n11355), .IN2(n10669), .QN(n11354) );
  NAND2X0 U11451 ( .IN1(n11356), .IN2(n10672), .QN(n10669) );
  NAND2X0 U11452 ( .IN1(n11357), .IN2(n11358), .QN(n11356) );
  NAND2X0 U11453 ( .IN1(n16102), .IN2(n9118), .QN(n11358) );
  NAND2X0 U11454 ( .IN1(TM1), .IN2(n8378), .QN(n11357) );
  NAND3X0 U11455 ( .IN1(n11359), .IN2(n11360), .IN3(n11361), .QN(n11355) );
  NAND2X0 U11456 ( .IN1(n9332), .IN2(n10672), .QN(n11361) );
  NAND2X0 U11457 ( .IN1(n11362), .IN2(n11363), .QN(n10672) );
  NAND2X0 U11458 ( .IN1(n7615), .IN2(n11364), .QN(n11363) );
  INVX0 U11459 ( .INP(n11365), .ZN(n11362) );
  NOR2X0 U11460 ( .IN1(n11364), .IN2(n7615), .QN(n11365) );
  NOR2X0 U11461 ( .IN1(n11366), .IN2(n11367), .QN(n11364) );
  NOR2X0 U11462 ( .IN1(WX8595), .IN2(n7616), .QN(n11367) );
  INVX0 U11463 ( .INP(n11368), .ZN(n11366) );
  NAND2X0 U11464 ( .IN1(n7616), .IN2(WX8595), .QN(n11368) );
  NAND2X0 U11465 ( .IN1(n9081), .IN2(n8378), .QN(n11360) );
  NAND2X0 U11466 ( .IN1(n16102), .IN2(n9791), .QN(n11359) );
  NAND2X0 U11467 ( .IN1(n11369), .IN2(n11370), .QN(n11353) );
  NAND2X0 U11468 ( .IN1(n11371), .IN2(n11372), .QN(n11369) );
  NAND2X0 U11469 ( .IN1(n9092), .IN2(n11373), .QN(n11372) );
  NAND2X0 U11470 ( .IN1(n9092), .IN2(n8437), .QN(n11371) );
  NAND2X0 U11471 ( .IN1(n9309), .IN2(CRC_OUT_4_31), .QN(n11352) );
  NAND2X0 U11472 ( .IN1(n2245), .IN2(WX6950), .QN(n11351) );
  NAND4X0 U11473 ( .IN1(n11374), .IN2(n11375), .IN3(n11376), .IN4(n11377), 
        .QN(WX706) );
  NAND3X0 U11474 ( .IN1(n11378), .IN2(n11379), .IN3(n9321), .QN(n11377) );
  NAND2X0 U11475 ( .IN1(n9093), .IN2(n11380), .QN(n11376) );
  NAND2X0 U11476 ( .IN1(WX544), .IN2(n9277), .QN(n11375) );
  NAND2X0 U11477 ( .IN1(n9310), .IN2(CRC_OUT_9_0), .QN(n11374) );
  NAND4X0 U11478 ( .IN1(n11381), .IN2(n11382), .IN3(n11383), .IN4(n11384), 
        .QN(WX704) );
  NAND2X0 U11479 ( .IN1(n9332), .IN2(n11385), .QN(n11384) );
  NAND2X0 U11480 ( .IN1(n9092), .IN2(n11386), .QN(n11383) );
  NAND2X0 U11481 ( .IN1(WX542), .IN2(n9277), .QN(n11382) );
  NAND2X0 U11482 ( .IN1(test_so9), .IN2(n9314), .QN(n11381) );
  NAND4X0 U11483 ( .IN1(n11387), .IN2(n11388), .IN3(n11389), .IN4(n11390), 
        .QN(WX702) );
  NAND2X0 U11484 ( .IN1(n9332), .IN2(n11391), .QN(n11390) );
  NAND2X0 U11485 ( .IN1(n11392), .IN2(n9109), .QN(n11389) );
  INVX0 U11486 ( .INP(n11393), .ZN(n11392) );
  NAND2X0 U11487 ( .IN1(WX540), .IN2(n9277), .QN(n11388) );
  NAND2X0 U11488 ( .IN1(n9310), .IN2(CRC_OUT_9_2), .QN(n11387) );
  NOR2X0 U11489 ( .IN1(n9225), .IN2(WX6950), .QN(WX7011) );
  NAND4X0 U11490 ( .IN1(n11394), .IN2(n11395), .IN3(n11396), .IN4(n11397), 
        .QN(WX700) );
  NAND2X0 U11491 ( .IN1(n9332), .IN2(n11398), .QN(n11397) );
  NAND2X0 U11492 ( .IN1(n9092), .IN2(n11399), .QN(n11396) );
  NAND2X0 U11493 ( .IN1(WX538), .IN2(n9277), .QN(n11395) );
  NAND2X0 U11494 ( .IN1(n9309), .IN2(CRC_OUT_9_3), .QN(n11394) );
  NAND4X0 U11495 ( .IN1(n11400), .IN2(n11401), .IN3(n11402), .IN4(n11403), 
        .QN(WX698) );
  NAND3X0 U11496 ( .IN1(n11404), .IN2(n11405), .IN3(n9321), .QN(n11403) );
  NAND2X0 U11497 ( .IN1(n9092), .IN2(n11406), .QN(n11402) );
  NAND2X0 U11498 ( .IN1(WX536), .IN2(n9277), .QN(n11401) );
  NAND2X0 U11499 ( .IN1(n9310), .IN2(CRC_OUT_9_4), .QN(n11400) );
  NAND4X0 U11500 ( .IN1(n11407), .IN2(n11408), .IN3(n11409), .IN4(n11410), 
        .QN(WX696) );
  NAND2X0 U11501 ( .IN1(n9332), .IN2(n11411), .QN(n11410) );
  NAND2X0 U11502 ( .IN1(n9093), .IN2(n11412), .QN(n11409) );
  NAND2X0 U11503 ( .IN1(WX534), .IN2(n9277), .QN(n11408) );
  NAND2X0 U11504 ( .IN1(n9311), .IN2(CRC_OUT_9_5), .QN(n11407) );
  NAND4X0 U11505 ( .IN1(n11413), .IN2(n11414), .IN3(n11415), .IN4(n11416), 
        .QN(WX694) );
  NAND2X0 U11506 ( .IN1(n9332), .IN2(n11417), .QN(n11416) );
  NAND2X0 U11507 ( .IN1(n11418), .IN2(n9111), .QN(n11415) );
  INVX0 U11508 ( .INP(n11419), .ZN(n11418) );
  NAND2X0 U11509 ( .IN1(WX532), .IN2(n9277), .QN(n11414) );
  NAND2X0 U11510 ( .IN1(n9310), .IN2(CRC_OUT_9_6), .QN(n11413) );
  NAND4X0 U11511 ( .IN1(n11420), .IN2(n11421), .IN3(n11422), .IN4(n11423), 
        .QN(WX692) );
  NAND2X0 U11512 ( .IN1(n9332), .IN2(n11424), .QN(n11423) );
  NAND2X0 U11513 ( .IN1(n9093), .IN2(n11425), .QN(n11422) );
  NAND2X0 U11514 ( .IN1(WX530), .IN2(n9277), .QN(n11421) );
  NAND2X0 U11515 ( .IN1(n9311), .IN2(CRC_OUT_9_7), .QN(n11420) );
  NAND4X0 U11516 ( .IN1(n11426), .IN2(n11427), .IN3(n11428), .IN4(n11429), 
        .QN(WX690) );
  NAND2X0 U11517 ( .IN1(n9332), .IN2(n11430), .QN(n11429) );
  NAND2X0 U11518 ( .IN1(n9093), .IN2(n11431), .QN(n11428) );
  NAND2X0 U11519 ( .IN1(WX528), .IN2(n9278), .QN(n11427) );
  NAND2X0 U11520 ( .IN1(n9309), .IN2(CRC_OUT_9_8), .QN(n11426) );
  NAND4X0 U11521 ( .IN1(n11432), .IN2(n11433), .IN3(n11434), .IN4(n11435), 
        .QN(WX688) );
  NAND2X0 U11522 ( .IN1(n9332), .IN2(n11436), .QN(n11435) );
  NAND2X0 U11523 ( .IN1(n9093), .IN2(n11437), .QN(n11434) );
  NAND2X0 U11524 ( .IN1(WX526), .IN2(n9278), .QN(n11433) );
  NAND2X0 U11525 ( .IN1(n9311), .IN2(CRC_OUT_9_9), .QN(n11432) );
  NAND4X0 U11526 ( .IN1(n11438), .IN2(n11439), .IN3(n11440), .IN4(n11441), 
        .QN(WX686) );
  NAND3X0 U11527 ( .IN1(n11442), .IN2(n11443), .IN3(n9321), .QN(n11441) );
  NAND2X0 U11528 ( .IN1(n11444), .IN2(n9110), .QN(n11440) );
  INVX0 U11529 ( .INP(n11445), .ZN(n11444) );
  NAND2X0 U11530 ( .IN1(WX524), .IN2(n9278), .QN(n11439) );
  NAND2X0 U11531 ( .IN1(n9311), .IN2(CRC_OUT_9_10), .QN(n11438) );
  NAND4X0 U11532 ( .IN1(n11446), .IN2(n11447), .IN3(n11448), .IN4(n11449), 
        .QN(WX684) );
  NAND2X0 U11533 ( .IN1(n9332), .IN2(n11450), .QN(n11449) );
  NAND2X0 U11534 ( .IN1(n9093), .IN2(n11451), .QN(n11448) );
  NAND2X0 U11535 ( .IN1(WX522), .IN2(n9278), .QN(n11447) );
  NAND2X0 U11536 ( .IN1(n9311), .IN2(CRC_OUT_9_11), .QN(n11446) );
  NAND4X0 U11537 ( .IN1(n11452), .IN2(n11453), .IN3(n11454), .IN4(n11455), 
        .QN(WX682) );
  NAND2X0 U11538 ( .IN1(n9331), .IN2(n11456), .QN(n11455) );
  NAND2X0 U11539 ( .IN1(n9093), .IN2(n11457), .QN(n11454) );
  NAND2X0 U11540 ( .IN1(WX520), .IN2(n9278), .QN(n11453) );
  NAND2X0 U11541 ( .IN1(n9310), .IN2(CRC_OUT_9_12), .QN(n11452) );
  NAND4X0 U11542 ( .IN1(n11458), .IN2(n11459), .IN3(n11460), .IN4(n11461), 
        .QN(WX680) );
  NAND2X0 U11543 ( .IN1(n9332), .IN2(n11462), .QN(n11461) );
  NAND2X0 U11544 ( .IN1(n9093), .IN2(n11463), .QN(n11460) );
  NAND2X0 U11545 ( .IN1(WX518), .IN2(n9278), .QN(n11459) );
  NAND2X0 U11546 ( .IN1(n9308), .IN2(CRC_OUT_9_13), .QN(n11458) );
  NAND4X0 U11547 ( .IN1(n11464), .IN2(n11465), .IN3(n11466), .IN4(n11467), 
        .QN(WX678) );
  NAND3X0 U11548 ( .IN1(n11468), .IN2(n11469), .IN3(n9321), .QN(n11467) );
  NAND2X0 U11549 ( .IN1(n9093), .IN2(n11470), .QN(n11466) );
  NAND2X0 U11550 ( .IN1(WX516), .IN2(n9278), .QN(n11465) );
  NAND2X0 U11551 ( .IN1(n9310), .IN2(CRC_OUT_9_14), .QN(n11464) );
  NAND4X0 U11552 ( .IN1(n11471), .IN2(n11472), .IN3(n11473), .IN4(n11474), 
        .QN(WX676) );
  NAND2X0 U11553 ( .IN1(n9332), .IN2(n11475), .QN(n11474) );
  NAND2X0 U11554 ( .IN1(n9093), .IN2(n11476), .QN(n11473) );
  NAND2X0 U11555 ( .IN1(WX514), .IN2(n9278), .QN(n11472) );
  NAND2X0 U11556 ( .IN1(n9312), .IN2(CRC_OUT_9_15), .QN(n11471) );
  NAND4X0 U11557 ( .IN1(n11477), .IN2(n11478), .IN3(n11479), .IN4(n11480), 
        .QN(WX674) );
  NAND2X0 U11558 ( .IN1(n11481), .IN2(n11482), .QN(n11480) );
  NAND3X0 U11559 ( .IN1(n11483), .IN2(n11484), .IN3(n11485), .QN(n11481) );
  NAND2X0 U11560 ( .IN1(n9332), .IN2(n11486), .QN(n11485) );
  NAND2X0 U11561 ( .IN1(n9790), .IN2(n8653), .QN(n11484) );
  NAND2X0 U11562 ( .IN1(n16041), .IN2(n9079), .QN(n11483) );
  NAND2X0 U11563 ( .IN1(n11487), .IN2(n9109), .QN(n11479) );
  INVX0 U11564 ( .INP(n11488), .ZN(n11487) );
  NAND2X0 U11565 ( .IN1(WX512), .IN2(n9278), .QN(n11478) );
  NAND2X0 U11566 ( .IN1(n9311), .IN2(CRC_OUT_9_16), .QN(n11477) );
  NAND4X0 U11567 ( .IN1(n11489), .IN2(n11490), .IN3(n11491), .IN4(n11492), 
        .QN(WX672) );
  NAND2X0 U11568 ( .IN1(n11493), .IN2(n11494), .QN(n11492) );
  NAND3X0 U11569 ( .IN1(n11495), .IN2(n11496), .IN3(n11497), .QN(n11493) );
  NAND2X0 U11570 ( .IN1(n9333), .IN2(n11498), .QN(n11497) );
  NAND2X0 U11571 ( .IN1(n9083), .IN2(n8654), .QN(n11496) );
  NAND2X0 U11572 ( .IN1(n16040), .IN2(n9078), .QN(n11495) );
  NAND2X0 U11573 ( .IN1(n9093), .IN2(n11499), .QN(n11491) );
  NAND2X0 U11574 ( .IN1(WX510), .IN2(n9278), .QN(n11490) );
  NAND2X0 U11575 ( .IN1(n9312), .IN2(CRC_OUT_9_17), .QN(n11489) );
  NAND4X0 U11576 ( .IN1(n11500), .IN2(n11501), .IN3(n11502), .IN4(n11503), 
        .QN(WX670) );
  NAND2X0 U11577 ( .IN1(n11504), .IN2(n9335), .QN(n11503) );
  NAND2X0 U11578 ( .IN1(n9093), .IN2(n11505), .QN(n11502) );
  NAND2X0 U11579 ( .IN1(WX508), .IN2(n9278), .QN(n11501) );
  NAND2X0 U11580 ( .IN1(n9310), .IN2(CRC_OUT_9_18), .QN(n11500) );
  NAND4X0 U11581 ( .IN1(n11506), .IN2(n11507), .IN3(n11508), .IN4(n11509), 
        .QN(WX668) );
  NAND2X0 U11582 ( .IN1(n11510), .IN2(n11511), .QN(n11509) );
  NAND3X0 U11583 ( .IN1(n11512), .IN2(n11513), .IN3(n11514), .QN(n11510) );
  NAND2X0 U11584 ( .IN1(n9333), .IN2(n11515), .QN(n11514) );
  NAND2X0 U11585 ( .IN1(n9082), .IN2(n8656), .QN(n11513) );
  NAND2X0 U11586 ( .IN1(n16038), .IN2(n9077), .QN(n11512) );
  NAND2X0 U11587 ( .IN1(n9093), .IN2(n11516), .QN(n11508) );
  NAND2X0 U11588 ( .IN1(WX506), .IN2(n9278), .QN(n11507) );
  NAND2X0 U11589 ( .IN1(test_so10), .IN2(n9313), .QN(n11506) );
  NAND4X0 U11590 ( .IN1(n11517), .IN2(n11518), .IN3(n11519), .IN4(n11520), 
        .QN(WX666) );
  NAND2X0 U11591 ( .IN1(n11521), .IN2(n11522), .QN(n11520) );
  NAND3X0 U11592 ( .IN1(n11523), .IN2(n11524), .IN3(n11525), .QN(n11521) );
  NAND2X0 U11593 ( .IN1(n9333), .IN2(n11526), .QN(n11525) );
  NAND2X0 U11594 ( .IN1(n9081), .IN2(n8657), .QN(n11524) );
  NAND2X0 U11595 ( .IN1(n16037), .IN2(n9791), .QN(n11523) );
  NAND2X0 U11596 ( .IN1(n11527), .IN2(n9109), .QN(n11519) );
  INVX0 U11597 ( .INP(n11528), .ZN(n11527) );
  NAND2X0 U11598 ( .IN1(WX504), .IN2(n9278), .QN(n11518) );
  NAND2X0 U11599 ( .IN1(n9312), .IN2(CRC_OUT_9_20), .QN(n11517) );
  NAND4X0 U11600 ( .IN1(n11529), .IN2(n11530), .IN3(n11531), .IN4(n11532), 
        .QN(WX664) );
  NAND2X0 U11601 ( .IN1(n11533), .IN2(n11534), .QN(n11532) );
  NAND3X0 U11602 ( .IN1(n11535), .IN2(n11536), .IN3(n11537), .QN(n11533) );
  NAND2X0 U11603 ( .IN1(n9332), .IN2(n11538), .QN(n11537) );
  NAND2X0 U11604 ( .IN1(n9790), .IN2(n8658), .QN(n11536) );
  NAND2X0 U11605 ( .IN1(n16036), .IN2(n9079), .QN(n11535) );
  NAND2X0 U11606 ( .IN1(n9093), .IN2(n11539), .QN(n11531) );
  NAND2X0 U11607 ( .IN1(WX502), .IN2(n9278), .QN(n11530) );
  NAND2X0 U11608 ( .IN1(n9311), .IN2(CRC_OUT_9_21), .QN(n11529) );
  NAND4X0 U11609 ( .IN1(n11540), .IN2(n11541), .IN3(n11542), .IN4(n11543), 
        .QN(WX662) );
  NAND2X0 U11610 ( .IN1(n11544), .IN2(n11545), .QN(n11543) );
  NAND3X0 U11611 ( .IN1(n11546), .IN2(n11547), .IN3(n11548), .QN(n11544) );
  NAND2X0 U11612 ( .IN1(n9333), .IN2(n11549), .QN(n11548) );
  NAND2X0 U11613 ( .IN1(n9078), .IN2(WX2148), .QN(n11547) );
  NAND2X0 U11614 ( .IN1(n9083), .IN2(n8592), .QN(n11546) );
  NAND2X0 U11615 ( .IN1(n9093), .IN2(n11550), .QN(n11542) );
  NAND2X0 U11616 ( .IN1(WX500), .IN2(n9278), .QN(n11541) );
  NAND2X0 U11617 ( .IN1(n9312), .IN2(CRC_OUT_9_22), .QN(n11540) );
  NAND4X0 U11618 ( .IN1(n11551), .IN2(n11552), .IN3(n11553), .IN4(n11554), 
        .QN(WX660) );
  NAND2X0 U11619 ( .IN1(n11555), .IN2(n11556), .QN(n11554) );
  NAND3X0 U11620 ( .IN1(n11557), .IN2(n11558), .IN3(n11559), .QN(n11555) );
  NAND2X0 U11621 ( .IN1(n9333), .IN2(n11560), .QN(n11559) );
  NAND2X0 U11622 ( .IN1(n9082), .IN2(n8661), .QN(n11558) );
  NAND2X0 U11623 ( .IN1(n16035), .IN2(n9078), .QN(n11557) );
  NAND2X0 U11624 ( .IN1(n9093), .IN2(n11561), .QN(n11553) );
  NAND2X0 U11625 ( .IN1(WX498), .IN2(n9278), .QN(n11552) );
  NAND2X0 U11626 ( .IN1(n9310), .IN2(CRC_OUT_9_23), .QN(n11551) );
  NAND4X0 U11627 ( .IN1(n11562), .IN2(n11563), .IN3(n11564), .IN4(n11565), 
        .QN(WX658) );
  NAND2X0 U11628 ( .IN1(n11566), .IN2(n11567), .QN(n11565) );
  NAND3X0 U11629 ( .IN1(n11568), .IN2(n11569), .IN3(n11570), .QN(n11566) );
  NAND2X0 U11630 ( .IN1(n9333), .IN2(n11571), .QN(n11570) );
  NAND2X0 U11631 ( .IN1(n9081), .IN2(n8662), .QN(n11569) );
  NAND2X0 U11632 ( .IN1(n16034), .IN2(n9077), .QN(n11568) );
  NAND2X0 U11633 ( .IN1(n11572), .IN2(n9110), .QN(n11564) );
  INVX0 U11634 ( .INP(n11573), .ZN(n11572) );
  NAND2X0 U11635 ( .IN1(WX496), .IN2(n9278), .QN(n11563) );
  NAND2X0 U11636 ( .IN1(n9312), .IN2(CRC_OUT_9_24), .QN(n11562) );
  NAND4X0 U11637 ( .IN1(n11574), .IN2(n11575), .IN3(n11576), .IN4(n11577), 
        .QN(WX656) );
  NAND2X0 U11638 ( .IN1(n11578), .IN2(n11579), .QN(n11577) );
  NAND3X0 U11639 ( .IN1(n11580), .IN2(n11581), .IN3(n11582), .QN(n11578) );
  NAND2X0 U11640 ( .IN1(n9333), .IN2(n11583), .QN(n11582) );
  NAND2X0 U11641 ( .IN1(n9790), .IN2(n8663), .QN(n11581) );
  NAND2X0 U11642 ( .IN1(n16033), .IN2(n9791), .QN(n11580) );
  NAND2X0 U11643 ( .IN1(n9093), .IN2(n11584), .QN(n11576) );
  NAND2X0 U11644 ( .IN1(WX494), .IN2(n9279), .QN(n11575) );
  NAND2X0 U11645 ( .IN1(n9311), .IN2(CRC_OUT_9_25), .QN(n11574) );
  NAND4X0 U11646 ( .IN1(n11585), .IN2(n11586), .IN3(n11587), .IN4(n11588), 
        .QN(WX654) );
  NAND2X0 U11647 ( .IN1(n11589), .IN2(n11590), .QN(n11588) );
  NAND3X0 U11648 ( .IN1(n11591), .IN2(n11592), .IN3(n11593), .QN(n11589) );
  NAND2X0 U11649 ( .IN1(n9333), .IN2(n11594), .QN(n11593) );
  NAND2X0 U11650 ( .IN1(n9083), .IN2(n8664), .QN(n11592) );
  NAND2X0 U11651 ( .IN1(n16032), .IN2(n9079), .QN(n11591) );
  NAND2X0 U11652 ( .IN1(n9094), .IN2(n11595), .QN(n11587) );
  NAND2X0 U11653 ( .IN1(WX492), .IN2(n9279), .QN(n11586) );
  NAND2X0 U11654 ( .IN1(n9312), .IN2(CRC_OUT_9_26), .QN(n11585) );
  NAND4X0 U11655 ( .IN1(n11596), .IN2(n11597), .IN3(n11598), .IN4(n11599), 
        .QN(WX652) );
  NAND2X0 U11656 ( .IN1(n11600), .IN2(n11601), .QN(n11599) );
  NAND3X0 U11657 ( .IN1(n11602), .IN2(n11603), .IN3(n11604), .QN(n11600) );
  NAND2X0 U11658 ( .IN1(n9333), .IN2(n11605), .QN(n11604) );
  NAND2X0 U11659 ( .IN1(n9082), .IN2(n8665), .QN(n11603) );
  NAND2X0 U11660 ( .IN1(n16031), .IN2(n9078), .QN(n11602) );
  NAND2X0 U11661 ( .IN1(n9094), .IN2(n11606), .QN(n11598) );
  NAND2X0 U11662 ( .IN1(WX490), .IN2(n9279), .QN(n11597) );
  NAND2X0 U11663 ( .IN1(n9311), .IN2(CRC_OUT_9_27), .QN(n11596) );
  NAND4X0 U11664 ( .IN1(n11607), .IN2(n11608), .IN3(n11609), .IN4(n11610), 
        .QN(WX650) );
  NAND2X0 U11665 ( .IN1(n11611), .IN2(n9335), .QN(n11610) );
  NAND2X0 U11666 ( .IN1(n11612), .IN2(n9109), .QN(n11609) );
  INVX0 U11667 ( .INP(n11613), .ZN(n11612) );
  NAND2X0 U11668 ( .IN1(WX488), .IN2(n9279), .QN(n11608) );
  NAND2X0 U11669 ( .IN1(n9311), .IN2(CRC_OUT_9_28), .QN(n11607) );
  NOR3X0 U11670 ( .IN1(n9142), .IN2(n11614), .IN3(n11615), .QN(WX6498) );
  NOR2X0 U11671 ( .IN1(n8238), .IN2(CRC_OUT_5_30), .QN(n11615) );
  NOR2X0 U11672 ( .IN1(DFF_958_n1), .IN2(WX6009), .QN(n11614) );
  NOR3X0 U11673 ( .IN1(n9142), .IN2(n11616), .IN3(n11617), .QN(WX6496) );
  NOR2X0 U11674 ( .IN1(n8239), .IN2(CRC_OUT_5_29), .QN(n11617) );
  NOR2X0 U11675 ( .IN1(DFF_957_n1), .IN2(WX6011), .QN(n11616) );
  NOR3X0 U11676 ( .IN1(n9141), .IN2(n11618), .IN3(n11619), .QN(WX6494) );
  NOR2X0 U11677 ( .IN1(n8240), .IN2(CRC_OUT_5_28), .QN(n11619) );
  NOR2X0 U11678 ( .IN1(DFF_956_n1), .IN2(WX6013), .QN(n11618) );
  NOR3X0 U11679 ( .IN1(n9141), .IN2(n11620), .IN3(n11621), .QN(WX6492) );
  NOR2X0 U11680 ( .IN1(n8241), .IN2(CRC_OUT_5_27), .QN(n11621) );
  NOR2X0 U11681 ( .IN1(DFF_955_n1), .IN2(WX6015), .QN(n11620) );
  NOR3X0 U11682 ( .IN1(n9141), .IN2(n11622), .IN3(n11623), .QN(WX6490) );
  NOR2X0 U11683 ( .IN1(n8242), .IN2(CRC_OUT_5_26), .QN(n11623) );
  NOR2X0 U11684 ( .IN1(DFF_954_n1), .IN2(WX6017), .QN(n11622) );
  NOR3X0 U11685 ( .IN1(n9141), .IN2(n11624), .IN3(n11625), .QN(WX6488) );
  NOR2X0 U11686 ( .IN1(n8243), .IN2(CRC_OUT_5_25), .QN(n11625) );
  NOR2X0 U11687 ( .IN1(DFF_953_n1), .IN2(WX6019), .QN(n11624) );
  NOR3X0 U11688 ( .IN1(n9141), .IN2(n11626), .IN3(n11627), .QN(WX6486) );
  NOR2X0 U11689 ( .IN1(n8244), .IN2(CRC_OUT_5_24), .QN(n11627) );
  NOR2X0 U11690 ( .IN1(DFF_952_n1), .IN2(WX6021), .QN(n11626) );
  NOR3X0 U11691 ( .IN1(n9141), .IN2(n11628), .IN3(n11629), .QN(WX6484) );
  NOR2X0 U11692 ( .IN1(n8245), .IN2(CRC_OUT_5_23), .QN(n11629) );
  NOR2X0 U11693 ( .IN1(DFF_951_n1), .IN2(WX6023), .QN(n11628) );
  NOR3X0 U11694 ( .IN1(n9141), .IN2(n11630), .IN3(n11631), .QN(WX6482) );
  NOR2X0 U11695 ( .IN1(n8255), .IN2(CRC_OUT_5_22), .QN(n11631) );
  NOR2X0 U11696 ( .IN1(DFF_950_n1), .IN2(WX6025), .QN(n11630) );
  NOR3X0 U11697 ( .IN1(n9141), .IN2(n11632), .IN3(n11633), .QN(WX6480) );
  NOR2X0 U11698 ( .IN1(n8256), .IN2(CRC_OUT_5_21), .QN(n11633) );
  NOR2X0 U11699 ( .IN1(DFF_949_n1), .IN2(WX6027), .QN(n11632) );
  NAND4X0 U11700 ( .IN1(n11634), .IN2(n11635), .IN3(n11636), .IN4(n11637), 
        .QN(WX648) );
  NAND2X0 U11701 ( .IN1(n11638), .IN2(n11639), .QN(n11637) );
  NAND3X0 U11702 ( .IN1(n11640), .IN2(n11641), .IN3(n11642), .QN(n11638) );
  NAND2X0 U11703 ( .IN1(n9333), .IN2(n11643), .QN(n11642) );
  NAND2X0 U11704 ( .IN1(n9081), .IN2(n8667), .QN(n11641) );
  NAND2X0 U11705 ( .IN1(n16029), .IN2(n9077), .QN(n11640) );
  NAND2X0 U11706 ( .IN1(n9094), .IN2(n11644), .QN(n11636) );
  NAND2X0 U11707 ( .IN1(WX486), .IN2(n9279), .QN(n11635) );
  NAND2X0 U11708 ( .IN1(n9312), .IN2(CRC_OUT_9_29), .QN(n11634) );
  NOR3X0 U11709 ( .IN1(n9141), .IN2(n11645), .IN3(n11646), .QN(WX6478) );
  NOR2X0 U11710 ( .IN1(n8273), .IN2(CRC_OUT_5_20), .QN(n11646) );
  NOR2X0 U11711 ( .IN1(DFF_948_n1), .IN2(WX6029), .QN(n11645) );
  NOR3X0 U11712 ( .IN1(n9141), .IN2(n11647), .IN3(n11648), .QN(WX6476) );
  NOR2X0 U11713 ( .IN1(n8274), .IN2(CRC_OUT_5_19), .QN(n11648) );
  NOR2X0 U11714 ( .IN1(DFF_947_n1), .IN2(WX6031), .QN(n11647) );
  NOR3X0 U11715 ( .IN1(n9141), .IN2(n11649), .IN3(n11650), .QN(WX6474) );
  NOR2X0 U11716 ( .IN1(n8291), .IN2(CRC_OUT_5_18), .QN(n11650) );
  NOR2X0 U11717 ( .IN1(DFF_946_n1), .IN2(WX6033), .QN(n11649) );
  NOR2X0 U11718 ( .IN1(n9225), .IN2(n11651), .QN(WX6472) );
  NOR2X0 U11719 ( .IN1(n11652), .IN2(n11653), .QN(n11651) );
  NOR2X0 U11720 ( .IN1(test_so54), .IN2(WX6035), .QN(n11653) );
  NOR2X0 U11721 ( .IN1(n8292), .IN2(n8827), .QN(n11652) );
  NOR3X0 U11722 ( .IN1(n9141), .IN2(n11654), .IN3(n11655), .QN(WX6470) );
  NOR2X0 U11723 ( .IN1(n8296), .IN2(CRC_OUT_5_16), .QN(n11655) );
  NOR2X0 U11724 ( .IN1(DFF_944_n1), .IN2(WX6037), .QN(n11654) );
  NOR3X0 U11725 ( .IN1(n9140), .IN2(n11656), .IN3(n11657), .QN(WX6468) );
  INVX0 U11726 ( .INP(n11658), .ZN(n11657) );
  NAND2X0 U11727 ( .IN1(CRC_OUT_5_15), .IN2(n11659), .QN(n11658) );
  NOR2X0 U11728 ( .IN1(n11659), .IN2(CRC_OUT_5_15), .QN(n11656) );
  NAND2X0 U11729 ( .IN1(n11660), .IN2(n11661), .QN(n11659) );
  NAND2X0 U11730 ( .IN1(test_so52), .IN2(CRC_OUT_5_31), .QN(n11661) );
  NAND2X0 U11731 ( .IN1(DFF_959_n1), .IN2(n8826), .QN(n11660) );
  NOR3X0 U11732 ( .IN1(n9140), .IN2(n11662), .IN3(n11663), .QN(WX6466) );
  NOR2X0 U11733 ( .IN1(n8297), .IN2(CRC_OUT_5_14), .QN(n11663) );
  NOR2X0 U11734 ( .IN1(DFF_942_n1), .IN2(WX6041), .QN(n11662) );
  NOR3X0 U11735 ( .IN1(n9140), .IN2(n11664), .IN3(n11665), .QN(WX6464) );
  NOR2X0 U11736 ( .IN1(n8298), .IN2(CRC_OUT_5_13), .QN(n11665) );
  NOR2X0 U11737 ( .IN1(DFF_941_n1), .IN2(WX6043), .QN(n11664) );
  NOR3X0 U11738 ( .IN1(n9140), .IN2(n11666), .IN3(n11667), .QN(WX6462) );
  NOR2X0 U11739 ( .IN1(n8299), .IN2(CRC_OUT_5_12), .QN(n11667) );
  NOR2X0 U11740 ( .IN1(DFF_940_n1), .IN2(WX6045), .QN(n11666) );
  NOR3X0 U11741 ( .IN1(n9140), .IN2(n11668), .IN3(n11669), .QN(WX6460) );
  NOR2X0 U11742 ( .IN1(n8300), .IN2(CRC_OUT_5_11), .QN(n11669) );
  NOR2X0 U11743 ( .IN1(DFF_939_n1), .IN2(WX6047), .QN(n11668) );
  NAND4X0 U11744 ( .IN1(n11670), .IN2(n11671), .IN3(n11672), .IN4(n11673), 
        .QN(WX646) );
  NAND2X0 U11745 ( .IN1(n11674), .IN2(n11675), .QN(n11673) );
  NAND3X0 U11746 ( .IN1(n11676), .IN2(n11677), .IN3(n11678), .QN(n11674) );
  NAND2X0 U11747 ( .IN1(n9333), .IN2(n11679), .QN(n11678) );
  NAND2X0 U11748 ( .IN1(n9790), .IN2(n8668), .QN(n11677) );
  NAND2X0 U11749 ( .IN1(n16028), .IN2(n9791), .QN(n11676) );
  NAND2X0 U11750 ( .IN1(n9094), .IN2(n11680), .QN(n11672) );
  NAND2X0 U11751 ( .IN1(WX484), .IN2(n9279), .QN(n11671) );
  NAND2X0 U11752 ( .IN1(n9313), .IN2(CRC_OUT_9_30), .QN(n11670) );
  NOR2X0 U11753 ( .IN1(n9240), .IN2(n11681), .QN(WX6458) );
  NOR2X0 U11754 ( .IN1(n11682), .IN2(n11683), .QN(n11681) );
  INVX0 U11755 ( .INP(n11684), .ZN(n11683) );
  NAND2X0 U11756 ( .IN1(CRC_OUT_5_10), .IN2(n11685), .QN(n11684) );
  NOR2X0 U11757 ( .IN1(n11685), .IN2(CRC_OUT_5_10), .QN(n11682) );
  NAND2X0 U11758 ( .IN1(n11686), .IN2(n11687), .QN(n11685) );
  NAND2X0 U11759 ( .IN1(n8115), .IN2(CRC_OUT_5_31), .QN(n11687) );
  NAND2X0 U11760 ( .IN1(DFF_959_n1), .IN2(WX6049), .QN(n11686) );
  NOR3X0 U11761 ( .IN1(n9140), .IN2(n11688), .IN3(n11689), .QN(WX6456) );
  NOR2X0 U11762 ( .IN1(n8301), .IN2(CRC_OUT_5_9), .QN(n11689) );
  NOR2X0 U11763 ( .IN1(DFF_937_n1), .IN2(WX6051), .QN(n11688) );
  NOR3X0 U11764 ( .IN1(n9140), .IN2(n11690), .IN3(n11691), .QN(WX6454) );
  NOR2X0 U11765 ( .IN1(n8302), .IN2(CRC_OUT_5_8), .QN(n11691) );
  NOR2X0 U11766 ( .IN1(DFF_936_n1), .IN2(WX6053), .QN(n11690) );
  NOR3X0 U11767 ( .IN1(n9140), .IN2(n11692), .IN3(n11693), .QN(WX6452) );
  NOR2X0 U11768 ( .IN1(n8303), .IN2(CRC_OUT_5_7), .QN(n11693) );
  NOR2X0 U11769 ( .IN1(DFF_935_n1), .IN2(WX6055), .QN(n11692) );
  NOR3X0 U11770 ( .IN1(n9140), .IN2(n11694), .IN3(n11695), .QN(WX6450) );
  NOR2X0 U11771 ( .IN1(n8308), .IN2(CRC_OUT_5_6), .QN(n11695) );
  NOR2X0 U11772 ( .IN1(DFF_934_n1), .IN2(WX6057), .QN(n11694) );
  NOR3X0 U11773 ( .IN1(n9140), .IN2(n11696), .IN3(n11697), .QN(WX6448) );
  NOR2X0 U11774 ( .IN1(n8309), .IN2(CRC_OUT_5_5), .QN(n11697) );
  NOR2X0 U11775 ( .IN1(DFF_933_n1), .IN2(WX6059), .QN(n11696) );
  NOR3X0 U11776 ( .IN1(n9140), .IN2(n11698), .IN3(n11699), .QN(WX6446) );
  NOR2X0 U11777 ( .IN1(n8326), .IN2(CRC_OUT_5_4), .QN(n11699) );
  NOR2X0 U11778 ( .IN1(DFF_932_n1), .IN2(WX6061), .QN(n11698) );
  NOR2X0 U11779 ( .IN1(n9240), .IN2(n11700), .QN(WX6444) );
  NOR2X0 U11780 ( .IN1(n11701), .IN2(n11702), .QN(n11700) );
  INVX0 U11781 ( .INP(n11703), .ZN(n11702) );
  NAND2X0 U11782 ( .IN1(CRC_OUT_5_3), .IN2(n11704), .QN(n11703) );
  NOR2X0 U11783 ( .IN1(n11704), .IN2(CRC_OUT_5_3), .QN(n11701) );
  NAND2X0 U11784 ( .IN1(n11705), .IN2(n11706), .QN(n11704) );
  NAND2X0 U11785 ( .IN1(n8116), .IN2(CRC_OUT_5_31), .QN(n11706) );
  NAND2X0 U11786 ( .IN1(DFF_959_n1), .IN2(WX6063), .QN(n11705) );
  NOR3X0 U11787 ( .IN1(n9139), .IN2(n11707), .IN3(n11708), .QN(WX6442) );
  NOR2X0 U11788 ( .IN1(n8327), .IN2(CRC_OUT_5_2), .QN(n11708) );
  NOR2X0 U11789 ( .IN1(DFF_930_n1), .IN2(WX6065), .QN(n11707) );
  NOR3X0 U11790 ( .IN1(n9139), .IN2(n11709), .IN3(n11710), .QN(WX6440) );
  NOR2X0 U11791 ( .IN1(n8344), .IN2(CRC_OUT_5_1), .QN(n11710) );
  NOR2X0 U11792 ( .IN1(DFF_929_n1), .IN2(WX6067), .QN(n11709) );
  NAND4X0 U11793 ( .IN1(n11711), .IN2(n11712), .IN3(n11713), .IN4(n11714), 
        .QN(WX644) );
  NAND2X0 U11794 ( .IN1(n11715), .IN2(n11716), .QN(n11714) );
  NAND3X0 U11795 ( .IN1(n11717), .IN2(n11718), .IN3(n11719), .QN(n11715) );
  NAND2X0 U11796 ( .IN1(n9333), .IN2(n11720), .QN(n11719) );
  NAND2X0 U11797 ( .IN1(n9083), .IN2(n8669), .QN(n11718) );
  NAND2X0 U11798 ( .IN1(n16027), .IN2(n9079), .QN(n11717) );
  NAND2X0 U11799 ( .IN1(n9094), .IN2(n11721), .QN(n11713) );
  NAND2X0 U11800 ( .IN1(n9312), .IN2(CRC_OUT_9_31), .QN(n11712) );
  NAND2X0 U11801 ( .IN1(n2245), .IN2(WX485), .QN(n11711) );
  NOR2X0 U11802 ( .IN1(n9240), .IN2(n11722), .QN(WX6438) );
  NOR2X0 U11803 ( .IN1(n11723), .IN2(n11724), .QN(n11722) );
  NOR2X0 U11804 ( .IN1(test_so53), .IN2(WX6069), .QN(n11724) );
  INVX0 U11805 ( .INP(n11725), .ZN(n11723) );
  NAND2X0 U11806 ( .IN1(WX6069), .IN2(test_so53), .QN(n11725) );
  NOR3X0 U11807 ( .IN1(n9139), .IN2(n11726), .IN3(n11727), .QN(WX6436) );
  NOR2X0 U11808 ( .IN1(n8129), .IN2(CRC_OUT_5_31), .QN(n11727) );
  NOR2X0 U11809 ( .IN1(DFF_959_n1), .IN2(WX6071), .QN(n11726) );
  NOR2X0 U11810 ( .IN1(n16086), .IN2(n9161), .QN(WX5910) );
  NOR2X0 U11811 ( .IN1(n16085), .IN2(n9163), .QN(WX5908) );
  NOR2X0 U11812 ( .IN1(n16084), .IN2(n9163), .QN(WX5906) );
  NOR2X0 U11813 ( .IN1(n16083), .IN2(n9162), .QN(WX5904) );
  NOR2X0 U11814 ( .IN1(n16082), .IN2(n9162), .QN(WX5902) );
  NOR2X0 U11815 ( .IN1(n16081), .IN2(n9162), .QN(WX5900) );
  NOR2X0 U11816 ( .IN1(n9240), .IN2(n8821), .QN(WX5898) );
  NOR2X0 U11817 ( .IN1(n16080), .IN2(n9162), .QN(WX5896) );
  NOR2X0 U11818 ( .IN1(n16079), .IN2(n9162), .QN(WX5894) );
  NOR2X0 U11819 ( .IN1(n16078), .IN2(n9162), .QN(WX5892) );
  NOR2X0 U11820 ( .IN1(n16077), .IN2(n9162), .QN(WX5890) );
  NOR2X0 U11821 ( .IN1(n16076), .IN2(n9162), .QN(WX5888) );
  NOR2X0 U11822 ( .IN1(n16075), .IN2(n9162), .QN(WX5886) );
  NOR2X0 U11823 ( .IN1(n16074), .IN2(n9162), .QN(WX5884) );
  NOR2X0 U11824 ( .IN1(n16073), .IN2(n9162), .QN(WX5882) );
  NOR2X0 U11825 ( .IN1(n16072), .IN2(n9162), .QN(WX5880) );
  NAND4X0 U11826 ( .IN1(n11728), .IN2(n11729), .IN3(n11730), .IN4(n11731), 
        .QN(WX5878) );
  NAND2X0 U11827 ( .IN1(n9333), .IN2(n10784), .QN(n11731) );
  NAND2X0 U11828 ( .IN1(n11732), .IN2(n11733), .QN(n10784) );
  INVX0 U11829 ( .INP(n11734), .ZN(n11733) );
  NOR2X0 U11830 ( .IN1(n11735), .IN2(n11736), .QN(n11734) );
  NAND2X0 U11831 ( .IN1(n11736), .IN2(n11735), .QN(n11732) );
  NOR2X0 U11832 ( .IN1(n11737), .IN2(n11738), .QN(n11735) );
  NOR2X0 U11833 ( .IN1(WX7364), .IN2(n7945), .QN(n11738) );
  INVX0 U11834 ( .INP(n11739), .ZN(n11737) );
  NAND2X0 U11835 ( .IN1(n7945), .IN2(WX7364), .QN(n11739) );
  NAND2X0 U11836 ( .IN1(n11740), .IN2(n11741), .QN(n11736) );
  NAND2X0 U11837 ( .IN1(n7944), .IN2(WX7236), .QN(n11741) );
  INVX0 U11838 ( .INP(n11742), .ZN(n11740) );
  NOR2X0 U11839 ( .IN1(WX7236), .IN2(n7944), .QN(n11742) );
  NAND2X0 U11840 ( .IN1(n9094), .IN2(n11743), .QN(n11730) );
  NAND2X0 U11841 ( .IN1(n1003), .IN2(n9279), .QN(n11729) );
  NOR2X0 U11842 ( .IN1(n9239), .IN2(n8915), .QN(n1003) );
  NAND2X0 U11843 ( .IN1(test_so53), .IN2(n9314), .QN(n11728) );
  NAND4X0 U11844 ( .IN1(n11744), .IN2(n11745), .IN3(n11746), .IN4(n11747), 
        .QN(WX5876) );
  NAND3X0 U11845 ( .IN1(n11748), .IN2(n11749), .IN3(n9089), .QN(n11747) );
  NAND2X0 U11846 ( .IN1(n9333), .IN2(n10800), .QN(n11746) );
  NAND2X0 U11847 ( .IN1(n11750), .IN2(n11751), .QN(n10800) );
  INVX0 U11848 ( .INP(n11752), .ZN(n11751) );
  NOR2X0 U11849 ( .IN1(n11753), .IN2(n11754), .QN(n11752) );
  NAND2X0 U11850 ( .IN1(n11754), .IN2(n11753), .QN(n11750) );
  NOR2X0 U11851 ( .IN1(n11755), .IN2(n11756), .QN(n11753) );
  NOR2X0 U11852 ( .IN1(WX7362), .IN2(n7947), .QN(n11756) );
  INVX0 U11853 ( .INP(n11757), .ZN(n11755) );
  NAND2X0 U11854 ( .IN1(n7947), .IN2(WX7362), .QN(n11757) );
  NAND2X0 U11855 ( .IN1(n11758), .IN2(n11759), .QN(n11754) );
  NAND2X0 U11856 ( .IN1(n7946), .IN2(WX7234), .QN(n11759) );
  INVX0 U11857 ( .INP(n11760), .ZN(n11758) );
  NOR2X0 U11858 ( .IN1(WX7234), .IN2(n7946), .QN(n11760) );
  NAND2X0 U11859 ( .IN1(n1002), .IN2(n9279), .QN(n11745) );
  NOR2X0 U11860 ( .IN1(n9239), .IN2(n8916), .QN(n1002) );
  NAND2X0 U11861 ( .IN1(n9311), .IN2(CRC_OUT_5_1), .QN(n11744) );
  NAND4X0 U11862 ( .IN1(n11761), .IN2(n11762), .IN3(n11763), .IN4(n11764), 
        .QN(WX5874) );
  NAND2X0 U11863 ( .IN1(n9324), .IN2(n10816), .QN(n11764) );
  NAND2X0 U11864 ( .IN1(n11765), .IN2(n11766), .QN(n10816) );
  INVX0 U11865 ( .INP(n11767), .ZN(n11766) );
  NOR2X0 U11866 ( .IN1(n11768), .IN2(n11769), .QN(n11767) );
  NAND2X0 U11867 ( .IN1(n11769), .IN2(n11768), .QN(n11765) );
  NOR2X0 U11868 ( .IN1(n11770), .IN2(n11771), .QN(n11768) );
  NOR2X0 U11869 ( .IN1(WX7360), .IN2(n7949), .QN(n11771) );
  INVX0 U11870 ( .INP(n11772), .ZN(n11770) );
  NAND2X0 U11871 ( .IN1(n7949), .IN2(WX7360), .QN(n11772) );
  NAND2X0 U11872 ( .IN1(n11773), .IN2(n11774), .QN(n11769) );
  NAND2X0 U11873 ( .IN1(n7948), .IN2(WX7232), .QN(n11774) );
  INVX0 U11874 ( .INP(n11775), .ZN(n11773) );
  NOR2X0 U11875 ( .IN1(WX7232), .IN2(n7948), .QN(n11775) );
  NAND2X0 U11876 ( .IN1(n9094), .IN2(n11776), .QN(n11763) );
  NAND2X0 U11877 ( .IN1(n1001), .IN2(n9279), .QN(n11762) );
  NOR2X0 U11878 ( .IN1(n9239), .IN2(n8917), .QN(n1001) );
  NAND2X0 U11879 ( .IN1(n9313), .IN2(CRC_OUT_5_2), .QN(n11761) );
  NAND4X0 U11880 ( .IN1(n11777), .IN2(n11778), .IN3(n11779), .IN4(n11780), 
        .QN(WX5872) );
  NAND3X0 U11881 ( .IN1(n11781), .IN2(n11782), .IN3(n9090), .QN(n11780) );
  NAND2X0 U11882 ( .IN1(n9322), .IN2(n10832), .QN(n11779) );
  NAND2X0 U11883 ( .IN1(n11783), .IN2(n11784), .QN(n10832) );
  INVX0 U11884 ( .INP(n11785), .ZN(n11784) );
  NOR2X0 U11885 ( .IN1(n11786), .IN2(n11787), .QN(n11785) );
  NAND2X0 U11886 ( .IN1(n11787), .IN2(n11786), .QN(n11783) );
  NOR2X0 U11887 ( .IN1(n11788), .IN2(n11789), .QN(n11786) );
  NOR2X0 U11888 ( .IN1(WX7358), .IN2(n7951), .QN(n11789) );
  INVX0 U11889 ( .INP(n11790), .ZN(n11788) );
  NAND2X0 U11890 ( .IN1(n7951), .IN2(WX7358), .QN(n11790) );
  NAND2X0 U11891 ( .IN1(n11791), .IN2(n11792), .QN(n11787) );
  NAND2X0 U11892 ( .IN1(n7950), .IN2(WX7230), .QN(n11792) );
  INVX0 U11893 ( .INP(n11793), .ZN(n11791) );
  NOR2X0 U11894 ( .IN1(WX7230), .IN2(n7950), .QN(n11793) );
  NAND2X0 U11895 ( .IN1(n1000), .IN2(n9279), .QN(n11778) );
  NOR2X0 U11896 ( .IN1(n9239), .IN2(n8918), .QN(n1000) );
  NAND2X0 U11897 ( .IN1(n9312), .IN2(CRC_OUT_5_3), .QN(n11777) );
  NAND4X0 U11898 ( .IN1(n11794), .IN2(n11795), .IN3(n11796), .IN4(n11797), 
        .QN(WX5870) );
  NAND3X0 U11899 ( .IN1(n10837), .IN2(n10838), .IN3(n9320), .QN(n11797) );
  NAND3X0 U11900 ( .IN1(n11798), .IN2(n11799), .IN3(n11800), .QN(n10838) );
  INVX0 U11901 ( .INP(n11801), .ZN(n11800) );
  NAND2X0 U11902 ( .IN1(n11801), .IN2(n11802), .QN(n10837) );
  NAND2X0 U11903 ( .IN1(n11798), .IN2(n11799), .QN(n11802) );
  NAND2X0 U11904 ( .IN1(n7953), .IN2(WX7228), .QN(n11799) );
  NAND2X0 U11905 ( .IN1(n3635), .IN2(WX7292), .QN(n11798) );
  NOR2X0 U11906 ( .IN1(n11803), .IN2(n11804), .QN(n11801) );
  NOR2X0 U11907 ( .IN1(n8795), .IN2(n7952), .QN(n11804) );
  INVX0 U11908 ( .INP(n11805), .ZN(n11803) );
  NAND2X0 U11909 ( .IN1(n7952), .IN2(n8795), .QN(n11805) );
  NAND2X0 U11910 ( .IN1(n9094), .IN2(n11806), .QN(n11796) );
  NAND2X0 U11911 ( .IN1(n999), .IN2(n9279), .QN(n11795) );
  NOR2X0 U11912 ( .IN1(n9239), .IN2(n8919), .QN(n999) );
  NAND2X0 U11913 ( .IN1(n9313), .IN2(CRC_OUT_5_4), .QN(n11794) );
  NAND4X0 U11914 ( .IN1(n11807), .IN2(n11808), .IN3(n11809), .IN4(n11810), 
        .QN(WX5868) );
  NAND3X0 U11915 ( .IN1(n11811), .IN2(n11812), .IN3(n9090), .QN(n11810) );
  NAND2X0 U11916 ( .IN1(n9323), .IN2(n10865), .QN(n11809) );
  NAND2X0 U11917 ( .IN1(n11813), .IN2(n11814), .QN(n10865) );
  INVX0 U11918 ( .INP(n11815), .ZN(n11814) );
  NOR2X0 U11919 ( .IN1(n11816), .IN2(n11817), .QN(n11815) );
  NAND2X0 U11920 ( .IN1(n11817), .IN2(n11816), .QN(n11813) );
  NOR2X0 U11921 ( .IN1(n11818), .IN2(n11819), .QN(n11816) );
  NOR2X0 U11922 ( .IN1(WX7354), .IN2(n7955), .QN(n11819) );
  INVX0 U11923 ( .INP(n11820), .ZN(n11818) );
  NAND2X0 U11924 ( .IN1(n7955), .IN2(WX7354), .QN(n11820) );
  NAND2X0 U11925 ( .IN1(n11821), .IN2(n11822), .QN(n11817) );
  NAND2X0 U11926 ( .IN1(n7954), .IN2(WX7226), .QN(n11822) );
  INVX0 U11927 ( .INP(n11823), .ZN(n11821) );
  NOR2X0 U11928 ( .IN1(WX7226), .IN2(n7954), .QN(n11823) );
  NAND2X0 U11929 ( .IN1(n998), .IN2(n9279), .QN(n11808) );
  NOR2X0 U11930 ( .IN1(n9239), .IN2(n8920), .QN(n998) );
  NAND2X0 U11931 ( .IN1(n9312), .IN2(CRC_OUT_5_5), .QN(n11807) );
  NAND4X0 U11932 ( .IN1(n11824), .IN2(n11825), .IN3(n11826), .IN4(n11827), 
        .QN(WX5866) );
  NAND3X0 U11933 ( .IN1(n10870), .IN2(n10871), .IN3(n9320), .QN(n11827) );
  NAND3X0 U11934 ( .IN1(n11828), .IN2(n11829), .IN3(n11830), .QN(n10871) );
  INVX0 U11935 ( .INP(n11831), .ZN(n11830) );
  NAND2X0 U11936 ( .IN1(n11831), .IN2(n11832), .QN(n10870) );
  NAND2X0 U11937 ( .IN1(n11828), .IN2(n11829), .QN(n11832) );
  NAND2X0 U11938 ( .IN1(n8233), .IN2(WX7224), .QN(n11829) );
  NAND2X0 U11939 ( .IN1(n3639), .IN2(WX7352), .QN(n11828) );
  NOR2X0 U11940 ( .IN1(n11833), .IN2(n11834), .QN(n11831) );
  INVX0 U11941 ( .INP(n11835), .ZN(n11834) );
  NAND2X0 U11942 ( .IN1(test_so62), .IN2(WX7160), .QN(n11835) );
  NOR2X0 U11943 ( .IN1(WX7160), .IN2(test_so62), .QN(n11833) );
  NAND2X0 U11944 ( .IN1(n9094), .IN2(n11836), .QN(n11826) );
  NAND2X0 U11945 ( .IN1(n997), .IN2(n9279), .QN(n11825) );
  NOR2X0 U11946 ( .IN1(n9238), .IN2(n8921), .QN(n997) );
  NAND2X0 U11947 ( .IN1(n9313), .IN2(CRC_OUT_5_6), .QN(n11824) );
  NAND4X0 U11948 ( .IN1(n11837), .IN2(n11838), .IN3(n11839), .IN4(n11840), 
        .QN(WX5864) );
  NAND2X0 U11949 ( .IN1(n9322), .IN2(n10898), .QN(n11840) );
  NAND2X0 U11950 ( .IN1(n11841), .IN2(n11842), .QN(n10898) );
  INVX0 U11951 ( .INP(n11843), .ZN(n11842) );
  NOR2X0 U11952 ( .IN1(n11844), .IN2(n11845), .QN(n11843) );
  NAND2X0 U11953 ( .IN1(n11845), .IN2(n11844), .QN(n11841) );
  NOR2X0 U11954 ( .IN1(n11846), .IN2(n11847), .QN(n11844) );
  NOR2X0 U11955 ( .IN1(WX7350), .IN2(n7958), .QN(n11847) );
  INVX0 U11956 ( .INP(n11848), .ZN(n11846) );
  NAND2X0 U11957 ( .IN1(n7958), .IN2(WX7350), .QN(n11848) );
  NAND2X0 U11958 ( .IN1(n11849), .IN2(n11850), .QN(n11845) );
  NAND2X0 U11959 ( .IN1(n7957), .IN2(WX7222), .QN(n11850) );
  INVX0 U11960 ( .INP(n11851), .ZN(n11849) );
  NOR2X0 U11961 ( .IN1(WX7222), .IN2(n7957), .QN(n11851) );
  NAND2X0 U11962 ( .IN1(n9094), .IN2(n11852), .QN(n11839) );
  NAND2X0 U11963 ( .IN1(n996), .IN2(n9279), .QN(n11838) );
  NOR2X0 U11964 ( .IN1(n9066), .IN2(n9162), .QN(n996) );
  NAND2X0 U11965 ( .IN1(n9313), .IN2(CRC_OUT_5_7), .QN(n11837) );
  NAND4X0 U11966 ( .IN1(n11853), .IN2(n11854), .IN3(n11855), .IN4(n11856), 
        .QN(WX5862) );
  NAND3X0 U11967 ( .IN1(n10903), .IN2(n10904), .IN3(n9320), .QN(n11856) );
  NAND3X0 U11968 ( .IN1(n11857), .IN2(n11858), .IN3(n11859), .QN(n10904) );
  INVX0 U11969 ( .INP(n11860), .ZN(n11859) );
  NAND2X0 U11970 ( .IN1(n11860), .IN2(n11861), .QN(n10903) );
  NAND2X0 U11971 ( .IN1(n11857), .IN2(n11858), .QN(n11861) );
  NAND2X0 U11972 ( .IN1(n8231), .IN2(WX7284), .QN(n11858) );
  NAND2X0 U11973 ( .IN1(n7960), .IN2(WX7348), .QN(n11857) );
  NOR2X0 U11974 ( .IN1(n11862), .IN2(n11863), .QN(n11860) );
  INVX0 U11975 ( .INP(n11864), .ZN(n11863) );
  NAND2X0 U11976 ( .IN1(test_so60), .IN2(WX7156), .QN(n11864) );
  NOR2X0 U11977 ( .IN1(WX7156), .IN2(test_so60), .QN(n11862) );
  NAND2X0 U11978 ( .IN1(n9094), .IN2(n11865), .QN(n11855) );
  NAND2X0 U11979 ( .IN1(n995), .IN2(n9279), .QN(n11854) );
  NOR2X0 U11980 ( .IN1(n9238), .IN2(n8922), .QN(n995) );
  NAND2X0 U11981 ( .IN1(n9312), .IN2(CRC_OUT_5_8), .QN(n11853) );
  NAND4X0 U11982 ( .IN1(n11866), .IN2(n11867), .IN3(n11868), .IN4(n11869), 
        .QN(WX5860) );
  NAND2X0 U11983 ( .IN1(n9323), .IN2(n10928), .QN(n11869) );
  NAND2X0 U11984 ( .IN1(n11870), .IN2(n11871), .QN(n10928) );
  INVX0 U11985 ( .INP(n11872), .ZN(n11871) );
  NOR2X0 U11986 ( .IN1(n11873), .IN2(n11874), .QN(n11872) );
  NAND2X0 U11987 ( .IN1(n11874), .IN2(n11873), .QN(n11870) );
  NOR2X0 U11988 ( .IN1(n11875), .IN2(n11876), .QN(n11873) );
  NOR2X0 U11989 ( .IN1(WX7346), .IN2(n7962), .QN(n11876) );
  INVX0 U11990 ( .INP(n11877), .ZN(n11875) );
  NAND2X0 U11991 ( .IN1(n7962), .IN2(WX7346), .QN(n11877) );
  NAND2X0 U11992 ( .IN1(n11878), .IN2(n11879), .QN(n11874) );
  NAND2X0 U11993 ( .IN1(n7961), .IN2(WX7218), .QN(n11879) );
  INVX0 U11994 ( .INP(n11880), .ZN(n11878) );
  NOR2X0 U11995 ( .IN1(WX7218), .IN2(n7961), .QN(n11880) );
  NAND2X0 U11996 ( .IN1(n9094), .IN2(n11881), .QN(n11868) );
  NAND2X0 U11997 ( .IN1(n994), .IN2(n9279), .QN(n11867) );
  NOR2X0 U11998 ( .IN1(n9238), .IN2(n8923), .QN(n994) );
  NAND2X0 U11999 ( .IN1(n9313), .IN2(CRC_OUT_5_9), .QN(n11866) );
  NAND4X0 U12000 ( .IN1(n11882), .IN2(n11883), .IN3(n11884), .IN4(n11885), 
        .QN(WX5858) );
  NAND3X0 U12001 ( .IN1(n10933), .IN2(n10934), .IN3(n9320), .QN(n11885) );
  NAND3X0 U12002 ( .IN1(n11886), .IN2(n11887), .IN3(n11888), .QN(n10934) );
  INVX0 U12003 ( .INP(n11889), .ZN(n11888) );
  NAND2X0 U12004 ( .IN1(n11889), .IN2(n11890), .QN(n10933) );
  NAND2X0 U12005 ( .IN1(n11886), .IN2(n11887), .QN(n11890) );
  NAND2X0 U12006 ( .IN1(n8229), .IN2(WX7216), .QN(n11887) );
  NAND2X0 U12007 ( .IN1(n3647), .IN2(WX7344), .QN(n11886) );
  NOR2X0 U12008 ( .IN1(n11891), .IN2(n11892), .QN(n11889) );
  INVX0 U12009 ( .INP(n11893), .ZN(n11892) );
  NAND2X0 U12010 ( .IN1(test_so58), .IN2(WX7280), .QN(n11893) );
  NOR2X0 U12011 ( .IN1(WX7280), .IN2(test_so58), .QN(n11891) );
  NAND2X0 U12012 ( .IN1(n9094), .IN2(n11894), .QN(n11884) );
  NAND2X0 U12013 ( .IN1(n993), .IN2(n9279), .QN(n11883) );
  NOR2X0 U12014 ( .IN1(n9236), .IN2(n8924), .QN(n993) );
  NAND2X0 U12015 ( .IN1(n9312), .IN2(CRC_OUT_5_10), .QN(n11882) );
  NAND4X0 U12016 ( .IN1(n11895), .IN2(n11896), .IN3(n11897), .IN4(n11898), 
        .QN(WX5856) );
  NAND2X0 U12017 ( .IN1(n9322), .IN2(n10958), .QN(n11898) );
  NAND2X0 U12018 ( .IN1(n11899), .IN2(n11900), .QN(n10958) );
  INVX0 U12019 ( .INP(n11901), .ZN(n11900) );
  NOR2X0 U12020 ( .IN1(n11902), .IN2(n11903), .QN(n11901) );
  NAND2X0 U12021 ( .IN1(n11903), .IN2(n11902), .QN(n11899) );
  NOR2X0 U12022 ( .IN1(n11904), .IN2(n11905), .QN(n11902) );
  NOR2X0 U12023 ( .IN1(WX7342), .IN2(n7965), .QN(n11905) );
  INVX0 U12024 ( .INP(n11906), .ZN(n11904) );
  NAND2X0 U12025 ( .IN1(n7965), .IN2(WX7342), .QN(n11906) );
  NAND2X0 U12026 ( .IN1(n11907), .IN2(n11908), .QN(n11903) );
  NAND2X0 U12027 ( .IN1(n7964), .IN2(WX7214), .QN(n11908) );
  INVX0 U12028 ( .INP(n11909), .ZN(n11907) );
  NOR2X0 U12029 ( .IN1(WX7214), .IN2(n7964), .QN(n11909) );
  NAND2X0 U12030 ( .IN1(n9094), .IN2(n11910), .QN(n11897) );
  NAND2X0 U12031 ( .IN1(n992), .IN2(n9280), .QN(n11896) );
  NOR2X0 U12032 ( .IN1(n9236), .IN2(n8925), .QN(n992) );
  NAND2X0 U12033 ( .IN1(n9311), .IN2(CRC_OUT_5_11), .QN(n11895) );
  NAND4X0 U12034 ( .IN1(n11911), .IN2(n11912), .IN3(n11913), .IN4(n11914), 
        .QN(WX5854) );
  NAND2X0 U12035 ( .IN1(n9322), .IN2(n10974), .QN(n11914) );
  NAND2X0 U12036 ( .IN1(n11915), .IN2(n11916), .QN(n10974) );
  INVX0 U12037 ( .INP(n11917), .ZN(n11916) );
  NOR2X0 U12038 ( .IN1(n11918), .IN2(n11919), .QN(n11917) );
  NAND2X0 U12039 ( .IN1(n11919), .IN2(n11918), .QN(n11915) );
  NOR2X0 U12040 ( .IN1(n11920), .IN2(n11921), .QN(n11918) );
  NOR2X0 U12041 ( .IN1(WX7340), .IN2(n7967), .QN(n11921) );
  INVX0 U12042 ( .INP(n11922), .ZN(n11920) );
  NAND2X0 U12043 ( .IN1(n7967), .IN2(WX7340), .QN(n11922) );
  NAND2X0 U12044 ( .IN1(n11923), .IN2(n11924), .QN(n11919) );
  NAND2X0 U12045 ( .IN1(n7966), .IN2(WX7212), .QN(n11924) );
  INVX0 U12046 ( .INP(n11925), .ZN(n11923) );
  NOR2X0 U12047 ( .IN1(WX7212), .IN2(n7966), .QN(n11925) );
  NAND2X0 U12048 ( .IN1(n9094), .IN2(n11926), .QN(n11913) );
  NAND2X0 U12049 ( .IN1(n991), .IN2(n9280), .QN(n11912) );
  NOR2X0 U12050 ( .IN1(n9236), .IN2(n8926), .QN(n991) );
  NAND2X0 U12051 ( .IN1(n9296), .IN2(CRC_OUT_5_12), .QN(n11911) );
  NAND4X0 U12052 ( .IN1(n11927), .IN2(n11928), .IN3(n11929), .IN4(n11930), 
        .QN(WX5852) );
  NAND2X0 U12053 ( .IN1(n9323), .IN2(n10987), .QN(n11930) );
  NAND2X0 U12054 ( .IN1(n11931), .IN2(n11932), .QN(n10987) );
  INVX0 U12055 ( .INP(n11933), .ZN(n11932) );
  NOR2X0 U12056 ( .IN1(n11934), .IN2(n11935), .QN(n11933) );
  NAND2X0 U12057 ( .IN1(n11935), .IN2(n11934), .QN(n11931) );
  NOR2X0 U12058 ( .IN1(n11936), .IN2(n11937), .QN(n11934) );
  NOR2X0 U12059 ( .IN1(WX7338), .IN2(n7969), .QN(n11937) );
  INVX0 U12060 ( .INP(n11938), .ZN(n11936) );
  NAND2X0 U12061 ( .IN1(n7969), .IN2(WX7338), .QN(n11938) );
  NAND2X0 U12062 ( .IN1(n11939), .IN2(n11940), .QN(n11935) );
  NAND2X0 U12063 ( .IN1(n7968), .IN2(WX7210), .QN(n11940) );
  INVX0 U12064 ( .INP(n11941), .ZN(n11939) );
  NOR2X0 U12065 ( .IN1(WX7210), .IN2(n7968), .QN(n11941) );
  NAND2X0 U12066 ( .IN1(n9094), .IN2(n11942), .QN(n11929) );
  NAND2X0 U12067 ( .IN1(n990), .IN2(n9280), .QN(n11928) );
  NOR2X0 U12068 ( .IN1(n9236), .IN2(n8927), .QN(n990) );
  NAND2X0 U12069 ( .IN1(n9291), .IN2(CRC_OUT_5_13), .QN(n11927) );
  NAND4X0 U12070 ( .IN1(n11943), .IN2(n11944), .IN3(n11945), .IN4(n11946), 
        .QN(WX5850) );
  NAND2X0 U12071 ( .IN1(n9322), .IN2(n11003), .QN(n11946) );
  NAND2X0 U12072 ( .IN1(n11947), .IN2(n11948), .QN(n11003) );
  INVX0 U12073 ( .INP(n11949), .ZN(n11948) );
  NOR2X0 U12074 ( .IN1(n11950), .IN2(n11951), .QN(n11949) );
  NAND2X0 U12075 ( .IN1(n11951), .IN2(n11950), .QN(n11947) );
  NOR2X0 U12076 ( .IN1(n11952), .IN2(n11953), .QN(n11950) );
  NOR2X0 U12077 ( .IN1(WX7336), .IN2(n7971), .QN(n11953) );
  INVX0 U12078 ( .INP(n11954), .ZN(n11952) );
  NAND2X0 U12079 ( .IN1(n7971), .IN2(WX7336), .QN(n11954) );
  NAND2X0 U12080 ( .IN1(n11955), .IN2(n11956), .QN(n11951) );
  NAND2X0 U12081 ( .IN1(n7970), .IN2(WX7208), .QN(n11956) );
  INVX0 U12082 ( .INP(n11957), .ZN(n11955) );
  NOR2X0 U12083 ( .IN1(WX7208), .IN2(n7970), .QN(n11957) );
  NAND2X0 U12084 ( .IN1(n9094), .IN2(n11958), .QN(n11945) );
  NAND2X0 U12085 ( .IN1(n989), .IN2(n9280), .QN(n11944) );
  NOR2X0 U12086 ( .IN1(n9236), .IN2(n8928), .QN(n989) );
  NAND2X0 U12087 ( .IN1(n9291), .IN2(CRC_OUT_5_14), .QN(n11943) );
  NAND4X0 U12088 ( .IN1(n11959), .IN2(n11960), .IN3(n11961), .IN4(n11962), 
        .QN(WX5848) );
  NAND2X0 U12089 ( .IN1(n9323), .IN2(n11016), .QN(n11962) );
  NAND2X0 U12090 ( .IN1(n11963), .IN2(n11964), .QN(n11016) );
  INVX0 U12091 ( .INP(n11965), .ZN(n11964) );
  NOR2X0 U12092 ( .IN1(n11966), .IN2(n11967), .QN(n11965) );
  NAND2X0 U12093 ( .IN1(n11967), .IN2(n11966), .QN(n11963) );
  NOR2X0 U12094 ( .IN1(n11968), .IN2(n11969), .QN(n11966) );
  NOR2X0 U12095 ( .IN1(WX7334), .IN2(n7973), .QN(n11969) );
  INVX0 U12096 ( .INP(n11970), .ZN(n11968) );
  NAND2X0 U12097 ( .IN1(n7973), .IN2(WX7334), .QN(n11970) );
  NAND2X0 U12098 ( .IN1(n11971), .IN2(n11972), .QN(n11967) );
  NAND2X0 U12099 ( .IN1(n7972), .IN2(WX7206), .QN(n11972) );
  INVX0 U12100 ( .INP(n11973), .ZN(n11971) );
  NOR2X0 U12101 ( .IN1(WX7206), .IN2(n7972), .QN(n11973) );
  NAND2X0 U12102 ( .IN1(n9094), .IN2(n11974), .QN(n11961) );
  NAND2X0 U12103 ( .IN1(n988), .IN2(n9280), .QN(n11960) );
  NOR2X0 U12104 ( .IN1(n9236), .IN2(n8929), .QN(n988) );
  NAND2X0 U12105 ( .IN1(n9291), .IN2(CRC_OUT_5_15), .QN(n11959) );
  NAND4X0 U12106 ( .IN1(n11975), .IN2(n11976), .IN3(n11977), .IN4(n11978), 
        .QN(WX5846) );
  NAND2X0 U12107 ( .IN1(n11979), .IN2(n11036), .QN(n11978) );
  NAND2X0 U12108 ( .IN1(n11980), .IN2(n11039), .QN(n11036) );
  NAND2X0 U12109 ( .IN1(n11981), .IN2(n11982), .QN(n11980) );
  NAND2X0 U12110 ( .IN1(n16101), .IN2(n9118), .QN(n11982) );
  NAND2X0 U12111 ( .IN1(TM1), .IN2(n8421), .QN(n11981) );
  NAND3X0 U12112 ( .IN1(n11983), .IN2(n11984), .IN3(n11985), .QN(n11979) );
  NAND2X0 U12113 ( .IN1(n9322), .IN2(n11039), .QN(n11985) );
  NAND2X0 U12114 ( .IN1(n11986), .IN2(n11987), .QN(n11039) );
  NAND2X0 U12115 ( .IN1(n7711), .IN2(n11988), .QN(n11987) );
  INVX0 U12116 ( .INP(n11989), .ZN(n11986) );
  NOR2X0 U12117 ( .IN1(n11988), .IN2(n7711), .QN(n11989) );
  NOR2X0 U12118 ( .IN1(n11990), .IN2(n11991), .QN(n11988) );
  NOR2X0 U12119 ( .IN1(WX7332), .IN2(n7712), .QN(n11991) );
  INVX0 U12120 ( .INP(n11992), .ZN(n11990) );
  NAND2X0 U12121 ( .IN1(n7712), .IN2(WX7332), .QN(n11992) );
  NAND2X0 U12122 ( .IN1(n9082), .IN2(n8421), .QN(n11984) );
  NAND2X0 U12123 ( .IN1(n16101), .IN2(n9078), .QN(n11983) );
  NAND2X0 U12124 ( .IN1(n11993), .IN2(n9110), .QN(n11977) );
  NAND2X0 U12125 ( .IN1(n987), .IN2(n9280), .QN(n11976) );
  NOR2X0 U12126 ( .IN1(n9236), .IN2(n8930), .QN(n987) );
  NAND2X0 U12127 ( .IN1(n9291), .IN2(CRC_OUT_5_16), .QN(n11975) );
  NAND4X0 U12128 ( .IN1(n11994), .IN2(n11995), .IN3(n11996), .IN4(n11997), 
        .QN(WX5844) );
  NAND2X0 U12129 ( .IN1(n11998), .IN2(n11059), .QN(n11997) );
  NAND2X0 U12130 ( .IN1(n11999), .IN2(n11062), .QN(n11059) );
  NAND2X0 U12131 ( .IN1(n12000), .IN2(n12001), .QN(n11999) );
  NAND2X0 U12132 ( .IN1(n16100), .IN2(n9118), .QN(n12001) );
  NAND2X0 U12133 ( .IN1(TM1), .IN2(n8422), .QN(n12000) );
  NAND3X0 U12134 ( .IN1(n12002), .IN2(n12003), .IN3(n12004), .QN(n11998) );
  NAND2X0 U12135 ( .IN1(n9323), .IN2(n11062), .QN(n12004) );
  NAND2X0 U12136 ( .IN1(n12005), .IN2(n12006), .QN(n11062) );
  NAND2X0 U12137 ( .IN1(n7713), .IN2(n12007), .QN(n12006) );
  INVX0 U12138 ( .INP(n12008), .ZN(n12005) );
  NOR2X0 U12139 ( .IN1(n12007), .IN2(n7713), .QN(n12008) );
  NOR2X0 U12140 ( .IN1(n12009), .IN2(n12010), .QN(n12007) );
  NOR2X0 U12141 ( .IN1(WX7330), .IN2(n7714), .QN(n12010) );
  INVX0 U12142 ( .INP(n12011), .ZN(n12009) );
  NAND2X0 U12143 ( .IN1(n7714), .IN2(WX7330), .QN(n12011) );
  NAND2X0 U12144 ( .IN1(n9081), .IN2(n8422), .QN(n12003) );
  NAND2X0 U12145 ( .IN1(n16100), .IN2(n9077), .QN(n12002) );
  NAND2X0 U12146 ( .IN1(n12012), .IN2(n12013), .QN(n11996) );
  NAND2X0 U12147 ( .IN1(n12014), .IN2(n12015), .QN(n12012) );
  NAND2X0 U12148 ( .IN1(n9095), .IN2(n12016), .QN(n12015) );
  NAND2X0 U12149 ( .IN1(n9095), .IN2(n8480), .QN(n12014) );
  NAND2X0 U12150 ( .IN1(n986), .IN2(n9280), .QN(n11995) );
  NOR2X0 U12151 ( .IN1(n9236), .IN2(n8931), .QN(n986) );
  NAND2X0 U12152 ( .IN1(test_so54), .IN2(n9314), .QN(n11994) );
  NAND4X0 U12153 ( .IN1(n12017), .IN2(n12018), .IN3(n12019), .IN4(n12020), 
        .QN(WX5842) );
  NAND2X0 U12154 ( .IN1(n12021), .IN2(n11082), .QN(n12020) );
  NAND2X0 U12155 ( .IN1(n12022), .IN2(n11085), .QN(n11082) );
  NAND2X0 U12156 ( .IN1(n12023), .IN2(n12024), .QN(n12022) );
  NAND2X0 U12157 ( .IN1(n16099), .IN2(n9118), .QN(n12024) );
  NAND2X0 U12158 ( .IN1(TM1), .IN2(n8423), .QN(n12023) );
  NAND3X0 U12159 ( .IN1(n12025), .IN2(n12026), .IN3(n12027), .QN(n12021) );
  NAND2X0 U12160 ( .IN1(n9322), .IN2(n11085), .QN(n12027) );
  NAND2X0 U12161 ( .IN1(n12028), .IN2(n12029), .QN(n11085) );
  NAND2X0 U12162 ( .IN1(n7715), .IN2(n12030), .QN(n12029) );
  INVX0 U12163 ( .INP(n12031), .ZN(n12028) );
  NOR2X0 U12164 ( .IN1(n12030), .IN2(n7715), .QN(n12031) );
  NOR2X0 U12165 ( .IN1(n12032), .IN2(n12033), .QN(n12030) );
  NOR2X0 U12166 ( .IN1(WX7328), .IN2(n7716), .QN(n12033) );
  INVX0 U12167 ( .INP(n12034), .ZN(n12032) );
  NAND2X0 U12168 ( .IN1(n7716), .IN2(WX7328), .QN(n12034) );
  NAND2X0 U12169 ( .IN1(n9790), .IN2(n8423), .QN(n12026) );
  NAND2X0 U12170 ( .IN1(n16099), .IN2(n9791), .QN(n12025) );
  NAND2X0 U12171 ( .IN1(n12035), .IN2(n9111), .QN(n12019) );
  NAND2X0 U12172 ( .IN1(n985), .IN2(n9280), .QN(n12018) );
  NOR2X0 U12173 ( .IN1(n9236), .IN2(n8932), .QN(n985) );
  NAND2X0 U12174 ( .IN1(n9291), .IN2(CRC_OUT_5_18), .QN(n12017) );
  NAND4X0 U12175 ( .IN1(n12036), .IN2(n12037), .IN3(n12038), .IN4(n12039), 
        .QN(WX5840) );
  NAND2X0 U12176 ( .IN1(n12040), .IN2(n11105), .QN(n12039) );
  NAND2X0 U12177 ( .IN1(n12041), .IN2(n11108), .QN(n11105) );
  NAND2X0 U12178 ( .IN1(n12042), .IN2(n12043), .QN(n12041) );
  NAND2X0 U12179 ( .IN1(n16098), .IN2(n9118), .QN(n12043) );
  NAND2X0 U12180 ( .IN1(TM1), .IN2(n8424), .QN(n12042) );
  NAND3X0 U12181 ( .IN1(n12044), .IN2(n12045), .IN3(n12046), .QN(n12040) );
  NAND2X0 U12182 ( .IN1(n9322), .IN2(n11108), .QN(n12046) );
  NAND2X0 U12183 ( .IN1(n12047), .IN2(n12048), .QN(n11108) );
  NAND2X0 U12184 ( .IN1(n7717), .IN2(n12049), .QN(n12048) );
  INVX0 U12185 ( .INP(n12050), .ZN(n12047) );
  NOR2X0 U12186 ( .IN1(n12049), .IN2(n7717), .QN(n12050) );
  NOR2X0 U12187 ( .IN1(n12051), .IN2(n12052), .QN(n12049) );
  NOR2X0 U12188 ( .IN1(WX7326), .IN2(n7718), .QN(n12052) );
  INVX0 U12189 ( .INP(n12053), .ZN(n12051) );
  NAND2X0 U12190 ( .IN1(n7718), .IN2(WX7326), .QN(n12053) );
  NAND2X0 U12191 ( .IN1(n9083), .IN2(n8424), .QN(n12045) );
  NAND2X0 U12192 ( .IN1(n16098), .IN2(n9079), .QN(n12044) );
  NAND2X0 U12193 ( .IN1(n12054), .IN2(n12055), .QN(n12038) );
  NAND2X0 U12194 ( .IN1(n12056), .IN2(n12057), .QN(n12054) );
  NAND2X0 U12195 ( .IN1(n9095), .IN2(n12058), .QN(n12057) );
  NAND2X0 U12196 ( .IN1(n9095), .IN2(n8482), .QN(n12056) );
  NAND2X0 U12197 ( .IN1(n984), .IN2(n9280), .QN(n12037) );
  NOR2X0 U12198 ( .IN1(n9236), .IN2(n8933), .QN(n984) );
  NAND2X0 U12199 ( .IN1(n9291), .IN2(CRC_OUT_5_19), .QN(n12036) );
  NAND4X0 U12200 ( .IN1(n12059), .IN2(n12060), .IN3(n12061), .IN4(n12062), 
        .QN(WX5838) );
  NAND2X0 U12201 ( .IN1(n12063), .IN2(n11128), .QN(n12062) );
  NAND2X0 U12202 ( .IN1(n12064), .IN2(n11131), .QN(n11128) );
  NAND2X0 U12203 ( .IN1(n12065), .IN2(n12066), .QN(n12064) );
  NAND2X0 U12204 ( .IN1(n16097), .IN2(n9118), .QN(n12066) );
  NAND2X0 U12205 ( .IN1(TM1), .IN2(n8425), .QN(n12065) );
  NAND3X0 U12206 ( .IN1(n12067), .IN2(n12068), .IN3(n12069), .QN(n12063) );
  NAND2X0 U12207 ( .IN1(n9323), .IN2(n11131), .QN(n12069) );
  NAND2X0 U12208 ( .IN1(n12070), .IN2(n12071), .QN(n11131) );
  NAND2X0 U12209 ( .IN1(n7719), .IN2(n12072), .QN(n12071) );
  INVX0 U12210 ( .INP(n12073), .ZN(n12070) );
  NOR2X0 U12211 ( .IN1(n12072), .IN2(n7719), .QN(n12073) );
  NOR2X0 U12212 ( .IN1(n12074), .IN2(n12075), .QN(n12072) );
  NOR2X0 U12213 ( .IN1(WX7324), .IN2(n7720), .QN(n12075) );
  INVX0 U12214 ( .INP(n12076), .ZN(n12074) );
  NAND2X0 U12215 ( .IN1(n7720), .IN2(WX7324), .QN(n12076) );
  NAND2X0 U12216 ( .IN1(n9082), .IN2(n8425), .QN(n12068) );
  NAND2X0 U12217 ( .IN1(n16097), .IN2(n9078), .QN(n12067) );
  NAND2X0 U12218 ( .IN1(n12077), .IN2(n9111), .QN(n12061) );
  NAND2X0 U12219 ( .IN1(n983), .IN2(n9280), .QN(n12060) );
  NOR2X0 U12220 ( .IN1(n9236), .IN2(n8934), .QN(n983) );
  NAND2X0 U12221 ( .IN1(n9291), .IN2(CRC_OUT_5_20), .QN(n12059) );
  NAND4X0 U12222 ( .IN1(n12078), .IN2(n12079), .IN3(n12080), .IN4(n12081), 
        .QN(WX5836) );
  NAND2X0 U12223 ( .IN1(n12082), .IN2(n12083), .QN(n12081) );
  NAND2X0 U12224 ( .IN1(n12084), .IN2(n12085), .QN(n12082) );
  NAND2X0 U12225 ( .IN1(n9095), .IN2(n12086), .QN(n12085) );
  NAND2X0 U12226 ( .IN1(n9095), .IN2(n8484), .QN(n12084) );
  NAND2X0 U12227 ( .IN1(n11150), .IN2(n9335), .QN(n12080) );
  NOR2X0 U12228 ( .IN1(n12087), .IN2(n12088), .QN(n11150) );
  INVX0 U12229 ( .INP(n12089), .ZN(n12088) );
  NAND2X0 U12230 ( .IN1(n12090), .IN2(n12091), .QN(n12089) );
  NOR2X0 U12231 ( .IN1(n12091), .IN2(n12090), .QN(n12087) );
  NAND2X0 U12232 ( .IN1(n12092), .IN2(n12093), .QN(n12090) );
  NAND2X0 U12233 ( .IN1(n12094), .IN2(WX7258), .QN(n12093) );
  NAND2X0 U12234 ( .IN1(n12095), .IN2(n12096), .QN(n12094) );
  NAND3X0 U12235 ( .IN1(n12095), .IN2(n12096), .IN3(n7722), .QN(n12092) );
  NAND2X0 U12236 ( .IN1(test_so63), .IN2(WX7194), .QN(n12096) );
  NAND2X0 U12237 ( .IN1(n7721), .IN2(n8799), .QN(n12095) );
  NOR2X0 U12238 ( .IN1(n12097), .IN2(n12098), .QN(n12091) );
  INVX0 U12239 ( .INP(n12099), .ZN(n12098) );
  NAND2X0 U12240 ( .IN1(n16096), .IN2(n9118), .QN(n12099) );
  NOR2X0 U12241 ( .IN1(n9116), .IN2(n16096), .QN(n12097) );
  NAND2X0 U12242 ( .IN1(n982), .IN2(n9280), .QN(n12079) );
  NOR2X0 U12243 ( .IN1(n9236), .IN2(n8935), .QN(n982) );
  NAND2X0 U12244 ( .IN1(n9291), .IN2(CRC_OUT_5_21), .QN(n12078) );
  NAND4X0 U12245 ( .IN1(n12100), .IN2(n12101), .IN3(n12102), .IN4(n12103), 
        .QN(WX5834) );
  NAND2X0 U12246 ( .IN1(n12104), .IN2(n11170), .QN(n12103) );
  NAND2X0 U12247 ( .IN1(n12105), .IN2(n11173), .QN(n11170) );
  NAND2X0 U12248 ( .IN1(n12106), .IN2(n12107), .QN(n12105) );
  NAND2X0 U12249 ( .IN1(n16095), .IN2(n9118), .QN(n12107) );
  NAND2X0 U12250 ( .IN1(TM1), .IN2(n8427), .QN(n12106) );
  NAND3X0 U12251 ( .IN1(n12108), .IN2(n12109), .IN3(n12110), .QN(n12104) );
  NAND2X0 U12252 ( .IN1(n9322), .IN2(n11173), .QN(n12110) );
  NAND2X0 U12253 ( .IN1(n12111), .IN2(n12112), .QN(n11173) );
  NAND2X0 U12254 ( .IN1(n7723), .IN2(n12113), .QN(n12112) );
  INVX0 U12255 ( .INP(n12114), .ZN(n12111) );
  NOR2X0 U12256 ( .IN1(n12113), .IN2(n7723), .QN(n12114) );
  NOR2X0 U12257 ( .IN1(n12115), .IN2(n12116), .QN(n12113) );
  NOR2X0 U12258 ( .IN1(WX7320), .IN2(n7724), .QN(n12116) );
  INVX0 U12259 ( .INP(n12117), .ZN(n12115) );
  NAND2X0 U12260 ( .IN1(n7724), .IN2(WX7320), .QN(n12117) );
  NAND2X0 U12261 ( .IN1(n9081), .IN2(n8427), .QN(n12109) );
  NAND2X0 U12262 ( .IN1(n16095), .IN2(n9077), .QN(n12108) );
  NAND2X0 U12263 ( .IN1(n12118), .IN2(n12119), .QN(n12102) );
  NAND2X0 U12264 ( .IN1(n12120), .IN2(n12121), .QN(n12118) );
  NAND2X0 U12265 ( .IN1(n9095), .IN2(n12122), .QN(n12121) );
  NAND2X0 U12266 ( .IN1(n8256), .IN2(n9111), .QN(n12120) );
  NAND2X0 U12267 ( .IN1(n981), .IN2(n9280), .QN(n12101) );
  NOR2X0 U12268 ( .IN1(n9236), .IN2(n8936), .QN(n981) );
  NAND2X0 U12269 ( .IN1(n9291), .IN2(CRC_OUT_5_22), .QN(n12100) );
  NAND4X0 U12270 ( .IN1(n12123), .IN2(n12124), .IN3(n12125), .IN4(n12126), 
        .QN(WX5832) );
  NAND2X0 U12271 ( .IN1(n12127), .IN2(n12128), .QN(n12126) );
  NAND2X0 U12272 ( .IN1(n12129), .IN2(n12130), .QN(n12127) );
  NAND2X0 U12273 ( .IN1(n9095), .IN2(n12131), .QN(n12130) );
  NAND2X0 U12274 ( .IN1(n9095), .IN2(n8487), .QN(n12129) );
  NAND2X0 U12275 ( .IN1(n11192), .IN2(n9335), .QN(n12125) );
  NOR2X0 U12276 ( .IN1(n12132), .IN2(n12133), .QN(n11192) );
  INVX0 U12277 ( .INP(n12134), .ZN(n12133) );
  NAND2X0 U12278 ( .IN1(n12135), .IN2(n12136), .QN(n12134) );
  NOR2X0 U12279 ( .IN1(n12136), .IN2(n12135), .QN(n12132) );
  NAND2X0 U12280 ( .IN1(n12137), .IN2(n12138), .QN(n12135) );
  NAND2X0 U12281 ( .IN1(n8219), .IN2(n12139), .QN(n12138) );
  INVX0 U12282 ( .INP(n12140), .ZN(n12139) );
  NAND2X0 U12283 ( .IN1(n12140), .IN2(WX7318), .QN(n12137) );
  NAND2X0 U12284 ( .IN1(n12141), .IN2(n12142), .QN(n12140) );
  INVX0 U12285 ( .INP(n12143), .ZN(n12142) );
  NOR2X0 U12286 ( .IN1(n8809), .IN2(n16094), .QN(n12143) );
  NAND2X0 U12287 ( .IN1(n16094), .IN2(n8809), .QN(n12141) );
  NOR2X0 U12288 ( .IN1(n12144), .IN2(n12145), .QN(n12136) );
  INVX0 U12289 ( .INP(n12146), .ZN(n12145) );
  NAND2X0 U12290 ( .IN1(n7725), .IN2(n9118), .QN(n12146) );
  NOR2X0 U12291 ( .IN1(n9116), .IN2(n7725), .QN(n12144) );
  NAND2X0 U12292 ( .IN1(n980), .IN2(n9280), .QN(n12124) );
  NOR2X0 U12293 ( .IN1(n9235), .IN2(n8937), .QN(n980) );
  NAND2X0 U12294 ( .IN1(n9291), .IN2(CRC_OUT_5_23), .QN(n12123) );
  NAND4X0 U12295 ( .IN1(n12147), .IN2(n12148), .IN3(n12149), .IN4(n12150), 
        .QN(WX5830) );
  NAND2X0 U12296 ( .IN1(n12151), .IN2(n11212), .QN(n12150) );
  NAND2X0 U12297 ( .IN1(n12152), .IN2(n11215), .QN(n11212) );
  NAND2X0 U12298 ( .IN1(n12153), .IN2(n12154), .QN(n12152) );
  NAND2X0 U12299 ( .IN1(n16093), .IN2(n9118), .QN(n12154) );
  NAND2X0 U12300 ( .IN1(TM1), .IN2(n8429), .QN(n12153) );
  NAND3X0 U12301 ( .IN1(n12155), .IN2(n12156), .IN3(n12157), .QN(n12151) );
  NAND2X0 U12302 ( .IN1(n9322), .IN2(n11215), .QN(n12157) );
  NAND2X0 U12303 ( .IN1(n12158), .IN2(n12159), .QN(n11215) );
  NAND2X0 U12304 ( .IN1(n7726), .IN2(n12160), .QN(n12159) );
  INVX0 U12305 ( .INP(n12161), .ZN(n12158) );
  NOR2X0 U12306 ( .IN1(n12160), .IN2(n7726), .QN(n12161) );
  NOR2X0 U12307 ( .IN1(n12162), .IN2(n12163), .QN(n12160) );
  NOR2X0 U12308 ( .IN1(WX7316), .IN2(n7727), .QN(n12163) );
  INVX0 U12309 ( .INP(n12164), .ZN(n12162) );
  NAND2X0 U12310 ( .IN1(n7727), .IN2(WX7316), .QN(n12164) );
  NAND2X0 U12311 ( .IN1(n9790), .IN2(n8429), .QN(n12156) );
  NAND2X0 U12312 ( .IN1(n16093), .IN2(n9791), .QN(n12155) );
  NAND2X0 U12313 ( .IN1(n12165), .IN2(n12166), .QN(n12149) );
  NAND2X0 U12314 ( .IN1(n12167), .IN2(n12168), .QN(n12165) );
  NAND2X0 U12315 ( .IN1(n9095), .IN2(n12169), .QN(n12168) );
  NAND2X0 U12316 ( .IN1(n9095), .IN2(n8488), .QN(n12167) );
  NAND2X0 U12317 ( .IN1(n979), .IN2(n9280), .QN(n12148) );
  NOR2X0 U12318 ( .IN1(n9067), .IN2(n9162), .QN(n979) );
  NAND2X0 U12319 ( .IN1(n9291), .IN2(CRC_OUT_5_24), .QN(n12147) );
  NAND4X0 U12320 ( .IN1(n12170), .IN2(n12171), .IN3(n12172), .IN4(n12173), 
        .QN(WX5828) );
  NAND2X0 U12321 ( .IN1(n12174), .IN2(n12175), .QN(n12173) );
  NAND2X0 U12322 ( .IN1(n12176), .IN2(n12177), .QN(n12174) );
  NAND2X0 U12323 ( .IN1(n9095), .IN2(n12178), .QN(n12177) );
  NAND2X0 U12324 ( .IN1(n9095), .IN2(n8489), .QN(n12176) );
  NAND2X0 U12325 ( .IN1(n11234), .IN2(n9335), .QN(n12172) );
  NOR2X0 U12326 ( .IN1(n12179), .IN2(n12180), .QN(n11234) );
  INVX0 U12327 ( .INP(n12181), .ZN(n12180) );
  NAND2X0 U12328 ( .IN1(n12182), .IN2(n12183), .QN(n12181) );
  NOR2X0 U12329 ( .IN1(n12183), .IN2(n12182), .QN(n12179) );
  NAND2X0 U12330 ( .IN1(n12184), .IN2(n12185), .QN(n12182) );
  NAND2X0 U12331 ( .IN1(n8217), .IN2(n12186), .QN(n12185) );
  INVX0 U12332 ( .INP(n12187), .ZN(n12186) );
  NAND2X0 U12333 ( .IN1(n12187), .IN2(WX7314), .QN(n12184) );
  NAND2X0 U12334 ( .IN1(n12188), .IN2(n12189), .QN(n12187) );
  INVX0 U12335 ( .INP(n12190), .ZN(n12189) );
  NOR2X0 U12336 ( .IN1(n8810), .IN2(n16092), .QN(n12190) );
  NAND2X0 U12337 ( .IN1(n16092), .IN2(n8810), .QN(n12188) );
  NOR2X0 U12338 ( .IN1(n12191), .IN2(n12192), .QN(n12183) );
  INVX0 U12339 ( .INP(n12193), .ZN(n12192) );
  NAND2X0 U12340 ( .IN1(n7728), .IN2(n9118), .QN(n12193) );
  NOR2X0 U12341 ( .IN1(n9116), .IN2(n7728), .QN(n12191) );
  NAND2X0 U12342 ( .IN1(n978), .IN2(n9280), .QN(n12171) );
  NOR2X0 U12343 ( .IN1(n9235), .IN2(n8938), .QN(n978) );
  NAND2X0 U12344 ( .IN1(n9292), .IN2(CRC_OUT_5_25), .QN(n12170) );
  NAND4X0 U12345 ( .IN1(n12194), .IN2(n12195), .IN3(n12196), .IN4(n12197), 
        .QN(WX5826) );
  NAND2X0 U12346 ( .IN1(n12198), .IN2(n11240), .QN(n12197) );
  NAND2X0 U12347 ( .IN1(n12199), .IN2(n11243), .QN(n11240) );
  NAND2X0 U12348 ( .IN1(n12200), .IN2(n12201), .QN(n12199) );
  NAND2X0 U12349 ( .IN1(n16091), .IN2(n9118), .QN(n12201) );
  NAND2X0 U12350 ( .IN1(TM1), .IN2(n8431), .QN(n12200) );
  NAND3X0 U12351 ( .IN1(n12202), .IN2(n12203), .IN3(n12204), .QN(n12198) );
  NAND2X0 U12352 ( .IN1(n9323), .IN2(n11243), .QN(n12204) );
  NAND2X0 U12353 ( .IN1(n12205), .IN2(n12206), .QN(n11243) );
  NAND2X0 U12354 ( .IN1(n7729), .IN2(n12207), .QN(n12206) );
  INVX0 U12355 ( .INP(n12208), .ZN(n12205) );
  NOR2X0 U12356 ( .IN1(n12207), .IN2(n7729), .QN(n12208) );
  NOR2X0 U12357 ( .IN1(n12209), .IN2(n12210), .QN(n12207) );
  NOR2X0 U12358 ( .IN1(WX7312), .IN2(n7730), .QN(n12210) );
  INVX0 U12359 ( .INP(n12211), .ZN(n12209) );
  NAND2X0 U12360 ( .IN1(n7730), .IN2(WX7312), .QN(n12211) );
  NAND2X0 U12361 ( .IN1(n9083), .IN2(n8431), .QN(n12203) );
  NAND2X0 U12362 ( .IN1(n16091), .IN2(n9079), .QN(n12202) );
  NAND2X0 U12363 ( .IN1(n12212), .IN2(n12213), .QN(n12196) );
  NAND2X0 U12364 ( .IN1(n12214), .IN2(n12215), .QN(n12212) );
  NAND2X0 U12365 ( .IN1(n9108), .IN2(n12216), .QN(n12215) );
  NAND2X0 U12366 ( .IN1(n9105), .IN2(n8490), .QN(n12214) );
  NAND2X0 U12367 ( .IN1(n977), .IN2(n9280), .QN(n12195) );
  NOR2X0 U12368 ( .IN1(n9235), .IN2(n8939), .QN(n977) );
  NAND2X0 U12369 ( .IN1(n9292), .IN2(CRC_OUT_5_26), .QN(n12194) );
  NAND4X0 U12370 ( .IN1(n12217), .IN2(n12218), .IN3(n12219), .IN4(n12220), 
        .QN(WX5824) );
  NAND2X0 U12371 ( .IN1(n12221), .IN2(n11276), .QN(n12220) );
  NAND3X0 U12372 ( .IN1(n12222), .IN2(n12223), .IN3(n11279), .QN(n11276) );
  NAND2X0 U12373 ( .IN1(n8215), .IN2(n9118), .QN(n12223) );
  NAND2X0 U12374 ( .IN1(TM1), .IN2(WX7310), .QN(n12222) );
  NAND3X0 U12375 ( .IN1(n12224), .IN2(n12225), .IN3(n12226), .QN(n12221) );
  NAND2X0 U12376 ( .IN1(n9323), .IN2(n11279), .QN(n12226) );
  NAND2X0 U12377 ( .IN1(n12227), .IN2(n12228), .QN(n11279) );
  NAND2X0 U12378 ( .IN1(n12229), .IN2(WX7246), .QN(n12228) );
  NAND2X0 U12379 ( .IN1(n12230), .IN2(n12231), .QN(n12229) );
  NAND3X0 U12380 ( .IN1(n12230), .IN2(n12231), .IN3(n7732), .QN(n12227) );
  NAND2X0 U12381 ( .IN1(test_so57), .IN2(WX7182), .QN(n12231) );
  NAND2X0 U12382 ( .IN1(n7731), .IN2(n8820), .QN(n12230) );
  NAND2X0 U12383 ( .IN1(n9077), .IN2(WX7310), .QN(n12225) );
  NAND2X0 U12384 ( .IN1(n9082), .IN2(n8215), .QN(n12224) );
  NAND2X0 U12385 ( .IN1(n12232), .IN2(n12233), .QN(n12219) );
  NAND2X0 U12386 ( .IN1(n12234), .IN2(n12235), .QN(n12232) );
  NAND2X0 U12387 ( .IN1(n9105), .IN2(n12236), .QN(n12235) );
  NAND2X0 U12388 ( .IN1(n9105), .IN2(n8491), .QN(n12234) );
  NAND2X0 U12389 ( .IN1(n976), .IN2(n9280), .QN(n12218) );
  NOR2X0 U12390 ( .IN1(n9235), .IN2(n8940), .QN(n976) );
  NAND2X0 U12391 ( .IN1(n9292), .IN2(CRC_OUT_5_27), .QN(n12217) );
  NAND4X0 U12392 ( .IN1(n12237), .IN2(n12238), .IN3(n12239), .IN4(n12240), 
        .QN(WX5822) );
  NAND2X0 U12393 ( .IN1(n12241), .IN2(n11285), .QN(n12240) );
  NAND2X0 U12394 ( .IN1(n12242), .IN2(n11288), .QN(n11285) );
  NAND2X0 U12395 ( .IN1(n12243), .IN2(n12244), .QN(n12242) );
  NAND2X0 U12396 ( .IN1(n16090), .IN2(n9118), .QN(n12244) );
  NAND2X0 U12397 ( .IN1(TM1), .IN2(n8434), .QN(n12243) );
  NAND3X0 U12398 ( .IN1(n12245), .IN2(n12246), .IN3(n12247), .QN(n12241) );
  NAND2X0 U12399 ( .IN1(n9323), .IN2(n11288), .QN(n12247) );
  NAND2X0 U12400 ( .IN1(n12248), .IN2(n12249), .QN(n11288) );
  NAND2X0 U12401 ( .IN1(n7733), .IN2(n12250), .QN(n12249) );
  INVX0 U12402 ( .INP(n12251), .ZN(n12248) );
  NOR2X0 U12403 ( .IN1(n12250), .IN2(n7733), .QN(n12251) );
  NOR2X0 U12404 ( .IN1(n12252), .IN2(n12253), .QN(n12250) );
  NOR2X0 U12405 ( .IN1(WX7308), .IN2(n7734), .QN(n12253) );
  INVX0 U12406 ( .INP(n12254), .ZN(n12252) );
  NAND2X0 U12407 ( .IN1(n7734), .IN2(WX7308), .QN(n12254) );
  NAND2X0 U12408 ( .IN1(n9081), .IN2(n8434), .QN(n12246) );
  NAND2X0 U12409 ( .IN1(n16090), .IN2(n9078), .QN(n12245) );
  NAND2X0 U12410 ( .IN1(n12255), .IN2(n12256), .QN(n12239) );
  NAND2X0 U12411 ( .IN1(n12257), .IN2(n12258), .QN(n12255) );
  NAND2X0 U12412 ( .IN1(n9105), .IN2(n12259), .QN(n12258) );
  NAND2X0 U12413 ( .IN1(n9105), .IN2(n8492), .QN(n12257) );
  NAND2X0 U12414 ( .IN1(n975), .IN2(n9281), .QN(n12238) );
  NOR2X0 U12415 ( .IN1(n9235), .IN2(n8941), .QN(n975) );
  NAND2X0 U12416 ( .IN1(n9292), .IN2(CRC_OUT_5_28), .QN(n12237) );
  NAND4X0 U12417 ( .IN1(n12260), .IN2(n12261), .IN3(n12262), .IN4(n12263), 
        .QN(WX5820) );
  NAND2X0 U12418 ( .IN1(n12264), .IN2(n11323), .QN(n12263) );
  NAND2X0 U12419 ( .IN1(n12265), .IN2(n11326), .QN(n11323) );
  NAND2X0 U12420 ( .IN1(n12266), .IN2(n12267), .QN(n12265) );
  NAND2X0 U12421 ( .IN1(n16089), .IN2(n9118), .QN(n12267) );
  NAND2X0 U12422 ( .IN1(TM1), .IN2(n8435), .QN(n12266) );
  NAND3X0 U12423 ( .IN1(n12268), .IN2(n12269), .IN3(n12270), .QN(n12264) );
  NAND2X0 U12424 ( .IN1(n9323), .IN2(n11326), .QN(n12270) );
  NAND2X0 U12425 ( .IN1(n12271), .IN2(n12272), .QN(n11326) );
  NAND2X0 U12426 ( .IN1(n7735), .IN2(n12273), .QN(n12272) );
  INVX0 U12427 ( .INP(n12274), .ZN(n12271) );
  NOR2X0 U12428 ( .IN1(n12273), .IN2(n7735), .QN(n12274) );
  NOR2X0 U12429 ( .IN1(n12275), .IN2(n12276), .QN(n12273) );
  NOR2X0 U12430 ( .IN1(WX7306), .IN2(n7736), .QN(n12276) );
  INVX0 U12431 ( .INP(n12277), .ZN(n12275) );
  NAND2X0 U12432 ( .IN1(n7736), .IN2(WX7306), .QN(n12277) );
  NAND2X0 U12433 ( .IN1(n9790), .IN2(n8435), .QN(n12269) );
  NAND2X0 U12434 ( .IN1(n16089), .IN2(n9077), .QN(n12268) );
  NAND2X0 U12435 ( .IN1(n12278), .IN2(n12279), .QN(n12262) );
  NAND2X0 U12436 ( .IN1(n12280), .IN2(n12281), .QN(n12278) );
  NAND2X0 U12437 ( .IN1(n9105), .IN2(n12282), .QN(n12281) );
  NAND2X0 U12438 ( .IN1(n9106), .IN2(n8493), .QN(n12280) );
  NAND2X0 U12439 ( .IN1(n974), .IN2(n9281), .QN(n12261) );
  NOR2X0 U12440 ( .IN1(n9235), .IN2(n8942), .QN(n974) );
  NAND2X0 U12441 ( .IN1(n9292), .IN2(CRC_OUT_5_29), .QN(n12260) );
  NAND4X0 U12442 ( .IN1(n12283), .IN2(n12284), .IN3(n12285), .IN4(n12286), 
        .QN(WX5818) );
  NAND2X0 U12443 ( .IN1(n12287), .IN2(n11332), .QN(n12286) );
  NAND2X0 U12444 ( .IN1(n12288), .IN2(n11335), .QN(n11332) );
  NAND2X0 U12445 ( .IN1(n12289), .IN2(n12290), .QN(n12288) );
  NAND2X0 U12446 ( .IN1(n16088), .IN2(n9117), .QN(n12290) );
  NAND2X0 U12447 ( .IN1(TM1), .IN2(n8436), .QN(n12289) );
  NAND3X0 U12448 ( .IN1(n12291), .IN2(n12292), .IN3(n12293), .QN(n12287) );
  NAND2X0 U12449 ( .IN1(n9323), .IN2(n11335), .QN(n12293) );
  NAND2X0 U12450 ( .IN1(n12294), .IN2(n12295), .QN(n11335) );
  NAND2X0 U12451 ( .IN1(n7737), .IN2(n12296), .QN(n12295) );
  INVX0 U12452 ( .INP(n12297), .ZN(n12294) );
  NOR2X0 U12453 ( .IN1(n12296), .IN2(n7737), .QN(n12297) );
  NOR2X0 U12454 ( .IN1(n12298), .IN2(n12299), .QN(n12296) );
  NOR2X0 U12455 ( .IN1(WX7304), .IN2(n7738), .QN(n12299) );
  INVX0 U12456 ( .INP(n12300), .ZN(n12298) );
  NAND2X0 U12457 ( .IN1(n7738), .IN2(WX7304), .QN(n12300) );
  NAND2X0 U12458 ( .IN1(n9083), .IN2(n8436), .QN(n12292) );
  NAND2X0 U12459 ( .IN1(n16088), .IN2(n9791), .QN(n12291) );
  NAND2X0 U12460 ( .IN1(n12301), .IN2(n12302), .QN(n12285) );
  NAND2X0 U12461 ( .IN1(n12303), .IN2(n12304), .QN(n12301) );
  NAND2X0 U12462 ( .IN1(n9106), .IN2(n12305), .QN(n12304) );
  NAND2X0 U12463 ( .IN1(n9106), .IN2(n8494), .QN(n12303) );
  NAND2X0 U12464 ( .IN1(n973), .IN2(n9281), .QN(n12284) );
  NOR2X0 U12465 ( .IN1(n9235), .IN2(n8943), .QN(n973) );
  NAND2X0 U12466 ( .IN1(n9292), .IN2(CRC_OUT_5_30), .QN(n12283) );
  NAND4X0 U12467 ( .IN1(n12306), .IN2(n12307), .IN3(n12308), .IN4(n12309), 
        .QN(WX5816) );
  NAND2X0 U12468 ( .IN1(n12310), .IN2(n11370), .QN(n12309) );
  NAND2X0 U12469 ( .IN1(n12311), .IN2(n11373), .QN(n11370) );
  NAND2X0 U12470 ( .IN1(n12312), .IN2(n12313), .QN(n12311) );
  NAND2X0 U12471 ( .IN1(n16087), .IN2(n9117), .QN(n12313) );
  NAND2X0 U12472 ( .IN1(TM1), .IN2(n8437), .QN(n12312) );
  NAND3X0 U12473 ( .IN1(n12314), .IN2(n12315), .IN3(n12316), .QN(n12310) );
  NAND2X0 U12474 ( .IN1(n9323), .IN2(n11373), .QN(n12316) );
  NAND2X0 U12475 ( .IN1(n12317), .IN2(n12318), .QN(n11373) );
  NAND2X0 U12476 ( .IN1(n7617), .IN2(n12319), .QN(n12318) );
  INVX0 U12477 ( .INP(n12320), .ZN(n12317) );
  NOR2X0 U12478 ( .IN1(n12319), .IN2(n7617), .QN(n12320) );
  NOR2X0 U12479 ( .IN1(n12321), .IN2(n12322), .QN(n12319) );
  NOR2X0 U12480 ( .IN1(WX7302), .IN2(n7618), .QN(n12322) );
  INVX0 U12481 ( .INP(n12323), .ZN(n12321) );
  NAND2X0 U12482 ( .IN1(n7618), .IN2(WX7302), .QN(n12323) );
  NAND2X0 U12483 ( .IN1(n9082), .IN2(n8437), .QN(n12315) );
  NAND2X0 U12484 ( .IN1(n16087), .IN2(n9079), .QN(n12314) );
  NAND2X0 U12485 ( .IN1(n12324), .IN2(n12325), .QN(n12308) );
  NAND2X0 U12486 ( .IN1(n12326), .IN2(n12327), .QN(n12324) );
  NAND2X0 U12487 ( .IN1(n9106), .IN2(n12328), .QN(n12327) );
  NAND2X0 U12488 ( .IN1(n9106), .IN2(n8495), .QN(n12326) );
  NAND2X0 U12489 ( .IN1(n9292), .IN2(CRC_OUT_5_31), .QN(n12307) );
  NAND2X0 U12490 ( .IN1(n2245), .IN2(WX5657), .QN(n12306) );
  NOR2X0 U12491 ( .IN1(n9235), .IN2(WX5657), .QN(WX5718) );
  NOR2X0 U12492 ( .IN1(n9235), .IN2(WX485), .QN(WX546) );
  NOR3X0 U12493 ( .IN1(n9139), .IN2(n12329), .IN3(n12330), .QN(WX5205) );
  NOR2X0 U12494 ( .IN1(n8354), .IN2(CRC_OUT_6_30), .QN(n12330) );
  NOR2X0 U12495 ( .IN1(DFF_766_n1), .IN2(WX4716), .QN(n12329) );
  NOR3X0 U12496 ( .IN1(n9139), .IN2(n12331), .IN3(n12332), .QN(WX5203) );
  NOR2X0 U12497 ( .IN1(n8355), .IN2(CRC_OUT_6_29), .QN(n12332) );
  NOR2X0 U12498 ( .IN1(DFF_765_n1), .IN2(WX4718), .QN(n12331) );
  NOR3X0 U12499 ( .IN1(n9139), .IN2(n12333), .IN3(n12334), .QN(WX5201) );
  NOR2X0 U12500 ( .IN1(n8356), .IN2(CRC_OUT_6_28), .QN(n12334) );
  NOR2X0 U12501 ( .IN1(DFF_764_n1), .IN2(WX4720), .QN(n12333) );
  NOR2X0 U12502 ( .IN1(n9234), .IN2(n12335), .QN(WX5199) );
  NOR2X0 U12503 ( .IN1(n12336), .IN2(n12337), .QN(n12335) );
  NOR2X0 U12504 ( .IN1(test_so40), .IN2(CRC_OUT_6_27), .QN(n12337) );
  NOR2X0 U12505 ( .IN1(DFF_763_n1), .IN2(n8800), .QN(n12336) );
  NOR3X0 U12506 ( .IN1(n9139), .IN2(n12338), .IN3(n12339), .QN(WX5197) );
  NOR2X0 U12507 ( .IN1(n8357), .IN2(CRC_OUT_6_26), .QN(n12339) );
  NOR2X0 U12508 ( .IN1(DFF_762_n1), .IN2(WX4724), .QN(n12338) );
  NOR3X0 U12509 ( .IN1(n9139), .IN2(n12340), .IN3(n12341), .QN(WX5195) );
  NOR2X0 U12510 ( .IN1(n8358), .IN2(CRC_OUT_6_25), .QN(n12341) );
  NOR2X0 U12511 ( .IN1(DFF_761_n1), .IN2(WX4726), .QN(n12340) );
  NOR3X0 U12512 ( .IN1(n9139), .IN2(n12342), .IN3(n12343), .QN(WX5193) );
  NOR2X0 U12513 ( .IN1(n8359), .IN2(CRC_OUT_6_24), .QN(n12343) );
  NOR2X0 U12514 ( .IN1(DFF_760_n1), .IN2(WX4728), .QN(n12342) );
  NOR3X0 U12515 ( .IN1(n9139), .IN2(n12344), .IN3(n12345), .QN(WX5191) );
  NOR2X0 U12516 ( .IN1(n8360), .IN2(CRC_OUT_6_23), .QN(n12345) );
  NOR2X0 U12517 ( .IN1(DFF_759_n1), .IN2(WX4730), .QN(n12344) );
  NOR2X0 U12518 ( .IN1(n9234), .IN2(n12346), .QN(WX5189) );
  NOR2X0 U12519 ( .IN1(n12347), .IN2(n12348), .QN(n12346) );
  NOR2X0 U12520 ( .IN1(test_so43), .IN2(WX4732), .QN(n12348) );
  INVX0 U12521 ( .INP(n12349), .ZN(n12347) );
  NAND2X0 U12522 ( .IN1(WX4732), .IN2(test_so43), .QN(n12349) );
  NOR3X0 U12523 ( .IN1(n9139), .IN2(n12350), .IN3(n12351), .QN(WX5187) );
  NOR2X0 U12524 ( .IN1(n8362), .IN2(CRC_OUT_6_21), .QN(n12351) );
  NOR2X0 U12525 ( .IN1(DFF_757_n1), .IN2(WX4734), .QN(n12350) );
  NOR3X0 U12526 ( .IN1(n9139), .IN2(n12352), .IN3(n12353), .QN(WX5185) );
  NOR2X0 U12527 ( .IN1(n8379), .IN2(CRC_OUT_6_20), .QN(n12353) );
  NOR2X0 U12528 ( .IN1(DFF_756_n1), .IN2(WX4736), .QN(n12352) );
  NOR3X0 U12529 ( .IN1(n9138), .IN2(n12354), .IN3(n12355), .QN(WX5183) );
  NOR2X0 U12530 ( .IN1(n8380), .IN2(CRC_OUT_6_19), .QN(n12355) );
  NOR2X0 U12531 ( .IN1(DFF_755_n1), .IN2(WX4738), .QN(n12354) );
  NOR3X0 U12532 ( .IN1(n9138), .IN2(n12356), .IN3(n12357), .QN(WX5181) );
  NOR2X0 U12533 ( .IN1(n8397), .IN2(CRC_OUT_6_18), .QN(n12357) );
  NOR2X0 U12534 ( .IN1(DFF_754_n1), .IN2(WX4740), .QN(n12356) );
  NOR3X0 U12535 ( .IN1(n9138), .IN2(n12358), .IN3(n12359), .QN(WX5179) );
  NOR2X0 U12536 ( .IN1(n8398), .IN2(CRC_OUT_6_17), .QN(n12359) );
  NOR2X0 U12537 ( .IN1(DFF_753_n1), .IN2(WX4742), .QN(n12358) );
  NOR3X0 U12538 ( .IN1(n9138), .IN2(n12360), .IN3(n12361), .QN(WX5177) );
  NOR2X0 U12539 ( .IN1(n8412), .IN2(CRC_OUT_6_16), .QN(n12361) );
  NOR2X0 U12540 ( .IN1(DFF_752_n1), .IN2(WX4744), .QN(n12360) );
  NOR2X0 U12541 ( .IN1(n9234), .IN2(n12362), .QN(WX5175) );
  NOR2X0 U12542 ( .IN1(n12363), .IN2(n12364), .QN(n12362) );
  INVX0 U12543 ( .INP(n12365), .ZN(n12364) );
  NAND2X0 U12544 ( .IN1(CRC_OUT_6_15), .IN2(n12366), .QN(n12365) );
  NOR2X0 U12545 ( .IN1(n12366), .IN2(CRC_OUT_6_15), .QN(n12363) );
  NAND2X0 U12546 ( .IN1(n12367), .IN2(n12368), .QN(n12366) );
  NAND2X0 U12547 ( .IN1(n8117), .IN2(CRC_OUT_6_31), .QN(n12368) );
  NAND2X0 U12548 ( .IN1(DFF_767_n1), .IN2(WX4746), .QN(n12367) );
  NOR3X0 U12549 ( .IN1(n9138), .IN2(n12369), .IN3(n12370), .QN(WX5173) );
  NOR2X0 U12550 ( .IN1(n8413), .IN2(CRC_OUT_6_14), .QN(n12370) );
  NOR2X0 U12551 ( .IN1(DFF_750_n1), .IN2(WX4748), .QN(n12369) );
  NOR3X0 U12552 ( .IN1(n9138), .IN2(n12371), .IN3(n12372), .QN(WX5171) );
  NOR2X0 U12553 ( .IN1(n8414), .IN2(CRC_OUT_6_13), .QN(n12372) );
  NOR2X0 U12554 ( .IN1(DFF_749_n1), .IN2(WX4750), .QN(n12371) );
  NOR3X0 U12555 ( .IN1(n9138), .IN2(n12373), .IN3(n12374), .QN(WX5169) );
  NOR2X0 U12556 ( .IN1(n8415), .IN2(CRC_OUT_6_12), .QN(n12374) );
  NOR2X0 U12557 ( .IN1(DFF_748_n1), .IN2(WX4752), .QN(n12373) );
  NOR3X0 U12558 ( .IN1(n9138), .IN2(n12375), .IN3(n12376), .QN(WX5167) );
  NOR2X0 U12559 ( .IN1(n8416), .IN2(CRC_OUT_6_11), .QN(n12376) );
  NOR2X0 U12560 ( .IN1(DFF_747_n1), .IN2(WX4754), .QN(n12375) );
  NOR3X0 U12561 ( .IN1(n9138), .IN2(n12377), .IN3(n12378), .QN(WX5165) );
  INVX0 U12562 ( .INP(n12379), .ZN(n12378) );
  NAND2X0 U12563 ( .IN1(CRC_OUT_6_10), .IN2(n12380), .QN(n12379) );
  NOR2X0 U12564 ( .IN1(n12380), .IN2(CRC_OUT_6_10), .QN(n12377) );
  NAND2X0 U12565 ( .IN1(n12381), .IN2(n12382), .QN(n12380) );
  NAND2X0 U12566 ( .IN1(test_so41), .IN2(CRC_OUT_6_31), .QN(n12382) );
  NAND2X0 U12567 ( .IN1(DFF_767_n1), .IN2(n8796), .QN(n12381) );
  NOR3X0 U12568 ( .IN1(n9138), .IN2(n12383), .IN3(n12384), .QN(WX5163) );
  NOR2X0 U12569 ( .IN1(n8417), .IN2(CRC_OUT_6_9), .QN(n12384) );
  NOR2X0 U12570 ( .IN1(DFF_745_n1), .IN2(WX4758), .QN(n12383) );
  NOR3X0 U12571 ( .IN1(n9138), .IN2(n12385), .IN3(n12386), .QN(WX5161) );
  NOR2X0 U12572 ( .IN1(n8418), .IN2(CRC_OUT_6_8), .QN(n12386) );
  NOR2X0 U12573 ( .IN1(DFF_744_n1), .IN2(WX4760), .QN(n12385) );
  NOR3X0 U12574 ( .IN1(n9138), .IN2(n12387), .IN3(n12388), .QN(WX5159) );
  NOR2X0 U12575 ( .IN1(n8419), .IN2(CRC_OUT_6_7), .QN(n12388) );
  NOR2X0 U12576 ( .IN1(DFF_743_n1), .IN2(WX4762), .QN(n12387) );
  NOR3X0 U12577 ( .IN1(n9137), .IN2(n12389), .IN3(n12390), .QN(WX5157) );
  NOR2X0 U12578 ( .IN1(n8420), .IN2(CRC_OUT_6_6), .QN(n12390) );
  NOR2X0 U12579 ( .IN1(DFF_742_n1), .IN2(WX4764), .QN(n12389) );
  NOR2X0 U12580 ( .IN1(n9231), .IN2(n12391), .QN(WX5155) );
  NOR2X0 U12581 ( .IN1(n12392), .IN2(n12393), .QN(n12391) );
  NOR2X0 U12582 ( .IN1(test_so42), .IN2(WX4766), .QN(n12393) );
  INVX0 U12583 ( .INP(n12394), .ZN(n12392) );
  NAND2X0 U12584 ( .IN1(WX4766), .IN2(test_so42), .QN(n12394) );
  NOR3X0 U12585 ( .IN1(n9137), .IN2(n12395), .IN3(n12396), .QN(WX5153) );
  NOR2X0 U12586 ( .IN1(n8433), .IN2(CRC_OUT_6_4), .QN(n12396) );
  NOR2X0 U12587 ( .IN1(DFF_740_n1), .IN2(WX4768), .QN(n12395) );
  NOR2X0 U12588 ( .IN1(n9231), .IN2(n12397), .QN(WX5151) );
  NOR2X0 U12589 ( .IN1(n12398), .IN2(n12399), .QN(n12397) );
  INVX0 U12590 ( .INP(n12400), .ZN(n12399) );
  NAND2X0 U12591 ( .IN1(CRC_OUT_6_3), .IN2(n12401), .QN(n12400) );
  NOR2X0 U12592 ( .IN1(n12401), .IN2(CRC_OUT_6_3), .QN(n12398) );
  NAND2X0 U12593 ( .IN1(n12402), .IN2(n12403), .QN(n12401) );
  NAND2X0 U12594 ( .IN1(n8118), .IN2(CRC_OUT_6_31), .QN(n12403) );
  NAND2X0 U12595 ( .IN1(DFF_767_n1), .IN2(WX4770), .QN(n12402) );
  NOR3X0 U12596 ( .IN1(n9137), .IN2(n12404), .IN3(n12405), .QN(WX5149) );
  NOR2X0 U12597 ( .IN1(n8450), .IN2(CRC_OUT_6_2), .QN(n12405) );
  NOR2X0 U12598 ( .IN1(DFF_738_n1), .IN2(WX4772), .QN(n12404) );
  NOR3X0 U12599 ( .IN1(n9137), .IN2(n12406), .IN3(n12407), .QN(WX5147) );
  NOR2X0 U12600 ( .IN1(n8451), .IN2(CRC_OUT_6_1), .QN(n12407) );
  NOR2X0 U12601 ( .IN1(DFF_737_n1), .IN2(WX4774), .QN(n12406) );
  NOR3X0 U12602 ( .IN1(n9137), .IN2(n12408), .IN3(n12409), .QN(WX5145) );
  NOR2X0 U12603 ( .IN1(n8468), .IN2(CRC_OUT_6_0), .QN(n12409) );
  NOR2X0 U12604 ( .IN1(DFF_736_n1), .IN2(WX4776), .QN(n12408) );
  NOR3X0 U12605 ( .IN1(n9137), .IN2(n12410), .IN3(n12411), .QN(WX5143) );
  NOR2X0 U12606 ( .IN1(n8130), .IN2(CRC_OUT_6_31), .QN(n12411) );
  NOR2X0 U12607 ( .IN1(DFF_767_n1), .IN2(WX4778), .QN(n12410) );
  NOR2X0 U12608 ( .IN1(n16071), .IN2(n9161), .QN(WX4617) );
  NOR2X0 U12609 ( .IN1(n9223), .IN2(n8822), .QN(WX4615) );
  NOR2X0 U12610 ( .IN1(n16070), .IN2(n9161), .QN(WX4613) );
  NOR2X0 U12611 ( .IN1(n16069), .IN2(n9161), .QN(WX4611) );
  NOR2X0 U12612 ( .IN1(n16068), .IN2(n9161), .QN(WX4609) );
  NOR2X0 U12613 ( .IN1(n16067), .IN2(n9161), .QN(WX4607) );
  NOR2X0 U12614 ( .IN1(n16066), .IN2(n9161), .QN(WX4605) );
  NOR2X0 U12615 ( .IN1(n16065), .IN2(n9160), .QN(WX4603) );
  NOR2X0 U12616 ( .IN1(n16064), .IN2(n9160), .QN(WX4601) );
  NOR2X0 U12617 ( .IN1(n16063), .IN2(n9160), .QN(WX4599) );
  NOR2X0 U12618 ( .IN1(n16062), .IN2(n9160), .QN(WX4597) );
  NOR2X0 U12619 ( .IN1(n16061), .IN2(n9160), .QN(WX4595) );
  NOR2X0 U12620 ( .IN1(n16060), .IN2(n9160), .QN(WX4593) );
  NOR2X0 U12621 ( .IN1(n16059), .IN2(n9160), .QN(WX4591) );
  NOR2X0 U12622 ( .IN1(n16058), .IN2(n9160), .QN(WX4589) );
  NOR2X0 U12623 ( .IN1(n16057), .IN2(n9160), .QN(WX4587) );
  NAND4X0 U12624 ( .IN1(n12412), .IN2(n12413), .IN3(n12414), .IN4(n12415), 
        .QN(WX4585) );
  NAND3X0 U12625 ( .IN1(n12416), .IN2(n12417), .IN3(n9089), .QN(n12415) );
  NAND2X0 U12626 ( .IN1(n9323), .IN2(n11743), .QN(n12414) );
  NAND2X0 U12627 ( .IN1(n12418), .IN2(n12419), .QN(n11743) );
  INVX0 U12628 ( .INP(n12420), .ZN(n12419) );
  NOR2X0 U12629 ( .IN1(n12421), .IN2(n12422), .QN(n12420) );
  NAND2X0 U12630 ( .IN1(n12422), .IN2(n12421), .QN(n12418) );
  NOR2X0 U12631 ( .IN1(n12423), .IN2(n12424), .QN(n12421) );
  NOR2X0 U12632 ( .IN1(WX6071), .IN2(n7975), .QN(n12424) );
  INVX0 U12633 ( .INP(n12425), .ZN(n12423) );
  NAND2X0 U12634 ( .IN1(n7975), .IN2(WX6071), .QN(n12425) );
  NAND2X0 U12635 ( .IN1(n12426), .IN2(n12427), .QN(n12422) );
  NAND2X0 U12636 ( .IN1(n7974), .IN2(WX5943), .QN(n12427) );
  INVX0 U12637 ( .INP(n12428), .ZN(n12426) );
  NOR2X0 U12638 ( .IN1(WX5943), .IN2(n7974), .QN(n12428) );
  NAND2X0 U12639 ( .IN1(n762), .IN2(n9281), .QN(n12413) );
  NOR2X0 U12640 ( .IN1(n9231), .IN2(n8944), .QN(n762) );
  NAND2X0 U12641 ( .IN1(n9292), .IN2(CRC_OUT_6_0), .QN(n12412) );
  NAND4X0 U12642 ( .IN1(n12429), .IN2(n12430), .IN3(n12431), .IN4(n12432), 
        .QN(WX4583) );
  NAND3X0 U12643 ( .IN1(n11748), .IN2(n11749), .IN3(n9321), .QN(n12432) );
  NAND3X0 U12644 ( .IN1(n12433), .IN2(n12434), .IN3(n12435), .QN(n11749) );
  INVX0 U12645 ( .INP(n12436), .ZN(n12435) );
  NAND2X0 U12646 ( .IN1(n12436), .IN2(n12437), .QN(n11748) );
  NAND2X0 U12647 ( .IN1(n12433), .IN2(n12434), .QN(n12437) );
  NAND2X0 U12648 ( .IN1(n8345), .IN2(WX5941), .QN(n12434) );
  NAND2X0 U12649 ( .IN1(n3661), .IN2(WX6069), .QN(n12433) );
  NOR2X0 U12650 ( .IN1(n12438), .IN2(n12439), .QN(n12436) );
  INVX0 U12651 ( .INP(n12440), .ZN(n12439) );
  NAND2X0 U12652 ( .IN1(test_so51), .IN2(WX5877), .QN(n12440) );
  NOR2X0 U12653 ( .IN1(WX5877), .IN2(test_so51), .QN(n12438) );
  NAND2X0 U12654 ( .IN1(n9106), .IN2(n12441), .QN(n12431) );
  NAND2X0 U12655 ( .IN1(n761), .IN2(n9281), .QN(n12430) );
  NOR2X0 U12656 ( .IN1(n9231), .IN2(n8945), .QN(n761) );
  NAND2X0 U12657 ( .IN1(n9292), .IN2(CRC_OUT_6_1), .QN(n12429) );
  NAND4X0 U12658 ( .IN1(n12442), .IN2(n12443), .IN3(n12444), .IN4(n12445), 
        .QN(WX4581) );
  NAND2X0 U12659 ( .IN1(n9323), .IN2(n11776), .QN(n12445) );
  NAND2X0 U12660 ( .IN1(n12446), .IN2(n12447), .QN(n11776) );
  INVX0 U12661 ( .INP(n12448), .ZN(n12447) );
  NOR2X0 U12662 ( .IN1(n12449), .IN2(n12450), .QN(n12448) );
  NAND2X0 U12663 ( .IN1(n12450), .IN2(n12449), .QN(n12446) );
  NOR2X0 U12664 ( .IN1(n12451), .IN2(n12452), .QN(n12449) );
  NOR2X0 U12665 ( .IN1(WX6067), .IN2(n7978), .QN(n12452) );
  INVX0 U12666 ( .INP(n12453), .ZN(n12451) );
  NAND2X0 U12667 ( .IN1(n7978), .IN2(WX6067), .QN(n12453) );
  NAND2X0 U12668 ( .IN1(n12454), .IN2(n12455), .QN(n12450) );
  NAND2X0 U12669 ( .IN1(n7977), .IN2(WX5939), .QN(n12455) );
  INVX0 U12670 ( .INP(n12456), .ZN(n12454) );
  NOR2X0 U12671 ( .IN1(WX5939), .IN2(n7977), .QN(n12456) );
  NAND2X0 U12672 ( .IN1(n9106), .IN2(n12457), .QN(n12444) );
  NAND2X0 U12673 ( .IN1(n760), .IN2(n9281), .QN(n12443) );
  NOR2X0 U12674 ( .IN1(n9068), .IN2(n9160), .QN(n760) );
  NAND2X0 U12675 ( .IN1(n9292), .IN2(CRC_OUT_6_2), .QN(n12442) );
  NAND4X0 U12676 ( .IN1(n12458), .IN2(n12459), .IN3(n12460), .IN4(n12461), 
        .QN(WX4579) );
  NAND3X0 U12677 ( .IN1(n11781), .IN2(n11782), .IN3(n9320), .QN(n12461) );
  NAND3X0 U12678 ( .IN1(n12462), .IN2(n12463), .IN3(n12464), .QN(n11782) );
  INVX0 U12679 ( .INP(n12465), .ZN(n12464) );
  NAND2X0 U12680 ( .IN1(n12465), .IN2(n12466), .QN(n11781) );
  NAND2X0 U12681 ( .IN1(n12462), .IN2(n12463), .QN(n12466) );
  NAND2X0 U12682 ( .IN1(n8327), .IN2(WX6001), .QN(n12463) );
  NAND2X0 U12683 ( .IN1(n7980), .IN2(WX6065), .QN(n12462) );
  NOR2X0 U12684 ( .IN1(n12467), .IN2(n12468), .QN(n12465) );
  INVX0 U12685 ( .INP(n12469), .ZN(n12468) );
  NAND2X0 U12686 ( .IN1(test_so49), .IN2(WX5873), .QN(n12469) );
  NOR2X0 U12687 ( .IN1(WX5873), .IN2(test_so49), .QN(n12467) );
  NAND2X0 U12688 ( .IN1(n9106), .IN2(n12470), .QN(n12460) );
  NAND2X0 U12689 ( .IN1(n759), .IN2(n9281), .QN(n12459) );
  NOR2X0 U12690 ( .IN1(n9232), .IN2(n8946), .QN(n759) );
  NAND2X0 U12691 ( .IN1(n9292), .IN2(CRC_OUT_6_3), .QN(n12458) );
  NAND4X0 U12692 ( .IN1(n12471), .IN2(n12472), .IN3(n12473), .IN4(n12474), 
        .QN(WX4577) );
  NAND2X0 U12693 ( .IN1(n9323), .IN2(n11806), .QN(n12474) );
  NAND2X0 U12694 ( .IN1(n12475), .IN2(n12476), .QN(n11806) );
  INVX0 U12695 ( .INP(n12477), .ZN(n12476) );
  NOR2X0 U12696 ( .IN1(n12478), .IN2(n12479), .QN(n12477) );
  NAND2X0 U12697 ( .IN1(n12479), .IN2(n12478), .QN(n12475) );
  NOR2X0 U12698 ( .IN1(n12480), .IN2(n12481), .QN(n12478) );
  NOR2X0 U12699 ( .IN1(WX6063), .IN2(n7982), .QN(n12481) );
  INVX0 U12700 ( .INP(n12482), .ZN(n12480) );
  NAND2X0 U12701 ( .IN1(n7982), .IN2(WX6063), .QN(n12482) );
  NAND2X0 U12702 ( .IN1(n12483), .IN2(n12484), .QN(n12479) );
  NAND2X0 U12703 ( .IN1(n7981), .IN2(WX5935), .QN(n12484) );
  INVX0 U12704 ( .INP(n12485), .ZN(n12483) );
  NOR2X0 U12705 ( .IN1(WX5935), .IN2(n7981), .QN(n12485) );
  NAND2X0 U12706 ( .IN1(n9106), .IN2(n12486), .QN(n12473) );
  NAND2X0 U12707 ( .IN1(n758), .IN2(n9281), .QN(n12472) );
  NOR2X0 U12708 ( .IN1(n9232), .IN2(n8947), .QN(n758) );
  NAND2X0 U12709 ( .IN1(n9292), .IN2(CRC_OUT_6_4), .QN(n12471) );
  NAND4X0 U12710 ( .IN1(n12487), .IN2(n12488), .IN3(n12489), .IN4(n12490), 
        .QN(WX4575) );
  NAND3X0 U12711 ( .IN1(n11811), .IN2(n11812), .IN3(n9321), .QN(n12490) );
  NAND3X0 U12712 ( .IN1(n12491), .IN2(n12492), .IN3(n12493), .QN(n11812) );
  INVX0 U12713 ( .INP(n12494), .ZN(n12493) );
  NAND2X0 U12714 ( .IN1(n12494), .IN2(n12495), .QN(n11811) );
  NAND2X0 U12715 ( .IN1(n12491), .IN2(n12492), .QN(n12495) );
  NAND2X0 U12716 ( .IN1(n8326), .IN2(WX5933), .QN(n12492) );
  NAND2X0 U12717 ( .IN1(n3669), .IN2(WX6061), .QN(n12491) );
  NOR2X0 U12718 ( .IN1(n12496), .IN2(n12497), .QN(n12494) );
  INVX0 U12719 ( .INP(n12498), .ZN(n12497) );
  NAND2X0 U12720 ( .IN1(test_so47), .IN2(WX5997), .QN(n12498) );
  NOR2X0 U12721 ( .IN1(WX5997), .IN2(test_so47), .QN(n12496) );
  NAND2X0 U12722 ( .IN1(n9106), .IN2(n12499), .QN(n12489) );
  NAND2X0 U12723 ( .IN1(n757), .IN2(n9281), .QN(n12488) );
  NOR2X0 U12724 ( .IN1(n9232), .IN2(n8948), .QN(n757) );
  NAND2X0 U12725 ( .IN1(test_so42), .IN2(n9314), .QN(n12487) );
  NAND4X0 U12726 ( .IN1(n12500), .IN2(n12501), .IN3(n12502), .IN4(n12503), 
        .QN(WX4573) );
  NAND2X0 U12727 ( .IN1(n9324), .IN2(n11836), .QN(n12503) );
  NAND2X0 U12728 ( .IN1(n12504), .IN2(n12505), .QN(n11836) );
  INVX0 U12729 ( .INP(n12506), .ZN(n12505) );
  NOR2X0 U12730 ( .IN1(n12507), .IN2(n12508), .QN(n12506) );
  NAND2X0 U12731 ( .IN1(n12508), .IN2(n12507), .QN(n12504) );
  NOR2X0 U12732 ( .IN1(n12509), .IN2(n12510), .QN(n12507) );
  NOR2X0 U12733 ( .IN1(WX6059), .IN2(n7985), .QN(n12510) );
  INVX0 U12734 ( .INP(n12511), .ZN(n12509) );
  NAND2X0 U12735 ( .IN1(n7985), .IN2(WX6059), .QN(n12511) );
  NAND2X0 U12736 ( .IN1(n12512), .IN2(n12513), .QN(n12508) );
  NAND2X0 U12737 ( .IN1(n7984), .IN2(WX5931), .QN(n12513) );
  INVX0 U12738 ( .INP(n12514), .ZN(n12512) );
  NOR2X0 U12739 ( .IN1(WX5931), .IN2(n7984), .QN(n12514) );
  NAND2X0 U12740 ( .IN1(n9106), .IN2(n12515), .QN(n12502) );
  NAND2X0 U12741 ( .IN1(n756), .IN2(n9281), .QN(n12501) );
  NOR2X0 U12742 ( .IN1(n9232), .IN2(n8949), .QN(n756) );
  NAND2X0 U12743 ( .IN1(n9293), .IN2(CRC_OUT_6_6), .QN(n12500) );
  NAND4X0 U12744 ( .IN1(n12516), .IN2(n12517), .IN3(n12518), .IN4(n12519), 
        .QN(WX4571) );
  NAND2X0 U12745 ( .IN1(n9323), .IN2(n11852), .QN(n12519) );
  NAND2X0 U12746 ( .IN1(n12520), .IN2(n12521), .QN(n11852) );
  INVX0 U12747 ( .INP(n12522), .ZN(n12521) );
  NOR2X0 U12748 ( .IN1(n12523), .IN2(n12524), .QN(n12522) );
  NAND2X0 U12749 ( .IN1(n12524), .IN2(n12523), .QN(n12520) );
  NOR2X0 U12750 ( .IN1(n12525), .IN2(n12526), .QN(n12523) );
  NOR2X0 U12751 ( .IN1(WX6057), .IN2(n7987), .QN(n12526) );
  INVX0 U12752 ( .INP(n12527), .ZN(n12525) );
  NAND2X0 U12753 ( .IN1(n7987), .IN2(WX6057), .QN(n12527) );
  NAND2X0 U12754 ( .IN1(n12528), .IN2(n12529), .QN(n12524) );
  NAND2X0 U12755 ( .IN1(n7986), .IN2(WX5929), .QN(n12529) );
  INVX0 U12756 ( .INP(n12530), .ZN(n12528) );
  NOR2X0 U12757 ( .IN1(WX5929), .IN2(n7986), .QN(n12530) );
  NAND2X0 U12758 ( .IN1(n9106), .IN2(n12531), .QN(n12518) );
  NAND2X0 U12759 ( .IN1(n755), .IN2(n9281), .QN(n12517) );
  NOR2X0 U12760 ( .IN1(n9232), .IN2(n8950), .QN(n755) );
  NAND2X0 U12761 ( .IN1(n9293), .IN2(CRC_OUT_6_7), .QN(n12516) );
  NAND4X0 U12762 ( .IN1(n12532), .IN2(n12533), .IN3(n12534), .IN4(n12535), 
        .QN(WX4569) );
  NAND2X0 U12763 ( .IN1(n9323), .IN2(n11865), .QN(n12535) );
  NAND2X0 U12764 ( .IN1(n12536), .IN2(n12537), .QN(n11865) );
  INVX0 U12765 ( .INP(n12538), .ZN(n12537) );
  NOR2X0 U12766 ( .IN1(n12539), .IN2(n12540), .QN(n12538) );
  NAND2X0 U12767 ( .IN1(n12540), .IN2(n12539), .QN(n12536) );
  NOR2X0 U12768 ( .IN1(n12541), .IN2(n12542), .QN(n12539) );
  NOR2X0 U12769 ( .IN1(WX6055), .IN2(n7989), .QN(n12542) );
  INVX0 U12770 ( .INP(n12543), .ZN(n12541) );
  NAND2X0 U12771 ( .IN1(n7989), .IN2(WX6055), .QN(n12543) );
  NAND2X0 U12772 ( .IN1(n12544), .IN2(n12545), .QN(n12540) );
  NAND2X0 U12773 ( .IN1(n7988), .IN2(WX5927), .QN(n12545) );
  INVX0 U12774 ( .INP(n12546), .ZN(n12544) );
  NOR2X0 U12775 ( .IN1(WX5927), .IN2(n7988), .QN(n12546) );
  NAND2X0 U12776 ( .IN1(n9106), .IN2(n12547), .QN(n12534) );
  NAND2X0 U12777 ( .IN1(n754), .IN2(n9281), .QN(n12533) );
  NOR2X0 U12778 ( .IN1(n9232), .IN2(n8951), .QN(n754) );
  NAND2X0 U12779 ( .IN1(n9293), .IN2(CRC_OUT_6_8), .QN(n12532) );
  NAND4X0 U12780 ( .IN1(n12548), .IN2(n12549), .IN3(n12550), .IN4(n12551), 
        .QN(WX4567) );
  NAND2X0 U12781 ( .IN1(n9323), .IN2(n11881), .QN(n12551) );
  NAND2X0 U12782 ( .IN1(n12552), .IN2(n12553), .QN(n11881) );
  INVX0 U12783 ( .INP(n12554), .ZN(n12553) );
  NOR2X0 U12784 ( .IN1(n12555), .IN2(n12556), .QN(n12554) );
  NAND2X0 U12785 ( .IN1(n12556), .IN2(n12555), .QN(n12552) );
  NOR2X0 U12786 ( .IN1(n12557), .IN2(n12558), .QN(n12555) );
  NOR2X0 U12787 ( .IN1(WX6053), .IN2(n7991), .QN(n12558) );
  INVX0 U12788 ( .INP(n12559), .ZN(n12557) );
  NAND2X0 U12789 ( .IN1(n7991), .IN2(WX6053), .QN(n12559) );
  NAND2X0 U12790 ( .IN1(n12560), .IN2(n12561), .QN(n12556) );
  NAND2X0 U12791 ( .IN1(n7990), .IN2(WX5925), .QN(n12561) );
  INVX0 U12792 ( .INP(n12562), .ZN(n12560) );
  NOR2X0 U12793 ( .IN1(WX5925), .IN2(n7990), .QN(n12562) );
  NAND2X0 U12794 ( .IN1(n9106), .IN2(n12563), .QN(n12550) );
  NAND2X0 U12795 ( .IN1(n753), .IN2(n9281), .QN(n12549) );
  NOR2X0 U12796 ( .IN1(n9232), .IN2(n8952), .QN(n753) );
  NAND2X0 U12797 ( .IN1(n9293), .IN2(CRC_OUT_6_9), .QN(n12548) );
  NAND4X0 U12798 ( .IN1(n12564), .IN2(n12565), .IN3(n12566), .IN4(n12567), 
        .QN(WX4565) );
  NAND2X0 U12799 ( .IN1(n9324), .IN2(n11894), .QN(n12567) );
  NAND2X0 U12800 ( .IN1(n12568), .IN2(n12569), .QN(n11894) );
  INVX0 U12801 ( .INP(n12570), .ZN(n12569) );
  NOR2X0 U12802 ( .IN1(n12571), .IN2(n12572), .QN(n12570) );
  NAND2X0 U12803 ( .IN1(n12572), .IN2(n12571), .QN(n12568) );
  NOR2X0 U12804 ( .IN1(n12573), .IN2(n12574), .QN(n12571) );
  NOR2X0 U12805 ( .IN1(WX6051), .IN2(n7993), .QN(n12574) );
  INVX0 U12806 ( .INP(n12575), .ZN(n12573) );
  NAND2X0 U12807 ( .IN1(n7993), .IN2(WX6051), .QN(n12575) );
  NAND2X0 U12808 ( .IN1(n12576), .IN2(n12577), .QN(n12572) );
  NAND2X0 U12809 ( .IN1(n7992), .IN2(WX5923), .QN(n12577) );
  INVX0 U12810 ( .INP(n12578), .ZN(n12576) );
  NOR2X0 U12811 ( .IN1(WX5923), .IN2(n7992), .QN(n12578) );
  NAND2X0 U12812 ( .IN1(n9106), .IN2(n12579), .QN(n12566) );
  NAND2X0 U12813 ( .IN1(n752), .IN2(n9281), .QN(n12565) );
  NOR2X0 U12814 ( .IN1(n9232), .IN2(n8953), .QN(n752) );
  NAND2X0 U12815 ( .IN1(n9293), .IN2(CRC_OUT_6_10), .QN(n12564) );
  NAND4X0 U12816 ( .IN1(n12580), .IN2(n12581), .IN3(n12582), .IN4(n12583), 
        .QN(WX4563) );
  NAND3X0 U12817 ( .IN1(n12584), .IN2(n12585), .IN3(n9090), .QN(n12583) );
  NAND2X0 U12818 ( .IN1(n9324), .IN2(n11910), .QN(n12582) );
  NAND2X0 U12819 ( .IN1(n12586), .IN2(n12587), .QN(n11910) );
  INVX0 U12820 ( .INP(n12588), .ZN(n12587) );
  NOR2X0 U12821 ( .IN1(n12589), .IN2(n12590), .QN(n12588) );
  NAND2X0 U12822 ( .IN1(n12590), .IN2(n12589), .QN(n12586) );
  NOR2X0 U12823 ( .IN1(n12591), .IN2(n12592), .QN(n12589) );
  NOR2X0 U12824 ( .IN1(WX6049), .IN2(n7995), .QN(n12592) );
  INVX0 U12825 ( .INP(n12593), .ZN(n12591) );
  NAND2X0 U12826 ( .IN1(n7995), .IN2(WX6049), .QN(n12593) );
  NAND2X0 U12827 ( .IN1(n12594), .IN2(n12595), .QN(n12590) );
  NAND2X0 U12828 ( .IN1(n7994), .IN2(WX5921), .QN(n12595) );
  INVX0 U12829 ( .INP(n12596), .ZN(n12594) );
  NOR2X0 U12830 ( .IN1(WX5921), .IN2(n7994), .QN(n12596) );
  NAND2X0 U12831 ( .IN1(n751), .IN2(n9281), .QN(n12581) );
  NOR2X0 U12832 ( .IN1(n9232), .IN2(n8954), .QN(n751) );
  NAND2X0 U12833 ( .IN1(n9293), .IN2(CRC_OUT_6_11), .QN(n12580) );
  NAND4X0 U12834 ( .IN1(n12597), .IN2(n12598), .IN3(n12599), .IN4(n12600), 
        .QN(WX4561) );
  NAND2X0 U12835 ( .IN1(n9324), .IN2(n11926), .QN(n12600) );
  NAND2X0 U12836 ( .IN1(n12601), .IN2(n12602), .QN(n11926) );
  INVX0 U12837 ( .INP(n12603), .ZN(n12602) );
  NOR2X0 U12838 ( .IN1(n12604), .IN2(n12605), .QN(n12603) );
  NAND2X0 U12839 ( .IN1(n12605), .IN2(n12604), .QN(n12601) );
  NOR2X0 U12840 ( .IN1(n12606), .IN2(n12607), .QN(n12604) );
  NOR2X0 U12841 ( .IN1(WX6047), .IN2(n7997), .QN(n12607) );
  INVX0 U12842 ( .INP(n12608), .ZN(n12606) );
  NAND2X0 U12843 ( .IN1(n7997), .IN2(WX6047), .QN(n12608) );
  NAND2X0 U12844 ( .IN1(n12609), .IN2(n12610), .QN(n12605) );
  NAND2X0 U12845 ( .IN1(n7996), .IN2(WX5919), .QN(n12610) );
  INVX0 U12846 ( .INP(n12611), .ZN(n12609) );
  NOR2X0 U12847 ( .IN1(WX5919), .IN2(n7996), .QN(n12611) );
  NAND2X0 U12848 ( .IN1(n9106), .IN2(n12612), .QN(n12599) );
  NAND2X0 U12849 ( .IN1(n750), .IN2(n9281), .QN(n12598) );
  NOR2X0 U12850 ( .IN1(n9232), .IN2(n8955), .QN(n750) );
  NAND2X0 U12851 ( .IN1(n9293), .IN2(CRC_OUT_6_12), .QN(n12597) );
  NAND4X0 U12852 ( .IN1(n12613), .IN2(n12614), .IN3(n12615), .IN4(n12616), 
        .QN(WX4559) );
  NAND3X0 U12853 ( .IN1(n12617), .IN2(n12618), .IN3(n9090), .QN(n12616) );
  NAND2X0 U12854 ( .IN1(n9324), .IN2(n11942), .QN(n12615) );
  NAND2X0 U12855 ( .IN1(n12619), .IN2(n12620), .QN(n11942) );
  INVX0 U12856 ( .INP(n12621), .ZN(n12620) );
  NOR2X0 U12857 ( .IN1(n12622), .IN2(n12623), .QN(n12621) );
  NAND2X0 U12858 ( .IN1(n12623), .IN2(n12622), .QN(n12619) );
  NOR2X0 U12859 ( .IN1(n12624), .IN2(n12625), .QN(n12622) );
  NOR2X0 U12860 ( .IN1(WX6045), .IN2(n7999), .QN(n12625) );
  INVX0 U12861 ( .INP(n12626), .ZN(n12624) );
  NAND2X0 U12862 ( .IN1(n7999), .IN2(WX6045), .QN(n12626) );
  NAND2X0 U12863 ( .IN1(n12627), .IN2(n12628), .QN(n12623) );
  NAND2X0 U12864 ( .IN1(n7998), .IN2(WX5917), .QN(n12628) );
  INVX0 U12865 ( .INP(n12629), .ZN(n12627) );
  NOR2X0 U12866 ( .IN1(WX5917), .IN2(n7998), .QN(n12629) );
  NAND2X0 U12867 ( .IN1(n749), .IN2(n9281), .QN(n12614) );
  NOR2X0 U12868 ( .IN1(n9232), .IN2(n8956), .QN(n749) );
  NAND2X0 U12869 ( .IN1(n9293), .IN2(CRC_OUT_6_13), .QN(n12613) );
  NAND4X0 U12870 ( .IN1(n12630), .IN2(n12631), .IN3(n12632), .IN4(n12633), 
        .QN(WX4557) );
  NAND2X0 U12871 ( .IN1(n9324), .IN2(n11958), .QN(n12633) );
  NAND2X0 U12872 ( .IN1(n12634), .IN2(n12635), .QN(n11958) );
  INVX0 U12873 ( .INP(n12636), .ZN(n12635) );
  NOR2X0 U12874 ( .IN1(n12637), .IN2(n12638), .QN(n12636) );
  NAND2X0 U12875 ( .IN1(n12638), .IN2(n12637), .QN(n12634) );
  NOR2X0 U12876 ( .IN1(n12639), .IN2(n12640), .QN(n12637) );
  NOR2X0 U12877 ( .IN1(WX6043), .IN2(n8001), .QN(n12640) );
  INVX0 U12878 ( .INP(n12641), .ZN(n12639) );
  NAND2X0 U12879 ( .IN1(n8001), .IN2(WX6043), .QN(n12641) );
  NAND2X0 U12880 ( .IN1(n12642), .IN2(n12643), .QN(n12638) );
  NAND2X0 U12881 ( .IN1(n8000), .IN2(WX5915), .QN(n12643) );
  INVX0 U12882 ( .INP(n12644), .ZN(n12642) );
  NOR2X0 U12883 ( .IN1(WX5915), .IN2(n8000), .QN(n12644) );
  NAND2X0 U12884 ( .IN1(n9106), .IN2(n12645), .QN(n12632) );
  NAND2X0 U12885 ( .IN1(n748), .IN2(n9282), .QN(n12631) );
  NOR2X0 U12886 ( .IN1(n9232), .IN2(n8957), .QN(n748) );
  NAND2X0 U12887 ( .IN1(n9293), .IN2(CRC_OUT_6_14), .QN(n12630) );
  NAND4X0 U12888 ( .IN1(n12646), .IN2(n12647), .IN3(n12648), .IN4(n12649), 
        .QN(WX4555) );
  NAND3X0 U12889 ( .IN1(n12650), .IN2(n12651), .IN3(n9090), .QN(n12649) );
  NAND2X0 U12890 ( .IN1(n9324), .IN2(n11974), .QN(n12648) );
  NAND2X0 U12891 ( .IN1(n12652), .IN2(n12653), .QN(n11974) );
  INVX0 U12892 ( .INP(n12654), .ZN(n12653) );
  NOR2X0 U12893 ( .IN1(n12655), .IN2(n12656), .QN(n12654) );
  NAND2X0 U12894 ( .IN1(n12656), .IN2(n12655), .QN(n12652) );
  NOR2X0 U12895 ( .IN1(n12657), .IN2(n12658), .QN(n12655) );
  NOR2X0 U12896 ( .IN1(WX6041), .IN2(n8003), .QN(n12658) );
  INVX0 U12897 ( .INP(n12659), .ZN(n12657) );
  NAND2X0 U12898 ( .IN1(n8003), .IN2(WX6041), .QN(n12659) );
  NAND2X0 U12899 ( .IN1(n12660), .IN2(n12661), .QN(n12656) );
  NAND2X0 U12900 ( .IN1(n8002), .IN2(WX5913), .QN(n12661) );
  INVX0 U12901 ( .INP(n12662), .ZN(n12660) );
  NOR2X0 U12902 ( .IN1(WX5913), .IN2(n8002), .QN(n12662) );
  NAND2X0 U12903 ( .IN1(n747), .IN2(n9282), .QN(n12647) );
  NOR2X0 U12904 ( .IN1(n9232), .IN2(n8958), .QN(n747) );
  NAND2X0 U12905 ( .IN1(n9293), .IN2(CRC_OUT_6_15), .QN(n12646) );
  NAND4X0 U12906 ( .IN1(n12663), .IN2(n12664), .IN3(n12665), .IN4(n12666), 
        .QN(WX4553) );
  NAND2X0 U12907 ( .IN1(n12667), .IN2(n12668), .QN(n12666) );
  NAND2X0 U12908 ( .IN1(n12669), .IN2(n12670), .QN(n12667) );
  NAND2X0 U12909 ( .IN1(n9106), .IN2(n12671), .QN(n12670) );
  NAND2X0 U12910 ( .IN1(n9107), .IN2(n8537), .QN(n12669) );
  NAND2X0 U12911 ( .IN1(n11993), .IN2(n2153), .QN(n12665) );
  NOR2X0 U12912 ( .IN1(n12672), .IN2(n12673), .QN(n11993) );
  INVX0 U12913 ( .INP(n12674), .ZN(n12673) );
  NAND2X0 U12914 ( .IN1(n12675), .IN2(n12676), .QN(n12674) );
  NOR2X0 U12915 ( .IN1(n12676), .IN2(n12675), .QN(n12672) );
  NAND2X0 U12916 ( .IN1(n12677), .IN2(n12678), .QN(n12675) );
  NAND2X0 U12917 ( .IN1(n12679), .IN2(WX5975), .QN(n12678) );
  NAND2X0 U12918 ( .IN1(n12680), .IN2(n12681), .QN(n12679) );
  NAND3X0 U12919 ( .IN1(n12680), .IN2(n12681), .IN3(n7740), .QN(n12677) );
  NAND2X0 U12920 ( .IN1(test_so52), .IN2(WX5911), .QN(n12681) );
  NAND2X0 U12921 ( .IN1(n7739), .IN2(n8826), .QN(n12680) );
  NOR2X0 U12922 ( .IN1(n12682), .IN2(n12683), .QN(n12676) );
  INVX0 U12923 ( .INP(n12684), .ZN(n12683) );
  NAND2X0 U12924 ( .IN1(n16086), .IN2(n9117), .QN(n12684) );
  NOR2X0 U12925 ( .IN1(n9116), .IN2(n16086), .QN(n12682) );
  NAND2X0 U12926 ( .IN1(n746), .IN2(n9282), .QN(n12664) );
  NOR2X0 U12927 ( .IN1(n9232), .IN2(n8959), .QN(n746) );
  NAND2X0 U12928 ( .IN1(n9293), .IN2(CRC_OUT_6_16), .QN(n12663) );
  NAND4X0 U12929 ( .IN1(n12685), .IN2(n12686), .IN3(n12687), .IN4(n12688), 
        .QN(WX4551) );
  NAND2X0 U12930 ( .IN1(n12689), .IN2(n12013), .QN(n12688) );
  NAND2X0 U12931 ( .IN1(n12690), .IN2(n12016), .QN(n12013) );
  NAND2X0 U12932 ( .IN1(n12691), .IN2(n12692), .QN(n12690) );
  NAND2X0 U12933 ( .IN1(n16085), .IN2(n9117), .QN(n12692) );
  NAND2X0 U12934 ( .IN1(TM1), .IN2(n8480), .QN(n12691) );
  NAND3X0 U12935 ( .IN1(n12693), .IN2(n12694), .IN3(n12695), .QN(n12689) );
  NAND2X0 U12936 ( .IN1(n9324), .IN2(n12016), .QN(n12695) );
  NAND2X0 U12937 ( .IN1(n12696), .IN2(n12697), .QN(n12016) );
  NAND2X0 U12938 ( .IN1(n7741), .IN2(n12698), .QN(n12697) );
  INVX0 U12939 ( .INP(n12699), .ZN(n12696) );
  NOR2X0 U12940 ( .IN1(n12698), .IN2(n7741), .QN(n12699) );
  NOR2X0 U12941 ( .IN1(n12700), .IN2(n12701), .QN(n12698) );
  NOR2X0 U12942 ( .IN1(WX6037), .IN2(n7742), .QN(n12701) );
  INVX0 U12943 ( .INP(n12702), .ZN(n12700) );
  NAND2X0 U12944 ( .IN1(n7742), .IN2(WX6037), .QN(n12702) );
  NAND2X0 U12945 ( .IN1(n9081), .IN2(n8480), .QN(n12694) );
  NAND2X0 U12946 ( .IN1(n16085), .IN2(n9078), .QN(n12693) );
  NAND2X0 U12947 ( .IN1(n12703), .IN2(n12704), .QN(n12687) );
  NAND2X0 U12948 ( .IN1(n12705), .IN2(n12706), .QN(n12703) );
  NAND2X0 U12949 ( .IN1(n9107), .IN2(n12707), .QN(n12706) );
  NAND2X0 U12950 ( .IN1(n8412), .IN2(n9110), .QN(n12705) );
  NAND2X0 U12951 ( .IN1(n745), .IN2(n9282), .QN(n12686) );
  NOR2X0 U12952 ( .IN1(n9232), .IN2(n8960), .QN(n745) );
  NAND2X0 U12953 ( .IN1(n9293), .IN2(CRC_OUT_6_17), .QN(n12685) );
  NAND4X0 U12954 ( .IN1(n12708), .IN2(n12709), .IN3(n12710), .IN4(n12711), 
        .QN(WX4549) );
  NAND2X0 U12955 ( .IN1(n12712), .IN2(n12713), .QN(n12711) );
  NAND2X0 U12956 ( .IN1(n12714), .IN2(n12715), .QN(n12712) );
  NAND2X0 U12957 ( .IN1(n9107), .IN2(n12716), .QN(n12715) );
  NAND2X0 U12958 ( .IN1(n9107), .IN2(n8540), .QN(n12714) );
  NAND2X0 U12959 ( .IN1(n12035), .IN2(n2153), .QN(n12710) );
  NOR2X0 U12960 ( .IN1(n12717), .IN2(n12718), .QN(n12035) );
  INVX0 U12961 ( .INP(n12719), .ZN(n12718) );
  NAND2X0 U12962 ( .IN1(n12720), .IN2(n12721), .QN(n12719) );
  NOR2X0 U12963 ( .IN1(n12721), .IN2(n12720), .QN(n12717) );
  NAND2X0 U12964 ( .IN1(n12722), .IN2(n12723), .QN(n12720) );
  NAND2X0 U12965 ( .IN1(n8292), .IN2(n12724), .QN(n12723) );
  INVX0 U12966 ( .INP(n12725), .ZN(n12724) );
  NAND2X0 U12967 ( .IN1(n12725), .IN2(WX6035), .QN(n12722) );
  NAND2X0 U12968 ( .IN1(n12726), .IN2(n12727), .QN(n12725) );
  INVX0 U12969 ( .INP(n12728), .ZN(n12727) );
  NOR2X0 U12970 ( .IN1(n8811), .IN2(n16084), .QN(n12728) );
  NAND2X0 U12971 ( .IN1(n16084), .IN2(n8811), .QN(n12726) );
  NOR2X0 U12972 ( .IN1(n12729), .IN2(n12730), .QN(n12721) );
  INVX0 U12973 ( .INP(n12731), .ZN(n12730) );
  NAND2X0 U12974 ( .IN1(n7743), .IN2(n9117), .QN(n12731) );
  NOR2X0 U12975 ( .IN1(n9115), .IN2(n7743), .QN(n12729) );
  NAND2X0 U12976 ( .IN1(n744), .IN2(n9282), .QN(n12709) );
  NOR2X0 U12977 ( .IN1(n9232), .IN2(n8961), .QN(n744) );
  NAND2X0 U12978 ( .IN1(n9294), .IN2(CRC_OUT_6_18), .QN(n12708) );
  NAND4X0 U12979 ( .IN1(n12732), .IN2(n12733), .IN3(n12734), .IN4(n12735), 
        .QN(WX4547) );
  NAND2X0 U12980 ( .IN1(n12736), .IN2(n12055), .QN(n12735) );
  NAND2X0 U12981 ( .IN1(n12737), .IN2(n12058), .QN(n12055) );
  NAND2X0 U12982 ( .IN1(n12738), .IN2(n12739), .QN(n12737) );
  NAND2X0 U12983 ( .IN1(n16083), .IN2(n9118), .QN(n12739) );
  NAND2X0 U12984 ( .IN1(TM1), .IN2(n8482), .QN(n12738) );
  NAND3X0 U12985 ( .IN1(n12740), .IN2(n12741), .IN3(n12742), .QN(n12736) );
  NAND2X0 U12986 ( .IN1(n9324), .IN2(n12058), .QN(n12742) );
  NAND2X0 U12987 ( .IN1(n12743), .IN2(n12744), .QN(n12058) );
  NAND2X0 U12988 ( .IN1(n7744), .IN2(n12745), .QN(n12744) );
  INVX0 U12989 ( .INP(n12746), .ZN(n12743) );
  NOR2X0 U12990 ( .IN1(n12745), .IN2(n7744), .QN(n12746) );
  NOR2X0 U12991 ( .IN1(n12747), .IN2(n12748), .QN(n12745) );
  NOR2X0 U12992 ( .IN1(WX6033), .IN2(n7745), .QN(n12748) );
  INVX0 U12993 ( .INP(n12749), .ZN(n12747) );
  NAND2X0 U12994 ( .IN1(n7745), .IN2(WX6033), .QN(n12749) );
  NAND2X0 U12995 ( .IN1(n9790), .IN2(n8482), .QN(n12741) );
  NAND2X0 U12996 ( .IN1(n16083), .IN2(n9077), .QN(n12740) );
  NAND2X0 U12997 ( .IN1(n12750), .IN2(n12751), .QN(n12734) );
  NAND2X0 U12998 ( .IN1(n12752), .IN2(n12753), .QN(n12750) );
  NAND2X0 U12999 ( .IN1(n9107), .IN2(n12754), .QN(n12753) );
  NAND2X0 U13000 ( .IN1(n9107), .IN2(n8541), .QN(n12752) );
  NAND2X0 U13001 ( .IN1(n743), .IN2(n9282), .QN(n12733) );
  NOR2X0 U13002 ( .IN1(n9069), .IN2(n9160), .QN(n743) );
  NAND2X0 U13003 ( .IN1(n9294), .IN2(CRC_OUT_6_19), .QN(n12732) );
  NAND4X0 U13004 ( .IN1(n12755), .IN2(n12756), .IN3(n12757), .IN4(n12758), 
        .QN(WX4545) );
  NAND2X0 U13005 ( .IN1(n12759), .IN2(n12760), .QN(n12758) );
  NAND2X0 U13006 ( .IN1(n12761), .IN2(n12762), .QN(n12759) );
  NAND2X0 U13007 ( .IN1(n9107), .IN2(n12763), .QN(n12762) );
  NAND2X0 U13008 ( .IN1(n9107), .IN2(n8542), .QN(n12761) );
  NAND2X0 U13009 ( .IN1(n12077), .IN2(n2153), .QN(n12757) );
  NOR2X0 U13010 ( .IN1(n12764), .IN2(n12765), .QN(n12077) );
  INVX0 U13011 ( .INP(n12766), .ZN(n12765) );
  NAND2X0 U13012 ( .IN1(n12767), .IN2(n12768), .QN(n12766) );
  NOR2X0 U13013 ( .IN1(n12768), .IN2(n12767), .QN(n12764) );
  NAND2X0 U13014 ( .IN1(n12769), .IN2(n12770), .QN(n12767) );
  NAND2X0 U13015 ( .IN1(n8274), .IN2(n12771), .QN(n12770) );
  INVX0 U13016 ( .INP(n12772), .ZN(n12771) );
  NAND2X0 U13017 ( .IN1(n12772), .IN2(WX6031), .QN(n12769) );
  NAND2X0 U13018 ( .IN1(n12773), .IN2(n12774), .QN(n12772) );
  INVX0 U13019 ( .INP(n12775), .ZN(n12774) );
  NOR2X0 U13020 ( .IN1(n8812), .IN2(n16082), .QN(n12775) );
  NAND2X0 U13021 ( .IN1(n16082), .IN2(n8812), .QN(n12773) );
  NOR2X0 U13022 ( .IN1(n12776), .IN2(n12777), .QN(n12768) );
  INVX0 U13023 ( .INP(n12778), .ZN(n12777) );
  NAND2X0 U13024 ( .IN1(n7746), .IN2(n9117), .QN(n12778) );
  NOR2X0 U13025 ( .IN1(n9116), .IN2(n7746), .QN(n12776) );
  NAND2X0 U13026 ( .IN1(n742), .IN2(n9282), .QN(n12756) );
  NOR2X0 U13027 ( .IN1(n9233), .IN2(n8962), .QN(n742) );
  NAND2X0 U13028 ( .IN1(n9294), .IN2(CRC_OUT_6_20), .QN(n12755) );
  NAND4X0 U13029 ( .IN1(n12779), .IN2(n12780), .IN3(n12781), .IN4(n12782), 
        .QN(WX4543) );
  NAND2X0 U13030 ( .IN1(n12783), .IN2(n12083), .QN(n12782) );
  NAND2X0 U13031 ( .IN1(n12784), .IN2(n12086), .QN(n12083) );
  NAND2X0 U13032 ( .IN1(n12785), .IN2(n12786), .QN(n12784) );
  NAND2X0 U13033 ( .IN1(n16081), .IN2(n9117), .QN(n12786) );
  NAND2X0 U13034 ( .IN1(TM1), .IN2(n8484), .QN(n12785) );
  NAND3X0 U13035 ( .IN1(n12787), .IN2(n12788), .IN3(n12789), .QN(n12783) );
  NAND2X0 U13036 ( .IN1(n9324), .IN2(n12086), .QN(n12789) );
  NAND2X0 U13037 ( .IN1(n12790), .IN2(n12791), .QN(n12086) );
  NAND2X0 U13038 ( .IN1(n7747), .IN2(n12792), .QN(n12791) );
  INVX0 U13039 ( .INP(n12793), .ZN(n12790) );
  NOR2X0 U13040 ( .IN1(n12792), .IN2(n7747), .QN(n12793) );
  NOR2X0 U13041 ( .IN1(n12794), .IN2(n12795), .QN(n12792) );
  NOR2X0 U13042 ( .IN1(WX6029), .IN2(n7748), .QN(n12795) );
  INVX0 U13043 ( .INP(n12796), .ZN(n12794) );
  NAND2X0 U13044 ( .IN1(n7748), .IN2(WX6029), .QN(n12796) );
  NAND2X0 U13045 ( .IN1(n9083), .IN2(n8484), .QN(n12788) );
  NAND2X0 U13046 ( .IN1(n16081), .IN2(n9791), .QN(n12787) );
  NAND2X0 U13047 ( .IN1(n12797), .IN2(n12798), .QN(n12781) );
  NAND2X0 U13048 ( .IN1(n12799), .IN2(n12800), .QN(n12797) );
  NAND2X0 U13049 ( .IN1(n9107), .IN2(n12801), .QN(n12800) );
  NAND2X0 U13050 ( .IN1(n9107), .IN2(n8543), .QN(n12799) );
  NAND2X0 U13051 ( .IN1(n741), .IN2(n9282), .QN(n12780) );
  NOR2X0 U13052 ( .IN1(n9233), .IN2(n8963), .QN(n741) );
  NAND2X0 U13053 ( .IN1(n9294), .IN2(CRC_OUT_6_21), .QN(n12779) );
  NAND4X0 U13054 ( .IN1(n12802), .IN2(n12803), .IN3(n12804), .IN4(n12805), 
        .QN(WX4541) );
  NAND2X0 U13055 ( .IN1(n12806), .IN2(n12119), .QN(n12805) );
  NAND3X0 U13056 ( .IN1(n12807), .IN2(n12808), .IN3(n12122), .QN(n12119) );
  NAND2X0 U13057 ( .IN1(n8256), .IN2(n9118), .QN(n12808) );
  NAND2X0 U13058 ( .IN1(TM1), .IN2(WX6027), .QN(n12807) );
  NAND3X0 U13059 ( .IN1(n12809), .IN2(n12810), .IN3(n12811), .QN(n12806) );
  NAND2X0 U13060 ( .IN1(n9324), .IN2(n12122), .QN(n12811) );
  NAND2X0 U13061 ( .IN1(n12812), .IN2(n12813), .QN(n12122) );
  NAND2X0 U13062 ( .IN1(n12814), .IN2(WX5963), .QN(n12813) );
  NAND2X0 U13063 ( .IN1(n12815), .IN2(n12816), .QN(n12814) );
  NAND3X0 U13064 ( .IN1(n12815), .IN2(n12816), .IN3(n7750), .QN(n12812) );
  NAND2X0 U13065 ( .IN1(test_so46), .IN2(WX5899), .QN(n12816) );
  NAND2X0 U13066 ( .IN1(n7749), .IN2(n8821), .QN(n12815) );
  NAND2X0 U13067 ( .IN1(n9791), .IN2(WX6027), .QN(n12810) );
  NAND2X0 U13068 ( .IN1(n9082), .IN2(n8256), .QN(n12809) );
  NAND2X0 U13069 ( .IN1(n12817), .IN2(n12818), .QN(n12804) );
  NAND2X0 U13070 ( .IN1(n12819), .IN2(n12820), .QN(n12817) );
  NAND2X0 U13071 ( .IN1(n9107), .IN2(n12821), .QN(n12820) );
  NAND2X0 U13072 ( .IN1(n9107), .IN2(n8544), .QN(n12819) );
  NAND2X0 U13073 ( .IN1(n740), .IN2(n9282), .QN(n12803) );
  NOR2X0 U13074 ( .IN1(n9233), .IN2(n8964), .QN(n740) );
  NAND2X0 U13075 ( .IN1(test_so43), .IN2(n9313), .QN(n12802) );
  NAND4X0 U13076 ( .IN1(n12822), .IN2(n12823), .IN3(n12824), .IN4(n12825), 
        .QN(WX4539) );
  NAND2X0 U13077 ( .IN1(n12826), .IN2(n12128), .QN(n12825) );
  NAND2X0 U13078 ( .IN1(n12827), .IN2(n12131), .QN(n12128) );
  NAND2X0 U13079 ( .IN1(n12828), .IN2(n12829), .QN(n12827) );
  NAND2X0 U13080 ( .IN1(n16080), .IN2(n9117), .QN(n12829) );
  NAND2X0 U13081 ( .IN1(TM1), .IN2(n8487), .QN(n12828) );
  NAND3X0 U13082 ( .IN1(n12830), .IN2(n12831), .IN3(n12832), .QN(n12826) );
  NAND2X0 U13083 ( .IN1(n9324), .IN2(n12131), .QN(n12832) );
  NAND2X0 U13084 ( .IN1(n12833), .IN2(n12834), .QN(n12131) );
  NAND2X0 U13085 ( .IN1(n7751), .IN2(n12835), .QN(n12834) );
  INVX0 U13086 ( .INP(n12836), .ZN(n12833) );
  NOR2X0 U13087 ( .IN1(n12835), .IN2(n7751), .QN(n12836) );
  NOR2X0 U13088 ( .IN1(n12837), .IN2(n12838), .QN(n12835) );
  NOR2X0 U13089 ( .IN1(WX6025), .IN2(n7752), .QN(n12838) );
  INVX0 U13090 ( .INP(n12839), .ZN(n12837) );
  NAND2X0 U13091 ( .IN1(n7752), .IN2(WX6025), .QN(n12839) );
  NAND2X0 U13092 ( .IN1(n9081), .IN2(n8487), .QN(n12831) );
  NAND2X0 U13093 ( .IN1(n16080), .IN2(n9079), .QN(n12830) );
  NAND2X0 U13094 ( .IN1(n12840), .IN2(n12841), .QN(n12824) );
  NAND2X0 U13095 ( .IN1(n12842), .IN2(n12843), .QN(n12840) );
  NAND2X0 U13096 ( .IN1(n9107), .IN2(n12844), .QN(n12843) );
  NAND2X0 U13097 ( .IN1(n9107), .IN2(n8545), .QN(n12842) );
  NAND2X0 U13098 ( .IN1(n739), .IN2(n9282), .QN(n12823) );
  NOR2X0 U13099 ( .IN1(n9233), .IN2(n8965), .QN(n739) );
  NAND2X0 U13100 ( .IN1(n9294), .IN2(CRC_OUT_6_23), .QN(n12822) );
  NAND4X0 U13101 ( .IN1(n12845), .IN2(n12846), .IN3(n12847), .IN4(n12848), 
        .QN(WX4537) );
  NAND2X0 U13102 ( .IN1(n12849), .IN2(n12166), .QN(n12848) );
  NAND2X0 U13103 ( .IN1(n12850), .IN2(n12169), .QN(n12166) );
  NAND2X0 U13104 ( .IN1(n12851), .IN2(n12852), .QN(n12850) );
  NAND2X0 U13105 ( .IN1(n16079), .IN2(n9117), .QN(n12852) );
  NAND2X0 U13106 ( .IN1(TM1), .IN2(n8488), .QN(n12851) );
  NAND3X0 U13107 ( .IN1(n12853), .IN2(n12854), .IN3(n12855), .QN(n12849) );
  NAND2X0 U13108 ( .IN1(n9324), .IN2(n12169), .QN(n12855) );
  NAND2X0 U13109 ( .IN1(n12856), .IN2(n12857), .QN(n12169) );
  NAND2X0 U13110 ( .IN1(n7753), .IN2(n12858), .QN(n12857) );
  INVX0 U13111 ( .INP(n12859), .ZN(n12856) );
  NOR2X0 U13112 ( .IN1(n12858), .IN2(n7753), .QN(n12859) );
  NOR2X0 U13113 ( .IN1(n12860), .IN2(n12861), .QN(n12858) );
  NOR2X0 U13114 ( .IN1(WX6023), .IN2(n7754), .QN(n12861) );
  INVX0 U13115 ( .INP(n12862), .ZN(n12860) );
  NAND2X0 U13116 ( .IN1(n7754), .IN2(WX6023), .QN(n12862) );
  NAND2X0 U13117 ( .IN1(n9790), .IN2(n8488), .QN(n12854) );
  NAND2X0 U13118 ( .IN1(n16079), .IN2(n9078), .QN(n12853) );
  NAND2X0 U13119 ( .IN1(n12863), .IN2(n12864), .QN(n12847) );
  NAND2X0 U13120 ( .IN1(n12865), .IN2(n12866), .QN(n12863) );
  NAND2X0 U13121 ( .IN1(n9107), .IN2(n12867), .QN(n12866) );
  NAND2X0 U13122 ( .IN1(n9107), .IN2(n8546), .QN(n12865) );
  NAND2X0 U13123 ( .IN1(n738), .IN2(n9282), .QN(n12846) );
  NOR2X0 U13124 ( .IN1(n9233), .IN2(n8966), .QN(n738) );
  NAND2X0 U13125 ( .IN1(n9294), .IN2(CRC_OUT_6_24), .QN(n12845) );
  NAND4X0 U13126 ( .IN1(n12868), .IN2(n12869), .IN3(n12870), .IN4(n12871), 
        .QN(WX4535) );
  NAND2X0 U13127 ( .IN1(n12872), .IN2(n12175), .QN(n12871) );
  NAND2X0 U13128 ( .IN1(n12873), .IN2(n12178), .QN(n12175) );
  NAND2X0 U13129 ( .IN1(n12874), .IN2(n12875), .QN(n12873) );
  NAND2X0 U13130 ( .IN1(n16078), .IN2(n9117), .QN(n12875) );
  NAND2X0 U13131 ( .IN1(TM1), .IN2(n8489), .QN(n12874) );
  NAND3X0 U13132 ( .IN1(n12876), .IN2(n12877), .IN3(n12878), .QN(n12872) );
  NAND2X0 U13133 ( .IN1(n9324), .IN2(n12178), .QN(n12878) );
  NAND2X0 U13134 ( .IN1(n12879), .IN2(n12880), .QN(n12178) );
  NAND2X0 U13135 ( .IN1(n7755), .IN2(n12881), .QN(n12880) );
  INVX0 U13136 ( .INP(n12882), .ZN(n12879) );
  NOR2X0 U13137 ( .IN1(n12881), .IN2(n7755), .QN(n12882) );
  NOR2X0 U13138 ( .IN1(n12883), .IN2(n12884), .QN(n12881) );
  NOR2X0 U13139 ( .IN1(WX6021), .IN2(n7756), .QN(n12884) );
  INVX0 U13140 ( .INP(n12885), .ZN(n12883) );
  NAND2X0 U13141 ( .IN1(n7756), .IN2(WX6021), .QN(n12885) );
  NAND2X0 U13142 ( .IN1(n9083), .IN2(n8489), .QN(n12877) );
  NAND2X0 U13143 ( .IN1(n16078), .IN2(n9077), .QN(n12876) );
  NAND2X0 U13144 ( .IN1(n12886), .IN2(n12887), .QN(n12870) );
  NAND2X0 U13145 ( .IN1(n12888), .IN2(n12889), .QN(n12886) );
  NAND2X0 U13146 ( .IN1(n9107), .IN2(n12890), .QN(n12889) );
  NAND2X0 U13147 ( .IN1(n9107), .IN2(n8547), .QN(n12888) );
  NAND2X0 U13148 ( .IN1(n737), .IN2(n9282), .QN(n12869) );
  NOR2X0 U13149 ( .IN1(n9233), .IN2(n8967), .QN(n737) );
  NAND2X0 U13150 ( .IN1(n9294), .IN2(CRC_OUT_6_25), .QN(n12868) );
  NAND4X0 U13151 ( .IN1(n12891), .IN2(n12892), .IN3(n12893), .IN4(n12894), 
        .QN(WX4533) );
  NAND2X0 U13152 ( .IN1(n12895), .IN2(n12213), .QN(n12894) );
  NAND2X0 U13153 ( .IN1(n12896), .IN2(n12216), .QN(n12213) );
  NAND2X0 U13154 ( .IN1(n12897), .IN2(n12898), .QN(n12896) );
  NAND2X0 U13155 ( .IN1(n16077), .IN2(n9117), .QN(n12898) );
  NAND2X0 U13156 ( .IN1(TM1), .IN2(n8490), .QN(n12897) );
  NAND3X0 U13157 ( .IN1(n12899), .IN2(n12900), .IN3(n12901), .QN(n12895) );
  NAND2X0 U13158 ( .IN1(n9324), .IN2(n12216), .QN(n12901) );
  NAND2X0 U13159 ( .IN1(n12902), .IN2(n12903), .QN(n12216) );
  NAND2X0 U13160 ( .IN1(n7757), .IN2(n12904), .QN(n12903) );
  INVX0 U13161 ( .INP(n12905), .ZN(n12902) );
  NOR2X0 U13162 ( .IN1(n12904), .IN2(n7757), .QN(n12905) );
  NOR2X0 U13163 ( .IN1(n12906), .IN2(n12907), .QN(n12904) );
  NOR2X0 U13164 ( .IN1(WX6019), .IN2(n7758), .QN(n12907) );
  INVX0 U13165 ( .INP(n12908), .ZN(n12906) );
  NAND2X0 U13166 ( .IN1(n7758), .IN2(WX6019), .QN(n12908) );
  NAND2X0 U13167 ( .IN1(n9082), .IN2(n8490), .QN(n12900) );
  NAND2X0 U13168 ( .IN1(n16077), .IN2(n9791), .QN(n12899) );
  NAND2X0 U13169 ( .IN1(n12909), .IN2(n12910), .QN(n12893) );
  NAND2X0 U13170 ( .IN1(n12911), .IN2(n12912), .QN(n12909) );
  NAND2X0 U13171 ( .IN1(n9108), .IN2(n12913), .QN(n12912) );
  NAND2X0 U13172 ( .IN1(n9108), .IN2(n8548), .QN(n12911) );
  NAND2X0 U13173 ( .IN1(n736), .IN2(n9282), .QN(n12892) );
  NOR2X0 U13174 ( .IN1(n9233), .IN2(n8968), .QN(n736) );
  NAND2X0 U13175 ( .IN1(n9294), .IN2(CRC_OUT_6_26), .QN(n12891) );
  NAND4X0 U13176 ( .IN1(n12914), .IN2(n12915), .IN3(n12916), .IN4(n12917), 
        .QN(WX4531) );
  NAND2X0 U13177 ( .IN1(n12918), .IN2(n12233), .QN(n12917) );
  NAND2X0 U13178 ( .IN1(n12919), .IN2(n12236), .QN(n12233) );
  NAND2X0 U13179 ( .IN1(n12920), .IN2(n12921), .QN(n12919) );
  NAND2X0 U13180 ( .IN1(n16076), .IN2(n9118), .QN(n12921) );
  NAND2X0 U13181 ( .IN1(TM1), .IN2(n8491), .QN(n12920) );
  NAND3X0 U13182 ( .IN1(n12922), .IN2(n12923), .IN3(n12924), .QN(n12918) );
  NAND2X0 U13183 ( .IN1(n9324), .IN2(n12236), .QN(n12924) );
  NAND2X0 U13184 ( .IN1(n12925), .IN2(n12926), .QN(n12236) );
  NAND2X0 U13185 ( .IN1(n7759), .IN2(n12927), .QN(n12926) );
  INVX0 U13186 ( .INP(n12928), .ZN(n12925) );
  NOR2X0 U13187 ( .IN1(n12927), .IN2(n7759), .QN(n12928) );
  NOR2X0 U13188 ( .IN1(n12929), .IN2(n12930), .QN(n12927) );
  NOR2X0 U13189 ( .IN1(WX6017), .IN2(n7760), .QN(n12930) );
  INVX0 U13190 ( .INP(n12931), .ZN(n12929) );
  NAND2X0 U13191 ( .IN1(n7760), .IN2(WX6017), .QN(n12931) );
  NAND2X0 U13192 ( .IN1(n9081), .IN2(n8491), .QN(n12923) );
  NAND2X0 U13193 ( .IN1(n16076), .IN2(n9079), .QN(n12922) );
  NAND2X0 U13194 ( .IN1(n12932), .IN2(n12933), .QN(n12916) );
  NAND2X0 U13195 ( .IN1(n12934), .IN2(n12935), .QN(n12932) );
  NAND2X0 U13196 ( .IN1(n9108), .IN2(n12936), .QN(n12935) );
  NAND2X0 U13197 ( .IN1(n9108), .IN2(n8549), .QN(n12934) );
  NAND2X0 U13198 ( .IN1(n735), .IN2(n9282), .QN(n12915) );
  NOR2X0 U13199 ( .IN1(n9233), .IN2(n8969), .QN(n735) );
  NAND2X0 U13200 ( .IN1(n9294), .IN2(CRC_OUT_6_27), .QN(n12914) );
  NAND4X0 U13201 ( .IN1(n12937), .IN2(n12938), .IN3(n12939), .IN4(n12940), 
        .QN(WX4529) );
  NAND2X0 U13202 ( .IN1(n12941), .IN2(n12256), .QN(n12940) );
  NAND2X0 U13203 ( .IN1(n12942), .IN2(n12259), .QN(n12256) );
  NAND2X0 U13204 ( .IN1(n12943), .IN2(n12944), .QN(n12942) );
  NAND2X0 U13205 ( .IN1(n16075), .IN2(n9117), .QN(n12944) );
  NAND2X0 U13206 ( .IN1(TM1), .IN2(n8492), .QN(n12943) );
  NAND3X0 U13207 ( .IN1(n12945), .IN2(n12946), .IN3(n12947), .QN(n12941) );
  NAND2X0 U13208 ( .IN1(n9324), .IN2(n12259), .QN(n12947) );
  NAND2X0 U13209 ( .IN1(n12948), .IN2(n12949), .QN(n12259) );
  NAND2X0 U13210 ( .IN1(n7761), .IN2(n12950), .QN(n12949) );
  INVX0 U13211 ( .INP(n12951), .ZN(n12948) );
  NOR2X0 U13212 ( .IN1(n12950), .IN2(n7761), .QN(n12951) );
  NOR2X0 U13213 ( .IN1(n12952), .IN2(n12953), .QN(n12950) );
  NOR2X0 U13214 ( .IN1(WX6015), .IN2(n7762), .QN(n12953) );
  INVX0 U13215 ( .INP(n12954), .ZN(n12952) );
  NAND2X0 U13216 ( .IN1(n7762), .IN2(WX6015), .QN(n12954) );
  NAND2X0 U13217 ( .IN1(n9790), .IN2(n8492), .QN(n12946) );
  NAND2X0 U13218 ( .IN1(n16075), .IN2(n9078), .QN(n12945) );
  NAND2X0 U13219 ( .IN1(n12955), .IN2(n9110), .QN(n12939) );
  NAND2X0 U13220 ( .IN1(n734), .IN2(n9282), .QN(n12938) );
  NOR2X0 U13221 ( .IN1(n9233), .IN2(n8970), .QN(n734) );
  NAND2X0 U13222 ( .IN1(n9294), .IN2(CRC_OUT_6_28), .QN(n12937) );
  NAND4X0 U13223 ( .IN1(n12956), .IN2(n12957), .IN3(n12958), .IN4(n12959), 
        .QN(WX4527) );
  NAND2X0 U13224 ( .IN1(n12960), .IN2(n12279), .QN(n12959) );
  NAND2X0 U13225 ( .IN1(n12961), .IN2(n12282), .QN(n12279) );
  NAND2X0 U13226 ( .IN1(n12962), .IN2(n12963), .QN(n12961) );
  NAND2X0 U13227 ( .IN1(n16074), .IN2(n9117), .QN(n12963) );
  NAND2X0 U13228 ( .IN1(TM1), .IN2(n8493), .QN(n12962) );
  NAND3X0 U13229 ( .IN1(n12964), .IN2(n12965), .IN3(n12966), .QN(n12960) );
  NAND2X0 U13230 ( .IN1(n9325), .IN2(n12282), .QN(n12966) );
  NAND2X0 U13231 ( .IN1(n12967), .IN2(n12968), .QN(n12282) );
  NAND2X0 U13232 ( .IN1(n7763), .IN2(n12969), .QN(n12968) );
  INVX0 U13233 ( .INP(n12970), .ZN(n12967) );
  NOR2X0 U13234 ( .IN1(n12969), .IN2(n7763), .QN(n12970) );
  NOR2X0 U13235 ( .IN1(n12971), .IN2(n12972), .QN(n12969) );
  NOR2X0 U13236 ( .IN1(WX6013), .IN2(n7764), .QN(n12972) );
  INVX0 U13237 ( .INP(n12973), .ZN(n12971) );
  NAND2X0 U13238 ( .IN1(n7764), .IN2(WX6013), .QN(n12973) );
  NAND2X0 U13239 ( .IN1(n9083), .IN2(n8493), .QN(n12965) );
  NAND2X0 U13240 ( .IN1(n16074), .IN2(n9077), .QN(n12964) );
  NAND2X0 U13241 ( .IN1(n12974), .IN2(n12975), .QN(n12958) );
  NAND2X0 U13242 ( .IN1(n12976), .IN2(n12977), .QN(n12974) );
  NAND2X0 U13243 ( .IN1(n9108), .IN2(n12978), .QN(n12977) );
  NAND2X0 U13244 ( .IN1(n9108), .IN2(n8551), .QN(n12976) );
  NAND2X0 U13245 ( .IN1(n733), .IN2(n9282), .QN(n12957) );
  NOR2X0 U13246 ( .IN1(n9233), .IN2(n8971), .QN(n733) );
  NAND2X0 U13247 ( .IN1(n9294), .IN2(CRC_OUT_6_29), .QN(n12956) );
  NAND4X0 U13248 ( .IN1(n12979), .IN2(n12980), .IN3(n12981), .IN4(n12982), 
        .QN(WX4525) );
  NAND2X0 U13249 ( .IN1(n12983), .IN2(n12302), .QN(n12982) );
  NAND2X0 U13250 ( .IN1(n12984), .IN2(n12305), .QN(n12302) );
  NAND2X0 U13251 ( .IN1(n12985), .IN2(n12986), .QN(n12984) );
  NAND2X0 U13252 ( .IN1(n16073), .IN2(n9118), .QN(n12986) );
  NAND2X0 U13253 ( .IN1(TM1), .IN2(n8494), .QN(n12985) );
  NAND3X0 U13254 ( .IN1(n12987), .IN2(n12988), .IN3(n12989), .QN(n12983) );
  NAND2X0 U13255 ( .IN1(n9325), .IN2(n12305), .QN(n12989) );
  NAND2X0 U13256 ( .IN1(n12990), .IN2(n12991), .QN(n12305) );
  NAND2X0 U13257 ( .IN1(n7765), .IN2(n12992), .QN(n12991) );
  INVX0 U13258 ( .INP(n12993), .ZN(n12990) );
  NOR2X0 U13259 ( .IN1(n12992), .IN2(n7765), .QN(n12993) );
  NOR2X0 U13260 ( .IN1(n12994), .IN2(n12995), .QN(n12992) );
  NOR2X0 U13261 ( .IN1(WX6011), .IN2(n7766), .QN(n12995) );
  INVX0 U13262 ( .INP(n12996), .ZN(n12994) );
  NAND2X0 U13263 ( .IN1(n7766), .IN2(WX6011), .QN(n12996) );
  NAND2X0 U13264 ( .IN1(n9082), .IN2(n8494), .QN(n12988) );
  NAND2X0 U13265 ( .IN1(n16073), .IN2(n9791), .QN(n12987) );
  NAND2X0 U13266 ( .IN1(n12997), .IN2(n9109), .QN(n12981) );
  NAND2X0 U13267 ( .IN1(n732), .IN2(n9282), .QN(n12980) );
  NOR2X0 U13268 ( .IN1(n9233), .IN2(n8972), .QN(n732) );
  NAND2X0 U13269 ( .IN1(n9294), .IN2(CRC_OUT_6_30), .QN(n12979) );
  NAND4X0 U13270 ( .IN1(n12998), .IN2(n12999), .IN3(n13000), .IN4(n13001), 
        .QN(WX4523) );
  NAND2X0 U13271 ( .IN1(n13002), .IN2(n12325), .QN(n13001) );
  NAND2X0 U13272 ( .IN1(n13003), .IN2(n12328), .QN(n12325) );
  NAND2X0 U13273 ( .IN1(n13004), .IN2(n13005), .QN(n13003) );
  NAND2X0 U13274 ( .IN1(n16072), .IN2(n9118), .QN(n13005) );
  NAND2X0 U13275 ( .IN1(TM1), .IN2(n8495), .QN(n13004) );
  NAND3X0 U13276 ( .IN1(n13006), .IN2(n13007), .IN3(n13008), .QN(n13002) );
  NAND2X0 U13277 ( .IN1(n9325), .IN2(n12328), .QN(n13008) );
  NAND2X0 U13278 ( .IN1(n13009), .IN2(n13010), .QN(n12328) );
  NAND2X0 U13279 ( .IN1(n7619), .IN2(n13011), .QN(n13010) );
  INVX0 U13280 ( .INP(n13012), .ZN(n13009) );
  NOR2X0 U13281 ( .IN1(n13011), .IN2(n7619), .QN(n13012) );
  NOR2X0 U13282 ( .IN1(n13013), .IN2(n13014), .QN(n13011) );
  NOR2X0 U13283 ( .IN1(WX6009), .IN2(n7620), .QN(n13014) );
  INVX0 U13284 ( .INP(n13015), .ZN(n13013) );
  NAND2X0 U13285 ( .IN1(n7620), .IN2(WX6009), .QN(n13015) );
  NAND2X0 U13286 ( .IN1(n9081), .IN2(n8495), .QN(n13007) );
  NAND2X0 U13287 ( .IN1(n16072), .IN2(n9079), .QN(n13006) );
  NAND2X0 U13288 ( .IN1(n13016), .IN2(n13017), .QN(n13000) );
  NAND2X0 U13289 ( .IN1(n13018), .IN2(n13019), .QN(n13016) );
  NAND2X0 U13290 ( .IN1(n9108), .IN2(n13020), .QN(n13019) );
  NAND2X0 U13291 ( .IN1(n9108), .IN2(n8553), .QN(n13018) );
  NAND2X0 U13292 ( .IN1(n9295), .IN2(CRC_OUT_6_31), .QN(n12999) );
  NAND2X0 U13293 ( .IN1(n2245), .IN2(WX4364), .QN(n12998) );
  NOR2X0 U13294 ( .IN1(n9233), .IN2(WX4364), .QN(WX4425) );
  NOR3X0 U13295 ( .IN1(n9137), .IN2(n13021), .IN3(n13022), .QN(WX3912) );
  NOR2X0 U13296 ( .IN1(n8469), .IN2(CRC_OUT_7_30), .QN(n13022) );
  NOR2X0 U13297 ( .IN1(DFF_574_n1), .IN2(WX3423), .QN(n13021) );
  NOR3X0 U13298 ( .IN1(n9137), .IN2(n13023), .IN3(n13024), .QN(WX3910) );
  NOR2X0 U13299 ( .IN1(n8471), .IN2(CRC_OUT_7_29), .QN(n13024) );
  NOR2X0 U13300 ( .IN1(DFF_573_n1), .IN2(WX3425), .QN(n13023) );
  NOR3X0 U13301 ( .IN1(n9137), .IN2(n13025), .IN3(n13026), .QN(WX3908) );
  NOR2X0 U13302 ( .IN1(n8472), .IN2(CRC_OUT_7_28), .QN(n13026) );
  NOR2X0 U13303 ( .IN1(DFF_572_n1), .IN2(WX3427), .QN(n13025) );
  NOR2X0 U13304 ( .IN1(n9234), .IN2(n13027), .QN(WX3906) );
  NOR2X0 U13305 ( .IN1(n13028), .IN2(n13029), .QN(n13027) );
  NOR2X0 U13306 ( .IN1(test_so32), .IN2(WX3429), .QN(n13029) );
  INVX0 U13307 ( .INP(n13030), .ZN(n13028) );
  NAND2X0 U13308 ( .IN1(WX3429), .IN2(test_so32), .QN(n13030) );
  NOR3X0 U13309 ( .IN1(n9137), .IN2(n13031), .IN3(n13032), .QN(WX3904) );
  NOR2X0 U13310 ( .IN1(n8474), .IN2(CRC_OUT_7_26), .QN(n13032) );
  NOR2X0 U13311 ( .IN1(DFF_570_n1), .IN2(WX3431), .QN(n13031) );
  NOR3X0 U13312 ( .IN1(n9137), .IN2(n13033), .IN3(n13034), .QN(WX3902) );
  NOR2X0 U13313 ( .IN1(n8475), .IN2(CRC_OUT_7_25), .QN(n13034) );
  NOR2X0 U13314 ( .IN1(DFF_569_n1), .IN2(WX3433), .QN(n13033) );
  NOR3X0 U13315 ( .IN1(n9137), .IN2(n13035), .IN3(n13036), .QN(WX3900) );
  NOR2X0 U13316 ( .IN1(n8476), .IN2(CRC_OUT_7_24), .QN(n13036) );
  NOR2X0 U13317 ( .IN1(DFF_568_n1), .IN2(WX3435), .QN(n13035) );
  NOR3X0 U13318 ( .IN1(n9136), .IN2(n13037), .IN3(n13038), .QN(WX3898) );
  NOR2X0 U13319 ( .IN1(n8477), .IN2(CRC_OUT_7_23), .QN(n13038) );
  NOR2X0 U13320 ( .IN1(DFF_567_n1), .IN2(WX3437), .QN(n13037) );
  NOR2X0 U13321 ( .IN1(n9234), .IN2(n13039), .QN(WX3896) );
  NOR2X0 U13322 ( .IN1(n13040), .IN2(n13041), .QN(n13039) );
  NOR2X0 U13323 ( .IN1(test_so29), .IN2(CRC_OUT_7_22), .QN(n13041) );
  NOR2X0 U13324 ( .IN1(DFF_566_n1), .IN2(n8801), .QN(n13040) );
  NOR3X0 U13325 ( .IN1(n9136), .IN2(n13042), .IN3(n13043), .QN(WX3894) );
  NOR2X0 U13326 ( .IN1(n8478), .IN2(CRC_OUT_7_21), .QN(n13043) );
  NOR2X0 U13327 ( .IN1(DFF_565_n1), .IN2(WX3441), .QN(n13042) );
  NOR3X0 U13328 ( .IN1(n9136), .IN2(n13044), .IN3(n13045), .QN(WX3892) );
  NOR2X0 U13329 ( .IN1(n8485), .IN2(CRC_OUT_7_20), .QN(n13045) );
  NOR2X0 U13330 ( .IN1(DFF_564_n1), .IN2(WX3443), .QN(n13044) );
  NOR3X0 U13331 ( .IN1(n9136), .IN2(n13046), .IN3(n13047), .QN(WX3890) );
  NOR2X0 U13332 ( .IN1(n8486), .IN2(CRC_OUT_7_19), .QN(n13047) );
  NOR2X0 U13333 ( .IN1(DFF_563_n1), .IN2(WX3445), .QN(n13046) );
  NOR3X0 U13334 ( .IN1(n9136), .IN2(n13048), .IN3(n13049), .QN(WX3888) );
  NOR2X0 U13335 ( .IN1(n8503), .IN2(CRC_OUT_7_18), .QN(n13049) );
  NOR2X0 U13336 ( .IN1(DFF_562_n1), .IN2(WX3447), .QN(n13048) );
  NOR3X0 U13337 ( .IN1(n9136), .IN2(n13050), .IN3(n13051), .QN(WX3886) );
  NOR2X0 U13338 ( .IN1(n8504), .IN2(CRC_OUT_7_17), .QN(n13051) );
  NOR2X0 U13339 ( .IN1(DFF_561_n1), .IN2(WX3449), .QN(n13050) );
  NOR3X0 U13340 ( .IN1(n9136), .IN2(n13052), .IN3(n13053), .QN(WX3884) );
  NOR2X0 U13341 ( .IN1(n8521), .IN2(CRC_OUT_7_16), .QN(n13053) );
  NOR2X0 U13342 ( .IN1(DFF_560_n1), .IN2(WX3451), .QN(n13052) );
  NOR2X0 U13343 ( .IN1(n9234), .IN2(n13054), .QN(WX3882) );
  NOR2X0 U13344 ( .IN1(n13055), .IN2(n13056), .QN(n13054) );
  INVX0 U13345 ( .INP(n13057), .ZN(n13056) );
  NAND2X0 U13346 ( .IN1(CRC_OUT_7_15), .IN2(n13058), .QN(n13057) );
  NOR2X0 U13347 ( .IN1(n13058), .IN2(CRC_OUT_7_15), .QN(n13055) );
  NAND2X0 U13348 ( .IN1(n13059), .IN2(n13060), .QN(n13058) );
  NAND2X0 U13349 ( .IN1(n8119), .IN2(CRC_OUT_7_31), .QN(n13060) );
  NAND2X0 U13350 ( .IN1(DFF_575_n1), .IN2(WX3453), .QN(n13059) );
  NOR3X0 U13351 ( .IN1(n9136), .IN2(n13061), .IN3(n13062), .QN(WX3880) );
  NOR2X0 U13352 ( .IN1(n8522), .IN2(CRC_OUT_7_14), .QN(n13062) );
  NOR2X0 U13353 ( .IN1(DFF_558_n1), .IN2(WX3455), .QN(n13061) );
  NOR3X0 U13354 ( .IN1(n9136), .IN2(n13063), .IN3(n13064), .QN(WX3878) );
  NOR2X0 U13355 ( .IN1(n8529), .IN2(CRC_OUT_7_13), .QN(n13064) );
  NOR2X0 U13356 ( .IN1(DFF_557_n1), .IN2(WX3457), .QN(n13063) );
  NOR3X0 U13357 ( .IN1(n9136), .IN2(n13065), .IN3(n13066), .QN(WX3876) );
  NOR2X0 U13358 ( .IN1(n8530), .IN2(CRC_OUT_7_12), .QN(n13066) );
  NOR2X0 U13359 ( .IN1(DFF_556_n1), .IN2(WX3459), .QN(n13065) );
  NOR3X0 U13360 ( .IN1(n9136), .IN2(n13067), .IN3(n13068), .QN(WX3874) );
  NOR2X0 U13361 ( .IN1(n8531), .IN2(CRC_OUT_7_11), .QN(n13068) );
  NOR2X0 U13362 ( .IN1(DFF_555_n1), .IN2(WX3461), .QN(n13067) );
  NOR3X0 U13363 ( .IN1(n9136), .IN2(n13069), .IN3(n13070), .QN(WX3872) );
  NOR2X0 U13364 ( .IN1(DFF_575_n1), .IN2(n13071), .QN(n13070) );
  INVX0 U13365 ( .INP(n13072), .ZN(n13069) );
  NAND2X0 U13366 ( .IN1(n13071), .IN2(DFF_575_n1), .QN(n13072) );
  NOR2X0 U13367 ( .IN1(n13073), .IN2(n13074), .QN(n13071) );
  INVX0 U13368 ( .INP(n13075), .ZN(n13074) );
  NAND2X0 U13369 ( .IN1(test_so31), .IN2(WX3463), .QN(n13075) );
  NOR2X0 U13370 ( .IN1(WX3463), .IN2(test_so31), .QN(n13073) );
  NOR3X0 U13371 ( .IN1(n9135), .IN2(n13076), .IN3(n13077), .QN(WX3870) );
  NOR2X0 U13372 ( .IN1(n8532), .IN2(CRC_OUT_7_9), .QN(n13077) );
  NOR2X0 U13373 ( .IN1(DFF_553_n1), .IN2(WX3465), .QN(n13076) );
  NOR3X0 U13374 ( .IN1(n9135), .IN2(n13078), .IN3(n13079), .QN(WX3868) );
  NOR2X0 U13375 ( .IN1(n8533), .IN2(CRC_OUT_7_8), .QN(n13079) );
  NOR2X0 U13376 ( .IN1(DFF_552_n1), .IN2(WX3467), .QN(n13078) );
  NOR3X0 U13377 ( .IN1(n9135), .IN2(n13080), .IN3(n13081), .QN(WX3866) );
  NOR2X0 U13378 ( .IN1(n8534), .IN2(CRC_OUT_7_7), .QN(n13081) );
  NOR2X0 U13379 ( .IN1(DFF_551_n1), .IN2(WX3469), .QN(n13080) );
  NOR3X0 U13380 ( .IN1(n9135), .IN2(n13082), .IN3(n13083), .QN(WX3864) );
  NOR2X0 U13381 ( .IN1(n8535), .IN2(CRC_OUT_7_6), .QN(n13083) );
  NOR2X0 U13382 ( .IN1(DFF_550_n1), .IN2(WX3471), .QN(n13082) );
  NOR2X0 U13383 ( .IN1(n9235), .IN2(n13084), .QN(WX3862) );
  NOR2X0 U13384 ( .IN1(n13085), .IN2(n13086), .QN(n13084) );
  NOR2X0 U13385 ( .IN1(test_so30), .IN2(CRC_OUT_7_5), .QN(n13086) );
  NOR2X0 U13386 ( .IN1(DFF_549_n1), .IN2(n8791), .QN(n13085) );
  NOR3X0 U13387 ( .IN1(n9135), .IN2(n13087), .IN3(n13088), .QN(WX3860) );
  NOR2X0 U13388 ( .IN1(n8536), .IN2(CRC_OUT_7_4), .QN(n13088) );
  NOR2X0 U13389 ( .IN1(DFF_548_n1), .IN2(WX3475), .QN(n13087) );
  NOR2X0 U13390 ( .IN1(n9235), .IN2(n13089), .QN(WX3858) );
  NOR2X0 U13391 ( .IN1(n13090), .IN2(n13091), .QN(n13089) );
  INVX0 U13392 ( .INP(n13092), .ZN(n13091) );
  NAND2X0 U13393 ( .IN1(CRC_OUT_7_3), .IN2(n13093), .QN(n13092) );
  NOR2X0 U13394 ( .IN1(n13093), .IN2(CRC_OUT_7_3), .QN(n13090) );
  NAND2X0 U13395 ( .IN1(n13094), .IN2(n13095), .QN(n13093) );
  NAND2X0 U13396 ( .IN1(n8121), .IN2(CRC_OUT_7_31), .QN(n13095) );
  NAND2X0 U13397 ( .IN1(DFF_575_n1), .IN2(WX3477), .QN(n13094) );
  NOR3X0 U13398 ( .IN1(n9135), .IN2(n13096), .IN3(n13097), .QN(WX3856) );
  NOR2X0 U13399 ( .IN1(n8538), .IN2(CRC_OUT_7_2), .QN(n13097) );
  NOR2X0 U13400 ( .IN1(DFF_546_n1), .IN2(WX3479), .QN(n13096) );
  NOR3X0 U13401 ( .IN1(n9135), .IN2(n13098), .IN3(n13099), .QN(WX3854) );
  NOR2X0 U13402 ( .IN1(n8539), .IN2(CRC_OUT_7_1), .QN(n13099) );
  NOR2X0 U13403 ( .IN1(DFF_545_n1), .IN2(WX3481), .QN(n13098) );
  NOR3X0 U13404 ( .IN1(n9135), .IN2(n13100), .IN3(n13101), .QN(WX3852) );
  NOR2X0 U13405 ( .IN1(n8556), .IN2(CRC_OUT_7_0), .QN(n13101) );
  NOR2X0 U13406 ( .IN1(DFF_544_n1), .IN2(WX3483), .QN(n13100) );
  NOR3X0 U13407 ( .IN1(n9135), .IN2(n13102), .IN3(n13103), .QN(WX3850) );
  NOR2X0 U13408 ( .IN1(n8131), .IN2(CRC_OUT_7_31), .QN(n13103) );
  NOR2X0 U13409 ( .IN1(DFF_575_n1), .IN2(WX3485), .QN(n13102) );
  NOR2X0 U13410 ( .IN1(n9235), .IN2(n8823), .QN(WX3324) );
  NOR2X0 U13411 ( .IN1(n16056), .IN2(n9159), .QN(WX3322) );
  NOR2X0 U13412 ( .IN1(n16055), .IN2(n9159), .QN(WX3320) );
  NOR2X0 U13413 ( .IN1(n16054), .IN2(n9159), .QN(WX3318) );
  NOR2X0 U13414 ( .IN1(n16053), .IN2(n9159), .QN(WX3316) );
  NOR2X0 U13415 ( .IN1(n16052), .IN2(n9159), .QN(WX3314) );
  NOR2X0 U13416 ( .IN1(n16051), .IN2(n9159), .QN(WX3312) );
  NOR2X0 U13417 ( .IN1(n16050), .IN2(n9159), .QN(WX3310) );
  NOR2X0 U13418 ( .IN1(n16049), .IN2(n9159), .QN(WX3308) );
  NOR2X0 U13419 ( .IN1(n16048), .IN2(n9159), .QN(WX3306) );
  NOR2X0 U13420 ( .IN1(n16047), .IN2(n9159), .QN(WX3304) );
  NOR2X0 U13421 ( .IN1(n16046), .IN2(n9159), .QN(WX3302) );
  NOR2X0 U13422 ( .IN1(n16045), .IN2(n9158), .QN(WX3300) );
  NOR2X0 U13423 ( .IN1(n16044), .IN2(n9158), .QN(WX3298) );
  NOR2X0 U13424 ( .IN1(n16043), .IN2(n9158), .QN(WX3296) );
  NOR2X0 U13425 ( .IN1(n16042), .IN2(n9158), .QN(WX3294) );
  NAND4X0 U13426 ( .IN1(n13104), .IN2(n13105), .IN3(n13106), .IN4(n13107), 
        .QN(WX3292) );
  NAND3X0 U13427 ( .IN1(n12416), .IN2(n12417), .IN3(n9320), .QN(n13107) );
  NAND3X0 U13428 ( .IN1(n13108), .IN2(n13109), .IN3(n13110), .QN(n12417) );
  INVX0 U13429 ( .INP(n13111), .ZN(n13110) );
  NAND2X0 U13430 ( .IN1(n13111), .IN2(n13112), .QN(n12416) );
  NAND2X0 U13431 ( .IN1(n13108), .IN2(n13109), .QN(n13112) );
  NAND2X0 U13432 ( .IN1(n8130), .IN2(WX4650), .QN(n13109) );
  NAND2X0 U13433 ( .IN1(n3691), .IN2(WX4778), .QN(n13108) );
  NOR2X0 U13434 ( .IN1(n13113), .IN2(n13114), .QN(n13111) );
  INVX0 U13435 ( .INP(n13115), .ZN(n13114) );
  NAND2X0 U13436 ( .IN1(test_so36), .IN2(WX4714), .QN(n13115) );
  NOR2X0 U13437 ( .IN1(WX4714), .IN2(test_so36), .QN(n13113) );
  NAND2X0 U13438 ( .IN1(n9108), .IN2(n13116), .QN(n13106) );
  NAND2X0 U13439 ( .IN1(n521), .IN2(n9283), .QN(n13105) );
  NOR2X0 U13440 ( .IN1(n9236), .IN2(n8973), .QN(n521) );
  NAND2X0 U13441 ( .IN1(n9295), .IN2(CRC_OUT_7_0), .QN(n13104) );
  NAND4X0 U13442 ( .IN1(n13117), .IN2(n13118), .IN3(n13119), .IN4(n13120), 
        .QN(WX3290) );
  NAND2X0 U13443 ( .IN1(n9325), .IN2(n12441), .QN(n13120) );
  NAND2X0 U13444 ( .IN1(n13121), .IN2(n13122), .QN(n12441) );
  INVX0 U13445 ( .INP(n13123), .ZN(n13122) );
  NOR2X0 U13446 ( .IN1(n13124), .IN2(n13125), .QN(n13123) );
  NAND2X0 U13447 ( .IN1(n13125), .IN2(n13124), .QN(n13121) );
  NOR2X0 U13448 ( .IN1(n13126), .IN2(n13127), .QN(n13124) );
  NOR2X0 U13449 ( .IN1(WX4776), .IN2(n8006), .QN(n13127) );
  INVX0 U13450 ( .INP(n13128), .ZN(n13126) );
  NAND2X0 U13451 ( .IN1(n8006), .IN2(WX4776), .QN(n13128) );
  NAND2X0 U13452 ( .IN1(n13129), .IN2(n13130), .QN(n13125) );
  NAND2X0 U13453 ( .IN1(n8005), .IN2(WX4648), .QN(n13130) );
  INVX0 U13454 ( .INP(n13131), .ZN(n13129) );
  NOR2X0 U13455 ( .IN1(WX4648), .IN2(n8005), .QN(n13131) );
  NAND2X0 U13456 ( .IN1(n9108), .IN2(n13132), .QN(n13119) );
  NAND2X0 U13457 ( .IN1(n520), .IN2(n9283), .QN(n13118) );
  NOR2X0 U13458 ( .IN1(n9236), .IN2(n8974), .QN(n520) );
  NAND2X0 U13459 ( .IN1(n9295), .IN2(CRC_OUT_7_1), .QN(n13117) );
  NAND4X0 U13460 ( .IN1(n13133), .IN2(n13134), .IN3(n13135), .IN4(n13136), 
        .QN(WX3288) );
  NAND2X0 U13461 ( .IN1(n9325), .IN2(n12457), .QN(n13136) );
  NAND2X0 U13462 ( .IN1(n13137), .IN2(n13138), .QN(n12457) );
  INVX0 U13463 ( .INP(n13139), .ZN(n13138) );
  NOR2X0 U13464 ( .IN1(n13140), .IN2(n13141), .QN(n13139) );
  NAND2X0 U13465 ( .IN1(n13141), .IN2(n13140), .QN(n13137) );
  NOR2X0 U13466 ( .IN1(n13142), .IN2(n13143), .QN(n13140) );
  NOR2X0 U13467 ( .IN1(WX4774), .IN2(n8008), .QN(n13143) );
  INVX0 U13468 ( .INP(n13144), .ZN(n13142) );
  NAND2X0 U13469 ( .IN1(n8008), .IN2(WX4774), .QN(n13144) );
  NAND2X0 U13470 ( .IN1(n13145), .IN2(n13146), .QN(n13141) );
  NAND2X0 U13471 ( .IN1(n8007), .IN2(WX4646), .QN(n13146) );
  INVX0 U13472 ( .INP(n13147), .ZN(n13145) );
  NOR2X0 U13473 ( .IN1(WX4646), .IN2(n8007), .QN(n13147) );
  NAND2X0 U13474 ( .IN1(n9109), .IN2(n13148), .QN(n13135) );
  NAND2X0 U13475 ( .IN1(n519), .IN2(n9283), .QN(n13134) );
  NOR2X0 U13476 ( .IN1(n9070), .IN2(n9158), .QN(n519) );
  NAND2X0 U13477 ( .IN1(n9295), .IN2(CRC_OUT_7_2), .QN(n13133) );
  NAND4X0 U13478 ( .IN1(n13149), .IN2(n13150), .IN3(n13151), .IN4(n13152), 
        .QN(WX3286) );
  NAND2X0 U13479 ( .IN1(n9325), .IN2(n12470), .QN(n13152) );
  NAND2X0 U13480 ( .IN1(n13153), .IN2(n13154), .QN(n12470) );
  INVX0 U13481 ( .INP(n13155), .ZN(n13154) );
  NOR2X0 U13482 ( .IN1(n13156), .IN2(n13157), .QN(n13155) );
  NAND2X0 U13483 ( .IN1(n13157), .IN2(n13156), .QN(n13153) );
  NOR2X0 U13484 ( .IN1(n13158), .IN2(n13159), .QN(n13156) );
  NOR2X0 U13485 ( .IN1(WX4772), .IN2(n8010), .QN(n13159) );
  INVX0 U13486 ( .INP(n13160), .ZN(n13158) );
  NAND2X0 U13487 ( .IN1(n8010), .IN2(WX4772), .QN(n13160) );
  NAND2X0 U13488 ( .IN1(n13161), .IN2(n13162), .QN(n13157) );
  NAND2X0 U13489 ( .IN1(n8009), .IN2(WX4644), .QN(n13162) );
  INVX0 U13490 ( .INP(n13163), .ZN(n13161) );
  NOR2X0 U13491 ( .IN1(WX4644), .IN2(n8009), .QN(n13163) );
  NAND2X0 U13492 ( .IN1(n9108), .IN2(n13164), .QN(n13151) );
  NAND2X0 U13493 ( .IN1(n518), .IN2(n9283), .QN(n13150) );
  NOR2X0 U13494 ( .IN1(n9237), .IN2(n8975), .QN(n518) );
  NAND2X0 U13495 ( .IN1(n9295), .IN2(CRC_OUT_7_3), .QN(n13149) );
  NAND4X0 U13496 ( .IN1(n13165), .IN2(n13166), .IN3(n13167), .IN4(n13168), 
        .QN(WX3284) );
  NAND2X0 U13497 ( .IN1(n9325), .IN2(n12486), .QN(n13168) );
  NAND2X0 U13498 ( .IN1(n13169), .IN2(n13170), .QN(n12486) );
  INVX0 U13499 ( .INP(n13171), .ZN(n13170) );
  NOR2X0 U13500 ( .IN1(n13172), .IN2(n13173), .QN(n13171) );
  NAND2X0 U13501 ( .IN1(n13173), .IN2(n13172), .QN(n13169) );
  NOR2X0 U13502 ( .IN1(n13174), .IN2(n13175), .QN(n13172) );
  NOR2X0 U13503 ( .IN1(WX4770), .IN2(n8012), .QN(n13175) );
  INVX0 U13504 ( .INP(n13176), .ZN(n13174) );
  NAND2X0 U13505 ( .IN1(n8012), .IN2(WX4770), .QN(n13176) );
  NAND2X0 U13506 ( .IN1(n13177), .IN2(n13178), .QN(n13173) );
  NAND2X0 U13507 ( .IN1(n8011), .IN2(WX4642), .QN(n13178) );
  INVX0 U13508 ( .INP(n13179), .ZN(n13177) );
  NOR2X0 U13509 ( .IN1(WX4642), .IN2(n8011), .QN(n13179) );
  NAND2X0 U13510 ( .IN1(n9109), .IN2(n13180), .QN(n13167) );
  NAND2X0 U13511 ( .IN1(n517), .IN2(n9283), .QN(n13166) );
  NOR2X0 U13512 ( .IN1(n9237), .IN2(n8976), .QN(n517) );
  NAND2X0 U13513 ( .IN1(n9295), .IN2(CRC_OUT_7_4), .QN(n13165) );
  NAND4X0 U13514 ( .IN1(n13181), .IN2(n13182), .IN3(n13183), .IN4(n13184), 
        .QN(WX3282) );
  NAND2X0 U13515 ( .IN1(n9325), .IN2(n12499), .QN(n13184) );
  NAND2X0 U13516 ( .IN1(n13185), .IN2(n13186), .QN(n12499) );
  INVX0 U13517 ( .INP(n13187), .ZN(n13186) );
  NOR2X0 U13518 ( .IN1(n13188), .IN2(n13189), .QN(n13187) );
  NAND2X0 U13519 ( .IN1(n13189), .IN2(n13188), .QN(n13185) );
  NOR2X0 U13520 ( .IN1(n13190), .IN2(n13191), .QN(n13188) );
  NOR2X0 U13521 ( .IN1(WX4768), .IN2(n8014), .QN(n13191) );
  INVX0 U13522 ( .INP(n13192), .ZN(n13190) );
  NAND2X0 U13523 ( .IN1(n8014), .IN2(WX4768), .QN(n13192) );
  NAND2X0 U13524 ( .IN1(n13193), .IN2(n13194), .QN(n13189) );
  NAND2X0 U13525 ( .IN1(n8013), .IN2(WX4640), .QN(n13194) );
  INVX0 U13526 ( .INP(n13195), .ZN(n13193) );
  NOR2X0 U13527 ( .IN1(WX4640), .IN2(n8013), .QN(n13195) );
  NAND2X0 U13528 ( .IN1(n9108), .IN2(n13196), .QN(n13183) );
  NAND2X0 U13529 ( .IN1(n516), .IN2(n9283), .QN(n13182) );
  NOR2X0 U13530 ( .IN1(n9237), .IN2(n8977), .QN(n516) );
  NAND2X0 U13531 ( .IN1(n9295), .IN2(CRC_OUT_7_5), .QN(n13181) );
  NAND4X0 U13532 ( .IN1(n13197), .IN2(n13198), .IN3(n13199), .IN4(n13200), 
        .QN(WX3280) );
  NAND3X0 U13533 ( .IN1(n13201), .IN2(n13202), .IN3(n9090), .QN(n13200) );
  NAND2X0 U13534 ( .IN1(n9325), .IN2(n12515), .QN(n13199) );
  NAND2X0 U13535 ( .IN1(n13203), .IN2(n13204), .QN(n12515) );
  INVX0 U13536 ( .INP(n13205), .ZN(n13204) );
  NOR2X0 U13537 ( .IN1(n13206), .IN2(n13207), .QN(n13205) );
  NAND2X0 U13538 ( .IN1(n13207), .IN2(n13206), .QN(n13203) );
  NOR2X0 U13539 ( .IN1(n13208), .IN2(n13209), .QN(n13206) );
  NOR2X0 U13540 ( .IN1(WX4766), .IN2(n8016), .QN(n13209) );
  INVX0 U13541 ( .INP(n13210), .ZN(n13208) );
  NAND2X0 U13542 ( .IN1(n8016), .IN2(WX4766), .QN(n13210) );
  NAND2X0 U13543 ( .IN1(n13211), .IN2(n13212), .QN(n13207) );
  NAND2X0 U13544 ( .IN1(n8015), .IN2(WX4638), .QN(n13212) );
  INVX0 U13545 ( .INP(n13213), .ZN(n13211) );
  NOR2X0 U13546 ( .IN1(WX4638), .IN2(n8015), .QN(n13213) );
  NAND2X0 U13547 ( .IN1(n515), .IN2(n9283), .QN(n13198) );
  NOR2X0 U13548 ( .IN1(n9237), .IN2(n8978), .QN(n515) );
  NAND2X0 U13549 ( .IN1(n9295), .IN2(CRC_OUT_7_6), .QN(n13197) );
  NAND4X0 U13550 ( .IN1(n13214), .IN2(n13215), .IN3(n13216), .IN4(n13217), 
        .QN(WX3278) );
  NAND2X0 U13551 ( .IN1(n9325), .IN2(n12531), .QN(n13217) );
  NAND2X0 U13552 ( .IN1(n13218), .IN2(n13219), .QN(n12531) );
  INVX0 U13553 ( .INP(n13220), .ZN(n13219) );
  NOR2X0 U13554 ( .IN1(n13221), .IN2(n13222), .QN(n13220) );
  NAND2X0 U13555 ( .IN1(n13222), .IN2(n13221), .QN(n13218) );
  NOR2X0 U13556 ( .IN1(n13223), .IN2(n13224), .QN(n13221) );
  NOR2X0 U13557 ( .IN1(WX4764), .IN2(n8018), .QN(n13224) );
  INVX0 U13558 ( .INP(n13225), .ZN(n13223) );
  NAND2X0 U13559 ( .IN1(n8018), .IN2(WX4764), .QN(n13225) );
  NAND2X0 U13560 ( .IN1(n13226), .IN2(n13227), .QN(n13222) );
  NAND2X0 U13561 ( .IN1(n8017), .IN2(WX4636), .QN(n13227) );
  INVX0 U13562 ( .INP(n13228), .ZN(n13226) );
  NOR2X0 U13563 ( .IN1(WX4636), .IN2(n8017), .QN(n13228) );
  NAND2X0 U13564 ( .IN1(n9108), .IN2(n13229), .QN(n13216) );
  NAND2X0 U13565 ( .IN1(n514), .IN2(n9283), .QN(n13215) );
  NOR2X0 U13566 ( .IN1(n9237), .IN2(n8979), .QN(n514) );
  NAND2X0 U13567 ( .IN1(n9295), .IN2(CRC_OUT_7_7), .QN(n13214) );
  NAND4X0 U13568 ( .IN1(n13230), .IN2(n13231), .IN3(n13232), .IN4(n13233), 
        .QN(WX3276) );
  NAND3X0 U13569 ( .IN1(n13234), .IN2(n13235), .IN3(n9089), .QN(n13233) );
  NAND2X0 U13570 ( .IN1(n9325), .IN2(n12547), .QN(n13232) );
  NAND2X0 U13571 ( .IN1(n13236), .IN2(n13237), .QN(n12547) );
  INVX0 U13572 ( .INP(n13238), .ZN(n13237) );
  NOR2X0 U13573 ( .IN1(n13239), .IN2(n13240), .QN(n13238) );
  NAND2X0 U13574 ( .IN1(n13240), .IN2(n13239), .QN(n13236) );
  NOR2X0 U13575 ( .IN1(n13241), .IN2(n13242), .QN(n13239) );
  NOR2X0 U13576 ( .IN1(WX4762), .IN2(n8020), .QN(n13242) );
  INVX0 U13577 ( .INP(n13243), .ZN(n13241) );
  NAND2X0 U13578 ( .IN1(n8020), .IN2(WX4762), .QN(n13243) );
  NAND2X0 U13579 ( .IN1(n13244), .IN2(n13245), .QN(n13240) );
  NAND2X0 U13580 ( .IN1(n8019), .IN2(WX4634), .QN(n13245) );
  INVX0 U13581 ( .INP(n13246), .ZN(n13244) );
  NOR2X0 U13582 ( .IN1(WX4634), .IN2(n8019), .QN(n13246) );
  NAND2X0 U13583 ( .IN1(n513), .IN2(n9283), .QN(n13231) );
  NOR2X0 U13584 ( .IN1(n9237), .IN2(n8980), .QN(n513) );
  NAND2X0 U13585 ( .IN1(n9295), .IN2(CRC_OUT_7_8), .QN(n13230) );
  NAND4X0 U13586 ( .IN1(n13247), .IN2(n13248), .IN3(n13249), .IN4(n13250), 
        .QN(WX3274) );
  NAND2X0 U13587 ( .IN1(n9325), .IN2(n12563), .QN(n13250) );
  NAND2X0 U13588 ( .IN1(n13251), .IN2(n13252), .QN(n12563) );
  INVX0 U13589 ( .INP(n13253), .ZN(n13252) );
  NOR2X0 U13590 ( .IN1(n13254), .IN2(n13255), .QN(n13253) );
  NAND2X0 U13591 ( .IN1(n13255), .IN2(n13254), .QN(n13251) );
  NOR2X0 U13592 ( .IN1(n13256), .IN2(n13257), .QN(n13254) );
  NOR2X0 U13593 ( .IN1(WX4760), .IN2(n8022), .QN(n13257) );
  INVX0 U13594 ( .INP(n13258), .ZN(n13256) );
  NAND2X0 U13595 ( .IN1(n8022), .IN2(WX4760), .QN(n13258) );
  NAND2X0 U13596 ( .IN1(n13259), .IN2(n13260), .QN(n13255) );
  NAND2X0 U13597 ( .IN1(n8021), .IN2(WX4632), .QN(n13260) );
  INVX0 U13598 ( .INP(n13261), .ZN(n13259) );
  NOR2X0 U13599 ( .IN1(WX4632), .IN2(n8021), .QN(n13261) );
  NAND2X0 U13600 ( .IN1(n9109), .IN2(n13262), .QN(n13249) );
  NAND2X0 U13601 ( .IN1(n512), .IN2(n9283), .QN(n13248) );
  NOR2X0 U13602 ( .IN1(n9237), .IN2(n8981), .QN(n512) );
  NAND2X0 U13603 ( .IN1(n9295), .IN2(CRC_OUT_7_9), .QN(n13247) );
  NAND4X0 U13604 ( .IN1(n13263), .IN2(n13264), .IN3(n13265), .IN4(n13266), 
        .QN(WX3272) );
  NAND2X0 U13605 ( .IN1(n9325), .IN2(n12579), .QN(n13266) );
  NAND2X0 U13606 ( .IN1(n13267), .IN2(n13268), .QN(n12579) );
  INVX0 U13607 ( .INP(n13269), .ZN(n13268) );
  NOR2X0 U13608 ( .IN1(n13270), .IN2(n13271), .QN(n13269) );
  NAND2X0 U13609 ( .IN1(n13271), .IN2(n13270), .QN(n13267) );
  NOR2X0 U13610 ( .IN1(n13272), .IN2(n13273), .QN(n13270) );
  NOR2X0 U13611 ( .IN1(WX4758), .IN2(n8024), .QN(n13273) );
  INVX0 U13612 ( .INP(n13274), .ZN(n13272) );
  NAND2X0 U13613 ( .IN1(n8024), .IN2(WX4758), .QN(n13274) );
  NAND2X0 U13614 ( .IN1(n13275), .IN2(n13276), .QN(n13271) );
  NAND2X0 U13615 ( .IN1(n8023), .IN2(WX4630), .QN(n13276) );
  INVX0 U13616 ( .INP(n13277), .ZN(n13275) );
  NOR2X0 U13617 ( .IN1(WX4630), .IN2(n8023), .QN(n13277) );
  NAND2X0 U13618 ( .IN1(n9108), .IN2(n13278), .QN(n13265) );
  NAND2X0 U13619 ( .IN1(n511), .IN2(n9283), .QN(n13264) );
  NOR2X0 U13620 ( .IN1(n9237), .IN2(n8982), .QN(n511) );
  NAND2X0 U13621 ( .IN1(test_so31), .IN2(n9314), .QN(n13263) );
  NAND4X0 U13622 ( .IN1(n13279), .IN2(n13280), .IN3(n13281), .IN4(n13282), 
        .QN(WX3270) );
  NAND3X0 U13623 ( .IN1(n12584), .IN2(n12585), .IN3(n9322), .QN(n13282) );
  NAND3X0 U13624 ( .IN1(n13283), .IN2(n13284), .IN3(n13285), .QN(n12585) );
  INVX0 U13625 ( .INP(n13286), .ZN(n13285) );
  NAND2X0 U13626 ( .IN1(n13286), .IN2(n13287), .QN(n12584) );
  NAND2X0 U13627 ( .IN1(n13283), .IN2(n13284), .QN(n13287) );
  NAND2X0 U13628 ( .IN1(n8026), .IN2(WX4628), .QN(n13284) );
  NAND2X0 U13629 ( .IN1(n3713), .IN2(WX4692), .QN(n13283) );
  NOR2X0 U13630 ( .IN1(n13288), .IN2(n13289), .QN(n13286) );
  NOR2X0 U13631 ( .IN1(n8796), .IN2(n8025), .QN(n13289) );
  INVX0 U13632 ( .INP(n13290), .ZN(n13288) );
  NAND2X0 U13633 ( .IN1(n8025), .IN2(n8796), .QN(n13290) );
  NAND2X0 U13634 ( .IN1(n9109), .IN2(n13291), .QN(n13281) );
  NAND2X0 U13635 ( .IN1(n510), .IN2(n9283), .QN(n13280) );
  NOR2X0 U13636 ( .IN1(n9237), .IN2(n8983), .QN(n510) );
  NAND2X0 U13637 ( .IN1(n9295), .IN2(CRC_OUT_7_11), .QN(n13279) );
  NAND4X0 U13638 ( .IN1(n13292), .IN2(n13293), .IN3(n13294), .IN4(n13295), 
        .QN(WX3268) );
  NAND3X0 U13639 ( .IN1(n13296), .IN2(n13297), .IN3(n9089), .QN(n13295) );
  NAND2X0 U13640 ( .IN1(n9325), .IN2(n12612), .QN(n13294) );
  NAND2X0 U13641 ( .IN1(n13298), .IN2(n13299), .QN(n12612) );
  INVX0 U13642 ( .INP(n13300), .ZN(n13299) );
  NOR2X0 U13643 ( .IN1(n13301), .IN2(n13302), .QN(n13300) );
  NAND2X0 U13644 ( .IN1(n13302), .IN2(n13301), .QN(n13298) );
  NOR2X0 U13645 ( .IN1(n13303), .IN2(n13304), .QN(n13301) );
  NOR2X0 U13646 ( .IN1(WX4754), .IN2(n8028), .QN(n13304) );
  INVX0 U13647 ( .INP(n13305), .ZN(n13303) );
  NAND2X0 U13648 ( .IN1(n8028), .IN2(WX4754), .QN(n13305) );
  NAND2X0 U13649 ( .IN1(n13306), .IN2(n13307), .QN(n13302) );
  NAND2X0 U13650 ( .IN1(n8027), .IN2(WX4626), .QN(n13307) );
  INVX0 U13651 ( .INP(n13308), .ZN(n13306) );
  NOR2X0 U13652 ( .IN1(WX4626), .IN2(n8027), .QN(n13308) );
  NAND2X0 U13653 ( .IN1(n509), .IN2(n9283), .QN(n13293) );
  NOR2X0 U13654 ( .IN1(n9237), .IN2(n8984), .QN(n509) );
  NAND2X0 U13655 ( .IN1(n9296), .IN2(CRC_OUT_7_12), .QN(n13292) );
  NAND4X0 U13656 ( .IN1(n13309), .IN2(n13310), .IN3(n13311), .IN4(n13312), 
        .QN(WX3266) );
  NAND3X0 U13657 ( .IN1(n12617), .IN2(n12618), .IN3(n9322), .QN(n13312) );
  NAND3X0 U13658 ( .IN1(n13313), .IN2(n13314), .IN3(n13315), .QN(n12618) );
  INVX0 U13659 ( .INP(n13316), .ZN(n13315) );
  NAND2X0 U13660 ( .IN1(n13316), .IN2(n13317), .QN(n12617) );
  NAND2X0 U13661 ( .IN1(n13313), .IN2(n13314), .QN(n13317) );
  NAND2X0 U13662 ( .IN1(n8415), .IN2(WX4624), .QN(n13314) );
  NAND2X0 U13663 ( .IN1(n3717), .IN2(WX4752), .QN(n13313) );
  NOR2X0 U13664 ( .IN1(n13318), .IN2(n13319), .QN(n13316) );
  INVX0 U13665 ( .INP(n13320), .ZN(n13319) );
  NAND2X0 U13666 ( .IN1(test_so39), .IN2(WX4560), .QN(n13320) );
  NOR2X0 U13667 ( .IN1(WX4560), .IN2(test_so39), .QN(n13318) );
  NAND2X0 U13668 ( .IN1(n9108), .IN2(n13321), .QN(n13311) );
  NAND2X0 U13669 ( .IN1(n508), .IN2(n9283), .QN(n13310) );
  NOR2X0 U13670 ( .IN1(n9237), .IN2(n8985), .QN(n508) );
  NAND2X0 U13671 ( .IN1(n9296), .IN2(CRC_OUT_7_13), .QN(n13309) );
  NAND4X0 U13672 ( .IN1(n13322), .IN2(n13323), .IN3(n13324), .IN4(n13325), 
        .QN(WX3264) );
  NAND2X0 U13673 ( .IN1(n9325), .IN2(n12645), .QN(n13325) );
  NAND2X0 U13674 ( .IN1(n13326), .IN2(n13327), .QN(n12645) );
  INVX0 U13675 ( .INP(n13328), .ZN(n13327) );
  NOR2X0 U13676 ( .IN1(n13329), .IN2(n13330), .QN(n13328) );
  NAND2X0 U13677 ( .IN1(n13330), .IN2(n13329), .QN(n13326) );
  NOR2X0 U13678 ( .IN1(n13331), .IN2(n13332), .QN(n13329) );
  NOR2X0 U13679 ( .IN1(WX4750), .IN2(n8031), .QN(n13332) );
  INVX0 U13680 ( .INP(n13333), .ZN(n13331) );
  NAND2X0 U13681 ( .IN1(n8031), .IN2(WX4750), .QN(n13333) );
  NAND2X0 U13682 ( .IN1(n13334), .IN2(n13335), .QN(n13330) );
  NAND2X0 U13683 ( .IN1(n8030), .IN2(WX4622), .QN(n13335) );
  INVX0 U13684 ( .INP(n13336), .ZN(n13334) );
  NOR2X0 U13685 ( .IN1(WX4622), .IN2(n8030), .QN(n13336) );
  NAND2X0 U13686 ( .IN1(n9109), .IN2(n13337), .QN(n13324) );
  NAND2X0 U13687 ( .IN1(n507), .IN2(n9283), .QN(n13323) );
  NOR2X0 U13688 ( .IN1(n9237), .IN2(n8986), .QN(n507) );
  NAND2X0 U13689 ( .IN1(n9296), .IN2(CRC_OUT_7_14), .QN(n13322) );
  NAND4X0 U13690 ( .IN1(n13338), .IN2(n13339), .IN3(n13340), .IN4(n13341), 
        .QN(WX3262) );
  NAND3X0 U13691 ( .IN1(n12650), .IN2(n12651), .IN3(n9321), .QN(n13341) );
  NAND3X0 U13692 ( .IN1(n13342), .IN2(n13343), .IN3(n13344), .QN(n12651) );
  INVX0 U13693 ( .INP(n13345), .ZN(n13344) );
  NAND2X0 U13694 ( .IN1(n13345), .IN2(n13346), .QN(n12650) );
  NAND2X0 U13695 ( .IN1(n13342), .IN2(n13343), .QN(n13346) );
  NAND2X0 U13696 ( .IN1(n8413), .IN2(WX4684), .QN(n13343) );
  NAND2X0 U13697 ( .IN1(n8033), .IN2(WX4748), .QN(n13342) );
  NOR2X0 U13698 ( .IN1(n13347), .IN2(n13348), .QN(n13345) );
  INVX0 U13699 ( .INP(n13349), .ZN(n13348) );
  NAND2X0 U13700 ( .IN1(test_so37), .IN2(WX4556), .QN(n13349) );
  NOR2X0 U13701 ( .IN1(WX4556), .IN2(test_so37), .QN(n13347) );
  NAND2X0 U13702 ( .IN1(n9109), .IN2(n13350), .QN(n13340) );
  NAND2X0 U13703 ( .IN1(n506), .IN2(n9283), .QN(n13339) );
  NOR2X0 U13704 ( .IN1(n9237), .IN2(n8987), .QN(n506) );
  NAND2X0 U13705 ( .IN1(n9296), .IN2(CRC_OUT_7_15), .QN(n13338) );
  NAND4X0 U13706 ( .IN1(n13351), .IN2(n13352), .IN3(n13353), .IN4(n13354), 
        .QN(WX3260) );
  NAND2X0 U13707 ( .IN1(n13355), .IN2(n12668), .QN(n13354) );
  NAND2X0 U13708 ( .IN1(n13356), .IN2(n12671), .QN(n12668) );
  NAND2X0 U13709 ( .IN1(n13357), .IN2(n13358), .QN(n13356) );
  NAND2X0 U13710 ( .IN1(n16071), .IN2(n9118), .QN(n13358) );
  NAND2X0 U13711 ( .IN1(TM1), .IN2(n8537), .QN(n13357) );
  NAND3X0 U13712 ( .IN1(n13359), .IN2(n13360), .IN3(n13361), .QN(n13355) );
  NAND2X0 U13713 ( .IN1(n9325), .IN2(n12671), .QN(n13361) );
  NAND2X0 U13714 ( .IN1(n13362), .IN2(n13363), .QN(n12671) );
  NAND2X0 U13715 ( .IN1(n7767), .IN2(n13364), .QN(n13363) );
  INVX0 U13716 ( .INP(n13365), .ZN(n13362) );
  NOR2X0 U13717 ( .IN1(n13364), .IN2(n7767), .QN(n13365) );
  NOR2X0 U13718 ( .IN1(n13366), .IN2(n13367), .QN(n13364) );
  NOR2X0 U13719 ( .IN1(WX4746), .IN2(n7768), .QN(n13367) );
  INVX0 U13720 ( .INP(n13368), .ZN(n13366) );
  NAND2X0 U13721 ( .IN1(n7768), .IN2(WX4746), .QN(n13368) );
  NAND2X0 U13722 ( .IN1(n9790), .IN2(n8537), .QN(n13360) );
  NAND2X0 U13723 ( .IN1(n16071), .IN2(n9078), .QN(n13359) );
  NAND2X0 U13724 ( .IN1(n13369), .IN2(n13370), .QN(n13353) );
  NAND2X0 U13725 ( .IN1(n13371), .IN2(n13372), .QN(n13369) );
  NAND2X0 U13726 ( .IN1(n9109), .IN2(n13373), .QN(n13372) );
  NAND2X0 U13727 ( .IN1(n8119), .IN2(n9110), .QN(n13371) );
  NAND2X0 U13728 ( .IN1(n505), .IN2(n9283), .QN(n13352) );
  NOR2X0 U13729 ( .IN1(n9237), .IN2(n8988), .QN(n505) );
  NAND2X0 U13730 ( .IN1(n9296), .IN2(CRC_OUT_7_16), .QN(n13351) );
  NAND4X0 U13731 ( .IN1(n13374), .IN2(n13375), .IN3(n13376), .IN4(n13377), 
        .QN(WX3258) );
  NAND2X0 U13732 ( .IN1(n13378), .IN2(n12704), .QN(n13377) );
  NAND3X0 U13733 ( .IN1(n13379), .IN2(n13380), .IN3(n12707), .QN(n12704) );
  NAND2X0 U13734 ( .IN1(n8412), .IN2(n9118), .QN(n13380) );
  NAND2X0 U13735 ( .IN1(TM1), .IN2(WX4744), .QN(n13379) );
  NAND3X0 U13736 ( .IN1(n13381), .IN2(n13382), .IN3(n13383), .QN(n13378) );
  NAND2X0 U13737 ( .IN1(n9325), .IN2(n12707), .QN(n13383) );
  NAND2X0 U13738 ( .IN1(n13384), .IN2(n13385), .QN(n12707) );
  NAND2X0 U13739 ( .IN1(n13386), .IN2(WX4680), .QN(n13385) );
  NAND2X0 U13740 ( .IN1(n13387), .IN2(n13388), .QN(n13386) );
  NAND3X0 U13741 ( .IN1(n13387), .IN2(n13388), .IN3(n7770), .QN(n13384) );
  NAND2X0 U13742 ( .IN1(test_so35), .IN2(WX4616), .QN(n13388) );
  NAND2X0 U13743 ( .IN1(n7769), .IN2(n8822), .QN(n13387) );
  NAND2X0 U13744 ( .IN1(n9079), .IN2(WX4744), .QN(n13382) );
  NAND2X0 U13745 ( .IN1(n9083), .IN2(n8412), .QN(n13381) );
  NAND2X0 U13746 ( .IN1(n13389), .IN2(n13390), .QN(n13376) );
  NAND2X0 U13747 ( .IN1(n13391), .IN2(n13392), .QN(n13389) );
  NAND2X0 U13748 ( .IN1(n9109), .IN2(n13393), .QN(n13392) );
  NAND2X0 U13749 ( .IN1(n9109), .IN2(n8597), .QN(n13391) );
  NAND2X0 U13750 ( .IN1(n504), .IN2(n9284), .QN(n13375) );
  NOR2X0 U13751 ( .IN1(n9237), .IN2(n8989), .QN(n504) );
  NAND2X0 U13752 ( .IN1(n9296), .IN2(CRC_OUT_7_17), .QN(n13374) );
  NAND4X0 U13753 ( .IN1(n13394), .IN2(n13395), .IN3(n13396), .IN4(n13397), 
        .QN(WX3256) );
  NAND2X0 U13754 ( .IN1(n13398), .IN2(n12713), .QN(n13397) );
  NAND2X0 U13755 ( .IN1(n13399), .IN2(n12716), .QN(n12713) );
  NAND2X0 U13756 ( .IN1(n13400), .IN2(n13401), .QN(n13399) );
  NAND2X0 U13757 ( .IN1(n16070), .IN2(n9120), .QN(n13401) );
  NAND2X0 U13758 ( .IN1(TM1), .IN2(n8540), .QN(n13400) );
  NAND3X0 U13759 ( .IN1(n13402), .IN2(n13403), .IN3(n13404), .QN(n13398) );
  NAND2X0 U13760 ( .IN1(n9325), .IN2(n12716), .QN(n13404) );
  NAND2X0 U13761 ( .IN1(n13405), .IN2(n13406), .QN(n12716) );
  NAND2X0 U13762 ( .IN1(n7771), .IN2(n13407), .QN(n13406) );
  INVX0 U13763 ( .INP(n13408), .ZN(n13405) );
  NOR2X0 U13764 ( .IN1(n13407), .IN2(n7771), .QN(n13408) );
  NOR2X0 U13765 ( .IN1(n13409), .IN2(n13410), .QN(n13407) );
  NOR2X0 U13766 ( .IN1(WX4742), .IN2(n7772), .QN(n13410) );
  INVX0 U13767 ( .INP(n13411), .ZN(n13409) );
  NAND2X0 U13768 ( .IN1(n7772), .IN2(WX4742), .QN(n13411) );
  NAND2X0 U13769 ( .IN1(n9082), .IN2(n8540), .QN(n13403) );
  NAND2X0 U13770 ( .IN1(n16070), .IN2(n9077), .QN(n13402) );
  NAND2X0 U13771 ( .IN1(n13412), .IN2(n13413), .QN(n13396) );
  NAND2X0 U13772 ( .IN1(n13414), .IN2(n13415), .QN(n13412) );
  NAND2X0 U13773 ( .IN1(n9108), .IN2(n13416), .QN(n13415) );
  NAND2X0 U13774 ( .IN1(n9109), .IN2(n8598), .QN(n13414) );
  NAND2X0 U13775 ( .IN1(n503), .IN2(n9284), .QN(n13395) );
  NOR2X0 U13776 ( .IN1(n9237), .IN2(n8990), .QN(n503) );
  NAND2X0 U13777 ( .IN1(n9296), .IN2(CRC_OUT_7_18), .QN(n13394) );
  NAND4X0 U13778 ( .IN1(n13417), .IN2(n13418), .IN3(n13419), .IN4(n13420), 
        .QN(WX3254) );
  NAND2X0 U13779 ( .IN1(n13421), .IN2(n12751), .QN(n13420) );
  NAND2X0 U13780 ( .IN1(n13422), .IN2(n12754), .QN(n12751) );
  NAND2X0 U13781 ( .IN1(n13423), .IN2(n13424), .QN(n13422) );
  NAND2X0 U13782 ( .IN1(n16069), .IN2(n9120), .QN(n13424) );
  NAND2X0 U13783 ( .IN1(TM1), .IN2(n8541), .QN(n13423) );
  NAND3X0 U13784 ( .IN1(n13425), .IN2(n13426), .IN3(n13427), .QN(n13421) );
  NAND2X0 U13785 ( .IN1(n9326), .IN2(n12754), .QN(n13427) );
  NAND2X0 U13786 ( .IN1(n13428), .IN2(n13429), .QN(n12754) );
  NAND2X0 U13787 ( .IN1(n7773), .IN2(n13430), .QN(n13429) );
  INVX0 U13788 ( .INP(n13431), .ZN(n13428) );
  NOR2X0 U13789 ( .IN1(n13430), .IN2(n7773), .QN(n13431) );
  NOR2X0 U13790 ( .IN1(n13432), .IN2(n13433), .QN(n13430) );
  NOR2X0 U13791 ( .IN1(WX4740), .IN2(n7774), .QN(n13433) );
  INVX0 U13792 ( .INP(n13434), .ZN(n13432) );
  NAND2X0 U13793 ( .IN1(n7774), .IN2(WX4740), .QN(n13434) );
  NAND2X0 U13794 ( .IN1(n9081), .IN2(n8541), .QN(n13426) );
  NAND2X0 U13795 ( .IN1(n16069), .IN2(n9791), .QN(n13425) );
  NAND2X0 U13796 ( .IN1(n13435), .IN2(n13436), .QN(n13419) );
  NAND2X0 U13797 ( .IN1(n13437), .IN2(n13438), .QN(n13435) );
  NAND2X0 U13798 ( .IN1(n9109), .IN2(n13439), .QN(n13438) );
  NAND2X0 U13799 ( .IN1(n9109), .IN2(n8599), .QN(n13437) );
  NAND2X0 U13800 ( .IN1(n502), .IN2(n9284), .QN(n13418) );
  NOR2X0 U13801 ( .IN1(n9238), .IN2(n8991), .QN(n502) );
  NAND2X0 U13802 ( .IN1(n9296), .IN2(CRC_OUT_7_19), .QN(n13417) );
  NAND4X0 U13803 ( .IN1(n13440), .IN2(n13441), .IN3(n13442), .IN4(n13443), 
        .QN(WX3252) );
  NAND2X0 U13804 ( .IN1(n13444), .IN2(n12760), .QN(n13443) );
  NAND2X0 U13805 ( .IN1(n13445), .IN2(n12763), .QN(n12760) );
  NAND2X0 U13806 ( .IN1(n13446), .IN2(n13447), .QN(n13445) );
  NAND2X0 U13807 ( .IN1(n16068), .IN2(n9120), .QN(n13447) );
  NAND2X0 U13808 ( .IN1(TM1), .IN2(n8542), .QN(n13446) );
  NAND3X0 U13809 ( .IN1(n13448), .IN2(n13449), .IN3(n13450), .QN(n13444) );
  NAND2X0 U13810 ( .IN1(n9326), .IN2(n12763), .QN(n13450) );
  NAND2X0 U13811 ( .IN1(n13451), .IN2(n13452), .QN(n12763) );
  NAND2X0 U13812 ( .IN1(n7775), .IN2(n13453), .QN(n13452) );
  INVX0 U13813 ( .INP(n13454), .ZN(n13451) );
  NOR2X0 U13814 ( .IN1(n13453), .IN2(n7775), .QN(n13454) );
  NOR2X0 U13815 ( .IN1(n13455), .IN2(n13456), .QN(n13453) );
  NOR2X0 U13816 ( .IN1(WX4738), .IN2(n7776), .QN(n13456) );
  INVX0 U13817 ( .INP(n13457), .ZN(n13455) );
  NAND2X0 U13818 ( .IN1(n7776), .IN2(WX4738), .QN(n13457) );
  NAND2X0 U13819 ( .IN1(n9790), .IN2(n8542), .QN(n13449) );
  NAND2X0 U13820 ( .IN1(n16068), .IN2(n9079), .QN(n13448) );
  NAND2X0 U13821 ( .IN1(n13458), .IN2(n13459), .QN(n13442) );
  NAND2X0 U13822 ( .IN1(n13460), .IN2(n13461), .QN(n13458) );
  NAND2X0 U13823 ( .IN1(n9108), .IN2(n13462), .QN(n13461) );
  NAND2X0 U13824 ( .IN1(n9105), .IN2(n8600), .QN(n13460) );
  NAND2X0 U13825 ( .IN1(n501), .IN2(n9284), .QN(n13441) );
  NOR2X0 U13826 ( .IN1(n9071), .IN2(n9158), .QN(n501) );
  NAND2X0 U13827 ( .IN1(n9296), .IN2(CRC_OUT_7_20), .QN(n13440) );
  NAND4X0 U13828 ( .IN1(n13463), .IN2(n13464), .IN3(n13465), .IN4(n13466), 
        .QN(WX3250) );
  NAND2X0 U13829 ( .IN1(n13467), .IN2(n12798), .QN(n13466) );
  NAND2X0 U13830 ( .IN1(n13468), .IN2(n12801), .QN(n12798) );
  NAND2X0 U13831 ( .IN1(n13469), .IN2(n13470), .QN(n13468) );
  NAND2X0 U13832 ( .IN1(n16067), .IN2(n9120), .QN(n13470) );
  NAND2X0 U13833 ( .IN1(TM1), .IN2(n8543), .QN(n13469) );
  NAND3X0 U13834 ( .IN1(n13471), .IN2(n13472), .IN3(n13473), .QN(n13467) );
  NAND2X0 U13835 ( .IN1(n9326), .IN2(n12801), .QN(n13473) );
  NAND2X0 U13836 ( .IN1(n13474), .IN2(n13475), .QN(n12801) );
  NAND2X0 U13837 ( .IN1(n7777), .IN2(n13476), .QN(n13475) );
  INVX0 U13838 ( .INP(n13477), .ZN(n13474) );
  NOR2X0 U13839 ( .IN1(n13476), .IN2(n7777), .QN(n13477) );
  NOR2X0 U13840 ( .IN1(n13478), .IN2(n13479), .QN(n13476) );
  NOR2X0 U13841 ( .IN1(WX4736), .IN2(n7778), .QN(n13479) );
  INVX0 U13842 ( .INP(n13480), .ZN(n13478) );
  NAND2X0 U13843 ( .IN1(n7778), .IN2(WX4736), .QN(n13480) );
  NAND2X0 U13844 ( .IN1(n9083), .IN2(n8543), .QN(n13472) );
  NAND2X0 U13845 ( .IN1(n16067), .IN2(n9078), .QN(n13471) );
  NAND2X0 U13846 ( .IN1(n13481), .IN2(n13482), .QN(n13465) );
  NAND2X0 U13847 ( .IN1(n13483), .IN2(n13484), .QN(n13481) );
  NAND2X0 U13848 ( .IN1(n9105), .IN2(n13485), .QN(n13484) );
  NAND2X0 U13849 ( .IN1(n9105), .IN2(n8601), .QN(n13483) );
  NAND2X0 U13850 ( .IN1(n500), .IN2(n9284), .QN(n13464) );
  NOR2X0 U13851 ( .IN1(n9238), .IN2(n8992), .QN(n500) );
  NAND2X0 U13852 ( .IN1(n9296), .IN2(CRC_OUT_7_21), .QN(n13463) );
  NAND4X0 U13853 ( .IN1(n13486), .IN2(n13487), .IN3(n13488), .IN4(n13489), 
        .QN(WX3248) );
  NAND2X0 U13854 ( .IN1(n13490), .IN2(n12818), .QN(n13489) );
  NAND2X0 U13855 ( .IN1(n13491), .IN2(n12821), .QN(n12818) );
  NAND2X0 U13856 ( .IN1(n13492), .IN2(n13493), .QN(n13491) );
  NAND2X0 U13857 ( .IN1(n16066), .IN2(n9120), .QN(n13493) );
  NAND2X0 U13858 ( .IN1(TM1), .IN2(n8544), .QN(n13492) );
  NAND3X0 U13859 ( .IN1(n13494), .IN2(n13495), .IN3(n13496), .QN(n13490) );
  NAND2X0 U13860 ( .IN1(n9326), .IN2(n12821), .QN(n13496) );
  NAND2X0 U13861 ( .IN1(n13497), .IN2(n13498), .QN(n12821) );
  NAND2X0 U13862 ( .IN1(n7779), .IN2(n13499), .QN(n13498) );
  INVX0 U13863 ( .INP(n13500), .ZN(n13497) );
  NOR2X0 U13864 ( .IN1(n13499), .IN2(n7779), .QN(n13500) );
  NOR2X0 U13865 ( .IN1(n13501), .IN2(n13502), .QN(n13499) );
  NOR2X0 U13866 ( .IN1(WX4734), .IN2(n7780), .QN(n13502) );
  INVX0 U13867 ( .INP(n13503), .ZN(n13501) );
  NAND2X0 U13868 ( .IN1(n7780), .IN2(WX4734), .QN(n13503) );
  NAND2X0 U13869 ( .IN1(n9082), .IN2(n8544), .QN(n13495) );
  NAND2X0 U13870 ( .IN1(n16066), .IN2(n9077), .QN(n13494) );
  NAND2X0 U13871 ( .IN1(n13504), .IN2(n13505), .QN(n13488) );
  NAND2X0 U13872 ( .IN1(n13506), .IN2(n13507), .QN(n13504) );
  NAND2X0 U13873 ( .IN1(n9105), .IN2(n13508), .QN(n13507) );
  NAND2X0 U13874 ( .IN1(n9105), .IN2(n8602), .QN(n13506) );
  NAND2X0 U13875 ( .IN1(n499), .IN2(n9284), .QN(n13487) );
  NOR2X0 U13876 ( .IN1(n9238), .IN2(n8993), .QN(n499) );
  NAND2X0 U13877 ( .IN1(n9296), .IN2(CRC_OUT_7_22), .QN(n13486) );
  NAND4X0 U13878 ( .IN1(n13509), .IN2(n13510), .IN3(n13511), .IN4(n13512), 
        .QN(WX3246) );
  NAND2X0 U13879 ( .IN1(n13513), .IN2(n12841), .QN(n13512) );
  NAND2X0 U13880 ( .IN1(n13514), .IN2(n12844), .QN(n12841) );
  NAND2X0 U13881 ( .IN1(n13515), .IN2(n13516), .QN(n13514) );
  NAND2X0 U13882 ( .IN1(n16065), .IN2(n9120), .QN(n13516) );
  NAND2X0 U13883 ( .IN1(TM1), .IN2(n8545), .QN(n13515) );
  NAND3X0 U13884 ( .IN1(n13517), .IN2(n13518), .IN3(n13519), .QN(n13513) );
  NAND2X0 U13885 ( .IN1(n9328), .IN2(n12844), .QN(n13519) );
  NAND2X0 U13886 ( .IN1(n13520), .IN2(n13521), .QN(n12844) );
  NAND2X0 U13887 ( .IN1(n7781), .IN2(n13522), .QN(n13521) );
  INVX0 U13888 ( .INP(n13523), .ZN(n13520) );
  NOR2X0 U13889 ( .IN1(n13522), .IN2(n7781), .QN(n13523) );
  NOR2X0 U13890 ( .IN1(n13524), .IN2(n13525), .QN(n13522) );
  NOR2X0 U13891 ( .IN1(WX4732), .IN2(n7782), .QN(n13525) );
  INVX0 U13892 ( .INP(n13526), .ZN(n13524) );
  NAND2X0 U13893 ( .IN1(n7782), .IN2(WX4732), .QN(n13526) );
  NAND2X0 U13894 ( .IN1(n9081), .IN2(n8545), .QN(n13518) );
  NAND2X0 U13895 ( .IN1(n16065), .IN2(n9791), .QN(n13517) );
  NAND2X0 U13896 ( .IN1(n13527), .IN2(n9111), .QN(n13511) );
  NAND2X0 U13897 ( .IN1(n498), .IN2(n9284), .QN(n13510) );
  NOR2X0 U13898 ( .IN1(n9238), .IN2(n8994), .QN(n498) );
  NAND2X0 U13899 ( .IN1(n9302), .IN2(CRC_OUT_7_23), .QN(n13509) );
  NAND4X0 U13900 ( .IN1(n13528), .IN2(n13529), .IN3(n13530), .IN4(n13531), 
        .QN(WX3244) );
  NAND2X0 U13901 ( .IN1(n13532), .IN2(n12864), .QN(n13531) );
  NAND2X0 U13902 ( .IN1(n13533), .IN2(n12867), .QN(n12864) );
  NAND2X0 U13903 ( .IN1(n13534), .IN2(n13535), .QN(n13533) );
  NAND2X0 U13904 ( .IN1(n16064), .IN2(n9120), .QN(n13535) );
  NAND2X0 U13905 ( .IN1(TM1), .IN2(n8546), .QN(n13534) );
  NAND3X0 U13906 ( .IN1(n13536), .IN2(n13537), .IN3(n13538), .QN(n13532) );
  NAND2X0 U13907 ( .IN1(n9326), .IN2(n12867), .QN(n13538) );
  NAND2X0 U13908 ( .IN1(n13539), .IN2(n13540), .QN(n12867) );
  NAND2X0 U13909 ( .IN1(n7783), .IN2(n13541), .QN(n13540) );
  INVX0 U13910 ( .INP(n13542), .ZN(n13539) );
  NOR2X0 U13911 ( .IN1(n13541), .IN2(n7783), .QN(n13542) );
  NOR2X0 U13912 ( .IN1(n13543), .IN2(n13544), .QN(n13541) );
  NOR2X0 U13913 ( .IN1(WX4730), .IN2(n7784), .QN(n13544) );
  INVX0 U13914 ( .INP(n13545), .ZN(n13543) );
  NAND2X0 U13915 ( .IN1(n7784), .IN2(WX4730), .QN(n13545) );
  NAND2X0 U13916 ( .IN1(n9790), .IN2(n8546), .QN(n13537) );
  NAND2X0 U13917 ( .IN1(n16064), .IN2(n9079), .QN(n13536) );
  NAND2X0 U13918 ( .IN1(n13546), .IN2(n13547), .QN(n13530) );
  NAND2X0 U13919 ( .IN1(n13548), .IN2(n13549), .QN(n13546) );
  NAND2X0 U13920 ( .IN1(n9105), .IN2(n13550), .QN(n13549) );
  NAND2X0 U13921 ( .IN1(n9105), .IN2(n8604), .QN(n13548) );
  NAND2X0 U13922 ( .IN1(n497), .IN2(n9284), .QN(n13529) );
  NOR2X0 U13923 ( .IN1(n9238), .IN2(n8995), .QN(n497) );
  NAND2X0 U13924 ( .IN1(n9297), .IN2(CRC_OUT_7_24), .QN(n13528) );
  NAND4X0 U13925 ( .IN1(n13551), .IN2(n13552), .IN3(n13553), .IN4(n13554), 
        .QN(WX3242) );
  NAND2X0 U13926 ( .IN1(n13555), .IN2(n12887), .QN(n13554) );
  NAND2X0 U13927 ( .IN1(n13556), .IN2(n12890), .QN(n12887) );
  NAND2X0 U13928 ( .IN1(n13557), .IN2(n13558), .QN(n13556) );
  NAND2X0 U13929 ( .IN1(n16063), .IN2(n9120), .QN(n13558) );
  NAND2X0 U13930 ( .IN1(TM1), .IN2(n8547), .QN(n13557) );
  NAND3X0 U13931 ( .IN1(n13559), .IN2(n13560), .IN3(n13561), .QN(n13555) );
  NAND2X0 U13932 ( .IN1(n9326), .IN2(n12890), .QN(n13561) );
  NAND2X0 U13933 ( .IN1(n13562), .IN2(n13563), .QN(n12890) );
  NAND2X0 U13934 ( .IN1(n7785), .IN2(n13564), .QN(n13563) );
  INVX0 U13935 ( .INP(n13565), .ZN(n13562) );
  NOR2X0 U13936 ( .IN1(n13564), .IN2(n7785), .QN(n13565) );
  NOR2X0 U13937 ( .IN1(n13566), .IN2(n13567), .QN(n13564) );
  NOR2X0 U13938 ( .IN1(WX4728), .IN2(n7786), .QN(n13567) );
  INVX0 U13939 ( .INP(n13568), .ZN(n13566) );
  NAND2X0 U13940 ( .IN1(n7786), .IN2(WX4728), .QN(n13568) );
  NAND2X0 U13941 ( .IN1(n9083), .IN2(n8547), .QN(n13560) );
  NAND2X0 U13942 ( .IN1(n16063), .IN2(n9078), .QN(n13559) );
  NAND2X0 U13943 ( .IN1(n13569), .IN2(n13570), .QN(n13553) );
  NAND2X0 U13944 ( .IN1(n13571), .IN2(n13572), .QN(n13569) );
  NAND2X0 U13945 ( .IN1(n9105), .IN2(n13573), .QN(n13572) );
  NAND2X0 U13946 ( .IN1(n9105), .IN2(n8605), .QN(n13571) );
  NAND2X0 U13947 ( .IN1(n496), .IN2(n9284), .QN(n13552) );
  NOR2X0 U13948 ( .IN1(n9238), .IN2(n8996), .QN(n496) );
  NAND2X0 U13949 ( .IN1(n9297), .IN2(CRC_OUT_7_25), .QN(n13551) );
  NAND4X0 U13950 ( .IN1(n13574), .IN2(n13575), .IN3(n13576), .IN4(n13577), 
        .QN(WX3240) );
  NAND2X0 U13951 ( .IN1(n13578), .IN2(n12910), .QN(n13577) );
  NAND2X0 U13952 ( .IN1(n13579), .IN2(n12913), .QN(n12910) );
  NAND2X0 U13953 ( .IN1(n13580), .IN2(n13581), .QN(n13579) );
  NAND2X0 U13954 ( .IN1(n16062), .IN2(n9120), .QN(n13581) );
  NAND2X0 U13955 ( .IN1(TM1), .IN2(n8548), .QN(n13580) );
  NAND3X0 U13956 ( .IN1(n13582), .IN2(n13583), .IN3(n13584), .QN(n13578) );
  NAND2X0 U13957 ( .IN1(n9326), .IN2(n12913), .QN(n13584) );
  NAND2X0 U13958 ( .IN1(n13585), .IN2(n13586), .QN(n12913) );
  NAND2X0 U13959 ( .IN1(n7787), .IN2(n13587), .QN(n13586) );
  INVX0 U13960 ( .INP(n13588), .ZN(n13585) );
  NOR2X0 U13961 ( .IN1(n13587), .IN2(n7787), .QN(n13588) );
  NOR2X0 U13962 ( .IN1(n13589), .IN2(n13590), .QN(n13587) );
  NOR2X0 U13963 ( .IN1(WX4726), .IN2(n7788), .QN(n13590) );
  INVX0 U13964 ( .INP(n13591), .ZN(n13589) );
  NAND2X0 U13965 ( .IN1(n7788), .IN2(WX4726), .QN(n13591) );
  NAND2X0 U13966 ( .IN1(n9082), .IN2(n8548), .QN(n13583) );
  NAND2X0 U13967 ( .IN1(n16062), .IN2(n9077), .QN(n13582) );
  NAND2X0 U13968 ( .IN1(n13592), .IN2(n9111), .QN(n13576) );
  NAND2X0 U13969 ( .IN1(n495), .IN2(n9284), .QN(n13575) );
  NOR2X0 U13970 ( .IN1(n9238), .IN2(n8997), .QN(n495) );
  NAND2X0 U13971 ( .IN1(n9297), .IN2(CRC_OUT_7_26), .QN(n13574) );
  NAND4X0 U13972 ( .IN1(n13593), .IN2(n13594), .IN3(n13595), .IN4(n13596), 
        .QN(WX3238) );
  NAND2X0 U13973 ( .IN1(n13597), .IN2(n12933), .QN(n13596) );
  NAND2X0 U13974 ( .IN1(n13598), .IN2(n12936), .QN(n12933) );
  NAND2X0 U13975 ( .IN1(n13599), .IN2(n13600), .QN(n13598) );
  NAND2X0 U13976 ( .IN1(n16061), .IN2(n9120), .QN(n13600) );
  NAND2X0 U13977 ( .IN1(TM1), .IN2(n8549), .QN(n13599) );
  NAND3X0 U13978 ( .IN1(n13601), .IN2(n13602), .IN3(n13603), .QN(n13597) );
  NAND2X0 U13979 ( .IN1(n9326), .IN2(n12936), .QN(n13603) );
  NAND2X0 U13980 ( .IN1(n13604), .IN2(n13605), .QN(n12936) );
  NAND2X0 U13981 ( .IN1(n7789), .IN2(n13606), .QN(n13605) );
  INVX0 U13982 ( .INP(n13607), .ZN(n13604) );
  NOR2X0 U13983 ( .IN1(n13606), .IN2(n7789), .QN(n13607) );
  NOR2X0 U13984 ( .IN1(n13608), .IN2(n13609), .QN(n13606) );
  NOR2X0 U13985 ( .IN1(WX4724), .IN2(n7790), .QN(n13609) );
  INVX0 U13986 ( .INP(n13610), .ZN(n13608) );
  NAND2X0 U13987 ( .IN1(n7790), .IN2(WX4724), .QN(n13610) );
  NAND2X0 U13988 ( .IN1(n9081), .IN2(n8549), .QN(n13602) );
  NAND2X0 U13989 ( .IN1(n16061), .IN2(n9791), .QN(n13601) );
  NAND2X0 U13990 ( .IN1(n13611), .IN2(n13612), .QN(n13595) );
  NAND2X0 U13991 ( .IN1(n13613), .IN2(n13614), .QN(n13611) );
  NAND2X0 U13992 ( .IN1(n9105), .IN2(n13615), .QN(n13614) );
  NAND2X0 U13993 ( .IN1(n9105), .IN2(n8607), .QN(n13613) );
  NAND2X0 U13994 ( .IN1(n494), .IN2(n9284), .QN(n13594) );
  NOR2X0 U13995 ( .IN1(n9238), .IN2(n8998), .QN(n494) );
  NAND2X0 U13996 ( .IN1(test_so32), .IN2(n9313), .QN(n13593) );
  NAND4X0 U13997 ( .IN1(n13616), .IN2(n13617), .IN3(n13618), .IN4(n13619), 
        .QN(WX3236) );
  NAND2X0 U13998 ( .IN1(n13620), .IN2(n13621), .QN(n13619) );
  NAND2X0 U13999 ( .IN1(n13622), .IN2(n13623), .QN(n13620) );
  NAND2X0 U14000 ( .IN1(n9104), .IN2(n13624), .QN(n13623) );
  NAND2X0 U14001 ( .IN1(n9104), .IN2(n8608), .QN(n13622) );
  NAND2X0 U14002 ( .IN1(n12955), .IN2(n9335), .QN(n13618) );
  NOR2X0 U14003 ( .IN1(n13625), .IN2(n13626), .QN(n12955) );
  INVX0 U14004 ( .INP(n13627), .ZN(n13626) );
  NAND2X0 U14005 ( .IN1(n13628), .IN2(n13629), .QN(n13627) );
  NOR2X0 U14006 ( .IN1(n13629), .IN2(n13628), .QN(n13625) );
  NAND2X0 U14007 ( .IN1(n13630), .IN2(n13631), .QN(n13628) );
  NAND2X0 U14008 ( .IN1(n13632), .IN2(WX4658), .QN(n13631) );
  NAND2X0 U14009 ( .IN1(n13633), .IN2(n13634), .QN(n13632) );
  NAND3X0 U14010 ( .IN1(n13633), .IN2(n13634), .IN3(n7792), .QN(n13630) );
  NAND2X0 U14011 ( .IN1(test_so40), .IN2(WX4594), .QN(n13634) );
  NAND2X0 U14012 ( .IN1(n7791), .IN2(n8800), .QN(n13633) );
  NOR2X0 U14013 ( .IN1(n13635), .IN2(n13636), .QN(n13629) );
  INVX0 U14014 ( .INP(n13637), .ZN(n13636) );
  NAND2X0 U14015 ( .IN1(n16060), .IN2(n9120), .QN(n13637) );
  NOR2X0 U14016 ( .IN1(n9116), .IN2(n16060), .QN(n13635) );
  NAND2X0 U14017 ( .IN1(n493), .IN2(n9284), .QN(n13617) );
  NOR2X0 U14018 ( .IN1(n9238), .IN2(n8999), .QN(n493) );
  NAND2X0 U14019 ( .IN1(n9297), .IN2(CRC_OUT_7_28), .QN(n13616) );
  NAND4X0 U14020 ( .IN1(n13638), .IN2(n13639), .IN3(n13640), .IN4(n13641), 
        .QN(WX3234) );
  NAND2X0 U14021 ( .IN1(n13642), .IN2(n12975), .QN(n13641) );
  NAND2X0 U14022 ( .IN1(n13643), .IN2(n12978), .QN(n12975) );
  NAND2X0 U14023 ( .IN1(n13644), .IN2(n13645), .QN(n13643) );
  NAND2X0 U14024 ( .IN1(n16059), .IN2(n9120), .QN(n13645) );
  NAND2X0 U14025 ( .IN1(TM1), .IN2(n8551), .QN(n13644) );
  NAND3X0 U14026 ( .IN1(n13646), .IN2(n13647), .IN3(n13648), .QN(n13642) );
  NAND2X0 U14027 ( .IN1(n9326), .IN2(n12978), .QN(n13648) );
  NAND2X0 U14028 ( .IN1(n13649), .IN2(n13650), .QN(n12978) );
  NAND2X0 U14029 ( .IN1(n7793), .IN2(n13651), .QN(n13650) );
  INVX0 U14030 ( .INP(n13652), .ZN(n13649) );
  NOR2X0 U14031 ( .IN1(n13651), .IN2(n7793), .QN(n13652) );
  NOR2X0 U14032 ( .IN1(n13653), .IN2(n13654), .QN(n13651) );
  NOR2X0 U14033 ( .IN1(WX4720), .IN2(n7794), .QN(n13654) );
  INVX0 U14034 ( .INP(n13655), .ZN(n13653) );
  NAND2X0 U14035 ( .IN1(n7794), .IN2(WX4720), .QN(n13655) );
  NAND2X0 U14036 ( .IN1(n9790), .IN2(n8551), .QN(n13647) );
  NAND2X0 U14037 ( .IN1(n16059), .IN2(n9079), .QN(n13646) );
  NAND2X0 U14038 ( .IN1(n13656), .IN2(n13657), .QN(n13640) );
  NAND2X0 U14039 ( .IN1(n13658), .IN2(n13659), .QN(n13656) );
  NAND2X0 U14040 ( .IN1(n9104), .IN2(n13660), .QN(n13659) );
  NAND2X0 U14041 ( .IN1(n9104), .IN2(n8609), .QN(n13658) );
  NAND2X0 U14042 ( .IN1(n492), .IN2(n9284), .QN(n13639) );
  NOR2X0 U14043 ( .IN1(n9238), .IN2(n9000), .QN(n492) );
  NAND2X0 U14044 ( .IN1(n9297), .IN2(CRC_OUT_7_29), .QN(n13638) );
  NAND4X0 U14045 ( .IN1(n13661), .IN2(n13662), .IN3(n13663), .IN4(n13664), 
        .QN(WX3232) );
  NAND2X0 U14046 ( .IN1(n12997), .IN2(n9335), .QN(n13664) );
  NOR2X0 U14047 ( .IN1(n13665), .IN2(n13666), .QN(n12997) );
  INVX0 U14048 ( .INP(n13667), .ZN(n13666) );
  NAND2X0 U14049 ( .IN1(n13668), .IN2(n13669), .QN(n13667) );
  NOR2X0 U14050 ( .IN1(n13669), .IN2(n13668), .QN(n13665) );
  NAND2X0 U14051 ( .IN1(n13670), .IN2(n13671), .QN(n13668) );
  NAND2X0 U14052 ( .IN1(n8355), .IN2(n13672), .QN(n13671) );
  INVX0 U14053 ( .INP(n13673), .ZN(n13672) );
  NAND2X0 U14054 ( .IN1(n13673), .IN2(WX4718), .QN(n13670) );
  NAND2X0 U14055 ( .IN1(n13674), .IN2(n13675), .QN(n13673) );
  INVX0 U14056 ( .INP(n13676), .ZN(n13675) );
  NOR2X0 U14057 ( .IN1(n8813), .IN2(n16058), .QN(n13676) );
  NAND2X0 U14058 ( .IN1(n16058), .IN2(n8813), .QN(n13674) );
  NOR2X0 U14059 ( .IN1(n13677), .IN2(n13678), .QN(n13669) );
  INVX0 U14060 ( .INP(n13679), .ZN(n13678) );
  NAND2X0 U14061 ( .IN1(n7795), .IN2(n9120), .QN(n13679) );
  NOR2X0 U14062 ( .IN1(n9116), .IN2(n7795), .QN(n13677) );
  NAND2X0 U14063 ( .IN1(n13680), .IN2(n9110), .QN(n13663) );
  NAND2X0 U14064 ( .IN1(n491), .IN2(n9284), .QN(n13662) );
  NOR2X0 U14065 ( .IN1(n9238), .IN2(n9001), .QN(n491) );
  NAND2X0 U14066 ( .IN1(n9297), .IN2(CRC_OUT_7_30), .QN(n13661) );
  NAND4X0 U14067 ( .IN1(n13681), .IN2(n13682), .IN3(n13683), .IN4(n13684), 
        .QN(WX3230) );
  NAND2X0 U14068 ( .IN1(n13685), .IN2(n13017), .QN(n13684) );
  NAND2X0 U14069 ( .IN1(n13686), .IN2(n13020), .QN(n13017) );
  NAND2X0 U14070 ( .IN1(n13687), .IN2(n13688), .QN(n13686) );
  NAND2X0 U14071 ( .IN1(n16057), .IN2(n9120), .QN(n13688) );
  NAND2X0 U14072 ( .IN1(TM1), .IN2(n8553), .QN(n13687) );
  NAND3X0 U14073 ( .IN1(n13689), .IN2(n13690), .IN3(n13691), .QN(n13685) );
  NAND2X0 U14074 ( .IN1(n9326), .IN2(n13020), .QN(n13691) );
  NAND2X0 U14075 ( .IN1(n13692), .IN2(n13693), .QN(n13020) );
  NAND2X0 U14076 ( .IN1(n7621), .IN2(n13694), .QN(n13693) );
  INVX0 U14077 ( .INP(n13695), .ZN(n13692) );
  NOR2X0 U14078 ( .IN1(n13694), .IN2(n7621), .QN(n13695) );
  NOR2X0 U14079 ( .IN1(n13696), .IN2(n13697), .QN(n13694) );
  NOR2X0 U14080 ( .IN1(WX4716), .IN2(n7622), .QN(n13697) );
  INVX0 U14081 ( .INP(n13698), .ZN(n13696) );
  NAND2X0 U14082 ( .IN1(n7622), .IN2(WX4716), .QN(n13698) );
  NAND2X0 U14083 ( .IN1(n9083), .IN2(n8553), .QN(n13690) );
  NAND2X0 U14084 ( .IN1(n16057), .IN2(n9078), .QN(n13689) );
  NAND2X0 U14085 ( .IN1(n13699), .IN2(n13700), .QN(n13683) );
  NAND2X0 U14086 ( .IN1(n13701), .IN2(n13702), .QN(n13699) );
  NAND2X0 U14087 ( .IN1(n9104), .IN2(n13703), .QN(n13702) );
  NAND2X0 U14088 ( .IN1(n9104), .IN2(n8611), .QN(n13701) );
  NAND2X0 U14089 ( .IN1(n9297), .IN2(CRC_OUT_7_31), .QN(n13682) );
  NAND2X0 U14090 ( .IN1(n2245), .IN2(WX3071), .QN(n13681) );
  NOR2X0 U14091 ( .IN1(n9238), .IN2(WX3071), .QN(WX3132) );
  NOR3X0 U14092 ( .IN1(n9135), .IN2(n13704), .IN3(n13705), .QN(WX2619) );
  NOR2X0 U14093 ( .IN1(n8557), .IN2(CRC_OUT_8_30), .QN(n13705) );
  NOR2X0 U14094 ( .IN1(DFF_382_n1), .IN2(WX2130), .QN(n13704) );
  NOR3X0 U14095 ( .IN1(n9135), .IN2(n13706), .IN3(n13707), .QN(WX2617) );
  NOR2X0 U14096 ( .IN1(n8574), .IN2(CRC_OUT_8_29), .QN(n13707) );
  NOR2X0 U14097 ( .IN1(DFF_381_n1), .IN2(WX2132), .QN(n13706) );
  NOR3X0 U14098 ( .IN1(n9140), .IN2(n13708), .IN3(n13709), .QN(WX2615) );
  NOR2X0 U14099 ( .IN1(n8575), .IN2(CRC_OUT_8_28), .QN(n13709) );
  NOR2X0 U14100 ( .IN1(DFF_380_n1), .IN2(WX2134), .QN(n13708) );
  NOR2X0 U14101 ( .IN1(n9239), .IN2(n13710), .QN(WX2613) );
  NOR2X0 U14102 ( .IN1(n13711), .IN2(n13712), .QN(n13710) );
  NOR2X0 U14103 ( .IN1(test_so18), .IN2(CRC_OUT_8_27), .QN(n13712) );
  NOR2X0 U14104 ( .IN1(DFF_379_n1), .IN2(n8802), .QN(n13711) );
  NOR3X0 U14105 ( .IN1(n9154), .IN2(n13713), .IN3(n13714), .QN(WX2611) );
  NOR2X0 U14106 ( .IN1(n8587), .IN2(CRC_OUT_8_26), .QN(n13714) );
  NOR2X0 U14107 ( .IN1(DFF_378_n1), .IN2(WX2138), .QN(n13713) );
  NOR2X0 U14108 ( .IN1(n9239), .IN2(n13715), .QN(WX2609) );
  NOR2X0 U14109 ( .IN1(n13716), .IN2(n13717), .QN(n13715) );
  NOR2X0 U14110 ( .IN1(test_so21), .IN2(WX2140), .QN(n13717) );
  INVX0 U14111 ( .INP(n13718), .ZN(n13716) );
  NAND2X0 U14112 ( .IN1(WX2140), .IN2(test_so21), .QN(n13718) );
  NOR3X0 U14113 ( .IN1(n9155), .IN2(n13719), .IN3(n13720), .QN(WX2607) );
  NOR2X0 U14114 ( .IN1(n8589), .IN2(CRC_OUT_8_24), .QN(n13720) );
  NOR2X0 U14115 ( .IN1(DFF_376_n1), .IN2(WX2142), .QN(n13719) );
  NOR3X0 U14116 ( .IN1(n9154), .IN2(n13721), .IN3(n13722), .QN(WX2605) );
  NOR2X0 U14117 ( .IN1(n8590), .IN2(CRC_OUT_8_23), .QN(n13722) );
  NOR2X0 U14118 ( .IN1(DFF_375_n1), .IN2(WX2144), .QN(n13721) );
  NOR3X0 U14119 ( .IN1(n9154), .IN2(n13723), .IN3(n13724), .QN(WX2603) );
  NOR2X0 U14120 ( .IN1(n8591), .IN2(CRC_OUT_8_22), .QN(n13724) );
  NOR2X0 U14121 ( .IN1(DFF_374_n1), .IN2(WX2146), .QN(n13723) );
  NOR3X0 U14122 ( .IN1(n9154), .IN2(n13725), .IN3(n13726), .QN(WX2601) );
  NOR2X0 U14123 ( .IN1(n8592), .IN2(CRC_OUT_8_21), .QN(n13726) );
  NOR2X0 U14124 ( .IN1(DFF_373_n1), .IN2(WX2148), .QN(n13725) );
  NOR3X0 U14125 ( .IN1(n9153), .IN2(n13727), .IN3(n13728), .QN(WX2599) );
  NOR2X0 U14126 ( .IN1(n8593), .IN2(CRC_OUT_8_20), .QN(n13728) );
  NOR2X0 U14127 ( .IN1(DFF_372_n1), .IN2(WX2150), .QN(n13727) );
  NOR3X0 U14128 ( .IN1(n9154), .IN2(n13729), .IN3(n13730), .QN(WX2597) );
  NOR2X0 U14129 ( .IN1(n8594), .IN2(CRC_OUT_8_19), .QN(n13730) );
  NOR2X0 U14130 ( .IN1(DFF_371_n1), .IN2(WX2152), .QN(n13729) );
  NOR3X0 U14131 ( .IN1(n9154), .IN2(n13731), .IN3(n13732), .QN(WX2595) );
  NOR2X0 U14132 ( .IN1(n8595), .IN2(CRC_OUT_8_18), .QN(n13732) );
  NOR2X0 U14133 ( .IN1(DFF_370_n1), .IN2(WX2154), .QN(n13731) );
  NOR3X0 U14134 ( .IN1(n9154), .IN2(n13733), .IN3(n13734), .QN(WX2593) );
  NOR2X0 U14135 ( .IN1(n8596), .IN2(CRC_OUT_8_17), .QN(n13734) );
  NOR2X0 U14136 ( .IN1(DFF_369_n1), .IN2(WX2156), .QN(n13733) );
  NOR3X0 U14137 ( .IN1(n9154), .IN2(n13735), .IN3(n13736), .QN(WX2591) );
  NOR2X0 U14138 ( .IN1(n8614), .IN2(CRC_OUT_8_16), .QN(n13736) );
  NOR2X0 U14139 ( .IN1(DFF_368_n1), .IN2(WX2158), .QN(n13735) );
  NOR2X0 U14140 ( .IN1(n9239), .IN2(n13737), .QN(WX2589) );
  NOR2X0 U14141 ( .IN1(n13738), .IN2(n13739), .QN(n13737) );
  INVX0 U14142 ( .INP(n13740), .ZN(n13739) );
  NAND2X0 U14143 ( .IN1(CRC_OUT_8_15), .IN2(n13741), .QN(n13740) );
  NOR2X0 U14144 ( .IN1(n13741), .IN2(CRC_OUT_8_15), .QN(n13738) );
  NAND2X0 U14145 ( .IN1(n13742), .IN2(n13743), .QN(n13741) );
  NAND2X0 U14146 ( .IN1(n8122), .IN2(CRC_OUT_8_31), .QN(n13743) );
  NAND2X0 U14147 ( .IN1(DFF_383_n1), .IN2(WX2160), .QN(n13742) );
  NOR3X0 U14148 ( .IN1(n9153), .IN2(n13744), .IN3(n13745), .QN(WX2587) );
  NOR2X0 U14149 ( .IN1(n8615), .IN2(CRC_OUT_8_14), .QN(n13745) );
  NOR2X0 U14150 ( .IN1(DFF_366_n1), .IN2(WX2162), .QN(n13744) );
  NOR3X0 U14151 ( .IN1(n9153), .IN2(n13746), .IN3(n13747), .QN(WX2585) );
  NOR2X0 U14152 ( .IN1(n8633), .IN2(CRC_OUT_8_13), .QN(n13747) );
  NOR2X0 U14153 ( .IN1(DFF_365_n1), .IN2(WX2164), .QN(n13746) );
  NOR3X0 U14154 ( .IN1(n9152), .IN2(n13748), .IN3(n13749), .QN(WX2583) );
  NOR2X0 U14155 ( .IN1(n8634), .IN2(CRC_OUT_8_12), .QN(n13749) );
  NOR2X0 U14156 ( .IN1(DFF_364_n1), .IN2(WX2166), .QN(n13748) );
  NOR3X0 U14157 ( .IN1(n9154), .IN2(n13750), .IN3(n13751), .QN(WX2581) );
  NOR2X0 U14158 ( .IN1(n8645), .IN2(CRC_OUT_8_11), .QN(n13751) );
  NOR2X0 U14159 ( .IN1(DFF_363_n1), .IN2(WX2168), .QN(n13750) );
  NOR2X0 U14160 ( .IN1(n9240), .IN2(n13752), .QN(WX2579) );
  NOR2X0 U14161 ( .IN1(n13753), .IN2(n13754), .QN(n13752) );
  INVX0 U14162 ( .INP(n13755), .ZN(n13754) );
  NAND2X0 U14163 ( .IN1(CRC_OUT_8_10), .IN2(n13756), .QN(n13755) );
  NOR2X0 U14164 ( .IN1(n13756), .IN2(CRC_OUT_8_10), .QN(n13753) );
  NAND2X0 U14165 ( .IN1(n13757), .IN2(n13758), .QN(n13756) );
  NAND2X0 U14166 ( .IN1(n8123), .IN2(CRC_OUT_8_31), .QN(n13758) );
  NAND2X0 U14167 ( .IN1(DFF_383_n1), .IN2(WX2170), .QN(n13757) );
  NOR2X0 U14168 ( .IN1(n9240), .IN2(n13759), .QN(WX2577) );
  NOR2X0 U14169 ( .IN1(n13760), .IN2(n13761), .QN(n13759) );
  NOR2X0 U14170 ( .IN1(test_so19), .IN2(CRC_OUT_8_9), .QN(n13761) );
  NOR2X0 U14171 ( .IN1(DFF_361_n1), .IN2(n8792), .QN(n13760) );
  NOR3X0 U14172 ( .IN1(n9153), .IN2(n13762), .IN3(n13763), .QN(WX2575) );
  NOR2X0 U14173 ( .IN1(n8646), .IN2(CRC_OUT_8_8), .QN(n13763) );
  NOR2X0 U14174 ( .IN1(DFF_360_n1), .IN2(WX2174), .QN(n13762) );
  NOR2X0 U14175 ( .IN1(n9240), .IN2(n13764), .QN(WX2573) );
  NOR2X0 U14176 ( .IN1(n13765), .IN2(n13766), .QN(n13764) );
  NOR2X0 U14177 ( .IN1(test_so20), .IN2(WX2176), .QN(n13766) );
  INVX0 U14178 ( .INP(n13767), .ZN(n13765) );
  NAND2X0 U14179 ( .IN1(WX2176), .IN2(test_so20), .QN(n13767) );
  NOR3X0 U14180 ( .IN1(n9152), .IN2(n13768), .IN3(n13769), .QN(WX2571) );
  NOR2X0 U14181 ( .IN1(n8648), .IN2(CRC_OUT_8_6), .QN(n13769) );
  NOR2X0 U14182 ( .IN1(DFF_358_n1), .IN2(WX2178), .QN(n13768) );
  NOR3X0 U14183 ( .IN1(n9154), .IN2(n13770), .IN3(n13771), .QN(WX2569) );
  NOR2X0 U14184 ( .IN1(n8649), .IN2(CRC_OUT_8_5), .QN(n13771) );
  NOR2X0 U14185 ( .IN1(DFF_357_n1), .IN2(WX2180), .QN(n13770) );
  NOR3X0 U14186 ( .IN1(n9153), .IN2(n13772), .IN3(n13773), .QN(WX2567) );
  NOR2X0 U14187 ( .IN1(n8650), .IN2(CRC_OUT_8_4), .QN(n13773) );
  NOR2X0 U14188 ( .IN1(DFF_356_n1), .IN2(WX2182), .QN(n13772) );
  NOR2X0 U14189 ( .IN1(n9240), .IN2(n13774), .QN(WX2565) );
  NOR2X0 U14190 ( .IN1(n13775), .IN2(n13776), .QN(n13774) );
  INVX0 U14191 ( .INP(n13777), .ZN(n13776) );
  NAND2X0 U14192 ( .IN1(CRC_OUT_8_3), .IN2(n13778), .QN(n13777) );
  NOR2X0 U14193 ( .IN1(n13778), .IN2(CRC_OUT_8_3), .QN(n13775) );
  NAND2X0 U14194 ( .IN1(n13779), .IN2(n13780), .QN(n13778) );
  NAND2X0 U14195 ( .IN1(n8124), .IN2(CRC_OUT_8_31), .QN(n13780) );
  NAND2X0 U14196 ( .IN1(DFF_383_n1), .IN2(WX2184), .QN(n13779) );
  NOR3X0 U14197 ( .IN1(n9154), .IN2(n13781), .IN3(n13782), .QN(WX2563) );
  NOR2X0 U14198 ( .IN1(n8651), .IN2(CRC_OUT_8_2), .QN(n13782) );
  NOR2X0 U14199 ( .IN1(DFF_354_n1), .IN2(WX2186), .QN(n13781) );
  NOR3X0 U14200 ( .IN1(n9154), .IN2(n13783), .IN3(n13784), .QN(WX2561) );
  NOR2X0 U14201 ( .IN1(n8652), .IN2(CRC_OUT_8_1), .QN(n13784) );
  NOR2X0 U14202 ( .IN1(DFF_353_n1), .IN2(WX2188), .QN(n13783) );
  NOR3X0 U14203 ( .IN1(n9153), .IN2(n13785), .IN3(n13786), .QN(WX2559) );
  NOR2X0 U14204 ( .IN1(n8659), .IN2(CRC_OUT_8_0), .QN(n13786) );
  NOR2X0 U14205 ( .IN1(DFF_352_n1), .IN2(WX2190), .QN(n13785) );
  NOR3X0 U14206 ( .IN1(n9153), .IN2(n13787), .IN3(n13788), .QN(WX2557) );
  NOR2X0 U14207 ( .IN1(n8132), .IN2(CRC_OUT_8_31), .QN(n13788) );
  NOR2X0 U14208 ( .IN1(DFF_383_n1), .IN2(WX2192), .QN(n13787) );
  NOR2X0 U14209 ( .IN1(n16041), .IN2(n9159), .QN(WX2031) );
  NOR2X0 U14210 ( .IN1(n16040), .IN2(n9159), .QN(WX2029) );
  NOR2X0 U14211 ( .IN1(n16039), .IN2(n9159), .QN(WX2027) );
  NOR2X0 U14212 ( .IN1(n16038), .IN2(n9159), .QN(WX2025) );
  NOR2X0 U14213 ( .IN1(n16037), .IN2(n9160), .QN(WX2023) );
  NOR2X0 U14214 ( .IN1(n16036), .IN2(n9160), .QN(WX2021) );
  NOR2X0 U14215 ( .IN1(n9240), .IN2(n8824), .QN(WX2019) );
  NOR2X0 U14216 ( .IN1(n16035), .IN2(n9160), .QN(WX2017) );
  NOR2X0 U14217 ( .IN1(n16034), .IN2(n9160), .QN(WX2015) );
  NOR2X0 U14218 ( .IN1(n16033), .IN2(n9161), .QN(WX2013) );
  NOR2X0 U14219 ( .IN1(n16032), .IN2(n9161), .QN(WX2011) );
  NOR2X0 U14220 ( .IN1(n16031), .IN2(n9161), .QN(WX2009) );
  NOR2X0 U14221 ( .IN1(n16030), .IN2(n9161), .QN(WX2007) );
  NOR2X0 U14222 ( .IN1(n16029), .IN2(n9161), .QN(WX2005) );
  NOR2X0 U14223 ( .IN1(n16028), .IN2(n9161), .QN(WX2003) );
  NOR2X0 U14224 ( .IN1(n16027), .IN2(n9161), .QN(WX2001) );
  NAND4X0 U14225 ( .IN1(n13789), .IN2(n13790), .IN3(n13791), .IN4(n13792), 
        .QN(WX1999) );
  NAND3X0 U14226 ( .IN1(n11378), .IN2(n11379), .IN3(n9089), .QN(n13792) );
  NAND3X0 U14227 ( .IN1(n13793), .IN2(n13794), .IN3(n13795), .QN(n11379) );
  INVX0 U14228 ( .INP(n13796), .ZN(n13795) );
  NAND2X0 U14229 ( .IN1(n13796), .IN2(n13797), .QN(n11378) );
  NAND2X0 U14230 ( .IN1(n13793), .IN2(n13794), .QN(n13797) );
  NAND2X0 U14231 ( .IN1(n8132), .IN2(WX2128), .QN(n13794) );
  NAND2X0 U14232 ( .IN1(n8066), .IN2(WX2192), .QN(n13793) );
  NOR2X0 U14233 ( .IN1(n13798), .IN2(n13799), .QN(n13796) );
  INVX0 U14234 ( .INP(n13800), .ZN(n13799) );
  NAND2X0 U14235 ( .IN1(test_so16), .IN2(WX2000), .QN(n13800) );
  NOR2X0 U14236 ( .IN1(WX2000), .IN2(test_so16), .QN(n13798) );
  NAND2X0 U14237 ( .IN1(n9326), .IN2(n13116), .QN(n13791) );
  NAND2X0 U14238 ( .IN1(n13801), .IN2(n13802), .QN(n13116) );
  INVX0 U14239 ( .INP(n13803), .ZN(n13802) );
  NOR2X0 U14240 ( .IN1(n13804), .IN2(n13805), .QN(n13803) );
  NAND2X0 U14241 ( .IN1(n13805), .IN2(n13804), .QN(n13801) );
  NOR2X0 U14242 ( .IN1(n13806), .IN2(n13807), .QN(n13804) );
  NOR2X0 U14243 ( .IN1(WX3485), .IN2(n8035), .QN(n13807) );
  INVX0 U14244 ( .INP(n13808), .ZN(n13806) );
  NAND2X0 U14245 ( .IN1(n8035), .IN2(WX3485), .QN(n13808) );
  NAND2X0 U14246 ( .IN1(n13809), .IN2(n13810), .QN(n13805) );
  NAND2X0 U14247 ( .IN1(n8034), .IN2(WX3357), .QN(n13810) );
  INVX0 U14248 ( .INP(n13811), .ZN(n13809) );
  NOR2X0 U14249 ( .IN1(WX3357), .IN2(n8034), .QN(n13811) );
  NAND2X0 U14250 ( .IN1(n280), .IN2(n9284), .QN(n13790) );
  NOR2X0 U14251 ( .IN1(n9240), .IN2(n9002), .QN(n280) );
  NAND2X0 U14252 ( .IN1(n9297), .IN2(CRC_OUT_8_0), .QN(n13789) );
  NAND4X0 U14253 ( .IN1(n13812), .IN2(n13813), .IN3(n13814), .IN4(n13815), 
        .QN(WX1997) );
  NAND2X0 U14254 ( .IN1(n9326), .IN2(n13132), .QN(n13815) );
  NAND2X0 U14255 ( .IN1(n13816), .IN2(n13817), .QN(n13132) );
  INVX0 U14256 ( .INP(n13818), .ZN(n13817) );
  NOR2X0 U14257 ( .IN1(n13819), .IN2(n13820), .QN(n13818) );
  NAND2X0 U14258 ( .IN1(n13820), .IN2(n13819), .QN(n13816) );
  NOR2X0 U14259 ( .IN1(n13821), .IN2(n13822), .QN(n13819) );
  NOR2X0 U14260 ( .IN1(WX3483), .IN2(n8037), .QN(n13822) );
  INVX0 U14261 ( .INP(n13823), .ZN(n13821) );
  NAND2X0 U14262 ( .IN1(n8037), .IN2(WX3483), .QN(n13823) );
  NAND2X0 U14263 ( .IN1(n13824), .IN2(n13825), .QN(n13820) );
  NAND2X0 U14264 ( .IN1(n8036), .IN2(WX3355), .QN(n13825) );
  INVX0 U14265 ( .INP(n13826), .ZN(n13824) );
  NOR2X0 U14266 ( .IN1(WX3355), .IN2(n8036), .QN(n13826) );
  NAND2X0 U14267 ( .IN1(n9104), .IN2(n11385), .QN(n13814) );
  NAND2X0 U14268 ( .IN1(n13827), .IN2(n13828), .QN(n11385) );
  INVX0 U14269 ( .INP(n13829), .ZN(n13828) );
  NOR2X0 U14270 ( .IN1(n13830), .IN2(n13831), .QN(n13829) );
  NAND2X0 U14271 ( .IN1(n13831), .IN2(n13830), .QN(n13827) );
  NOR2X0 U14272 ( .IN1(n13832), .IN2(n13833), .QN(n13830) );
  NOR2X0 U14273 ( .IN1(WX2190), .IN2(n8068), .QN(n13833) );
  INVX0 U14274 ( .INP(n13834), .ZN(n13832) );
  NAND2X0 U14275 ( .IN1(n8068), .IN2(WX2190), .QN(n13834) );
  NAND2X0 U14276 ( .IN1(n13835), .IN2(n13836), .QN(n13831) );
  NAND2X0 U14277 ( .IN1(n8067), .IN2(WX2062), .QN(n13836) );
  INVX0 U14278 ( .INP(n13837), .ZN(n13835) );
  NOR2X0 U14279 ( .IN1(WX2062), .IN2(n8067), .QN(n13837) );
  NAND2X0 U14280 ( .IN1(n279), .IN2(n9284), .QN(n13813) );
  NOR2X0 U14281 ( .IN1(n9241), .IN2(n9003), .QN(n279) );
  NAND2X0 U14282 ( .IN1(n9297), .IN2(CRC_OUT_8_1), .QN(n13812) );
  NAND4X0 U14283 ( .IN1(n13838), .IN2(n13839), .IN3(n13840), .IN4(n13841), 
        .QN(WX1995) );
  NAND2X0 U14284 ( .IN1(n9326), .IN2(n13148), .QN(n13841) );
  NAND2X0 U14285 ( .IN1(n13842), .IN2(n13843), .QN(n13148) );
  INVX0 U14286 ( .INP(n13844), .ZN(n13843) );
  NOR2X0 U14287 ( .IN1(n13845), .IN2(n13846), .QN(n13844) );
  NAND2X0 U14288 ( .IN1(n13846), .IN2(n13845), .QN(n13842) );
  NOR2X0 U14289 ( .IN1(n13847), .IN2(n13848), .QN(n13845) );
  NOR2X0 U14290 ( .IN1(WX3481), .IN2(n8039), .QN(n13848) );
  INVX0 U14291 ( .INP(n13849), .ZN(n13847) );
  NAND2X0 U14292 ( .IN1(n8039), .IN2(WX3481), .QN(n13849) );
  NAND2X0 U14293 ( .IN1(n13850), .IN2(n13851), .QN(n13846) );
  NAND2X0 U14294 ( .IN1(n8038), .IN2(WX3353), .QN(n13851) );
  INVX0 U14295 ( .INP(n13852), .ZN(n13850) );
  NOR2X0 U14296 ( .IN1(WX3353), .IN2(n8038), .QN(n13852) );
  NAND2X0 U14297 ( .IN1(n9104), .IN2(n11391), .QN(n13840) );
  NAND2X0 U14298 ( .IN1(n13853), .IN2(n13854), .QN(n11391) );
  INVX0 U14299 ( .INP(n13855), .ZN(n13854) );
  NOR2X0 U14300 ( .IN1(n13856), .IN2(n13857), .QN(n13855) );
  NAND2X0 U14301 ( .IN1(n13857), .IN2(n13856), .QN(n13853) );
  NOR2X0 U14302 ( .IN1(n13858), .IN2(n13859), .QN(n13856) );
  NOR2X0 U14303 ( .IN1(WX2188), .IN2(n8070), .QN(n13859) );
  INVX0 U14304 ( .INP(n13860), .ZN(n13858) );
  NAND2X0 U14305 ( .IN1(n8070), .IN2(WX2188), .QN(n13860) );
  NAND2X0 U14306 ( .IN1(n13861), .IN2(n13862), .QN(n13857) );
  NAND2X0 U14307 ( .IN1(n8069), .IN2(WX2060), .QN(n13862) );
  INVX0 U14308 ( .INP(n13863), .ZN(n13861) );
  NOR2X0 U14309 ( .IN1(WX2060), .IN2(n8069), .QN(n13863) );
  NAND2X0 U14310 ( .IN1(n278), .IN2(n9284), .QN(n13839) );
  NOR2X0 U14311 ( .IN1(n9241), .IN2(n9004), .QN(n278) );
  NAND2X0 U14312 ( .IN1(n9297), .IN2(CRC_OUT_8_2), .QN(n13838) );
  NAND4X0 U14313 ( .IN1(n13864), .IN2(n13865), .IN3(n13866), .IN4(n13867), 
        .QN(WX1993) );
  NAND2X0 U14314 ( .IN1(n9326), .IN2(n13164), .QN(n13867) );
  NAND2X0 U14315 ( .IN1(n13868), .IN2(n13869), .QN(n13164) );
  INVX0 U14316 ( .INP(n13870), .ZN(n13869) );
  NOR2X0 U14317 ( .IN1(n13871), .IN2(n13872), .QN(n13870) );
  NAND2X0 U14318 ( .IN1(n13872), .IN2(n13871), .QN(n13868) );
  NOR2X0 U14319 ( .IN1(n13873), .IN2(n13874), .QN(n13871) );
  NOR2X0 U14320 ( .IN1(WX3479), .IN2(n8041), .QN(n13874) );
  INVX0 U14321 ( .INP(n13875), .ZN(n13873) );
  NAND2X0 U14322 ( .IN1(n8041), .IN2(WX3479), .QN(n13875) );
  NAND2X0 U14323 ( .IN1(n13876), .IN2(n13877), .QN(n13872) );
  NAND2X0 U14324 ( .IN1(n8040), .IN2(WX3351), .QN(n13877) );
  INVX0 U14325 ( .INP(n13878), .ZN(n13876) );
  NOR2X0 U14326 ( .IN1(WX3351), .IN2(n8040), .QN(n13878) );
  NAND2X0 U14327 ( .IN1(n9104), .IN2(n11398), .QN(n13866) );
  NAND2X0 U14328 ( .IN1(n13879), .IN2(n13880), .QN(n11398) );
  INVX0 U14329 ( .INP(n13881), .ZN(n13880) );
  NOR2X0 U14330 ( .IN1(n13882), .IN2(n13883), .QN(n13881) );
  NAND2X0 U14331 ( .IN1(n13883), .IN2(n13882), .QN(n13879) );
  NOR2X0 U14332 ( .IN1(n13884), .IN2(n13885), .QN(n13882) );
  NOR2X0 U14333 ( .IN1(WX2186), .IN2(n8072), .QN(n13885) );
  INVX0 U14334 ( .INP(n13886), .ZN(n13884) );
  NAND2X0 U14335 ( .IN1(n8072), .IN2(WX2186), .QN(n13886) );
  NAND2X0 U14336 ( .IN1(n13887), .IN2(n13888), .QN(n13883) );
  NAND2X0 U14337 ( .IN1(n8071), .IN2(WX2058), .QN(n13888) );
  INVX0 U14338 ( .INP(n13889), .ZN(n13887) );
  NOR2X0 U14339 ( .IN1(WX2058), .IN2(n8071), .QN(n13889) );
  NAND2X0 U14340 ( .IN1(n277), .IN2(n9285), .QN(n13865) );
  NOR2X0 U14341 ( .IN1(n9241), .IN2(n9005), .QN(n277) );
  NAND2X0 U14342 ( .IN1(n9297), .IN2(CRC_OUT_8_3), .QN(n13864) );
  NAND4X0 U14343 ( .IN1(n13890), .IN2(n13891), .IN3(n13892), .IN4(n13893), 
        .QN(WX1991) );
  NAND3X0 U14344 ( .IN1(n11404), .IN2(n11405), .IN3(n9090), .QN(n13893) );
  NAND3X0 U14345 ( .IN1(n13894), .IN2(n13895), .IN3(n13896), .QN(n11405) );
  INVX0 U14346 ( .INP(n13897), .ZN(n13896) );
  NAND2X0 U14347 ( .IN1(n13897), .IN2(n13898), .QN(n11404) );
  NAND2X0 U14348 ( .IN1(n13894), .IN2(n13895), .QN(n13898) );
  NAND2X0 U14349 ( .IN1(n8124), .IN2(WX2056), .QN(n13895) );
  NAND2X0 U14350 ( .IN1(n3763), .IN2(WX2184), .QN(n13894) );
  NOR2X0 U14351 ( .IN1(n13899), .IN2(n13900), .QN(n13897) );
  INVX0 U14352 ( .INP(n13901), .ZN(n13900) );
  NAND2X0 U14353 ( .IN1(test_so14), .IN2(WX2120), .QN(n13901) );
  NOR2X0 U14354 ( .IN1(WX2120), .IN2(test_so14), .QN(n13899) );
  NAND2X0 U14355 ( .IN1(n9326), .IN2(n13180), .QN(n13892) );
  NAND2X0 U14356 ( .IN1(n13902), .IN2(n13903), .QN(n13180) );
  INVX0 U14357 ( .INP(n13904), .ZN(n13903) );
  NOR2X0 U14358 ( .IN1(n13905), .IN2(n13906), .QN(n13904) );
  NAND2X0 U14359 ( .IN1(n13906), .IN2(n13905), .QN(n13902) );
  NOR2X0 U14360 ( .IN1(n13907), .IN2(n13908), .QN(n13905) );
  NOR2X0 U14361 ( .IN1(WX3477), .IN2(n8043), .QN(n13908) );
  INVX0 U14362 ( .INP(n13909), .ZN(n13907) );
  NAND2X0 U14363 ( .IN1(n8043), .IN2(WX3477), .QN(n13909) );
  NAND2X0 U14364 ( .IN1(n13910), .IN2(n13911), .QN(n13906) );
  NAND2X0 U14365 ( .IN1(n8042), .IN2(WX3349), .QN(n13911) );
  INVX0 U14366 ( .INP(n13912), .ZN(n13910) );
  NOR2X0 U14367 ( .IN1(WX3349), .IN2(n8042), .QN(n13912) );
  NAND2X0 U14368 ( .IN1(n276), .IN2(n9285), .QN(n13891) );
  NOR2X0 U14369 ( .IN1(n9241), .IN2(n9006), .QN(n276) );
  NAND2X0 U14370 ( .IN1(n9297), .IN2(CRC_OUT_8_4), .QN(n13890) );
  NAND4X0 U14371 ( .IN1(n13913), .IN2(n13914), .IN3(n13915), .IN4(n13916), 
        .QN(WX1989) );
  NAND2X0 U14372 ( .IN1(n9326), .IN2(n13196), .QN(n13916) );
  NAND2X0 U14373 ( .IN1(n13917), .IN2(n13918), .QN(n13196) );
  INVX0 U14374 ( .INP(n13919), .ZN(n13918) );
  NOR2X0 U14375 ( .IN1(n13920), .IN2(n13921), .QN(n13919) );
  NAND2X0 U14376 ( .IN1(n13921), .IN2(n13920), .QN(n13917) );
  NOR2X0 U14377 ( .IN1(n13922), .IN2(n13923), .QN(n13920) );
  NOR2X0 U14378 ( .IN1(WX3475), .IN2(n8045), .QN(n13923) );
  INVX0 U14379 ( .INP(n13924), .ZN(n13922) );
  NAND2X0 U14380 ( .IN1(n8045), .IN2(WX3475), .QN(n13924) );
  NAND2X0 U14381 ( .IN1(n13925), .IN2(n13926), .QN(n13921) );
  NAND2X0 U14382 ( .IN1(n8044), .IN2(WX3347), .QN(n13926) );
  INVX0 U14383 ( .INP(n13927), .ZN(n13925) );
  NOR2X0 U14384 ( .IN1(WX3347), .IN2(n8044), .QN(n13927) );
  NAND2X0 U14385 ( .IN1(n9104), .IN2(n11411), .QN(n13915) );
  NAND2X0 U14386 ( .IN1(n13928), .IN2(n13929), .QN(n11411) );
  INVX0 U14387 ( .INP(n13930), .ZN(n13929) );
  NOR2X0 U14388 ( .IN1(n13931), .IN2(n13932), .QN(n13930) );
  NAND2X0 U14389 ( .IN1(n13932), .IN2(n13931), .QN(n13928) );
  NOR2X0 U14390 ( .IN1(n13933), .IN2(n13934), .QN(n13931) );
  NOR2X0 U14391 ( .IN1(WX2182), .IN2(n8075), .QN(n13934) );
  INVX0 U14392 ( .INP(n13935), .ZN(n13933) );
  NAND2X0 U14393 ( .IN1(n8075), .IN2(WX2182), .QN(n13935) );
  NAND2X0 U14394 ( .IN1(n13936), .IN2(n13937), .QN(n13932) );
  NAND2X0 U14395 ( .IN1(n8074), .IN2(WX2054), .QN(n13937) );
  INVX0 U14396 ( .INP(n13938), .ZN(n13936) );
  NOR2X0 U14397 ( .IN1(WX2054), .IN2(n8074), .QN(n13938) );
  NAND2X0 U14398 ( .IN1(n275), .IN2(n9285), .QN(n13914) );
  NOR2X0 U14399 ( .IN1(n9241), .IN2(n9007), .QN(n275) );
  NAND2X0 U14400 ( .IN1(n9298), .IN2(CRC_OUT_8_5), .QN(n13913) );
  NAND4X0 U14401 ( .IN1(n13939), .IN2(n13940), .IN3(n13941), .IN4(n13942), 
        .QN(WX1987) );
  NAND3X0 U14402 ( .IN1(n13201), .IN2(n13202), .IN3(n9321), .QN(n13942) );
  NAND3X0 U14403 ( .IN1(n13943), .IN2(n13944), .IN3(n13945), .QN(n13202) );
  INVX0 U14404 ( .INP(n13946), .ZN(n13945) );
  NAND2X0 U14405 ( .IN1(n13946), .IN2(n13947), .QN(n13201) );
  NAND2X0 U14406 ( .IN1(n13943), .IN2(n13944), .QN(n13947) );
  NAND2X0 U14407 ( .IN1(n8047), .IN2(WX3345), .QN(n13944) );
  NAND2X0 U14408 ( .IN1(n3735), .IN2(WX3409), .QN(n13943) );
  NOR2X0 U14409 ( .IN1(n13948), .IN2(n13949), .QN(n13946) );
  NOR2X0 U14410 ( .IN1(n8791), .IN2(n8046), .QN(n13949) );
  INVX0 U14411 ( .INP(n13950), .ZN(n13948) );
  NAND2X0 U14412 ( .IN1(n8046), .IN2(n8791), .QN(n13950) );
  NAND2X0 U14413 ( .IN1(n9104), .IN2(n11417), .QN(n13941) );
  NAND2X0 U14414 ( .IN1(n13951), .IN2(n13952), .QN(n11417) );
  INVX0 U14415 ( .INP(n13953), .ZN(n13952) );
  NOR2X0 U14416 ( .IN1(n13954), .IN2(n13955), .QN(n13953) );
  NAND2X0 U14417 ( .IN1(n13955), .IN2(n13954), .QN(n13951) );
  NOR2X0 U14418 ( .IN1(n13956), .IN2(n13957), .QN(n13954) );
  NOR2X0 U14419 ( .IN1(WX2180), .IN2(n8077), .QN(n13957) );
  INVX0 U14420 ( .INP(n13958), .ZN(n13956) );
  NAND2X0 U14421 ( .IN1(n8077), .IN2(WX2180), .QN(n13958) );
  NAND2X0 U14422 ( .IN1(n13959), .IN2(n13960), .QN(n13955) );
  NAND2X0 U14423 ( .IN1(n8076), .IN2(WX2052), .QN(n13960) );
  INVX0 U14424 ( .INP(n13961), .ZN(n13959) );
  NOR2X0 U14425 ( .IN1(WX2052), .IN2(n8076), .QN(n13961) );
  NAND2X0 U14426 ( .IN1(n274), .IN2(n9285), .QN(n13940) );
  NOR2X0 U14427 ( .IN1(n9241), .IN2(n9008), .QN(n274) );
  NAND2X0 U14428 ( .IN1(n9298), .IN2(CRC_OUT_8_6), .QN(n13939) );
  NAND4X0 U14429 ( .IN1(n13962), .IN2(n13963), .IN3(n13964), .IN4(n13965), 
        .QN(WX1985) );
  NAND2X0 U14430 ( .IN1(n9326), .IN2(n13229), .QN(n13965) );
  NAND2X0 U14431 ( .IN1(n13966), .IN2(n13967), .QN(n13229) );
  INVX0 U14432 ( .INP(n13968), .ZN(n13967) );
  NOR2X0 U14433 ( .IN1(n13969), .IN2(n13970), .QN(n13968) );
  NAND2X0 U14434 ( .IN1(n13970), .IN2(n13969), .QN(n13966) );
  NOR2X0 U14435 ( .IN1(n13971), .IN2(n13972), .QN(n13969) );
  NOR2X0 U14436 ( .IN1(WX3471), .IN2(n8049), .QN(n13972) );
  INVX0 U14437 ( .INP(n13973), .ZN(n13971) );
  NAND2X0 U14438 ( .IN1(n8049), .IN2(WX3471), .QN(n13973) );
  NAND2X0 U14439 ( .IN1(n13974), .IN2(n13975), .QN(n13970) );
  NAND2X0 U14440 ( .IN1(n8048), .IN2(WX3343), .QN(n13975) );
  INVX0 U14441 ( .INP(n13976), .ZN(n13974) );
  NOR2X0 U14442 ( .IN1(WX3343), .IN2(n8048), .QN(n13976) );
  NAND2X0 U14443 ( .IN1(n9104), .IN2(n11424), .QN(n13964) );
  NAND2X0 U14444 ( .IN1(n13977), .IN2(n13978), .QN(n11424) );
  INVX0 U14445 ( .INP(n13979), .ZN(n13978) );
  NOR2X0 U14446 ( .IN1(n13980), .IN2(n13981), .QN(n13979) );
  NAND2X0 U14447 ( .IN1(n13981), .IN2(n13980), .QN(n13977) );
  NOR2X0 U14448 ( .IN1(n13982), .IN2(n13983), .QN(n13980) );
  NOR2X0 U14449 ( .IN1(WX2178), .IN2(n8079), .QN(n13983) );
  INVX0 U14450 ( .INP(n13984), .ZN(n13982) );
  NAND2X0 U14451 ( .IN1(n8079), .IN2(WX2178), .QN(n13984) );
  NAND2X0 U14452 ( .IN1(n13985), .IN2(n13986), .QN(n13981) );
  NAND2X0 U14453 ( .IN1(n8078), .IN2(WX2050), .QN(n13986) );
  INVX0 U14454 ( .INP(n13987), .ZN(n13985) );
  NOR2X0 U14455 ( .IN1(WX2050), .IN2(n8078), .QN(n13987) );
  NAND2X0 U14456 ( .IN1(n273), .IN2(n9285), .QN(n13963) );
  NOR2X0 U14457 ( .IN1(n9241), .IN2(n9009), .QN(n273) );
  NAND2X0 U14458 ( .IN1(test_so20), .IN2(n9314), .QN(n13962) );
  NAND4X0 U14459 ( .IN1(n13988), .IN2(n13989), .IN3(n13990), .IN4(n13991), 
        .QN(WX1983) );
  NAND3X0 U14460 ( .IN1(n13234), .IN2(n13235), .IN3(n9321), .QN(n13991) );
  NAND3X0 U14461 ( .IN1(n13992), .IN2(n13993), .IN3(n13994), .QN(n13235) );
  INVX0 U14462 ( .INP(n13995), .ZN(n13994) );
  NAND2X0 U14463 ( .IN1(n13995), .IN2(n13996), .QN(n13234) );
  NAND2X0 U14464 ( .IN1(n13992), .IN2(n13993), .QN(n13996) );
  NAND2X0 U14465 ( .IN1(n8534), .IN2(WX3341), .QN(n13993) );
  NAND2X0 U14466 ( .IN1(n3739), .IN2(WX3469), .QN(n13992) );
  NOR2X0 U14467 ( .IN1(n13997), .IN2(n13998), .QN(n13995) );
  INVX0 U14468 ( .INP(n13999), .ZN(n13998) );
  NAND2X0 U14469 ( .IN1(test_so28), .IN2(WX3277), .QN(n13999) );
  NOR2X0 U14470 ( .IN1(WX3277), .IN2(test_so28), .QN(n13997) );
  NAND2X0 U14471 ( .IN1(n9104), .IN2(n11430), .QN(n13990) );
  NAND2X0 U14472 ( .IN1(n14000), .IN2(n14001), .QN(n11430) );
  INVX0 U14473 ( .INP(n14002), .ZN(n14001) );
  NOR2X0 U14474 ( .IN1(n14003), .IN2(n14004), .QN(n14002) );
  NAND2X0 U14475 ( .IN1(n14004), .IN2(n14003), .QN(n14000) );
  NOR2X0 U14476 ( .IN1(n14005), .IN2(n14006), .QN(n14003) );
  NOR2X0 U14477 ( .IN1(WX2176), .IN2(n8081), .QN(n14006) );
  INVX0 U14478 ( .INP(n14007), .ZN(n14005) );
  NAND2X0 U14479 ( .IN1(n8081), .IN2(WX2176), .QN(n14007) );
  NAND2X0 U14480 ( .IN1(n14008), .IN2(n14009), .QN(n14004) );
  NAND2X0 U14481 ( .IN1(n8080), .IN2(WX2048), .QN(n14009) );
  INVX0 U14482 ( .INP(n14010), .ZN(n14008) );
  NOR2X0 U14483 ( .IN1(WX2048), .IN2(n8080), .QN(n14010) );
  NAND2X0 U14484 ( .IN1(n272), .IN2(n9285), .QN(n13989) );
  NOR2X0 U14485 ( .IN1(n9072), .IN2(n9161), .QN(n272) );
  NAND2X0 U14486 ( .IN1(n9298), .IN2(CRC_OUT_8_8), .QN(n13988) );
  NAND4X0 U14487 ( .IN1(n14011), .IN2(n14012), .IN3(n14013), .IN4(n14014), 
        .QN(WX1981) );
  NAND2X0 U14488 ( .IN1(n9326), .IN2(n13262), .QN(n14014) );
  NAND2X0 U14489 ( .IN1(n14015), .IN2(n14016), .QN(n13262) );
  INVX0 U14490 ( .INP(n14017), .ZN(n14016) );
  NOR2X0 U14491 ( .IN1(n14018), .IN2(n14019), .QN(n14017) );
  NAND2X0 U14492 ( .IN1(n14019), .IN2(n14018), .QN(n14015) );
  NOR2X0 U14493 ( .IN1(n14020), .IN2(n14021), .QN(n14018) );
  NOR2X0 U14494 ( .IN1(WX3467), .IN2(n8052), .QN(n14021) );
  INVX0 U14495 ( .INP(n14022), .ZN(n14020) );
  NAND2X0 U14496 ( .IN1(n8052), .IN2(WX3467), .QN(n14022) );
  NAND2X0 U14497 ( .IN1(n14023), .IN2(n14024), .QN(n14019) );
  NAND2X0 U14498 ( .IN1(n8051), .IN2(WX3339), .QN(n14024) );
  INVX0 U14499 ( .INP(n14025), .ZN(n14023) );
  NOR2X0 U14500 ( .IN1(WX3339), .IN2(n8051), .QN(n14025) );
  NAND2X0 U14501 ( .IN1(n9104), .IN2(n11436), .QN(n14013) );
  NAND2X0 U14502 ( .IN1(n14026), .IN2(n14027), .QN(n11436) );
  INVX0 U14503 ( .INP(n14028), .ZN(n14027) );
  NOR2X0 U14504 ( .IN1(n14029), .IN2(n14030), .QN(n14028) );
  NAND2X0 U14505 ( .IN1(n14030), .IN2(n14029), .QN(n14026) );
  NOR2X0 U14506 ( .IN1(n14031), .IN2(n14032), .QN(n14029) );
  NOR2X0 U14507 ( .IN1(WX2174), .IN2(n8083), .QN(n14032) );
  INVX0 U14508 ( .INP(n14033), .ZN(n14031) );
  NAND2X0 U14509 ( .IN1(n8083), .IN2(WX2174), .QN(n14033) );
  NAND2X0 U14510 ( .IN1(n14034), .IN2(n14035), .QN(n14030) );
  NAND2X0 U14511 ( .IN1(n8082), .IN2(WX2046), .QN(n14035) );
  INVX0 U14512 ( .INP(n14036), .ZN(n14034) );
  NOR2X0 U14513 ( .IN1(WX2046), .IN2(n8082), .QN(n14036) );
  NAND2X0 U14514 ( .IN1(n271), .IN2(n9285), .QN(n14012) );
  NOR2X0 U14515 ( .IN1(n9241), .IN2(n9010), .QN(n271) );
  NAND2X0 U14516 ( .IN1(n9298), .IN2(CRC_OUT_8_9), .QN(n14011) );
  NAND4X0 U14517 ( .IN1(n14037), .IN2(n14038), .IN3(n14039), .IN4(n14040), 
        .QN(WX1979) );
  NAND3X0 U14518 ( .IN1(n11442), .IN2(n11443), .IN3(n9090), .QN(n14040) );
  NAND3X0 U14519 ( .IN1(n14041), .IN2(n14042), .IN3(n14043), .QN(n11443) );
  INVX0 U14520 ( .INP(n14044), .ZN(n14043) );
  NAND2X0 U14521 ( .IN1(n14044), .IN2(n14045), .QN(n11442) );
  NAND2X0 U14522 ( .IN1(n14041), .IN2(n14042), .QN(n14045) );
  NAND2X0 U14523 ( .IN1(n8085), .IN2(WX2044), .QN(n14042) );
  NAND2X0 U14524 ( .IN1(n3775), .IN2(WX2108), .QN(n14041) );
  NOR2X0 U14525 ( .IN1(n14046), .IN2(n14047), .QN(n14044) );
  NOR2X0 U14526 ( .IN1(n8792), .IN2(n8084), .QN(n14047) );
  INVX0 U14527 ( .INP(n14048), .ZN(n14046) );
  NAND2X0 U14528 ( .IN1(n8084), .IN2(n8792), .QN(n14048) );
  NAND2X0 U14529 ( .IN1(n9327), .IN2(n13278), .QN(n14039) );
  NAND2X0 U14530 ( .IN1(n14049), .IN2(n14050), .QN(n13278) );
  INVX0 U14531 ( .INP(n14051), .ZN(n14050) );
  NOR2X0 U14532 ( .IN1(n14052), .IN2(n14053), .QN(n14051) );
  NAND2X0 U14533 ( .IN1(n14053), .IN2(n14052), .QN(n14049) );
  NOR2X0 U14534 ( .IN1(n14054), .IN2(n14055), .QN(n14052) );
  NOR2X0 U14535 ( .IN1(WX3465), .IN2(n8054), .QN(n14055) );
  INVX0 U14536 ( .INP(n14056), .ZN(n14054) );
  NAND2X0 U14537 ( .IN1(n8054), .IN2(WX3465), .QN(n14056) );
  NAND2X0 U14538 ( .IN1(n14057), .IN2(n14058), .QN(n14053) );
  NAND2X0 U14539 ( .IN1(n8053), .IN2(WX3337), .QN(n14058) );
  INVX0 U14540 ( .INP(n14059), .ZN(n14057) );
  NOR2X0 U14541 ( .IN1(WX3337), .IN2(n8053), .QN(n14059) );
  NAND2X0 U14542 ( .IN1(n270), .IN2(n9285), .QN(n14038) );
  NOR2X0 U14543 ( .IN1(n9241), .IN2(n9011), .QN(n270) );
  NAND2X0 U14544 ( .IN1(n9298), .IN2(CRC_OUT_8_10), .QN(n14037) );
  NAND4X0 U14545 ( .IN1(n14060), .IN2(n14061), .IN3(n14062), .IN4(n14063), 
        .QN(WX1977) );
  NAND2X0 U14546 ( .IN1(n9327), .IN2(n13291), .QN(n14063) );
  NAND2X0 U14547 ( .IN1(n14064), .IN2(n14065), .QN(n13291) );
  INVX0 U14548 ( .INP(n14066), .ZN(n14065) );
  NOR2X0 U14549 ( .IN1(n14067), .IN2(n14068), .QN(n14066) );
  NAND2X0 U14550 ( .IN1(n14068), .IN2(n14067), .QN(n14064) );
  NOR2X0 U14551 ( .IN1(n14069), .IN2(n14070), .QN(n14067) );
  NOR2X0 U14552 ( .IN1(WX3463), .IN2(n8056), .QN(n14070) );
  INVX0 U14553 ( .INP(n14071), .ZN(n14069) );
  NAND2X0 U14554 ( .IN1(n8056), .IN2(WX3463), .QN(n14071) );
  NAND2X0 U14555 ( .IN1(n14072), .IN2(n14073), .QN(n14068) );
  NAND2X0 U14556 ( .IN1(n8055), .IN2(WX3335), .QN(n14073) );
  INVX0 U14557 ( .INP(n14074), .ZN(n14072) );
  NOR2X0 U14558 ( .IN1(WX3335), .IN2(n8055), .QN(n14074) );
  NAND2X0 U14559 ( .IN1(n9104), .IN2(n11450), .QN(n14062) );
  NAND2X0 U14560 ( .IN1(n14075), .IN2(n14076), .QN(n11450) );
  INVX0 U14561 ( .INP(n14077), .ZN(n14076) );
  NOR2X0 U14562 ( .IN1(n14078), .IN2(n14079), .QN(n14077) );
  NAND2X0 U14563 ( .IN1(n14079), .IN2(n14078), .QN(n14075) );
  NOR2X0 U14564 ( .IN1(n14080), .IN2(n14081), .QN(n14078) );
  NOR2X0 U14565 ( .IN1(WX2170), .IN2(n8087), .QN(n14081) );
  INVX0 U14566 ( .INP(n14082), .ZN(n14080) );
  NAND2X0 U14567 ( .IN1(n8087), .IN2(WX2170), .QN(n14082) );
  NAND2X0 U14568 ( .IN1(n14083), .IN2(n14084), .QN(n14079) );
  NAND2X0 U14569 ( .IN1(n8086), .IN2(WX2042), .QN(n14084) );
  INVX0 U14570 ( .INP(n14085), .ZN(n14083) );
  NOR2X0 U14571 ( .IN1(WX2042), .IN2(n8086), .QN(n14085) );
  NAND2X0 U14572 ( .IN1(n269), .IN2(n9285), .QN(n14061) );
  NOR2X0 U14573 ( .IN1(n9241), .IN2(n9012), .QN(n269) );
  NAND2X0 U14574 ( .IN1(n9298), .IN2(CRC_OUT_8_11), .QN(n14060) );
  NAND4X0 U14575 ( .IN1(n14086), .IN2(n14087), .IN3(n14088), .IN4(n14089), 
        .QN(WX1975) );
  NAND3X0 U14576 ( .IN1(n13296), .IN2(n13297), .IN3(n9320), .QN(n14089) );
  NAND3X0 U14577 ( .IN1(n14090), .IN2(n14091), .IN3(n14092), .QN(n13297) );
  INVX0 U14578 ( .INP(n14093), .ZN(n14092) );
  NAND2X0 U14579 ( .IN1(n14093), .IN2(n14094), .QN(n13296) );
  NAND2X0 U14580 ( .IN1(n14090), .IN2(n14091), .QN(n14094) );
  NAND2X0 U14581 ( .IN1(n8531), .IN2(WX3397), .QN(n14091) );
  NAND2X0 U14582 ( .IN1(n8058), .IN2(WX3461), .QN(n14090) );
  NOR2X0 U14583 ( .IN1(n14095), .IN2(n14096), .QN(n14093) );
  INVX0 U14584 ( .INP(n14097), .ZN(n14096) );
  NAND2X0 U14585 ( .IN1(test_so26), .IN2(WX3269), .QN(n14097) );
  NOR2X0 U14586 ( .IN1(WX3269), .IN2(test_so26), .QN(n14095) );
  NAND2X0 U14587 ( .IN1(n9104), .IN2(n11456), .QN(n14088) );
  NAND2X0 U14588 ( .IN1(n14098), .IN2(n14099), .QN(n11456) );
  INVX0 U14589 ( .INP(n14100), .ZN(n14099) );
  NOR2X0 U14590 ( .IN1(n14101), .IN2(n14102), .QN(n14100) );
  NAND2X0 U14591 ( .IN1(n14102), .IN2(n14101), .QN(n14098) );
  NOR2X0 U14592 ( .IN1(n14103), .IN2(n14104), .QN(n14101) );
  NOR2X0 U14593 ( .IN1(WX2168), .IN2(n8089), .QN(n14104) );
  INVX0 U14594 ( .INP(n14105), .ZN(n14103) );
  NAND2X0 U14595 ( .IN1(n8089), .IN2(WX2168), .QN(n14105) );
  NAND2X0 U14596 ( .IN1(n14106), .IN2(n14107), .QN(n14102) );
  NAND2X0 U14597 ( .IN1(n8088), .IN2(WX2040), .QN(n14107) );
  INVX0 U14598 ( .INP(n14108), .ZN(n14106) );
  NOR2X0 U14599 ( .IN1(WX2040), .IN2(n8088), .QN(n14108) );
  NAND2X0 U14600 ( .IN1(n268), .IN2(n9285), .QN(n14087) );
  NOR2X0 U14601 ( .IN1(n9241), .IN2(n9013), .QN(n268) );
  NAND2X0 U14602 ( .IN1(n9298), .IN2(CRC_OUT_8_12), .QN(n14086) );
  NAND4X0 U14603 ( .IN1(n14109), .IN2(n14110), .IN3(n14111), .IN4(n14112), 
        .QN(WX1973) );
  NAND2X0 U14604 ( .IN1(n9327), .IN2(n13321), .QN(n14112) );
  NAND2X0 U14605 ( .IN1(n14113), .IN2(n14114), .QN(n13321) );
  INVX0 U14606 ( .INP(n14115), .ZN(n14114) );
  NOR2X0 U14607 ( .IN1(n14116), .IN2(n14117), .QN(n14115) );
  NAND2X0 U14608 ( .IN1(n14117), .IN2(n14116), .QN(n14113) );
  NOR2X0 U14609 ( .IN1(n14118), .IN2(n14119), .QN(n14116) );
  NOR2X0 U14610 ( .IN1(WX3459), .IN2(n8060), .QN(n14119) );
  INVX0 U14611 ( .INP(n14120), .ZN(n14118) );
  NAND2X0 U14612 ( .IN1(n8060), .IN2(WX3459), .QN(n14120) );
  NAND2X0 U14613 ( .IN1(n14121), .IN2(n14122), .QN(n14117) );
  NAND2X0 U14614 ( .IN1(n8059), .IN2(WX3331), .QN(n14122) );
  INVX0 U14615 ( .INP(n14123), .ZN(n14121) );
  NOR2X0 U14616 ( .IN1(WX3331), .IN2(n8059), .QN(n14123) );
  NAND2X0 U14617 ( .IN1(n9104), .IN2(n11462), .QN(n14111) );
  NAND2X0 U14618 ( .IN1(n14124), .IN2(n14125), .QN(n11462) );
  INVX0 U14619 ( .INP(n14126), .ZN(n14125) );
  NOR2X0 U14620 ( .IN1(n14127), .IN2(n14128), .QN(n14126) );
  NAND2X0 U14621 ( .IN1(n14128), .IN2(n14127), .QN(n14124) );
  NOR2X0 U14622 ( .IN1(n14129), .IN2(n14130), .QN(n14127) );
  NOR2X0 U14623 ( .IN1(WX2166), .IN2(n8091), .QN(n14130) );
  INVX0 U14624 ( .INP(n14131), .ZN(n14129) );
  NAND2X0 U14625 ( .IN1(n8091), .IN2(WX2166), .QN(n14131) );
  NAND2X0 U14626 ( .IN1(n14132), .IN2(n14133), .QN(n14128) );
  NAND2X0 U14627 ( .IN1(n8090), .IN2(WX2038), .QN(n14133) );
  INVX0 U14628 ( .INP(n14134), .ZN(n14132) );
  NOR2X0 U14629 ( .IN1(WX2038), .IN2(n8090), .QN(n14134) );
  NAND2X0 U14630 ( .IN1(n267), .IN2(n9285), .QN(n14110) );
  NOR2X0 U14631 ( .IN1(n9241), .IN2(n9014), .QN(n267) );
  NAND2X0 U14632 ( .IN1(n9298), .IN2(CRC_OUT_8_13), .QN(n14109) );
  NAND4X0 U14633 ( .IN1(n14135), .IN2(n14136), .IN3(n14137), .IN4(n14138), 
        .QN(WX1971) );
  NAND3X0 U14634 ( .IN1(n11468), .IN2(n11469), .IN3(n9090), .QN(n14138) );
  NAND3X0 U14635 ( .IN1(n14139), .IN2(n14140), .IN3(n14141), .QN(n11469) );
  INVX0 U14636 ( .INP(n14142), .ZN(n14141) );
  NAND2X0 U14637 ( .IN1(n14142), .IN2(n14143), .QN(n11468) );
  NAND2X0 U14638 ( .IN1(n14139), .IN2(n14140), .QN(n14143) );
  NAND2X0 U14639 ( .IN1(n8633), .IN2(WX2036), .QN(n14140) );
  NAND2X0 U14640 ( .IN1(n3783), .IN2(WX2164), .QN(n14139) );
  NOR2X0 U14641 ( .IN1(n14144), .IN2(n14145), .QN(n14142) );
  INVX0 U14642 ( .INP(n14146), .ZN(n14145) );
  NAND2X0 U14643 ( .IN1(test_so17), .IN2(WX1972), .QN(n14146) );
  NOR2X0 U14644 ( .IN1(WX1972), .IN2(test_so17), .QN(n14144) );
  NAND2X0 U14645 ( .IN1(n9327), .IN2(n13337), .QN(n14137) );
  NAND2X0 U14646 ( .IN1(n14147), .IN2(n14148), .QN(n13337) );
  INVX0 U14647 ( .INP(n14149), .ZN(n14148) );
  NOR2X0 U14648 ( .IN1(n14150), .IN2(n14151), .QN(n14149) );
  NAND2X0 U14649 ( .IN1(n14151), .IN2(n14150), .QN(n14147) );
  NOR2X0 U14650 ( .IN1(n14152), .IN2(n14153), .QN(n14150) );
  NOR2X0 U14651 ( .IN1(WX3457), .IN2(n8062), .QN(n14153) );
  INVX0 U14652 ( .INP(n14154), .ZN(n14152) );
  NAND2X0 U14653 ( .IN1(n8062), .IN2(WX3457), .QN(n14154) );
  NAND2X0 U14654 ( .IN1(n14155), .IN2(n14156), .QN(n14151) );
  NAND2X0 U14655 ( .IN1(n8061), .IN2(WX3329), .QN(n14156) );
  INVX0 U14656 ( .INP(n14157), .ZN(n14155) );
  NOR2X0 U14657 ( .IN1(WX3329), .IN2(n8061), .QN(n14157) );
  NAND2X0 U14658 ( .IN1(n266), .IN2(n9285), .QN(n14136) );
  NOR2X0 U14659 ( .IN1(n9241), .IN2(n9015), .QN(n266) );
  NAND2X0 U14660 ( .IN1(n9298), .IN2(CRC_OUT_8_14), .QN(n14135) );
  NAND4X0 U14661 ( .IN1(n14158), .IN2(n14159), .IN3(n14160), .IN4(n14161), 
        .QN(WX1969) );
  NAND2X0 U14662 ( .IN1(n9327), .IN2(n13350), .QN(n14161) );
  NAND2X0 U14663 ( .IN1(n14162), .IN2(n14163), .QN(n13350) );
  INVX0 U14664 ( .INP(n14164), .ZN(n14163) );
  NOR2X0 U14665 ( .IN1(n14165), .IN2(n14166), .QN(n14164) );
  NAND2X0 U14666 ( .IN1(n14166), .IN2(n14165), .QN(n14162) );
  NOR2X0 U14667 ( .IN1(n14167), .IN2(n14168), .QN(n14165) );
  NOR2X0 U14668 ( .IN1(WX3455), .IN2(n8064), .QN(n14168) );
  INVX0 U14669 ( .INP(n14169), .ZN(n14167) );
  NAND2X0 U14670 ( .IN1(n8064), .IN2(WX3455), .QN(n14169) );
  NAND2X0 U14671 ( .IN1(n14170), .IN2(n14171), .QN(n14166) );
  NAND2X0 U14672 ( .IN1(n8063), .IN2(WX3327), .QN(n14171) );
  INVX0 U14673 ( .INP(n14172), .ZN(n14170) );
  NOR2X0 U14674 ( .IN1(WX3327), .IN2(n8063), .QN(n14172) );
  NAND2X0 U14675 ( .IN1(n9104), .IN2(n11475), .QN(n14160) );
  NAND2X0 U14676 ( .IN1(n14173), .IN2(n14174), .QN(n11475) );
  INVX0 U14677 ( .INP(n14175), .ZN(n14174) );
  NOR2X0 U14678 ( .IN1(n14176), .IN2(n14177), .QN(n14175) );
  NAND2X0 U14679 ( .IN1(n14177), .IN2(n14176), .QN(n14173) );
  NOR2X0 U14680 ( .IN1(n14178), .IN2(n14179), .QN(n14176) );
  NOR2X0 U14681 ( .IN1(WX2162), .IN2(n8094), .QN(n14179) );
  INVX0 U14682 ( .INP(n14180), .ZN(n14178) );
  NAND2X0 U14683 ( .IN1(n8094), .IN2(WX2162), .QN(n14180) );
  NAND2X0 U14684 ( .IN1(n14181), .IN2(n14182), .QN(n14177) );
  NAND2X0 U14685 ( .IN1(n8093), .IN2(WX2034), .QN(n14182) );
  INVX0 U14686 ( .INP(n14183), .ZN(n14181) );
  NOR2X0 U14687 ( .IN1(WX2034), .IN2(n8093), .QN(n14183) );
  NAND2X0 U14688 ( .IN1(n265), .IN2(n9285), .QN(n14159) );
  NOR2X0 U14689 ( .IN1(n9226), .IN2(n9016), .QN(n265) );
  NAND2X0 U14690 ( .IN1(n9298), .IN2(CRC_OUT_8_15), .QN(n14158) );
  NAND4X0 U14691 ( .IN1(n14184), .IN2(n14185), .IN3(n14186), .IN4(n14187), 
        .QN(WX1967) );
  NAND2X0 U14692 ( .IN1(n14188), .IN2(n13370), .QN(n14187) );
  NAND3X0 U14693 ( .IN1(n14189), .IN2(n14190), .IN3(n13373), .QN(n13370) );
  NAND2X0 U14694 ( .IN1(n8119), .IN2(n9120), .QN(n14190) );
  NAND2X0 U14695 ( .IN1(TM1), .IN2(WX3453), .QN(n14189) );
  NAND3X0 U14696 ( .IN1(n14191), .IN2(n14192), .IN3(n14193), .QN(n14188) );
  NAND2X0 U14697 ( .IN1(n9327), .IN2(n13373), .QN(n14193) );
  NAND2X0 U14698 ( .IN1(n14194), .IN2(n14195), .QN(n13373) );
  NAND2X0 U14699 ( .IN1(n14196), .IN2(WX3389), .QN(n14195) );
  NAND2X0 U14700 ( .IN1(n14197), .IN2(n14198), .QN(n14196) );
  NAND3X0 U14701 ( .IN1(n14197), .IN2(n14198), .IN3(n7797), .QN(n14194) );
  NAND2X0 U14702 ( .IN1(test_so24), .IN2(WX3325), .QN(n14198) );
  NAND2X0 U14703 ( .IN1(n7796), .IN2(n8823), .QN(n14197) );
  NAND2X0 U14704 ( .IN1(n9078), .IN2(WX3453), .QN(n14192) );
  NAND2X0 U14705 ( .IN1(n9082), .IN2(n8119), .QN(n14191) );
  NAND2X0 U14706 ( .IN1(n14199), .IN2(n11482), .QN(n14186) );
  NAND2X0 U14707 ( .IN1(n14200), .IN2(n11486), .QN(n11482) );
  NAND2X0 U14708 ( .IN1(n14201), .IN2(n14202), .QN(n14200) );
  NAND2X0 U14709 ( .IN1(n16041), .IN2(n9120), .QN(n14202) );
  NAND2X0 U14710 ( .IN1(TM1), .IN2(n8653), .QN(n14201) );
  NAND2X0 U14711 ( .IN1(n14203), .IN2(n14204), .QN(n14199) );
  NAND2X0 U14712 ( .IN1(n9103), .IN2(n11486), .QN(n14204) );
  NAND2X0 U14713 ( .IN1(n14205), .IN2(n14206), .QN(n11486) );
  NAND2X0 U14714 ( .IN1(n7824), .IN2(n14207), .QN(n14206) );
  INVX0 U14715 ( .INP(n14208), .ZN(n14205) );
  NOR2X0 U14716 ( .IN1(n14207), .IN2(n7824), .QN(n14208) );
  NOR2X0 U14717 ( .IN1(n14209), .IN2(n14210), .QN(n14207) );
  NOR2X0 U14718 ( .IN1(WX2160), .IN2(n7825), .QN(n14210) );
  INVX0 U14719 ( .INP(n14211), .ZN(n14209) );
  NAND2X0 U14720 ( .IN1(n7825), .IN2(WX2160), .QN(n14211) );
  NAND2X0 U14721 ( .IN1(n9103), .IN2(n8653), .QN(n14203) );
  NAND2X0 U14722 ( .IN1(n264), .IN2(n9285), .QN(n14185) );
  NOR2X0 U14723 ( .IN1(n9226), .IN2(n9017), .QN(n264) );
  NAND2X0 U14724 ( .IN1(n9298), .IN2(CRC_OUT_8_16), .QN(n14184) );
  NAND4X0 U14725 ( .IN1(n14212), .IN2(n14213), .IN3(n14214), .IN4(n14215), 
        .QN(WX1965) );
  NAND2X0 U14726 ( .IN1(n14216), .IN2(n13390), .QN(n14215) );
  NAND2X0 U14727 ( .IN1(n14217), .IN2(n13393), .QN(n13390) );
  NAND2X0 U14728 ( .IN1(n14218), .IN2(n14219), .QN(n14217) );
  NAND2X0 U14729 ( .IN1(n16056), .IN2(n9121), .QN(n14219) );
  NAND2X0 U14730 ( .IN1(TM1), .IN2(n8597), .QN(n14218) );
  NAND3X0 U14731 ( .IN1(n14220), .IN2(n14221), .IN3(n14222), .QN(n14216) );
  NAND2X0 U14732 ( .IN1(n9327), .IN2(n13393), .QN(n14222) );
  NAND2X0 U14733 ( .IN1(n14223), .IN2(n14224), .QN(n13393) );
  NAND2X0 U14734 ( .IN1(n7798), .IN2(n14225), .QN(n14224) );
  INVX0 U14735 ( .INP(n14226), .ZN(n14223) );
  NOR2X0 U14736 ( .IN1(n14225), .IN2(n7798), .QN(n14226) );
  NOR2X0 U14737 ( .IN1(n14227), .IN2(n14228), .QN(n14225) );
  NOR2X0 U14738 ( .IN1(WX3451), .IN2(n7799), .QN(n14228) );
  INVX0 U14739 ( .INP(n14229), .ZN(n14227) );
  NAND2X0 U14740 ( .IN1(n7799), .IN2(WX3451), .QN(n14229) );
  NAND2X0 U14741 ( .IN1(n9081), .IN2(n8597), .QN(n14221) );
  NAND2X0 U14742 ( .IN1(n16056), .IN2(n9077), .QN(n14220) );
  NAND2X0 U14743 ( .IN1(n14230), .IN2(n11494), .QN(n14214) );
  NAND2X0 U14744 ( .IN1(n14231), .IN2(n11498), .QN(n11494) );
  NAND2X0 U14745 ( .IN1(n14232), .IN2(n14233), .QN(n14231) );
  NAND2X0 U14746 ( .IN1(n16040), .IN2(n9121), .QN(n14233) );
  NAND2X0 U14747 ( .IN1(TM1), .IN2(n8654), .QN(n14232) );
  NAND2X0 U14748 ( .IN1(n14234), .IN2(n14235), .QN(n14230) );
  NAND2X0 U14749 ( .IN1(n9103), .IN2(n11498), .QN(n14235) );
  NAND2X0 U14750 ( .IN1(n14236), .IN2(n14237), .QN(n11498) );
  NAND2X0 U14751 ( .IN1(n7826), .IN2(n14238), .QN(n14237) );
  INVX0 U14752 ( .INP(n14239), .ZN(n14236) );
  NOR2X0 U14753 ( .IN1(n14238), .IN2(n7826), .QN(n14239) );
  NOR2X0 U14754 ( .IN1(n14240), .IN2(n14241), .QN(n14238) );
  NOR2X0 U14755 ( .IN1(WX2158), .IN2(n7827), .QN(n14241) );
  INVX0 U14756 ( .INP(n14242), .ZN(n14240) );
  NAND2X0 U14757 ( .IN1(n7827), .IN2(WX2158), .QN(n14242) );
  NAND2X0 U14758 ( .IN1(n9103), .IN2(n8654), .QN(n14234) );
  NAND2X0 U14759 ( .IN1(n263), .IN2(n9285), .QN(n14213) );
  NOR2X0 U14760 ( .IN1(n9226), .IN2(n9018), .QN(n263) );
  NAND2X0 U14761 ( .IN1(n9298), .IN2(CRC_OUT_8_17), .QN(n14212) );
  NAND4X0 U14762 ( .IN1(n14243), .IN2(n14244), .IN3(n14245), .IN4(n14246), 
        .QN(WX1963) );
  NAND2X0 U14763 ( .IN1(n14247), .IN2(n13413), .QN(n14246) );
  NAND2X0 U14764 ( .IN1(n14248), .IN2(n13416), .QN(n13413) );
  NAND2X0 U14765 ( .IN1(n14249), .IN2(n14250), .QN(n14248) );
  NAND2X0 U14766 ( .IN1(n16055), .IN2(n9121), .QN(n14250) );
  NAND2X0 U14767 ( .IN1(TM1), .IN2(n8598), .QN(n14249) );
  NAND3X0 U14768 ( .IN1(n14251), .IN2(n14252), .IN3(n14253), .QN(n14247) );
  NAND2X0 U14769 ( .IN1(n9327), .IN2(n13416), .QN(n14253) );
  NAND2X0 U14770 ( .IN1(n14254), .IN2(n14255), .QN(n13416) );
  NAND2X0 U14771 ( .IN1(n7800), .IN2(n14256), .QN(n14255) );
  INVX0 U14772 ( .INP(n14257), .ZN(n14254) );
  NOR2X0 U14773 ( .IN1(n14256), .IN2(n7800), .QN(n14257) );
  NOR2X0 U14774 ( .IN1(n14258), .IN2(n14259), .QN(n14256) );
  NOR2X0 U14775 ( .IN1(WX3449), .IN2(n7801), .QN(n14259) );
  INVX0 U14776 ( .INP(n14260), .ZN(n14258) );
  NAND2X0 U14777 ( .IN1(n7801), .IN2(WX3449), .QN(n14260) );
  NAND2X0 U14778 ( .IN1(n9790), .IN2(n8598), .QN(n14252) );
  NAND2X0 U14779 ( .IN1(n16055), .IN2(n9791), .QN(n14251) );
  NAND2X0 U14780 ( .IN1(n11504), .IN2(n9110), .QN(n14245) );
  NOR2X0 U14781 ( .IN1(n14261), .IN2(n14262), .QN(n11504) );
  INVX0 U14782 ( .INP(n14263), .ZN(n14262) );
  NAND2X0 U14783 ( .IN1(n14264), .IN2(n14265), .QN(n14263) );
  NOR2X0 U14784 ( .IN1(n14265), .IN2(n14264), .QN(n14261) );
  NAND2X0 U14785 ( .IN1(n14266), .IN2(n14267), .QN(n14264) );
  NAND2X0 U14786 ( .IN1(n8596), .IN2(n14268), .QN(n14267) );
  INVX0 U14787 ( .INP(n14269), .ZN(n14268) );
  NAND2X0 U14788 ( .IN1(n14269), .IN2(WX2156), .QN(n14266) );
  NAND2X0 U14789 ( .IN1(n14270), .IN2(n14271), .QN(n14269) );
  INVX0 U14790 ( .INP(n14272), .ZN(n14271) );
  NOR2X0 U14791 ( .IN1(n8814), .IN2(n16039), .QN(n14272) );
  NAND2X0 U14792 ( .IN1(n16039), .IN2(n8814), .QN(n14270) );
  NOR2X0 U14793 ( .IN1(n14273), .IN2(n14274), .QN(n14265) );
  INVX0 U14794 ( .INP(n14275), .ZN(n14274) );
  NAND2X0 U14795 ( .IN1(n7828), .IN2(n9121), .QN(n14275) );
  NOR2X0 U14796 ( .IN1(n9116), .IN2(n7828), .QN(n14273) );
  NAND2X0 U14797 ( .IN1(n262), .IN2(n9285), .QN(n14244) );
  NOR2X0 U14798 ( .IN1(n9226), .IN2(n9019), .QN(n262) );
  NAND2X0 U14799 ( .IN1(n9299), .IN2(CRC_OUT_8_18), .QN(n14243) );
  NAND4X0 U14800 ( .IN1(n14276), .IN2(n14277), .IN3(n14278), .IN4(n14279), 
        .QN(WX1961) );
  NAND2X0 U14801 ( .IN1(n14280), .IN2(n13436), .QN(n14279) );
  NAND2X0 U14802 ( .IN1(n14281), .IN2(n13439), .QN(n13436) );
  NAND2X0 U14803 ( .IN1(n14282), .IN2(n14283), .QN(n14281) );
  NAND2X0 U14804 ( .IN1(n16054), .IN2(n9121), .QN(n14283) );
  NAND2X0 U14805 ( .IN1(TM1), .IN2(n8599), .QN(n14282) );
  NAND3X0 U14806 ( .IN1(n14284), .IN2(n14285), .IN3(n14286), .QN(n14280) );
  NAND2X0 U14807 ( .IN1(n9327), .IN2(n13439), .QN(n14286) );
  NAND2X0 U14808 ( .IN1(n14287), .IN2(n14288), .QN(n13439) );
  NAND2X0 U14809 ( .IN1(n7802), .IN2(n14289), .QN(n14288) );
  INVX0 U14810 ( .INP(n14290), .ZN(n14287) );
  NOR2X0 U14811 ( .IN1(n14289), .IN2(n7802), .QN(n14290) );
  NOR2X0 U14812 ( .IN1(n14291), .IN2(n14292), .QN(n14289) );
  NOR2X0 U14813 ( .IN1(WX3447), .IN2(n7803), .QN(n14292) );
  INVX0 U14814 ( .INP(n14293), .ZN(n14291) );
  NAND2X0 U14815 ( .IN1(n7803), .IN2(WX3447), .QN(n14293) );
  NAND2X0 U14816 ( .IN1(n9083), .IN2(n8599), .QN(n14285) );
  NAND2X0 U14817 ( .IN1(n16054), .IN2(n9079), .QN(n14284) );
  NAND2X0 U14818 ( .IN1(n14294), .IN2(n11511), .QN(n14278) );
  NAND2X0 U14819 ( .IN1(n14295), .IN2(n11515), .QN(n11511) );
  NAND2X0 U14820 ( .IN1(n14296), .IN2(n14297), .QN(n14295) );
  NAND2X0 U14821 ( .IN1(n16038), .IN2(n9121), .QN(n14297) );
  NAND2X0 U14822 ( .IN1(TM1), .IN2(n8656), .QN(n14296) );
  NAND2X0 U14823 ( .IN1(n14298), .IN2(n14299), .QN(n14294) );
  NAND2X0 U14824 ( .IN1(n9103), .IN2(n11515), .QN(n14299) );
  NAND2X0 U14825 ( .IN1(n14300), .IN2(n14301), .QN(n11515) );
  NAND2X0 U14826 ( .IN1(n7829), .IN2(n14302), .QN(n14301) );
  INVX0 U14827 ( .INP(n14303), .ZN(n14300) );
  NOR2X0 U14828 ( .IN1(n14302), .IN2(n7829), .QN(n14303) );
  NOR2X0 U14829 ( .IN1(n14304), .IN2(n14305), .QN(n14302) );
  NOR2X0 U14830 ( .IN1(WX2154), .IN2(n7830), .QN(n14305) );
  INVX0 U14831 ( .INP(n14306), .ZN(n14304) );
  NAND2X0 U14832 ( .IN1(n7830), .IN2(WX2154), .QN(n14306) );
  NAND2X0 U14833 ( .IN1(n9103), .IN2(n8656), .QN(n14298) );
  NAND2X0 U14834 ( .IN1(n261), .IN2(n9285), .QN(n14277) );
  NOR2X0 U14835 ( .IN1(n9226), .IN2(n9020), .QN(n261) );
  NAND2X0 U14836 ( .IN1(n9299), .IN2(CRC_OUT_8_19), .QN(n14276) );
  NAND4X0 U14837 ( .IN1(n14307), .IN2(n14308), .IN3(n14309), .IN4(n14310), 
        .QN(WX1959) );
  NAND2X0 U14838 ( .IN1(n14311), .IN2(n13459), .QN(n14310) );
  NAND2X0 U14839 ( .IN1(n14312), .IN2(n13462), .QN(n13459) );
  NAND2X0 U14840 ( .IN1(n14313), .IN2(n14314), .QN(n14312) );
  NAND2X0 U14841 ( .IN1(n16053), .IN2(n9121), .QN(n14314) );
  NAND2X0 U14842 ( .IN1(TM1), .IN2(n8600), .QN(n14313) );
  NAND3X0 U14843 ( .IN1(n14315), .IN2(n14316), .IN3(n14317), .QN(n14311) );
  NAND2X0 U14844 ( .IN1(n9327), .IN2(n13462), .QN(n14317) );
  NAND2X0 U14845 ( .IN1(n14318), .IN2(n14319), .QN(n13462) );
  NAND2X0 U14846 ( .IN1(n7804), .IN2(n14320), .QN(n14319) );
  INVX0 U14847 ( .INP(n14321), .ZN(n14318) );
  NOR2X0 U14848 ( .IN1(n14320), .IN2(n7804), .QN(n14321) );
  NOR2X0 U14849 ( .IN1(n14322), .IN2(n14323), .QN(n14320) );
  NOR2X0 U14850 ( .IN1(WX3445), .IN2(n7805), .QN(n14323) );
  INVX0 U14851 ( .INP(n14324), .ZN(n14322) );
  NAND2X0 U14852 ( .IN1(n7805), .IN2(WX3445), .QN(n14324) );
  NAND2X0 U14853 ( .IN1(n9082), .IN2(n8600), .QN(n14316) );
  NAND2X0 U14854 ( .IN1(n16053), .IN2(n9078), .QN(n14315) );
  NAND2X0 U14855 ( .IN1(n14325), .IN2(n11522), .QN(n14309) );
  NAND2X0 U14856 ( .IN1(n14326), .IN2(n11526), .QN(n11522) );
  NAND2X0 U14857 ( .IN1(n14327), .IN2(n14328), .QN(n14326) );
  NAND2X0 U14858 ( .IN1(n16037), .IN2(n9121), .QN(n14328) );
  NAND2X0 U14859 ( .IN1(TM1), .IN2(n8657), .QN(n14327) );
  NAND2X0 U14860 ( .IN1(n14329), .IN2(n14330), .QN(n14325) );
  NAND2X0 U14861 ( .IN1(n9103), .IN2(n11526), .QN(n14330) );
  NAND2X0 U14862 ( .IN1(n14331), .IN2(n14332), .QN(n11526) );
  NAND2X0 U14863 ( .IN1(n7831), .IN2(n14333), .QN(n14332) );
  INVX0 U14864 ( .INP(n14334), .ZN(n14331) );
  NOR2X0 U14865 ( .IN1(n14333), .IN2(n7831), .QN(n14334) );
  NOR2X0 U14866 ( .IN1(n14335), .IN2(n14336), .QN(n14333) );
  NOR2X0 U14867 ( .IN1(WX2152), .IN2(n7832), .QN(n14336) );
  INVX0 U14868 ( .INP(n14337), .ZN(n14335) );
  NAND2X0 U14869 ( .IN1(n7832), .IN2(WX2152), .QN(n14337) );
  NAND2X0 U14870 ( .IN1(n9103), .IN2(n8657), .QN(n14329) );
  NAND2X0 U14871 ( .IN1(n260), .IN2(n9286), .QN(n14308) );
  NOR2X0 U14872 ( .IN1(n9226), .IN2(n9021), .QN(n260) );
  NAND2X0 U14873 ( .IN1(n9299), .IN2(CRC_OUT_8_20), .QN(n14307) );
  NAND4X0 U14874 ( .IN1(n14338), .IN2(n14339), .IN3(n14340), .IN4(n14341), 
        .QN(WX1957) );
  NAND2X0 U14875 ( .IN1(n14342), .IN2(n13482), .QN(n14341) );
  NAND2X0 U14876 ( .IN1(n14343), .IN2(n13485), .QN(n13482) );
  NAND2X0 U14877 ( .IN1(n14344), .IN2(n14345), .QN(n14343) );
  NAND2X0 U14878 ( .IN1(n16052), .IN2(n9121), .QN(n14345) );
  NAND2X0 U14879 ( .IN1(TM1), .IN2(n8601), .QN(n14344) );
  NAND3X0 U14880 ( .IN1(n14346), .IN2(n14347), .IN3(n14348), .QN(n14342) );
  NAND2X0 U14881 ( .IN1(n9327), .IN2(n13485), .QN(n14348) );
  NAND2X0 U14882 ( .IN1(n14349), .IN2(n14350), .QN(n13485) );
  NAND2X0 U14883 ( .IN1(n7806), .IN2(n14351), .QN(n14350) );
  INVX0 U14884 ( .INP(n14352), .ZN(n14349) );
  NOR2X0 U14885 ( .IN1(n14351), .IN2(n7806), .QN(n14352) );
  NOR2X0 U14886 ( .IN1(n14353), .IN2(n14354), .QN(n14351) );
  NOR2X0 U14887 ( .IN1(WX3443), .IN2(n7807), .QN(n14354) );
  INVX0 U14888 ( .INP(n14355), .ZN(n14353) );
  NAND2X0 U14889 ( .IN1(n7807), .IN2(WX3443), .QN(n14355) );
  NAND2X0 U14890 ( .IN1(n9081), .IN2(n8601), .QN(n14347) );
  NAND2X0 U14891 ( .IN1(n16052), .IN2(n9077), .QN(n14346) );
  NAND2X0 U14892 ( .IN1(n14356), .IN2(n11534), .QN(n14340) );
  NAND2X0 U14893 ( .IN1(n14357), .IN2(n11538), .QN(n11534) );
  NAND2X0 U14894 ( .IN1(n14358), .IN2(n14359), .QN(n14357) );
  NAND2X0 U14895 ( .IN1(n16036), .IN2(n9121), .QN(n14359) );
  NAND2X0 U14896 ( .IN1(TM1), .IN2(n8658), .QN(n14358) );
  NAND2X0 U14897 ( .IN1(n14360), .IN2(n14361), .QN(n14356) );
  NAND2X0 U14898 ( .IN1(n9103), .IN2(n11538), .QN(n14361) );
  NAND2X0 U14899 ( .IN1(n14362), .IN2(n14363), .QN(n11538) );
  NAND2X0 U14900 ( .IN1(n7833), .IN2(n14364), .QN(n14363) );
  INVX0 U14901 ( .INP(n14365), .ZN(n14362) );
  NOR2X0 U14902 ( .IN1(n14364), .IN2(n7833), .QN(n14365) );
  NOR2X0 U14903 ( .IN1(n14366), .IN2(n14367), .QN(n14364) );
  NOR2X0 U14904 ( .IN1(WX2150), .IN2(n7834), .QN(n14367) );
  INVX0 U14905 ( .INP(n14368), .ZN(n14366) );
  NAND2X0 U14906 ( .IN1(n7834), .IN2(WX2150), .QN(n14368) );
  NAND2X0 U14907 ( .IN1(n9103), .IN2(n8658), .QN(n14360) );
  NAND2X0 U14908 ( .IN1(n259), .IN2(n9286), .QN(n14339) );
  NOR2X0 U14909 ( .IN1(n9226), .IN2(n9022), .QN(n259) );
  NAND2X0 U14910 ( .IN1(n9299), .IN2(CRC_OUT_8_21), .QN(n14338) );
  NAND4X0 U14911 ( .IN1(n14369), .IN2(n14370), .IN3(n14371), .IN4(n14372), 
        .QN(WX1955) );
  NAND2X0 U14912 ( .IN1(n14373), .IN2(n13505), .QN(n14372) );
  NAND2X0 U14913 ( .IN1(n14374), .IN2(n13508), .QN(n13505) );
  NAND2X0 U14914 ( .IN1(n14375), .IN2(n14376), .QN(n14374) );
  NAND2X0 U14915 ( .IN1(n16051), .IN2(n9121), .QN(n14376) );
  NAND2X0 U14916 ( .IN1(TM1), .IN2(n8602), .QN(n14375) );
  NAND3X0 U14917 ( .IN1(n14377), .IN2(n14378), .IN3(n14379), .QN(n14373) );
  NAND2X0 U14918 ( .IN1(n9327), .IN2(n13508), .QN(n14379) );
  NAND2X0 U14919 ( .IN1(n14380), .IN2(n14381), .QN(n13508) );
  NAND2X0 U14920 ( .IN1(n7808), .IN2(n14382), .QN(n14381) );
  INVX0 U14921 ( .INP(n14383), .ZN(n14380) );
  NOR2X0 U14922 ( .IN1(n14382), .IN2(n7808), .QN(n14383) );
  NOR2X0 U14923 ( .IN1(n14384), .IN2(n14385), .QN(n14382) );
  NOR2X0 U14924 ( .IN1(WX3441), .IN2(n7809), .QN(n14385) );
  INVX0 U14925 ( .INP(n14386), .ZN(n14384) );
  NAND2X0 U14926 ( .IN1(n7809), .IN2(WX3441), .QN(n14386) );
  NAND2X0 U14927 ( .IN1(n9790), .IN2(n8602), .QN(n14378) );
  NAND2X0 U14928 ( .IN1(n16051), .IN2(n9791), .QN(n14377) );
  NAND2X0 U14929 ( .IN1(n14387), .IN2(n11545), .QN(n14371) );
  NAND3X0 U14930 ( .IN1(n14388), .IN2(n14389), .IN3(n11549), .QN(n11545) );
  NAND2X0 U14931 ( .IN1(n8592), .IN2(n9121), .QN(n14389) );
  NAND2X0 U14932 ( .IN1(TM1), .IN2(WX2148), .QN(n14388) );
  NAND2X0 U14933 ( .IN1(n14390), .IN2(n14391), .QN(n14387) );
  NAND2X0 U14934 ( .IN1(n9103), .IN2(n11549), .QN(n14391) );
  NAND2X0 U14935 ( .IN1(n14392), .IN2(n14393), .QN(n11549) );
  NAND2X0 U14936 ( .IN1(n14394), .IN2(WX2084), .QN(n14393) );
  NAND2X0 U14937 ( .IN1(n14395), .IN2(n14396), .QN(n14394) );
  NAND3X0 U14938 ( .IN1(n14395), .IN2(n14396), .IN3(n7836), .QN(n14392) );
  NAND2X0 U14939 ( .IN1(test_so13), .IN2(WX2020), .QN(n14396) );
  NAND2X0 U14940 ( .IN1(n7835), .IN2(n8824), .QN(n14395) );
  NAND2X0 U14941 ( .IN1(n8592), .IN2(n9109), .QN(n14390) );
  NAND2X0 U14942 ( .IN1(n258), .IN2(n9286), .QN(n14370) );
  NOR2X0 U14943 ( .IN1(n9226), .IN2(n9023), .QN(n258) );
  NAND2X0 U14944 ( .IN1(n9299), .IN2(CRC_OUT_8_22), .QN(n14369) );
  NAND4X0 U14945 ( .IN1(n14397), .IN2(n14398), .IN3(n14399), .IN4(n14400), 
        .QN(WX1953) );
  NAND2X0 U14946 ( .IN1(n14401), .IN2(n11556), .QN(n14400) );
  NAND2X0 U14947 ( .IN1(n14402), .IN2(n11560), .QN(n11556) );
  NAND2X0 U14948 ( .IN1(n14403), .IN2(n14404), .QN(n14402) );
  NAND2X0 U14949 ( .IN1(n16035), .IN2(n9121), .QN(n14404) );
  NAND2X0 U14950 ( .IN1(TM1), .IN2(n8661), .QN(n14403) );
  NAND2X0 U14951 ( .IN1(n14405), .IN2(n14406), .QN(n14401) );
  NAND2X0 U14952 ( .IN1(n9103), .IN2(n11560), .QN(n14406) );
  NAND2X0 U14953 ( .IN1(n14407), .IN2(n14408), .QN(n11560) );
  NAND2X0 U14954 ( .IN1(n7837), .IN2(n14409), .QN(n14408) );
  INVX0 U14955 ( .INP(n14410), .ZN(n14407) );
  NOR2X0 U14956 ( .IN1(n14409), .IN2(n7837), .QN(n14410) );
  NOR2X0 U14957 ( .IN1(n14411), .IN2(n14412), .QN(n14409) );
  NOR2X0 U14958 ( .IN1(WX2146), .IN2(n7838), .QN(n14412) );
  INVX0 U14959 ( .INP(n14413), .ZN(n14411) );
  NAND2X0 U14960 ( .IN1(n7838), .IN2(WX2146), .QN(n14413) );
  NAND2X0 U14961 ( .IN1(n9103), .IN2(n8661), .QN(n14405) );
  NAND2X0 U14962 ( .IN1(n13527), .IN2(n9335), .QN(n14399) );
  NOR2X0 U14963 ( .IN1(n14414), .IN2(n14415), .QN(n13527) );
  INVX0 U14964 ( .INP(n14416), .ZN(n14415) );
  NAND2X0 U14965 ( .IN1(n14417), .IN2(n14418), .QN(n14416) );
  NOR2X0 U14966 ( .IN1(n14418), .IN2(n14417), .QN(n14414) );
  NAND2X0 U14967 ( .IN1(n14419), .IN2(n14420), .QN(n14417) );
  NAND2X0 U14968 ( .IN1(n14421), .IN2(WX3375), .QN(n14420) );
  NAND2X0 U14969 ( .IN1(n14422), .IN2(n14423), .QN(n14421) );
  NAND3X0 U14970 ( .IN1(n14422), .IN2(n14423), .IN3(n7811), .QN(n14419) );
  NAND2X0 U14971 ( .IN1(test_so29), .IN2(WX3311), .QN(n14423) );
  NAND2X0 U14972 ( .IN1(n7810), .IN2(n8801), .QN(n14422) );
  NOR2X0 U14973 ( .IN1(n14424), .IN2(n14425), .QN(n14418) );
  INVX0 U14974 ( .INP(n14426), .ZN(n14425) );
  NAND2X0 U14975 ( .IN1(n16050), .IN2(n9121), .QN(n14426) );
  NOR2X0 U14976 ( .IN1(n9117), .IN2(n16050), .QN(n14424) );
  NAND2X0 U14977 ( .IN1(n257), .IN2(n9286), .QN(n14398) );
  NOR2X0 U14978 ( .IN1(n9226), .IN2(n9024), .QN(n257) );
  NAND2X0 U14979 ( .IN1(n9299), .IN2(CRC_OUT_8_23), .QN(n14397) );
  NAND4X0 U14980 ( .IN1(n14427), .IN2(n14428), .IN3(n14429), .IN4(n14430), 
        .QN(WX1951) );
  NAND2X0 U14981 ( .IN1(n14431), .IN2(n13547), .QN(n14430) );
  NAND2X0 U14982 ( .IN1(n14432), .IN2(n13550), .QN(n13547) );
  NAND2X0 U14983 ( .IN1(n14433), .IN2(n14434), .QN(n14432) );
  NAND2X0 U14984 ( .IN1(n16049), .IN2(n9121), .QN(n14434) );
  NAND2X0 U14985 ( .IN1(TM1), .IN2(n8604), .QN(n14433) );
  NAND3X0 U14986 ( .IN1(n14435), .IN2(n14436), .IN3(n14437), .QN(n14431) );
  NAND2X0 U14987 ( .IN1(n9327), .IN2(n13550), .QN(n14437) );
  NAND2X0 U14988 ( .IN1(n14438), .IN2(n14439), .QN(n13550) );
  NAND2X0 U14989 ( .IN1(n7812), .IN2(n14440), .QN(n14439) );
  INVX0 U14990 ( .INP(n14441), .ZN(n14438) );
  NOR2X0 U14991 ( .IN1(n14440), .IN2(n7812), .QN(n14441) );
  NOR2X0 U14992 ( .IN1(n14442), .IN2(n14443), .QN(n14440) );
  NOR2X0 U14993 ( .IN1(WX3437), .IN2(n7813), .QN(n14443) );
  INVX0 U14994 ( .INP(n14444), .ZN(n14442) );
  NAND2X0 U14995 ( .IN1(n7813), .IN2(WX3437), .QN(n14444) );
  NAND2X0 U14996 ( .IN1(n9083), .IN2(n8604), .QN(n14436) );
  NAND2X0 U14997 ( .IN1(n16049), .IN2(n9079), .QN(n14435) );
  NAND2X0 U14998 ( .IN1(n14445), .IN2(n11567), .QN(n14429) );
  NAND2X0 U14999 ( .IN1(n14446), .IN2(n11571), .QN(n11567) );
  NAND2X0 U15000 ( .IN1(n14447), .IN2(n14448), .QN(n14446) );
  NAND2X0 U15001 ( .IN1(n16034), .IN2(n9121), .QN(n14448) );
  NAND2X0 U15002 ( .IN1(TM1), .IN2(n8662), .QN(n14447) );
  NAND2X0 U15003 ( .IN1(n14449), .IN2(n14450), .QN(n14445) );
  NAND2X0 U15004 ( .IN1(n9103), .IN2(n11571), .QN(n14450) );
  NAND2X0 U15005 ( .IN1(n14451), .IN2(n14452), .QN(n11571) );
  NAND2X0 U15006 ( .IN1(n7839), .IN2(n14453), .QN(n14452) );
  INVX0 U15007 ( .INP(n14454), .ZN(n14451) );
  NOR2X0 U15008 ( .IN1(n14453), .IN2(n7839), .QN(n14454) );
  NOR2X0 U15009 ( .IN1(n14455), .IN2(n14456), .QN(n14453) );
  NOR2X0 U15010 ( .IN1(WX2144), .IN2(n7840), .QN(n14456) );
  INVX0 U15011 ( .INP(n14457), .ZN(n14455) );
  NAND2X0 U15012 ( .IN1(n7840), .IN2(WX2144), .QN(n14457) );
  NAND2X0 U15013 ( .IN1(n9103), .IN2(n8662), .QN(n14449) );
  NAND2X0 U15014 ( .IN1(n256), .IN2(n9286), .QN(n14428) );
  NOR2X0 U15015 ( .IN1(n9226), .IN2(n9025), .QN(n256) );
  NAND2X0 U15016 ( .IN1(n9299), .IN2(CRC_OUT_8_24), .QN(n14427) );
  NAND4X0 U15017 ( .IN1(n14458), .IN2(n14459), .IN3(n14460), .IN4(n14461), 
        .QN(WX1949) );
  NAND2X0 U15018 ( .IN1(n14462), .IN2(n13570), .QN(n14461) );
  NAND2X0 U15019 ( .IN1(n14463), .IN2(n13573), .QN(n13570) );
  NAND2X0 U15020 ( .IN1(n14464), .IN2(n14465), .QN(n14463) );
  NAND2X0 U15021 ( .IN1(n16048), .IN2(n9121), .QN(n14465) );
  NAND2X0 U15022 ( .IN1(TM1), .IN2(n8605), .QN(n14464) );
  NAND3X0 U15023 ( .IN1(n14466), .IN2(n14467), .IN3(n14468), .QN(n14462) );
  NAND2X0 U15024 ( .IN1(n9327), .IN2(n13573), .QN(n14468) );
  NAND2X0 U15025 ( .IN1(n14469), .IN2(n14470), .QN(n13573) );
  NAND2X0 U15026 ( .IN1(n7814), .IN2(n14471), .QN(n14470) );
  INVX0 U15027 ( .INP(n14472), .ZN(n14469) );
  NOR2X0 U15028 ( .IN1(n14471), .IN2(n7814), .QN(n14472) );
  NOR2X0 U15029 ( .IN1(n14473), .IN2(n14474), .QN(n14471) );
  NOR2X0 U15030 ( .IN1(WX3435), .IN2(n7815), .QN(n14474) );
  INVX0 U15031 ( .INP(n14475), .ZN(n14473) );
  NAND2X0 U15032 ( .IN1(n7815), .IN2(WX3435), .QN(n14475) );
  NAND2X0 U15033 ( .IN1(n9082), .IN2(n8605), .QN(n14467) );
  NAND2X0 U15034 ( .IN1(n16048), .IN2(n9078), .QN(n14466) );
  NAND2X0 U15035 ( .IN1(n14476), .IN2(n11579), .QN(n14460) );
  NAND2X0 U15036 ( .IN1(n14477), .IN2(n11583), .QN(n11579) );
  NAND2X0 U15037 ( .IN1(n14478), .IN2(n14479), .QN(n14477) );
  NAND2X0 U15038 ( .IN1(n16033), .IN2(n9121), .QN(n14479) );
  NAND2X0 U15039 ( .IN1(TM1), .IN2(n8663), .QN(n14478) );
  NAND2X0 U15040 ( .IN1(n14480), .IN2(n14481), .QN(n14476) );
  NAND2X0 U15041 ( .IN1(n9103), .IN2(n11583), .QN(n14481) );
  NAND2X0 U15042 ( .IN1(n14482), .IN2(n14483), .QN(n11583) );
  NAND2X0 U15043 ( .IN1(n7841), .IN2(n14484), .QN(n14483) );
  INVX0 U15044 ( .INP(n14485), .ZN(n14482) );
  NOR2X0 U15045 ( .IN1(n14484), .IN2(n7841), .QN(n14485) );
  NOR2X0 U15046 ( .IN1(n14486), .IN2(n14487), .QN(n14484) );
  NOR2X0 U15047 ( .IN1(WX2142), .IN2(n7842), .QN(n14487) );
  INVX0 U15048 ( .INP(n14488), .ZN(n14486) );
  NAND2X0 U15049 ( .IN1(n7842), .IN2(WX2142), .QN(n14488) );
  NAND2X0 U15050 ( .IN1(n9103), .IN2(n8663), .QN(n14480) );
  NAND2X0 U15051 ( .IN1(n255), .IN2(n9286), .QN(n14459) );
  NOR2X0 U15052 ( .IN1(n9225), .IN2(n9026), .QN(n255) );
  NAND2X0 U15053 ( .IN1(test_so21), .IN2(n9314), .QN(n14458) );
  NAND4X0 U15054 ( .IN1(n14489), .IN2(n14490), .IN3(n14491), .IN4(n14492), 
        .QN(WX1947) );
  NAND2X0 U15055 ( .IN1(n14493), .IN2(n11590), .QN(n14492) );
  NAND2X0 U15056 ( .IN1(n14494), .IN2(n11594), .QN(n11590) );
  NAND2X0 U15057 ( .IN1(n14495), .IN2(n14496), .QN(n14494) );
  NAND2X0 U15058 ( .IN1(n16032), .IN2(n9121), .QN(n14496) );
  NAND2X0 U15059 ( .IN1(TM1), .IN2(n8664), .QN(n14495) );
  NAND2X0 U15060 ( .IN1(n14497), .IN2(n14498), .QN(n14493) );
  NAND2X0 U15061 ( .IN1(n9103), .IN2(n11594), .QN(n14498) );
  NAND2X0 U15062 ( .IN1(n14499), .IN2(n14500), .QN(n11594) );
  NAND2X0 U15063 ( .IN1(n7843), .IN2(n14501), .QN(n14500) );
  INVX0 U15064 ( .INP(n14502), .ZN(n14499) );
  NOR2X0 U15065 ( .IN1(n14501), .IN2(n7843), .QN(n14502) );
  NOR2X0 U15066 ( .IN1(n14503), .IN2(n14504), .QN(n14501) );
  NOR2X0 U15067 ( .IN1(WX2140), .IN2(n7844), .QN(n14504) );
  INVX0 U15068 ( .INP(n14505), .ZN(n14503) );
  NAND2X0 U15069 ( .IN1(n7844), .IN2(WX2140), .QN(n14505) );
  NAND2X0 U15070 ( .IN1(n9102), .IN2(n8664), .QN(n14497) );
  NAND2X0 U15071 ( .IN1(n13592), .IN2(n9335), .QN(n14491) );
  NOR2X0 U15072 ( .IN1(n14506), .IN2(n14507), .QN(n13592) );
  INVX0 U15073 ( .INP(n14508), .ZN(n14507) );
  NAND2X0 U15074 ( .IN1(n14509), .IN2(n14510), .QN(n14508) );
  NOR2X0 U15075 ( .IN1(n14510), .IN2(n14509), .QN(n14506) );
  NAND2X0 U15076 ( .IN1(n14511), .IN2(n14512), .QN(n14509) );
  NAND2X0 U15077 ( .IN1(n8475), .IN2(n14513), .QN(n14512) );
  INVX0 U15078 ( .INP(n14514), .ZN(n14513) );
  NAND2X0 U15079 ( .IN1(n14514), .IN2(WX3433), .QN(n14511) );
  NAND2X0 U15080 ( .IN1(n14515), .IN2(n14516), .QN(n14514) );
  INVX0 U15081 ( .INP(n14517), .ZN(n14516) );
  NOR2X0 U15082 ( .IN1(n8815), .IN2(n16047), .QN(n14517) );
  NAND2X0 U15083 ( .IN1(n16047), .IN2(n8815), .QN(n14515) );
  NOR2X0 U15084 ( .IN1(n14518), .IN2(n14519), .QN(n14510) );
  INVX0 U15085 ( .INP(n14520), .ZN(n14519) );
  NAND2X0 U15086 ( .IN1(n7816), .IN2(n9121), .QN(n14520) );
  NOR2X0 U15087 ( .IN1(n9117), .IN2(n7816), .QN(n14518) );
  NAND2X0 U15088 ( .IN1(n254), .IN2(n9286), .QN(n14490) );
  NOR2X0 U15089 ( .IN1(n9073), .IN2(n9162), .QN(n254) );
  NAND2X0 U15090 ( .IN1(n9299), .IN2(CRC_OUT_8_26), .QN(n14489) );
  NAND4X0 U15091 ( .IN1(n14521), .IN2(n14522), .IN3(n14523), .IN4(n14524), 
        .QN(WX1945) );
  NAND2X0 U15092 ( .IN1(n14525), .IN2(n13612), .QN(n14524) );
  NAND2X0 U15093 ( .IN1(n14526), .IN2(n13615), .QN(n13612) );
  NAND2X0 U15094 ( .IN1(n14527), .IN2(n14528), .QN(n14526) );
  NAND2X0 U15095 ( .IN1(n16046), .IN2(n9121), .QN(n14528) );
  NAND2X0 U15096 ( .IN1(TM1), .IN2(n8607), .QN(n14527) );
  NAND3X0 U15097 ( .IN1(n14529), .IN2(n14530), .IN3(n14531), .QN(n14525) );
  NAND2X0 U15098 ( .IN1(n9327), .IN2(n13615), .QN(n14531) );
  NAND2X0 U15099 ( .IN1(n14532), .IN2(n14533), .QN(n13615) );
  NAND2X0 U15100 ( .IN1(n7817), .IN2(n14534), .QN(n14533) );
  INVX0 U15101 ( .INP(n14535), .ZN(n14532) );
  NOR2X0 U15102 ( .IN1(n14534), .IN2(n7817), .QN(n14535) );
  NOR2X0 U15103 ( .IN1(n14536), .IN2(n14537), .QN(n14534) );
  NOR2X0 U15104 ( .IN1(WX3431), .IN2(n7818), .QN(n14537) );
  INVX0 U15105 ( .INP(n14538), .ZN(n14536) );
  NAND2X0 U15106 ( .IN1(n7818), .IN2(WX3431), .QN(n14538) );
  NAND2X0 U15107 ( .IN1(n9081), .IN2(n8607), .QN(n14530) );
  NAND2X0 U15108 ( .IN1(n16046), .IN2(n9077), .QN(n14529) );
  NAND2X0 U15109 ( .IN1(n14539), .IN2(n11601), .QN(n14523) );
  NAND2X0 U15110 ( .IN1(n14540), .IN2(n11605), .QN(n11601) );
  NAND2X0 U15111 ( .IN1(n14541), .IN2(n14542), .QN(n14540) );
  NAND2X0 U15112 ( .IN1(n16031), .IN2(n9121), .QN(n14542) );
  NAND2X0 U15113 ( .IN1(TM1), .IN2(n8665), .QN(n14541) );
  NAND2X0 U15114 ( .IN1(n14543), .IN2(n14544), .QN(n14539) );
  NAND2X0 U15115 ( .IN1(n9102), .IN2(n11605), .QN(n14544) );
  NAND2X0 U15116 ( .IN1(n14545), .IN2(n14546), .QN(n11605) );
  NAND2X0 U15117 ( .IN1(n7845), .IN2(n14547), .QN(n14546) );
  INVX0 U15118 ( .INP(n14548), .ZN(n14545) );
  NOR2X0 U15119 ( .IN1(n14547), .IN2(n7845), .QN(n14548) );
  NOR2X0 U15120 ( .IN1(n14549), .IN2(n14550), .QN(n14547) );
  NOR2X0 U15121 ( .IN1(WX2138), .IN2(n7846), .QN(n14550) );
  INVX0 U15122 ( .INP(n14551), .ZN(n14549) );
  NAND2X0 U15123 ( .IN1(n7846), .IN2(WX2138), .QN(n14551) );
  NAND2X0 U15124 ( .IN1(n9102), .IN2(n8665), .QN(n14543) );
  NAND2X0 U15125 ( .IN1(n253), .IN2(n9286), .QN(n14522) );
  NOR2X0 U15126 ( .IN1(n9225), .IN2(n9027), .QN(n253) );
  NAND2X0 U15127 ( .IN1(n9299), .IN2(CRC_OUT_8_27), .QN(n14521) );
  NAND4X0 U15128 ( .IN1(n14552), .IN2(n14553), .IN3(n14554), .IN4(n14555), 
        .QN(WX1943) );
  NAND2X0 U15129 ( .IN1(n14556), .IN2(n13621), .QN(n14555) );
  NAND2X0 U15130 ( .IN1(n14557), .IN2(n13624), .QN(n13621) );
  NAND2X0 U15131 ( .IN1(n14558), .IN2(n14559), .QN(n14557) );
  NAND2X0 U15132 ( .IN1(n16045), .IN2(n9121), .QN(n14559) );
  NAND2X0 U15133 ( .IN1(TM1), .IN2(n8608), .QN(n14558) );
  NAND3X0 U15134 ( .IN1(n14560), .IN2(n14561), .IN3(n14562), .QN(n14556) );
  NAND2X0 U15135 ( .IN1(n9327), .IN2(n13624), .QN(n14562) );
  NAND2X0 U15136 ( .IN1(n14563), .IN2(n14564), .QN(n13624) );
  NAND2X0 U15137 ( .IN1(n7819), .IN2(n14565), .QN(n14564) );
  INVX0 U15138 ( .INP(n14566), .ZN(n14563) );
  NOR2X0 U15139 ( .IN1(n14565), .IN2(n7819), .QN(n14566) );
  NOR2X0 U15140 ( .IN1(n14567), .IN2(n14568), .QN(n14565) );
  NOR2X0 U15141 ( .IN1(WX3429), .IN2(n7820), .QN(n14568) );
  INVX0 U15142 ( .INP(n14569), .ZN(n14567) );
  NAND2X0 U15143 ( .IN1(n7820), .IN2(WX3429), .QN(n14569) );
  NAND2X0 U15144 ( .IN1(n9790), .IN2(n8608), .QN(n14561) );
  NAND2X0 U15145 ( .IN1(n16045), .IN2(n9791), .QN(n14560) );
  NAND2X0 U15146 ( .IN1(n11611), .IN2(n9110), .QN(n14554) );
  NOR2X0 U15147 ( .IN1(n14570), .IN2(n14571), .QN(n11611) );
  INVX0 U15148 ( .INP(n14572), .ZN(n14571) );
  NAND2X0 U15149 ( .IN1(n14573), .IN2(n14574), .QN(n14572) );
  NOR2X0 U15150 ( .IN1(n14574), .IN2(n14573), .QN(n14570) );
  NAND2X0 U15151 ( .IN1(n14575), .IN2(n14576), .QN(n14573) );
  NAND2X0 U15152 ( .IN1(n14577), .IN2(WX2072), .QN(n14576) );
  NAND2X0 U15153 ( .IN1(n14578), .IN2(n14579), .QN(n14577) );
  NAND3X0 U15154 ( .IN1(n14578), .IN2(n14579), .IN3(n7848), .QN(n14575) );
  NAND2X0 U15155 ( .IN1(test_so18), .IN2(WX2008), .QN(n14579) );
  NAND2X0 U15156 ( .IN1(n7847), .IN2(n8802), .QN(n14578) );
  NOR2X0 U15157 ( .IN1(n14580), .IN2(n14581), .QN(n14574) );
  INVX0 U15158 ( .INP(n14582), .ZN(n14581) );
  NAND2X0 U15159 ( .IN1(n16030), .IN2(n9122), .QN(n14582) );
  NOR2X0 U15160 ( .IN1(n9117), .IN2(n16030), .QN(n14580) );
  NAND2X0 U15161 ( .IN1(n252), .IN2(n9286), .QN(n14553) );
  NOR2X0 U15162 ( .IN1(n9225), .IN2(n9028), .QN(n252) );
  NAND2X0 U15163 ( .IN1(n9299), .IN2(CRC_OUT_8_28), .QN(n14552) );
  NAND4X0 U15164 ( .IN1(n14583), .IN2(n14584), .IN3(n14585), .IN4(n14586), 
        .QN(WX1941) );
  NAND2X0 U15165 ( .IN1(n14587), .IN2(n13657), .QN(n14586) );
  NAND2X0 U15166 ( .IN1(n14588), .IN2(n13660), .QN(n13657) );
  NAND2X0 U15167 ( .IN1(n14589), .IN2(n14590), .QN(n14588) );
  NAND2X0 U15168 ( .IN1(n16044), .IN2(n9122), .QN(n14590) );
  NAND2X0 U15169 ( .IN1(TM1), .IN2(n8609), .QN(n14589) );
  NAND3X0 U15170 ( .IN1(n14591), .IN2(n14592), .IN3(n14593), .QN(n14587) );
  NAND2X0 U15171 ( .IN1(n9327), .IN2(n13660), .QN(n14593) );
  NAND2X0 U15172 ( .IN1(n14594), .IN2(n14595), .QN(n13660) );
  NAND2X0 U15173 ( .IN1(n7821), .IN2(n14596), .QN(n14595) );
  INVX0 U15174 ( .INP(n14597), .ZN(n14594) );
  NOR2X0 U15175 ( .IN1(n14596), .IN2(n7821), .QN(n14597) );
  NOR2X0 U15176 ( .IN1(n14598), .IN2(n14599), .QN(n14596) );
  NOR2X0 U15177 ( .IN1(WX3427), .IN2(n7822), .QN(n14599) );
  INVX0 U15178 ( .INP(n14600), .ZN(n14598) );
  NAND2X0 U15179 ( .IN1(n7822), .IN2(WX3427), .QN(n14600) );
  NAND2X0 U15180 ( .IN1(n9083), .IN2(n8609), .QN(n14592) );
  NAND2X0 U15181 ( .IN1(n16044), .IN2(n9079), .QN(n14591) );
  NAND2X0 U15182 ( .IN1(n14601), .IN2(n11639), .QN(n14585) );
  NAND2X0 U15183 ( .IN1(n14602), .IN2(n11643), .QN(n11639) );
  NAND2X0 U15184 ( .IN1(n14603), .IN2(n14604), .QN(n14602) );
  NAND2X0 U15185 ( .IN1(n16029), .IN2(n9122), .QN(n14604) );
  NAND2X0 U15186 ( .IN1(TM1), .IN2(n8667), .QN(n14603) );
  NAND2X0 U15187 ( .IN1(n14605), .IN2(n14606), .QN(n14601) );
  NAND2X0 U15188 ( .IN1(n9102), .IN2(n11643), .QN(n14606) );
  NAND2X0 U15189 ( .IN1(n14607), .IN2(n14608), .QN(n11643) );
  NAND2X0 U15190 ( .IN1(n7849), .IN2(n14609), .QN(n14608) );
  INVX0 U15191 ( .INP(n14610), .ZN(n14607) );
  NOR2X0 U15192 ( .IN1(n14609), .IN2(n7849), .QN(n14610) );
  NOR2X0 U15193 ( .IN1(n14611), .IN2(n14612), .QN(n14609) );
  NOR2X0 U15194 ( .IN1(WX2134), .IN2(n7850), .QN(n14612) );
  INVX0 U15195 ( .INP(n14613), .ZN(n14611) );
  NAND2X0 U15196 ( .IN1(n7850), .IN2(WX2134), .QN(n14613) );
  NAND2X0 U15197 ( .IN1(n9102), .IN2(n8667), .QN(n14605) );
  NAND2X0 U15198 ( .IN1(n251), .IN2(n9286), .QN(n14584) );
  NOR2X0 U15199 ( .IN1(n9225), .IN2(n9029), .QN(n251) );
  NAND2X0 U15200 ( .IN1(n9299), .IN2(CRC_OUT_8_29), .QN(n14583) );
  NAND4X0 U15201 ( .IN1(n14614), .IN2(n14615), .IN3(n14616), .IN4(n14617), 
        .QN(WX1939) );
  NAND2X0 U15202 ( .IN1(n14618), .IN2(n11675), .QN(n14617) );
  NAND2X0 U15203 ( .IN1(n14619), .IN2(n11679), .QN(n11675) );
  NAND2X0 U15204 ( .IN1(n14620), .IN2(n14621), .QN(n14619) );
  NAND2X0 U15205 ( .IN1(n16028), .IN2(n9122), .QN(n14621) );
  NAND2X0 U15206 ( .IN1(TM1), .IN2(n8668), .QN(n14620) );
  NAND2X0 U15207 ( .IN1(n14622), .IN2(n14623), .QN(n14618) );
  NAND2X0 U15208 ( .IN1(n9102), .IN2(n11679), .QN(n14623) );
  NAND2X0 U15209 ( .IN1(n14624), .IN2(n14625), .QN(n11679) );
  NAND2X0 U15210 ( .IN1(n7851), .IN2(n14626), .QN(n14625) );
  INVX0 U15211 ( .INP(n14627), .ZN(n14624) );
  NOR2X0 U15212 ( .IN1(n14626), .IN2(n7851), .QN(n14627) );
  NOR2X0 U15213 ( .IN1(n14628), .IN2(n14629), .QN(n14626) );
  NOR2X0 U15214 ( .IN1(WX2132), .IN2(n7852), .QN(n14629) );
  INVX0 U15215 ( .INP(n14630), .ZN(n14628) );
  NAND2X0 U15216 ( .IN1(n7852), .IN2(WX2132), .QN(n14630) );
  NAND2X0 U15217 ( .IN1(n9102), .IN2(n8668), .QN(n14622) );
  NAND2X0 U15218 ( .IN1(n13680), .IN2(n9335), .QN(n14616) );
  NOR2X0 U15219 ( .IN1(n14631), .IN2(n14632), .QN(n13680) );
  INVX0 U15220 ( .INP(n14633), .ZN(n14632) );
  NAND2X0 U15221 ( .IN1(n14634), .IN2(n14635), .QN(n14633) );
  NOR2X0 U15222 ( .IN1(n14635), .IN2(n14634), .QN(n14631) );
  NAND2X0 U15223 ( .IN1(n14636), .IN2(n14637), .QN(n14634) );
  NAND2X0 U15224 ( .IN1(n8471), .IN2(n14638), .QN(n14637) );
  INVX0 U15225 ( .INP(n14639), .ZN(n14638) );
  NAND2X0 U15226 ( .IN1(n14639), .IN2(WX3425), .QN(n14636) );
  NAND2X0 U15227 ( .IN1(n14640), .IN2(n14641), .QN(n14639) );
  INVX0 U15228 ( .INP(n14642), .ZN(n14641) );
  NOR2X0 U15229 ( .IN1(n8816), .IN2(n16043), .QN(n14642) );
  NAND2X0 U15230 ( .IN1(n16043), .IN2(n8816), .QN(n14640) );
  NOR2X0 U15231 ( .IN1(n14643), .IN2(n14644), .QN(n14635) );
  INVX0 U15232 ( .INP(n14645), .ZN(n14644) );
  NAND2X0 U15233 ( .IN1(n7823), .IN2(n9122), .QN(n14645) );
  NOR2X0 U15234 ( .IN1(n9116), .IN2(n7823), .QN(n14643) );
  NAND2X0 U15235 ( .IN1(n250), .IN2(n9286), .QN(n14615) );
  NOR2X0 U15236 ( .IN1(n9225), .IN2(n9030), .QN(n250) );
  NAND2X0 U15237 ( .IN1(n9299), .IN2(CRC_OUT_8_30), .QN(n14614) );
  NAND4X0 U15238 ( .IN1(n14646), .IN2(n14647), .IN3(n14648), .IN4(n14649), 
        .QN(WX1937) );
  NAND2X0 U15239 ( .IN1(n14650), .IN2(n11716), .QN(n14649) );
  NAND2X0 U15240 ( .IN1(n14651), .IN2(n11720), .QN(n11716) );
  NAND2X0 U15241 ( .IN1(n14652), .IN2(n14653), .QN(n14651) );
  NAND2X0 U15242 ( .IN1(n16027), .IN2(n9122), .QN(n14653) );
  NAND2X0 U15243 ( .IN1(TM1), .IN2(n8669), .QN(n14652) );
  NAND2X0 U15244 ( .IN1(n14654), .IN2(n14655), .QN(n14650) );
  NAND2X0 U15245 ( .IN1(n9102), .IN2(n11720), .QN(n14655) );
  NAND2X0 U15246 ( .IN1(n14656), .IN2(n14657), .QN(n11720) );
  NAND2X0 U15247 ( .IN1(n7625), .IN2(n14658), .QN(n14657) );
  INVX0 U15248 ( .INP(n14659), .ZN(n14656) );
  NOR2X0 U15249 ( .IN1(n14658), .IN2(n7625), .QN(n14659) );
  NOR2X0 U15250 ( .IN1(n14660), .IN2(n14661), .QN(n14658) );
  NOR2X0 U15251 ( .IN1(WX2130), .IN2(n7626), .QN(n14661) );
  INVX0 U15252 ( .INP(n14662), .ZN(n14660) );
  NAND2X0 U15253 ( .IN1(n7626), .IN2(WX2130), .QN(n14662) );
  NAND2X0 U15254 ( .IN1(n9102), .IN2(n8669), .QN(n14654) );
  NAND2X0 U15255 ( .IN1(n14663), .IN2(n13700), .QN(n14648) );
  NAND2X0 U15256 ( .IN1(n14664), .IN2(n13703), .QN(n13700) );
  NAND2X0 U15257 ( .IN1(n14665), .IN2(n14666), .QN(n14664) );
  NAND2X0 U15258 ( .IN1(n16042), .IN2(n9122), .QN(n14666) );
  NAND2X0 U15259 ( .IN1(TM1), .IN2(n8611), .QN(n14665) );
  NAND3X0 U15260 ( .IN1(n14667), .IN2(n14668), .IN3(n14669), .QN(n14663) );
  NAND2X0 U15261 ( .IN1(n9327), .IN2(n13703), .QN(n14669) );
  NAND2X0 U15262 ( .IN1(n14670), .IN2(n14671), .QN(n13703) );
  NAND2X0 U15263 ( .IN1(n7623), .IN2(n14672), .QN(n14671) );
  INVX0 U15264 ( .INP(n14673), .ZN(n14670) );
  NOR2X0 U15265 ( .IN1(n14672), .IN2(n7623), .QN(n14673) );
  NOR2X0 U15266 ( .IN1(n14674), .IN2(n14675), .QN(n14672) );
  NOR2X0 U15267 ( .IN1(WX3423), .IN2(n7624), .QN(n14675) );
  INVX0 U15268 ( .INP(n14676), .ZN(n14674) );
  NAND2X0 U15269 ( .IN1(n7624), .IN2(WX3423), .QN(n14676) );
  NAND2X0 U15270 ( .IN1(n9082), .IN2(n8611), .QN(n14668) );
  NOR2X0 U15271 ( .IN1(n9336), .IN2(n9115), .QN(n9790) );
  NAND2X0 U15272 ( .IN1(n16042), .IN2(n9078), .QN(n14667) );
  NOR2X0 U15273 ( .IN1(n9336), .IN2(TM1), .QN(n9791) );
  NAND2X0 U15274 ( .IN1(n9300), .IN2(CRC_OUT_8_31), .QN(n14647) );
  NAND2X0 U15275 ( .IN1(n2245), .IN2(WX1778), .QN(n14646) );
  NOR2X0 U15276 ( .IN1(n9225), .IN2(WX1778), .QN(WX1839) );
  NOR3X0 U15277 ( .IN1(n9151), .IN2(n14677), .IN3(n14678), .QN(WX1326) );
  NOR2X0 U15278 ( .IN1(n8774), .IN2(CRC_OUT_9_30), .QN(n14678) );
  NOR2X0 U15279 ( .IN1(DFF_190_n1), .IN2(WX837), .QN(n14677) );
  NOR3X0 U15280 ( .IN1(n9150), .IN2(n14679), .IN3(n14680), .QN(WX1324) );
  NOR2X0 U15281 ( .IN1(n8679), .IN2(CRC_OUT_9_29), .QN(n14680) );
  NOR2X0 U15282 ( .IN1(DFF_189_n1), .IN2(WX839), .QN(n14679) );
  NOR3X0 U15283 ( .IN1(n9150), .IN2(n14681), .IN3(n14682), .QN(WX1322) );
  NOR2X0 U15284 ( .IN1(n8708), .IN2(CRC_OUT_9_28), .QN(n14682) );
  NOR2X0 U15285 ( .IN1(DFF_188_n1), .IN2(WX841), .QN(n14681) );
  NOR3X0 U15286 ( .IN1(n9150), .IN2(n14683), .IN3(n14684), .QN(WX1320) );
  NOR2X0 U15287 ( .IN1(n8717), .IN2(CRC_OUT_9_27), .QN(n14684) );
  NOR2X0 U15288 ( .IN1(DFF_187_n1), .IN2(WX843), .QN(n14683) );
  NOR3X0 U15289 ( .IN1(n9150), .IN2(n14685), .IN3(n14686), .QN(WX1318) );
  NOR2X0 U15290 ( .IN1(n8723), .IN2(CRC_OUT_9_26), .QN(n14686) );
  NOR2X0 U15291 ( .IN1(DFF_186_n1), .IN2(WX845), .QN(n14685) );
  NOR3X0 U15292 ( .IN1(n9150), .IN2(n14687), .IN3(n14688), .QN(WX1316) );
  NOR2X0 U15293 ( .IN1(n8726), .IN2(CRC_OUT_9_25), .QN(n14688) );
  NOR2X0 U15294 ( .IN1(DFF_185_n1), .IN2(WX847), .QN(n14687) );
  NOR3X0 U15295 ( .IN1(n9150), .IN2(n14689), .IN3(n14690), .QN(WX1314) );
  NOR2X0 U15296 ( .IN1(n8735), .IN2(CRC_OUT_9_24), .QN(n14690) );
  NOR2X0 U15297 ( .IN1(DFF_184_n1), .IN2(WX849), .QN(n14689) );
  NOR3X0 U15298 ( .IN1(n9150), .IN2(n14691), .IN3(n14692), .QN(WX1312) );
  NOR2X0 U15299 ( .IN1(n8744), .IN2(CRC_OUT_9_23), .QN(n14692) );
  NOR2X0 U15300 ( .IN1(DFF_183_n1), .IN2(WX851), .QN(n14691) );
  NOR3X0 U15301 ( .IN1(n9150), .IN2(n14693), .IN3(n14694), .QN(WX1310) );
  NOR2X0 U15302 ( .IN1(n8746), .IN2(CRC_OUT_9_22), .QN(n14694) );
  NOR2X0 U15303 ( .IN1(DFF_182_n1), .IN2(WX853), .QN(n14693) );
  NOR3X0 U15304 ( .IN1(n9150), .IN2(n14695), .IN3(n14696), .QN(WX1308) );
  NOR2X0 U15305 ( .IN1(n8761), .IN2(CRC_OUT_9_21), .QN(n14696) );
  NOR2X0 U15306 ( .IN1(DFF_181_n1), .IN2(WX855), .QN(n14695) );
  NOR3X0 U15307 ( .IN1(n9150), .IN2(n14697), .IN3(n14698), .QN(WX1306) );
  NOR2X0 U15308 ( .IN1(n8767), .IN2(CRC_OUT_9_20), .QN(n14698) );
  NOR2X0 U15309 ( .IN1(DFF_180_n1), .IN2(WX857), .QN(n14697) );
  NOR2X0 U15310 ( .IN1(n9225), .IN2(n14699), .QN(WX1304) );
  NOR2X0 U15311 ( .IN1(n14700), .IN2(n14701), .QN(n14699) );
  NOR2X0 U15312 ( .IN1(test_so10), .IN2(WX859), .QN(n14701) );
  INVX0 U15313 ( .INP(n14702), .ZN(n14700) );
  NAND2X0 U15314 ( .IN1(WX859), .IN2(test_so10), .QN(n14702) );
  NOR3X0 U15315 ( .IN1(n9150), .IN2(n14703), .IN3(n14704), .QN(WX1302) );
  NOR2X0 U15316 ( .IN1(n8705), .IN2(CRC_OUT_9_18), .QN(n14704) );
  NOR2X0 U15317 ( .IN1(DFF_178_n1), .IN2(WX861), .QN(n14703) );
  NOR3X0 U15318 ( .IN1(n9150), .IN2(n14705), .IN3(n14706), .QN(WX1300) );
  NOR2X0 U15319 ( .IN1(n8720), .IN2(CRC_OUT_9_17), .QN(n14706) );
  NOR2X0 U15320 ( .IN1(DFF_177_n1), .IN2(WX863), .QN(n14705) );
  NOR3X0 U15321 ( .IN1(n9149), .IN2(n14707), .IN3(n14708), .QN(WX1298) );
  NOR2X0 U15322 ( .IN1(n8732), .IN2(CRC_OUT_9_16), .QN(n14708) );
  NOR2X0 U15323 ( .IN1(DFF_176_n1), .IN2(WX865), .QN(n14707) );
  NOR3X0 U15324 ( .IN1(n9149), .IN2(n14709), .IN3(n14710), .QN(WX1296) );
  INVX0 U15325 ( .INP(n14711), .ZN(n14710) );
  NAND2X0 U15326 ( .IN1(CRC_OUT_9_15), .IN2(n14712), .QN(n14711) );
  NOR2X0 U15327 ( .IN1(n14712), .IN2(CRC_OUT_9_15), .QN(n14709) );
  NAND2X0 U15328 ( .IN1(n14713), .IN2(n14714), .QN(n14712) );
  NAND2X0 U15329 ( .IN1(test_so8), .IN2(CRC_OUT_9_31), .QN(n14714) );
  NAND2X0 U15330 ( .IN1(DFF_191_n1), .IN2(n8797), .QN(n14713) );
  NOR3X0 U15331 ( .IN1(n9149), .IN2(n14715), .IN3(n14716), .QN(WX1294) );
  NOR2X0 U15332 ( .IN1(n8764), .IN2(CRC_OUT_9_14), .QN(n14716) );
  NOR2X0 U15333 ( .IN1(DFF_174_n1), .IN2(WX869), .QN(n14715) );
  NOR3X0 U15334 ( .IN1(n9149), .IN2(n14717), .IN3(n14718), .QN(WX1292) );
  NOR2X0 U15335 ( .IN1(n8776), .IN2(CRC_OUT_9_13), .QN(n14718) );
  NOR2X0 U15336 ( .IN1(DFF_173_n1), .IN2(WX871), .QN(n14717) );
  NOR3X0 U15337 ( .IN1(n9149), .IN2(n14719), .IN3(n14720), .QN(WX1290) );
  NOR2X0 U15338 ( .IN1(n8711), .IN2(CRC_OUT_9_12), .QN(n14720) );
  NOR2X0 U15339 ( .IN1(DFF_172_n1), .IN2(WX873), .QN(n14719) );
  NOR3X0 U15340 ( .IN1(n9149), .IN2(n14721), .IN3(n14722), .QN(WX1288) );
  NOR2X0 U15341 ( .IN1(n8738), .IN2(CRC_OUT_9_11), .QN(n14722) );
  NOR2X0 U15342 ( .IN1(DFF_171_n1), .IN2(WX875), .QN(n14721) );
  NOR2X0 U15343 ( .IN1(n9225), .IN2(n14723), .QN(WX1286) );
  NOR2X0 U15344 ( .IN1(n14724), .IN2(n14725), .QN(n14723) );
  INVX0 U15345 ( .INP(n14726), .ZN(n14725) );
  NAND2X0 U15346 ( .IN1(CRC_OUT_9_10), .IN2(n14727), .QN(n14726) );
  NOR2X0 U15347 ( .IN1(n14727), .IN2(CRC_OUT_9_10), .QN(n14724) );
  NAND2X0 U15348 ( .IN1(n14728), .IN2(n14729), .QN(n14727) );
  NAND2X0 U15349 ( .IN1(n8784), .IN2(CRC_OUT_9_31), .QN(n14729) );
  NAND2X0 U15350 ( .IN1(DFF_191_n1), .IN2(WX877), .QN(n14728) );
  NOR3X0 U15351 ( .IN1(n9149), .IN2(n14730), .IN3(n14731), .QN(WX1284) );
  NOR2X0 U15352 ( .IN1(n8729), .IN2(CRC_OUT_9_9), .QN(n14731) );
  NOR2X0 U15353 ( .IN1(DFF_169_n1), .IN2(WX879), .QN(n14730) );
  NOR3X0 U15354 ( .IN1(n9149), .IN2(n14732), .IN3(n14733), .QN(WX1282) );
  NOR2X0 U15355 ( .IN1(n8742), .IN2(CRC_OUT_9_8), .QN(n14733) );
  NOR2X0 U15356 ( .IN1(DFF_168_n1), .IN2(WX881), .QN(n14732) );
  NOR3X0 U15357 ( .IN1(n9149), .IN2(n14734), .IN3(n14735), .QN(WX1280) );
  NOR2X0 U15358 ( .IN1(n8751), .IN2(CRC_OUT_9_7), .QN(n14735) );
  NOR2X0 U15359 ( .IN1(DFF_167_n1), .IN2(WX883), .QN(n14734) );
  NOR3X0 U15360 ( .IN1(n9149), .IN2(n14736), .IN3(n14737), .QN(WX1278) );
  NOR2X0 U15361 ( .IN1(n8782), .IN2(CRC_OUT_9_6), .QN(n14737) );
  NOR2X0 U15362 ( .IN1(DFF_166_n1), .IN2(WX885), .QN(n14736) );
  NOR3X0 U15363 ( .IN1(n9149), .IN2(n14738), .IN3(n14739), .QN(WX1276) );
  NOR2X0 U15364 ( .IN1(n8769), .IN2(CRC_OUT_9_5), .QN(n14739) );
  NOR2X0 U15365 ( .IN1(DFF_165_n1), .IN2(WX887), .QN(n14738) );
  NOR3X0 U15366 ( .IN1(n9149), .IN2(n14740), .IN3(n14741), .QN(WX1274) );
  NOR2X0 U15367 ( .IN1(n8754), .IN2(CRC_OUT_9_4), .QN(n14741) );
  NOR2X0 U15368 ( .IN1(DFF_164_n1), .IN2(WX889), .QN(n14740) );
  NOR2X0 U15369 ( .IN1(n9224), .IN2(n14742), .QN(WX1272) );
  NOR2X0 U15370 ( .IN1(n14743), .IN2(n14744), .QN(n14742) );
  INVX0 U15371 ( .INP(n14745), .ZN(n14744) );
  NAND2X0 U15372 ( .IN1(CRC_OUT_9_3), .IN2(n14746), .QN(n14745) );
  NOR2X0 U15373 ( .IN1(n14746), .IN2(CRC_OUT_9_3), .QN(n14743) );
  NAND2X0 U15374 ( .IN1(n14747), .IN2(n14748), .QN(n14746) );
  NAND2X0 U15375 ( .IN1(n8757), .IN2(CRC_OUT_9_31), .QN(n14748) );
  NAND2X0 U15376 ( .IN1(DFF_191_n1), .IN2(WX891), .QN(n14747) );
  NOR3X0 U15377 ( .IN1(n9148), .IN2(n14749), .IN3(n14750), .QN(WX1270) );
  NOR2X0 U15378 ( .IN1(n8698), .IN2(CRC_OUT_9_2), .QN(n14750) );
  NOR2X0 U15379 ( .IN1(DFF_162_n1), .IN2(WX893), .QN(n14749) );
  NOR2X0 U15380 ( .IN1(n9224), .IN2(n14751), .QN(WX1268) );
  NOR2X0 U15381 ( .IN1(n14752), .IN2(n14753), .QN(n14751) );
  NOR2X0 U15382 ( .IN1(test_so9), .IN2(WX895), .QN(n14753) );
  INVX0 U15383 ( .INP(n14754), .ZN(n14752) );
  NAND2X0 U15384 ( .IN1(WX895), .IN2(test_so9), .QN(n14754) );
  NOR3X0 U15385 ( .IN1(n9148), .IN2(n14755), .IN3(n14756), .QN(WX1266) );
  NOR2X0 U15386 ( .IN1(n8713), .IN2(CRC_OUT_9_0), .QN(n14756) );
  NOR2X0 U15387 ( .IN1(DFF_160_n1), .IN2(WX897), .QN(n14755) );
  NOR3X0 U15388 ( .IN1(n9148), .IN2(n14757), .IN3(n14758), .QN(WX1264) );
  NOR2X0 U15389 ( .IN1(n8788), .IN2(CRC_OUT_9_31), .QN(n14758) );
  NOR2X0 U15390 ( .IN1(DFF_191_n1), .IN2(WX899), .QN(n14757) );
  NOR3X0 U15391 ( .IN1(n9146), .IN2(n14759), .IN3(n14760), .QN(WX11670) );
  NOR2X0 U15392 ( .IN1(n8133), .IN2(CRC_OUT_1_30), .QN(n14760) );
  NOR2X0 U15393 ( .IN1(DFF_1726_n1), .IN2(WX11181), .QN(n14759) );
  NOR3X0 U15394 ( .IN1(n9148), .IN2(n14761), .IN3(n14762), .QN(WX11668) );
  NOR2X0 U15395 ( .IN1(n8134), .IN2(CRC_OUT_1_29), .QN(n14762) );
  NOR2X0 U15396 ( .IN1(DFF_1725_n1), .IN2(WX11183), .QN(n14761) );
  NOR3X0 U15397 ( .IN1(n9148), .IN2(n14763), .IN3(n14764), .QN(WX11666) );
  NOR2X0 U15398 ( .IN1(n8135), .IN2(CRC_OUT_1_28), .QN(n14764) );
  NOR2X0 U15399 ( .IN1(DFF_1724_n1), .IN2(WX11185), .QN(n14763) );
  NOR3X0 U15400 ( .IN1(n9148), .IN2(n14765), .IN3(n14766), .QN(WX11664) );
  NOR2X0 U15401 ( .IN1(n8136), .IN2(CRC_OUT_1_27), .QN(n14766) );
  NOR2X0 U15402 ( .IN1(DFF_1723_n1), .IN2(WX11187), .QN(n14765) );
  NOR3X0 U15403 ( .IN1(n9148), .IN2(n14767), .IN3(n14768), .QN(WX11662) );
  NOR2X0 U15404 ( .IN1(n8137), .IN2(CRC_OUT_1_26), .QN(n14768) );
  NOR2X0 U15405 ( .IN1(DFF_1722_n1), .IN2(WX11189), .QN(n14767) );
  NOR3X0 U15406 ( .IN1(n9148), .IN2(n14769), .IN3(n14770), .QN(WX11660) );
  NOR2X0 U15407 ( .IN1(n8138), .IN2(CRC_OUT_1_25), .QN(n14770) );
  NOR2X0 U15408 ( .IN1(DFF_1721_n1), .IN2(WX11191), .QN(n14769) );
  NOR3X0 U15409 ( .IN1(n9148), .IN2(n14771), .IN3(n14772), .QN(WX11658) );
  NOR2X0 U15410 ( .IN1(n8139), .IN2(CRC_OUT_1_24), .QN(n14772) );
  NOR2X0 U15411 ( .IN1(DFF_1720_n1), .IN2(WX11193), .QN(n14771) );
  NOR3X0 U15412 ( .IN1(n9148), .IN2(n14773), .IN3(n14774), .QN(WX11656) );
  NOR2X0 U15413 ( .IN1(n8140), .IN2(CRC_OUT_1_23), .QN(n14774) );
  NOR2X0 U15414 ( .IN1(DFF_1719_n1), .IN2(WX11195), .QN(n14773) );
  NOR3X0 U15415 ( .IN1(n9148), .IN2(n14775), .IN3(n14776), .QN(WX11654) );
  NOR2X0 U15416 ( .IN1(n8141), .IN2(CRC_OUT_1_22), .QN(n14776) );
  NOR2X0 U15417 ( .IN1(DFF_1718_n1), .IN2(WX11197), .QN(n14775) );
  NOR3X0 U15418 ( .IN1(n9148), .IN2(n14777), .IN3(n14778), .QN(WX11652) );
  NOR2X0 U15419 ( .IN1(n8142), .IN2(CRC_OUT_1_21), .QN(n14778) );
  NOR2X0 U15420 ( .IN1(DFF_1717_n1), .IN2(WX11199), .QN(n14777) );
  NOR3X0 U15421 ( .IN1(n9147), .IN2(n14779), .IN3(n14780), .QN(WX11650) );
  NOR2X0 U15422 ( .IN1(n8143), .IN2(CRC_OUT_1_20), .QN(n14780) );
  NOR2X0 U15423 ( .IN1(DFF_1716_n1), .IN2(WX11201), .QN(n14779) );
  NOR3X0 U15424 ( .IN1(n9147), .IN2(n14781), .IN3(n14782), .QN(WX11648) );
  NOR2X0 U15425 ( .IN1(n8144), .IN2(CRC_OUT_1_19), .QN(n14782) );
  NOR2X0 U15426 ( .IN1(DFF_1715_n1), .IN2(WX11203), .QN(n14781) );
  NOR2X0 U15427 ( .IN1(n9223), .IN2(n14783), .QN(WX11646) );
  NOR2X0 U15428 ( .IN1(n14784), .IN2(n14785), .QN(n14783) );
  NOR2X0 U15429 ( .IN1(test_so97), .IN2(CRC_OUT_1_18), .QN(n14785) );
  NOR2X0 U15430 ( .IN1(DFF_1714_n1), .IN2(n8803), .QN(n14784) );
  NOR3X0 U15431 ( .IN1(n9147), .IN2(n14786), .IN3(n14787), .QN(WX11644) );
  NOR2X0 U15432 ( .IN1(n8145), .IN2(CRC_OUT_1_17), .QN(n14787) );
  NOR2X0 U15433 ( .IN1(DFF_1713_n1), .IN2(WX11207), .QN(n14786) );
  NOR3X0 U15434 ( .IN1(n9147), .IN2(n14788), .IN3(n14789), .QN(WX11642) );
  NOR2X0 U15435 ( .IN1(n8146), .IN2(CRC_OUT_1_16), .QN(n14789) );
  NOR2X0 U15436 ( .IN1(DFF_1712_n1), .IN2(WX11209), .QN(n14788) );
  NOR3X0 U15437 ( .IN1(n9147), .IN2(n14790), .IN3(n14791), .QN(WX11640) );
  INVX0 U15438 ( .INP(n14792), .ZN(n14791) );
  NAND2X0 U15439 ( .IN1(CRC_OUT_1_15), .IN2(n14793), .QN(n14792) );
  NOR2X0 U15440 ( .IN1(n14793), .IN2(CRC_OUT_1_15), .QN(n14790) );
  NAND2X0 U15441 ( .IN1(n14794), .IN2(n14795), .QN(n14793) );
  NAND2X0 U15442 ( .IN1(test_so100), .IN2(WX11211), .QN(n14795) );
  NAND2X0 U15443 ( .IN1(n8104), .IN2(n8789), .QN(n14794) );
  NOR2X0 U15444 ( .IN1(n9226), .IN2(n14796), .QN(WX11638) );
  NOR2X0 U15445 ( .IN1(n14797), .IN2(n14798), .QN(n14796) );
  NOR2X0 U15446 ( .IN1(test_so99), .IN2(WX11213), .QN(n14798) );
  INVX0 U15447 ( .INP(n14799), .ZN(n14797) );
  NAND2X0 U15448 ( .IN1(WX11213), .IN2(test_so99), .QN(n14799) );
  NOR3X0 U15449 ( .IN1(n9147), .IN2(n14800), .IN3(n14801), .QN(WX11636) );
  NOR2X0 U15450 ( .IN1(n8148), .IN2(CRC_OUT_1_13), .QN(n14801) );
  NOR2X0 U15451 ( .IN1(DFF_1709_n1), .IN2(WX11215), .QN(n14800) );
  NOR3X0 U15452 ( .IN1(n9147), .IN2(n14802), .IN3(n14803), .QN(WX11634) );
  NOR2X0 U15453 ( .IN1(n8149), .IN2(CRC_OUT_1_12), .QN(n14803) );
  NOR2X0 U15454 ( .IN1(DFF_1708_n1), .IN2(WX11217), .QN(n14802) );
  NOR3X0 U15455 ( .IN1(n9147), .IN2(n14804), .IN3(n14805), .QN(WX11632) );
  NOR2X0 U15456 ( .IN1(n8150), .IN2(CRC_OUT_1_11), .QN(n14805) );
  NOR2X0 U15457 ( .IN1(DFF_1707_n1), .IN2(WX11219), .QN(n14804) );
  NOR3X0 U15458 ( .IN1(n9146), .IN2(n14806), .IN3(n14807), .QN(WX11630) );
  INVX0 U15459 ( .INP(n14808), .ZN(n14807) );
  NAND2X0 U15460 ( .IN1(CRC_OUT_1_10), .IN2(n14809), .QN(n14808) );
  NOR2X0 U15461 ( .IN1(n14809), .IN2(CRC_OUT_1_10), .QN(n14806) );
  NAND2X0 U15462 ( .IN1(n14810), .IN2(n14811), .QN(n14809) );
  NAND2X0 U15463 ( .IN1(test_so100), .IN2(WX11221), .QN(n14811) );
  NAND2X0 U15464 ( .IN1(n8105), .IN2(n8789), .QN(n14810) );
  NOR3X0 U15465 ( .IN1(n9146), .IN2(n14812), .IN3(n14813), .QN(WX11628) );
  NOR2X0 U15466 ( .IN1(n8151), .IN2(CRC_OUT_1_9), .QN(n14813) );
  NOR2X0 U15467 ( .IN1(DFF_1705_n1), .IN2(WX11223), .QN(n14812) );
  NOR3X0 U15468 ( .IN1(n9151), .IN2(n14814), .IN3(n14815), .QN(WX11626) );
  NOR2X0 U15469 ( .IN1(n8152), .IN2(CRC_OUT_1_8), .QN(n14815) );
  NOR2X0 U15470 ( .IN1(DFF_1704_n1), .IN2(WX11225), .QN(n14814) );
  NOR3X0 U15471 ( .IN1(n9146), .IN2(n14816), .IN3(n14817), .QN(WX11624) );
  NOR2X0 U15472 ( .IN1(n8153), .IN2(CRC_OUT_1_7), .QN(n14817) );
  NOR2X0 U15473 ( .IN1(DFF_1703_n1), .IN2(WX11227), .QN(n14816) );
  NOR3X0 U15474 ( .IN1(n9146), .IN2(n14818), .IN3(n14819), .QN(WX11622) );
  NOR2X0 U15475 ( .IN1(n8154), .IN2(CRC_OUT_1_6), .QN(n14819) );
  NOR2X0 U15476 ( .IN1(DFF_1702_n1), .IN2(WX11229), .QN(n14818) );
  NOR3X0 U15477 ( .IN1(n9146), .IN2(n14820), .IN3(n14821), .QN(WX11620) );
  NOR2X0 U15478 ( .IN1(n8155), .IN2(CRC_OUT_1_5), .QN(n14821) );
  NOR2X0 U15479 ( .IN1(DFF_1701_n1), .IN2(WX11231), .QN(n14820) );
  NOR3X0 U15480 ( .IN1(n9147), .IN2(n14822), .IN3(n14823), .QN(WX11618) );
  NOR2X0 U15481 ( .IN1(n8156), .IN2(CRC_OUT_1_4), .QN(n14823) );
  NOR2X0 U15482 ( .IN1(DFF_1700_n1), .IN2(WX11233), .QN(n14822) );
  NOR3X0 U15483 ( .IN1(n9147), .IN2(n14824), .IN3(n14825), .QN(WX11616) );
  INVX0 U15484 ( .INP(n14826), .ZN(n14825) );
  NAND2X0 U15485 ( .IN1(CRC_OUT_1_3), .IN2(n14827), .QN(n14826) );
  NOR2X0 U15486 ( .IN1(n14827), .IN2(CRC_OUT_1_3), .QN(n14824) );
  NAND2X0 U15487 ( .IN1(n14828), .IN2(n14829), .QN(n14827) );
  NAND2X0 U15488 ( .IN1(test_so100), .IN2(WX11235), .QN(n14829) );
  NAND2X0 U15489 ( .IN1(n8106), .IN2(n8789), .QN(n14828) );
  NOR3X0 U15490 ( .IN1(n9147), .IN2(n14830), .IN3(n14831), .QN(WX11614) );
  NOR2X0 U15491 ( .IN1(n8157), .IN2(CRC_OUT_1_2), .QN(n14831) );
  NOR2X0 U15492 ( .IN1(DFF_1698_n1), .IN2(WX11237), .QN(n14830) );
  NOR2X0 U15493 ( .IN1(n9227), .IN2(n14832), .QN(WX11612) );
  NOR2X0 U15494 ( .IN1(n14833), .IN2(n14834), .QN(n14832) );
  NOR2X0 U15495 ( .IN1(test_so98), .IN2(CRC_OUT_1_1), .QN(n14834) );
  NOR2X0 U15496 ( .IN1(DFF_1697_n1), .IN2(n8793), .QN(n14833) );
  NOR3X0 U15497 ( .IN1(n9147), .IN2(n14835), .IN3(n14836), .QN(WX11610) );
  NOR2X0 U15498 ( .IN1(n8158), .IN2(CRC_OUT_1_0), .QN(n14836) );
  NOR2X0 U15499 ( .IN1(DFF_1696_n1), .IN2(WX11241), .QN(n14835) );
  NOR2X0 U15500 ( .IN1(n9227), .IN2(n14837), .QN(WX11608) );
  NOR2X0 U15501 ( .IN1(n14838), .IN2(n14839), .QN(n14837) );
  NOR2X0 U15502 ( .IN1(test_so100), .IN2(WX11243), .QN(n14839) );
  NOR2X0 U15503 ( .IN1(n8125), .IN2(n8789), .QN(n14838) );
  NOR2X0 U15504 ( .IN1(n16147), .IN2(n9158), .QN(WX11082) );
  NOR2X0 U15505 ( .IN1(n16146), .IN2(n9158), .QN(WX11080) );
  NOR2X0 U15506 ( .IN1(n16145), .IN2(n9157), .QN(WX11078) );
  NOR2X0 U15507 ( .IN1(n16144), .IN2(n9157), .QN(WX11076) );
  NOR2X0 U15508 ( .IN1(n16143), .IN2(n9157), .QN(WX11074) );
  NOR2X0 U15509 ( .IN1(n16142), .IN2(n9157), .QN(WX11072) );
  NOR2X0 U15510 ( .IN1(n16141), .IN2(n9157), .QN(WX11070) );
  NOR2X0 U15511 ( .IN1(n16140), .IN2(n9157), .QN(WX11068) );
  NOR2X0 U15512 ( .IN1(n16139), .IN2(n9157), .QN(WX11066) );
  NOR2X0 U15513 ( .IN1(n9227), .IN2(n8825), .QN(WX11064) );
  NOR2X0 U15514 ( .IN1(n16138), .IN2(n9157), .QN(WX11062) );
  NOR2X0 U15515 ( .IN1(n16137), .IN2(n9156), .QN(WX11060) );
  NOR2X0 U15516 ( .IN1(n16136), .IN2(n9156), .QN(WX11058) );
  NOR2X0 U15517 ( .IN1(n16135), .IN2(n9156), .QN(WX11056) );
  NOR2X0 U15518 ( .IN1(n16134), .IN2(n9155), .QN(WX11054) );
  NOR2X0 U15519 ( .IN1(n16133), .IN2(n9156), .QN(WX11052) );
  NAND4X0 U15520 ( .IN1(n14840), .IN2(n14841), .IN3(n14842), .IN4(n14843), 
        .QN(WX11050) );
  NAND2X0 U15521 ( .IN1(n9102), .IN2(n9682), .QN(n14843) );
  NAND2X0 U15522 ( .IN1(n14844), .IN2(n14845), .QN(n9682) );
  INVX0 U15523 ( .INP(n14846), .ZN(n14845) );
  NOR2X0 U15524 ( .IN1(n14847), .IN2(n14848), .QN(n14846) );
  NAND2X0 U15525 ( .IN1(n14848), .IN2(n14847), .QN(n14844) );
  NOR2X0 U15526 ( .IN1(n14849), .IN2(n14850), .QN(n14847) );
  NOR2X0 U15527 ( .IN1(WX11243), .IN2(n7854), .QN(n14850) );
  INVX0 U15528 ( .INP(n14851), .ZN(n14849) );
  NAND2X0 U15529 ( .IN1(n7854), .IN2(WX11243), .QN(n14851) );
  NAND2X0 U15530 ( .IN1(n14852), .IN2(n14853), .QN(n14848) );
  NAND2X0 U15531 ( .IN1(n7853), .IN2(WX11115), .QN(n14853) );
  INVX0 U15532 ( .INP(n14854), .ZN(n14852) );
  NOR2X0 U15533 ( .IN1(WX11115), .IN2(n7853), .QN(n14854) );
  NAND2X0 U15534 ( .IN1(n1968), .IN2(n9286), .QN(n14842) );
  NOR2X0 U15535 ( .IN1(n9227), .IN2(n9031), .QN(n1968) );
  NAND2X0 U15536 ( .IN1(DATA_0_0), .IN2(n9335), .QN(n14841) );
  NAND2X0 U15537 ( .IN1(n9300), .IN2(CRC_OUT_1_0), .QN(n14840) );
  NAND4X0 U15538 ( .IN1(n14855), .IN2(n14856), .IN3(n14857), .IN4(n14858), 
        .QN(WX11048) );
  NAND2X0 U15539 ( .IN1(n9102), .IN2(n9689), .QN(n14858) );
  NAND2X0 U15540 ( .IN1(n14859), .IN2(n14860), .QN(n9689) );
  INVX0 U15541 ( .INP(n14861), .ZN(n14860) );
  NOR2X0 U15542 ( .IN1(n14862), .IN2(n14863), .QN(n14861) );
  NAND2X0 U15543 ( .IN1(n14863), .IN2(n14862), .QN(n14859) );
  NOR2X0 U15544 ( .IN1(n14864), .IN2(n14865), .QN(n14862) );
  NOR2X0 U15545 ( .IN1(WX11241), .IN2(n7856), .QN(n14865) );
  INVX0 U15546 ( .INP(n14866), .ZN(n14864) );
  NAND2X0 U15547 ( .IN1(n7856), .IN2(WX11241), .QN(n14866) );
  NAND2X0 U15548 ( .IN1(n14867), .IN2(n14868), .QN(n14863) );
  NAND2X0 U15549 ( .IN1(n7855), .IN2(WX11113), .QN(n14868) );
  INVX0 U15550 ( .INP(n14869), .ZN(n14867) );
  NOR2X0 U15551 ( .IN1(WX11113), .IN2(n7855), .QN(n14869) );
  NAND2X0 U15552 ( .IN1(n1967), .IN2(n9286), .QN(n14857) );
  NOR2X0 U15553 ( .IN1(n9227), .IN2(n9032), .QN(n1967) );
  NAND2X0 U15554 ( .IN1(DATA_0_1), .IN2(n9335), .QN(n14856) );
  NAND2X0 U15555 ( .IN1(n9300), .IN2(CRC_OUT_1_1), .QN(n14855) );
  NAND4X0 U15556 ( .IN1(n14870), .IN2(n14871), .IN3(n14872), .IN4(n14873), 
        .QN(WX11046) );
  NAND3X0 U15557 ( .IN1(n9694), .IN2(n9695), .IN3(n9091), .QN(n14873) );
  NAND3X0 U15558 ( .IN1(n14874), .IN2(n14875), .IN3(n14876), .QN(n9695) );
  INVX0 U15559 ( .INP(n14877), .ZN(n14876) );
  NAND2X0 U15560 ( .IN1(n14877), .IN2(n14878), .QN(n9694) );
  NAND2X0 U15561 ( .IN1(n14874), .IN2(n14875), .QN(n14878) );
  NAND2X0 U15562 ( .IN1(n7858), .IN2(WX11111), .QN(n14875) );
  NAND2X0 U15563 ( .IN1(n3535), .IN2(WX11175), .QN(n14874) );
  NOR2X0 U15564 ( .IN1(n14879), .IN2(n14880), .QN(n14877) );
  NOR2X0 U15565 ( .IN1(n8793), .IN2(n7857), .QN(n14880) );
  INVX0 U15566 ( .INP(n14881), .ZN(n14879) );
  NAND2X0 U15567 ( .IN1(n7857), .IN2(n8793), .QN(n14881) );
  NAND2X0 U15568 ( .IN1(n1966), .IN2(n9286), .QN(n14872) );
  NOR2X0 U15569 ( .IN1(n9227), .IN2(n9033), .QN(n1966) );
  NAND2X0 U15570 ( .IN1(DATA_0_2), .IN2(n9335), .QN(n14871) );
  NAND2X0 U15571 ( .IN1(n9300), .IN2(CRC_OUT_1_2), .QN(n14870) );
  NAND4X0 U15572 ( .IN1(n14882), .IN2(n14883), .IN3(n14884), .IN4(n14885), 
        .QN(WX11044) );
  NAND2X0 U15573 ( .IN1(n9102), .IN2(n9703), .QN(n14885) );
  NAND2X0 U15574 ( .IN1(n14886), .IN2(n14887), .QN(n9703) );
  INVX0 U15575 ( .INP(n14888), .ZN(n14887) );
  NOR2X0 U15576 ( .IN1(n14889), .IN2(n14890), .QN(n14888) );
  NAND2X0 U15577 ( .IN1(n14890), .IN2(n14889), .QN(n14886) );
  NOR2X0 U15578 ( .IN1(n14891), .IN2(n14892), .QN(n14889) );
  NOR2X0 U15579 ( .IN1(WX11237), .IN2(n7860), .QN(n14892) );
  INVX0 U15580 ( .INP(n14893), .ZN(n14891) );
  NAND2X0 U15581 ( .IN1(n7860), .IN2(WX11237), .QN(n14893) );
  NAND2X0 U15582 ( .IN1(n14894), .IN2(n14895), .QN(n14890) );
  NAND2X0 U15583 ( .IN1(n7859), .IN2(WX11109), .QN(n14895) );
  INVX0 U15584 ( .INP(n14896), .ZN(n14894) );
  NOR2X0 U15585 ( .IN1(WX11109), .IN2(n7859), .QN(n14896) );
  NAND2X0 U15586 ( .IN1(n1965), .IN2(n9286), .QN(n14884) );
  NOR2X0 U15587 ( .IN1(n9227), .IN2(n9034), .QN(n1965) );
  NAND2X0 U15588 ( .IN1(DATA_0_3), .IN2(n9335), .QN(n14883) );
  NAND2X0 U15589 ( .IN1(n9300), .IN2(CRC_OUT_1_3), .QN(n14882) );
  NAND4X0 U15590 ( .IN1(n14897), .IN2(n14898), .IN3(n14899), .IN4(n14900), 
        .QN(WX11042) );
  NAND3X0 U15591 ( .IN1(n9708), .IN2(n9709), .IN3(n9091), .QN(n14900) );
  NAND3X0 U15592 ( .IN1(n14901), .IN2(n14902), .IN3(n14903), .QN(n9709) );
  INVX0 U15593 ( .INP(n14904), .ZN(n14903) );
  NAND2X0 U15594 ( .IN1(n14904), .IN2(n14905), .QN(n9708) );
  NAND2X0 U15595 ( .IN1(n14901), .IN2(n14902), .QN(n14905) );
  NAND2X0 U15596 ( .IN1(n8106), .IN2(WX11107), .QN(n14902) );
  NAND2X0 U15597 ( .IN1(n3539), .IN2(WX11235), .QN(n14901) );
  NOR2X0 U15598 ( .IN1(n14906), .IN2(n14907), .QN(n14904) );
  INVX0 U15599 ( .INP(n14908), .ZN(n14907) );
  NAND2X0 U15600 ( .IN1(test_so96), .IN2(WX11043), .QN(n14908) );
  NOR2X0 U15601 ( .IN1(WX11043), .IN2(test_so96), .QN(n14906) );
  NAND2X0 U15602 ( .IN1(n1964), .IN2(n9286), .QN(n14899) );
  NOR2X0 U15603 ( .IN1(n9227), .IN2(n9035), .QN(n1964) );
  NAND2X0 U15604 ( .IN1(DATA_0_4), .IN2(n9335), .QN(n14898) );
  NAND2X0 U15605 ( .IN1(n9300), .IN2(CRC_OUT_1_4), .QN(n14897) );
  NAND4X0 U15606 ( .IN1(n14909), .IN2(n14910), .IN3(n14911), .IN4(n14912), 
        .QN(WX11040) );
  NAND2X0 U15607 ( .IN1(n9102), .IN2(n9716), .QN(n14912) );
  NAND2X0 U15608 ( .IN1(n14913), .IN2(n14914), .QN(n9716) );
  INVX0 U15609 ( .INP(n14915), .ZN(n14914) );
  NOR2X0 U15610 ( .IN1(n14916), .IN2(n14917), .QN(n14915) );
  NAND2X0 U15611 ( .IN1(n14917), .IN2(n14916), .QN(n14913) );
  NOR2X0 U15612 ( .IN1(n14918), .IN2(n14919), .QN(n14916) );
  NOR2X0 U15613 ( .IN1(WX11233), .IN2(n7863), .QN(n14919) );
  INVX0 U15614 ( .INP(n14920), .ZN(n14918) );
  NAND2X0 U15615 ( .IN1(n7863), .IN2(WX11233), .QN(n14920) );
  NAND2X0 U15616 ( .IN1(n14921), .IN2(n14922), .QN(n14917) );
  NAND2X0 U15617 ( .IN1(n7862), .IN2(WX11105), .QN(n14922) );
  INVX0 U15618 ( .INP(n14923), .ZN(n14921) );
  NOR2X0 U15619 ( .IN1(WX11105), .IN2(n7862), .QN(n14923) );
  NAND2X0 U15620 ( .IN1(n1963), .IN2(n9286), .QN(n14911) );
  NOR2X0 U15621 ( .IN1(n9228), .IN2(n9036), .QN(n1963) );
  NAND2X0 U15622 ( .IN1(DATA_0_5), .IN2(n9335), .QN(n14910) );
  NAND2X0 U15623 ( .IN1(n9300), .IN2(CRC_OUT_1_5), .QN(n14909) );
  NAND4X0 U15624 ( .IN1(n14924), .IN2(n14925), .IN3(n14926), .IN4(n14927), 
        .QN(WX11038) );
  NAND3X0 U15625 ( .IN1(n9721), .IN2(n9722), .IN3(n9090), .QN(n14927) );
  NAND3X0 U15626 ( .IN1(n14928), .IN2(n14929), .IN3(n14930), .QN(n9722) );
  INVX0 U15627 ( .INP(n14931), .ZN(n14930) );
  NAND2X0 U15628 ( .IN1(n14931), .IN2(n14932), .QN(n9721) );
  NAND2X0 U15629 ( .IN1(n14928), .IN2(n14929), .QN(n14932) );
  NAND2X0 U15630 ( .IN1(n8155), .IN2(WX11167), .QN(n14929) );
  NAND2X0 U15631 ( .IN1(n7865), .IN2(WX11231), .QN(n14928) );
  NOR2X0 U15632 ( .IN1(n14933), .IN2(n14934), .QN(n14931) );
  INVX0 U15633 ( .INP(n14935), .ZN(n14934) );
  NAND2X0 U15634 ( .IN1(test_so94), .IN2(WX11039), .QN(n14935) );
  NOR2X0 U15635 ( .IN1(WX11039), .IN2(test_so94), .QN(n14933) );
  NAND2X0 U15636 ( .IN1(n1962), .IN2(n9287), .QN(n14926) );
  NOR2X0 U15637 ( .IN1(n9228), .IN2(n9037), .QN(n1962) );
  NAND2X0 U15638 ( .IN1(DATA_0_6), .IN2(n9334), .QN(n14925) );
  NAND2X0 U15639 ( .IN1(n9300), .IN2(CRC_OUT_1_6), .QN(n14924) );
  NAND4X0 U15640 ( .IN1(n14936), .IN2(n14937), .IN3(n14938), .IN4(n14939), 
        .QN(WX11036) );
  NAND2X0 U15641 ( .IN1(n9102), .IN2(n9729), .QN(n14939) );
  NAND2X0 U15642 ( .IN1(n14940), .IN2(n14941), .QN(n9729) );
  INVX0 U15643 ( .INP(n14942), .ZN(n14941) );
  NOR2X0 U15644 ( .IN1(n14943), .IN2(n14944), .QN(n14942) );
  NAND2X0 U15645 ( .IN1(n14944), .IN2(n14943), .QN(n14940) );
  NOR2X0 U15646 ( .IN1(n14945), .IN2(n14946), .QN(n14943) );
  NOR2X0 U15647 ( .IN1(WX11229), .IN2(n7867), .QN(n14946) );
  INVX0 U15648 ( .INP(n14947), .ZN(n14945) );
  NAND2X0 U15649 ( .IN1(n7867), .IN2(WX11229), .QN(n14947) );
  NAND2X0 U15650 ( .IN1(n14948), .IN2(n14949), .QN(n14944) );
  NAND2X0 U15651 ( .IN1(n7866), .IN2(WX11101), .QN(n14949) );
  INVX0 U15652 ( .INP(n14950), .ZN(n14948) );
  NOR2X0 U15653 ( .IN1(WX11101), .IN2(n7866), .QN(n14950) );
  NAND2X0 U15654 ( .IN1(n1961), .IN2(n9287), .QN(n14938) );
  NOR2X0 U15655 ( .IN1(n9228), .IN2(n9038), .QN(n1961) );
  NAND2X0 U15656 ( .IN1(DATA_0_7), .IN2(n9335), .QN(n14937) );
  NAND2X0 U15657 ( .IN1(n9300), .IN2(CRC_OUT_1_7), .QN(n14936) );
  NAND4X0 U15658 ( .IN1(n14951), .IN2(n14952), .IN3(n14953), .IN4(n14954), 
        .QN(WX11034) );
  NAND3X0 U15659 ( .IN1(n9734), .IN2(n9735), .IN3(n9090), .QN(n14954) );
  NAND3X0 U15660 ( .IN1(n14955), .IN2(n14956), .IN3(n14957), .QN(n9735) );
  INVX0 U15661 ( .INP(n14958), .ZN(n14957) );
  NAND2X0 U15662 ( .IN1(n14958), .IN2(n14959), .QN(n9734) );
  NAND2X0 U15663 ( .IN1(n14955), .IN2(n14956), .QN(n14959) );
  NAND2X0 U15664 ( .IN1(n8153), .IN2(WX11099), .QN(n14956) );
  NAND2X0 U15665 ( .IN1(n3547), .IN2(WX11227), .QN(n14955) );
  NOR2X0 U15666 ( .IN1(n14960), .IN2(n14961), .QN(n14958) );
  INVX0 U15667 ( .INP(n14962), .ZN(n14961) );
  NAND2X0 U15668 ( .IN1(test_so92), .IN2(WX11163), .QN(n14962) );
  NOR2X0 U15669 ( .IN1(WX11163), .IN2(test_so92), .QN(n14960) );
  NAND2X0 U15670 ( .IN1(n1960), .IN2(n9287), .QN(n14953) );
  NOR2X0 U15671 ( .IN1(n9228), .IN2(n9039), .QN(n1960) );
  NAND2X0 U15672 ( .IN1(DATA_0_8), .IN2(n9334), .QN(n14952) );
  NAND2X0 U15673 ( .IN1(n9300), .IN2(CRC_OUT_1_8), .QN(n14951) );
  NAND4X0 U15674 ( .IN1(n14963), .IN2(n14964), .IN3(n14965), .IN4(n14966), 
        .QN(WX11032) );
  NAND2X0 U15675 ( .IN1(n9102), .IN2(n9742), .QN(n14966) );
  NAND2X0 U15676 ( .IN1(n14967), .IN2(n14968), .QN(n9742) );
  INVX0 U15677 ( .INP(n14969), .ZN(n14968) );
  NOR2X0 U15678 ( .IN1(n14970), .IN2(n14971), .QN(n14969) );
  NAND2X0 U15679 ( .IN1(n14971), .IN2(n14970), .QN(n14967) );
  NOR2X0 U15680 ( .IN1(n14972), .IN2(n14973), .QN(n14970) );
  NOR2X0 U15681 ( .IN1(WX11225), .IN2(n7870), .QN(n14973) );
  INVX0 U15682 ( .INP(n14974), .ZN(n14972) );
  NAND2X0 U15683 ( .IN1(n7870), .IN2(WX11225), .QN(n14974) );
  NAND2X0 U15684 ( .IN1(n14975), .IN2(n14976), .QN(n14971) );
  NAND2X0 U15685 ( .IN1(n7869), .IN2(WX11097), .QN(n14976) );
  INVX0 U15686 ( .INP(n14977), .ZN(n14975) );
  NOR2X0 U15687 ( .IN1(WX11097), .IN2(n7869), .QN(n14977) );
  NAND2X0 U15688 ( .IN1(n1959), .IN2(n9287), .QN(n14965) );
  NOR2X0 U15689 ( .IN1(n9228), .IN2(n9040), .QN(n1959) );
  NAND2X0 U15690 ( .IN1(DATA_0_9), .IN2(n9334), .QN(n14964) );
  NAND2X0 U15691 ( .IN1(n9300), .IN2(CRC_OUT_1_9), .QN(n14963) );
  NAND4X0 U15692 ( .IN1(n14978), .IN2(n14979), .IN3(n14980), .IN4(n14981), 
        .QN(WX11030) );
  NAND2X0 U15693 ( .IN1(n9102), .IN2(n9748), .QN(n14981) );
  NAND2X0 U15694 ( .IN1(n14982), .IN2(n14983), .QN(n9748) );
  INVX0 U15695 ( .INP(n14984), .ZN(n14983) );
  NOR2X0 U15696 ( .IN1(n14985), .IN2(n14986), .QN(n14984) );
  NAND2X0 U15697 ( .IN1(n14986), .IN2(n14985), .QN(n14982) );
  NOR2X0 U15698 ( .IN1(n14987), .IN2(n14988), .QN(n14985) );
  NOR2X0 U15699 ( .IN1(WX11223), .IN2(n7872), .QN(n14988) );
  INVX0 U15700 ( .INP(n14989), .ZN(n14987) );
  NAND2X0 U15701 ( .IN1(n7872), .IN2(WX11223), .QN(n14989) );
  NAND2X0 U15702 ( .IN1(n14990), .IN2(n14991), .QN(n14986) );
  NAND2X0 U15703 ( .IN1(n7871), .IN2(WX11095), .QN(n14991) );
  INVX0 U15704 ( .INP(n14992), .ZN(n14990) );
  NOR2X0 U15705 ( .IN1(WX11095), .IN2(n7871), .QN(n14992) );
  NAND2X0 U15706 ( .IN1(n1958), .IN2(n9287), .QN(n14980) );
  NOR2X0 U15707 ( .IN1(n9074), .IN2(n9155), .QN(n1958) );
  NAND2X0 U15708 ( .IN1(DATA_0_10), .IN2(n9334), .QN(n14979) );
  NAND2X0 U15709 ( .IN1(n9300), .IN2(CRC_OUT_1_10), .QN(n14978) );
  NAND4X0 U15710 ( .IN1(n14993), .IN2(n14994), .IN3(n14995), .IN4(n14996), 
        .QN(WX11028) );
  NAND2X0 U15711 ( .IN1(n9102), .IN2(n9754), .QN(n14996) );
  NAND2X0 U15712 ( .IN1(n14997), .IN2(n14998), .QN(n9754) );
  INVX0 U15713 ( .INP(n14999), .ZN(n14998) );
  NOR2X0 U15714 ( .IN1(n15000), .IN2(n15001), .QN(n14999) );
  NAND2X0 U15715 ( .IN1(n15001), .IN2(n15000), .QN(n14997) );
  NOR2X0 U15716 ( .IN1(n15002), .IN2(n15003), .QN(n15000) );
  NOR2X0 U15717 ( .IN1(WX11221), .IN2(n7874), .QN(n15003) );
  INVX0 U15718 ( .INP(n15004), .ZN(n15002) );
  NAND2X0 U15719 ( .IN1(n7874), .IN2(WX11221), .QN(n15004) );
  NAND2X0 U15720 ( .IN1(n15005), .IN2(n15006), .QN(n15001) );
  NAND2X0 U15721 ( .IN1(n7873), .IN2(WX11093), .QN(n15006) );
  INVX0 U15722 ( .INP(n15007), .ZN(n15005) );
  NOR2X0 U15723 ( .IN1(WX11093), .IN2(n7873), .QN(n15007) );
  NAND2X0 U15724 ( .IN1(n1957), .IN2(n9287), .QN(n14995) );
  NOR2X0 U15725 ( .IN1(n9228), .IN2(n9041), .QN(n1957) );
  NAND2X0 U15726 ( .IN1(DATA_0_11), .IN2(n9334), .QN(n14994) );
  NAND2X0 U15727 ( .IN1(n9301), .IN2(CRC_OUT_1_11), .QN(n14993) );
  NAND4X0 U15728 ( .IN1(n15008), .IN2(n15009), .IN3(n15010), .IN4(n15011), 
        .QN(WX11026) );
  NAND2X0 U15729 ( .IN1(n9102), .IN2(n9760), .QN(n15011) );
  NAND2X0 U15730 ( .IN1(n15012), .IN2(n15013), .QN(n9760) );
  INVX0 U15731 ( .INP(n15014), .ZN(n15013) );
  NOR2X0 U15732 ( .IN1(n15015), .IN2(n15016), .QN(n15014) );
  NAND2X0 U15733 ( .IN1(n15016), .IN2(n15015), .QN(n15012) );
  NOR2X0 U15734 ( .IN1(n15017), .IN2(n15018), .QN(n15015) );
  NOR2X0 U15735 ( .IN1(WX11219), .IN2(n7876), .QN(n15018) );
  INVX0 U15736 ( .INP(n15019), .ZN(n15017) );
  NAND2X0 U15737 ( .IN1(n7876), .IN2(WX11219), .QN(n15019) );
  NAND2X0 U15738 ( .IN1(n15020), .IN2(n15021), .QN(n15016) );
  NAND2X0 U15739 ( .IN1(n7875), .IN2(WX11091), .QN(n15021) );
  INVX0 U15740 ( .INP(n15022), .ZN(n15020) );
  NOR2X0 U15741 ( .IN1(WX11091), .IN2(n7875), .QN(n15022) );
  NAND2X0 U15742 ( .IN1(n1956), .IN2(n9287), .QN(n15010) );
  NOR2X0 U15743 ( .IN1(n9228), .IN2(n9042), .QN(n1956) );
  NAND2X0 U15744 ( .IN1(DATA_0_12), .IN2(n9334), .QN(n15009) );
  NAND2X0 U15745 ( .IN1(n9301), .IN2(CRC_OUT_1_12), .QN(n15008) );
  NAND4X0 U15746 ( .IN1(n15023), .IN2(n15024), .IN3(n15025), .IN4(n15026), 
        .QN(WX11024) );
  NAND2X0 U15747 ( .IN1(n9101), .IN2(n9766), .QN(n15026) );
  NAND2X0 U15748 ( .IN1(n15027), .IN2(n15028), .QN(n9766) );
  INVX0 U15749 ( .INP(n15029), .ZN(n15028) );
  NOR2X0 U15750 ( .IN1(n15030), .IN2(n15031), .QN(n15029) );
  NAND2X0 U15751 ( .IN1(n15031), .IN2(n15030), .QN(n15027) );
  NOR2X0 U15752 ( .IN1(n15032), .IN2(n15033), .QN(n15030) );
  NOR2X0 U15753 ( .IN1(WX11217), .IN2(n7878), .QN(n15033) );
  INVX0 U15754 ( .INP(n15034), .ZN(n15032) );
  NAND2X0 U15755 ( .IN1(n7878), .IN2(WX11217), .QN(n15034) );
  NAND2X0 U15756 ( .IN1(n15035), .IN2(n15036), .QN(n15031) );
  NAND2X0 U15757 ( .IN1(n7877), .IN2(WX11089), .QN(n15036) );
  INVX0 U15758 ( .INP(n15037), .ZN(n15035) );
  NOR2X0 U15759 ( .IN1(WX11089), .IN2(n7877), .QN(n15037) );
  NAND2X0 U15760 ( .IN1(n1955), .IN2(n9287), .QN(n15025) );
  NOR2X0 U15761 ( .IN1(n9228), .IN2(n9043), .QN(n1955) );
  NAND2X0 U15762 ( .IN1(DATA_0_13), .IN2(n9334), .QN(n15024) );
  NAND2X0 U15763 ( .IN1(n9301), .IN2(CRC_OUT_1_13), .QN(n15023) );
  NAND4X0 U15764 ( .IN1(n15038), .IN2(n15039), .IN3(n15040), .IN4(n15041), 
        .QN(WX11022) );
  NAND2X0 U15765 ( .IN1(n9101), .IN2(n9773), .QN(n15041) );
  NAND2X0 U15766 ( .IN1(n15042), .IN2(n15043), .QN(n9773) );
  INVX0 U15767 ( .INP(n15044), .ZN(n15043) );
  NOR2X0 U15768 ( .IN1(n15045), .IN2(n15046), .QN(n15044) );
  NAND2X0 U15769 ( .IN1(n15046), .IN2(n15045), .QN(n15042) );
  NOR2X0 U15770 ( .IN1(n15047), .IN2(n15048), .QN(n15045) );
  NOR2X0 U15771 ( .IN1(WX11215), .IN2(n7880), .QN(n15048) );
  INVX0 U15772 ( .INP(n15049), .ZN(n15047) );
  NAND2X0 U15773 ( .IN1(n7880), .IN2(WX11215), .QN(n15049) );
  NAND2X0 U15774 ( .IN1(n15050), .IN2(n15051), .QN(n15046) );
  NAND2X0 U15775 ( .IN1(n7879), .IN2(WX11087), .QN(n15051) );
  INVX0 U15776 ( .INP(n15052), .ZN(n15050) );
  NOR2X0 U15777 ( .IN1(WX11087), .IN2(n7879), .QN(n15052) );
  NAND2X0 U15778 ( .IN1(n1954), .IN2(n9287), .QN(n15040) );
  NOR2X0 U15779 ( .IN1(n9228), .IN2(n9044), .QN(n1954) );
  NAND2X0 U15780 ( .IN1(DATA_0_14), .IN2(n9334), .QN(n15039) );
  NAND2X0 U15781 ( .IN1(test_so99), .IN2(n9313), .QN(n15038) );
  NAND4X0 U15782 ( .IN1(n15053), .IN2(n15054), .IN3(n15055), .IN4(n15056), 
        .QN(WX11020) );
  NAND2X0 U15783 ( .IN1(n9101), .IN2(n9779), .QN(n15056) );
  NAND2X0 U15784 ( .IN1(n15057), .IN2(n15058), .QN(n9779) );
  INVX0 U15785 ( .INP(n15059), .ZN(n15058) );
  NOR2X0 U15786 ( .IN1(n15060), .IN2(n15061), .QN(n15059) );
  NAND2X0 U15787 ( .IN1(n15061), .IN2(n15060), .QN(n15057) );
  NOR2X0 U15788 ( .IN1(n15062), .IN2(n15063), .QN(n15060) );
  NOR2X0 U15789 ( .IN1(WX11213), .IN2(n7882), .QN(n15063) );
  INVX0 U15790 ( .INP(n15064), .ZN(n15062) );
  NAND2X0 U15791 ( .IN1(n7882), .IN2(WX11213), .QN(n15064) );
  NAND2X0 U15792 ( .IN1(n15065), .IN2(n15066), .QN(n15061) );
  NAND2X0 U15793 ( .IN1(n7881), .IN2(WX11085), .QN(n15066) );
  INVX0 U15794 ( .INP(n15067), .ZN(n15065) );
  NOR2X0 U15795 ( .IN1(WX11085), .IN2(n7881), .QN(n15067) );
  NAND2X0 U15796 ( .IN1(n1953), .IN2(n9287), .QN(n15055) );
  NOR2X0 U15797 ( .IN1(n9228), .IN2(n9045), .QN(n1953) );
  NAND2X0 U15798 ( .IN1(DATA_0_15), .IN2(n9334), .QN(n15054) );
  NAND2X0 U15799 ( .IN1(n9301), .IN2(CRC_OUT_1_15), .QN(n15053) );
  NAND4X0 U15800 ( .IN1(n15068), .IN2(n15069), .IN3(n15070), .IN4(n15071), 
        .QN(WX11018) );
  NAND2X0 U15801 ( .IN1(n15072), .IN2(n9785), .QN(n15071) );
  NAND2X0 U15802 ( .IN1(n15073), .IN2(n9789), .QN(n9785) );
  NAND2X0 U15803 ( .IN1(n15074), .IN2(n15075), .QN(n15073) );
  NAND2X0 U15804 ( .IN1(n16147), .IN2(n9122), .QN(n15075) );
  NAND2X0 U15805 ( .IN1(TM1), .IN2(n8246), .QN(n15074) );
  NAND2X0 U15806 ( .IN1(n15076), .IN2(n15077), .QN(n15072) );
  NAND2X0 U15807 ( .IN1(n9101), .IN2(n9789), .QN(n15077) );
  NAND2X0 U15808 ( .IN1(n15078), .IN2(n15079), .QN(n9789) );
  NAND2X0 U15809 ( .IN1(n7627), .IN2(n15080), .QN(n15079) );
  INVX0 U15810 ( .INP(n15081), .ZN(n15078) );
  NOR2X0 U15811 ( .IN1(n15080), .IN2(n7627), .QN(n15081) );
  NOR2X0 U15812 ( .IN1(n15082), .IN2(n15083), .QN(n15080) );
  NOR2X0 U15813 ( .IN1(WX11211), .IN2(n7628), .QN(n15083) );
  INVX0 U15814 ( .INP(n15084), .ZN(n15082) );
  NAND2X0 U15815 ( .IN1(n7628), .IN2(WX11211), .QN(n15084) );
  NAND2X0 U15816 ( .IN1(n9101), .IN2(n8246), .QN(n15076) );
  NAND2X0 U15817 ( .IN1(n1952), .IN2(n9287), .QN(n15070) );
  NOR2X0 U15818 ( .IN1(n9228), .IN2(n9046), .QN(n1952) );
  NAND2X0 U15819 ( .IN1(DATA_0_16), .IN2(n9334), .QN(n15069) );
  NAND2X0 U15820 ( .IN1(n9301), .IN2(CRC_OUT_1_16), .QN(n15068) );
  NAND4X0 U15821 ( .IN1(n15085), .IN2(n15086), .IN3(n15087), .IN4(n15088), 
        .QN(WX11016) );
  NAND2X0 U15822 ( .IN1(n15089), .IN2(n9803), .QN(n15088) );
  NAND2X0 U15823 ( .IN1(n15090), .IN2(n9807), .QN(n9803) );
  NAND2X0 U15824 ( .IN1(n15091), .IN2(n15092), .QN(n15090) );
  NAND2X0 U15825 ( .IN1(n16146), .IN2(n9122), .QN(n15092) );
  NAND2X0 U15826 ( .IN1(TM1), .IN2(n8247), .QN(n15091) );
  NAND2X0 U15827 ( .IN1(n15093), .IN2(n15094), .QN(n15089) );
  NAND2X0 U15828 ( .IN1(n9101), .IN2(n9807), .QN(n15094) );
  NAND2X0 U15829 ( .IN1(n15095), .IN2(n15096), .QN(n9807) );
  NAND2X0 U15830 ( .IN1(n7629), .IN2(n15097), .QN(n15096) );
  INVX0 U15831 ( .INP(n15098), .ZN(n15095) );
  NOR2X0 U15832 ( .IN1(n15097), .IN2(n7629), .QN(n15098) );
  NOR2X0 U15833 ( .IN1(n15099), .IN2(n15100), .QN(n15097) );
  NOR2X0 U15834 ( .IN1(WX11209), .IN2(n7630), .QN(n15100) );
  INVX0 U15835 ( .INP(n15101), .ZN(n15099) );
  NAND2X0 U15836 ( .IN1(n7630), .IN2(WX11209), .QN(n15101) );
  NAND2X0 U15837 ( .IN1(n9101), .IN2(n8247), .QN(n15093) );
  NAND2X0 U15838 ( .IN1(n1951), .IN2(n9287), .QN(n15087) );
  NOR2X0 U15839 ( .IN1(n9228), .IN2(n9047), .QN(n1951) );
  NAND2X0 U15840 ( .IN1(DATA_0_17), .IN2(n9334), .QN(n15086) );
  NAND2X0 U15841 ( .IN1(n9301), .IN2(CRC_OUT_1_17), .QN(n15085) );
  NAND4X0 U15842 ( .IN1(n15102), .IN2(n15103), .IN3(n15104), .IN4(n15105), 
        .QN(WX11014) );
  NAND2X0 U15843 ( .IN1(n15106), .IN2(n9813), .QN(n15105) );
  NAND2X0 U15844 ( .IN1(n15107), .IN2(n9817), .QN(n9813) );
  NAND2X0 U15845 ( .IN1(n15108), .IN2(n15109), .QN(n15107) );
  NAND2X0 U15846 ( .IN1(n16145), .IN2(n9122), .QN(n15109) );
  NAND2X0 U15847 ( .IN1(TM1), .IN2(n8248), .QN(n15108) );
  NAND2X0 U15848 ( .IN1(n15110), .IN2(n15111), .QN(n15106) );
  NAND2X0 U15849 ( .IN1(n9101), .IN2(n9817), .QN(n15111) );
  NAND2X0 U15850 ( .IN1(n15112), .IN2(n15113), .QN(n9817) );
  NAND2X0 U15851 ( .IN1(n7631), .IN2(n15114), .QN(n15113) );
  INVX0 U15852 ( .INP(n15115), .ZN(n15112) );
  NOR2X0 U15853 ( .IN1(n15114), .IN2(n7631), .QN(n15115) );
  NOR2X0 U15854 ( .IN1(n15116), .IN2(n15117), .QN(n15114) );
  NOR2X0 U15855 ( .IN1(WX11207), .IN2(n7632), .QN(n15117) );
  INVX0 U15856 ( .INP(n15118), .ZN(n15116) );
  NAND2X0 U15857 ( .IN1(n7632), .IN2(WX11207), .QN(n15118) );
  NAND2X0 U15858 ( .IN1(n9105), .IN2(n8248), .QN(n15110) );
  NAND2X0 U15859 ( .IN1(n1950), .IN2(n9287), .QN(n15104) );
  NOR2X0 U15860 ( .IN1(n9228), .IN2(n9048), .QN(n1950) );
  NAND2X0 U15861 ( .IN1(DATA_0_18), .IN2(n9334), .QN(n15103) );
  NAND2X0 U15862 ( .IN1(n9301), .IN2(CRC_OUT_1_18), .QN(n15102) );
  NAND4X0 U15863 ( .IN1(n15119), .IN2(n15120), .IN3(n15121), .IN4(n15122), 
        .QN(WX11012) );
  NAND2X0 U15864 ( .IN1(n9828), .IN2(n9110), .QN(n15122) );
  NOR2X0 U15865 ( .IN1(n15123), .IN2(n15124), .QN(n9828) );
  INVX0 U15866 ( .INP(n15125), .ZN(n15124) );
  NAND2X0 U15867 ( .IN1(n15126), .IN2(n15127), .QN(n15125) );
  NOR2X0 U15868 ( .IN1(n15127), .IN2(n15126), .QN(n15123) );
  NAND2X0 U15869 ( .IN1(n15128), .IN2(n15129), .QN(n15126) );
  NAND2X0 U15870 ( .IN1(n15130), .IN2(WX11141), .QN(n15129) );
  NAND2X0 U15871 ( .IN1(n15131), .IN2(n15132), .QN(n15130) );
  NAND3X0 U15872 ( .IN1(n15131), .IN2(n15132), .IN3(n7634), .QN(n15128) );
  NAND2X0 U15873 ( .IN1(test_so97), .IN2(WX11077), .QN(n15132) );
  NAND2X0 U15874 ( .IN1(n7633), .IN2(n8803), .QN(n15131) );
  NOR2X0 U15875 ( .IN1(n15133), .IN2(n15134), .QN(n15127) );
  INVX0 U15876 ( .INP(n15135), .ZN(n15134) );
  NAND2X0 U15877 ( .IN1(n16144), .IN2(n9122), .QN(n15135) );
  NOR2X0 U15878 ( .IN1(n9116), .IN2(n16144), .QN(n15133) );
  NAND2X0 U15879 ( .IN1(n1949), .IN2(n9287), .QN(n15121) );
  NOR2X0 U15880 ( .IN1(n9228), .IN2(n9049), .QN(n1949) );
  NAND2X0 U15881 ( .IN1(DATA_0_19), .IN2(n9334), .QN(n15120) );
  NAND2X0 U15882 ( .IN1(n9301), .IN2(CRC_OUT_1_19), .QN(n15119) );
  NAND4X0 U15883 ( .IN1(n15136), .IN2(n15137), .IN3(n15138), .IN4(n15139), 
        .QN(WX11010) );
  NAND2X0 U15884 ( .IN1(n15140), .IN2(n9839), .QN(n15139) );
  NAND2X0 U15885 ( .IN1(n15141), .IN2(n9843), .QN(n9839) );
  NAND2X0 U15886 ( .IN1(n15142), .IN2(n15143), .QN(n15141) );
  NAND2X0 U15887 ( .IN1(n16143), .IN2(n9122), .QN(n15143) );
  NAND2X0 U15888 ( .IN1(TM1), .IN2(n8250), .QN(n15142) );
  NAND2X0 U15889 ( .IN1(n15144), .IN2(n15145), .QN(n15140) );
  NAND2X0 U15890 ( .IN1(n9101), .IN2(n9843), .QN(n15145) );
  NAND2X0 U15891 ( .IN1(n15146), .IN2(n15147), .QN(n9843) );
  NAND2X0 U15892 ( .IN1(n7635), .IN2(n15148), .QN(n15147) );
  INVX0 U15893 ( .INP(n15149), .ZN(n15146) );
  NOR2X0 U15894 ( .IN1(n15148), .IN2(n7635), .QN(n15149) );
  NOR2X0 U15895 ( .IN1(n15150), .IN2(n15151), .QN(n15148) );
  NOR2X0 U15896 ( .IN1(WX11203), .IN2(n7636), .QN(n15151) );
  INVX0 U15897 ( .INP(n15152), .ZN(n15150) );
  NAND2X0 U15898 ( .IN1(n7636), .IN2(WX11203), .QN(n15152) );
  NAND2X0 U15899 ( .IN1(n9101), .IN2(n8250), .QN(n15144) );
  NAND2X0 U15900 ( .IN1(n1948), .IN2(n9287), .QN(n15138) );
  NOR2X0 U15901 ( .IN1(n9228), .IN2(n9050), .QN(n1948) );
  NAND2X0 U15902 ( .IN1(DATA_0_20), .IN2(n9334), .QN(n15137) );
  NAND2X0 U15903 ( .IN1(n9301), .IN2(CRC_OUT_1_20), .QN(n15136) );
  NAND4X0 U15904 ( .IN1(n15153), .IN2(n15154), .IN3(n15155), .IN4(n15156), 
        .QN(WX11008) );
  NAND2X0 U15905 ( .IN1(n9853), .IN2(n9110), .QN(n15156) );
  NOR2X0 U15906 ( .IN1(n15157), .IN2(n15158), .QN(n9853) );
  INVX0 U15907 ( .INP(n15159), .ZN(n15158) );
  NAND2X0 U15908 ( .IN1(n15160), .IN2(n15161), .QN(n15159) );
  NOR2X0 U15909 ( .IN1(n15161), .IN2(n15160), .QN(n15157) );
  NAND2X0 U15910 ( .IN1(n15162), .IN2(n15163), .QN(n15160) );
  NAND2X0 U15911 ( .IN1(n8143), .IN2(n15164), .QN(n15163) );
  INVX0 U15912 ( .INP(n15165), .ZN(n15164) );
  NAND2X0 U15913 ( .IN1(n15165), .IN2(WX11201), .QN(n15162) );
  NAND2X0 U15914 ( .IN1(n15166), .IN2(n15167), .QN(n15165) );
  INVX0 U15915 ( .INP(n15168), .ZN(n15167) );
  NOR2X0 U15916 ( .IN1(n8817), .IN2(n16142), .QN(n15168) );
  NAND2X0 U15917 ( .IN1(n16142), .IN2(n8817), .QN(n15166) );
  NOR2X0 U15918 ( .IN1(n15169), .IN2(n15170), .QN(n15161) );
  INVX0 U15919 ( .INP(n15171), .ZN(n15170) );
  NAND2X0 U15920 ( .IN1(n7637), .IN2(n9122), .QN(n15171) );
  NOR2X0 U15921 ( .IN1(n9117), .IN2(n7637), .QN(n15169) );
  NAND2X0 U15922 ( .IN1(n1947), .IN2(n9287), .QN(n15155) );
  NOR2X0 U15923 ( .IN1(n9229), .IN2(n9051), .QN(n1947) );
  NAND2X0 U15924 ( .IN1(DATA_0_21), .IN2(n9334), .QN(n15154) );
  NAND2X0 U15925 ( .IN1(n9301), .IN2(CRC_OUT_1_21), .QN(n15153) );
  NAND4X0 U15926 ( .IN1(n15172), .IN2(n15173), .IN3(n15174), .IN4(n15175), 
        .QN(WX11006) );
  NAND2X0 U15927 ( .IN1(n15176), .IN2(n9864), .QN(n15175) );
  NAND2X0 U15928 ( .IN1(n15177), .IN2(n9868), .QN(n9864) );
  NAND2X0 U15929 ( .IN1(n15178), .IN2(n15179), .QN(n15177) );
  NAND2X0 U15930 ( .IN1(n16141), .IN2(n9122), .QN(n15179) );
  NAND2X0 U15931 ( .IN1(TM1), .IN2(n8252), .QN(n15178) );
  NAND2X0 U15932 ( .IN1(n15180), .IN2(n15181), .QN(n15176) );
  NAND2X0 U15933 ( .IN1(n9101), .IN2(n9868), .QN(n15181) );
  NAND2X0 U15934 ( .IN1(n15182), .IN2(n15183), .QN(n9868) );
  NAND2X0 U15935 ( .IN1(n7638), .IN2(n15184), .QN(n15183) );
  INVX0 U15936 ( .INP(n15185), .ZN(n15182) );
  NOR2X0 U15937 ( .IN1(n15184), .IN2(n7638), .QN(n15185) );
  NOR2X0 U15938 ( .IN1(n15186), .IN2(n15187), .QN(n15184) );
  NOR2X0 U15939 ( .IN1(WX11199), .IN2(n7639), .QN(n15187) );
  INVX0 U15940 ( .INP(n15188), .ZN(n15186) );
  NAND2X0 U15941 ( .IN1(n7639), .IN2(WX11199), .QN(n15188) );
  NAND2X0 U15942 ( .IN1(n9101), .IN2(n8252), .QN(n15180) );
  NAND2X0 U15943 ( .IN1(n1946), .IN2(n9287), .QN(n15174) );
  NOR2X0 U15944 ( .IN1(n9229), .IN2(n9052), .QN(n1946) );
  NAND2X0 U15945 ( .IN1(DATA_0_22), .IN2(n9334), .QN(n15173) );
  NAND2X0 U15946 ( .IN1(n9301), .IN2(CRC_OUT_1_22), .QN(n15172) );
  NAND4X0 U15947 ( .IN1(n15189), .IN2(n15190), .IN3(n15191), .IN4(n15192), 
        .QN(WX11004) );
  NAND2X0 U15948 ( .IN1(n9878), .IN2(n9111), .QN(n15192) );
  NOR2X0 U15949 ( .IN1(n15193), .IN2(n15194), .QN(n9878) );
  INVX0 U15950 ( .INP(n15195), .ZN(n15194) );
  NAND2X0 U15951 ( .IN1(n15196), .IN2(n15197), .QN(n15195) );
  NOR2X0 U15952 ( .IN1(n15197), .IN2(n15196), .QN(n15193) );
  NAND2X0 U15953 ( .IN1(n15198), .IN2(n15199), .QN(n15196) );
  NAND2X0 U15954 ( .IN1(n8141), .IN2(n15200), .QN(n15199) );
  INVX0 U15955 ( .INP(n15201), .ZN(n15200) );
  NAND2X0 U15956 ( .IN1(n15201), .IN2(WX11197), .QN(n15198) );
  NAND2X0 U15957 ( .IN1(n15202), .IN2(n15203), .QN(n15201) );
  INVX0 U15958 ( .INP(n15204), .ZN(n15203) );
  NOR2X0 U15959 ( .IN1(n8818), .IN2(n16140), .QN(n15204) );
  NAND2X0 U15960 ( .IN1(n16140), .IN2(n8818), .QN(n15202) );
  NOR2X0 U15961 ( .IN1(n15205), .IN2(n15206), .QN(n15197) );
  INVX0 U15962 ( .INP(n15207), .ZN(n15206) );
  NAND2X0 U15963 ( .IN1(n7640), .IN2(n9122), .QN(n15207) );
  NOR2X0 U15964 ( .IN1(n9116), .IN2(n7640), .QN(n15205) );
  NAND2X0 U15965 ( .IN1(n1945), .IN2(n9288), .QN(n15191) );
  NOR2X0 U15966 ( .IN1(n9229), .IN2(n9053), .QN(n1945) );
  NAND2X0 U15967 ( .IN1(DATA_0_23), .IN2(n9334), .QN(n15190) );
  NAND2X0 U15968 ( .IN1(n9301), .IN2(CRC_OUT_1_23), .QN(n15189) );
  NAND4X0 U15969 ( .IN1(n15208), .IN2(n15209), .IN3(n15210), .IN4(n15211), 
        .QN(WX11002) );
  NAND2X0 U15970 ( .IN1(n15212), .IN2(n9889), .QN(n15211) );
  NAND2X0 U15971 ( .IN1(n15213), .IN2(n9893), .QN(n9889) );
  NAND2X0 U15972 ( .IN1(n15214), .IN2(n15215), .QN(n15213) );
  NAND2X0 U15973 ( .IN1(n16139), .IN2(n9122), .QN(n15215) );
  NAND2X0 U15974 ( .IN1(TM1), .IN2(n8254), .QN(n15214) );
  NAND2X0 U15975 ( .IN1(n15216), .IN2(n15217), .QN(n15212) );
  NAND2X0 U15976 ( .IN1(n9101), .IN2(n9893), .QN(n15217) );
  NAND2X0 U15977 ( .IN1(n15218), .IN2(n15219), .QN(n9893) );
  NAND2X0 U15978 ( .IN1(n7641), .IN2(n15220), .QN(n15219) );
  INVX0 U15979 ( .INP(n15221), .ZN(n15218) );
  NOR2X0 U15980 ( .IN1(n15220), .IN2(n7641), .QN(n15221) );
  NOR2X0 U15981 ( .IN1(n15222), .IN2(n15223), .QN(n15220) );
  NOR2X0 U15982 ( .IN1(WX11195), .IN2(n7642), .QN(n15223) );
  INVX0 U15983 ( .INP(n15224), .ZN(n15222) );
  NAND2X0 U15984 ( .IN1(n7642), .IN2(WX11195), .QN(n15224) );
  NAND2X0 U15985 ( .IN1(n9101), .IN2(n8254), .QN(n15216) );
  NAND2X0 U15986 ( .IN1(n1944), .IN2(n9288), .QN(n15210) );
  NOR2X0 U15987 ( .IN1(n9229), .IN2(n9054), .QN(n1944) );
  NAND2X0 U15988 ( .IN1(DATA_0_24), .IN2(n9334), .QN(n15209) );
  NAND2X0 U15989 ( .IN1(n9302), .IN2(CRC_OUT_1_24), .QN(n15208) );
  NAND4X0 U15990 ( .IN1(n15225), .IN2(n15226), .IN3(n15227), .IN4(n15228), 
        .QN(WX11000) );
  NAND2X0 U15991 ( .IN1(n15229), .IN2(n9904), .QN(n15228) );
  NAND3X0 U15992 ( .IN1(n15230), .IN2(n15231), .IN3(n9908), .QN(n9904) );
  NAND2X0 U15993 ( .IN1(n8139), .IN2(n9122), .QN(n15231) );
  NAND2X0 U15994 ( .IN1(TM1), .IN2(WX11193), .QN(n15230) );
  NAND2X0 U15995 ( .IN1(n15232), .IN2(n15233), .QN(n15229) );
  NAND2X0 U15996 ( .IN1(n9101), .IN2(n9908), .QN(n15233) );
  NAND2X0 U15997 ( .IN1(n15234), .IN2(n15235), .QN(n9908) );
  NAND2X0 U15998 ( .IN1(n15236), .IN2(WX11129), .QN(n15235) );
  NAND2X0 U15999 ( .IN1(n15237), .IN2(n15238), .QN(n15236) );
  NAND3X0 U16000 ( .IN1(n15237), .IN2(n15238), .IN3(n7644), .QN(n15234) );
  NAND2X0 U16001 ( .IN1(test_so91), .IN2(WX11065), .QN(n15238) );
  NAND2X0 U16002 ( .IN1(n7643), .IN2(n8825), .QN(n15237) );
  NAND2X0 U16003 ( .IN1(n8139), .IN2(n9111), .QN(n15232) );
  NAND2X0 U16004 ( .IN1(n1943), .IN2(n9288), .QN(n15227) );
  NOR2X0 U16005 ( .IN1(n9229), .IN2(n9055), .QN(n1943) );
  NAND2X0 U16006 ( .IN1(DATA_0_25), .IN2(n9333), .QN(n15226) );
  NAND2X0 U16007 ( .IN1(n9302), .IN2(CRC_OUT_1_25), .QN(n15225) );
  NAND4X0 U16008 ( .IN1(n15239), .IN2(n15240), .IN3(n15241), .IN4(n15242), 
        .QN(WX10998) );
  NAND2X0 U16009 ( .IN1(n15243), .IN2(n9919), .QN(n15242) );
  NAND2X0 U16010 ( .IN1(n15244), .IN2(n9923), .QN(n9919) );
  NAND2X0 U16011 ( .IN1(n15245), .IN2(n15246), .QN(n15244) );
  NAND2X0 U16012 ( .IN1(n16138), .IN2(n9122), .QN(n15246) );
  NAND2X0 U16013 ( .IN1(TM1), .IN2(n8257), .QN(n15245) );
  NAND2X0 U16014 ( .IN1(n15247), .IN2(n15248), .QN(n15243) );
  NAND2X0 U16015 ( .IN1(n9101), .IN2(n9923), .QN(n15248) );
  NAND2X0 U16016 ( .IN1(n15249), .IN2(n15250), .QN(n9923) );
  NAND2X0 U16017 ( .IN1(n7645), .IN2(n15251), .QN(n15250) );
  INVX0 U16018 ( .INP(n15252), .ZN(n15249) );
  NOR2X0 U16019 ( .IN1(n15251), .IN2(n7645), .QN(n15252) );
  NOR2X0 U16020 ( .IN1(n15253), .IN2(n15254), .QN(n15251) );
  NOR2X0 U16021 ( .IN1(WX11191), .IN2(n7646), .QN(n15254) );
  INVX0 U16022 ( .INP(n15255), .ZN(n15253) );
  NAND2X0 U16023 ( .IN1(n7646), .IN2(WX11191), .QN(n15255) );
  NAND2X0 U16024 ( .IN1(n9101), .IN2(n8257), .QN(n15247) );
  NAND2X0 U16025 ( .IN1(n1942), .IN2(n9288), .QN(n15241) );
  NOR2X0 U16026 ( .IN1(n9229), .IN2(n9056), .QN(n1942) );
  NAND2X0 U16027 ( .IN1(DATA_0_26), .IN2(n9333), .QN(n15240) );
  NAND2X0 U16028 ( .IN1(n9302), .IN2(CRC_OUT_1_26), .QN(n15239) );
  NAND4X0 U16029 ( .IN1(n15256), .IN2(n15257), .IN3(n15258), .IN4(n15259), 
        .QN(WX10996) );
  NAND2X0 U16030 ( .IN1(n15260), .IN2(n9934), .QN(n15259) );
  NAND2X0 U16031 ( .IN1(n15261), .IN2(n9938), .QN(n9934) );
  NAND2X0 U16032 ( .IN1(n15262), .IN2(n15263), .QN(n15261) );
  NAND2X0 U16033 ( .IN1(n16137), .IN2(n9122), .QN(n15263) );
  NAND2X0 U16034 ( .IN1(TM1), .IN2(n8258), .QN(n15262) );
  NAND2X0 U16035 ( .IN1(n15264), .IN2(n15265), .QN(n15260) );
  NAND2X0 U16036 ( .IN1(n9100), .IN2(n9938), .QN(n15265) );
  NAND2X0 U16037 ( .IN1(n15266), .IN2(n15267), .QN(n9938) );
  NAND2X0 U16038 ( .IN1(n7647), .IN2(n15268), .QN(n15267) );
  INVX0 U16039 ( .INP(n15269), .ZN(n15266) );
  NOR2X0 U16040 ( .IN1(n15268), .IN2(n7647), .QN(n15269) );
  NOR2X0 U16041 ( .IN1(n15270), .IN2(n15271), .QN(n15268) );
  NOR2X0 U16042 ( .IN1(WX11189), .IN2(n7648), .QN(n15271) );
  INVX0 U16043 ( .INP(n15272), .ZN(n15270) );
  NAND2X0 U16044 ( .IN1(n7648), .IN2(WX11189), .QN(n15272) );
  NAND2X0 U16045 ( .IN1(n9100), .IN2(n8258), .QN(n15264) );
  NAND2X0 U16046 ( .IN1(n1941), .IN2(n9288), .QN(n15258) );
  NOR2X0 U16047 ( .IN1(n9075), .IN2(n9155), .QN(n1941) );
  NAND2X0 U16048 ( .IN1(DATA_0_27), .IN2(n9334), .QN(n15257) );
  NAND2X0 U16049 ( .IN1(n9302), .IN2(CRC_OUT_1_27), .QN(n15256) );
  NAND4X0 U16050 ( .IN1(n15273), .IN2(n15274), .IN3(n15275), .IN4(n15276), 
        .QN(WX10994) );
  NAND2X0 U16051 ( .IN1(n15277), .IN2(n9949), .QN(n15276) );
  NAND2X0 U16052 ( .IN1(n15278), .IN2(n9953), .QN(n9949) );
  NAND2X0 U16053 ( .IN1(n15279), .IN2(n15280), .QN(n15278) );
  NAND2X0 U16054 ( .IN1(n16136), .IN2(n9122), .QN(n15280) );
  NAND2X0 U16055 ( .IN1(TM1), .IN2(n8259), .QN(n15279) );
  NAND2X0 U16056 ( .IN1(n15281), .IN2(n15282), .QN(n15277) );
  NAND2X0 U16057 ( .IN1(n9100), .IN2(n9953), .QN(n15282) );
  NAND2X0 U16058 ( .IN1(n15283), .IN2(n15284), .QN(n9953) );
  NAND2X0 U16059 ( .IN1(n7649), .IN2(n15285), .QN(n15284) );
  INVX0 U16060 ( .INP(n15286), .ZN(n15283) );
  NOR2X0 U16061 ( .IN1(n15285), .IN2(n7649), .QN(n15286) );
  NOR2X0 U16062 ( .IN1(n15287), .IN2(n15288), .QN(n15285) );
  NOR2X0 U16063 ( .IN1(WX11187), .IN2(n7650), .QN(n15288) );
  INVX0 U16064 ( .INP(n15289), .ZN(n15287) );
  NAND2X0 U16065 ( .IN1(n7650), .IN2(WX11187), .QN(n15289) );
  NAND2X0 U16066 ( .IN1(n9100), .IN2(n8259), .QN(n15281) );
  NAND2X0 U16067 ( .IN1(n1940), .IN2(n9288), .QN(n15275) );
  NOR2X0 U16068 ( .IN1(n9229), .IN2(n9057), .QN(n1940) );
  NAND2X0 U16069 ( .IN1(DATA_0_28), .IN2(n9333), .QN(n15274) );
  NAND2X0 U16070 ( .IN1(n9302), .IN2(CRC_OUT_1_28), .QN(n15273) );
  NAND4X0 U16071 ( .IN1(n15290), .IN2(n15291), .IN3(n15292), .IN4(n15293), 
        .QN(WX10992) );
  NAND2X0 U16072 ( .IN1(n15294), .IN2(n9964), .QN(n15293) );
  NAND2X0 U16073 ( .IN1(n15295), .IN2(n9968), .QN(n9964) );
  NAND2X0 U16074 ( .IN1(n15296), .IN2(n15297), .QN(n15295) );
  NAND2X0 U16075 ( .IN1(n16135), .IN2(n9122), .QN(n15297) );
  NAND2X0 U16076 ( .IN1(TM1), .IN2(n8260), .QN(n15296) );
  NAND2X0 U16077 ( .IN1(n15298), .IN2(n15299), .QN(n15294) );
  NAND2X0 U16078 ( .IN1(n9100), .IN2(n9968), .QN(n15299) );
  NAND2X0 U16079 ( .IN1(n15300), .IN2(n15301), .QN(n9968) );
  NAND2X0 U16080 ( .IN1(n7651), .IN2(n15302), .QN(n15301) );
  INVX0 U16081 ( .INP(n15303), .ZN(n15300) );
  NOR2X0 U16082 ( .IN1(n15302), .IN2(n7651), .QN(n15303) );
  NOR2X0 U16083 ( .IN1(n15304), .IN2(n15305), .QN(n15302) );
  NOR2X0 U16084 ( .IN1(WX11185), .IN2(n7652), .QN(n15305) );
  INVX0 U16085 ( .INP(n15306), .ZN(n15304) );
  NAND2X0 U16086 ( .IN1(n7652), .IN2(WX11185), .QN(n15306) );
  NAND2X0 U16087 ( .IN1(n9100), .IN2(n8260), .QN(n15298) );
  NAND2X0 U16088 ( .IN1(n1939), .IN2(n9288), .QN(n15292) );
  NOR2X0 U16089 ( .IN1(n9229), .IN2(n9058), .QN(n1939) );
  NAND2X0 U16090 ( .IN1(DATA_0_29), .IN2(n9333), .QN(n15291) );
  NAND2X0 U16091 ( .IN1(n9302), .IN2(CRC_OUT_1_29), .QN(n15290) );
  NAND4X0 U16092 ( .IN1(n15307), .IN2(n15308), .IN3(n15309), .IN4(n15310), 
        .QN(WX10990) );
  NAND2X0 U16093 ( .IN1(n15311), .IN2(n9979), .QN(n15310) );
  NAND2X0 U16094 ( .IN1(n15312), .IN2(n9983), .QN(n9979) );
  NAND2X0 U16095 ( .IN1(n15313), .IN2(n15314), .QN(n15312) );
  NAND2X0 U16096 ( .IN1(n16134), .IN2(n9122), .QN(n15314) );
  NAND2X0 U16097 ( .IN1(TM1), .IN2(n8261), .QN(n15313) );
  NAND2X0 U16098 ( .IN1(n15315), .IN2(n15316), .QN(n15311) );
  NAND2X0 U16099 ( .IN1(n9100), .IN2(n9983), .QN(n15316) );
  NAND2X0 U16100 ( .IN1(n15317), .IN2(n15318), .QN(n9983) );
  NAND2X0 U16101 ( .IN1(n7653), .IN2(n15319), .QN(n15318) );
  INVX0 U16102 ( .INP(n15320), .ZN(n15317) );
  NOR2X0 U16103 ( .IN1(n15319), .IN2(n7653), .QN(n15320) );
  NOR2X0 U16104 ( .IN1(n15321), .IN2(n15322), .QN(n15319) );
  NOR2X0 U16105 ( .IN1(WX11183), .IN2(n7654), .QN(n15322) );
  INVX0 U16106 ( .INP(n15323), .ZN(n15321) );
  NAND2X0 U16107 ( .IN1(n7654), .IN2(WX11183), .QN(n15323) );
  NAND2X0 U16108 ( .IN1(n9100), .IN2(n8261), .QN(n15315) );
  NAND2X0 U16109 ( .IN1(n1938), .IN2(n9288), .QN(n15309) );
  NOR2X0 U16110 ( .IN1(n9116), .IN2(n2182), .QN(n2148) );
  NOR2X0 U16111 ( .IN1(n9229), .IN2(n9059), .QN(n1938) );
  NAND2X0 U16112 ( .IN1(DATA_0_30), .IN2(n9333), .QN(n15308) );
  NAND2X0 U16113 ( .IN1(n9302), .IN2(CRC_OUT_1_30), .QN(n15307) );
  NAND4X0 U16114 ( .IN1(n15324), .IN2(n15325), .IN3(n15326), .IN4(n15327), 
        .QN(WX10988) );
  NAND2X0 U16115 ( .IN1(n15328), .IN2(n9989), .QN(n15327) );
  NAND2X0 U16116 ( .IN1(n15329), .IN2(n9993), .QN(n9989) );
  NAND2X0 U16117 ( .IN1(n15330), .IN2(n15331), .QN(n15329) );
  NAND2X0 U16118 ( .IN1(n16133), .IN2(n9122), .QN(n15331) );
  NAND2X0 U16119 ( .IN1(TM1), .IN2(n8262), .QN(n15330) );
  NAND2X0 U16120 ( .IN1(n15332), .IN2(n15333), .QN(n15328) );
  NAND2X0 U16121 ( .IN1(n9101), .IN2(n9993), .QN(n15333) );
  NAND2X0 U16122 ( .IN1(n15334), .IN2(n15335), .QN(n9993) );
  NAND2X0 U16123 ( .IN1(n7611), .IN2(n15336), .QN(n15335) );
  INVX0 U16124 ( .INP(n15337), .ZN(n15334) );
  NOR2X0 U16125 ( .IN1(n15336), .IN2(n7611), .QN(n15337) );
  NOR2X0 U16126 ( .IN1(n15338), .IN2(n15339), .QN(n15336) );
  NOR2X0 U16127 ( .IN1(WX11181), .IN2(n7612), .QN(n15339) );
  INVX0 U16128 ( .INP(n15340), .ZN(n15338) );
  NAND2X0 U16129 ( .IN1(n7612), .IN2(WX11181), .QN(n15340) );
  NAND2X0 U16130 ( .IN1(n9091), .IN2(n8262), .QN(n15332) );
  NOR3X0 U16131 ( .IN1(n9151), .IN2(TM0), .IN3(n9115), .QN(n9680) );
  NAND2X0 U16132 ( .IN1(DATA_0_31), .IN2(n2153), .QN(n15326) );
  NAND2X0 U16133 ( .IN1(test_so100), .IN2(n9314), .QN(n15325) );
  NAND2X0 U16134 ( .IN1(n2245), .IN2(WX10829), .QN(n15324) );
  NOR2X0 U16135 ( .IN1(n9229), .IN2(WX10829), .QN(WX10890) );
  NOR2X0 U16136 ( .IN1(n9229), .IN2(n15341), .QN(WX10377) );
  NOR2X0 U16137 ( .IN1(n15342), .IN2(n15343), .QN(n15341) );
  NOR2X0 U16138 ( .IN1(test_so85), .IN2(CRC_OUT_2_30), .QN(n15343) );
  NOR2X0 U16139 ( .IN1(DFF_1534_n1), .IN2(n8804), .QN(n15342) );
  NOR3X0 U16140 ( .IN1(n9151), .IN2(n15344), .IN3(n15345), .QN(WX10375) );
  NOR2X0 U16141 ( .IN1(n8159), .IN2(CRC_OUT_2_29), .QN(n15345) );
  NOR2X0 U16142 ( .IN1(DFF_1533_n1), .IN2(WX9890), .QN(n15344) );
  NOR3X0 U16143 ( .IN1(n9151), .IN2(n15346), .IN3(n15347), .QN(WX10373) );
  NOR2X0 U16144 ( .IN1(n8160), .IN2(CRC_OUT_2_28), .QN(n15347) );
  NOR2X0 U16145 ( .IN1(DFF_1532_n1), .IN2(WX9892), .QN(n15346) );
  NOR3X0 U16146 ( .IN1(n9151), .IN2(n15348), .IN3(n15349), .QN(WX10371) );
  NOR2X0 U16147 ( .IN1(n8161), .IN2(CRC_OUT_2_27), .QN(n15349) );
  NOR2X0 U16148 ( .IN1(DFF_1531_n1), .IN2(WX9894), .QN(n15348) );
  NOR3X0 U16149 ( .IN1(n9151), .IN2(n15350), .IN3(n15351), .QN(WX10369) );
  NOR2X0 U16150 ( .IN1(n8162), .IN2(CRC_OUT_2_26), .QN(n15351) );
  NOR2X0 U16151 ( .IN1(DFF_1530_n1), .IN2(WX9896), .QN(n15350) );
  NOR3X0 U16152 ( .IN1(n9151), .IN2(n15352), .IN3(n15353), .QN(WX10367) );
  NOR2X0 U16153 ( .IN1(n8163), .IN2(CRC_OUT_2_25), .QN(n15353) );
  NOR2X0 U16154 ( .IN1(DFF_1529_n1), .IN2(WX9898), .QN(n15352) );
  NOR3X0 U16155 ( .IN1(n9151), .IN2(n15354), .IN3(n15355), .QN(WX10365) );
  NOR2X0 U16156 ( .IN1(n8164), .IN2(CRC_OUT_2_24), .QN(n15355) );
  NOR2X0 U16157 ( .IN1(DFF_1528_n1), .IN2(WX9900), .QN(n15354) );
  NOR3X0 U16158 ( .IN1(n9151), .IN2(n15356), .IN3(n15357), .QN(WX10363) );
  NOR2X0 U16159 ( .IN1(n8165), .IN2(CRC_OUT_2_23), .QN(n15357) );
  NOR2X0 U16160 ( .IN1(DFF_1527_n1), .IN2(WX9902), .QN(n15356) );
  NOR3X0 U16161 ( .IN1(n9151), .IN2(n15358), .IN3(n15359), .QN(WX10361) );
  NOR2X0 U16162 ( .IN1(n8166), .IN2(CRC_OUT_2_22), .QN(n15359) );
  NOR2X0 U16163 ( .IN1(DFF_1526_n1), .IN2(WX9904), .QN(n15358) );
  NOR3X0 U16164 ( .IN1(n9151), .IN2(n15360), .IN3(n15361), .QN(WX10359) );
  NOR2X0 U16165 ( .IN1(n8167), .IN2(CRC_OUT_2_21), .QN(n15361) );
  NOR2X0 U16166 ( .IN1(DFF_1525_n1), .IN2(WX9906), .QN(n15360) );
  NOR3X0 U16167 ( .IN1(n9152), .IN2(n15362), .IN3(n15363), .QN(WX10357) );
  NOR2X0 U16168 ( .IN1(n8168), .IN2(CRC_OUT_2_20), .QN(n15363) );
  NOR2X0 U16169 ( .IN1(DFF_1524_n1), .IN2(WX9908), .QN(n15362) );
  NOR2X0 U16170 ( .IN1(n9230), .IN2(n15364), .QN(WX10355) );
  NOR2X0 U16171 ( .IN1(n15365), .IN2(n15366), .QN(n15364) );
  NOR2X0 U16172 ( .IN1(test_so88), .IN2(WX9910), .QN(n15366) );
  INVX0 U16173 ( .INP(n15367), .ZN(n15365) );
  NAND2X0 U16174 ( .IN1(WX9910), .IN2(test_so88), .QN(n15367) );
  NOR3X0 U16175 ( .IN1(n9152), .IN2(n15368), .IN3(n15369), .QN(WX10353) );
  NOR2X0 U16176 ( .IN1(n8170), .IN2(CRC_OUT_2_18), .QN(n15369) );
  NOR2X0 U16177 ( .IN1(DFF_1522_n1), .IN2(WX9912), .QN(n15368) );
  NOR3X0 U16178 ( .IN1(n9152), .IN2(n15370), .IN3(n15371), .QN(WX10351) );
  NOR2X0 U16179 ( .IN1(n8171), .IN2(CRC_OUT_2_17), .QN(n15371) );
  NOR2X0 U16180 ( .IN1(DFF_1521_n1), .IN2(WX9914), .QN(n15370) );
  NOR3X0 U16181 ( .IN1(n9152), .IN2(n15372), .IN3(n15373), .QN(WX10349) );
  NOR2X0 U16182 ( .IN1(n8172), .IN2(CRC_OUT_2_16), .QN(n15373) );
  NOR2X0 U16183 ( .IN1(DFF_1520_n1), .IN2(WX9916), .QN(n15372) );
  NOR2X0 U16184 ( .IN1(n9230), .IN2(n15374), .QN(WX10347) );
  NOR2X0 U16185 ( .IN1(n15375), .IN2(n15376), .QN(n15374) );
  NOR2X0 U16186 ( .IN1(DFF_1519_n1), .IN2(n15377), .QN(n15376) );
  INVX0 U16187 ( .INP(n15378), .ZN(n15375) );
  NAND2X0 U16188 ( .IN1(n15377), .IN2(DFF_1519_n1), .QN(n15378) );
  NOR2X0 U16189 ( .IN1(n15379), .IN2(n15380), .QN(n15377) );
  NOR2X0 U16190 ( .IN1(WX9918), .IN2(DFF_1535_n1), .QN(n15380) );
  NOR2X0 U16191 ( .IN1(CRC_OUT_2_31), .IN2(n8107), .QN(n15379) );
  NOR3X0 U16192 ( .IN1(n9152), .IN2(n15381), .IN3(n15382), .QN(WX10345) );
  NOR2X0 U16193 ( .IN1(n8173), .IN2(CRC_OUT_2_14), .QN(n15382) );
  NOR2X0 U16194 ( .IN1(DFF_1518_n1), .IN2(WX9920), .QN(n15381) );
  NOR2X0 U16195 ( .IN1(n9230), .IN2(n15383), .QN(WX10343) );
  NOR2X0 U16196 ( .IN1(n15384), .IN2(n15385), .QN(n15383) );
  NOR2X0 U16197 ( .IN1(test_so86), .IN2(CRC_OUT_2_13), .QN(n15385) );
  NOR2X0 U16198 ( .IN1(DFF_1517_n1), .IN2(n8794), .QN(n15384) );
  NOR3X0 U16199 ( .IN1(n9152), .IN2(n15386), .IN3(n15387), .QN(WX10341) );
  NOR2X0 U16200 ( .IN1(n8174), .IN2(CRC_OUT_2_12), .QN(n15387) );
  NOR2X0 U16201 ( .IN1(DFF_1516_n1), .IN2(WX9924), .QN(n15386) );
  NOR3X0 U16202 ( .IN1(n9152), .IN2(n15388), .IN3(n15389), .QN(WX10339) );
  NOR2X0 U16203 ( .IN1(n8175), .IN2(CRC_OUT_2_11), .QN(n15389) );
  NOR2X0 U16204 ( .IN1(DFF_1515_n1), .IN2(WX9926), .QN(n15388) );
  NOR2X0 U16205 ( .IN1(n9230), .IN2(n15390), .QN(WX10337) );
  NOR2X0 U16206 ( .IN1(n15391), .IN2(n15392), .QN(n15390) );
  INVX0 U16207 ( .INP(n15393), .ZN(n15392) );
  NAND2X0 U16208 ( .IN1(CRC_OUT_2_10), .IN2(n15394), .QN(n15393) );
  NOR2X0 U16209 ( .IN1(n15394), .IN2(CRC_OUT_2_10), .QN(n15391) );
  NAND2X0 U16210 ( .IN1(n15395), .IN2(n15396), .QN(n15394) );
  NAND2X0 U16211 ( .IN1(n8108), .IN2(CRC_OUT_2_31), .QN(n15396) );
  NAND2X0 U16212 ( .IN1(DFF_1535_n1), .IN2(WX9928), .QN(n15395) );
  NOR3X0 U16213 ( .IN1(n9152), .IN2(n15397), .IN3(n15398), .QN(WX10335) );
  NOR2X0 U16214 ( .IN1(n8176), .IN2(CRC_OUT_2_9), .QN(n15398) );
  NOR2X0 U16215 ( .IN1(DFF_1513_n1), .IN2(WX9930), .QN(n15397) );
  NOR3X0 U16216 ( .IN1(n9152), .IN2(n15399), .IN3(n15400), .QN(WX10333) );
  NOR2X0 U16217 ( .IN1(n8177), .IN2(CRC_OUT_2_8), .QN(n15400) );
  NOR2X0 U16218 ( .IN1(DFF_1512_n1), .IN2(WX9932), .QN(n15399) );
  NOR3X0 U16219 ( .IN1(n9153), .IN2(n15401), .IN3(n15402), .QN(WX10331) );
  NOR2X0 U16220 ( .IN1(n8178), .IN2(CRC_OUT_2_7), .QN(n15402) );
  NOR2X0 U16221 ( .IN1(DFF_1511_n1), .IN2(WX9934), .QN(n15401) );
  NOR3X0 U16222 ( .IN1(n9153), .IN2(n15403), .IN3(n15404), .QN(WX10329) );
  NOR2X0 U16223 ( .IN1(n8179), .IN2(CRC_OUT_2_6), .QN(n15404) );
  NOR2X0 U16224 ( .IN1(DFF_1510_n1), .IN2(WX9936), .QN(n15403) );
  NOR3X0 U16225 ( .IN1(n9152), .IN2(n15405), .IN3(n15406), .QN(WX10327) );
  NOR2X0 U16226 ( .IN1(n8180), .IN2(CRC_OUT_2_5), .QN(n15406) );
  NOR2X0 U16227 ( .IN1(DFF_1509_n1), .IN2(WX9938), .QN(n15405) );
  NOR3X0 U16228 ( .IN1(n9153), .IN2(n15407), .IN3(n15408), .QN(WX10325) );
  NOR2X0 U16229 ( .IN1(n8181), .IN2(CRC_OUT_2_4), .QN(n15408) );
  NOR2X0 U16230 ( .IN1(DFF_1508_n1), .IN2(WX9940), .QN(n15407) );
  NOR2X0 U16231 ( .IN1(n9231), .IN2(n15409), .QN(WX10323) );
  NOR2X0 U16232 ( .IN1(n15410), .IN2(n15411), .QN(n15409) );
  INVX0 U16233 ( .INP(n15412), .ZN(n15411) );
  NAND2X0 U16234 ( .IN1(CRC_OUT_2_3), .IN2(n15413), .QN(n15412) );
  NOR2X0 U16235 ( .IN1(n15413), .IN2(CRC_OUT_2_3), .QN(n15410) );
  NAND2X0 U16236 ( .IN1(n15414), .IN2(n15415), .QN(n15413) );
  NAND2X0 U16237 ( .IN1(n8109), .IN2(CRC_OUT_2_31), .QN(n15415) );
  NAND2X0 U16238 ( .IN1(DFF_1535_n1), .IN2(WX9942), .QN(n15414) );
  NOR2X0 U16239 ( .IN1(n9231), .IN2(n15416), .QN(WX10321) );
  NOR2X0 U16240 ( .IN1(n15417), .IN2(n15418), .QN(n15416) );
  NOR2X0 U16241 ( .IN1(test_so87), .IN2(WX9944), .QN(n15418) );
  INVX0 U16242 ( .INP(n15419), .ZN(n15417) );
  NAND2X0 U16243 ( .IN1(WX9944), .IN2(test_so87), .QN(n15419) );
  NOR3X0 U16244 ( .IN1(n9153), .IN2(n15420), .IN3(n15421), .QN(WX10319) );
  NOR2X0 U16245 ( .IN1(n8183), .IN2(CRC_OUT_2_1), .QN(n15421) );
  NOR2X0 U16246 ( .IN1(DFF_1505_n1), .IN2(WX9946), .QN(n15420) );
  NOR3X0 U16247 ( .IN1(n9153), .IN2(n15422), .IN3(n15423), .QN(WX10317) );
  NOR2X0 U16248 ( .IN1(n8184), .IN2(CRC_OUT_2_0), .QN(n15423) );
  NOR2X0 U16249 ( .IN1(DFF_1504_n1), .IN2(WX9948), .QN(n15422) );
  NOR3X0 U16250 ( .IN1(n9135), .IN2(n15424), .IN3(n15425), .QN(WX10315) );
  NOR2X0 U16251 ( .IN1(n8126), .IN2(CRC_OUT_2_31), .QN(n15425) );
  NOR2X0 U16252 ( .IN1(DFF_1535_n1), .IN2(WX9950), .QN(n15424) );
  INVX0 U16253 ( .INP(RESET), .ZN(n2181) );
  NAND2X0 U16254 ( .IN1(n15426), .IN2(n15427), .QN(DATA_9_9) );
  INVX0 U16255 ( .INP(n15428), .ZN(n15427) );
  NOR2X0 U16256 ( .IN1(n15429), .IN2(n11437), .QN(n15428) );
  NAND2X0 U16257 ( .IN1(n11437), .IN2(n15429), .QN(n15426) );
  NAND2X0 U16258 ( .IN1(TM0), .IN2(WX529), .QN(n15429) );
  NAND2X0 U16259 ( .IN1(n15430), .IN2(n15431), .QN(n11437) );
  NAND2X0 U16260 ( .IN1(n15432), .IN2(n15433), .QN(n15431) );
  INVX0 U16261 ( .INP(n15434), .ZN(n15430) );
  NOR2X0 U16262 ( .IN1(n15433), .IN2(n15432), .QN(n15434) );
  NAND2X0 U16263 ( .IN1(n15435), .IN2(n15436), .QN(n15432) );
  NAND2X0 U16264 ( .IN1(n8740), .IN2(n15437), .QN(n15436) );
  INVX0 U16265 ( .INP(n15438), .ZN(n15435) );
  NOR2X0 U16266 ( .IN1(n15437), .IN2(n8740), .QN(n15438) );
  NOR2X0 U16267 ( .IN1(n15439), .IN2(n15440), .QN(n15437) );
  NOR2X0 U16268 ( .IN1(WX881), .IN2(n8741), .QN(n15440) );
  INVX0 U16269 ( .INP(n15441), .ZN(n15439) );
  NAND2X0 U16270 ( .IN1(n8741), .IN2(WX881), .QN(n15441) );
  NOR2X0 U16271 ( .IN1(n15442), .IN2(n15443), .QN(n15433) );
  INVX0 U16272 ( .INP(n15444), .ZN(n15443) );
  NAND2X0 U16273 ( .IN1(n3485), .IN2(n2182), .QN(n15444) );
  NOR2X0 U16274 ( .IN1(n2182), .IN2(n3485), .QN(n15442) );
  NAND2X0 U16275 ( .IN1(n15445), .IN2(n15446), .QN(DATA_9_8) );
  INVX0 U16276 ( .INP(n15447), .ZN(n15446) );
  NOR2X0 U16277 ( .IN1(n15448), .IN2(n11431), .QN(n15447) );
  NAND2X0 U16278 ( .IN1(n11431), .IN2(n15448), .QN(n15445) );
  NAND2X0 U16279 ( .IN1(TM0), .IN2(WX531), .QN(n15448) );
  NAND2X0 U16280 ( .IN1(n15449), .IN2(n15450), .QN(n11431) );
  NAND2X0 U16281 ( .IN1(n15451), .IN2(n15452), .QN(n15450) );
  INVX0 U16282 ( .INP(n15453), .ZN(n15449) );
  NOR2X0 U16283 ( .IN1(n15452), .IN2(n15451), .QN(n15453) );
  NAND2X0 U16284 ( .IN1(n15454), .IN2(n15455), .QN(n15451) );
  NAND2X0 U16285 ( .IN1(n8750), .IN2(n15456), .QN(n15455) );
  INVX0 U16286 ( .INP(n15457), .ZN(n15454) );
  NOR2X0 U16287 ( .IN1(n15456), .IN2(n8750), .QN(n15457) );
  NOR2X0 U16288 ( .IN1(n15458), .IN2(n15459), .QN(n15456) );
  INVX0 U16289 ( .INP(n15460), .ZN(n15459) );
  NAND2X0 U16290 ( .IN1(n8752), .IN2(WX883), .QN(n15460) );
  NOR2X0 U16291 ( .IN1(WX883), .IN2(n8752), .QN(n15458) );
  NOR2X0 U16292 ( .IN1(n15461), .IN2(n15462), .QN(n15452) );
  INVX0 U16293 ( .INP(n15463), .ZN(n15462) );
  NAND2X0 U16294 ( .IN1(n3483), .IN2(n2182), .QN(n15463) );
  NOR2X0 U16295 ( .IN1(n2182), .IN2(n3483), .QN(n15461) );
  NAND2X0 U16296 ( .IN1(n15464), .IN2(n15465), .QN(DATA_9_7) );
  INVX0 U16297 ( .INP(n15466), .ZN(n15465) );
  NOR2X0 U16298 ( .IN1(n15467), .IN2(n11425), .QN(n15466) );
  NAND2X0 U16299 ( .IN1(n11425), .IN2(n15467), .QN(n15464) );
  NAND2X0 U16300 ( .IN1(TM0), .IN2(WX533), .QN(n15467) );
  NAND2X0 U16301 ( .IN1(n15468), .IN2(n15469), .QN(n11425) );
  NAND2X0 U16302 ( .IN1(n15470), .IN2(n15471), .QN(n15469) );
  INVX0 U16303 ( .INP(n15472), .ZN(n15468) );
  NOR2X0 U16304 ( .IN1(n15471), .IN2(n15470), .QN(n15472) );
  NAND2X0 U16305 ( .IN1(n15473), .IN2(n15474), .QN(n15470) );
  NAND2X0 U16306 ( .IN1(n8780), .IN2(n15475), .QN(n15474) );
  INVX0 U16307 ( .INP(n15476), .ZN(n15473) );
  NOR2X0 U16308 ( .IN1(n15475), .IN2(n8780), .QN(n15476) );
  NOR2X0 U16309 ( .IN1(n15477), .IN2(n15478), .QN(n15475) );
  NOR2X0 U16310 ( .IN1(WX885), .IN2(n8781), .QN(n15478) );
  INVX0 U16311 ( .INP(n15479), .ZN(n15477) );
  NAND2X0 U16312 ( .IN1(n8781), .IN2(WX885), .QN(n15479) );
  NOR2X0 U16313 ( .IN1(n15480), .IN2(n15481), .QN(n15471) );
  INVX0 U16314 ( .INP(n15482), .ZN(n15481) );
  NAND2X0 U16315 ( .IN1(n3481), .IN2(n2182), .QN(n15482) );
  NOR2X0 U16316 ( .IN1(n2182), .IN2(n3481), .QN(n15480) );
  NOR2X0 U16317 ( .IN1(n15483), .IN2(n15484), .QN(DATA_9_6) );
  INVX0 U16318 ( .INP(n15485), .ZN(n15484) );
  NAND2X0 U16319 ( .IN1(n15486), .IN2(n11419), .QN(n15485) );
  NOR2X0 U16320 ( .IN1(n11419), .IN2(n15486), .QN(n15483) );
  NAND2X0 U16321 ( .IN1(TM0), .IN2(WX535), .QN(n15486) );
  NAND2X0 U16322 ( .IN1(n15487), .IN2(n15488), .QN(n11419) );
  NAND2X0 U16323 ( .IN1(n15489), .IN2(n15490), .QN(n15488) );
  NAND2X0 U16324 ( .IN1(n15491), .IN2(n15492), .QN(n15489) );
  NAND3X0 U16325 ( .IN1(n15491), .IN2(n15492), .IN3(n15493), .QN(n15487) );
  INVX0 U16326 ( .INP(n15490), .ZN(n15493) );
  NOR2X0 U16327 ( .IN1(n15494), .IN2(n15495), .QN(n15490) );
  INVX0 U16328 ( .INP(n15496), .ZN(n15495) );
  NAND2X0 U16329 ( .IN1(n8768), .IN2(n15497), .QN(n15496) );
  NOR2X0 U16330 ( .IN1(n15497), .IN2(n8768), .QN(n15494) );
  NOR2X0 U16331 ( .IN1(n15498), .IN2(n15499), .QN(n15497) );
  INVX0 U16332 ( .INP(n15500), .ZN(n15499) );
  NAND2X0 U16333 ( .IN1(test_so5), .IN2(WX887), .QN(n15500) );
  NOR2X0 U16334 ( .IN1(WX887), .IN2(test_so5), .QN(n15498) );
  NAND2X0 U16335 ( .IN1(n3479), .IN2(n2182), .QN(n15492) );
  NAND2X0 U16336 ( .IN1(TM0), .IN2(WX695), .QN(n15491) );
  NAND2X0 U16337 ( .IN1(n15501), .IN2(n15502), .QN(DATA_9_5) );
  INVX0 U16338 ( .INP(n15503), .ZN(n15502) );
  NOR2X0 U16339 ( .IN1(n15504), .IN2(n11412), .QN(n15503) );
  NAND2X0 U16340 ( .IN1(n11412), .IN2(n15504), .QN(n15501) );
  NAND2X0 U16341 ( .IN1(TM0), .IN2(WX537), .QN(n15504) );
  NAND2X0 U16342 ( .IN1(n15505), .IN2(n15506), .QN(n11412) );
  NAND2X0 U16343 ( .IN1(n15507), .IN2(n15508), .QN(n15506) );
  INVX0 U16344 ( .INP(n15509), .ZN(n15505) );
  NOR2X0 U16345 ( .IN1(n15508), .IN2(n15507), .QN(n15509) );
  NAND2X0 U16346 ( .IN1(n15510), .IN2(n15511), .QN(n15507) );
  NAND2X0 U16347 ( .IN1(n8753), .IN2(n15512), .QN(n15511) );
  INVX0 U16348 ( .INP(n15513), .ZN(n15510) );
  NOR2X0 U16349 ( .IN1(n15512), .IN2(n8753), .QN(n15513) );
  NOR2X0 U16350 ( .IN1(n15514), .IN2(n15515), .QN(n15512) );
  INVX0 U16351 ( .INP(n15516), .ZN(n15515) );
  NAND2X0 U16352 ( .IN1(n8755), .IN2(WX889), .QN(n15516) );
  NOR2X0 U16353 ( .IN1(WX889), .IN2(n8755), .QN(n15514) );
  NOR2X0 U16354 ( .IN1(n15517), .IN2(n15518), .QN(n15508) );
  INVX0 U16355 ( .INP(n15519), .ZN(n15518) );
  NAND2X0 U16356 ( .IN1(n3477), .IN2(n2182), .QN(n15519) );
  NOR2X0 U16357 ( .IN1(n2182), .IN2(n3477), .QN(n15517) );
  NAND2X0 U16358 ( .IN1(n15520), .IN2(n15521), .QN(DATA_9_4) );
  INVX0 U16359 ( .INP(n15522), .ZN(n15521) );
  NOR2X0 U16360 ( .IN1(n15523), .IN2(n11406), .QN(n15522) );
  NAND2X0 U16361 ( .IN1(n11406), .IN2(n15523), .QN(n15520) );
  NAND2X0 U16362 ( .IN1(TM0), .IN2(WX539), .QN(n15523) );
  NAND2X0 U16363 ( .IN1(n15524), .IN2(n15525), .QN(n11406) );
  NAND2X0 U16364 ( .IN1(n15526), .IN2(n15527), .QN(n15525) );
  INVX0 U16365 ( .INP(n15528), .ZN(n15524) );
  NOR2X0 U16366 ( .IN1(n15527), .IN2(n15526), .QN(n15528) );
  NAND2X0 U16367 ( .IN1(n15529), .IN2(n15530), .QN(n15526) );
  NAND2X0 U16368 ( .IN1(n8756), .IN2(n15531), .QN(n15530) );
  INVX0 U16369 ( .INP(n15532), .ZN(n15529) );
  NOR2X0 U16370 ( .IN1(n15531), .IN2(n8756), .QN(n15532) );
  NOR2X0 U16371 ( .IN1(n15533), .IN2(n15534), .QN(n15531) );
  INVX0 U16372 ( .INP(n15535), .ZN(n15534) );
  NAND2X0 U16373 ( .IN1(n8758), .IN2(WX891), .QN(n15535) );
  NOR2X0 U16374 ( .IN1(WX891), .IN2(n8758), .QN(n15533) );
  NOR2X0 U16375 ( .IN1(n15536), .IN2(n15537), .QN(n15527) );
  INVX0 U16376 ( .INP(n15538), .ZN(n15537) );
  NAND2X0 U16377 ( .IN1(n3475), .IN2(n2182), .QN(n15538) );
  NOR2X0 U16378 ( .IN1(n2182), .IN2(n3475), .QN(n15536) );
  NAND2X0 U16379 ( .IN1(n15539), .IN2(n15540), .QN(DATA_9_31) );
  INVX0 U16380 ( .INP(n15541), .ZN(n15540) );
  NOR2X0 U16381 ( .IN1(n15542), .IN2(n11721), .QN(n15541) );
  NAND2X0 U16382 ( .IN1(n11721), .IN2(n15542), .QN(n15539) );
  NAND2X0 U16383 ( .IN1(TM0), .IN2(WX485), .QN(n15542) );
  NAND2X0 U16384 ( .IN1(n15543), .IN2(n15544), .QN(n11721) );
  NAND2X0 U16385 ( .IN1(n15545), .IN2(n15546), .QN(n15544) );
  INVX0 U16386 ( .INP(n15547), .ZN(n15543) );
  NOR2X0 U16387 ( .IN1(n15546), .IN2(n15545), .QN(n15547) );
  NAND2X0 U16388 ( .IN1(n15548), .IN2(n15549), .QN(n15545) );
  NAND2X0 U16389 ( .IN1(n8772), .IN2(n15550), .QN(n15549) );
  INVX0 U16390 ( .INP(n15551), .ZN(n15548) );
  NOR2X0 U16391 ( .IN1(n15550), .IN2(n8772), .QN(n15551) );
  NOR2X0 U16392 ( .IN1(n15552), .IN2(n15553), .QN(n15550) );
  NOR2X0 U16393 ( .IN1(WX837), .IN2(n8773), .QN(n15553) );
  INVX0 U16394 ( .INP(n15554), .ZN(n15552) );
  NAND2X0 U16395 ( .IN1(n8773), .IN2(WX837), .QN(n15554) );
  NOR2X0 U16396 ( .IN1(n15555), .IN2(n15556), .QN(n15546) );
  INVX0 U16397 ( .INP(n15557), .ZN(n15556) );
  NAND2X0 U16398 ( .IN1(n3529), .IN2(n9123), .QN(n15557) );
  NOR2X0 U16399 ( .IN1(n9116), .IN2(n3529), .QN(n15555) );
  NAND2X0 U16400 ( .IN1(n15558), .IN2(n15559), .QN(DATA_9_30) );
  INVX0 U16401 ( .INP(n15560), .ZN(n15559) );
  NOR2X0 U16402 ( .IN1(n15561), .IN2(n11680), .QN(n15560) );
  NAND2X0 U16403 ( .IN1(n11680), .IN2(n15561), .QN(n15558) );
  NAND2X0 U16404 ( .IN1(TM0), .IN2(WX487), .QN(n15561) );
  NAND2X0 U16405 ( .IN1(n15562), .IN2(n15563), .QN(n11680) );
  NAND2X0 U16406 ( .IN1(n15564), .IN2(n15565), .QN(n15563) );
  INVX0 U16407 ( .INP(n15566), .ZN(n15562) );
  NOR2X0 U16408 ( .IN1(n15565), .IN2(n15564), .QN(n15566) );
  NAND2X0 U16409 ( .IN1(n15567), .IN2(n15568), .QN(n15564) );
  NAND2X0 U16410 ( .IN1(n8660), .IN2(n15569), .QN(n15568) );
  INVX0 U16411 ( .INP(n15570), .ZN(n15567) );
  NOR2X0 U16412 ( .IN1(n15569), .IN2(n8660), .QN(n15570) );
  NOR2X0 U16413 ( .IN1(n15571), .IN2(n15572), .QN(n15569) );
  NOR2X0 U16414 ( .IN1(WX839), .IN2(n8678), .QN(n15572) );
  INVX0 U16415 ( .INP(n15573), .ZN(n15571) );
  NAND2X0 U16416 ( .IN1(n8678), .IN2(WX839), .QN(n15573) );
  NOR2X0 U16417 ( .IN1(n15574), .IN2(n15575), .QN(n15565) );
  INVX0 U16418 ( .INP(n15576), .ZN(n15575) );
  NAND2X0 U16419 ( .IN1(n3527), .IN2(n9123), .QN(n15576) );
  NOR2X0 U16420 ( .IN1(n9115), .IN2(n3527), .QN(n15574) );
  NAND2X0 U16421 ( .IN1(n15577), .IN2(n15578), .QN(DATA_9_3) );
  INVX0 U16422 ( .INP(n15579), .ZN(n15578) );
  NOR2X0 U16423 ( .IN1(n15580), .IN2(n11399), .QN(n15579) );
  NAND2X0 U16424 ( .IN1(n11399), .IN2(n15580), .QN(n15577) );
  NAND2X0 U16425 ( .IN1(TM0), .IN2(WX541), .QN(n15580) );
  NAND2X0 U16426 ( .IN1(n15581), .IN2(n15582), .QN(n11399) );
  NAND2X0 U16427 ( .IN1(n15583), .IN2(n15584), .QN(n15582) );
  INVX0 U16428 ( .INP(n15585), .ZN(n15581) );
  NOR2X0 U16429 ( .IN1(n15584), .IN2(n15583), .QN(n15585) );
  NAND2X0 U16430 ( .IN1(n15586), .IN2(n15587), .QN(n15583) );
  NAND2X0 U16431 ( .IN1(n8697), .IN2(n15588), .QN(n15587) );
  INVX0 U16432 ( .INP(n15589), .ZN(n15586) );
  NOR2X0 U16433 ( .IN1(n15588), .IN2(n8697), .QN(n15589) );
  NOR2X0 U16434 ( .IN1(n15590), .IN2(n15591), .QN(n15588) );
  INVX0 U16435 ( .INP(n15592), .ZN(n15591) );
  NAND2X0 U16436 ( .IN1(n8703), .IN2(WX893), .QN(n15592) );
  NOR2X0 U16437 ( .IN1(WX893), .IN2(n8703), .QN(n15590) );
  NOR2X0 U16438 ( .IN1(n15593), .IN2(n15594), .QN(n15584) );
  INVX0 U16439 ( .INP(n15595), .ZN(n15594) );
  NAND2X0 U16440 ( .IN1(n3473), .IN2(n2182), .QN(n15595) );
  NOR2X0 U16441 ( .IN1(n2182), .IN2(n3473), .QN(n15593) );
  NAND2X0 U16442 ( .IN1(n15596), .IN2(n15597), .QN(DATA_9_29) );
  INVX0 U16443 ( .INP(n15598), .ZN(n15597) );
  NOR2X0 U16444 ( .IN1(n15599), .IN2(n11644), .QN(n15598) );
  NAND2X0 U16445 ( .IN1(n11644), .IN2(n15599), .QN(n15596) );
  NAND2X0 U16446 ( .IN1(TM0), .IN2(WX489), .QN(n15599) );
  NAND2X0 U16447 ( .IN1(n15600), .IN2(n15601), .QN(n11644) );
  NAND2X0 U16448 ( .IN1(n15602), .IN2(n15603), .QN(n15601) );
  INVX0 U16449 ( .INP(n15604), .ZN(n15600) );
  NOR2X0 U16450 ( .IN1(n15603), .IN2(n15602), .QN(n15604) );
  NAND2X0 U16451 ( .IN1(n15605), .IN2(n15606), .QN(n15602) );
  NAND2X0 U16452 ( .IN1(n8707), .IN2(n15607), .QN(n15606) );
  INVX0 U16453 ( .INP(n15608), .ZN(n15605) );
  NOR2X0 U16454 ( .IN1(n15607), .IN2(n8707), .QN(n15608) );
  NOR2X0 U16455 ( .IN1(n15609), .IN2(n15610), .QN(n15607) );
  INVX0 U16456 ( .INP(n15611), .ZN(n15610) );
  NAND2X0 U16457 ( .IN1(n8709), .IN2(WX841), .QN(n15611) );
  NOR2X0 U16458 ( .IN1(WX841), .IN2(n8709), .QN(n15609) );
  NOR2X0 U16459 ( .IN1(n15612), .IN2(n15613), .QN(n15603) );
  INVX0 U16460 ( .INP(n15614), .ZN(n15613) );
  NAND2X0 U16461 ( .IN1(n3525), .IN2(n9123), .QN(n15614) );
  NOR2X0 U16462 ( .IN1(n9115), .IN2(n3525), .QN(n15612) );
  NOR2X0 U16463 ( .IN1(n15615), .IN2(n15616), .QN(DATA_9_28) );
  INVX0 U16464 ( .INP(n15617), .ZN(n15616) );
  NAND2X0 U16465 ( .IN1(n15618), .IN2(n11613), .QN(n15617) );
  NOR2X0 U16466 ( .IN1(n11613), .IN2(n15618), .QN(n15615) );
  NAND2X0 U16467 ( .IN1(TM0), .IN2(WX491), .QN(n15618) );
  NAND2X0 U16468 ( .IN1(n15619), .IN2(n15620), .QN(n11613) );
  NAND2X0 U16469 ( .IN1(n15621), .IN2(n15622), .QN(n15620) );
  NAND2X0 U16470 ( .IN1(n15623), .IN2(n15624), .QN(n15621) );
  NAND3X0 U16471 ( .IN1(n15623), .IN2(n15624), .IN3(n15625), .QN(n15619) );
  INVX0 U16472 ( .INP(n15622), .ZN(n15625) );
  NOR2X0 U16473 ( .IN1(n15626), .IN2(n15627), .QN(n15622) );
  INVX0 U16474 ( .INP(n15628), .ZN(n15627) );
  NAND2X0 U16475 ( .IN1(n8716), .IN2(n15629), .QN(n15628) );
  NOR2X0 U16476 ( .IN1(n15629), .IN2(n8716), .QN(n15626) );
  NOR2X0 U16477 ( .IN1(n15630), .IN2(n15631), .QN(n15629) );
  INVX0 U16478 ( .INP(n15632), .ZN(n15631) );
  NAND2X0 U16479 ( .IN1(test_so2), .IN2(WX843), .QN(n15632) );
  NOR2X0 U16480 ( .IN1(WX843), .IN2(test_so2), .QN(n15630) );
  NAND2X0 U16481 ( .IN1(n8718), .IN2(n9123), .QN(n15624) );
  NAND2X0 U16482 ( .IN1(TM1), .IN2(WX715), .QN(n15623) );
  NAND2X0 U16483 ( .IN1(n15633), .IN2(n15634), .QN(DATA_9_27) );
  INVX0 U16484 ( .INP(n15635), .ZN(n15634) );
  NOR2X0 U16485 ( .IN1(n15636), .IN2(n11606), .QN(n15635) );
  NAND2X0 U16486 ( .IN1(n11606), .IN2(n15636), .QN(n15633) );
  NAND2X0 U16487 ( .IN1(TM0), .IN2(WX493), .QN(n15636) );
  NAND2X0 U16488 ( .IN1(n15637), .IN2(n15638), .QN(n11606) );
  NAND2X0 U16489 ( .IN1(n15639), .IN2(n15640), .QN(n15638) );
  INVX0 U16490 ( .INP(n15641), .ZN(n15637) );
  NOR2X0 U16491 ( .IN1(n15640), .IN2(n15639), .QN(n15641) );
  NAND2X0 U16492 ( .IN1(n15642), .IN2(n15643), .QN(n15639) );
  NAND2X0 U16493 ( .IN1(n8722), .IN2(n15644), .QN(n15643) );
  INVX0 U16494 ( .INP(n15645), .ZN(n15642) );
  NOR2X0 U16495 ( .IN1(n15644), .IN2(n8722), .QN(n15645) );
  NOR2X0 U16496 ( .IN1(n15646), .IN2(n15647), .QN(n15644) );
  INVX0 U16497 ( .INP(n15648), .ZN(n15647) );
  NAND2X0 U16498 ( .IN1(n8724), .IN2(WX845), .QN(n15648) );
  NOR2X0 U16499 ( .IN1(WX845), .IN2(n8724), .QN(n15646) );
  NOR2X0 U16500 ( .IN1(n15649), .IN2(n15650), .QN(n15640) );
  INVX0 U16501 ( .INP(n15651), .ZN(n15650) );
  NAND2X0 U16502 ( .IN1(n3521), .IN2(n9123), .QN(n15651) );
  NOR2X0 U16503 ( .IN1(n9115), .IN2(n3521), .QN(n15649) );
  NAND2X0 U16504 ( .IN1(n15652), .IN2(n15653), .QN(DATA_9_26) );
  INVX0 U16505 ( .INP(n15654), .ZN(n15653) );
  NOR2X0 U16506 ( .IN1(n15655), .IN2(n11595), .QN(n15654) );
  NAND2X0 U16507 ( .IN1(n11595), .IN2(n15655), .QN(n15652) );
  NAND2X0 U16508 ( .IN1(TM0), .IN2(WX495), .QN(n15655) );
  NAND2X0 U16509 ( .IN1(n15656), .IN2(n15657), .QN(n11595) );
  NAND2X0 U16510 ( .IN1(n15658), .IN2(n15659), .QN(n15657) );
  INVX0 U16511 ( .INP(n15660), .ZN(n15656) );
  NOR2X0 U16512 ( .IN1(n15659), .IN2(n15658), .QN(n15660) );
  NAND2X0 U16513 ( .IN1(n15661), .IN2(n15662), .QN(n15658) );
  NAND2X0 U16514 ( .IN1(n8725), .IN2(n15663), .QN(n15662) );
  INVX0 U16515 ( .INP(n15664), .ZN(n15661) );
  NOR2X0 U16516 ( .IN1(n15663), .IN2(n8725), .QN(n15664) );
  NOR2X0 U16517 ( .IN1(n15665), .IN2(n15666), .QN(n15663) );
  INVX0 U16518 ( .INP(n15667), .ZN(n15666) );
  NAND2X0 U16519 ( .IN1(n8727), .IN2(WX847), .QN(n15667) );
  NOR2X0 U16520 ( .IN1(WX847), .IN2(n8727), .QN(n15665) );
  NOR2X0 U16521 ( .IN1(n15668), .IN2(n15669), .QN(n15659) );
  INVX0 U16522 ( .INP(n15670), .ZN(n15669) );
  NAND2X0 U16523 ( .IN1(n3519), .IN2(n9123), .QN(n15670) );
  NOR2X0 U16524 ( .IN1(n9116), .IN2(n3519), .QN(n15668) );
  NAND2X0 U16525 ( .IN1(n15671), .IN2(n15672), .QN(DATA_9_25) );
  INVX0 U16526 ( .INP(n15673), .ZN(n15672) );
  NOR2X0 U16527 ( .IN1(n15674), .IN2(n11584), .QN(n15673) );
  NAND2X0 U16528 ( .IN1(n11584), .IN2(n15674), .QN(n15671) );
  NAND2X0 U16529 ( .IN1(TM0), .IN2(WX497), .QN(n15674) );
  NAND2X0 U16530 ( .IN1(n15675), .IN2(n15676), .QN(n11584) );
  NAND2X0 U16531 ( .IN1(n15677), .IN2(n15678), .QN(n15676) );
  INVX0 U16532 ( .INP(n15679), .ZN(n15675) );
  NOR2X0 U16533 ( .IN1(n15678), .IN2(n15677), .QN(n15679) );
  NAND2X0 U16534 ( .IN1(n15680), .IN2(n15681), .QN(n15677) );
  NAND2X0 U16535 ( .IN1(n8734), .IN2(n15682), .QN(n15681) );
  INVX0 U16536 ( .INP(n15683), .ZN(n15680) );
  NOR2X0 U16537 ( .IN1(n15682), .IN2(n8734), .QN(n15683) );
  NOR2X0 U16538 ( .IN1(n15684), .IN2(n15685), .QN(n15682) );
  INVX0 U16539 ( .INP(n15686), .ZN(n15685) );
  NAND2X0 U16540 ( .IN1(n8736), .IN2(WX849), .QN(n15686) );
  NOR2X0 U16541 ( .IN1(WX849), .IN2(n8736), .QN(n15684) );
  NOR2X0 U16542 ( .IN1(n15687), .IN2(n15688), .QN(n15678) );
  INVX0 U16543 ( .INP(n15689), .ZN(n15688) );
  NAND2X0 U16544 ( .IN1(n3517), .IN2(n9123), .QN(n15689) );
  NOR2X0 U16545 ( .IN1(n9115), .IN2(n3517), .QN(n15687) );
  NOR2X0 U16546 ( .IN1(n15690), .IN2(n15691), .QN(DATA_9_24) );
  INVX0 U16547 ( .INP(n15692), .ZN(n15691) );
  NAND2X0 U16548 ( .IN1(n15693), .IN2(n11573), .QN(n15692) );
  NOR2X0 U16549 ( .IN1(n11573), .IN2(n15693), .QN(n15690) );
  NAND2X0 U16550 ( .IN1(TM0), .IN2(WX499), .QN(n15693) );
  NAND2X0 U16551 ( .IN1(n15694), .IN2(n15695), .QN(n11573) );
  NAND2X0 U16552 ( .IN1(n15696), .IN2(n15697), .QN(n15695) );
  NAND2X0 U16553 ( .IN1(n15698), .IN2(n15699), .QN(n15696) );
  NAND3X0 U16554 ( .IN1(n15698), .IN2(n15699), .IN3(n15700), .QN(n15694) );
  INVX0 U16555 ( .INP(n15697), .ZN(n15700) );
  NOR2X0 U16556 ( .IN1(n15701), .IN2(n15702), .QN(n15697) );
  INVX0 U16557 ( .INP(n15703), .ZN(n15702) );
  NAND2X0 U16558 ( .IN1(n8743), .IN2(n15704), .QN(n15703) );
  NOR2X0 U16559 ( .IN1(n15704), .IN2(n8743), .QN(n15701) );
  NOR2X0 U16560 ( .IN1(n15705), .IN2(n15706), .QN(n15704) );
  INVX0 U16561 ( .INP(n15707), .ZN(n15706) );
  NAND2X0 U16562 ( .IN1(test_so4), .IN2(WX851), .QN(n15707) );
  NOR2X0 U16563 ( .IN1(WX851), .IN2(test_so4), .QN(n15705) );
  NAND2X0 U16564 ( .IN1(n3515), .IN2(n9123), .QN(n15699) );
  NAND2X0 U16565 ( .IN1(TM1), .IN2(WX659), .QN(n15698) );
  NAND2X0 U16566 ( .IN1(n15708), .IN2(n15709), .QN(DATA_9_23) );
  INVX0 U16567 ( .INP(n15710), .ZN(n15709) );
  NOR2X0 U16568 ( .IN1(n15711), .IN2(n11561), .QN(n15710) );
  NAND2X0 U16569 ( .IN1(n11561), .IN2(n15711), .QN(n15708) );
  NAND2X0 U16570 ( .IN1(TM0), .IN2(WX501), .QN(n15711) );
  NAND2X0 U16571 ( .IN1(n15712), .IN2(n15713), .QN(n11561) );
  NAND2X0 U16572 ( .IN1(n15714), .IN2(n15715), .QN(n15713) );
  INVX0 U16573 ( .INP(n15716), .ZN(n15712) );
  NOR2X0 U16574 ( .IN1(n15715), .IN2(n15714), .QN(n15716) );
  NAND2X0 U16575 ( .IN1(n15717), .IN2(n15718), .QN(n15714) );
  NAND2X0 U16576 ( .IN1(n8745), .IN2(n15719), .QN(n15718) );
  INVX0 U16577 ( .INP(n15720), .ZN(n15717) );
  NOR2X0 U16578 ( .IN1(n15719), .IN2(n8745), .QN(n15720) );
  NOR2X0 U16579 ( .IN1(n15721), .IN2(n15722), .QN(n15719) );
  INVX0 U16580 ( .INP(n15723), .ZN(n15722) );
  NAND2X0 U16581 ( .IN1(n8747), .IN2(WX853), .QN(n15723) );
  NOR2X0 U16582 ( .IN1(WX853), .IN2(n8747), .QN(n15721) );
  NOR2X0 U16583 ( .IN1(n15724), .IN2(n15725), .QN(n15715) );
  INVX0 U16584 ( .INP(n15726), .ZN(n15725) );
  NAND2X0 U16585 ( .IN1(n3513), .IN2(n9123), .QN(n15726) );
  NOR2X0 U16586 ( .IN1(n9115), .IN2(n3513), .QN(n15724) );
  NAND2X0 U16587 ( .IN1(n15727), .IN2(n15728), .QN(DATA_9_22) );
  INVX0 U16588 ( .INP(n15729), .ZN(n15728) );
  NOR2X0 U16589 ( .IN1(n15730), .IN2(n11550), .QN(n15729) );
  NAND2X0 U16590 ( .IN1(n11550), .IN2(n15730), .QN(n15727) );
  NAND2X0 U16591 ( .IN1(TM0), .IN2(WX503), .QN(n15730) );
  NAND2X0 U16592 ( .IN1(n15731), .IN2(n15732), .QN(n11550) );
  NAND2X0 U16593 ( .IN1(n15733), .IN2(n15734), .QN(n15732) );
  INVX0 U16594 ( .INP(n15735), .ZN(n15731) );
  NOR2X0 U16595 ( .IN1(n15734), .IN2(n15733), .QN(n15735) );
  NAND2X0 U16596 ( .IN1(n15736), .IN2(n15737), .QN(n15733) );
  NAND2X0 U16597 ( .IN1(n8759), .IN2(n15738), .QN(n15737) );
  INVX0 U16598 ( .INP(n15739), .ZN(n15736) );
  NOR2X0 U16599 ( .IN1(n15738), .IN2(n8759), .QN(n15739) );
  NOR2X0 U16600 ( .IN1(n15740), .IN2(n15741), .QN(n15738) );
  NOR2X0 U16601 ( .IN1(WX855), .IN2(n8760), .QN(n15741) );
  INVX0 U16602 ( .INP(n15742), .ZN(n15740) );
  NAND2X0 U16603 ( .IN1(n8760), .IN2(WX855), .QN(n15742) );
  NOR2X0 U16604 ( .IN1(n15743), .IN2(n15744), .QN(n15734) );
  INVX0 U16605 ( .INP(n15745), .ZN(n15744) );
  NAND2X0 U16606 ( .IN1(n3511), .IN2(n9123), .QN(n15745) );
  NOR2X0 U16607 ( .IN1(n9115), .IN2(n3511), .QN(n15743) );
  NAND2X0 U16608 ( .IN1(n15746), .IN2(n15747), .QN(DATA_9_21) );
  INVX0 U16609 ( .INP(n15748), .ZN(n15747) );
  NOR2X0 U16610 ( .IN1(n15749), .IN2(n11539), .QN(n15748) );
  NAND2X0 U16611 ( .IN1(n11539), .IN2(n15749), .QN(n15746) );
  NAND2X0 U16612 ( .IN1(TM0), .IN2(WX505), .QN(n15749) );
  NAND2X0 U16613 ( .IN1(n15750), .IN2(n15751), .QN(n11539) );
  NAND2X0 U16614 ( .IN1(n15752), .IN2(n15753), .QN(n15751) );
  INVX0 U16615 ( .INP(n15754), .ZN(n15750) );
  NOR2X0 U16616 ( .IN1(n15753), .IN2(n15752), .QN(n15754) );
  NAND2X0 U16617 ( .IN1(n15755), .IN2(n15756), .QN(n15752) );
  NAND2X0 U16618 ( .IN1(n8765), .IN2(n15757), .QN(n15756) );
  INVX0 U16619 ( .INP(n15758), .ZN(n15755) );
  NOR2X0 U16620 ( .IN1(n15757), .IN2(n8765), .QN(n15758) );
  NOR2X0 U16621 ( .IN1(n15759), .IN2(n15760), .QN(n15757) );
  NOR2X0 U16622 ( .IN1(WX857), .IN2(n8766), .QN(n15760) );
  INVX0 U16623 ( .INP(n15761), .ZN(n15759) );
  NAND2X0 U16624 ( .IN1(n8766), .IN2(WX857), .QN(n15761) );
  NOR2X0 U16625 ( .IN1(n15762), .IN2(n15763), .QN(n15753) );
  INVX0 U16626 ( .INP(n15764), .ZN(n15763) );
  NAND2X0 U16627 ( .IN1(n3509), .IN2(n9123), .QN(n15764) );
  NOR2X0 U16628 ( .IN1(n9115), .IN2(n3509), .QN(n15762) );
  NOR2X0 U16629 ( .IN1(n15765), .IN2(n15766), .QN(DATA_9_20) );
  INVX0 U16630 ( .INP(n15767), .ZN(n15766) );
  NAND2X0 U16631 ( .IN1(n15768), .IN2(n11528), .QN(n15767) );
  NOR2X0 U16632 ( .IN1(n11528), .IN2(n15768), .QN(n15765) );
  NAND2X0 U16633 ( .IN1(TM0), .IN2(WX507), .QN(n15768) );
  NAND2X0 U16634 ( .IN1(n15769), .IN2(n15770), .QN(n11528) );
  NAND2X0 U16635 ( .IN1(n15771), .IN2(n15772), .QN(n15770) );
  NAND2X0 U16636 ( .IN1(n15773), .IN2(n15774), .QN(n15771) );
  NAND3X0 U16637 ( .IN1(n15773), .IN2(n15774), .IN3(n15775), .QN(n15769) );
  INVX0 U16638 ( .INP(n15772), .ZN(n15775) );
  NOR2X0 U16639 ( .IN1(n15776), .IN2(n15777), .QN(n15772) );
  INVX0 U16640 ( .INP(n15778), .ZN(n15777) );
  NAND2X0 U16641 ( .IN1(n8770), .IN2(n15779), .QN(n15778) );
  NOR2X0 U16642 ( .IN1(n15779), .IN2(n8770), .QN(n15776) );
  NOR2X0 U16643 ( .IN1(n15780), .IN2(n15781), .QN(n15779) );
  INVX0 U16644 ( .INP(n15782), .ZN(n15781) );
  NAND2X0 U16645 ( .IN1(test_so6), .IN2(WX731), .QN(n15782) );
  NOR2X0 U16646 ( .IN1(WX731), .IN2(test_so6), .QN(n15780) );
  NAND2X0 U16647 ( .IN1(n3507), .IN2(n9123), .QN(n15774) );
  NAND2X0 U16648 ( .IN1(TM1), .IN2(WX667), .QN(n15773) );
  NOR2X0 U16649 ( .IN1(n15783), .IN2(n15784), .QN(DATA_9_2) );
  INVX0 U16650 ( .INP(n15785), .ZN(n15784) );
  NAND2X0 U16651 ( .IN1(n15786), .IN2(n11393), .QN(n15785) );
  NOR2X0 U16652 ( .IN1(n11393), .IN2(n15786), .QN(n15783) );
  NAND2X0 U16653 ( .IN1(TM0), .IN2(WX543), .QN(n15786) );
  NAND2X0 U16654 ( .IN1(n15787), .IN2(n15788), .QN(n11393) );
  NAND2X0 U16655 ( .IN1(n15789), .IN2(n15790), .QN(n15788) );
  NAND2X0 U16656 ( .IN1(n15791), .IN2(n15792), .QN(n15789) );
  NAND3X0 U16657 ( .IN1(n15791), .IN2(n15792), .IN3(n15793), .QN(n15787) );
  INVX0 U16658 ( .INP(n15790), .ZN(n15793) );
  NOR2X0 U16659 ( .IN1(n15794), .IN2(n15795), .QN(n15790) );
  INVX0 U16660 ( .INP(n15796), .ZN(n15795) );
  NAND2X0 U16661 ( .IN1(n8778), .IN2(n15797), .QN(n15796) );
  NOR2X0 U16662 ( .IN1(n15797), .IN2(n8778), .QN(n15794) );
  NOR2X0 U16663 ( .IN1(n15798), .IN2(n15799), .QN(n15797) );
  INVX0 U16664 ( .INP(n15800), .ZN(n15799) );
  NAND2X0 U16665 ( .IN1(test_so7), .IN2(WX895), .QN(n15800) );
  NOR2X0 U16666 ( .IN1(WX895), .IN2(test_so7), .QN(n15798) );
  NAND2X0 U16667 ( .IN1(n3471), .IN2(n2182), .QN(n15792) );
  NAND2X0 U16668 ( .IN1(TM0), .IN2(WX703), .QN(n15791) );
  NAND2X0 U16669 ( .IN1(n15801), .IN2(n15802), .QN(DATA_9_19) );
  INVX0 U16670 ( .INP(n15803), .ZN(n15802) );
  NOR2X0 U16671 ( .IN1(n15804), .IN2(n11516), .QN(n15803) );
  NAND2X0 U16672 ( .IN1(n11516), .IN2(n15804), .QN(n15801) );
  NAND2X0 U16673 ( .IN1(TM0), .IN2(WX509), .QN(n15804) );
  NAND2X0 U16674 ( .IN1(n15805), .IN2(n15806), .QN(n11516) );
  NAND2X0 U16675 ( .IN1(n15807), .IN2(n15808), .QN(n15806) );
  INVX0 U16676 ( .INP(n15809), .ZN(n15805) );
  NOR2X0 U16677 ( .IN1(n15808), .IN2(n15807), .QN(n15809) );
  NAND2X0 U16678 ( .IN1(n15810), .IN2(n15811), .QN(n15807) );
  NAND2X0 U16679 ( .IN1(n8704), .IN2(n15812), .QN(n15811) );
  INVX0 U16680 ( .INP(n15813), .ZN(n15810) );
  NOR2X0 U16681 ( .IN1(n15812), .IN2(n8704), .QN(n15813) );
  NOR2X0 U16682 ( .IN1(n15814), .IN2(n15815), .QN(n15812) );
  INVX0 U16683 ( .INP(n15816), .ZN(n15815) );
  NAND2X0 U16684 ( .IN1(n8706), .IN2(WX861), .QN(n15816) );
  NOR2X0 U16685 ( .IN1(WX861), .IN2(n8706), .QN(n15814) );
  NOR2X0 U16686 ( .IN1(n15817), .IN2(n15818), .QN(n15808) );
  INVX0 U16687 ( .INP(n15819), .ZN(n15818) );
  NAND2X0 U16688 ( .IN1(n3505), .IN2(n9123), .QN(n15819) );
  NOR2X0 U16689 ( .IN1(n9115), .IN2(n3505), .QN(n15817) );
  NAND2X0 U16690 ( .IN1(n15820), .IN2(n15821), .QN(DATA_9_18) );
  INVX0 U16691 ( .INP(n15822), .ZN(n15821) );
  NOR2X0 U16692 ( .IN1(n15823), .IN2(n11505), .QN(n15822) );
  NAND2X0 U16693 ( .IN1(n11505), .IN2(n15823), .QN(n15820) );
  NAND2X0 U16694 ( .IN1(TM0), .IN2(WX511), .QN(n15823) );
  NAND2X0 U16695 ( .IN1(n15824), .IN2(n15825), .QN(n11505) );
  NAND2X0 U16696 ( .IN1(n15826), .IN2(n15827), .QN(n15825) );
  INVX0 U16697 ( .INP(n15828), .ZN(n15824) );
  NOR2X0 U16698 ( .IN1(n15827), .IN2(n15826), .QN(n15828) );
  NAND2X0 U16699 ( .IN1(n15829), .IN2(n15830), .QN(n15826) );
  NAND2X0 U16700 ( .IN1(n8719), .IN2(n15831), .QN(n15830) );
  INVX0 U16701 ( .INP(n15832), .ZN(n15829) );
  NOR2X0 U16702 ( .IN1(n15831), .IN2(n8719), .QN(n15832) );
  NOR2X0 U16703 ( .IN1(n15833), .IN2(n15834), .QN(n15831) );
  INVX0 U16704 ( .INP(n15835), .ZN(n15834) );
  NAND2X0 U16705 ( .IN1(n8721), .IN2(WX863), .QN(n15835) );
  NOR2X0 U16706 ( .IN1(WX863), .IN2(n8721), .QN(n15833) );
  NOR2X0 U16707 ( .IN1(n15836), .IN2(n15837), .QN(n15827) );
  INVX0 U16708 ( .INP(n15838), .ZN(n15837) );
  NAND2X0 U16709 ( .IN1(n3503), .IN2(n9123), .QN(n15838) );
  NOR2X0 U16710 ( .IN1(n9115), .IN2(n3503), .QN(n15836) );
  NAND2X0 U16711 ( .IN1(n15839), .IN2(n15840), .QN(DATA_9_17) );
  INVX0 U16712 ( .INP(n15841), .ZN(n15840) );
  NOR2X0 U16713 ( .IN1(n15842), .IN2(n11499), .QN(n15841) );
  NAND2X0 U16714 ( .IN1(n11499), .IN2(n15842), .QN(n15839) );
  NAND2X0 U16715 ( .IN1(TM0), .IN2(WX513), .QN(n15842) );
  NAND2X0 U16716 ( .IN1(n15843), .IN2(n15844), .QN(n11499) );
  NAND2X0 U16717 ( .IN1(n15845), .IN2(n15846), .QN(n15844) );
  INVX0 U16718 ( .INP(n15847), .ZN(n15843) );
  NOR2X0 U16719 ( .IN1(n15846), .IN2(n15845), .QN(n15847) );
  NAND2X0 U16720 ( .IN1(n15848), .IN2(n15849), .QN(n15845) );
  NAND2X0 U16721 ( .IN1(n8731), .IN2(n15850), .QN(n15849) );
  INVX0 U16722 ( .INP(n15851), .ZN(n15848) );
  NOR2X0 U16723 ( .IN1(n15850), .IN2(n8731), .QN(n15851) );
  NOR2X0 U16724 ( .IN1(n15852), .IN2(n15853), .QN(n15850) );
  INVX0 U16725 ( .INP(n15854), .ZN(n15853) );
  NAND2X0 U16726 ( .IN1(n8733), .IN2(WX865), .QN(n15854) );
  NOR2X0 U16727 ( .IN1(WX865), .IN2(n8733), .QN(n15852) );
  NOR2X0 U16728 ( .IN1(n15855), .IN2(n15856), .QN(n15846) );
  INVX0 U16729 ( .INP(n15857), .ZN(n15856) );
  NAND2X0 U16730 ( .IN1(n3501), .IN2(n9123), .QN(n15857) );
  NOR2X0 U16731 ( .IN1(n9115), .IN2(n3501), .QN(n15855) );
  NOR2X0 U16732 ( .IN1(n15858), .IN2(n15859), .QN(DATA_9_16) );
  INVX0 U16733 ( .INP(n15860), .ZN(n15859) );
  NAND2X0 U16734 ( .IN1(n15861), .IN2(n11488), .QN(n15860) );
  NOR2X0 U16735 ( .IN1(n11488), .IN2(n15861), .QN(n15858) );
  NAND2X0 U16736 ( .IN1(TM0), .IN2(WX515), .QN(n15861) );
  NAND2X0 U16737 ( .IN1(n15862), .IN2(n15863), .QN(n11488) );
  NAND2X0 U16738 ( .IN1(n15864), .IN2(n15865), .QN(n15863) );
  NAND2X0 U16739 ( .IN1(n15866), .IN2(n15867), .QN(n15864) );
  NAND3X0 U16740 ( .IN1(n15866), .IN2(n15867), .IN3(n15868), .QN(n15862) );
  INVX0 U16741 ( .INP(n15865), .ZN(n15868) );
  NOR2X0 U16742 ( .IN1(n15869), .IN2(n15870), .QN(n15865) );
  INVX0 U16743 ( .INP(n15871), .ZN(n15870) );
  NAND2X0 U16744 ( .IN1(n8748), .IN2(n15872), .QN(n15871) );
  NOR2X0 U16745 ( .IN1(n15872), .IN2(n8748), .QN(n15869) );
  NOR2X0 U16746 ( .IN1(n15873), .IN2(n15874), .QN(n15872) );
  NOR2X0 U16747 ( .IN1(n8797), .IN2(n8749), .QN(n15874) );
  INVX0 U16748 ( .INP(n15875), .ZN(n15873) );
  NAND2X0 U16749 ( .IN1(n8749), .IN2(n8797), .QN(n15875) );
  NAND2X0 U16750 ( .IN1(n3499), .IN2(n9117), .QN(n15867) );
  INVX0 U16751 ( .INP(TM1), .ZN(n10355) );
  NAND2X0 U16752 ( .IN1(TM1), .IN2(WX675), .QN(n15866) );
  NAND2X0 U16753 ( .IN1(n15876), .IN2(n15877), .QN(DATA_9_15) );
  INVX0 U16754 ( .INP(n15878), .ZN(n15877) );
  NOR2X0 U16755 ( .IN1(n15879), .IN2(n11476), .QN(n15878) );
  NAND2X0 U16756 ( .IN1(n11476), .IN2(n15879), .QN(n15876) );
  NAND2X0 U16757 ( .IN1(TM0), .IN2(WX517), .QN(n15879) );
  NAND2X0 U16758 ( .IN1(n15880), .IN2(n15881), .QN(n11476) );
  NAND2X0 U16759 ( .IN1(n15882), .IN2(n15883), .QN(n15881) );
  INVX0 U16760 ( .INP(n15884), .ZN(n15880) );
  NOR2X0 U16761 ( .IN1(n15883), .IN2(n15882), .QN(n15884) );
  NAND2X0 U16762 ( .IN1(n15885), .IN2(n15886), .QN(n15882) );
  NAND2X0 U16763 ( .IN1(n8762), .IN2(n15887), .QN(n15886) );
  INVX0 U16764 ( .INP(n15888), .ZN(n15885) );
  NOR2X0 U16765 ( .IN1(n15887), .IN2(n8762), .QN(n15888) );
  NOR2X0 U16766 ( .IN1(n15889), .IN2(n15890), .QN(n15887) );
  NOR2X0 U16767 ( .IN1(WX869), .IN2(n8763), .QN(n15890) );
  INVX0 U16768 ( .INP(n15891), .ZN(n15889) );
  NAND2X0 U16769 ( .IN1(n8763), .IN2(WX869), .QN(n15891) );
  NOR2X0 U16770 ( .IN1(n15892), .IN2(n15893), .QN(n15883) );
  INVX0 U16771 ( .INP(n15894), .ZN(n15893) );
  NAND2X0 U16772 ( .IN1(n3497), .IN2(n2182), .QN(n15894) );
  NOR2X0 U16773 ( .IN1(n2182), .IN2(n3497), .QN(n15892) );
  NAND2X0 U16774 ( .IN1(n15895), .IN2(n15896), .QN(DATA_9_14) );
  INVX0 U16775 ( .INP(n15897), .ZN(n15896) );
  NOR2X0 U16776 ( .IN1(n15898), .IN2(n11470), .QN(n15897) );
  NAND2X0 U16777 ( .IN1(n11470), .IN2(n15898), .QN(n15895) );
  NAND2X0 U16778 ( .IN1(test_so1), .IN2(TM0), .QN(n15898) );
  NAND2X0 U16779 ( .IN1(n15899), .IN2(n15900), .QN(n11470) );
  NAND2X0 U16780 ( .IN1(n15901), .IN2(n15902), .QN(n15900) );
  INVX0 U16781 ( .INP(n15903), .ZN(n15899) );
  NOR2X0 U16782 ( .IN1(n15902), .IN2(n15901), .QN(n15903) );
  NAND2X0 U16783 ( .IN1(n15904), .IN2(n15905), .QN(n15901) );
  NAND2X0 U16784 ( .IN1(n8775), .IN2(n15906), .QN(n15905) );
  INVX0 U16785 ( .INP(n15907), .ZN(n15904) );
  NOR2X0 U16786 ( .IN1(n15906), .IN2(n8775), .QN(n15907) );
  NOR2X0 U16787 ( .IN1(n15908), .IN2(n15909), .QN(n15906) );
  INVX0 U16788 ( .INP(n15910), .ZN(n15909) );
  NAND2X0 U16789 ( .IN1(n8777), .IN2(WX871), .QN(n15910) );
  NOR2X0 U16790 ( .IN1(WX871), .IN2(n8777), .QN(n15908) );
  NOR2X0 U16791 ( .IN1(n15911), .IN2(n15912), .QN(n15902) );
  INVX0 U16792 ( .INP(n15913), .ZN(n15912) );
  NAND2X0 U16793 ( .IN1(n3495), .IN2(n2182), .QN(n15913) );
  NOR2X0 U16794 ( .IN1(n2182), .IN2(n3495), .QN(n15911) );
  NAND2X0 U16795 ( .IN1(n15914), .IN2(n15915), .QN(DATA_9_13) );
  INVX0 U16796 ( .INP(n15916), .ZN(n15915) );
  NOR2X0 U16797 ( .IN1(n15917), .IN2(n11463), .QN(n15916) );
  NAND2X0 U16798 ( .IN1(n11463), .IN2(n15917), .QN(n15914) );
  NAND2X0 U16799 ( .IN1(TM0), .IN2(WX521), .QN(n15917) );
  NAND2X0 U16800 ( .IN1(n15918), .IN2(n15919), .QN(n11463) );
  NAND2X0 U16801 ( .IN1(n15920), .IN2(n15921), .QN(n15919) );
  INVX0 U16802 ( .INP(n15922), .ZN(n15918) );
  NOR2X0 U16803 ( .IN1(n15921), .IN2(n15920), .QN(n15922) );
  NAND2X0 U16804 ( .IN1(n15923), .IN2(n15924), .QN(n15920) );
  NAND2X0 U16805 ( .IN1(n8710), .IN2(n15925), .QN(n15924) );
  INVX0 U16806 ( .INP(n15926), .ZN(n15923) );
  NOR2X0 U16807 ( .IN1(n15925), .IN2(n8710), .QN(n15926) );
  NOR2X0 U16808 ( .IN1(n15927), .IN2(n15928), .QN(n15925) );
  INVX0 U16809 ( .INP(n15929), .ZN(n15928) );
  NAND2X0 U16810 ( .IN1(n8712), .IN2(WX873), .QN(n15929) );
  NOR2X0 U16811 ( .IN1(WX873), .IN2(n8712), .QN(n15927) );
  NOR2X0 U16812 ( .IN1(n15930), .IN2(n15931), .QN(n15921) );
  INVX0 U16813 ( .INP(n15932), .ZN(n15931) );
  NAND2X0 U16814 ( .IN1(n3493), .IN2(n2182), .QN(n15932) );
  NOR2X0 U16815 ( .IN1(n2182), .IN2(n3493), .QN(n15930) );
  NAND2X0 U16816 ( .IN1(n15933), .IN2(n15934), .QN(DATA_9_12) );
  INVX0 U16817 ( .INP(n15935), .ZN(n15934) );
  NOR2X0 U16818 ( .IN1(n15936), .IN2(n11457), .QN(n15935) );
  NAND2X0 U16819 ( .IN1(n11457), .IN2(n15936), .QN(n15933) );
  NAND2X0 U16820 ( .IN1(TM0), .IN2(WX523), .QN(n15936) );
  NAND2X0 U16821 ( .IN1(n15937), .IN2(n15938), .QN(n11457) );
  NAND2X0 U16822 ( .IN1(n15939), .IN2(n15940), .QN(n15938) );
  INVX0 U16823 ( .INP(n15941), .ZN(n15937) );
  NOR2X0 U16824 ( .IN1(n15940), .IN2(n15939), .QN(n15941) );
  NAND2X0 U16825 ( .IN1(n15942), .IN2(n15943), .QN(n15939) );
  NAND2X0 U16826 ( .IN1(n8737), .IN2(n15944), .QN(n15943) );
  INVX0 U16827 ( .INP(n15945), .ZN(n15942) );
  NOR2X0 U16828 ( .IN1(n15944), .IN2(n8737), .QN(n15945) );
  NOR2X0 U16829 ( .IN1(n15946), .IN2(n15947), .QN(n15944) );
  INVX0 U16830 ( .INP(n15948), .ZN(n15947) );
  NAND2X0 U16831 ( .IN1(n8739), .IN2(WX875), .QN(n15948) );
  NOR2X0 U16832 ( .IN1(WX875), .IN2(n8739), .QN(n15946) );
  NOR2X0 U16833 ( .IN1(n15949), .IN2(n15950), .QN(n15940) );
  INVX0 U16834 ( .INP(n15951), .ZN(n15950) );
  NAND2X0 U16835 ( .IN1(n3491), .IN2(n2182), .QN(n15951) );
  NOR2X0 U16836 ( .IN1(n2182), .IN2(n3491), .QN(n15949) );
  NAND2X0 U16837 ( .IN1(n15952), .IN2(n15953), .QN(DATA_9_11) );
  INVX0 U16838 ( .INP(n15954), .ZN(n15953) );
  NOR2X0 U16839 ( .IN1(n15955), .IN2(n11451), .QN(n15954) );
  NAND2X0 U16840 ( .IN1(n11451), .IN2(n15955), .QN(n15952) );
  NAND2X0 U16841 ( .IN1(TM0), .IN2(WX525), .QN(n15955) );
  NAND2X0 U16842 ( .IN1(n15956), .IN2(n15957), .QN(n11451) );
  NAND2X0 U16843 ( .IN1(n15958), .IN2(n15959), .QN(n15957) );
  INVX0 U16844 ( .INP(n15960), .ZN(n15956) );
  NOR2X0 U16845 ( .IN1(n15959), .IN2(n15958), .QN(n15960) );
  NAND2X0 U16846 ( .IN1(n15961), .IN2(n15962), .QN(n15958) );
  NAND2X0 U16847 ( .IN1(n8783), .IN2(n15963), .QN(n15962) );
  INVX0 U16848 ( .INP(n15964), .ZN(n15961) );
  NOR2X0 U16849 ( .IN1(n15963), .IN2(n8783), .QN(n15964) );
  NOR2X0 U16850 ( .IN1(n15965), .IN2(n15966), .QN(n15963) );
  INVX0 U16851 ( .INP(n15967), .ZN(n15966) );
  NAND2X0 U16852 ( .IN1(n8785), .IN2(WX877), .QN(n15967) );
  NOR2X0 U16853 ( .IN1(WX877), .IN2(n8785), .QN(n15965) );
  NOR2X0 U16854 ( .IN1(n15968), .IN2(n15969), .QN(n15959) );
  INVX0 U16855 ( .INP(n15970), .ZN(n15969) );
  NAND2X0 U16856 ( .IN1(n3489), .IN2(n2182), .QN(n15970) );
  NOR2X0 U16857 ( .IN1(n2182), .IN2(n3489), .QN(n15968) );
  NOR2X0 U16858 ( .IN1(n15971), .IN2(n15972), .QN(DATA_9_10) );
  INVX0 U16859 ( .INP(n15973), .ZN(n15972) );
  NAND2X0 U16860 ( .IN1(n15974), .IN2(n11445), .QN(n15973) );
  NOR2X0 U16861 ( .IN1(n11445), .IN2(n15974), .QN(n15971) );
  NAND2X0 U16862 ( .IN1(TM0), .IN2(WX527), .QN(n15974) );
  NAND2X0 U16863 ( .IN1(n15975), .IN2(n15976), .QN(n11445) );
  NAND2X0 U16864 ( .IN1(n15977), .IN2(n15978), .QN(n15976) );
  NAND2X0 U16865 ( .IN1(n15979), .IN2(n15980), .QN(n15977) );
  NAND3X0 U16866 ( .IN1(n15979), .IN2(n15980), .IN3(n15981), .QN(n15975) );
  INVX0 U16867 ( .INP(n15978), .ZN(n15981) );
  NOR2X0 U16868 ( .IN1(n15982), .IN2(n15983), .QN(n15978) );
  INVX0 U16869 ( .INP(n15984), .ZN(n15983) );
  NAND2X0 U16870 ( .IN1(n8728), .IN2(n15985), .QN(n15984) );
  NOR2X0 U16871 ( .IN1(n15985), .IN2(n8728), .QN(n15982) );
  NOR2X0 U16872 ( .IN1(n15986), .IN2(n15987), .QN(n15985) );
  INVX0 U16873 ( .INP(n15988), .ZN(n15987) );
  NAND2X0 U16874 ( .IN1(test_so3), .IN2(WX879), .QN(n15988) );
  NOR2X0 U16875 ( .IN1(WX879), .IN2(test_so3), .QN(n15986) );
  NAND2X0 U16876 ( .IN1(n8730), .IN2(n2182), .QN(n15980) );
  NAND2X0 U16877 ( .IN1(TM0), .IN2(WX751), .QN(n15979) );
  NAND2X0 U16878 ( .IN1(n15989), .IN2(n15990), .QN(DATA_9_1) );
  INVX0 U16879 ( .INP(n15991), .ZN(n15990) );
  NOR2X0 U16880 ( .IN1(n15992), .IN2(n11386), .QN(n15991) );
  NAND2X0 U16881 ( .IN1(n11386), .IN2(n15992), .QN(n15989) );
  NAND2X0 U16882 ( .IN1(TM0), .IN2(WX545), .QN(n15992) );
  NAND2X0 U16883 ( .IN1(n15993), .IN2(n15994), .QN(n11386) );
  NAND2X0 U16884 ( .IN1(n15995), .IN2(n15996), .QN(n15994) );
  INVX0 U16885 ( .INP(n15997), .ZN(n15993) );
  NOR2X0 U16886 ( .IN1(n15996), .IN2(n15995), .QN(n15997) );
  NAND2X0 U16887 ( .IN1(n15998), .IN2(n15999), .QN(n15995) );
  NAND2X0 U16888 ( .IN1(n8713), .IN2(n16000), .QN(n15999) );
  INVX0 U16889 ( .INP(n16001), .ZN(n16000) );
  NAND2X0 U16890 ( .IN1(n16001), .IN2(WX897), .QN(n15998) );
  NAND2X0 U16891 ( .IN1(n16002), .IN2(n16003), .QN(n16001) );
  INVX0 U16892 ( .INP(n16004), .ZN(n16003) );
  NOR2X0 U16893 ( .IN1(WX833), .IN2(n8714), .QN(n16004) );
  NAND2X0 U16894 ( .IN1(n8714), .IN2(WX833), .QN(n16002) );
  NOR2X0 U16895 ( .IN1(n16005), .IN2(n16006), .QN(n15996) );
  INVX0 U16896 ( .INP(n16007), .ZN(n16006) );
  NAND2X0 U16897 ( .IN1(n3469), .IN2(n2182), .QN(n16007) );
  NOR2X0 U16898 ( .IN1(n2182), .IN2(n3469), .QN(n16005) );
  NAND2X0 U16899 ( .IN1(n16008), .IN2(n16009), .QN(DATA_9_0) );
  INVX0 U16900 ( .INP(n16010), .ZN(n16009) );
  NOR2X0 U16901 ( .IN1(n16011), .IN2(n11380), .QN(n16010) );
  NAND2X0 U16902 ( .IN1(n11380), .IN2(n16011), .QN(n16008) );
  NAND2X0 U16903 ( .IN1(TM0), .IN2(WX547), .QN(n16011) );
  NAND2X0 U16904 ( .IN1(n16012), .IN2(n16013), .QN(n11380) );
  NAND2X0 U16905 ( .IN1(n16014), .IN2(n16015), .QN(n16013) );
  INVX0 U16906 ( .INP(n16016), .ZN(n16012) );
  NOR2X0 U16907 ( .IN1(n16015), .IN2(n16014), .QN(n16016) );
  NAND2X0 U16908 ( .IN1(n16017), .IN2(n16018), .QN(n16014) );
  NAND2X0 U16909 ( .IN1(n8786), .IN2(n16019), .QN(n16018) );
  INVX0 U16910 ( .INP(n16020), .ZN(n16017) );
  NOR2X0 U16911 ( .IN1(n16019), .IN2(n8786), .QN(n16020) );
  NOR2X0 U16912 ( .IN1(n16021), .IN2(n16022), .QN(n16019) );
  NOR2X0 U16913 ( .IN1(WX899), .IN2(n8787), .QN(n16022) );
  INVX0 U16914 ( .INP(n16023), .ZN(n16021) );
  NAND2X0 U16915 ( .IN1(n8787), .IN2(WX899), .QN(n16023) );
  NOR2X0 U16916 ( .IN1(n16024), .IN2(n16025), .QN(n16015) );
  INVX0 U16917 ( .INP(n16026), .ZN(n16025) );
  NAND2X0 U16918 ( .IN1(n3467), .IN2(n2182), .QN(n16026) );
  NOR2X0 U16919 ( .IN1(n2182), .IN2(n3467), .QN(n16024) );
  INVX0 U16920 ( .INP(TM0), .ZN(n2182) );
  NOR2X0 U3558_U2 ( .IN1(n9179), .IN2(U3558_n1), .QN(n2245) );
  INVX0 U3558_U1 ( .INP(n9272), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(n3278), .ZN(U3871_n1) );
  NOR2X0 U3871_U1 ( .IN1(TM0), .IN2(U3871_n1), .QN(n2153) );
  INVX0 U3991_U2 ( .INP(n3278), .ZN(U3991_n1) );
  NOR2X0 U3991_U1 ( .IN1(n2182), .IN2(U3991_n1), .QN(n2152) );
  INVX0 U5716_U2 ( .INP(WX547), .ZN(U5716_n1) );
  NOR2X0 U5716_U1 ( .IN1(n9179), .IN2(U5716_n1), .QN(WX544) );
  INVX0 U5717_U2 ( .INP(WX545), .ZN(U5717_n1) );
  NOR2X0 U5717_U1 ( .IN1(n9179), .IN2(U5717_n1), .QN(WX542) );
  INVX0 U5718_U2 ( .INP(WX543), .ZN(U5718_n1) );
  NOR2X0 U5718_U1 ( .IN1(n9203), .IN2(U5718_n1), .QN(WX540) );
  INVX0 U5719_U2 ( .INP(WX541), .ZN(U5719_n1) );
  NOR2X0 U5719_U1 ( .IN1(n9197), .IN2(U5719_n1), .QN(WX538) );
  INVX0 U5720_U2 ( .INP(WX539), .ZN(U5720_n1) );
  NOR2X0 U5720_U1 ( .IN1(n9191), .IN2(U5720_n1), .QN(WX536) );
  INVX0 U5721_U2 ( .INP(WX537), .ZN(U5721_n1) );
  NOR2X0 U5721_U1 ( .IN1(n9191), .IN2(U5721_n1), .QN(WX534) );
  INVX0 U5722_U2 ( .INP(WX535), .ZN(U5722_n1) );
  NOR2X0 U5722_U1 ( .IN1(n9191), .IN2(U5722_n1), .QN(WX532) );
  INVX0 U5723_U2 ( .INP(WX533), .ZN(U5723_n1) );
  NOR2X0 U5723_U1 ( .IN1(n9191), .IN2(U5723_n1), .QN(WX530) );
  INVX0 U5724_U2 ( .INP(WX531), .ZN(U5724_n1) );
  NOR2X0 U5724_U1 ( .IN1(n9191), .IN2(U5724_n1), .QN(WX528) );
  INVX0 U5725_U2 ( .INP(WX529), .ZN(U5725_n1) );
  NOR2X0 U5725_U1 ( .IN1(n9192), .IN2(U5725_n1), .QN(WX526) );
  INVX0 U5726_U2 ( .INP(WX527), .ZN(U5726_n1) );
  NOR2X0 U5726_U1 ( .IN1(n9192), .IN2(U5726_n1), .QN(WX524) );
  INVX0 U5727_U2 ( .INP(WX525), .ZN(U5727_n1) );
  NOR2X0 U5727_U1 ( .IN1(n9192), .IN2(U5727_n1), .QN(WX522) );
  INVX0 U5728_U2 ( .INP(WX523), .ZN(U5728_n1) );
  NOR2X0 U5728_U1 ( .IN1(n9192), .IN2(U5728_n1), .QN(WX520) );
  INVX0 U5729_U2 ( .INP(WX521), .ZN(U5729_n1) );
  NOR2X0 U5729_U1 ( .IN1(n9192), .IN2(U5729_n1), .QN(WX518) );
  INVX0 U5730_U2 ( .INP(test_so1), .ZN(U5730_n1) );
  NOR2X0 U5730_U1 ( .IN1(n9192), .IN2(U5730_n1), .QN(WX516) );
  INVX0 U5731_U2 ( .INP(WX517), .ZN(U5731_n1) );
  NOR2X0 U5731_U1 ( .IN1(n9192), .IN2(U5731_n1), .QN(WX514) );
  INVX0 U5732_U2 ( .INP(WX515), .ZN(U5732_n1) );
  NOR2X0 U5732_U1 ( .IN1(n9192), .IN2(U5732_n1), .QN(WX512) );
  INVX0 U5733_U2 ( .INP(WX513), .ZN(U5733_n1) );
  NOR2X0 U5733_U1 ( .IN1(n9192), .IN2(U5733_n1), .QN(WX510) );
  INVX0 U5734_U2 ( .INP(WX511), .ZN(U5734_n1) );
  NOR2X0 U5734_U1 ( .IN1(n9192), .IN2(U5734_n1), .QN(WX508) );
  INVX0 U5735_U2 ( .INP(WX509), .ZN(U5735_n1) );
  NOR2X0 U5735_U1 ( .IN1(n9192), .IN2(U5735_n1), .QN(WX506) );
  INVX0 U5736_U2 ( .INP(WX507), .ZN(U5736_n1) );
  NOR2X0 U5736_U1 ( .IN1(n9192), .IN2(U5736_n1), .QN(WX504) );
  INVX0 U5737_U2 ( .INP(WX505), .ZN(U5737_n1) );
  NOR2X0 U5737_U1 ( .IN1(n9192), .IN2(U5737_n1), .QN(WX502) );
  INVX0 U5738_U2 ( .INP(WX503), .ZN(U5738_n1) );
  NOR2X0 U5738_U1 ( .IN1(n9193), .IN2(U5738_n1), .QN(WX500) );
  INVX0 U5739_U2 ( .INP(WX501), .ZN(U5739_n1) );
  NOR2X0 U5739_U1 ( .IN1(n9193), .IN2(U5739_n1), .QN(WX498) );
  INVX0 U5740_U2 ( .INP(WX499), .ZN(U5740_n1) );
  NOR2X0 U5740_U1 ( .IN1(n9193), .IN2(U5740_n1), .QN(WX496) );
  INVX0 U5741_U2 ( .INP(WX497), .ZN(U5741_n1) );
  NOR2X0 U5741_U1 ( .IN1(n9193), .IN2(U5741_n1), .QN(WX494) );
  INVX0 U5742_U2 ( .INP(WX495), .ZN(U5742_n1) );
  NOR2X0 U5742_U1 ( .IN1(n9193), .IN2(U5742_n1), .QN(WX492) );
  INVX0 U5743_U2 ( .INP(WX493), .ZN(U5743_n1) );
  NOR2X0 U5743_U1 ( .IN1(n9193), .IN2(U5743_n1), .QN(WX490) );
  INVX0 U5744_U2 ( .INP(WX491), .ZN(U5744_n1) );
  NOR2X0 U5744_U1 ( .IN1(n9193), .IN2(U5744_n1), .QN(WX488) );
  INVX0 U5745_U2 ( .INP(WX489), .ZN(U5745_n1) );
  NOR2X0 U5745_U1 ( .IN1(n9193), .IN2(U5745_n1), .QN(WX486) );
  INVX0 U5746_U2 ( .INP(WX487), .ZN(U5746_n1) );
  NOR2X0 U5746_U1 ( .IN1(n9193), .IN2(U5746_n1), .QN(WX484) );
  INVX0 U5747_U2 ( .INP(WX5939), .ZN(U5747_n1) );
  NOR2X0 U5747_U1 ( .IN1(n9193), .IN2(U5747_n1), .QN(WX6002) );
  INVX0 U5748_U2 ( .INP(test_so49), .ZN(U5748_n1) );
  NOR2X0 U5748_U1 ( .IN1(n9193), .IN2(U5748_n1), .QN(WX6000) );
  INVX0 U5749_U2 ( .INP(WX5935), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n9193), .IN2(U5749_n1), .QN(WX5998) );
  INVX0 U5750_U2 ( .INP(WX5933), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n9193), .IN2(U5750_n1), .QN(WX5996) );
  INVX0 U5751_U2 ( .INP(WX5931), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n9194), .IN2(U5751_n1), .QN(WX5994) );
  INVX0 U5752_U2 ( .INP(WX3269), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n9194), .IN2(U5752_n1), .QN(WX3332) );
  INVX0 U5753_U2 ( .INP(WX3265), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n9194), .IN2(U5753_n1), .QN(WX3328) );
  INVX0 U5754_U2 ( .INP(WX3263), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n9194), .IN2(U5754_n1), .QN(WX3326) );
  INVX0 U5755_U2 ( .INP(WX11179), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n9194), .IN2(U5755_n1), .QN(WX11242) );
  INVX0 U5756_U2 ( .INP(WX11177), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n9194), .IN2(U5756_n1), .QN(WX11240) );
  INVX0 U5757_U2 ( .INP(WX11175), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n9194), .IN2(U5757_n1), .QN(WX11238) );
  INVX0 U5758_U2 ( .INP(WX11173), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n9194), .IN2(U5758_n1), .QN(WX11236) );
  INVX0 U5759_U2 ( .INP(test_so96), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n9194), .IN2(U5759_n1), .QN(WX11234) );
  INVX0 U5760_U2 ( .INP(WX11169), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n9194), .IN2(U5760_n1), .QN(WX11232) );
  INVX0 U5761_U2 ( .INP(WX11167), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n9194), .IN2(U5761_n1), .QN(WX11230) );
  INVX0 U5762_U2 ( .INP(WX11165), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n9194), .IN2(U5762_n1), .QN(WX11228) );
  INVX0 U5763_U2 ( .INP(WX11163), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n9194), .IN2(U5763_n1), .QN(WX11226) );
  INVX0 U5764_U2 ( .INP(WX11161), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n9195), .IN2(U5764_n1), .QN(WX11224) );
  INVX0 U5765_U2 ( .INP(WX11159), .ZN(U5765_n1) );
  NOR2X0 U5765_U1 ( .IN1(n9195), .IN2(U5765_n1), .QN(WX11222) );
  INVX0 U5766_U2 ( .INP(WX11157), .ZN(U5766_n1) );
  NOR2X0 U5766_U1 ( .IN1(n9195), .IN2(U5766_n1), .QN(WX11220) );
  INVX0 U5767_U2 ( .INP(WX11155), .ZN(U5767_n1) );
  NOR2X0 U5767_U1 ( .IN1(n9195), .IN2(U5767_n1), .QN(WX11218) );
  INVX0 U5768_U2 ( .INP(WX11153), .ZN(U5768_n1) );
  NOR2X0 U5768_U1 ( .IN1(n9195), .IN2(U5768_n1), .QN(WX11216) );
  INVX0 U5769_U2 ( .INP(WX11151), .ZN(U5769_n1) );
  NOR2X0 U5769_U1 ( .IN1(n9195), .IN2(U5769_n1), .QN(WX11214) );
  INVX0 U5770_U2 ( .INP(WX11149), .ZN(U5770_n1) );
  NOR2X0 U5770_U1 ( .IN1(n9195), .IN2(U5770_n1), .QN(WX11212) );
  INVX0 U5771_U2 ( .INP(WX11147), .ZN(U5771_n1) );
  NOR2X0 U5771_U1 ( .IN1(n9195), .IN2(U5771_n1), .QN(WX11210) );
  INVX0 U5772_U2 ( .INP(WX11145), .ZN(U5772_n1) );
  NOR2X0 U5772_U1 ( .IN1(n9195), .IN2(U5772_n1), .QN(WX11208) );
  INVX0 U5773_U2 ( .INP(WX11143), .ZN(U5773_n1) );
  NOR2X0 U5773_U1 ( .IN1(n9195), .IN2(U5773_n1), .QN(WX11206) );
  INVX0 U5774_U2 ( .INP(WX11141), .ZN(U5774_n1) );
  NOR2X0 U5774_U1 ( .IN1(n9195), .IN2(U5774_n1), .QN(WX11204) );
  INVX0 U5775_U2 ( .INP(WX11139), .ZN(U5775_n1) );
  NOR2X0 U5775_U1 ( .IN1(n9195), .IN2(U5775_n1), .QN(WX11202) );
  INVX0 U5776_U2 ( .INP(test_so95), .ZN(U5776_n1) );
  NOR2X0 U5776_U1 ( .IN1(n9195), .IN2(U5776_n1), .QN(WX11200) );
  INVX0 U5777_U2 ( .INP(WX11135), .ZN(U5777_n1) );
  NOR2X0 U5777_U1 ( .IN1(n9196), .IN2(U5777_n1), .QN(WX11198) );
  INVX0 U5778_U2 ( .INP(WX11133), .ZN(U5778_n1) );
  NOR2X0 U5778_U1 ( .IN1(n9196), .IN2(U5778_n1), .QN(WX11196) );
  INVX0 U5779_U2 ( .INP(WX11131), .ZN(U5779_n1) );
  NOR2X0 U5779_U1 ( .IN1(n9196), .IN2(U5779_n1), .QN(WX11194) );
  INVX0 U5780_U2 ( .INP(WX11129), .ZN(U5780_n1) );
  NOR2X0 U5780_U1 ( .IN1(n9196), .IN2(U5780_n1), .QN(WX11192) );
  INVX0 U5781_U2 ( .INP(WX11127), .ZN(U5781_n1) );
  NOR2X0 U5781_U1 ( .IN1(n9196), .IN2(U5781_n1), .QN(WX11190) );
  INVX0 U5782_U2 ( .INP(WX11125), .ZN(U5782_n1) );
  NOR2X0 U5782_U1 ( .IN1(n9196), .IN2(U5782_n1), .QN(WX11188) );
  INVX0 U5783_U2 ( .INP(WX11123), .ZN(U5783_n1) );
  NOR2X0 U5783_U1 ( .IN1(n9196), .IN2(U5783_n1), .QN(WX11186) );
  INVX0 U5784_U2 ( .INP(WX11121), .ZN(U5784_n1) );
  NOR2X0 U5784_U1 ( .IN1(n9196), .IN2(U5784_n1), .QN(WX11184) );
  INVX0 U5785_U2 ( .INP(WX11119), .ZN(U5785_n1) );
  NOR2X0 U5785_U1 ( .IN1(n9196), .IN2(U5785_n1), .QN(WX11182) );
  INVX0 U5786_U2 ( .INP(WX11117), .ZN(U5786_n1) );
  NOR2X0 U5786_U1 ( .IN1(n9196), .IN2(U5786_n1), .QN(WX11180) );
  INVX0 U5787_U2 ( .INP(WX11115), .ZN(U5787_n1) );
  NOR2X0 U5787_U1 ( .IN1(n9196), .IN2(U5787_n1), .QN(WX11178) );
  INVX0 U5788_U2 ( .INP(WX11113), .ZN(U5788_n1) );
  NOR2X0 U5788_U1 ( .IN1(n9196), .IN2(U5788_n1), .QN(WX11176) );
  INVX0 U5789_U2 ( .INP(WX11111), .ZN(U5789_n1) );
  NOR2X0 U5789_U1 ( .IN1(n9196), .IN2(U5789_n1), .QN(WX11174) );
  INVX0 U5790_U2 ( .INP(WX11109), .ZN(U5790_n1) );
  NOR2X0 U5790_U1 ( .IN1(n9197), .IN2(U5790_n1), .QN(WX11172) );
  INVX0 U5791_U2 ( .INP(WX11107), .ZN(U5791_n1) );
  NOR2X0 U5791_U1 ( .IN1(n9197), .IN2(U5791_n1), .QN(WX11170) );
  INVX0 U5792_U2 ( .INP(WX11105), .ZN(U5792_n1) );
  NOR2X0 U5792_U1 ( .IN1(n9197), .IN2(U5792_n1), .QN(WX11168) );
  INVX0 U5793_U2 ( .INP(test_so94), .ZN(U5793_n1) );
  NOR2X0 U5793_U1 ( .IN1(n9197), .IN2(U5793_n1), .QN(WX11166) );
  INVX0 U5794_U2 ( .INP(WX11101), .ZN(U5794_n1) );
  NOR2X0 U5794_U1 ( .IN1(n9197), .IN2(U5794_n1), .QN(WX11164) );
  INVX0 U5795_U2 ( .INP(WX11099), .ZN(U5795_n1) );
  NOR2X0 U5795_U1 ( .IN1(n9197), .IN2(U5795_n1), .QN(WX11162) );
  INVX0 U5796_U2 ( .INP(WX11097), .ZN(U5796_n1) );
  NOR2X0 U5796_U1 ( .IN1(n9197), .IN2(U5796_n1), .QN(WX11160) );
  INVX0 U5797_U2 ( .INP(WX11095), .ZN(U5797_n1) );
  NOR2X0 U5797_U1 ( .IN1(n9197), .IN2(U5797_n1), .QN(WX11158) );
  INVX0 U5798_U2 ( .INP(WX11093), .ZN(U5798_n1) );
  NOR2X0 U5798_U1 ( .IN1(n9197), .IN2(U5798_n1), .QN(WX11156) );
  INVX0 U5799_U2 ( .INP(WX11091), .ZN(U5799_n1) );
  NOR2X0 U5799_U1 ( .IN1(n9197), .IN2(U5799_n1), .QN(WX11154) );
  INVX0 U5800_U2 ( .INP(WX11089), .ZN(U5800_n1) );
  NOR2X0 U5800_U1 ( .IN1(n9197), .IN2(U5800_n1), .QN(WX11152) );
  INVX0 U5801_U2 ( .INP(WX11087), .ZN(U5801_n1) );
  NOR2X0 U5801_U1 ( .IN1(n9197), .IN2(U5801_n1), .QN(WX11150) );
  INVX0 U5802_U2 ( .INP(WX11085), .ZN(U5802_n1) );
  NOR2X0 U5802_U1 ( .IN1(n9198), .IN2(U5802_n1), .QN(WX11148) );
  INVX0 U5803_U2 ( .INP(WX11083), .ZN(U5803_n1) );
  NOR2X0 U5803_U1 ( .IN1(n9198), .IN2(U5803_n1), .QN(WX11146) );
  INVX0 U5804_U2 ( .INP(WX11081), .ZN(U5804_n1) );
  NOR2X0 U5804_U1 ( .IN1(n9198), .IN2(U5804_n1), .QN(WX11144) );
  INVX0 U5805_U2 ( .INP(WX11079), .ZN(U5805_n1) );
  NOR2X0 U5805_U1 ( .IN1(n9198), .IN2(U5805_n1), .QN(WX11142) );
  INVX0 U5806_U2 ( .INP(WX11077), .ZN(U5806_n1) );
  NOR2X0 U5806_U1 ( .IN1(n9198), .IN2(U5806_n1), .QN(WX11140) );
  INVX0 U5807_U2 ( .INP(WX11075), .ZN(U5807_n1) );
  NOR2X0 U5807_U1 ( .IN1(n9198), .IN2(U5807_n1), .QN(WX11138) );
  INVX0 U5808_U2 ( .INP(WX11073), .ZN(U5808_n1) );
  NOR2X0 U5808_U1 ( .IN1(n9198), .IN2(U5808_n1), .QN(WX11136) );
  INVX0 U5809_U2 ( .INP(WX11071), .ZN(U5809_n1) );
  NOR2X0 U5809_U1 ( .IN1(n9198), .IN2(U5809_n1), .QN(WX11134) );
  INVX0 U5810_U2 ( .INP(test_so93), .ZN(U5810_n1) );
  NOR2X0 U5810_U1 ( .IN1(n9198), .IN2(U5810_n1), .QN(WX11132) );
  INVX0 U5811_U2 ( .INP(WX11067), .ZN(U5811_n1) );
  NOR2X0 U5811_U1 ( .IN1(n9198), .IN2(U5811_n1), .QN(WX11130) );
  INVX0 U5812_U2 ( .INP(WX11065), .ZN(U5812_n1) );
  NOR2X0 U5812_U1 ( .IN1(n9198), .IN2(U5812_n1), .QN(WX11128) );
  INVX0 U5813_U2 ( .INP(WX11063), .ZN(U5813_n1) );
  NOR2X0 U5813_U1 ( .IN1(n9198), .IN2(U5813_n1), .QN(WX11126) );
  INVX0 U5814_U2 ( .INP(WX11061), .ZN(U5814_n1) );
  NOR2X0 U5814_U1 ( .IN1(n9198), .IN2(U5814_n1), .QN(WX11124) );
  INVX0 U5815_U2 ( .INP(WX11059), .ZN(U5815_n1) );
  NOR2X0 U5815_U1 ( .IN1(n9199), .IN2(U5815_n1), .QN(WX11122) );
  INVX0 U5816_U2 ( .INP(WX11057), .ZN(U5816_n1) );
  NOR2X0 U5816_U1 ( .IN1(n9199), .IN2(U5816_n1), .QN(WX11120) );
  INVX0 U5817_U2 ( .INP(WX11055), .ZN(U5817_n1) );
  NOR2X0 U5817_U1 ( .IN1(n9199), .IN2(U5817_n1), .QN(WX11118) );
  INVX0 U5818_U2 ( .INP(WX11053), .ZN(U5818_n1) );
  NOR2X0 U5818_U1 ( .IN1(n9199), .IN2(U5818_n1), .QN(WX11116) );
  INVX0 U5819_U2 ( .INP(WX11051), .ZN(U5819_n1) );
  NOR2X0 U5819_U1 ( .IN1(n9199), .IN2(U5819_n1), .QN(WX11114) );
  INVX0 U5820_U2 ( .INP(WX11049), .ZN(U5820_n1) );
  NOR2X0 U5820_U1 ( .IN1(n9199), .IN2(U5820_n1), .QN(WX11112) );
  INVX0 U5821_U2 ( .INP(WX11047), .ZN(U5821_n1) );
  NOR2X0 U5821_U1 ( .IN1(n9199), .IN2(U5821_n1), .QN(WX11110) );
  INVX0 U5822_U2 ( .INP(WX11045), .ZN(U5822_n1) );
  NOR2X0 U5822_U1 ( .IN1(n9199), .IN2(U5822_n1), .QN(WX11108) );
  INVX0 U5823_U2 ( .INP(WX11043), .ZN(U5823_n1) );
  NOR2X0 U5823_U1 ( .IN1(n9199), .IN2(U5823_n1), .QN(WX11106) );
  INVX0 U5824_U2 ( .INP(WX11041), .ZN(U5824_n1) );
  NOR2X0 U5824_U1 ( .IN1(n9199), .IN2(U5824_n1), .QN(WX11104) );
  INVX0 U5825_U2 ( .INP(WX11039), .ZN(U5825_n1) );
  NOR2X0 U5825_U1 ( .IN1(n9199), .IN2(U5825_n1), .QN(WX11102) );
  INVX0 U5826_U2 ( .INP(WX11037), .ZN(U5826_n1) );
  NOR2X0 U5826_U1 ( .IN1(n9199), .IN2(U5826_n1), .QN(WX11100) );
  INVX0 U5827_U2 ( .INP(test_so92), .ZN(U5827_n1) );
  NOR2X0 U5827_U1 ( .IN1(n9199), .IN2(U5827_n1), .QN(WX11098) );
  INVX0 U5828_U2 ( .INP(WX11033), .ZN(U5828_n1) );
  NOR2X0 U5828_U1 ( .IN1(n9200), .IN2(U5828_n1), .QN(WX11096) );
  INVX0 U5829_U2 ( .INP(WX11031), .ZN(U5829_n1) );
  NOR2X0 U5829_U1 ( .IN1(n9200), .IN2(U5829_n1), .QN(WX11094) );
  INVX0 U5830_U2 ( .INP(WX11029), .ZN(U5830_n1) );
  NOR2X0 U5830_U1 ( .IN1(n9200), .IN2(U5830_n1), .QN(WX11092) );
  INVX0 U5831_U2 ( .INP(WX11027), .ZN(U5831_n1) );
  NOR2X0 U5831_U1 ( .IN1(n9200), .IN2(U5831_n1), .QN(WX11090) );
  INVX0 U5832_U2 ( .INP(WX11025), .ZN(U5832_n1) );
  NOR2X0 U5832_U1 ( .IN1(n9200), .IN2(U5832_n1), .QN(WX11088) );
  INVX0 U5833_U2 ( .INP(WX11023), .ZN(U5833_n1) );
  NOR2X0 U5833_U1 ( .IN1(n9200), .IN2(U5833_n1), .QN(WX11086) );
  INVX0 U5834_U2 ( .INP(WX11021), .ZN(U5834_n1) );
  NOR2X0 U5834_U1 ( .IN1(n9200), .IN2(U5834_n1), .QN(WX11084) );
  INVX0 U5835_U2 ( .INP(WX9886), .ZN(U5835_n1) );
  NOR2X0 U5835_U1 ( .IN1(n9200), .IN2(U5835_n1), .QN(WX9949) );
  INVX0 U5836_U2 ( .INP(WX9884), .ZN(U5836_n1) );
  NOR2X0 U5836_U1 ( .IN1(n9200), .IN2(U5836_n1), .QN(WX9947) );
  INVX0 U5837_U2 ( .INP(WX9882), .ZN(U5837_n1) );
  NOR2X0 U5837_U1 ( .IN1(n9200), .IN2(U5837_n1), .QN(WX9945) );
  INVX0 U5838_U2 ( .INP(WX9880), .ZN(U5838_n1) );
  NOR2X0 U5838_U1 ( .IN1(n9200), .IN2(U5838_n1), .QN(WX9943) );
  INVX0 U5839_U2 ( .INP(WX9878), .ZN(U5839_n1) );
  NOR2X0 U5839_U1 ( .IN1(n9200), .IN2(U5839_n1), .QN(WX9941) );
  INVX0 U5840_U2 ( .INP(WX9876), .ZN(U5840_n1) );
  NOR2X0 U5840_U1 ( .IN1(n9200), .IN2(U5840_n1), .QN(WX9939) );
  INVX0 U5841_U2 ( .INP(WX9874), .ZN(U5841_n1) );
  NOR2X0 U5841_U1 ( .IN1(n9201), .IN2(U5841_n1), .QN(WX9937) );
  INVX0 U5842_U2 ( .INP(WX9872), .ZN(U5842_n1) );
  NOR2X0 U5842_U1 ( .IN1(n9201), .IN2(U5842_n1), .QN(WX9935) );
  INVX0 U5843_U2 ( .INP(WX9870), .ZN(U5843_n1) );
  NOR2X0 U5843_U1 ( .IN1(n9201), .IN2(U5843_n1), .QN(WX9933) );
  INVX0 U5844_U2 ( .INP(WX9868), .ZN(U5844_n1) );
  NOR2X0 U5844_U1 ( .IN1(n9201), .IN2(U5844_n1), .QN(WX9931) );
  INVX0 U5845_U2 ( .INP(WX9866), .ZN(U5845_n1) );
  NOR2X0 U5845_U1 ( .IN1(n9201), .IN2(U5845_n1), .QN(WX9929) );
  INVX0 U5846_U2 ( .INP(WX9864), .ZN(U5846_n1) );
  NOR2X0 U5846_U1 ( .IN1(n9201), .IN2(U5846_n1), .QN(WX9927) );
  INVX0 U5847_U2 ( .INP(WX9862), .ZN(U5847_n1) );
  NOR2X0 U5847_U1 ( .IN1(n9201), .IN2(U5847_n1), .QN(WX9925) );
  INVX0 U5848_U2 ( .INP(WX9860), .ZN(U5848_n1) );
  NOR2X0 U5848_U1 ( .IN1(n9201), .IN2(U5848_n1), .QN(WX9923) );
  INVX0 U5849_U2 ( .INP(WX9858), .ZN(U5849_n1) );
  NOR2X0 U5849_U1 ( .IN1(n9201), .IN2(U5849_n1), .QN(WX9921) );
  INVX0 U5850_U2 ( .INP(WX9856), .ZN(U5850_n1) );
  NOR2X0 U5850_U1 ( .IN1(n9201), .IN2(U5850_n1), .QN(WX9919) );
  INVX0 U5851_U2 ( .INP(test_so84), .ZN(U5851_n1) );
  NOR2X0 U5851_U1 ( .IN1(n9201), .IN2(U5851_n1), .QN(WX9917) );
  INVX0 U5852_U2 ( .INP(WX9852), .ZN(U5852_n1) );
  NOR2X0 U5852_U1 ( .IN1(n9201), .IN2(U5852_n1), .QN(WX9915) );
  INVX0 U5853_U2 ( .INP(WX9850), .ZN(U5853_n1) );
  NOR2X0 U5853_U1 ( .IN1(n9201), .IN2(U5853_n1), .QN(WX9913) );
  INVX0 U5854_U2 ( .INP(WX9848), .ZN(U5854_n1) );
  NOR2X0 U5854_U1 ( .IN1(n9202), .IN2(U5854_n1), .QN(WX9911) );
  INVX0 U5855_U2 ( .INP(WX9846), .ZN(U5855_n1) );
  NOR2X0 U5855_U1 ( .IN1(n9202), .IN2(U5855_n1), .QN(WX9909) );
  INVX0 U5856_U2 ( .INP(WX9844), .ZN(U5856_n1) );
  NOR2X0 U5856_U1 ( .IN1(n9202), .IN2(U5856_n1), .QN(WX9907) );
  INVX0 U5857_U2 ( .INP(WX9842), .ZN(U5857_n1) );
  NOR2X0 U5857_U1 ( .IN1(n9202), .IN2(U5857_n1), .QN(WX9905) );
  INVX0 U5858_U2 ( .INP(WX9840), .ZN(U5858_n1) );
  NOR2X0 U5858_U1 ( .IN1(n9202), .IN2(U5858_n1), .QN(WX9903) );
  INVX0 U5859_U2 ( .INP(WX9838), .ZN(U5859_n1) );
  NOR2X0 U5859_U1 ( .IN1(n9202), .IN2(U5859_n1), .QN(WX9901) );
  INVX0 U5860_U2 ( .INP(WX9836), .ZN(U5860_n1) );
  NOR2X0 U5860_U1 ( .IN1(n9202), .IN2(U5860_n1), .QN(WX9899) );
  INVX0 U5861_U2 ( .INP(WX9834), .ZN(U5861_n1) );
  NOR2X0 U5861_U1 ( .IN1(n9202), .IN2(U5861_n1), .QN(WX9897) );
  INVX0 U5862_U2 ( .INP(WX9832), .ZN(U5862_n1) );
  NOR2X0 U5862_U1 ( .IN1(n9202), .IN2(U5862_n1), .QN(WX9895) );
  INVX0 U5863_U2 ( .INP(WX9830), .ZN(U5863_n1) );
  NOR2X0 U5863_U1 ( .IN1(n9202), .IN2(U5863_n1), .QN(WX9893) );
  INVX0 U5864_U2 ( .INP(WX9828), .ZN(U5864_n1) );
  NOR2X0 U5864_U1 ( .IN1(n9202), .IN2(U5864_n1), .QN(WX9891) );
  INVX0 U5865_U2 ( .INP(WX9826), .ZN(U5865_n1) );
  NOR2X0 U5865_U1 ( .IN1(n9202), .IN2(U5865_n1), .QN(WX9889) );
  INVX0 U5866_U2 ( .INP(WX9824), .ZN(U5866_n1) );
  NOR2X0 U5866_U1 ( .IN1(n9202), .IN2(U5866_n1), .QN(WX9887) );
  INVX0 U5867_U2 ( .INP(WX9822), .ZN(U5867_n1) );
  NOR2X0 U5867_U1 ( .IN1(n9203), .IN2(U5867_n1), .QN(WX9885) );
  INVX0 U5868_U2 ( .INP(test_so83), .ZN(U5868_n1) );
  NOR2X0 U5868_U1 ( .IN1(n9203), .IN2(U5868_n1), .QN(WX9883) );
  INVX0 U5869_U2 ( .INP(WX9818), .ZN(U5869_n1) );
  NOR2X0 U5869_U1 ( .IN1(n9203), .IN2(U5869_n1), .QN(WX9881) );
  INVX0 U5870_U2 ( .INP(WX9816), .ZN(U5870_n1) );
  NOR2X0 U5870_U1 ( .IN1(n9203), .IN2(U5870_n1), .QN(WX9879) );
  INVX0 U5871_U2 ( .INP(WX9814), .ZN(U5871_n1) );
  NOR2X0 U5871_U1 ( .IN1(n9203), .IN2(U5871_n1), .QN(WX9877) );
  INVX0 U5872_U2 ( .INP(WX9812), .ZN(U5872_n1) );
  NOR2X0 U5872_U1 ( .IN1(n9203), .IN2(U5872_n1), .QN(WX9875) );
  INVX0 U5873_U2 ( .INP(WX9810), .ZN(U5873_n1) );
  NOR2X0 U5873_U1 ( .IN1(n9203), .IN2(U5873_n1), .QN(WX9873) );
  INVX0 U5874_U2 ( .INP(WX9808), .ZN(U5874_n1) );
  NOR2X0 U5874_U1 ( .IN1(n9203), .IN2(U5874_n1), .QN(WX9871) );
  INVX0 U5875_U2 ( .INP(WX9806), .ZN(U5875_n1) );
  NOR2X0 U5875_U1 ( .IN1(n9203), .IN2(U5875_n1), .QN(WX9869) );
  INVX0 U5876_U2 ( .INP(WX9804), .ZN(U5876_n1) );
  NOR2X0 U5876_U1 ( .IN1(n9203), .IN2(U5876_n1), .QN(WX9867) );
  INVX0 U5877_U2 ( .INP(WX9802), .ZN(U5877_n1) );
  NOR2X0 U5877_U1 ( .IN1(n9185), .IN2(U5877_n1), .QN(WX9865) );
  INVX0 U5878_U2 ( .INP(WX9800), .ZN(U5878_n1) );
  NOR2X0 U5878_U1 ( .IN1(n9179), .IN2(U5878_n1), .QN(WX9863) );
  INVX0 U5879_U2 ( .INP(WX9798), .ZN(U5879_n1) );
  NOR2X0 U5879_U1 ( .IN1(n9179), .IN2(U5879_n1), .QN(WX9861) );
  INVX0 U5880_U2 ( .INP(WX9796), .ZN(U5880_n1) );
  NOR2X0 U5880_U1 ( .IN1(n9179), .IN2(U5880_n1), .QN(WX9859) );
  INVX0 U5881_U2 ( .INP(WX9794), .ZN(U5881_n1) );
  NOR2X0 U5881_U1 ( .IN1(n9179), .IN2(U5881_n1), .QN(WX9857) );
  INVX0 U5882_U2 ( .INP(WX9792), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(n9179), .IN2(U5882_n1), .QN(WX9855) );
  INVX0 U5883_U2 ( .INP(WX9790), .ZN(U5883_n1) );
  NOR2X0 U5883_U1 ( .IN1(n9179), .IN2(U5883_n1), .QN(WX9853) );
  INVX0 U5884_U2 ( .INP(WX9788), .ZN(U5884_n1) );
  NOR2X0 U5884_U1 ( .IN1(n9179), .IN2(U5884_n1), .QN(WX9851) );
  INVX0 U5885_U2 ( .INP(test_so82), .ZN(U5885_n1) );
  NOR2X0 U5885_U1 ( .IN1(n9179), .IN2(U5885_n1), .QN(WX9849) );
  INVX0 U5886_U2 ( .INP(WX9784), .ZN(U5886_n1) );
  NOR2X0 U5886_U1 ( .IN1(n9180), .IN2(U5886_n1), .QN(WX9847) );
  INVX0 U5887_U2 ( .INP(WX9782), .ZN(U5887_n1) );
  NOR2X0 U5887_U1 ( .IN1(n9180), .IN2(U5887_n1), .QN(WX9845) );
  INVX0 U5888_U2 ( .INP(WX9780), .ZN(U5888_n1) );
  NOR2X0 U5888_U1 ( .IN1(n9180), .IN2(U5888_n1), .QN(WX9843) );
  INVX0 U5889_U2 ( .INP(WX9778), .ZN(U5889_n1) );
  NOR2X0 U5889_U1 ( .IN1(n9180), .IN2(U5889_n1), .QN(WX9841) );
  INVX0 U5890_U2 ( .INP(WX9776), .ZN(U5890_n1) );
  NOR2X0 U5890_U1 ( .IN1(n9180), .IN2(U5890_n1), .QN(WX9839) );
  INVX0 U5891_U2 ( .INP(WX9774), .ZN(U5891_n1) );
  NOR2X0 U5891_U1 ( .IN1(n9180), .IN2(U5891_n1), .QN(WX9837) );
  INVX0 U5892_U2 ( .INP(WX9772), .ZN(U5892_n1) );
  NOR2X0 U5892_U1 ( .IN1(n9180), .IN2(U5892_n1), .QN(WX9835) );
  INVX0 U5893_U2 ( .INP(WX9770), .ZN(U5893_n1) );
  NOR2X0 U5893_U1 ( .IN1(n9180), .IN2(U5893_n1), .QN(WX9833) );
  INVX0 U5894_U2 ( .INP(WX9768), .ZN(U5894_n1) );
  NOR2X0 U5894_U1 ( .IN1(n9180), .IN2(U5894_n1), .QN(WX9831) );
  INVX0 U5895_U2 ( .INP(WX9766), .ZN(U5895_n1) );
  NOR2X0 U5895_U1 ( .IN1(n9180), .IN2(U5895_n1), .QN(WX9829) );
  INVX0 U5896_U2 ( .INP(WX9764), .ZN(U5896_n1) );
  NOR2X0 U5896_U1 ( .IN1(n9180), .IN2(U5896_n1), .QN(WX9827) );
  INVX0 U5897_U2 ( .INP(WX9762), .ZN(U5897_n1) );
  NOR2X0 U5897_U1 ( .IN1(n9180), .IN2(U5897_n1), .QN(WX9825) );
  INVX0 U5898_U2 ( .INP(WX9760), .ZN(U5898_n1) );
  NOR2X0 U5898_U1 ( .IN1(n9180), .IN2(U5898_n1), .QN(WX9823) );
  INVX0 U5899_U2 ( .INP(WX9758), .ZN(U5899_n1) );
  NOR2X0 U5899_U1 ( .IN1(n9181), .IN2(U5899_n1), .QN(WX9821) );
  INVX0 U5900_U2 ( .INP(WX9756), .ZN(U5900_n1) );
  NOR2X0 U5900_U1 ( .IN1(n9181), .IN2(U5900_n1), .QN(WX9819) );
  INVX0 U5901_U2 ( .INP(WX9754), .ZN(U5901_n1) );
  NOR2X0 U5901_U1 ( .IN1(n9181), .IN2(U5901_n1), .QN(WX9817) );
  INVX0 U5902_U2 ( .INP(test_so81), .ZN(U5902_n1) );
  NOR2X0 U5902_U1 ( .IN1(n9181), .IN2(U5902_n1), .QN(WX9815) );
  INVX0 U5903_U2 ( .INP(WX9750), .ZN(U5903_n1) );
  NOR2X0 U5903_U1 ( .IN1(n9181), .IN2(U5903_n1), .QN(WX9813) );
  INVX0 U5904_U2 ( .INP(WX9748), .ZN(U5904_n1) );
  NOR2X0 U5904_U1 ( .IN1(n9181), .IN2(U5904_n1), .QN(WX9811) );
  INVX0 U5905_U2 ( .INP(WX9746), .ZN(U5905_n1) );
  NOR2X0 U5905_U1 ( .IN1(n9181), .IN2(U5905_n1), .QN(WX9809) );
  INVX0 U5906_U2 ( .INP(WX9744), .ZN(U5906_n1) );
  NOR2X0 U5906_U1 ( .IN1(n9181), .IN2(U5906_n1), .QN(WX9807) );
  INVX0 U5907_U2 ( .INP(WX9742), .ZN(U5907_n1) );
  NOR2X0 U5907_U1 ( .IN1(n9181), .IN2(U5907_n1), .QN(WX9805) );
  INVX0 U5908_U2 ( .INP(WX9740), .ZN(U5908_n1) );
  NOR2X0 U5908_U1 ( .IN1(n9181), .IN2(U5908_n1), .QN(WX9803) );
  INVX0 U5909_U2 ( .INP(WX9738), .ZN(U5909_n1) );
  NOR2X0 U5909_U1 ( .IN1(n9181), .IN2(U5909_n1), .QN(WX9801) );
  INVX0 U5910_U2 ( .INP(WX9736), .ZN(U5910_n1) );
  NOR2X0 U5910_U1 ( .IN1(n9181), .IN2(U5910_n1), .QN(WX9799) );
  INVX0 U5911_U2 ( .INP(WX9734), .ZN(U5911_n1) );
  NOR2X0 U5911_U1 ( .IN1(n9181), .IN2(U5911_n1), .QN(WX9797) );
  INVX0 U5912_U2 ( .INP(WX9732), .ZN(U5912_n1) );
  NOR2X0 U5912_U1 ( .IN1(n9182), .IN2(U5912_n1), .QN(WX9795) );
  INVX0 U5913_U2 ( .INP(WX9730), .ZN(U5913_n1) );
  NOR2X0 U5913_U1 ( .IN1(n9182), .IN2(U5913_n1), .QN(WX9793) );
  INVX0 U5914_U2 ( .INP(WX9728), .ZN(U5914_n1) );
  NOR2X0 U5914_U1 ( .IN1(n9182), .IN2(U5914_n1), .QN(WX9791) );
  INVX0 U5915_U2 ( .INP(WX8593), .ZN(U5915_n1) );
  NOR2X0 U5915_U1 ( .IN1(n9182), .IN2(U5915_n1), .QN(WX8656) );
  INVX0 U5916_U2 ( .INP(WX8591), .ZN(U5916_n1) );
  NOR2X0 U5916_U1 ( .IN1(n9182), .IN2(U5916_n1), .QN(WX8654) );
  INVX0 U5917_U2 ( .INP(WX8589), .ZN(U5917_n1) );
  NOR2X0 U5917_U1 ( .IN1(n9182), .IN2(U5917_n1), .QN(WX8652) );
  INVX0 U5918_U2 ( .INP(WX8587), .ZN(U5918_n1) );
  NOR2X0 U5918_U1 ( .IN1(n9182), .IN2(U5918_n1), .QN(WX8650) );
  INVX0 U5919_U2 ( .INP(WX8585), .ZN(U5919_n1) );
  NOR2X0 U5919_U1 ( .IN1(n9182), .IN2(U5919_n1), .QN(WX8648) );
  INVX0 U5920_U2 ( .INP(WX8583), .ZN(U5920_n1) );
  NOR2X0 U5920_U1 ( .IN1(n9182), .IN2(U5920_n1), .QN(WX8646) );
  INVX0 U5921_U2 ( .INP(WX8581), .ZN(U5921_n1) );
  NOR2X0 U5921_U1 ( .IN1(n9182), .IN2(U5921_n1), .QN(WX8644) );
  INVX0 U5922_U2 ( .INP(WX8579), .ZN(U5922_n1) );
  NOR2X0 U5922_U1 ( .IN1(n9182), .IN2(U5922_n1), .QN(WX8642) );
  INVX0 U5923_U2 ( .INP(WX8577), .ZN(U5923_n1) );
  NOR2X0 U5923_U1 ( .IN1(n9182), .IN2(U5923_n1), .QN(WX8640) );
  INVX0 U5924_U2 ( .INP(WX8575), .ZN(U5924_n1) );
  NOR2X0 U5924_U1 ( .IN1(n9182), .IN2(U5924_n1), .QN(WX8638) );
  INVX0 U5925_U2 ( .INP(WX8573), .ZN(U5925_n1) );
  NOR2X0 U5925_U1 ( .IN1(n9183), .IN2(U5925_n1), .QN(WX8636) );
  INVX0 U5926_U2 ( .INP(test_so73), .ZN(U5926_n1) );
  NOR2X0 U5926_U1 ( .IN1(n9183), .IN2(U5926_n1), .QN(WX8634) );
  INVX0 U5927_U2 ( .INP(WX8569), .ZN(U5927_n1) );
  NOR2X0 U5927_U1 ( .IN1(n9183), .IN2(U5927_n1), .QN(WX8632) );
  INVX0 U5928_U2 ( .INP(WX8567), .ZN(U5928_n1) );
  NOR2X0 U5928_U1 ( .IN1(n9183), .IN2(U5928_n1), .QN(WX8630) );
  INVX0 U5929_U2 ( .INP(WX8565), .ZN(U5929_n1) );
  NOR2X0 U5929_U1 ( .IN1(n9183), .IN2(U5929_n1), .QN(WX8628) );
  INVX0 U5930_U2 ( .INP(WX8563), .ZN(U5930_n1) );
  NOR2X0 U5930_U1 ( .IN1(n9183), .IN2(U5930_n1), .QN(WX8626) );
  INVX0 U5931_U2 ( .INP(WX8561), .ZN(U5931_n1) );
  NOR2X0 U5931_U1 ( .IN1(n9183), .IN2(U5931_n1), .QN(WX8624) );
  INVX0 U5932_U2 ( .INP(WX8559), .ZN(U5932_n1) );
  NOR2X0 U5932_U1 ( .IN1(n9183), .IN2(U5932_n1), .QN(WX8622) );
  INVX0 U5933_U2 ( .INP(WX8557), .ZN(U5933_n1) );
  NOR2X0 U5933_U1 ( .IN1(n9183), .IN2(U5933_n1), .QN(WX8620) );
  INVX0 U5934_U2 ( .INP(WX8555), .ZN(U5934_n1) );
  NOR2X0 U5934_U1 ( .IN1(n9183), .IN2(U5934_n1), .QN(WX8618) );
  INVX0 U5935_U2 ( .INP(WX8553), .ZN(U5935_n1) );
  NOR2X0 U5935_U1 ( .IN1(n9183), .IN2(U5935_n1), .QN(WX8616) );
  INVX0 U5936_U2 ( .INP(WX8551), .ZN(U5936_n1) );
  NOR2X0 U5936_U1 ( .IN1(n9183), .IN2(U5936_n1), .QN(WX8614) );
  INVX0 U5937_U2 ( .INP(WX8549), .ZN(U5937_n1) );
  NOR2X0 U5937_U1 ( .IN1(n9183), .IN2(U5937_n1), .QN(WX8612) );
  INVX0 U5938_U2 ( .INP(WX8547), .ZN(U5938_n1) );
  NOR2X0 U5938_U1 ( .IN1(n9184), .IN2(U5938_n1), .QN(WX8610) );
  INVX0 U5939_U2 ( .INP(WX8545), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n9184), .IN2(U5939_n1), .QN(WX8608) );
  INVX0 U5940_U2 ( .INP(WX8543), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n9184), .IN2(U5940_n1), .QN(WX8606) );
  INVX0 U5941_U2 ( .INP(WX8541), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n9184), .IN2(U5941_n1), .QN(WX8604) );
  INVX0 U5942_U2 ( .INP(WX8539), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n9184), .IN2(U5942_n1), .QN(WX8602) );
  INVX0 U5943_U2 ( .INP(test_so72), .ZN(U5943_n1) );
  NOR2X0 U5943_U1 ( .IN1(n9184), .IN2(U5943_n1), .QN(WX8600) );
  INVX0 U5944_U2 ( .INP(WX8535), .ZN(U5944_n1) );
  NOR2X0 U5944_U1 ( .IN1(n9184), .IN2(U5944_n1), .QN(WX8598) );
  INVX0 U5945_U2 ( .INP(WX8533), .ZN(U5945_n1) );
  NOR2X0 U5945_U1 ( .IN1(n9184), .IN2(U5945_n1), .QN(WX8596) );
  INVX0 U5946_U2 ( .INP(WX8531), .ZN(U5946_n1) );
  NOR2X0 U5946_U1 ( .IN1(n9184), .IN2(U5946_n1), .QN(WX8594) );
  INVX0 U5947_U2 ( .INP(WX8529), .ZN(U5947_n1) );
  NOR2X0 U5947_U1 ( .IN1(n9184), .IN2(U5947_n1), .QN(WX8592) );
  INVX0 U5948_U2 ( .INP(WX8527), .ZN(U5948_n1) );
  NOR2X0 U5948_U1 ( .IN1(n9184), .IN2(U5948_n1), .QN(WX8590) );
  INVX0 U5949_U2 ( .INP(WX8525), .ZN(U5949_n1) );
  NOR2X0 U5949_U1 ( .IN1(n9184), .IN2(U5949_n1), .QN(WX8588) );
  INVX0 U5950_U2 ( .INP(WX8523), .ZN(U5950_n1) );
  NOR2X0 U5950_U1 ( .IN1(n9184), .IN2(U5950_n1), .QN(WX8586) );
  INVX0 U5951_U2 ( .INP(WX8521), .ZN(U5951_n1) );
  NOR2X0 U5951_U1 ( .IN1(n9185), .IN2(U5951_n1), .QN(WX8584) );
  INVX0 U5952_U2 ( .INP(WX8519), .ZN(U5952_n1) );
  NOR2X0 U5952_U1 ( .IN1(n9185), .IN2(U5952_n1), .QN(WX8582) );
  INVX0 U5953_U2 ( .INP(WX8517), .ZN(U5953_n1) );
  NOR2X0 U5953_U1 ( .IN1(n9185), .IN2(U5953_n1), .QN(WX8580) );
  INVX0 U5954_U2 ( .INP(WX8515), .ZN(U5954_n1) );
  NOR2X0 U5954_U1 ( .IN1(n9185), .IN2(U5954_n1), .QN(WX8578) );
  INVX0 U5955_U2 ( .INP(WX8513), .ZN(U5955_n1) );
  NOR2X0 U5955_U1 ( .IN1(n9185), .IN2(U5955_n1), .QN(WX8576) );
  INVX0 U5956_U2 ( .INP(WX8511), .ZN(U5956_n1) );
  NOR2X0 U5956_U1 ( .IN1(n9185), .IN2(U5956_n1), .QN(WX8574) );
  INVX0 U5957_U2 ( .INP(WX8509), .ZN(U5957_n1) );
  NOR2X0 U5957_U1 ( .IN1(n9185), .IN2(U5957_n1), .QN(WX8572) );
  INVX0 U5958_U2 ( .INP(WX8507), .ZN(U5958_n1) );
  NOR2X0 U5958_U1 ( .IN1(n9185), .IN2(U5958_n1), .QN(WX8570) );
  INVX0 U5959_U2 ( .INP(WX8505), .ZN(U5959_n1) );
  NOR2X0 U5959_U1 ( .IN1(n9185), .IN2(U5959_n1), .QN(WX8568) );
  INVX0 U5960_U2 ( .INP(test_so71), .ZN(U5960_n1) );
  NOR2X0 U5960_U1 ( .IN1(n9185), .IN2(U5960_n1), .QN(WX8566) );
  INVX0 U5961_U2 ( .INP(WX8501), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n9185), .IN2(U5961_n1), .QN(WX8564) );
  INVX0 U5962_U2 ( .INP(WX8499), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n9185), .IN2(U5962_n1), .QN(WX8562) );
  INVX0 U5963_U2 ( .INP(WX8497), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n9186), .IN2(U5963_n1), .QN(WX8560) );
  INVX0 U5964_U2 ( .INP(WX8495), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n9186), .IN2(U5964_n1), .QN(WX8558) );
  INVX0 U5965_U2 ( .INP(WX8493), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n9186), .IN2(U5965_n1), .QN(WX8556) );
  INVX0 U5966_U2 ( .INP(WX8491), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n9186), .IN2(U5966_n1), .QN(WX8554) );
  INVX0 U5967_U2 ( .INP(WX8489), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n9186), .IN2(U5967_n1), .QN(WX8552) );
  INVX0 U5968_U2 ( .INP(WX8487), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n9186), .IN2(U5968_n1), .QN(WX8550) );
  INVX0 U5969_U2 ( .INP(WX8485), .ZN(U5969_n1) );
  NOR2X0 U5969_U1 ( .IN1(n9186), .IN2(U5969_n1), .QN(WX8548) );
  INVX0 U5970_U2 ( .INP(WX8483), .ZN(U5970_n1) );
  NOR2X0 U5970_U1 ( .IN1(n9186), .IN2(U5970_n1), .QN(WX8546) );
  INVX0 U5971_U2 ( .INP(WX8481), .ZN(U5971_n1) );
  NOR2X0 U5971_U1 ( .IN1(n9186), .IN2(U5971_n1), .QN(WX8544) );
  INVX0 U5972_U2 ( .INP(WX8479), .ZN(U5972_n1) );
  NOR2X0 U5972_U1 ( .IN1(n9186), .IN2(U5972_n1), .QN(WX8542) );
  INVX0 U5973_U2 ( .INP(WX8477), .ZN(U5973_n1) );
  NOR2X0 U5973_U1 ( .IN1(n9186), .IN2(U5973_n1), .QN(WX8540) );
  INVX0 U5974_U2 ( .INP(WX8475), .ZN(U5974_n1) );
  NOR2X0 U5974_U1 ( .IN1(n9186), .IN2(U5974_n1), .QN(WX8538) );
  INVX0 U5975_U2 ( .INP(WX8473), .ZN(U5975_n1) );
  NOR2X0 U5975_U1 ( .IN1(n9186), .IN2(U5975_n1), .QN(WX8536) );
  INVX0 U5976_U2 ( .INP(WX8471), .ZN(U5976_n1) );
  NOR2X0 U5976_U1 ( .IN1(n9187), .IN2(U5976_n1), .QN(WX8534) );
  INVX0 U5977_U2 ( .INP(test_so70), .ZN(U5977_n1) );
  NOR2X0 U5977_U1 ( .IN1(n9187), .IN2(U5977_n1), .QN(WX8532) );
  INVX0 U5978_U2 ( .INP(WX8467), .ZN(U5978_n1) );
  NOR2X0 U5978_U1 ( .IN1(n9187), .IN2(U5978_n1), .QN(WX8530) );
  INVX0 U5979_U2 ( .INP(WX8465), .ZN(U5979_n1) );
  NOR2X0 U5979_U1 ( .IN1(n9187), .IN2(U5979_n1), .QN(WX8528) );
  INVX0 U5980_U2 ( .INP(WX8463), .ZN(U5980_n1) );
  NOR2X0 U5980_U1 ( .IN1(n9187), .IN2(U5980_n1), .QN(WX8526) );
  INVX0 U5981_U2 ( .INP(WX8461), .ZN(U5981_n1) );
  NOR2X0 U5981_U1 ( .IN1(n9187), .IN2(U5981_n1), .QN(WX8524) );
  INVX0 U5982_U2 ( .INP(WX8459), .ZN(U5982_n1) );
  NOR2X0 U5982_U1 ( .IN1(n9187), .IN2(U5982_n1), .QN(WX8522) );
  INVX0 U5983_U2 ( .INP(WX8457), .ZN(U5983_n1) );
  NOR2X0 U5983_U1 ( .IN1(n9187), .IN2(U5983_n1), .QN(WX8520) );
  INVX0 U5984_U2 ( .INP(WX8455), .ZN(U5984_n1) );
  NOR2X0 U5984_U1 ( .IN1(n9187), .IN2(U5984_n1), .QN(WX8518) );
  INVX0 U5985_U2 ( .INP(WX8453), .ZN(U5985_n1) );
  NOR2X0 U5985_U1 ( .IN1(n9187), .IN2(U5985_n1), .QN(WX8516) );
  INVX0 U5986_U2 ( .INP(WX8451), .ZN(U5986_n1) );
  NOR2X0 U5986_U1 ( .IN1(n9187), .IN2(U5986_n1), .QN(WX8514) );
  INVX0 U5987_U2 ( .INP(WX8449), .ZN(U5987_n1) );
  NOR2X0 U5987_U1 ( .IN1(n9187), .IN2(U5987_n1), .QN(WX8512) );
  INVX0 U5988_U2 ( .INP(WX8447), .ZN(U5988_n1) );
  NOR2X0 U5988_U1 ( .IN1(n9187), .IN2(U5988_n1), .QN(WX8510) );
  INVX0 U5989_U2 ( .INP(WX8445), .ZN(U5989_n1) );
  NOR2X0 U5989_U1 ( .IN1(n9188), .IN2(U5989_n1), .QN(WX8508) );
  INVX0 U5990_U2 ( .INP(WX8443), .ZN(U5990_n1) );
  NOR2X0 U5990_U1 ( .IN1(n9188), .IN2(U5990_n1), .QN(WX8506) );
  INVX0 U5991_U2 ( .INP(WX8441), .ZN(U5991_n1) );
  NOR2X0 U5991_U1 ( .IN1(n9188), .IN2(U5991_n1), .QN(WX8504) );
  INVX0 U5992_U2 ( .INP(WX8439), .ZN(U5992_n1) );
  NOR2X0 U5992_U1 ( .IN1(n9188), .IN2(U5992_n1), .QN(WX8502) );
  INVX0 U5993_U2 ( .INP(WX8437), .ZN(U5993_n1) );
  NOR2X0 U5993_U1 ( .IN1(n9188), .IN2(U5993_n1), .QN(WX8500) );
  INVX0 U5994_U2 ( .INP(test_so69), .ZN(U5994_n1) );
  NOR2X0 U5994_U1 ( .IN1(n9188), .IN2(U5994_n1), .QN(WX8498) );
  INVX0 U5995_U2 ( .INP(WX7300), .ZN(U5995_n1) );
  NOR2X0 U5995_U1 ( .IN1(n9188), .IN2(U5995_n1), .QN(WX7363) );
  INVX0 U5996_U2 ( .INP(WX7298), .ZN(U5996_n1) );
  NOR2X0 U5996_U1 ( .IN1(n9188), .IN2(U5996_n1), .QN(WX7361) );
  INVX0 U5997_U2 ( .INP(WX7296), .ZN(U5997_n1) );
  NOR2X0 U5997_U1 ( .IN1(n9188), .IN2(U5997_n1), .QN(WX7359) );
  INVX0 U5998_U2 ( .INP(WX7294), .ZN(U5998_n1) );
  NOR2X0 U5998_U1 ( .IN1(n9188), .IN2(U5998_n1), .QN(WX7357) );
  INVX0 U5999_U2 ( .INP(WX7292), .ZN(U5999_n1) );
  NOR2X0 U5999_U1 ( .IN1(n9188), .IN2(U5999_n1), .QN(WX7355) );
  INVX0 U6000_U2 ( .INP(WX7290), .ZN(U6000_n1) );
  NOR2X0 U6000_U1 ( .IN1(n9188), .IN2(U6000_n1), .QN(WX7353) );
  INVX0 U6001_U2 ( .INP(test_so62), .ZN(U6001_n1) );
  NOR2X0 U6001_U1 ( .IN1(n9188), .IN2(U6001_n1), .QN(WX7351) );
  INVX0 U6002_U2 ( .INP(WX7286), .ZN(U6002_n1) );
  NOR2X0 U6002_U1 ( .IN1(n9189), .IN2(U6002_n1), .QN(WX7349) );
  INVX0 U6003_U2 ( .INP(WX7284), .ZN(U6003_n1) );
  NOR2X0 U6003_U1 ( .IN1(n9189), .IN2(U6003_n1), .QN(WX7347) );
  INVX0 U6004_U2 ( .INP(WX7282), .ZN(U6004_n1) );
  NOR2X0 U6004_U1 ( .IN1(n9189), .IN2(U6004_n1), .QN(WX7345) );
  INVX0 U6005_U2 ( .INP(WX7280), .ZN(U6005_n1) );
  NOR2X0 U6005_U1 ( .IN1(n9189), .IN2(U6005_n1), .QN(WX7343) );
  INVX0 U6006_U2 ( .INP(WX7278), .ZN(U6006_n1) );
  NOR2X0 U6006_U1 ( .IN1(n9189), .IN2(U6006_n1), .QN(WX7341) );
  INVX0 U6007_U2 ( .INP(WX7276), .ZN(U6007_n1) );
  NOR2X0 U6007_U1 ( .IN1(n9189), .IN2(U6007_n1), .QN(WX7339) );
  INVX0 U6008_U2 ( .INP(WX7274), .ZN(U6008_n1) );
  NOR2X0 U6008_U1 ( .IN1(n9189), .IN2(U6008_n1), .QN(WX7337) );
  INVX0 U6009_U2 ( .INP(WX7272), .ZN(U6009_n1) );
  NOR2X0 U6009_U1 ( .IN1(n9189), .IN2(U6009_n1), .QN(WX7335) );
  INVX0 U6010_U2 ( .INP(WX7270), .ZN(U6010_n1) );
  NOR2X0 U6010_U1 ( .IN1(n9189), .IN2(U6010_n1), .QN(WX7333) );
  INVX0 U6011_U2 ( .INP(WX7268), .ZN(U6011_n1) );
  NOR2X0 U6011_U1 ( .IN1(n9189), .IN2(U6011_n1), .QN(WX7331) );
  INVX0 U6012_U2 ( .INP(WX7266), .ZN(U6012_n1) );
  NOR2X0 U6012_U1 ( .IN1(n9189), .IN2(U6012_n1), .QN(WX7329) );
  INVX0 U6013_U2 ( .INP(WX7264), .ZN(U6013_n1) );
  NOR2X0 U6013_U1 ( .IN1(n9189), .IN2(U6013_n1), .QN(WX7327) );
  INVX0 U6014_U2 ( .INP(WX7262), .ZN(U6014_n1) );
  NOR2X0 U6014_U1 ( .IN1(n9189), .IN2(U6014_n1), .QN(WX7325) );
  INVX0 U6015_U2 ( .INP(WX7260), .ZN(U6015_n1) );
  NOR2X0 U6015_U1 ( .IN1(n9190), .IN2(U6015_n1), .QN(WX7323) );
  INVX0 U6016_U2 ( .INP(WX7258), .ZN(U6016_n1) );
  NOR2X0 U6016_U1 ( .IN1(n9190), .IN2(U6016_n1), .QN(WX7321) );
  INVX0 U6017_U2 ( .INP(WX7256), .ZN(U6017_n1) );
  NOR2X0 U6017_U1 ( .IN1(n9190), .IN2(U6017_n1), .QN(WX7319) );
  INVX0 U6018_U2 ( .INP(test_so61), .ZN(U6018_n1) );
  NOR2X0 U6018_U1 ( .IN1(n9190), .IN2(U6018_n1), .QN(WX7317) );
  INVX0 U6019_U2 ( .INP(WX7252), .ZN(U6019_n1) );
  NOR2X0 U6019_U1 ( .IN1(n9190), .IN2(U6019_n1), .QN(WX7315) );
  INVX0 U6020_U2 ( .INP(WX7250), .ZN(U6020_n1) );
  NOR2X0 U6020_U1 ( .IN1(n9190), .IN2(U6020_n1), .QN(WX7313) );
  INVX0 U6021_U2 ( .INP(WX7248), .ZN(U6021_n1) );
  NOR2X0 U6021_U1 ( .IN1(n9190), .IN2(U6021_n1), .QN(WX7311) );
  INVX0 U6022_U2 ( .INP(WX7246), .ZN(U6022_n1) );
  NOR2X0 U6022_U1 ( .IN1(n9190), .IN2(U6022_n1), .QN(WX7309) );
  INVX0 U6023_U2 ( .INP(WX7244), .ZN(U6023_n1) );
  NOR2X0 U6023_U1 ( .IN1(n9190), .IN2(U6023_n1), .QN(WX7307) );
  INVX0 U6024_U2 ( .INP(WX7242), .ZN(U6024_n1) );
  NOR2X0 U6024_U1 ( .IN1(n9190), .IN2(U6024_n1), .QN(WX7305) );
  INVX0 U6025_U2 ( .INP(WX7240), .ZN(U6025_n1) );
  NOR2X0 U6025_U1 ( .IN1(n9190), .IN2(U6025_n1), .QN(WX7303) );
  INVX0 U6026_U2 ( .INP(WX7238), .ZN(U6026_n1) );
  NOR2X0 U6026_U1 ( .IN1(n9190), .IN2(U6026_n1), .QN(WX7301) );
  INVX0 U6027_U2 ( .INP(WX7236), .ZN(U6027_n1) );
  NOR2X0 U6027_U1 ( .IN1(n9190), .IN2(U6027_n1), .QN(WX7299) );
  INVX0 U6028_U2 ( .INP(WX7234), .ZN(U6028_n1) );
  NOR2X0 U6028_U1 ( .IN1(n9191), .IN2(U6028_n1), .QN(WX7297) );
  INVX0 U6029_U2 ( .INP(WX7232), .ZN(U6029_n1) );
  NOR2X0 U6029_U1 ( .IN1(n9191), .IN2(U6029_n1), .QN(WX7295) );
  INVX0 U6030_U2 ( .INP(WX7230), .ZN(U6030_n1) );
  NOR2X0 U6030_U1 ( .IN1(n9191), .IN2(U6030_n1), .QN(WX7293) );
  INVX0 U6031_U2 ( .INP(WX7228), .ZN(U6031_n1) );
  NOR2X0 U6031_U1 ( .IN1(n9191), .IN2(U6031_n1), .QN(WX7291) );
  INVX0 U6032_U2 ( .INP(WX7226), .ZN(U6032_n1) );
  NOR2X0 U6032_U1 ( .IN1(n9191), .IN2(U6032_n1), .QN(WX7289) );
  INVX0 U6033_U2 ( .INP(WX7224), .ZN(U6033_n1) );
  NOR2X0 U6033_U1 ( .IN1(n9191), .IN2(U6033_n1), .QN(WX7287) );
  INVX0 U6034_U2 ( .INP(WX7222), .ZN(U6034_n1) );
  NOR2X0 U6034_U1 ( .IN1(n9191), .IN2(U6034_n1), .QN(WX7285) );
  INVX0 U6035_U2 ( .INP(test_so60), .ZN(U6035_n1) );
  NOR2X0 U6035_U1 ( .IN1(n9191), .IN2(U6035_n1), .QN(WX7283) );
  INVX0 U6036_U2 ( .INP(WX7218), .ZN(U6036_n1) );
  NOR2X0 U6036_U1 ( .IN1(n9221), .IN2(U6036_n1), .QN(WX7281) );
  INVX0 U6037_U2 ( .INP(WX7216), .ZN(U6037_n1) );
  NOR2X0 U6037_U1 ( .IN1(n9222), .IN2(U6037_n1), .QN(WX7279) );
  INVX0 U6038_U2 ( .INP(WX7214), .ZN(U6038_n1) );
  NOR2X0 U6038_U1 ( .IN1(n9223), .IN2(U6038_n1), .QN(WX7277) );
  INVX0 U6039_U2 ( .INP(WX7212), .ZN(U6039_n1) );
  NOR2X0 U6039_U1 ( .IN1(n9221), .IN2(U6039_n1), .QN(WX7275) );
  INVX0 U6040_U2 ( .INP(WX7210), .ZN(U6040_n1) );
  NOR2X0 U6040_U1 ( .IN1(n9222), .IN2(U6040_n1), .QN(WX7273) );
  INVX0 U6041_U2 ( .INP(WX7208), .ZN(U6041_n1) );
  NOR2X0 U6041_U1 ( .IN1(n9222), .IN2(U6041_n1), .QN(WX7271) );
  INVX0 U6042_U2 ( .INP(WX7206), .ZN(U6042_n1) );
  NOR2X0 U6042_U1 ( .IN1(n9221), .IN2(U6042_n1), .QN(WX7269) );
  INVX0 U6043_U2 ( .INP(WX7204), .ZN(U6043_n1) );
  NOR2X0 U6043_U1 ( .IN1(n9221), .IN2(U6043_n1), .QN(WX7267) );
  INVX0 U6044_U2 ( .INP(WX7202), .ZN(U6044_n1) );
  NOR2X0 U6044_U1 ( .IN1(n9221), .IN2(U6044_n1), .QN(WX7265) );
  INVX0 U6045_U2 ( .INP(WX7200), .ZN(U6045_n1) );
  NOR2X0 U6045_U1 ( .IN1(n9220), .IN2(U6045_n1), .QN(WX7263) );
  INVX0 U6046_U2 ( .INP(WX7198), .ZN(U6046_n1) );
  NOR2X0 U6046_U1 ( .IN1(n9220), .IN2(U6046_n1), .QN(WX7261) );
  INVX0 U6047_U2 ( .INP(WX7196), .ZN(U6047_n1) );
  NOR2X0 U6047_U1 ( .IN1(n9220), .IN2(U6047_n1), .QN(WX7259) );
  INVX0 U6048_U2 ( .INP(WX7194), .ZN(U6048_n1) );
  NOR2X0 U6048_U1 ( .IN1(n9220), .IN2(U6048_n1), .QN(WX7257) );
  INVX0 U6049_U2 ( .INP(WX7192), .ZN(U6049_n1) );
  NOR2X0 U6049_U1 ( .IN1(n9220), .IN2(U6049_n1), .QN(WX7255) );
  INVX0 U6050_U2 ( .INP(WX7190), .ZN(U6050_n1) );
  NOR2X0 U6050_U1 ( .IN1(n9219), .IN2(U6050_n1), .QN(WX7253) );
  INVX0 U6051_U2 ( .INP(WX7188), .ZN(U6051_n1) );
  NOR2X0 U6051_U1 ( .IN1(n9220), .IN2(U6051_n1), .QN(WX7251) );
  INVX0 U6052_U2 ( .INP(test_so59), .ZN(U6052_n1) );
  NOR2X0 U6052_U1 ( .IN1(n9223), .IN2(U6052_n1), .QN(WX7249) );
  INVX0 U6053_U2 ( .INP(WX7184), .ZN(U6053_n1) );
  NOR2X0 U6053_U1 ( .IN1(n9222), .IN2(U6053_n1), .QN(WX7247) );
  INVX0 U6054_U2 ( .INP(WX7182), .ZN(U6054_n1) );
  NOR2X0 U6054_U1 ( .IN1(n9221), .IN2(U6054_n1), .QN(WX7245) );
  INVX0 U6055_U2 ( .INP(WX7180), .ZN(U6055_n1) );
  NOR2X0 U6055_U1 ( .IN1(n9223), .IN2(U6055_n1), .QN(WX7243) );
  INVX0 U6056_U2 ( .INP(WX7178), .ZN(U6056_n1) );
  NOR2X0 U6056_U1 ( .IN1(n9222), .IN2(U6056_n1), .QN(WX7241) );
  INVX0 U6057_U2 ( .INP(WX7176), .ZN(U6057_n1) );
  NOR2X0 U6057_U1 ( .IN1(n9223), .IN2(U6057_n1), .QN(WX7239) );
  INVX0 U6058_U2 ( .INP(WX7174), .ZN(U6058_n1) );
  NOR2X0 U6058_U1 ( .IN1(n9222), .IN2(U6058_n1), .QN(WX7237) );
  INVX0 U6059_U2 ( .INP(WX7172), .ZN(U6059_n1) );
  NOR2X0 U6059_U1 ( .IN1(n9222), .IN2(U6059_n1), .QN(WX7235) );
  INVX0 U6060_U2 ( .INP(WX7170), .ZN(U6060_n1) );
  NOR2X0 U6060_U1 ( .IN1(n9222), .IN2(U6060_n1), .QN(WX7233) );
  INVX0 U6061_U2 ( .INP(WX7168), .ZN(U6061_n1) );
  NOR2X0 U6061_U1 ( .IN1(n9222), .IN2(U6061_n1), .QN(WX7231) );
  INVX0 U6062_U2 ( .INP(WX7166), .ZN(U6062_n1) );
  NOR2X0 U6062_U1 ( .IN1(n9222), .IN2(U6062_n1), .QN(WX7229) );
  INVX0 U6063_U2 ( .INP(WX7164), .ZN(U6063_n1) );
  NOR2X0 U6063_U1 ( .IN1(n9221), .IN2(U6063_n1), .QN(WX7227) );
  INVX0 U6064_U2 ( .INP(WX7162), .ZN(U6064_n1) );
  NOR2X0 U6064_U1 ( .IN1(n9220), .IN2(U6064_n1), .QN(WX7225) );
  INVX0 U6065_U2 ( .INP(WX7160), .ZN(U6065_n1) );
  NOR2X0 U6065_U1 ( .IN1(n9220), .IN2(U6065_n1), .QN(WX7223) );
  INVX0 U6066_U2 ( .INP(WX7158), .ZN(U6066_n1) );
  NOR2X0 U6066_U1 ( .IN1(n9220), .IN2(U6066_n1), .QN(WX7221) );
  INVX0 U6067_U2 ( .INP(WX7156), .ZN(U6067_n1) );
  NOR2X0 U6067_U1 ( .IN1(n9220), .IN2(U6067_n1), .QN(WX7219) );
  INVX0 U6068_U2 ( .INP(WX7154), .ZN(U6068_n1) );
  NOR2X0 U6068_U1 ( .IN1(n9221), .IN2(U6068_n1), .QN(WX7217) );
  INVX0 U6069_U2 ( .INP(test_so58), .ZN(U6069_n1) );
  NOR2X0 U6069_U1 ( .IN1(n9221), .IN2(U6069_n1), .QN(WX7215) );
  INVX0 U6070_U2 ( .INP(WX7150), .ZN(U6070_n1) );
  NOR2X0 U6070_U1 ( .IN1(n9220), .IN2(U6070_n1), .QN(WX7213) );
  INVX0 U6071_U2 ( .INP(WX7148), .ZN(U6071_n1) );
  NOR2X0 U6071_U1 ( .IN1(n9221), .IN2(U6071_n1), .QN(WX7211) );
  INVX0 U6072_U2 ( .INP(WX7146), .ZN(U6072_n1) );
  NOR2X0 U6072_U1 ( .IN1(n9221), .IN2(U6072_n1), .QN(WX7209) );
  INVX0 U6073_U2 ( .INP(WX7144), .ZN(U6073_n1) );
  NOR2X0 U6073_U1 ( .IN1(n9221), .IN2(U6073_n1), .QN(WX7207) );
  INVX0 U6074_U2 ( .INP(WX7142), .ZN(U6074_n1) );
  NOR2X0 U6074_U1 ( .IN1(n9219), .IN2(U6074_n1), .QN(WX7205) );
  INVX0 U6075_U2 ( .INP(WX6007), .ZN(U6075_n1) );
  NOR2X0 U6075_U1 ( .IN1(n9222), .IN2(U6075_n1), .QN(WX6070) );
  INVX0 U6076_U2 ( .INP(test_so51), .ZN(U6076_n1) );
  NOR2X0 U6076_U1 ( .IN1(n9221), .IN2(U6076_n1), .QN(WX6068) );
  INVX0 U6077_U2 ( .INP(WX6003), .ZN(U6077_n1) );
  NOR2X0 U6077_U1 ( .IN1(n9222), .IN2(U6077_n1), .QN(WX6066) );
  INVX0 U6078_U2 ( .INP(WX6001), .ZN(U6078_n1) );
  NOR2X0 U6078_U1 ( .IN1(n9220), .IN2(U6078_n1), .QN(WX6064) );
  INVX0 U6079_U2 ( .INP(WX5999), .ZN(U6079_n1) );
  NOR2X0 U6079_U1 ( .IN1(n9223), .IN2(U6079_n1), .QN(WX6062) );
  INVX0 U6080_U2 ( .INP(WX5997), .ZN(U6080_n1) );
  NOR2X0 U6080_U1 ( .IN1(n9222), .IN2(U6080_n1), .QN(WX6060) );
  INVX0 U6081_U2 ( .INP(WX5995), .ZN(U6081_n1) );
  NOR2X0 U6081_U1 ( .IN1(n9220), .IN2(U6081_n1), .QN(WX6058) );
  INVX0 U6082_U2 ( .INP(WX5993), .ZN(U6082_n1) );
  NOR2X0 U6082_U1 ( .IN1(n9219), .IN2(U6082_n1), .QN(WX6056) );
  INVX0 U6083_U2 ( .INP(WX5991), .ZN(U6083_n1) );
  NOR2X0 U6083_U1 ( .IN1(n9219), .IN2(U6083_n1), .QN(WX6054) );
  INVX0 U6084_U2 ( .INP(WX5989), .ZN(U6084_n1) );
  NOR2X0 U6084_U1 ( .IN1(n9219), .IN2(U6084_n1), .QN(WX6052) );
  INVX0 U6085_U2 ( .INP(WX5987), .ZN(U6085_n1) );
  NOR2X0 U6085_U1 ( .IN1(n9219), .IN2(U6085_n1), .QN(WX6050) );
  INVX0 U6086_U2 ( .INP(WX5985), .ZN(U6086_n1) );
  NOR2X0 U6086_U1 ( .IN1(n9219), .IN2(U6086_n1), .QN(WX6048) );
  INVX0 U6087_U2 ( .INP(WX5983), .ZN(U6087_n1) );
  NOR2X0 U6087_U1 ( .IN1(n9219), .IN2(U6087_n1), .QN(WX6046) );
  INVX0 U6088_U2 ( .INP(WX5981), .ZN(U6088_n1) );
  NOR2X0 U6088_U1 ( .IN1(n9219), .IN2(U6088_n1), .QN(WX6044) );
  INVX0 U6089_U2 ( .INP(WX5979), .ZN(U6089_n1) );
  NOR2X0 U6089_U1 ( .IN1(n9219), .IN2(U6089_n1), .QN(WX6042) );
  INVX0 U6090_U2 ( .INP(WX5977), .ZN(U6090_n1) );
  NOR2X0 U6090_U1 ( .IN1(n9211), .IN2(U6090_n1), .QN(WX6040) );
  INVX0 U6091_U2 ( .INP(WX5975), .ZN(U6091_n1) );
  NOR2X0 U6091_U1 ( .IN1(n9211), .IN2(U6091_n1), .QN(WX6038) );
  INVX0 U6092_U2 ( .INP(WX5973), .ZN(U6092_n1) );
  NOR2X0 U6092_U1 ( .IN1(n9211), .IN2(U6092_n1), .QN(WX6036) );
  INVX0 U6093_U2 ( .INP(test_so50), .ZN(U6093_n1) );
  NOR2X0 U6093_U1 ( .IN1(n9211), .IN2(U6093_n1), .QN(WX6034) );
  INVX0 U6094_U2 ( .INP(WX5969), .ZN(U6094_n1) );
  NOR2X0 U6094_U1 ( .IN1(n9211), .IN2(U6094_n1), .QN(WX6032) );
  INVX0 U6095_U2 ( .INP(WX5967), .ZN(U6095_n1) );
  NOR2X0 U6095_U1 ( .IN1(n9211), .IN2(U6095_n1), .QN(WX6030) );
  INVX0 U6096_U2 ( .INP(WX5965), .ZN(U6096_n1) );
  NOR2X0 U6096_U1 ( .IN1(n9211), .IN2(U6096_n1), .QN(WX6028) );
  INVX0 U6097_U2 ( .INP(WX5963), .ZN(U6097_n1) );
  NOR2X0 U6097_U1 ( .IN1(n9210), .IN2(U6097_n1), .QN(WX6026) );
  INVX0 U6098_U2 ( .INP(WX5961), .ZN(U6098_n1) );
  NOR2X0 U6098_U1 ( .IN1(n9210), .IN2(U6098_n1), .QN(WX6024) );
  INVX0 U6099_U2 ( .INP(WX5959), .ZN(U6099_n1) );
  NOR2X0 U6099_U1 ( .IN1(n9210), .IN2(U6099_n1), .QN(WX6022) );
  INVX0 U6100_U2 ( .INP(WX5957), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n9210), .IN2(U6100_n1), .QN(WX6020) );
  INVX0 U6101_U2 ( .INP(WX5955), .ZN(U6101_n1) );
  NOR2X0 U6101_U1 ( .IN1(n9210), .IN2(U6101_n1), .QN(WX6018) );
  INVX0 U6102_U2 ( .INP(WX5953), .ZN(U6102_n1) );
  NOR2X0 U6102_U1 ( .IN1(n9210), .IN2(U6102_n1), .QN(WX6016) );
  INVX0 U6103_U2 ( .INP(WX5951), .ZN(U6103_n1) );
  NOR2X0 U6103_U1 ( .IN1(n9210), .IN2(U6103_n1), .QN(WX6014) );
  INVX0 U6104_U2 ( .INP(WX5949), .ZN(U6104_n1) );
  NOR2X0 U6104_U1 ( .IN1(n9210), .IN2(U6104_n1), .QN(WX6012) );
  INVX0 U6105_U2 ( .INP(WX5947), .ZN(U6105_n1) );
  NOR2X0 U6105_U1 ( .IN1(n9210), .IN2(U6105_n1), .QN(WX6010) );
  INVX0 U6106_U2 ( .INP(WX5945), .ZN(U6106_n1) );
  NOR2X0 U6106_U1 ( .IN1(n9210), .IN2(U6106_n1), .QN(WX6008) );
  INVX0 U6107_U2 ( .INP(WX5943), .ZN(U6107_n1) );
  NOR2X0 U6107_U1 ( .IN1(n9210), .IN2(U6107_n1), .QN(WX6006) );
  INVX0 U6108_U2 ( .INP(WX5941), .ZN(U6108_n1) );
  NOR2X0 U6108_U1 ( .IN1(n9210), .IN2(U6108_n1), .QN(WX6004) );
  INVX0 U6109_U2 ( .INP(WX5929), .ZN(U6109_n1) );
  NOR2X0 U6109_U1 ( .IN1(n9210), .IN2(U6109_n1), .QN(WX5992) );
  INVX0 U6110_U2 ( .INP(WX5927), .ZN(U6110_n1) );
  NOR2X0 U6110_U1 ( .IN1(n9209), .IN2(U6110_n1), .QN(WX5990) );
  INVX0 U6111_U2 ( .INP(WX5925), .ZN(U6111_n1) );
  NOR2X0 U6111_U1 ( .IN1(n9209), .IN2(U6111_n1), .QN(WX5988) );
  INVX0 U6112_U2 ( .INP(WX5923), .ZN(U6112_n1) );
  NOR2X0 U6112_U1 ( .IN1(n9209), .IN2(U6112_n1), .QN(WX5986) );
  INVX0 U6113_U2 ( .INP(WX5921), .ZN(U6113_n1) );
  NOR2X0 U6113_U1 ( .IN1(n9209), .IN2(U6113_n1), .QN(WX5984) );
  INVX0 U6114_U2 ( .INP(WX5919), .ZN(U6114_n1) );
  NOR2X0 U6114_U1 ( .IN1(n9209), .IN2(U6114_n1), .QN(WX5982) );
  INVX0 U6115_U2 ( .INP(WX5917), .ZN(U6115_n1) );
  NOR2X0 U6115_U1 ( .IN1(n9209), .IN2(U6115_n1), .QN(WX5980) );
  INVX0 U6116_U2 ( .INP(WX5915), .ZN(U6116_n1) );
  NOR2X0 U6116_U1 ( .IN1(n9209), .IN2(U6116_n1), .QN(WX5978) );
  INVX0 U6117_U2 ( .INP(WX5913), .ZN(U6117_n1) );
  NOR2X0 U6117_U1 ( .IN1(n9209), .IN2(U6117_n1), .QN(WX5976) );
  INVX0 U6118_U2 ( .INP(WX5911), .ZN(U6118_n1) );
  NOR2X0 U6118_U1 ( .IN1(n9209), .IN2(U6118_n1), .QN(WX5974) );
  INVX0 U6119_U2 ( .INP(WX5909), .ZN(U6119_n1) );
  NOR2X0 U6119_U1 ( .IN1(n9209), .IN2(U6119_n1), .QN(WX5972) );
  INVX0 U6120_U2 ( .INP(WX5907), .ZN(U6120_n1) );
  NOR2X0 U6120_U1 ( .IN1(n9209), .IN2(U6120_n1), .QN(WX5970) );
  INVX0 U6121_U2 ( .INP(WX5905), .ZN(U6121_n1) );
  NOR2X0 U6121_U1 ( .IN1(n9209), .IN2(U6121_n1), .QN(WX5968) );
  INVX0 U6122_U2 ( .INP(test_so48), .ZN(U6122_n1) );
  NOR2X0 U6122_U1 ( .IN1(n9209), .IN2(U6122_n1), .QN(WX5966) );
  INVX0 U6123_U2 ( .INP(WX5901), .ZN(U6123_n1) );
  NOR2X0 U6123_U1 ( .IN1(n9208), .IN2(U6123_n1), .QN(WX5964) );
  INVX0 U6124_U2 ( .INP(WX5899), .ZN(U6124_n1) );
  NOR2X0 U6124_U1 ( .IN1(n9208), .IN2(U6124_n1), .QN(WX5962) );
  INVX0 U6125_U2 ( .INP(WX5897), .ZN(U6125_n1) );
  NOR2X0 U6125_U1 ( .IN1(n9208), .IN2(U6125_n1), .QN(WX5960) );
  INVX0 U6126_U2 ( .INP(WX5895), .ZN(U6126_n1) );
  NOR2X0 U6126_U1 ( .IN1(n9208), .IN2(U6126_n1), .QN(WX5958) );
  INVX0 U6127_U2 ( .INP(WX5893), .ZN(U6127_n1) );
  NOR2X0 U6127_U1 ( .IN1(n9208), .IN2(U6127_n1), .QN(WX5956) );
  INVX0 U6128_U2 ( .INP(WX5891), .ZN(U6128_n1) );
  NOR2X0 U6128_U1 ( .IN1(n9208), .IN2(U6128_n1), .QN(WX5954) );
  INVX0 U6129_U2 ( .INP(WX5889), .ZN(U6129_n1) );
  NOR2X0 U6129_U1 ( .IN1(n9219), .IN2(U6129_n1), .QN(WX5952) );
  INVX0 U6130_U2 ( .INP(WX5887), .ZN(U6130_n1) );
  NOR2X0 U6130_U1 ( .IN1(n9208), .IN2(U6130_n1), .QN(WX5950) );
  INVX0 U6131_U2 ( .INP(WX5885), .ZN(U6131_n1) );
  NOR2X0 U6131_U1 ( .IN1(n9208), .IN2(U6131_n1), .QN(WX5948) );
  INVX0 U6132_U2 ( .INP(WX5883), .ZN(U6132_n1) );
  NOR2X0 U6132_U1 ( .IN1(n9208), .IN2(U6132_n1), .QN(WX5946) );
  INVX0 U6133_U2 ( .INP(WX5881), .ZN(U6133_n1) );
  NOR2X0 U6133_U1 ( .IN1(n9208), .IN2(U6133_n1), .QN(WX5944) );
  INVX0 U6134_U2 ( .INP(WX5879), .ZN(U6134_n1) );
  NOR2X0 U6134_U1 ( .IN1(n9208), .IN2(U6134_n1), .QN(WX5942) );
  INVX0 U6135_U2 ( .INP(WX5877), .ZN(U6135_n1) );
  NOR2X0 U6135_U1 ( .IN1(n9208), .IN2(U6135_n1), .QN(WX5940) );
  INVX0 U6136_U2 ( .INP(WX5875), .ZN(U6136_n1) );
  NOR2X0 U6136_U1 ( .IN1(n9207), .IN2(U6136_n1), .QN(WX5938) );
  INVX0 U6137_U2 ( .INP(WX5873), .ZN(U6137_n1) );
  NOR2X0 U6137_U1 ( .IN1(n9207), .IN2(U6137_n1), .QN(WX5936) );
  INVX0 U6138_U2 ( .INP(WX5871), .ZN(U6138_n1) );
  NOR2X0 U6138_U1 ( .IN1(n9207), .IN2(U6138_n1), .QN(WX5934) );
  INVX0 U6139_U2 ( .INP(test_so47), .ZN(U6139_n1) );
  NOR2X0 U6139_U1 ( .IN1(n9207), .IN2(U6139_n1), .QN(WX5932) );
  INVX0 U6140_U2 ( .INP(WX5867), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n9207), .IN2(U6140_n1), .QN(WX5930) );
  INVX0 U6141_U2 ( .INP(WX5865), .ZN(U6141_n1) );
  NOR2X0 U6141_U1 ( .IN1(n9207), .IN2(U6141_n1), .QN(WX5928) );
  INVX0 U6142_U2 ( .INP(WX5863), .ZN(U6142_n1) );
  NOR2X0 U6142_U1 ( .IN1(n9207), .IN2(U6142_n1), .QN(WX5926) );
  INVX0 U6143_U2 ( .INP(WX5861), .ZN(U6143_n1) );
  NOR2X0 U6143_U1 ( .IN1(n9207), .IN2(U6143_n1), .QN(WX5924) );
  INVX0 U6144_U2 ( .INP(WX5859), .ZN(U6144_n1) );
  NOR2X0 U6144_U1 ( .IN1(n9207), .IN2(U6144_n1), .QN(WX5922) );
  INVX0 U6145_U2 ( .INP(WX5857), .ZN(U6145_n1) );
  NOR2X0 U6145_U1 ( .IN1(n9207), .IN2(U6145_n1), .QN(WX5920) );
  INVX0 U6146_U2 ( .INP(WX5855), .ZN(U6146_n1) );
  NOR2X0 U6146_U1 ( .IN1(n9207), .IN2(U6146_n1), .QN(WX5918) );
  INVX0 U6147_U2 ( .INP(WX5853), .ZN(U6147_n1) );
  NOR2X0 U6147_U1 ( .IN1(n9207), .IN2(U6147_n1), .QN(WX5916) );
  INVX0 U6148_U2 ( .INP(WX5851), .ZN(U6148_n1) );
  NOR2X0 U6148_U1 ( .IN1(n9206), .IN2(U6148_n1), .QN(WX5914) );
  INVX0 U6149_U2 ( .INP(WX5849), .ZN(U6149_n1) );
  NOR2X0 U6149_U1 ( .IN1(n9206), .IN2(U6149_n1), .QN(WX5912) );
  INVX0 U6150_U2 ( .INP(WX4714), .ZN(U6150_n1) );
  NOR2X0 U6150_U1 ( .IN1(n9206), .IN2(U6150_n1), .QN(WX4777) );
  INVX0 U6151_U2 ( .INP(WX4712), .ZN(U6151_n1) );
  NOR2X0 U6151_U1 ( .IN1(n9206), .IN2(U6151_n1), .QN(WX4775) );
  INVX0 U6152_U2 ( .INP(WX4710), .ZN(U6152_n1) );
  NOR2X0 U6152_U1 ( .IN1(n9206), .IN2(U6152_n1), .QN(WX4773) );
  INVX0 U6153_U2 ( .INP(WX4708), .ZN(U6153_n1) );
  NOR2X0 U6153_U1 ( .IN1(n9206), .IN2(U6153_n1), .QN(WX4771) );
  INVX0 U6154_U2 ( .INP(WX4706), .ZN(U6154_n1) );
  NOR2X0 U6154_U1 ( .IN1(n9206), .IN2(U6154_n1), .QN(WX4769) );
  INVX0 U6155_U2 ( .INP(WX4704), .ZN(U6155_n1) );
  NOR2X0 U6155_U1 ( .IN1(n9206), .IN2(U6155_n1), .QN(WX4767) );
  INVX0 U6156_U2 ( .INP(WX4702), .ZN(U6156_n1) );
  NOR2X0 U6156_U1 ( .IN1(n9206), .IN2(U6156_n1), .QN(WX4765) );
  INVX0 U6157_U2 ( .INP(WX4700), .ZN(U6157_n1) );
  NOR2X0 U6157_U1 ( .IN1(n9206), .IN2(U6157_n1), .QN(WX4763) );
  INVX0 U6158_U2 ( .INP(WX4698), .ZN(U6158_n1) );
  NOR2X0 U6158_U1 ( .IN1(n9206), .IN2(U6158_n1), .QN(WX4761) );
  INVX0 U6159_U2 ( .INP(WX4696), .ZN(U6159_n1) );
  NOR2X0 U6159_U1 ( .IN1(n9206), .IN2(U6159_n1), .QN(WX4759) );
  INVX0 U6160_U2 ( .INP(WX4694), .ZN(U6160_n1) );
  NOR2X0 U6160_U1 ( .IN1(n9206), .IN2(U6160_n1), .QN(WX4757) );
  INVX0 U6161_U2 ( .INP(WX4692), .ZN(U6161_n1) );
  NOR2X0 U6161_U1 ( .IN1(n9205), .IN2(U6161_n1), .QN(WX4755) );
  INVX0 U6162_U2 ( .INP(WX4690), .ZN(U6162_n1) );
  NOR2X0 U6162_U1 ( .IN1(n9205), .IN2(U6162_n1), .QN(WX4753) );
  INVX0 U6163_U2 ( .INP(test_so39), .ZN(U6163_n1) );
  NOR2X0 U6163_U1 ( .IN1(n9205), .IN2(U6163_n1), .QN(WX4751) );
  INVX0 U6164_U2 ( .INP(WX4686), .ZN(U6164_n1) );
  NOR2X0 U6164_U1 ( .IN1(n9205), .IN2(U6164_n1), .QN(WX4749) );
  INVX0 U6165_U2 ( .INP(WX4684), .ZN(U6165_n1) );
  NOR2X0 U6165_U1 ( .IN1(n9205), .IN2(U6165_n1), .QN(WX4747) );
  INVX0 U6166_U2 ( .INP(WX4682), .ZN(U6166_n1) );
  NOR2X0 U6166_U1 ( .IN1(n9205), .IN2(U6166_n1), .QN(WX4745) );
  INVX0 U6167_U2 ( .INP(WX4680), .ZN(U6167_n1) );
  NOR2X0 U6167_U1 ( .IN1(n9205), .IN2(U6167_n1), .QN(WX4743) );
  INVX0 U6168_U2 ( .INP(WX4678), .ZN(U6168_n1) );
  NOR2X0 U6168_U1 ( .IN1(n9205), .IN2(U6168_n1), .QN(WX4741) );
  INVX0 U6169_U2 ( .INP(WX4676), .ZN(U6169_n1) );
  NOR2X0 U6169_U1 ( .IN1(n9205), .IN2(U6169_n1), .QN(WX4739) );
  INVX0 U6170_U2 ( .INP(WX4674), .ZN(U6170_n1) );
  NOR2X0 U6170_U1 ( .IN1(n9205), .IN2(U6170_n1), .QN(WX4737) );
  INVX0 U6171_U2 ( .INP(WX4672), .ZN(U6171_n1) );
  NOR2X0 U6171_U1 ( .IN1(n9205), .IN2(U6171_n1), .QN(WX4735) );
  INVX0 U6172_U2 ( .INP(WX4670), .ZN(U6172_n1) );
  NOR2X0 U6172_U1 ( .IN1(n9205), .IN2(U6172_n1), .QN(WX4733) );
  INVX0 U6173_U2 ( .INP(WX4668), .ZN(U6173_n1) );
  NOR2X0 U6173_U1 ( .IN1(n9205), .IN2(U6173_n1), .QN(WX4731) );
  INVX0 U6174_U2 ( .INP(WX4666), .ZN(U6174_n1) );
  NOR2X0 U6174_U1 ( .IN1(n9204), .IN2(U6174_n1), .QN(WX4729) );
  INVX0 U6175_U2 ( .INP(WX4664), .ZN(U6175_n1) );
  NOR2X0 U6175_U1 ( .IN1(n9204), .IN2(U6175_n1), .QN(WX4727) );
  INVX0 U6176_U2 ( .INP(WX4662), .ZN(U6176_n1) );
  NOR2X0 U6176_U1 ( .IN1(n9204), .IN2(U6176_n1), .QN(WX4725) );
  INVX0 U6177_U2 ( .INP(WX4660), .ZN(U6177_n1) );
  NOR2X0 U6177_U1 ( .IN1(n9204), .IN2(U6177_n1), .QN(WX4723) );
  INVX0 U6178_U2 ( .INP(WX4658), .ZN(U6178_n1) );
  NOR2X0 U6178_U1 ( .IN1(n9204), .IN2(U6178_n1), .QN(WX4721) );
  INVX0 U6179_U2 ( .INP(WX4656), .ZN(U6179_n1) );
  NOR2X0 U6179_U1 ( .IN1(n9204), .IN2(U6179_n1), .QN(WX4719) );
  INVX0 U6180_U2 ( .INP(test_so38), .ZN(U6180_n1) );
  NOR2X0 U6180_U1 ( .IN1(n9204), .IN2(U6180_n1), .QN(WX4717) );
  INVX0 U6181_U2 ( .INP(WX4652), .ZN(U6181_n1) );
  NOR2X0 U6181_U1 ( .IN1(n9204), .IN2(U6181_n1), .QN(WX4715) );
  INVX0 U6182_U2 ( .INP(WX4650), .ZN(U6182_n1) );
  NOR2X0 U6182_U1 ( .IN1(n9204), .IN2(U6182_n1), .QN(WX4713) );
  INVX0 U6183_U2 ( .INP(WX4648), .ZN(U6183_n1) );
  NOR2X0 U6183_U1 ( .IN1(n9204), .IN2(U6183_n1), .QN(WX4711) );
  INVX0 U6184_U2 ( .INP(WX4646), .ZN(U6184_n1) );
  NOR2X0 U6184_U1 ( .IN1(n9204), .IN2(U6184_n1), .QN(WX4709) );
  INVX0 U6185_U2 ( .INP(WX4644), .ZN(U6185_n1) );
  NOR2X0 U6185_U1 ( .IN1(n9204), .IN2(U6185_n1), .QN(WX4707) );
  INVX0 U6186_U2 ( .INP(WX4642), .ZN(U6186_n1) );
  NOR2X0 U6186_U1 ( .IN1(n9204), .IN2(U6186_n1), .QN(WX4705) );
  INVX0 U6187_U2 ( .INP(WX4640), .ZN(U6187_n1) );
  NOR2X0 U6187_U1 ( .IN1(n9203), .IN2(U6187_n1), .QN(WX4703) );
  INVX0 U6188_U2 ( .INP(WX4638), .ZN(U6188_n1) );
  NOR2X0 U6188_U1 ( .IN1(n9203), .IN2(U6188_n1), .QN(WX4701) );
  INVX0 U6189_U2 ( .INP(WX4636), .ZN(U6189_n1) );
  NOR2X0 U6189_U1 ( .IN1(n9207), .IN2(U6189_n1), .QN(WX4699) );
  INVX0 U6190_U2 ( .INP(WX4634), .ZN(U6190_n1) );
  NOR2X0 U6190_U1 ( .IN1(n9219), .IN2(U6190_n1), .QN(WX4697) );
  INVX0 U6191_U2 ( .INP(WX4632), .ZN(U6191_n1) );
  NOR2X0 U6191_U1 ( .IN1(n9219), .IN2(U6191_n1), .QN(WX4695) );
  INVX0 U6192_U2 ( .INP(WX4630), .ZN(U6192_n1) );
  NOR2X0 U6192_U1 ( .IN1(n9218), .IN2(U6192_n1), .QN(WX4693) );
  INVX0 U6193_U2 ( .INP(WX4628), .ZN(U6193_n1) );
  NOR2X0 U6193_U1 ( .IN1(n9218), .IN2(U6193_n1), .QN(WX4691) );
  INVX0 U6194_U2 ( .INP(WX4626), .ZN(U6194_n1) );
  NOR2X0 U6194_U1 ( .IN1(n9218), .IN2(U6194_n1), .QN(WX4689) );
  INVX0 U6195_U2 ( .INP(WX4624), .ZN(U6195_n1) );
  NOR2X0 U6195_U1 ( .IN1(n9218), .IN2(U6195_n1), .QN(WX4687) );
  INVX0 U6196_U2 ( .INP(WX4622), .ZN(U6196_n1) );
  NOR2X0 U6196_U1 ( .IN1(n9218), .IN2(U6196_n1), .QN(WX4685) );
  INVX0 U6197_U2 ( .INP(test_so37), .ZN(U6197_n1) );
  NOR2X0 U6197_U1 ( .IN1(n9218), .IN2(U6197_n1), .QN(WX4683) );
  INVX0 U6198_U2 ( .INP(WX4618), .ZN(U6198_n1) );
  NOR2X0 U6198_U1 ( .IN1(n9218), .IN2(U6198_n1), .QN(WX4681) );
  INVX0 U6199_U2 ( .INP(WX4616), .ZN(U6199_n1) );
  NOR2X0 U6199_U1 ( .IN1(n9218), .IN2(U6199_n1), .QN(WX4679) );
  INVX0 U6200_U2 ( .INP(WX4614), .ZN(U6200_n1) );
  NOR2X0 U6200_U1 ( .IN1(n9218), .IN2(U6200_n1), .QN(WX4677) );
  INVX0 U6201_U2 ( .INP(WX4612), .ZN(U6201_n1) );
  NOR2X0 U6201_U1 ( .IN1(n9218), .IN2(U6201_n1), .QN(WX4675) );
  INVX0 U6202_U2 ( .INP(WX4610), .ZN(U6202_n1) );
  NOR2X0 U6202_U1 ( .IN1(n9218), .IN2(U6202_n1), .QN(WX4673) );
  INVX0 U6203_U2 ( .INP(WX4608), .ZN(U6203_n1) );
  NOR2X0 U6203_U1 ( .IN1(n9218), .IN2(U6203_n1), .QN(WX4671) );
  INVX0 U6204_U2 ( .INP(WX4606), .ZN(U6204_n1) );
  NOR2X0 U6204_U1 ( .IN1(n9218), .IN2(U6204_n1), .QN(WX4669) );
  INVX0 U6205_U2 ( .INP(WX4604), .ZN(U6205_n1) );
  NOR2X0 U6205_U1 ( .IN1(n9217), .IN2(U6205_n1), .QN(WX4667) );
  INVX0 U6206_U2 ( .INP(WX4602), .ZN(U6206_n1) );
  NOR2X0 U6206_U1 ( .IN1(n9217), .IN2(U6206_n1), .QN(WX4665) );
  INVX0 U6207_U2 ( .INP(WX4600), .ZN(U6207_n1) );
  NOR2X0 U6207_U1 ( .IN1(n9217), .IN2(U6207_n1), .QN(WX4663) );
  INVX0 U6208_U2 ( .INP(WX4598), .ZN(U6208_n1) );
  NOR2X0 U6208_U1 ( .IN1(n9217), .IN2(U6208_n1), .QN(WX4661) );
  INVX0 U6209_U2 ( .INP(WX4596), .ZN(U6209_n1) );
  NOR2X0 U6209_U1 ( .IN1(n9217), .IN2(U6209_n1), .QN(WX4659) );
  INVX0 U6210_U2 ( .INP(WX4594), .ZN(U6210_n1) );
  NOR2X0 U6210_U1 ( .IN1(n9217), .IN2(U6210_n1), .QN(WX4657) );
  INVX0 U6211_U2 ( .INP(WX4592), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n9217), .IN2(U6211_n1), .QN(WX4655) );
  INVX0 U6212_U2 ( .INP(WX4590), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n9217), .IN2(U6212_n1), .QN(WX4653) );
  INVX0 U6213_U2 ( .INP(WX4588), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n9217), .IN2(U6213_n1), .QN(WX4651) );
  INVX0 U6214_U2 ( .INP(test_so36), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n9217), .IN2(U6214_n1), .QN(WX4649) );
  INVX0 U6215_U2 ( .INP(WX4584), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n9217), .IN2(U6215_n1), .QN(WX4647) );
  INVX0 U6216_U2 ( .INP(WX4582), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n9217), .IN2(U6216_n1), .QN(WX4645) );
  INVX0 U6217_U2 ( .INP(WX4580), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n9217), .IN2(U6217_n1), .QN(WX4643) );
  INVX0 U6218_U2 ( .INP(WX4578), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n9216), .IN2(U6218_n1), .QN(WX4641) );
  INVX0 U6219_U2 ( .INP(WX4576), .ZN(U6219_n1) );
  NOR2X0 U6219_U1 ( .IN1(n9216), .IN2(U6219_n1), .QN(WX4639) );
  INVX0 U6220_U2 ( .INP(WX4574), .ZN(U6220_n1) );
  NOR2X0 U6220_U1 ( .IN1(n9216), .IN2(U6220_n1), .QN(WX4637) );
  INVX0 U6221_U2 ( .INP(WX4572), .ZN(U6221_n1) );
  NOR2X0 U6221_U1 ( .IN1(n9216), .IN2(U6221_n1), .QN(WX4635) );
  INVX0 U6222_U2 ( .INP(WX4570), .ZN(U6222_n1) );
  NOR2X0 U6222_U1 ( .IN1(n9216), .IN2(U6222_n1), .QN(WX4633) );
  INVX0 U6223_U2 ( .INP(WX4568), .ZN(U6223_n1) );
  NOR2X0 U6223_U1 ( .IN1(n9216), .IN2(U6223_n1), .QN(WX4631) );
  INVX0 U6224_U2 ( .INP(WX4566), .ZN(U6224_n1) );
  NOR2X0 U6224_U1 ( .IN1(n9216), .IN2(U6224_n1), .QN(WX4629) );
  INVX0 U6225_U2 ( .INP(WX4564), .ZN(U6225_n1) );
  NOR2X0 U6225_U1 ( .IN1(n9216), .IN2(U6225_n1), .QN(WX4627) );
  INVX0 U6226_U2 ( .INP(WX4562), .ZN(U6226_n1) );
  NOR2X0 U6226_U1 ( .IN1(n9216), .IN2(U6226_n1), .QN(WX4625) );
  INVX0 U6227_U2 ( .INP(WX4560), .ZN(U6227_n1) );
  NOR2X0 U6227_U1 ( .IN1(n9216), .IN2(U6227_n1), .QN(WX4623) );
  INVX0 U6228_U2 ( .INP(WX4558), .ZN(U6228_n1) );
  NOR2X0 U6228_U1 ( .IN1(n9216), .IN2(U6228_n1), .QN(WX4621) );
  INVX0 U6229_U2 ( .INP(WX4556), .ZN(U6229_n1) );
  NOR2X0 U6229_U1 ( .IN1(n9216), .IN2(U6229_n1), .QN(WX4619) );
  INVX0 U6230_U2 ( .INP(WX3421), .ZN(U6230_n1) );
  NOR2X0 U6230_U1 ( .IN1(n9216), .IN2(U6230_n1), .QN(WX3484) );
  INVX0 U6231_U2 ( .INP(WX3419), .ZN(U6231_n1) );
  NOR2X0 U6231_U1 ( .IN1(n9215), .IN2(U6231_n1), .QN(WX3482) );
  INVX0 U6232_U2 ( .INP(WX3417), .ZN(U6232_n1) );
  NOR2X0 U6232_U1 ( .IN1(n9215), .IN2(U6232_n1), .QN(WX3480) );
  INVX0 U6233_U2 ( .INP(WX3415), .ZN(U6233_n1) );
  NOR2X0 U6233_U1 ( .IN1(n9215), .IN2(U6233_n1), .QN(WX3478) );
  INVX0 U6234_U2 ( .INP(WX3413), .ZN(U6234_n1) );
  NOR2X0 U6234_U1 ( .IN1(n9215), .IN2(U6234_n1), .QN(WX3476) );
  INVX0 U6235_U2 ( .INP(WX3411), .ZN(U6235_n1) );
  NOR2X0 U6235_U1 ( .IN1(n9215), .IN2(U6235_n1), .QN(WX3474) );
  INVX0 U6236_U2 ( .INP(WX3409), .ZN(U6236_n1) );
  NOR2X0 U6236_U1 ( .IN1(n9215), .IN2(U6236_n1), .QN(WX3472) );
  INVX0 U6237_U2 ( .INP(WX3407), .ZN(U6237_n1) );
  NOR2X0 U6237_U1 ( .IN1(n9215), .IN2(U6237_n1), .QN(WX3470) );
  INVX0 U6238_U2 ( .INP(test_so28), .ZN(U6238_n1) );
  NOR2X0 U6238_U1 ( .IN1(n9215), .IN2(U6238_n1), .QN(WX3468) );
  INVX0 U6239_U2 ( .INP(WX3403), .ZN(U6239_n1) );
  NOR2X0 U6239_U1 ( .IN1(n9215), .IN2(U6239_n1), .QN(WX3466) );
  INVX0 U6240_U2 ( .INP(WX3401), .ZN(U6240_n1) );
  NOR2X0 U6240_U1 ( .IN1(n9215), .IN2(U6240_n1), .QN(WX3464) );
  INVX0 U6241_U2 ( .INP(WX3399), .ZN(U6241_n1) );
  NOR2X0 U6241_U1 ( .IN1(n9215), .IN2(U6241_n1), .QN(WX3462) );
  INVX0 U6242_U2 ( .INP(WX3397), .ZN(U6242_n1) );
  NOR2X0 U6242_U1 ( .IN1(n9215), .IN2(U6242_n1), .QN(WX3460) );
  INVX0 U6243_U2 ( .INP(WX3395), .ZN(U6243_n1) );
  NOR2X0 U6243_U1 ( .IN1(n9214), .IN2(U6243_n1), .QN(WX3458) );
  INVX0 U6244_U2 ( .INP(WX3393), .ZN(U6244_n1) );
  NOR2X0 U6244_U1 ( .IN1(n9214), .IN2(U6244_n1), .QN(WX3456) );
  INVX0 U6245_U2 ( .INP(WX3391), .ZN(U6245_n1) );
  NOR2X0 U6245_U1 ( .IN1(n9214), .IN2(U6245_n1), .QN(WX3454) );
  INVX0 U6246_U2 ( .INP(WX3389), .ZN(U6246_n1) );
  NOR2X0 U6246_U1 ( .IN1(n9214), .IN2(U6246_n1), .QN(WX3452) );
  INVX0 U6247_U2 ( .INP(WX3387), .ZN(U6247_n1) );
  NOR2X0 U6247_U1 ( .IN1(n9214), .IN2(U6247_n1), .QN(WX3450) );
  INVX0 U6248_U2 ( .INP(WX3385), .ZN(U6248_n1) );
  NOR2X0 U6248_U1 ( .IN1(n9214), .IN2(U6248_n1), .QN(WX3448) );
  INVX0 U6249_U2 ( .INP(WX3383), .ZN(U6249_n1) );
  NOR2X0 U6249_U1 ( .IN1(n9214), .IN2(U6249_n1), .QN(WX3446) );
  INVX0 U6250_U2 ( .INP(WX3381), .ZN(U6250_n1) );
  NOR2X0 U6250_U1 ( .IN1(n9214), .IN2(U6250_n1), .QN(WX3444) );
  INVX0 U6251_U2 ( .INP(WX3379), .ZN(U6251_n1) );
  NOR2X0 U6251_U1 ( .IN1(n9214), .IN2(U6251_n1), .QN(WX3442) );
  INVX0 U6252_U2 ( .INP(WX3377), .ZN(U6252_n1) );
  NOR2X0 U6252_U1 ( .IN1(n9214), .IN2(U6252_n1), .QN(WX3440) );
  INVX0 U6253_U2 ( .INP(WX3375), .ZN(U6253_n1) );
  NOR2X0 U6253_U1 ( .IN1(n9214), .IN2(U6253_n1), .QN(WX3438) );
  INVX0 U6254_U2 ( .INP(WX3373), .ZN(U6254_n1) );
  NOR2X0 U6254_U1 ( .IN1(n9214), .IN2(U6254_n1), .QN(WX3436) );
  INVX0 U6255_U2 ( .INP(WX3371), .ZN(U6255_n1) );
  NOR2X0 U6255_U1 ( .IN1(n9214), .IN2(U6255_n1), .QN(WX3434) );
  INVX0 U6256_U2 ( .INP(test_so27), .ZN(U6256_n1) );
  NOR2X0 U6256_U1 ( .IN1(n9213), .IN2(U6256_n1), .QN(WX3432) );
  INVX0 U6257_U2 ( .INP(WX3367), .ZN(U6257_n1) );
  NOR2X0 U6257_U1 ( .IN1(n9213), .IN2(U6257_n1), .QN(WX3430) );
  INVX0 U6258_U2 ( .INP(WX3365), .ZN(U6258_n1) );
  NOR2X0 U6258_U1 ( .IN1(n9213), .IN2(U6258_n1), .QN(WX3428) );
  INVX0 U6259_U2 ( .INP(WX3363), .ZN(U6259_n1) );
  NOR2X0 U6259_U1 ( .IN1(n9213), .IN2(U6259_n1), .QN(WX3426) );
  INVX0 U6260_U2 ( .INP(WX3361), .ZN(U6260_n1) );
  NOR2X0 U6260_U1 ( .IN1(n9213), .IN2(U6260_n1), .QN(WX3424) );
  INVX0 U6261_U2 ( .INP(WX3359), .ZN(U6261_n1) );
  NOR2X0 U6261_U1 ( .IN1(n9213), .IN2(U6261_n1), .QN(WX3422) );
  INVX0 U6262_U2 ( .INP(WX3357), .ZN(U6262_n1) );
  NOR2X0 U6262_U1 ( .IN1(n9213), .IN2(U6262_n1), .QN(WX3420) );
  INVX0 U6263_U2 ( .INP(WX3355), .ZN(U6263_n1) );
  NOR2X0 U6263_U1 ( .IN1(n9213), .IN2(U6263_n1), .QN(WX3418) );
  INVX0 U6264_U2 ( .INP(WX3353), .ZN(U6264_n1) );
  NOR2X0 U6264_U1 ( .IN1(n9213), .IN2(U6264_n1), .QN(WX3416) );
  INVX0 U6265_U2 ( .INP(WX3351), .ZN(U6265_n1) );
  NOR2X0 U6265_U1 ( .IN1(n9213), .IN2(U6265_n1), .QN(WX3414) );
  INVX0 U6266_U2 ( .INP(WX3349), .ZN(U6266_n1) );
  NOR2X0 U6266_U1 ( .IN1(n9213), .IN2(U6266_n1), .QN(WX3412) );
  INVX0 U6267_U2 ( .INP(WX3347), .ZN(U6267_n1) );
  NOR2X0 U6267_U1 ( .IN1(n9213), .IN2(U6267_n1), .QN(WX3410) );
  INVX0 U6268_U2 ( .INP(WX3345), .ZN(U6268_n1) );
  NOR2X0 U6268_U1 ( .IN1(n9213), .IN2(U6268_n1), .QN(WX3408) );
  INVX0 U6269_U2 ( .INP(WX3343), .ZN(U6269_n1) );
  NOR2X0 U6269_U1 ( .IN1(n9212), .IN2(U6269_n1), .QN(WX3406) );
  INVX0 U6270_U2 ( .INP(WX3341), .ZN(U6270_n1) );
  NOR2X0 U6270_U1 ( .IN1(n9212), .IN2(U6270_n1), .QN(WX3404) );
  INVX0 U6271_U2 ( .INP(WX3339), .ZN(U6271_n1) );
  NOR2X0 U6271_U1 ( .IN1(n9212), .IN2(U6271_n1), .QN(WX3402) );
  INVX0 U6272_U2 ( .INP(WX3337), .ZN(U6272_n1) );
  NOR2X0 U6272_U1 ( .IN1(n9212), .IN2(U6272_n1), .QN(WX3400) );
  INVX0 U6273_U2 ( .INP(WX3335), .ZN(U6273_n1) );
  NOR2X0 U6273_U1 ( .IN1(n9212), .IN2(U6273_n1), .QN(WX3398) );
  INVX0 U6274_U2 ( .INP(test_so26), .ZN(U6274_n1) );
  NOR2X0 U6274_U1 ( .IN1(n9212), .IN2(U6274_n1), .QN(WX3396) );
  INVX0 U6275_U2 ( .INP(WX3331), .ZN(U6275_n1) );
  NOR2X0 U6275_U1 ( .IN1(n9212), .IN2(U6275_n1), .QN(WX3394) );
  INVX0 U6276_U2 ( .INP(WX3329), .ZN(U6276_n1) );
  NOR2X0 U6276_U1 ( .IN1(n9212), .IN2(U6276_n1), .QN(WX3392) );
  INVX0 U6277_U2 ( .INP(WX3327), .ZN(U6277_n1) );
  NOR2X0 U6277_U1 ( .IN1(n9212), .IN2(U6277_n1), .QN(WX3390) );
  INVX0 U6278_U2 ( .INP(WX3325), .ZN(U6278_n1) );
  NOR2X0 U6278_U1 ( .IN1(n9212), .IN2(U6278_n1), .QN(WX3388) );
  INVX0 U6279_U2 ( .INP(WX3323), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n9212), .IN2(U6279_n1), .QN(WX3386) );
  INVX0 U6280_U2 ( .INP(WX3321), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n9212), .IN2(U6280_n1), .QN(WX3384) );
  INVX0 U6281_U2 ( .INP(WX3319), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n9212), .IN2(U6281_n1), .QN(WX3382) );
  INVX0 U6282_U2 ( .INP(WX3317), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n9211), .IN2(U6282_n1), .QN(WX3380) );
  INVX0 U6283_U2 ( .INP(WX3315), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n9211), .IN2(U6283_n1), .QN(WX3378) );
  INVX0 U6284_U2 ( .INP(WX3313), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n9211), .IN2(U6284_n1), .QN(WX3376) );
  INVX0 U6285_U2 ( .INP(WX3311), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n9211), .IN2(U6285_n1), .QN(WX3374) );
  INVX0 U6286_U2 ( .INP(WX3309), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n9211), .IN2(U6286_n1), .QN(WX3372) );
  INVX0 U6287_U2 ( .INP(WX3307), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n9211), .IN2(U6287_n1), .QN(WX3370) );
  INVX0 U6288_U2 ( .INP(WX3305), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n9215), .IN2(U6288_n1), .QN(WX3368) );
  INVX0 U6289_U2 ( .INP(WX3303), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n9208), .IN2(U6289_n1), .QN(WX3366) );
  INVX0 U6290_U2 ( .INP(WX3301), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n9164), .IN2(U6290_n1), .QN(WX3364) );
  INVX0 U6291_U2 ( .INP(WX3299), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n9171), .IN2(U6291_n1), .QN(WX3362) );
  INVX0 U6292_U2 ( .INP(test_so25), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n9171), .IN2(U6292_n1), .QN(WX3360) );
  INVX0 U6293_U2 ( .INP(WX3295), .ZN(U6293_n1) );
  NOR2X0 U6293_U1 ( .IN1(n9171), .IN2(U6293_n1), .QN(WX3358) );
  INVX0 U6294_U2 ( .INP(WX3293), .ZN(U6294_n1) );
  NOR2X0 U6294_U1 ( .IN1(n9171), .IN2(U6294_n1), .QN(WX3356) );
  INVX0 U6295_U2 ( .INP(WX3291), .ZN(U6295_n1) );
  NOR2X0 U6295_U1 ( .IN1(n9171), .IN2(U6295_n1), .QN(WX3354) );
  INVX0 U6296_U2 ( .INP(WX3289), .ZN(U6296_n1) );
  NOR2X0 U6296_U1 ( .IN1(n9171), .IN2(U6296_n1), .QN(WX3352) );
  INVX0 U6297_U2 ( .INP(WX3287), .ZN(U6297_n1) );
  NOR2X0 U6297_U1 ( .IN1(n9171), .IN2(U6297_n1), .QN(WX3350) );
  INVX0 U6298_U2 ( .INP(WX3285), .ZN(U6298_n1) );
  NOR2X0 U6298_U1 ( .IN1(n9171), .IN2(U6298_n1), .QN(WX3348) );
  INVX0 U6299_U2 ( .INP(WX3283), .ZN(U6299_n1) );
  NOR2X0 U6299_U1 ( .IN1(n9171), .IN2(U6299_n1), .QN(WX3346) );
  INVX0 U6300_U2 ( .INP(WX3281), .ZN(U6300_n1) );
  NOR2X0 U6300_U1 ( .IN1(n9171), .IN2(U6300_n1), .QN(WX3344) );
  INVX0 U6301_U2 ( .INP(WX3279), .ZN(U6301_n1) );
  NOR2X0 U6301_U1 ( .IN1(n9170), .IN2(U6301_n1), .QN(WX3342) );
  INVX0 U6302_U2 ( .INP(WX3277), .ZN(U6302_n1) );
  NOR2X0 U6302_U1 ( .IN1(n9170), .IN2(U6302_n1), .QN(WX3340) );
  INVX0 U6303_U2 ( .INP(WX3275), .ZN(U6303_n1) );
  NOR2X0 U6303_U1 ( .IN1(n9170), .IN2(U6303_n1), .QN(WX3338) );
  INVX0 U6304_U2 ( .INP(WX3273), .ZN(U6304_n1) );
  NOR2X0 U6304_U1 ( .IN1(n9170), .IN2(U6304_n1), .QN(WX3336) );
  INVX0 U6305_U2 ( .INP(WX3271), .ZN(U6305_n1) );
  NOR2X0 U6305_U1 ( .IN1(n9170), .IN2(U6305_n1), .QN(WX3334) );
  INVX0 U6306_U2 ( .INP(WX3267), .ZN(U6306_n1) );
  NOR2X0 U6306_U1 ( .IN1(n9170), .IN2(U6306_n1), .QN(WX3330) );
  INVX0 U6307_U2 ( .INP(WX2128), .ZN(U6307_n1) );
  NOR2X0 U6307_U1 ( .IN1(n9170), .IN2(U6307_n1), .QN(WX2191) );
  INVX0 U6308_U2 ( .INP(WX2126), .ZN(U6308_n1) );
  NOR2X0 U6308_U1 ( .IN1(n9170), .IN2(U6308_n1), .QN(WX2189) );
  INVX0 U6309_U2 ( .INP(WX2124), .ZN(U6309_n1) );
  NOR2X0 U6309_U1 ( .IN1(n9170), .IN2(U6309_n1), .QN(WX2187) );
  INVX0 U6310_U2 ( .INP(WX2122), .ZN(U6310_n1) );
  NOR2X0 U6310_U1 ( .IN1(n9170), .IN2(U6310_n1), .QN(WX2185) );
  INVX0 U6311_U2 ( .INP(WX2120), .ZN(U6311_n1) );
  NOR2X0 U6311_U1 ( .IN1(n9170), .IN2(U6311_n1), .QN(WX2183) );
  INVX0 U6312_U2 ( .INP(WX2118), .ZN(U6312_n1) );
  NOR2X0 U6312_U1 ( .IN1(n9170), .IN2(U6312_n1), .QN(WX2181) );
  INVX0 U6313_U2 ( .INP(WX2116), .ZN(U6313_n1) );
  NOR2X0 U6313_U1 ( .IN1(n9170), .IN2(U6313_n1), .QN(WX2179) );
  INVX0 U6314_U2 ( .INP(WX2114), .ZN(U6314_n1) );
  NOR2X0 U6314_U1 ( .IN1(n9169), .IN2(U6314_n1), .QN(WX2177) );
  INVX0 U6315_U2 ( .INP(WX2112), .ZN(U6315_n1) );
  NOR2X0 U6315_U1 ( .IN1(n9169), .IN2(U6315_n1), .QN(WX2175) );
  INVX0 U6316_U2 ( .INP(WX2110), .ZN(U6316_n1) );
  NOR2X0 U6316_U1 ( .IN1(n9169), .IN2(U6316_n1), .QN(WX2173) );
  INVX0 U6317_U2 ( .INP(WX2108), .ZN(U6317_n1) );
  NOR2X0 U6317_U1 ( .IN1(n9169), .IN2(U6317_n1), .QN(WX2171) );
  INVX0 U6318_U2 ( .INP(WX2106), .ZN(U6318_n1) );
  NOR2X0 U6318_U1 ( .IN1(n9169), .IN2(U6318_n1), .QN(WX2169) );
  INVX0 U6319_U2 ( .INP(WX2104), .ZN(U6319_n1) );
  NOR2X0 U6319_U1 ( .IN1(n9169), .IN2(U6319_n1), .QN(WX2167) );
  INVX0 U6320_U2 ( .INP(WX2102), .ZN(U6320_n1) );
  NOR2X0 U6320_U1 ( .IN1(n9169), .IN2(U6320_n1), .QN(WX2165) );
  INVX0 U6321_U2 ( .INP(test_so17), .ZN(U6321_n1) );
  NOR2X0 U6321_U1 ( .IN1(n9169), .IN2(U6321_n1), .QN(WX2163) );
  INVX0 U6322_U2 ( .INP(WX2098), .ZN(U6322_n1) );
  NOR2X0 U6322_U1 ( .IN1(n9169), .IN2(U6322_n1), .QN(WX2161) );
  INVX0 U6323_U2 ( .INP(WX2096), .ZN(U6323_n1) );
  NOR2X0 U6323_U1 ( .IN1(n9169), .IN2(U6323_n1), .QN(WX2159) );
  INVX0 U6324_U2 ( .INP(WX2094), .ZN(U6324_n1) );
  NOR2X0 U6324_U1 ( .IN1(n9169), .IN2(U6324_n1), .QN(WX2157) );
  INVX0 U6325_U2 ( .INP(WX2092), .ZN(U6325_n1) );
  NOR2X0 U6325_U1 ( .IN1(n9169), .IN2(U6325_n1), .QN(WX2155) );
  INVX0 U6326_U2 ( .INP(WX2090), .ZN(U6326_n1) );
  NOR2X0 U6326_U1 ( .IN1(n9169), .IN2(U6326_n1), .QN(WX2153) );
  INVX0 U6327_U2 ( .INP(WX2088), .ZN(U6327_n1) );
  NOR2X0 U6327_U1 ( .IN1(n9168), .IN2(U6327_n1), .QN(WX2151) );
  INVX0 U6328_U2 ( .INP(WX2086), .ZN(U6328_n1) );
  NOR2X0 U6328_U1 ( .IN1(n9168), .IN2(U6328_n1), .QN(WX2149) );
  INVX0 U6329_U2 ( .INP(WX2084), .ZN(U6329_n1) );
  NOR2X0 U6329_U1 ( .IN1(n9168), .IN2(U6329_n1), .QN(WX2147) );
  INVX0 U6330_U2 ( .INP(WX2082), .ZN(U6330_n1) );
  NOR2X0 U6330_U1 ( .IN1(n9168), .IN2(U6330_n1), .QN(WX2145) );
  INVX0 U6331_U2 ( .INP(WX2080), .ZN(U6331_n1) );
  NOR2X0 U6331_U1 ( .IN1(n9168), .IN2(U6331_n1), .QN(WX2143) );
  INVX0 U6332_U2 ( .INP(WX2078), .ZN(U6332_n1) );
  NOR2X0 U6332_U1 ( .IN1(n9168), .IN2(U6332_n1), .QN(WX2141) );
  INVX0 U6333_U2 ( .INP(WX2076), .ZN(U6333_n1) );
  NOR2X0 U6333_U1 ( .IN1(n9168), .IN2(U6333_n1), .QN(WX2139) );
  INVX0 U6334_U2 ( .INP(WX2074), .ZN(U6334_n1) );
  NOR2X0 U6334_U1 ( .IN1(n9168), .IN2(U6334_n1), .QN(WX2137) );
  INVX0 U6335_U2 ( .INP(WX2072), .ZN(U6335_n1) );
  NOR2X0 U6335_U1 ( .IN1(n9168), .IN2(U6335_n1), .QN(WX2135) );
  INVX0 U6336_U2 ( .INP(WX2070), .ZN(U6336_n1) );
  NOR2X0 U6336_U1 ( .IN1(n9168), .IN2(U6336_n1), .QN(WX2133) );
  INVX0 U6337_U2 ( .INP(WX2068), .ZN(U6337_n1) );
  NOR2X0 U6337_U1 ( .IN1(n9168), .IN2(U6337_n1), .QN(WX2131) );
  INVX0 U6338_U2 ( .INP(WX2066), .ZN(U6338_n1) );
  NOR2X0 U6338_U1 ( .IN1(n9168), .IN2(U6338_n1), .QN(WX2129) );
  INVX0 U6339_U2 ( .INP(test_so16), .ZN(U6339_n1) );
  NOR2X0 U6339_U1 ( .IN1(n9167), .IN2(U6339_n1), .QN(WX2127) );
  INVX0 U6340_U2 ( .INP(WX2062), .ZN(U6340_n1) );
  NOR2X0 U6340_U1 ( .IN1(n9167), .IN2(U6340_n1), .QN(WX2125) );
  INVX0 U6341_U2 ( .INP(WX2060), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n9167), .IN2(U6341_n1), .QN(WX2123) );
  INVX0 U6342_U2 ( .INP(WX2058), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n9167), .IN2(U6342_n1), .QN(WX2121) );
  INVX0 U6343_U2 ( .INP(WX2056), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n9167), .IN2(U6343_n1), .QN(WX2119) );
  INVX0 U6344_U2 ( .INP(WX2054), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n9167), .IN2(U6344_n1), .QN(WX2117) );
  INVX0 U6345_U2 ( .INP(WX2052), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n9167), .IN2(U6345_n1), .QN(WX2115) );
  INVX0 U6346_U2 ( .INP(WX2050), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n9167), .IN2(U6346_n1), .QN(WX2113) );
  INVX0 U6347_U2 ( .INP(WX2048), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n9167), .IN2(U6347_n1), .QN(WX2111) );
  INVX0 U6348_U2 ( .INP(WX2046), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n9167), .IN2(U6348_n1), .QN(WX2109) );
  INVX0 U6349_U2 ( .INP(WX2044), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n9167), .IN2(U6349_n1), .QN(WX2107) );
  INVX0 U6350_U2 ( .INP(WX2042), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n9167), .IN2(U6350_n1), .QN(WX2105) );
  INVX0 U6351_U2 ( .INP(WX2040), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n9167), .IN2(U6351_n1), .QN(WX2103) );
  INVX0 U6352_U2 ( .INP(WX2038), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n9166), .IN2(U6352_n1), .QN(WX2101) );
  INVX0 U6353_U2 ( .INP(WX2036), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n9166), .IN2(U6353_n1), .QN(WX2099) );
  INVX0 U6354_U2 ( .INP(WX2034), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n9166), .IN2(U6354_n1), .QN(WX2097) );
  INVX0 U6355_U2 ( .INP(WX2032), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n9166), .IN2(U6355_n1), .QN(WX2095) );
  INVX0 U6356_U2 ( .INP(WX2030), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n9166), .IN2(U6356_n1), .QN(WX2093) );
  INVX0 U6357_U2 ( .INP(test_so15), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n9166), .IN2(U6357_n1), .QN(WX2091) );
  INVX0 U6358_U2 ( .INP(WX2026), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n9171), .IN2(U6358_n1), .QN(WX2089) );
  INVX0 U6359_U2 ( .INP(WX2024), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n9166), .IN2(U6359_n1), .QN(WX2087) );
  INVX0 U6360_U2 ( .INP(WX2022), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n9166), .IN2(U6360_n1), .QN(WX2085) );
  INVX0 U6361_U2 ( .INP(WX2020), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n9166), .IN2(U6361_n1), .QN(WX2083) );
  INVX0 U6362_U2 ( .INP(WX2018), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n9166), .IN2(U6362_n1), .QN(WX2081) );
  INVX0 U6363_U2 ( .INP(WX2016), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n9166), .IN2(U6363_n1), .QN(WX2079) );
  INVX0 U6364_U2 ( .INP(WX2014), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n9166), .IN2(U6364_n1), .QN(WX2077) );
  INVX0 U6365_U2 ( .INP(WX2012), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n9166), .IN2(U6365_n1), .QN(WX2075) );
  INVX0 U6366_U2 ( .INP(WX2010), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n9165), .IN2(U6366_n1), .QN(WX2073) );
  INVX0 U6367_U2 ( .INP(WX2008), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n9165), .IN2(U6367_n1), .QN(WX2071) );
  INVX0 U6368_U2 ( .INP(WX2006), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n9165), .IN2(U6368_n1), .QN(WX2069) );
  INVX0 U6369_U2 ( .INP(WX2004), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n9165), .IN2(U6369_n1), .QN(WX2067) );
  INVX0 U6370_U2 ( .INP(WX2002), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n9165), .IN2(U6370_n1), .QN(WX2065) );
  INVX0 U6371_U2 ( .INP(WX2000), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n9165), .IN2(U6371_n1), .QN(WX2063) );
  INVX0 U6372_U2 ( .INP(WX1998), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n9165), .IN2(U6372_n1), .QN(WX2061) );
  INVX0 U6373_U2 ( .INP(WX1996), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n9165), .IN2(U6373_n1), .QN(WX2059) );
  INVX0 U6374_U2 ( .INP(WX1994), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n9165), .IN2(U6374_n1), .QN(WX2057) );
  INVX0 U6375_U2 ( .INP(test_so14), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n9165), .IN2(U6375_n1), .QN(WX2055) );
  INVX0 U6376_U2 ( .INP(WX1990), .ZN(U6376_n1) );
  NOR2X0 U6376_U1 ( .IN1(n9165), .IN2(U6376_n1), .QN(WX2053) );
  INVX0 U6377_U2 ( .INP(WX1988), .ZN(U6377_n1) );
  NOR2X0 U6377_U1 ( .IN1(n9165), .IN2(U6377_n1), .QN(WX2051) );
  INVX0 U6378_U2 ( .INP(WX1986), .ZN(U6378_n1) );
  NOR2X0 U6378_U1 ( .IN1(n9165), .IN2(U6378_n1), .QN(WX2049) );
  INVX0 U6379_U2 ( .INP(WX1984), .ZN(U6379_n1) );
  NOR2X0 U6379_U1 ( .IN1(n9164), .IN2(U6379_n1), .QN(WX2047) );
  INVX0 U6380_U2 ( .INP(WX1982), .ZN(U6380_n1) );
  NOR2X0 U6380_U1 ( .IN1(n9164), .IN2(U6380_n1), .QN(WX2045) );
  INVX0 U6381_U2 ( .INP(WX1980), .ZN(U6381_n1) );
  NOR2X0 U6381_U1 ( .IN1(n9164), .IN2(U6381_n1), .QN(WX2043) );
  INVX0 U6382_U2 ( .INP(WX1978), .ZN(U6382_n1) );
  NOR2X0 U6382_U1 ( .IN1(n9164), .IN2(U6382_n1), .QN(WX2041) );
  INVX0 U6383_U2 ( .INP(WX1976), .ZN(U6383_n1) );
  NOR2X0 U6383_U1 ( .IN1(n9164), .IN2(U6383_n1), .QN(WX2039) );
  INVX0 U6384_U2 ( .INP(WX1974), .ZN(U6384_n1) );
  NOR2X0 U6384_U1 ( .IN1(n9164), .IN2(U6384_n1), .QN(WX2037) );
  INVX0 U6385_U2 ( .INP(WX1972), .ZN(U6385_n1) );
  NOR2X0 U6385_U1 ( .IN1(n9164), .IN2(U6385_n1), .QN(WX2035) );
  INVX0 U6386_U2 ( .INP(WX1970), .ZN(U6386_n1) );
  NOR2X0 U6386_U1 ( .IN1(n9164), .IN2(U6386_n1), .QN(WX2033) );
  INVX0 U6387_U2 ( .INP(WX835), .ZN(U6387_n1) );
  NOR2X0 U6387_U1 ( .IN1(n9168), .IN2(U6387_n1), .QN(WX898) );
  INVX0 U6388_U2 ( .INP(WX833), .ZN(U6388_n1) );
  NOR2X0 U6388_U1 ( .IN1(n9171), .IN2(U6388_n1), .QN(WX896) );
  INVX0 U6389_U2 ( .INP(test_so7), .ZN(U6389_n1) );
  NOR2X0 U6389_U1 ( .IN1(n9171), .IN2(U6389_n1), .QN(WX894) );
  INVX0 U6390_U2 ( .INP(WX829), .ZN(U6390_n1) );
  NOR2X0 U6390_U1 ( .IN1(n9172), .IN2(U6390_n1), .QN(WX892) );
  INVX0 U6391_U2 ( .INP(WX827), .ZN(U6391_n1) );
  NOR2X0 U6391_U1 ( .IN1(n9172), .IN2(U6391_n1), .QN(WX890) );
  INVX0 U6392_U2 ( .INP(WX825), .ZN(U6392_n1) );
  NOR2X0 U6392_U1 ( .IN1(n9172), .IN2(U6392_n1), .QN(WX888) );
  INVX0 U6393_U2 ( .INP(WX823), .ZN(U6393_n1) );
  NOR2X0 U6393_U1 ( .IN1(n9172), .IN2(U6393_n1), .QN(WX886) );
  INVX0 U6394_U2 ( .INP(WX821), .ZN(U6394_n1) );
  NOR2X0 U6394_U1 ( .IN1(n9172), .IN2(U6394_n1), .QN(WX884) );
  INVX0 U6395_U2 ( .INP(WX819), .ZN(U6395_n1) );
  NOR2X0 U6395_U1 ( .IN1(n9172), .IN2(U6395_n1), .QN(WX882) );
  INVX0 U6396_U2 ( .INP(WX817), .ZN(U6396_n1) );
  NOR2X0 U6396_U1 ( .IN1(n9172), .IN2(U6396_n1), .QN(WX880) );
  INVX0 U6397_U2 ( .INP(WX815), .ZN(U6397_n1) );
  NOR2X0 U6397_U1 ( .IN1(n9172), .IN2(U6397_n1), .QN(WX878) );
  INVX0 U6398_U2 ( .INP(WX813), .ZN(U6398_n1) );
  NOR2X0 U6398_U1 ( .IN1(n9172), .IN2(U6398_n1), .QN(WX876) );
  INVX0 U6399_U2 ( .INP(WX811), .ZN(U6399_n1) );
  NOR2X0 U6399_U1 ( .IN1(n9172), .IN2(U6399_n1), .QN(WX874) );
  INVX0 U6400_U2 ( .INP(WX809), .ZN(U6400_n1) );
  NOR2X0 U6400_U1 ( .IN1(n9172), .IN2(U6400_n1), .QN(WX872) );
  INVX0 U6401_U2 ( .INP(WX807), .ZN(U6401_n1) );
  NOR2X0 U6401_U1 ( .IN1(n9172), .IN2(U6401_n1), .QN(WX870) );
  INVX0 U6402_U2 ( .INP(WX805), .ZN(U6402_n1) );
  NOR2X0 U6402_U1 ( .IN1(n9172), .IN2(U6402_n1), .QN(WX868) );
  INVX0 U6403_U2 ( .INP(WX803), .ZN(U6403_n1) );
  NOR2X0 U6403_U1 ( .IN1(n9173), .IN2(U6403_n1), .QN(WX866) );
  INVX0 U6404_U2 ( .INP(WX801), .ZN(U6404_n1) );
  NOR2X0 U6404_U1 ( .IN1(n9173), .IN2(U6404_n1), .QN(WX864) );
  INVX0 U6405_U2 ( .INP(WX799), .ZN(U6405_n1) );
  NOR2X0 U6405_U1 ( .IN1(n9173), .IN2(U6405_n1), .QN(WX862) );
  INVX0 U6406_U2 ( .INP(WX797), .ZN(U6406_n1) );
  NOR2X0 U6406_U1 ( .IN1(n9173), .IN2(U6406_n1), .QN(WX860) );
  INVX0 U6407_U2 ( .INP(test_so6), .ZN(U6407_n1) );
  NOR2X0 U6407_U1 ( .IN1(n9173), .IN2(U6407_n1), .QN(WX858) );
  INVX0 U6408_U2 ( .INP(WX793), .ZN(U6408_n1) );
  NOR2X0 U6408_U1 ( .IN1(n9173), .IN2(U6408_n1), .QN(WX856) );
  INVX0 U6409_U2 ( .INP(WX791), .ZN(U6409_n1) );
  NOR2X0 U6409_U1 ( .IN1(n9173), .IN2(U6409_n1), .QN(WX854) );
  INVX0 U6410_U2 ( .INP(WX789), .ZN(U6410_n1) );
  NOR2X0 U6410_U1 ( .IN1(n9173), .IN2(U6410_n1), .QN(WX852) );
  INVX0 U6411_U2 ( .INP(WX787), .ZN(U6411_n1) );
  NOR2X0 U6411_U1 ( .IN1(n9173), .IN2(U6411_n1), .QN(WX850) );
  INVX0 U6412_U2 ( .INP(WX785), .ZN(U6412_n1) );
  NOR2X0 U6412_U1 ( .IN1(n9173), .IN2(U6412_n1), .QN(WX848) );
  INVX0 U6413_U2 ( .INP(WX783), .ZN(U6413_n1) );
  NOR2X0 U6413_U1 ( .IN1(n9173), .IN2(U6413_n1), .QN(WX846) );
  INVX0 U6414_U2 ( .INP(WX781), .ZN(U6414_n1) );
  NOR2X0 U6414_U1 ( .IN1(n9173), .IN2(U6414_n1), .QN(WX844) );
  INVX0 U6415_U2 ( .INP(WX779), .ZN(U6415_n1) );
  NOR2X0 U6415_U1 ( .IN1(n9173), .IN2(U6415_n1), .QN(WX842) );
  INVX0 U6416_U2 ( .INP(WX777), .ZN(U6416_n1) );
  NOR2X0 U6416_U1 ( .IN1(n9174), .IN2(U6416_n1), .QN(WX840) );
  INVX0 U6417_U2 ( .INP(WX775), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n9174), .IN2(U6417_n1), .QN(WX838) );
  INVX0 U6418_U2 ( .INP(WX773), .ZN(U6418_n1) );
  NOR2X0 U6418_U1 ( .IN1(n9174), .IN2(U6418_n1), .QN(WX836) );
  INVX0 U6419_U2 ( .INP(WX771), .ZN(U6419_n1) );
  NOR2X0 U6419_U1 ( .IN1(n9174), .IN2(U6419_n1), .QN(WX834) );
  INVX0 U6420_U2 ( .INP(WX769), .ZN(U6420_n1) );
  NOR2X0 U6420_U1 ( .IN1(n9174), .IN2(U6420_n1), .QN(WX832) );
  INVX0 U6421_U2 ( .INP(WX767), .ZN(U6421_n1) );
  NOR2X0 U6421_U1 ( .IN1(n9174), .IN2(U6421_n1), .QN(WX830) );
  INVX0 U6422_U2 ( .INP(WX765), .ZN(U6422_n1) );
  NOR2X0 U6422_U1 ( .IN1(n9174), .IN2(U6422_n1), .QN(WX828) );
  INVX0 U6423_U2 ( .INP(WX763), .ZN(U6423_n1) );
  NOR2X0 U6423_U1 ( .IN1(n9174), .IN2(U6423_n1), .QN(WX826) );
  INVX0 U6424_U2 ( .INP(WX761), .ZN(U6424_n1) );
  NOR2X0 U6424_U1 ( .IN1(n9174), .IN2(U6424_n1), .QN(WX824) );
  INVX0 U6425_U2 ( .INP(test_so5), .ZN(U6425_n1) );
  NOR2X0 U6425_U1 ( .IN1(n9174), .IN2(U6425_n1), .QN(WX822) );
  INVX0 U6426_U2 ( .INP(WX757), .ZN(U6426_n1) );
  NOR2X0 U6426_U1 ( .IN1(n9174), .IN2(U6426_n1), .QN(WX820) );
  INVX0 U6427_U2 ( .INP(WX755), .ZN(U6427_n1) );
  NOR2X0 U6427_U1 ( .IN1(n9174), .IN2(U6427_n1), .QN(WX818) );
  INVX0 U6428_U2 ( .INP(WX753), .ZN(U6428_n1) );
  NOR2X0 U6428_U1 ( .IN1(n9174), .IN2(U6428_n1), .QN(WX816) );
  INVX0 U6429_U2 ( .INP(WX751), .ZN(U6429_n1) );
  NOR2X0 U6429_U1 ( .IN1(n9175), .IN2(U6429_n1), .QN(WX814) );
  INVX0 U6430_U2 ( .INP(WX749), .ZN(U6430_n1) );
  NOR2X0 U6430_U1 ( .IN1(n9175), .IN2(U6430_n1), .QN(WX812) );
  INVX0 U6431_U2 ( .INP(WX747), .ZN(U6431_n1) );
  NOR2X0 U6431_U1 ( .IN1(n9175), .IN2(U6431_n1), .QN(WX810) );
  INVX0 U6432_U2 ( .INP(WX745), .ZN(U6432_n1) );
  NOR2X0 U6432_U1 ( .IN1(n9175), .IN2(U6432_n1), .QN(WX808) );
  INVX0 U6433_U2 ( .INP(WX743), .ZN(U6433_n1) );
  NOR2X0 U6433_U1 ( .IN1(n9175), .IN2(U6433_n1), .QN(WX806) );
  INVX0 U6434_U2 ( .INP(WX741), .ZN(U6434_n1) );
  NOR2X0 U6434_U1 ( .IN1(n9175), .IN2(U6434_n1), .QN(WX804) );
  INVX0 U6435_U2 ( .INP(WX739), .ZN(U6435_n1) );
  NOR2X0 U6435_U1 ( .IN1(n9175), .IN2(U6435_n1), .QN(WX802) );
  INVX0 U6436_U2 ( .INP(WX737), .ZN(U6436_n1) );
  NOR2X0 U6436_U1 ( .IN1(n9175), .IN2(U6436_n1), .QN(WX800) );
  INVX0 U6437_U2 ( .INP(WX735), .ZN(U6437_n1) );
  NOR2X0 U6437_U1 ( .IN1(n9175), .IN2(U6437_n1), .QN(WX798) );
  INVX0 U6438_U2 ( .INP(WX733), .ZN(U6438_n1) );
  NOR2X0 U6438_U1 ( .IN1(n9175), .IN2(U6438_n1), .QN(WX796) );
  INVX0 U6439_U2 ( .INP(WX731), .ZN(U6439_n1) );
  NOR2X0 U6439_U1 ( .IN1(n9175), .IN2(U6439_n1), .QN(WX794) );
  INVX0 U6440_U2 ( .INP(WX729), .ZN(U6440_n1) );
  NOR2X0 U6440_U1 ( .IN1(n9175), .IN2(U6440_n1), .QN(WX792) );
  INVX0 U6441_U2 ( .INP(WX727), .ZN(U6441_n1) );
  NOR2X0 U6441_U1 ( .IN1(n9175), .IN2(U6441_n1), .QN(WX790) );
  INVX0 U6442_U2 ( .INP(WX725), .ZN(U6442_n1) );
  NOR2X0 U6442_U1 ( .IN1(n9176), .IN2(U6442_n1), .QN(WX788) );
  INVX0 U6443_U2 ( .INP(test_so4), .ZN(U6443_n1) );
  NOR2X0 U6443_U1 ( .IN1(n9176), .IN2(U6443_n1), .QN(WX786) );
  INVX0 U6444_U2 ( .INP(WX721), .ZN(U6444_n1) );
  NOR2X0 U6444_U1 ( .IN1(n9176), .IN2(U6444_n1), .QN(WX784) );
  INVX0 U6445_U2 ( .INP(WX719), .ZN(U6445_n1) );
  NOR2X0 U6445_U1 ( .IN1(n9176), .IN2(U6445_n1), .QN(WX782) );
  INVX0 U6446_U2 ( .INP(WX717), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n9176), .IN2(U6446_n1), .QN(WX780) );
  INVX0 U6447_U2 ( .INP(WX715), .ZN(U6447_n1) );
  NOR2X0 U6447_U1 ( .IN1(n9176), .IN2(U6447_n1), .QN(WX778) );
  INVX0 U6448_U2 ( .INP(WX713), .ZN(U6448_n1) );
  NOR2X0 U6448_U1 ( .IN1(n9176), .IN2(U6448_n1), .QN(WX776) );
  INVX0 U6449_U2 ( .INP(WX711), .ZN(U6449_n1) );
  NOR2X0 U6449_U1 ( .IN1(n9176), .IN2(U6449_n1), .QN(WX774) );
  INVX0 U6450_U2 ( .INP(WX709), .ZN(U6450_n1) );
  NOR2X0 U6450_U1 ( .IN1(n9176), .IN2(U6450_n1), .QN(WX772) );
  INVX0 U6451_U2 ( .INP(WX707), .ZN(U6451_n1) );
  NOR2X0 U6451_U1 ( .IN1(n9176), .IN2(U6451_n1), .QN(WX770) );
  INVX0 U6452_U2 ( .INP(WX705), .ZN(U6452_n1) );
  NOR2X0 U6452_U1 ( .IN1(n9176), .IN2(U6452_n1), .QN(WX768) );
  INVX0 U6453_U2 ( .INP(WX703), .ZN(U6453_n1) );
  NOR2X0 U6453_U1 ( .IN1(n9176), .IN2(U6453_n1), .QN(WX766) );
  INVX0 U6454_U2 ( .INP(WX701), .ZN(U6454_n1) );
  NOR2X0 U6454_U1 ( .IN1(n9176), .IN2(U6454_n1), .QN(WX764) );
  INVX0 U6455_U2 ( .INP(WX699), .ZN(U6455_n1) );
  NOR2X0 U6455_U1 ( .IN1(n9177), .IN2(U6455_n1), .QN(WX762) );
  INVX0 U6456_U2 ( .INP(WX697), .ZN(U6456_n1) );
  NOR2X0 U6456_U1 ( .IN1(n9177), .IN2(U6456_n1), .QN(WX760) );
  INVX0 U6457_U2 ( .INP(WX695), .ZN(U6457_n1) );
  NOR2X0 U6457_U1 ( .IN1(n9177), .IN2(U6457_n1), .QN(WX758) );
  INVX0 U6458_U2 ( .INP(WX693), .ZN(U6458_n1) );
  NOR2X0 U6458_U1 ( .IN1(n9177), .IN2(U6458_n1), .QN(WX756) );
  INVX0 U6459_U2 ( .INP(WX691), .ZN(U6459_n1) );
  NOR2X0 U6459_U1 ( .IN1(n9177), .IN2(U6459_n1), .QN(WX754) );
  INVX0 U6460_U2 ( .INP(WX689), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(n9177), .IN2(U6460_n1), .QN(WX752) );
  INVX0 U6461_U2 ( .INP(test_so3), .ZN(U6461_n1) );
  NOR2X0 U6461_U1 ( .IN1(n9177), .IN2(U6461_n1), .QN(WX750) );
  INVX0 U6462_U2 ( .INP(WX685), .ZN(U6462_n1) );
  NOR2X0 U6462_U1 ( .IN1(n9177), .IN2(U6462_n1), .QN(WX748) );
  INVX0 U6463_U2 ( .INP(WX683), .ZN(U6463_n1) );
  NOR2X0 U6463_U1 ( .IN1(n9177), .IN2(U6463_n1), .QN(WX746) );
  INVX0 U6464_U2 ( .INP(WX681), .ZN(U6464_n1) );
  NOR2X0 U6464_U1 ( .IN1(n9177), .IN2(U6464_n1), .QN(WX744) );
  INVX0 U6465_U2 ( .INP(WX679), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n9177), .IN2(U6465_n1), .QN(WX742) );
  INVX0 U6466_U2 ( .INP(WX677), .ZN(U6466_n1) );
  NOR2X0 U6466_U1 ( .IN1(n9177), .IN2(U6466_n1), .QN(WX740) );
  INVX0 U6467_U2 ( .INP(WX675), .ZN(U6467_n1) );
  NOR2X0 U6467_U1 ( .IN1(n9177), .IN2(U6467_n1), .QN(WX738) );
  INVX0 U6468_U2 ( .INP(WX673), .ZN(U6468_n1) );
  NOR2X0 U6468_U1 ( .IN1(n9178), .IN2(U6468_n1), .QN(WX736) );
  INVX0 U6469_U2 ( .INP(WX671), .ZN(U6469_n1) );
  NOR2X0 U6469_U1 ( .IN1(n9178), .IN2(U6469_n1), .QN(WX734) );
  INVX0 U6470_U2 ( .INP(WX669), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n9178), .IN2(U6470_n1), .QN(WX732) );
  INVX0 U6471_U2 ( .INP(WX667), .ZN(U6471_n1) );
  NOR2X0 U6471_U1 ( .IN1(n9178), .IN2(U6471_n1), .QN(WX730) );
  INVX0 U6472_U2 ( .INP(WX665), .ZN(U6472_n1) );
  NOR2X0 U6472_U1 ( .IN1(n9178), .IN2(U6472_n1), .QN(WX728) );
  INVX0 U6473_U2 ( .INP(WX663), .ZN(U6473_n1) );
  NOR2X0 U6473_U1 ( .IN1(n9178), .IN2(U6473_n1), .QN(WX726) );
  INVX0 U6474_U2 ( .INP(WX661), .ZN(U6474_n1) );
  NOR2X0 U6474_U1 ( .IN1(n9178), .IN2(U6474_n1), .QN(WX724) );
  INVX0 U6475_U2 ( .INP(WX659), .ZN(U6475_n1) );
  NOR2X0 U6475_U1 ( .IN1(n9178), .IN2(U6475_n1), .QN(WX722) );
  INVX0 U6476_U2 ( .INP(WX657), .ZN(U6476_n1) );
  NOR2X0 U6476_U1 ( .IN1(n9178), .IN2(U6476_n1), .QN(WX720) );
  INVX0 U6477_U2 ( .INP(WX655), .ZN(U6477_n1) );
  NOR2X0 U6477_U1 ( .IN1(n9178), .IN2(U6477_n1), .QN(WX718) );
  INVX0 U6478_U2 ( .INP(WX653), .ZN(U6478_n1) );
  NOR2X0 U6478_U1 ( .IN1(n9178), .IN2(U6478_n1), .QN(WX716) );
  INVX0 U6479_U2 ( .INP(test_so2), .ZN(U6479_n1) );
  NOR2X0 U6479_U1 ( .IN1(n9178), .IN2(U6479_n1), .QN(WX714) );
  INVX0 U6480_U2 ( .INP(WX649), .ZN(U6480_n1) );
  NOR2X0 U6480_U1 ( .IN1(n9178), .IN2(U6480_n1), .QN(WX712) );
  INVX0 U6481_U2 ( .INP(WX647), .ZN(U6481_n1) );
  NOR2X0 U6481_U1 ( .IN1(n9179), .IN2(U6481_n1), .QN(WX710) );
  INVX0 U6482_U2 ( .INP(WX645), .ZN(U6482_n1) );
  NOR2X0 U6482_U1 ( .IN1(n9179), .IN2(U6482_n1), .QN(WX708) );
endmodule

