module add_mul_mix_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_, 
        c_9_, c_10_, c_11_, c_12_, c_13_, c_14_, c_15_, d_0_, d_1_, d_2_, d_3_, 
        d_4_, d_5_, d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, 
        d_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_, c_9_, c_10_,
         c_11_, c_12_, c_13_, c_14_, c_15_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_,
         d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, d_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319;

  XNOR2_X2 U2188 ( .A(n4180), .B(n4181), .ZN(n2525) );
  XNOR2_X2 U2189 ( .A(n4198), .B(n4199), .ZN(n3990) );
  XOR2_X2 U2190 ( .A(n4171), .B(n4172), .Z(n2542) );
  XNOR2_X2 U2191 ( .A(n3575), .B(n3576), .ZN(n3317) );
  XNOR2_X2 U2192 ( .A(n3699), .B(n3700), .ZN(n3432) );
  XNOR2_X2 U2193 ( .A(n3321), .B(n3322), .ZN(n3062) );
  XNOR2_X2 U2194 ( .A(n4195), .B(n4196), .ZN(n2497) );
  XNOR2_X2 U2195 ( .A(n2941), .B(n2942), .ZN(n2688) );
  XNOR2_X2 U2196 ( .A(n4049), .B(n4050), .ZN(n3748) );
  XNOR2_X2 U2197 ( .A(n4183), .B(n4184), .ZN(n2406) );
  XNOR2_X2 U2198 ( .A(n3824), .B(n3825), .ZN(n3571) );
  XNOR2_X2 U2199 ( .A(n3436), .B(n3437), .ZN(n3185) );
  XNOR2_X2 U2200 ( .A(n4188), .B(n4189), .ZN(n2388) );
  NOR2_X2 U2201 ( .A1(n4167), .A2(n4165), .ZN(n2210) );
  XNOR2_X2 U2202 ( .A(n4175), .B(n4176), .ZN(n2429) );
  XNOR2_X2 U2203 ( .A(n4178), .B(n4179), .ZN(n2424) );
  XNOR2_X2 U2204 ( .A(n4190), .B(n4191), .ZN(n2508) );
  XNOR2_X2 U2205 ( .A(n4193), .B(n4194), .ZN(n2369) );
  XNOR2_X2 U2206 ( .A(n3189), .B(n3190), .ZN(n2937) );
  XNOR2_X2 U2207 ( .A(n2692), .B(n2693), .ZN(n2454) );
  XNOR2_X2 U2208 ( .A(n3934), .B(n3935), .ZN(n3695) );
  XNOR2_X2 U2209 ( .A(n2810), .B(n2811), .ZN(n2551) );
  XNOR2_X2 U2210 ( .A(n4185), .B(n4186), .ZN(n2396) );
  XNOR2_X2 U2211 ( .A(n4204), .B(n4267), .ZN(n3929) );
  XOR2_X2 U2212 ( .A(n4165), .B(n4166), .Z(n2205) );
  XNOR2_X2 U2213 ( .A(n3066), .B(n3067), .ZN(n2806) );
  XNOR2_X2 U2214 ( .A(n4208), .B(n4209), .ZN(n2303) );
  XOR2_X1 U2215 ( .A(n2156), .B(n2157), .Z(Result_9_) );
  NAND2_X1 U2216 ( .A1(n2158), .A2(n2159), .ZN(n2157) );
  NAND2_X1 U2217 ( .A1(n2160), .A2(n2161), .ZN(n2156) );
  NAND2_X1 U2218 ( .A1(n2162), .A2(n2163), .ZN(n2161) );
  NAND2_X1 U2219 ( .A1(n2164), .A2(n2165), .ZN(n2162) );
  XOR2_X1 U2220 ( .A(n2166), .B(n2167), .Z(Result_8_) );
  XOR2_X1 U2221 ( .A(n2168), .B(n2169), .Z(Result_7_) );
  NAND2_X1 U2222 ( .A1(n2170), .A2(n2171), .ZN(n2169) );
  NAND2_X1 U2223 ( .A1(n2172), .A2(n2173), .ZN(n2171) );
  NAND2_X1 U2224 ( .A1(n2174), .A2(n2175), .ZN(n2172) );
  XOR2_X1 U2225 ( .A(n2176), .B(n2177), .Z(Result_6_) );
  XOR2_X1 U2226 ( .A(n2178), .B(n2179), .Z(Result_5_) );
  NAND2_X1 U2227 ( .A1(n2177), .A2(n2176), .ZN(n2179) );
  NAND2_X1 U2228 ( .A1(n2180), .A2(n2181), .ZN(n2178) );
  NAND2_X1 U2229 ( .A1(n2182), .A2(n2183), .ZN(n2180) );
  NAND2_X1 U2230 ( .A1(n2184), .A2(n2185), .ZN(n2183) );
  XOR2_X1 U2231 ( .A(n2186), .B(n2187), .Z(Result_4_) );
  XNOR2_X1 U2232 ( .A(n2188), .B(n2189), .ZN(Result_3_) );
  NAND2_X1 U2233 ( .A1(n2186), .A2(n2187), .ZN(n2189) );
  NOR2_X1 U2234 ( .A1(n2190), .A2(n2191), .ZN(n2188) );
  NOR2_X1 U2235 ( .A1(n2192), .A2(n2193), .ZN(n2190) );
  NOR2_X1 U2236 ( .A1(n2194), .A2(n2195), .ZN(n2192) );
  NOR2_X1 U2237 ( .A1(n2196), .A2(n2197), .ZN(Result_31_) );
  NAND2_X1 U2238 ( .A1(n2198), .A2(n2199), .ZN(Result_30_) );
  NAND2_X1 U2239 ( .A1(n2200), .A2(n2201), .ZN(n2199) );
  NAND2_X1 U2240 ( .A1(n2202), .A2(n2203), .ZN(n2201) );
  NAND2_X1 U2241 ( .A1(n2204), .A2(n2205), .ZN(n2203) );
  NAND2_X1 U2242 ( .A1(n2206), .A2(n2207), .ZN(n2198) );
  NAND2_X1 U2243 ( .A1(n2208), .A2(n2209), .ZN(n2207) );
  NAND2_X1 U2244 ( .A1(n2196), .A2(n2210), .ZN(n2209) );
  XOR2_X1 U2245 ( .A(n2211), .B(n2212), .Z(Result_2_) );
  XNOR2_X1 U2246 ( .A(n2213), .B(n2214), .ZN(Result_29_) );
  XOR2_X1 U2247 ( .A(n2215), .B(n2216), .Z(n2214) );
  XNOR2_X1 U2248 ( .A(n2217), .B(n2218), .ZN(Result_28_) );
  NAND2_X1 U2249 ( .A1(n2219), .A2(n2220), .ZN(n2217) );
  XOR2_X1 U2250 ( .A(n2221), .B(n2222), .Z(Result_27_) );
  XOR2_X1 U2251 ( .A(n2223), .B(n2224), .Z(n2221) );
  XOR2_X1 U2252 ( .A(n2225), .B(n2226), .Z(Result_26_) );
  XOR2_X1 U2253 ( .A(n2227), .B(n2228), .Z(n2226) );
  XOR2_X1 U2254 ( .A(n2229), .B(n2230), .Z(Result_25_) );
  XOR2_X1 U2255 ( .A(n2231), .B(n2232), .Z(n2229) );
  XOR2_X1 U2256 ( .A(n2233), .B(n2234), .Z(Result_24_) );
  XNOR2_X1 U2257 ( .A(n2235), .B(n2236), .ZN(n2234) );
  XOR2_X1 U2258 ( .A(n2237), .B(n2238), .Z(Result_23_) );
  XOR2_X1 U2259 ( .A(n2239), .B(n2240), .Z(n2238) );
  XOR2_X1 U2260 ( .A(n2241), .B(n2242), .Z(Result_22_) );
  XOR2_X1 U2261 ( .A(n2243), .B(n2244), .Z(n2242) );
  XNOR2_X1 U2262 ( .A(n2245), .B(n2246), .ZN(Result_21_) );
  XNOR2_X1 U2263 ( .A(n2247), .B(n2248), .ZN(n2246) );
  XOR2_X1 U2264 ( .A(n2249), .B(n2250), .Z(Result_20_) );
  XNOR2_X1 U2265 ( .A(n2251), .B(n2252), .ZN(n2250) );
  XOR2_X1 U2266 ( .A(n2253), .B(n2254), .Z(Result_1_) );
  NAND2_X1 U2267 ( .A1(n2212), .A2(n2211), .ZN(n2254) );
  NAND2_X1 U2268 ( .A1(n2255), .A2(n2256), .ZN(n2253) );
  INV_X1 U2269 ( .A(n2257), .ZN(n2256) );
  NOR2_X1 U2270 ( .A1(n2258), .A2(n2259), .ZN(n2257) );
  XNOR2_X1 U2271 ( .A(n2260), .B(n2261), .ZN(Result_19_) );
  XNOR2_X1 U2272 ( .A(n2262), .B(n2263), .ZN(n2261) );
  XNOR2_X1 U2273 ( .A(n2264), .B(n2265), .ZN(Result_18_) );
  NAND2_X1 U2274 ( .A1(n2266), .A2(n2267), .ZN(n2264) );
  XOR2_X1 U2275 ( .A(n2268), .B(n2269), .Z(Result_17_) );
  XOR2_X1 U2276 ( .A(n2270), .B(n2271), .Z(n2268) );
  XNOR2_X1 U2277 ( .A(n2272), .B(n2273), .ZN(Result_16_) );
  XNOR2_X1 U2278 ( .A(n2274), .B(n2275), .ZN(n2273) );
  XNOR2_X1 U2279 ( .A(n2276), .B(n2277), .ZN(Result_15_) );
  NOR2_X1 U2280 ( .A1(n2278), .A2(n2279), .ZN(Result_14_) );
  NOR2_X1 U2281 ( .A1(n2280), .A2(n2281), .ZN(n2279) );
  NOR2_X1 U2282 ( .A1(n2282), .A2(n2277), .ZN(n2280) );
  XOR2_X1 U2283 ( .A(n2278), .B(n2283), .Z(Result_13_) );
  NOR2_X1 U2284 ( .A1(n2284), .A2(n2285), .ZN(n2283) );
  NOR2_X1 U2285 ( .A1(n2286), .A2(n2287), .ZN(n2284) );
  NOR2_X1 U2286 ( .A1(n2288), .A2(n2289), .ZN(n2287) );
  XOR2_X1 U2287 ( .A(n2290), .B(n2291), .Z(Result_12_) );
  XOR2_X1 U2288 ( .A(n2292), .B(n2293), .Z(Result_11_) );
  NAND2_X1 U2289 ( .A1(n2291), .A2(n2290), .ZN(n2293) );
  NAND2_X1 U2290 ( .A1(n2294), .A2(n2295), .ZN(n2292) );
  NAND2_X1 U2291 ( .A1(n2296), .A2(n2297), .ZN(n2295) );
  INV_X1 U2292 ( .A(n2298), .ZN(n2297) );
  NAND2_X1 U2293 ( .A1(n2299), .A2(n2300), .ZN(n2296) );
  XOR2_X1 U2294 ( .A(n2159), .B(n2158), .Z(Result_10_) );
  NAND3_X1 U2295 ( .A1(n2301), .A2(n2258), .A3(n2302), .ZN(Result_0_) );
  NAND2_X1 U2296 ( .A1(n2303), .A2(n2259), .ZN(n2302) );
  NAND4_X1 U2297 ( .A1(n2304), .A2(n2305), .A3(n2303), .A4(n2306), .ZN(n2258)
         );
  NAND3_X1 U2298 ( .A1(n2255), .A2(n2211), .A3(n2212), .ZN(n2301) );
  XOR2_X1 U2299 ( .A(n2306), .B(n2304), .Z(n2212) );
  NAND3_X1 U2300 ( .A1(n2307), .A2(n2308), .A3(n2309), .ZN(n2211) );
  NAND2_X1 U2301 ( .A1(n2310), .A2(n2311), .ZN(n2309) );
  INV_X1 U2302 ( .A(n2191), .ZN(n2308) );
  NOR3_X1 U2303 ( .A1(n2312), .A2(n2194), .A3(n2195), .ZN(n2191) );
  INV_X1 U2304 ( .A(n2193), .ZN(n2312) );
  NAND3_X1 U2305 ( .A1(n2187), .A2(n2186), .A3(n2193), .ZN(n2307) );
  XOR2_X1 U2306 ( .A(n2311), .B(n2310), .Z(n2193) );
  XNOR2_X1 U2307 ( .A(n2313), .B(n2314), .ZN(n2310) );
  NAND2_X1 U2308 ( .A1(n2315), .A2(n2316), .ZN(n2313) );
  NAND2_X1 U2309 ( .A1(n2317), .A2(n2318), .ZN(n2311) );
  NAND2_X1 U2310 ( .A1(n2319), .A2(n2320), .ZN(n2318) );
  NAND2_X1 U2311 ( .A1(n2321), .A2(n2322), .ZN(n2320) );
  INV_X1 U2312 ( .A(n2323), .ZN(n2317) );
  NOR2_X1 U2313 ( .A1(n2321), .A2(n2322), .ZN(n2323) );
  NAND3_X1 U2314 ( .A1(n2324), .A2(n2181), .A3(n2325), .ZN(n2186) );
  NAND3_X1 U2315 ( .A1(n2176), .A2(n2177), .A3(n2326), .ZN(n2325) );
  NAND3_X1 U2316 ( .A1(n2327), .A2(n2170), .A3(n2328), .ZN(n2177) );
  NAND2_X1 U2317 ( .A1(n2329), .A2(n2330), .ZN(n2328) );
  INV_X1 U2318 ( .A(n2168), .ZN(n2329) );
  NAND2_X1 U2319 ( .A1(n2167), .A2(n2166), .ZN(n2168) );
  NAND3_X1 U2320 ( .A1(n2331), .A2(n2160), .A3(n2332), .ZN(n2166) );
  NAND3_X1 U2321 ( .A1(n2158), .A2(n2159), .A3(n2333), .ZN(n2332) );
  NAND3_X1 U2322 ( .A1(n2334), .A2(n2294), .A3(n2335), .ZN(n2159) );
  NAND3_X1 U2323 ( .A1(n2291), .A2(n2290), .A3(n2298), .ZN(n2335) );
  NAND3_X1 U2324 ( .A1(n2336), .A2(n2337), .A3(n2338), .ZN(n2290) );
  NAND2_X1 U2325 ( .A1(n2278), .A2(n2286), .ZN(n2338) );
  INV_X1 U2326 ( .A(n2339), .ZN(n2286) );
  NOR3_X1 U2327 ( .A1(n2340), .A2(n2282), .A3(n2277), .ZN(n2278) );
  XOR2_X1 U2328 ( .A(n2341), .B(n2342), .Z(n2277) );
  XNOR2_X1 U2329 ( .A(n2343), .B(n2344), .ZN(n2341) );
  NOR2_X1 U2330 ( .A1(n2345), .A2(n2204), .ZN(n2344) );
  INV_X1 U2331 ( .A(n2276), .ZN(n2282) );
  NAND2_X1 U2332 ( .A1(n2346), .A2(n2347), .ZN(n2276) );
  NAND2_X1 U2333 ( .A1(n2275), .A2(n2348), .ZN(n2347) );
  INV_X1 U2334 ( .A(n2349), .ZN(n2348) );
  NOR2_X1 U2335 ( .A1(n2274), .A2(n2272), .ZN(n2349) );
  NOR2_X1 U2336 ( .A1(n2196), .A2(n2345), .ZN(n2275) );
  NAND2_X1 U2337 ( .A1(n2272), .A2(n2274), .ZN(n2346) );
  NAND2_X1 U2338 ( .A1(n2350), .A2(n2351), .ZN(n2274) );
  NAND2_X1 U2339 ( .A1(n2271), .A2(n2352), .ZN(n2351) );
  INV_X1 U2340 ( .A(n2353), .ZN(n2352) );
  NOR2_X1 U2341 ( .A1(n2270), .A2(n2269), .ZN(n2353) );
  NOR2_X1 U2342 ( .A1(n2354), .A2(n2196), .ZN(n2271) );
  NAND2_X1 U2343 ( .A1(n2269), .A2(n2270), .ZN(n2350) );
  NAND2_X1 U2344 ( .A1(n2266), .A2(n2355), .ZN(n2270) );
  NAND2_X1 U2345 ( .A1(n2265), .A2(n2267), .ZN(n2355) );
  NAND2_X1 U2346 ( .A1(n2356), .A2(n2357), .ZN(n2267) );
  NAND2_X1 U2347 ( .A1(n2358), .A2(n2200), .ZN(n2357) );
  INV_X1 U2348 ( .A(n2359), .ZN(n2356) );
  XNOR2_X1 U2349 ( .A(n2360), .B(n2361), .ZN(n2265) );
  XNOR2_X1 U2350 ( .A(n2362), .B(n2363), .ZN(n2360) );
  NAND2_X1 U2351 ( .A1(n2358), .A2(n2359), .ZN(n2266) );
  NAND2_X1 U2352 ( .A1(n2364), .A2(n2365), .ZN(n2359) );
  NAND2_X1 U2353 ( .A1(n2263), .A2(n2366), .ZN(n2365) );
  NAND2_X1 U2354 ( .A1(n2367), .A2(n2368), .ZN(n2366) );
  INV_X1 U2355 ( .A(n2262), .ZN(n2368) );
  INV_X1 U2356 ( .A(n2260), .ZN(n2367) );
  NOR2_X1 U2357 ( .A1(n2369), .A2(n2196), .ZN(n2263) );
  NAND2_X1 U2358 ( .A1(n2262), .A2(n2260), .ZN(n2364) );
  XNOR2_X1 U2359 ( .A(n2370), .B(n2371), .ZN(n2260) );
  XNOR2_X1 U2360 ( .A(n2372), .B(n2373), .ZN(n2370) );
  NOR2_X1 U2361 ( .A1(n2374), .A2(n2375), .ZN(n2262) );
  INV_X1 U2362 ( .A(n2376), .ZN(n2375) );
  NAND2_X1 U2363 ( .A1(n2377), .A2(n2252), .ZN(n2376) );
  NAND2_X1 U2364 ( .A1(n2378), .A2(n2200), .ZN(n2252) );
  NAND2_X1 U2365 ( .A1(n2249), .A2(n2251), .ZN(n2377) );
  NOR2_X1 U2366 ( .A1(n2251), .A2(n2249), .ZN(n2374) );
  XOR2_X1 U2367 ( .A(n2379), .B(n2380), .Z(n2249) );
  XOR2_X1 U2368 ( .A(n2381), .B(n2382), .Z(n2380) );
  NAND2_X1 U2369 ( .A1(n2383), .A2(n2384), .ZN(n2251) );
  NAND2_X1 U2370 ( .A1(n2248), .A2(n2385), .ZN(n2384) );
  NAND2_X1 U2371 ( .A1(n2386), .A2(n2387), .ZN(n2385) );
  INV_X1 U2372 ( .A(n2247), .ZN(n2387) );
  INV_X1 U2373 ( .A(n2245), .ZN(n2386) );
  NOR2_X1 U2374 ( .A1(n2388), .A2(n2196), .ZN(n2248) );
  NAND2_X1 U2375 ( .A1(n2247), .A2(n2245), .ZN(n2383) );
  XNOR2_X1 U2376 ( .A(n2389), .B(n2390), .ZN(n2245) );
  XNOR2_X1 U2377 ( .A(n2391), .B(n2392), .ZN(n2389) );
  NOR2_X1 U2378 ( .A1(n2393), .A2(n2394), .ZN(n2247) );
  NOR2_X1 U2379 ( .A1(n2395), .A2(n2243), .ZN(n2394) );
  NOR2_X1 U2380 ( .A1(n2396), .A2(n2196), .ZN(n2243) );
  NOR2_X1 U2381 ( .A1(n2241), .A2(n2244), .ZN(n2395) );
  INV_X1 U2382 ( .A(n2397), .ZN(n2393) );
  NAND2_X1 U2383 ( .A1(n2244), .A2(n2241), .ZN(n2397) );
  XOR2_X1 U2384 ( .A(n2398), .B(n2399), .Z(n2241) );
  XNOR2_X1 U2385 ( .A(n2400), .B(n2401), .ZN(n2398) );
  NOR2_X1 U2386 ( .A1(n2402), .A2(n2403), .ZN(n2244) );
  INV_X1 U2387 ( .A(n2404), .ZN(n2403) );
  NAND2_X1 U2388 ( .A1(n2240), .A2(n2405), .ZN(n2404) );
  NAND2_X1 U2389 ( .A1(n2237), .A2(n2239), .ZN(n2405) );
  NOR2_X1 U2390 ( .A1(n2406), .A2(n2196), .ZN(n2240) );
  NOR2_X1 U2391 ( .A1(n2239), .A2(n2237), .ZN(n2402) );
  XOR2_X1 U2392 ( .A(n2407), .B(n2408), .Z(n2237) );
  XNOR2_X1 U2393 ( .A(n2409), .B(n2410), .ZN(n2407) );
  NAND2_X1 U2394 ( .A1(n2411), .A2(n2412), .ZN(n2239) );
  NAND2_X1 U2395 ( .A1(n2413), .A2(n2235), .ZN(n2412) );
  NAND2_X1 U2396 ( .A1(n2414), .A2(n2200), .ZN(n2235) );
  NAND2_X1 U2397 ( .A1(n2233), .A2(n2236), .ZN(n2413) );
  INV_X1 U2398 ( .A(n2415), .ZN(n2411) );
  NOR2_X1 U2399 ( .A1(n2236), .A2(n2233), .ZN(n2415) );
  XNOR2_X1 U2400 ( .A(n2416), .B(n2417), .ZN(n2233) );
  XNOR2_X1 U2401 ( .A(n2418), .B(n2419), .ZN(n2416) );
  NAND2_X1 U2402 ( .A1(n2420), .A2(n2421), .ZN(n2236) );
  NAND2_X1 U2403 ( .A1(n2232), .A2(n2422), .ZN(n2421) );
  INV_X1 U2404 ( .A(n2423), .ZN(n2422) );
  NOR2_X1 U2405 ( .A1(n2231), .A2(n2230), .ZN(n2423) );
  NOR2_X1 U2406 ( .A1(n2424), .A2(n2196), .ZN(n2232) );
  NAND2_X1 U2407 ( .A1(n2230), .A2(n2231), .ZN(n2420) );
  NAND2_X1 U2408 ( .A1(n2425), .A2(n2426), .ZN(n2231) );
  NAND2_X1 U2409 ( .A1(n2227), .A2(n2427), .ZN(n2426) );
  INV_X1 U2410 ( .A(n2428), .ZN(n2427) );
  NOR2_X1 U2411 ( .A1(n2228), .A2(n2225), .ZN(n2428) );
  NOR2_X1 U2412 ( .A1(n2429), .A2(n2196), .ZN(n2227) );
  NAND2_X1 U2413 ( .A1(n2225), .A2(n2228), .ZN(n2425) );
  NAND2_X1 U2414 ( .A1(n2430), .A2(n2431), .ZN(n2228) );
  NAND2_X1 U2415 ( .A1(n2224), .A2(n2432), .ZN(n2431) );
  INV_X1 U2416 ( .A(n2433), .ZN(n2432) );
  NOR2_X1 U2417 ( .A1(n2223), .A2(n2222), .ZN(n2433) );
  NOR2_X1 U2418 ( .A1(n2434), .A2(n2196), .ZN(n2224) );
  NAND2_X1 U2419 ( .A1(n2222), .A2(n2223), .ZN(n2430) );
  NAND2_X1 U2420 ( .A1(n2219), .A2(n2435), .ZN(n2223) );
  NAND2_X1 U2421 ( .A1(n2218), .A2(n2220), .ZN(n2435) );
  NAND2_X1 U2422 ( .A1(n2436), .A2(n2437), .ZN(n2220) );
  NAND2_X1 U2423 ( .A1(n2438), .A2(n2200), .ZN(n2436) );
  XOR2_X1 U2424 ( .A(n2439), .B(n2440), .Z(n2218) );
  XNOR2_X1 U2425 ( .A(n2441), .B(n2442), .ZN(n2440) );
  NAND2_X1 U2426 ( .A1(n2443), .A2(n2438), .ZN(n2219) );
  INV_X1 U2427 ( .A(n2437), .ZN(n2443) );
  NAND2_X1 U2428 ( .A1(n2444), .A2(n2445), .ZN(n2437) );
  NAND2_X1 U2429 ( .A1(n2446), .A2(n2215), .ZN(n2445) );
  NAND2_X1 U2430 ( .A1(n2447), .A2(n2200), .ZN(n2215) );
  NAND2_X1 U2431 ( .A1(n2213), .A2(n2216), .ZN(n2446) );
  INV_X1 U2432 ( .A(n2448), .ZN(n2444) );
  NOR2_X1 U2433 ( .A1(n2216), .A2(n2213), .ZN(n2448) );
  NOR3_X1 U2434 ( .A1(n2196), .A2(n2204), .A3(n2449), .ZN(n2213) );
  INV_X1 U2435 ( .A(n2200), .ZN(n2196) );
  XOR2_X1 U2436 ( .A(c_15_), .B(d_15_), .Z(n2200) );
  NAND2_X1 U2437 ( .A1(n2450), .A2(n2451), .ZN(n2216) );
  NAND2_X1 U2438 ( .A1(n2206), .A2(n2452), .ZN(n2451) );
  NAND2_X1 U2439 ( .A1(n2202), .A2(n2453), .ZN(n2452) );
  NAND2_X1 U2440 ( .A1(n2454), .A2(n2205), .ZN(n2453) );
  NAND2_X1 U2441 ( .A1(n2455), .A2(n2456), .ZN(n2450) );
  NAND2_X1 U2442 ( .A1(n2208), .A2(n2457), .ZN(n2456) );
  NAND2_X1 U2443 ( .A1(n2204), .A2(n2210), .ZN(n2457) );
  XNOR2_X1 U2444 ( .A(n2458), .B(n2459), .ZN(n2222) );
  XNOR2_X1 U2445 ( .A(n2460), .B(n2461), .ZN(n2458) );
  XNOR2_X1 U2446 ( .A(n2462), .B(n2463), .ZN(n2225) );
  XNOR2_X1 U2447 ( .A(n2464), .B(n2465), .ZN(n2462) );
  XNOR2_X1 U2448 ( .A(n2466), .B(n2467), .ZN(n2230) );
  XNOR2_X1 U2449 ( .A(n2468), .B(n2469), .ZN(n2466) );
  XNOR2_X1 U2450 ( .A(n2470), .B(n2471), .ZN(n2269) );
  XNOR2_X1 U2451 ( .A(n2472), .B(n2473), .ZN(n2470) );
  XOR2_X1 U2452 ( .A(n2474), .B(n2475), .Z(n2272) );
  XOR2_X1 U2453 ( .A(n2476), .B(n2477), .Z(n2475) );
  NOR2_X1 U2454 ( .A1(n2204), .A2(n2354), .ZN(n2477) );
  INV_X1 U2455 ( .A(n2281), .ZN(n2340) );
  XOR2_X1 U2456 ( .A(n2288), .B(n2289), .Z(n2281) );
  INV_X1 U2457 ( .A(n2285), .ZN(n2337) );
  NOR3_X1 U2458 ( .A1(n2289), .A2(n2288), .A3(n2339), .ZN(n2285) );
  NAND2_X1 U2459 ( .A1(n2478), .A2(n2336), .ZN(n2339) );
  NAND2_X1 U2460 ( .A1(n2479), .A2(n2480), .ZN(n2478) );
  INV_X1 U2461 ( .A(n2481), .ZN(n2480) );
  XNOR2_X1 U2462 ( .A(n2482), .B(n2483), .ZN(n2479) );
  NOR2_X1 U2463 ( .A1(n2484), .A2(n2485), .ZN(n2288) );
  NOR3_X1 U2464 ( .A1(n2345), .A2(n2486), .A3(n2204), .ZN(n2485) );
  INV_X1 U2465 ( .A(n2487), .ZN(n2486) );
  NAND2_X1 U2466 ( .A1(n2343), .A2(n2342), .ZN(n2487) );
  NOR2_X1 U2467 ( .A1(n2342), .A2(n2343), .ZN(n2484) );
  NOR2_X1 U2468 ( .A1(n2488), .A2(n2489), .ZN(n2343) );
  INV_X1 U2469 ( .A(n2490), .ZN(n2489) );
  NAND3_X1 U2470 ( .A1(n2206), .A2(n2491), .A3(n2492), .ZN(n2490) );
  NAND2_X1 U2471 ( .A1(n2476), .A2(n2474), .ZN(n2491) );
  NOR2_X1 U2472 ( .A1(n2474), .A2(n2476), .ZN(n2488) );
  NOR2_X1 U2473 ( .A1(n2493), .A2(n2494), .ZN(n2476) );
  INV_X1 U2474 ( .A(n2495), .ZN(n2494) );
  NAND2_X1 U2475 ( .A1(n2472), .A2(n2496), .ZN(n2495) );
  NAND2_X1 U2476 ( .A1(n2473), .A2(n2471), .ZN(n2496) );
  NOR2_X1 U2477 ( .A1(n2497), .A2(n2204), .ZN(n2472) );
  NOR2_X1 U2478 ( .A1(n2471), .A2(n2473), .ZN(n2493) );
  INV_X1 U2479 ( .A(n2498), .ZN(n2473) );
  NAND2_X1 U2480 ( .A1(n2499), .A2(n2500), .ZN(n2498) );
  NAND2_X1 U2481 ( .A1(n2363), .A2(n2501), .ZN(n2500) );
  NAND2_X1 U2482 ( .A1(n2362), .A2(n2361), .ZN(n2501) );
  NOR2_X1 U2483 ( .A1(n2369), .A2(n2204), .ZN(n2363) );
  NAND2_X1 U2484 ( .A1(n2502), .A2(n2503), .ZN(n2499) );
  INV_X1 U2485 ( .A(n2362), .ZN(n2503) );
  NOR2_X1 U2486 ( .A1(n2504), .A2(n2505), .ZN(n2362) );
  INV_X1 U2487 ( .A(n2506), .ZN(n2505) );
  NAND2_X1 U2488 ( .A1(n2373), .A2(n2507), .ZN(n2506) );
  NAND2_X1 U2489 ( .A1(n2372), .A2(n2371), .ZN(n2507) );
  NOR2_X1 U2490 ( .A1(n2508), .A2(n2204), .ZN(n2373) );
  NOR2_X1 U2491 ( .A1(n2371), .A2(n2372), .ZN(n2504) );
  NOR2_X1 U2492 ( .A1(n2509), .A2(n2510), .ZN(n2372) );
  INV_X1 U2493 ( .A(n2511), .ZN(n2510) );
  NAND2_X1 U2494 ( .A1(n2382), .A2(n2512), .ZN(n2511) );
  NAND2_X1 U2495 ( .A1(n2381), .A2(n2379), .ZN(n2512) );
  NOR2_X1 U2496 ( .A1(n2388), .A2(n2204), .ZN(n2382) );
  NOR2_X1 U2497 ( .A1(n2379), .A2(n2381), .ZN(n2509) );
  NOR2_X1 U2498 ( .A1(n2513), .A2(n2514), .ZN(n2381) );
  INV_X1 U2499 ( .A(n2515), .ZN(n2514) );
  NAND2_X1 U2500 ( .A1(n2392), .A2(n2516), .ZN(n2515) );
  NAND2_X1 U2501 ( .A1(n2391), .A2(n2390), .ZN(n2516) );
  NOR2_X1 U2502 ( .A1(n2396), .A2(n2204), .ZN(n2392) );
  NOR2_X1 U2503 ( .A1(n2390), .A2(n2391), .ZN(n2513) );
  NOR2_X1 U2504 ( .A1(n2517), .A2(n2518), .ZN(n2391) );
  INV_X1 U2505 ( .A(n2519), .ZN(n2518) );
  NAND2_X1 U2506 ( .A1(n2400), .A2(n2520), .ZN(n2519) );
  NAND2_X1 U2507 ( .A1(n2401), .A2(n2399), .ZN(n2520) );
  NOR2_X1 U2508 ( .A1(n2406), .A2(n2204), .ZN(n2400) );
  NOR2_X1 U2509 ( .A1(n2399), .A2(n2401), .ZN(n2517) );
  NOR2_X1 U2510 ( .A1(n2521), .A2(n2522), .ZN(n2401) );
  INV_X1 U2511 ( .A(n2523), .ZN(n2522) );
  NAND2_X1 U2512 ( .A1(n2410), .A2(n2524), .ZN(n2523) );
  NAND2_X1 U2513 ( .A1(n2409), .A2(n2408), .ZN(n2524) );
  NOR2_X1 U2514 ( .A1(n2525), .A2(n2204), .ZN(n2410) );
  NOR2_X1 U2515 ( .A1(n2408), .A2(n2409), .ZN(n2521) );
  NOR2_X1 U2516 ( .A1(n2526), .A2(n2527), .ZN(n2409) );
  INV_X1 U2517 ( .A(n2528), .ZN(n2527) );
  NAND2_X1 U2518 ( .A1(n2418), .A2(n2529), .ZN(n2528) );
  NAND2_X1 U2519 ( .A1(n2419), .A2(n2417), .ZN(n2529) );
  NOR2_X1 U2520 ( .A1(n2424), .A2(n2204), .ZN(n2418) );
  NOR2_X1 U2521 ( .A1(n2417), .A2(n2419), .ZN(n2526) );
  NOR2_X1 U2522 ( .A1(n2530), .A2(n2531), .ZN(n2419) );
  INV_X1 U2523 ( .A(n2532), .ZN(n2531) );
  NAND2_X1 U2524 ( .A1(n2468), .A2(n2533), .ZN(n2532) );
  NAND2_X1 U2525 ( .A1(n2469), .A2(n2467), .ZN(n2533) );
  NOR2_X1 U2526 ( .A1(n2429), .A2(n2204), .ZN(n2468) );
  NOR2_X1 U2527 ( .A1(n2467), .A2(n2469), .ZN(n2530) );
  NOR2_X1 U2528 ( .A1(n2534), .A2(n2535), .ZN(n2469) );
  INV_X1 U2529 ( .A(n2536), .ZN(n2535) );
  NAND2_X1 U2530 ( .A1(n2464), .A2(n2537), .ZN(n2536) );
  NAND2_X1 U2531 ( .A1(n2465), .A2(n2463), .ZN(n2537) );
  NOR2_X1 U2532 ( .A1(n2434), .A2(n2204), .ZN(n2464) );
  NOR2_X1 U2533 ( .A1(n2463), .A2(n2465), .ZN(n2534) );
  NOR2_X1 U2534 ( .A1(n2538), .A2(n2539), .ZN(n2465) );
  INV_X1 U2535 ( .A(n2540), .ZN(n2539) );
  NAND2_X1 U2536 ( .A1(n2460), .A2(n2541), .ZN(n2540) );
  NAND2_X1 U2537 ( .A1(n2461), .A2(n2459), .ZN(n2541) );
  NOR2_X1 U2538 ( .A1(n2542), .A2(n2204), .ZN(n2460) );
  NOR2_X1 U2539 ( .A1(n2459), .A2(n2461), .ZN(n2538) );
  NOR2_X1 U2540 ( .A1(n2543), .A2(n2544), .ZN(n2461) );
  NOR2_X1 U2541 ( .A1(n2439), .A2(n2545), .ZN(n2544) );
  NOR2_X1 U2542 ( .A1(n2442), .A2(n2441), .ZN(n2545) );
  NAND2_X1 U2543 ( .A1(n2447), .A2(n2206), .ZN(n2439) );
  INV_X1 U2544 ( .A(n2546), .ZN(n2543) );
  NAND2_X1 U2545 ( .A1(n2441), .A2(n2442), .ZN(n2546) );
  NAND2_X1 U2546 ( .A1(n2547), .A2(n2548), .ZN(n2442) );
  NAND2_X1 U2547 ( .A1(n2455), .A2(n2549), .ZN(n2548) );
  NAND2_X1 U2548 ( .A1(n2202), .A2(n2550), .ZN(n2549) );
  NAND2_X1 U2549 ( .A1(n2551), .A2(n2205), .ZN(n2550) );
  NAND2_X1 U2550 ( .A1(n2552), .A2(n2553), .ZN(n2547) );
  NAND2_X1 U2551 ( .A1(n2208), .A2(n2554), .ZN(n2553) );
  NAND2_X1 U2552 ( .A1(n2210), .A2(n2454), .ZN(n2554) );
  NOR3_X1 U2553 ( .A1(n2449), .A2(n2204), .A3(n2454), .ZN(n2441) );
  INV_X1 U2554 ( .A(n2206), .ZN(n2204) );
  XNOR2_X1 U2555 ( .A(n2555), .B(n2556), .ZN(n2206) );
  XOR2_X1 U2556 ( .A(d_14_), .B(c_14_), .Z(n2556) );
  NAND2_X1 U2557 ( .A1(d_15_), .A2(c_15_), .ZN(n2555) );
  XNOR2_X1 U2558 ( .A(n2557), .B(n2558), .ZN(n2459) );
  XNOR2_X1 U2559 ( .A(n2559), .B(n2560), .ZN(n2558) );
  XOR2_X1 U2560 ( .A(n2561), .B(n2562), .Z(n2463) );
  XNOR2_X1 U2561 ( .A(n2563), .B(n2564), .ZN(n2561) );
  XOR2_X1 U2562 ( .A(n2565), .B(n2566), .Z(n2467) );
  XNOR2_X1 U2563 ( .A(n2567), .B(n2568), .ZN(n2565) );
  XOR2_X1 U2564 ( .A(n2569), .B(n2570), .Z(n2417) );
  XNOR2_X1 U2565 ( .A(n2571), .B(n2572), .ZN(n2569) );
  XOR2_X1 U2566 ( .A(n2573), .B(n2574), .Z(n2408) );
  XNOR2_X1 U2567 ( .A(n2575), .B(n2576), .ZN(n2573) );
  XNOR2_X1 U2568 ( .A(n2577), .B(n2578), .ZN(n2399) );
  XOR2_X1 U2569 ( .A(n2579), .B(n2580), .Z(n2577) );
  XNOR2_X1 U2570 ( .A(n2581), .B(n2582), .ZN(n2390) );
  XOR2_X1 U2571 ( .A(n2583), .B(n2584), .Z(n2581) );
  NOR2_X1 U2572 ( .A1(n2406), .A2(n2454), .ZN(n2584) );
  XOR2_X1 U2573 ( .A(n2585), .B(n2586), .Z(n2379) );
  XNOR2_X1 U2574 ( .A(n2587), .B(n2588), .ZN(n2585) );
  NOR2_X1 U2575 ( .A1(n2396), .A2(n2454), .ZN(n2588) );
  XNOR2_X1 U2576 ( .A(n2589), .B(n2590), .ZN(n2371) );
  XNOR2_X1 U2577 ( .A(n2591), .B(n2592), .ZN(n2590) );
  NAND2_X1 U2578 ( .A1(n2455), .A2(n2593), .ZN(n2592) );
  INV_X1 U2579 ( .A(n2361), .ZN(n2502) );
  XOR2_X1 U2580 ( .A(n2594), .B(n2595), .Z(n2361) );
  XNOR2_X1 U2581 ( .A(n2596), .B(n2597), .ZN(n2594) );
  NOR2_X1 U2582 ( .A1(n2508), .A2(n2454), .ZN(n2597) );
  XOR2_X1 U2583 ( .A(n2598), .B(n2599), .Z(n2471) );
  XNOR2_X1 U2584 ( .A(n2600), .B(n2601), .ZN(n2598) );
  NOR2_X1 U2585 ( .A1(n2369), .A2(n2454), .ZN(n2601) );
  XOR2_X1 U2586 ( .A(n2602), .B(n2603), .Z(n2474) );
  XNOR2_X1 U2587 ( .A(n2604), .B(n2605), .ZN(n2602) );
  NOR2_X1 U2588 ( .A1(n2497), .A2(n2454), .ZN(n2605) );
  XOR2_X1 U2589 ( .A(n2606), .B(n2607), .Z(n2342) );
  NAND2_X1 U2590 ( .A1(n2608), .A2(n2609), .ZN(n2606) );
  XNOR2_X1 U2591 ( .A(n2610), .B(n2611), .ZN(n2289) );
  NOR2_X1 U2592 ( .A1(n2612), .A2(n2613), .ZN(n2611) );
  INV_X1 U2593 ( .A(n2614), .ZN(n2613) );
  NOR2_X1 U2594 ( .A1(n2615), .A2(n2616), .ZN(n2612) );
  NOR2_X1 U2595 ( .A1(n2345), .A2(n2454), .ZN(n2615) );
  NAND2_X1 U2596 ( .A1(n2617), .A2(n2481), .ZN(n2336) );
  NAND2_X1 U2597 ( .A1(n2614), .A2(n2618), .ZN(n2481) );
  NAND2_X1 U2598 ( .A1(n2610), .A2(n2619), .ZN(n2618) );
  NAND2_X1 U2599 ( .A1(n2620), .A2(n2621), .ZN(n2619) );
  NAND2_X1 U2600 ( .A1(n2455), .A2(n2303), .ZN(n2621) );
  INV_X1 U2601 ( .A(n2616), .ZN(n2620) );
  XOR2_X1 U2602 ( .A(n2622), .B(n2623), .Z(n2610) );
  XOR2_X1 U2603 ( .A(n2624), .B(n2625), .Z(n2622) );
  NAND2_X1 U2604 ( .A1(n2303), .A2(n2616), .ZN(n2614) );
  NAND2_X1 U2605 ( .A1(n2608), .A2(n2626), .ZN(n2616) );
  NAND2_X1 U2606 ( .A1(n2607), .A2(n2609), .ZN(n2626) );
  NAND2_X1 U2607 ( .A1(n2627), .A2(n2628), .ZN(n2609) );
  NAND2_X1 U2608 ( .A1(n2455), .A2(n2492), .ZN(n2628) );
  INV_X1 U2609 ( .A(n2629), .ZN(n2627) );
  XOR2_X1 U2610 ( .A(n2630), .B(n2631), .Z(n2607) );
  XNOR2_X1 U2611 ( .A(n2632), .B(n2633), .ZN(n2631) );
  NAND2_X1 U2612 ( .A1(n2552), .A2(n2358), .ZN(n2633) );
  NAND2_X1 U2613 ( .A1(n2492), .A2(n2629), .ZN(n2608) );
  NAND2_X1 U2614 ( .A1(n2634), .A2(n2635), .ZN(n2629) );
  NAND3_X1 U2615 ( .A1(n2358), .A2(n2636), .A3(n2455), .ZN(n2635) );
  NAND2_X1 U2616 ( .A1(n2604), .A2(n2603), .ZN(n2636) );
  INV_X1 U2617 ( .A(n2637), .ZN(n2634) );
  NOR2_X1 U2618 ( .A1(n2603), .A2(n2604), .ZN(n2637) );
  NOR2_X1 U2619 ( .A1(n2638), .A2(n2639), .ZN(n2604) );
  INV_X1 U2620 ( .A(n2640), .ZN(n2639) );
  NAND3_X1 U2621 ( .A1(n2641), .A2(n2642), .A3(n2455), .ZN(n2640) );
  NAND2_X1 U2622 ( .A1(n2600), .A2(n2599), .ZN(n2642) );
  NOR2_X1 U2623 ( .A1(n2599), .A2(n2600), .ZN(n2638) );
  NOR2_X1 U2624 ( .A1(n2643), .A2(n2644), .ZN(n2600) );
  INV_X1 U2625 ( .A(n2645), .ZN(n2644) );
  NAND3_X1 U2626 ( .A1(n2378), .A2(n2646), .A3(n2455), .ZN(n2645) );
  NAND2_X1 U2627 ( .A1(n2596), .A2(n2595), .ZN(n2646) );
  NOR2_X1 U2628 ( .A1(n2595), .A2(n2596), .ZN(n2643) );
  NOR2_X1 U2629 ( .A1(n2647), .A2(n2648), .ZN(n2596) );
  NOR3_X1 U2630 ( .A1(n2388), .A2(n2649), .A3(n2454), .ZN(n2648) );
  INV_X1 U2631 ( .A(n2650), .ZN(n2649) );
  NAND2_X1 U2632 ( .A1(n2591), .A2(n2589), .ZN(n2650) );
  NOR2_X1 U2633 ( .A1(n2589), .A2(n2591), .ZN(n2647) );
  NOR2_X1 U2634 ( .A1(n2651), .A2(n2652), .ZN(n2591) );
  INV_X1 U2635 ( .A(n2653), .ZN(n2652) );
  NAND3_X1 U2636 ( .A1(n2654), .A2(n2655), .A3(n2455), .ZN(n2653) );
  NAND2_X1 U2637 ( .A1(n2587), .A2(n2586), .ZN(n2655) );
  NOR2_X1 U2638 ( .A1(n2586), .A2(n2587), .ZN(n2651) );
  NOR2_X1 U2639 ( .A1(n2656), .A2(n2657), .ZN(n2587) );
  NOR3_X1 U2640 ( .A1(n2406), .A2(n2658), .A3(n2454), .ZN(n2657) );
  NOR2_X1 U2641 ( .A1(n2583), .A2(n2582), .ZN(n2658) );
  INV_X1 U2642 ( .A(n2659), .ZN(n2656) );
  NAND2_X1 U2643 ( .A1(n2582), .A2(n2583), .ZN(n2659) );
  NAND2_X1 U2644 ( .A1(n2660), .A2(n2661), .ZN(n2583) );
  NAND2_X1 U2645 ( .A1(n2579), .A2(n2662), .ZN(n2661) );
  INV_X1 U2646 ( .A(n2663), .ZN(n2662) );
  NOR2_X1 U2647 ( .A1(n2580), .A2(n2578), .ZN(n2663) );
  NOR2_X1 U2648 ( .A1(n2454), .A2(n2525), .ZN(n2579) );
  NAND2_X1 U2649 ( .A1(n2578), .A2(n2580), .ZN(n2660) );
  NAND2_X1 U2650 ( .A1(n2664), .A2(n2665), .ZN(n2580) );
  NAND2_X1 U2651 ( .A1(n2576), .A2(n2666), .ZN(n2665) );
  NAND2_X1 U2652 ( .A1(n2575), .A2(n2574), .ZN(n2666) );
  NOR2_X1 U2653 ( .A1(n2454), .A2(n2424), .ZN(n2576) );
  INV_X1 U2654 ( .A(n2667), .ZN(n2664) );
  NOR2_X1 U2655 ( .A1(n2574), .A2(n2575), .ZN(n2667) );
  NOR2_X1 U2656 ( .A1(n2668), .A2(n2669), .ZN(n2575) );
  INV_X1 U2657 ( .A(n2670), .ZN(n2669) );
  NAND2_X1 U2658 ( .A1(n2571), .A2(n2671), .ZN(n2670) );
  NAND2_X1 U2659 ( .A1(n2572), .A2(n2570), .ZN(n2671) );
  NOR2_X1 U2660 ( .A1(n2454), .A2(n2429), .ZN(n2571) );
  NOR2_X1 U2661 ( .A1(n2570), .A2(n2572), .ZN(n2668) );
  NOR2_X1 U2662 ( .A1(n2672), .A2(n2673), .ZN(n2572) );
  INV_X1 U2663 ( .A(n2674), .ZN(n2673) );
  NAND2_X1 U2664 ( .A1(n2567), .A2(n2675), .ZN(n2674) );
  NAND2_X1 U2665 ( .A1(n2568), .A2(n2566), .ZN(n2675) );
  NOR2_X1 U2666 ( .A1(n2454), .A2(n2434), .ZN(n2567) );
  NOR2_X1 U2667 ( .A1(n2566), .A2(n2568), .ZN(n2672) );
  NOR2_X1 U2668 ( .A1(n2676), .A2(n2677), .ZN(n2568) );
  INV_X1 U2669 ( .A(n2678), .ZN(n2677) );
  NAND2_X1 U2670 ( .A1(n2563), .A2(n2679), .ZN(n2678) );
  NAND2_X1 U2671 ( .A1(n2564), .A2(n2562), .ZN(n2679) );
  NOR2_X1 U2672 ( .A1(n2454), .A2(n2542), .ZN(n2563) );
  NOR2_X1 U2673 ( .A1(n2562), .A2(n2564), .ZN(n2676) );
  NOR2_X1 U2674 ( .A1(n2680), .A2(n2681), .ZN(n2564) );
  NOR2_X1 U2675 ( .A1(n2557), .A2(n2682), .ZN(n2681) );
  NOR2_X1 U2676 ( .A1(n2560), .A2(n2559), .ZN(n2682) );
  NAND2_X1 U2677 ( .A1(n2455), .A2(n2447), .ZN(n2557) );
  INV_X1 U2678 ( .A(n2454), .ZN(n2455) );
  INV_X1 U2679 ( .A(n2683), .ZN(n2680) );
  NAND2_X1 U2680 ( .A1(n2559), .A2(n2560), .ZN(n2683) );
  NAND2_X1 U2681 ( .A1(n2684), .A2(n2685), .ZN(n2560) );
  NAND2_X1 U2682 ( .A1(n2552), .A2(n2686), .ZN(n2685) );
  NAND2_X1 U2683 ( .A1(n2202), .A2(n2687), .ZN(n2686) );
  NAND2_X1 U2684 ( .A1(n2688), .A2(n2205), .ZN(n2687) );
  NAND2_X1 U2685 ( .A1(n2689), .A2(n2690), .ZN(n2684) );
  NAND2_X1 U2686 ( .A1(n2208), .A2(n2691), .ZN(n2690) );
  NAND2_X1 U2687 ( .A1(n2210), .A2(n2551), .ZN(n2691) );
  NOR3_X1 U2688 ( .A1(n2551), .A2(n2449), .A3(n2454), .ZN(n2559) );
  XOR2_X1 U2689 ( .A(d_13_), .B(c_13_), .Z(n2693) );
  XNOR2_X1 U2690 ( .A(n2694), .B(n2695), .ZN(n2562) );
  XNOR2_X1 U2691 ( .A(n2696), .B(n2697), .ZN(n2695) );
  XOR2_X1 U2692 ( .A(n2698), .B(n2699), .Z(n2566) );
  XNOR2_X1 U2693 ( .A(n2700), .B(n2701), .ZN(n2698) );
  XOR2_X1 U2694 ( .A(n2702), .B(n2703), .Z(n2570) );
  XNOR2_X1 U2695 ( .A(n2704), .B(n2705), .ZN(n2702) );
  XOR2_X1 U2696 ( .A(n2706), .B(n2707), .Z(n2574) );
  XNOR2_X1 U2697 ( .A(n2708), .B(n2709), .ZN(n2706) );
  XNOR2_X1 U2698 ( .A(n2710), .B(n2711), .ZN(n2578) );
  XNOR2_X1 U2699 ( .A(n2712), .B(n2713), .ZN(n2710) );
  XNOR2_X1 U2700 ( .A(n2714), .B(n2715), .ZN(n2582) );
  XNOR2_X1 U2701 ( .A(n2716), .B(n2717), .ZN(n2714) );
  XOR2_X1 U2702 ( .A(n2718), .B(n2719), .Z(n2586) );
  XNOR2_X1 U2703 ( .A(n2720), .B(n2721), .ZN(n2718) );
  XOR2_X1 U2704 ( .A(n2722), .B(n2723), .Z(n2589) );
  XNOR2_X1 U2705 ( .A(n2724), .B(n2725), .ZN(n2722) );
  XNOR2_X1 U2706 ( .A(n2726), .B(n2727), .ZN(n2595) );
  XNOR2_X1 U2707 ( .A(n2728), .B(n2729), .ZN(n2726) );
  XOR2_X1 U2708 ( .A(n2730), .B(n2731), .Z(n2599) );
  XNOR2_X1 U2709 ( .A(n2732), .B(n2733), .ZN(n2730) );
  XNOR2_X1 U2710 ( .A(n2734), .B(n2735), .ZN(n2603) );
  XOR2_X1 U2711 ( .A(n2736), .B(n2737), .Z(n2735) );
  NOR2_X1 U2712 ( .A1(n2369), .A2(n2551), .ZN(n2737) );
  XOR2_X1 U2713 ( .A(n2483), .B(n2482), .Z(n2617) );
  XOR2_X1 U2714 ( .A(n2738), .B(n2739), .Z(n2482) );
  NOR2_X1 U2715 ( .A1(n2345), .A2(n2551), .ZN(n2739) );
  XOR2_X1 U2716 ( .A(n2300), .B(n2299), .Z(n2291) );
  NAND3_X1 U2717 ( .A1(n2299), .A2(n2300), .A3(n2298), .ZN(n2294) );
  NOR2_X1 U2718 ( .A1(n2740), .A2(n2741), .ZN(n2298) );
  NOR2_X1 U2719 ( .A1(n2742), .A2(n2743), .ZN(n2741) );
  INV_X1 U2720 ( .A(n2334), .ZN(n2740) );
  NAND2_X1 U2721 ( .A1(n2744), .A2(n2745), .ZN(n2300) );
  INV_X1 U2722 ( .A(n2746), .ZN(n2745) );
  NOR3_X1 U2723 ( .A1(n2345), .A2(n2747), .A3(n2551), .ZN(n2746) );
  NOR2_X1 U2724 ( .A1(n2738), .A2(n2483), .ZN(n2747) );
  NAND2_X1 U2725 ( .A1(n2483), .A2(n2738), .ZN(n2744) );
  NAND2_X1 U2726 ( .A1(n2748), .A2(n2749), .ZN(n2738) );
  NAND2_X1 U2727 ( .A1(n2625), .A2(n2750), .ZN(n2749) );
  INV_X1 U2728 ( .A(n2751), .ZN(n2750) );
  NOR2_X1 U2729 ( .A1(n2624), .A2(n2623), .ZN(n2751) );
  NOR2_X1 U2730 ( .A1(n2551), .A2(n2354), .ZN(n2625) );
  NAND2_X1 U2731 ( .A1(n2623), .A2(n2624), .ZN(n2748) );
  NAND2_X1 U2732 ( .A1(n2752), .A2(n2753), .ZN(n2624) );
  NAND3_X1 U2733 ( .A1(n2358), .A2(n2754), .A3(n2552), .ZN(n2753) );
  NAND2_X1 U2734 ( .A1(n2632), .A2(n2630), .ZN(n2754) );
  INV_X1 U2735 ( .A(n2755), .ZN(n2752) );
  NOR2_X1 U2736 ( .A1(n2630), .A2(n2632), .ZN(n2755) );
  NOR2_X1 U2737 ( .A1(n2756), .A2(n2757), .ZN(n2632) );
  INV_X1 U2738 ( .A(n2758), .ZN(n2757) );
  NAND3_X1 U2739 ( .A1(n2641), .A2(n2759), .A3(n2552), .ZN(n2758) );
  NAND2_X1 U2740 ( .A1(n2736), .A2(n2734), .ZN(n2759) );
  NOR2_X1 U2741 ( .A1(n2734), .A2(n2736), .ZN(n2756) );
  NOR2_X1 U2742 ( .A1(n2760), .A2(n2761), .ZN(n2736) );
  INV_X1 U2743 ( .A(n2762), .ZN(n2761) );
  NAND2_X1 U2744 ( .A1(n2732), .A2(n2763), .ZN(n2762) );
  NAND2_X1 U2745 ( .A1(n2733), .A2(n2731), .ZN(n2763) );
  NOR2_X1 U2746 ( .A1(n2551), .A2(n2508), .ZN(n2732) );
  NOR2_X1 U2747 ( .A1(n2731), .A2(n2733), .ZN(n2760) );
  INV_X1 U2748 ( .A(n2764), .ZN(n2733) );
  NAND2_X1 U2749 ( .A1(n2765), .A2(n2766), .ZN(n2764) );
  NAND2_X1 U2750 ( .A1(n2729), .A2(n2767), .ZN(n2766) );
  NAND2_X1 U2751 ( .A1(n2728), .A2(n2768), .ZN(n2767) );
  INV_X1 U2752 ( .A(n2727), .ZN(n2768) );
  NOR2_X1 U2753 ( .A1(n2551), .A2(n2388), .ZN(n2729) );
  NAND2_X1 U2754 ( .A1(n2727), .A2(n2769), .ZN(n2765) );
  INV_X1 U2755 ( .A(n2728), .ZN(n2769) );
  NOR2_X1 U2756 ( .A1(n2770), .A2(n2771), .ZN(n2728) );
  INV_X1 U2757 ( .A(n2772), .ZN(n2771) );
  NAND2_X1 U2758 ( .A1(n2725), .A2(n2773), .ZN(n2772) );
  NAND2_X1 U2759 ( .A1(n2724), .A2(n2723), .ZN(n2773) );
  NOR2_X1 U2760 ( .A1(n2551), .A2(n2396), .ZN(n2725) );
  NOR2_X1 U2761 ( .A1(n2723), .A2(n2724), .ZN(n2770) );
  NOR2_X1 U2762 ( .A1(n2774), .A2(n2775), .ZN(n2724) );
  INV_X1 U2763 ( .A(n2776), .ZN(n2775) );
  NAND2_X1 U2764 ( .A1(n2720), .A2(n2777), .ZN(n2776) );
  NAND2_X1 U2765 ( .A1(n2721), .A2(n2719), .ZN(n2777) );
  NOR2_X1 U2766 ( .A1(n2551), .A2(n2406), .ZN(n2720) );
  NOR2_X1 U2767 ( .A1(n2719), .A2(n2721), .ZN(n2774) );
  NOR2_X1 U2768 ( .A1(n2778), .A2(n2779), .ZN(n2721) );
  INV_X1 U2769 ( .A(n2780), .ZN(n2779) );
  NAND2_X1 U2770 ( .A1(n2717), .A2(n2781), .ZN(n2780) );
  NAND2_X1 U2771 ( .A1(n2716), .A2(n2715), .ZN(n2781) );
  NOR2_X1 U2772 ( .A1(n2551), .A2(n2525), .ZN(n2717) );
  NOR2_X1 U2773 ( .A1(n2715), .A2(n2716), .ZN(n2778) );
  NOR2_X1 U2774 ( .A1(n2782), .A2(n2783), .ZN(n2716) );
  INV_X1 U2775 ( .A(n2784), .ZN(n2783) );
  NAND2_X1 U2776 ( .A1(n2712), .A2(n2785), .ZN(n2784) );
  NAND2_X1 U2777 ( .A1(n2713), .A2(n2711), .ZN(n2785) );
  NOR2_X1 U2778 ( .A1(n2551), .A2(n2424), .ZN(n2712) );
  NOR2_X1 U2779 ( .A1(n2711), .A2(n2713), .ZN(n2782) );
  NOR2_X1 U2780 ( .A1(n2786), .A2(n2787), .ZN(n2713) );
  INV_X1 U2781 ( .A(n2788), .ZN(n2787) );
  NAND2_X1 U2782 ( .A1(n2708), .A2(n2789), .ZN(n2788) );
  NAND2_X1 U2783 ( .A1(n2709), .A2(n2707), .ZN(n2789) );
  NOR2_X1 U2784 ( .A1(n2551), .A2(n2429), .ZN(n2708) );
  NOR2_X1 U2785 ( .A1(n2707), .A2(n2709), .ZN(n2786) );
  NOR2_X1 U2786 ( .A1(n2790), .A2(n2791), .ZN(n2709) );
  INV_X1 U2787 ( .A(n2792), .ZN(n2791) );
  NAND2_X1 U2788 ( .A1(n2704), .A2(n2793), .ZN(n2792) );
  NAND2_X1 U2789 ( .A1(n2705), .A2(n2703), .ZN(n2793) );
  NOR2_X1 U2790 ( .A1(n2551), .A2(n2434), .ZN(n2704) );
  NOR2_X1 U2791 ( .A1(n2703), .A2(n2705), .ZN(n2790) );
  NOR2_X1 U2792 ( .A1(n2794), .A2(n2795), .ZN(n2705) );
  INV_X1 U2793 ( .A(n2796), .ZN(n2795) );
  NAND2_X1 U2794 ( .A1(n2700), .A2(n2797), .ZN(n2796) );
  NAND2_X1 U2795 ( .A1(n2701), .A2(n2699), .ZN(n2797) );
  NOR2_X1 U2796 ( .A1(n2551), .A2(n2542), .ZN(n2700) );
  NOR2_X1 U2797 ( .A1(n2699), .A2(n2701), .ZN(n2794) );
  NOR2_X1 U2798 ( .A1(n2798), .A2(n2799), .ZN(n2701) );
  NOR2_X1 U2799 ( .A1(n2694), .A2(n2800), .ZN(n2799) );
  NOR2_X1 U2800 ( .A1(n2697), .A2(n2696), .ZN(n2800) );
  NAND2_X1 U2801 ( .A1(n2552), .A2(n2447), .ZN(n2694) );
  INV_X1 U2802 ( .A(n2551), .ZN(n2552) );
  INV_X1 U2803 ( .A(n2801), .ZN(n2798) );
  NAND2_X1 U2804 ( .A1(n2696), .A2(n2697), .ZN(n2801) );
  NAND2_X1 U2805 ( .A1(n2802), .A2(n2803), .ZN(n2697) );
  NAND2_X1 U2806 ( .A1(n2689), .A2(n2804), .ZN(n2803) );
  NAND2_X1 U2807 ( .A1(n2202), .A2(n2805), .ZN(n2804) );
  NAND2_X1 U2808 ( .A1(n2806), .A2(n2205), .ZN(n2805) );
  NAND2_X1 U2809 ( .A1(n2807), .A2(n2808), .ZN(n2802) );
  NAND2_X1 U2810 ( .A1(n2208), .A2(n2809), .ZN(n2808) );
  NAND2_X1 U2811 ( .A1(n2210), .A2(n2688), .ZN(n2809) );
  NOR3_X1 U2812 ( .A1(n2688), .A2(n2449), .A3(n2551), .ZN(n2696) );
  XOR2_X1 U2813 ( .A(d_12_), .B(c_12_), .Z(n2811) );
  XNOR2_X1 U2814 ( .A(n2812), .B(n2813), .ZN(n2699) );
  XNOR2_X1 U2815 ( .A(n2814), .B(n2815), .ZN(n2813) );
  XOR2_X1 U2816 ( .A(n2816), .B(n2817), .Z(n2703) );
  XNOR2_X1 U2817 ( .A(n2818), .B(n2819), .ZN(n2816) );
  XOR2_X1 U2818 ( .A(n2820), .B(n2821), .Z(n2707) );
  XNOR2_X1 U2819 ( .A(n2822), .B(n2823), .ZN(n2820) );
  XOR2_X1 U2820 ( .A(n2824), .B(n2825), .Z(n2711) );
  XNOR2_X1 U2821 ( .A(n2826), .B(n2827), .ZN(n2824) );
  XOR2_X1 U2822 ( .A(n2828), .B(n2829), .Z(n2715) );
  XNOR2_X1 U2823 ( .A(n2830), .B(n2831), .ZN(n2828) );
  XNOR2_X1 U2824 ( .A(n2832), .B(n2833), .ZN(n2719) );
  XOR2_X1 U2825 ( .A(n2834), .B(n2835), .Z(n2832) );
  XOR2_X1 U2826 ( .A(n2836), .B(n2837), .Z(n2723) );
  XOR2_X1 U2827 ( .A(n2838), .B(n2839), .Z(n2837) );
  NAND2_X1 U2828 ( .A1(n2689), .A2(n2840), .ZN(n2839) );
  XOR2_X1 U2829 ( .A(n2841), .B(n2842), .Z(n2727) );
  XOR2_X1 U2830 ( .A(n2843), .B(n2844), .Z(n2841) );
  NOR2_X1 U2831 ( .A1(n2396), .A2(n2688), .ZN(n2844) );
  XOR2_X1 U2832 ( .A(n2845), .B(n2846), .Z(n2731) );
  XNOR2_X1 U2833 ( .A(n2847), .B(n2848), .ZN(n2845) );
  NOR2_X1 U2834 ( .A1(n2388), .A2(n2688), .ZN(n2848) );
  XOR2_X1 U2835 ( .A(n2849), .B(n2850), .Z(n2734) );
  XNOR2_X1 U2836 ( .A(n2851), .B(n2852), .ZN(n2849) );
  NOR2_X1 U2837 ( .A1(n2508), .A2(n2688), .ZN(n2852) );
  XOR2_X1 U2838 ( .A(n2853), .B(n2854), .Z(n2630) );
  NAND2_X1 U2839 ( .A1(n2855), .A2(n2856), .ZN(n2853) );
  XNOR2_X1 U2840 ( .A(n2857), .B(n2858), .ZN(n2623) );
  XOR2_X1 U2841 ( .A(n2859), .B(n2860), .Z(n2858) );
  NAND2_X1 U2842 ( .A1(n2689), .A2(n2358), .ZN(n2860) );
  XNOR2_X1 U2843 ( .A(n2861), .B(n2862), .ZN(n2483) );
  XOR2_X1 U2844 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND2_X1 U2845 ( .A1(n2689), .A2(n2492), .ZN(n2864) );
  XNOR2_X1 U2846 ( .A(n2865), .B(n2866), .ZN(n2299) );
  NAND2_X1 U2847 ( .A1(n2867), .A2(n2868), .ZN(n2865) );
  NAND2_X1 U2848 ( .A1(n2743), .A2(n2742), .ZN(n2334) );
  NAND2_X1 U2849 ( .A1(n2867), .A2(n2869), .ZN(n2742) );
  NAND2_X1 U2850 ( .A1(n2866), .A2(n2868), .ZN(n2869) );
  NAND2_X1 U2851 ( .A1(n2870), .A2(n2871), .ZN(n2868) );
  NAND2_X1 U2852 ( .A1(n2689), .A2(n2303), .ZN(n2871) );
  INV_X1 U2853 ( .A(n2872), .ZN(n2870) );
  XOR2_X1 U2854 ( .A(n2873), .B(n2874), .Z(n2866) );
  XOR2_X1 U2855 ( .A(n2875), .B(n2876), .Z(n2873) );
  NAND2_X1 U2856 ( .A1(n2303), .A2(n2872), .ZN(n2867) );
  NAND2_X1 U2857 ( .A1(n2877), .A2(n2878), .ZN(n2872) );
  INV_X1 U2858 ( .A(n2879), .ZN(n2878) );
  NOR3_X1 U2859 ( .A1(n2354), .A2(n2880), .A3(n2688), .ZN(n2879) );
  NOR2_X1 U2860 ( .A1(n2863), .A2(n2861), .ZN(n2880) );
  NAND2_X1 U2861 ( .A1(n2861), .A2(n2863), .ZN(n2877) );
  NAND2_X1 U2862 ( .A1(n2881), .A2(n2882), .ZN(n2863) );
  NAND3_X1 U2863 ( .A1(n2358), .A2(n2883), .A3(n2689), .ZN(n2882) );
  INV_X1 U2864 ( .A(n2884), .ZN(n2883) );
  NOR2_X1 U2865 ( .A1(n2859), .A2(n2857), .ZN(n2884) );
  NAND2_X1 U2866 ( .A1(n2857), .A2(n2859), .ZN(n2881) );
  NAND2_X1 U2867 ( .A1(n2855), .A2(n2885), .ZN(n2859) );
  NAND2_X1 U2868 ( .A1(n2854), .A2(n2856), .ZN(n2885) );
  NAND2_X1 U2869 ( .A1(n2886), .A2(n2887), .ZN(n2856) );
  NAND2_X1 U2870 ( .A1(n2689), .A2(n2641), .ZN(n2887) );
  INV_X1 U2871 ( .A(n2888), .ZN(n2886) );
  XNOR2_X1 U2872 ( .A(n2889), .B(n2890), .ZN(n2854) );
  XNOR2_X1 U2873 ( .A(n2891), .B(n2892), .ZN(n2889) );
  NOR2_X1 U2874 ( .A1(n2508), .A2(n2806), .ZN(n2892) );
  NAND2_X1 U2875 ( .A1(n2641), .A2(n2888), .ZN(n2855) );
  NAND2_X1 U2876 ( .A1(n2893), .A2(n2894), .ZN(n2888) );
  NAND3_X1 U2877 ( .A1(n2378), .A2(n2895), .A3(n2689), .ZN(n2894) );
  NAND2_X1 U2878 ( .A1(n2851), .A2(n2850), .ZN(n2895) );
  INV_X1 U2879 ( .A(n2896), .ZN(n2893) );
  NOR2_X1 U2880 ( .A1(n2850), .A2(n2851), .ZN(n2896) );
  NOR2_X1 U2881 ( .A1(n2897), .A2(n2898), .ZN(n2851) );
  INV_X1 U2882 ( .A(n2899), .ZN(n2898) );
  NAND3_X1 U2883 ( .A1(n2593), .A2(n2900), .A3(n2689), .ZN(n2899) );
  NAND2_X1 U2884 ( .A1(n2847), .A2(n2846), .ZN(n2900) );
  NOR2_X1 U2885 ( .A1(n2846), .A2(n2847), .ZN(n2897) );
  NOR2_X1 U2886 ( .A1(n2901), .A2(n2902), .ZN(n2847) );
  NOR3_X1 U2887 ( .A1(n2396), .A2(n2903), .A3(n2688), .ZN(n2902) );
  NOR2_X1 U2888 ( .A1(n2843), .A2(n2842), .ZN(n2903) );
  INV_X1 U2889 ( .A(n2904), .ZN(n2901) );
  NAND2_X1 U2890 ( .A1(n2842), .A2(n2843), .ZN(n2904) );
  NAND2_X1 U2891 ( .A1(n2905), .A2(n2906), .ZN(n2843) );
  NAND3_X1 U2892 ( .A1(n2840), .A2(n2907), .A3(n2689), .ZN(n2906) );
  INV_X1 U2893 ( .A(n2908), .ZN(n2907) );
  NOR2_X1 U2894 ( .A1(n2838), .A2(n2836), .ZN(n2908) );
  NAND2_X1 U2895 ( .A1(n2836), .A2(n2838), .ZN(n2905) );
  NAND2_X1 U2896 ( .A1(n2909), .A2(n2910), .ZN(n2838) );
  NAND2_X1 U2897 ( .A1(n2834), .A2(n2911), .ZN(n2910) );
  INV_X1 U2898 ( .A(n2912), .ZN(n2911) );
  NOR2_X1 U2899 ( .A1(n2835), .A2(n2833), .ZN(n2912) );
  NOR2_X1 U2900 ( .A1(n2688), .A2(n2525), .ZN(n2834) );
  NAND2_X1 U2901 ( .A1(n2833), .A2(n2835), .ZN(n2909) );
  NAND2_X1 U2902 ( .A1(n2913), .A2(n2914), .ZN(n2835) );
  NAND2_X1 U2903 ( .A1(n2831), .A2(n2915), .ZN(n2914) );
  NAND2_X1 U2904 ( .A1(n2830), .A2(n2829), .ZN(n2915) );
  NOR2_X1 U2905 ( .A1(n2688), .A2(n2424), .ZN(n2831) );
  INV_X1 U2906 ( .A(n2916), .ZN(n2913) );
  NOR2_X1 U2907 ( .A1(n2829), .A2(n2830), .ZN(n2916) );
  NOR2_X1 U2908 ( .A1(n2917), .A2(n2918), .ZN(n2830) );
  INV_X1 U2909 ( .A(n2919), .ZN(n2918) );
  NAND2_X1 U2910 ( .A1(n2826), .A2(n2920), .ZN(n2919) );
  NAND2_X1 U2911 ( .A1(n2827), .A2(n2825), .ZN(n2920) );
  NOR2_X1 U2912 ( .A1(n2688), .A2(n2429), .ZN(n2826) );
  NOR2_X1 U2913 ( .A1(n2825), .A2(n2827), .ZN(n2917) );
  NOR2_X1 U2914 ( .A1(n2921), .A2(n2922), .ZN(n2827) );
  INV_X1 U2915 ( .A(n2923), .ZN(n2922) );
  NAND2_X1 U2916 ( .A1(n2822), .A2(n2924), .ZN(n2923) );
  NAND2_X1 U2917 ( .A1(n2823), .A2(n2821), .ZN(n2924) );
  NOR2_X1 U2918 ( .A1(n2688), .A2(n2434), .ZN(n2822) );
  NOR2_X1 U2919 ( .A1(n2821), .A2(n2823), .ZN(n2921) );
  NOR2_X1 U2920 ( .A1(n2925), .A2(n2926), .ZN(n2823) );
  INV_X1 U2921 ( .A(n2927), .ZN(n2926) );
  NAND2_X1 U2922 ( .A1(n2818), .A2(n2928), .ZN(n2927) );
  NAND2_X1 U2923 ( .A1(n2819), .A2(n2817), .ZN(n2928) );
  NOR2_X1 U2924 ( .A1(n2688), .A2(n2542), .ZN(n2818) );
  NOR2_X1 U2925 ( .A1(n2817), .A2(n2819), .ZN(n2925) );
  NOR2_X1 U2926 ( .A1(n2929), .A2(n2930), .ZN(n2819) );
  NOR2_X1 U2927 ( .A1(n2812), .A2(n2931), .ZN(n2930) );
  NOR2_X1 U2928 ( .A1(n2815), .A2(n2814), .ZN(n2931) );
  NAND2_X1 U2929 ( .A1(n2689), .A2(n2447), .ZN(n2812) );
  INV_X1 U2930 ( .A(n2688), .ZN(n2689) );
  INV_X1 U2931 ( .A(n2932), .ZN(n2929) );
  NAND2_X1 U2932 ( .A1(n2814), .A2(n2815), .ZN(n2932) );
  NAND2_X1 U2933 ( .A1(n2933), .A2(n2934), .ZN(n2815) );
  NAND2_X1 U2934 ( .A1(n2807), .A2(n2935), .ZN(n2934) );
  NAND2_X1 U2935 ( .A1(n2202), .A2(n2936), .ZN(n2935) );
  NAND2_X1 U2936 ( .A1(n2205), .A2(n2937), .ZN(n2936) );
  NAND2_X1 U2937 ( .A1(n2938), .A2(n2939), .ZN(n2933) );
  NAND2_X1 U2938 ( .A1(n2208), .A2(n2940), .ZN(n2939) );
  NAND2_X1 U2939 ( .A1(n2210), .A2(n2806), .ZN(n2940) );
  NOR3_X1 U2940 ( .A1(n2806), .A2(n2449), .A3(n2688), .ZN(n2814) );
  XOR2_X1 U2941 ( .A(d_11_), .B(c_11_), .Z(n2942) );
  XNOR2_X1 U2942 ( .A(n2943), .B(n2944), .ZN(n2817) );
  XNOR2_X1 U2943 ( .A(n2945), .B(n2946), .ZN(n2944) );
  XOR2_X1 U2944 ( .A(n2947), .B(n2948), .Z(n2821) );
  XNOR2_X1 U2945 ( .A(n2949), .B(n2950), .ZN(n2947) );
  XOR2_X1 U2946 ( .A(n2951), .B(n2952), .Z(n2825) );
  XNOR2_X1 U2947 ( .A(n2953), .B(n2954), .ZN(n2951) );
  XOR2_X1 U2948 ( .A(n2955), .B(n2956), .Z(n2829) );
  XNOR2_X1 U2949 ( .A(n2957), .B(n2958), .ZN(n2955) );
  XNOR2_X1 U2950 ( .A(n2959), .B(n2960), .ZN(n2833) );
  XNOR2_X1 U2951 ( .A(n2961), .B(n2962), .ZN(n2959) );
  XNOR2_X1 U2952 ( .A(n2963), .B(n2964), .ZN(n2836) );
  XNOR2_X1 U2953 ( .A(n2965), .B(n2966), .ZN(n2963) );
  XNOR2_X1 U2954 ( .A(n2967), .B(n2968), .ZN(n2842) );
  XNOR2_X1 U2955 ( .A(n2969), .B(n2970), .ZN(n2967) );
  XOR2_X1 U2956 ( .A(n2971), .B(n2972), .Z(n2846) );
  XNOR2_X1 U2957 ( .A(n2973), .B(n2974), .ZN(n2971) );
  XNOR2_X1 U2958 ( .A(n2975), .B(n2976), .ZN(n2850) );
  XOR2_X1 U2959 ( .A(n2977), .B(n2978), .Z(n2976) );
  NOR2_X1 U2960 ( .A1(n2388), .A2(n2806), .ZN(n2978) );
  XOR2_X1 U2961 ( .A(n2979), .B(n2980), .Z(n2857) );
  XOR2_X1 U2962 ( .A(n2981), .B(n2982), .Z(n2979) );
  NOR2_X1 U2963 ( .A1(n2369), .A2(n2806), .ZN(n2982) );
  XNOR2_X1 U2964 ( .A(n2983), .B(n2984), .ZN(n2861) );
  NAND2_X1 U2965 ( .A1(n2985), .A2(n2986), .ZN(n2983) );
  XOR2_X1 U2966 ( .A(n2987), .B(n2988), .Z(n2743) );
  XOR2_X1 U2967 ( .A(n2989), .B(n2990), .Z(n2987) );
  NOR2_X1 U2968 ( .A1(n2345), .A2(n2806), .ZN(n2990) );
  XOR2_X1 U2969 ( .A(n2165), .B(n2164), .Z(n2158) );
  NAND3_X1 U2970 ( .A1(n2164), .A2(n2165), .A3(n2333), .ZN(n2160) );
  INV_X1 U2971 ( .A(n2163), .ZN(n2333) );
  NAND2_X1 U2972 ( .A1(n2991), .A2(n2331), .ZN(n2163) );
  NAND2_X1 U2973 ( .A1(n2992), .A2(n2993), .ZN(n2991) );
  INV_X1 U2974 ( .A(n2994), .ZN(n2993) );
  XNOR2_X1 U2975 ( .A(n2995), .B(n2996), .ZN(n2992) );
  INV_X1 U2976 ( .A(n2997), .ZN(n2996) );
  NAND2_X1 U2977 ( .A1(n2998), .A2(n2999), .ZN(n2165) );
  INV_X1 U2978 ( .A(n3000), .ZN(n2999) );
  NOR3_X1 U2979 ( .A1(n2345), .A2(n3001), .A3(n2806), .ZN(n3000) );
  NOR2_X1 U2980 ( .A1(n2989), .A2(n2988), .ZN(n3001) );
  NAND2_X1 U2981 ( .A1(n2988), .A2(n2989), .ZN(n2998) );
  NAND2_X1 U2982 ( .A1(n3002), .A2(n3003), .ZN(n2989) );
  NAND2_X1 U2983 ( .A1(n2876), .A2(n3004), .ZN(n3003) );
  INV_X1 U2984 ( .A(n3005), .ZN(n3004) );
  NOR2_X1 U2985 ( .A1(n2875), .A2(n2874), .ZN(n3005) );
  NOR2_X1 U2986 ( .A1(n2806), .A2(n2354), .ZN(n2876) );
  NAND2_X1 U2987 ( .A1(n2874), .A2(n2875), .ZN(n3002) );
  NAND2_X1 U2988 ( .A1(n2985), .A2(n3006), .ZN(n2875) );
  NAND2_X1 U2989 ( .A1(n2984), .A2(n2986), .ZN(n3006) );
  NAND2_X1 U2990 ( .A1(n3007), .A2(n3008), .ZN(n2986) );
  NAND2_X1 U2991 ( .A1(n2807), .A2(n2358), .ZN(n3008) );
  XNOR2_X1 U2992 ( .A(n3009), .B(n3010), .ZN(n2984) );
  XNOR2_X1 U2993 ( .A(n3011), .B(n3012), .ZN(n3009) );
  NOR2_X1 U2994 ( .A1(n2937), .A2(n2369), .ZN(n3012) );
  INV_X1 U2995 ( .A(n3013), .ZN(n2985) );
  NOR2_X1 U2996 ( .A1(n2497), .A2(n3007), .ZN(n3013) );
  NOR2_X1 U2997 ( .A1(n3014), .A2(n3015), .ZN(n3007) );
  NOR3_X1 U2998 ( .A1(n2369), .A2(n3016), .A3(n2806), .ZN(n3015) );
  NOR2_X1 U2999 ( .A1(n2981), .A2(n2980), .ZN(n3016) );
  INV_X1 U3000 ( .A(n3017), .ZN(n3014) );
  NAND2_X1 U3001 ( .A1(n2980), .A2(n2981), .ZN(n3017) );
  NAND2_X1 U3002 ( .A1(n3018), .A2(n3019), .ZN(n2981) );
  NAND3_X1 U3003 ( .A1(n2378), .A2(n3020), .A3(n2807), .ZN(n3019) );
  NAND2_X1 U3004 ( .A1(n2891), .A2(n2890), .ZN(n3020) );
  INV_X1 U3005 ( .A(n3021), .ZN(n3018) );
  NOR2_X1 U3006 ( .A1(n2890), .A2(n2891), .ZN(n3021) );
  NOR2_X1 U3007 ( .A1(n3022), .A2(n3023), .ZN(n2891) );
  NOR3_X1 U3008 ( .A1(n2388), .A2(n3024), .A3(n2806), .ZN(n3023) );
  INV_X1 U3009 ( .A(n3025), .ZN(n3024) );
  NAND2_X1 U3010 ( .A1(n2977), .A2(n2975), .ZN(n3025) );
  NOR2_X1 U3011 ( .A1(n2975), .A2(n2977), .ZN(n3022) );
  NOR2_X1 U3012 ( .A1(n3026), .A2(n3027), .ZN(n2977) );
  INV_X1 U3013 ( .A(n3028), .ZN(n3027) );
  NAND2_X1 U3014 ( .A1(n2973), .A2(n3029), .ZN(n3028) );
  NAND2_X1 U3015 ( .A1(n2974), .A2(n2972), .ZN(n3029) );
  NOR2_X1 U3016 ( .A1(n2806), .A2(n2396), .ZN(n2973) );
  NOR2_X1 U3017 ( .A1(n2972), .A2(n2974), .ZN(n3026) );
  NOR2_X1 U3018 ( .A1(n3030), .A2(n3031), .ZN(n2974) );
  INV_X1 U3019 ( .A(n3032), .ZN(n3031) );
  NAND2_X1 U3020 ( .A1(n2970), .A2(n3033), .ZN(n3032) );
  NAND2_X1 U3021 ( .A1(n2969), .A2(n2968), .ZN(n3033) );
  NOR2_X1 U3022 ( .A1(n2806), .A2(n2406), .ZN(n2970) );
  NOR2_X1 U3023 ( .A1(n2968), .A2(n2969), .ZN(n3030) );
  NOR2_X1 U3024 ( .A1(n3034), .A2(n3035), .ZN(n2969) );
  INV_X1 U3025 ( .A(n3036), .ZN(n3035) );
  NAND2_X1 U3026 ( .A1(n2966), .A2(n3037), .ZN(n3036) );
  NAND2_X1 U3027 ( .A1(n2965), .A2(n2964), .ZN(n3037) );
  NOR2_X1 U3028 ( .A1(n2806), .A2(n2525), .ZN(n2966) );
  NOR2_X1 U3029 ( .A1(n2964), .A2(n2965), .ZN(n3034) );
  NOR2_X1 U3030 ( .A1(n3038), .A2(n3039), .ZN(n2965) );
  INV_X1 U3031 ( .A(n3040), .ZN(n3039) );
  NAND2_X1 U3032 ( .A1(n2961), .A2(n3041), .ZN(n3040) );
  NAND2_X1 U3033 ( .A1(n2962), .A2(n2960), .ZN(n3041) );
  NOR2_X1 U3034 ( .A1(n2806), .A2(n2424), .ZN(n2961) );
  NOR2_X1 U3035 ( .A1(n2960), .A2(n2962), .ZN(n3038) );
  NOR2_X1 U3036 ( .A1(n3042), .A2(n3043), .ZN(n2962) );
  INV_X1 U3037 ( .A(n3044), .ZN(n3043) );
  NAND2_X1 U3038 ( .A1(n2957), .A2(n3045), .ZN(n3044) );
  NAND2_X1 U3039 ( .A1(n2958), .A2(n2956), .ZN(n3045) );
  NOR2_X1 U3040 ( .A1(n2806), .A2(n2429), .ZN(n2957) );
  NOR2_X1 U3041 ( .A1(n2956), .A2(n2958), .ZN(n3042) );
  NOR2_X1 U3042 ( .A1(n3046), .A2(n3047), .ZN(n2958) );
  INV_X1 U3043 ( .A(n3048), .ZN(n3047) );
  NAND2_X1 U3044 ( .A1(n2953), .A2(n3049), .ZN(n3048) );
  NAND2_X1 U3045 ( .A1(n2954), .A2(n2952), .ZN(n3049) );
  NOR2_X1 U3046 ( .A1(n2806), .A2(n2434), .ZN(n2953) );
  NOR2_X1 U3047 ( .A1(n2952), .A2(n2954), .ZN(n3046) );
  NOR2_X1 U3048 ( .A1(n3050), .A2(n3051), .ZN(n2954) );
  INV_X1 U3049 ( .A(n3052), .ZN(n3051) );
  NAND2_X1 U3050 ( .A1(n2949), .A2(n3053), .ZN(n3052) );
  NAND2_X1 U3051 ( .A1(n2950), .A2(n2948), .ZN(n3053) );
  NOR2_X1 U3052 ( .A1(n2806), .A2(n2542), .ZN(n2949) );
  NOR2_X1 U3053 ( .A1(n2948), .A2(n2950), .ZN(n3050) );
  NOR2_X1 U3054 ( .A1(n3054), .A2(n3055), .ZN(n2950) );
  NOR2_X1 U3055 ( .A1(n2943), .A2(n3056), .ZN(n3055) );
  NOR2_X1 U3056 ( .A1(n2946), .A2(n2945), .ZN(n3056) );
  NAND2_X1 U3057 ( .A1(n2807), .A2(n2447), .ZN(n2943) );
  INV_X1 U3058 ( .A(n2806), .ZN(n2807) );
  INV_X1 U3059 ( .A(n3057), .ZN(n3054) );
  NAND2_X1 U3060 ( .A1(n2945), .A2(n2946), .ZN(n3057) );
  NAND2_X1 U3061 ( .A1(n3058), .A2(n3059), .ZN(n2946) );
  NAND2_X1 U3062 ( .A1(n2938), .A2(n3060), .ZN(n3059) );
  NAND2_X1 U3063 ( .A1(n2202), .A2(n3061), .ZN(n3060) );
  NAND2_X1 U3064 ( .A1(n3062), .A2(n2205), .ZN(n3061) );
  NAND2_X1 U3065 ( .A1(n3063), .A2(n3064), .ZN(n3058) );
  NAND2_X1 U3066 ( .A1(n2208), .A2(n3065), .ZN(n3064) );
  NAND2_X1 U3067 ( .A1(n2210), .A2(n2937), .ZN(n3065) );
  NOR3_X1 U3068 ( .A1(n2937), .A2(n2449), .A3(n2806), .ZN(n2945) );
  XOR2_X1 U3069 ( .A(d_10_), .B(c_10_), .Z(n3067) );
  XNOR2_X1 U3070 ( .A(n3068), .B(n3069), .ZN(n2948) );
  XNOR2_X1 U3071 ( .A(n3070), .B(n3071), .ZN(n3069) );
  XOR2_X1 U3072 ( .A(n3072), .B(n3073), .Z(n2952) );
  XNOR2_X1 U3073 ( .A(n3074), .B(n3075), .ZN(n3072) );
  XOR2_X1 U3074 ( .A(n3076), .B(n3077), .Z(n2956) );
  XNOR2_X1 U3075 ( .A(n3078), .B(n3079), .ZN(n3076) );
  XOR2_X1 U3076 ( .A(n3080), .B(n3081), .Z(n2960) );
  XNOR2_X1 U3077 ( .A(n3082), .B(n3083), .ZN(n3080) );
  XNOR2_X1 U3078 ( .A(n3084), .B(n3085), .ZN(n2964) );
  XOR2_X1 U3079 ( .A(n3086), .B(n3087), .Z(n3085) );
  XOR2_X1 U3080 ( .A(n3088), .B(n3089), .Z(n2968) );
  XNOR2_X1 U3081 ( .A(n3090), .B(n3091), .ZN(n3088) );
  XOR2_X1 U3082 ( .A(n3092), .B(n3093), .Z(n2972) );
  XOR2_X1 U3083 ( .A(n3094), .B(n3095), .Z(n3092) );
  NAND2_X1 U3084 ( .A1(n2840), .A2(n2938), .ZN(n3094) );
  XOR2_X1 U3085 ( .A(n3096), .B(n3097), .Z(n2975) );
  XNOR2_X1 U3086 ( .A(n3098), .B(n3099), .ZN(n3096) );
  NOR2_X1 U3087 ( .A1(n2937), .A2(n2396), .ZN(n3099) );
  XOR2_X1 U3088 ( .A(n3100), .B(n3101), .Z(n2890) );
  NAND2_X1 U3089 ( .A1(n3102), .A2(n3103), .ZN(n3100) );
  XOR2_X1 U3090 ( .A(n3104), .B(n3105), .Z(n2980) );
  XOR2_X1 U3091 ( .A(n3106), .B(n3107), .Z(n3104) );
  NOR2_X1 U3092 ( .A1(n2937), .A2(n2508), .ZN(n3107) );
  XOR2_X1 U3093 ( .A(n3108), .B(n3109), .Z(n2874) );
  XNOR2_X1 U3094 ( .A(n3110), .B(n3111), .ZN(n3109) );
  NAND2_X1 U3095 ( .A1(n2358), .A2(n2938), .ZN(n3111) );
  XNOR2_X1 U3096 ( .A(n3112), .B(n3113), .ZN(n2988) );
  XOR2_X1 U3097 ( .A(n3114), .B(n3115), .Z(n3113) );
  NAND2_X1 U3098 ( .A1(n2492), .A2(n2938), .ZN(n3115) );
  XOR2_X1 U3099 ( .A(n3116), .B(n3117), .Z(n2164) );
  XNOR2_X1 U3100 ( .A(n3118), .B(n3119), .ZN(n3117) );
  NAND2_X1 U3101 ( .A1(n2938), .A2(n2303), .ZN(n3119) );
  NAND2_X1 U3102 ( .A1(n3120), .A2(n2994), .ZN(n2331) );
  NAND2_X1 U3103 ( .A1(n3121), .A2(n3122), .ZN(n2994) );
  NAND3_X1 U3104 ( .A1(n2303), .A2(n3123), .A3(n2938), .ZN(n3122) );
  NAND2_X1 U3105 ( .A1(n3118), .A2(n3116), .ZN(n3123) );
  INV_X1 U3106 ( .A(n3124), .ZN(n3121) );
  NOR2_X1 U3107 ( .A1(n3116), .A2(n3118), .ZN(n3124) );
  NOR2_X1 U3108 ( .A1(n3125), .A2(n3126), .ZN(n3118) );
  NOR3_X1 U3109 ( .A1(n2937), .A2(n3127), .A3(n2354), .ZN(n3126) );
  NOR2_X1 U3110 ( .A1(n3114), .A2(n3112), .ZN(n3127) );
  INV_X1 U3111 ( .A(n3128), .ZN(n3125) );
  NAND2_X1 U3112 ( .A1(n3112), .A2(n3114), .ZN(n3128) );
  NAND2_X1 U3113 ( .A1(n3129), .A2(n3130), .ZN(n3114) );
  NAND3_X1 U3114 ( .A1(n2938), .A2(n3131), .A3(n2358), .ZN(n3130) );
  NAND2_X1 U3115 ( .A1(n3110), .A2(n3108), .ZN(n3131) );
  INV_X1 U3116 ( .A(n3132), .ZN(n3129) );
  NOR2_X1 U3117 ( .A1(n3108), .A2(n3110), .ZN(n3132) );
  NOR2_X1 U3118 ( .A1(n3133), .A2(n3134), .ZN(n3110) );
  NOR3_X1 U3119 ( .A1(n2937), .A2(n3135), .A3(n2369), .ZN(n3134) );
  INV_X1 U3120 ( .A(n3136), .ZN(n3135) );
  NAND2_X1 U3121 ( .A1(n3011), .A2(n3010), .ZN(n3136) );
  NOR2_X1 U3122 ( .A1(n3010), .A2(n3011), .ZN(n3133) );
  NOR2_X1 U3123 ( .A1(n3137), .A2(n3138), .ZN(n3011) );
  NOR3_X1 U3124 ( .A1(n2937), .A2(n3139), .A3(n2508), .ZN(n3138) );
  NOR2_X1 U3125 ( .A1(n3106), .A2(n3105), .ZN(n3139) );
  INV_X1 U3126 ( .A(n3140), .ZN(n3137) );
  NAND2_X1 U3127 ( .A1(n3105), .A2(n3106), .ZN(n3140) );
  NAND2_X1 U3128 ( .A1(n3102), .A2(n3141), .ZN(n3106) );
  NAND2_X1 U3129 ( .A1(n3101), .A2(n3103), .ZN(n3141) );
  NAND2_X1 U3130 ( .A1(n3142), .A2(n3143), .ZN(n3103) );
  NAND2_X1 U3131 ( .A1(n2593), .A2(n2938), .ZN(n3143) );
  XOR2_X1 U3132 ( .A(n3144), .B(n3145), .Z(n3101) );
  XNOR2_X1 U3133 ( .A(n3146), .B(n3147), .ZN(n3145) );
  NAND2_X1 U3134 ( .A1(n2654), .A2(n3063), .ZN(n3147) );
  INV_X1 U3135 ( .A(n3148), .ZN(n3102) );
  NOR2_X1 U3136 ( .A1(n2388), .A2(n3142), .ZN(n3148) );
  NOR2_X1 U3137 ( .A1(n3149), .A2(n3150), .ZN(n3142) );
  NOR3_X1 U3138 ( .A1(n2937), .A2(n3151), .A3(n2396), .ZN(n3150) );
  INV_X1 U3139 ( .A(n3152), .ZN(n3151) );
  NAND2_X1 U3140 ( .A1(n3098), .A2(n3097), .ZN(n3152) );
  NOR2_X1 U3141 ( .A1(n3097), .A2(n3098), .ZN(n3149) );
  NOR2_X1 U3142 ( .A1(n3153), .A2(n3154), .ZN(n3098) );
  INV_X1 U3143 ( .A(n3155), .ZN(n3154) );
  NAND3_X1 U3144 ( .A1(n2938), .A2(n3156), .A3(n2840), .ZN(n3155) );
  NAND2_X1 U3145 ( .A1(n3095), .A2(n3093), .ZN(n3156) );
  NOR2_X1 U3146 ( .A1(n3093), .A2(n3095), .ZN(n3153) );
  NOR2_X1 U3147 ( .A1(n3157), .A2(n3158), .ZN(n3095) );
  INV_X1 U3148 ( .A(n3159), .ZN(n3158) );
  NAND2_X1 U3149 ( .A1(n3091), .A2(n3160), .ZN(n3159) );
  NAND2_X1 U3150 ( .A1(n3090), .A2(n3089), .ZN(n3160) );
  NOR2_X1 U3151 ( .A1(n2937), .A2(n2525), .ZN(n3091) );
  NOR2_X1 U3152 ( .A1(n3089), .A2(n3090), .ZN(n3157) );
  NOR2_X1 U3153 ( .A1(n3161), .A2(n3162), .ZN(n3090) );
  INV_X1 U3154 ( .A(n3163), .ZN(n3162) );
  NAND2_X1 U3155 ( .A1(n3087), .A2(n3164), .ZN(n3163) );
  NAND2_X1 U3156 ( .A1(n3086), .A2(n3084), .ZN(n3164) );
  NOR2_X1 U3157 ( .A1(n2424), .A2(n2937), .ZN(n3087) );
  NOR2_X1 U3158 ( .A1(n3084), .A2(n3086), .ZN(n3161) );
  NOR2_X1 U3159 ( .A1(n3165), .A2(n3166), .ZN(n3086) );
  INV_X1 U3160 ( .A(n3167), .ZN(n3166) );
  NAND2_X1 U3161 ( .A1(n3082), .A2(n3168), .ZN(n3167) );
  NAND2_X1 U3162 ( .A1(n3083), .A2(n3081), .ZN(n3168) );
  NOR2_X1 U3163 ( .A1(n2429), .A2(n2937), .ZN(n3082) );
  NOR2_X1 U3164 ( .A1(n3081), .A2(n3083), .ZN(n3165) );
  NOR2_X1 U3165 ( .A1(n3169), .A2(n3170), .ZN(n3083) );
  INV_X1 U3166 ( .A(n3171), .ZN(n3170) );
  NAND2_X1 U3167 ( .A1(n3078), .A2(n3172), .ZN(n3171) );
  NAND2_X1 U3168 ( .A1(n3079), .A2(n3077), .ZN(n3172) );
  NOR2_X1 U3169 ( .A1(n2434), .A2(n2937), .ZN(n3078) );
  NOR2_X1 U3170 ( .A1(n3077), .A2(n3079), .ZN(n3169) );
  NOR2_X1 U3171 ( .A1(n3173), .A2(n3174), .ZN(n3079) );
  INV_X1 U3172 ( .A(n3175), .ZN(n3174) );
  NAND2_X1 U3173 ( .A1(n3074), .A2(n3176), .ZN(n3175) );
  NAND2_X1 U3174 ( .A1(n3075), .A2(n3073), .ZN(n3176) );
  NOR2_X1 U3175 ( .A1(n2542), .A2(n2937), .ZN(n3074) );
  NOR2_X1 U3176 ( .A1(n3073), .A2(n3075), .ZN(n3173) );
  NOR2_X1 U3177 ( .A1(n3177), .A2(n3178), .ZN(n3075) );
  NOR2_X1 U3178 ( .A1(n3068), .A2(n3179), .ZN(n3178) );
  NOR2_X1 U3179 ( .A1(n3071), .A2(n3070), .ZN(n3179) );
  NAND2_X1 U3180 ( .A1(n2447), .A2(n2938), .ZN(n3068) );
  INV_X1 U3181 ( .A(n2937), .ZN(n2938) );
  INV_X1 U3182 ( .A(n3180), .ZN(n3177) );
  NAND2_X1 U3183 ( .A1(n3070), .A2(n3071), .ZN(n3180) );
  NAND2_X1 U3184 ( .A1(n3181), .A2(n3182), .ZN(n3071) );
  NAND2_X1 U3185 ( .A1(n3063), .A2(n3183), .ZN(n3182) );
  NAND2_X1 U3186 ( .A1(n2202), .A2(n3184), .ZN(n3183) );
  NAND2_X1 U3187 ( .A1(n3185), .A2(n2205), .ZN(n3184) );
  NAND2_X1 U3188 ( .A1(n3186), .A2(n3187), .ZN(n3181) );
  NAND2_X1 U3189 ( .A1(n2208), .A2(n3188), .ZN(n3187) );
  NAND2_X1 U3190 ( .A1(n2210), .A2(n3062), .ZN(n3188) );
  NOR3_X1 U3191 ( .A1(n2937), .A2(n3062), .A3(n2449), .ZN(n3070) );
  XOR2_X1 U3192 ( .A(d_9_), .B(c_9_), .Z(n3190) );
  XNOR2_X1 U3193 ( .A(n3191), .B(n3192), .ZN(n3073) );
  XNOR2_X1 U3194 ( .A(n3193), .B(n3194), .ZN(n3192) );
  XOR2_X1 U3195 ( .A(n3195), .B(n3196), .Z(n3077) );
  XNOR2_X1 U3196 ( .A(n3197), .B(n3198), .ZN(n3195) );
  XOR2_X1 U3197 ( .A(n3199), .B(n3200), .Z(n3081) );
  XNOR2_X1 U3198 ( .A(n3201), .B(n3202), .ZN(n3199) );
  XOR2_X1 U3199 ( .A(n3203), .B(n3204), .Z(n3084) );
  XNOR2_X1 U3200 ( .A(n3205), .B(n3206), .ZN(n3203) );
  XOR2_X1 U3201 ( .A(n3207), .B(n3208), .Z(n3089) );
  XNOR2_X1 U3202 ( .A(n3209), .B(n3210), .ZN(n3207) );
  XOR2_X1 U3203 ( .A(n3211), .B(n3212), .Z(n3093) );
  XNOR2_X1 U3204 ( .A(n3213), .B(n3214), .ZN(n3211) );
  XOR2_X1 U3205 ( .A(n3215), .B(n3216), .Z(n3097) );
  XOR2_X1 U3206 ( .A(n3217), .B(n3218), .Z(n3215) );
  NAND2_X1 U3207 ( .A1(n2840), .A2(n3063), .ZN(n3217) );
  XNOR2_X1 U3208 ( .A(n3219), .B(n3220), .ZN(n3105) );
  XOR2_X1 U3209 ( .A(n3221), .B(n3222), .Z(n3220) );
  NAND2_X1 U3210 ( .A1(n2593), .A2(n3063), .ZN(n3222) );
  XOR2_X1 U3211 ( .A(n3223), .B(n3224), .Z(n3010) );
  NAND2_X1 U3212 ( .A1(n3225), .A2(n3226), .ZN(n3223) );
  XNOR2_X1 U3213 ( .A(n3227), .B(n3228), .ZN(n3108) );
  XOR2_X1 U3214 ( .A(n3229), .B(n3230), .Z(n3227) );
  XNOR2_X1 U3215 ( .A(n3231), .B(n3232), .ZN(n3112) );
  XNOR2_X1 U3216 ( .A(n3233), .B(n3234), .ZN(n3231) );
  XOR2_X1 U3217 ( .A(n3235), .B(n3236), .Z(n3116) );
  XNOR2_X1 U3218 ( .A(n3237), .B(n3238), .ZN(n3235) );
  XNOR2_X1 U3219 ( .A(n2995), .B(n2997), .ZN(n3120) );
  NAND2_X1 U3220 ( .A1(n3239), .A2(n3240), .ZN(n2995) );
  XOR2_X1 U3221 ( .A(n2174), .B(n2175), .Z(n2167) );
  NAND3_X1 U3222 ( .A1(n2174), .A2(n2175), .A3(n2330), .ZN(n2170) );
  INV_X1 U3223 ( .A(n2173), .ZN(n2330) );
  NAND2_X1 U3224 ( .A1(n3241), .A2(n2327), .ZN(n2173) );
  NAND2_X1 U3225 ( .A1(n3242), .A2(n3243), .ZN(n3241) );
  INV_X1 U3226 ( .A(n3244), .ZN(n3243) );
  XNOR2_X1 U3227 ( .A(n3245), .B(n3246), .ZN(n3242) );
  INV_X1 U3228 ( .A(n3247), .ZN(n3246) );
  NAND2_X1 U3229 ( .A1(n3239), .A2(n3248), .ZN(n2175) );
  NAND2_X1 U3230 ( .A1(n2997), .A2(n3240), .ZN(n3248) );
  NAND2_X1 U3231 ( .A1(n3249), .A2(n3250), .ZN(n3240) );
  NAND2_X1 U3232 ( .A1(n3063), .A2(n2303), .ZN(n3250) );
  INV_X1 U3233 ( .A(n3251), .ZN(n3249) );
  XOR2_X1 U3234 ( .A(n3252), .B(n3253), .Z(n2997) );
  XNOR2_X1 U3235 ( .A(n3254), .B(n3255), .ZN(n3253) );
  NAND2_X1 U3236 ( .A1(n2492), .A2(n3186), .ZN(n3255) );
  NAND2_X1 U3237 ( .A1(n2303), .A2(n3251), .ZN(n3239) );
  NAND2_X1 U3238 ( .A1(n3256), .A2(n3257), .ZN(n3251) );
  NAND2_X1 U3239 ( .A1(n3238), .A2(n3258), .ZN(n3257) );
  NAND2_X1 U3240 ( .A1(n3237), .A2(n3236), .ZN(n3258) );
  NOR2_X1 U3241 ( .A1(n2354), .A2(n3062), .ZN(n3238) );
  INV_X1 U3242 ( .A(n3259), .ZN(n3256) );
  NOR2_X1 U3243 ( .A1(n3236), .A2(n3237), .ZN(n3259) );
  NOR2_X1 U3244 ( .A1(n3260), .A2(n3261), .ZN(n3237) );
  INV_X1 U3245 ( .A(n3262), .ZN(n3261) );
  NAND2_X1 U3246 ( .A1(n3234), .A2(n3263), .ZN(n3262) );
  NAND2_X1 U3247 ( .A1(n3233), .A2(n3232), .ZN(n3263) );
  NOR2_X1 U3248 ( .A1(n2497), .A2(n3062), .ZN(n3234) );
  NOR2_X1 U3249 ( .A1(n3232), .A2(n3233), .ZN(n3260) );
  INV_X1 U3250 ( .A(n3264), .ZN(n3233) );
  NAND2_X1 U3251 ( .A1(n3265), .A2(n3266), .ZN(n3264) );
  NAND2_X1 U3252 ( .A1(n3230), .A2(n3267), .ZN(n3266) );
  INV_X1 U3253 ( .A(n3268), .ZN(n3267) );
  NOR2_X1 U3254 ( .A1(n3228), .A2(n3229), .ZN(n3268) );
  NOR2_X1 U3255 ( .A1(n2369), .A2(n3062), .ZN(n3230) );
  NAND2_X1 U3256 ( .A1(n3228), .A2(n3229), .ZN(n3265) );
  NAND2_X1 U3257 ( .A1(n3225), .A2(n3269), .ZN(n3229) );
  NAND2_X1 U3258 ( .A1(n3224), .A2(n3226), .ZN(n3269) );
  NAND2_X1 U3259 ( .A1(n3270), .A2(n3271), .ZN(n3226) );
  NAND2_X1 U3260 ( .A1(n2378), .A2(n3063), .ZN(n3271) );
  XOR2_X1 U3261 ( .A(n3272), .B(n3273), .Z(n3224) );
  XOR2_X1 U3262 ( .A(n3274), .B(n3275), .Z(n3272) );
  NOR2_X1 U3263 ( .A1(n3185), .A2(n2388), .ZN(n3275) );
  INV_X1 U3264 ( .A(n3276), .ZN(n3225) );
  NOR2_X1 U3265 ( .A1(n2508), .A2(n3270), .ZN(n3276) );
  NOR2_X1 U3266 ( .A1(n3277), .A2(n3278), .ZN(n3270) );
  NOR3_X1 U3267 ( .A1(n3062), .A2(n3279), .A3(n2388), .ZN(n3278) );
  NOR2_X1 U3268 ( .A1(n3219), .A2(n3221), .ZN(n3279) );
  INV_X1 U3269 ( .A(n3280), .ZN(n3277) );
  NAND2_X1 U3270 ( .A1(n3219), .A2(n3221), .ZN(n3280) );
  NAND2_X1 U3271 ( .A1(n3281), .A2(n3282), .ZN(n3221) );
  NAND3_X1 U3272 ( .A1(n3063), .A2(n3283), .A3(n2654), .ZN(n3282) );
  NAND2_X1 U3273 ( .A1(n3146), .A2(n3144), .ZN(n3283) );
  INV_X1 U3274 ( .A(n3284), .ZN(n3281) );
  NOR2_X1 U3275 ( .A1(n3144), .A2(n3146), .ZN(n3284) );
  NOR2_X1 U3276 ( .A1(n3285), .A2(n3286), .ZN(n3146) );
  INV_X1 U3277 ( .A(n3287), .ZN(n3286) );
  NAND3_X1 U3278 ( .A1(n3063), .A2(n3288), .A3(n2840), .ZN(n3287) );
  NAND2_X1 U3279 ( .A1(n3218), .A2(n3216), .ZN(n3288) );
  NOR2_X1 U3280 ( .A1(n3216), .A2(n3218), .ZN(n3285) );
  NOR2_X1 U3281 ( .A1(n3289), .A2(n3290), .ZN(n3218) );
  INV_X1 U3282 ( .A(n3291), .ZN(n3290) );
  NAND2_X1 U3283 ( .A1(n3214), .A2(n3292), .ZN(n3291) );
  NAND2_X1 U3284 ( .A1(n3213), .A2(n3212), .ZN(n3292) );
  NOR2_X1 U3285 ( .A1(n3062), .A2(n2525), .ZN(n3214) );
  NOR2_X1 U3286 ( .A1(n3212), .A2(n3213), .ZN(n3289) );
  NOR2_X1 U3287 ( .A1(n3293), .A2(n3294), .ZN(n3213) );
  INV_X1 U3288 ( .A(n3295), .ZN(n3294) );
  NAND2_X1 U3289 ( .A1(n3210), .A2(n3296), .ZN(n3295) );
  NAND2_X1 U3290 ( .A1(n3208), .A2(n3209), .ZN(n3296) );
  NOR2_X1 U3291 ( .A1(n3062), .A2(n2424), .ZN(n3210) );
  NOR2_X1 U3292 ( .A1(n3208), .A2(n3209), .ZN(n3293) );
  NOR2_X1 U3293 ( .A1(n3297), .A2(n3298), .ZN(n3209) );
  INV_X1 U3294 ( .A(n3299), .ZN(n3298) );
  NAND2_X1 U3295 ( .A1(n3206), .A2(n3300), .ZN(n3299) );
  NAND2_X1 U3296 ( .A1(n3205), .A2(n3204), .ZN(n3300) );
  NOR2_X1 U3297 ( .A1(n3062), .A2(n2429), .ZN(n3206) );
  NOR2_X1 U3298 ( .A1(n3204), .A2(n3205), .ZN(n3297) );
  NOR2_X1 U3299 ( .A1(n3301), .A2(n3302), .ZN(n3205) );
  INV_X1 U3300 ( .A(n3303), .ZN(n3302) );
  NAND2_X1 U3301 ( .A1(n3201), .A2(n3304), .ZN(n3303) );
  NAND2_X1 U3302 ( .A1(n3200), .A2(n3202), .ZN(n3304) );
  NOR2_X1 U3303 ( .A1(n3062), .A2(n2434), .ZN(n3201) );
  NOR2_X1 U3304 ( .A1(n3200), .A2(n3202), .ZN(n3301) );
  NOR2_X1 U3305 ( .A1(n3305), .A2(n3306), .ZN(n3202) );
  INV_X1 U3306 ( .A(n3307), .ZN(n3306) );
  NAND2_X1 U3307 ( .A1(n3197), .A2(n3308), .ZN(n3307) );
  NAND2_X1 U3308 ( .A1(n3198), .A2(n3196), .ZN(n3308) );
  NOR2_X1 U3309 ( .A1(n3062), .A2(n2542), .ZN(n3197) );
  NOR2_X1 U3310 ( .A1(n3196), .A2(n3198), .ZN(n3305) );
  NOR2_X1 U3311 ( .A1(n3309), .A2(n3310), .ZN(n3198) );
  NOR2_X1 U3312 ( .A1(n3191), .A2(n3311), .ZN(n3310) );
  NOR2_X1 U3313 ( .A1(n3194), .A2(n3193), .ZN(n3311) );
  NAND2_X1 U3314 ( .A1(n3063), .A2(n2447), .ZN(n3191) );
  INV_X1 U3315 ( .A(n3062), .ZN(n3063) );
  INV_X1 U3316 ( .A(n3312), .ZN(n3309) );
  NAND2_X1 U3317 ( .A1(n3193), .A2(n3194), .ZN(n3312) );
  NAND2_X1 U3318 ( .A1(n3313), .A2(n3314), .ZN(n3194) );
  NAND2_X1 U3319 ( .A1(n3186), .A2(n3315), .ZN(n3314) );
  NAND2_X1 U3320 ( .A1(n2202), .A2(n3316), .ZN(n3315) );
  NAND2_X1 U3321 ( .A1(n3317), .A2(n2205), .ZN(n3316) );
  NAND2_X1 U3322 ( .A1(n3318), .A2(n3319), .ZN(n3313) );
  NAND2_X1 U3323 ( .A1(n2208), .A2(n3320), .ZN(n3319) );
  NAND2_X1 U3324 ( .A1(n2210), .A2(n3185), .ZN(n3320) );
  NOR3_X1 U3325 ( .A1(n3062), .A2(n2449), .A3(n3185), .ZN(n3193) );
  XOR2_X1 U3326 ( .A(d_8_), .B(c_8_), .Z(n3322) );
  XNOR2_X1 U3327 ( .A(n3323), .B(n3324), .ZN(n3196) );
  XNOR2_X1 U3328 ( .A(n3325), .B(n3326), .ZN(n3324) );
  XOR2_X1 U3329 ( .A(n3327), .B(n3328), .Z(n3200) );
  XNOR2_X1 U3330 ( .A(n3329), .B(n3330), .ZN(n3327) );
  XOR2_X1 U3331 ( .A(n3331), .B(n3332), .Z(n3204) );
  XNOR2_X1 U3332 ( .A(n3333), .B(n3334), .ZN(n3331) );
  XOR2_X1 U3333 ( .A(n3335), .B(n3336), .Z(n3208) );
  XNOR2_X1 U3334 ( .A(n3337), .B(n3338), .ZN(n3335) );
  XOR2_X1 U3335 ( .A(n3339), .B(n3340), .Z(n3212) );
  XNOR2_X1 U3336 ( .A(n3341), .B(n3342), .ZN(n3339) );
  XOR2_X1 U3337 ( .A(n3343), .B(n3344), .Z(n3216) );
  XNOR2_X1 U3338 ( .A(n3345), .B(n3346), .ZN(n3343) );
  XNOR2_X1 U3339 ( .A(n3347), .B(n3348), .ZN(n3144) );
  XOR2_X1 U3340 ( .A(n3349), .B(n3350), .Z(n3347) );
  XOR2_X1 U3341 ( .A(n3351), .B(n3352), .Z(n3219) );
  XOR2_X1 U3342 ( .A(n3353), .B(n3354), .Z(n3351) );
  NOR2_X1 U3343 ( .A1(n3185), .A2(n2396), .ZN(n3354) );
  XNOR2_X1 U3344 ( .A(n3355), .B(n3356), .ZN(n3228) );
  XOR2_X1 U3345 ( .A(n3357), .B(n3358), .Z(n3356) );
  NAND2_X1 U3346 ( .A1(n2378), .A2(n3186), .ZN(n3358) );
  XOR2_X1 U3347 ( .A(n3359), .B(n3360), .Z(n3232) );
  XOR2_X1 U3348 ( .A(n3361), .B(n3362), .Z(n3360) );
  NAND2_X1 U3349 ( .A1(n2641), .A2(n3186), .ZN(n3362) );
  XNOR2_X1 U3350 ( .A(n3363), .B(n3364), .ZN(n3236) );
  XNOR2_X1 U3351 ( .A(n3365), .B(n3366), .ZN(n3364) );
  NAND2_X1 U3352 ( .A1(n2358), .A2(n3186), .ZN(n3366) );
  XNOR2_X1 U3353 ( .A(n3367), .B(n3368), .ZN(n2174) );
  XNOR2_X1 U3354 ( .A(n3369), .B(n3370), .ZN(n3367) );
  NOR2_X1 U3355 ( .A1(n2345), .A2(n3185), .ZN(n3370) );
  NAND2_X1 U3356 ( .A1(n3371), .A2(n3244), .ZN(n2327) );
  NAND2_X1 U3357 ( .A1(n3372), .A2(n3373), .ZN(n3244) );
  NAND3_X1 U3358 ( .A1(n2303), .A2(n3374), .A3(n3186), .ZN(n3373) );
  NAND2_X1 U3359 ( .A1(n3368), .A2(n3369), .ZN(n3374) );
  INV_X1 U3360 ( .A(n3375), .ZN(n3372) );
  NOR2_X1 U3361 ( .A1(n3368), .A2(n3369), .ZN(n3375) );
  NOR2_X1 U3362 ( .A1(n3376), .A2(n3377), .ZN(n3369) );
  INV_X1 U3363 ( .A(n3378), .ZN(n3377) );
  NAND3_X1 U3364 ( .A1(n3186), .A2(n3379), .A3(n2492), .ZN(n3378) );
  NAND2_X1 U3365 ( .A1(n3254), .A2(n3252), .ZN(n3379) );
  NOR2_X1 U3366 ( .A1(n3252), .A2(n3254), .ZN(n3376) );
  NOR2_X1 U3367 ( .A1(n3380), .A2(n3381), .ZN(n3254) );
  INV_X1 U3368 ( .A(n3382), .ZN(n3381) );
  NAND3_X1 U3369 ( .A1(n3186), .A2(n3383), .A3(n2358), .ZN(n3382) );
  NAND2_X1 U3370 ( .A1(n3363), .A2(n3365), .ZN(n3383) );
  NOR2_X1 U3371 ( .A1(n3363), .A2(n3365), .ZN(n3380) );
  NOR2_X1 U3372 ( .A1(n3384), .A2(n3385), .ZN(n3365) );
  NOR3_X1 U3373 ( .A1(n3185), .A2(n3386), .A3(n2369), .ZN(n3385) );
  NOR2_X1 U3374 ( .A1(n3359), .A2(n3361), .ZN(n3386) );
  INV_X1 U3375 ( .A(n3387), .ZN(n3384) );
  NAND2_X1 U3376 ( .A1(n3359), .A2(n3361), .ZN(n3387) );
  NAND2_X1 U3377 ( .A1(n3388), .A2(n3389), .ZN(n3361) );
  INV_X1 U3378 ( .A(n3390), .ZN(n3389) );
  NOR3_X1 U3379 ( .A1(n3185), .A2(n3391), .A3(n2508), .ZN(n3390) );
  NOR2_X1 U3380 ( .A1(n3357), .A2(n3355), .ZN(n3391) );
  NAND2_X1 U3381 ( .A1(n3355), .A2(n3357), .ZN(n3388) );
  NAND2_X1 U3382 ( .A1(n3392), .A2(n3393), .ZN(n3357) );
  NAND3_X1 U3383 ( .A1(n3186), .A2(n3394), .A3(n2593), .ZN(n3393) );
  INV_X1 U3384 ( .A(n3395), .ZN(n3394) );
  NOR2_X1 U3385 ( .A1(n3273), .A2(n3274), .ZN(n3395) );
  NAND2_X1 U3386 ( .A1(n3273), .A2(n3274), .ZN(n3392) );
  NAND2_X1 U3387 ( .A1(n3396), .A2(n3397), .ZN(n3274) );
  NAND3_X1 U3388 ( .A1(n3186), .A2(n3398), .A3(n2654), .ZN(n3397) );
  INV_X1 U3389 ( .A(n3399), .ZN(n3398) );
  NOR2_X1 U3390 ( .A1(n3353), .A2(n3352), .ZN(n3399) );
  NAND2_X1 U3391 ( .A1(n3352), .A2(n3353), .ZN(n3396) );
  NAND2_X1 U3392 ( .A1(n3400), .A2(n3401), .ZN(n3353) );
  NAND2_X1 U3393 ( .A1(n3350), .A2(n3402), .ZN(n3401) );
  INV_X1 U3394 ( .A(n3403), .ZN(n3402) );
  NOR2_X1 U3395 ( .A1(n3348), .A2(n3349), .ZN(n3403) );
  NOR2_X1 U3396 ( .A1(n2406), .A2(n3185), .ZN(n3350) );
  NAND2_X1 U3397 ( .A1(n3348), .A2(n3349), .ZN(n3400) );
  NAND2_X1 U3398 ( .A1(n3404), .A2(n3405), .ZN(n3349) );
  NAND2_X1 U3399 ( .A1(n3346), .A2(n3406), .ZN(n3405) );
  NAND2_X1 U3400 ( .A1(n3344), .A2(n3345), .ZN(n3406) );
  NOR2_X1 U3401 ( .A1(n3185), .A2(n2525), .ZN(n3346) );
  INV_X1 U3402 ( .A(n3407), .ZN(n3404) );
  NOR2_X1 U3403 ( .A1(n3344), .A2(n3345), .ZN(n3407) );
  NOR2_X1 U3404 ( .A1(n3408), .A2(n3409), .ZN(n3345) );
  INV_X1 U3405 ( .A(n3410), .ZN(n3409) );
  NAND2_X1 U3406 ( .A1(n3341), .A2(n3411), .ZN(n3410) );
  NAND2_X1 U3407 ( .A1(n3340), .A2(n3342), .ZN(n3411) );
  NOR2_X1 U3408 ( .A1(n3185), .A2(n2424), .ZN(n3341) );
  NOR2_X1 U3409 ( .A1(n3340), .A2(n3342), .ZN(n3408) );
  NOR2_X1 U3410 ( .A1(n3412), .A2(n3413), .ZN(n3342) );
  INV_X1 U3411 ( .A(n3414), .ZN(n3413) );
  NAND2_X1 U3412 ( .A1(n3338), .A2(n3415), .ZN(n3414) );
  NAND2_X1 U3413 ( .A1(n3337), .A2(n3336), .ZN(n3415) );
  NOR2_X1 U3414 ( .A1(n3185), .A2(n2429), .ZN(n3338) );
  NOR2_X1 U3415 ( .A1(n3336), .A2(n3337), .ZN(n3412) );
  NOR2_X1 U3416 ( .A1(n3416), .A2(n3417), .ZN(n3337) );
  INV_X1 U3417 ( .A(n3418), .ZN(n3417) );
  NAND2_X1 U3418 ( .A1(n3333), .A2(n3419), .ZN(n3418) );
  NAND2_X1 U3419 ( .A1(n3332), .A2(n3334), .ZN(n3419) );
  NOR2_X1 U3420 ( .A1(n3185), .A2(n2434), .ZN(n3333) );
  NOR2_X1 U3421 ( .A1(n3332), .A2(n3334), .ZN(n3416) );
  NOR2_X1 U3422 ( .A1(n3420), .A2(n3421), .ZN(n3334) );
  INV_X1 U3423 ( .A(n3422), .ZN(n3421) );
  NAND2_X1 U3424 ( .A1(n3329), .A2(n3423), .ZN(n3422) );
  NAND2_X1 U3425 ( .A1(n3330), .A2(n3328), .ZN(n3423) );
  NOR2_X1 U3426 ( .A1(n3185), .A2(n2542), .ZN(n3329) );
  NOR2_X1 U3427 ( .A1(n3328), .A2(n3330), .ZN(n3420) );
  NOR2_X1 U3428 ( .A1(n3424), .A2(n3425), .ZN(n3330) );
  NOR2_X1 U3429 ( .A1(n3323), .A2(n3426), .ZN(n3425) );
  NOR2_X1 U3430 ( .A1(n3326), .A2(n3325), .ZN(n3426) );
  NAND2_X1 U3431 ( .A1(n3186), .A2(n2447), .ZN(n3323) );
  INV_X1 U3432 ( .A(n3185), .ZN(n3186) );
  INV_X1 U3433 ( .A(n3427), .ZN(n3424) );
  NAND2_X1 U3434 ( .A1(n3325), .A2(n3326), .ZN(n3427) );
  NAND2_X1 U3435 ( .A1(n3428), .A2(n3429), .ZN(n3326) );
  NAND2_X1 U3436 ( .A1(n3318), .A2(n3430), .ZN(n3429) );
  NAND2_X1 U3437 ( .A1(n2202), .A2(n3431), .ZN(n3430) );
  NAND2_X1 U3438 ( .A1(n3432), .A2(n2205), .ZN(n3431) );
  NAND2_X1 U3439 ( .A1(n3433), .A2(n3434), .ZN(n3428) );
  NAND2_X1 U3440 ( .A1(n2208), .A2(n3435), .ZN(n3434) );
  NAND2_X1 U3441 ( .A1(n2210), .A2(n3317), .ZN(n3435) );
  NOR3_X1 U3442 ( .A1(n3185), .A2(n2449), .A3(n3317), .ZN(n3325) );
  XOR2_X1 U3443 ( .A(d_7_), .B(c_7_), .Z(n3437) );
  XNOR2_X1 U3444 ( .A(n3438), .B(n3439), .ZN(n3328) );
  XNOR2_X1 U3445 ( .A(n3440), .B(n3441), .ZN(n3439) );
  XOR2_X1 U3446 ( .A(n3442), .B(n3443), .Z(n3332) );
  XNOR2_X1 U3447 ( .A(n3444), .B(n3445), .ZN(n3442) );
  XOR2_X1 U3448 ( .A(n3446), .B(n3447), .Z(n3336) );
  XNOR2_X1 U3449 ( .A(n3448), .B(n3449), .ZN(n3446) );
  XOR2_X1 U3450 ( .A(n3450), .B(n3451), .Z(n3340) );
  XNOR2_X1 U3451 ( .A(n3452), .B(n3453), .ZN(n3450) );
  XOR2_X1 U3452 ( .A(n3454), .B(n3455), .Z(n3344) );
  XNOR2_X1 U3453 ( .A(n3456), .B(n3457), .ZN(n3454) );
  XOR2_X1 U3454 ( .A(n3458), .B(n3459), .Z(n3348) );
  XNOR2_X1 U3455 ( .A(n3460), .B(n3461), .ZN(n3459) );
  NAND2_X1 U3456 ( .A1(n3318), .A2(n2414), .ZN(n3461) );
  XNOR2_X1 U3457 ( .A(n3462), .B(n3463), .ZN(n3352) );
  XOR2_X1 U3458 ( .A(n3464), .B(n3465), .Z(n3463) );
  NAND2_X1 U3459 ( .A1(n2840), .A2(n3318), .ZN(n3465) );
  XNOR2_X1 U3460 ( .A(n3466), .B(n3467), .ZN(n3273) );
  NAND2_X1 U3461 ( .A1(n3468), .A2(n3469), .ZN(n3466) );
  XNOR2_X1 U3462 ( .A(n3470), .B(n3471), .ZN(n3355) );
  NAND2_X1 U3463 ( .A1(n3472), .A2(n3473), .ZN(n3470) );
  XOR2_X1 U3464 ( .A(n3474), .B(n3475), .Z(n3359) );
  XOR2_X1 U3465 ( .A(n3476), .B(n3477), .Z(n3474) );
  XNOR2_X1 U3466 ( .A(n3478), .B(n3479), .ZN(n3363) );
  XOR2_X1 U3467 ( .A(n3480), .B(n3481), .Z(n3478) );
  XOR2_X1 U3468 ( .A(n3482), .B(n3483), .Z(n3252) );
  XNOR2_X1 U3469 ( .A(n3484), .B(n3485), .ZN(n3483) );
  XNOR2_X1 U3470 ( .A(n3486), .B(n3487), .ZN(n3368) );
  XOR2_X1 U3471 ( .A(n3488), .B(n3489), .Z(n3486) );
  XNOR2_X1 U3472 ( .A(n3245), .B(n3247), .ZN(n3371) );
  NAND2_X1 U3473 ( .A1(n3490), .A2(n3491), .ZN(n3245) );
  XOR2_X1 U3474 ( .A(n2185), .B(n2184), .Z(n2176) );
  NAND3_X1 U3475 ( .A1(n2185), .A2(n2184), .A3(n2326), .ZN(n2181) );
  INV_X1 U3476 ( .A(n2182), .ZN(n2326) );
  NAND2_X1 U3477 ( .A1(n3492), .A2(n2324), .ZN(n2182) );
  NAND2_X1 U3478 ( .A1(n3493), .A2(n3494), .ZN(n3492) );
  INV_X1 U3479 ( .A(n3495), .ZN(n3494) );
  XNOR2_X1 U3480 ( .A(n3496), .B(n3497), .ZN(n3493) );
  NAND2_X1 U3481 ( .A1(n3490), .A2(n3498), .ZN(n2184) );
  NAND2_X1 U3482 ( .A1(n3247), .A2(n3491), .ZN(n3498) );
  NAND2_X1 U3483 ( .A1(n3499), .A2(n3500), .ZN(n3491) );
  NAND2_X1 U3484 ( .A1(n3318), .A2(n2303), .ZN(n3500) );
  INV_X1 U3485 ( .A(n3501), .ZN(n3499) );
  XNOR2_X1 U3486 ( .A(n3502), .B(n3503), .ZN(n3247) );
  NAND2_X1 U3487 ( .A1(n3504), .A2(n3505), .ZN(n3502) );
  NAND2_X1 U3488 ( .A1(n2303), .A2(n3501), .ZN(n3490) );
  NAND2_X1 U3489 ( .A1(n3506), .A2(n3507), .ZN(n3501) );
  NAND2_X1 U3490 ( .A1(n3489), .A2(n3508), .ZN(n3507) );
  INV_X1 U3491 ( .A(n3509), .ZN(n3508) );
  NOR2_X1 U3492 ( .A1(n3488), .A2(n3487), .ZN(n3509) );
  NOR2_X1 U3493 ( .A1(n2354), .A2(n3317), .ZN(n3489) );
  NAND2_X1 U3494 ( .A1(n3487), .A2(n3488), .ZN(n3506) );
  NAND2_X1 U3495 ( .A1(n3510), .A2(n3511), .ZN(n3488) );
  NAND2_X1 U3496 ( .A1(n3485), .A2(n3512), .ZN(n3511) );
  INV_X1 U3497 ( .A(n3513), .ZN(n3512) );
  NOR2_X1 U3498 ( .A1(n3482), .A2(n3484), .ZN(n3513) );
  NOR2_X1 U3499 ( .A1(n2497), .A2(n3317), .ZN(n3485) );
  NAND2_X1 U3500 ( .A1(n3482), .A2(n3484), .ZN(n3510) );
  NAND2_X1 U3501 ( .A1(n3514), .A2(n3515), .ZN(n3484) );
  NAND2_X1 U3502 ( .A1(n3481), .A2(n3516), .ZN(n3515) );
  INV_X1 U3503 ( .A(n3517), .ZN(n3516) );
  NOR2_X1 U3504 ( .A1(n3480), .A2(n3479), .ZN(n3517) );
  NOR2_X1 U3505 ( .A1(n2369), .A2(n3317), .ZN(n3481) );
  NAND2_X1 U3506 ( .A1(n3479), .A2(n3480), .ZN(n3514) );
  NAND2_X1 U3507 ( .A1(n3518), .A2(n3519), .ZN(n3480) );
  NAND2_X1 U3508 ( .A1(n3477), .A2(n3520), .ZN(n3519) );
  INV_X1 U3509 ( .A(n3521), .ZN(n3520) );
  NOR2_X1 U3510 ( .A1(n3476), .A2(n3475), .ZN(n3521) );
  NOR2_X1 U3511 ( .A1(n2508), .A2(n3317), .ZN(n3477) );
  NAND2_X1 U3512 ( .A1(n3475), .A2(n3476), .ZN(n3518) );
  NAND2_X1 U3513 ( .A1(n3472), .A2(n3522), .ZN(n3476) );
  NAND2_X1 U3514 ( .A1(n3471), .A2(n3473), .ZN(n3522) );
  NAND2_X1 U3515 ( .A1(n3523), .A2(n3524), .ZN(n3473) );
  NAND2_X1 U3516 ( .A1(n2593), .A2(n3318), .ZN(n3524) );
  INV_X1 U3517 ( .A(n3525), .ZN(n3523) );
  XOR2_X1 U3518 ( .A(n3526), .B(n3527), .Z(n3471) );
  XNOR2_X1 U3519 ( .A(n3528), .B(n3529), .ZN(n3527) );
  NAND2_X1 U3520 ( .A1(n2654), .A2(n3433), .ZN(n3529) );
  NAND2_X1 U3521 ( .A1(n2593), .A2(n3525), .ZN(n3472) );
  NAND2_X1 U3522 ( .A1(n3468), .A2(n3530), .ZN(n3525) );
  NAND2_X1 U3523 ( .A1(n3467), .A2(n3469), .ZN(n3530) );
  NAND2_X1 U3524 ( .A1(n3531), .A2(n3532), .ZN(n3469) );
  NAND2_X1 U3525 ( .A1(n2654), .A2(n3318), .ZN(n3532) );
  XNOR2_X1 U3526 ( .A(n3533), .B(n3534), .ZN(n3467) );
  XOR2_X1 U3527 ( .A(n3535), .B(n3536), .Z(n3534) );
  NAND2_X1 U3528 ( .A1(n2840), .A2(n3433), .ZN(n3536) );
  INV_X1 U3529 ( .A(n3537), .ZN(n3468) );
  NOR2_X1 U3530 ( .A1(n2396), .A2(n3531), .ZN(n3537) );
  NOR2_X1 U3531 ( .A1(n3538), .A2(n3539), .ZN(n3531) );
  NOR3_X1 U3532 ( .A1(n3317), .A2(n3540), .A3(n2406), .ZN(n3539) );
  NOR2_X1 U3533 ( .A1(n3462), .A2(n3464), .ZN(n3540) );
  INV_X1 U3534 ( .A(n3541), .ZN(n3538) );
  NAND2_X1 U3535 ( .A1(n3462), .A2(n3464), .ZN(n3541) );
  NAND2_X1 U3536 ( .A1(n3542), .A2(n3543), .ZN(n3464) );
  NAND3_X1 U3537 ( .A1(n2414), .A2(n3544), .A3(n3318), .ZN(n3543) );
  NAND2_X1 U3538 ( .A1(n3460), .A2(n3458), .ZN(n3544) );
  NAND2_X1 U3539 ( .A1(n3545), .A2(n3546), .ZN(n3542) );
  INV_X1 U3540 ( .A(n3460), .ZN(n3546) );
  NOR2_X1 U3541 ( .A1(n3547), .A2(n3548), .ZN(n3460) );
  INV_X1 U3542 ( .A(n3549), .ZN(n3548) );
  NAND2_X1 U3543 ( .A1(n3456), .A2(n3550), .ZN(n3549) );
  NAND2_X1 U3544 ( .A1(n3457), .A2(n3455), .ZN(n3550) );
  NOR2_X1 U3545 ( .A1(n3317), .A2(n2424), .ZN(n3456) );
  NOR2_X1 U3546 ( .A1(n3455), .A2(n3457), .ZN(n3547) );
  NOR2_X1 U3547 ( .A1(n3551), .A2(n3552), .ZN(n3457) );
  INV_X1 U3548 ( .A(n3553), .ZN(n3552) );
  NAND2_X1 U3549 ( .A1(n3453), .A2(n3554), .ZN(n3553) );
  NAND2_X1 U3550 ( .A1(n3452), .A2(n3451), .ZN(n3554) );
  NOR2_X1 U3551 ( .A1(n3317), .A2(n2429), .ZN(n3453) );
  NOR2_X1 U3552 ( .A1(n3451), .A2(n3452), .ZN(n3551) );
  NOR2_X1 U3553 ( .A1(n3555), .A2(n3556), .ZN(n3452) );
  INV_X1 U3554 ( .A(n3557), .ZN(n3556) );
  NAND2_X1 U3555 ( .A1(n3448), .A2(n3558), .ZN(n3557) );
  NAND2_X1 U3556 ( .A1(n3447), .A2(n3449), .ZN(n3558) );
  NOR2_X1 U3557 ( .A1(n3317), .A2(n2434), .ZN(n3448) );
  NOR2_X1 U3558 ( .A1(n3447), .A2(n3449), .ZN(n3555) );
  NOR2_X1 U3559 ( .A1(n3559), .A2(n3560), .ZN(n3449) );
  INV_X1 U3560 ( .A(n3561), .ZN(n3560) );
  NAND2_X1 U3561 ( .A1(n3444), .A2(n3562), .ZN(n3561) );
  NAND2_X1 U3562 ( .A1(n3445), .A2(n3443), .ZN(n3562) );
  NOR2_X1 U3563 ( .A1(n3317), .A2(n2542), .ZN(n3444) );
  NOR2_X1 U3564 ( .A1(n3443), .A2(n3445), .ZN(n3559) );
  NOR2_X1 U3565 ( .A1(n3563), .A2(n3564), .ZN(n3445) );
  NOR2_X1 U3566 ( .A1(n3438), .A2(n3565), .ZN(n3564) );
  NOR2_X1 U3567 ( .A1(n3441), .A2(n3440), .ZN(n3565) );
  NAND2_X1 U3568 ( .A1(n3318), .A2(n2447), .ZN(n3438) );
  INV_X1 U3569 ( .A(n3317), .ZN(n3318) );
  INV_X1 U3570 ( .A(n3566), .ZN(n3563) );
  NAND2_X1 U3571 ( .A1(n3440), .A2(n3441), .ZN(n3566) );
  NAND2_X1 U3572 ( .A1(n3567), .A2(n3568), .ZN(n3441) );
  NAND2_X1 U3573 ( .A1(n3433), .A2(n3569), .ZN(n3568) );
  NAND2_X1 U3574 ( .A1(n2202), .A2(n3570), .ZN(n3569) );
  NAND2_X1 U3575 ( .A1(n3571), .A2(n2205), .ZN(n3570) );
  NAND2_X1 U3576 ( .A1(n3572), .A2(n3573), .ZN(n3567) );
  NAND2_X1 U3577 ( .A1(n2208), .A2(n3574), .ZN(n3573) );
  NAND2_X1 U3578 ( .A1(n2210), .A2(n3432), .ZN(n3574) );
  NOR3_X1 U3579 ( .A1(n3317), .A2(n2449), .A3(n3432), .ZN(n3440) );
  XOR2_X1 U3580 ( .A(d_6_), .B(c_6_), .Z(n3576) );
  XNOR2_X1 U3581 ( .A(n3577), .B(n3578), .ZN(n3443) );
  XNOR2_X1 U3582 ( .A(n3579), .B(n3580), .ZN(n3578) );
  XOR2_X1 U3583 ( .A(n3581), .B(n3582), .Z(n3447) );
  XNOR2_X1 U3584 ( .A(n3583), .B(n3584), .ZN(n3581) );
  XOR2_X1 U3585 ( .A(n3585), .B(n3586), .Z(n3451) );
  XNOR2_X1 U3586 ( .A(n3587), .B(n3588), .ZN(n3585) );
  XOR2_X1 U3587 ( .A(n3589), .B(n3590), .Z(n3455) );
  XNOR2_X1 U3588 ( .A(n3591), .B(n3592), .ZN(n3589) );
  INV_X1 U3589 ( .A(n3458), .ZN(n3545) );
  XNOR2_X1 U3590 ( .A(n3593), .B(n3594), .ZN(n3458) );
  XOR2_X1 U3591 ( .A(n3595), .B(n3596), .Z(n3593) );
  XNOR2_X1 U3592 ( .A(n3597), .B(n3598), .ZN(n3462) );
  NAND2_X1 U3593 ( .A1(n3599), .A2(n3600), .ZN(n3597) );
  XOR2_X1 U3594 ( .A(n3601), .B(n3602), .Z(n3475) );
  XNOR2_X1 U3595 ( .A(n3603), .B(n3604), .ZN(n3602) );
  NAND2_X1 U3596 ( .A1(n2593), .A2(n3433), .ZN(n3604) );
  XNOR2_X1 U3597 ( .A(n3605), .B(n3606), .ZN(n3479) );
  XNOR2_X1 U3598 ( .A(n3607), .B(n3608), .ZN(n3605) );
  NOR2_X1 U3599 ( .A1(n3432), .A2(n2508), .ZN(n3608) );
  XNOR2_X1 U3600 ( .A(n3609), .B(n3610), .ZN(n3482) );
  NAND2_X1 U3601 ( .A1(n3611), .A2(n3612), .ZN(n3609) );
  XOR2_X1 U3602 ( .A(n3613), .B(n3614), .Z(n3487) );
  XOR2_X1 U3603 ( .A(n3615), .B(n3616), .Z(n3613) );
  NOR2_X1 U3604 ( .A1(n3432), .A2(n2497), .ZN(n3616) );
  XOR2_X1 U3605 ( .A(n3617), .B(n3618), .Z(n2185) );
  XOR2_X1 U3606 ( .A(n3619), .B(n3620), .Z(n3617) );
  NOR2_X1 U3607 ( .A1(n2345), .A2(n3432), .ZN(n3620) );
  NAND2_X1 U3608 ( .A1(n3621), .A2(n3495), .ZN(n2324) );
  NAND2_X1 U3609 ( .A1(n3622), .A2(n3623), .ZN(n3495) );
  INV_X1 U3610 ( .A(n3624), .ZN(n3623) );
  NOR3_X1 U3611 ( .A1(n2345), .A2(n3625), .A3(n3432), .ZN(n3624) );
  NOR2_X1 U3612 ( .A1(n3618), .A2(n3619), .ZN(n3625) );
  NAND2_X1 U3613 ( .A1(n3618), .A2(n3619), .ZN(n3622) );
  NAND2_X1 U3614 ( .A1(n3504), .A2(n3626), .ZN(n3619) );
  NAND2_X1 U3615 ( .A1(n3503), .A2(n3505), .ZN(n3626) );
  NAND2_X1 U3616 ( .A1(n3627), .A2(n3628), .ZN(n3505) );
  NAND2_X1 U3617 ( .A1(n2492), .A2(n3433), .ZN(n3628) );
  INV_X1 U3618 ( .A(n3629), .ZN(n3627) );
  XNOR2_X1 U3619 ( .A(n3630), .B(n3631), .ZN(n3503) );
  XNOR2_X1 U3620 ( .A(n3632), .B(n3633), .ZN(n3630) );
  NAND2_X1 U3621 ( .A1(n2492), .A2(n3629), .ZN(n3504) );
  NAND2_X1 U3622 ( .A1(n3634), .A2(n3635), .ZN(n3629) );
  NAND3_X1 U3623 ( .A1(n3433), .A2(n3636), .A3(n2358), .ZN(n3635) );
  INV_X1 U3624 ( .A(n3637), .ZN(n3636) );
  NOR2_X1 U3625 ( .A1(n3614), .A2(n3615), .ZN(n3637) );
  NAND2_X1 U3626 ( .A1(n3614), .A2(n3615), .ZN(n3634) );
  NAND2_X1 U3627 ( .A1(n3611), .A2(n3638), .ZN(n3615) );
  NAND2_X1 U3628 ( .A1(n3610), .A2(n3612), .ZN(n3638) );
  NAND2_X1 U3629 ( .A1(n3639), .A2(n3640), .ZN(n3612) );
  NAND2_X1 U3630 ( .A1(n2641), .A2(n3433), .ZN(n3640) );
  INV_X1 U3631 ( .A(n3641), .ZN(n3639) );
  XNOR2_X1 U3632 ( .A(n3642), .B(n3643), .ZN(n3610) );
  XNOR2_X1 U3633 ( .A(n3644), .B(n3645), .ZN(n3642) );
  NAND2_X1 U3634 ( .A1(n2641), .A2(n3641), .ZN(n3611) );
  NAND2_X1 U3635 ( .A1(n3646), .A2(n3647), .ZN(n3641) );
  NAND3_X1 U3636 ( .A1(n3433), .A2(n3648), .A3(n2378), .ZN(n3647) );
  NAND2_X1 U3637 ( .A1(n3606), .A2(n3607), .ZN(n3648) );
  INV_X1 U3638 ( .A(n3649), .ZN(n3646) );
  NOR2_X1 U3639 ( .A1(n3606), .A2(n3607), .ZN(n3649) );
  NOR2_X1 U3640 ( .A1(n3650), .A2(n3651), .ZN(n3607) );
  INV_X1 U3641 ( .A(n3652), .ZN(n3651) );
  NAND3_X1 U3642 ( .A1(n3433), .A2(n3653), .A3(n2593), .ZN(n3652) );
  NAND2_X1 U3643 ( .A1(n3601), .A2(n3603), .ZN(n3653) );
  NOR2_X1 U3644 ( .A1(n3601), .A2(n3603), .ZN(n3650) );
  NOR2_X1 U3645 ( .A1(n3654), .A2(n3655), .ZN(n3603) );
  INV_X1 U3646 ( .A(n3656), .ZN(n3655) );
  NAND3_X1 U3647 ( .A1(n3433), .A2(n3657), .A3(n2654), .ZN(n3656) );
  NAND2_X1 U3648 ( .A1(n3526), .A2(n3528), .ZN(n3657) );
  NOR2_X1 U3649 ( .A1(n3526), .A2(n3528), .ZN(n3654) );
  NOR2_X1 U3650 ( .A1(n3658), .A2(n3659), .ZN(n3528) );
  NOR3_X1 U3651 ( .A1(n3432), .A2(n3660), .A3(n2406), .ZN(n3659) );
  NOR2_X1 U3652 ( .A1(n3535), .A2(n3533), .ZN(n3660) );
  INV_X1 U3653 ( .A(n3661), .ZN(n3658) );
  NAND2_X1 U3654 ( .A1(n3533), .A2(n3535), .ZN(n3661) );
  NAND2_X1 U3655 ( .A1(n3599), .A2(n3662), .ZN(n3535) );
  NAND2_X1 U3656 ( .A1(n3598), .A2(n3600), .ZN(n3662) );
  NAND2_X1 U3657 ( .A1(n3663), .A2(n3664), .ZN(n3600) );
  NAND2_X1 U3658 ( .A1(n3433), .A2(n2414), .ZN(n3664) );
  INV_X1 U3659 ( .A(n3665), .ZN(n3663) );
  XOR2_X1 U3660 ( .A(n3666), .B(n3667), .Z(n3598) );
  XNOR2_X1 U3661 ( .A(n3668), .B(n3669), .ZN(n3667) );
  NAND2_X1 U3662 ( .A1(n3572), .A2(n3670), .ZN(n3669) );
  NAND2_X1 U3663 ( .A1(n2414), .A2(n3665), .ZN(n3599) );
  NAND2_X1 U3664 ( .A1(n3671), .A2(n3672), .ZN(n3665) );
  NAND2_X1 U3665 ( .A1(n3596), .A2(n3673), .ZN(n3672) );
  INV_X1 U3666 ( .A(n3674), .ZN(n3673) );
  NOR2_X1 U3667 ( .A1(n3594), .A2(n3595), .ZN(n3674) );
  NOR2_X1 U3668 ( .A1(n3432), .A2(n2424), .ZN(n3596) );
  NAND2_X1 U3669 ( .A1(n3594), .A2(n3595), .ZN(n3671) );
  NAND2_X1 U3670 ( .A1(n3675), .A2(n3676), .ZN(n3595) );
  NAND2_X1 U3671 ( .A1(n3592), .A2(n3677), .ZN(n3676) );
  NAND2_X1 U3672 ( .A1(n3590), .A2(n3591), .ZN(n3677) );
  NOR2_X1 U3673 ( .A1(n3432), .A2(n2429), .ZN(n3592) );
  INV_X1 U3674 ( .A(n3678), .ZN(n3675) );
  NOR2_X1 U3675 ( .A1(n3590), .A2(n3591), .ZN(n3678) );
  NOR2_X1 U3676 ( .A1(n3679), .A2(n3680), .ZN(n3591) );
  INV_X1 U3677 ( .A(n3681), .ZN(n3680) );
  NAND2_X1 U3678 ( .A1(n3587), .A2(n3682), .ZN(n3681) );
  NAND2_X1 U3679 ( .A1(n3586), .A2(n3588), .ZN(n3682) );
  NOR2_X1 U3680 ( .A1(n3432), .A2(n2434), .ZN(n3587) );
  NOR2_X1 U3681 ( .A1(n3586), .A2(n3588), .ZN(n3679) );
  NOR2_X1 U3682 ( .A1(n3683), .A2(n3684), .ZN(n3588) );
  INV_X1 U3683 ( .A(n3685), .ZN(n3684) );
  NAND2_X1 U3684 ( .A1(n3583), .A2(n3686), .ZN(n3685) );
  NAND2_X1 U3685 ( .A1(n3584), .A2(n3582), .ZN(n3686) );
  NOR2_X1 U3686 ( .A1(n3432), .A2(n2542), .ZN(n3583) );
  NOR2_X1 U3687 ( .A1(n3582), .A2(n3584), .ZN(n3683) );
  NOR2_X1 U3688 ( .A1(n3687), .A2(n3688), .ZN(n3584) );
  NOR2_X1 U3689 ( .A1(n3577), .A2(n3689), .ZN(n3688) );
  NOR2_X1 U3690 ( .A1(n3580), .A2(n3579), .ZN(n3689) );
  NAND2_X1 U3691 ( .A1(n3433), .A2(n2447), .ZN(n3577) );
  INV_X1 U3692 ( .A(n3432), .ZN(n3433) );
  INV_X1 U3693 ( .A(n3690), .ZN(n3687) );
  NAND2_X1 U3694 ( .A1(n3579), .A2(n3580), .ZN(n3690) );
  NAND2_X1 U3695 ( .A1(n3691), .A2(n3692), .ZN(n3580) );
  NAND2_X1 U3696 ( .A1(n3572), .A2(n3693), .ZN(n3692) );
  NAND2_X1 U3697 ( .A1(n2202), .A2(n3694), .ZN(n3693) );
  NAND2_X1 U3698 ( .A1(n3695), .A2(n2205), .ZN(n3694) );
  NAND2_X1 U3699 ( .A1(n3696), .A2(n3697), .ZN(n3691) );
  NAND2_X1 U3700 ( .A1(n2208), .A2(n3698), .ZN(n3697) );
  NAND2_X1 U3701 ( .A1(n2210), .A2(n3571), .ZN(n3698) );
  NOR3_X1 U3702 ( .A1(n3432), .A2(n2449), .A3(n3571), .ZN(n3579) );
  XOR2_X1 U3703 ( .A(d_5_), .B(c_5_), .Z(n3700) );
  XNOR2_X1 U3704 ( .A(n3701), .B(n3702), .ZN(n3582) );
  XNOR2_X1 U3705 ( .A(n3703), .B(n3704), .ZN(n3702) );
  XOR2_X1 U3706 ( .A(n3705), .B(n3706), .Z(n3586) );
  XNOR2_X1 U3707 ( .A(n3707), .B(n3708), .ZN(n3705) );
  XOR2_X1 U3708 ( .A(n3709), .B(n3710), .Z(n3590) );
  XNOR2_X1 U3709 ( .A(n3711), .B(n3712), .ZN(n3709) );
  XNOR2_X1 U3710 ( .A(n3713), .B(n3714), .ZN(n3594) );
  XNOR2_X1 U3711 ( .A(n3715), .B(n3716), .ZN(n3713) );
  XNOR2_X1 U3712 ( .A(n3717), .B(n3718), .ZN(n3533) );
  NAND2_X1 U3713 ( .A1(n3719), .A2(n3720), .ZN(n3717) );
  XNOR2_X1 U3714 ( .A(n3721), .B(n3722), .ZN(n3526) );
  XOR2_X1 U3715 ( .A(n3723), .B(n3724), .Z(n3721) );
  XNOR2_X1 U3716 ( .A(n3725), .B(n3726), .ZN(n3601) );
  XOR2_X1 U3717 ( .A(n3727), .B(n3728), .Z(n3725) );
  XNOR2_X1 U3718 ( .A(n3729), .B(n3730), .ZN(n3606) );
  XNOR2_X1 U3719 ( .A(n3731), .B(n3732), .ZN(n3730) );
  XOR2_X1 U3720 ( .A(n3733), .B(n3734), .Z(n3614) );
  XOR2_X1 U3721 ( .A(n3735), .B(n3736), .Z(n3734) );
  XOR2_X1 U3722 ( .A(n3737), .B(n3738), .Z(n3618) );
  XNOR2_X1 U3723 ( .A(n3739), .B(n3740), .ZN(n3738) );
  NAND2_X1 U3724 ( .A1(n2492), .A2(n3572), .ZN(n3740) );
  XOR2_X1 U3725 ( .A(n3496), .B(n3497), .Z(n3621) );
  XOR2_X1 U3726 ( .A(n3741), .B(n3742), .Z(n3497) );
  NOR2_X1 U3727 ( .A1(n2345), .A2(n3571), .ZN(n3742) );
  XOR2_X1 U3728 ( .A(n2194), .B(n2195), .Z(n2187) );
  XOR2_X1 U3729 ( .A(n3743), .B(n2321), .Z(n2195) );
  XNOR2_X1 U3730 ( .A(n3744), .B(n3745), .ZN(n2321) );
  XOR2_X1 U3731 ( .A(n3746), .B(n3747), .Z(n3744) );
  NOR2_X1 U3732 ( .A1(n3748), .A2(n2354), .ZN(n3747) );
  XNOR2_X1 U3733 ( .A(n2322), .B(n2319), .ZN(n3743) );
  NOR2_X1 U3734 ( .A1(n3695), .A2(n2345), .ZN(n2319) );
  NOR2_X1 U3735 ( .A1(n3749), .A2(n3750), .ZN(n2322) );
  INV_X1 U3736 ( .A(n3751), .ZN(n3750) );
  NAND2_X1 U3737 ( .A1(n3752), .A2(n3753), .ZN(n3751) );
  NAND2_X1 U3738 ( .A1(n3754), .A2(n3755), .ZN(n3753) );
  NOR2_X1 U3739 ( .A1(n3754), .A2(n3755), .ZN(n3749) );
  NOR2_X1 U3740 ( .A1(n3756), .A2(n3757), .ZN(n2194) );
  NOR3_X1 U3741 ( .A1(n2345), .A2(n3758), .A3(n3571), .ZN(n3757) );
  INV_X1 U3742 ( .A(n3759), .ZN(n3758) );
  NAND2_X1 U3743 ( .A1(n3741), .A2(n3496), .ZN(n3759) );
  NOR2_X1 U3744 ( .A1(n3496), .A2(n3741), .ZN(n3756) );
  NOR2_X1 U3745 ( .A1(n3760), .A2(n3761), .ZN(n3741) );
  INV_X1 U3746 ( .A(n3762), .ZN(n3761) );
  NAND3_X1 U3747 ( .A1(n3572), .A2(n3763), .A3(n2492), .ZN(n3762) );
  NAND2_X1 U3748 ( .A1(n3739), .A2(n3737), .ZN(n3763) );
  NOR2_X1 U3749 ( .A1(n3737), .A2(n3739), .ZN(n3760) );
  NOR2_X1 U3750 ( .A1(n3764), .A2(n3765), .ZN(n3739) );
  INV_X1 U3751 ( .A(n3766), .ZN(n3765) );
  NAND2_X1 U3752 ( .A1(n3633), .A2(n3767), .ZN(n3766) );
  NAND2_X1 U3753 ( .A1(n3632), .A2(n3631), .ZN(n3767) );
  NOR2_X1 U3754 ( .A1(n2497), .A2(n3571), .ZN(n3633) );
  NOR2_X1 U3755 ( .A1(n3631), .A2(n3632), .ZN(n3764) );
  NOR2_X1 U3756 ( .A1(n3768), .A2(n3769), .ZN(n3632) );
  INV_X1 U3757 ( .A(n3770), .ZN(n3769) );
  NAND2_X1 U3758 ( .A1(n3736), .A2(n3771), .ZN(n3770) );
  NAND2_X1 U3759 ( .A1(n3735), .A2(n3733), .ZN(n3771) );
  NOR2_X1 U3760 ( .A1(n2369), .A2(n3571), .ZN(n3736) );
  NOR2_X1 U3761 ( .A1(n3733), .A2(n3735), .ZN(n3768) );
  NOR2_X1 U3762 ( .A1(n3772), .A2(n3773), .ZN(n3735) );
  INV_X1 U3763 ( .A(n3774), .ZN(n3773) );
  NAND2_X1 U3764 ( .A1(n3645), .A2(n3775), .ZN(n3774) );
  NAND2_X1 U3765 ( .A1(n3644), .A2(n3643), .ZN(n3775) );
  NOR2_X1 U3766 ( .A1(n2508), .A2(n3571), .ZN(n3645) );
  NOR2_X1 U3767 ( .A1(n3643), .A2(n3644), .ZN(n3772) );
  NOR2_X1 U3768 ( .A1(n3776), .A2(n3777), .ZN(n3644) );
  INV_X1 U3769 ( .A(n3778), .ZN(n3777) );
  NAND2_X1 U3770 ( .A1(n3732), .A2(n3779), .ZN(n3778) );
  NAND2_X1 U3771 ( .A1(n3780), .A2(n3729), .ZN(n3779) );
  NOR2_X1 U3772 ( .A1(n2388), .A2(n3571), .ZN(n3732) );
  NOR2_X1 U3773 ( .A1(n3729), .A2(n3780), .ZN(n3776) );
  INV_X1 U3774 ( .A(n3731), .ZN(n3780) );
  NAND2_X1 U3775 ( .A1(n3781), .A2(n3782), .ZN(n3731) );
  NAND2_X1 U3776 ( .A1(n3728), .A2(n3783), .ZN(n3782) );
  INV_X1 U3777 ( .A(n3784), .ZN(n3783) );
  NOR2_X1 U3778 ( .A1(n3727), .A2(n3726), .ZN(n3784) );
  NOR2_X1 U3779 ( .A1(n2396), .A2(n3571), .ZN(n3728) );
  NAND2_X1 U3780 ( .A1(n3726), .A2(n3727), .ZN(n3781) );
  NAND2_X1 U3781 ( .A1(n3785), .A2(n3786), .ZN(n3727) );
  NAND2_X1 U3782 ( .A1(n3724), .A2(n3787), .ZN(n3786) );
  INV_X1 U3783 ( .A(n3788), .ZN(n3787) );
  NOR2_X1 U3784 ( .A1(n3723), .A2(n3722), .ZN(n3788) );
  NOR2_X1 U3785 ( .A1(n2406), .A2(n3571), .ZN(n3724) );
  NAND2_X1 U3786 ( .A1(n3722), .A2(n3723), .ZN(n3785) );
  NAND2_X1 U3787 ( .A1(n3719), .A2(n3789), .ZN(n3723) );
  NAND2_X1 U3788 ( .A1(n3718), .A2(n3720), .ZN(n3789) );
  NAND2_X1 U3789 ( .A1(n3790), .A2(n3791), .ZN(n3720) );
  NAND2_X1 U3790 ( .A1(n3572), .A2(n2414), .ZN(n3791) );
  INV_X1 U3791 ( .A(n3792), .ZN(n3790) );
  XNOR2_X1 U3792 ( .A(n3793), .B(n3794), .ZN(n3718) );
  XNOR2_X1 U3793 ( .A(n3795), .B(n3796), .ZN(n3793) );
  NAND2_X1 U3794 ( .A1(n2414), .A2(n3792), .ZN(n3719) );
  NAND2_X1 U3795 ( .A1(n3797), .A2(n3798), .ZN(n3792) );
  NAND3_X1 U3796 ( .A1(n3670), .A2(n3799), .A3(n3572), .ZN(n3798) );
  NAND2_X1 U3797 ( .A1(n3668), .A2(n3666), .ZN(n3799) );
  INV_X1 U3798 ( .A(n2424), .ZN(n3670) );
  INV_X1 U3799 ( .A(n3800), .ZN(n3797) );
  NOR2_X1 U3800 ( .A1(n3666), .A2(n3668), .ZN(n3800) );
  NOR2_X1 U3801 ( .A1(n3801), .A2(n3802), .ZN(n3668) );
  INV_X1 U3802 ( .A(n3803), .ZN(n3802) );
  NAND2_X1 U3803 ( .A1(n3716), .A2(n3804), .ZN(n3803) );
  NAND2_X1 U3804 ( .A1(n3715), .A2(n3714), .ZN(n3804) );
  NOR2_X1 U3805 ( .A1(n3571), .A2(n2429), .ZN(n3716) );
  NOR2_X1 U3806 ( .A1(n3714), .A2(n3715), .ZN(n3801) );
  NOR2_X1 U3807 ( .A1(n3805), .A2(n3806), .ZN(n3715) );
  INV_X1 U3808 ( .A(n3807), .ZN(n3806) );
  NAND2_X1 U3809 ( .A1(n3711), .A2(n3808), .ZN(n3807) );
  NAND2_X1 U3810 ( .A1(n3712), .A2(n3710), .ZN(n3808) );
  NOR2_X1 U3811 ( .A1(n3571), .A2(n2434), .ZN(n3711) );
  NOR2_X1 U3812 ( .A1(n3710), .A2(n3712), .ZN(n3805) );
  NOR2_X1 U3813 ( .A1(n3809), .A2(n3810), .ZN(n3712) );
  INV_X1 U3814 ( .A(n3811), .ZN(n3810) );
  NAND2_X1 U3815 ( .A1(n3707), .A2(n3812), .ZN(n3811) );
  NAND2_X1 U3816 ( .A1(n3708), .A2(n3706), .ZN(n3812) );
  NOR2_X1 U3817 ( .A1(n3571), .A2(n2542), .ZN(n3707) );
  NOR2_X1 U3818 ( .A1(n3706), .A2(n3708), .ZN(n3809) );
  NOR2_X1 U3819 ( .A1(n3813), .A2(n3814), .ZN(n3708) );
  NOR2_X1 U3820 ( .A1(n3701), .A2(n3815), .ZN(n3814) );
  NOR2_X1 U3821 ( .A1(n3704), .A2(n3703), .ZN(n3815) );
  NAND2_X1 U3822 ( .A1(n3572), .A2(n2447), .ZN(n3701) );
  INV_X1 U3823 ( .A(n3571), .ZN(n3572) );
  INV_X1 U3824 ( .A(n3816), .ZN(n3813) );
  NAND2_X1 U3825 ( .A1(n3703), .A2(n3704), .ZN(n3816) );
  NAND2_X1 U3826 ( .A1(n3817), .A2(n3818), .ZN(n3704) );
  NAND2_X1 U3827 ( .A1(n3696), .A2(n3819), .ZN(n3818) );
  NAND2_X1 U3828 ( .A1(n2202), .A2(n3820), .ZN(n3819) );
  NAND2_X1 U3829 ( .A1(n3748), .A2(n2205), .ZN(n3820) );
  NAND2_X1 U3830 ( .A1(n3821), .A2(n3822), .ZN(n3817) );
  NAND2_X1 U3831 ( .A1(n2208), .A2(n3823), .ZN(n3822) );
  NAND2_X1 U3832 ( .A1(n2210), .A2(n3695), .ZN(n3823) );
  NOR3_X1 U3833 ( .A1(n3571), .A2(n2449), .A3(n3695), .ZN(n3703) );
  XOR2_X1 U3834 ( .A(d_4_), .B(c_4_), .Z(n3825) );
  XOR2_X1 U3835 ( .A(n3826), .B(n3827), .Z(n3706) );
  XNOR2_X1 U3836 ( .A(n3828), .B(n3829), .ZN(n3827) );
  XOR2_X1 U3837 ( .A(n3830), .B(n3831), .Z(n3710) );
  XNOR2_X1 U3838 ( .A(n3832), .B(n3833), .ZN(n3830) );
  XOR2_X1 U3839 ( .A(n3834), .B(n3835), .Z(n3714) );
  XNOR2_X1 U3840 ( .A(n3836), .B(n3837), .ZN(n3834) );
  XOR2_X1 U3841 ( .A(n3838), .B(n3839), .Z(n3666) );
  XNOR2_X1 U3842 ( .A(n3840), .B(n3841), .ZN(n3838) );
  XNOR2_X1 U3843 ( .A(n3842), .B(n3843), .ZN(n3722) );
  XNOR2_X1 U3844 ( .A(n3844), .B(n3845), .ZN(n3842) );
  XNOR2_X1 U3845 ( .A(n3846), .B(n3847), .ZN(n3726) );
  XNOR2_X1 U3846 ( .A(n3848), .B(n3849), .ZN(n3846) );
  XOR2_X1 U3847 ( .A(n3850), .B(n3851), .Z(n3729) );
  XNOR2_X1 U3848 ( .A(n3852), .B(n3853), .ZN(n3850) );
  XOR2_X1 U3849 ( .A(n3854), .B(n3855), .Z(n3643) );
  XNOR2_X1 U3850 ( .A(n3856), .B(n3857), .ZN(n3854) );
  XOR2_X1 U3851 ( .A(n3858), .B(n3859), .Z(n3733) );
  XNOR2_X1 U3852 ( .A(n3860), .B(n3861), .ZN(n3858) );
  XOR2_X1 U3853 ( .A(n3862), .B(n3863), .Z(n3631) );
  XNOR2_X1 U3854 ( .A(n3864), .B(n3865), .ZN(n3862) );
  XOR2_X1 U3855 ( .A(n3866), .B(n3867), .Z(n3737) );
  XNOR2_X1 U3856 ( .A(n3868), .B(n3869), .ZN(n3866) );
  XOR2_X1 U3857 ( .A(n3870), .B(n3754), .Z(n3496) );
  XNOR2_X1 U3858 ( .A(n3871), .B(n3872), .ZN(n3754) );
  XOR2_X1 U3859 ( .A(n3873), .B(n3874), .Z(n3871) );
  XNOR2_X1 U3860 ( .A(n3755), .B(n3752), .ZN(n3870) );
  NOR2_X1 U3861 ( .A1(n2354), .A2(n3695), .ZN(n3752) );
  NOR2_X1 U3862 ( .A1(n3875), .A2(n3876), .ZN(n3755) );
  INV_X1 U3863 ( .A(n3877), .ZN(n3876) );
  NAND2_X1 U3864 ( .A1(n3869), .A2(n3878), .ZN(n3877) );
  NAND2_X1 U3865 ( .A1(n3867), .A2(n3868), .ZN(n3878) );
  NOR2_X1 U3866 ( .A1(n2497), .A2(n3695), .ZN(n3869) );
  NOR2_X1 U3867 ( .A1(n3867), .A2(n3868), .ZN(n3875) );
  NOR2_X1 U3868 ( .A1(n3879), .A2(n3880), .ZN(n3868) );
  INV_X1 U3869 ( .A(n3881), .ZN(n3880) );
  NAND2_X1 U3870 ( .A1(n3865), .A2(n3882), .ZN(n3881) );
  NAND2_X1 U3871 ( .A1(n3863), .A2(n3864), .ZN(n3882) );
  NOR2_X1 U3872 ( .A1(n2369), .A2(n3695), .ZN(n3865) );
  NOR2_X1 U3873 ( .A1(n3863), .A2(n3864), .ZN(n3879) );
  NOR2_X1 U3874 ( .A1(n3883), .A2(n3884), .ZN(n3864) );
  INV_X1 U3875 ( .A(n3885), .ZN(n3884) );
  NAND2_X1 U3876 ( .A1(n3861), .A2(n3886), .ZN(n3885) );
  NAND2_X1 U3877 ( .A1(n3859), .A2(n3860), .ZN(n3886) );
  NOR2_X1 U3878 ( .A1(n2508), .A2(n3695), .ZN(n3861) );
  NOR2_X1 U3879 ( .A1(n3859), .A2(n3860), .ZN(n3883) );
  NOR2_X1 U3880 ( .A1(n3887), .A2(n3888), .ZN(n3860) );
  INV_X1 U3881 ( .A(n3889), .ZN(n3888) );
  NAND2_X1 U3882 ( .A1(n3857), .A2(n3890), .ZN(n3889) );
  NAND2_X1 U3883 ( .A1(n3855), .A2(n3856), .ZN(n3890) );
  NOR2_X1 U3884 ( .A1(n2388), .A2(n3695), .ZN(n3857) );
  NOR2_X1 U3885 ( .A1(n3855), .A2(n3856), .ZN(n3887) );
  NOR2_X1 U3886 ( .A1(n3891), .A2(n3892), .ZN(n3856) );
  INV_X1 U3887 ( .A(n3893), .ZN(n3892) );
  NAND2_X1 U3888 ( .A1(n3853), .A2(n3894), .ZN(n3893) );
  NAND2_X1 U3889 ( .A1(n3851), .A2(n3852), .ZN(n3894) );
  NOR2_X1 U3890 ( .A1(n2396), .A2(n3695), .ZN(n3853) );
  NOR2_X1 U3891 ( .A1(n3851), .A2(n3852), .ZN(n3891) );
  NOR2_X1 U3892 ( .A1(n3895), .A2(n3896), .ZN(n3852) );
  INV_X1 U3893 ( .A(n3897), .ZN(n3896) );
  NAND2_X1 U3894 ( .A1(n3849), .A2(n3898), .ZN(n3897) );
  NAND2_X1 U3895 ( .A1(n3847), .A2(n3848), .ZN(n3898) );
  NOR2_X1 U3896 ( .A1(n2406), .A2(n3695), .ZN(n3849) );
  NOR2_X1 U3897 ( .A1(n3847), .A2(n3848), .ZN(n3895) );
  NOR2_X1 U3898 ( .A1(n3899), .A2(n3900), .ZN(n3848) );
  INV_X1 U3899 ( .A(n3901), .ZN(n3900) );
  NAND2_X1 U3900 ( .A1(n3845), .A2(n3902), .ZN(n3901) );
  NAND2_X1 U3901 ( .A1(n3843), .A2(n3844), .ZN(n3902) );
  NOR2_X1 U3902 ( .A1(n3695), .A2(n2525), .ZN(n3845) );
  NOR2_X1 U3903 ( .A1(n3843), .A2(n3844), .ZN(n3899) );
  NOR2_X1 U3904 ( .A1(n3903), .A2(n3904), .ZN(n3844) );
  INV_X1 U3905 ( .A(n3905), .ZN(n3904) );
  NAND2_X1 U3906 ( .A1(n3796), .A2(n3906), .ZN(n3905) );
  NAND2_X1 U3907 ( .A1(n3794), .A2(n3795), .ZN(n3906) );
  NOR2_X1 U3908 ( .A1(n3695), .A2(n2424), .ZN(n3796) );
  NOR2_X1 U3909 ( .A1(n3794), .A2(n3795), .ZN(n3903) );
  NOR2_X1 U3910 ( .A1(n3907), .A2(n3908), .ZN(n3795) );
  INV_X1 U3911 ( .A(n3909), .ZN(n3908) );
  NAND2_X1 U3912 ( .A1(n3841), .A2(n3910), .ZN(n3909) );
  NAND2_X1 U3913 ( .A1(n3839), .A2(n3840), .ZN(n3910) );
  NOR2_X1 U3914 ( .A1(n3695), .A2(n2429), .ZN(n3841) );
  NOR2_X1 U3915 ( .A1(n3839), .A2(n3840), .ZN(n3907) );
  NOR2_X1 U3916 ( .A1(n3911), .A2(n3912), .ZN(n3840) );
  INV_X1 U3917 ( .A(n3913), .ZN(n3912) );
  NAND2_X1 U3918 ( .A1(n3836), .A2(n3914), .ZN(n3913) );
  NAND2_X1 U3919 ( .A1(n3835), .A2(n3837), .ZN(n3914) );
  NOR2_X1 U3920 ( .A1(n3695), .A2(n2434), .ZN(n3836) );
  NOR2_X1 U3921 ( .A1(n3835), .A2(n3837), .ZN(n3911) );
  NOR2_X1 U3922 ( .A1(n3915), .A2(n3916), .ZN(n3837) );
  INV_X1 U3923 ( .A(n3917), .ZN(n3916) );
  NAND2_X1 U3924 ( .A1(n3832), .A2(n3918), .ZN(n3917) );
  NAND2_X1 U3925 ( .A1(n3831), .A2(n3833), .ZN(n3918) );
  NOR2_X1 U3926 ( .A1(n3695), .A2(n2542), .ZN(n3832) );
  NOR2_X1 U3927 ( .A1(n3831), .A2(n3833), .ZN(n3915) );
  NOR2_X1 U3928 ( .A1(n3919), .A2(n3920), .ZN(n3833) );
  INV_X1 U3929 ( .A(n3921), .ZN(n3920) );
  NAND2_X1 U3930 ( .A1(n3826), .A2(n3922), .ZN(n3921) );
  NAND2_X1 U3931 ( .A1(n3829), .A2(n3828), .ZN(n3922) );
  NOR2_X1 U3932 ( .A1(n3695), .A2(n3923), .ZN(n3826) );
  NOR2_X1 U3933 ( .A1(n3828), .A2(n3829), .ZN(n3919) );
  INV_X1 U3934 ( .A(n3924), .ZN(n3829) );
  NAND2_X1 U3935 ( .A1(n3925), .A2(n3926), .ZN(n3924) );
  NAND2_X1 U3936 ( .A1(n3821), .A2(n3927), .ZN(n3926) );
  NAND2_X1 U3937 ( .A1(n2202), .A2(n3928), .ZN(n3927) );
  NAND2_X1 U3938 ( .A1(n3929), .A2(n2205), .ZN(n3928) );
  NAND2_X1 U3939 ( .A1(n3930), .A2(n3931), .ZN(n3925) );
  NAND2_X1 U3940 ( .A1(n2208), .A2(n3932), .ZN(n3931) );
  NAND2_X1 U3941 ( .A1(n2210), .A2(n3748), .ZN(n3932) );
  NAND3_X1 U3942 ( .A1(n3696), .A2(n3933), .A3(n3821), .ZN(n3828) );
  INV_X1 U3943 ( .A(n3695), .ZN(n3696) );
  XOR2_X1 U3944 ( .A(d_3_), .B(c_3_), .Z(n3935) );
  XOR2_X1 U3945 ( .A(n3936), .B(n3937), .Z(n3831) );
  NAND2_X1 U3946 ( .A1(n3938), .A2(n3939), .ZN(n3936) );
  NAND2_X1 U3947 ( .A1(n3940), .A2(n3941), .ZN(n3939) );
  NAND2_X1 U3948 ( .A1(n3821), .A2(n2447), .ZN(n3941) );
  XOR2_X1 U3949 ( .A(n3942), .B(n3943), .Z(n3835) );
  NAND2_X1 U3950 ( .A1(n3944), .A2(n3945), .ZN(n3942) );
  XNOR2_X1 U3951 ( .A(n3946), .B(n3947), .ZN(n3839) );
  XOR2_X1 U3952 ( .A(n3948), .B(n3949), .Z(n3946) );
  NOR2_X1 U3953 ( .A1(n2434), .A2(n3748), .ZN(n3949) );
  XNOR2_X1 U3954 ( .A(n3950), .B(n3951), .ZN(n3794) );
  XOR2_X1 U3955 ( .A(n3952), .B(n3953), .Z(n3950) );
  XNOR2_X1 U3956 ( .A(n3954), .B(n3955), .ZN(n3843) );
  XOR2_X1 U3957 ( .A(n3956), .B(n3957), .Z(n3954) );
  XNOR2_X1 U3958 ( .A(n3958), .B(n3959), .ZN(n3847) );
  XOR2_X1 U3959 ( .A(n3960), .B(n3961), .Z(n3958) );
  XNOR2_X1 U3960 ( .A(n3962), .B(n3963), .ZN(n3851) );
  XOR2_X1 U3961 ( .A(n3964), .B(n3965), .Z(n3962) );
  XNOR2_X1 U3962 ( .A(n3966), .B(n3967), .ZN(n3855) );
  XOR2_X1 U3963 ( .A(n3968), .B(n3969), .Z(n3966) );
  XNOR2_X1 U3964 ( .A(n3970), .B(n3971), .ZN(n3859) );
  XOR2_X1 U3965 ( .A(n3972), .B(n3973), .Z(n3970) );
  XNOR2_X1 U3966 ( .A(n3974), .B(n3975), .ZN(n3863) );
  XOR2_X1 U3967 ( .A(n3976), .B(n3977), .Z(n3974) );
  XNOR2_X1 U3968 ( .A(n3978), .B(n3979), .ZN(n3867) );
  XOR2_X1 U3969 ( .A(n3980), .B(n3981), .Z(n3978) );
  NAND2_X1 U3970 ( .A1(n3982), .A2(n3983), .ZN(n2255) );
  NAND2_X1 U3971 ( .A1(n2304), .A2(n2306), .ZN(n3983) );
  NAND2_X1 U3972 ( .A1(n2315), .A2(n3984), .ZN(n2306) );
  NAND2_X1 U3973 ( .A1(n2314), .A2(n2316), .ZN(n3984) );
  NAND2_X1 U3974 ( .A1(n3985), .A2(n3986), .ZN(n2316) );
  NAND2_X1 U3975 ( .A1(n3821), .A2(n2303), .ZN(n3986) );
  INV_X1 U3976 ( .A(n3987), .ZN(n3985) );
  XOR2_X1 U3977 ( .A(n3988), .B(n3989), .Z(n2314) );
  NOR2_X1 U3978 ( .A1(n3990), .A2(n2497), .ZN(n3989) );
  XOR2_X1 U3979 ( .A(n3991), .B(n3992), .Z(n3988) );
  NAND2_X1 U3980 ( .A1(n2303), .A2(n3987), .ZN(n2315) );
  NAND2_X1 U3981 ( .A1(n3993), .A2(n3994), .ZN(n3987) );
  NAND3_X1 U3982 ( .A1(n3821), .A2(n3995), .A3(n2492), .ZN(n3994) );
  INV_X1 U3983 ( .A(n3996), .ZN(n3995) );
  NOR2_X1 U3984 ( .A1(n3746), .A2(n3745), .ZN(n3996) );
  NAND2_X1 U3985 ( .A1(n3745), .A2(n3746), .ZN(n3993) );
  NAND2_X1 U3986 ( .A1(n3997), .A2(n3998), .ZN(n3746) );
  NAND2_X1 U3987 ( .A1(n3874), .A2(n3999), .ZN(n3998) );
  INV_X1 U3988 ( .A(n4000), .ZN(n3999) );
  NOR2_X1 U3989 ( .A1(n3873), .A2(n3872), .ZN(n4000) );
  NOR2_X1 U3990 ( .A1(n2497), .A2(n3748), .ZN(n3874) );
  NAND2_X1 U3991 ( .A1(n3872), .A2(n3873), .ZN(n3997) );
  NAND2_X1 U3992 ( .A1(n4001), .A2(n4002), .ZN(n3873) );
  NAND2_X1 U3993 ( .A1(n3981), .A2(n4003), .ZN(n4002) );
  INV_X1 U3994 ( .A(n4004), .ZN(n4003) );
  NOR2_X1 U3995 ( .A1(n3980), .A2(n3979), .ZN(n4004) );
  NOR2_X1 U3996 ( .A1(n2369), .A2(n3748), .ZN(n3981) );
  NAND2_X1 U3997 ( .A1(n3979), .A2(n3980), .ZN(n4001) );
  NAND2_X1 U3998 ( .A1(n4005), .A2(n4006), .ZN(n3980) );
  NAND2_X1 U3999 ( .A1(n3977), .A2(n4007), .ZN(n4006) );
  INV_X1 U4000 ( .A(n4008), .ZN(n4007) );
  NOR2_X1 U4001 ( .A1(n3976), .A2(n3975), .ZN(n4008) );
  NOR2_X1 U4002 ( .A1(n2508), .A2(n3748), .ZN(n3977) );
  NAND2_X1 U4003 ( .A1(n3975), .A2(n3976), .ZN(n4005) );
  NAND2_X1 U4004 ( .A1(n4009), .A2(n4010), .ZN(n3976) );
  NAND2_X1 U4005 ( .A1(n3973), .A2(n4011), .ZN(n4010) );
  INV_X1 U4006 ( .A(n4012), .ZN(n4011) );
  NOR2_X1 U4007 ( .A1(n3972), .A2(n3971), .ZN(n4012) );
  NOR2_X1 U4008 ( .A1(n2388), .A2(n3748), .ZN(n3973) );
  NAND2_X1 U4009 ( .A1(n3971), .A2(n3972), .ZN(n4009) );
  NAND2_X1 U4010 ( .A1(n4013), .A2(n4014), .ZN(n3972) );
  NAND2_X1 U4011 ( .A1(n3969), .A2(n4015), .ZN(n4014) );
  INV_X1 U4012 ( .A(n4016), .ZN(n4015) );
  NOR2_X1 U4013 ( .A1(n3968), .A2(n3967), .ZN(n4016) );
  NOR2_X1 U4014 ( .A1(n2396), .A2(n3748), .ZN(n3969) );
  NAND2_X1 U4015 ( .A1(n3967), .A2(n3968), .ZN(n4013) );
  NAND2_X1 U4016 ( .A1(n4017), .A2(n4018), .ZN(n3968) );
  NAND2_X1 U4017 ( .A1(n3965), .A2(n4019), .ZN(n4018) );
  INV_X1 U4018 ( .A(n4020), .ZN(n4019) );
  NOR2_X1 U4019 ( .A1(n3964), .A2(n3963), .ZN(n4020) );
  NOR2_X1 U4020 ( .A1(n2406), .A2(n3748), .ZN(n3965) );
  NAND2_X1 U4021 ( .A1(n3963), .A2(n3964), .ZN(n4017) );
  NAND2_X1 U4022 ( .A1(n4021), .A2(n4022), .ZN(n3964) );
  NAND2_X1 U4023 ( .A1(n3961), .A2(n4023), .ZN(n4022) );
  INV_X1 U4024 ( .A(n4024), .ZN(n4023) );
  NOR2_X1 U4025 ( .A1(n3960), .A2(n3959), .ZN(n4024) );
  NOR2_X1 U4026 ( .A1(n3748), .A2(n2525), .ZN(n3961) );
  NAND2_X1 U4027 ( .A1(n3959), .A2(n3960), .ZN(n4021) );
  NAND2_X1 U4028 ( .A1(n4025), .A2(n4026), .ZN(n3960) );
  NAND2_X1 U4029 ( .A1(n3957), .A2(n4027), .ZN(n4026) );
  INV_X1 U4030 ( .A(n4028), .ZN(n4027) );
  NOR2_X1 U4031 ( .A1(n3956), .A2(n3955), .ZN(n4028) );
  NOR2_X1 U4032 ( .A1(n3748), .A2(n2424), .ZN(n3957) );
  NAND2_X1 U4033 ( .A1(n3955), .A2(n3956), .ZN(n4025) );
  NAND2_X1 U4034 ( .A1(n4029), .A2(n4030), .ZN(n3956) );
  NAND2_X1 U4035 ( .A1(n3953), .A2(n4031), .ZN(n4030) );
  INV_X1 U4036 ( .A(n4032), .ZN(n4031) );
  NOR2_X1 U4037 ( .A1(n3952), .A2(n3951), .ZN(n4032) );
  NOR2_X1 U4038 ( .A1(n3748), .A2(n2429), .ZN(n3953) );
  NAND2_X1 U4039 ( .A1(n3951), .A2(n3952), .ZN(n4029) );
  NAND2_X1 U4040 ( .A1(n4033), .A2(n4034), .ZN(n3952) );
  NAND3_X1 U4041 ( .A1(n4035), .A2(n4036), .A3(n3821), .ZN(n4034) );
  INV_X1 U4042 ( .A(n4037), .ZN(n4036) );
  NOR2_X1 U4043 ( .A1(n3948), .A2(n3947), .ZN(n4037) );
  NAND2_X1 U4044 ( .A1(n3947), .A2(n3948), .ZN(n4033) );
  NAND2_X1 U4045 ( .A1(n3944), .A2(n4038), .ZN(n3948) );
  NAND2_X1 U4046 ( .A1(n3943), .A2(n3945), .ZN(n4038) );
  NAND2_X1 U4047 ( .A1(n4039), .A2(n4040), .ZN(n3945) );
  NAND2_X1 U4048 ( .A1(n3821), .A2(n2438), .ZN(n4040) );
  INV_X1 U4049 ( .A(n4041), .ZN(n4039) );
  XNOR2_X1 U4050 ( .A(n4042), .B(n4043), .ZN(n3943) );
  XNOR2_X1 U4051 ( .A(n4044), .B(n4045), .ZN(n4043) );
  NAND2_X1 U4052 ( .A1(n2305), .A2(n2205), .ZN(n4042) );
  NAND2_X1 U4053 ( .A1(n2438), .A2(n4041), .ZN(n3944) );
  NAND2_X1 U4054 ( .A1(n3938), .A2(n4046), .ZN(n4041) );
  NAND2_X1 U4055 ( .A1(n3937), .A2(n4047), .ZN(n4046) );
  NAND2_X1 U4056 ( .A1(n3940), .A2(n3923), .ZN(n4047) );
  INV_X1 U4057 ( .A(n4048), .ZN(n3940) );
  NOR3_X1 U4058 ( .A1(n3748), .A2(n2449), .A3(n3929), .ZN(n3937) );
  INV_X1 U4059 ( .A(n3933), .ZN(n2449) );
  NAND3_X1 U4060 ( .A1(n2447), .A2(n4048), .A3(n3821), .ZN(n3938) );
  INV_X1 U4061 ( .A(n3748), .ZN(n3821) );
  XOR2_X1 U4062 ( .A(d_2_), .B(c_2_), .Z(n4050) );
  NAND2_X1 U4063 ( .A1(n4051), .A2(n4052), .ZN(n4048) );
  NAND2_X1 U4064 ( .A1(n3930), .A2(n4053), .ZN(n4052) );
  NAND2_X1 U4065 ( .A1(n2202), .A2(n4054), .ZN(n4053) );
  NAND2_X1 U4066 ( .A1(n3990), .A2(n2205), .ZN(n4054) );
  NAND2_X1 U4067 ( .A1(n2205), .A2(n2197), .ZN(n2202) );
  NAND2_X1 U4068 ( .A1(n2305), .A2(n4055), .ZN(n4051) );
  NAND2_X1 U4069 ( .A1(n2208), .A2(n4056), .ZN(n4055) );
  NAND2_X1 U4070 ( .A1(n2210), .A2(n3929), .ZN(n4056) );
  NAND2_X1 U4071 ( .A1(n4057), .A2(n2210), .ZN(n2208) );
  INV_X1 U4072 ( .A(n3923), .ZN(n2447) );
  XOR2_X1 U4073 ( .A(n4058), .B(n4059), .Z(n3947) );
  XNOR2_X1 U4074 ( .A(n4060), .B(n4061), .ZN(n4059) );
  NAND2_X1 U4075 ( .A1(n3930), .A2(n2438), .ZN(n4058) );
  XNOR2_X1 U4076 ( .A(n4062), .B(n4063), .ZN(n3951) );
  NAND2_X1 U4077 ( .A1(n4064), .A2(n4065), .ZN(n4062) );
  NAND2_X1 U4078 ( .A1(n4066), .A2(n4067), .ZN(n4065) );
  NAND2_X1 U4079 ( .A1(n3930), .A2(n4035), .ZN(n4066) );
  XNOR2_X1 U4080 ( .A(n4068), .B(n4069), .ZN(n3955) );
  XNOR2_X1 U4081 ( .A(n4070), .B(n4071), .ZN(n4069) );
  NOR2_X1 U4082 ( .A1(n3929), .A2(n2429), .ZN(n4068) );
  XOR2_X1 U4083 ( .A(n4072), .B(n4073), .Z(n3959) );
  NOR2_X1 U4084 ( .A1(n2424), .A2(n3929), .ZN(n4073) );
  XOR2_X1 U4085 ( .A(n4074), .B(n4075), .Z(n4072) );
  XOR2_X1 U4086 ( .A(n4076), .B(n4077), .Z(n3963) );
  NOR2_X1 U4087 ( .A1(n4078), .A2(n4079), .ZN(n4077) );
  INV_X1 U4088 ( .A(n4080), .ZN(n4079) );
  NOR2_X1 U4089 ( .A1(n4081), .A2(n4082), .ZN(n4078) );
  NOR2_X1 U4090 ( .A1(n2525), .A2(n3929), .ZN(n4082) );
  XOR2_X1 U4091 ( .A(n4083), .B(n4084), .Z(n3967) );
  XNOR2_X1 U4092 ( .A(n4085), .B(n4086), .ZN(n4084) );
  NAND2_X1 U4093 ( .A1(n2840), .A2(n3930), .ZN(n4083) );
  INV_X1 U4094 ( .A(n2406), .ZN(n2840) );
  XOR2_X1 U4095 ( .A(n4087), .B(n4088), .Z(n3971) );
  NOR2_X1 U4096 ( .A1(n4089), .A2(n4090), .ZN(n4088) );
  NOR2_X1 U4097 ( .A1(n4091), .A2(n4092), .ZN(n4089) );
  NOR2_X1 U4098 ( .A1(n3929), .A2(n2396), .ZN(n4092) );
  XOR2_X1 U4099 ( .A(n4093), .B(n4094), .Z(n3975) );
  NOR2_X1 U4100 ( .A1(n3929), .A2(n2388), .ZN(n4094) );
  XOR2_X1 U4101 ( .A(n4095), .B(n4096), .Z(n4093) );
  XOR2_X1 U4102 ( .A(n4097), .B(n4098), .Z(n3979) );
  NOR2_X1 U4103 ( .A1(n4099), .A2(n4100), .ZN(n4098) );
  INV_X1 U4104 ( .A(n4101), .ZN(n4100) );
  NOR2_X1 U4105 ( .A1(n4102), .A2(n4103), .ZN(n4099) );
  NOR2_X1 U4106 ( .A1(n3929), .A2(n2508), .ZN(n4103) );
  XOR2_X1 U4107 ( .A(n4104), .B(n4105), .Z(n3872) );
  XNOR2_X1 U4108 ( .A(n4106), .B(n4107), .ZN(n4105) );
  NAND2_X1 U4109 ( .A1(n2641), .A2(n3930), .ZN(n4104) );
  INV_X1 U4110 ( .A(n2369), .ZN(n2641) );
  XOR2_X1 U4111 ( .A(n4108), .B(n4109), .Z(n3745) );
  NOR2_X1 U4112 ( .A1(n4110), .A2(n4111), .ZN(n4109) );
  NOR2_X1 U4113 ( .A1(n4112), .A2(n4113), .ZN(n4110) );
  NOR2_X1 U4114 ( .A1(n3929), .A2(n2497), .ZN(n4113) );
  XOR2_X1 U4115 ( .A(n4114), .B(n4115), .Z(n2304) );
  NOR2_X1 U4116 ( .A1(n4116), .A2(n4117), .ZN(n4115) );
  INV_X1 U4117 ( .A(n4118), .ZN(n4117) );
  NOR2_X1 U4118 ( .A1(n4119), .A2(n4120), .ZN(n4116) );
  NOR2_X1 U4119 ( .A1(n2345), .A2(n3929), .ZN(n4120) );
  INV_X1 U4120 ( .A(n2303), .ZN(n2345) );
  XOR2_X1 U4121 ( .A(n2259), .B(n4121), .Z(n3982) );
  NAND2_X1 U4122 ( .A1(n2305), .A2(n2303), .ZN(n4121) );
  NAND2_X1 U4123 ( .A1(n4118), .A2(n4122), .ZN(n2259) );
  NAND2_X1 U4124 ( .A1(n4123), .A2(n4114), .ZN(n4122) );
  NAND2_X1 U4125 ( .A1(n4124), .A2(n4125), .ZN(n4114) );
  NAND3_X1 U4126 ( .A1(n2305), .A2(n4126), .A3(n2358), .ZN(n4125) );
  INV_X1 U4127 ( .A(n2497), .ZN(n2358) );
  NAND2_X1 U4128 ( .A1(n3991), .A2(n3992), .ZN(n4126) );
  INV_X1 U4129 ( .A(n4127), .ZN(n4124) );
  NOR2_X1 U4130 ( .A1(n3992), .A2(n3991), .ZN(n4127) );
  NOR2_X1 U4131 ( .A1(n4111), .A2(n4128), .ZN(n3991) );
  INV_X1 U4132 ( .A(n4129), .ZN(n4128) );
  NAND2_X1 U4133 ( .A1(n4130), .A2(n4108), .ZN(n4129) );
  NAND2_X1 U4134 ( .A1(n4131), .A2(n4132), .ZN(n4108) );
  INV_X1 U4135 ( .A(n4133), .ZN(n4132) );
  NOR3_X1 U4136 ( .A1(n3929), .A2(n4134), .A3(n2369), .ZN(n4133) );
  NOR2_X1 U4137 ( .A1(n4107), .A2(n4106), .ZN(n4134) );
  NAND2_X1 U4138 ( .A1(n4106), .A2(n4107), .ZN(n4131) );
  NAND2_X1 U4139 ( .A1(n4101), .A2(n4135), .ZN(n4107) );
  NAND2_X1 U4140 ( .A1(n4136), .A2(n4097), .ZN(n4135) );
  NAND2_X1 U4141 ( .A1(n4137), .A2(n4138), .ZN(n4097) );
  NAND3_X1 U4142 ( .A1(n3930), .A2(n4139), .A3(n2593), .ZN(n4138) );
  INV_X1 U4143 ( .A(n2388), .ZN(n2593) );
  NAND2_X1 U4144 ( .A1(n4095), .A2(n4096), .ZN(n4139) );
  INV_X1 U4145 ( .A(n4140), .ZN(n4137) );
  NOR2_X1 U4146 ( .A1(n4096), .A2(n4095), .ZN(n4140) );
  NOR2_X1 U4147 ( .A1(n4090), .A2(n4141), .ZN(n4095) );
  INV_X1 U4148 ( .A(n4142), .ZN(n4141) );
  NAND2_X1 U4149 ( .A1(n4143), .A2(n4087), .ZN(n4142) );
  NAND2_X1 U4150 ( .A1(n4144), .A2(n4145), .ZN(n4087) );
  INV_X1 U4151 ( .A(n4146), .ZN(n4145) );
  NOR3_X1 U4152 ( .A1(n3929), .A2(n4147), .A3(n2406), .ZN(n4146) );
  NOR2_X1 U4153 ( .A1(n4086), .A2(n4085), .ZN(n4147) );
  NAND2_X1 U4154 ( .A1(n4085), .A2(n4086), .ZN(n4144) );
  NAND2_X1 U4155 ( .A1(n4080), .A2(n4148), .ZN(n4086) );
  NAND2_X1 U4156 ( .A1(n4149), .A2(n4076), .ZN(n4148) );
  NAND2_X1 U4157 ( .A1(n4150), .A2(n4151), .ZN(n4076) );
  INV_X1 U4158 ( .A(n4152), .ZN(n4151) );
  NOR3_X1 U4159 ( .A1(n2424), .A2(n4153), .A3(n3929), .ZN(n4152) );
  NOR2_X1 U4160 ( .A1(n4074), .A2(n4075), .ZN(n4153) );
  NAND2_X1 U4161 ( .A1(n4075), .A2(n4074), .ZN(n4150) );
  NAND2_X1 U4162 ( .A1(n4154), .A2(n4155), .ZN(n4074) );
  INV_X1 U4163 ( .A(n4156), .ZN(n4155) );
  NOR3_X1 U4164 ( .A1(n2429), .A2(n4157), .A3(n3929), .ZN(n4156) );
  NOR2_X1 U4165 ( .A1(n4071), .A2(n4070), .ZN(n4157) );
  NAND2_X1 U4166 ( .A1(n4070), .A2(n4071), .ZN(n4154) );
  NAND2_X1 U4167 ( .A1(n4064), .A2(n4158), .ZN(n4071) );
  NAND2_X1 U4168 ( .A1(n4159), .A2(n4063), .ZN(n4158) );
  NAND2_X1 U4169 ( .A1(n4160), .A2(n4161), .ZN(n4063) );
  NAND3_X1 U4170 ( .A1(n2438), .A2(n4162), .A3(n3930), .ZN(n4161) );
  INV_X1 U4171 ( .A(n4163), .ZN(n4162) );
  NOR2_X1 U4172 ( .A1(n4061), .A2(n4060), .ZN(n4163) );
  NAND2_X1 U4173 ( .A1(n4060), .A2(n4061), .ZN(n4160) );
  NAND2_X1 U4174 ( .A1(n4045), .A2(n4164), .ZN(n4061) );
  NAND3_X1 U4175 ( .A1(n2305), .A2(n2205), .A3(n4044), .ZN(n4164) );
  NOR2_X1 U4176 ( .A1(n3929), .A2(n3923), .ZN(n4044) );
  NAND3_X1 U4177 ( .A1(n3930), .A2(n3933), .A3(n2305), .ZN(n4045) );
  NOR2_X1 U4178 ( .A1(n2197), .A2(n4057), .ZN(n3933) );
  INV_X1 U4179 ( .A(n2205), .ZN(n4057) );
  XOR2_X1 U4180 ( .A(b_14_), .B(a_14_), .Z(n4166) );
  INV_X1 U4181 ( .A(n2210), .ZN(n2197) );
  NOR2_X1 U4182 ( .A1(b_15_), .A2(a_15_), .ZN(n4167) );
  NOR2_X1 U4183 ( .A1(n3990), .A2(n3923), .ZN(n4060) );
  XNOR2_X1 U4184 ( .A(n4168), .B(n4169), .ZN(n3923) );
  XOR2_X1 U4185 ( .A(b_13_), .B(a_13_), .Z(n4169) );
  NAND2_X1 U4186 ( .A1(n2434), .A2(n4067), .ZN(n4159) );
  NAND3_X1 U4187 ( .A1(n3930), .A2(n4035), .A3(n4170), .ZN(n4064) );
  INV_X1 U4188 ( .A(n4067), .ZN(n4170) );
  NAND2_X1 U4189 ( .A1(n2305), .A2(n2438), .ZN(n4067) );
  INV_X1 U4190 ( .A(n2542), .ZN(n2438) );
  XNOR2_X1 U4191 ( .A(a_12_), .B(b_12_), .ZN(n4171) );
  NOR2_X1 U4192 ( .A1(n3990), .A2(n2434), .ZN(n4070) );
  INV_X1 U4193 ( .A(n4035), .ZN(n2434) );
  XOR2_X1 U4194 ( .A(n4173), .B(n4174), .Z(n4035) );
  XOR2_X1 U4195 ( .A(b_11_), .B(a_11_), .Z(n4174) );
  NOR2_X1 U4196 ( .A1(n3990), .A2(n2429), .ZN(n4075) );
  XOR2_X1 U4197 ( .A(b_10_), .B(a_10_), .Z(n4176) );
  INV_X1 U4198 ( .A(n4177), .ZN(n4149) );
  NOR2_X1 U4199 ( .A1(n2414), .A2(n4081), .ZN(n4177) );
  NAND3_X1 U4200 ( .A1(n2414), .A2(n3930), .A3(n4081), .ZN(n4080) );
  NOR2_X1 U4201 ( .A1(n3990), .A2(n2424), .ZN(n4081) );
  XOR2_X1 U4202 ( .A(b_9_), .B(a_9_), .Z(n4179) );
  INV_X1 U4203 ( .A(n2525), .ZN(n2414) );
  NOR2_X1 U4204 ( .A1(n3990), .A2(n2525), .ZN(n4085) );
  XOR2_X1 U4205 ( .A(b_8_), .B(a_8_), .Z(n4181) );
  NAND2_X1 U4206 ( .A1(n2396), .A2(n4182), .ZN(n4143) );
  NOR3_X1 U4207 ( .A1(n2396), .A2(n3929), .A3(n4182), .ZN(n4090) );
  INV_X1 U4208 ( .A(n4091), .ZN(n4182) );
  NOR2_X1 U4209 ( .A1(n3990), .A2(n2406), .ZN(n4091) );
  XOR2_X1 U4210 ( .A(b_7_), .B(a_7_), .Z(n4184) );
  NAND2_X1 U4211 ( .A1(n2654), .A2(n2305), .ZN(n4096) );
  INV_X1 U4212 ( .A(n3990), .ZN(n2305) );
  INV_X1 U4213 ( .A(n2396), .ZN(n2654) );
  XOR2_X1 U4214 ( .A(b_6_), .B(a_6_), .Z(n4186) );
  INV_X1 U4215 ( .A(n4187), .ZN(n4136) );
  NOR2_X1 U4216 ( .A1(n2378), .A2(n4102), .ZN(n4187) );
  NAND3_X1 U4217 ( .A1(n2378), .A2(n3930), .A3(n4102), .ZN(n4101) );
  NOR2_X1 U4218 ( .A1(n2388), .A2(n3990), .ZN(n4102) );
  XOR2_X1 U4219 ( .A(b_5_), .B(a_5_), .Z(n4189) );
  INV_X1 U4220 ( .A(n2508), .ZN(n2378) );
  NOR2_X1 U4221 ( .A1(n2508), .A2(n3990), .ZN(n4106) );
  XOR2_X1 U4222 ( .A(b_4_), .B(a_4_), .Z(n4191) );
  NAND2_X1 U4223 ( .A1(n2497), .A2(n4192), .ZN(n4130) );
  NOR3_X1 U4224 ( .A1(n2497), .A2(n3929), .A3(n4192), .ZN(n4111) );
  INV_X1 U4225 ( .A(n4112), .ZN(n4192) );
  NOR2_X1 U4226 ( .A1(n2369), .A2(n3990), .ZN(n4112) );
  XOR2_X1 U4227 ( .A(b_3_), .B(a_3_), .Z(n4194) );
  XOR2_X1 U4228 ( .A(b_2_), .B(a_2_), .Z(n4196) );
  NAND2_X1 U4229 ( .A1(n2492), .A2(n3930), .ZN(n3992) );
  INV_X1 U4230 ( .A(n2354), .ZN(n2492) );
  INV_X1 U4231 ( .A(n4197), .ZN(n4123) );
  NOR2_X1 U4232 ( .A1(n2303), .A2(n4119), .ZN(n4197) );
  NAND3_X1 U4233 ( .A1(n3930), .A2(n2303), .A3(n4119), .ZN(n4118) );
  NOR2_X1 U4234 ( .A1(n2354), .A2(n3990), .ZN(n4119) );
  XOR2_X1 U4235 ( .A(d_0_), .B(c_0_), .Z(n4199) );
  NAND2_X1 U4236 ( .A1(n4200), .A2(n4201), .ZN(n4198) );
  NAND2_X1 U4237 ( .A1(d_1_), .A2(n4202), .ZN(n4201) );
  INV_X1 U4238 ( .A(n4203), .ZN(n4202) );
  NOR2_X1 U4239 ( .A1(n4204), .A2(c_1_), .ZN(n4203) );
  NAND2_X1 U4240 ( .A1(c_1_), .A2(n4204), .ZN(n4200) );
  XNOR2_X1 U4241 ( .A(n4205), .B(n4206), .ZN(n2354) );
  XNOR2_X1 U4242 ( .A(n4207), .B(a_1_), .ZN(n4206) );
  XOR2_X1 U4243 ( .A(b_0_), .B(a_0_), .Z(n4209) );
  NAND2_X1 U4244 ( .A1(n4210), .A2(n4211), .ZN(n4208) );
  NAND2_X1 U4245 ( .A1(n4212), .A2(n4207), .ZN(n4211) );
  INV_X1 U4246 ( .A(b_1_), .ZN(n4207) );
  NAND2_X1 U4247 ( .A1(a_1_), .A2(n4205), .ZN(n4212) );
  INV_X1 U4248 ( .A(n4213), .ZN(n4210) );
  NOR2_X1 U4249 ( .A1(n4205), .A2(a_1_), .ZN(n4213) );
  NAND2_X1 U4250 ( .A1(n4214), .A2(n4215), .ZN(n4205) );
  NAND2_X1 U4251 ( .A1(b_2_), .A2(n4216), .ZN(n4215) );
  INV_X1 U4252 ( .A(n4217), .ZN(n4216) );
  NOR2_X1 U4253 ( .A1(n4195), .A2(a_2_), .ZN(n4217) );
  NAND2_X1 U4254 ( .A1(a_2_), .A2(n4195), .ZN(n4214) );
  NAND2_X1 U4255 ( .A1(n4218), .A2(n4219), .ZN(n4195) );
  NAND2_X1 U4256 ( .A1(b_3_), .A2(n4220), .ZN(n4219) );
  INV_X1 U4257 ( .A(n4221), .ZN(n4220) );
  NOR2_X1 U4258 ( .A1(n4193), .A2(a_3_), .ZN(n4221) );
  NAND2_X1 U4259 ( .A1(a_3_), .A2(n4193), .ZN(n4218) );
  NAND2_X1 U4260 ( .A1(n4222), .A2(n4223), .ZN(n4193) );
  NAND2_X1 U4261 ( .A1(b_4_), .A2(n4224), .ZN(n4223) );
  INV_X1 U4262 ( .A(n4225), .ZN(n4224) );
  NOR2_X1 U4263 ( .A1(n4190), .A2(a_4_), .ZN(n4225) );
  NAND2_X1 U4264 ( .A1(a_4_), .A2(n4190), .ZN(n4222) );
  NAND2_X1 U4265 ( .A1(n4226), .A2(n4227), .ZN(n4190) );
  NAND2_X1 U4266 ( .A1(b_5_), .A2(n4228), .ZN(n4227) );
  INV_X1 U4267 ( .A(n4229), .ZN(n4228) );
  NOR2_X1 U4268 ( .A1(n4188), .A2(a_5_), .ZN(n4229) );
  NAND2_X1 U4269 ( .A1(a_5_), .A2(n4188), .ZN(n4226) );
  NAND2_X1 U4270 ( .A1(n4230), .A2(n4231), .ZN(n4188) );
  NAND2_X1 U4271 ( .A1(b_6_), .A2(n4232), .ZN(n4231) );
  INV_X1 U4272 ( .A(n4233), .ZN(n4232) );
  NOR2_X1 U4273 ( .A1(n4185), .A2(a_6_), .ZN(n4233) );
  NAND2_X1 U4274 ( .A1(a_6_), .A2(n4185), .ZN(n4230) );
  NAND2_X1 U4275 ( .A1(n4234), .A2(n4235), .ZN(n4185) );
  NAND2_X1 U4276 ( .A1(b_7_), .A2(n4236), .ZN(n4235) );
  INV_X1 U4277 ( .A(n4237), .ZN(n4236) );
  NOR2_X1 U4278 ( .A1(n4183), .A2(a_7_), .ZN(n4237) );
  NAND2_X1 U4279 ( .A1(a_7_), .A2(n4183), .ZN(n4234) );
  NAND2_X1 U4280 ( .A1(n4238), .A2(n4239), .ZN(n4183) );
  NAND2_X1 U4281 ( .A1(b_8_), .A2(n4240), .ZN(n4239) );
  INV_X1 U4282 ( .A(n4241), .ZN(n4240) );
  NOR2_X1 U4283 ( .A1(n4180), .A2(a_8_), .ZN(n4241) );
  NAND2_X1 U4284 ( .A1(a_8_), .A2(n4180), .ZN(n4238) );
  NAND2_X1 U4285 ( .A1(n4242), .A2(n4243), .ZN(n4180) );
  NAND2_X1 U4286 ( .A1(b_9_), .A2(n4244), .ZN(n4243) );
  INV_X1 U4287 ( .A(n4245), .ZN(n4244) );
  NOR2_X1 U4288 ( .A1(n4178), .A2(a_9_), .ZN(n4245) );
  NAND2_X1 U4289 ( .A1(a_9_), .A2(n4178), .ZN(n4242) );
  NAND2_X1 U4290 ( .A1(n4246), .A2(n4247), .ZN(n4178) );
  NAND2_X1 U4291 ( .A1(b_10_), .A2(n4248), .ZN(n4247) );
  INV_X1 U4292 ( .A(n4249), .ZN(n4248) );
  NOR2_X1 U4293 ( .A1(n4175), .A2(a_10_), .ZN(n4249) );
  NAND2_X1 U4294 ( .A1(a_10_), .A2(n4175), .ZN(n4246) );
  NAND2_X1 U4295 ( .A1(n4250), .A2(n4251), .ZN(n4175) );
  NAND2_X1 U4296 ( .A1(b_11_), .A2(n4252), .ZN(n4251) );
  INV_X1 U4297 ( .A(n4253), .ZN(n4252) );
  NOR2_X1 U4298 ( .A1(n4173), .A2(a_11_), .ZN(n4253) );
  NAND2_X1 U4299 ( .A1(a_11_), .A2(n4173), .ZN(n4250) );
  NAND2_X1 U4300 ( .A1(n4254), .A2(n4255), .ZN(n4173) );
  NAND2_X1 U4301 ( .A1(b_12_), .A2(n4256), .ZN(n4255) );
  INV_X1 U4302 ( .A(n4257), .ZN(n4256) );
  NOR2_X1 U4303 ( .A1(n4172), .A2(a_12_), .ZN(n4257) );
  NAND2_X1 U4304 ( .A1(a_12_), .A2(n4172), .ZN(n4254) );
  NAND2_X1 U4305 ( .A1(n4258), .A2(n4259), .ZN(n4172) );
  NAND2_X1 U4306 ( .A1(b_13_), .A2(n4260), .ZN(n4259) );
  INV_X1 U4307 ( .A(n4261), .ZN(n4260) );
  NOR2_X1 U4308 ( .A1(n4168), .A2(a_13_), .ZN(n4261) );
  NAND2_X1 U4309 ( .A1(a_13_), .A2(n4168), .ZN(n4258) );
  NAND2_X1 U4310 ( .A1(n4262), .A2(n4263), .ZN(n4168) );
  NAND2_X1 U4311 ( .A1(b_14_), .A2(n4264), .ZN(n4263) );
  NAND2_X1 U4312 ( .A1(n4265), .A2(n4266), .ZN(n4264) );
  INV_X1 U4313 ( .A(a_14_), .ZN(n4265) );
  NAND2_X1 U4314 ( .A1(a_14_), .A2(n4165), .ZN(n4262) );
  INV_X1 U4315 ( .A(n4266), .ZN(n4165) );
  NAND2_X1 U4316 ( .A1(b_15_), .A2(a_15_), .ZN(n4266) );
  INV_X1 U4317 ( .A(n3929), .ZN(n3930) );
  XOR2_X1 U4318 ( .A(d_1_), .B(c_1_), .Z(n4267) );
  NAND2_X1 U4319 ( .A1(n4268), .A2(n4269), .ZN(n4204) );
  NAND2_X1 U4320 ( .A1(d_2_), .A2(n4270), .ZN(n4269) );
  INV_X1 U4321 ( .A(n4271), .ZN(n4270) );
  NOR2_X1 U4322 ( .A1(n4049), .A2(c_2_), .ZN(n4271) );
  NAND2_X1 U4323 ( .A1(c_2_), .A2(n4049), .ZN(n4268) );
  NAND2_X1 U4324 ( .A1(n4272), .A2(n4273), .ZN(n4049) );
  NAND2_X1 U4325 ( .A1(d_3_), .A2(n4274), .ZN(n4273) );
  INV_X1 U4326 ( .A(n4275), .ZN(n4274) );
  NOR2_X1 U4327 ( .A1(n3934), .A2(c_3_), .ZN(n4275) );
  NAND2_X1 U4328 ( .A1(c_3_), .A2(n3934), .ZN(n4272) );
  NAND2_X1 U4329 ( .A1(n4276), .A2(n4277), .ZN(n3934) );
  NAND2_X1 U4330 ( .A1(d_4_), .A2(n4278), .ZN(n4277) );
  INV_X1 U4331 ( .A(n4279), .ZN(n4278) );
  NOR2_X1 U4332 ( .A1(n3824), .A2(c_4_), .ZN(n4279) );
  NAND2_X1 U4333 ( .A1(c_4_), .A2(n3824), .ZN(n4276) );
  NAND2_X1 U4334 ( .A1(n4280), .A2(n4281), .ZN(n3824) );
  NAND2_X1 U4335 ( .A1(d_5_), .A2(n4282), .ZN(n4281) );
  INV_X1 U4336 ( .A(n4283), .ZN(n4282) );
  NOR2_X1 U4337 ( .A1(n3699), .A2(c_5_), .ZN(n4283) );
  NAND2_X1 U4338 ( .A1(c_5_), .A2(n3699), .ZN(n4280) );
  NAND2_X1 U4339 ( .A1(n4284), .A2(n4285), .ZN(n3699) );
  NAND2_X1 U4340 ( .A1(d_6_), .A2(n4286), .ZN(n4285) );
  INV_X1 U4341 ( .A(n4287), .ZN(n4286) );
  NOR2_X1 U4342 ( .A1(n3575), .A2(c_6_), .ZN(n4287) );
  NAND2_X1 U4343 ( .A1(c_6_), .A2(n3575), .ZN(n4284) );
  NAND2_X1 U4344 ( .A1(n4288), .A2(n4289), .ZN(n3575) );
  NAND2_X1 U4345 ( .A1(d_7_), .A2(n4290), .ZN(n4289) );
  INV_X1 U4346 ( .A(n4291), .ZN(n4290) );
  NOR2_X1 U4347 ( .A1(n3436), .A2(c_7_), .ZN(n4291) );
  NAND2_X1 U4348 ( .A1(c_7_), .A2(n3436), .ZN(n4288) );
  NAND2_X1 U4349 ( .A1(n4292), .A2(n4293), .ZN(n3436) );
  NAND2_X1 U4350 ( .A1(d_8_), .A2(n4294), .ZN(n4293) );
  INV_X1 U4351 ( .A(n4295), .ZN(n4294) );
  NOR2_X1 U4352 ( .A1(n3321), .A2(c_8_), .ZN(n4295) );
  NAND2_X1 U4353 ( .A1(c_8_), .A2(n3321), .ZN(n4292) );
  NAND2_X1 U4354 ( .A1(n4296), .A2(n4297), .ZN(n3321) );
  NAND2_X1 U4355 ( .A1(d_9_), .A2(n4298), .ZN(n4297) );
  INV_X1 U4356 ( .A(n4299), .ZN(n4298) );
  NOR2_X1 U4357 ( .A1(n3189), .A2(c_9_), .ZN(n4299) );
  NAND2_X1 U4358 ( .A1(c_9_), .A2(n3189), .ZN(n4296) );
  NAND2_X1 U4359 ( .A1(n4300), .A2(n4301), .ZN(n3189) );
  NAND2_X1 U4360 ( .A1(d_10_), .A2(n4302), .ZN(n4301) );
  INV_X1 U4361 ( .A(n4303), .ZN(n4302) );
  NOR2_X1 U4362 ( .A1(n3066), .A2(c_10_), .ZN(n4303) );
  NAND2_X1 U4363 ( .A1(c_10_), .A2(n3066), .ZN(n4300) );
  NAND2_X1 U4364 ( .A1(n4304), .A2(n4305), .ZN(n3066) );
  NAND2_X1 U4365 ( .A1(d_11_), .A2(n4306), .ZN(n4305) );
  INV_X1 U4366 ( .A(n4307), .ZN(n4306) );
  NOR2_X1 U4367 ( .A1(n2941), .A2(c_11_), .ZN(n4307) );
  NAND2_X1 U4368 ( .A1(c_11_), .A2(n2941), .ZN(n4304) );
  NAND2_X1 U4369 ( .A1(n4308), .A2(n4309), .ZN(n2941) );
  NAND2_X1 U4370 ( .A1(d_12_), .A2(n4310), .ZN(n4309) );
  INV_X1 U4371 ( .A(n4311), .ZN(n4310) );
  NOR2_X1 U4372 ( .A1(n2810), .A2(c_12_), .ZN(n4311) );
  NAND2_X1 U4373 ( .A1(c_12_), .A2(n2810), .ZN(n4308) );
  NAND2_X1 U4374 ( .A1(n4312), .A2(n4313), .ZN(n2810) );
  NAND2_X1 U4375 ( .A1(d_13_), .A2(n4314), .ZN(n4313) );
  INV_X1 U4376 ( .A(n4315), .ZN(n4314) );
  NOR2_X1 U4377 ( .A1(n2692), .A2(c_13_), .ZN(n4315) );
  NAND2_X1 U4378 ( .A1(c_13_), .A2(n2692), .ZN(n4312) );
  NAND2_X1 U4379 ( .A1(n4316), .A2(n4317), .ZN(n2692) );
  NAND3_X1 U4380 ( .A1(c_15_), .A2(n4318), .A3(d_15_), .ZN(n4317) );
  INV_X1 U4381 ( .A(n4319), .ZN(n4318) );
  NOR2_X1 U4382 ( .A1(d_14_), .A2(c_14_), .ZN(n4319) );
  NAND2_X1 U4383 ( .A1(d_14_), .A2(c_14_), .ZN(n4316) );
endmodule

