module add_mul_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, 
        b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, 
        b_15_, operation, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874;

  AND2_X1 U1962 ( .A1(n1930), .A2(operation), .ZN(Result_9_) );
  XOR2_X1 U1963 ( .A(n1931), .B(n1932), .Z(n1930) );
  AND2_X1 U1964 ( .A1(operation), .A2(n1933), .ZN(Result_8_) );
  XOR2_X1 U1965 ( .A(n1934), .B(n1935), .Z(n1933) );
  AND2_X1 U1966 ( .A1(operation), .A2(n1936), .ZN(Result_7_) );
  XOR2_X1 U1967 ( .A(n1937), .B(n1938), .Z(n1936) );
  AND2_X1 U1968 ( .A1(operation), .A2(n1939), .ZN(Result_6_) );
  XOR2_X1 U1969 ( .A(n1940), .B(n1941), .Z(n1939) );
  AND2_X1 U1970 ( .A1(operation), .A2(n1942), .ZN(Result_5_) );
  XOR2_X1 U1971 ( .A(n1943), .B(n1944), .Z(n1942) );
  AND2_X1 U1972 ( .A1(operation), .A2(n1945), .ZN(Result_4_) );
  XOR2_X1 U1973 ( .A(n1946), .B(n1947), .Z(n1945) );
  AND2_X1 U1974 ( .A1(operation), .A2(n1948), .ZN(Result_3_) );
  XOR2_X1 U1975 ( .A(n1949), .B(n1950), .Z(n1948) );
  OR2_X1 U1976 ( .A1(n1951), .A2(n1952), .ZN(Result_31_) );
  AND2_X1 U1977 ( .A1(n1953), .A2(operation), .ZN(n1952) );
  AND2_X1 U1978 ( .A1(n1954), .A2(n1955), .ZN(n1951) );
  XOR2_X1 U1979 ( .A(b_15_), .B(a_15_), .Z(n1954) );
  OR2_X1 U1980 ( .A1(n1956), .A2(n1957), .ZN(Result_30_) );
  AND2_X1 U1981 ( .A1(n1958), .A2(n1955), .ZN(n1957) );
  XOR2_X1 U1982 ( .A(n1953), .B(n1959), .Z(n1958) );
  XOR2_X1 U1983 ( .A(b_14_), .B(a_14_), .Z(n1959) );
  AND2_X1 U1984 ( .A1(operation), .A2(n1960), .ZN(n1956) );
  OR2_X1 U1985 ( .A1(n1961), .A2(n1962), .ZN(n1960) );
  AND2_X1 U1986 ( .A1(b_15_), .A2(n1963), .ZN(n1962) );
  OR2_X1 U1987 ( .A1(n1964), .A2(n1965), .ZN(n1963) );
  AND2_X1 U1988 ( .A1(a_14_), .A2(n1966), .ZN(n1964) );
  AND2_X1 U1989 ( .A1(b_14_), .A2(n1967), .ZN(n1961) );
  OR2_X1 U1990 ( .A1(n1968), .A2(n1969), .ZN(n1967) );
  AND2_X1 U1991 ( .A1(a_15_), .A2(n1970), .ZN(n1968) );
  AND2_X1 U1992 ( .A1(operation), .A2(n1971), .ZN(Result_2_) );
  XOR2_X1 U1993 ( .A(n1972), .B(n1973), .Z(n1971) );
  OR2_X1 U1994 ( .A1(n1974), .A2(n1975), .ZN(Result_29_) );
  AND2_X1 U1995 ( .A1(n1976), .A2(operation), .ZN(n1975) );
  XOR2_X1 U1996 ( .A(n1977), .B(n1978), .Z(n1976) );
  XOR2_X1 U1997 ( .A(n1979), .B(n1980), .Z(n1978) );
  AND2_X1 U1998 ( .A1(n1981), .A2(n1955), .ZN(n1974) );
  OR2_X1 U1999 ( .A1(n1982), .A2(n1983), .ZN(n1981) );
  OR2_X1 U2000 ( .A1(n1984), .A2(n1985), .ZN(n1983) );
  AND2_X1 U2001 ( .A1(n1986), .A2(n1987), .ZN(n1985) );
  XOR2_X1 U2002 ( .A(n1988), .B(n1989), .Z(n1986) );
  AND2_X1 U2003 ( .A1(n1990), .A2(b_13_), .ZN(n1984) );
  AND2_X1 U2004 ( .A1(n1988), .A2(n1989), .ZN(n1990) );
  INV_X1 U2005 ( .A(n1991), .ZN(n1982) );
  OR2_X1 U2006 ( .A1(n1992), .A2(n1988), .ZN(n1991) );
  OR2_X1 U2007 ( .A1(n1993), .A2(n1994), .ZN(Result_28_) );
  AND2_X1 U2008 ( .A1(n1995), .A2(operation), .ZN(n1994) );
  XNOR2_X1 U2009 ( .A(n1996), .B(n1997), .ZN(n1995) );
  XOR2_X1 U2010 ( .A(n1998), .B(n1999), .Z(n1997) );
  AND2_X1 U2011 ( .A1(n2000), .A2(n1955), .ZN(n1993) );
  XOR2_X1 U2012 ( .A(n2001), .B(n2002), .Z(n2000) );
  OR2_X1 U2013 ( .A1(n2003), .A2(n2004), .ZN(n2002) );
  INV_X1 U2014 ( .A(n2005), .ZN(n2003) );
  OR2_X1 U2015 ( .A1(n2006), .A2(n2007), .ZN(Result_27_) );
  AND2_X1 U2016 ( .A1(n2008), .A2(operation), .ZN(n2007) );
  XNOR2_X1 U2017 ( .A(n2009), .B(n2010), .ZN(n2008) );
  XOR2_X1 U2018 ( .A(n2011), .B(n2012), .Z(n2010) );
  AND2_X1 U2019 ( .A1(n2013), .A2(n1955), .ZN(n2006) );
  OR2_X1 U2020 ( .A1(n2014), .A2(n2015), .ZN(n2013) );
  OR2_X1 U2021 ( .A1(n2016), .A2(n2017), .ZN(n2015) );
  AND2_X1 U2022 ( .A1(n2018), .A2(n2019), .ZN(n2017) );
  XOR2_X1 U2023 ( .A(n2020), .B(n2021), .Z(n2018) );
  AND2_X1 U2024 ( .A1(n2022), .A2(b_11_), .ZN(n2016) );
  AND2_X1 U2025 ( .A1(n2021), .A2(n2020), .ZN(n2022) );
  INV_X1 U2026 ( .A(n2023), .ZN(n2014) );
  OR2_X1 U2027 ( .A1(n2021), .A2(n2024), .ZN(n2023) );
  OR2_X1 U2028 ( .A1(n2025), .A2(n2026), .ZN(Result_26_) );
  AND2_X1 U2029 ( .A1(n2027), .A2(operation), .ZN(n2026) );
  XNOR2_X1 U2030 ( .A(n2028), .B(n2029), .ZN(n2027) );
  XOR2_X1 U2031 ( .A(n2030), .B(n2031), .Z(n2029) );
  AND2_X1 U2032 ( .A1(n2032), .A2(n1955), .ZN(n2025) );
  XOR2_X1 U2033 ( .A(n2033), .B(n2034), .Z(n2032) );
  OR2_X1 U2034 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
  INV_X1 U2035 ( .A(n2037), .ZN(n2035) );
  OR2_X1 U2036 ( .A1(n2038), .A2(n2039), .ZN(Result_25_) );
  AND2_X1 U2037 ( .A1(n2040), .A2(operation), .ZN(n2039) );
  XNOR2_X1 U2038 ( .A(n2041), .B(n2042), .ZN(n2040) );
  XOR2_X1 U2039 ( .A(n2043), .B(n2044), .Z(n2042) );
  AND2_X1 U2040 ( .A1(n2045), .A2(n1955), .ZN(n2038) );
  OR2_X1 U2041 ( .A1(n2046), .A2(n2047), .ZN(n2045) );
  OR2_X1 U2042 ( .A1(n2048), .A2(n2049), .ZN(n2047) );
  AND2_X1 U2043 ( .A1(n2050), .A2(n2051), .ZN(n2049) );
  XOR2_X1 U2044 ( .A(n2052), .B(n2053), .Z(n2050) );
  AND2_X1 U2045 ( .A1(n2054), .A2(b_9_), .ZN(n2048) );
  AND2_X1 U2046 ( .A1(n2053), .A2(n2052), .ZN(n2054) );
  INV_X1 U2047 ( .A(n2055), .ZN(n2046) );
  OR2_X1 U2048 ( .A1(n2053), .A2(n2056), .ZN(n2055) );
  OR2_X1 U2049 ( .A1(n2057), .A2(n2058), .ZN(Result_24_) );
  AND2_X1 U2050 ( .A1(n2059), .A2(operation), .ZN(n2058) );
  XNOR2_X1 U2051 ( .A(n2060), .B(n2061), .ZN(n2059) );
  XOR2_X1 U2052 ( .A(n2062), .B(n2063), .Z(n2061) );
  AND2_X1 U2053 ( .A1(n2064), .A2(n1955), .ZN(n2057) );
  XOR2_X1 U2054 ( .A(n2065), .B(n2066), .Z(n2064) );
  OR2_X1 U2055 ( .A1(n2067), .A2(n2068), .ZN(n2066) );
  INV_X1 U2056 ( .A(n2069), .ZN(n2068) );
  OR2_X1 U2057 ( .A1(n2070), .A2(n2071), .ZN(Result_23_) );
  AND2_X1 U2058 ( .A1(n2072), .A2(operation), .ZN(n2071) );
  XNOR2_X1 U2059 ( .A(n2073), .B(n2074), .ZN(n2072) );
  XOR2_X1 U2060 ( .A(n2075), .B(n2076), .Z(n2074) );
  AND2_X1 U2061 ( .A1(n2077), .A2(n1955), .ZN(n2070) );
  OR2_X1 U2062 ( .A1(n2078), .A2(n2079), .ZN(n2077) );
  OR2_X1 U2063 ( .A1(n2080), .A2(n2081), .ZN(n2079) );
  AND2_X1 U2064 ( .A1(n2082), .A2(n2083), .ZN(n2081) );
  XOR2_X1 U2065 ( .A(n2084), .B(n2085), .Z(n2082) );
  AND2_X1 U2066 ( .A1(n2086), .A2(b_7_), .ZN(n2080) );
  AND2_X1 U2067 ( .A1(n2085), .A2(n2084), .ZN(n2086) );
  INV_X1 U2068 ( .A(n2087), .ZN(n2078) );
  OR2_X1 U2069 ( .A1(n2085), .A2(n2088), .ZN(n2087) );
  OR2_X1 U2070 ( .A1(n2089), .A2(n2090), .ZN(Result_22_) );
  AND2_X1 U2071 ( .A1(n2091), .A2(operation), .ZN(n2090) );
  XNOR2_X1 U2072 ( .A(n2092), .B(n2093), .ZN(n2091) );
  XOR2_X1 U2073 ( .A(n2094), .B(n2095), .Z(n2093) );
  AND2_X1 U2074 ( .A1(n2096), .A2(n1955), .ZN(n2089) );
  XOR2_X1 U2075 ( .A(n2097), .B(n2098), .Z(n2096) );
  OR2_X1 U2076 ( .A1(n2099), .A2(n2100), .ZN(n2098) );
  INV_X1 U2077 ( .A(n2101), .ZN(n2100) );
  OR2_X1 U2078 ( .A1(n2102), .A2(n2103), .ZN(Result_21_) );
  AND2_X1 U2079 ( .A1(n2104), .A2(operation), .ZN(n2103) );
  XNOR2_X1 U2080 ( .A(n2105), .B(n2106), .ZN(n2104) );
  XOR2_X1 U2081 ( .A(n2107), .B(n2108), .Z(n2106) );
  AND2_X1 U2082 ( .A1(n2109), .A2(n1955), .ZN(n2102) );
  OR2_X1 U2083 ( .A1(n2110), .A2(n2111), .ZN(n2109) );
  OR2_X1 U2084 ( .A1(n2112), .A2(n2113), .ZN(n2111) );
  AND2_X1 U2085 ( .A1(n2114), .A2(n2115), .ZN(n2113) );
  XOR2_X1 U2086 ( .A(n2116), .B(n2117), .Z(n2114) );
  AND2_X1 U2087 ( .A1(n2118), .A2(b_5_), .ZN(n2112) );
  AND2_X1 U2088 ( .A1(n2117), .A2(n2116), .ZN(n2118) );
  INV_X1 U2089 ( .A(n2119), .ZN(n2110) );
  OR2_X1 U2090 ( .A1(n2117), .A2(n2120), .ZN(n2119) );
  OR2_X1 U2091 ( .A1(n2121), .A2(n2122), .ZN(Result_20_) );
  AND2_X1 U2092 ( .A1(n2123), .A2(operation), .ZN(n2122) );
  XNOR2_X1 U2093 ( .A(n2124), .B(n2125), .ZN(n2123) );
  XOR2_X1 U2094 ( .A(n2126), .B(n2127), .Z(n2125) );
  AND2_X1 U2095 ( .A1(n2128), .A2(n1955), .ZN(n2121) );
  XOR2_X1 U2096 ( .A(n2129), .B(n2130), .Z(n2128) );
  OR2_X1 U2097 ( .A1(n2131), .A2(n2132), .ZN(n2130) );
  INV_X1 U2098 ( .A(n2133), .ZN(n2132) );
  AND2_X1 U2099 ( .A1(operation), .A2(n2134), .ZN(Result_1_) );
  XOR2_X1 U2100 ( .A(n2135), .B(n2136), .Z(n2134) );
  OR2_X1 U2101 ( .A1(n2137), .A2(n2138), .ZN(n2136) );
  INV_X1 U2102 ( .A(n2139), .ZN(n2138) );
  AND2_X1 U2103 ( .A1(n2140), .A2(n2141), .ZN(n2137) );
  OR2_X1 U2104 ( .A1(n2142), .A2(n2143), .ZN(n2141) );
  OR2_X1 U2105 ( .A1(n2144), .A2(n2145), .ZN(Result_19_) );
  AND2_X1 U2106 ( .A1(n2146), .A2(operation), .ZN(n2145) );
  XNOR2_X1 U2107 ( .A(n2147), .B(n2148), .ZN(n2146) );
  XOR2_X1 U2108 ( .A(n2149), .B(n2150), .Z(n2148) );
  AND2_X1 U2109 ( .A1(n2151), .A2(n1955), .ZN(n2144) );
  OR2_X1 U2110 ( .A1(n2152), .A2(n2153), .ZN(n2151) );
  OR2_X1 U2111 ( .A1(n2154), .A2(n2155), .ZN(n2153) );
  AND2_X1 U2112 ( .A1(n2156), .A2(n2157), .ZN(n2155) );
  XOR2_X1 U2113 ( .A(n2158), .B(n2159), .Z(n2156) );
  AND2_X1 U2114 ( .A1(n2160), .A2(b_3_), .ZN(n2154) );
  AND2_X1 U2115 ( .A1(n2159), .A2(n2158), .ZN(n2160) );
  INV_X1 U2116 ( .A(n2161), .ZN(n2152) );
  OR2_X1 U2117 ( .A1(n2159), .A2(n2162), .ZN(n2161) );
  OR2_X1 U2118 ( .A1(n2163), .A2(n2164), .ZN(Result_18_) );
  AND2_X1 U2119 ( .A1(n2165), .A2(operation), .ZN(n2164) );
  XNOR2_X1 U2120 ( .A(n2166), .B(n2167), .ZN(n2165) );
  XOR2_X1 U2121 ( .A(n2168), .B(n2169), .Z(n2167) );
  AND2_X1 U2122 ( .A1(n2170), .A2(n1955), .ZN(n2163) );
  XOR2_X1 U2123 ( .A(n2171), .B(n2172), .Z(n2170) );
  OR2_X1 U2124 ( .A1(n2173), .A2(n2174), .ZN(n2172) );
  INV_X1 U2125 ( .A(n2175), .ZN(n2174) );
  OR2_X1 U2126 ( .A1(n2176), .A2(n2177), .ZN(Result_17_) );
  AND2_X1 U2127 ( .A1(n2178), .A2(operation), .ZN(n2177) );
  XNOR2_X1 U2128 ( .A(n2179), .B(n2180), .ZN(n2178) );
  XOR2_X1 U2129 ( .A(n2181), .B(n2182), .Z(n2180) );
  AND2_X1 U2130 ( .A1(n2183), .A2(n1955), .ZN(n2176) );
  OR2_X1 U2131 ( .A1(n2184), .A2(n2185), .ZN(n2183) );
  OR2_X1 U2132 ( .A1(n2186), .A2(n2187), .ZN(n2185) );
  AND2_X1 U2133 ( .A1(n2188), .A2(n2189), .ZN(n2187) );
  XOR2_X1 U2134 ( .A(n2190), .B(n2191), .Z(n2188) );
  AND2_X1 U2135 ( .A1(n2192), .A2(b_1_), .ZN(n2186) );
  AND2_X1 U2136 ( .A1(n2191), .A2(n2190), .ZN(n2192) );
  INV_X1 U2137 ( .A(n2193), .ZN(n2184) );
  OR2_X1 U2138 ( .A1(n2191), .A2(n2194), .ZN(n2193) );
  OR2_X1 U2139 ( .A1(n2195), .A2(n2196), .ZN(Result_16_) );
  AND2_X1 U2140 ( .A1(n2197), .A2(operation), .ZN(n2196) );
  XNOR2_X1 U2141 ( .A(n2198), .B(n2199), .ZN(n2197) );
  XOR2_X1 U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  AND2_X1 U2143 ( .A1(n2202), .A2(n1955), .ZN(n2195) );
  XOR2_X1 U2144 ( .A(n2203), .B(n2204), .Z(n2202) );
  XOR2_X1 U2145 ( .A(n2205), .B(b_0_), .Z(n2204) );
  OR2_X1 U2146 ( .A1(n2206), .A2(n2207), .ZN(n2203) );
  AND2_X1 U2147 ( .A1(n2190), .A2(n2189), .ZN(n2207) );
  AND2_X1 U2148 ( .A1(n2191), .A2(n2194), .ZN(n2206) );
  OR2_X1 U2149 ( .A1(n2208), .A2(n2173), .ZN(n2191) );
  AND2_X1 U2150 ( .A1(n2209), .A2(n2210), .ZN(n2173) );
  AND2_X1 U2151 ( .A1(n2171), .A2(n2175), .ZN(n2208) );
  OR2_X1 U2152 ( .A1(n2211), .A2(n2212), .ZN(n2171) );
  AND2_X1 U2153 ( .A1(n2158), .A2(n2157), .ZN(n2212) );
  AND2_X1 U2154 ( .A1(n2159), .A2(n2162), .ZN(n2211) );
  OR2_X1 U2155 ( .A1(n2213), .A2(n2131), .ZN(n2159) );
  AND2_X1 U2156 ( .A1(n2214), .A2(n2215), .ZN(n2131) );
  AND2_X1 U2157 ( .A1(n2129), .A2(n2133), .ZN(n2213) );
  OR2_X1 U2158 ( .A1(n2216), .A2(n2217), .ZN(n2129) );
  AND2_X1 U2159 ( .A1(n2116), .A2(n2115), .ZN(n2217) );
  AND2_X1 U2160 ( .A1(n2117), .A2(n2120), .ZN(n2216) );
  OR2_X1 U2161 ( .A1(n2218), .A2(n2099), .ZN(n2117) );
  AND2_X1 U2162 ( .A1(n2219), .A2(n2220), .ZN(n2099) );
  AND2_X1 U2163 ( .A1(n2097), .A2(n2101), .ZN(n2218) );
  OR2_X1 U2164 ( .A1(n2221), .A2(n2222), .ZN(n2097) );
  AND2_X1 U2165 ( .A1(n2084), .A2(n2083), .ZN(n2222) );
  AND2_X1 U2166 ( .A1(n2085), .A2(n2088), .ZN(n2221) );
  OR2_X1 U2167 ( .A1(n2223), .A2(n2067), .ZN(n2085) );
  AND2_X1 U2168 ( .A1(n2224), .A2(n2225), .ZN(n2067) );
  AND2_X1 U2169 ( .A1(n2065), .A2(n2069), .ZN(n2223) );
  OR2_X1 U2170 ( .A1(n2226), .A2(n2227), .ZN(n2065) );
  AND2_X1 U2171 ( .A1(n2052), .A2(n2051), .ZN(n2227) );
  AND2_X1 U2172 ( .A1(n2053), .A2(n2056), .ZN(n2226) );
  OR2_X1 U2173 ( .A1(n2228), .A2(n2036), .ZN(n2053) );
  AND2_X1 U2174 ( .A1(n2229), .A2(n2230), .ZN(n2036) );
  AND2_X1 U2175 ( .A1(n2033), .A2(n2037), .ZN(n2228) );
  OR2_X1 U2176 ( .A1(n2231), .A2(n2232), .ZN(n2033) );
  AND2_X1 U2177 ( .A1(n2020), .A2(n2019), .ZN(n2232) );
  AND2_X1 U2178 ( .A1(n2021), .A2(n2024), .ZN(n2231) );
  OR2_X1 U2179 ( .A1(n2233), .A2(n2004), .ZN(n2021) );
  AND2_X1 U2180 ( .A1(n2234), .A2(n2235), .ZN(n2004) );
  AND2_X1 U2181 ( .A1(n2001), .A2(n2005), .ZN(n2233) );
  OR2_X1 U2182 ( .A1(n2236), .A2(n2237), .ZN(n2001) );
  AND2_X1 U2183 ( .A1(n1989), .A2(n1987), .ZN(n2237) );
  AND2_X1 U2184 ( .A1(n1988), .A2(n1992), .ZN(n2236) );
  AND2_X1 U2185 ( .A1(n2238), .A2(n2239), .ZN(n1988) );
  OR2_X1 U2186 ( .A1(n1966), .A2(n2240), .ZN(n2239) );
  INV_X1 U2187 ( .A(n2241), .ZN(n2240) );
  OR2_X1 U2188 ( .A1(a_14_), .A2(n1953), .ZN(n2241) );
  AND2_X1 U2189 ( .A1(a_15_), .A2(b_15_), .ZN(n1953) );
  AND2_X1 U2190 ( .A1(operation), .A2(n2242), .ZN(Result_15_) );
  XOR2_X1 U2191 ( .A(n2243), .B(n2244), .Z(n2242) );
  AND2_X1 U2192 ( .A1(n2245), .A2(operation), .ZN(Result_14_) );
  AND2_X1 U2193 ( .A1(n2246), .A2(n2247), .ZN(n2245) );
  INV_X1 U2194 ( .A(n2248), .ZN(n2247) );
  OR2_X1 U2195 ( .A1(n2249), .A2(n2250), .ZN(n2246) );
  AND2_X1 U2196 ( .A1(n2243), .A2(n2244), .ZN(n2249) );
  AND2_X1 U2197 ( .A1(operation), .A2(n2251), .ZN(Result_13_) );
  XNOR2_X1 U2198 ( .A(n2248), .B(n2252), .ZN(n2251) );
  OR2_X1 U2199 ( .A1(n2253), .A2(n2254), .ZN(n2252) );
  AND2_X1 U2200 ( .A1(n2255), .A2(n2256), .ZN(n2254) );
  AND2_X1 U2201 ( .A1(n2257), .A2(operation), .ZN(Result_12_) );
  XOR2_X1 U2202 ( .A(n2258), .B(n2259), .Z(n2257) );
  AND2_X1 U2203 ( .A1(n2260), .A2(n2261), .ZN(n2259) );
  OR2_X1 U2204 ( .A1(n2262), .A2(n2263), .ZN(n2261) );
  INV_X1 U2205 ( .A(n2264), .ZN(n2260) );
  AND2_X1 U2206 ( .A1(n2265), .A2(operation), .ZN(Result_11_) );
  XOR2_X1 U2207 ( .A(n2266), .B(n2267), .Z(n2265) );
  AND2_X1 U2208 ( .A1(n2268), .A2(n2269), .ZN(n2267) );
  OR2_X1 U2209 ( .A1(n2270), .A2(n2271), .ZN(n2269) );
  AND2_X1 U2210 ( .A1(n2272), .A2(n2273), .ZN(n2270) );
  INV_X1 U2211 ( .A(n2274), .ZN(n2268) );
  AND2_X1 U2212 ( .A1(n2275), .A2(operation), .ZN(Result_10_) );
  XOR2_X1 U2213 ( .A(n2276), .B(n2277), .Z(n2275) );
  AND2_X1 U2214 ( .A1(n2278), .A2(n2279), .ZN(n2277) );
  OR2_X1 U2215 ( .A1(n2280), .A2(n2281), .ZN(n2279) );
  INV_X1 U2216 ( .A(n2282), .ZN(n2278) );
  INV_X1 U2217 ( .A(n2283), .ZN(Result_0_) );
  OR2_X1 U2218 ( .A1(n1955), .A2(n2284), .ZN(n2283) );
  AND2_X1 U2219 ( .A1(n2285), .A2(n2286), .ZN(n2284) );
  AND2_X1 U2220 ( .A1(n2139), .A2(n2287), .ZN(n2286) );
  OR2_X1 U2221 ( .A1(n2135), .A2(n2140), .ZN(n2287) );
  OR2_X1 U2222 ( .A1(n1973), .A2(n1972), .ZN(n2135) );
  XNOR2_X1 U2223 ( .A(n2142), .B(n2143), .ZN(n1972) );
  AND2_X1 U2224 ( .A1(n2288), .A2(n2289), .ZN(n1973) );
  OR2_X1 U2225 ( .A1(n1950), .A2(n1949), .ZN(n2289) );
  OR2_X1 U2226 ( .A1(n2290), .A2(n2291), .ZN(n1949) );
  INV_X1 U2227 ( .A(n2288), .ZN(n2291) );
  AND2_X1 U2228 ( .A1(n2292), .A2(n2293), .ZN(n2290) );
  AND2_X1 U2229 ( .A1(n2294), .A2(n2295), .ZN(n1950) );
  OR2_X1 U2230 ( .A1(n1947), .A2(n1946), .ZN(n2294) );
  OR2_X1 U2231 ( .A1(n2296), .A2(n2297), .ZN(n1946) );
  INV_X1 U2232 ( .A(n2295), .ZN(n2297) );
  OR2_X1 U2233 ( .A1(n2298), .A2(n2299), .ZN(n2295) );
  AND2_X1 U2234 ( .A1(n2298), .A2(n2299), .ZN(n2296) );
  OR2_X1 U2235 ( .A1(n2300), .A2(n2301), .ZN(n2299) );
  AND2_X1 U2236 ( .A1(n2302), .A2(n2303), .ZN(n2301) );
  AND2_X1 U2237 ( .A1(n2304), .A2(n2305), .ZN(n2300) );
  OR2_X1 U2238 ( .A1(n2303), .A2(n2302), .ZN(n2305) );
  XOR2_X1 U2239 ( .A(n2306), .B(n2307), .Z(n2298) );
  XOR2_X1 U2240 ( .A(n2308), .B(n2309), .Z(n2307) );
  AND2_X1 U2241 ( .A1(n2310), .A2(n2311), .ZN(n1947) );
  OR2_X1 U2242 ( .A1(n1944), .A2(n1943), .ZN(n2311) );
  OR2_X1 U2243 ( .A1(n2312), .A2(n2313), .ZN(n1943) );
  INV_X1 U2244 ( .A(n2310), .ZN(n2313) );
  AND2_X1 U2245 ( .A1(n2314), .A2(n2315), .ZN(n2312) );
  AND2_X1 U2246 ( .A1(n2316), .A2(n2317), .ZN(n1944) );
  OR2_X1 U2247 ( .A1(n1941), .A2(n1940), .ZN(n2316) );
  OR2_X1 U2248 ( .A1(n2318), .A2(n2319), .ZN(n1940) );
  INV_X1 U2249 ( .A(n2317), .ZN(n2319) );
  OR2_X1 U2250 ( .A1(n2320), .A2(n2321), .ZN(n2317) );
  AND2_X1 U2251 ( .A1(n2320), .A2(n2321), .ZN(n2318) );
  OR2_X1 U2252 ( .A1(n2322), .A2(n2323), .ZN(n2321) );
  AND2_X1 U2253 ( .A1(n2324), .A2(n2325), .ZN(n2323) );
  AND2_X1 U2254 ( .A1(n2326), .A2(n2327), .ZN(n2322) );
  OR2_X1 U2255 ( .A1(n2325), .A2(n2324), .ZN(n2327) );
  XOR2_X1 U2256 ( .A(n2328), .B(n2329), .Z(n2320) );
  XOR2_X1 U2257 ( .A(n2330), .B(n2331), .Z(n2329) );
  AND2_X1 U2258 ( .A1(n2332), .A2(n2333), .ZN(n1941) );
  OR2_X1 U2259 ( .A1(n1938), .A2(n1937), .ZN(n2333) );
  OR2_X1 U2260 ( .A1(n2334), .A2(n2335), .ZN(n1937) );
  INV_X1 U2261 ( .A(n2332), .ZN(n2335) );
  AND2_X1 U2262 ( .A1(n2336), .A2(n2337), .ZN(n2334) );
  AND2_X1 U2263 ( .A1(n2338), .A2(n2339), .ZN(n1938) );
  OR2_X1 U2264 ( .A1(n1935), .A2(n1934), .ZN(n2338) );
  OR2_X1 U2265 ( .A1(n2340), .A2(n2341), .ZN(n1934) );
  INV_X1 U2266 ( .A(n2339), .ZN(n2341) );
  OR2_X1 U2267 ( .A1(n2342), .A2(n2343), .ZN(n2339) );
  AND2_X1 U2268 ( .A1(n2342), .A2(n2343), .ZN(n2340) );
  OR2_X1 U2269 ( .A1(n2344), .A2(n2345), .ZN(n2343) );
  AND2_X1 U2270 ( .A1(n2346), .A2(n2347), .ZN(n2345) );
  AND2_X1 U2271 ( .A1(n2348), .A2(n2349), .ZN(n2344) );
  OR2_X1 U2272 ( .A1(n2347), .A2(n2346), .ZN(n2349) );
  XOR2_X1 U2273 ( .A(n2350), .B(n2351), .Z(n2342) );
  XOR2_X1 U2274 ( .A(n2352), .B(n2353), .Z(n2351) );
  AND2_X1 U2275 ( .A1(n2354), .A2(n2355), .ZN(n1935) );
  OR2_X1 U2276 ( .A1(n1932), .A2(n1931), .ZN(n2355) );
  OR2_X1 U2277 ( .A1(n2356), .A2(n2357), .ZN(n1931) );
  INV_X1 U2278 ( .A(n2354), .ZN(n2357) );
  AND2_X1 U2279 ( .A1(n2358), .A2(n2359), .ZN(n2356) );
  AND2_X1 U2280 ( .A1(n2360), .A2(n2361), .ZN(n1932) );
  INV_X1 U2281 ( .A(n2362), .ZN(n2360) );
  OR2_X1 U2282 ( .A1(n2363), .A2(n2282), .ZN(n2362) );
  AND2_X1 U2283 ( .A1(n2280), .A2(n2281), .ZN(n2282) );
  AND2_X1 U2284 ( .A1(n2364), .A2(n2365), .ZN(n2281) );
  AND2_X1 U2285 ( .A1(n2280), .A2(n2276), .ZN(n2363) );
  OR2_X1 U2286 ( .A1(n2366), .A2(n2274), .ZN(n2276) );
  AND2_X1 U2287 ( .A1(n2272), .A2(n2367), .ZN(n2274) );
  AND2_X1 U2288 ( .A1(n2273), .A2(n2271), .ZN(n2367) );
  AND2_X1 U2289 ( .A1(n2271), .A2(n2266), .ZN(n2366) );
  OR2_X1 U2290 ( .A1(n2368), .A2(n2264), .ZN(n2266) );
  AND2_X1 U2291 ( .A1(n2263), .A2(n2262), .ZN(n2264) );
  AND2_X1 U2292 ( .A1(n2263), .A2(n2258), .ZN(n2368) );
  OR2_X1 U2293 ( .A1(n2369), .A2(n2253), .ZN(n2258) );
  INV_X1 U2294 ( .A(n2370), .ZN(n2253) );
  OR2_X1 U2295 ( .A1(n2255), .A2(n2256), .ZN(n2370) );
  OR2_X1 U2296 ( .A1(n2371), .A2(n2372), .ZN(n2256) );
  AND2_X1 U2297 ( .A1(n2248), .A2(n2373), .ZN(n2369) );
  INV_X1 U2298 ( .A(n2255), .ZN(n2373) );
  OR2_X1 U2299 ( .A1(n2374), .A2(n2262), .ZN(n2255) );
  INV_X1 U2300 ( .A(n2375), .ZN(n2262) );
  OR2_X1 U2301 ( .A1(n2376), .A2(n2377), .ZN(n2375) );
  AND2_X1 U2302 ( .A1(n2376), .A2(n2377), .ZN(n2374) );
  OR2_X1 U2303 ( .A1(n2378), .A2(n2379), .ZN(n2377) );
  AND2_X1 U2304 ( .A1(n2380), .A2(n2381), .ZN(n2379) );
  AND2_X1 U2305 ( .A1(n2382), .A2(n2383), .ZN(n2378) );
  OR2_X1 U2306 ( .A1(n2381), .A2(n2380), .ZN(n2383) );
  XOR2_X1 U2307 ( .A(n2384), .B(n2385), .Z(n2376) );
  XOR2_X1 U2308 ( .A(n2386), .B(n2387), .Z(n2385) );
  AND2_X1 U2309 ( .A1(n2243), .A2(n2388), .ZN(n2248) );
  AND2_X1 U2310 ( .A1(n2244), .A2(n2250), .ZN(n2388) );
  XOR2_X1 U2311 ( .A(n2372), .B(n2371), .Z(n2250) );
  OR2_X1 U2312 ( .A1(n2389), .A2(n2390), .ZN(n2371) );
  AND2_X1 U2313 ( .A1(n2391), .A2(n2392), .ZN(n2390) );
  AND2_X1 U2314 ( .A1(n2393), .A2(n2394), .ZN(n2389) );
  OR2_X1 U2315 ( .A1(n2391), .A2(n2392), .ZN(n2394) );
  XOR2_X1 U2316 ( .A(n2382), .B(n2395), .Z(n2372) );
  XOR2_X1 U2317 ( .A(n2381), .B(n2380), .Z(n2395) );
  OR2_X1 U2318 ( .A1(n2205), .A2(n1987), .ZN(n2380) );
  OR2_X1 U2319 ( .A1(n2396), .A2(n2397), .ZN(n2381) );
  AND2_X1 U2320 ( .A1(n2398), .A2(n2399), .ZN(n2397) );
  AND2_X1 U2321 ( .A1(n2400), .A2(n2401), .ZN(n2396) );
  OR2_X1 U2322 ( .A1(n2399), .A2(n2398), .ZN(n2401) );
  XOR2_X1 U2323 ( .A(n2402), .B(n2403), .Z(n2382) );
  XOR2_X1 U2324 ( .A(n2404), .B(n2405), .Z(n2403) );
  XNOR2_X1 U2325 ( .A(n2393), .B(n2406), .ZN(n2244) );
  XOR2_X1 U2326 ( .A(n2392), .B(n2391), .Z(n2406) );
  OR2_X1 U2327 ( .A1(n2205), .A2(n1966), .ZN(n2391) );
  OR2_X1 U2328 ( .A1(n2407), .A2(n2408), .ZN(n2392) );
  AND2_X1 U2329 ( .A1(n2409), .A2(n2410), .ZN(n2408) );
  AND2_X1 U2330 ( .A1(n2411), .A2(n2412), .ZN(n2407) );
  OR2_X1 U2331 ( .A1(n2410), .A2(n2409), .ZN(n2412) );
  XOR2_X1 U2332 ( .A(n2400), .B(n2413), .Z(n2393) );
  XOR2_X1 U2333 ( .A(n2399), .B(n2398), .Z(n2413) );
  OR2_X1 U2334 ( .A1(n2190), .A2(n1987), .ZN(n2398) );
  OR2_X1 U2335 ( .A1(n2414), .A2(n2415), .ZN(n2399) );
  AND2_X1 U2336 ( .A1(n2416), .A2(n2417), .ZN(n2415) );
  AND2_X1 U2337 ( .A1(n2418), .A2(n2419), .ZN(n2414) );
  OR2_X1 U2338 ( .A1(n2417), .A2(n2416), .ZN(n2419) );
  XOR2_X1 U2339 ( .A(n2420), .B(n2421), .Z(n2400) );
  XOR2_X1 U2340 ( .A(n2422), .B(n2423), .Z(n2421) );
  INV_X1 U2341 ( .A(n2424), .ZN(n2243) );
  OR2_X1 U2342 ( .A1(n2425), .A2(n2426), .ZN(n2424) );
  AND2_X1 U2343 ( .A1(n2201), .A2(n2200), .ZN(n2426) );
  AND2_X1 U2344 ( .A1(n2198), .A2(n2427), .ZN(n2425) );
  OR2_X1 U2345 ( .A1(n2201), .A2(n2200), .ZN(n2427) );
  OR2_X1 U2346 ( .A1(n2428), .A2(n2429), .ZN(n2200) );
  AND2_X1 U2347 ( .A1(n2182), .A2(n2181), .ZN(n2429) );
  AND2_X1 U2348 ( .A1(n2179), .A2(n2430), .ZN(n2428) );
  OR2_X1 U2349 ( .A1(n2182), .A2(n2181), .ZN(n2430) );
  OR2_X1 U2350 ( .A1(n2431), .A2(n2432), .ZN(n2181) );
  AND2_X1 U2351 ( .A1(n2169), .A2(n2168), .ZN(n2432) );
  AND2_X1 U2352 ( .A1(n2166), .A2(n2433), .ZN(n2431) );
  OR2_X1 U2353 ( .A1(n2169), .A2(n2168), .ZN(n2433) );
  OR2_X1 U2354 ( .A1(n2434), .A2(n2435), .ZN(n2168) );
  AND2_X1 U2355 ( .A1(n2150), .A2(n2149), .ZN(n2435) );
  AND2_X1 U2356 ( .A1(n2147), .A2(n2436), .ZN(n2434) );
  OR2_X1 U2357 ( .A1(n2150), .A2(n2149), .ZN(n2436) );
  OR2_X1 U2358 ( .A1(n2437), .A2(n2438), .ZN(n2149) );
  AND2_X1 U2359 ( .A1(n2127), .A2(n2126), .ZN(n2438) );
  AND2_X1 U2360 ( .A1(n2124), .A2(n2439), .ZN(n2437) );
  OR2_X1 U2361 ( .A1(n2127), .A2(n2126), .ZN(n2439) );
  OR2_X1 U2362 ( .A1(n2440), .A2(n2441), .ZN(n2126) );
  AND2_X1 U2363 ( .A1(n2108), .A2(n2107), .ZN(n2441) );
  AND2_X1 U2364 ( .A1(n2105), .A2(n2442), .ZN(n2440) );
  OR2_X1 U2365 ( .A1(n2108), .A2(n2107), .ZN(n2442) );
  OR2_X1 U2366 ( .A1(n2443), .A2(n2444), .ZN(n2107) );
  AND2_X1 U2367 ( .A1(n2095), .A2(n2094), .ZN(n2444) );
  AND2_X1 U2368 ( .A1(n2092), .A2(n2445), .ZN(n2443) );
  OR2_X1 U2369 ( .A1(n2095), .A2(n2094), .ZN(n2445) );
  OR2_X1 U2370 ( .A1(n2446), .A2(n2447), .ZN(n2094) );
  AND2_X1 U2371 ( .A1(n2076), .A2(n2075), .ZN(n2447) );
  AND2_X1 U2372 ( .A1(n2073), .A2(n2448), .ZN(n2446) );
  OR2_X1 U2373 ( .A1(n2076), .A2(n2075), .ZN(n2448) );
  OR2_X1 U2374 ( .A1(n2449), .A2(n2450), .ZN(n2075) );
  AND2_X1 U2375 ( .A1(n2063), .A2(n2062), .ZN(n2450) );
  AND2_X1 U2376 ( .A1(n2060), .A2(n2451), .ZN(n2449) );
  OR2_X1 U2377 ( .A1(n2063), .A2(n2062), .ZN(n2451) );
  OR2_X1 U2378 ( .A1(n2452), .A2(n2453), .ZN(n2062) );
  AND2_X1 U2379 ( .A1(n2044), .A2(n2043), .ZN(n2453) );
  AND2_X1 U2380 ( .A1(n2041), .A2(n2454), .ZN(n2452) );
  OR2_X1 U2381 ( .A1(n2044), .A2(n2043), .ZN(n2454) );
  OR2_X1 U2382 ( .A1(n2455), .A2(n2456), .ZN(n2043) );
  AND2_X1 U2383 ( .A1(n2031), .A2(n2030), .ZN(n2456) );
  AND2_X1 U2384 ( .A1(n2028), .A2(n2457), .ZN(n2455) );
  OR2_X1 U2385 ( .A1(n2031), .A2(n2030), .ZN(n2457) );
  OR2_X1 U2386 ( .A1(n2458), .A2(n2459), .ZN(n2030) );
  AND2_X1 U2387 ( .A1(n2012), .A2(n2011), .ZN(n2459) );
  AND2_X1 U2388 ( .A1(n2009), .A2(n2460), .ZN(n2458) );
  OR2_X1 U2389 ( .A1(n2012), .A2(n2011), .ZN(n2460) );
  OR2_X1 U2390 ( .A1(n2461), .A2(n2462), .ZN(n2011) );
  AND2_X1 U2391 ( .A1(n1999), .A2(n1998), .ZN(n2462) );
  AND2_X1 U2392 ( .A1(n1996), .A2(n2463), .ZN(n2461) );
  OR2_X1 U2393 ( .A1(n1999), .A2(n1998), .ZN(n2463) );
  OR2_X1 U2394 ( .A1(n2464), .A2(n2465), .ZN(n1998) );
  AND2_X1 U2395 ( .A1(n1977), .A2(n1980), .ZN(n2465) );
  AND2_X1 U2396 ( .A1(n2466), .A2(n2467), .ZN(n2464) );
  OR2_X1 U2397 ( .A1(n1977), .A2(n1980), .ZN(n2467) );
  OR2_X1 U2398 ( .A1(n1989), .A2(n1970), .ZN(n1980) );
  OR2_X1 U2399 ( .A1(n1966), .A2(n2238), .ZN(n1977) );
  OR2_X1 U2400 ( .A1(n2468), .A2(n1970), .ZN(n2238) );
  INV_X1 U2401 ( .A(n1979), .ZN(n2466) );
  OR2_X1 U2402 ( .A1(n2469), .A2(n2470), .ZN(n1979) );
  AND2_X1 U2403 ( .A1(b_14_), .A2(n2471), .ZN(n2470) );
  OR2_X1 U2404 ( .A1(n2472), .A2(n1965), .ZN(n2471) );
  AND2_X1 U2405 ( .A1(a_14_), .A2(n1987), .ZN(n2472) );
  AND2_X1 U2406 ( .A1(b_13_), .A2(n2473), .ZN(n2469) );
  OR2_X1 U2407 ( .A1(n2474), .A2(n1969), .ZN(n2473) );
  AND2_X1 U2408 ( .A1(a_15_), .A2(n1966), .ZN(n2474) );
  OR2_X1 U2409 ( .A1(n2234), .A2(n1970), .ZN(n1999) );
  XNOR2_X1 U2410 ( .A(n2475), .B(n2476), .ZN(n1996) );
  XOR2_X1 U2411 ( .A(n2477), .B(n2478), .Z(n2476) );
  OR2_X1 U2412 ( .A1(n2020), .A2(n1970), .ZN(n2012) );
  XOR2_X1 U2413 ( .A(n2479), .B(n2480), .Z(n2009) );
  XOR2_X1 U2414 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR2_X1 U2415 ( .A1(n2229), .A2(n1970), .ZN(n2031) );
  XOR2_X1 U2416 ( .A(n2483), .B(n2484), .Z(n2028) );
  XOR2_X1 U2417 ( .A(n2485), .B(n2486), .Z(n2484) );
  OR2_X1 U2418 ( .A1(n2052), .A2(n1970), .ZN(n2044) );
  XOR2_X1 U2419 ( .A(n2487), .B(n2488), .Z(n2041) );
  XOR2_X1 U2420 ( .A(n2489), .B(n2490), .Z(n2488) );
  OR2_X1 U2421 ( .A1(n2224), .A2(n1970), .ZN(n2063) );
  XOR2_X1 U2422 ( .A(n2491), .B(n2492), .Z(n2060) );
  XOR2_X1 U2423 ( .A(n2493), .B(n2494), .Z(n2492) );
  OR2_X1 U2424 ( .A1(n2084), .A2(n1970), .ZN(n2076) );
  XOR2_X1 U2425 ( .A(n2495), .B(n2496), .Z(n2073) );
  XOR2_X1 U2426 ( .A(n2497), .B(n2498), .Z(n2496) );
  OR2_X1 U2427 ( .A1(n2219), .A2(n1970), .ZN(n2095) );
  XOR2_X1 U2428 ( .A(n2499), .B(n2500), .Z(n2092) );
  XOR2_X1 U2429 ( .A(n2501), .B(n2502), .Z(n2500) );
  OR2_X1 U2430 ( .A1(n2116), .A2(n1970), .ZN(n2108) );
  XOR2_X1 U2431 ( .A(n2503), .B(n2504), .Z(n2105) );
  XOR2_X1 U2432 ( .A(n2505), .B(n2506), .Z(n2504) );
  OR2_X1 U2433 ( .A1(n2214), .A2(n1970), .ZN(n2127) );
  XOR2_X1 U2434 ( .A(n2507), .B(n2508), .Z(n2124) );
  XOR2_X1 U2435 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR2_X1 U2436 ( .A1(n2158), .A2(n1970), .ZN(n2150) );
  XOR2_X1 U2437 ( .A(n2511), .B(n2512), .Z(n2147) );
  XOR2_X1 U2438 ( .A(n2513), .B(n2514), .Z(n2512) );
  OR2_X1 U2439 ( .A1(n2209), .A2(n1970), .ZN(n2169) );
  XOR2_X1 U2440 ( .A(n2515), .B(n2516), .Z(n2166) );
  XOR2_X1 U2441 ( .A(n2517), .B(n2518), .Z(n2516) );
  OR2_X1 U2442 ( .A1(n2190), .A2(n1970), .ZN(n2182) );
  XOR2_X1 U2443 ( .A(n2519), .B(n2520), .Z(n2179) );
  XOR2_X1 U2444 ( .A(n2521), .B(n2522), .Z(n2520) );
  OR2_X1 U2445 ( .A1(n2205), .A2(n1970), .ZN(n2201) );
  INV_X1 U2446 ( .A(b_15_), .ZN(n1970) );
  XOR2_X1 U2447 ( .A(n2411), .B(n2523), .Z(n2198) );
  XOR2_X1 U2448 ( .A(n2410), .B(n2409), .Z(n2523) );
  OR2_X1 U2449 ( .A1(n2190), .A2(n1966), .ZN(n2409) );
  OR2_X1 U2450 ( .A1(n2524), .A2(n2525), .ZN(n2410) );
  AND2_X1 U2451 ( .A1(n2522), .A2(n2521), .ZN(n2525) );
  AND2_X1 U2452 ( .A1(n2519), .A2(n2526), .ZN(n2524) );
  OR2_X1 U2453 ( .A1(n2521), .A2(n2522), .ZN(n2526) );
  OR2_X1 U2454 ( .A1(n2209), .A2(n1966), .ZN(n2522) );
  OR2_X1 U2455 ( .A1(n2527), .A2(n2528), .ZN(n2521) );
  AND2_X1 U2456 ( .A1(n2518), .A2(n2517), .ZN(n2528) );
  AND2_X1 U2457 ( .A1(n2515), .A2(n2529), .ZN(n2527) );
  OR2_X1 U2458 ( .A1(n2517), .A2(n2518), .ZN(n2529) );
  OR2_X1 U2459 ( .A1(n2158), .A2(n1966), .ZN(n2518) );
  OR2_X1 U2460 ( .A1(n2530), .A2(n2531), .ZN(n2517) );
  AND2_X1 U2461 ( .A1(n2514), .A2(n2513), .ZN(n2531) );
  AND2_X1 U2462 ( .A1(n2511), .A2(n2532), .ZN(n2530) );
  OR2_X1 U2463 ( .A1(n2513), .A2(n2514), .ZN(n2532) );
  OR2_X1 U2464 ( .A1(n2214), .A2(n1966), .ZN(n2514) );
  OR2_X1 U2465 ( .A1(n2533), .A2(n2534), .ZN(n2513) );
  AND2_X1 U2466 ( .A1(n2510), .A2(n2509), .ZN(n2534) );
  AND2_X1 U2467 ( .A1(n2507), .A2(n2535), .ZN(n2533) );
  OR2_X1 U2468 ( .A1(n2509), .A2(n2510), .ZN(n2535) );
  OR2_X1 U2469 ( .A1(n2116), .A2(n1966), .ZN(n2510) );
  OR2_X1 U2470 ( .A1(n2536), .A2(n2537), .ZN(n2509) );
  AND2_X1 U2471 ( .A1(n2506), .A2(n2505), .ZN(n2537) );
  AND2_X1 U2472 ( .A1(n2503), .A2(n2538), .ZN(n2536) );
  OR2_X1 U2473 ( .A1(n2505), .A2(n2506), .ZN(n2538) );
  OR2_X1 U2474 ( .A1(n2219), .A2(n1966), .ZN(n2506) );
  OR2_X1 U2475 ( .A1(n2539), .A2(n2540), .ZN(n2505) );
  AND2_X1 U2476 ( .A1(n2502), .A2(n2501), .ZN(n2540) );
  AND2_X1 U2477 ( .A1(n2499), .A2(n2541), .ZN(n2539) );
  OR2_X1 U2478 ( .A1(n2501), .A2(n2502), .ZN(n2541) );
  OR2_X1 U2479 ( .A1(n2084), .A2(n1966), .ZN(n2502) );
  OR2_X1 U2480 ( .A1(n2542), .A2(n2543), .ZN(n2501) );
  AND2_X1 U2481 ( .A1(n2498), .A2(n2497), .ZN(n2543) );
  AND2_X1 U2482 ( .A1(n2495), .A2(n2544), .ZN(n2542) );
  OR2_X1 U2483 ( .A1(n2497), .A2(n2498), .ZN(n2544) );
  OR2_X1 U2484 ( .A1(n2224), .A2(n1966), .ZN(n2498) );
  OR2_X1 U2485 ( .A1(n2545), .A2(n2546), .ZN(n2497) );
  AND2_X1 U2486 ( .A1(n2494), .A2(n2493), .ZN(n2546) );
  AND2_X1 U2487 ( .A1(n2491), .A2(n2547), .ZN(n2545) );
  OR2_X1 U2488 ( .A1(n2493), .A2(n2494), .ZN(n2547) );
  OR2_X1 U2489 ( .A1(n2052), .A2(n1966), .ZN(n2494) );
  OR2_X1 U2490 ( .A1(n2548), .A2(n2549), .ZN(n2493) );
  AND2_X1 U2491 ( .A1(n2490), .A2(n2489), .ZN(n2549) );
  AND2_X1 U2492 ( .A1(n2487), .A2(n2550), .ZN(n2548) );
  OR2_X1 U2493 ( .A1(n2489), .A2(n2490), .ZN(n2550) );
  OR2_X1 U2494 ( .A1(n2229), .A2(n1966), .ZN(n2490) );
  OR2_X1 U2495 ( .A1(n2551), .A2(n2552), .ZN(n2489) );
  AND2_X1 U2496 ( .A1(n2486), .A2(n2485), .ZN(n2552) );
  AND2_X1 U2497 ( .A1(n2483), .A2(n2553), .ZN(n2551) );
  OR2_X1 U2498 ( .A1(n2485), .A2(n2486), .ZN(n2553) );
  OR2_X1 U2499 ( .A1(n2020), .A2(n1966), .ZN(n2486) );
  OR2_X1 U2500 ( .A1(n2554), .A2(n2555), .ZN(n2485) );
  AND2_X1 U2501 ( .A1(n2482), .A2(n2481), .ZN(n2555) );
  AND2_X1 U2502 ( .A1(n2479), .A2(n2556), .ZN(n2554) );
  OR2_X1 U2503 ( .A1(n2481), .A2(n2482), .ZN(n2556) );
  OR2_X1 U2504 ( .A1(n2234), .A2(n1966), .ZN(n2482) );
  OR2_X1 U2505 ( .A1(n2557), .A2(n2558), .ZN(n2481) );
  AND2_X1 U2506 ( .A1(n2475), .A2(n2478), .ZN(n2558) );
  AND2_X1 U2507 ( .A1(n2559), .A2(n2560), .ZN(n2557) );
  OR2_X1 U2508 ( .A1(n2478), .A2(n2475), .ZN(n2560) );
  OR2_X1 U2509 ( .A1(n1989), .A2(n1966), .ZN(n2475) );
  OR2_X1 U2510 ( .A1(n1966), .A2(n2561), .ZN(n2478) );
  INV_X1 U2511 ( .A(b_14_), .ZN(n1966) );
  INV_X1 U2512 ( .A(n2477), .ZN(n2559) );
  OR2_X1 U2513 ( .A1(n2562), .A2(n2563), .ZN(n2477) );
  AND2_X1 U2514 ( .A1(b_13_), .A2(n2564), .ZN(n2563) );
  OR2_X1 U2515 ( .A1(n2565), .A2(n1965), .ZN(n2564) );
  AND2_X1 U2516 ( .A1(a_14_), .A2(n2235), .ZN(n2565) );
  AND2_X1 U2517 ( .A1(b_12_), .A2(n2566), .ZN(n2562) );
  OR2_X1 U2518 ( .A1(n2567), .A2(n1969), .ZN(n2566) );
  AND2_X1 U2519 ( .A1(a_15_), .A2(n1987), .ZN(n2567) );
  XNOR2_X1 U2520 ( .A(n1992), .B(n2568), .ZN(n2479) );
  XOR2_X1 U2521 ( .A(n2569), .B(n2570), .Z(n2568) );
  XOR2_X1 U2522 ( .A(n2571), .B(n2572), .Z(n2483) );
  XOR2_X1 U2523 ( .A(n2573), .B(n2574), .Z(n2572) );
  XOR2_X1 U2524 ( .A(n2575), .B(n2576), .Z(n2487) );
  XOR2_X1 U2525 ( .A(n2577), .B(n2578), .Z(n2576) );
  XOR2_X1 U2526 ( .A(n2579), .B(n2580), .Z(n2491) );
  XOR2_X1 U2527 ( .A(n2581), .B(n2582), .Z(n2580) );
  XOR2_X1 U2528 ( .A(n2583), .B(n2584), .Z(n2495) );
  XOR2_X1 U2529 ( .A(n2585), .B(n2586), .Z(n2584) );
  XOR2_X1 U2530 ( .A(n2587), .B(n2588), .Z(n2499) );
  XOR2_X1 U2531 ( .A(n2589), .B(n2590), .Z(n2588) );
  XOR2_X1 U2532 ( .A(n2591), .B(n2592), .Z(n2503) );
  XOR2_X1 U2533 ( .A(n2593), .B(n2594), .Z(n2592) );
  XOR2_X1 U2534 ( .A(n2595), .B(n2596), .Z(n2507) );
  XOR2_X1 U2535 ( .A(n2597), .B(n2598), .Z(n2596) );
  XOR2_X1 U2536 ( .A(n2599), .B(n2600), .Z(n2511) );
  XOR2_X1 U2537 ( .A(n2601), .B(n2602), .Z(n2600) );
  XOR2_X1 U2538 ( .A(n2603), .B(n2604), .Z(n2515) );
  XOR2_X1 U2539 ( .A(n2605), .B(n2606), .Z(n2604) );
  XOR2_X1 U2540 ( .A(n2607), .B(n2608), .Z(n2519) );
  XOR2_X1 U2541 ( .A(n2609), .B(n2610), .Z(n2608) );
  XOR2_X1 U2542 ( .A(n2418), .B(n2611), .Z(n2411) );
  XOR2_X1 U2543 ( .A(n2417), .B(n2416), .Z(n2611) );
  OR2_X1 U2544 ( .A1(n2209), .A2(n1987), .ZN(n2416) );
  OR2_X1 U2545 ( .A1(n2612), .A2(n2613), .ZN(n2417) );
  AND2_X1 U2546 ( .A1(n2610), .A2(n2609), .ZN(n2613) );
  AND2_X1 U2547 ( .A1(n2607), .A2(n2614), .ZN(n2612) );
  OR2_X1 U2548 ( .A1(n2609), .A2(n2610), .ZN(n2614) );
  OR2_X1 U2549 ( .A1(n2158), .A2(n1987), .ZN(n2610) );
  OR2_X1 U2550 ( .A1(n2615), .A2(n2616), .ZN(n2609) );
  AND2_X1 U2551 ( .A1(n2606), .A2(n2605), .ZN(n2616) );
  AND2_X1 U2552 ( .A1(n2603), .A2(n2617), .ZN(n2615) );
  OR2_X1 U2553 ( .A1(n2605), .A2(n2606), .ZN(n2617) );
  OR2_X1 U2554 ( .A1(n2214), .A2(n1987), .ZN(n2606) );
  OR2_X1 U2555 ( .A1(n2618), .A2(n2619), .ZN(n2605) );
  AND2_X1 U2556 ( .A1(n2602), .A2(n2601), .ZN(n2619) );
  AND2_X1 U2557 ( .A1(n2599), .A2(n2620), .ZN(n2618) );
  OR2_X1 U2558 ( .A1(n2601), .A2(n2602), .ZN(n2620) );
  OR2_X1 U2559 ( .A1(n2116), .A2(n1987), .ZN(n2602) );
  OR2_X1 U2560 ( .A1(n2621), .A2(n2622), .ZN(n2601) );
  AND2_X1 U2561 ( .A1(n2598), .A2(n2597), .ZN(n2622) );
  AND2_X1 U2562 ( .A1(n2595), .A2(n2623), .ZN(n2621) );
  OR2_X1 U2563 ( .A1(n2597), .A2(n2598), .ZN(n2623) );
  OR2_X1 U2564 ( .A1(n2219), .A2(n1987), .ZN(n2598) );
  OR2_X1 U2565 ( .A1(n2624), .A2(n2625), .ZN(n2597) );
  AND2_X1 U2566 ( .A1(n2594), .A2(n2593), .ZN(n2625) );
  AND2_X1 U2567 ( .A1(n2591), .A2(n2626), .ZN(n2624) );
  OR2_X1 U2568 ( .A1(n2593), .A2(n2594), .ZN(n2626) );
  OR2_X1 U2569 ( .A1(n2084), .A2(n1987), .ZN(n2594) );
  OR2_X1 U2570 ( .A1(n2627), .A2(n2628), .ZN(n2593) );
  AND2_X1 U2571 ( .A1(n2590), .A2(n2589), .ZN(n2628) );
  AND2_X1 U2572 ( .A1(n2587), .A2(n2629), .ZN(n2627) );
  OR2_X1 U2573 ( .A1(n2589), .A2(n2590), .ZN(n2629) );
  OR2_X1 U2574 ( .A1(n2224), .A2(n1987), .ZN(n2590) );
  OR2_X1 U2575 ( .A1(n2630), .A2(n2631), .ZN(n2589) );
  AND2_X1 U2576 ( .A1(n2586), .A2(n2585), .ZN(n2631) );
  AND2_X1 U2577 ( .A1(n2583), .A2(n2632), .ZN(n2630) );
  OR2_X1 U2578 ( .A1(n2585), .A2(n2586), .ZN(n2632) );
  OR2_X1 U2579 ( .A1(n2052), .A2(n1987), .ZN(n2586) );
  OR2_X1 U2580 ( .A1(n2633), .A2(n2634), .ZN(n2585) );
  AND2_X1 U2581 ( .A1(n2582), .A2(n2581), .ZN(n2634) );
  AND2_X1 U2582 ( .A1(n2579), .A2(n2635), .ZN(n2633) );
  OR2_X1 U2583 ( .A1(n2581), .A2(n2582), .ZN(n2635) );
  OR2_X1 U2584 ( .A1(n2229), .A2(n1987), .ZN(n2582) );
  OR2_X1 U2585 ( .A1(n2636), .A2(n2637), .ZN(n2581) );
  AND2_X1 U2586 ( .A1(n2578), .A2(n2577), .ZN(n2637) );
  AND2_X1 U2587 ( .A1(n2575), .A2(n2638), .ZN(n2636) );
  OR2_X1 U2588 ( .A1(n2577), .A2(n2578), .ZN(n2638) );
  OR2_X1 U2589 ( .A1(n2020), .A2(n1987), .ZN(n2578) );
  OR2_X1 U2590 ( .A1(n2639), .A2(n2640), .ZN(n2577) );
  AND2_X1 U2591 ( .A1(n2574), .A2(n2573), .ZN(n2640) );
  AND2_X1 U2592 ( .A1(n2571), .A2(n2641), .ZN(n2639) );
  OR2_X1 U2593 ( .A1(n2573), .A2(n2574), .ZN(n2641) );
  OR2_X1 U2594 ( .A1(n2234), .A2(n1987), .ZN(n2574) );
  OR2_X1 U2595 ( .A1(n2642), .A2(n2643), .ZN(n2573) );
  AND2_X1 U2596 ( .A1(n1992), .A2(n2570), .ZN(n2643) );
  AND2_X1 U2597 ( .A1(n2644), .A2(n2645), .ZN(n2642) );
  OR2_X1 U2598 ( .A1(n2570), .A2(n1992), .ZN(n2645) );
  OR2_X1 U2599 ( .A1(n1989), .A2(n1987), .ZN(n1992) );
  OR2_X1 U2600 ( .A1(n2235), .A2(n2561), .ZN(n2570) );
  OR2_X1 U2601 ( .A1(n2468), .A2(n1987), .ZN(n2561) );
  INV_X1 U2602 ( .A(b_13_), .ZN(n1987) );
  INV_X1 U2603 ( .A(n2569), .ZN(n2644) );
  OR2_X1 U2604 ( .A1(n2646), .A2(n2647), .ZN(n2569) );
  AND2_X1 U2605 ( .A1(b_12_), .A2(n2648), .ZN(n2647) );
  OR2_X1 U2606 ( .A1(n2649), .A2(n1965), .ZN(n2648) );
  AND2_X1 U2607 ( .A1(a_14_), .A2(n2019), .ZN(n2649) );
  AND2_X1 U2608 ( .A1(b_11_), .A2(n2650), .ZN(n2646) );
  OR2_X1 U2609 ( .A1(n2651), .A2(n1969), .ZN(n2650) );
  AND2_X1 U2610 ( .A1(a_15_), .A2(n2235), .ZN(n2651) );
  XNOR2_X1 U2611 ( .A(n2652), .B(n2653), .ZN(n2571) );
  XOR2_X1 U2612 ( .A(n2654), .B(n2655), .Z(n2653) );
  XOR2_X1 U2613 ( .A(n2656), .B(n2657), .Z(n2575) );
  XOR2_X1 U2614 ( .A(n2658), .B(n2005), .Z(n2657) );
  XOR2_X1 U2615 ( .A(n2659), .B(n2660), .Z(n2579) );
  XOR2_X1 U2616 ( .A(n2661), .B(n2662), .Z(n2660) );
  XOR2_X1 U2617 ( .A(n2663), .B(n2664), .Z(n2583) );
  XOR2_X1 U2618 ( .A(n2665), .B(n2666), .Z(n2664) );
  XOR2_X1 U2619 ( .A(n2667), .B(n2668), .Z(n2587) );
  XOR2_X1 U2620 ( .A(n2669), .B(n2670), .Z(n2668) );
  XOR2_X1 U2621 ( .A(n2671), .B(n2672), .Z(n2591) );
  XOR2_X1 U2622 ( .A(n2673), .B(n2674), .Z(n2672) );
  XOR2_X1 U2623 ( .A(n2675), .B(n2676), .Z(n2595) );
  XOR2_X1 U2624 ( .A(n2677), .B(n2678), .Z(n2676) );
  XOR2_X1 U2625 ( .A(n2679), .B(n2680), .Z(n2599) );
  XOR2_X1 U2626 ( .A(n2681), .B(n2682), .Z(n2680) );
  XOR2_X1 U2627 ( .A(n2683), .B(n2684), .Z(n2603) );
  XOR2_X1 U2628 ( .A(n2685), .B(n2686), .Z(n2684) );
  XOR2_X1 U2629 ( .A(n2687), .B(n2688), .Z(n2607) );
  XOR2_X1 U2630 ( .A(n2689), .B(n2690), .Z(n2688) );
  XOR2_X1 U2631 ( .A(n2691), .B(n2692), .Z(n2418) );
  XOR2_X1 U2632 ( .A(n2693), .B(n2694), .Z(n2692) );
  XOR2_X1 U2633 ( .A(n2273), .B(n2272), .Z(n2263) );
  INV_X1 U2634 ( .A(n2695), .ZN(n2272) );
  OR2_X1 U2635 ( .A1(n2696), .A2(n2697), .ZN(n2695) );
  AND2_X1 U2636 ( .A1(n2387), .A2(n2386), .ZN(n2697) );
  AND2_X1 U2637 ( .A1(n2384), .A2(n2698), .ZN(n2696) );
  OR2_X1 U2638 ( .A1(n2386), .A2(n2387), .ZN(n2698) );
  OR2_X1 U2639 ( .A1(n2205), .A2(n2235), .ZN(n2387) );
  OR2_X1 U2640 ( .A1(n2699), .A2(n2700), .ZN(n2386) );
  AND2_X1 U2641 ( .A1(n2405), .A2(n2404), .ZN(n2700) );
  AND2_X1 U2642 ( .A1(n2402), .A2(n2701), .ZN(n2699) );
  OR2_X1 U2643 ( .A1(n2404), .A2(n2405), .ZN(n2701) );
  OR2_X1 U2644 ( .A1(n2190), .A2(n2235), .ZN(n2405) );
  OR2_X1 U2645 ( .A1(n2702), .A2(n2703), .ZN(n2404) );
  AND2_X1 U2646 ( .A1(n2423), .A2(n2422), .ZN(n2703) );
  AND2_X1 U2647 ( .A1(n2420), .A2(n2704), .ZN(n2702) );
  OR2_X1 U2648 ( .A1(n2422), .A2(n2423), .ZN(n2704) );
  OR2_X1 U2649 ( .A1(n2209), .A2(n2235), .ZN(n2423) );
  OR2_X1 U2650 ( .A1(n2705), .A2(n2706), .ZN(n2422) );
  AND2_X1 U2651 ( .A1(n2694), .A2(n2693), .ZN(n2706) );
  AND2_X1 U2652 ( .A1(n2691), .A2(n2707), .ZN(n2705) );
  OR2_X1 U2653 ( .A1(n2693), .A2(n2694), .ZN(n2707) );
  OR2_X1 U2654 ( .A1(n2158), .A2(n2235), .ZN(n2694) );
  OR2_X1 U2655 ( .A1(n2708), .A2(n2709), .ZN(n2693) );
  AND2_X1 U2656 ( .A1(n2690), .A2(n2689), .ZN(n2709) );
  AND2_X1 U2657 ( .A1(n2687), .A2(n2710), .ZN(n2708) );
  OR2_X1 U2658 ( .A1(n2689), .A2(n2690), .ZN(n2710) );
  OR2_X1 U2659 ( .A1(n2214), .A2(n2235), .ZN(n2690) );
  OR2_X1 U2660 ( .A1(n2711), .A2(n2712), .ZN(n2689) );
  AND2_X1 U2661 ( .A1(n2686), .A2(n2685), .ZN(n2712) );
  AND2_X1 U2662 ( .A1(n2683), .A2(n2713), .ZN(n2711) );
  OR2_X1 U2663 ( .A1(n2685), .A2(n2686), .ZN(n2713) );
  OR2_X1 U2664 ( .A1(n2116), .A2(n2235), .ZN(n2686) );
  OR2_X1 U2665 ( .A1(n2714), .A2(n2715), .ZN(n2685) );
  AND2_X1 U2666 ( .A1(n2682), .A2(n2681), .ZN(n2715) );
  AND2_X1 U2667 ( .A1(n2679), .A2(n2716), .ZN(n2714) );
  OR2_X1 U2668 ( .A1(n2681), .A2(n2682), .ZN(n2716) );
  OR2_X1 U2669 ( .A1(n2219), .A2(n2235), .ZN(n2682) );
  OR2_X1 U2670 ( .A1(n2717), .A2(n2718), .ZN(n2681) );
  AND2_X1 U2671 ( .A1(n2678), .A2(n2677), .ZN(n2718) );
  AND2_X1 U2672 ( .A1(n2675), .A2(n2719), .ZN(n2717) );
  OR2_X1 U2673 ( .A1(n2677), .A2(n2678), .ZN(n2719) );
  OR2_X1 U2674 ( .A1(n2084), .A2(n2235), .ZN(n2678) );
  OR2_X1 U2675 ( .A1(n2720), .A2(n2721), .ZN(n2677) );
  AND2_X1 U2676 ( .A1(n2674), .A2(n2673), .ZN(n2721) );
  AND2_X1 U2677 ( .A1(n2671), .A2(n2722), .ZN(n2720) );
  OR2_X1 U2678 ( .A1(n2673), .A2(n2674), .ZN(n2722) );
  OR2_X1 U2679 ( .A1(n2224), .A2(n2235), .ZN(n2674) );
  OR2_X1 U2680 ( .A1(n2723), .A2(n2724), .ZN(n2673) );
  AND2_X1 U2681 ( .A1(n2670), .A2(n2669), .ZN(n2724) );
  AND2_X1 U2682 ( .A1(n2667), .A2(n2725), .ZN(n2723) );
  OR2_X1 U2683 ( .A1(n2669), .A2(n2670), .ZN(n2725) );
  OR2_X1 U2684 ( .A1(n2052), .A2(n2235), .ZN(n2670) );
  OR2_X1 U2685 ( .A1(n2726), .A2(n2727), .ZN(n2669) );
  AND2_X1 U2686 ( .A1(n2666), .A2(n2665), .ZN(n2727) );
  AND2_X1 U2687 ( .A1(n2663), .A2(n2728), .ZN(n2726) );
  OR2_X1 U2688 ( .A1(n2665), .A2(n2666), .ZN(n2728) );
  OR2_X1 U2689 ( .A1(n2229), .A2(n2235), .ZN(n2666) );
  OR2_X1 U2690 ( .A1(n2729), .A2(n2730), .ZN(n2665) );
  AND2_X1 U2691 ( .A1(n2662), .A2(n2661), .ZN(n2730) );
  AND2_X1 U2692 ( .A1(n2659), .A2(n2731), .ZN(n2729) );
  OR2_X1 U2693 ( .A1(n2661), .A2(n2662), .ZN(n2731) );
  OR2_X1 U2694 ( .A1(n2020), .A2(n2235), .ZN(n2662) );
  OR2_X1 U2695 ( .A1(n2732), .A2(n2733), .ZN(n2661) );
  AND2_X1 U2696 ( .A1(n2005), .A2(n2658), .ZN(n2733) );
  AND2_X1 U2697 ( .A1(n2656), .A2(n2734), .ZN(n2732) );
  OR2_X1 U2698 ( .A1(n2658), .A2(n2005), .ZN(n2734) );
  OR2_X1 U2699 ( .A1(n2234), .A2(n2235), .ZN(n2005) );
  OR2_X1 U2700 ( .A1(n2735), .A2(n2736), .ZN(n2658) );
  AND2_X1 U2701 ( .A1(n2652), .A2(n2655), .ZN(n2736) );
  AND2_X1 U2702 ( .A1(n2737), .A2(n2738), .ZN(n2735) );
  OR2_X1 U2703 ( .A1(n2655), .A2(n2652), .ZN(n2738) );
  OR2_X1 U2704 ( .A1(n1989), .A2(n2235), .ZN(n2652) );
  OR2_X1 U2705 ( .A1(n2019), .A2(n2739), .ZN(n2655) );
  OR2_X1 U2706 ( .A1(n2468), .A2(n2235), .ZN(n2739) );
  INV_X1 U2707 ( .A(b_12_), .ZN(n2235) );
  INV_X1 U2708 ( .A(n2654), .ZN(n2737) );
  OR2_X1 U2709 ( .A1(n2740), .A2(n2741), .ZN(n2654) );
  AND2_X1 U2710 ( .A1(b_11_), .A2(n2742), .ZN(n2741) );
  OR2_X1 U2711 ( .A1(n2743), .A2(n1965), .ZN(n2742) );
  AND2_X1 U2712 ( .A1(a_14_), .A2(n2230), .ZN(n2743) );
  AND2_X1 U2713 ( .A1(b_10_), .A2(n2744), .ZN(n2740) );
  OR2_X1 U2714 ( .A1(n2745), .A2(n1969), .ZN(n2744) );
  AND2_X1 U2715 ( .A1(a_15_), .A2(n2019), .ZN(n2745) );
  XNOR2_X1 U2716 ( .A(n2746), .B(n2747), .ZN(n2656) );
  XOR2_X1 U2717 ( .A(n2748), .B(n2749), .Z(n2747) );
  XOR2_X1 U2718 ( .A(n2750), .B(n2751), .Z(n2659) );
  XOR2_X1 U2719 ( .A(n2752), .B(n2753), .Z(n2751) );
  XOR2_X1 U2720 ( .A(n2754), .B(n2755), .Z(n2663) );
  XOR2_X1 U2721 ( .A(n2756), .B(n2024), .Z(n2755) );
  XOR2_X1 U2722 ( .A(n2757), .B(n2758), .Z(n2667) );
  XOR2_X1 U2723 ( .A(n2759), .B(n2760), .Z(n2758) );
  XOR2_X1 U2724 ( .A(n2761), .B(n2762), .Z(n2671) );
  XOR2_X1 U2725 ( .A(n2763), .B(n2764), .Z(n2762) );
  XOR2_X1 U2726 ( .A(n2765), .B(n2766), .Z(n2675) );
  XOR2_X1 U2727 ( .A(n2767), .B(n2768), .Z(n2766) );
  XOR2_X1 U2728 ( .A(n2769), .B(n2770), .Z(n2679) );
  XOR2_X1 U2729 ( .A(n2771), .B(n2772), .Z(n2770) );
  XOR2_X1 U2730 ( .A(n2773), .B(n2774), .Z(n2683) );
  XOR2_X1 U2731 ( .A(n2775), .B(n2776), .Z(n2774) );
  XOR2_X1 U2732 ( .A(n2777), .B(n2778), .Z(n2687) );
  XOR2_X1 U2733 ( .A(n2779), .B(n2780), .Z(n2778) );
  XOR2_X1 U2734 ( .A(n2781), .B(n2782), .Z(n2691) );
  XOR2_X1 U2735 ( .A(n2783), .B(n2784), .Z(n2782) );
  XOR2_X1 U2736 ( .A(n2785), .B(n2786), .Z(n2420) );
  XOR2_X1 U2737 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR2_X1 U2738 ( .A(n2789), .B(n2790), .Z(n2402) );
  XOR2_X1 U2739 ( .A(n2791), .B(n2792), .Z(n2790) );
  XOR2_X1 U2740 ( .A(n2793), .B(n2794), .Z(n2384) );
  XOR2_X1 U2741 ( .A(n2795), .B(n2796), .Z(n2794) );
  XNOR2_X1 U2742 ( .A(n2797), .B(n2798), .ZN(n2273) );
  XOR2_X1 U2743 ( .A(n2799), .B(n2800), .Z(n2798) );
  XOR2_X1 U2744 ( .A(n2365), .B(n2364), .Z(n2271) );
  INV_X1 U2745 ( .A(n2801), .ZN(n2364) );
  OR2_X1 U2746 ( .A1(n2802), .A2(n2803), .ZN(n2801) );
  AND2_X1 U2747 ( .A1(n2800), .A2(n2799), .ZN(n2803) );
  AND2_X1 U2748 ( .A1(n2797), .A2(n2804), .ZN(n2802) );
  OR2_X1 U2749 ( .A1(n2799), .A2(n2800), .ZN(n2804) );
  OR2_X1 U2750 ( .A1(n2205), .A2(n2019), .ZN(n2800) );
  OR2_X1 U2751 ( .A1(n2805), .A2(n2806), .ZN(n2799) );
  AND2_X1 U2752 ( .A1(n2796), .A2(n2795), .ZN(n2806) );
  AND2_X1 U2753 ( .A1(n2793), .A2(n2807), .ZN(n2805) );
  OR2_X1 U2754 ( .A1(n2795), .A2(n2796), .ZN(n2807) );
  OR2_X1 U2755 ( .A1(n2190), .A2(n2019), .ZN(n2796) );
  OR2_X1 U2756 ( .A1(n2808), .A2(n2809), .ZN(n2795) );
  AND2_X1 U2757 ( .A1(n2792), .A2(n2791), .ZN(n2809) );
  AND2_X1 U2758 ( .A1(n2789), .A2(n2810), .ZN(n2808) );
  OR2_X1 U2759 ( .A1(n2791), .A2(n2792), .ZN(n2810) );
  OR2_X1 U2760 ( .A1(n2209), .A2(n2019), .ZN(n2792) );
  OR2_X1 U2761 ( .A1(n2811), .A2(n2812), .ZN(n2791) );
  AND2_X1 U2762 ( .A1(n2788), .A2(n2787), .ZN(n2812) );
  AND2_X1 U2763 ( .A1(n2785), .A2(n2813), .ZN(n2811) );
  OR2_X1 U2764 ( .A1(n2787), .A2(n2788), .ZN(n2813) );
  OR2_X1 U2765 ( .A1(n2158), .A2(n2019), .ZN(n2788) );
  OR2_X1 U2766 ( .A1(n2814), .A2(n2815), .ZN(n2787) );
  AND2_X1 U2767 ( .A1(n2784), .A2(n2783), .ZN(n2815) );
  AND2_X1 U2768 ( .A1(n2781), .A2(n2816), .ZN(n2814) );
  OR2_X1 U2769 ( .A1(n2783), .A2(n2784), .ZN(n2816) );
  OR2_X1 U2770 ( .A1(n2214), .A2(n2019), .ZN(n2784) );
  OR2_X1 U2771 ( .A1(n2817), .A2(n2818), .ZN(n2783) );
  AND2_X1 U2772 ( .A1(n2780), .A2(n2779), .ZN(n2818) );
  AND2_X1 U2773 ( .A1(n2777), .A2(n2819), .ZN(n2817) );
  OR2_X1 U2774 ( .A1(n2779), .A2(n2780), .ZN(n2819) );
  OR2_X1 U2775 ( .A1(n2116), .A2(n2019), .ZN(n2780) );
  OR2_X1 U2776 ( .A1(n2820), .A2(n2821), .ZN(n2779) );
  AND2_X1 U2777 ( .A1(n2776), .A2(n2775), .ZN(n2821) );
  AND2_X1 U2778 ( .A1(n2773), .A2(n2822), .ZN(n2820) );
  OR2_X1 U2779 ( .A1(n2775), .A2(n2776), .ZN(n2822) );
  OR2_X1 U2780 ( .A1(n2219), .A2(n2019), .ZN(n2776) );
  OR2_X1 U2781 ( .A1(n2823), .A2(n2824), .ZN(n2775) );
  AND2_X1 U2782 ( .A1(n2772), .A2(n2771), .ZN(n2824) );
  AND2_X1 U2783 ( .A1(n2769), .A2(n2825), .ZN(n2823) );
  OR2_X1 U2784 ( .A1(n2771), .A2(n2772), .ZN(n2825) );
  OR2_X1 U2785 ( .A1(n2084), .A2(n2019), .ZN(n2772) );
  OR2_X1 U2786 ( .A1(n2826), .A2(n2827), .ZN(n2771) );
  AND2_X1 U2787 ( .A1(n2768), .A2(n2767), .ZN(n2827) );
  AND2_X1 U2788 ( .A1(n2765), .A2(n2828), .ZN(n2826) );
  OR2_X1 U2789 ( .A1(n2767), .A2(n2768), .ZN(n2828) );
  OR2_X1 U2790 ( .A1(n2224), .A2(n2019), .ZN(n2768) );
  OR2_X1 U2791 ( .A1(n2829), .A2(n2830), .ZN(n2767) );
  AND2_X1 U2792 ( .A1(n2764), .A2(n2763), .ZN(n2830) );
  AND2_X1 U2793 ( .A1(n2761), .A2(n2831), .ZN(n2829) );
  OR2_X1 U2794 ( .A1(n2763), .A2(n2764), .ZN(n2831) );
  OR2_X1 U2795 ( .A1(n2052), .A2(n2019), .ZN(n2764) );
  OR2_X1 U2796 ( .A1(n2832), .A2(n2833), .ZN(n2763) );
  AND2_X1 U2797 ( .A1(n2760), .A2(n2759), .ZN(n2833) );
  AND2_X1 U2798 ( .A1(n2757), .A2(n2834), .ZN(n2832) );
  OR2_X1 U2799 ( .A1(n2759), .A2(n2760), .ZN(n2834) );
  OR2_X1 U2800 ( .A1(n2229), .A2(n2019), .ZN(n2760) );
  OR2_X1 U2801 ( .A1(n2835), .A2(n2836), .ZN(n2759) );
  AND2_X1 U2802 ( .A1(n2024), .A2(n2756), .ZN(n2836) );
  AND2_X1 U2803 ( .A1(n2754), .A2(n2837), .ZN(n2835) );
  OR2_X1 U2804 ( .A1(n2756), .A2(n2024), .ZN(n2837) );
  OR2_X1 U2805 ( .A1(n2020), .A2(n2019), .ZN(n2024) );
  OR2_X1 U2806 ( .A1(n2838), .A2(n2839), .ZN(n2756) );
  AND2_X1 U2807 ( .A1(n2753), .A2(n2752), .ZN(n2839) );
  AND2_X1 U2808 ( .A1(n2750), .A2(n2840), .ZN(n2838) );
  OR2_X1 U2809 ( .A1(n2752), .A2(n2753), .ZN(n2840) );
  OR2_X1 U2810 ( .A1(n2234), .A2(n2019), .ZN(n2753) );
  OR2_X1 U2811 ( .A1(n2841), .A2(n2842), .ZN(n2752) );
  AND2_X1 U2812 ( .A1(n2746), .A2(n2749), .ZN(n2842) );
  AND2_X1 U2813 ( .A1(n2843), .A2(n2844), .ZN(n2841) );
  OR2_X1 U2814 ( .A1(n2749), .A2(n2746), .ZN(n2844) );
  OR2_X1 U2815 ( .A1(n1989), .A2(n2019), .ZN(n2746) );
  OR2_X1 U2816 ( .A1(n2019), .A2(n2845), .ZN(n2749) );
  OR2_X1 U2817 ( .A1(n2468), .A2(n2230), .ZN(n2845) );
  INV_X1 U2818 ( .A(b_11_), .ZN(n2019) );
  INV_X1 U2819 ( .A(n2748), .ZN(n2843) );
  OR2_X1 U2820 ( .A1(n2846), .A2(n2847), .ZN(n2748) );
  AND2_X1 U2821 ( .A1(b_9_), .A2(n2848), .ZN(n2847) );
  OR2_X1 U2822 ( .A1(n2849), .A2(n1969), .ZN(n2848) );
  AND2_X1 U2823 ( .A1(a_15_), .A2(n2230), .ZN(n2849) );
  AND2_X1 U2824 ( .A1(b_10_), .A2(n2850), .ZN(n2846) );
  OR2_X1 U2825 ( .A1(n2851), .A2(n1965), .ZN(n2850) );
  AND2_X1 U2826 ( .A1(a_14_), .A2(n2051), .ZN(n2851) );
  XNOR2_X1 U2827 ( .A(n2852), .B(n2853), .ZN(n2750) );
  XOR2_X1 U2828 ( .A(n2854), .B(n2855), .Z(n2853) );
  XOR2_X1 U2829 ( .A(n2856), .B(n2857), .Z(n2754) );
  XOR2_X1 U2830 ( .A(n2858), .B(n2859), .Z(n2857) );
  XOR2_X1 U2831 ( .A(n2860), .B(n2861), .Z(n2757) );
  XOR2_X1 U2832 ( .A(n2862), .B(n2863), .Z(n2861) );
  XOR2_X1 U2833 ( .A(n2864), .B(n2865), .Z(n2761) );
  XOR2_X1 U2834 ( .A(n2866), .B(n2037), .Z(n2865) );
  XOR2_X1 U2835 ( .A(n2867), .B(n2868), .Z(n2765) );
  XOR2_X1 U2836 ( .A(n2869), .B(n2870), .Z(n2868) );
  XOR2_X1 U2837 ( .A(n2871), .B(n2872), .Z(n2769) );
  XOR2_X1 U2838 ( .A(n2873), .B(n2874), .Z(n2872) );
  XOR2_X1 U2839 ( .A(n2875), .B(n2876), .Z(n2773) );
  XOR2_X1 U2840 ( .A(n2877), .B(n2878), .Z(n2876) );
  XOR2_X1 U2841 ( .A(n2879), .B(n2880), .Z(n2777) );
  XOR2_X1 U2842 ( .A(n2881), .B(n2882), .Z(n2880) );
  XOR2_X1 U2843 ( .A(n2883), .B(n2884), .Z(n2781) );
  XOR2_X1 U2844 ( .A(n2885), .B(n2886), .Z(n2884) );
  XOR2_X1 U2845 ( .A(n2887), .B(n2888), .Z(n2785) );
  XOR2_X1 U2846 ( .A(n2889), .B(n2890), .Z(n2888) );
  XOR2_X1 U2847 ( .A(n2891), .B(n2892), .Z(n2789) );
  XOR2_X1 U2848 ( .A(n2893), .B(n2894), .Z(n2892) );
  XOR2_X1 U2849 ( .A(n2895), .B(n2896), .Z(n2793) );
  XOR2_X1 U2850 ( .A(n2897), .B(n2898), .Z(n2896) );
  XOR2_X1 U2851 ( .A(n2899), .B(n2900), .Z(n2797) );
  XOR2_X1 U2852 ( .A(n2901), .B(n2902), .Z(n2900) );
  XNOR2_X1 U2853 ( .A(n2903), .B(n2904), .ZN(n2365) );
  XOR2_X1 U2854 ( .A(n2905), .B(n2906), .Z(n2904) );
  AND2_X1 U2855 ( .A1(n2907), .A2(n2361), .ZN(n2280) );
  OR2_X1 U2856 ( .A1(n2908), .A2(n2909), .ZN(n2361) );
  INV_X1 U2857 ( .A(n2910), .ZN(n2907) );
  AND2_X1 U2858 ( .A1(n2908), .A2(n2909), .ZN(n2910) );
  OR2_X1 U2859 ( .A1(n2911), .A2(n2912), .ZN(n2909) );
  AND2_X1 U2860 ( .A1(n2906), .A2(n2905), .ZN(n2912) );
  AND2_X1 U2861 ( .A1(n2903), .A2(n2913), .ZN(n2911) );
  OR2_X1 U2862 ( .A1(n2906), .A2(n2905), .ZN(n2913) );
  OR2_X1 U2863 ( .A1(n2914), .A2(n2915), .ZN(n2905) );
  AND2_X1 U2864 ( .A1(n2902), .A2(n2901), .ZN(n2915) );
  AND2_X1 U2865 ( .A1(n2899), .A2(n2916), .ZN(n2914) );
  OR2_X1 U2866 ( .A1(n2902), .A2(n2901), .ZN(n2916) );
  OR2_X1 U2867 ( .A1(n2917), .A2(n2918), .ZN(n2901) );
  AND2_X1 U2868 ( .A1(n2898), .A2(n2897), .ZN(n2918) );
  AND2_X1 U2869 ( .A1(n2895), .A2(n2919), .ZN(n2917) );
  OR2_X1 U2870 ( .A1(n2898), .A2(n2897), .ZN(n2919) );
  OR2_X1 U2871 ( .A1(n2920), .A2(n2921), .ZN(n2897) );
  AND2_X1 U2872 ( .A1(n2891), .A2(n2894), .ZN(n2921) );
  AND2_X1 U2873 ( .A1(n2922), .A2(n2893), .ZN(n2920) );
  OR2_X1 U2874 ( .A1(n2923), .A2(n2924), .ZN(n2893) );
  AND2_X1 U2875 ( .A1(n2890), .A2(n2889), .ZN(n2924) );
  AND2_X1 U2876 ( .A1(n2887), .A2(n2925), .ZN(n2923) );
  OR2_X1 U2877 ( .A1(n2890), .A2(n2889), .ZN(n2925) );
  OR2_X1 U2878 ( .A1(n2926), .A2(n2927), .ZN(n2889) );
  AND2_X1 U2879 ( .A1(n2883), .A2(n2886), .ZN(n2927) );
  AND2_X1 U2880 ( .A1(n2928), .A2(n2885), .ZN(n2926) );
  OR2_X1 U2881 ( .A1(n2929), .A2(n2930), .ZN(n2885) );
  AND2_X1 U2882 ( .A1(n2879), .A2(n2882), .ZN(n2930) );
  AND2_X1 U2883 ( .A1(n2931), .A2(n2881), .ZN(n2929) );
  OR2_X1 U2884 ( .A1(n2932), .A2(n2933), .ZN(n2881) );
  AND2_X1 U2885 ( .A1(n2875), .A2(n2878), .ZN(n2933) );
  AND2_X1 U2886 ( .A1(n2934), .A2(n2877), .ZN(n2932) );
  OR2_X1 U2887 ( .A1(n2935), .A2(n2936), .ZN(n2877) );
  AND2_X1 U2888 ( .A1(n2871), .A2(n2874), .ZN(n2936) );
  AND2_X1 U2889 ( .A1(n2937), .A2(n2873), .ZN(n2935) );
  OR2_X1 U2890 ( .A1(n2938), .A2(n2939), .ZN(n2873) );
  AND2_X1 U2891 ( .A1(n2867), .A2(n2870), .ZN(n2939) );
  AND2_X1 U2892 ( .A1(n2940), .A2(n2869), .ZN(n2938) );
  OR2_X1 U2893 ( .A1(n2941), .A2(n2942), .ZN(n2869) );
  AND2_X1 U2894 ( .A1(n2864), .A2(n2037), .ZN(n2942) );
  AND2_X1 U2895 ( .A1(n2943), .A2(n2866), .ZN(n2941) );
  OR2_X1 U2896 ( .A1(n2944), .A2(n2945), .ZN(n2866) );
  AND2_X1 U2897 ( .A1(n2860), .A2(n2863), .ZN(n2945) );
  AND2_X1 U2898 ( .A1(n2946), .A2(n2862), .ZN(n2944) );
  OR2_X1 U2899 ( .A1(n2947), .A2(n2948), .ZN(n2862) );
  AND2_X1 U2900 ( .A1(n2856), .A2(n2859), .ZN(n2948) );
  AND2_X1 U2901 ( .A1(n2949), .A2(n2858), .ZN(n2947) );
  OR2_X1 U2902 ( .A1(n2950), .A2(n2951), .ZN(n2858) );
  AND2_X1 U2903 ( .A1(n2852), .A2(n2855), .ZN(n2951) );
  AND2_X1 U2904 ( .A1(n2952), .A2(n2953), .ZN(n2950) );
  OR2_X1 U2905 ( .A1(n2852), .A2(n2855), .ZN(n2953) );
  OR2_X1 U2906 ( .A1(n2230), .A2(n2954), .ZN(n2855) );
  OR2_X1 U2907 ( .A1(n2468), .A2(n2051), .ZN(n2954) );
  OR2_X1 U2908 ( .A1(n1989), .A2(n2230), .ZN(n2852) );
  INV_X1 U2909 ( .A(n2854), .ZN(n2952) );
  OR2_X1 U2910 ( .A1(n2955), .A2(n2956), .ZN(n2854) );
  AND2_X1 U2911 ( .A1(b_9_), .A2(n2957), .ZN(n2956) );
  OR2_X1 U2912 ( .A1(n2958), .A2(n1965), .ZN(n2957) );
  AND2_X1 U2913 ( .A1(a_14_), .A2(n2225), .ZN(n2958) );
  AND2_X1 U2914 ( .A1(b_8_), .A2(n2959), .ZN(n2955) );
  OR2_X1 U2915 ( .A1(n2960), .A2(n1969), .ZN(n2959) );
  AND2_X1 U2916 ( .A1(a_15_), .A2(n2051), .ZN(n2960) );
  OR2_X1 U2917 ( .A1(n2856), .A2(n2859), .ZN(n2949) );
  OR2_X1 U2918 ( .A1(n2234), .A2(n2230), .ZN(n2859) );
  XNOR2_X1 U2919 ( .A(n2961), .B(n2962), .ZN(n2856) );
  XOR2_X1 U2920 ( .A(n2963), .B(n2964), .Z(n2962) );
  OR2_X1 U2921 ( .A1(n2860), .A2(n2863), .ZN(n2946) );
  OR2_X1 U2922 ( .A1(n2020), .A2(n2230), .ZN(n2863) );
  XOR2_X1 U2923 ( .A(n2965), .B(n2966), .Z(n2860) );
  XOR2_X1 U2924 ( .A(n2967), .B(n2968), .Z(n2966) );
  OR2_X1 U2925 ( .A1(n2864), .A2(n2037), .ZN(n2943) );
  OR2_X1 U2926 ( .A1(n2229), .A2(n2230), .ZN(n2037) );
  XOR2_X1 U2927 ( .A(n2969), .B(n2970), .Z(n2864) );
  XOR2_X1 U2928 ( .A(n2971), .B(n2972), .Z(n2970) );
  OR2_X1 U2929 ( .A1(n2867), .A2(n2870), .ZN(n2940) );
  OR2_X1 U2930 ( .A1(n2052), .A2(n2230), .ZN(n2870) );
  XOR2_X1 U2931 ( .A(n2973), .B(n2974), .Z(n2867) );
  XOR2_X1 U2932 ( .A(n2975), .B(n2976), .Z(n2974) );
  OR2_X1 U2933 ( .A1(n2871), .A2(n2874), .ZN(n2937) );
  OR2_X1 U2934 ( .A1(n2224), .A2(n2230), .ZN(n2874) );
  XOR2_X1 U2935 ( .A(n2977), .B(n2978), .Z(n2871) );
  XOR2_X1 U2936 ( .A(n2979), .B(n2056), .Z(n2978) );
  OR2_X1 U2937 ( .A1(n2875), .A2(n2878), .ZN(n2934) );
  OR2_X1 U2938 ( .A1(n2084), .A2(n2230), .ZN(n2878) );
  XOR2_X1 U2939 ( .A(n2980), .B(n2981), .Z(n2875) );
  XOR2_X1 U2940 ( .A(n2982), .B(n2983), .Z(n2981) );
  OR2_X1 U2941 ( .A1(n2879), .A2(n2882), .ZN(n2931) );
  OR2_X1 U2942 ( .A1(n2219), .A2(n2230), .ZN(n2882) );
  XOR2_X1 U2943 ( .A(n2984), .B(n2985), .Z(n2879) );
  XOR2_X1 U2944 ( .A(n2986), .B(n2987), .Z(n2985) );
  OR2_X1 U2945 ( .A1(n2883), .A2(n2886), .ZN(n2928) );
  OR2_X1 U2946 ( .A1(n2116), .A2(n2230), .ZN(n2886) );
  XOR2_X1 U2947 ( .A(n2988), .B(n2989), .Z(n2883) );
  XOR2_X1 U2948 ( .A(n2990), .B(n2991), .Z(n2989) );
  OR2_X1 U2949 ( .A1(n2214), .A2(n2230), .ZN(n2890) );
  XOR2_X1 U2950 ( .A(n2992), .B(n2993), .Z(n2887) );
  XOR2_X1 U2951 ( .A(n2994), .B(n2995), .Z(n2993) );
  OR2_X1 U2952 ( .A1(n2891), .A2(n2894), .ZN(n2922) );
  OR2_X1 U2953 ( .A1(n2158), .A2(n2230), .ZN(n2894) );
  XOR2_X1 U2954 ( .A(n2996), .B(n2997), .Z(n2891) );
  XOR2_X1 U2955 ( .A(n2998), .B(n2999), .Z(n2997) );
  OR2_X1 U2956 ( .A1(n2209), .A2(n2230), .ZN(n2898) );
  XOR2_X1 U2957 ( .A(n3000), .B(n3001), .Z(n2895) );
  XOR2_X1 U2958 ( .A(n3002), .B(n3003), .Z(n3001) );
  OR2_X1 U2959 ( .A1(n2190), .A2(n2230), .ZN(n2902) );
  XOR2_X1 U2960 ( .A(n3004), .B(n3005), .Z(n2899) );
  XOR2_X1 U2961 ( .A(n3006), .B(n3007), .Z(n3005) );
  OR2_X1 U2962 ( .A1(n2205), .A2(n2230), .ZN(n2906) );
  INV_X1 U2963 ( .A(b_10_), .ZN(n2230) );
  XOR2_X1 U2964 ( .A(n3008), .B(n3009), .Z(n2903) );
  XOR2_X1 U2965 ( .A(n3010), .B(n3011), .Z(n3009) );
  XOR2_X1 U2966 ( .A(n3012), .B(n3013), .Z(n2908) );
  XOR2_X1 U2967 ( .A(n3014), .B(n3015), .Z(n3013) );
  OR2_X1 U2968 ( .A1(n2358), .A2(n2359), .ZN(n2354) );
  OR2_X1 U2969 ( .A1(n3016), .A2(n3017), .ZN(n2359) );
  AND2_X1 U2970 ( .A1(n3015), .A2(n3014), .ZN(n3017) );
  AND2_X1 U2971 ( .A1(n3012), .A2(n3018), .ZN(n3016) );
  OR2_X1 U2972 ( .A1(n3015), .A2(n3014), .ZN(n3018) );
  OR2_X1 U2973 ( .A1(n3019), .A2(n3020), .ZN(n3014) );
  AND2_X1 U2974 ( .A1(n3011), .A2(n3010), .ZN(n3020) );
  AND2_X1 U2975 ( .A1(n3008), .A2(n3021), .ZN(n3019) );
  OR2_X1 U2976 ( .A1(n3011), .A2(n3010), .ZN(n3021) );
  OR2_X1 U2977 ( .A1(n3022), .A2(n3023), .ZN(n3010) );
  AND2_X1 U2978 ( .A1(n3007), .A2(n3006), .ZN(n3023) );
  AND2_X1 U2979 ( .A1(n3004), .A2(n3024), .ZN(n3022) );
  OR2_X1 U2980 ( .A1(n3007), .A2(n3006), .ZN(n3024) );
  OR2_X1 U2981 ( .A1(n3025), .A2(n3026), .ZN(n3006) );
  AND2_X1 U2982 ( .A1(n3003), .A2(n3002), .ZN(n3026) );
  AND2_X1 U2983 ( .A1(n3000), .A2(n3027), .ZN(n3025) );
  OR2_X1 U2984 ( .A1(n3003), .A2(n3002), .ZN(n3027) );
  OR2_X1 U2985 ( .A1(n3028), .A2(n3029), .ZN(n3002) );
  AND2_X1 U2986 ( .A1(n2996), .A2(n2999), .ZN(n3029) );
  AND2_X1 U2987 ( .A1(n3030), .A2(n2998), .ZN(n3028) );
  OR2_X1 U2988 ( .A1(n3031), .A2(n3032), .ZN(n2998) );
  AND2_X1 U2989 ( .A1(n2995), .A2(n2994), .ZN(n3032) );
  AND2_X1 U2990 ( .A1(n2992), .A2(n3033), .ZN(n3031) );
  OR2_X1 U2991 ( .A1(n2995), .A2(n2994), .ZN(n3033) );
  OR2_X1 U2992 ( .A1(n3034), .A2(n3035), .ZN(n2994) );
  AND2_X1 U2993 ( .A1(n2988), .A2(n2991), .ZN(n3035) );
  AND2_X1 U2994 ( .A1(n3036), .A2(n2990), .ZN(n3034) );
  OR2_X1 U2995 ( .A1(n3037), .A2(n3038), .ZN(n2990) );
  AND2_X1 U2996 ( .A1(n2984), .A2(n2987), .ZN(n3038) );
  AND2_X1 U2997 ( .A1(n3039), .A2(n2986), .ZN(n3037) );
  OR2_X1 U2998 ( .A1(n3040), .A2(n3041), .ZN(n2986) );
  AND2_X1 U2999 ( .A1(n2980), .A2(n2983), .ZN(n3041) );
  AND2_X1 U3000 ( .A1(n3042), .A2(n2982), .ZN(n3040) );
  OR2_X1 U3001 ( .A1(n3043), .A2(n3044), .ZN(n2982) );
  AND2_X1 U3002 ( .A1(n2977), .A2(n2056), .ZN(n3044) );
  AND2_X1 U3003 ( .A1(n3045), .A2(n2979), .ZN(n3043) );
  OR2_X1 U3004 ( .A1(n3046), .A2(n3047), .ZN(n2979) );
  AND2_X1 U3005 ( .A1(n2973), .A2(n2976), .ZN(n3047) );
  AND2_X1 U3006 ( .A1(n3048), .A2(n2975), .ZN(n3046) );
  OR2_X1 U3007 ( .A1(n3049), .A2(n3050), .ZN(n2975) );
  AND2_X1 U3008 ( .A1(n2969), .A2(n2972), .ZN(n3050) );
  AND2_X1 U3009 ( .A1(n3051), .A2(n2971), .ZN(n3049) );
  OR2_X1 U3010 ( .A1(n3052), .A2(n3053), .ZN(n2971) );
  AND2_X1 U3011 ( .A1(n2965), .A2(n2968), .ZN(n3053) );
  AND2_X1 U3012 ( .A1(n3054), .A2(n2967), .ZN(n3052) );
  OR2_X1 U3013 ( .A1(n3055), .A2(n3056), .ZN(n2967) );
  AND2_X1 U3014 ( .A1(n2961), .A2(n2964), .ZN(n3056) );
  AND2_X1 U3015 ( .A1(n3057), .A2(n3058), .ZN(n3055) );
  OR2_X1 U3016 ( .A1(n2961), .A2(n2964), .ZN(n3058) );
  OR2_X1 U3017 ( .A1(n2051), .A2(n3059), .ZN(n2964) );
  OR2_X1 U3018 ( .A1(n2225), .A2(n2468), .ZN(n3059) );
  OR2_X1 U3019 ( .A1(n2051), .A2(n1989), .ZN(n2961) );
  INV_X1 U3020 ( .A(n2963), .ZN(n3057) );
  OR2_X1 U3021 ( .A1(n3060), .A2(n3061), .ZN(n2963) );
  AND2_X1 U3022 ( .A1(b_8_), .A2(n3062), .ZN(n3061) );
  OR2_X1 U3023 ( .A1(n3063), .A2(n1965), .ZN(n3062) );
  AND2_X1 U3024 ( .A1(a_14_), .A2(n2083), .ZN(n3063) );
  AND2_X1 U3025 ( .A1(b_7_), .A2(n3064), .ZN(n3060) );
  OR2_X1 U3026 ( .A1(n3065), .A2(n1969), .ZN(n3064) );
  AND2_X1 U3027 ( .A1(a_15_), .A2(n2225), .ZN(n3065) );
  OR2_X1 U3028 ( .A1(n2965), .A2(n2968), .ZN(n3054) );
  OR2_X1 U3029 ( .A1(n2051), .A2(n2234), .ZN(n2968) );
  XNOR2_X1 U3030 ( .A(n3066), .B(n3067), .ZN(n2965) );
  XOR2_X1 U3031 ( .A(n3068), .B(n3069), .Z(n3067) );
  OR2_X1 U3032 ( .A1(n2969), .A2(n2972), .ZN(n3051) );
  OR2_X1 U3033 ( .A1(n2051), .A2(n2020), .ZN(n2972) );
  XNOR2_X1 U3034 ( .A(n3070), .B(n3071), .ZN(n2969) );
  XNOR2_X1 U3035 ( .A(n3072), .B(n3073), .ZN(n3070) );
  OR2_X1 U3036 ( .A1(n2973), .A2(n2976), .ZN(n3048) );
  OR2_X1 U3037 ( .A1(n2051), .A2(n2229), .ZN(n2976) );
  XOR2_X1 U3038 ( .A(n3074), .B(n3075), .Z(n2973) );
  XOR2_X1 U3039 ( .A(n3076), .B(n3077), .Z(n3075) );
  OR2_X1 U3040 ( .A1(n2977), .A2(n2056), .ZN(n3045) );
  OR2_X1 U3041 ( .A1(n2051), .A2(n2052), .ZN(n2056) );
  XOR2_X1 U3042 ( .A(n3078), .B(n3079), .Z(n2977) );
  XOR2_X1 U3043 ( .A(n3080), .B(n3081), .Z(n3079) );
  OR2_X1 U3044 ( .A1(n2980), .A2(n2983), .ZN(n3042) );
  OR2_X1 U3045 ( .A1(n2051), .A2(n2224), .ZN(n2983) );
  XOR2_X1 U3046 ( .A(n3082), .B(n3083), .Z(n2980) );
  XOR2_X1 U3047 ( .A(n3084), .B(n3085), .Z(n3083) );
  OR2_X1 U3048 ( .A1(n2984), .A2(n2987), .ZN(n3039) );
  OR2_X1 U3049 ( .A1(n2051), .A2(n2084), .ZN(n2987) );
  XOR2_X1 U3050 ( .A(n3086), .B(n3087), .Z(n2984) );
  XOR2_X1 U3051 ( .A(n3088), .B(n2069), .Z(n3087) );
  OR2_X1 U3052 ( .A1(n2988), .A2(n2991), .ZN(n3036) );
  OR2_X1 U3053 ( .A1(n2051), .A2(n2219), .ZN(n2991) );
  XOR2_X1 U3054 ( .A(n3089), .B(n3090), .Z(n2988) );
  XOR2_X1 U3055 ( .A(n3091), .B(n3092), .Z(n3090) );
  OR2_X1 U3056 ( .A1(n2051), .A2(n2116), .ZN(n2995) );
  XOR2_X1 U3057 ( .A(n3093), .B(n3094), .Z(n2992) );
  XOR2_X1 U3058 ( .A(n3095), .B(n3096), .Z(n3094) );
  OR2_X1 U3059 ( .A1(n2996), .A2(n2999), .ZN(n3030) );
  OR2_X1 U3060 ( .A1(n2051), .A2(n2214), .ZN(n2999) );
  XOR2_X1 U3061 ( .A(n3097), .B(n3098), .Z(n2996) );
  XOR2_X1 U3062 ( .A(n3099), .B(n3100), .Z(n3098) );
  OR2_X1 U3063 ( .A1(n2051), .A2(n2158), .ZN(n3003) );
  XOR2_X1 U3064 ( .A(n3101), .B(n3102), .Z(n3000) );
  XOR2_X1 U3065 ( .A(n3103), .B(n3104), .Z(n3102) );
  OR2_X1 U3066 ( .A1(n2051), .A2(n2209), .ZN(n3007) );
  XOR2_X1 U3067 ( .A(n3105), .B(n3106), .Z(n3004) );
  XOR2_X1 U3068 ( .A(n3107), .B(n3108), .Z(n3106) );
  OR2_X1 U3069 ( .A1(n2051), .A2(n2190), .ZN(n3011) );
  XOR2_X1 U3070 ( .A(n3109), .B(n3110), .Z(n3008) );
  XOR2_X1 U3071 ( .A(n3111), .B(n3112), .Z(n3110) );
  OR2_X1 U3072 ( .A1(n2051), .A2(n2205), .ZN(n3015) );
  INV_X1 U3073 ( .A(b_9_), .ZN(n2051) );
  XOR2_X1 U3074 ( .A(n3113), .B(n3114), .Z(n3012) );
  XOR2_X1 U3075 ( .A(n3115), .B(n3116), .Z(n3114) );
  XOR2_X1 U3076 ( .A(n2348), .B(n3117), .Z(n2358) );
  XOR2_X1 U3077 ( .A(n2347), .B(n2346), .Z(n3117) );
  OR2_X1 U3078 ( .A1(n2225), .A2(n2205), .ZN(n2346) );
  OR2_X1 U3079 ( .A1(n3118), .A2(n3119), .ZN(n2347) );
  AND2_X1 U3080 ( .A1(n3116), .A2(n3115), .ZN(n3119) );
  AND2_X1 U3081 ( .A1(n3113), .A2(n3120), .ZN(n3118) );
  OR2_X1 U3082 ( .A1(n3115), .A2(n3116), .ZN(n3120) );
  OR2_X1 U3083 ( .A1(n2225), .A2(n2190), .ZN(n3116) );
  OR2_X1 U3084 ( .A1(n3121), .A2(n3122), .ZN(n3115) );
  AND2_X1 U3085 ( .A1(n3112), .A2(n3111), .ZN(n3122) );
  AND2_X1 U3086 ( .A1(n3109), .A2(n3123), .ZN(n3121) );
  OR2_X1 U3087 ( .A1(n3111), .A2(n3112), .ZN(n3123) );
  OR2_X1 U3088 ( .A1(n2225), .A2(n2209), .ZN(n3112) );
  OR2_X1 U3089 ( .A1(n3124), .A2(n3125), .ZN(n3111) );
  AND2_X1 U3090 ( .A1(n3108), .A2(n3107), .ZN(n3125) );
  AND2_X1 U3091 ( .A1(n3105), .A2(n3126), .ZN(n3124) );
  OR2_X1 U3092 ( .A1(n3107), .A2(n3108), .ZN(n3126) );
  OR2_X1 U3093 ( .A1(n2225), .A2(n2158), .ZN(n3108) );
  OR2_X1 U3094 ( .A1(n3127), .A2(n3128), .ZN(n3107) );
  AND2_X1 U3095 ( .A1(n3104), .A2(n3103), .ZN(n3128) );
  AND2_X1 U3096 ( .A1(n3101), .A2(n3129), .ZN(n3127) );
  OR2_X1 U3097 ( .A1(n3103), .A2(n3104), .ZN(n3129) );
  OR2_X1 U3098 ( .A1(n2225), .A2(n2214), .ZN(n3104) );
  OR2_X1 U3099 ( .A1(n3130), .A2(n3131), .ZN(n3103) );
  AND2_X1 U3100 ( .A1(n3097), .A2(n3100), .ZN(n3131) );
  AND2_X1 U3101 ( .A1(n3132), .A2(n3099), .ZN(n3130) );
  OR2_X1 U3102 ( .A1(n3133), .A2(n3134), .ZN(n3099) );
  AND2_X1 U3103 ( .A1(n3096), .A2(n3095), .ZN(n3134) );
  AND2_X1 U3104 ( .A1(n3093), .A2(n3135), .ZN(n3133) );
  OR2_X1 U3105 ( .A1(n3095), .A2(n3096), .ZN(n3135) );
  OR2_X1 U3106 ( .A1(n2225), .A2(n2219), .ZN(n3096) );
  OR2_X1 U3107 ( .A1(n3136), .A2(n3137), .ZN(n3095) );
  AND2_X1 U3108 ( .A1(n3089), .A2(n3092), .ZN(n3137) );
  AND2_X1 U3109 ( .A1(n3138), .A2(n3091), .ZN(n3136) );
  OR2_X1 U3110 ( .A1(n3139), .A2(n3140), .ZN(n3091) );
  AND2_X1 U3111 ( .A1(n3086), .A2(n2069), .ZN(n3140) );
  AND2_X1 U3112 ( .A1(n3141), .A2(n3088), .ZN(n3139) );
  OR2_X1 U3113 ( .A1(n3142), .A2(n3143), .ZN(n3088) );
  AND2_X1 U3114 ( .A1(n3082), .A2(n3085), .ZN(n3143) );
  AND2_X1 U3115 ( .A1(n3144), .A2(n3084), .ZN(n3142) );
  OR2_X1 U3116 ( .A1(n3145), .A2(n3146), .ZN(n3084) );
  AND2_X1 U3117 ( .A1(n3078), .A2(n3081), .ZN(n3146) );
  AND2_X1 U3118 ( .A1(n3147), .A2(n3080), .ZN(n3145) );
  OR2_X1 U3119 ( .A1(n3148), .A2(n3149), .ZN(n3080) );
  AND2_X1 U3120 ( .A1(n3074), .A2(n3077), .ZN(n3149) );
  AND2_X1 U3121 ( .A1(n3150), .A2(n3076), .ZN(n3148) );
  OR2_X1 U3122 ( .A1(n3151), .A2(n3152), .ZN(n3076) );
  AND2_X1 U3123 ( .A1(n3071), .A2(n3073), .ZN(n3152) );
  AND2_X1 U3124 ( .A1(n3153), .A2(n3072), .ZN(n3151) );
  OR2_X1 U3125 ( .A1(n3154), .A2(n3155), .ZN(n3072) );
  AND2_X1 U3126 ( .A1(n3066), .A2(n3069), .ZN(n3155) );
  AND2_X1 U3127 ( .A1(n3156), .A2(n3157), .ZN(n3154) );
  OR2_X1 U3128 ( .A1(n3069), .A2(n3066), .ZN(n3157) );
  OR2_X1 U3129 ( .A1(n2225), .A2(n1989), .ZN(n3066) );
  OR2_X1 U3130 ( .A1(n2468), .A2(n3158), .ZN(n3069) );
  OR2_X1 U3131 ( .A1(n2083), .A2(n2225), .ZN(n3158) );
  INV_X1 U3132 ( .A(n3068), .ZN(n3156) );
  OR2_X1 U3133 ( .A1(n3159), .A2(n3160), .ZN(n3068) );
  AND2_X1 U3134 ( .A1(b_7_), .A2(n3161), .ZN(n3160) );
  OR2_X1 U3135 ( .A1(n3162), .A2(n1965), .ZN(n3161) );
  AND2_X1 U3136 ( .A1(a_14_), .A2(n2220), .ZN(n3162) );
  AND2_X1 U3137 ( .A1(b_6_), .A2(n3163), .ZN(n3159) );
  OR2_X1 U3138 ( .A1(n3164), .A2(n1969), .ZN(n3163) );
  AND2_X1 U3139 ( .A1(a_15_), .A2(n2083), .ZN(n3164) );
  OR2_X1 U3140 ( .A1(n3073), .A2(n3071), .ZN(n3153) );
  XNOR2_X1 U3141 ( .A(n3165), .B(n3166), .ZN(n3071) );
  XOR2_X1 U3142 ( .A(n3167), .B(n3168), .Z(n3166) );
  OR2_X1 U3143 ( .A1(n2225), .A2(n2234), .ZN(n3073) );
  OR2_X1 U3144 ( .A1(n3077), .A2(n3074), .ZN(n3150) );
  XOR2_X1 U3145 ( .A(n3169), .B(n3170), .Z(n3074) );
  XOR2_X1 U3146 ( .A(n3171), .B(n3172), .Z(n3170) );
  OR2_X1 U3147 ( .A1(n2225), .A2(n2020), .ZN(n3077) );
  OR2_X1 U3148 ( .A1(n3081), .A2(n3078), .ZN(n3147) );
  XOR2_X1 U3149 ( .A(n3173), .B(n3174), .Z(n3078) );
  XOR2_X1 U3150 ( .A(n3175), .B(n3176), .Z(n3174) );
  OR2_X1 U3151 ( .A1(n2225), .A2(n2229), .ZN(n3081) );
  OR2_X1 U3152 ( .A1(n3085), .A2(n3082), .ZN(n3144) );
  XOR2_X1 U3153 ( .A(n3177), .B(n3178), .Z(n3082) );
  XOR2_X1 U3154 ( .A(n3179), .B(n3180), .Z(n3178) );
  OR2_X1 U3155 ( .A1(n2225), .A2(n2052), .ZN(n3085) );
  OR2_X1 U3156 ( .A1(n2069), .A2(n3086), .ZN(n3141) );
  XOR2_X1 U3157 ( .A(n3181), .B(n3182), .Z(n3086) );
  XOR2_X1 U3158 ( .A(n3183), .B(n3184), .Z(n3182) );
  OR2_X1 U3159 ( .A1(n2225), .A2(n2224), .ZN(n2069) );
  OR2_X1 U3160 ( .A1(n3092), .A2(n3089), .ZN(n3138) );
  XOR2_X1 U3161 ( .A(n3185), .B(n3186), .Z(n3089) );
  XOR2_X1 U3162 ( .A(n3187), .B(n3188), .Z(n3186) );
  OR2_X1 U3163 ( .A1(n2225), .A2(n2084), .ZN(n3092) );
  XOR2_X1 U3164 ( .A(n3189), .B(n3190), .Z(n3093) );
  XOR2_X1 U3165 ( .A(n3191), .B(n2088), .Z(n3190) );
  OR2_X1 U3166 ( .A1(n3100), .A2(n3097), .ZN(n3132) );
  XOR2_X1 U3167 ( .A(n3192), .B(n3193), .Z(n3097) );
  XOR2_X1 U3168 ( .A(n3194), .B(n3195), .Z(n3193) );
  OR2_X1 U3169 ( .A1(n2225), .A2(n2116), .ZN(n3100) );
  INV_X1 U3170 ( .A(b_8_), .ZN(n2225) );
  XOR2_X1 U3171 ( .A(n3196), .B(n3197), .Z(n3101) );
  XOR2_X1 U3172 ( .A(n3198), .B(n3199), .Z(n3197) );
  XOR2_X1 U3173 ( .A(n3200), .B(n3201), .Z(n3105) );
  XOR2_X1 U3174 ( .A(n3202), .B(n3203), .Z(n3201) );
  XOR2_X1 U3175 ( .A(n3204), .B(n3205), .Z(n3109) );
  XOR2_X1 U3176 ( .A(n3206), .B(n3207), .Z(n3205) );
  XOR2_X1 U3177 ( .A(n3208), .B(n3209), .Z(n3113) );
  XOR2_X1 U3178 ( .A(n3210), .B(n3211), .Z(n3209) );
  XOR2_X1 U3179 ( .A(n3212), .B(n3213), .Z(n2348) );
  XOR2_X1 U3180 ( .A(n3214), .B(n3215), .Z(n3213) );
  OR2_X1 U3181 ( .A1(n2336), .A2(n2337), .ZN(n2332) );
  OR2_X1 U3182 ( .A1(n3216), .A2(n3217), .ZN(n2337) );
  AND2_X1 U3183 ( .A1(n2353), .A2(n2352), .ZN(n3217) );
  AND2_X1 U3184 ( .A1(n2350), .A2(n3218), .ZN(n3216) );
  OR2_X1 U3185 ( .A1(n2352), .A2(n2353), .ZN(n3218) );
  OR2_X1 U3186 ( .A1(n2083), .A2(n2205), .ZN(n2353) );
  OR2_X1 U3187 ( .A1(n3219), .A2(n3220), .ZN(n2352) );
  AND2_X1 U3188 ( .A1(n3215), .A2(n3214), .ZN(n3220) );
  AND2_X1 U3189 ( .A1(n3212), .A2(n3221), .ZN(n3219) );
  OR2_X1 U3190 ( .A1(n3214), .A2(n3215), .ZN(n3221) );
  OR2_X1 U3191 ( .A1(n2083), .A2(n2190), .ZN(n3215) );
  OR2_X1 U3192 ( .A1(n3222), .A2(n3223), .ZN(n3214) );
  AND2_X1 U3193 ( .A1(n3211), .A2(n3210), .ZN(n3223) );
  AND2_X1 U3194 ( .A1(n3208), .A2(n3224), .ZN(n3222) );
  OR2_X1 U3195 ( .A1(n3210), .A2(n3211), .ZN(n3224) );
  OR2_X1 U3196 ( .A1(n2083), .A2(n2209), .ZN(n3211) );
  OR2_X1 U3197 ( .A1(n3225), .A2(n3226), .ZN(n3210) );
  AND2_X1 U3198 ( .A1(n3207), .A2(n3206), .ZN(n3226) );
  AND2_X1 U3199 ( .A1(n3204), .A2(n3227), .ZN(n3225) );
  OR2_X1 U3200 ( .A1(n3206), .A2(n3207), .ZN(n3227) );
  OR2_X1 U3201 ( .A1(n2083), .A2(n2158), .ZN(n3207) );
  OR2_X1 U3202 ( .A1(n3228), .A2(n3229), .ZN(n3206) );
  AND2_X1 U3203 ( .A1(n3203), .A2(n3202), .ZN(n3229) );
  AND2_X1 U3204 ( .A1(n3200), .A2(n3230), .ZN(n3228) );
  OR2_X1 U3205 ( .A1(n3202), .A2(n3203), .ZN(n3230) );
  OR2_X1 U3206 ( .A1(n2083), .A2(n2214), .ZN(n3203) );
  OR2_X1 U3207 ( .A1(n3231), .A2(n3232), .ZN(n3202) );
  AND2_X1 U3208 ( .A1(n3199), .A2(n3198), .ZN(n3232) );
  AND2_X1 U3209 ( .A1(n3196), .A2(n3233), .ZN(n3231) );
  OR2_X1 U3210 ( .A1(n3198), .A2(n3199), .ZN(n3233) );
  OR2_X1 U3211 ( .A1(n2083), .A2(n2116), .ZN(n3199) );
  OR2_X1 U3212 ( .A1(n3234), .A2(n3235), .ZN(n3198) );
  AND2_X1 U3213 ( .A1(n3192), .A2(n3195), .ZN(n3235) );
  AND2_X1 U3214 ( .A1(n3236), .A2(n3194), .ZN(n3234) );
  OR2_X1 U3215 ( .A1(n3237), .A2(n3238), .ZN(n3194) );
  AND2_X1 U3216 ( .A1(n2088), .A2(n3191), .ZN(n3238) );
  AND2_X1 U3217 ( .A1(n3189), .A2(n3239), .ZN(n3237) );
  OR2_X1 U3218 ( .A1(n3191), .A2(n2088), .ZN(n3239) );
  OR2_X1 U3219 ( .A1(n2083), .A2(n2084), .ZN(n2088) );
  OR2_X1 U3220 ( .A1(n3240), .A2(n3241), .ZN(n3191) );
  AND2_X1 U3221 ( .A1(n3185), .A2(n3188), .ZN(n3241) );
  AND2_X1 U3222 ( .A1(n3242), .A2(n3187), .ZN(n3240) );
  OR2_X1 U3223 ( .A1(n3243), .A2(n3244), .ZN(n3187) );
  AND2_X1 U3224 ( .A1(n3181), .A2(n3184), .ZN(n3244) );
  AND2_X1 U3225 ( .A1(n3245), .A2(n3183), .ZN(n3243) );
  OR2_X1 U3226 ( .A1(n3246), .A2(n3247), .ZN(n3183) );
  AND2_X1 U3227 ( .A1(n3177), .A2(n3180), .ZN(n3247) );
  AND2_X1 U3228 ( .A1(n3248), .A2(n3179), .ZN(n3246) );
  OR2_X1 U3229 ( .A1(n3249), .A2(n3250), .ZN(n3179) );
  AND2_X1 U3230 ( .A1(n3173), .A2(n3176), .ZN(n3250) );
  AND2_X1 U3231 ( .A1(n3251), .A2(n3175), .ZN(n3249) );
  OR2_X1 U3232 ( .A1(n3252), .A2(n3253), .ZN(n3175) );
  AND2_X1 U3233 ( .A1(n3169), .A2(n3172), .ZN(n3253) );
  AND2_X1 U3234 ( .A1(n3254), .A2(n3171), .ZN(n3252) );
  OR2_X1 U3235 ( .A1(n3255), .A2(n3256), .ZN(n3171) );
  AND2_X1 U3236 ( .A1(n3165), .A2(n3168), .ZN(n3256) );
  AND2_X1 U3237 ( .A1(n3257), .A2(n3258), .ZN(n3255) );
  OR2_X1 U3238 ( .A1(n3168), .A2(n3165), .ZN(n3258) );
  OR2_X1 U3239 ( .A1(n2083), .A2(n1989), .ZN(n3165) );
  OR2_X1 U3240 ( .A1(n2220), .A2(n3259), .ZN(n3168) );
  OR2_X1 U3241 ( .A1(n2083), .A2(n2468), .ZN(n3259) );
  INV_X1 U3242 ( .A(n3167), .ZN(n3257) );
  OR2_X1 U3243 ( .A1(n3260), .A2(n3261), .ZN(n3167) );
  AND2_X1 U3244 ( .A1(b_6_), .A2(n3262), .ZN(n3261) );
  OR2_X1 U3245 ( .A1(n3263), .A2(n1965), .ZN(n3262) );
  AND2_X1 U3246 ( .A1(a_14_), .A2(n2115), .ZN(n3263) );
  AND2_X1 U3247 ( .A1(b_5_), .A2(n3264), .ZN(n3260) );
  OR2_X1 U3248 ( .A1(n3265), .A2(n1969), .ZN(n3264) );
  AND2_X1 U3249 ( .A1(a_15_), .A2(n2220), .ZN(n3265) );
  OR2_X1 U3250 ( .A1(n3172), .A2(n3169), .ZN(n3254) );
  XNOR2_X1 U3251 ( .A(n3266), .B(n3267), .ZN(n3169) );
  XOR2_X1 U3252 ( .A(n3268), .B(n3269), .Z(n3267) );
  OR2_X1 U3253 ( .A1(n2083), .A2(n2234), .ZN(n3172) );
  OR2_X1 U3254 ( .A1(n3176), .A2(n3173), .ZN(n3251) );
  XOR2_X1 U3255 ( .A(n3270), .B(n3271), .Z(n3173) );
  XOR2_X1 U3256 ( .A(n3272), .B(n3273), .Z(n3271) );
  OR2_X1 U3257 ( .A1(n2083), .A2(n2020), .ZN(n3176) );
  OR2_X1 U3258 ( .A1(n3180), .A2(n3177), .ZN(n3248) );
  XOR2_X1 U3259 ( .A(n3274), .B(n3275), .Z(n3177) );
  XOR2_X1 U3260 ( .A(n3276), .B(n3277), .Z(n3275) );
  OR2_X1 U3261 ( .A1(n2083), .A2(n2229), .ZN(n3180) );
  OR2_X1 U3262 ( .A1(n3184), .A2(n3181), .ZN(n3245) );
  XOR2_X1 U3263 ( .A(n3278), .B(n3279), .Z(n3181) );
  XOR2_X1 U3264 ( .A(n3280), .B(n3281), .Z(n3279) );
  OR2_X1 U3265 ( .A1(n2083), .A2(n2052), .ZN(n3184) );
  OR2_X1 U3266 ( .A1(n3188), .A2(n3185), .ZN(n3242) );
  XOR2_X1 U3267 ( .A(n3282), .B(n3283), .Z(n3185) );
  XOR2_X1 U3268 ( .A(n3284), .B(n3285), .Z(n3283) );
  OR2_X1 U3269 ( .A1(n2083), .A2(n2224), .ZN(n3188) );
  XOR2_X1 U3270 ( .A(n3286), .B(n3287), .Z(n3189) );
  XOR2_X1 U3271 ( .A(n3288), .B(n3289), .Z(n3287) );
  OR2_X1 U3272 ( .A1(n3195), .A2(n3192), .ZN(n3236) );
  XOR2_X1 U3273 ( .A(n3290), .B(n3291), .Z(n3192) );
  XOR2_X1 U3274 ( .A(n3292), .B(n3293), .Z(n3291) );
  OR2_X1 U3275 ( .A1(n2083), .A2(n2219), .ZN(n3195) );
  INV_X1 U3276 ( .A(b_7_), .ZN(n2083) );
  XOR2_X1 U3277 ( .A(n3294), .B(n3295), .Z(n3196) );
  XOR2_X1 U3278 ( .A(n3296), .B(n2101), .Z(n3295) );
  XOR2_X1 U3279 ( .A(n3297), .B(n3298), .Z(n3200) );
  XOR2_X1 U3280 ( .A(n3299), .B(n3300), .Z(n3298) );
  XOR2_X1 U3281 ( .A(n3301), .B(n3302), .Z(n3204) );
  XOR2_X1 U3282 ( .A(n3303), .B(n3304), .Z(n3302) );
  XOR2_X1 U3283 ( .A(n3305), .B(n3306), .Z(n3208) );
  XOR2_X1 U3284 ( .A(n3307), .B(n3308), .Z(n3306) );
  XOR2_X1 U3285 ( .A(n3309), .B(n3310), .Z(n3212) );
  XOR2_X1 U3286 ( .A(n3311), .B(n3312), .Z(n3310) );
  XOR2_X1 U3287 ( .A(n3313), .B(n3314), .Z(n2350) );
  XOR2_X1 U3288 ( .A(n3315), .B(n3316), .Z(n3314) );
  XOR2_X1 U3289 ( .A(n2326), .B(n3317), .Z(n2336) );
  XOR2_X1 U3290 ( .A(n2325), .B(n2324), .Z(n3317) );
  OR2_X1 U3291 ( .A1(n2220), .A2(n2205), .ZN(n2324) );
  OR2_X1 U3292 ( .A1(n3318), .A2(n3319), .ZN(n2325) );
  AND2_X1 U3293 ( .A1(n3316), .A2(n3315), .ZN(n3319) );
  AND2_X1 U3294 ( .A1(n3313), .A2(n3320), .ZN(n3318) );
  OR2_X1 U3295 ( .A1(n3315), .A2(n3316), .ZN(n3320) );
  OR2_X1 U3296 ( .A1(n2220), .A2(n2190), .ZN(n3316) );
  OR2_X1 U3297 ( .A1(n3321), .A2(n3322), .ZN(n3315) );
  AND2_X1 U3298 ( .A1(n3312), .A2(n3311), .ZN(n3322) );
  AND2_X1 U3299 ( .A1(n3309), .A2(n3323), .ZN(n3321) );
  OR2_X1 U3300 ( .A1(n3311), .A2(n3312), .ZN(n3323) );
  OR2_X1 U3301 ( .A1(n2220), .A2(n2209), .ZN(n3312) );
  OR2_X1 U3302 ( .A1(n3324), .A2(n3325), .ZN(n3311) );
  AND2_X1 U3303 ( .A1(n3308), .A2(n3307), .ZN(n3325) );
  AND2_X1 U3304 ( .A1(n3305), .A2(n3326), .ZN(n3324) );
  OR2_X1 U3305 ( .A1(n3307), .A2(n3308), .ZN(n3326) );
  OR2_X1 U3306 ( .A1(n2220), .A2(n2158), .ZN(n3308) );
  OR2_X1 U3307 ( .A1(n3327), .A2(n3328), .ZN(n3307) );
  AND2_X1 U3308 ( .A1(n3304), .A2(n3303), .ZN(n3328) );
  AND2_X1 U3309 ( .A1(n3301), .A2(n3329), .ZN(n3327) );
  OR2_X1 U3310 ( .A1(n3303), .A2(n3304), .ZN(n3329) );
  OR2_X1 U3311 ( .A1(n2220), .A2(n2214), .ZN(n3304) );
  OR2_X1 U3312 ( .A1(n3330), .A2(n3331), .ZN(n3303) );
  AND2_X1 U3313 ( .A1(n3300), .A2(n3299), .ZN(n3331) );
  AND2_X1 U3314 ( .A1(n3297), .A2(n3332), .ZN(n3330) );
  OR2_X1 U3315 ( .A1(n3299), .A2(n3300), .ZN(n3332) );
  OR2_X1 U3316 ( .A1(n2220), .A2(n2116), .ZN(n3300) );
  OR2_X1 U3317 ( .A1(n3333), .A2(n3334), .ZN(n3299) );
  AND2_X1 U3318 ( .A1(n2101), .A2(n3296), .ZN(n3334) );
  AND2_X1 U3319 ( .A1(n3294), .A2(n3335), .ZN(n3333) );
  OR2_X1 U3320 ( .A1(n3296), .A2(n2101), .ZN(n3335) );
  OR2_X1 U3321 ( .A1(n2220), .A2(n2219), .ZN(n2101) );
  OR2_X1 U3322 ( .A1(n3336), .A2(n3337), .ZN(n3296) );
  AND2_X1 U3323 ( .A1(n3290), .A2(n3293), .ZN(n3337) );
  AND2_X1 U3324 ( .A1(n3338), .A2(n3292), .ZN(n3336) );
  OR2_X1 U3325 ( .A1(n3339), .A2(n3340), .ZN(n3292) );
  AND2_X1 U3326 ( .A1(n3289), .A2(n3288), .ZN(n3340) );
  AND2_X1 U3327 ( .A1(n3286), .A2(n3341), .ZN(n3339) );
  OR2_X1 U3328 ( .A1(n3288), .A2(n3289), .ZN(n3341) );
  OR2_X1 U3329 ( .A1(n2220), .A2(n2224), .ZN(n3289) );
  OR2_X1 U3330 ( .A1(n3342), .A2(n3343), .ZN(n3288) );
  AND2_X1 U3331 ( .A1(n3282), .A2(n3285), .ZN(n3343) );
  AND2_X1 U3332 ( .A1(n3344), .A2(n3284), .ZN(n3342) );
  OR2_X1 U3333 ( .A1(n3345), .A2(n3346), .ZN(n3284) );
  AND2_X1 U3334 ( .A1(n3278), .A2(n3281), .ZN(n3346) );
  AND2_X1 U3335 ( .A1(n3347), .A2(n3280), .ZN(n3345) );
  OR2_X1 U3336 ( .A1(n3348), .A2(n3349), .ZN(n3280) );
  AND2_X1 U3337 ( .A1(n3274), .A2(n3277), .ZN(n3349) );
  AND2_X1 U3338 ( .A1(n3350), .A2(n3276), .ZN(n3348) );
  OR2_X1 U3339 ( .A1(n3351), .A2(n3352), .ZN(n3276) );
  AND2_X1 U3340 ( .A1(n3270), .A2(n3273), .ZN(n3352) );
  AND2_X1 U3341 ( .A1(n3353), .A2(n3272), .ZN(n3351) );
  OR2_X1 U3342 ( .A1(n3354), .A2(n3355), .ZN(n3272) );
  AND2_X1 U3343 ( .A1(n3266), .A2(n3269), .ZN(n3355) );
  AND2_X1 U3344 ( .A1(n3356), .A2(n3357), .ZN(n3354) );
  OR2_X1 U3345 ( .A1(n3269), .A2(n3266), .ZN(n3357) );
  OR2_X1 U3346 ( .A1(n1989), .A2(n2220), .ZN(n3266) );
  OR2_X1 U3347 ( .A1(n2115), .A2(n3358), .ZN(n3269) );
  OR2_X1 U3348 ( .A1(n2468), .A2(n2220), .ZN(n3358) );
  INV_X1 U3349 ( .A(n3268), .ZN(n3356) );
  OR2_X1 U3350 ( .A1(n3359), .A2(n3360), .ZN(n3268) );
  AND2_X1 U3351 ( .A1(b_5_), .A2(n3361), .ZN(n3360) );
  OR2_X1 U3352 ( .A1(n3362), .A2(n1965), .ZN(n3361) );
  AND2_X1 U3353 ( .A1(a_14_), .A2(n2215), .ZN(n3362) );
  AND2_X1 U3354 ( .A1(b_4_), .A2(n3363), .ZN(n3359) );
  OR2_X1 U3355 ( .A1(n3364), .A2(n1969), .ZN(n3363) );
  AND2_X1 U3356 ( .A1(a_15_), .A2(n2115), .ZN(n3364) );
  OR2_X1 U3357 ( .A1(n3273), .A2(n3270), .ZN(n3353) );
  XNOR2_X1 U3358 ( .A(n3365), .B(n3366), .ZN(n3270) );
  XOR2_X1 U3359 ( .A(n3367), .B(n3368), .Z(n3366) );
  OR2_X1 U3360 ( .A1(n2234), .A2(n2220), .ZN(n3273) );
  OR2_X1 U3361 ( .A1(n3277), .A2(n3274), .ZN(n3350) );
  XOR2_X1 U3362 ( .A(n3369), .B(n3370), .Z(n3274) );
  XOR2_X1 U3363 ( .A(n3371), .B(n3372), .Z(n3370) );
  OR2_X1 U3364 ( .A1(n2220), .A2(n2020), .ZN(n3277) );
  OR2_X1 U3365 ( .A1(n3281), .A2(n3278), .ZN(n3347) );
  XOR2_X1 U3366 ( .A(n3373), .B(n3374), .Z(n3278) );
  XOR2_X1 U3367 ( .A(n3375), .B(n3376), .Z(n3374) );
  OR2_X1 U3368 ( .A1(n2220), .A2(n2229), .ZN(n3281) );
  OR2_X1 U3369 ( .A1(n3285), .A2(n3282), .ZN(n3344) );
  XOR2_X1 U3370 ( .A(n3377), .B(n3378), .Z(n3282) );
  XOR2_X1 U3371 ( .A(n3379), .B(n3380), .Z(n3378) );
  OR2_X1 U3372 ( .A1(n2220), .A2(n2052), .ZN(n3285) );
  XOR2_X1 U3373 ( .A(n3381), .B(n3382), .Z(n3286) );
  XOR2_X1 U3374 ( .A(n3383), .B(n3384), .Z(n3382) );
  OR2_X1 U3375 ( .A1(n3293), .A2(n3290), .ZN(n3338) );
  XOR2_X1 U3376 ( .A(n3385), .B(n3386), .Z(n3290) );
  XOR2_X1 U3377 ( .A(n3387), .B(n3388), .Z(n3386) );
  OR2_X1 U3378 ( .A1(n2220), .A2(n2084), .ZN(n3293) );
  INV_X1 U3379 ( .A(b_6_), .ZN(n2220) );
  XOR2_X1 U3380 ( .A(n3389), .B(n3390), .Z(n3294) );
  XOR2_X1 U3381 ( .A(n3391), .B(n3392), .Z(n3390) );
  XOR2_X1 U3382 ( .A(n3393), .B(n3394), .Z(n3297) );
  XOR2_X1 U3383 ( .A(n3395), .B(n3396), .Z(n3394) );
  XOR2_X1 U3384 ( .A(n3397), .B(n3398), .Z(n3301) );
  XOR2_X1 U3385 ( .A(n3399), .B(n2120), .Z(n3398) );
  XOR2_X1 U3386 ( .A(n3400), .B(n3401), .Z(n3305) );
  XOR2_X1 U3387 ( .A(n3402), .B(n3403), .Z(n3401) );
  XOR2_X1 U3388 ( .A(n3404), .B(n3405), .Z(n3309) );
  XOR2_X1 U3389 ( .A(n3406), .B(n3407), .Z(n3405) );
  XOR2_X1 U3390 ( .A(n3408), .B(n3409), .Z(n3313) );
  XOR2_X1 U3391 ( .A(n3410), .B(n3411), .Z(n3409) );
  XOR2_X1 U3392 ( .A(n3412), .B(n3413), .Z(n2326) );
  XOR2_X1 U3393 ( .A(n3414), .B(n3415), .Z(n3413) );
  OR2_X1 U3394 ( .A1(n2314), .A2(n2315), .ZN(n2310) );
  OR2_X1 U3395 ( .A1(n3416), .A2(n3417), .ZN(n2315) );
  AND2_X1 U3396 ( .A1(n2331), .A2(n2330), .ZN(n3417) );
  AND2_X1 U3397 ( .A1(n2328), .A2(n3418), .ZN(n3416) );
  OR2_X1 U3398 ( .A1(n2330), .A2(n2331), .ZN(n3418) );
  OR2_X1 U3399 ( .A1(n2115), .A2(n2205), .ZN(n2331) );
  OR2_X1 U3400 ( .A1(n3419), .A2(n3420), .ZN(n2330) );
  AND2_X1 U3401 ( .A1(n3415), .A2(n3414), .ZN(n3420) );
  AND2_X1 U3402 ( .A1(n3412), .A2(n3421), .ZN(n3419) );
  OR2_X1 U3403 ( .A1(n3414), .A2(n3415), .ZN(n3421) );
  OR2_X1 U3404 ( .A1(n2115), .A2(n2190), .ZN(n3415) );
  OR2_X1 U3405 ( .A1(n3422), .A2(n3423), .ZN(n3414) );
  AND2_X1 U3406 ( .A1(n3411), .A2(n3410), .ZN(n3423) );
  AND2_X1 U3407 ( .A1(n3408), .A2(n3424), .ZN(n3422) );
  OR2_X1 U3408 ( .A1(n3410), .A2(n3411), .ZN(n3424) );
  OR2_X1 U3409 ( .A1(n2115), .A2(n2209), .ZN(n3411) );
  OR2_X1 U3410 ( .A1(n3425), .A2(n3426), .ZN(n3410) );
  AND2_X1 U3411 ( .A1(n3407), .A2(n3406), .ZN(n3426) );
  AND2_X1 U3412 ( .A1(n3404), .A2(n3427), .ZN(n3425) );
  OR2_X1 U3413 ( .A1(n3406), .A2(n3407), .ZN(n3427) );
  OR2_X1 U3414 ( .A1(n2115), .A2(n2158), .ZN(n3407) );
  OR2_X1 U3415 ( .A1(n3428), .A2(n3429), .ZN(n3406) );
  AND2_X1 U3416 ( .A1(n3403), .A2(n3402), .ZN(n3429) );
  AND2_X1 U3417 ( .A1(n3400), .A2(n3430), .ZN(n3428) );
  OR2_X1 U3418 ( .A1(n3402), .A2(n3403), .ZN(n3430) );
  OR2_X1 U3419 ( .A1(n2115), .A2(n2214), .ZN(n3403) );
  OR2_X1 U3420 ( .A1(n3431), .A2(n3432), .ZN(n3402) );
  AND2_X1 U3421 ( .A1(n2120), .A2(n3399), .ZN(n3432) );
  AND2_X1 U3422 ( .A1(n3397), .A2(n3433), .ZN(n3431) );
  OR2_X1 U3423 ( .A1(n3399), .A2(n2120), .ZN(n3433) );
  OR2_X1 U3424 ( .A1(n2115), .A2(n2116), .ZN(n2120) );
  OR2_X1 U3425 ( .A1(n3434), .A2(n3435), .ZN(n3399) );
  AND2_X1 U3426 ( .A1(n3396), .A2(n3395), .ZN(n3435) );
  AND2_X1 U3427 ( .A1(n3393), .A2(n3436), .ZN(n3434) );
  OR2_X1 U3428 ( .A1(n3395), .A2(n3396), .ZN(n3436) );
  OR2_X1 U3429 ( .A1(n2115), .A2(n2219), .ZN(n3396) );
  OR2_X1 U3430 ( .A1(n3437), .A2(n3438), .ZN(n3395) );
  AND2_X1 U3431 ( .A1(n3392), .A2(n3391), .ZN(n3438) );
  AND2_X1 U3432 ( .A1(n3389), .A2(n3439), .ZN(n3437) );
  OR2_X1 U3433 ( .A1(n3391), .A2(n3392), .ZN(n3439) );
  OR2_X1 U3434 ( .A1(n2115), .A2(n2084), .ZN(n3392) );
  OR2_X1 U3435 ( .A1(n3440), .A2(n3441), .ZN(n3391) );
  AND2_X1 U3436 ( .A1(n3385), .A2(n3388), .ZN(n3441) );
  AND2_X1 U3437 ( .A1(n3442), .A2(n3387), .ZN(n3440) );
  OR2_X1 U3438 ( .A1(n3443), .A2(n3444), .ZN(n3387) );
  AND2_X1 U3439 ( .A1(n3384), .A2(n3383), .ZN(n3444) );
  AND2_X1 U3440 ( .A1(n3381), .A2(n3445), .ZN(n3443) );
  OR2_X1 U3441 ( .A1(n3383), .A2(n3384), .ZN(n3445) );
  OR2_X1 U3442 ( .A1(n2115), .A2(n2052), .ZN(n3384) );
  OR2_X1 U3443 ( .A1(n3446), .A2(n3447), .ZN(n3383) );
  AND2_X1 U3444 ( .A1(n3377), .A2(n3380), .ZN(n3447) );
  AND2_X1 U3445 ( .A1(n3448), .A2(n3379), .ZN(n3446) );
  OR2_X1 U3446 ( .A1(n3449), .A2(n3450), .ZN(n3379) );
  AND2_X1 U3447 ( .A1(n3373), .A2(n3376), .ZN(n3450) );
  AND2_X1 U3448 ( .A1(n3451), .A2(n3375), .ZN(n3449) );
  OR2_X1 U3449 ( .A1(n3452), .A2(n3453), .ZN(n3375) );
  AND2_X1 U3450 ( .A1(n3369), .A2(n3372), .ZN(n3453) );
  AND2_X1 U3451 ( .A1(n3454), .A2(n3371), .ZN(n3452) );
  OR2_X1 U3452 ( .A1(n3455), .A2(n3456), .ZN(n3371) );
  AND2_X1 U3453 ( .A1(n3365), .A2(n3368), .ZN(n3456) );
  AND2_X1 U3454 ( .A1(n3457), .A2(n3458), .ZN(n3455) );
  OR2_X1 U3455 ( .A1(n3368), .A2(n3365), .ZN(n3458) );
  OR2_X1 U3456 ( .A1(n1989), .A2(n2115), .ZN(n3365) );
  OR2_X1 U3457 ( .A1(n2215), .A2(n3459), .ZN(n3368) );
  OR2_X1 U3458 ( .A1(n2468), .A2(n2115), .ZN(n3459) );
  INV_X1 U3459 ( .A(n3367), .ZN(n3457) );
  OR2_X1 U3460 ( .A1(n3460), .A2(n3461), .ZN(n3367) );
  AND2_X1 U3461 ( .A1(b_4_), .A2(n3462), .ZN(n3461) );
  OR2_X1 U3462 ( .A1(n3463), .A2(n1965), .ZN(n3462) );
  AND2_X1 U3463 ( .A1(a_14_), .A2(n2157), .ZN(n3463) );
  AND2_X1 U3464 ( .A1(b_3_), .A2(n3464), .ZN(n3460) );
  OR2_X1 U3465 ( .A1(n3465), .A2(n1969), .ZN(n3464) );
  AND2_X1 U3466 ( .A1(a_15_), .A2(n2215), .ZN(n3465) );
  OR2_X1 U3467 ( .A1(n3372), .A2(n3369), .ZN(n3454) );
  XNOR2_X1 U3468 ( .A(n3466), .B(n3467), .ZN(n3369) );
  XOR2_X1 U3469 ( .A(n3468), .B(n3469), .Z(n3467) );
  OR2_X1 U3470 ( .A1(n2234), .A2(n2115), .ZN(n3372) );
  OR2_X1 U3471 ( .A1(n3376), .A2(n3373), .ZN(n3451) );
  XOR2_X1 U3472 ( .A(n3470), .B(n3471), .Z(n3373) );
  XOR2_X1 U3473 ( .A(n3472), .B(n3473), .Z(n3471) );
  OR2_X1 U3474 ( .A1(n2020), .A2(n2115), .ZN(n3376) );
  OR2_X1 U3475 ( .A1(n3380), .A2(n3377), .ZN(n3448) );
  XOR2_X1 U3476 ( .A(n3474), .B(n3475), .Z(n3377) );
  XOR2_X1 U3477 ( .A(n3476), .B(n3477), .Z(n3475) );
  OR2_X1 U3478 ( .A1(n2115), .A2(n2229), .ZN(n3380) );
  XOR2_X1 U3479 ( .A(n3478), .B(n3479), .Z(n3381) );
  XOR2_X1 U3480 ( .A(n3480), .B(n3481), .Z(n3479) );
  OR2_X1 U3481 ( .A1(n3388), .A2(n3385), .ZN(n3442) );
  XOR2_X1 U3482 ( .A(n3482), .B(n3483), .Z(n3385) );
  XOR2_X1 U3483 ( .A(n3484), .B(n3485), .Z(n3483) );
  OR2_X1 U3484 ( .A1(n2115), .A2(n2224), .ZN(n3388) );
  INV_X1 U3485 ( .A(b_5_), .ZN(n2115) );
  XOR2_X1 U3486 ( .A(n3486), .B(n3487), .Z(n3389) );
  XOR2_X1 U3487 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR2_X1 U3488 ( .A(n3490), .B(n3491), .Z(n3393) );
  XOR2_X1 U3489 ( .A(n3492), .B(n3493), .Z(n3491) );
  XOR2_X1 U3490 ( .A(n3494), .B(n3495), .Z(n3397) );
  XOR2_X1 U3491 ( .A(n3496), .B(n3497), .Z(n3495) );
  XOR2_X1 U3492 ( .A(n3498), .B(n3499), .Z(n3400) );
  XOR2_X1 U3493 ( .A(n3500), .B(n3501), .Z(n3499) );
  XOR2_X1 U3494 ( .A(n3502), .B(n3503), .Z(n3404) );
  XOR2_X1 U3495 ( .A(n3504), .B(n2133), .Z(n3503) );
  XOR2_X1 U3496 ( .A(n3505), .B(n3506), .Z(n3408) );
  XOR2_X1 U3497 ( .A(n3507), .B(n3508), .Z(n3506) );
  XOR2_X1 U3498 ( .A(n3509), .B(n3510), .Z(n3412) );
  XOR2_X1 U3499 ( .A(n3511), .B(n3512), .Z(n3510) );
  XOR2_X1 U3500 ( .A(n3513), .B(n3514), .Z(n2328) );
  XOR2_X1 U3501 ( .A(n3515), .B(n3516), .Z(n3514) );
  XOR2_X1 U3502 ( .A(n2304), .B(n3517), .Z(n2314) );
  XOR2_X1 U3503 ( .A(n2303), .B(n2302), .Z(n3517) );
  OR2_X1 U3504 ( .A1(n2215), .A2(n2205), .ZN(n2302) );
  OR2_X1 U3505 ( .A1(n3518), .A2(n3519), .ZN(n2303) );
  AND2_X1 U3506 ( .A1(n3516), .A2(n3515), .ZN(n3519) );
  AND2_X1 U3507 ( .A1(n3513), .A2(n3520), .ZN(n3518) );
  OR2_X1 U3508 ( .A1(n3515), .A2(n3516), .ZN(n3520) );
  OR2_X1 U3509 ( .A1(n2215), .A2(n2190), .ZN(n3516) );
  OR2_X1 U3510 ( .A1(n3521), .A2(n3522), .ZN(n3515) );
  AND2_X1 U3511 ( .A1(n3512), .A2(n3511), .ZN(n3522) );
  AND2_X1 U3512 ( .A1(n3509), .A2(n3523), .ZN(n3521) );
  OR2_X1 U3513 ( .A1(n3511), .A2(n3512), .ZN(n3523) );
  OR2_X1 U3514 ( .A1(n2215), .A2(n2209), .ZN(n3512) );
  OR2_X1 U3515 ( .A1(n3524), .A2(n3525), .ZN(n3511) );
  AND2_X1 U3516 ( .A1(n3508), .A2(n3507), .ZN(n3525) );
  AND2_X1 U3517 ( .A1(n3505), .A2(n3526), .ZN(n3524) );
  OR2_X1 U3518 ( .A1(n3507), .A2(n3508), .ZN(n3526) );
  OR2_X1 U3519 ( .A1(n2215), .A2(n2158), .ZN(n3508) );
  OR2_X1 U3520 ( .A1(n3527), .A2(n3528), .ZN(n3507) );
  AND2_X1 U3521 ( .A1(n2133), .A2(n3504), .ZN(n3528) );
  AND2_X1 U3522 ( .A1(n3502), .A2(n3529), .ZN(n3527) );
  OR2_X1 U3523 ( .A1(n3504), .A2(n2133), .ZN(n3529) );
  OR2_X1 U3524 ( .A1(n2215), .A2(n2214), .ZN(n2133) );
  OR2_X1 U3525 ( .A1(n3530), .A2(n3531), .ZN(n3504) );
  AND2_X1 U3526 ( .A1(n3501), .A2(n3500), .ZN(n3531) );
  AND2_X1 U3527 ( .A1(n3498), .A2(n3532), .ZN(n3530) );
  OR2_X1 U3528 ( .A1(n3500), .A2(n3501), .ZN(n3532) );
  OR2_X1 U3529 ( .A1(n2215), .A2(n2116), .ZN(n3501) );
  OR2_X1 U3530 ( .A1(n3533), .A2(n3534), .ZN(n3500) );
  AND2_X1 U3531 ( .A1(n3497), .A2(n3496), .ZN(n3534) );
  AND2_X1 U3532 ( .A1(n3494), .A2(n3535), .ZN(n3533) );
  OR2_X1 U3533 ( .A1(n3496), .A2(n3497), .ZN(n3535) );
  OR2_X1 U3534 ( .A1(n2215), .A2(n2219), .ZN(n3497) );
  OR2_X1 U3535 ( .A1(n3536), .A2(n3537), .ZN(n3496) );
  AND2_X1 U3536 ( .A1(n3493), .A2(n3492), .ZN(n3537) );
  AND2_X1 U3537 ( .A1(n3490), .A2(n3538), .ZN(n3536) );
  OR2_X1 U3538 ( .A1(n3492), .A2(n3493), .ZN(n3538) );
  OR2_X1 U3539 ( .A1(n2215), .A2(n2084), .ZN(n3493) );
  OR2_X1 U3540 ( .A1(n3539), .A2(n3540), .ZN(n3492) );
  AND2_X1 U3541 ( .A1(n3489), .A2(n3488), .ZN(n3540) );
  AND2_X1 U3542 ( .A1(n3486), .A2(n3541), .ZN(n3539) );
  OR2_X1 U3543 ( .A1(n3488), .A2(n3489), .ZN(n3541) );
  OR2_X1 U3544 ( .A1(n2215), .A2(n2224), .ZN(n3489) );
  OR2_X1 U3545 ( .A1(n3542), .A2(n3543), .ZN(n3488) );
  AND2_X1 U3546 ( .A1(n3482), .A2(n3485), .ZN(n3543) );
  AND2_X1 U3547 ( .A1(n3544), .A2(n3484), .ZN(n3542) );
  OR2_X1 U3548 ( .A1(n3545), .A2(n3546), .ZN(n3484) );
  AND2_X1 U3549 ( .A1(n3481), .A2(n3480), .ZN(n3546) );
  AND2_X1 U3550 ( .A1(n3478), .A2(n3547), .ZN(n3545) );
  OR2_X1 U3551 ( .A1(n3480), .A2(n3481), .ZN(n3547) );
  OR2_X1 U3552 ( .A1(n2229), .A2(n2215), .ZN(n3481) );
  OR2_X1 U3553 ( .A1(n3548), .A2(n3549), .ZN(n3480) );
  AND2_X1 U3554 ( .A1(n3474), .A2(n3477), .ZN(n3549) );
  AND2_X1 U3555 ( .A1(n3550), .A2(n3476), .ZN(n3548) );
  OR2_X1 U3556 ( .A1(n3551), .A2(n3552), .ZN(n3476) );
  AND2_X1 U3557 ( .A1(n3470), .A2(n3473), .ZN(n3552) );
  AND2_X1 U3558 ( .A1(n3553), .A2(n3472), .ZN(n3551) );
  OR2_X1 U3559 ( .A1(n3554), .A2(n3555), .ZN(n3472) );
  AND2_X1 U3560 ( .A1(n3466), .A2(n3469), .ZN(n3555) );
  AND2_X1 U3561 ( .A1(n3556), .A2(n3557), .ZN(n3554) );
  OR2_X1 U3562 ( .A1(n3469), .A2(n3466), .ZN(n3557) );
  OR2_X1 U3563 ( .A1(n1989), .A2(n2215), .ZN(n3466) );
  OR2_X1 U3564 ( .A1(n2157), .A2(n3558), .ZN(n3469) );
  OR2_X1 U3565 ( .A1(n2468), .A2(n2215), .ZN(n3558) );
  INV_X1 U3566 ( .A(n3468), .ZN(n3556) );
  OR2_X1 U3567 ( .A1(n3559), .A2(n3560), .ZN(n3468) );
  AND2_X1 U3568 ( .A1(b_3_), .A2(n3561), .ZN(n3560) );
  OR2_X1 U3569 ( .A1(n3562), .A2(n1965), .ZN(n3561) );
  AND2_X1 U3570 ( .A1(a_14_), .A2(n2210), .ZN(n3562) );
  AND2_X1 U3571 ( .A1(b_2_), .A2(n3563), .ZN(n3559) );
  OR2_X1 U3572 ( .A1(n3564), .A2(n1969), .ZN(n3563) );
  AND2_X1 U3573 ( .A1(a_15_), .A2(n2157), .ZN(n3564) );
  OR2_X1 U3574 ( .A1(n3473), .A2(n3470), .ZN(n3553) );
  XNOR2_X1 U3575 ( .A(n3565), .B(n3566), .ZN(n3470) );
  XOR2_X1 U3576 ( .A(n3567), .B(n3568), .Z(n3566) );
  OR2_X1 U3577 ( .A1(n2234), .A2(n2215), .ZN(n3473) );
  OR2_X1 U3578 ( .A1(n3477), .A2(n3474), .ZN(n3550) );
  XOR2_X1 U3579 ( .A(n3569), .B(n3570), .Z(n3474) );
  XOR2_X1 U3580 ( .A(n3571), .B(n3572), .Z(n3570) );
  OR2_X1 U3581 ( .A1(n2020), .A2(n2215), .ZN(n3477) );
  XOR2_X1 U3582 ( .A(n3573), .B(n3574), .Z(n3478) );
  XOR2_X1 U3583 ( .A(n3575), .B(n3576), .Z(n3574) );
  OR2_X1 U3584 ( .A1(n3485), .A2(n3482), .ZN(n3544) );
  XOR2_X1 U3585 ( .A(n3577), .B(n3578), .Z(n3482) );
  XOR2_X1 U3586 ( .A(n3579), .B(n3580), .Z(n3578) );
  OR2_X1 U3587 ( .A1(n2215), .A2(n2052), .ZN(n3485) );
  INV_X1 U3588 ( .A(b_4_), .ZN(n2215) );
  XOR2_X1 U3589 ( .A(n3581), .B(n3582), .Z(n3486) );
  XOR2_X1 U3590 ( .A(n3583), .B(n3584), .Z(n3582) );
  XOR2_X1 U3591 ( .A(n3585), .B(n3586), .Z(n3490) );
  XOR2_X1 U3592 ( .A(n3587), .B(n3588), .Z(n3586) );
  XOR2_X1 U3593 ( .A(n3589), .B(n3590), .Z(n3494) );
  XOR2_X1 U3594 ( .A(n3591), .B(n3592), .Z(n3590) );
  XOR2_X1 U3595 ( .A(n3593), .B(n3594), .Z(n3498) );
  XOR2_X1 U3596 ( .A(n3595), .B(n3596), .Z(n3594) );
  XOR2_X1 U3597 ( .A(n3597), .B(n3598), .Z(n3502) );
  XOR2_X1 U3598 ( .A(n3599), .B(n3600), .Z(n3598) );
  XOR2_X1 U3599 ( .A(n3601), .B(n3602), .Z(n3505) );
  XOR2_X1 U3600 ( .A(n3603), .B(n3604), .Z(n3602) );
  XOR2_X1 U3601 ( .A(n3605), .B(n3606), .Z(n3509) );
  XOR2_X1 U3602 ( .A(n3607), .B(n2162), .Z(n3606) );
  XOR2_X1 U3603 ( .A(n3608), .B(n3609), .Z(n3513) );
  XOR2_X1 U3604 ( .A(n3610), .B(n3611), .Z(n3609) );
  XOR2_X1 U3605 ( .A(n3612), .B(n3613), .Z(n2304) );
  XOR2_X1 U3606 ( .A(n3614), .B(n3615), .Z(n3613) );
  OR2_X1 U3607 ( .A1(n2292), .A2(n2293), .ZN(n2288) );
  OR2_X1 U3608 ( .A1(n3616), .A2(n3617), .ZN(n2293) );
  AND2_X1 U3609 ( .A1(n2309), .A2(n2308), .ZN(n3617) );
  AND2_X1 U3610 ( .A1(n2306), .A2(n3618), .ZN(n3616) );
  OR2_X1 U3611 ( .A1(n2308), .A2(n2309), .ZN(n3618) );
  OR2_X1 U3612 ( .A1(n2157), .A2(n2205), .ZN(n2309) );
  OR2_X1 U3613 ( .A1(n3619), .A2(n3620), .ZN(n2308) );
  AND2_X1 U3614 ( .A1(n3615), .A2(n3614), .ZN(n3620) );
  AND2_X1 U3615 ( .A1(n3612), .A2(n3621), .ZN(n3619) );
  OR2_X1 U3616 ( .A1(n3614), .A2(n3615), .ZN(n3621) );
  OR2_X1 U3617 ( .A1(n2157), .A2(n2190), .ZN(n3615) );
  OR2_X1 U3618 ( .A1(n3622), .A2(n3623), .ZN(n3614) );
  AND2_X1 U3619 ( .A1(n3611), .A2(n3610), .ZN(n3623) );
  AND2_X1 U3620 ( .A1(n3608), .A2(n3624), .ZN(n3622) );
  OR2_X1 U3621 ( .A1(n3610), .A2(n3611), .ZN(n3624) );
  OR2_X1 U3622 ( .A1(n2157), .A2(n2209), .ZN(n3611) );
  OR2_X1 U3623 ( .A1(n3625), .A2(n3626), .ZN(n3610) );
  AND2_X1 U3624 ( .A1(n2162), .A2(n3607), .ZN(n3626) );
  AND2_X1 U3625 ( .A1(n3605), .A2(n3627), .ZN(n3625) );
  OR2_X1 U3626 ( .A1(n3607), .A2(n2162), .ZN(n3627) );
  OR2_X1 U3627 ( .A1(n2157), .A2(n2158), .ZN(n2162) );
  OR2_X1 U3628 ( .A1(n3628), .A2(n3629), .ZN(n3607) );
  AND2_X1 U3629 ( .A1(n3604), .A2(n3603), .ZN(n3629) );
  AND2_X1 U3630 ( .A1(n3601), .A2(n3630), .ZN(n3628) );
  OR2_X1 U3631 ( .A1(n3603), .A2(n3604), .ZN(n3630) );
  OR2_X1 U3632 ( .A1(n2157), .A2(n2214), .ZN(n3604) );
  OR2_X1 U3633 ( .A1(n3631), .A2(n3632), .ZN(n3603) );
  AND2_X1 U3634 ( .A1(n3600), .A2(n3599), .ZN(n3632) );
  AND2_X1 U3635 ( .A1(n3597), .A2(n3633), .ZN(n3631) );
  OR2_X1 U3636 ( .A1(n3599), .A2(n3600), .ZN(n3633) );
  OR2_X1 U3637 ( .A1(n2157), .A2(n2116), .ZN(n3600) );
  OR2_X1 U3638 ( .A1(n3634), .A2(n3635), .ZN(n3599) );
  AND2_X1 U3639 ( .A1(n3596), .A2(n3595), .ZN(n3635) );
  AND2_X1 U3640 ( .A1(n3593), .A2(n3636), .ZN(n3634) );
  OR2_X1 U3641 ( .A1(n3595), .A2(n3596), .ZN(n3636) );
  OR2_X1 U3642 ( .A1(n2157), .A2(n2219), .ZN(n3596) );
  OR2_X1 U3643 ( .A1(n3637), .A2(n3638), .ZN(n3595) );
  AND2_X1 U3644 ( .A1(n3592), .A2(n3591), .ZN(n3638) );
  AND2_X1 U3645 ( .A1(n3589), .A2(n3639), .ZN(n3637) );
  OR2_X1 U3646 ( .A1(n3591), .A2(n3592), .ZN(n3639) );
  OR2_X1 U3647 ( .A1(n2157), .A2(n2084), .ZN(n3592) );
  OR2_X1 U3648 ( .A1(n3640), .A2(n3641), .ZN(n3591) );
  AND2_X1 U3649 ( .A1(n3588), .A2(n3587), .ZN(n3641) );
  AND2_X1 U3650 ( .A1(n3585), .A2(n3642), .ZN(n3640) );
  OR2_X1 U3651 ( .A1(n3587), .A2(n3588), .ZN(n3642) );
  OR2_X1 U3652 ( .A1(n2157), .A2(n2224), .ZN(n3588) );
  OR2_X1 U3653 ( .A1(n3643), .A2(n3644), .ZN(n3587) );
  AND2_X1 U3654 ( .A1(n3584), .A2(n3583), .ZN(n3644) );
  AND2_X1 U3655 ( .A1(n3581), .A2(n3645), .ZN(n3643) );
  OR2_X1 U3656 ( .A1(n3583), .A2(n3584), .ZN(n3645) );
  OR2_X1 U3657 ( .A1(n2052), .A2(n2157), .ZN(n3584) );
  OR2_X1 U3658 ( .A1(n3646), .A2(n3647), .ZN(n3583) );
  AND2_X1 U3659 ( .A1(n3577), .A2(n3580), .ZN(n3647) );
  AND2_X1 U3660 ( .A1(n3648), .A2(n3579), .ZN(n3646) );
  OR2_X1 U3661 ( .A1(n3649), .A2(n3650), .ZN(n3579) );
  AND2_X1 U3662 ( .A1(n3576), .A2(n3575), .ZN(n3650) );
  AND2_X1 U3663 ( .A1(n3573), .A2(n3651), .ZN(n3649) );
  OR2_X1 U3664 ( .A1(n3575), .A2(n3576), .ZN(n3651) );
  OR2_X1 U3665 ( .A1(n2020), .A2(n2157), .ZN(n3576) );
  OR2_X1 U3666 ( .A1(n3652), .A2(n3653), .ZN(n3575) );
  AND2_X1 U3667 ( .A1(n3569), .A2(n3572), .ZN(n3653) );
  AND2_X1 U3668 ( .A1(n3654), .A2(n3571), .ZN(n3652) );
  OR2_X1 U3669 ( .A1(n3655), .A2(n3656), .ZN(n3571) );
  AND2_X1 U3670 ( .A1(n3565), .A2(n3568), .ZN(n3656) );
  AND2_X1 U3671 ( .A1(n3657), .A2(n3658), .ZN(n3655) );
  OR2_X1 U3672 ( .A1(n3568), .A2(n3565), .ZN(n3658) );
  OR2_X1 U3673 ( .A1(n1989), .A2(n2157), .ZN(n3565) );
  OR2_X1 U3674 ( .A1(n2210), .A2(n3659), .ZN(n3568) );
  OR2_X1 U3675 ( .A1(n2468), .A2(n2157), .ZN(n3659) );
  INV_X1 U3676 ( .A(n3567), .ZN(n3657) );
  OR2_X1 U3677 ( .A1(n3660), .A2(n3661), .ZN(n3567) );
  AND2_X1 U3678 ( .A1(b_2_), .A2(n3662), .ZN(n3661) );
  OR2_X1 U3679 ( .A1(n3663), .A2(n1965), .ZN(n3662) );
  AND2_X1 U3680 ( .A1(a_14_), .A2(n2189), .ZN(n3663) );
  AND2_X1 U3681 ( .A1(b_1_), .A2(n3664), .ZN(n3660) );
  OR2_X1 U3682 ( .A1(n3665), .A2(n1969), .ZN(n3664) );
  AND2_X1 U3683 ( .A1(a_15_), .A2(n2210), .ZN(n3665) );
  OR2_X1 U3684 ( .A1(n3572), .A2(n3569), .ZN(n3654) );
  XNOR2_X1 U3685 ( .A(n3666), .B(n3667), .ZN(n3569) );
  XOR2_X1 U3686 ( .A(n3668), .B(n3669), .Z(n3667) );
  OR2_X1 U3687 ( .A1(n2234), .A2(n2157), .ZN(n3572) );
  XOR2_X1 U3688 ( .A(n3670), .B(n3671), .Z(n3573) );
  XOR2_X1 U3689 ( .A(n3672), .B(n3673), .Z(n3671) );
  OR2_X1 U3690 ( .A1(n3580), .A2(n3577), .ZN(n3648) );
  XOR2_X1 U3691 ( .A(n3674), .B(n3675), .Z(n3577) );
  XOR2_X1 U3692 ( .A(n3676), .B(n3677), .Z(n3675) );
  OR2_X1 U3693 ( .A1(n2229), .A2(n2157), .ZN(n3580) );
  INV_X1 U3694 ( .A(b_3_), .ZN(n2157) );
  XOR2_X1 U3695 ( .A(n3678), .B(n3679), .Z(n3581) );
  XOR2_X1 U3696 ( .A(n3680), .B(n3681), .Z(n3679) );
  XOR2_X1 U3697 ( .A(n3682), .B(n3683), .Z(n3585) );
  XOR2_X1 U3698 ( .A(n3684), .B(n3685), .Z(n3683) );
  XOR2_X1 U3699 ( .A(n3686), .B(n3687), .Z(n3589) );
  XOR2_X1 U3700 ( .A(n3688), .B(n3689), .Z(n3687) );
  XOR2_X1 U3701 ( .A(n3690), .B(n3691), .Z(n3593) );
  XOR2_X1 U3702 ( .A(n3692), .B(n3693), .Z(n3691) );
  XOR2_X1 U3703 ( .A(n3694), .B(n3695), .Z(n3597) );
  XOR2_X1 U3704 ( .A(n3696), .B(n3697), .Z(n3695) );
  XOR2_X1 U3705 ( .A(n3698), .B(n3699), .Z(n3601) );
  XOR2_X1 U3706 ( .A(n3700), .B(n3701), .Z(n3699) );
  XOR2_X1 U3707 ( .A(n3702), .B(n3703), .Z(n3605) );
  XOR2_X1 U3708 ( .A(n3704), .B(n3705), .Z(n3703) );
  XOR2_X1 U3709 ( .A(n3706), .B(n3707), .Z(n3608) );
  XOR2_X1 U3710 ( .A(n3708), .B(n3709), .Z(n3707) );
  XOR2_X1 U3711 ( .A(n3710), .B(n3711), .Z(n3612) );
  XOR2_X1 U3712 ( .A(n3712), .B(n2175), .Z(n3711) );
  XOR2_X1 U3713 ( .A(n3713), .B(n3714), .Z(n2306) );
  XOR2_X1 U3714 ( .A(n3715), .B(n3716), .Z(n3714) );
  XOR2_X1 U3715 ( .A(n3717), .B(n3718), .Z(n2292) );
  XOR2_X1 U3716 ( .A(n3719), .B(n3720), .Z(n3718) );
  OR2_X1 U3717 ( .A1(n2143), .A2(n3721), .ZN(n2139) );
  OR2_X1 U3718 ( .A1(n2142), .A2(n2140), .ZN(n3721) );
  XNOR2_X1 U3719 ( .A(n3722), .B(n3723), .ZN(n2140) );
  OR2_X1 U3720 ( .A1(n3724), .A2(n2205), .ZN(n3722) );
  XOR2_X1 U3721 ( .A(n3725), .B(n3726), .Z(n2142) );
  XOR2_X1 U3722 ( .A(n3727), .B(n3728), .Z(n3726) );
  OR2_X1 U3723 ( .A1(n3729), .A2(n3730), .ZN(n2143) );
  AND2_X1 U3724 ( .A1(n3720), .A2(n3719), .ZN(n3730) );
  AND2_X1 U3725 ( .A1(n3717), .A2(n3731), .ZN(n3729) );
  OR2_X1 U3726 ( .A1(n3719), .A2(n3720), .ZN(n3731) );
  OR2_X1 U3727 ( .A1(n2210), .A2(n2205), .ZN(n3720) );
  OR2_X1 U3728 ( .A1(n3732), .A2(n3733), .ZN(n3719) );
  AND2_X1 U3729 ( .A1(n3716), .A2(n3715), .ZN(n3733) );
  AND2_X1 U3730 ( .A1(n3713), .A2(n3734), .ZN(n3732) );
  OR2_X1 U3731 ( .A1(n3715), .A2(n3716), .ZN(n3734) );
  OR2_X1 U3732 ( .A1(n2210), .A2(n2190), .ZN(n3716) );
  OR2_X1 U3733 ( .A1(n3735), .A2(n3736), .ZN(n3715) );
  AND2_X1 U3734 ( .A1(n2175), .A2(n3712), .ZN(n3736) );
  AND2_X1 U3735 ( .A1(n3710), .A2(n3737), .ZN(n3735) );
  OR2_X1 U3736 ( .A1(n3712), .A2(n2175), .ZN(n3737) );
  OR2_X1 U3737 ( .A1(n2210), .A2(n2209), .ZN(n2175) );
  OR2_X1 U3738 ( .A1(n3738), .A2(n3739), .ZN(n3712) );
  AND2_X1 U3739 ( .A1(n3709), .A2(n3708), .ZN(n3739) );
  AND2_X1 U3740 ( .A1(n3706), .A2(n3740), .ZN(n3738) );
  OR2_X1 U3741 ( .A1(n3708), .A2(n3709), .ZN(n3740) );
  OR2_X1 U3742 ( .A1(n2210), .A2(n2158), .ZN(n3709) );
  OR2_X1 U3743 ( .A1(n3741), .A2(n3742), .ZN(n3708) );
  AND2_X1 U3744 ( .A1(n3705), .A2(n3704), .ZN(n3742) );
  AND2_X1 U3745 ( .A1(n3702), .A2(n3743), .ZN(n3741) );
  OR2_X1 U3746 ( .A1(n3704), .A2(n3705), .ZN(n3743) );
  OR2_X1 U3747 ( .A1(n2210), .A2(n2214), .ZN(n3705) );
  OR2_X1 U3748 ( .A1(n3744), .A2(n3745), .ZN(n3704) );
  AND2_X1 U3749 ( .A1(n3701), .A2(n3700), .ZN(n3745) );
  AND2_X1 U3750 ( .A1(n3698), .A2(n3746), .ZN(n3744) );
  OR2_X1 U3751 ( .A1(n3700), .A2(n3701), .ZN(n3746) );
  OR2_X1 U3752 ( .A1(n2210), .A2(n2116), .ZN(n3701) );
  OR2_X1 U3753 ( .A1(n3747), .A2(n3748), .ZN(n3700) );
  AND2_X1 U3754 ( .A1(n3697), .A2(n3696), .ZN(n3748) );
  AND2_X1 U3755 ( .A1(n3694), .A2(n3749), .ZN(n3747) );
  OR2_X1 U3756 ( .A1(n3696), .A2(n3697), .ZN(n3749) );
  OR2_X1 U3757 ( .A1(n2210), .A2(n2219), .ZN(n3697) );
  OR2_X1 U3758 ( .A1(n3750), .A2(n3751), .ZN(n3696) );
  AND2_X1 U3759 ( .A1(n3693), .A2(n3692), .ZN(n3751) );
  AND2_X1 U3760 ( .A1(n3690), .A2(n3752), .ZN(n3750) );
  OR2_X1 U3761 ( .A1(n3692), .A2(n3693), .ZN(n3752) );
  OR2_X1 U3762 ( .A1(n2210), .A2(n2084), .ZN(n3693) );
  OR2_X1 U3763 ( .A1(n3753), .A2(n3754), .ZN(n3692) );
  AND2_X1 U3764 ( .A1(n3689), .A2(n3688), .ZN(n3754) );
  AND2_X1 U3765 ( .A1(n3686), .A2(n3755), .ZN(n3753) );
  OR2_X1 U3766 ( .A1(n3688), .A2(n3689), .ZN(n3755) );
  OR2_X1 U3767 ( .A1(n2224), .A2(n2210), .ZN(n3689) );
  OR2_X1 U3768 ( .A1(n3756), .A2(n3757), .ZN(n3688) );
  AND2_X1 U3769 ( .A1(n3685), .A2(n3684), .ZN(n3757) );
  AND2_X1 U3770 ( .A1(n3682), .A2(n3758), .ZN(n3756) );
  OR2_X1 U3771 ( .A1(n3684), .A2(n3685), .ZN(n3758) );
  OR2_X1 U3772 ( .A1(n2052), .A2(n2210), .ZN(n3685) );
  OR2_X1 U3773 ( .A1(n3759), .A2(n3760), .ZN(n3684) );
  AND2_X1 U3774 ( .A1(n3681), .A2(n3680), .ZN(n3760) );
  AND2_X1 U3775 ( .A1(n3678), .A2(n3761), .ZN(n3759) );
  OR2_X1 U3776 ( .A1(n3680), .A2(n3681), .ZN(n3761) );
  OR2_X1 U3777 ( .A1(n2229), .A2(n2210), .ZN(n3681) );
  OR2_X1 U3778 ( .A1(n3762), .A2(n3763), .ZN(n3680) );
  AND2_X1 U3779 ( .A1(n3674), .A2(n3677), .ZN(n3763) );
  AND2_X1 U3780 ( .A1(n3764), .A2(n3676), .ZN(n3762) );
  OR2_X1 U3781 ( .A1(n3765), .A2(n3766), .ZN(n3676) );
  AND2_X1 U3782 ( .A1(n3673), .A2(n3672), .ZN(n3766) );
  AND2_X1 U3783 ( .A1(n3670), .A2(n3767), .ZN(n3765) );
  OR2_X1 U3784 ( .A1(n3672), .A2(n3673), .ZN(n3767) );
  OR2_X1 U3785 ( .A1(n2234), .A2(n2210), .ZN(n3673) );
  OR2_X1 U3786 ( .A1(n3768), .A2(n3769), .ZN(n3672) );
  AND2_X1 U3787 ( .A1(n3666), .A2(n3669), .ZN(n3769) );
  AND2_X1 U3788 ( .A1(n3770), .A2(n3771), .ZN(n3768) );
  OR2_X1 U3789 ( .A1(n3669), .A2(n3666), .ZN(n3771) );
  OR2_X1 U3790 ( .A1(n1989), .A2(n2210), .ZN(n3666) );
  OR2_X1 U3791 ( .A1(n2189), .A2(n3772), .ZN(n3669) );
  OR2_X1 U3792 ( .A1(n2468), .A2(n2210), .ZN(n3772) );
  INV_X1 U3793 ( .A(n3668), .ZN(n3770) );
  OR2_X1 U3794 ( .A1(n3773), .A2(n3774), .ZN(n3668) );
  AND2_X1 U3795 ( .A1(b_1_), .A2(n3775), .ZN(n3774) );
  OR2_X1 U3796 ( .A1(n3776), .A2(n1965), .ZN(n3775) );
  AND2_X1 U3797 ( .A1(n3777), .A2(a_14_), .ZN(n1965) );
  AND2_X1 U3798 ( .A1(a_14_), .A2(n3724), .ZN(n3776) );
  AND2_X1 U3799 ( .A1(b_0_), .A2(n3778), .ZN(n3773) );
  OR2_X1 U3800 ( .A1(n3779), .A2(n1969), .ZN(n3778) );
  AND2_X1 U3801 ( .A1(n3780), .A2(a_15_), .ZN(n1969) );
  AND2_X1 U3802 ( .A1(a_15_), .A2(n2189), .ZN(n3779) );
  XNOR2_X1 U3803 ( .A(n3781), .B(n3782), .ZN(n3670) );
  OR2_X1 U3804 ( .A1(n3783), .A2(n3784), .ZN(n3781) );
  INV_X1 U3805 ( .A(n3785), .ZN(n3784) );
  AND2_X1 U3806 ( .A1(n3786), .A2(n3787), .ZN(n3783) );
  OR2_X1 U3807 ( .A1(n3677), .A2(n3674), .ZN(n3764) );
  XOR2_X1 U3808 ( .A(n3788), .B(n3789), .Z(n3674) );
  XOR2_X1 U3809 ( .A(n3790), .B(n3791), .Z(n3788) );
  OR2_X1 U3810 ( .A1(n2020), .A2(n2210), .ZN(n3677) );
  INV_X1 U3811 ( .A(b_2_), .ZN(n2210) );
  XNOR2_X1 U3812 ( .A(n3792), .B(n3793), .ZN(n3678) );
  XNOR2_X1 U3813 ( .A(n3794), .B(n3795), .ZN(n3792) );
  XNOR2_X1 U3814 ( .A(n3796), .B(n3797), .ZN(n3682) );
  XNOR2_X1 U3815 ( .A(n3798), .B(n3799), .ZN(n3796) );
  XNOR2_X1 U3816 ( .A(n3800), .B(n3801), .ZN(n3686) );
  XNOR2_X1 U3817 ( .A(n3802), .B(n3803), .ZN(n3800) );
  XOR2_X1 U3818 ( .A(n3804), .B(n3805), .Z(n3690) );
  XOR2_X1 U3819 ( .A(n3806), .B(n3807), .Z(n3805) );
  XOR2_X1 U3820 ( .A(n3808), .B(n3809), .Z(n3694) );
  XOR2_X1 U3821 ( .A(n3810), .B(n3811), .Z(n3809) );
  XOR2_X1 U3822 ( .A(n3812), .B(n3813), .Z(n3698) );
  XOR2_X1 U3823 ( .A(n3814), .B(n3815), .Z(n3813) );
  XOR2_X1 U3824 ( .A(n3816), .B(n3817), .Z(n3702) );
  XOR2_X1 U3825 ( .A(n3818), .B(n3819), .Z(n3817) );
  XOR2_X1 U3826 ( .A(n3820), .B(n3821), .Z(n3706) );
  XOR2_X1 U3827 ( .A(n3822), .B(n3823), .Z(n3821) );
  XOR2_X1 U3828 ( .A(n3824), .B(n3825), .Z(n3710) );
  XOR2_X1 U3829 ( .A(n3826), .B(n3827), .Z(n3825) );
  XOR2_X1 U3830 ( .A(n3828), .B(n3829), .Z(n3713) );
  XOR2_X1 U3831 ( .A(n3830), .B(n3831), .Z(n3829) );
  XOR2_X1 U3832 ( .A(n3832), .B(n3833), .Z(n3717) );
  XOR2_X1 U3833 ( .A(n3834), .B(n2194), .Z(n3833) );
  OR2_X1 U3834 ( .A1(n3723), .A2(n2205), .ZN(n2285) );
  OR2_X1 U3835 ( .A1(n3835), .A2(n3836), .ZN(n3723) );
  AND2_X1 U3836 ( .A1(n3725), .A2(n3727), .ZN(n3836) );
  AND2_X1 U3837 ( .A1(n3837), .A2(n3728), .ZN(n3835) );
  OR2_X1 U3838 ( .A1(n2189), .A2(n2205), .ZN(n3728) );
  INV_X1 U3839 ( .A(a_0_), .ZN(n2205) );
  OR2_X1 U3840 ( .A1(n3727), .A2(n3725), .ZN(n3837) );
  OR2_X1 U3841 ( .A1(n3724), .A2(n2190), .ZN(n3725) );
  OR2_X1 U3842 ( .A1(n3838), .A2(n3839), .ZN(n3727) );
  AND2_X1 U3843 ( .A1(n3832), .A2(n3834), .ZN(n3839) );
  AND2_X1 U3844 ( .A1(n3840), .A2(n2194), .ZN(n3838) );
  OR2_X1 U3845 ( .A1(n2189), .A2(n2190), .ZN(n2194) );
  INV_X1 U3846 ( .A(a_1_), .ZN(n2190) );
  OR2_X1 U3847 ( .A1(n3834), .A2(n3832), .ZN(n3840) );
  OR2_X1 U3848 ( .A1(n3724), .A2(n2209), .ZN(n3832) );
  OR2_X1 U3849 ( .A1(n3841), .A2(n3842), .ZN(n3834) );
  AND2_X1 U3850 ( .A1(n3828), .A2(n3830), .ZN(n3842) );
  AND2_X1 U3851 ( .A1(n3843), .A2(n3831), .ZN(n3841) );
  OR2_X1 U3852 ( .A1(n3724), .A2(n2158), .ZN(n3831) );
  OR2_X1 U3853 ( .A1(n3830), .A2(n3828), .ZN(n3843) );
  OR2_X1 U3854 ( .A1(n2189), .A2(n2209), .ZN(n3828) );
  INV_X1 U3855 ( .A(a_2_), .ZN(n2209) );
  OR2_X1 U3856 ( .A1(n3844), .A2(n3845), .ZN(n3830) );
  AND2_X1 U3857 ( .A1(n3824), .A2(n3826), .ZN(n3845) );
  AND2_X1 U3858 ( .A1(n3846), .A2(n3827), .ZN(n3844) );
  OR2_X1 U3859 ( .A1(n3724), .A2(n2214), .ZN(n3827) );
  OR2_X1 U3860 ( .A1(n3826), .A2(n3824), .ZN(n3846) );
  OR2_X1 U3861 ( .A1(n2189), .A2(n2158), .ZN(n3824) );
  INV_X1 U3862 ( .A(a_3_), .ZN(n2158) );
  OR2_X1 U3863 ( .A1(n3847), .A2(n3848), .ZN(n3826) );
  AND2_X1 U3864 ( .A1(n3820), .A2(n3822), .ZN(n3848) );
  AND2_X1 U3865 ( .A1(n3849), .A2(n3823), .ZN(n3847) );
  OR2_X1 U3866 ( .A1(n3724), .A2(n2116), .ZN(n3823) );
  OR2_X1 U3867 ( .A1(n3822), .A2(n3820), .ZN(n3849) );
  OR2_X1 U3868 ( .A1(n2189), .A2(n2214), .ZN(n3820) );
  INV_X1 U3869 ( .A(a_4_), .ZN(n2214) );
  OR2_X1 U3870 ( .A1(n3850), .A2(n3851), .ZN(n3822) );
  AND2_X1 U3871 ( .A1(n3816), .A2(n3818), .ZN(n3851) );
  AND2_X1 U3872 ( .A1(n3852), .A2(n3819), .ZN(n3850) );
  OR2_X1 U3873 ( .A1(n2219), .A2(n3724), .ZN(n3819) );
  OR2_X1 U3874 ( .A1(n3818), .A2(n3816), .ZN(n3852) );
  OR2_X1 U3875 ( .A1(n2189), .A2(n2116), .ZN(n3816) );
  INV_X1 U3876 ( .A(a_5_), .ZN(n2116) );
  OR2_X1 U3877 ( .A1(n3853), .A2(n3854), .ZN(n3818) );
  AND2_X1 U3878 ( .A1(n3812), .A2(n3814), .ZN(n3854) );
  AND2_X1 U3879 ( .A1(n3855), .A2(n3815), .ZN(n3853) );
  OR2_X1 U3880 ( .A1(n2084), .A2(n3724), .ZN(n3815) );
  OR2_X1 U3881 ( .A1(n3814), .A2(n3812), .ZN(n3855) );
  OR2_X1 U3882 ( .A1(n2189), .A2(n2219), .ZN(n3812) );
  INV_X1 U3883 ( .A(a_6_), .ZN(n2219) );
  OR2_X1 U3884 ( .A1(n3856), .A2(n3857), .ZN(n3814) );
  AND2_X1 U3885 ( .A1(n3808), .A2(n3810), .ZN(n3857) );
  AND2_X1 U3886 ( .A1(n3858), .A2(n3811), .ZN(n3856) );
  OR2_X1 U3887 ( .A1(n2224), .A2(n3724), .ZN(n3811) );
  OR2_X1 U3888 ( .A1(n3810), .A2(n3808), .ZN(n3858) );
  OR2_X1 U3889 ( .A1(n2084), .A2(n2189), .ZN(n3808) );
  INV_X1 U3890 ( .A(a_7_), .ZN(n2084) );
  OR2_X1 U3891 ( .A1(n3859), .A2(n3860), .ZN(n3810) );
  AND2_X1 U3892 ( .A1(n3804), .A2(n3806), .ZN(n3860) );
  AND2_X1 U3893 ( .A1(n3861), .A2(n3807), .ZN(n3859) );
  OR2_X1 U3894 ( .A1(n2052), .A2(n3724), .ZN(n3807) );
  OR2_X1 U3895 ( .A1(n3806), .A2(n3804), .ZN(n3861) );
  OR2_X1 U3896 ( .A1(n2224), .A2(n2189), .ZN(n3804) );
  INV_X1 U3897 ( .A(a_8_), .ZN(n2224) );
  OR2_X1 U3898 ( .A1(n3862), .A2(n3863), .ZN(n3806) );
  AND2_X1 U3899 ( .A1(n3801), .A2(n3803), .ZN(n3863) );
  AND2_X1 U3900 ( .A1(n3864), .A2(n3802), .ZN(n3862) );
  OR2_X1 U3901 ( .A1(n2229), .A2(n3724), .ZN(n3802) );
  OR2_X1 U3902 ( .A1(n3803), .A2(n3801), .ZN(n3864) );
  OR2_X1 U3903 ( .A1(n2052), .A2(n2189), .ZN(n3801) );
  INV_X1 U3904 ( .A(a_9_), .ZN(n2052) );
  OR2_X1 U3905 ( .A1(n3865), .A2(n3866), .ZN(n3803) );
  AND2_X1 U3906 ( .A1(n3797), .A2(n3799), .ZN(n3866) );
  AND2_X1 U3907 ( .A1(n3867), .A2(n3798), .ZN(n3865) );
  OR2_X1 U3908 ( .A1(n2020), .A2(n3724), .ZN(n3798) );
  OR2_X1 U3909 ( .A1(n3799), .A2(n3797), .ZN(n3867) );
  OR2_X1 U3910 ( .A1(n2229), .A2(n2189), .ZN(n3797) );
  INV_X1 U3911 ( .A(a_10_), .ZN(n2229) );
  OR2_X1 U3912 ( .A1(n3868), .A2(n3869), .ZN(n3799) );
  AND2_X1 U3913 ( .A1(n3793), .A2(n3795), .ZN(n3869) );
  AND2_X1 U3914 ( .A1(n3870), .A2(n3794), .ZN(n3868) );
  OR2_X1 U3915 ( .A1(n2234), .A2(n3724), .ZN(n3794) );
  OR2_X1 U3916 ( .A1(n3795), .A2(n3793), .ZN(n3870) );
  OR2_X1 U3917 ( .A1(n2020), .A2(n2189), .ZN(n3793) );
  INV_X1 U3918 ( .A(a_11_), .ZN(n2020) );
  OR2_X1 U3919 ( .A1(n3871), .A2(n3872), .ZN(n3795) );
  AND2_X1 U3920 ( .A1(n3789), .A2(n3791), .ZN(n3872) );
  AND2_X1 U3921 ( .A1(n3790), .A2(n3873), .ZN(n3871) );
  OR2_X1 U3922 ( .A1(n3791), .A2(n3789), .ZN(n3873) );
  OR2_X1 U3923 ( .A1(n2234), .A2(n2189), .ZN(n3789) );
  INV_X1 U3924 ( .A(a_12_), .ZN(n2234) );
  OR2_X1 U3925 ( .A1(n1989), .A2(n3724), .ZN(n3791) );
  AND2_X1 U3926 ( .A1(n3785), .A2(n3782), .ZN(n3790) );
  OR2_X1 U3927 ( .A1(n3724), .A2(n3874), .ZN(n3782) );
  OR2_X1 U3928 ( .A1(n2468), .A2(n2189), .ZN(n3874) );
  OR2_X1 U3929 ( .A1(n3777), .A2(n3780), .ZN(n2468) );
  INV_X1 U3930 ( .A(a_15_), .ZN(n3777) );
  OR2_X1 U3931 ( .A1(n3787), .A2(n3786), .ZN(n3785) );
  OR2_X1 U3932 ( .A1(n3780), .A2(n3724), .ZN(n3786) );
  INV_X1 U3933 ( .A(b_0_), .ZN(n3724) );
  INV_X1 U3934 ( .A(a_14_), .ZN(n3780) );
  OR2_X1 U3935 ( .A1(n1989), .A2(n2189), .ZN(n3787) );
  INV_X1 U3936 ( .A(b_1_), .ZN(n2189) );
  INV_X1 U3937 ( .A(a_13_), .ZN(n1989) );
  INV_X1 U3938 ( .A(operation), .ZN(n1955) );
endmodule

