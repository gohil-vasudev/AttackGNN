module add_mul_combine_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_mul_0_, Result_mul_1_, Result_mul_2_, 
        Result_mul_3_, Result_mul_4_, Result_mul_5_, Result_mul_6_, 
        Result_mul_7_, Result_mul_8_, Result_mul_9_, Result_mul_10_, 
        Result_mul_11_, Result_mul_12_, Result_mul_13_, Result_mul_14_, 
        Result_mul_15_, Result_mul_16_, Result_mul_17_, Result_mul_18_, 
        Result_mul_19_, Result_mul_20_, Result_mul_21_, Result_mul_22_, 
        Result_mul_23_, Result_mul_24_, Result_mul_25_, Result_mul_26_, 
        Result_mul_27_, Result_mul_28_, Result_mul_29_, Result_mul_30_, 
        Result_mul_31_, Result_add_0_, Result_add_1_, Result_add_2_, 
        Result_add_3_, Result_add_4_, Result_add_5_, Result_add_6_, 
        Result_add_7_, Result_add_8_, Result_add_9_, Result_add_10_, 
        Result_add_11_, Result_add_12_, Result_add_13_, Result_add_14_, 
        Result_add_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_;
  wire   n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080;

  XOR2_X1 U2081 ( .A(n2034), .B(n2035), .Z(Result_mul_9_) );
  NAND2_X1 U2082 ( .A1(n2036), .A2(n2037), .ZN(n2035) );
  NAND2_X1 U2083 ( .A1(n2038), .A2(n2039), .ZN(n2034) );
  NAND2_X1 U2084 ( .A1(n2040), .A2(n2041), .ZN(n2039) );
  NAND2_X1 U2085 ( .A1(n2042), .A2(n2043), .ZN(n2040) );
  XOR2_X1 U2086 ( .A(n2044), .B(n2045), .Z(Result_mul_8_) );
  XOR2_X1 U2087 ( .A(n2046), .B(n2047), .Z(Result_mul_7_) );
  NAND2_X1 U2088 ( .A1(n2045), .A2(n2044), .ZN(n2047) );
  NAND2_X1 U2089 ( .A1(n2048), .A2(n2049), .ZN(n2046) );
  NAND2_X1 U2090 ( .A1(n2050), .A2(n2051), .ZN(n2049) );
  NAND2_X1 U2091 ( .A1(n2052), .A2(n2053), .ZN(n2050) );
  XOR2_X1 U2092 ( .A(n2054), .B(n2055), .Z(Result_mul_6_) );
  XOR2_X1 U2093 ( .A(n2056), .B(n2057), .Z(Result_mul_5_) );
  NAND2_X1 U2094 ( .A1(n2055), .A2(n2054), .ZN(n2057) );
  NAND2_X1 U2095 ( .A1(n2058), .A2(n2059), .ZN(n2056) );
  NAND2_X1 U2096 ( .A1(n2060), .A2(n2061), .ZN(n2059) );
  NAND2_X1 U2097 ( .A1(n2062), .A2(n2063), .ZN(n2060) );
  XOR2_X1 U2098 ( .A(n2064), .B(n2065), .Z(Result_mul_4_) );
  XOR2_X1 U2099 ( .A(n2066), .B(n2067), .Z(Result_mul_3_) );
  NAND2_X1 U2100 ( .A1(n2065), .A2(n2064), .ZN(n2067) );
  NAND2_X1 U2101 ( .A1(n2068), .A2(n2069), .ZN(n2066) );
  NAND2_X1 U2102 ( .A1(n2070), .A2(n2071), .ZN(n2069) );
  NAND2_X1 U2103 ( .A1(n2072), .A2(n2073), .ZN(n2070) );
  NAND2_X1 U2104 ( .A1(n2074), .A2(n2075), .ZN(Result_mul_30_) );
  NAND2_X1 U2105 ( .A1(b_14_), .A2(n2076), .ZN(n2075) );
  NAND2_X1 U2106 ( .A1(n2077), .A2(n2078), .ZN(n2076) );
  NAND2_X1 U2107 ( .A1(a_15_), .A2(n2079), .ZN(n2078) );
  NAND2_X1 U2108 ( .A1(b_15_), .A2(n2080), .ZN(n2074) );
  NAND2_X1 U2109 ( .A1(n2081), .A2(n2082), .ZN(n2080) );
  NAND2_X1 U2110 ( .A1(a_14_), .A2(n2083), .ZN(n2082) );
  XOR2_X1 U2111 ( .A(n2084), .B(n2085), .Z(Result_mul_2_) );
  XOR2_X1 U2112 ( .A(n2086), .B(n2087), .Z(Result_mul_29_) );
  XOR2_X1 U2113 ( .A(n2088), .B(n2089), .Z(n2087) );
  XOR2_X1 U2114 ( .A(n2090), .B(n2091), .Z(Result_mul_28_) );
  XOR2_X1 U2115 ( .A(n2092), .B(n2093), .Z(n2090) );
  NOR2_X1 U2116 ( .A1(n2094), .A2(n2079), .ZN(n2093) );
  XNOR2_X1 U2117 ( .A(n2095), .B(n2096), .ZN(Result_mul_27_) );
  XNOR2_X1 U2118 ( .A(n2097), .B(n2098), .ZN(n2095) );
  XNOR2_X1 U2119 ( .A(n2099), .B(n2100), .ZN(Result_mul_26_) );
  XOR2_X1 U2120 ( .A(n2101), .B(n2102), .Z(n2100) );
  XNOR2_X1 U2121 ( .A(n2103), .B(n2104), .ZN(Result_mul_25_) );
  XNOR2_X1 U2122 ( .A(n2105), .B(n2106), .ZN(n2103) );
  XOR2_X1 U2123 ( .A(n2107), .B(n2108), .Z(Result_mul_24_) );
  XNOR2_X1 U2124 ( .A(n2109), .B(n2110), .ZN(n2107) );
  XNOR2_X1 U2125 ( .A(n2111), .B(n2112), .ZN(Result_mul_23_) );
  NAND2_X1 U2126 ( .A1(n2113), .A2(n2114), .ZN(n2111) );
  XNOR2_X1 U2127 ( .A(n2115), .B(n2116), .ZN(Result_mul_22_) );
  XOR2_X1 U2128 ( .A(n2117), .B(n2118), .Z(n2116) );
  XNOR2_X1 U2129 ( .A(n2119), .B(n2120), .ZN(Result_mul_21_) );
  NAND2_X1 U2130 ( .A1(n2121), .A2(n2122), .ZN(n2119) );
  XOR2_X1 U2131 ( .A(n2123), .B(n2124), .Z(Result_mul_20_) );
  XNOR2_X1 U2132 ( .A(n2125), .B(n2126), .ZN(n2124) );
  XOR2_X1 U2133 ( .A(n2127), .B(n2128), .Z(Result_mul_1_) );
  NAND2_X1 U2134 ( .A1(n2129), .A2(n2130), .ZN(n2128) );
  XNOR2_X1 U2135 ( .A(n2131), .B(n2132), .ZN(Result_mul_19_) );
  NAND2_X1 U2136 ( .A1(n2133), .A2(n2134), .ZN(n2131) );
  XOR2_X1 U2137 ( .A(n2135), .B(n2136), .Z(Result_mul_18_) );
  XOR2_X1 U2138 ( .A(n2137), .B(n2138), .Z(n2136) );
  NOR2_X1 U2139 ( .A1(n2139), .A2(n2079), .ZN(n2138) );
  XNOR2_X1 U2140 ( .A(n2140), .B(n2141), .ZN(Result_mul_17_) );
  XOR2_X1 U2141 ( .A(n2142), .B(n2143), .Z(n2141) );
  NAND2_X1 U2142 ( .A1(b_15_), .A2(a_1_), .ZN(n2143) );
  XNOR2_X1 U2143 ( .A(n2144), .B(n2145), .ZN(Result_mul_16_) );
  XOR2_X1 U2144 ( .A(n2146), .B(n2147), .Z(n2145) );
  NAND2_X1 U2145 ( .A1(b_15_), .A2(a_0_), .ZN(n2147) );
  XOR2_X1 U2146 ( .A(n2148), .B(n2149), .Z(Result_mul_15_) );
  NOR2_X1 U2147 ( .A1(n2150), .A2(n2151), .ZN(Result_mul_14_) );
  NOR2_X1 U2148 ( .A1(n2152), .A2(n2153), .ZN(n2151) );
  INV_X1 U2149 ( .A(n2154), .ZN(n2152) );
  NAND2_X1 U2150 ( .A1(n2148), .A2(n2149), .ZN(n2154) );
  XOR2_X1 U2151 ( .A(n2155), .B(n2156), .Z(Result_mul_13_) );
  NAND2_X1 U2152 ( .A1(n2157), .A2(n2158), .ZN(n2156) );
  NAND2_X1 U2153 ( .A1(n2159), .A2(n2160), .ZN(n2158) );
  NAND2_X1 U2154 ( .A1(n2161), .A2(n2162), .ZN(n2160) );
  XOR2_X1 U2155 ( .A(n2163), .B(n2164), .Z(Result_mul_12_) );
  XOR2_X1 U2156 ( .A(n2165), .B(n2166), .Z(Result_mul_11_) );
  NOR2_X1 U2157 ( .A1(n2163), .A2(n2164), .ZN(n2166) );
  NOR2_X1 U2158 ( .A1(n2167), .A2(n2168), .ZN(n2165) );
  NOR2_X1 U2159 ( .A1(n2169), .A2(n2170), .ZN(n2167) );
  NOR2_X1 U2160 ( .A1(n2171), .A2(n2172), .ZN(n2170) );
  XOR2_X1 U2161 ( .A(n2037), .B(n2036), .Z(Result_mul_10_) );
  NAND3_X1 U2162 ( .A1(n2173), .A2(n2129), .A3(n2174), .ZN(Result_mul_0_) );
  NAND2_X1 U2163 ( .A1(a_0_), .A2(n2175), .ZN(n2174) );
  INV_X1 U2164 ( .A(n2176), .ZN(n2175) );
  NAND4_X1 U2165 ( .A1(n2176), .A2(n2177), .A3(n2178), .A4(n2179), .ZN(n2129)
         );
  NAND2_X1 U2166 ( .A1(n2180), .A2(n2130), .ZN(n2173) );
  NAND2_X1 U2167 ( .A1(n2181), .A2(n2182), .ZN(n2130) );
  NAND2_X1 U2168 ( .A1(n2178), .A2(n2179), .ZN(n2182) );
  XOR2_X1 U2169 ( .A(n2177), .B(n2176), .Z(n2181) );
  NOR2_X1 U2170 ( .A1(n2183), .A2(n2184), .ZN(n2176) );
  INV_X1 U2171 ( .A(n2185), .ZN(n2184) );
  NAND3_X1 U2172 ( .A1(b_0_), .A2(n2186), .A3(a_1_), .ZN(n2185) );
  NAND2_X1 U2173 ( .A1(n2187), .A2(n2188), .ZN(n2186) );
  NOR2_X1 U2174 ( .A1(n2188), .A2(n2187), .ZN(n2183) );
  INV_X1 U2175 ( .A(n2127), .ZN(n2180) );
  NAND2_X1 U2176 ( .A1(n2085), .A2(n2084), .ZN(n2127) );
  NAND3_X1 U2177 ( .A1(n2189), .A2(n2068), .A3(n2190), .ZN(n2084) );
  NAND3_X1 U2178 ( .A1(n2065), .A2(n2064), .A3(n2191), .ZN(n2190) );
  NAND3_X1 U2179 ( .A1(n2192), .A2(n2058), .A3(n2193), .ZN(n2064) );
  NAND3_X1 U2180 ( .A1(n2055), .A2(n2054), .A3(n2194), .ZN(n2193) );
  NAND3_X1 U2181 ( .A1(n2195), .A2(n2048), .A3(n2196), .ZN(n2054) );
  NAND3_X1 U2182 ( .A1(n2045), .A2(n2044), .A3(n2197), .ZN(n2196) );
  NAND3_X1 U2183 ( .A1(n2198), .A2(n2038), .A3(n2199), .ZN(n2044) );
  NAND3_X1 U2184 ( .A1(n2200), .A2(n2037), .A3(n2036), .ZN(n2199) );
  XOR2_X1 U2185 ( .A(n2043), .B(n2042), .Z(n2036) );
  INV_X1 U2186 ( .A(n2201), .ZN(n2037) );
  NOR3_X1 U2187 ( .A1(n2202), .A2(n2168), .A3(n2203), .ZN(n2201) );
  NOR3_X1 U2188 ( .A1(n2204), .A2(n2163), .A3(n2164), .ZN(n2203) );
  XNOR2_X1 U2189 ( .A(n2171), .B(n2172), .ZN(n2164) );
  INV_X1 U2190 ( .A(n2205), .ZN(n2163) );
  NAND3_X1 U2191 ( .A1(n2206), .A2(n2157), .A3(n2207), .ZN(n2205) );
  NAND2_X1 U2192 ( .A1(n2150), .A2(n2208), .ZN(n2207) );
  INV_X1 U2193 ( .A(n2155), .ZN(n2150) );
  NAND3_X1 U2194 ( .A1(n2149), .A2(n2148), .A3(n2153), .ZN(n2155) );
  XOR2_X1 U2195 ( .A(n2162), .B(n2161), .Z(n2153) );
  NAND2_X1 U2196 ( .A1(n2209), .A2(n2210), .ZN(n2148) );
  INV_X1 U2197 ( .A(n2211), .ZN(n2210) );
  NOR3_X1 U2198 ( .A1(n2212), .A2(n2213), .A3(n2079), .ZN(n2211) );
  NOR2_X1 U2199 ( .A1(n2146), .A2(n2144), .ZN(n2213) );
  NAND2_X1 U2200 ( .A1(n2144), .A2(n2146), .ZN(n2209) );
  NAND2_X1 U2201 ( .A1(n2214), .A2(n2215), .ZN(n2146) );
  NAND3_X1 U2202 ( .A1(a_1_), .A2(n2216), .A3(b_15_), .ZN(n2215) );
  INV_X1 U2203 ( .A(n2217), .ZN(n2216) );
  NOR2_X1 U2204 ( .A1(n2142), .A2(n2140), .ZN(n2217) );
  NAND2_X1 U2205 ( .A1(n2140), .A2(n2142), .ZN(n2214) );
  NAND2_X1 U2206 ( .A1(n2218), .A2(n2219), .ZN(n2142) );
  INV_X1 U2207 ( .A(n2220), .ZN(n2219) );
  NOR3_X1 U2208 ( .A1(n2139), .A2(n2221), .A3(n2079), .ZN(n2220) );
  NOR2_X1 U2209 ( .A1(n2137), .A2(n2135), .ZN(n2221) );
  NAND2_X1 U2210 ( .A1(n2135), .A2(n2137), .ZN(n2218) );
  NAND2_X1 U2211 ( .A1(n2133), .A2(n2222), .ZN(n2137) );
  NAND2_X1 U2212 ( .A1(n2132), .A2(n2134), .ZN(n2222) );
  NAND2_X1 U2213 ( .A1(n2223), .A2(n2224), .ZN(n2134) );
  INV_X1 U2214 ( .A(n2225), .ZN(n2224) );
  NAND2_X1 U2215 ( .A1(b_15_), .A2(a_3_), .ZN(n2223) );
  XOR2_X1 U2216 ( .A(n2226), .B(n2227), .Z(n2132) );
  XOR2_X1 U2217 ( .A(n2228), .B(n2229), .Z(n2226) );
  NOR2_X1 U2218 ( .A1(n2230), .A2(n2083), .ZN(n2229) );
  NAND2_X1 U2219 ( .A1(n2225), .A2(a_3_), .ZN(n2133) );
  NOR2_X1 U2220 ( .A1(n2231), .A2(n2232), .ZN(n2225) );
  INV_X1 U2221 ( .A(n2233), .ZN(n2232) );
  NAND2_X1 U2222 ( .A1(n2234), .A2(n2126), .ZN(n2233) );
  NAND2_X1 U2223 ( .A1(b_15_), .A2(a_4_), .ZN(n2126) );
  NAND2_X1 U2224 ( .A1(n2123), .A2(n2125), .ZN(n2234) );
  NOR2_X1 U2225 ( .A1(n2125), .A2(n2123), .ZN(n2231) );
  XNOR2_X1 U2226 ( .A(n2235), .B(n2236), .ZN(n2123) );
  NAND2_X1 U2227 ( .A1(n2237), .A2(n2238), .ZN(n2235) );
  NAND2_X1 U2228 ( .A1(n2121), .A2(n2239), .ZN(n2125) );
  NAND2_X1 U2229 ( .A1(n2120), .A2(n2122), .ZN(n2239) );
  NAND2_X1 U2230 ( .A1(n2240), .A2(n2241), .ZN(n2122) );
  INV_X1 U2231 ( .A(n2242), .ZN(n2241) );
  NAND2_X1 U2232 ( .A1(b_15_), .A2(a_5_), .ZN(n2240) );
  XNOR2_X1 U2233 ( .A(n2243), .B(n2244), .ZN(n2120) );
  XNOR2_X1 U2234 ( .A(n2245), .B(n2246), .ZN(n2243) );
  NOR2_X1 U2235 ( .A1(n2247), .A2(n2083), .ZN(n2246) );
  NAND2_X1 U2236 ( .A1(n2242), .A2(a_5_), .ZN(n2121) );
  NOR2_X1 U2237 ( .A1(n2248), .A2(n2249), .ZN(n2242) );
  INV_X1 U2238 ( .A(n2250), .ZN(n2249) );
  NAND2_X1 U2239 ( .A1(n2251), .A2(n2117), .ZN(n2250) );
  NAND2_X1 U2240 ( .A1(b_15_), .A2(a_6_), .ZN(n2117) );
  NAND2_X1 U2241 ( .A1(n2115), .A2(n2118), .ZN(n2251) );
  NOR2_X1 U2242 ( .A1(n2118), .A2(n2115), .ZN(n2248) );
  XOR2_X1 U2243 ( .A(n2252), .B(n2253), .Z(n2115) );
  XNOR2_X1 U2244 ( .A(n2254), .B(n2255), .ZN(n2253) );
  NAND2_X1 U2245 ( .A1(b_14_), .A2(a_7_), .ZN(n2255) );
  NAND2_X1 U2246 ( .A1(n2113), .A2(n2256), .ZN(n2118) );
  NAND2_X1 U2247 ( .A1(n2112), .A2(n2114), .ZN(n2256) );
  NAND2_X1 U2248 ( .A1(n2257), .A2(n2258), .ZN(n2114) );
  INV_X1 U2249 ( .A(n2259), .ZN(n2258) );
  NAND2_X1 U2250 ( .A1(b_15_), .A2(a_7_), .ZN(n2257) );
  XNOR2_X1 U2251 ( .A(n2260), .B(n2261), .ZN(n2112) );
  XOR2_X1 U2252 ( .A(n2262), .B(n2263), .Z(n2261) );
  NAND2_X1 U2253 ( .A1(b_14_), .A2(a_8_), .ZN(n2263) );
  NAND2_X1 U2254 ( .A1(n2259), .A2(a_7_), .ZN(n2113) );
  NOR2_X1 U2255 ( .A1(n2264), .A2(n2265), .ZN(n2259) );
  INV_X1 U2256 ( .A(n2266), .ZN(n2265) );
  NAND2_X1 U2257 ( .A1(n2267), .A2(n2110), .ZN(n2266) );
  NAND2_X1 U2258 ( .A1(b_15_), .A2(a_8_), .ZN(n2110) );
  NAND2_X1 U2259 ( .A1(n2108), .A2(n2109), .ZN(n2267) );
  NOR2_X1 U2260 ( .A1(n2109), .A2(n2108), .ZN(n2264) );
  XNOR2_X1 U2261 ( .A(n2268), .B(n2269), .ZN(n2108) );
  NAND2_X1 U2262 ( .A1(n2270), .A2(n2271), .ZN(n2268) );
  NAND2_X1 U2263 ( .A1(n2272), .A2(n2273), .ZN(n2109) );
  NAND2_X1 U2264 ( .A1(n2106), .A2(n2274), .ZN(n2273) );
  NAND2_X1 U2265 ( .A1(n2105), .A2(n2104), .ZN(n2274) );
  NOR2_X1 U2266 ( .A1(n2079), .A2(n2275), .ZN(n2106) );
  INV_X1 U2267 ( .A(n2276), .ZN(n2272) );
  NOR2_X1 U2268 ( .A1(n2104), .A2(n2105), .ZN(n2276) );
  NOR2_X1 U2269 ( .A1(n2277), .A2(n2278), .ZN(n2105) );
  NOR2_X1 U2270 ( .A1(n2101), .A2(n2279), .ZN(n2278) );
  NOR2_X1 U2271 ( .A1(n2102), .A2(n2099), .ZN(n2279) );
  NAND2_X1 U2272 ( .A1(b_15_), .A2(a_10_), .ZN(n2101) );
  INV_X1 U2273 ( .A(n2280), .ZN(n2277) );
  NAND2_X1 U2274 ( .A1(n2099), .A2(n2102), .ZN(n2280) );
  NAND2_X1 U2275 ( .A1(n2281), .A2(n2282), .ZN(n2102) );
  NAND2_X1 U2276 ( .A1(n2098), .A2(n2283), .ZN(n2282) );
  NAND2_X1 U2277 ( .A1(n2097), .A2(n2096), .ZN(n2283) );
  NOR2_X1 U2278 ( .A1(n2079), .A2(n2284), .ZN(n2098) );
  INV_X1 U2279 ( .A(b_15_), .ZN(n2079) );
  INV_X1 U2280 ( .A(n2285), .ZN(n2281) );
  NOR2_X1 U2281 ( .A1(n2096), .A2(n2097), .ZN(n2285) );
  NOR2_X1 U2282 ( .A1(n2286), .A2(n2287), .ZN(n2097) );
  INV_X1 U2283 ( .A(n2288), .ZN(n2287) );
  NAND3_X1 U2284 ( .A1(a_12_), .A2(n2289), .A3(b_15_), .ZN(n2288) );
  NAND2_X1 U2285 ( .A1(n2091), .A2(n2092), .ZN(n2289) );
  NOR2_X1 U2286 ( .A1(n2092), .A2(n2091), .ZN(n2286) );
  XNOR2_X1 U2287 ( .A(n2290), .B(n2291), .ZN(n2091) );
  XOR2_X1 U2288 ( .A(n2292), .B(n2293), .Z(n2290) );
  NAND2_X1 U2289 ( .A1(n2294), .A2(n2295), .ZN(n2092) );
  NAND2_X1 U2290 ( .A1(n2296), .A2(n2088), .ZN(n2295) );
  NAND2_X1 U2291 ( .A1(b_15_), .A2(a_13_), .ZN(n2088) );
  NAND2_X1 U2292 ( .A1(n2297), .A2(n2089), .ZN(n2296) );
  INV_X1 U2293 ( .A(n2086), .ZN(n2297) );
  NAND2_X1 U2294 ( .A1(n2298), .A2(n2086), .ZN(n2294) );
  INV_X1 U2295 ( .A(n2089), .ZN(n2298) );
  NAND2_X1 U2296 ( .A1(n2299), .A2(n2300), .ZN(n2089) );
  NAND2_X1 U2297 ( .A1(b_13_), .A2(n2301), .ZN(n2300) );
  NAND2_X1 U2298 ( .A1(n2077), .A2(n2302), .ZN(n2301) );
  NAND2_X1 U2299 ( .A1(a_15_), .A2(n2083), .ZN(n2302) );
  NAND2_X1 U2300 ( .A1(b_14_), .A2(n2303), .ZN(n2299) );
  NAND2_X1 U2301 ( .A1(n2081), .A2(n2304), .ZN(n2303) );
  NAND2_X1 U2302 ( .A1(a_14_), .A2(n2305), .ZN(n2304) );
  XOR2_X1 U2303 ( .A(n2306), .B(n2307), .Z(n2096) );
  XNOR2_X1 U2304 ( .A(n2308), .B(n2309), .ZN(n2306) );
  XNOR2_X1 U2305 ( .A(n2310), .B(n2311), .ZN(n2099) );
  XOR2_X1 U2306 ( .A(n2312), .B(n2313), .Z(n2310) );
  NAND2_X1 U2307 ( .A1(b_14_), .A2(a_11_), .ZN(n2312) );
  XNOR2_X1 U2308 ( .A(n2314), .B(n2315), .ZN(n2104) );
  XNOR2_X1 U2309 ( .A(n2316), .B(n2317), .ZN(n2315) );
  XNOR2_X1 U2310 ( .A(n2318), .B(n2319), .ZN(n2135) );
  XNOR2_X1 U2311 ( .A(n2320), .B(n2321), .ZN(n2318) );
  NOR2_X1 U2312 ( .A1(n2322), .A2(n2083), .ZN(n2321) );
  XOR2_X1 U2313 ( .A(n2323), .B(n2324), .Z(n2140) );
  XNOR2_X1 U2314 ( .A(n2325), .B(n2326), .ZN(n2324) );
  NAND2_X1 U2315 ( .A1(b_14_), .A2(a_2_), .ZN(n2326) );
  XOR2_X1 U2316 ( .A(n2327), .B(n2328), .Z(n2144) );
  XNOR2_X1 U2317 ( .A(n2329), .B(n2330), .ZN(n2328) );
  NAND2_X1 U2318 ( .A1(b_14_), .A2(a_1_), .ZN(n2330) );
  XNOR2_X1 U2319 ( .A(n2331), .B(n2332), .ZN(n2149) );
  XNOR2_X1 U2320 ( .A(n2333), .B(n2334), .ZN(n2331) );
  NOR2_X1 U2321 ( .A1(n2212), .A2(n2083), .ZN(n2334) );
  NAND3_X1 U2322 ( .A1(n2161), .A2(n2162), .A3(n2208), .ZN(n2157) );
  INV_X1 U2323 ( .A(n2159), .ZN(n2208) );
  XNOR2_X1 U2324 ( .A(n2335), .B(n2336), .ZN(n2159) );
  NAND2_X1 U2325 ( .A1(n2337), .A2(n2338), .ZN(n2162) );
  NAND3_X1 U2326 ( .A1(a_0_), .A2(n2339), .A3(b_14_), .ZN(n2338) );
  NAND2_X1 U2327 ( .A1(n2333), .A2(n2332), .ZN(n2339) );
  INV_X1 U2328 ( .A(n2340), .ZN(n2337) );
  NOR2_X1 U2329 ( .A1(n2332), .A2(n2333), .ZN(n2340) );
  NOR2_X1 U2330 ( .A1(n2341), .A2(n2342), .ZN(n2333) );
  NOR3_X1 U2331 ( .A1(n2343), .A2(n2344), .A3(n2083), .ZN(n2342) );
  INV_X1 U2332 ( .A(n2345), .ZN(n2344) );
  NAND2_X1 U2333 ( .A1(n2329), .A2(n2327), .ZN(n2345) );
  NOR2_X1 U2334 ( .A1(n2327), .A2(n2329), .ZN(n2341) );
  NOR2_X1 U2335 ( .A1(n2346), .A2(n2347), .ZN(n2329) );
  INV_X1 U2336 ( .A(n2348), .ZN(n2347) );
  NAND3_X1 U2337 ( .A1(a_2_), .A2(n2349), .A3(b_14_), .ZN(n2348) );
  NAND2_X1 U2338 ( .A1(n2325), .A2(n2323), .ZN(n2349) );
  NOR2_X1 U2339 ( .A1(n2323), .A2(n2325), .ZN(n2346) );
  NOR2_X1 U2340 ( .A1(n2350), .A2(n2351), .ZN(n2325) );
  NOR3_X1 U2341 ( .A1(n2322), .A2(n2352), .A3(n2083), .ZN(n2351) );
  INV_X1 U2342 ( .A(n2353), .ZN(n2352) );
  NAND2_X1 U2343 ( .A1(n2320), .A2(n2319), .ZN(n2353) );
  NOR2_X1 U2344 ( .A1(n2319), .A2(n2320), .ZN(n2350) );
  NOR2_X1 U2345 ( .A1(n2354), .A2(n2355), .ZN(n2320) );
  NOR3_X1 U2346 ( .A1(n2230), .A2(n2356), .A3(n2083), .ZN(n2355) );
  NOR2_X1 U2347 ( .A1(n2228), .A2(n2227), .ZN(n2356) );
  INV_X1 U2348 ( .A(n2357), .ZN(n2354) );
  NAND2_X1 U2349 ( .A1(n2227), .A2(n2228), .ZN(n2357) );
  NAND2_X1 U2350 ( .A1(n2237), .A2(n2358), .ZN(n2228) );
  NAND2_X1 U2351 ( .A1(n2236), .A2(n2238), .ZN(n2358) );
  NAND2_X1 U2352 ( .A1(n2359), .A2(n2360), .ZN(n2238) );
  NAND2_X1 U2353 ( .A1(b_14_), .A2(a_5_), .ZN(n2360) );
  XNOR2_X1 U2354 ( .A(n2361), .B(n2362), .ZN(n2236) );
  XOR2_X1 U2355 ( .A(n2363), .B(n2364), .Z(n2362) );
  NAND2_X1 U2356 ( .A1(b_13_), .A2(a_6_), .ZN(n2364) );
  INV_X1 U2357 ( .A(n2365), .ZN(n2237) );
  NOR2_X1 U2358 ( .A1(n2366), .A2(n2359), .ZN(n2365) );
  NOR2_X1 U2359 ( .A1(n2367), .A2(n2368), .ZN(n2359) );
  INV_X1 U2360 ( .A(n2369), .ZN(n2368) );
  NAND3_X1 U2361 ( .A1(a_6_), .A2(n2370), .A3(b_14_), .ZN(n2369) );
  NAND2_X1 U2362 ( .A1(n2245), .A2(n2244), .ZN(n2370) );
  NOR2_X1 U2363 ( .A1(n2244), .A2(n2245), .ZN(n2367) );
  NOR2_X1 U2364 ( .A1(n2371), .A2(n2372), .ZN(n2245) );
  INV_X1 U2365 ( .A(n2373), .ZN(n2372) );
  NAND3_X1 U2366 ( .A1(a_7_), .A2(n2374), .A3(b_14_), .ZN(n2373) );
  NAND2_X1 U2367 ( .A1(n2254), .A2(n2252), .ZN(n2374) );
  NOR2_X1 U2368 ( .A1(n2252), .A2(n2254), .ZN(n2371) );
  NOR2_X1 U2369 ( .A1(n2375), .A2(n2376), .ZN(n2254) );
  NOR3_X1 U2370 ( .A1(n2377), .A2(n2378), .A3(n2083), .ZN(n2376) );
  NOR2_X1 U2371 ( .A1(n2262), .A2(n2260), .ZN(n2378) );
  INV_X1 U2372 ( .A(n2379), .ZN(n2375) );
  NAND2_X1 U2373 ( .A1(n2260), .A2(n2262), .ZN(n2379) );
  NAND2_X1 U2374 ( .A1(n2270), .A2(n2380), .ZN(n2262) );
  NAND2_X1 U2375 ( .A1(n2269), .A2(n2271), .ZN(n2380) );
  NAND2_X1 U2376 ( .A1(n2381), .A2(n2382), .ZN(n2271) );
  NAND2_X1 U2377 ( .A1(b_14_), .A2(a_9_), .ZN(n2381) );
  XNOR2_X1 U2378 ( .A(n2383), .B(n2384), .ZN(n2269) );
  NAND2_X1 U2379 ( .A1(n2385), .A2(n2386), .ZN(n2383) );
  NAND2_X1 U2380 ( .A1(n2387), .A2(a_9_), .ZN(n2270) );
  INV_X1 U2381 ( .A(n2382), .ZN(n2387) );
  NAND2_X1 U2382 ( .A1(n2388), .A2(n2389), .ZN(n2382) );
  NAND2_X1 U2383 ( .A1(n2314), .A2(n2390), .ZN(n2389) );
  INV_X1 U2384 ( .A(n2391), .ZN(n2390) );
  NOR2_X1 U2385 ( .A1(n2317), .A2(n2316), .ZN(n2391) );
  XOR2_X1 U2386 ( .A(n2392), .B(n2393), .Z(n2314) );
  XNOR2_X1 U2387 ( .A(n2394), .B(n2395), .ZN(n2392) );
  NOR2_X1 U2388 ( .A1(n2284), .A2(n2305), .ZN(n2395) );
  NAND2_X1 U2389 ( .A1(n2316), .A2(n2317), .ZN(n2388) );
  NAND2_X1 U2390 ( .A1(b_14_), .A2(a_10_), .ZN(n2317) );
  NOR2_X1 U2391 ( .A1(n2396), .A2(n2397), .ZN(n2316) );
  NOR3_X1 U2392 ( .A1(n2284), .A2(n2398), .A3(n2083), .ZN(n2397) );
  INV_X1 U2393 ( .A(n2399), .ZN(n2398) );
  NAND2_X1 U2394 ( .A1(n2313), .A2(n2311), .ZN(n2399) );
  NOR2_X1 U2395 ( .A1(n2311), .A2(n2313), .ZN(n2396) );
  NOR2_X1 U2396 ( .A1(n2400), .A2(n2401), .ZN(n2313) );
  INV_X1 U2397 ( .A(n2402), .ZN(n2401) );
  NAND2_X1 U2398 ( .A1(n2308), .A2(n2403), .ZN(n2402) );
  NAND2_X1 U2399 ( .A1(n2309), .A2(n2307), .ZN(n2403) );
  NOR2_X1 U2400 ( .A1(n2083), .A2(n2094), .ZN(n2308) );
  NOR2_X1 U2401 ( .A1(n2307), .A2(n2309), .ZN(n2400) );
  NOR2_X1 U2402 ( .A1(n2404), .A2(n2405), .ZN(n2309) );
  INV_X1 U2403 ( .A(n2406), .ZN(n2405) );
  NAND2_X1 U2404 ( .A1(n2291), .A2(n2407), .ZN(n2406) );
  NAND2_X1 U2405 ( .A1(n2292), .A2(n2293), .ZN(n2407) );
  NOR2_X1 U2406 ( .A1(n2083), .A2(n2408), .ZN(n2291) );
  NOR2_X1 U2407 ( .A1(n2293), .A2(n2292), .ZN(n2404) );
  INV_X1 U2408 ( .A(n2409), .ZN(n2292) );
  NAND2_X1 U2409 ( .A1(n2410), .A2(n2411), .ZN(n2409) );
  NAND2_X1 U2410 ( .A1(b_12_), .A2(n2412), .ZN(n2411) );
  NAND2_X1 U2411 ( .A1(n2077), .A2(n2413), .ZN(n2412) );
  NAND2_X1 U2412 ( .A1(a_15_), .A2(n2305), .ZN(n2413) );
  NAND2_X1 U2413 ( .A1(b_13_), .A2(n2414), .ZN(n2410) );
  NAND2_X1 U2414 ( .A1(n2081), .A2(n2415), .ZN(n2414) );
  NAND2_X1 U2415 ( .A1(a_14_), .A2(n2416), .ZN(n2415) );
  NAND3_X1 U2416 ( .A1(b_14_), .A2(n2417), .A3(b_13_), .ZN(n2293) );
  XNOR2_X1 U2417 ( .A(n2418), .B(n2419), .ZN(n2307) );
  XNOR2_X1 U2418 ( .A(n2420), .B(n2421), .ZN(n2418) );
  XNOR2_X1 U2419 ( .A(n2422), .B(n2423), .ZN(n2311) );
  XOR2_X1 U2420 ( .A(n2424), .B(n2425), .Z(n2422) );
  XNOR2_X1 U2421 ( .A(n2426), .B(n2427), .ZN(n2260) );
  NAND2_X1 U2422 ( .A1(n2428), .A2(n2429), .ZN(n2426) );
  XOR2_X1 U2423 ( .A(n2430), .B(n2431), .Z(n2252) );
  XOR2_X1 U2424 ( .A(n2432), .B(n2433), .Z(n2431) );
  NAND2_X1 U2425 ( .A1(b_13_), .A2(a_8_), .ZN(n2433) );
  XNOR2_X1 U2426 ( .A(n2434), .B(n2435), .ZN(n2244) );
  XNOR2_X1 U2427 ( .A(n2436), .B(n2437), .ZN(n2435) );
  NAND2_X1 U2428 ( .A1(b_13_), .A2(a_7_), .ZN(n2437) );
  XNOR2_X1 U2429 ( .A(n2438), .B(n2439), .ZN(n2227) );
  NAND2_X1 U2430 ( .A1(n2440), .A2(n2441), .ZN(n2438) );
  XNOR2_X1 U2431 ( .A(n2442), .B(n2443), .ZN(n2319) );
  XNOR2_X1 U2432 ( .A(n2444), .B(n2445), .ZN(n2442) );
  NAND2_X1 U2433 ( .A1(b_13_), .A2(a_4_), .ZN(n2444) );
  XOR2_X1 U2434 ( .A(n2446), .B(n2447), .Z(n2323) );
  NAND2_X1 U2435 ( .A1(n2448), .A2(n2449), .ZN(n2446) );
  XOR2_X1 U2436 ( .A(n2450), .B(n2451), .Z(n2327) );
  XOR2_X1 U2437 ( .A(n2452), .B(n2453), .Z(n2451) );
  XOR2_X1 U2438 ( .A(n2454), .B(n2455), .Z(n2332) );
  XOR2_X1 U2439 ( .A(n2456), .B(n2457), .Z(n2454) );
  XOR2_X1 U2440 ( .A(n2458), .B(n2459), .Z(n2161) );
  XOR2_X1 U2441 ( .A(n2460), .B(n2461), .Z(n2458) );
  NAND2_X1 U2442 ( .A1(n2335), .A2(n2336), .ZN(n2206) );
  NAND2_X1 U2443 ( .A1(n2462), .A2(n2463), .ZN(n2336) );
  NAND2_X1 U2444 ( .A1(n2461), .A2(n2464), .ZN(n2463) );
  INV_X1 U2445 ( .A(n2465), .ZN(n2464) );
  NOR2_X1 U2446 ( .A1(n2460), .A2(n2459), .ZN(n2465) );
  NOR2_X1 U2447 ( .A1(n2305), .A2(n2212), .ZN(n2461) );
  NAND2_X1 U2448 ( .A1(n2459), .A2(n2460), .ZN(n2462) );
  NAND2_X1 U2449 ( .A1(n2466), .A2(n2467), .ZN(n2460) );
  NAND2_X1 U2450 ( .A1(n2457), .A2(n2468), .ZN(n2467) );
  NAND2_X1 U2451 ( .A1(n2455), .A2(n2469), .ZN(n2468) );
  INV_X1 U2452 ( .A(n2456), .ZN(n2469) );
  NOR2_X1 U2453 ( .A1(n2305), .A2(n2343), .ZN(n2457) );
  NAND2_X1 U2454 ( .A1(n2470), .A2(n2456), .ZN(n2466) );
  NAND2_X1 U2455 ( .A1(n2471), .A2(n2472), .ZN(n2456) );
  INV_X1 U2456 ( .A(n2473), .ZN(n2472) );
  NOR2_X1 U2457 ( .A1(n2453), .A2(n2474), .ZN(n2473) );
  NOR2_X1 U2458 ( .A1(n2450), .A2(n2452), .ZN(n2474) );
  NAND2_X1 U2459 ( .A1(b_13_), .A2(a_2_), .ZN(n2453) );
  NAND2_X1 U2460 ( .A1(n2450), .A2(n2452), .ZN(n2471) );
  NAND2_X1 U2461 ( .A1(n2448), .A2(n2475), .ZN(n2452) );
  NAND2_X1 U2462 ( .A1(n2447), .A2(n2449), .ZN(n2475) );
  NAND2_X1 U2463 ( .A1(n2476), .A2(n2477), .ZN(n2449) );
  NAND2_X1 U2464 ( .A1(b_13_), .A2(a_3_), .ZN(n2477) );
  INV_X1 U2465 ( .A(n2478), .ZN(n2476) );
  XOR2_X1 U2466 ( .A(n2479), .B(n2480), .Z(n2447) );
  XNOR2_X1 U2467 ( .A(n2481), .B(n2482), .ZN(n2479) );
  NAND2_X1 U2468 ( .A1(b_12_), .A2(a_4_), .ZN(n2481) );
  NAND2_X1 U2469 ( .A1(a_3_), .A2(n2478), .ZN(n2448) );
  NAND2_X1 U2470 ( .A1(n2483), .A2(n2484), .ZN(n2478) );
  NAND3_X1 U2471 ( .A1(a_4_), .A2(n2485), .A3(b_13_), .ZN(n2484) );
  INV_X1 U2472 ( .A(n2486), .ZN(n2485) );
  NOR2_X1 U2473 ( .A1(n2445), .A2(n2443), .ZN(n2486) );
  NAND2_X1 U2474 ( .A1(n2443), .A2(n2445), .ZN(n2483) );
  NAND2_X1 U2475 ( .A1(n2440), .A2(n2487), .ZN(n2445) );
  NAND2_X1 U2476 ( .A1(n2439), .A2(n2441), .ZN(n2487) );
  NAND2_X1 U2477 ( .A1(n2488), .A2(n2489), .ZN(n2441) );
  NAND2_X1 U2478 ( .A1(b_13_), .A2(a_5_), .ZN(n2489) );
  XOR2_X1 U2479 ( .A(n2490), .B(n2491), .Z(n2439) );
  XOR2_X1 U2480 ( .A(n2492), .B(n2493), .Z(n2490) );
  NOR2_X1 U2481 ( .A1(n2247), .A2(n2416), .ZN(n2493) );
  NAND2_X1 U2482 ( .A1(a_5_), .A2(n2494), .ZN(n2440) );
  INV_X1 U2483 ( .A(n2488), .ZN(n2494) );
  NOR2_X1 U2484 ( .A1(n2495), .A2(n2496), .ZN(n2488) );
  NOR3_X1 U2485 ( .A1(n2247), .A2(n2497), .A3(n2305), .ZN(n2496) );
  NOR2_X1 U2486 ( .A1(n2361), .A2(n2363), .ZN(n2497) );
  INV_X1 U2487 ( .A(n2498), .ZN(n2495) );
  NAND2_X1 U2488 ( .A1(n2361), .A2(n2363), .ZN(n2498) );
  NAND2_X1 U2489 ( .A1(n2499), .A2(n2500), .ZN(n2363) );
  NAND3_X1 U2490 ( .A1(a_7_), .A2(n2501), .A3(b_13_), .ZN(n2500) );
  NAND2_X1 U2491 ( .A1(n2434), .A2(n2436), .ZN(n2501) );
  INV_X1 U2492 ( .A(n2502), .ZN(n2499) );
  NOR2_X1 U2493 ( .A1(n2434), .A2(n2436), .ZN(n2502) );
  NOR2_X1 U2494 ( .A1(n2503), .A2(n2504), .ZN(n2436) );
  NOR3_X1 U2495 ( .A1(n2377), .A2(n2505), .A3(n2305), .ZN(n2504) );
  NOR2_X1 U2496 ( .A1(n2432), .A2(n2430), .ZN(n2505) );
  INV_X1 U2497 ( .A(n2506), .ZN(n2503) );
  NAND2_X1 U2498 ( .A1(n2430), .A2(n2432), .ZN(n2506) );
  NAND2_X1 U2499 ( .A1(n2428), .A2(n2507), .ZN(n2432) );
  NAND2_X1 U2500 ( .A1(n2427), .A2(n2429), .ZN(n2507) );
  NAND2_X1 U2501 ( .A1(n2508), .A2(n2509), .ZN(n2429) );
  NAND2_X1 U2502 ( .A1(b_13_), .A2(a_9_), .ZN(n2509) );
  INV_X1 U2503 ( .A(n2510), .ZN(n2508) );
  XNOR2_X1 U2504 ( .A(n2511), .B(n2512), .ZN(n2427) );
  NAND2_X1 U2505 ( .A1(n2513), .A2(n2514), .ZN(n2511) );
  NAND2_X1 U2506 ( .A1(a_9_), .A2(n2510), .ZN(n2428) );
  NAND2_X1 U2507 ( .A1(n2385), .A2(n2515), .ZN(n2510) );
  NAND2_X1 U2508 ( .A1(n2384), .A2(n2386), .ZN(n2515) );
  NAND2_X1 U2509 ( .A1(n2516), .A2(n2517), .ZN(n2386) );
  NAND2_X1 U2510 ( .A1(b_13_), .A2(a_10_), .ZN(n2517) );
  XNOR2_X1 U2511 ( .A(n2518), .B(n2519), .ZN(n2384) );
  XNOR2_X1 U2512 ( .A(n2520), .B(n2521), .ZN(n2518) );
  NOR2_X1 U2513 ( .A1(n2284), .A2(n2416), .ZN(n2521) );
  INV_X1 U2514 ( .A(n2522), .ZN(n2385) );
  NOR2_X1 U2515 ( .A1(n2523), .A2(n2516), .ZN(n2522) );
  NOR2_X1 U2516 ( .A1(n2524), .A2(n2525), .ZN(n2516) );
  INV_X1 U2517 ( .A(n2526), .ZN(n2525) );
  NAND3_X1 U2518 ( .A1(a_11_), .A2(n2527), .A3(b_13_), .ZN(n2526) );
  NAND2_X1 U2519 ( .A1(n2393), .A2(n2394), .ZN(n2527) );
  NOR2_X1 U2520 ( .A1(n2393), .A2(n2394), .ZN(n2524) );
  NOR2_X1 U2521 ( .A1(n2528), .A2(n2529), .ZN(n2394) );
  INV_X1 U2522 ( .A(n2530), .ZN(n2529) );
  NAND2_X1 U2523 ( .A1(n2425), .A2(n2531), .ZN(n2530) );
  NAND2_X1 U2524 ( .A1(n2423), .A2(n2424), .ZN(n2531) );
  NOR2_X1 U2525 ( .A1(n2305), .A2(n2094), .ZN(n2425) );
  NOR2_X1 U2526 ( .A1(n2423), .A2(n2424), .ZN(n2528) );
  NAND2_X1 U2527 ( .A1(n2532), .A2(n2533), .ZN(n2424) );
  NAND2_X1 U2528 ( .A1(n2534), .A2(n2421), .ZN(n2533) );
  NAND3_X1 U2529 ( .A1(b_12_), .A2(n2417), .A3(b_13_), .ZN(n2421) );
  NAND2_X1 U2530 ( .A1(n2419), .A2(n2420), .ZN(n2534) );
  INV_X1 U2531 ( .A(n2535), .ZN(n2532) );
  NOR2_X1 U2532 ( .A1(n2420), .A2(n2419), .ZN(n2535) );
  NAND2_X1 U2533 ( .A1(n2536), .A2(n2537), .ZN(n2420) );
  NAND2_X1 U2534 ( .A1(b_11_), .A2(n2538), .ZN(n2537) );
  NAND2_X1 U2535 ( .A1(n2077), .A2(n2539), .ZN(n2538) );
  NAND2_X1 U2536 ( .A1(a_15_), .A2(n2416), .ZN(n2539) );
  NAND2_X1 U2537 ( .A1(b_12_), .A2(n2540), .ZN(n2536) );
  NAND2_X1 U2538 ( .A1(n2081), .A2(n2541), .ZN(n2540) );
  NAND2_X1 U2539 ( .A1(a_14_), .A2(n2542), .ZN(n2541) );
  XNOR2_X1 U2540 ( .A(n2543), .B(n2544), .ZN(n2423) );
  XOR2_X1 U2541 ( .A(n2545), .B(n2546), .Z(n2543) );
  XNOR2_X1 U2542 ( .A(n2547), .B(n2548), .ZN(n2393) );
  XOR2_X1 U2543 ( .A(n2549), .B(n2550), .Z(n2547) );
  XNOR2_X1 U2544 ( .A(n2551), .B(n2552), .ZN(n2430) );
  NAND2_X1 U2545 ( .A1(n2553), .A2(n2554), .ZN(n2551) );
  XOR2_X1 U2546 ( .A(n2555), .B(n2556), .Z(n2434) );
  XOR2_X1 U2547 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND2_X1 U2548 ( .A1(b_12_), .A2(a_8_), .ZN(n2558) );
  XNOR2_X1 U2549 ( .A(n2559), .B(n2560), .ZN(n2361) );
  XOR2_X1 U2550 ( .A(n2561), .B(n2562), .Z(n2560) );
  NAND2_X1 U2551 ( .A1(b_12_), .A2(a_7_), .ZN(n2562) );
  XNOR2_X1 U2552 ( .A(n2563), .B(n2564), .ZN(n2443) );
  NAND2_X1 U2553 ( .A1(n2565), .A2(n2566), .ZN(n2563) );
  XNOR2_X1 U2554 ( .A(n2567), .B(n2568), .ZN(n2450) );
  NAND2_X1 U2555 ( .A1(n2569), .A2(n2570), .ZN(n2567) );
  INV_X1 U2556 ( .A(n2455), .ZN(n2470) );
  XNOR2_X1 U2557 ( .A(n2571), .B(n2572), .ZN(n2455) );
  XNOR2_X1 U2558 ( .A(n2573), .B(n2574), .ZN(n2571) );
  NAND2_X1 U2559 ( .A1(b_12_), .A2(a_2_), .ZN(n2573) );
  XOR2_X1 U2560 ( .A(n2575), .B(n2576), .Z(n2459) );
  XOR2_X1 U2561 ( .A(n2577), .B(n2578), .Z(n2576) );
  XOR2_X1 U2562 ( .A(n2579), .B(n2580), .Z(n2335) );
  XOR2_X1 U2563 ( .A(n2581), .B(n2582), .Z(n2579) );
  NOR2_X1 U2564 ( .A1(n2212), .A2(n2416), .ZN(n2582) );
  NOR3_X1 U2565 ( .A1(n2172), .A2(n2171), .A3(n2204), .ZN(n2168) );
  INV_X1 U2566 ( .A(n2169), .ZN(n2204) );
  NOR2_X1 U2567 ( .A1(n2583), .A2(n2202), .ZN(n2169) );
  INV_X1 U2568 ( .A(n2584), .ZN(n2583) );
  NAND2_X1 U2569 ( .A1(n2585), .A2(n2586), .ZN(n2584) );
  NOR2_X1 U2570 ( .A1(n2587), .A2(n2588), .ZN(n2171) );
  NOR3_X1 U2571 ( .A1(n2212), .A2(n2589), .A3(n2416), .ZN(n2588) );
  NOR2_X1 U2572 ( .A1(n2581), .A2(n2580), .ZN(n2589) );
  INV_X1 U2573 ( .A(n2590), .ZN(n2587) );
  NAND2_X1 U2574 ( .A1(n2580), .A2(n2581), .ZN(n2590) );
  NAND2_X1 U2575 ( .A1(n2591), .A2(n2592), .ZN(n2581) );
  NAND2_X1 U2576 ( .A1(n2578), .A2(n2593), .ZN(n2592) );
  NAND2_X1 U2577 ( .A1(n2577), .A2(n2575), .ZN(n2593) );
  NOR2_X1 U2578 ( .A1(n2416), .A2(n2343), .ZN(n2578) );
  INV_X1 U2579 ( .A(n2594), .ZN(n2591) );
  NOR2_X1 U2580 ( .A1(n2575), .A2(n2577), .ZN(n2594) );
  NOR2_X1 U2581 ( .A1(n2595), .A2(n2596), .ZN(n2577) );
  NOR3_X1 U2582 ( .A1(n2139), .A2(n2597), .A3(n2416), .ZN(n2596) );
  NOR2_X1 U2583 ( .A1(n2574), .A2(n2572), .ZN(n2597) );
  INV_X1 U2584 ( .A(n2598), .ZN(n2595) );
  NAND2_X1 U2585 ( .A1(n2572), .A2(n2574), .ZN(n2598) );
  NAND2_X1 U2586 ( .A1(n2569), .A2(n2599), .ZN(n2574) );
  NAND2_X1 U2587 ( .A1(n2568), .A2(n2570), .ZN(n2599) );
  NAND2_X1 U2588 ( .A1(n2600), .A2(n2601), .ZN(n2570) );
  NAND2_X1 U2589 ( .A1(b_12_), .A2(a_3_), .ZN(n2601) );
  XNOR2_X1 U2590 ( .A(n2602), .B(n2603), .ZN(n2568) );
  XOR2_X1 U2591 ( .A(n2604), .B(n2605), .Z(n2603) );
  NAND2_X1 U2592 ( .A1(b_11_), .A2(a_4_), .ZN(n2605) );
  NAND2_X1 U2593 ( .A1(a_3_), .A2(n2606), .ZN(n2569) );
  INV_X1 U2594 ( .A(n2600), .ZN(n2606) );
  NOR2_X1 U2595 ( .A1(n2607), .A2(n2608), .ZN(n2600) );
  NOR3_X1 U2596 ( .A1(n2230), .A2(n2609), .A3(n2416), .ZN(n2608) );
  NOR2_X1 U2597 ( .A1(n2482), .A2(n2480), .ZN(n2609) );
  INV_X1 U2598 ( .A(n2610), .ZN(n2607) );
  NAND2_X1 U2599 ( .A1(n2480), .A2(n2482), .ZN(n2610) );
  NAND2_X1 U2600 ( .A1(n2565), .A2(n2611), .ZN(n2482) );
  NAND2_X1 U2601 ( .A1(n2564), .A2(n2566), .ZN(n2611) );
  NAND2_X1 U2602 ( .A1(n2612), .A2(n2613), .ZN(n2566) );
  NAND2_X1 U2603 ( .A1(b_12_), .A2(a_5_), .ZN(n2613) );
  XOR2_X1 U2604 ( .A(n2614), .B(n2615), .Z(n2564) );
  XNOR2_X1 U2605 ( .A(n2616), .B(n2617), .ZN(n2615) );
  NAND2_X1 U2606 ( .A1(b_11_), .A2(a_6_), .ZN(n2617) );
  NAND2_X1 U2607 ( .A1(a_5_), .A2(n2618), .ZN(n2565) );
  INV_X1 U2608 ( .A(n2612), .ZN(n2618) );
  NOR2_X1 U2609 ( .A1(n2619), .A2(n2620), .ZN(n2612) );
  NOR3_X1 U2610 ( .A1(n2247), .A2(n2621), .A3(n2416), .ZN(n2620) );
  NOR2_X1 U2611 ( .A1(n2492), .A2(n2491), .ZN(n2621) );
  INV_X1 U2612 ( .A(n2622), .ZN(n2619) );
  NAND2_X1 U2613 ( .A1(n2491), .A2(n2492), .ZN(n2622) );
  NAND2_X1 U2614 ( .A1(n2623), .A2(n2624), .ZN(n2492) );
  INV_X1 U2615 ( .A(n2625), .ZN(n2624) );
  NOR3_X1 U2616 ( .A1(n2626), .A2(n2627), .A3(n2416), .ZN(n2625) );
  NOR2_X1 U2617 ( .A1(n2561), .A2(n2559), .ZN(n2627) );
  NAND2_X1 U2618 ( .A1(n2559), .A2(n2561), .ZN(n2623) );
  NAND2_X1 U2619 ( .A1(n2628), .A2(n2629), .ZN(n2561) );
  INV_X1 U2620 ( .A(n2630), .ZN(n2629) );
  NOR3_X1 U2621 ( .A1(n2377), .A2(n2631), .A3(n2416), .ZN(n2630) );
  NOR2_X1 U2622 ( .A1(n2557), .A2(n2555), .ZN(n2631) );
  NAND2_X1 U2623 ( .A1(n2555), .A2(n2557), .ZN(n2628) );
  NAND2_X1 U2624 ( .A1(n2553), .A2(n2632), .ZN(n2557) );
  NAND2_X1 U2625 ( .A1(n2552), .A2(n2554), .ZN(n2632) );
  NAND2_X1 U2626 ( .A1(n2633), .A2(n2634), .ZN(n2554) );
  NAND2_X1 U2627 ( .A1(b_12_), .A2(a_9_), .ZN(n2634) );
  INV_X1 U2628 ( .A(n2635), .ZN(n2633) );
  XNOR2_X1 U2629 ( .A(n2636), .B(n2637), .ZN(n2552) );
  NAND2_X1 U2630 ( .A1(n2638), .A2(n2639), .ZN(n2636) );
  NAND2_X1 U2631 ( .A1(a_9_), .A2(n2635), .ZN(n2553) );
  NAND2_X1 U2632 ( .A1(n2513), .A2(n2640), .ZN(n2635) );
  NAND2_X1 U2633 ( .A1(n2512), .A2(n2514), .ZN(n2640) );
  NAND2_X1 U2634 ( .A1(n2641), .A2(n2642), .ZN(n2514) );
  NAND2_X1 U2635 ( .A1(b_12_), .A2(a_10_), .ZN(n2642) );
  XOR2_X1 U2636 ( .A(n2643), .B(n2644), .Z(n2512) );
  XOR2_X1 U2637 ( .A(n2645), .B(n2646), .Z(n2643) );
  NAND2_X1 U2638 ( .A1(a_10_), .A2(n2647), .ZN(n2513) );
  INV_X1 U2639 ( .A(n2641), .ZN(n2647) );
  NOR2_X1 U2640 ( .A1(n2648), .A2(n2649), .ZN(n2641) );
  NOR3_X1 U2641 ( .A1(n2284), .A2(n2650), .A3(n2416), .ZN(n2649) );
  NOR2_X1 U2642 ( .A1(n2519), .A2(n2520), .ZN(n2650) );
  INV_X1 U2643 ( .A(n2651), .ZN(n2648) );
  NAND2_X1 U2644 ( .A1(n2520), .A2(n2519), .ZN(n2651) );
  XNOR2_X1 U2645 ( .A(n2652), .B(n2653), .ZN(n2519) );
  XNOR2_X1 U2646 ( .A(n2654), .B(n2655), .ZN(n2652) );
  NOR2_X1 U2647 ( .A1(n2656), .A2(n2657), .ZN(n2520) );
  NOR2_X1 U2648 ( .A1(n2658), .A2(n2549), .ZN(n2657) );
  INV_X1 U2649 ( .A(n2659), .ZN(n2658) );
  NAND2_X1 U2650 ( .A1(n2548), .A2(n2550), .ZN(n2659) );
  NOR2_X1 U2651 ( .A1(n2550), .A2(n2548), .ZN(n2656) );
  XOR2_X1 U2652 ( .A(n2660), .B(n2661), .Z(n2548) );
  XOR2_X1 U2653 ( .A(n2662), .B(n2663), .Z(n2660) );
  NAND2_X1 U2654 ( .A1(n2664), .A2(n2665), .ZN(n2550) );
  NAND2_X1 U2655 ( .A1(n2544), .A2(n2666), .ZN(n2665) );
  INV_X1 U2656 ( .A(n2667), .ZN(n2666) );
  NOR2_X1 U2657 ( .A1(n2545), .A2(n2546), .ZN(n2667) );
  NOR2_X1 U2658 ( .A1(n2416), .A2(n2408), .ZN(n2544) );
  NAND2_X1 U2659 ( .A1(n2546), .A2(n2545), .ZN(n2664) );
  NAND2_X1 U2660 ( .A1(n2668), .A2(n2669), .ZN(n2545) );
  NAND2_X1 U2661 ( .A1(b_10_), .A2(n2670), .ZN(n2669) );
  NAND2_X1 U2662 ( .A1(n2077), .A2(n2671), .ZN(n2670) );
  NAND2_X1 U2663 ( .A1(a_15_), .A2(n2542), .ZN(n2671) );
  NAND2_X1 U2664 ( .A1(b_11_), .A2(n2672), .ZN(n2668) );
  NAND2_X1 U2665 ( .A1(n2081), .A2(n2673), .ZN(n2672) );
  NAND2_X1 U2666 ( .A1(a_14_), .A2(n2674), .ZN(n2673) );
  NOR3_X1 U2667 ( .A1(n2542), .A2(n2675), .A3(n2416), .ZN(n2546) );
  XOR2_X1 U2668 ( .A(n2676), .B(n2677), .Z(n2555) );
  XNOR2_X1 U2669 ( .A(n2678), .B(n2679), .ZN(n2677) );
  XOR2_X1 U2670 ( .A(n2680), .B(n2681), .Z(n2559) );
  XOR2_X1 U2671 ( .A(n2682), .B(n2683), .Z(n2680) );
  XNOR2_X1 U2672 ( .A(n2684), .B(n2685), .ZN(n2491) );
  XNOR2_X1 U2673 ( .A(n2686), .B(n2687), .ZN(n2684) );
  NOR2_X1 U2674 ( .A1(n2626), .A2(n2542), .ZN(n2687) );
  XNOR2_X1 U2675 ( .A(n2688), .B(n2689), .ZN(n2480) );
  NAND2_X1 U2676 ( .A1(n2690), .A2(n2691), .ZN(n2688) );
  XNOR2_X1 U2677 ( .A(n2692), .B(n2693), .ZN(n2572) );
  NAND2_X1 U2678 ( .A1(n2694), .A2(n2695), .ZN(n2692) );
  XOR2_X1 U2679 ( .A(n2696), .B(n2697), .Z(n2575) );
  XOR2_X1 U2680 ( .A(n2698), .B(n2699), .Z(n2697) );
  NAND2_X1 U2681 ( .A1(b_11_), .A2(a_2_), .ZN(n2699) );
  XNOR2_X1 U2682 ( .A(n2700), .B(n2701), .ZN(n2580) );
  XOR2_X1 U2683 ( .A(n2702), .B(n2703), .Z(n2701) );
  NAND2_X1 U2684 ( .A1(b_11_), .A2(a_1_), .ZN(n2703) );
  XNOR2_X1 U2685 ( .A(n2704), .B(n2705), .ZN(n2172) );
  XOR2_X1 U2686 ( .A(n2706), .B(n2707), .Z(n2704) );
  NOR2_X1 U2687 ( .A1(n2212), .A2(n2542), .ZN(n2707) );
  NOR2_X1 U2688 ( .A1(n2586), .A2(n2585), .ZN(n2202) );
  NOR2_X1 U2689 ( .A1(n2708), .A2(n2709), .ZN(n2585) );
  NOR3_X1 U2690 ( .A1(n2212), .A2(n2710), .A3(n2542), .ZN(n2709) );
  NOR2_X1 U2691 ( .A1(n2706), .A2(n2705), .ZN(n2710) );
  INV_X1 U2692 ( .A(n2711), .ZN(n2708) );
  NAND2_X1 U2693 ( .A1(n2705), .A2(n2706), .ZN(n2711) );
  NAND2_X1 U2694 ( .A1(n2712), .A2(n2713), .ZN(n2706) );
  INV_X1 U2695 ( .A(n2714), .ZN(n2713) );
  NOR3_X1 U2696 ( .A1(n2343), .A2(n2715), .A3(n2542), .ZN(n2714) );
  NOR2_X1 U2697 ( .A1(n2702), .A2(n2700), .ZN(n2715) );
  NAND2_X1 U2698 ( .A1(n2700), .A2(n2702), .ZN(n2712) );
  NAND2_X1 U2699 ( .A1(n2716), .A2(n2717), .ZN(n2702) );
  INV_X1 U2700 ( .A(n2718), .ZN(n2717) );
  NOR3_X1 U2701 ( .A1(n2139), .A2(n2719), .A3(n2542), .ZN(n2718) );
  NOR2_X1 U2702 ( .A1(n2698), .A2(n2696), .ZN(n2719) );
  NAND2_X1 U2703 ( .A1(n2696), .A2(n2698), .ZN(n2716) );
  NAND2_X1 U2704 ( .A1(n2694), .A2(n2720), .ZN(n2698) );
  NAND2_X1 U2705 ( .A1(n2693), .A2(n2695), .ZN(n2720) );
  NAND2_X1 U2706 ( .A1(n2721), .A2(n2722), .ZN(n2695) );
  NAND2_X1 U2707 ( .A1(b_11_), .A2(a_3_), .ZN(n2722) );
  XOR2_X1 U2708 ( .A(n2723), .B(n2724), .Z(n2693) );
  XOR2_X1 U2709 ( .A(n2725), .B(n2726), .Z(n2723) );
  NOR2_X1 U2710 ( .A1(n2230), .A2(n2674), .ZN(n2726) );
  NAND2_X1 U2711 ( .A1(a_3_), .A2(n2727), .ZN(n2694) );
  INV_X1 U2712 ( .A(n2721), .ZN(n2727) );
  NOR2_X1 U2713 ( .A1(n2728), .A2(n2729), .ZN(n2721) );
  NOR3_X1 U2714 ( .A1(n2230), .A2(n2730), .A3(n2542), .ZN(n2729) );
  NOR2_X1 U2715 ( .A1(n2604), .A2(n2602), .ZN(n2730) );
  INV_X1 U2716 ( .A(n2731), .ZN(n2728) );
  NAND2_X1 U2717 ( .A1(n2602), .A2(n2604), .ZN(n2731) );
  NAND2_X1 U2718 ( .A1(n2690), .A2(n2732), .ZN(n2604) );
  NAND2_X1 U2719 ( .A1(n2689), .A2(n2691), .ZN(n2732) );
  NAND2_X1 U2720 ( .A1(n2733), .A2(n2734), .ZN(n2691) );
  NAND2_X1 U2721 ( .A1(b_11_), .A2(a_5_), .ZN(n2734) );
  INV_X1 U2722 ( .A(n2735), .ZN(n2733) );
  XNOR2_X1 U2723 ( .A(n2736), .B(n2737), .ZN(n2689) );
  XNOR2_X1 U2724 ( .A(n2738), .B(n2739), .ZN(n2736) );
  NOR2_X1 U2725 ( .A1(n2247), .A2(n2674), .ZN(n2739) );
  NAND2_X1 U2726 ( .A1(a_5_), .A2(n2735), .ZN(n2690) );
  NAND2_X1 U2727 ( .A1(n2740), .A2(n2741), .ZN(n2735) );
  NAND3_X1 U2728 ( .A1(a_6_), .A2(n2742), .A3(b_11_), .ZN(n2741) );
  NAND2_X1 U2729 ( .A1(n2616), .A2(n2614), .ZN(n2742) );
  INV_X1 U2730 ( .A(n2743), .ZN(n2740) );
  NOR2_X1 U2731 ( .A1(n2614), .A2(n2616), .ZN(n2743) );
  NOR2_X1 U2732 ( .A1(n2744), .A2(n2745), .ZN(n2616) );
  NOR3_X1 U2733 ( .A1(n2626), .A2(n2746), .A3(n2542), .ZN(n2745) );
  INV_X1 U2734 ( .A(n2747), .ZN(n2746) );
  NAND2_X1 U2735 ( .A1(n2686), .A2(n2685), .ZN(n2747) );
  NOR2_X1 U2736 ( .A1(n2685), .A2(n2686), .ZN(n2744) );
  NOR2_X1 U2737 ( .A1(n2748), .A2(n2749), .ZN(n2686) );
  INV_X1 U2738 ( .A(n2750), .ZN(n2749) );
  NAND2_X1 U2739 ( .A1(n2683), .A2(n2751), .ZN(n2750) );
  NAND2_X1 U2740 ( .A1(n2681), .A2(n2682), .ZN(n2751) );
  NOR2_X1 U2741 ( .A1(n2542), .A2(n2377), .ZN(n2683) );
  NOR2_X1 U2742 ( .A1(n2682), .A2(n2681), .ZN(n2748) );
  XOR2_X1 U2743 ( .A(n2752), .B(n2753), .Z(n2681) );
  NAND2_X1 U2744 ( .A1(n2754), .A2(n2755), .ZN(n2752) );
  NAND2_X1 U2745 ( .A1(n2756), .A2(n2757), .ZN(n2682) );
  NAND2_X1 U2746 ( .A1(n2676), .A2(n2758), .ZN(n2757) );
  NAND2_X1 U2747 ( .A1(n2679), .A2(n2678), .ZN(n2758) );
  XOR2_X1 U2748 ( .A(n2759), .B(n2760), .Z(n2676) );
  XOR2_X1 U2749 ( .A(n2761), .B(n2762), .Z(n2760) );
  INV_X1 U2750 ( .A(n2763), .ZN(n2756) );
  NOR2_X1 U2751 ( .A1(n2678), .A2(n2679), .ZN(n2763) );
  NOR2_X1 U2752 ( .A1(n2542), .A2(n2275), .ZN(n2679) );
  NAND2_X1 U2753 ( .A1(n2638), .A2(n2764), .ZN(n2678) );
  NAND2_X1 U2754 ( .A1(n2637), .A2(n2639), .ZN(n2764) );
  NAND2_X1 U2755 ( .A1(n2765), .A2(n2766), .ZN(n2639) );
  NAND2_X1 U2756 ( .A1(b_11_), .A2(a_10_), .ZN(n2765) );
  XNOR2_X1 U2757 ( .A(n2767), .B(n2768), .ZN(n2637) );
  XOR2_X1 U2758 ( .A(n2769), .B(n2770), .Z(n2767) );
  NAND2_X1 U2759 ( .A1(b_10_), .A2(a_11_), .ZN(n2769) );
  NAND2_X1 U2760 ( .A1(n2771), .A2(a_10_), .ZN(n2638) );
  INV_X1 U2761 ( .A(n2766), .ZN(n2771) );
  NAND2_X1 U2762 ( .A1(n2772), .A2(n2773), .ZN(n2766) );
  INV_X1 U2763 ( .A(n2774), .ZN(n2773) );
  NOR2_X1 U2764 ( .A1(n2644), .A2(n2775), .ZN(n2774) );
  NOR2_X1 U2765 ( .A1(n2645), .A2(n2646), .ZN(n2775) );
  XNOR2_X1 U2766 ( .A(n2776), .B(n2777), .ZN(n2644) );
  XNOR2_X1 U2767 ( .A(n2778), .B(n2779), .ZN(n2776) );
  NAND2_X1 U2768 ( .A1(n2646), .A2(n2645), .ZN(n2772) );
  NOR2_X1 U2769 ( .A1(n2780), .A2(n2781), .ZN(n2646) );
  INV_X1 U2770 ( .A(n2782), .ZN(n2781) );
  NAND2_X1 U2771 ( .A1(n2654), .A2(n2783), .ZN(n2782) );
  NAND2_X1 U2772 ( .A1(n2655), .A2(n2653), .ZN(n2783) );
  NOR2_X1 U2773 ( .A1(n2542), .A2(n2094), .ZN(n2654) );
  NOR2_X1 U2774 ( .A1(n2653), .A2(n2655), .ZN(n2780) );
  NOR2_X1 U2775 ( .A1(n2784), .A2(n2785), .ZN(n2655) );
  INV_X1 U2776 ( .A(n2786), .ZN(n2785) );
  NAND2_X1 U2777 ( .A1(n2661), .A2(n2787), .ZN(n2786) );
  NAND2_X1 U2778 ( .A1(n2662), .A2(n2663), .ZN(n2787) );
  NOR2_X1 U2779 ( .A1(n2542), .A2(n2408), .ZN(n2661) );
  NOR2_X1 U2780 ( .A1(n2663), .A2(n2662), .ZN(n2784) );
  INV_X1 U2781 ( .A(n2788), .ZN(n2662) );
  NAND2_X1 U2782 ( .A1(n2789), .A2(n2790), .ZN(n2788) );
  NAND2_X1 U2783 ( .A1(b_10_), .A2(n2791), .ZN(n2790) );
  NAND2_X1 U2784 ( .A1(n2081), .A2(n2792), .ZN(n2791) );
  NAND2_X1 U2785 ( .A1(a_14_), .A2(n2793), .ZN(n2792) );
  NAND2_X1 U2786 ( .A1(b_9_), .A2(n2794), .ZN(n2789) );
  NAND2_X1 U2787 ( .A1(n2077), .A2(n2795), .ZN(n2794) );
  NAND2_X1 U2788 ( .A1(a_15_), .A2(n2674), .ZN(n2795) );
  NAND3_X1 U2789 ( .A1(b_10_), .A2(n2417), .A3(b_11_), .ZN(n2663) );
  XNOR2_X1 U2790 ( .A(n2796), .B(n2797), .ZN(n2653) );
  XOR2_X1 U2791 ( .A(n2798), .B(n2799), .Z(n2796) );
  XOR2_X1 U2792 ( .A(n2800), .B(n2801), .Z(n2685) );
  XOR2_X1 U2793 ( .A(n2802), .B(n2803), .Z(n2801) );
  NAND2_X1 U2794 ( .A1(b_10_), .A2(a_8_), .ZN(n2803) );
  XOR2_X1 U2795 ( .A(n2804), .B(n2805), .Z(n2614) );
  XOR2_X1 U2796 ( .A(n2806), .B(n2807), .Z(n2805) );
  NAND2_X1 U2797 ( .A1(b_10_), .A2(a_7_), .ZN(n2807) );
  XNOR2_X1 U2798 ( .A(n2808), .B(n2809), .ZN(n2602) );
  NAND2_X1 U2799 ( .A1(n2810), .A2(n2811), .ZN(n2808) );
  XNOR2_X1 U2800 ( .A(n2812), .B(n2813), .ZN(n2696) );
  XNOR2_X1 U2801 ( .A(n2814), .B(n2815), .ZN(n2812) );
  XOR2_X1 U2802 ( .A(n2816), .B(n2817), .Z(n2700) );
  XNOR2_X1 U2803 ( .A(n2818), .B(n2819), .ZN(n2817) );
  NAND2_X1 U2804 ( .A1(b_10_), .A2(a_2_), .ZN(n2819) );
  XNOR2_X1 U2805 ( .A(n2820), .B(n2821), .ZN(n2705) );
  NAND2_X1 U2806 ( .A1(n2822), .A2(n2823), .ZN(n2820) );
  XOR2_X1 U2807 ( .A(n2824), .B(n2825), .Z(n2586) );
  NAND2_X1 U2808 ( .A1(n2826), .A2(n2827), .ZN(n2824) );
  NAND3_X1 U2809 ( .A1(n2042), .A2(n2043), .A3(n2200), .ZN(n2038) );
  INV_X1 U2810 ( .A(n2041), .ZN(n2200) );
  NAND2_X1 U2811 ( .A1(n2828), .A2(n2198), .ZN(n2041) );
  NAND2_X1 U2812 ( .A1(n2829), .A2(n2830), .ZN(n2828) );
  XOR2_X1 U2813 ( .A(n2831), .B(n2832), .Z(n2830) );
  NAND2_X1 U2814 ( .A1(n2826), .A2(n2833), .ZN(n2043) );
  NAND2_X1 U2815 ( .A1(n2825), .A2(n2827), .ZN(n2833) );
  NAND2_X1 U2816 ( .A1(n2834), .A2(n2835), .ZN(n2827) );
  NAND2_X1 U2817 ( .A1(b_10_), .A2(a_0_), .ZN(n2835) );
  INV_X1 U2818 ( .A(n2836), .ZN(n2834) );
  XOR2_X1 U2819 ( .A(n2837), .B(n2838), .Z(n2825) );
  XOR2_X1 U2820 ( .A(n2839), .B(n2840), .Z(n2837) );
  NOR2_X1 U2821 ( .A1(n2793), .A2(n2343), .ZN(n2840) );
  NAND2_X1 U2822 ( .A1(a_0_), .A2(n2836), .ZN(n2826) );
  NAND2_X1 U2823 ( .A1(n2822), .A2(n2841), .ZN(n2836) );
  NAND2_X1 U2824 ( .A1(n2821), .A2(n2823), .ZN(n2841) );
  NAND2_X1 U2825 ( .A1(n2842), .A2(n2843), .ZN(n2823) );
  NAND2_X1 U2826 ( .A1(b_10_), .A2(a_1_), .ZN(n2843) );
  XOR2_X1 U2827 ( .A(n2844), .B(n2845), .Z(n2821) );
  XNOR2_X1 U2828 ( .A(n2846), .B(n2847), .ZN(n2845) );
  NAND2_X1 U2829 ( .A1(a_2_), .A2(b_9_), .ZN(n2847) );
  INV_X1 U2830 ( .A(n2848), .ZN(n2822) );
  NOR2_X1 U2831 ( .A1(n2343), .A2(n2842), .ZN(n2848) );
  NOR2_X1 U2832 ( .A1(n2849), .A2(n2850), .ZN(n2842) );
  INV_X1 U2833 ( .A(n2851), .ZN(n2850) );
  NAND3_X1 U2834 ( .A1(a_2_), .A2(n2852), .A3(b_10_), .ZN(n2851) );
  NAND2_X1 U2835 ( .A1(n2818), .A2(n2816), .ZN(n2852) );
  NOR2_X1 U2836 ( .A1(n2816), .A2(n2818), .ZN(n2849) );
  NOR2_X1 U2837 ( .A1(n2853), .A2(n2854), .ZN(n2818) );
  INV_X1 U2838 ( .A(n2855), .ZN(n2854) );
  NAND2_X1 U2839 ( .A1(n2815), .A2(n2856), .ZN(n2855) );
  NAND2_X1 U2840 ( .A1(n2814), .A2(n2813), .ZN(n2856) );
  NOR2_X1 U2841 ( .A1(n2674), .A2(n2322), .ZN(n2815) );
  NOR2_X1 U2842 ( .A1(n2813), .A2(n2814), .ZN(n2853) );
  NOR2_X1 U2843 ( .A1(n2857), .A2(n2858), .ZN(n2814) );
  NOR3_X1 U2844 ( .A1(n2230), .A2(n2859), .A3(n2674), .ZN(n2858) );
  NOR2_X1 U2845 ( .A1(n2725), .A2(n2724), .ZN(n2859) );
  INV_X1 U2846 ( .A(n2860), .ZN(n2857) );
  NAND2_X1 U2847 ( .A1(n2724), .A2(n2725), .ZN(n2860) );
  NAND2_X1 U2848 ( .A1(n2810), .A2(n2861), .ZN(n2725) );
  NAND2_X1 U2849 ( .A1(n2809), .A2(n2811), .ZN(n2861) );
  NAND2_X1 U2850 ( .A1(n2862), .A2(n2863), .ZN(n2811) );
  NAND2_X1 U2851 ( .A1(b_10_), .A2(a_5_), .ZN(n2863) );
  XOR2_X1 U2852 ( .A(n2864), .B(n2865), .Z(n2809) );
  XOR2_X1 U2853 ( .A(n2866), .B(n2867), .Z(n2864) );
  NOR2_X1 U2854 ( .A1(n2793), .A2(n2247), .ZN(n2867) );
  NAND2_X1 U2855 ( .A1(a_5_), .A2(n2868), .ZN(n2810) );
  INV_X1 U2856 ( .A(n2862), .ZN(n2868) );
  NOR2_X1 U2857 ( .A1(n2869), .A2(n2870), .ZN(n2862) );
  INV_X1 U2858 ( .A(n2871), .ZN(n2870) );
  NAND3_X1 U2859 ( .A1(a_6_), .A2(n2872), .A3(b_10_), .ZN(n2871) );
  NAND2_X1 U2860 ( .A1(n2738), .A2(n2737), .ZN(n2872) );
  NOR2_X1 U2861 ( .A1(n2737), .A2(n2738), .ZN(n2869) );
  NOR2_X1 U2862 ( .A1(n2873), .A2(n2874), .ZN(n2738) );
  NOR3_X1 U2863 ( .A1(n2626), .A2(n2875), .A3(n2674), .ZN(n2874) );
  NOR2_X1 U2864 ( .A1(n2806), .A2(n2804), .ZN(n2875) );
  INV_X1 U2865 ( .A(n2876), .ZN(n2873) );
  NAND2_X1 U2866 ( .A1(n2804), .A2(n2806), .ZN(n2876) );
  NAND2_X1 U2867 ( .A1(n2877), .A2(n2878), .ZN(n2806) );
  NAND3_X1 U2868 ( .A1(a_8_), .A2(n2879), .A3(b_10_), .ZN(n2878) );
  INV_X1 U2869 ( .A(n2880), .ZN(n2879) );
  NOR2_X1 U2870 ( .A1(n2802), .A2(n2800), .ZN(n2880) );
  NAND2_X1 U2871 ( .A1(n2800), .A2(n2802), .ZN(n2877) );
  NAND2_X1 U2872 ( .A1(n2754), .A2(n2881), .ZN(n2802) );
  NAND2_X1 U2873 ( .A1(n2753), .A2(n2755), .ZN(n2881) );
  NAND2_X1 U2874 ( .A1(n2882), .A2(n2883), .ZN(n2755) );
  NAND2_X1 U2875 ( .A1(b_10_), .A2(a_9_), .ZN(n2882) );
  XNOR2_X1 U2876 ( .A(n2884), .B(n2885), .ZN(n2753) );
  NAND2_X1 U2877 ( .A1(n2886), .A2(n2887), .ZN(n2884) );
  INV_X1 U2878 ( .A(n2888), .ZN(n2754) );
  NOR2_X1 U2879 ( .A1(n2883), .A2(n2275), .ZN(n2888) );
  NAND2_X1 U2880 ( .A1(n2889), .A2(n2890), .ZN(n2883) );
  NAND2_X1 U2881 ( .A1(n2891), .A2(n2761), .ZN(n2890) );
  NAND2_X1 U2882 ( .A1(n2759), .A2(n2762), .ZN(n2891) );
  INV_X1 U2883 ( .A(n2892), .ZN(n2889) );
  NOR2_X1 U2884 ( .A1(n2762), .A2(n2759), .ZN(n2892) );
  XNOR2_X1 U2885 ( .A(n2893), .B(n2894), .ZN(n2759) );
  XOR2_X1 U2886 ( .A(n2895), .B(n2896), .Z(n2893) );
  NAND2_X1 U2887 ( .A1(a_11_), .A2(b_9_), .ZN(n2895) );
  NAND2_X1 U2888 ( .A1(n2897), .A2(n2898), .ZN(n2762) );
  NAND3_X1 U2889 ( .A1(a_11_), .A2(n2899), .A3(b_10_), .ZN(n2898) );
  NAND2_X1 U2890 ( .A1(n2770), .A2(n2768), .ZN(n2899) );
  INV_X1 U2891 ( .A(n2900), .ZN(n2897) );
  NOR2_X1 U2892 ( .A1(n2768), .A2(n2770), .ZN(n2900) );
  NOR2_X1 U2893 ( .A1(n2901), .A2(n2902), .ZN(n2770) );
  INV_X1 U2894 ( .A(n2903), .ZN(n2902) );
  NAND2_X1 U2895 ( .A1(n2778), .A2(n2904), .ZN(n2903) );
  NAND2_X1 U2896 ( .A1(n2779), .A2(n2777), .ZN(n2904) );
  NOR2_X1 U2897 ( .A1(n2674), .A2(n2094), .ZN(n2778) );
  NOR2_X1 U2898 ( .A1(n2777), .A2(n2779), .ZN(n2901) );
  NOR2_X1 U2899 ( .A1(n2905), .A2(n2906), .ZN(n2779) );
  INV_X1 U2900 ( .A(n2907), .ZN(n2906) );
  NAND2_X1 U2901 ( .A1(n2797), .A2(n2908), .ZN(n2907) );
  NAND2_X1 U2902 ( .A1(n2798), .A2(n2799), .ZN(n2908) );
  NOR2_X1 U2903 ( .A1(n2674), .A2(n2408), .ZN(n2797) );
  NOR2_X1 U2904 ( .A1(n2799), .A2(n2798), .ZN(n2905) );
  INV_X1 U2905 ( .A(n2909), .ZN(n2798) );
  NAND2_X1 U2906 ( .A1(n2910), .A2(n2911), .ZN(n2909) );
  NAND2_X1 U2907 ( .A1(b_8_), .A2(n2912), .ZN(n2911) );
  NAND2_X1 U2908 ( .A1(n2077), .A2(n2913), .ZN(n2912) );
  NAND2_X1 U2909 ( .A1(a_15_), .A2(n2793), .ZN(n2913) );
  NAND2_X1 U2910 ( .A1(b_9_), .A2(n2914), .ZN(n2910) );
  NAND2_X1 U2911 ( .A1(n2081), .A2(n2915), .ZN(n2914) );
  NAND2_X1 U2912 ( .A1(a_14_), .A2(n2916), .ZN(n2915) );
  NAND3_X1 U2913 ( .A1(n2417), .A2(b_9_), .A3(b_10_), .ZN(n2799) );
  XNOR2_X1 U2914 ( .A(n2917), .B(n2918), .ZN(n2777) );
  XOR2_X1 U2915 ( .A(n2919), .B(n2920), .Z(n2917) );
  XOR2_X1 U2916 ( .A(n2921), .B(n2922), .Z(n2768) );
  XNOR2_X1 U2917 ( .A(n2923), .B(n2924), .ZN(n2921) );
  XOR2_X1 U2918 ( .A(n2925), .B(n2926), .Z(n2800) );
  XOR2_X1 U2919 ( .A(n2927), .B(n2928), .Z(n2926) );
  XNOR2_X1 U2920 ( .A(n2929), .B(n2930), .ZN(n2804) );
  XNOR2_X1 U2921 ( .A(n2931), .B(n2932), .ZN(n2930) );
  XNOR2_X1 U2922 ( .A(n2933), .B(n2934), .ZN(n2737) );
  XOR2_X1 U2923 ( .A(n2935), .B(n2936), .Z(n2933) );
  NOR2_X1 U2924 ( .A1(n2793), .A2(n2626), .ZN(n2936) );
  XNOR2_X1 U2925 ( .A(n2937), .B(n2938), .ZN(n2724) );
  NAND2_X1 U2926 ( .A1(n2939), .A2(n2940), .ZN(n2937) );
  XOR2_X1 U2927 ( .A(n2941), .B(n2942), .Z(n2813) );
  XOR2_X1 U2928 ( .A(n2943), .B(n2944), .Z(n2941) );
  XOR2_X1 U2929 ( .A(n2945), .B(n2946), .Z(n2816) );
  XOR2_X1 U2930 ( .A(n2947), .B(n2948), .Z(n2946) );
  NAND2_X1 U2931 ( .A1(a_3_), .A2(b_9_), .ZN(n2948) );
  XOR2_X1 U2932 ( .A(n2949), .B(n2950), .Z(n2042) );
  XNOR2_X1 U2933 ( .A(n2951), .B(n2952), .ZN(n2950) );
  NAND2_X1 U2934 ( .A1(a_0_), .A2(b_9_), .ZN(n2952) );
  NAND2_X1 U2935 ( .A1(n2953), .A2(n2954), .ZN(n2198) );
  INV_X1 U2936 ( .A(n2829), .ZN(n2954) );
  NOR2_X1 U2937 ( .A1(n2955), .A2(n2956), .ZN(n2829) );
  INV_X1 U2938 ( .A(n2957), .ZN(n2956) );
  NAND3_X1 U2939 ( .A1(b_9_), .A2(n2958), .A3(a_0_), .ZN(n2957) );
  NAND2_X1 U2940 ( .A1(n2951), .A2(n2949), .ZN(n2958) );
  NOR2_X1 U2941 ( .A1(n2949), .A2(n2951), .ZN(n2955) );
  NOR2_X1 U2942 ( .A1(n2959), .A2(n2960), .ZN(n2951) );
  NOR3_X1 U2943 ( .A1(n2793), .A2(n2961), .A3(n2343), .ZN(n2960) );
  NOR2_X1 U2944 ( .A1(n2839), .A2(n2838), .ZN(n2961) );
  INV_X1 U2945 ( .A(n2962), .ZN(n2959) );
  NAND2_X1 U2946 ( .A1(n2838), .A2(n2839), .ZN(n2962) );
  NAND2_X1 U2947 ( .A1(n2963), .A2(n2964), .ZN(n2839) );
  NAND3_X1 U2948 ( .A1(b_9_), .A2(n2965), .A3(a_2_), .ZN(n2964) );
  NAND2_X1 U2949 ( .A1(n2846), .A2(n2844), .ZN(n2965) );
  INV_X1 U2950 ( .A(n2966), .ZN(n2963) );
  NOR2_X1 U2951 ( .A1(n2844), .A2(n2846), .ZN(n2966) );
  NOR2_X1 U2952 ( .A1(n2967), .A2(n2968), .ZN(n2846) );
  NOR3_X1 U2953 ( .A1(n2793), .A2(n2969), .A3(n2322), .ZN(n2968) );
  INV_X1 U2954 ( .A(n2970), .ZN(n2969) );
  NAND2_X1 U2955 ( .A1(n2945), .A2(n2947), .ZN(n2970) );
  NOR2_X1 U2956 ( .A1(n2947), .A2(n2945), .ZN(n2967) );
  XOR2_X1 U2957 ( .A(n2971), .B(n2972), .Z(n2945) );
  XOR2_X1 U2958 ( .A(n2973), .B(n2974), .Z(n2972) );
  NAND2_X1 U2959 ( .A1(a_4_), .A2(b_8_), .ZN(n2974) );
  NAND2_X1 U2960 ( .A1(n2975), .A2(n2976), .ZN(n2947) );
  NAND2_X1 U2961 ( .A1(n2942), .A2(n2977), .ZN(n2976) );
  NAND2_X1 U2962 ( .A1(n2978), .A2(n2979), .ZN(n2977) );
  INV_X1 U2963 ( .A(n2943), .ZN(n2978) );
  XNOR2_X1 U2964 ( .A(n2980), .B(n2981), .ZN(n2942) );
  XOR2_X1 U2965 ( .A(n2982), .B(n2983), .Z(n2981) );
  NAND2_X1 U2966 ( .A1(n2944), .A2(n2943), .ZN(n2975) );
  NAND2_X1 U2967 ( .A1(a_4_), .A2(b_9_), .ZN(n2943) );
  INV_X1 U2968 ( .A(n2979), .ZN(n2944) );
  NAND2_X1 U2969 ( .A1(n2939), .A2(n2984), .ZN(n2979) );
  NAND2_X1 U2970 ( .A1(n2938), .A2(n2940), .ZN(n2984) );
  NAND2_X1 U2971 ( .A1(n2985), .A2(n2986), .ZN(n2940) );
  NAND2_X1 U2972 ( .A1(a_5_), .A2(b_9_), .ZN(n2986) );
  XNOR2_X1 U2973 ( .A(n2987), .B(n2988), .ZN(n2938) );
  XNOR2_X1 U2974 ( .A(n2989), .B(n2990), .ZN(n2987) );
  NOR2_X1 U2975 ( .A1(n2916), .A2(n2247), .ZN(n2990) );
  NAND2_X1 U2976 ( .A1(a_5_), .A2(n2991), .ZN(n2939) );
  INV_X1 U2977 ( .A(n2985), .ZN(n2991) );
  NOR2_X1 U2978 ( .A1(n2992), .A2(n2993), .ZN(n2985) );
  NOR3_X1 U2979 ( .A1(n2793), .A2(n2994), .A3(n2247), .ZN(n2993) );
  NOR2_X1 U2980 ( .A1(n2866), .A2(n2865), .ZN(n2994) );
  INV_X1 U2981 ( .A(n2995), .ZN(n2992) );
  NAND2_X1 U2982 ( .A1(n2865), .A2(n2866), .ZN(n2995) );
  NAND2_X1 U2983 ( .A1(n2996), .A2(n2997), .ZN(n2866) );
  INV_X1 U2984 ( .A(n2998), .ZN(n2997) );
  NOR3_X1 U2985 ( .A1(n2793), .A2(n2999), .A3(n2626), .ZN(n2998) );
  NOR2_X1 U2986 ( .A1(n2935), .A2(n2934), .ZN(n2999) );
  NAND2_X1 U2987 ( .A1(n2934), .A2(n2935), .ZN(n2996) );
  NAND2_X1 U2988 ( .A1(n3000), .A2(n3001), .ZN(n2935) );
  NAND2_X1 U2989 ( .A1(n2932), .A2(n3002), .ZN(n3001) );
  NAND2_X1 U2990 ( .A1(n2929), .A2(n2931), .ZN(n3002) );
  NOR2_X1 U2991 ( .A1(n2793), .A2(n2377), .ZN(n2932) );
  INV_X1 U2992 ( .A(n3003), .ZN(n3000) );
  NOR2_X1 U2993 ( .A1(n2931), .A2(n2929), .ZN(n3003) );
  XOR2_X1 U2994 ( .A(n3004), .B(n3005), .Z(n2929) );
  NAND2_X1 U2995 ( .A1(n3006), .A2(n3007), .ZN(n3004) );
  NAND2_X1 U2996 ( .A1(n3008), .A2(n3009), .ZN(n2931) );
  NAND2_X1 U2997 ( .A1(n2925), .A2(n3010), .ZN(n3009) );
  NAND2_X1 U2998 ( .A1(n2928), .A2(n3011), .ZN(n3010) );
  XOR2_X1 U2999 ( .A(n3012), .B(n3013), .Z(n2925) );
  NAND2_X1 U3000 ( .A1(n3014), .A2(n3015), .ZN(n3012) );
  NAND2_X1 U3001 ( .A1(n2927), .A2(n3016), .ZN(n3008) );
  INV_X1 U3002 ( .A(n3011), .ZN(n2927) );
  NAND2_X1 U3003 ( .A1(n2886), .A2(n3017), .ZN(n3011) );
  NAND2_X1 U3004 ( .A1(n2885), .A2(n2887), .ZN(n3017) );
  NAND2_X1 U3005 ( .A1(n3018), .A2(n3019), .ZN(n2887) );
  NAND2_X1 U3006 ( .A1(a_10_), .A2(b_9_), .ZN(n3019) );
  XNOR2_X1 U3007 ( .A(n3020), .B(n3021), .ZN(n2885) );
  XOR2_X1 U3008 ( .A(n3022), .B(n3023), .Z(n3020) );
  NAND2_X1 U3009 ( .A1(a_11_), .A2(b_8_), .ZN(n3022) );
  INV_X1 U3010 ( .A(n3024), .ZN(n2886) );
  NOR2_X1 U3011 ( .A1(n2523), .A2(n3018), .ZN(n3024) );
  NOR2_X1 U3012 ( .A1(n3025), .A2(n3026), .ZN(n3018) );
  INV_X1 U3013 ( .A(n3027), .ZN(n3026) );
  NAND3_X1 U3014 ( .A1(b_9_), .A2(n3028), .A3(a_11_), .ZN(n3027) );
  NAND2_X1 U3015 ( .A1(n2896), .A2(n2894), .ZN(n3028) );
  NOR2_X1 U3016 ( .A1(n2894), .A2(n2896), .ZN(n3025) );
  NOR2_X1 U3017 ( .A1(n3029), .A2(n3030), .ZN(n2896) );
  INV_X1 U3018 ( .A(n3031), .ZN(n3030) );
  NAND2_X1 U3019 ( .A1(n2923), .A2(n3032), .ZN(n3031) );
  NAND2_X1 U3020 ( .A1(n2924), .A2(n2922), .ZN(n3032) );
  NOR2_X1 U3021 ( .A1(n2094), .A2(n2793), .ZN(n2923) );
  NOR2_X1 U3022 ( .A1(n2922), .A2(n2924), .ZN(n3029) );
  NOR2_X1 U3023 ( .A1(n3033), .A2(n3034), .ZN(n2924) );
  INV_X1 U3024 ( .A(n3035), .ZN(n3034) );
  NAND2_X1 U3025 ( .A1(n2918), .A2(n3036), .ZN(n3035) );
  NAND2_X1 U3026 ( .A1(n2919), .A2(n2920), .ZN(n3036) );
  NOR2_X1 U3027 ( .A1(n2408), .A2(n2793), .ZN(n2918) );
  NOR2_X1 U3028 ( .A1(n2920), .A2(n2919), .ZN(n3033) );
  INV_X1 U3029 ( .A(n3037), .ZN(n2919) );
  NAND2_X1 U3030 ( .A1(n3038), .A2(n3039), .ZN(n3037) );
  NAND2_X1 U3031 ( .A1(b_7_), .A2(n3040), .ZN(n3039) );
  NAND2_X1 U3032 ( .A1(n2077), .A2(n3041), .ZN(n3040) );
  NAND2_X1 U3033 ( .A1(a_15_), .A2(n2916), .ZN(n3041) );
  NAND2_X1 U3034 ( .A1(b_8_), .A2(n3042), .ZN(n3038) );
  NAND2_X1 U3035 ( .A1(n2081), .A2(n3043), .ZN(n3042) );
  NAND2_X1 U3036 ( .A1(a_14_), .A2(n3044), .ZN(n3043) );
  NAND3_X1 U3037 ( .A1(n2417), .A2(b_9_), .A3(b_8_), .ZN(n2920) );
  XNOR2_X1 U3038 ( .A(n3045), .B(n3046), .ZN(n2922) );
  XOR2_X1 U3039 ( .A(n3047), .B(n3048), .Z(n3045) );
  XOR2_X1 U3040 ( .A(n3049), .B(n3050), .Z(n2894) );
  XNOR2_X1 U3041 ( .A(n3051), .B(n3052), .ZN(n3049) );
  XNOR2_X1 U3042 ( .A(n3053), .B(n3054), .ZN(n2934) );
  XOR2_X1 U3043 ( .A(n3055), .B(n3056), .Z(n3054) );
  XNOR2_X1 U3044 ( .A(n3057), .B(n3058), .ZN(n2865) );
  XNOR2_X1 U3045 ( .A(n3059), .B(n3060), .ZN(n3057) );
  NOR2_X1 U3046 ( .A1(n2916), .A2(n2626), .ZN(n3060) );
  XOR2_X1 U3047 ( .A(n3061), .B(n3062), .Z(n2844) );
  NAND2_X1 U3048 ( .A1(n3063), .A2(n3064), .ZN(n3061) );
  XNOR2_X1 U3049 ( .A(n3065), .B(n3066), .ZN(n2838) );
  NAND2_X1 U3050 ( .A1(n3067), .A2(n3068), .ZN(n3065) );
  XOR2_X1 U3051 ( .A(n3069), .B(n3070), .Z(n2949) );
  NAND2_X1 U3052 ( .A1(n3071), .A2(n3072), .ZN(n3069) );
  XNOR2_X1 U3053 ( .A(n2831), .B(n2832), .ZN(n2953) );
  NAND2_X1 U3054 ( .A1(n3073), .A2(n3074), .ZN(n2831) );
  XOR2_X1 U3055 ( .A(n2053), .B(n2052), .Z(n2045) );
  NAND3_X1 U3056 ( .A1(n2052), .A2(n2053), .A3(n2197), .ZN(n2048) );
  INV_X1 U3057 ( .A(n2051), .ZN(n2197) );
  NAND2_X1 U3058 ( .A1(n3075), .A2(n2195), .ZN(n2051) );
  NAND2_X1 U3059 ( .A1(n3076), .A2(n3077), .ZN(n3075) );
  XOR2_X1 U3060 ( .A(n3078), .B(n3079), .Z(n3076) );
  NAND2_X1 U3061 ( .A1(n3073), .A2(n3080), .ZN(n2053) );
  NAND2_X1 U3062 ( .A1(n2832), .A2(n3074), .ZN(n3080) );
  NAND2_X1 U3063 ( .A1(n3081), .A2(n3082), .ZN(n3074) );
  NAND2_X1 U3064 ( .A1(a_0_), .A2(b_8_), .ZN(n3082) );
  INV_X1 U3065 ( .A(n3083), .ZN(n3081) );
  XNOR2_X1 U3066 ( .A(n3084), .B(n3085), .ZN(n2832) );
  XNOR2_X1 U3067 ( .A(n3086), .B(n3087), .ZN(n3084) );
  NOR2_X1 U3068 ( .A1(n3044), .A2(n2343), .ZN(n3087) );
  NAND2_X1 U3069 ( .A1(a_0_), .A2(n3083), .ZN(n3073) );
  NAND2_X1 U3070 ( .A1(n3071), .A2(n3088), .ZN(n3083) );
  NAND2_X1 U3071 ( .A1(n3070), .A2(n3072), .ZN(n3088) );
  NAND2_X1 U3072 ( .A1(n3089), .A2(n3090), .ZN(n3072) );
  NAND2_X1 U3073 ( .A1(a_1_), .A2(b_8_), .ZN(n3090) );
  INV_X1 U3074 ( .A(n3091), .ZN(n3089) );
  XOR2_X1 U3075 ( .A(n3092), .B(n3093), .Z(n3070) );
  XNOR2_X1 U3076 ( .A(n3094), .B(n3095), .ZN(n3093) );
  NAND2_X1 U3077 ( .A1(a_2_), .A2(b_7_), .ZN(n3095) );
  NAND2_X1 U3078 ( .A1(a_1_), .A2(n3091), .ZN(n3071) );
  NAND2_X1 U3079 ( .A1(n3067), .A2(n3096), .ZN(n3091) );
  NAND2_X1 U3080 ( .A1(n3066), .A2(n3068), .ZN(n3096) );
  NAND2_X1 U3081 ( .A1(n3097), .A2(n3098), .ZN(n3068) );
  NAND2_X1 U3082 ( .A1(a_2_), .A2(b_8_), .ZN(n3098) );
  INV_X1 U3083 ( .A(n3099), .ZN(n3097) );
  XOR2_X1 U3084 ( .A(n3100), .B(n3101), .Z(n3066) );
  XNOR2_X1 U3085 ( .A(n3102), .B(n3103), .ZN(n3101) );
  NAND2_X1 U3086 ( .A1(a_3_), .A2(b_7_), .ZN(n3103) );
  NAND2_X1 U3087 ( .A1(a_2_), .A2(n3099), .ZN(n3067) );
  NAND2_X1 U3088 ( .A1(n3063), .A2(n3104), .ZN(n3099) );
  NAND2_X1 U3089 ( .A1(n3062), .A2(n3064), .ZN(n3104) );
  NAND2_X1 U3090 ( .A1(n3105), .A2(n3106), .ZN(n3064) );
  NAND2_X1 U3091 ( .A1(a_3_), .A2(b_8_), .ZN(n3106) );
  XOR2_X1 U3092 ( .A(n3107), .B(n3108), .Z(n3062) );
  XNOR2_X1 U3093 ( .A(n3109), .B(n3110), .ZN(n3108) );
  NAND2_X1 U3094 ( .A1(a_4_), .A2(b_7_), .ZN(n3110) );
  NAND2_X1 U3095 ( .A1(a_3_), .A2(n3111), .ZN(n3063) );
  INV_X1 U3096 ( .A(n3105), .ZN(n3111) );
  NOR2_X1 U3097 ( .A1(n3112), .A2(n3113), .ZN(n3105) );
  NOR3_X1 U3098 ( .A1(n2916), .A2(n3114), .A3(n2230), .ZN(n3113) );
  NOR2_X1 U3099 ( .A1(n2971), .A2(n2973), .ZN(n3114) );
  INV_X1 U3100 ( .A(n3115), .ZN(n3112) );
  NAND2_X1 U3101 ( .A1(n2971), .A2(n2973), .ZN(n3115) );
  NAND2_X1 U3102 ( .A1(n3116), .A2(n3117), .ZN(n2973) );
  NAND2_X1 U3103 ( .A1(n2983), .A2(n3118), .ZN(n3117) );
  NAND2_X1 U3104 ( .A1(n2980), .A2(n2982), .ZN(n3118) );
  NOR2_X1 U3105 ( .A1(n2366), .A2(n2916), .ZN(n2983) );
  INV_X1 U3106 ( .A(n3119), .ZN(n3116) );
  NOR2_X1 U3107 ( .A1(n2980), .A2(n2982), .ZN(n3119) );
  NOR2_X1 U3108 ( .A1(n3120), .A2(n3121), .ZN(n2982) );
  NOR3_X1 U3109 ( .A1(n2916), .A2(n3122), .A3(n2247), .ZN(n3121) );
  INV_X1 U3110 ( .A(n3123), .ZN(n3122) );
  NAND2_X1 U3111 ( .A1(n2989), .A2(n2988), .ZN(n3123) );
  NOR2_X1 U3112 ( .A1(n2988), .A2(n2989), .ZN(n3120) );
  NOR2_X1 U3113 ( .A1(n3124), .A2(n3125), .ZN(n2989) );
  NOR3_X1 U3114 ( .A1(n2916), .A2(n3126), .A3(n2626), .ZN(n3125) );
  NOR2_X1 U3115 ( .A1(n3058), .A2(n3059), .ZN(n3126) );
  INV_X1 U3116 ( .A(n3127), .ZN(n3124) );
  NAND2_X1 U3117 ( .A1(n3059), .A2(n3058), .ZN(n3127) );
  XNOR2_X1 U3118 ( .A(n3128), .B(n3129), .ZN(n3058) );
  XOR2_X1 U3119 ( .A(n3130), .B(n3131), .Z(n3129) );
  NOR2_X1 U3120 ( .A1(n3132), .A2(n3133), .ZN(n3059) );
  NOR2_X1 U3121 ( .A1(n3134), .A2(n3135), .ZN(n3133) );
  INV_X1 U3122 ( .A(n3055), .ZN(n3135) );
  INV_X1 U3123 ( .A(n3136), .ZN(n3134) );
  NAND2_X1 U3124 ( .A1(n3053), .A2(n3056), .ZN(n3136) );
  NOR2_X1 U3125 ( .A1(n3056), .A2(n3053), .ZN(n3132) );
  XNOR2_X1 U3126 ( .A(n3137), .B(n3138), .ZN(n3053) );
  NAND2_X1 U3127 ( .A1(n3139), .A2(n3140), .ZN(n3137) );
  NAND2_X1 U3128 ( .A1(n3006), .A2(n3141), .ZN(n3056) );
  NAND2_X1 U3129 ( .A1(n3005), .A2(n3007), .ZN(n3141) );
  NAND2_X1 U3130 ( .A1(n3142), .A2(n3143), .ZN(n3007) );
  NAND2_X1 U3131 ( .A1(a_9_), .A2(b_8_), .ZN(n3143) );
  INV_X1 U3132 ( .A(n3144), .ZN(n3142) );
  XNOR2_X1 U3133 ( .A(n3145), .B(n3146), .ZN(n3005) );
  NAND2_X1 U3134 ( .A1(n3147), .A2(n3148), .ZN(n3145) );
  NAND2_X1 U3135 ( .A1(a_9_), .A2(n3144), .ZN(n3006) );
  NAND2_X1 U3136 ( .A1(n3014), .A2(n3149), .ZN(n3144) );
  NAND2_X1 U3137 ( .A1(n3013), .A2(n3015), .ZN(n3149) );
  NAND2_X1 U3138 ( .A1(n3150), .A2(n3151), .ZN(n3015) );
  NAND2_X1 U3139 ( .A1(a_10_), .A2(b_8_), .ZN(n3151) );
  XNOR2_X1 U3140 ( .A(n3152), .B(n3153), .ZN(n3013) );
  XOR2_X1 U3141 ( .A(n3154), .B(n3155), .Z(n3152) );
  NAND2_X1 U3142 ( .A1(a_11_), .A2(b_7_), .ZN(n3154) );
  INV_X1 U3143 ( .A(n3156), .ZN(n3014) );
  NOR2_X1 U3144 ( .A1(n2523), .A2(n3150), .ZN(n3156) );
  NOR2_X1 U3145 ( .A1(n3157), .A2(n3158), .ZN(n3150) );
  INV_X1 U3146 ( .A(n3159), .ZN(n3158) );
  NAND3_X1 U3147 ( .A1(b_8_), .A2(n3160), .A3(a_11_), .ZN(n3159) );
  NAND2_X1 U3148 ( .A1(n3021), .A2(n3023), .ZN(n3160) );
  NOR2_X1 U3149 ( .A1(n3021), .A2(n3023), .ZN(n3157) );
  NOR2_X1 U3150 ( .A1(n3161), .A2(n3162), .ZN(n3023) );
  INV_X1 U3151 ( .A(n3163), .ZN(n3162) );
  NAND2_X1 U3152 ( .A1(n3051), .A2(n3164), .ZN(n3163) );
  NAND2_X1 U3153 ( .A1(n3052), .A2(n3050), .ZN(n3164) );
  NOR2_X1 U3154 ( .A1(n2916), .A2(n2094), .ZN(n3051) );
  NOR2_X1 U3155 ( .A1(n3050), .A2(n3052), .ZN(n3161) );
  NOR2_X1 U3156 ( .A1(n3165), .A2(n3166), .ZN(n3052) );
  INV_X1 U3157 ( .A(n3167), .ZN(n3166) );
  NAND2_X1 U3158 ( .A1(n3046), .A2(n3168), .ZN(n3167) );
  NAND2_X1 U3159 ( .A1(n3047), .A2(n3048), .ZN(n3168) );
  NOR2_X1 U3160 ( .A1(n2916), .A2(n2408), .ZN(n3046) );
  NOR2_X1 U3161 ( .A1(n3048), .A2(n3047), .ZN(n3165) );
  INV_X1 U3162 ( .A(n3169), .ZN(n3047) );
  NAND2_X1 U3163 ( .A1(n3170), .A2(n3171), .ZN(n3169) );
  NAND2_X1 U3164 ( .A1(b_6_), .A2(n3172), .ZN(n3171) );
  NAND2_X1 U3165 ( .A1(n2077), .A2(n3173), .ZN(n3172) );
  NAND2_X1 U3166 ( .A1(a_15_), .A2(n3044), .ZN(n3173) );
  NAND2_X1 U3167 ( .A1(b_7_), .A2(n3174), .ZN(n3170) );
  NAND2_X1 U3168 ( .A1(n2081), .A2(n3175), .ZN(n3174) );
  NAND2_X1 U3169 ( .A1(a_14_), .A2(n3176), .ZN(n3175) );
  NAND3_X1 U3170 ( .A1(b_8_), .A2(n2417), .A3(b_7_), .ZN(n3048) );
  XNOR2_X1 U3171 ( .A(n3177), .B(n3178), .ZN(n3050) );
  XOR2_X1 U3172 ( .A(n3179), .B(n3180), .Z(n3177) );
  XOR2_X1 U3173 ( .A(n3181), .B(n3182), .Z(n3021) );
  XNOR2_X1 U3174 ( .A(n3183), .B(n3184), .ZN(n3181) );
  XOR2_X1 U3175 ( .A(n3185), .B(n3186), .Z(n2988) );
  XOR2_X1 U3176 ( .A(n3187), .B(n3188), .Z(n3185) );
  XNOR2_X1 U3177 ( .A(n3189), .B(n3190), .ZN(n2980) );
  NOR2_X1 U3178 ( .A1(n3191), .A2(n3192), .ZN(n3190) );
  NOR2_X1 U3179 ( .A1(n3193), .A2(n3194), .ZN(n3191) );
  NOR2_X1 U3180 ( .A1(n3044), .A2(n2247), .ZN(n3194) );
  INV_X1 U3181 ( .A(n3195), .ZN(n3193) );
  XOR2_X1 U3182 ( .A(n3196), .B(n3197), .Z(n2971) );
  XNOR2_X1 U3183 ( .A(n3198), .B(n3199), .ZN(n3197) );
  NAND2_X1 U3184 ( .A1(a_5_), .A2(b_7_), .ZN(n3199) );
  XOR2_X1 U3185 ( .A(n3200), .B(n3201), .Z(n2052) );
  XNOR2_X1 U3186 ( .A(n3202), .B(n3203), .ZN(n3201) );
  NAND2_X1 U3187 ( .A1(a_0_), .A2(b_7_), .ZN(n3203) );
  NAND2_X1 U3188 ( .A1(n3204), .A2(n3205), .ZN(n2195) );
  INV_X1 U3189 ( .A(n3077), .ZN(n3205) );
  NOR2_X1 U3190 ( .A1(n3206), .A2(n3207), .ZN(n3077) );
  INV_X1 U3191 ( .A(n3208), .ZN(n3207) );
  NAND3_X1 U3192 ( .A1(b_7_), .A2(n3209), .A3(a_0_), .ZN(n3208) );
  NAND2_X1 U3193 ( .A1(n3202), .A2(n3200), .ZN(n3209) );
  NOR2_X1 U3194 ( .A1(n3200), .A2(n3202), .ZN(n3206) );
  NOR2_X1 U3195 ( .A1(n3210), .A2(n3211), .ZN(n3202) );
  NOR3_X1 U3196 ( .A1(n3044), .A2(n3212), .A3(n2343), .ZN(n3211) );
  INV_X1 U3197 ( .A(n3213), .ZN(n3212) );
  NAND2_X1 U3198 ( .A1(n3085), .A2(n3086), .ZN(n3213) );
  NOR2_X1 U3199 ( .A1(n3085), .A2(n3086), .ZN(n3210) );
  NOR2_X1 U3200 ( .A1(n3214), .A2(n3215), .ZN(n3086) );
  NOR3_X1 U3201 ( .A1(n3044), .A2(n3216), .A3(n2139), .ZN(n3215) );
  INV_X1 U3202 ( .A(n3217), .ZN(n3216) );
  NAND2_X1 U3203 ( .A1(n3092), .A2(n3094), .ZN(n3217) );
  NOR2_X1 U3204 ( .A1(n3092), .A2(n3094), .ZN(n3214) );
  NOR2_X1 U3205 ( .A1(n3218), .A2(n3219), .ZN(n3094) );
  NOR3_X1 U3206 ( .A1(n3044), .A2(n3220), .A3(n2322), .ZN(n3219) );
  INV_X1 U3207 ( .A(n3221), .ZN(n3220) );
  NAND2_X1 U3208 ( .A1(n3102), .A2(n3100), .ZN(n3221) );
  NOR2_X1 U3209 ( .A1(n3100), .A2(n3102), .ZN(n3218) );
  NOR2_X1 U3210 ( .A1(n3222), .A2(n3223), .ZN(n3102) );
  NOR3_X1 U3211 ( .A1(n3044), .A2(n3224), .A3(n2230), .ZN(n3223) );
  INV_X1 U3212 ( .A(n3225), .ZN(n3224) );
  NAND2_X1 U3213 ( .A1(n3109), .A2(n3107), .ZN(n3225) );
  NOR2_X1 U3214 ( .A1(n3107), .A2(n3109), .ZN(n3222) );
  NOR2_X1 U3215 ( .A1(n3226), .A2(n3227), .ZN(n3109) );
  NOR3_X1 U3216 ( .A1(n3044), .A2(n3228), .A3(n2366), .ZN(n3227) );
  INV_X1 U3217 ( .A(n3229), .ZN(n3228) );
  NAND2_X1 U3218 ( .A1(n3198), .A2(n3196), .ZN(n3229) );
  NOR2_X1 U3219 ( .A1(n3196), .A2(n3198), .ZN(n3226) );
  NOR2_X1 U3220 ( .A1(n3192), .A2(n3230), .ZN(n3198) );
  INV_X1 U3221 ( .A(n3231), .ZN(n3230) );
  NAND2_X1 U3222 ( .A1(n3189), .A2(n3232), .ZN(n3231) );
  NAND2_X1 U3223 ( .A1(n3195), .A2(n3233), .ZN(n3232) );
  NAND2_X1 U3224 ( .A1(a_6_), .A2(b_7_), .ZN(n3233) );
  XNOR2_X1 U3225 ( .A(n3234), .B(n3235), .ZN(n3189) );
  XNOR2_X1 U3226 ( .A(n3236), .B(n3237), .ZN(n3235) );
  NOR2_X1 U3227 ( .A1(n3195), .A2(n2247), .ZN(n3192) );
  NAND2_X1 U3228 ( .A1(n3238), .A2(n3239), .ZN(n3195) );
  NAND2_X1 U3229 ( .A1(n3186), .A2(n3240), .ZN(n3239) );
  INV_X1 U3230 ( .A(n3241), .ZN(n3240) );
  NOR2_X1 U3231 ( .A1(n3188), .A2(n3187), .ZN(n3241) );
  XOR2_X1 U3232 ( .A(n3242), .B(n3243), .Z(n3186) );
  XOR2_X1 U3233 ( .A(n3244), .B(n3245), .Z(n3243) );
  NAND2_X1 U3234 ( .A1(b_6_), .A2(a_8_), .ZN(n3245) );
  NAND2_X1 U3235 ( .A1(n3187), .A2(n3188), .ZN(n3238) );
  NOR2_X1 U3236 ( .A1(n3246), .A2(n3247), .ZN(n3187) );
  NOR2_X1 U3237 ( .A1(n3131), .A2(n3248), .ZN(n3247) );
  NOR2_X1 U3238 ( .A1(n3130), .A2(n3128), .ZN(n3248) );
  NAND2_X1 U3239 ( .A1(b_7_), .A2(a_8_), .ZN(n3131) );
  INV_X1 U3240 ( .A(n3249), .ZN(n3246) );
  NAND2_X1 U3241 ( .A1(n3128), .A2(n3130), .ZN(n3249) );
  NAND2_X1 U3242 ( .A1(n3139), .A2(n3250), .ZN(n3130) );
  NAND2_X1 U3243 ( .A1(n3138), .A2(n3140), .ZN(n3250) );
  NAND2_X1 U3244 ( .A1(n3251), .A2(n3252), .ZN(n3140) );
  NAND2_X1 U3245 ( .A1(a_9_), .A2(b_7_), .ZN(n3252) );
  INV_X1 U3246 ( .A(n3253), .ZN(n3251) );
  XNOR2_X1 U3247 ( .A(n3254), .B(n3255), .ZN(n3138) );
  NAND2_X1 U3248 ( .A1(n3256), .A2(n3257), .ZN(n3254) );
  NAND2_X1 U3249 ( .A1(a_9_), .A2(n3253), .ZN(n3139) );
  NAND2_X1 U3250 ( .A1(n3147), .A2(n3258), .ZN(n3253) );
  NAND2_X1 U3251 ( .A1(n3146), .A2(n3148), .ZN(n3258) );
  NAND2_X1 U3252 ( .A1(n3259), .A2(n3260), .ZN(n3148) );
  NAND2_X1 U3253 ( .A1(a_10_), .A2(b_7_), .ZN(n3260) );
  XNOR2_X1 U3254 ( .A(n3261), .B(n3262), .ZN(n3146) );
  XOR2_X1 U3255 ( .A(n3263), .B(n3264), .Z(n3261) );
  NAND2_X1 U3256 ( .A1(a_11_), .A2(b_6_), .ZN(n3263) );
  INV_X1 U3257 ( .A(n3265), .ZN(n3147) );
  NOR2_X1 U3258 ( .A1(n2523), .A2(n3259), .ZN(n3265) );
  NOR2_X1 U3259 ( .A1(n3266), .A2(n3267), .ZN(n3259) );
  INV_X1 U3260 ( .A(n3268), .ZN(n3267) );
  NAND3_X1 U3261 ( .A1(b_7_), .A2(n3269), .A3(a_11_), .ZN(n3268) );
  NAND2_X1 U3262 ( .A1(n3153), .A2(n3155), .ZN(n3269) );
  NOR2_X1 U3263 ( .A1(n3153), .A2(n3155), .ZN(n3266) );
  NOR2_X1 U3264 ( .A1(n3270), .A2(n3271), .ZN(n3155) );
  INV_X1 U3265 ( .A(n3272), .ZN(n3271) );
  NAND2_X1 U3266 ( .A1(n3183), .A2(n3273), .ZN(n3272) );
  NAND2_X1 U3267 ( .A1(n3184), .A2(n3182), .ZN(n3273) );
  NOR2_X1 U3268 ( .A1(n3044), .A2(n2094), .ZN(n3183) );
  NOR2_X1 U3269 ( .A1(n3182), .A2(n3184), .ZN(n3270) );
  NOR2_X1 U3270 ( .A1(n3274), .A2(n3275), .ZN(n3184) );
  INV_X1 U3271 ( .A(n3276), .ZN(n3275) );
  NAND2_X1 U3272 ( .A1(n3178), .A2(n3277), .ZN(n3276) );
  NAND2_X1 U3273 ( .A1(n3179), .A2(n3180), .ZN(n3277) );
  NOR2_X1 U3274 ( .A1(n3044), .A2(n2408), .ZN(n3178) );
  NOR2_X1 U3275 ( .A1(n3180), .A2(n3179), .ZN(n3274) );
  INV_X1 U3276 ( .A(n3278), .ZN(n3179) );
  NAND2_X1 U3277 ( .A1(n3279), .A2(n3280), .ZN(n3278) );
  NAND2_X1 U3278 ( .A1(b_5_), .A2(n3281), .ZN(n3280) );
  NAND2_X1 U3279 ( .A1(n2077), .A2(n3282), .ZN(n3281) );
  NAND2_X1 U3280 ( .A1(a_15_), .A2(n3176), .ZN(n3282) );
  NAND2_X1 U3281 ( .A1(b_6_), .A2(n3283), .ZN(n3279) );
  NAND2_X1 U3282 ( .A1(n2081), .A2(n3284), .ZN(n3283) );
  NAND2_X1 U3283 ( .A1(a_14_), .A2(n3285), .ZN(n3284) );
  NAND3_X1 U3284 ( .A1(b_7_), .A2(n2417), .A3(b_6_), .ZN(n3180) );
  XNOR2_X1 U3285 ( .A(n3286), .B(n3287), .ZN(n3182) );
  XOR2_X1 U3286 ( .A(n3288), .B(n3289), .Z(n3286) );
  XOR2_X1 U3287 ( .A(n3290), .B(n3291), .Z(n3153) );
  XNOR2_X1 U3288 ( .A(n3292), .B(n3293), .ZN(n3290) );
  XNOR2_X1 U3289 ( .A(n3294), .B(n3295), .ZN(n3128) );
  NAND2_X1 U3290 ( .A1(n3296), .A2(n3297), .ZN(n3294) );
  XNOR2_X1 U3291 ( .A(n3298), .B(n3299), .ZN(n3196) );
  XNOR2_X1 U3292 ( .A(n3300), .B(n3301), .ZN(n3298) );
  XNOR2_X1 U3293 ( .A(n3302), .B(n3303), .ZN(n3107) );
  XOR2_X1 U3294 ( .A(n3304), .B(n3305), .Z(n3302) );
  XNOR2_X1 U3295 ( .A(n3306), .B(n3307), .ZN(n3100) );
  XOR2_X1 U3296 ( .A(n3308), .B(n3309), .Z(n3306) );
  XNOR2_X1 U3297 ( .A(n3310), .B(n3311), .ZN(n3092) );
  XOR2_X1 U3298 ( .A(n3312), .B(n3313), .Z(n3311) );
  XOR2_X1 U3299 ( .A(n3314), .B(n3315), .Z(n3085) );
  XNOR2_X1 U3300 ( .A(n3316), .B(n3317), .ZN(n3314) );
  XNOR2_X1 U3301 ( .A(n3318), .B(n3319), .ZN(n3200) );
  XNOR2_X1 U3302 ( .A(n3320), .B(n3321), .ZN(n3319) );
  NAND2_X1 U3303 ( .A1(a_1_), .A2(b_6_), .ZN(n3321) );
  XNOR2_X1 U3304 ( .A(n3078), .B(n3079), .ZN(n3204) );
  XNOR2_X1 U3305 ( .A(n3322), .B(n3323), .ZN(n3078) );
  NOR2_X1 U3306 ( .A1(n3176), .A2(n2212), .ZN(n3323) );
  XOR2_X1 U3307 ( .A(n2063), .B(n2062), .Z(n2055) );
  NAND3_X1 U3308 ( .A1(n2062), .A2(n2063), .A3(n2194), .ZN(n2058) );
  INV_X1 U3309 ( .A(n2061), .ZN(n2194) );
  NAND2_X1 U3310 ( .A1(n3324), .A2(n2192), .ZN(n2061) );
  NAND2_X1 U3311 ( .A1(n3325), .A2(n3326), .ZN(n3324) );
  XOR2_X1 U3312 ( .A(n3327), .B(n3328), .Z(n3325) );
  NAND2_X1 U3313 ( .A1(n3329), .A2(n3330), .ZN(n2063) );
  NAND3_X1 U3314 ( .A1(b_6_), .A2(n3331), .A3(a_0_), .ZN(n3330) );
  INV_X1 U3315 ( .A(n3332), .ZN(n3331) );
  NOR2_X1 U3316 ( .A1(n3322), .A2(n3079), .ZN(n3332) );
  NAND2_X1 U3317 ( .A1(n3079), .A2(n3322), .ZN(n3329) );
  NAND2_X1 U3318 ( .A1(n3333), .A2(n3334), .ZN(n3322) );
  NAND3_X1 U3319 ( .A1(b_6_), .A2(n3335), .A3(a_1_), .ZN(n3334) );
  NAND2_X1 U3320 ( .A1(n3318), .A2(n3320), .ZN(n3335) );
  INV_X1 U3321 ( .A(n3336), .ZN(n3333) );
  NOR2_X1 U3322 ( .A1(n3318), .A2(n3320), .ZN(n3336) );
  NOR2_X1 U3323 ( .A1(n3337), .A2(n3338), .ZN(n3320) );
  INV_X1 U3324 ( .A(n3339), .ZN(n3338) );
  NAND2_X1 U3325 ( .A1(n3317), .A2(n3340), .ZN(n3339) );
  NAND2_X1 U3326 ( .A1(n3316), .A2(n3315), .ZN(n3340) );
  NOR2_X1 U3327 ( .A1(n2139), .A2(n3176), .ZN(n3317) );
  NOR2_X1 U3328 ( .A1(n3315), .A2(n3316), .ZN(n3337) );
  NOR2_X1 U3329 ( .A1(n3341), .A2(n3342), .ZN(n3316) );
  INV_X1 U3330 ( .A(n3343), .ZN(n3342) );
  NAND2_X1 U3331 ( .A1(n3313), .A2(n3344), .ZN(n3343) );
  NAND2_X1 U3332 ( .A1(n3312), .A2(n3310), .ZN(n3344) );
  NOR2_X1 U3333 ( .A1(n2322), .A2(n3176), .ZN(n3313) );
  NOR2_X1 U3334 ( .A1(n3310), .A2(n3312), .ZN(n3341) );
  INV_X1 U3335 ( .A(n3345), .ZN(n3312) );
  NAND2_X1 U3336 ( .A1(n3346), .A2(n3347), .ZN(n3345) );
  NAND2_X1 U3337 ( .A1(n3309), .A2(n3348), .ZN(n3347) );
  INV_X1 U3338 ( .A(n3349), .ZN(n3348) );
  NOR2_X1 U3339 ( .A1(n3307), .A2(n3308), .ZN(n3349) );
  NOR2_X1 U3340 ( .A1(n2230), .A2(n3176), .ZN(n3309) );
  NAND2_X1 U3341 ( .A1(n3307), .A2(n3308), .ZN(n3346) );
  NAND2_X1 U3342 ( .A1(n3350), .A2(n3351), .ZN(n3308) );
  NAND2_X1 U3343 ( .A1(n3305), .A2(n3352), .ZN(n3351) );
  NAND2_X1 U3344 ( .A1(n3303), .A2(n3304), .ZN(n3352) );
  NOR2_X1 U3345 ( .A1(n2366), .A2(n3176), .ZN(n3305) );
  INV_X1 U3346 ( .A(n3353), .ZN(n3350) );
  NOR2_X1 U3347 ( .A1(n3303), .A2(n3304), .ZN(n3353) );
  NAND2_X1 U3348 ( .A1(n3354), .A2(n3355), .ZN(n3304) );
  NAND2_X1 U3349 ( .A1(n3356), .A2(n3301), .ZN(n3355) );
  NAND2_X1 U3350 ( .A1(n3299), .A2(n3300), .ZN(n3356) );
  INV_X1 U3351 ( .A(n3357), .ZN(n3354) );
  NOR2_X1 U3352 ( .A1(n3299), .A2(n3300), .ZN(n3357) );
  NAND2_X1 U3353 ( .A1(n3358), .A2(n3359), .ZN(n3300) );
  NAND2_X1 U3354 ( .A1(n3237), .A2(n3360), .ZN(n3359) );
  INV_X1 U3355 ( .A(n3361), .ZN(n3360) );
  NOR2_X1 U3356 ( .A1(n3236), .A2(n3234), .ZN(n3361) );
  NOR2_X1 U3357 ( .A1(n2626), .A2(n3176), .ZN(n3237) );
  NAND2_X1 U3358 ( .A1(n3234), .A2(n3236), .ZN(n3358) );
  NAND2_X1 U3359 ( .A1(n3362), .A2(n3363), .ZN(n3236) );
  NAND3_X1 U3360 ( .A1(a_8_), .A2(n3364), .A3(b_6_), .ZN(n3363) );
  INV_X1 U3361 ( .A(n3365), .ZN(n3364) );
  NOR2_X1 U3362 ( .A1(n3244), .A2(n3242), .ZN(n3365) );
  NAND2_X1 U3363 ( .A1(n3242), .A2(n3244), .ZN(n3362) );
  NAND2_X1 U3364 ( .A1(n3296), .A2(n3366), .ZN(n3244) );
  NAND2_X1 U3365 ( .A1(n3295), .A2(n3297), .ZN(n3366) );
  NAND2_X1 U3366 ( .A1(n3367), .A2(n3368), .ZN(n3297) );
  NAND2_X1 U3367 ( .A1(a_9_), .A2(b_6_), .ZN(n3368) );
  INV_X1 U3368 ( .A(n3369), .ZN(n3367) );
  XNOR2_X1 U3369 ( .A(n3370), .B(n3371), .ZN(n3295) );
  NAND2_X1 U3370 ( .A1(n3372), .A2(n3373), .ZN(n3370) );
  NAND2_X1 U3371 ( .A1(a_9_), .A2(n3369), .ZN(n3296) );
  NAND2_X1 U3372 ( .A1(n3256), .A2(n3374), .ZN(n3369) );
  NAND2_X1 U3373 ( .A1(n3255), .A2(n3257), .ZN(n3374) );
  NAND2_X1 U3374 ( .A1(n3375), .A2(n3376), .ZN(n3257) );
  NAND2_X1 U3375 ( .A1(a_10_), .A2(b_6_), .ZN(n3376) );
  XNOR2_X1 U3376 ( .A(n3377), .B(n3378), .ZN(n3255) );
  XOR2_X1 U3377 ( .A(n3379), .B(n3380), .Z(n3377) );
  NAND2_X1 U3378 ( .A1(a_11_), .A2(b_5_), .ZN(n3379) );
  INV_X1 U3379 ( .A(n3381), .ZN(n3256) );
  NOR2_X1 U3380 ( .A1(n2523), .A2(n3375), .ZN(n3381) );
  NOR2_X1 U3381 ( .A1(n3382), .A2(n3383), .ZN(n3375) );
  INV_X1 U3382 ( .A(n3384), .ZN(n3383) );
  NAND3_X1 U3383 ( .A1(b_6_), .A2(n3385), .A3(a_11_), .ZN(n3384) );
  NAND2_X1 U3384 ( .A1(n3262), .A2(n3264), .ZN(n3385) );
  NOR2_X1 U3385 ( .A1(n3262), .A2(n3264), .ZN(n3382) );
  NOR2_X1 U3386 ( .A1(n3386), .A2(n3387), .ZN(n3264) );
  INV_X1 U3387 ( .A(n3388), .ZN(n3387) );
  NAND2_X1 U3388 ( .A1(n3292), .A2(n3389), .ZN(n3388) );
  NAND2_X1 U3389 ( .A1(n3293), .A2(n3291), .ZN(n3389) );
  NOR2_X1 U3390 ( .A1(n3176), .A2(n2094), .ZN(n3292) );
  NOR2_X1 U3391 ( .A1(n3291), .A2(n3293), .ZN(n3386) );
  NOR2_X1 U3392 ( .A1(n3390), .A2(n3391), .ZN(n3293) );
  INV_X1 U3393 ( .A(n3392), .ZN(n3391) );
  NAND2_X1 U3394 ( .A1(n3287), .A2(n3393), .ZN(n3392) );
  NAND2_X1 U3395 ( .A1(n3288), .A2(n3289), .ZN(n3393) );
  NOR2_X1 U3396 ( .A1(n3176), .A2(n2408), .ZN(n3287) );
  NOR2_X1 U3397 ( .A1(n3289), .A2(n3288), .ZN(n3390) );
  INV_X1 U3398 ( .A(n3394), .ZN(n3288) );
  NAND2_X1 U3399 ( .A1(n3395), .A2(n3396), .ZN(n3394) );
  NAND2_X1 U3400 ( .A1(b_4_), .A2(n3397), .ZN(n3396) );
  NAND2_X1 U3401 ( .A1(n2077), .A2(n3398), .ZN(n3397) );
  NAND2_X1 U3402 ( .A1(a_15_), .A2(n3285), .ZN(n3398) );
  NAND2_X1 U3403 ( .A1(b_5_), .A2(n3399), .ZN(n3395) );
  NAND2_X1 U3404 ( .A1(n2081), .A2(n3400), .ZN(n3399) );
  NAND2_X1 U3405 ( .A1(a_14_), .A2(n3401), .ZN(n3400) );
  NAND3_X1 U3406 ( .A1(b_6_), .A2(n2417), .A3(b_5_), .ZN(n3289) );
  XNOR2_X1 U3407 ( .A(n3402), .B(n3403), .ZN(n3291) );
  XOR2_X1 U3408 ( .A(n3404), .B(n3405), .Z(n3402) );
  XOR2_X1 U3409 ( .A(n3406), .B(n3407), .Z(n3262) );
  XNOR2_X1 U3410 ( .A(n3408), .B(n3409), .ZN(n3406) );
  XNOR2_X1 U3411 ( .A(n3410), .B(n3411), .ZN(n3242) );
  NAND2_X1 U3412 ( .A1(n3412), .A2(n3413), .ZN(n3410) );
  XNOR2_X1 U3413 ( .A(n3414), .B(n3415), .ZN(n3234) );
  XOR2_X1 U3414 ( .A(n3416), .B(n3417), .Z(n3415) );
  NAND2_X1 U3415 ( .A1(b_5_), .A2(a_8_), .ZN(n3417) );
  XOR2_X1 U3416 ( .A(n3418), .B(n3419), .Z(n3299) );
  XNOR2_X1 U3417 ( .A(n3420), .B(n3421), .ZN(n3419) );
  NAND2_X1 U3418 ( .A1(a_7_), .A2(b_5_), .ZN(n3421) );
  XNOR2_X1 U3419 ( .A(n3422), .B(n3423), .ZN(n3303) );
  XNOR2_X1 U3420 ( .A(n3424), .B(n3425), .ZN(n3423) );
  NAND2_X1 U3421 ( .A1(a_6_), .A2(b_5_), .ZN(n3425) );
  XOR2_X1 U3422 ( .A(n3426), .B(n3427), .Z(n3307) );
  XOR2_X1 U3423 ( .A(n3428), .B(n3429), .Z(n3426) );
  XOR2_X1 U3424 ( .A(n3430), .B(n3431), .Z(n3310) );
  XNOR2_X1 U3425 ( .A(n3432), .B(n3433), .ZN(n3430) );
  NOR2_X1 U3426 ( .A1(n3285), .A2(n2230), .ZN(n3433) );
  XOR2_X1 U3427 ( .A(n3434), .B(n3435), .Z(n3315) );
  XNOR2_X1 U3428 ( .A(n3436), .B(n3437), .ZN(n3434) );
  NOR2_X1 U3429 ( .A1(n3285), .A2(n2322), .ZN(n3437) );
  XOR2_X1 U3430 ( .A(n3438), .B(n3439), .Z(n3318) );
  XNOR2_X1 U3431 ( .A(n3440), .B(n3441), .ZN(n3438) );
  NOR2_X1 U3432 ( .A1(n3285), .A2(n2139), .ZN(n3441) );
  XNOR2_X1 U3433 ( .A(n3442), .B(n3443), .ZN(n3079) );
  XNOR2_X1 U3434 ( .A(n3444), .B(n3445), .ZN(n3442) );
  NOR2_X1 U3435 ( .A1(n3285), .A2(n2343), .ZN(n3445) );
  XNOR2_X1 U3436 ( .A(n3446), .B(n3447), .ZN(n2062) );
  XNOR2_X1 U3437 ( .A(n3448), .B(n3449), .ZN(n3446) );
  NOR2_X1 U3438 ( .A1(n3285), .A2(n2212), .ZN(n3449) );
  NAND2_X1 U3439 ( .A1(n3450), .A2(n3451), .ZN(n2192) );
  INV_X1 U3440 ( .A(n3326), .ZN(n3451) );
  NOR2_X1 U3441 ( .A1(n3452), .A2(n3453), .ZN(n3326) );
  INV_X1 U3442 ( .A(n3454), .ZN(n3453) );
  NAND3_X1 U3443 ( .A1(b_5_), .A2(n3455), .A3(a_0_), .ZN(n3454) );
  NAND2_X1 U3444 ( .A1(n3448), .A2(n3447), .ZN(n3455) );
  NOR2_X1 U3445 ( .A1(n3447), .A2(n3448), .ZN(n3452) );
  NOR2_X1 U3446 ( .A1(n3456), .A2(n3457), .ZN(n3448) );
  NOR3_X1 U3447 ( .A1(n3285), .A2(n3458), .A3(n2343), .ZN(n3457) );
  INV_X1 U3448 ( .A(n3459), .ZN(n3458) );
  NAND2_X1 U3449 ( .A1(n3443), .A2(n3444), .ZN(n3459) );
  NOR2_X1 U3450 ( .A1(n3443), .A2(n3444), .ZN(n3456) );
  NOR2_X1 U3451 ( .A1(n3460), .A2(n3461), .ZN(n3444) );
  NOR3_X1 U3452 ( .A1(n3285), .A2(n3462), .A3(n2139), .ZN(n3461) );
  INV_X1 U3453 ( .A(n3463), .ZN(n3462) );
  NAND2_X1 U3454 ( .A1(n3440), .A2(n3439), .ZN(n3463) );
  NOR2_X1 U3455 ( .A1(n3439), .A2(n3440), .ZN(n3460) );
  NOR2_X1 U3456 ( .A1(n3464), .A2(n3465), .ZN(n3440) );
  NOR3_X1 U3457 ( .A1(n3285), .A2(n3466), .A3(n2322), .ZN(n3465) );
  INV_X1 U3458 ( .A(n3467), .ZN(n3466) );
  NAND2_X1 U3459 ( .A1(n3435), .A2(n3436), .ZN(n3467) );
  NOR2_X1 U3460 ( .A1(n3435), .A2(n3436), .ZN(n3464) );
  NOR2_X1 U3461 ( .A1(n3468), .A2(n3469), .ZN(n3436) );
  NOR3_X1 U3462 ( .A1(n3285), .A2(n3470), .A3(n2230), .ZN(n3469) );
  INV_X1 U3463 ( .A(n3471), .ZN(n3470) );
  NAND2_X1 U3464 ( .A1(n3431), .A2(n3432), .ZN(n3471) );
  NOR2_X1 U3465 ( .A1(n3431), .A2(n3432), .ZN(n3468) );
  NOR2_X1 U3466 ( .A1(n3472), .A2(n3473), .ZN(n3432) );
  INV_X1 U3467 ( .A(n3474), .ZN(n3473) );
  NAND2_X1 U3468 ( .A1(n3427), .A2(n3475), .ZN(n3474) );
  NAND2_X1 U3469 ( .A1(n3428), .A2(n3429), .ZN(n3475) );
  XNOR2_X1 U3470 ( .A(n3476), .B(n3477), .ZN(n3427) );
  XNOR2_X1 U3471 ( .A(n3478), .B(n3479), .ZN(n3476) );
  NOR2_X1 U3472 ( .A1(n3429), .A2(n3428), .ZN(n3472) );
  NOR2_X1 U3473 ( .A1(n3480), .A2(n3481), .ZN(n3428) );
  NOR3_X1 U3474 ( .A1(n3285), .A2(n3482), .A3(n2247), .ZN(n3481) );
  INV_X1 U3475 ( .A(n3483), .ZN(n3482) );
  NAND2_X1 U3476 ( .A1(n3422), .A2(n3424), .ZN(n3483) );
  NOR2_X1 U3477 ( .A1(n3422), .A2(n3424), .ZN(n3480) );
  NOR2_X1 U3478 ( .A1(n3484), .A2(n3485), .ZN(n3424) );
  NOR3_X1 U3479 ( .A1(n3285), .A2(n3486), .A3(n2626), .ZN(n3485) );
  INV_X1 U3480 ( .A(n3487), .ZN(n3486) );
  NAND2_X1 U3481 ( .A1(n3420), .A2(n3418), .ZN(n3487) );
  NOR2_X1 U3482 ( .A1(n3418), .A2(n3420), .ZN(n3484) );
  NOR2_X1 U3483 ( .A1(n3488), .A2(n3489), .ZN(n3420) );
  NOR3_X1 U3484 ( .A1(n2377), .A2(n3490), .A3(n3285), .ZN(n3489) );
  NOR2_X1 U3485 ( .A1(n3414), .A2(n3416), .ZN(n3490) );
  INV_X1 U3486 ( .A(n3491), .ZN(n3488) );
  NAND2_X1 U3487 ( .A1(n3414), .A2(n3416), .ZN(n3491) );
  NAND2_X1 U3488 ( .A1(n3412), .A2(n3492), .ZN(n3416) );
  NAND2_X1 U3489 ( .A1(n3411), .A2(n3413), .ZN(n3492) );
  NAND2_X1 U3490 ( .A1(n3493), .A2(n3494), .ZN(n3413) );
  NAND2_X1 U3491 ( .A1(a_9_), .A2(b_5_), .ZN(n3494) );
  INV_X1 U3492 ( .A(n3495), .ZN(n3493) );
  XOR2_X1 U3493 ( .A(n3496), .B(n3497), .Z(n3411) );
  XNOR2_X1 U3494 ( .A(n3498), .B(n3499), .ZN(n3497) );
  NAND2_X1 U3495 ( .A1(a_9_), .A2(n3495), .ZN(n3412) );
  NAND2_X1 U3496 ( .A1(n3372), .A2(n3500), .ZN(n3495) );
  NAND2_X1 U3497 ( .A1(n3371), .A2(n3373), .ZN(n3500) );
  NAND2_X1 U3498 ( .A1(n3501), .A2(n3502), .ZN(n3373) );
  NAND2_X1 U3499 ( .A1(a_10_), .A2(b_5_), .ZN(n3502) );
  XNOR2_X1 U3500 ( .A(n3503), .B(n3504), .ZN(n3371) );
  XOR2_X1 U3501 ( .A(n3505), .B(n3506), .Z(n3503) );
  NAND2_X1 U3502 ( .A1(b_4_), .A2(a_11_), .ZN(n3505) );
  INV_X1 U3503 ( .A(n3507), .ZN(n3372) );
  NOR2_X1 U3504 ( .A1(n2523), .A2(n3501), .ZN(n3507) );
  NOR2_X1 U3505 ( .A1(n3508), .A2(n3509), .ZN(n3501) );
  INV_X1 U3506 ( .A(n3510), .ZN(n3509) );
  NAND3_X1 U3507 ( .A1(b_5_), .A2(n3511), .A3(a_11_), .ZN(n3510) );
  NAND2_X1 U3508 ( .A1(n3378), .A2(n3380), .ZN(n3511) );
  NOR2_X1 U3509 ( .A1(n3378), .A2(n3380), .ZN(n3508) );
  NOR2_X1 U3510 ( .A1(n3512), .A2(n3513), .ZN(n3380) );
  INV_X1 U3511 ( .A(n3514), .ZN(n3513) );
  NAND2_X1 U3512 ( .A1(n3408), .A2(n3515), .ZN(n3514) );
  NAND2_X1 U3513 ( .A1(n3409), .A2(n3407), .ZN(n3515) );
  NOR2_X1 U3514 ( .A1(n3285), .A2(n2094), .ZN(n3408) );
  NOR2_X1 U3515 ( .A1(n3407), .A2(n3409), .ZN(n3512) );
  NOR2_X1 U3516 ( .A1(n3516), .A2(n3517), .ZN(n3409) );
  INV_X1 U3517 ( .A(n3518), .ZN(n3517) );
  NAND2_X1 U3518 ( .A1(n3403), .A2(n3519), .ZN(n3518) );
  NAND2_X1 U3519 ( .A1(n3404), .A2(n3405), .ZN(n3519) );
  NOR2_X1 U3520 ( .A1(n3285), .A2(n2408), .ZN(n3403) );
  NOR2_X1 U3521 ( .A1(n3405), .A2(n3404), .ZN(n3516) );
  INV_X1 U3522 ( .A(n3520), .ZN(n3404) );
  NAND2_X1 U3523 ( .A1(n3521), .A2(n3522), .ZN(n3520) );
  NAND2_X1 U3524 ( .A1(b_3_), .A2(n3523), .ZN(n3522) );
  NAND2_X1 U3525 ( .A1(n2077), .A2(n3524), .ZN(n3523) );
  NAND2_X1 U3526 ( .A1(a_15_), .A2(n3401), .ZN(n3524) );
  NAND2_X1 U3527 ( .A1(b_4_), .A2(n3525), .ZN(n3521) );
  NAND2_X1 U3528 ( .A1(n2081), .A2(n3526), .ZN(n3525) );
  NAND2_X1 U3529 ( .A1(a_14_), .A2(n3527), .ZN(n3526) );
  NAND3_X1 U3530 ( .A1(b_5_), .A2(n2417), .A3(b_4_), .ZN(n3405) );
  XNOR2_X1 U3531 ( .A(n3528), .B(n3529), .ZN(n3407) );
  XOR2_X1 U3532 ( .A(n3530), .B(n3531), .Z(n3528) );
  XOR2_X1 U3533 ( .A(n3532), .B(n3533), .Z(n3378) );
  XNOR2_X1 U3534 ( .A(n3534), .B(n3535), .ZN(n3532) );
  XNOR2_X1 U3535 ( .A(n3536), .B(n3537), .ZN(n3414) );
  XNOR2_X1 U3536 ( .A(n3538), .B(n3539), .ZN(n3537) );
  XOR2_X1 U3537 ( .A(n3540), .B(n3541), .Z(n3418) );
  XNOR2_X1 U3538 ( .A(n3542), .B(n3543), .ZN(n3540) );
  XOR2_X1 U3539 ( .A(n3544), .B(n3545), .Z(n3422) );
  XNOR2_X1 U3540 ( .A(n3546), .B(n3547), .ZN(n3544) );
  XOR2_X1 U3541 ( .A(n3548), .B(n3549), .Z(n3431) );
  XNOR2_X1 U3542 ( .A(n3550), .B(n3551), .ZN(n3548) );
  XNOR2_X1 U3543 ( .A(n3552), .B(n3553), .ZN(n3435) );
  XOR2_X1 U3544 ( .A(n3554), .B(n3555), .Z(n3552) );
  XOR2_X1 U3545 ( .A(n3556), .B(n3557), .Z(n3439) );
  XNOR2_X1 U3546 ( .A(n3558), .B(n3559), .ZN(n3556) );
  XOR2_X1 U3547 ( .A(n3560), .B(n3561), .Z(n3443) );
  XNOR2_X1 U3548 ( .A(n3562), .B(n3563), .ZN(n3561) );
  XNOR2_X1 U3549 ( .A(n3564), .B(n3565), .ZN(n3447) );
  XNOR2_X1 U3550 ( .A(n3566), .B(n3567), .ZN(n3564) );
  NAND2_X1 U3551 ( .A1(a_1_), .A2(b_4_), .ZN(n3566) );
  XNOR2_X1 U3552 ( .A(n3328), .B(n3327), .ZN(n3450) );
  XNOR2_X1 U3553 ( .A(n3568), .B(n3569), .ZN(n3328) );
  NOR2_X1 U3554 ( .A1(n3401), .A2(n2212), .ZN(n3569) );
  XOR2_X1 U3555 ( .A(n2073), .B(n2072), .Z(n2065) );
  NAND3_X1 U3556 ( .A1(n2072), .A2(n2073), .A3(n2191), .ZN(n2068) );
  INV_X1 U3557 ( .A(n2071), .ZN(n2191) );
  NAND2_X1 U3558 ( .A1(n3570), .A2(n2189), .ZN(n2071) );
  NAND2_X1 U3559 ( .A1(n3571), .A2(n3572), .ZN(n3570) );
  XOR2_X1 U3560 ( .A(n3573), .B(n3574), .Z(n3572) );
  NAND2_X1 U3561 ( .A1(n3575), .A2(n3576), .ZN(n2073) );
  NAND3_X1 U3562 ( .A1(b_4_), .A2(n3577), .A3(a_0_), .ZN(n3576) );
  INV_X1 U3563 ( .A(n3578), .ZN(n3577) );
  NOR2_X1 U3564 ( .A1(n3568), .A2(n3327), .ZN(n3578) );
  NAND2_X1 U3565 ( .A1(n3327), .A2(n3568), .ZN(n3575) );
  NAND2_X1 U3566 ( .A1(n3579), .A2(n3580), .ZN(n3568) );
  NAND3_X1 U3567 ( .A1(b_4_), .A2(n3581), .A3(a_1_), .ZN(n3580) );
  INV_X1 U3568 ( .A(n3582), .ZN(n3581) );
  NOR2_X1 U3569 ( .A1(n3565), .A2(n3567), .ZN(n3582) );
  NAND2_X1 U3570 ( .A1(n3565), .A2(n3567), .ZN(n3579) );
  NAND2_X1 U3571 ( .A1(n3583), .A2(n3584), .ZN(n3567) );
  NAND2_X1 U3572 ( .A1(n3563), .A2(n3585), .ZN(n3584) );
  INV_X1 U3573 ( .A(n3586), .ZN(n3585) );
  NOR2_X1 U3574 ( .A1(n3562), .A2(n3560), .ZN(n3586) );
  NOR2_X1 U3575 ( .A1(n2139), .A2(n3401), .ZN(n3563) );
  NAND2_X1 U3576 ( .A1(n3560), .A2(n3562), .ZN(n3583) );
  NAND2_X1 U3577 ( .A1(n3587), .A2(n3588), .ZN(n3562) );
  NAND2_X1 U3578 ( .A1(n3559), .A2(n3589), .ZN(n3588) );
  INV_X1 U3579 ( .A(n3590), .ZN(n3589) );
  NOR2_X1 U3580 ( .A1(n3557), .A2(n3558), .ZN(n3590) );
  NOR2_X1 U3581 ( .A1(n2322), .A2(n3401), .ZN(n3559) );
  NAND2_X1 U3582 ( .A1(n3557), .A2(n3558), .ZN(n3587) );
  NOR2_X1 U3583 ( .A1(n3591), .A2(n3592), .ZN(n3558) );
  NOR2_X1 U3584 ( .A1(n3593), .A2(n3555), .ZN(n3592) );
  INV_X1 U3585 ( .A(n3594), .ZN(n3593) );
  NAND2_X1 U3586 ( .A1(n3553), .A2(n3554), .ZN(n3594) );
  NOR2_X1 U3587 ( .A1(n3554), .A2(n3553), .ZN(n3591) );
  XOR2_X1 U3588 ( .A(n3595), .B(n3596), .Z(n3553) );
  XNOR2_X1 U3589 ( .A(n3597), .B(n3598), .ZN(n3595) );
  NAND2_X1 U3590 ( .A1(a_5_), .A2(b_3_), .ZN(n3597) );
  NAND2_X1 U3591 ( .A1(n3599), .A2(n3600), .ZN(n3554) );
  NAND2_X1 U3592 ( .A1(n3551), .A2(n3601), .ZN(n3600) );
  NAND2_X1 U3593 ( .A1(n3550), .A2(n3549), .ZN(n3601) );
  NOR2_X1 U3594 ( .A1(n2366), .A2(n3401), .ZN(n3551) );
  INV_X1 U3595 ( .A(n3602), .ZN(n3599) );
  NOR2_X1 U3596 ( .A1(n3549), .A2(n3550), .ZN(n3602) );
  NOR2_X1 U3597 ( .A1(n3603), .A2(n3604), .ZN(n3550) );
  INV_X1 U3598 ( .A(n3605), .ZN(n3604) );
  NAND2_X1 U3599 ( .A1(n3479), .A2(n3606), .ZN(n3605) );
  NAND2_X1 U3600 ( .A1(n3477), .A2(n3478), .ZN(n3606) );
  NOR2_X1 U3601 ( .A1(n2247), .A2(n3401), .ZN(n3479) );
  NOR2_X1 U3602 ( .A1(n3477), .A2(n3478), .ZN(n3603) );
  NOR2_X1 U3603 ( .A1(n3607), .A2(n3608), .ZN(n3478) );
  INV_X1 U3604 ( .A(n3609), .ZN(n3608) );
  NAND2_X1 U3605 ( .A1(n3547), .A2(n3610), .ZN(n3609) );
  NAND2_X1 U3606 ( .A1(n3546), .A2(n3545), .ZN(n3610) );
  NOR2_X1 U3607 ( .A1(n2626), .A2(n3401), .ZN(n3547) );
  NOR2_X1 U3608 ( .A1(n3545), .A2(n3546), .ZN(n3607) );
  NOR2_X1 U3609 ( .A1(n3611), .A2(n3612), .ZN(n3546) );
  INV_X1 U3610 ( .A(n3613), .ZN(n3612) );
  NAND2_X1 U3611 ( .A1(n3543), .A2(n3614), .ZN(n3613) );
  NAND2_X1 U3612 ( .A1(n3541), .A2(n3542), .ZN(n3614) );
  NOR2_X1 U3613 ( .A1(n3401), .A2(n2377), .ZN(n3543) );
  NOR2_X1 U3614 ( .A1(n3541), .A2(n3542), .ZN(n3611) );
  NOR2_X1 U3615 ( .A1(n3615), .A2(n3616), .ZN(n3542) );
  INV_X1 U3616 ( .A(n3617), .ZN(n3616) );
  NAND2_X1 U3617 ( .A1(n3539), .A2(n3618), .ZN(n3617) );
  NAND2_X1 U3618 ( .A1(n3536), .A2(n3538), .ZN(n3618) );
  NOR2_X1 U3619 ( .A1(n2275), .A2(n3401), .ZN(n3539) );
  NOR2_X1 U3620 ( .A1(n3538), .A2(n3536), .ZN(n3615) );
  XOR2_X1 U3621 ( .A(n3619), .B(n3620), .Z(n3536) );
  NAND2_X1 U3622 ( .A1(n3621), .A2(n3622), .ZN(n3619) );
  NAND2_X1 U3623 ( .A1(n3623), .A2(n3624), .ZN(n3538) );
  NAND2_X1 U3624 ( .A1(n3496), .A2(n3625), .ZN(n3624) );
  INV_X1 U3625 ( .A(n3626), .ZN(n3625) );
  NOR2_X1 U3626 ( .A1(n3499), .A2(n3498), .ZN(n3626) );
  XOR2_X1 U3627 ( .A(n3627), .B(n3628), .Z(n3496) );
  XOR2_X1 U3628 ( .A(n3629), .B(n3630), .Z(n3627) );
  NAND2_X1 U3629 ( .A1(b_3_), .A2(a_11_), .ZN(n3629) );
  NAND2_X1 U3630 ( .A1(n3498), .A2(n3499), .ZN(n3623) );
  NAND2_X1 U3631 ( .A1(b_4_), .A2(a_10_), .ZN(n3499) );
  NOR2_X1 U3632 ( .A1(n3631), .A2(n3632), .ZN(n3498) );
  NOR3_X1 U3633 ( .A1(n2284), .A2(n3633), .A3(n3401), .ZN(n3632) );
  INV_X1 U3634 ( .A(n3634), .ZN(n3633) );
  NAND2_X1 U3635 ( .A1(n3504), .A2(n3506), .ZN(n3634) );
  NOR2_X1 U3636 ( .A1(n3504), .A2(n3506), .ZN(n3631) );
  NOR2_X1 U3637 ( .A1(n3635), .A2(n3636), .ZN(n3506) );
  INV_X1 U3638 ( .A(n3637), .ZN(n3636) );
  NAND2_X1 U3639 ( .A1(n3534), .A2(n3638), .ZN(n3637) );
  NAND2_X1 U3640 ( .A1(n3535), .A2(n3533), .ZN(n3638) );
  NOR2_X1 U3641 ( .A1(n3401), .A2(n2094), .ZN(n3534) );
  NOR2_X1 U3642 ( .A1(n3533), .A2(n3535), .ZN(n3635) );
  NOR2_X1 U3643 ( .A1(n3639), .A2(n3640), .ZN(n3535) );
  INV_X1 U3644 ( .A(n3641), .ZN(n3640) );
  NAND2_X1 U3645 ( .A1(n3529), .A2(n3642), .ZN(n3641) );
  NAND2_X1 U3646 ( .A1(n3530), .A2(n3531), .ZN(n3642) );
  NOR2_X1 U3647 ( .A1(n3401), .A2(n2408), .ZN(n3529) );
  NOR2_X1 U3648 ( .A1(n3531), .A2(n3530), .ZN(n3639) );
  INV_X1 U3649 ( .A(n3643), .ZN(n3530) );
  NAND2_X1 U3650 ( .A1(n3644), .A2(n3645), .ZN(n3643) );
  NAND2_X1 U3651 ( .A1(b_2_), .A2(n3646), .ZN(n3645) );
  NAND2_X1 U3652 ( .A1(n2077), .A2(n3647), .ZN(n3646) );
  NAND2_X1 U3653 ( .A1(a_15_), .A2(n3527), .ZN(n3647) );
  NAND2_X1 U3654 ( .A1(b_3_), .A2(n3648), .ZN(n3644) );
  NAND2_X1 U3655 ( .A1(n2081), .A2(n3649), .ZN(n3648) );
  NAND2_X1 U3656 ( .A1(a_14_), .A2(n3650), .ZN(n3649) );
  NAND3_X1 U3657 ( .A1(b_4_), .A2(n2417), .A3(b_3_), .ZN(n3531) );
  XNOR2_X1 U3658 ( .A(n3651), .B(n3652), .ZN(n3533) );
  XOR2_X1 U3659 ( .A(n3653), .B(n3654), .Z(n3651) );
  XOR2_X1 U3660 ( .A(n3655), .B(n3656), .Z(n3504) );
  XNOR2_X1 U3661 ( .A(n3657), .B(n3658), .ZN(n3655) );
  XOR2_X1 U3662 ( .A(n3659), .B(n3660), .Z(n3541) );
  NAND2_X1 U3663 ( .A1(n3661), .A2(n3662), .ZN(n3659) );
  XNOR2_X1 U3664 ( .A(n3663), .B(n3664), .ZN(n3545) );
  XOR2_X1 U3665 ( .A(n3665), .B(n3666), .Z(n3663) );
  NOR2_X1 U3666 ( .A1(n2377), .A2(n3527), .ZN(n3666) );
  XOR2_X1 U3667 ( .A(n3667), .B(n3668), .Z(n3477) );
  NAND2_X1 U3668 ( .A1(n3669), .A2(n3670), .ZN(n3667) );
  XNOR2_X1 U3669 ( .A(n3671), .B(n3672), .ZN(n3549) );
  XOR2_X1 U3670 ( .A(n3673), .B(n3674), .Z(n3671) );
  NOR2_X1 U3671 ( .A1(n3527), .A2(n2247), .ZN(n3674) );
  XNOR2_X1 U3672 ( .A(n3675), .B(n3676), .ZN(n3557) );
  XNOR2_X1 U3673 ( .A(n3677), .B(n3678), .ZN(n3675) );
  NOR2_X1 U3674 ( .A1(n3527), .A2(n2230), .ZN(n3678) );
  XOR2_X1 U3675 ( .A(n3679), .B(n3680), .Z(n3560) );
  XOR2_X1 U3676 ( .A(n3681), .B(n3682), .Z(n3679) );
  XNOR2_X1 U3677 ( .A(n3683), .B(n3684), .ZN(n3565) );
  XOR2_X1 U3678 ( .A(n3685), .B(n3686), .Z(n3683) );
  NAND2_X1 U3679 ( .A1(a_2_), .A2(b_3_), .ZN(n3685) );
  XOR2_X1 U3680 ( .A(n3687), .B(n3688), .Z(n3327) );
  XNOR2_X1 U3681 ( .A(n3689), .B(n3690), .ZN(n3688) );
  NAND2_X1 U3682 ( .A1(a_1_), .A2(b_3_), .ZN(n3690) );
  XOR2_X1 U3683 ( .A(n3691), .B(n3692), .Z(n2072) );
  XNOR2_X1 U3684 ( .A(n3693), .B(n3694), .ZN(n3692) );
  NAND2_X1 U3685 ( .A1(a_0_), .A2(b_3_), .ZN(n3694) );
  NAND2_X1 U3686 ( .A1(n3695), .A2(n3696), .ZN(n2189) );
  INV_X1 U3687 ( .A(n3571), .ZN(n3696) );
  NOR2_X1 U3688 ( .A1(n3697), .A2(n3698), .ZN(n3571) );
  INV_X1 U3689 ( .A(n3699), .ZN(n3698) );
  NAND3_X1 U3690 ( .A1(b_3_), .A2(n3700), .A3(a_0_), .ZN(n3699) );
  NAND2_X1 U3691 ( .A1(n3693), .A2(n3691), .ZN(n3700) );
  NOR2_X1 U3692 ( .A1(n3691), .A2(n3693), .ZN(n3697) );
  NOR2_X1 U3693 ( .A1(n3701), .A2(n3702), .ZN(n3693) );
  NOR3_X1 U3694 ( .A1(n3527), .A2(n3703), .A3(n2343), .ZN(n3702) );
  INV_X1 U3695 ( .A(n3704), .ZN(n3703) );
  NAND2_X1 U3696 ( .A1(n3687), .A2(n3689), .ZN(n3704) );
  NOR2_X1 U3697 ( .A1(n3687), .A2(n3689), .ZN(n3701) );
  NOR2_X1 U3698 ( .A1(n3705), .A2(n3706), .ZN(n3689) );
  NOR3_X1 U3699 ( .A1(n3527), .A2(n3707), .A3(n2139), .ZN(n3706) );
  NOR2_X1 U3700 ( .A1(n3684), .A2(n3686), .ZN(n3707) );
  INV_X1 U3701 ( .A(n3708), .ZN(n3705) );
  NAND2_X1 U3702 ( .A1(n3686), .A2(n3684), .ZN(n3708) );
  XNOR2_X1 U3703 ( .A(n3709), .B(n3710), .ZN(n3684) );
  XNOR2_X1 U3704 ( .A(n3711), .B(n3712), .ZN(n3709) );
  NOR2_X1 U3705 ( .A1(n3713), .A2(n3714), .ZN(n3686) );
  NOR2_X1 U3706 ( .A1(n3680), .A2(n3715), .ZN(n3714) );
  NOR2_X1 U3707 ( .A1(n3681), .A2(n3682), .ZN(n3715) );
  INV_X1 U3708 ( .A(n3716), .ZN(n3682) );
  XNOR2_X1 U3709 ( .A(n3717), .B(n3718), .ZN(n3680) );
  XNOR2_X1 U3710 ( .A(n3719), .B(n3720), .ZN(n3717) );
  NOR2_X1 U3711 ( .A1(n3716), .A2(n3721), .ZN(n3713) );
  NAND2_X1 U3712 ( .A1(n3722), .A2(n3723), .ZN(n3716) );
  NAND3_X1 U3713 ( .A1(b_3_), .A2(n3724), .A3(a_4_), .ZN(n3723) );
  NAND2_X1 U3714 ( .A1(n3676), .A2(n3677), .ZN(n3724) );
  INV_X1 U3715 ( .A(n3725), .ZN(n3722) );
  NOR2_X1 U3716 ( .A1(n3676), .A2(n3677), .ZN(n3725) );
  NOR2_X1 U3717 ( .A1(n3726), .A2(n3727), .ZN(n3677) );
  NOR3_X1 U3718 ( .A1(n3527), .A2(n3728), .A3(n2366), .ZN(n3727) );
  NOR2_X1 U3719 ( .A1(n3596), .A2(n3598), .ZN(n3728) );
  INV_X1 U3720 ( .A(n3729), .ZN(n3726) );
  NAND2_X1 U3721 ( .A1(n3596), .A2(n3598), .ZN(n3729) );
  NAND2_X1 U3722 ( .A1(n3730), .A2(n3731), .ZN(n3598) );
  NAND3_X1 U3723 ( .A1(b_3_), .A2(n3732), .A3(a_6_), .ZN(n3731) );
  INV_X1 U3724 ( .A(n3733), .ZN(n3732) );
  NOR2_X1 U3725 ( .A1(n3672), .A2(n3673), .ZN(n3733) );
  NAND2_X1 U3726 ( .A1(n3672), .A2(n3673), .ZN(n3730) );
  NAND2_X1 U3727 ( .A1(n3669), .A2(n3734), .ZN(n3673) );
  NAND2_X1 U3728 ( .A1(n3668), .A2(n3670), .ZN(n3734) );
  NAND2_X1 U3729 ( .A1(n3735), .A2(n3736), .ZN(n3670) );
  NAND2_X1 U3730 ( .A1(a_7_), .A2(b_3_), .ZN(n3736) );
  XNOR2_X1 U3731 ( .A(n3737), .B(n3738), .ZN(n3668) );
  XNOR2_X1 U3732 ( .A(n3739), .B(n3740), .ZN(n3737) );
  INV_X1 U3733 ( .A(n3741), .ZN(n3669) );
  NOR2_X1 U3734 ( .A1(n2626), .A2(n3735), .ZN(n3741) );
  NOR2_X1 U3735 ( .A1(n3742), .A2(n3743), .ZN(n3735) );
  NOR3_X1 U3736 ( .A1(n2377), .A2(n3744), .A3(n3527), .ZN(n3743) );
  NOR2_X1 U3737 ( .A1(n3664), .A2(n3665), .ZN(n3744) );
  INV_X1 U3738 ( .A(n3745), .ZN(n3742) );
  NAND2_X1 U3739 ( .A1(n3664), .A2(n3665), .ZN(n3745) );
  NAND2_X1 U3740 ( .A1(n3661), .A2(n3746), .ZN(n3665) );
  NAND2_X1 U3741 ( .A1(n3660), .A2(n3662), .ZN(n3746) );
  NAND2_X1 U3742 ( .A1(n3747), .A2(n3748), .ZN(n3662) );
  NAND2_X1 U3743 ( .A1(b_3_), .A2(a_9_), .ZN(n3748) );
  INV_X1 U3744 ( .A(n3749), .ZN(n3747) );
  XNOR2_X1 U3745 ( .A(n3750), .B(n3751), .ZN(n3660) );
  XOR2_X1 U3746 ( .A(n3752), .B(n3753), .Z(n3750) );
  NAND2_X1 U3747 ( .A1(a_9_), .A2(n3749), .ZN(n3661) );
  NAND2_X1 U3748 ( .A1(n3621), .A2(n3754), .ZN(n3749) );
  NAND2_X1 U3749 ( .A1(n3620), .A2(n3622), .ZN(n3754) );
  NAND2_X1 U3750 ( .A1(n3755), .A2(n3756), .ZN(n3622) );
  NAND2_X1 U3751 ( .A1(b_3_), .A2(a_10_), .ZN(n3756) );
  XNOR2_X1 U3752 ( .A(n3757), .B(n3758), .ZN(n3620) );
  XNOR2_X1 U3753 ( .A(n3759), .B(n3760), .ZN(n3758) );
  INV_X1 U3754 ( .A(n3761), .ZN(n3621) );
  NOR2_X1 U3755 ( .A1(n2523), .A2(n3755), .ZN(n3761) );
  NOR2_X1 U3756 ( .A1(n3762), .A2(n3763), .ZN(n3755) );
  INV_X1 U3757 ( .A(n3764), .ZN(n3763) );
  NAND3_X1 U3758 ( .A1(a_11_), .A2(n3765), .A3(b_3_), .ZN(n3764) );
  NAND2_X1 U3759 ( .A1(n3630), .A2(n3628), .ZN(n3765) );
  NOR2_X1 U3760 ( .A1(n3628), .A2(n3630), .ZN(n3762) );
  NOR2_X1 U3761 ( .A1(n3766), .A2(n3767), .ZN(n3630) );
  INV_X1 U3762 ( .A(n3768), .ZN(n3767) );
  NAND2_X1 U3763 ( .A1(n3657), .A2(n3769), .ZN(n3768) );
  NAND2_X1 U3764 ( .A1(n3658), .A2(n3656), .ZN(n3769) );
  NOR2_X1 U3765 ( .A1(n3527), .A2(n2094), .ZN(n3657) );
  NOR2_X1 U3766 ( .A1(n3656), .A2(n3658), .ZN(n3766) );
  NOR2_X1 U3767 ( .A1(n3770), .A2(n3771), .ZN(n3658) );
  INV_X1 U3768 ( .A(n3772), .ZN(n3771) );
  NAND2_X1 U3769 ( .A1(n3652), .A2(n3773), .ZN(n3772) );
  NAND2_X1 U3770 ( .A1(n3653), .A2(n3654), .ZN(n3773) );
  NOR2_X1 U3771 ( .A1(n3527), .A2(n2408), .ZN(n3652) );
  NOR2_X1 U3772 ( .A1(n3654), .A2(n3653), .ZN(n3770) );
  INV_X1 U3773 ( .A(n3774), .ZN(n3653) );
  NAND2_X1 U3774 ( .A1(n3775), .A2(n3776), .ZN(n3774) );
  NAND2_X1 U3775 ( .A1(b_1_), .A2(n3777), .ZN(n3776) );
  NAND2_X1 U3776 ( .A1(n2077), .A2(n3778), .ZN(n3777) );
  NAND2_X1 U3777 ( .A1(a_15_), .A2(n3650), .ZN(n3778) );
  NAND2_X1 U3778 ( .A1(b_2_), .A2(n3779), .ZN(n3775) );
  NAND2_X1 U3779 ( .A1(n2081), .A2(n3780), .ZN(n3779) );
  NAND2_X1 U3780 ( .A1(a_14_), .A2(n3781), .ZN(n3780) );
  NAND3_X1 U3781 ( .A1(b_3_), .A2(n2417), .A3(b_2_), .ZN(n3654) );
  XNOR2_X1 U3782 ( .A(n3782), .B(n3783), .ZN(n3656) );
  XOR2_X1 U3783 ( .A(n3784), .B(n3785), .Z(n3782) );
  XNOR2_X1 U3784 ( .A(n3786), .B(n3787), .ZN(n3628) );
  XOR2_X1 U3785 ( .A(n3788), .B(n3789), .Z(n3786) );
  XNOR2_X1 U3786 ( .A(n3790), .B(n3791), .ZN(n3664) );
  XNOR2_X1 U3787 ( .A(n3792), .B(n3793), .ZN(n3790) );
  XNOR2_X1 U3788 ( .A(n3794), .B(n3795), .ZN(n3672) );
  XNOR2_X1 U3789 ( .A(n3796), .B(n3797), .ZN(n3794) );
  XNOR2_X1 U3790 ( .A(n3798), .B(n3799), .ZN(n3596) );
  XNOR2_X1 U3791 ( .A(n3800), .B(n3801), .ZN(n3798) );
  XOR2_X1 U3792 ( .A(n3802), .B(n3803), .Z(n3676) );
  XNOR2_X1 U3793 ( .A(n3804), .B(n3805), .ZN(n3802) );
  XNOR2_X1 U3794 ( .A(n3806), .B(n3807), .ZN(n3687) );
  XNOR2_X1 U3795 ( .A(n3808), .B(n3809), .ZN(n3807) );
  XOR2_X1 U3796 ( .A(n3810), .B(n3811), .Z(n3691) );
  XNOR2_X1 U3797 ( .A(n3812), .B(n3813), .ZN(n3811) );
  NOR2_X1 U3798 ( .A1(n3650), .A2(n2343), .ZN(n3813) );
  XNOR2_X1 U3799 ( .A(n3573), .B(n3574), .ZN(n3695) );
  NAND2_X1 U3800 ( .A1(n3814), .A2(n3815), .ZN(n3573) );
  XOR2_X1 U3801 ( .A(n2179), .B(n2178), .Z(n2085) );
  XOR2_X1 U3802 ( .A(n3816), .B(n3817), .Z(n2178) );
  XNOR2_X1 U3803 ( .A(n2188), .B(n2187), .ZN(n3817) );
  NOR2_X1 U3804 ( .A1(n3818), .A2(n3819), .ZN(n2187) );
  INV_X1 U3805 ( .A(n3820), .ZN(n3819) );
  NAND3_X1 U3806 ( .A1(b_0_), .A2(n3821), .A3(a_2_), .ZN(n3820) );
  NAND2_X1 U3807 ( .A1(n3822), .A2(n3823), .ZN(n3821) );
  NOR2_X1 U3808 ( .A1(n3823), .A2(n3822), .ZN(n3818) );
  NAND2_X1 U3809 ( .A1(a_0_), .A2(b_1_), .ZN(n2188) );
  NAND2_X1 U3810 ( .A1(a_1_), .A2(b_0_), .ZN(n3816) );
  NAND2_X1 U3811 ( .A1(n3814), .A2(n3824), .ZN(n2179) );
  NAND2_X1 U3812 ( .A1(n3574), .A2(n3815), .ZN(n3824) );
  NAND2_X1 U3813 ( .A1(n3825), .A2(n3826), .ZN(n3815) );
  NAND2_X1 U3814 ( .A1(a_0_), .A2(b_2_), .ZN(n3826) );
  XOR2_X1 U3815 ( .A(n3827), .B(n3828), .Z(n3574) );
  NOR2_X1 U3816 ( .A1(n3829), .A2(n2139), .ZN(n3828) );
  XOR2_X1 U3817 ( .A(n3823), .B(n3822), .Z(n3827) );
  NOR2_X1 U3818 ( .A1(n3830), .A2(n3831), .ZN(n3822) );
  NOR3_X1 U3819 ( .A1(n3781), .A2(n3832), .A3(n2139), .ZN(n3831) );
  INV_X1 U3820 ( .A(n3833), .ZN(n3832) );
  NAND2_X1 U3821 ( .A1(n3834), .A2(n3835), .ZN(n3833) );
  NOR2_X1 U3822 ( .A1(n3835), .A2(n3834), .ZN(n3830) );
  INV_X1 U3823 ( .A(n3836), .ZN(n3814) );
  NOR2_X1 U3824 ( .A1(n2212), .A2(n3825), .ZN(n3836) );
  NOR2_X1 U3825 ( .A1(n3837), .A2(n3838), .ZN(n3825) );
  INV_X1 U3826 ( .A(n3839), .ZN(n3838) );
  NAND3_X1 U3827 ( .A1(b_2_), .A2(n3840), .A3(a_1_), .ZN(n3839) );
  NAND2_X1 U3828 ( .A1(n3810), .A2(n3812), .ZN(n3840) );
  NOR2_X1 U3829 ( .A1(n3810), .A2(n3812), .ZN(n3837) );
  NAND2_X1 U3830 ( .A1(n3841), .A2(n3842), .ZN(n3812) );
  NAND2_X1 U3831 ( .A1(n3843), .A2(n3808), .ZN(n3842) );
  INV_X1 U3832 ( .A(n3844), .ZN(n3843) );
  NOR2_X1 U3833 ( .A1(n3806), .A2(n3809), .ZN(n3844) );
  NAND2_X1 U3834 ( .A1(n3809), .A2(n3806), .ZN(n3841) );
  XNOR2_X1 U3835 ( .A(n3845), .B(n3846), .ZN(n3806) );
  NOR2_X1 U3836 ( .A1(n3781), .A2(n2322), .ZN(n3846) );
  XOR2_X1 U3837 ( .A(n3847), .B(n3848), .Z(n3845) );
  NOR2_X1 U3838 ( .A1(n3849), .A2(n3850), .ZN(n3809) );
  INV_X1 U3839 ( .A(n3851), .ZN(n3850) );
  NAND2_X1 U3840 ( .A1(n3712), .A2(n3852), .ZN(n3851) );
  NAND2_X1 U3841 ( .A1(n3711), .A2(n3710), .ZN(n3852) );
  NOR2_X1 U3842 ( .A1(n2322), .A2(n3650), .ZN(n3712) );
  NOR2_X1 U3843 ( .A1(n3710), .A2(n3711), .ZN(n3849) );
  NOR2_X1 U3844 ( .A1(n3853), .A2(n3854), .ZN(n3711) );
  INV_X1 U3845 ( .A(n3855), .ZN(n3854) );
  NAND2_X1 U3846 ( .A1(n3719), .A2(n3856), .ZN(n3855) );
  NAND2_X1 U3847 ( .A1(n3720), .A2(n3718), .ZN(n3856) );
  NOR2_X1 U3848 ( .A1(n2230), .A2(n3650), .ZN(n3719) );
  NOR2_X1 U3849 ( .A1(n3718), .A2(n3720), .ZN(n3853) );
  NOR2_X1 U3850 ( .A1(n3857), .A2(n3858), .ZN(n3720) );
  INV_X1 U3851 ( .A(n3859), .ZN(n3858) );
  NAND2_X1 U3852 ( .A1(n3805), .A2(n3860), .ZN(n3859) );
  NAND2_X1 U3853 ( .A1(n3804), .A2(n3803), .ZN(n3860) );
  NOR2_X1 U3854 ( .A1(n2366), .A2(n3650), .ZN(n3805) );
  NOR2_X1 U3855 ( .A1(n3803), .A2(n3804), .ZN(n3857) );
  NOR2_X1 U3856 ( .A1(n3861), .A2(n3862), .ZN(n3804) );
  INV_X1 U3857 ( .A(n3863), .ZN(n3862) );
  NAND2_X1 U3858 ( .A1(n3800), .A2(n3864), .ZN(n3863) );
  NAND2_X1 U3859 ( .A1(n3801), .A2(n3799), .ZN(n3864) );
  NOR2_X1 U3860 ( .A1(n2247), .A2(n3650), .ZN(n3800) );
  NOR2_X1 U3861 ( .A1(n3799), .A2(n3801), .ZN(n3861) );
  NOR2_X1 U3862 ( .A1(n3865), .A2(n3866), .ZN(n3801) );
  INV_X1 U3863 ( .A(n3867), .ZN(n3866) );
  NAND2_X1 U3864 ( .A1(n3797), .A2(n3868), .ZN(n3867) );
  NAND2_X1 U3865 ( .A1(n3796), .A2(n3795), .ZN(n3868) );
  NOR2_X1 U3866 ( .A1(n2626), .A2(n3650), .ZN(n3797) );
  NOR2_X1 U3867 ( .A1(n3795), .A2(n3796), .ZN(n3865) );
  NOR2_X1 U3868 ( .A1(n3869), .A2(n3870), .ZN(n3796) );
  INV_X1 U3869 ( .A(n3871), .ZN(n3870) );
  NAND2_X1 U3870 ( .A1(n3739), .A2(n3872), .ZN(n3871) );
  NAND2_X1 U3871 ( .A1(n3740), .A2(n3738), .ZN(n3872) );
  NOR2_X1 U3872 ( .A1(n3650), .A2(n2377), .ZN(n3739) );
  NOR2_X1 U3873 ( .A1(n3738), .A2(n3740), .ZN(n3869) );
  NOR2_X1 U3874 ( .A1(n3873), .A2(n3874), .ZN(n3740) );
  INV_X1 U3875 ( .A(n3875), .ZN(n3874) );
  NAND2_X1 U3876 ( .A1(n3793), .A2(n3876), .ZN(n3875) );
  NAND2_X1 U3877 ( .A1(n3792), .A2(n3791), .ZN(n3876) );
  NOR2_X1 U3878 ( .A1(n3650), .A2(n2275), .ZN(n3793) );
  NOR2_X1 U3879 ( .A1(n3791), .A2(n3792), .ZN(n3873) );
  NOR2_X1 U3880 ( .A1(n3877), .A2(n3878), .ZN(n3792) );
  INV_X1 U3881 ( .A(n3879), .ZN(n3878) );
  NAND2_X1 U3882 ( .A1(n3752), .A2(n3880), .ZN(n3879) );
  NAND2_X1 U3883 ( .A1(n3881), .A2(n3751), .ZN(n3880) );
  NOR2_X1 U3884 ( .A1(n3650), .A2(n2523), .ZN(n3752) );
  NOR2_X1 U3885 ( .A1(n3751), .A2(n3881), .ZN(n3877) );
  INV_X1 U3886 ( .A(n3753), .ZN(n3881) );
  NAND2_X1 U3887 ( .A1(n3882), .A2(n3883), .ZN(n3753) );
  NAND2_X1 U3888 ( .A1(n3760), .A2(n3884), .ZN(n3883) );
  INV_X1 U3889 ( .A(n3885), .ZN(n3884) );
  NOR2_X1 U3890 ( .A1(n3759), .A2(n3757), .ZN(n3885) );
  NOR2_X1 U3891 ( .A1(n3650), .A2(n2284), .ZN(n3760) );
  NAND2_X1 U3892 ( .A1(n3757), .A2(n3759), .ZN(n3882) );
  NAND2_X1 U3893 ( .A1(n3886), .A2(n3887), .ZN(n3759) );
  NAND2_X1 U3894 ( .A1(n3788), .A2(n3888), .ZN(n3887) );
  INV_X1 U3895 ( .A(n3889), .ZN(n3888) );
  NOR2_X1 U3896 ( .A1(n3787), .A2(n3789), .ZN(n3889) );
  NOR2_X1 U3897 ( .A1(n3650), .A2(n2094), .ZN(n3788) );
  NAND2_X1 U3898 ( .A1(n3787), .A2(n3789), .ZN(n3886) );
  NAND2_X1 U3899 ( .A1(n3890), .A2(n3891), .ZN(n3789) );
  NAND2_X1 U3900 ( .A1(n3783), .A2(n3892), .ZN(n3891) );
  INV_X1 U3901 ( .A(n3893), .ZN(n3892) );
  NOR2_X1 U3902 ( .A1(n3784), .A2(n3785), .ZN(n3893) );
  NOR2_X1 U3903 ( .A1(n3650), .A2(n2408), .ZN(n3783) );
  NAND2_X1 U3904 ( .A1(n3785), .A2(n3784), .ZN(n3890) );
  NAND2_X1 U3905 ( .A1(n3894), .A2(n3895), .ZN(n3784) );
  NAND2_X1 U3906 ( .A1(b_0_), .A2(n3896), .ZN(n3895) );
  NAND2_X1 U3907 ( .A1(n2077), .A2(n3897), .ZN(n3896) );
  NAND2_X1 U3908 ( .A1(a_15_), .A2(n3781), .ZN(n3897) );
  NAND2_X1 U3909 ( .A1(a_15_), .A2(n3898), .ZN(n2077) );
  NAND2_X1 U3910 ( .A1(b_1_), .A2(n3899), .ZN(n3894) );
  NAND2_X1 U3911 ( .A1(n2081), .A2(n3900), .ZN(n3899) );
  NAND2_X1 U3912 ( .A1(a_14_), .A2(n3829), .ZN(n3900) );
  NAND2_X1 U3913 ( .A1(a_14_), .A2(n3901), .ZN(n2081) );
  INV_X1 U3914 ( .A(a_15_), .ZN(n3901) );
  NOR3_X1 U3915 ( .A1(n3650), .A2(n2675), .A3(n3781), .ZN(n3785) );
  XNOR2_X1 U3916 ( .A(n3902), .B(n3903), .ZN(n3787) );
  XNOR2_X1 U3917 ( .A(n3904), .B(n3905), .ZN(n3903) );
  NAND2_X1 U3918 ( .A1(b_0_), .A2(a_14_), .ZN(n3902) );
  XNOR2_X1 U3919 ( .A(n3906), .B(n3907), .ZN(n3757) );
  NAND2_X1 U3920 ( .A1(n3908), .A2(n3909), .ZN(n3906) );
  NAND2_X1 U3921 ( .A1(n3910), .A2(n3911), .ZN(n3909) );
  NAND2_X1 U3922 ( .A1(b_1_), .A2(a_12_), .ZN(n3910) );
  XNOR2_X1 U3923 ( .A(n3912), .B(n3913), .ZN(n3751) );
  XOR2_X1 U3924 ( .A(n3914), .B(n3915), .Z(n3913) );
  NAND2_X1 U3925 ( .A1(b_1_), .A2(a_11_), .ZN(n3912) );
  XNOR2_X1 U3926 ( .A(n3916), .B(n3917), .ZN(n3791) );
  XNOR2_X1 U3927 ( .A(n3918), .B(n3919), .ZN(n3917) );
  NAND2_X1 U3928 ( .A1(b_1_), .A2(a_10_), .ZN(n3916) );
  XNOR2_X1 U3929 ( .A(n3920), .B(n3921), .ZN(n3738) );
  NOR2_X1 U3930 ( .A1(n2275), .A2(n3781), .ZN(n3921) );
  XOR2_X1 U3931 ( .A(n3922), .B(n3923), .Z(n3920) );
  XNOR2_X1 U3932 ( .A(n3924), .B(n3925), .ZN(n3795) );
  XNOR2_X1 U3933 ( .A(n3926), .B(n3927), .ZN(n3925) );
  NAND2_X1 U3934 ( .A1(b_1_), .A2(a_8_), .ZN(n3924) );
  XNOR2_X1 U3935 ( .A(n3928), .B(n3929), .ZN(n3799) );
  NOR2_X1 U3936 ( .A1(n3781), .A2(n2626), .ZN(n3929) );
  XOR2_X1 U3937 ( .A(n3930), .B(n3931), .Z(n3928) );
  XNOR2_X1 U3938 ( .A(n3932), .B(n3933), .ZN(n3803) );
  XNOR2_X1 U3939 ( .A(n3934), .B(n3935), .ZN(n3933) );
  NAND2_X1 U3940 ( .A1(a_6_), .A2(b_1_), .ZN(n3932) );
  XNOR2_X1 U3941 ( .A(n3936), .B(n3937), .ZN(n3718) );
  NOR2_X1 U3942 ( .A1(n3781), .A2(n2366), .ZN(n3937) );
  XOR2_X1 U3943 ( .A(n3938), .B(n3939), .Z(n3936) );
  XNOR2_X1 U3944 ( .A(n3940), .B(n3941), .ZN(n3710) );
  XNOR2_X1 U3945 ( .A(n3942), .B(n3943), .ZN(n3941) );
  NAND2_X1 U3946 ( .A1(a_4_), .A2(b_1_), .ZN(n3940) );
  XNOR2_X1 U3947 ( .A(n3944), .B(n3945), .ZN(n3810) );
  XNOR2_X1 U3948 ( .A(n3835), .B(n3834), .ZN(n3945) );
  NOR2_X1 U3949 ( .A1(n3946), .A2(n3947), .ZN(n3834) );
  NOR3_X1 U3950 ( .A1(n3781), .A2(n3948), .A3(n2322), .ZN(n3947) );
  INV_X1 U3951 ( .A(n3949), .ZN(n3948) );
  NAND2_X1 U3952 ( .A1(n3848), .A2(n3847), .ZN(n3949) );
  NOR2_X1 U3953 ( .A1(n3847), .A2(n3848), .ZN(n3946) );
  NOR2_X1 U3954 ( .A1(n3950), .A2(n3951), .ZN(n3848) );
  INV_X1 U3955 ( .A(n3952), .ZN(n3951) );
  NAND3_X1 U3956 ( .A1(b_1_), .A2(n3953), .A3(a_4_), .ZN(n3952) );
  NAND2_X1 U3957 ( .A1(n3943), .A2(n3942), .ZN(n3953) );
  NOR2_X1 U3958 ( .A1(n3942), .A2(n3943), .ZN(n3950) );
  NOR2_X1 U3959 ( .A1(n3954), .A2(n3955), .ZN(n3943) );
  NOR3_X1 U3960 ( .A1(n3781), .A2(n3956), .A3(n2366), .ZN(n3955) );
  INV_X1 U3961 ( .A(n3957), .ZN(n3956) );
  NAND2_X1 U3962 ( .A1(n3939), .A2(n3938), .ZN(n3957) );
  NOR2_X1 U3963 ( .A1(n3938), .A2(n3939), .ZN(n3954) );
  NOR2_X1 U3964 ( .A1(n3958), .A2(n3959), .ZN(n3939) );
  INV_X1 U3965 ( .A(n3960), .ZN(n3959) );
  NAND3_X1 U3966 ( .A1(b_1_), .A2(n3961), .A3(a_6_), .ZN(n3960) );
  NAND2_X1 U3967 ( .A1(n3935), .A2(n3934), .ZN(n3961) );
  NOR2_X1 U3968 ( .A1(n3934), .A2(n3935), .ZN(n3958) );
  NOR2_X1 U3969 ( .A1(n3962), .A2(n3963), .ZN(n3935) );
  NOR3_X1 U3970 ( .A1(n3781), .A2(n3964), .A3(n2626), .ZN(n3963) );
  INV_X1 U3971 ( .A(n3965), .ZN(n3964) );
  NAND2_X1 U3972 ( .A1(n3931), .A2(n3930), .ZN(n3965) );
  NOR2_X1 U3973 ( .A1(n3930), .A2(n3931), .ZN(n3962) );
  NOR2_X1 U3974 ( .A1(n3966), .A2(n3967), .ZN(n3931) );
  INV_X1 U3975 ( .A(n3968), .ZN(n3967) );
  NAND3_X1 U3976 ( .A1(a_8_), .A2(n3969), .A3(b_1_), .ZN(n3968) );
  NAND2_X1 U3977 ( .A1(n3927), .A2(n3926), .ZN(n3969) );
  NOR2_X1 U3978 ( .A1(n3926), .A2(n3927), .ZN(n3966) );
  NOR2_X1 U3979 ( .A1(n3970), .A2(n3971), .ZN(n3927) );
  NOR3_X1 U3980 ( .A1(n2275), .A2(n3972), .A3(n3781), .ZN(n3971) );
  INV_X1 U3981 ( .A(n3973), .ZN(n3972) );
  NAND2_X1 U3982 ( .A1(n3923), .A2(n3922), .ZN(n3973) );
  NOR2_X1 U3983 ( .A1(n3922), .A2(n3923), .ZN(n3970) );
  NOR2_X1 U3984 ( .A1(n3974), .A2(n3975), .ZN(n3923) );
  NOR3_X1 U3985 ( .A1(n2523), .A2(n3976), .A3(n3781), .ZN(n3975) );
  NOR2_X1 U3986 ( .A1(n3919), .A2(n3918), .ZN(n3976) );
  INV_X1 U3987 ( .A(n3977), .ZN(n3974) );
  NAND2_X1 U3988 ( .A1(n3918), .A2(n3919), .ZN(n3977) );
  NAND2_X1 U3989 ( .A1(n3978), .A2(n3979), .ZN(n3919) );
  NAND3_X1 U3990 ( .A1(a_11_), .A2(n3980), .A3(b_1_), .ZN(n3979) );
  NAND2_X1 U3991 ( .A1(n3915), .A2(n3981), .ZN(n3980) );
  INV_X1 U3992 ( .A(n3982), .ZN(n3915) );
  NAND2_X1 U3993 ( .A1(n3914), .A2(n3982), .ZN(n3978) );
  NAND2_X1 U3994 ( .A1(n3908), .A2(n3983), .ZN(n3982) );
  NAND2_X1 U3995 ( .A1(n3984), .A2(n3907), .ZN(n3983) );
  NAND2_X1 U3996 ( .A1(n3905), .A2(n3985), .ZN(n3907) );
  NAND3_X1 U3997 ( .A1(b_0_), .A2(a_14_), .A3(n3904), .ZN(n3985) );
  NOR2_X1 U3998 ( .A1(n3781), .A2(n2408), .ZN(n3904) );
  NAND3_X1 U3999 ( .A1(b_1_), .A2(n2417), .A3(b_0_), .ZN(n3905) );
  INV_X1 U4000 ( .A(n2675), .ZN(n2417) );
  NAND2_X1 U4001 ( .A1(a_15_), .A2(a_14_), .ZN(n2675) );
  NAND2_X1 U4002 ( .A1(n3911), .A2(n2094), .ZN(n3984) );
  INV_X1 U4003 ( .A(n3986), .ZN(n3911) );
  NAND3_X1 U4004 ( .A1(b_1_), .A2(a_12_), .A3(n3986), .ZN(n3908) );
  NOR2_X1 U4005 ( .A1(n3829), .A2(n2408), .ZN(n3986) );
  INV_X1 U4006 ( .A(n3981), .ZN(n3914) );
  NAND2_X1 U4007 ( .A1(b_0_), .A2(a_12_), .ZN(n3981) );
  NOR2_X1 U4008 ( .A1(n3829), .A2(n2284), .ZN(n3918) );
  NAND2_X1 U4009 ( .A1(b_0_), .A2(a_10_), .ZN(n3922) );
  NAND2_X1 U4010 ( .A1(b_0_), .A2(a_9_), .ZN(n3926) );
  NAND2_X1 U4011 ( .A1(b_0_), .A2(a_8_), .ZN(n3930) );
  NAND2_X1 U4012 ( .A1(b_0_), .A2(a_7_), .ZN(n3934) );
  NAND2_X1 U4013 ( .A1(a_6_), .A2(b_0_), .ZN(n3938) );
  NAND2_X1 U4014 ( .A1(a_5_), .A2(b_0_), .ZN(n3942) );
  NAND2_X1 U4015 ( .A1(a_4_), .A2(b_0_), .ZN(n3847) );
  NAND2_X1 U4016 ( .A1(a_3_), .A2(b_0_), .ZN(n3835) );
  NAND2_X1 U4017 ( .A1(a_2_), .A2(b_1_), .ZN(n3944) );
  NAND3_X1 U4018 ( .A1(n3987), .A2(n3988), .A3(n3989), .ZN(Result_add_9_) );
  NAND2_X1 U4019 ( .A1(n2928), .A2(n3990), .ZN(n3989) );
  INV_X1 U4020 ( .A(n3016), .ZN(n2928) );
  NAND3_X1 U4021 ( .A1(n3991), .A2(n2275), .A3(b_9_), .ZN(n3988) );
  NAND2_X1 U4022 ( .A1(n3992), .A2(n2793), .ZN(n3987) );
  XOR2_X1 U4023 ( .A(n3991), .B(n2275), .Z(n3992) );
  INV_X1 U4024 ( .A(n3990), .ZN(n3991) );
  XNOR2_X1 U4025 ( .A(n3993), .B(n3994), .ZN(Result_add_8_) );
  NAND2_X1 U4026 ( .A1(n3995), .A2(n3055), .ZN(n3994) );
  NAND3_X1 U4027 ( .A1(n3996), .A2(n3997), .A3(n3998), .ZN(Result_add_7_) );
  INV_X1 U4028 ( .A(n3999), .ZN(n3998) );
  NOR2_X1 U4029 ( .A1(n3188), .A2(n4000), .ZN(n3999) );
  NAND3_X1 U4030 ( .A1(n4000), .A2(n2626), .A3(b_7_), .ZN(n3997) );
  NAND2_X1 U4031 ( .A1(n4001), .A2(n3044), .ZN(n3996) );
  XOR2_X1 U4032 ( .A(n4000), .B(n2626), .Z(n4001) );
  INV_X1 U4033 ( .A(n4002), .ZN(n4000) );
  XNOR2_X1 U4034 ( .A(n4003), .B(n4004), .ZN(Result_add_6_) );
  NAND2_X1 U4035 ( .A1(n4005), .A2(n3301), .ZN(n4004) );
  NAND3_X1 U4036 ( .A1(n4006), .A2(n4007), .A3(n4008), .ZN(Result_add_5_) );
  NAND2_X1 U4037 ( .A1(n4009), .A2(n4010), .ZN(n4008) );
  INV_X1 U4038 ( .A(n3429), .ZN(n4009) );
  NAND3_X1 U4039 ( .A1(n4011), .A2(n2366), .A3(b_5_), .ZN(n4007) );
  INV_X1 U4040 ( .A(n4010), .ZN(n4011) );
  NAND2_X1 U4041 ( .A1(n4012), .A2(n3285), .ZN(n4006) );
  XOR2_X1 U4042 ( .A(n4010), .B(a_5_), .Z(n4012) );
  XNOR2_X1 U4043 ( .A(n4013), .B(n4014), .ZN(Result_add_4_) );
  NOR2_X1 U4044 ( .A1(n4015), .A2(n3555), .ZN(n4014) );
  NAND3_X1 U4045 ( .A1(n4016), .A2(n4017), .A3(n4018), .ZN(Result_add_3_) );
  NAND2_X1 U4046 ( .A1(n3721), .A2(n4019), .ZN(n4018) );
  INV_X1 U4047 ( .A(n3681), .ZN(n3721) );
  NAND3_X1 U4048 ( .A1(n4020), .A2(n2322), .A3(b_3_), .ZN(n4017) );
  NAND2_X1 U4049 ( .A1(n4021), .A2(n3527), .ZN(n4016) );
  XOR2_X1 U4050 ( .A(n4019), .B(a_3_), .Z(n4021) );
  XNOR2_X1 U4051 ( .A(n4022), .B(n4023), .ZN(Result_add_2_) );
  NAND2_X1 U4052 ( .A1(n4024), .A2(n3808), .ZN(n4023) );
  NAND2_X1 U4053 ( .A1(n4025), .A2(n4026), .ZN(Result_add_1_) );
  NAND2_X1 U4054 ( .A1(n4027), .A2(n4028), .ZN(n4026) );
  NAND2_X1 U4055 ( .A1(n3823), .A2(n4029), .ZN(n4027) );
  NAND2_X1 U4056 ( .A1(n4030), .A2(n4031), .ZN(n4025) );
  XOR2_X1 U4057 ( .A(b_1_), .B(a_1_), .Z(n4030) );
  XOR2_X1 U4058 ( .A(b_15_), .B(a_15_), .Z(Result_add_15_) );
  NAND3_X1 U4059 ( .A1(n4032), .A2(n4033), .A3(n2086), .ZN(Result_add_14_) );
  NAND3_X1 U4060 ( .A1(b_14_), .A2(a_14_), .A3(Result_mul_31_), .ZN(n2086) );
  NAND2_X1 U4061 ( .A1(n4034), .A2(n2083), .ZN(n4033) );
  INV_X1 U4062 ( .A(b_14_), .ZN(n2083) );
  XOR2_X1 U4063 ( .A(n3898), .B(n4035), .Z(n4034) );
  NAND3_X1 U4064 ( .A1(n4035), .A2(n3898), .A3(b_14_), .ZN(n4032) );
  NAND3_X1 U4065 ( .A1(n4036), .A2(n4037), .A3(n4038), .ZN(Result_add_13_) );
  NAND2_X1 U4066 ( .A1(n2419), .A2(n4039), .ZN(n4038) );
  NAND3_X1 U4067 ( .A1(n4040), .A2(n2408), .A3(b_13_), .ZN(n4037) );
  NAND2_X1 U4068 ( .A1(n4041), .A2(n2305), .ZN(n4036) );
  XOR2_X1 U4069 ( .A(n4040), .B(n2408), .Z(n4041) );
  XNOR2_X1 U4070 ( .A(n4042), .B(n4043), .ZN(Result_add_12_) );
  NOR2_X1 U4071 ( .A1(n4044), .A2(n2549), .ZN(n4043) );
  NAND3_X1 U4072 ( .A1(n4045), .A2(n4046), .A3(n4047), .ZN(Result_add_11_) );
  NAND2_X1 U4073 ( .A1(n4048), .A2(n4049), .ZN(n4047) );
  INV_X1 U4074 ( .A(n2645), .ZN(n4048) );
  NAND3_X1 U4075 ( .A1(n4050), .A2(n2284), .A3(b_11_), .ZN(n4046) );
  NAND2_X1 U4076 ( .A1(n4051), .A2(n2542), .ZN(n4045) );
  XOR2_X1 U4077 ( .A(n4049), .B(a_11_), .Z(n4051) );
  XNOR2_X1 U4078 ( .A(n4052), .B(n4053), .ZN(Result_add_10_) );
  NAND2_X1 U4079 ( .A1(n4054), .A2(n2761), .ZN(n4053) );
  XNOR2_X1 U4080 ( .A(n4055), .B(n4056), .ZN(Result_add_0_) );
  NOR2_X1 U4081 ( .A1(n4057), .A2(n2177), .ZN(n4056) );
  NOR2_X1 U4082 ( .A1(n2212), .A2(n3829), .ZN(n2177) );
  INV_X1 U4083 ( .A(b_0_), .ZN(n3829) );
  INV_X1 U4084 ( .A(a_0_), .ZN(n2212) );
  NOR2_X1 U4085 ( .A1(b_0_), .A2(a_0_), .ZN(n4057) );
  NAND2_X1 U4086 ( .A1(n4029), .A2(n4058), .ZN(n4055) );
  NAND2_X1 U4087 ( .A1(n3823), .A2(n4031), .ZN(n4058) );
  INV_X1 U4088 ( .A(n4028), .ZN(n4031) );
  NAND2_X1 U4089 ( .A1(n3808), .A2(n4059), .ZN(n4028) );
  NAND2_X1 U4090 ( .A1(n4024), .A2(n4022), .ZN(n4059) );
  NAND2_X1 U4091 ( .A1(n3681), .A2(n4060), .ZN(n4022) );
  NAND2_X1 U4092 ( .A1(n4061), .A2(n4019), .ZN(n4060) );
  INV_X1 U4093 ( .A(n4020), .ZN(n4019) );
  NOR2_X1 U4094 ( .A1(n3555), .A2(n4062), .ZN(n4020) );
  NOR2_X1 U4095 ( .A1(n4015), .A2(n4013), .ZN(n4062) );
  INV_X1 U4096 ( .A(n4063), .ZN(n4013) );
  NAND2_X1 U4097 ( .A1(n3429), .A2(n4064), .ZN(n4063) );
  NAND2_X1 U4098 ( .A1(n4065), .A2(n4010), .ZN(n4064) );
  NAND2_X1 U4099 ( .A1(n3301), .A2(n4066), .ZN(n4010) );
  NAND2_X1 U4100 ( .A1(n4005), .A2(n4003), .ZN(n4066) );
  NAND2_X1 U4101 ( .A1(n3188), .A2(n4067), .ZN(n4003) );
  NAND2_X1 U4102 ( .A1(n4068), .A2(n4002), .ZN(n4067) );
  NAND2_X1 U4103 ( .A1(n3055), .A2(n4069), .ZN(n4002) );
  NAND2_X1 U4104 ( .A1(n3995), .A2(n3993), .ZN(n4069) );
  NAND2_X1 U4105 ( .A1(n3016), .A2(n4070), .ZN(n3993) );
  NAND2_X1 U4106 ( .A1(n4071), .A2(n3990), .ZN(n4070) );
  NAND2_X1 U4107 ( .A1(n2761), .A2(n4072), .ZN(n3990) );
  NAND2_X1 U4108 ( .A1(n4054), .A2(n4052), .ZN(n4072) );
  NAND2_X1 U4109 ( .A1(n2645), .A2(n4073), .ZN(n4052) );
  NAND2_X1 U4110 ( .A1(n4074), .A2(n4049), .ZN(n4073) );
  INV_X1 U4111 ( .A(n4050), .ZN(n4049) );
  NOR2_X1 U4112 ( .A1(n2549), .A2(n4075), .ZN(n4050) );
  NOR2_X1 U4113 ( .A1(n4044), .A2(n4042), .ZN(n4075) );
  NOR2_X1 U4114 ( .A1(n2419), .A2(n4076), .ZN(n4042) );
  NOR2_X1 U4115 ( .A1(n4077), .A2(n4040), .ZN(n4076) );
  INV_X1 U4116 ( .A(n4039), .ZN(n4040) );
  NAND2_X1 U4117 ( .A1(n4078), .A2(n4079), .ZN(n4039) );
  NAND2_X1 U4118 ( .A1(b_14_), .A2(n4080), .ZN(n4079) );
  NAND2_X1 U4119 ( .A1(n3898), .A2(n4035), .ZN(n4080) );
  INV_X1 U4120 ( .A(a_14_), .ZN(n3898) );
  NAND2_X1 U4121 ( .A1(Result_mul_31_), .A2(a_14_), .ZN(n4078) );
  INV_X1 U4122 ( .A(n4035), .ZN(Result_mul_31_) );
  NAND2_X1 U4123 ( .A1(b_15_), .A2(a_15_), .ZN(n4035) );
  NOR2_X1 U4124 ( .A1(b_13_), .A2(a_13_), .ZN(n4077) );
  NOR2_X1 U4125 ( .A1(n2305), .A2(n2408), .ZN(n2419) );
  INV_X1 U4126 ( .A(a_13_), .ZN(n2408) );
  INV_X1 U4127 ( .A(b_13_), .ZN(n2305) );
  NOR2_X1 U4128 ( .A1(b_12_), .A2(a_12_), .ZN(n4044) );
  NOR2_X1 U4129 ( .A1(n2416), .A2(n2094), .ZN(n2549) );
  INV_X1 U4130 ( .A(a_12_), .ZN(n2094) );
  INV_X1 U4131 ( .A(b_12_), .ZN(n2416) );
  NAND2_X1 U4132 ( .A1(n2542), .A2(n2284), .ZN(n4074) );
  INV_X1 U4133 ( .A(a_11_), .ZN(n2284) );
  INV_X1 U4134 ( .A(b_11_), .ZN(n2542) );
  NAND2_X1 U4135 ( .A1(b_11_), .A2(a_11_), .ZN(n2645) );
  NAND2_X1 U4136 ( .A1(n2674), .A2(n2523), .ZN(n4054) );
  INV_X1 U4137 ( .A(a_10_), .ZN(n2523) );
  INV_X1 U4138 ( .A(b_10_), .ZN(n2674) );
  NAND2_X1 U4139 ( .A1(b_10_), .A2(a_10_), .ZN(n2761) );
  NAND2_X1 U4140 ( .A1(n2793), .A2(n2275), .ZN(n4071) );
  INV_X1 U4141 ( .A(a_9_), .ZN(n2275) );
  INV_X1 U4142 ( .A(b_9_), .ZN(n2793) );
  NAND2_X1 U4143 ( .A1(a_9_), .A2(b_9_), .ZN(n3016) );
  NAND2_X1 U4144 ( .A1(n2916), .A2(n2377), .ZN(n3995) );
  INV_X1 U4145 ( .A(a_8_), .ZN(n2377) );
  INV_X1 U4146 ( .A(b_8_), .ZN(n2916) );
  NAND2_X1 U4147 ( .A1(b_8_), .A2(a_8_), .ZN(n3055) );
  NAND2_X1 U4148 ( .A1(n3044), .A2(n2626), .ZN(n4068) );
  INV_X1 U4149 ( .A(a_7_), .ZN(n2626) );
  INV_X1 U4150 ( .A(b_7_), .ZN(n3044) );
  NAND2_X1 U4151 ( .A1(a_7_), .A2(b_7_), .ZN(n3188) );
  NAND2_X1 U4152 ( .A1(n3176), .A2(n2247), .ZN(n4005) );
  INV_X1 U4153 ( .A(a_6_), .ZN(n2247) );
  INV_X1 U4154 ( .A(b_6_), .ZN(n3176) );
  NAND2_X1 U4155 ( .A1(a_6_), .A2(b_6_), .ZN(n3301) );
  NAND2_X1 U4156 ( .A1(n3285), .A2(n2366), .ZN(n4065) );
  INV_X1 U4157 ( .A(a_5_), .ZN(n2366) );
  INV_X1 U4158 ( .A(b_5_), .ZN(n3285) );
  NAND2_X1 U4159 ( .A1(a_5_), .A2(b_5_), .ZN(n3429) );
  NOR2_X1 U4160 ( .A1(b_4_), .A2(a_4_), .ZN(n4015) );
  NOR2_X1 U4161 ( .A1(n2230), .A2(n3401), .ZN(n3555) );
  INV_X1 U4162 ( .A(b_4_), .ZN(n3401) );
  INV_X1 U4163 ( .A(a_4_), .ZN(n2230) );
  NAND2_X1 U4164 ( .A1(n3527), .A2(n2322), .ZN(n4061) );
  INV_X1 U4165 ( .A(a_3_), .ZN(n2322) );
  INV_X1 U4166 ( .A(b_3_), .ZN(n3527) );
  NAND2_X1 U4167 ( .A1(a_3_), .A2(b_3_), .ZN(n3681) );
  NAND2_X1 U4168 ( .A1(n3650), .A2(n2139), .ZN(n4024) );
  INV_X1 U4169 ( .A(a_2_), .ZN(n2139) );
  INV_X1 U4170 ( .A(b_2_), .ZN(n3650) );
  NAND2_X1 U4171 ( .A1(a_2_), .A2(b_2_), .ZN(n3808) );
  NAND2_X1 U4172 ( .A1(a_1_), .A2(b_1_), .ZN(n3823) );
  NAND2_X1 U4173 ( .A1(n3781), .A2(n2343), .ZN(n4029) );
  INV_X1 U4174 ( .A(a_1_), .ZN(n2343) );
  INV_X1 U4175 ( .A(b_1_), .ZN(n3781) );
endmodule

