module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n641_, new_n339_, new_n365_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n170_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n716_, new_n153_, new_n701_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n496_, new_n498_, new_n650_, new_n708_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n632_, new_n671_, new_n528_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n717_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n662_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n711_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n573_, new_n405_;

not g000 ( new_n151_, keyIn_0_3 );
nand g001 ( new_n152_, N29, N42, N75 );
nand g002 ( new_n153_, new_n152_, new_n151_ );
nand g003 ( new_n154_, keyIn_0_3, N29, N42, N75 );
nand g004 ( N388, new_n153_, new_n154_ );
nand g005 ( new_n156_, N29, N36, N80 );
not g006 ( N389, new_n156_ );
not g007 ( new_n158_, keyIn_0_4 );
nand g008 ( new_n159_, N29, N36, N42 );
not g009 ( new_n160_, new_n159_ );
nand g010 ( new_n161_, new_n160_, new_n158_ );
nand g011 ( new_n162_, new_n159_, keyIn_0_4 );
nand g012 ( N390, new_n161_, new_n162_ );
nand g013 ( new_n164_, N85, N86 );
not g014 ( N391, new_n164_ );
nand g015 ( new_n166_, N1, N8 );
not g016 ( new_n167_, new_n166_ );
nand g017 ( new_n168_, new_n167_, N13, N17 );
nand g018 ( new_n169_, new_n168_, keyIn_0_0 );
not g019 ( new_n170_, keyIn_0_0 );
nand g020 ( new_n171_, new_n167_, new_n170_, N13, N17 );
nand g021 ( N418, new_n169_, new_n171_ );
nand g022 ( new_n173_, N1, N26 );
nand g023 ( new_n174_, N13, N17 );
nor g024 ( new_n175_, new_n173_, new_n174_ );
nand g025 ( new_n176_, new_n160_, keyIn_0_1 );
not g026 ( new_n177_, keyIn_0_1 );
nand g027 ( new_n178_, new_n159_, new_n177_ );
nand g028 ( N419, new_n176_, new_n175_, new_n178_ );
nand g029 ( N420, N59, N75, N80 );
nand g030 ( N421, N36, N59, N80 );
not g031 ( new_n182_, keyIn_0_5 );
nand g032 ( new_n183_, N36, N42, N59 );
nand g033 ( new_n184_, new_n183_, new_n182_ );
nand g034 ( new_n185_, keyIn_0_5, N36, N42, N59 );
nand g035 ( N422, new_n184_, new_n185_ );
not g036 ( new_n187_, N90 );
nor g037 ( new_n188_, N87, N88 );
nor g038 ( N423, new_n188_, new_n187_ );
nand g039 ( new_n190_, new_n176_, new_n178_ );
nand g040 ( N446, new_n190_, new_n175_ );
not g041 ( new_n192_, keyIn_0_2 );
nand g042 ( new_n193_, N1, N26, N51 );
nand g043 ( new_n194_, new_n193_, new_n192_ );
nand g044 ( new_n195_, keyIn_0_2, N1, N26, N51 );
nand g045 ( new_n196_, new_n194_, new_n195_ );
not g046 ( N447, new_n196_ );
nand g047 ( new_n198_, new_n167_, N13, N55 );
nand g048 ( new_n199_, N29, N68 );
nor g049 ( N448, new_n198_, new_n199_ );
not g050 ( new_n201_, keyIn_0_12 );
not g051 ( new_n202_, new_n198_ );
nand g052 ( new_n203_, N59, N68 );
not g053 ( new_n204_, new_n203_ );
nand g054 ( new_n205_, new_n202_, N74, new_n204_ );
nand g055 ( new_n206_, new_n205_, new_n201_ );
nand g056 ( new_n207_, new_n202_, keyIn_0_12, N74, new_n204_ );
nand g057 ( N449, new_n206_, new_n207_ );
not g058 ( new_n209_, keyIn_0_9 );
not g059 ( new_n210_, new_n188_ );
nand g060 ( new_n211_, new_n210_, N89 );
nand g061 ( new_n212_, new_n211_, new_n209_ );
nand g062 ( new_n213_, new_n210_, keyIn_0_9, N89 );
nand g063 ( N450, new_n212_, new_n213_ );
not g064 ( new_n215_, N91 );
not g065 ( new_n216_, N96 );
nand g066 ( new_n217_, new_n215_, new_n216_ );
nand g067 ( new_n218_, N91, N96 );
nand g068 ( new_n219_, new_n217_, new_n218_ );
not g069 ( new_n220_, N101 );
not g070 ( new_n221_, N106 );
nand g071 ( new_n222_, new_n220_, new_n221_ );
nand g072 ( new_n223_, N101, N106 );
nand g073 ( new_n224_, new_n222_, new_n223_ );
nand g074 ( new_n225_, new_n219_, new_n224_ );
nand g075 ( new_n226_, new_n217_, new_n222_, new_n218_, new_n223_ );
nand g076 ( new_n227_, new_n225_, new_n226_ );
nand g077 ( new_n228_, new_n227_, N130 );
not g078 ( new_n229_, N130 );
nand g079 ( new_n230_, new_n225_, new_n229_, new_n226_ );
nand g080 ( new_n231_, new_n228_, new_n230_ );
not g081 ( new_n232_, keyIn_0_19 );
not g082 ( new_n233_, N135 );
nor g083 ( new_n234_, N111, N116 );
nor g084 ( new_n235_, new_n234_, keyIn_0_6 );
not g085 ( new_n236_, keyIn_0_6 );
nor g086 ( new_n237_, new_n236_, N111, N116 );
nor g087 ( new_n238_, new_n235_, new_n237_ );
nand g088 ( new_n239_, N111, N116 );
not g089 ( new_n240_, new_n239_ );
nor g090 ( new_n241_, new_n238_, new_n240_ );
not g091 ( new_n242_, new_n241_ );
not g092 ( new_n243_, N126 );
nor g093 ( new_n244_, new_n243_, N121 );
nand g094 ( new_n245_, new_n243_, N121 );
not g095 ( new_n246_, new_n245_ );
nor g096 ( new_n247_, new_n246_, new_n244_ );
not g097 ( new_n248_, new_n247_ );
nand g098 ( new_n249_, new_n242_, new_n248_ );
nand g099 ( new_n250_, new_n241_, new_n247_ );
nand g100 ( new_n251_, new_n249_, new_n232_, new_n233_, new_n250_ );
nand g101 ( new_n252_, new_n249_, new_n233_, new_n250_ );
nand g102 ( new_n253_, new_n252_, keyIn_0_19 );
nand g103 ( new_n254_, new_n249_, new_n250_ );
nand g104 ( new_n255_, new_n254_, N135 );
nand g105 ( new_n256_, new_n253_, new_n255_, new_n231_, new_n251_ );
nor g106 ( new_n257_, new_n256_, keyIn_0_32 );
nand g107 ( new_n258_, new_n256_, keyIn_0_32 );
nand g108 ( new_n259_, new_n253_, new_n251_, new_n255_ );
nand g109 ( new_n260_, new_n259_, new_n228_, new_n230_ );
nand g110 ( new_n261_, new_n260_, new_n258_ );
nor g111 ( N767, new_n261_, new_n257_ );
not g112 ( new_n263_, keyIn_0_25 );
nor g113 ( new_n264_, N159, N165 );
nand g114 ( new_n265_, N159, N165 );
not g115 ( new_n266_, new_n265_ );
nor g116 ( new_n267_, new_n266_, new_n264_, keyIn_0_13 );
not g117 ( new_n268_, new_n267_ );
not g118 ( new_n269_, N171 );
nor g119 ( new_n270_, new_n269_, N177 );
not g120 ( new_n271_, N177 );
nor g121 ( new_n272_, new_n271_, N171 );
nor g122 ( new_n273_, new_n268_, new_n270_, new_n272_ );
nor g123 ( new_n274_, new_n270_, new_n272_ );
nor g124 ( new_n275_, new_n267_, new_n274_ );
nor g125 ( new_n276_, new_n273_, new_n275_ );
nand g126 ( new_n277_, new_n276_, new_n263_, new_n229_ );
nand g127 ( new_n278_, new_n276_, new_n229_ );
nand g128 ( new_n279_, new_n278_, keyIn_0_25 );
not g129 ( new_n280_, new_n276_ );
nand g130 ( new_n281_, new_n280_, N130 );
nand g131 ( new_n282_, new_n279_, new_n281_, keyIn_0_31, new_n277_ );
not g132 ( new_n283_, new_n282_ );
not g133 ( new_n284_, keyIn_0_26 );
not g134 ( new_n285_, N207 );
not g135 ( new_n286_, N183 );
not g136 ( new_n287_, N189 );
nand g137 ( new_n288_, new_n286_, new_n287_ );
nand g138 ( new_n289_, N183, N189 );
nand g139 ( new_n290_, new_n288_, new_n289_ );
not g140 ( new_n291_, N195 );
not g141 ( new_n292_, N201 );
nand g142 ( new_n293_, new_n291_, new_n292_ );
nand g143 ( new_n294_, N195, N201 );
nand g144 ( new_n295_, new_n293_, new_n294_ );
nand g145 ( new_n296_, new_n290_, new_n295_ );
nand g146 ( new_n297_, new_n288_, new_n293_, new_n289_, new_n294_ );
nand g147 ( new_n298_, new_n296_, new_n297_ );
nand g148 ( new_n299_, new_n298_, new_n284_, new_n285_ );
nand g149 ( new_n300_, new_n298_, new_n285_ );
nand g150 ( new_n301_, new_n300_, keyIn_0_26 );
nand g151 ( new_n302_, new_n296_, N207, new_n297_ );
nand g152 ( new_n303_, new_n301_, new_n299_, new_n302_ );
nand g153 ( new_n304_, new_n283_, new_n303_ );
not g154 ( new_n305_, new_n303_ );
nand g155 ( new_n306_, new_n282_, new_n305_ );
nand g156 ( N768, new_n304_, new_n306_ );
not g157 ( new_n308_, keyIn_0_52 );
not g158 ( new_n309_, keyIn_0_24 );
nand g159 ( new_n310_, N59, N156 );
not g160 ( new_n311_, new_n310_ );
nor g161 ( new_n312_, N17, N42 );
nand g162 ( new_n313_, N17, N42 );
not g163 ( new_n314_, new_n313_ );
nor g164 ( new_n315_, new_n314_, new_n312_ );
nand g165 ( new_n316_, new_n315_, new_n194_, new_n195_, new_n311_ );
nand g166 ( new_n317_, N42, N59, N75 );
nand g167 ( new_n318_, new_n167_, N17, N51, new_n317_ );
nand g168 ( new_n319_, new_n316_, new_n318_ );
nand g169 ( new_n320_, new_n319_, N126 );
nand g170 ( new_n321_, new_n320_, new_n309_ );
not g171 ( new_n322_, keyIn_0_15 );
nand g172 ( new_n323_, N29, N55, N75, N80 );
not g173 ( new_n324_, new_n323_ );
nand g174 ( new_n325_, new_n324_, new_n194_, new_n195_ );
nand g175 ( new_n326_, new_n325_, new_n322_ );
nand g176 ( new_n327_, new_n324_, new_n194_, keyIn_0_15, new_n195_ );
nand g177 ( new_n328_, new_n326_, new_n327_ );
not g178 ( new_n329_, N268 );
nand g179 ( new_n330_, new_n329_, keyIn_0_10 );
not g180 ( new_n331_, keyIn_0_10 );
nand g181 ( new_n332_, new_n331_, N268 );
nand g182 ( new_n333_, new_n330_, new_n332_ );
nand g183 ( new_n334_, new_n328_, new_n333_ );
nand g184 ( new_n335_, new_n194_, N17, new_n195_, new_n310_ );
nand g185 ( new_n336_, new_n335_, N1 );
nand g186 ( new_n337_, new_n336_, N153 );
nand g187 ( new_n338_, new_n319_, keyIn_0_24, N126 );
nand g188 ( new_n339_, new_n321_, new_n334_, new_n337_, new_n338_ );
nand g189 ( new_n340_, new_n339_, N201 );
nand g190 ( new_n341_, new_n340_, keyIn_0_37 );
not g191 ( new_n342_, keyIn_0_37 );
nand g192 ( new_n343_, new_n339_, new_n342_, N201 );
nand g193 ( new_n344_, new_n341_, new_n343_ );
nand g194 ( new_n345_, new_n338_, new_n337_ );
not g195 ( new_n346_, new_n345_ );
nand g196 ( new_n347_, new_n346_, new_n292_, new_n321_, new_n334_ );
nor g197 ( new_n348_, new_n347_, keyIn_0_38 );
not g198 ( new_n349_, keyIn_0_38 );
nor g199 ( new_n350_, new_n339_, N201 );
nor g200 ( new_n351_, new_n350_, new_n349_ );
nor g201 ( new_n352_, new_n351_, new_n348_ );
nand g202 ( new_n353_, new_n352_, new_n344_ );
not g203 ( new_n354_, new_n353_ );
nand g204 ( new_n355_, new_n354_, N261 );
not g205 ( new_n356_, N261 );
nand g206 ( new_n357_, new_n353_, new_n356_ );
nand g207 ( new_n358_, new_n355_, new_n308_, new_n357_ );
nand g208 ( new_n359_, new_n355_, new_n357_ );
nand g209 ( new_n360_, new_n359_, keyIn_0_52 );
nand g210 ( new_n361_, new_n360_, N219, new_n358_ );
nand g211 ( new_n362_, N121, N210 );
nand g212 ( new_n363_, new_n361_, new_n362_ );
nand g213 ( new_n364_, new_n363_, keyIn_0_56 );
not g214 ( new_n365_, keyIn_0_56 );
nand g215 ( new_n366_, new_n361_, new_n365_, new_n362_ );
nand g216 ( new_n367_, new_n364_, new_n366_ );
not g217 ( new_n368_, keyIn_0_11 );
nand g218 ( new_n369_, new_n202_, N42, N72, new_n204_ );
not g219 ( new_n370_, new_n369_ );
nand g220 ( new_n371_, new_n370_, keyIn_0_8 );
not g221 ( new_n372_, keyIn_0_8 );
nand g222 ( new_n373_, new_n369_, new_n372_ );
nand g223 ( new_n374_, new_n371_, N73, new_n373_ );
nand g224 ( new_n375_, new_n374_, new_n368_ );
nand g225 ( new_n376_, new_n371_, keyIn_0_11, N73, new_n373_ );
nand g226 ( new_n377_, new_n375_, new_n376_ );
nand g227 ( new_n378_, new_n377_, keyIn_0_14 );
not g228 ( new_n379_, keyIn_0_14 );
nand g229 ( new_n380_, new_n375_, new_n379_, new_n376_ );
nand g230 ( new_n381_, new_n378_, new_n380_ );
nand g231 ( new_n382_, new_n381_, keyIn_0_16 );
not g232 ( new_n383_, keyIn_0_16 );
nand g233 ( new_n384_, new_n378_, new_n383_, new_n380_ );
nand g234 ( new_n385_, new_n382_, new_n384_ );
not g235 ( new_n386_, new_n385_ );
nand g236 ( new_n387_, new_n386_, N201 );
nand g237 ( new_n388_, new_n387_, keyIn_0_28 );
not g238 ( new_n389_, keyIn_0_28 );
nand g239 ( new_n390_, new_n386_, new_n389_, N201 );
nand g240 ( new_n391_, new_n388_, new_n390_ );
nand g241 ( new_n392_, new_n354_, N228 );
nand g242 ( new_n393_, N255, N267 );
nand g243 ( new_n394_, new_n339_, N246 );
nand g244 ( new_n395_, new_n392_, new_n393_, new_n394_ );
not g245 ( new_n396_, new_n344_ );
nand g246 ( new_n397_, new_n396_, N237 );
nand g247 ( new_n398_, new_n397_, keyIn_0_50 );
not g248 ( new_n399_, keyIn_0_50 );
nand g249 ( new_n400_, new_n396_, new_n399_, N237 );
nand g250 ( new_n401_, new_n398_, new_n400_ );
nor g251 ( new_n402_, new_n395_, new_n401_ );
nand g252 ( N850, new_n367_, new_n391_, new_n402_ );
not g253 ( new_n404_, keyIn_0_51 );
nand g254 ( new_n405_, new_n336_, N146 );
nand g255 ( new_n406_, new_n319_, keyIn_0_23, N116 );
not g256 ( new_n407_, keyIn_0_23 );
nand g257 ( new_n408_, new_n319_, N116 );
nand g258 ( new_n409_, new_n408_, new_n407_ );
nand g259 ( new_n410_, new_n409_, new_n334_, new_n405_, new_n406_ );
nand g260 ( new_n411_, new_n410_, keyIn_0_30 );
not g261 ( new_n412_, keyIn_0_30 );
nand g262 ( new_n413_, new_n406_, new_n405_ );
not g263 ( new_n414_, new_n413_ );
nand g264 ( new_n415_, new_n414_, new_n412_, new_n334_, new_n409_ );
nand g265 ( new_n416_, new_n415_, new_n411_ );
nand g266 ( new_n417_, new_n416_, new_n287_ );
nand g267 ( new_n418_, new_n336_, N149 );
nand g268 ( new_n419_, new_n319_, N121 );
nand g269 ( new_n420_, new_n334_, new_n419_, new_n291_, new_n418_ );
nand g270 ( new_n421_, new_n417_, new_n341_, new_n343_, new_n420_ );
nand g271 ( new_n422_, new_n421_, new_n404_ );
nand g272 ( new_n423_, new_n396_, keyIn_0_51, new_n417_, new_n420_ );
nand g273 ( new_n424_, new_n422_, new_n423_ );
not g274 ( new_n425_, keyIn_0_42 );
nand g275 ( new_n426_, new_n350_, new_n349_ );
nand g276 ( new_n427_, new_n347_, keyIn_0_38 );
nand g277 ( new_n428_, new_n426_, new_n427_, N261 );
not g278 ( new_n429_, new_n428_ );
nand g279 ( new_n430_, new_n429_, new_n425_, new_n417_, new_n420_ );
nand g280 ( new_n431_, new_n352_, N261, new_n417_, new_n420_ );
nand g281 ( new_n432_, new_n431_, keyIn_0_42 );
nand g282 ( new_n433_, new_n334_, new_n418_, new_n419_ );
nand g283 ( new_n434_, new_n433_, N195 );
not g284 ( new_n435_, new_n434_ );
nand g285 ( new_n436_, new_n417_, new_n435_ );
not g286 ( new_n437_, new_n416_ );
nand g287 ( new_n438_, new_n437_, N189 );
nand g288 ( new_n439_, new_n436_, new_n438_ );
not g289 ( new_n440_, new_n439_ );
nand g290 ( new_n441_, new_n424_, new_n430_, new_n432_, new_n440_ );
not g291 ( new_n442_, keyIn_0_29 );
nand g292 ( new_n443_, new_n336_, N143 );
nand g293 ( new_n444_, new_n319_, N111 );
nand g294 ( new_n445_, new_n444_, keyIn_0_22 );
not g295 ( new_n446_, keyIn_0_22 );
nand g296 ( new_n447_, new_n319_, new_n446_, N111 );
nand g297 ( new_n448_, new_n445_, new_n334_, new_n443_, new_n447_ );
nand g298 ( new_n449_, new_n448_, new_n442_ );
nand g299 ( new_n450_, new_n334_, new_n443_ );
not g300 ( new_n451_, new_n450_ );
nand g301 ( new_n452_, new_n451_, keyIn_0_29, new_n445_, new_n447_ );
nand g302 ( new_n453_, new_n452_, new_n449_ );
nand g303 ( new_n454_, new_n453_, N183 );
nand g304 ( new_n455_, new_n454_, keyIn_0_36 );
not g305 ( new_n456_, keyIn_0_36 );
nand g306 ( new_n457_, new_n453_, new_n456_, N183 );
nand g307 ( new_n458_, new_n455_, new_n457_ );
not g308 ( new_n459_, new_n458_ );
nand g309 ( new_n460_, new_n452_, new_n449_, new_n286_ );
nand g310 ( new_n461_, new_n459_, new_n460_ );
not g311 ( new_n462_, new_n461_ );
nand g312 ( new_n463_, new_n441_, keyIn_0_53, new_n462_ );
not g313 ( new_n464_, keyIn_0_53 );
nand g314 ( new_n465_, new_n441_, new_n462_ );
nand g315 ( new_n466_, new_n465_, new_n464_ );
not g316 ( new_n467_, new_n441_ );
nand g317 ( new_n468_, new_n467_, new_n461_ );
nand g318 ( new_n469_, new_n466_, new_n468_, keyIn_0_55, new_n463_ );
not g319 ( new_n470_, keyIn_0_55 );
nand g320 ( new_n471_, new_n466_, new_n463_, new_n468_ );
nand g321 ( new_n472_, new_n471_, new_n470_ );
nand g322 ( new_n473_, new_n472_, N219, new_n469_ );
not g323 ( new_n474_, keyIn_0_47 );
nand g324 ( new_n475_, new_n462_, N228 );
nand g325 ( new_n476_, new_n475_, new_n474_ );
nand g326 ( new_n477_, new_n386_, keyIn_0_27, N183 );
not g327 ( new_n478_, keyIn_0_27 );
nand g328 ( new_n479_, new_n386_, N183 );
nand g329 ( new_n480_, new_n479_, new_n478_ );
nand g330 ( new_n481_, new_n453_, N246 );
nand g331 ( new_n482_, N106, N210 );
nand g332 ( new_n483_, new_n481_, new_n482_ );
not g333 ( new_n484_, new_n483_ );
nand g334 ( new_n485_, new_n476_, new_n477_, new_n480_, new_n484_ );
not g335 ( new_n486_, new_n485_ );
nand g336 ( new_n487_, new_n462_, keyIn_0_47, N228 );
not g337 ( new_n488_, keyIn_0_40 );
nand g338 ( new_n489_, new_n458_, new_n488_ );
nand g339 ( new_n490_, new_n455_, keyIn_0_40, new_n457_ );
nand g340 ( new_n491_, new_n489_, N237, new_n490_ );
nand g341 ( N863, new_n473_, new_n486_, new_n487_, new_n491_ );
nand g342 ( new_n493_, new_n438_, new_n417_ );
nand g343 ( new_n494_, new_n428_, new_n344_ );
nand g344 ( new_n495_, new_n494_, new_n420_ );
not g345 ( new_n496_, keyIn_0_49 );
nand g346 ( new_n497_, new_n435_, new_n496_ );
nand g347 ( new_n498_, new_n434_, keyIn_0_49 );
nand g348 ( new_n499_, new_n497_, new_n498_ );
nand g349 ( new_n500_, new_n495_, new_n493_, new_n499_ );
not g350 ( new_n501_, new_n493_ );
nand g351 ( new_n502_, new_n495_, new_n499_ );
nand g352 ( new_n503_, new_n502_, new_n501_ );
nand g353 ( new_n504_, new_n503_, N219, new_n500_ );
nand g354 ( new_n505_, new_n437_, N189, N237 );
nand g355 ( new_n506_, N111, N210 );
nand g356 ( new_n507_, new_n386_, N189 );
nand g357 ( new_n508_, new_n507_, new_n505_, new_n506_ );
not g358 ( new_n509_, keyIn_0_41 );
nand g359 ( new_n510_, new_n437_, N246 );
nand g360 ( new_n511_, N255, N259 );
nand g361 ( new_n512_, new_n510_, new_n511_ );
nand g362 ( new_n513_, new_n512_, new_n509_ );
nand g363 ( new_n514_, new_n510_, keyIn_0_41, new_n511_ );
nand g364 ( new_n515_, new_n513_, new_n514_ );
nor g365 ( new_n516_, new_n508_, new_n515_ );
not g366 ( new_n517_, keyIn_0_48 );
nand g367 ( new_n518_, new_n501_, N228 );
nand g368 ( new_n519_, new_n518_, new_n517_ );
nand g369 ( new_n520_, new_n501_, keyIn_0_48, N228 );
nand g370 ( N864, new_n516_, new_n504_, new_n519_, new_n520_ );
nand g371 ( new_n522_, new_n434_, new_n420_ );
not g372 ( new_n523_, new_n522_ );
nand g373 ( new_n524_, new_n494_, new_n523_ );
nand g374 ( new_n525_, new_n428_, new_n344_, new_n522_ );
nand g375 ( new_n526_, new_n524_, N219, new_n525_ );
nand g376 ( new_n527_, new_n386_, N195 );
nand g377 ( new_n528_, new_n523_, N228 );
nand g378 ( new_n529_, new_n435_, N237 );
nand g379 ( new_n530_, new_n433_, N246 );
nand g380 ( new_n531_, N116, N210 );
nand g381 ( new_n532_, N255, N260 );
nand g382 ( new_n533_, new_n529_, new_n530_, new_n531_, new_n532_ );
not g383 ( new_n534_, new_n533_ );
nand g384 ( N865, new_n527_, new_n526_, new_n528_, new_n534_ );
nand g385 ( new_n536_, new_n489_, new_n490_ );
nand g386 ( new_n537_, new_n536_, keyIn_0_46 );
not g387 ( new_n538_, keyIn_0_46 );
nand g388 ( new_n539_, new_n489_, new_n538_, new_n490_ );
nand g389 ( new_n540_, new_n537_, new_n539_ );
nand g390 ( new_n541_, new_n441_, new_n460_ );
nand g391 ( new_n542_, new_n540_, new_n541_ );
nand g392 ( new_n543_, new_n542_, keyIn_0_54 );
not g393 ( new_n544_, keyIn_0_54 );
nand g394 ( new_n545_, new_n540_, new_n541_, new_n544_ );
nand g395 ( new_n546_, new_n543_, new_n545_ );
nand g396 ( new_n547_, N29, N75, N80 );
not g397 ( new_n548_, new_n547_ );
nand g398 ( new_n549_, N447, N17, new_n329_, new_n548_ );
not g399 ( new_n550_, new_n549_ );
nand g400 ( new_n551_, new_n550_, keyIn_0_18 );
not g401 ( new_n552_, keyIn_0_18 );
nand g402 ( new_n553_, new_n549_, new_n552_ );
nand g403 ( new_n554_, new_n551_, new_n553_ );
nand g404 ( new_n555_, new_n319_, N106 );
not g405 ( new_n556_, N55 );
nor g406 ( new_n557_, new_n196_, new_n556_, new_n311_ );
nand g407 ( new_n558_, new_n557_, N153 );
nand g408 ( new_n559_, N138, N152 );
nand g409 ( new_n560_, new_n558_, new_n559_ );
not g410 ( new_n561_, new_n560_ );
nand g411 ( new_n562_, new_n554_, new_n271_, new_n555_, new_n561_ );
nand g412 ( new_n563_, new_n546_, new_n562_ );
nand g413 ( new_n564_, new_n554_, new_n555_, new_n561_ );
nand g414 ( new_n565_, new_n564_, N177 );
nand g415 ( new_n566_, new_n563_, new_n565_ );
not g416 ( new_n567_, keyIn_0_17 );
nand g417 ( new_n568_, new_n557_, N149 );
nand g418 ( new_n569_, new_n568_, new_n567_ );
nand g419 ( new_n570_, new_n557_, keyIn_0_17, N149 );
nand g420 ( new_n571_, new_n569_, new_n570_ );
nand g421 ( new_n572_, new_n319_, N101 );
nand g422 ( new_n573_, N17, N138 );
nand g423 ( new_n574_, new_n571_, new_n549_, new_n572_, new_n573_ );
not g424 ( new_n575_, new_n574_ );
nand g425 ( new_n576_, new_n575_, new_n269_ );
nand g426 ( new_n577_, new_n566_, new_n576_ );
nand g427 ( new_n578_, new_n574_, N171 );
nand g428 ( new_n579_, new_n578_, keyIn_0_35 );
not g429 ( new_n580_, keyIn_0_35 );
nand g430 ( new_n581_, new_n574_, new_n580_, N171 );
nand g431 ( new_n582_, new_n579_, new_n581_ );
nand g432 ( new_n583_, new_n577_, new_n582_ );
nand g433 ( new_n584_, new_n557_, N146 );
nand g434 ( new_n585_, new_n584_, keyIn_0_21, new_n549_ );
not g435 ( new_n586_, keyIn_0_21 );
nand g436 ( new_n587_, new_n584_, new_n549_ );
nand g437 ( new_n588_, new_n587_, new_n586_ );
nand g438 ( new_n589_, N51, N138 );
nand g439 ( new_n590_, new_n319_, N96 );
nand g440 ( new_n591_, new_n588_, new_n585_, new_n589_, new_n590_ );
nor g441 ( new_n592_, new_n591_, N165 );
not g442 ( new_n593_, new_n592_ );
nand g443 ( new_n594_, new_n583_, new_n593_ );
nand g444 ( new_n595_, new_n591_, N165 );
nand g445 ( new_n596_, new_n594_, new_n595_ );
not g446 ( new_n597_, keyIn_0_20 );
nand g447 ( new_n598_, new_n557_, N143 );
nand g448 ( new_n599_, new_n598_, new_n597_, new_n549_ );
nand g449 ( new_n600_, new_n598_, new_n549_ );
nand g450 ( new_n601_, new_n600_, keyIn_0_20 );
nand g451 ( new_n602_, N8, N138 );
nand g452 ( new_n603_, new_n319_, N91 );
nand g453 ( new_n604_, new_n601_, new_n599_, new_n602_, new_n603_ );
nor g454 ( new_n605_, new_n604_, N159 );
nor g455 ( new_n606_, new_n605_, keyIn_0_33 );
not g456 ( new_n607_, keyIn_0_33 );
nor g457 ( new_n608_, new_n604_, new_n607_, N159 );
nor g458 ( new_n609_, new_n606_, new_n608_ );
nand g459 ( new_n610_, new_n596_, new_n609_ );
not g460 ( new_n611_, keyIn_0_43 );
nand g461 ( new_n612_, new_n604_, N159 );
not g462 ( new_n613_, new_n612_ );
nand g463 ( new_n614_, new_n613_, new_n611_ );
nand g464 ( new_n615_, new_n612_, keyIn_0_43 );
nand g465 ( new_n616_, new_n614_, new_n615_ );
nand g466 ( new_n617_, new_n610_, new_n616_ );
nand g467 ( new_n618_, new_n617_, keyIn_0_59 );
not g468 ( new_n619_, keyIn_0_59 );
nand g469 ( new_n620_, new_n610_, new_n619_, new_n616_ );
nand g470 ( N866, new_n618_, new_n620_ );
not g471 ( new_n622_, keyIn_0_62 );
not g472 ( new_n623_, new_n546_ );
nand g473 ( new_n624_, new_n565_, new_n562_ );
nand g474 ( new_n625_, new_n623_, keyIn_0_57, new_n624_ );
not g475 ( new_n626_, keyIn_0_57 );
nand g476 ( new_n627_, new_n623_, new_n624_ );
nand g477 ( new_n628_, new_n627_, new_n626_ );
not g478 ( new_n629_, new_n624_ );
nand g479 ( new_n630_, new_n546_, new_n629_ );
nand g480 ( new_n631_, new_n628_, N219, new_n625_, new_n630_ );
nand g481 ( new_n632_, new_n386_, N177 );
nand g482 ( new_n633_, new_n629_, N228 );
nand g483 ( new_n634_, new_n564_, N177, N237 );
nand g484 ( new_n635_, N101, N210 );
nand g485 ( new_n636_, new_n564_, N246 );
nand g486 ( new_n637_, new_n634_, new_n635_, new_n636_ );
not g487 ( new_n638_, new_n637_ );
nand g488 ( new_n639_, new_n632_, new_n633_, new_n638_ );
not g489 ( new_n640_, new_n639_ );
nand g490 ( new_n641_, new_n631_, new_n640_ );
nand g491 ( new_n642_, new_n641_, new_n622_ );
nand g492 ( new_n643_, new_n631_, keyIn_0_62, new_n640_ );
nand g493 ( N874, new_n642_, new_n643_ );
nand g494 ( new_n645_, new_n596_, new_n609_, new_n612_ );
nand g495 ( new_n646_, new_n609_, new_n612_ );
nand g496 ( new_n647_, new_n594_, new_n595_, new_n646_ );
nand g497 ( new_n648_, new_n645_, N219, new_n647_ );
not g498 ( new_n649_, keyIn_0_39 );
nand g499 ( new_n650_, new_n386_, N159 );
not g500 ( new_n651_, keyIn_0_34 );
nand g501 ( new_n652_, new_n604_, N246 );
nand g502 ( new_n653_, new_n652_, new_n651_ );
nand g503 ( new_n654_, new_n604_, keyIn_0_34, N246 );
nand g504 ( new_n655_, new_n653_, new_n654_ );
nand g505 ( new_n656_, new_n650_, new_n649_, new_n655_ );
nand g506 ( new_n657_, new_n650_, new_n655_ );
nand g507 ( new_n658_, new_n657_, keyIn_0_39 );
not g508 ( new_n659_, N228 );
nor g509 ( new_n660_, new_n646_, new_n659_ );
nand g510 ( new_n661_, new_n613_, N237 );
nand g511 ( new_n662_, new_n330_, new_n332_, N210 );
nand g512 ( new_n663_, new_n661_, new_n662_ );
nor g513 ( new_n664_, new_n660_, new_n663_ );
nand g514 ( N878, new_n648_, new_n656_, new_n658_, new_n664_ );
not g515 ( new_n666_, keyIn_0_60 );
not g516 ( new_n667_, new_n595_ );
nor g517 ( new_n668_, new_n667_, new_n592_ );
not g518 ( new_n669_, new_n668_ );
not g519 ( new_n670_, new_n582_ );
nand g520 ( new_n671_, new_n670_, keyIn_0_44 );
not g521 ( new_n672_, keyIn_0_44 );
nand g522 ( new_n673_, new_n582_, new_n672_ );
nand g523 ( new_n674_, new_n671_, new_n673_ );
not g524 ( new_n675_, new_n674_ );
nand g525 ( new_n676_, new_n577_, new_n669_, new_n675_ );
nand g526 ( new_n677_, new_n676_, keyIn_0_58 );
not g527 ( new_n678_, keyIn_0_58 );
nand g528 ( new_n679_, new_n577_, new_n678_, new_n669_, new_n675_ );
nand g529 ( new_n680_, new_n677_, new_n679_ );
nand g530 ( new_n681_, new_n577_, new_n675_ );
nand g531 ( new_n682_, new_n681_, new_n668_ );
nand g532 ( new_n683_, new_n680_, N219, new_n682_ );
not g533 ( new_n684_, keyIn_0_7 );
nand g534 ( new_n685_, N91, N210 );
nand g535 ( new_n686_, new_n685_, new_n684_ );
nand g536 ( new_n687_, keyIn_0_7, N91, N210 );
nand g537 ( new_n688_, new_n686_, new_n687_ );
nand g538 ( new_n689_, new_n683_, new_n688_ );
nand g539 ( new_n690_, new_n689_, new_n666_ );
nand g540 ( new_n691_, new_n683_, keyIn_0_60, new_n688_ );
nand g541 ( new_n692_, new_n690_, new_n691_ );
nand g542 ( new_n693_, new_n386_, N165 );
not g543 ( new_n694_, new_n693_ );
nand g544 ( new_n695_, new_n668_, N228 );
nand g545 ( new_n696_, new_n591_, N246 );
nand g546 ( new_n697_, new_n667_, N237 );
nand g547 ( new_n698_, new_n695_, new_n696_, new_n697_ );
nor g548 ( new_n699_, new_n694_, new_n698_ );
nand g549 ( N879, new_n692_, new_n699_ );
not g550 ( new_n701_, keyIn_0_61 );
nand g551 ( new_n702_, new_n582_, new_n576_ );
not g552 ( new_n703_, new_n702_ );
nand g553 ( new_n704_, new_n566_, new_n703_ );
nand g554 ( new_n705_, new_n563_, new_n565_, new_n702_ );
nand g555 ( new_n706_, new_n704_, N219, new_n705_ );
nand g556 ( new_n707_, N96, N210 );
nand g557 ( new_n708_, new_n706_, new_n707_ );
nand g558 ( new_n709_, new_n708_, new_n701_ );
nand g559 ( new_n710_, new_n706_, keyIn_0_61, new_n707_ );
nand g560 ( new_n711_, new_n709_, new_n710_ );
nand g561 ( new_n712_, new_n386_, N171 );
nand g562 ( new_n713_, new_n574_, N246 );
nand g563 ( new_n714_, new_n712_, new_n713_ );
not g564 ( new_n715_, keyIn_0_45 );
nand g565 ( new_n716_, new_n670_, N237 );
nand g566 ( new_n717_, new_n716_, new_n715_ );
nand g567 ( new_n718_, new_n703_, N228 );
nand g568 ( new_n719_, new_n670_, keyIn_0_45, N237 );
nand g569 ( new_n720_, new_n717_, new_n718_, new_n719_ );
nor g570 ( new_n721_, new_n714_, new_n720_ );
nand g571 ( new_n722_, new_n711_, new_n721_ );
nand g572 ( new_n723_, new_n722_, keyIn_0_63 );
not g573 ( new_n724_, keyIn_0_63 );
nand g574 ( new_n725_, new_n711_, new_n724_, new_n721_ );
nand g575 ( N880, new_n723_, new_n725_ );
endmodule