module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n170_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n959_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n759_, new_n630_, new_n167_, new_n385_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n158_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n970_, new_n466_, new_n262_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n940_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n824_, new_n143_, new_n520_, new_n1001_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n968_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n913_, new_n327_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_;

and g000 ( new_n138_, N73, N77 );
not g001 ( new_n139_, N73 );
not g002 ( new_n140_, N77 );
and g003 ( new_n141_, new_n139_, new_n140_ );
or g004 ( new_n142_, new_n141_, new_n138_ );
not g005 ( new_n143_, new_n142_ );
and g006 ( new_n144_, N65, N69 );
not g007 ( new_n145_, N65 );
not g008 ( new_n146_, N69 );
and g009 ( new_n147_, new_n145_, new_n146_ );
or g010 ( new_n148_, new_n147_, new_n144_ );
not g011 ( new_n149_, new_n148_ );
and g012 ( new_n150_, new_n143_, new_n149_ );
and g013 ( new_n151_, new_n142_, new_n148_ );
or g014 ( new_n152_, new_n150_, new_n151_ );
and g015 ( new_n153_, N89, N93 );
not g016 ( new_n154_, N89 );
not g017 ( new_n155_, N93 );
and g018 ( new_n156_, new_n154_, new_n155_ );
or g019 ( new_n157_, new_n156_, new_n153_ );
not g020 ( new_n158_, new_n157_ );
and g021 ( new_n159_, N81, N85 );
not g022 ( new_n160_, N81 );
not g023 ( new_n161_, N85 );
and g024 ( new_n162_, new_n160_, new_n161_ );
or g025 ( new_n163_, new_n162_, new_n159_ );
not g026 ( new_n164_, new_n163_ );
and g027 ( new_n165_, new_n158_, new_n164_ );
and g028 ( new_n166_, new_n157_, new_n163_ );
or g029 ( new_n167_, new_n165_, new_n166_ );
not g030 ( new_n168_, new_n167_ );
and g031 ( new_n169_, new_n168_, new_n152_ );
not g032 ( new_n170_, new_n152_ );
and g033 ( new_n171_, new_n170_, new_n167_ );
or g034 ( new_n172_, new_n169_, new_n171_ );
and g035 ( new_n173_, N129, N137 );
and g036 ( new_n174_, new_n172_, new_n173_ );
not g037 ( new_n175_, new_n174_ );
or g038 ( new_n176_, new_n172_, new_n173_ );
and g039 ( new_n177_, new_n175_, new_n176_ );
and g040 ( new_n178_, N33, N49 );
not g041 ( new_n179_, N33 );
not g042 ( new_n180_, N49 );
and g043 ( new_n181_, new_n179_, new_n180_ );
or g044 ( new_n182_, new_n181_, new_n178_ );
not g045 ( new_n183_, new_n182_ );
and g046 ( new_n184_, N1, N17 );
not g047 ( new_n185_, N1 );
not g048 ( new_n186_, N17 );
and g049 ( new_n187_, new_n185_, new_n186_ );
or g050 ( new_n188_, new_n187_, new_n184_ );
not g051 ( new_n189_, new_n188_ );
and g052 ( new_n190_, new_n183_, new_n189_ );
and g053 ( new_n191_, new_n182_, new_n188_ );
or g054 ( new_n192_, new_n190_, new_n191_ );
not g055 ( new_n193_, new_n192_ );
and g056 ( new_n194_, new_n177_, new_n193_ );
not g057 ( new_n195_, new_n194_ );
or g058 ( new_n196_, new_n177_, new_n193_ );
and g059 ( new_n197_, new_n195_, new_n196_ );
not g060 ( new_n198_, keyIn_0_19 );
not g061 ( new_n199_, keyIn_0_14 );
not g062 ( new_n200_, N37 );
and g063 ( new_n201_, new_n179_, new_n200_ );
and g064 ( new_n202_, N33, N37 );
or g065 ( new_n203_, new_n201_, new_n202_ );
and g066 ( new_n204_, new_n203_, keyIn_0_4 );
not g067 ( new_n205_, keyIn_0_4 );
or g068 ( new_n206_, N33, N37 );
not g069 ( new_n207_, new_n202_ );
and g070 ( new_n208_, new_n207_, new_n206_ );
and g071 ( new_n209_, new_n208_, new_n205_ );
or g072 ( new_n210_, new_n204_, new_n209_ );
not g073 ( new_n211_, keyIn_0_5 );
and g074 ( new_n212_, N41, N45 );
not g075 ( new_n213_, new_n212_ );
or g076 ( new_n214_, N41, N45 );
and g077 ( new_n215_, new_n213_, new_n214_ );
and g078 ( new_n216_, new_n215_, new_n211_ );
not g079 ( new_n217_, N41 );
not g080 ( new_n218_, N45 );
and g081 ( new_n219_, new_n217_, new_n218_ );
or g082 ( new_n220_, new_n219_, new_n212_ );
and g083 ( new_n221_, new_n220_, keyIn_0_5 );
or g084 ( new_n222_, new_n221_, new_n216_ );
and g085 ( new_n223_, new_n210_, new_n222_ );
or g086 ( new_n224_, new_n208_, new_n205_ );
or g087 ( new_n225_, new_n203_, keyIn_0_4 );
or g088 ( new_n226_, new_n220_, keyIn_0_5 );
or g089 ( new_n227_, new_n215_, new_n211_ );
and g090 ( new_n228_, new_n225_, new_n226_, new_n224_, new_n227_ );
or g091 ( new_n229_, new_n223_, new_n228_ );
or g092 ( new_n230_, new_n229_, new_n199_ );
and g093 ( new_n231_, new_n229_, new_n199_ );
not g094 ( new_n232_, new_n231_ );
and g095 ( new_n233_, new_n232_, new_n230_ );
not g096 ( new_n234_, keyIn_0_12 );
not g097 ( new_n235_, keyIn_0_0 );
and g098 ( new_n236_, N1, N5 );
not g099 ( new_n237_, new_n236_ );
or g100 ( new_n238_, N1, N5 );
and g101 ( new_n239_, new_n237_, new_n238_ );
and g102 ( new_n240_, new_n239_, new_n235_ );
not g103 ( new_n241_, new_n240_ );
or g104 ( new_n242_, new_n239_, new_n235_ );
and g105 ( new_n243_, new_n241_, new_n242_ );
not g106 ( new_n244_, keyIn_0_1 );
and g107 ( new_n245_, N9, N13 );
not g108 ( new_n246_, N9 );
not g109 ( new_n247_, N13 );
and g110 ( new_n248_, new_n246_, new_n247_ );
or g111 ( new_n249_, new_n248_, new_n245_ );
or g112 ( new_n250_, new_n249_, new_n244_ );
not g113 ( new_n251_, new_n245_ );
or g114 ( new_n252_, N9, N13 );
and g115 ( new_n253_, new_n251_, new_n252_ );
or g116 ( new_n254_, new_n253_, keyIn_0_1 );
and g117 ( new_n255_, new_n250_, new_n254_ );
or g118 ( new_n256_, new_n243_, new_n255_ );
and g119 ( new_n257_, new_n241_, new_n250_, new_n242_, new_n254_ );
not g120 ( new_n258_, new_n257_ );
and g121 ( new_n259_, new_n256_, new_n234_, new_n258_ );
not g122 ( new_n260_, new_n259_ );
and g123 ( new_n261_, new_n256_, new_n258_ );
or g124 ( new_n262_, new_n261_, new_n234_ );
and g125 ( new_n263_, new_n262_, new_n260_ );
or g126 ( new_n264_, new_n233_, new_n263_ );
and g127 ( new_n265_, new_n232_, new_n262_, new_n230_, new_n260_ );
not g128 ( new_n266_, new_n265_ );
and g129 ( new_n267_, new_n264_, new_n266_ );
or g130 ( new_n268_, new_n267_, new_n198_ );
and g131 ( new_n269_, new_n264_, new_n198_, new_n266_ );
not g132 ( new_n270_, new_n269_ );
and g133 ( new_n271_, new_n268_, new_n270_ );
and g134 ( new_n272_, N135, N137 );
or g135 ( new_n273_, new_n272_, keyIn_0_7 );
and g136 ( new_n274_, new_n272_, keyIn_0_7 );
not g137 ( new_n275_, new_n274_ );
and g138 ( new_n276_, new_n275_, new_n273_ );
or g139 ( new_n277_, new_n271_, new_n276_ );
and g140 ( new_n278_, new_n268_, new_n270_, new_n276_ );
not g141 ( new_n279_, new_n278_ );
and g142 ( new_n280_, new_n277_, new_n279_ );
or g143 ( new_n281_, new_n280_, keyIn_0_21 );
and g144 ( new_n282_, new_n277_, new_n279_, keyIn_0_21 );
not g145 ( new_n283_, new_n282_ );
and g146 ( new_n284_, new_n281_, new_n283_ );
not g147 ( new_n285_, keyIn_0_17 );
and g148 ( new_n286_, new_n154_, N73 );
and g149 ( new_n287_, new_n139_, N89 );
or g150 ( new_n288_, new_n286_, new_n287_ );
and g151 ( new_n289_, new_n288_, keyIn_0_10 );
not g152 ( new_n290_, new_n289_ );
or g153 ( new_n291_, new_n288_, keyIn_0_10 );
and g154 ( new_n292_, new_n290_, new_n291_ );
not g155 ( new_n293_, keyIn_0_11 );
and g156 ( new_n294_, N105, N121 );
not g157 ( new_n295_, N105 );
not g158 ( new_n296_, N121 );
and g159 ( new_n297_, new_n295_, new_n296_ );
or g160 ( new_n298_, new_n297_, new_n294_ );
not g161 ( new_n299_, new_n298_ );
and g162 ( new_n300_, new_n299_, new_n293_ );
and g163 ( new_n301_, new_n298_, keyIn_0_11 );
or g164 ( new_n302_, new_n300_, new_n301_ );
not g165 ( new_n303_, new_n302_ );
and g166 ( new_n304_, new_n303_, new_n292_ );
not g167 ( new_n305_, new_n304_ );
or g168 ( new_n306_, new_n303_, new_n292_ );
and g169 ( new_n307_, new_n305_, new_n306_ );
and g170 ( new_n308_, new_n307_, new_n285_ );
not g171 ( new_n309_, new_n308_ );
or g172 ( new_n310_, new_n307_, new_n285_ );
and g173 ( new_n311_, new_n309_, new_n310_ );
or g174 ( new_n312_, new_n284_, new_n311_ );
and g175 ( new_n313_, new_n281_, new_n283_, new_n311_ );
not g176 ( new_n314_, new_n313_ );
and g177 ( new_n315_, new_n312_, new_n314_, keyIn_0_23 );
not g178 ( new_n316_, keyIn_0_23 );
not g179 ( new_n317_, keyIn_0_21 );
and g180 ( new_n318_, new_n225_, new_n224_ );
and g181 ( new_n319_, new_n226_, new_n227_ );
or g182 ( new_n320_, new_n318_, new_n319_ );
not g183 ( new_n321_, new_n228_ );
and g184 ( new_n322_, new_n320_, new_n321_ );
and g185 ( new_n323_, new_n322_, keyIn_0_14 );
or g186 ( new_n324_, new_n323_, new_n231_ );
not g187 ( new_n325_, N5 );
and g188 ( new_n326_, new_n185_, new_n325_ );
or g189 ( new_n327_, new_n326_, new_n236_ );
and g190 ( new_n328_, new_n327_, keyIn_0_0 );
or g191 ( new_n329_, new_n328_, new_n240_ );
and g192 ( new_n330_, new_n253_, keyIn_0_1 );
and g193 ( new_n331_, new_n249_, new_n244_ );
or g194 ( new_n332_, new_n331_, new_n330_ );
and g195 ( new_n333_, new_n329_, new_n332_ );
or g196 ( new_n334_, new_n333_, new_n257_ );
and g197 ( new_n335_, new_n334_, keyIn_0_12 );
or g198 ( new_n336_, new_n335_, new_n259_ );
and g199 ( new_n337_, new_n324_, new_n336_ );
or g200 ( new_n338_, new_n337_, new_n265_ );
and g201 ( new_n339_, new_n338_, keyIn_0_19 );
or g202 ( new_n340_, new_n339_, new_n269_ );
not g203 ( new_n341_, new_n276_ );
and g204 ( new_n342_, new_n340_, new_n341_ );
or g205 ( new_n343_, new_n342_, new_n278_ );
and g206 ( new_n344_, new_n343_, new_n317_ );
or g207 ( new_n345_, new_n344_, new_n282_ );
not g208 ( new_n346_, new_n311_ );
and g209 ( new_n347_, new_n345_, new_n346_ );
or g210 ( new_n348_, new_n347_, new_n313_ );
and g211 ( new_n349_, new_n348_, new_n316_ );
or g212 ( new_n350_, new_n349_, new_n315_ );
not g213 ( new_n351_, keyIn_0_13 );
and g214 ( new_n352_, N17, N21 );
not g215 ( new_n353_, N21 );
and g216 ( new_n354_, new_n186_, new_n353_ );
or g217 ( new_n355_, new_n354_, new_n352_ );
or g218 ( new_n356_, new_n355_, keyIn_0_2 );
not g219 ( new_n357_, keyIn_0_2 );
not g220 ( new_n358_, new_n352_ );
or g221 ( new_n359_, N17, N21 );
and g222 ( new_n360_, new_n358_, new_n359_ );
or g223 ( new_n361_, new_n360_, new_n357_ );
and g224 ( new_n362_, new_n356_, new_n361_ );
and g225 ( new_n363_, N25, N29 );
not g226 ( new_n364_, new_n363_ );
or g227 ( new_n365_, N25, N29 );
and g228 ( new_n366_, new_n364_, keyIn_0_3, new_n365_ );
not g229 ( new_n367_, new_n366_ );
and g230 ( new_n368_, new_n364_, new_n365_ );
or g231 ( new_n369_, new_n368_, keyIn_0_3 );
and g232 ( new_n370_, new_n369_, new_n367_ );
or g233 ( new_n371_, new_n362_, new_n370_ );
and g234 ( new_n372_, new_n356_, new_n361_, new_n369_, new_n367_ );
not g235 ( new_n373_, new_n372_ );
and g236 ( new_n374_, new_n371_, new_n351_, new_n373_ );
and g237 ( new_n375_, new_n360_, new_n357_ );
and g238 ( new_n376_, new_n355_, keyIn_0_2 );
or g239 ( new_n377_, new_n376_, new_n375_ );
not g240 ( new_n378_, keyIn_0_3 );
not g241 ( new_n379_, N25 );
not g242 ( new_n380_, N29 );
and g243 ( new_n381_, new_n379_, new_n380_ );
or g244 ( new_n382_, new_n381_, new_n363_ );
and g245 ( new_n383_, new_n382_, new_n378_ );
or g246 ( new_n384_, new_n383_, new_n366_ );
and g247 ( new_n385_, new_n377_, new_n384_ );
or g248 ( new_n386_, new_n385_, new_n372_ );
and g249 ( new_n387_, new_n386_, keyIn_0_13 );
or g250 ( new_n388_, new_n387_, new_n374_ );
and g251 ( new_n389_, N57, N61 );
not g252 ( new_n390_, N57 );
not g253 ( new_n391_, N61 );
and g254 ( new_n392_, new_n390_, new_n391_ );
or g255 ( new_n393_, new_n392_, new_n389_ );
not g256 ( new_n394_, new_n393_ );
and g257 ( new_n395_, N49, N53 );
not g258 ( new_n396_, N53 );
and g259 ( new_n397_, new_n180_, new_n396_ );
or g260 ( new_n398_, new_n397_, new_n395_ );
not g261 ( new_n399_, new_n398_ );
and g262 ( new_n400_, new_n394_, new_n399_ );
and g263 ( new_n401_, new_n393_, new_n398_ );
or g264 ( new_n402_, new_n400_, new_n401_ );
and g265 ( new_n403_, new_n388_, new_n402_ );
not g266 ( new_n404_, new_n374_ );
and g267 ( new_n405_, new_n371_, new_n373_ );
or g268 ( new_n406_, new_n405_, new_n351_ );
and g269 ( new_n407_, new_n406_, new_n404_ );
not g270 ( new_n408_, new_n402_ );
and g271 ( new_n409_, new_n407_, new_n408_ );
or g272 ( new_n410_, new_n403_, new_n409_ );
not g273 ( new_n411_, new_n410_ );
and g274 ( new_n412_, N136, N137 );
and g275 ( new_n413_, new_n411_, new_n412_ );
not g276 ( new_n414_, new_n413_ );
or g277 ( new_n415_, new_n411_, new_n412_ );
and g278 ( new_n416_, new_n414_, new_n415_ );
and g279 ( new_n417_, N109, N125 );
not g280 ( new_n418_, N109 );
not g281 ( new_n419_, N125 );
and g282 ( new_n420_, new_n418_, new_n419_ );
or g283 ( new_n421_, new_n420_, new_n417_ );
not g284 ( new_n422_, new_n421_ );
and g285 ( new_n423_, N77, N93 );
and g286 ( new_n424_, new_n140_, new_n155_ );
or g287 ( new_n425_, new_n424_, new_n423_ );
not g288 ( new_n426_, new_n425_ );
and g289 ( new_n427_, new_n422_, new_n426_ );
and g290 ( new_n428_, new_n421_, new_n425_ );
or g291 ( new_n429_, new_n427_, new_n428_ );
not g292 ( new_n430_, new_n429_ );
and g293 ( new_n431_, new_n416_, new_n430_ );
not g294 ( new_n432_, new_n431_ );
or g295 ( new_n433_, new_n416_, new_n430_ );
and g296 ( new_n434_, new_n432_, new_n433_ );
not g297 ( new_n435_, new_n434_ );
not g298 ( new_n436_, new_n197_ );
and g299 ( new_n437_, N105, N109 );
and g300 ( new_n438_, new_n295_, new_n418_ );
or g301 ( new_n439_, new_n438_, new_n437_ );
not g302 ( new_n440_, new_n439_ );
and g303 ( new_n441_, N97, N101 );
not g304 ( new_n442_, N97 );
not g305 ( new_n443_, N101 );
and g306 ( new_n444_, new_n442_, new_n443_ );
or g307 ( new_n445_, new_n444_, new_n441_ );
not g308 ( new_n446_, new_n445_ );
and g309 ( new_n447_, new_n440_, new_n446_ );
and g310 ( new_n448_, new_n439_, new_n445_ );
or g311 ( new_n449_, new_n447_, new_n448_ );
not g312 ( new_n450_, new_n449_ );
and g313 ( new_n451_, new_n450_, new_n152_ );
and g314 ( new_n452_, new_n170_, new_n449_ );
or g315 ( new_n453_, new_n451_, new_n452_ );
and g316 ( new_n454_, N131, N137 );
and g317 ( new_n455_, new_n453_, new_n454_ );
not g318 ( new_n456_, new_n455_ );
or g319 ( new_n457_, new_n453_, new_n454_ );
and g320 ( new_n458_, new_n456_, new_n457_ );
and g321 ( new_n459_, N41, N57 );
and g322 ( new_n460_, new_n217_, new_n390_ );
or g323 ( new_n461_, new_n460_, new_n459_ );
not g324 ( new_n462_, new_n461_ );
and g325 ( new_n463_, N9, N25 );
and g326 ( new_n464_, new_n246_, new_n379_ );
or g327 ( new_n465_, new_n464_, new_n463_ );
not g328 ( new_n466_, new_n465_ );
and g329 ( new_n467_, new_n462_, new_n466_ );
and g330 ( new_n468_, new_n461_, new_n465_ );
or g331 ( new_n469_, new_n467_, new_n468_ );
not g332 ( new_n470_, new_n469_ );
and g333 ( new_n471_, new_n458_, new_n470_ );
not g334 ( new_n472_, new_n471_ );
or g335 ( new_n473_, new_n458_, new_n470_ );
and g336 ( new_n474_, new_n472_, new_n473_ );
and g337 ( new_n475_, new_n474_, keyIn_0_24 );
not g338 ( new_n476_, new_n475_ );
or g339 ( new_n477_, new_n476_, new_n436_ );
or g340 ( new_n478_, new_n475_, new_n197_ );
and g341 ( new_n479_, N121, N125 );
and g342 ( new_n480_, new_n296_, new_n419_ );
or g343 ( new_n481_, new_n480_, new_n479_ );
not g344 ( new_n482_, new_n481_ );
and g345 ( new_n483_, N113, N117 );
not g346 ( new_n484_, N113 );
not g347 ( new_n485_, N117 );
and g348 ( new_n486_, new_n484_, new_n485_ );
or g349 ( new_n487_, new_n486_, new_n483_ );
not g350 ( new_n488_, new_n487_ );
and g351 ( new_n489_, new_n482_, new_n488_ );
and g352 ( new_n490_, new_n481_, new_n487_ );
or g353 ( new_n491_, new_n489_, new_n490_ );
not g354 ( new_n492_, new_n491_ );
and g355 ( new_n493_, new_n492_, new_n449_ );
and g356 ( new_n494_, new_n450_, new_n491_ );
or g357 ( new_n495_, new_n493_, new_n494_ );
and g358 ( new_n496_, N130, N137 );
and g359 ( new_n497_, new_n495_, new_n496_ );
not g360 ( new_n498_, new_n497_ );
or g361 ( new_n499_, new_n495_, new_n496_ );
and g362 ( new_n500_, new_n498_, new_n499_ );
and g363 ( new_n501_, N37, N53 );
and g364 ( new_n502_, new_n200_, new_n396_ );
or g365 ( new_n503_, new_n502_, new_n501_ );
not g366 ( new_n504_, new_n503_ );
and g367 ( new_n505_, N5, N21 );
and g368 ( new_n506_, new_n325_, new_n353_ );
or g369 ( new_n507_, new_n506_, new_n505_ );
not g370 ( new_n508_, new_n507_ );
and g371 ( new_n509_, new_n504_, new_n508_ );
and g372 ( new_n510_, new_n503_, new_n507_ );
or g373 ( new_n511_, new_n509_, new_n510_ );
not g374 ( new_n512_, new_n511_ );
and g375 ( new_n513_, new_n500_, new_n512_ );
not g376 ( new_n514_, new_n513_ );
or g377 ( new_n515_, new_n500_, new_n512_ );
and g378 ( new_n516_, new_n514_, new_n515_ );
not g379 ( new_n517_, new_n516_ );
and g380 ( new_n518_, new_n477_, new_n478_, new_n517_ );
not g381 ( new_n519_, new_n474_ );
and g382 ( new_n520_, new_n436_, new_n516_ );
and g383 ( new_n521_, new_n520_, new_n519_ );
or g384 ( new_n522_, new_n518_, new_n521_ );
and g385 ( new_n523_, new_n492_, new_n167_ );
and g386 ( new_n524_, new_n168_, new_n491_ );
or g387 ( new_n525_, new_n523_, new_n524_ );
and g388 ( new_n526_, N132, N137 );
and g389 ( new_n527_, new_n525_, new_n526_ );
not g390 ( new_n528_, new_n527_ );
or g391 ( new_n529_, new_n525_, new_n526_ );
and g392 ( new_n530_, new_n528_, new_n529_ );
and g393 ( new_n531_, N45, N61 );
and g394 ( new_n532_, new_n218_, new_n391_ );
or g395 ( new_n533_, new_n532_, new_n531_ );
not g396 ( new_n534_, new_n533_ );
and g397 ( new_n535_, N13, N29 );
and g398 ( new_n536_, new_n247_, new_n380_ );
or g399 ( new_n537_, new_n536_, new_n535_ );
not g400 ( new_n538_, new_n537_ );
and g401 ( new_n539_, new_n534_, new_n538_ );
and g402 ( new_n540_, new_n533_, new_n537_ );
or g403 ( new_n541_, new_n539_, new_n540_ );
and g404 ( new_n542_, new_n541_, keyIn_0_15 );
not g405 ( new_n543_, new_n542_ );
or g406 ( new_n544_, new_n541_, keyIn_0_15 );
and g407 ( new_n545_, new_n543_, new_n544_ );
and g408 ( new_n546_, new_n530_, new_n545_ );
not g409 ( new_n547_, new_n546_ );
or g410 ( new_n548_, new_n530_, new_n545_ );
and g411 ( new_n549_, new_n547_, new_n548_ );
not g412 ( new_n550_, new_n549_ );
and g413 ( new_n551_, new_n522_, new_n550_ );
and g414 ( new_n552_, new_n519_, new_n549_ );
and g415 ( new_n553_, new_n552_, new_n436_, new_n517_ );
or g416 ( new_n554_, new_n551_, new_n553_ );
and g417 ( new_n555_, new_n350_, new_n435_, new_n554_ );
not g418 ( new_n556_, keyIn_0_20 );
not g419 ( new_n557_, keyIn_0_18 );
or g420 ( new_n558_, new_n263_, new_n407_ );
and g421 ( new_n559_, new_n262_, new_n406_, new_n260_, new_n404_ );
not g422 ( new_n560_, new_n559_ );
and g423 ( new_n561_, new_n558_, new_n560_ );
or g424 ( new_n562_, new_n561_, new_n557_ );
and g425 ( new_n563_, new_n558_, new_n557_, new_n560_ );
not g426 ( new_n564_, new_n563_ );
and g427 ( new_n565_, new_n562_, new_n564_ );
and g428 ( new_n566_, N133, N137 );
or g429 ( new_n567_, new_n566_, keyIn_0_6 );
and g430 ( new_n568_, new_n566_, keyIn_0_6 );
not g431 ( new_n569_, new_n568_ );
and g432 ( new_n570_, new_n569_, new_n567_ );
or g433 ( new_n571_, new_n565_, new_n570_ );
and g434 ( new_n572_, new_n562_, new_n564_, new_n570_ );
not g435 ( new_n573_, new_n572_ );
and g436 ( new_n574_, new_n571_, new_n573_ );
or g437 ( new_n575_, new_n574_, new_n556_ );
and g438 ( new_n576_, new_n571_, new_n556_, new_n573_ );
not g439 ( new_n577_, new_n576_ );
and g440 ( new_n578_, new_n575_, new_n577_ );
not g441 ( new_n579_, keyIn_0_8 );
and g442 ( new_n580_, N65, N81 );
and g443 ( new_n581_, new_n145_, new_n160_ );
or g444 ( new_n582_, new_n581_, new_n580_ );
not g445 ( new_n583_, new_n582_ );
and g446 ( new_n584_, new_n583_, new_n579_ );
and g447 ( new_n585_, new_n582_, keyIn_0_8 );
or g448 ( new_n586_, new_n584_, new_n585_ );
not g449 ( new_n587_, keyIn_0_9 );
and g450 ( new_n588_, N97, N113 );
and g451 ( new_n589_, new_n442_, new_n484_ );
or g452 ( new_n590_, new_n589_, new_n588_ );
not g453 ( new_n591_, new_n590_ );
and g454 ( new_n592_, new_n591_, new_n587_ );
and g455 ( new_n593_, new_n590_, keyIn_0_9 );
or g456 ( new_n594_, new_n592_, new_n593_ );
not g457 ( new_n595_, new_n594_ );
and g458 ( new_n596_, new_n595_, new_n586_ );
not g459 ( new_n597_, new_n596_ );
or g460 ( new_n598_, new_n595_, new_n586_ );
and g461 ( new_n599_, new_n597_, new_n598_ );
not g462 ( new_n600_, new_n599_ );
and g463 ( new_n601_, new_n600_, keyIn_0_16 );
not g464 ( new_n602_, new_n601_ );
or g465 ( new_n603_, new_n600_, keyIn_0_16 );
and g466 ( new_n604_, new_n602_, new_n603_ );
or g467 ( new_n605_, new_n578_, new_n604_ );
and g468 ( new_n606_, new_n575_, new_n577_, new_n604_ );
not g469 ( new_n607_, new_n606_ );
and g470 ( new_n608_, new_n605_, new_n607_ );
or g471 ( new_n609_, new_n608_, keyIn_0_22 );
and g472 ( new_n610_, new_n605_, keyIn_0_22, new_n607_ );
not g473 ( new_n611_, new_n610_ );
and g474 ( new_n612_, new_n609_, new_n611_ );
and g475 ( new_n613_, new_n324_, new_n408_ );
and g476 ( new_n614_, new_n233_, new_n402_ );
or g477 ( new_n615_, new_n614_, new_n613_ );
not g478 ( new_n616_, new_n615_ );
and g479 ( new_n617_, N134, N137 );
and g480 ( new_n618_, new_n616_, new_n617_ );
not g481 ( new_n619_, new_n618_ );
or g482 ( new_n620_, new_n616_, new_n617_ );
and g483 ( new_n621_, new_n619_, new_n620_ );
and g484 ( new_n622_, N101, N117 );
and g485 ( new_n623_, new_n443_, new_n485_ );
or g486 ( new_n624_, new_n623_, new_n622_ );
not g487 ( new_n625_, new_n624_ );
and g488 ( new_n626_, N69, N85 );
and g489 ( new_n627_, new_n146_, new_n161_ );
or g490 ( new_n628_, new_n627_, new_n626_ );
not g491 ( new_n629_, new_n628_ );
and g492 ( new_n630_, new_n625_, new_n629_ );
and g493 ( new_n631_, new_n624_, new_n628_ );
or g494 ( new_n632_, new_n630_, new_n631_ );
not g495 ( new_n633_, new_n632_ );
and g496 ( new_n634_, new_n621_, new_n633_ );
not g497 ( new_n635_, new_n634_ );
or g498 ( new_n636_, new_n621_, new_n633_ );
and g499 ( new_n637_, new_n635_, new_n636_ );
not g500 ( new_n638_, new_n637_ );
and g501 ( new_n639_, new_n612_, new_n638_ );
and g502 ( new_n640_, new_n555_, new_n639_ );
and g503 ( new_n641_, new_n640_, new_n197_ );
not g504 ( new_n642_, new_n641_ );
and g505 ( new_n643_, new_n642_, N1 );
and g506 ( new_n644_, new_n641_, new_n185_ );
or g507 ( N724, new_n643_, new_n644_ );
and g508 ( new_n646_, new_n640_, new_n516_ );
not g509 ( new_n647_, new_n646_ );
and g510 ( new_n648_, new_n647_, N5 );
and g511 ( new_n649_, new_n646_, new_n325_ );
or g512 ( N725, new_n648_, new_n649_ );
and g513 ( new_n651_, new_n640_, new_n474_ );
not g514 ( new_n652_, new_n651_ );
and g515 ( new_n653_, new_n652_, N9 );
and g516 ( new_n654_, new_n651_, new_n246_ );
or g517 ( N726, new_n653_, new_n654_ );
and g518 ( new_n656_, new_n640_, new_n549_ );
not g519 ( new_n657_, new_n656_ );
and g520 ( new_n658_, new_n657_, N13 );
and g521 ( new_n659_, new_n656_, new_n247_ );
or g522 ( N727, new_n658_, new_n659_ );
not g523 ( new_n661_, new_n315_ );
and g524 ( new_n662_, new_n312_, new_n314_ );
or g525 ( new_n663_, new_n662_, keyIn_0_23 );
and g526 ( new_n664_, new_n663_, new_n661_ );
and g527 ( new_n665_, new_n664_, new_n434_, new_n554_ );
and g528 ( new_n666_, new_n665_, new_n639_ );
and g529 ( new_n667_, new_n666_, new_n197_ );
not g530 ( new_n668_, new_n667_ );
and g531 ( new_n669_, new_n668_, N17 );
and g532 ( new_n670_, new_n667_, new_n186_ );
or g533 ( N728, new_n669_, new_n670_ );
and g534 ( new_n672_, new_n666_, new_n516_ );
not g535 ( new_n673_, new_n672_ );
and g536 ( new_n674_, new_n673_, N21 );
and g537 ( new_n675_, new_n672_, new_n353_ );
or g538 ( N729, new_n674_, new_n675_ );
and g539 ( new_n677_, new_n666_, new_n474_ );
not g540 ( new_n678_, new_n677_ );
and g541 ( new_n679_, new_n678_, N25 );
and g542 ( new_n680_, new_n677_, new_n379_ );
or g543 ( N730, new_n679_, new_n680_ );
and g544 ( new_n682_, new_n666_, new_n549_ );
not g545 ( new_n683_, new_n682_ );
and g546 ( new_n684_, new_n683_, N29 );
and g547 ( new_n685_, new_n682_, new_n380_ );
or g548 ( N731, new_n684_, new_n685_ );
not g549 ( new_n687_, keyIn_0_22 );
and g550 ( new_n688_, new_n336_, new_n388_ );
or g551 ( new_n689_, new_n688_, new_n559_ );
and g552 ( new_n690_, new_n689_, keyIn_0_18 );
or g553 ( new_n691_, new_n690_, new_n563_ );
not g554 ( new_n692_, new_n570_ );
and g555 ( new_n693_, new_n691_, new_n692_ );
or g556 ( new_n694_, new_n693_, new_n572_ );
and g557 ( new_n695_, new_n694_, keyIn_0_20 );
or g558 ( new_n696_, new_n695_, new_n576_ );
not g559 ( new_n697_, new_n604_ );
and g560 ( new_n698_, new_n696_, new_n697_ );
or g561 ( new_n699_, new_n698_, new_n606_ );
and g562 ( new_n700_, new_n699_, new_n687_ );
or g563 ( new_n701_, new_n700_, new_n610_ );
and g564 ( new_n702_, new_n701_, new_n637_ );
and g565 ( new_n703_, new_n555_, new_n702_ );
and g566 ( new_n704_, new_n703_, new_n197_ );
not g567 ( new_n705_, new_n704_ );
and g568 ( new_n706_, new_n705_, N33 );
and g569 ( new_n707_, new_n704_, new_n179_ );
or g570 ( N732, new_n706_, new_n707_ );
and g571 ( new_n709_, new_n703_, new_n516_ );
not g572 ( new_n710_, new_n709_ );
and g573 ( new_n711_, new_n710_, N37 );
and g574 ( new_n712_, new_n709_, new_n200_ );
or g575 ( N733, new_n711_, new_n712_ );
and g576 ( new_n714_, new_n703_, new_n474_ );
not g577 ( new_n715_, new_n714_ );
and g578 ( new_n716_, new_n715_, N41 );
and g579 ( new_n717_, new_n714_, new_n217_ );
or g580 ( N734, new_n716_, new_n717_ );
and g581 ( new_n719_, new_n703_, new_n549_ );
not g582 ( new_n720_, new_n719_ );
and g583 ( new_n721_, new_n720_, N45 );
and g584 ( new_n722_, new_n719_, new_n218_ );
or g585 ( N735, new_n721_, new_n722_ );
and g586 ( new_n724_, new_n665_, new_n702_ );
and g587 ( new_n725_, new_n724_, new_n197_ );
not g588 ( new_n726_, new_n725_ );
and g589 ( new_n727_, new_n726_, N49 );
and g590 ( new_n728_, new_n725_, new_n180_ );
or g591 ( N736, new_n727_, new_n728_ );
and g592 ( new_n730_, new_n724_, new_n516_ );
not g593 ( new_n731_, new_n730_ );
and g594 ( new_n732_, new_n731_, N53 );
and g595 ( new_n733_, new_n730_, new_n396_ );
or g596 ( N737, new_n732_, new_n733_ );
and g597 ( new_n735_, new_n724_, new_n474_ );
not g598 ( new_n736_, new_n735_ );
and g599 ( new_n737_, new_n736_, N57 );
and g600 ( new_n738_, new_n735_, new_n390_ );
or g601 ( N738, new_n737_, new_n738_ );
and g602 ( new_n740_, new_n724_, new_n549_ );
not g603 ( new_n741_, new_n740_ );
and g604 ( new_n742_, new_n741_, N61 );
and g605 ( new_n743_, new_n740_, new_n391_ );
or g606 ( N739, new_n742_, new_n743_ );
not g607 ( new_n745_, keyIn_0_52 );
not g608 ( new_n746_, keyIn_0_40 );
not g609 ( new_n747_, keyIn_0_37 );
not g610 ( new_n748_, keyIn_0_36 );
not g611 ( new_n749_, keyIn_0_32 );
not g612 ( new_n750_, keyIn_0_27 );
or g613 ( new_n751_, new_n349_, new_n750_, new_n315_ );
and g614 ( new_n752_, new_n637_, keyIn_0_26 );
not g615 ( new_n753_, new_n752_ );
or g616 ( new_n754_, new_n637_, keyIn_0_26 );
and g617 ( new_n755_, new_n751_, new_n434_, new_n753_, new_n754_ );
or g618 ( new_n756_, new_n701_, keyIn_0_25 );
and g619 ( new_n757_, new_n701_, keyIn_0_25 );
not g620 ( new_n758_, new_n757_ );
or g621 ( new_n759_, new_n664_, keyIn_0_27 );
and g622 ( new_n760_, new_n755_, new_n756_, new_n758_, new_n759_ );
or g623 ( new_n761_, new_n760_, new_n749_ );
and g624 ( new_n762_, new_n663_, new_n661_, keyIn_0_27 );
not g625 ( new_n763_, new_n754_ );
or g626 ( new_n764_, new_n763_, new_n435_, new_n752_ );
or g627 ( new_n765_, new_n762_, new_n764_ );
not g628 ( new_n766_, new_n756_ );
and g629 ( new_n767_, new_n350_, new_n750_ );
or g630 ( new_n768_, new_n767_, new_n757_ );
or g631 ( new_n769_, new_n768_, keyIn_0_32, new_n765_, new_n766_ );
and g632 ( new_n770_, new_n761_, new_n769_ );
not g633 ( new_n771_, new_n770_ );
not g634 ( new_n772_, keyIn_0_29 );
and g635 ( new_n773_, new_n612_, new_n772_ );
and g636 ( new_n774_, new_n701_, keyIn_0_29 );
or g637 ( new_n775_, new_n773_, new_n774_ );
not g638 ( new_n776_, new_n775_ );
not g639 ( new_n777_, keyIn_0_30 );
and g640 ( new_n778_, new_n664_, new_n777_ );
and g641 ( new_n779_, new_n350_, keyIn_0_30 );
or g642 ( new_n780_, new_n778_, new_n779_, new_n434_, new_n638_ );
or g643 ( new_n781_, new_n780_, keyIn_0_34, new_n776_ );
not g644 ( new_n782_, keyIn_0_34 );
not g645 ( new_n783_, new_n778_ );
not g646 ( new_n784_, new_n779_ );
and g647 ( new_n785_, new_n435_, new_n637_ );
and g648 ( new_n786_, new_n775_, new_n783_, new_n784_, new_n785_ );
or g649 ( new_n787_, new_n786_, new_n782_ );
and g650 ( new_n788_, new_n787_, new_n781_ );
not g651 ( new_n789_, new_n788_ );
not g652 ( new_n790_, keyIn_0_35 );
not g653 ( new_n791_, keyIn_0_31 );
and g654 ( new_n792_, new_n350_, new_n791_ );
and g655 ( new_n793_, new_n663_, new_n661_, keyIn_0_31 );
or g656 ( new_n794_, new_n792_, new_n793_ );
or g657 ( new_n795_, new_n701_, new_n434_, new_n637_ );
not g658 ( new_n796_, new_n795_ );
and g659 ( new_n797_, new_n794_, new_n796_ );
or g660 ( new_n798_, new_n797_, new_n790_ );
not g661 ( new_n799_, new_n792_ );
not g662 ( new_n800_, new_n793_ );
and g663 ( new_n801_, new_n799_, new_n800_ );
or g664 ( new_n802_, new_n801_, new_n795_, keyIn_0_35 );
and g665 ( new_n803_, new_n798_, new_n802_ );
not g666 ( new_n804_, new_n803_ );
not g667 ( new_n805_, keyIn_0_28 );
and g668 ( new_n806_, new_n609_, new_n805_, new_n611_ );
and g669 ( new_n807_, new_n701_, keyIn_0_28 );
or g670 ( new_n808_, new_n807_, new_n806_ );
and g671 ( new_n809_, new_n350_, new_n435_, new_n638_ );
and g672 ( new_n810_, new_n808_, new_n809_ );
or g673 ( new_n811_, new_n810_, keyIn_0_33 );
not g674 ( new_n812_, keyIn_0_33 );
not g675 ( new_n813_, new_n808_ );
not g676 ( new_n814_, new_n809_ );
or g677 ( new_n815_, new_n813_, new_n812_, new_n814_ );
and g678 ( new_n816_, new_n811_, new_n815_ );
not g679 ( new_n817_, new_n816_ );
and g680 ( new_n818_, new_n804_, new_n817_ );
and g681 ( new_n819_, new_n818_, new_n748_, new_n771_, new_n789_ );
or g682 ( new_n820_, new_n788_, new_n803_, new_n816_, new_n770_ );
and g683 ( new_n821_, new_n820_, keyIn_0_36 );
or g684 ( new_n822_, new_n821_, new_n819_ );
and g685 ( new_n823_, new_n517_, new_n197_ );
and g686 ( new_n824_, new_n550_, new_n474_ );
and g687 ( new_n825_, new_n823_, new_n824_ );
and g688 ( new_n826_, new_n822_, new_n825_ );
or g689 ( new_n827_, new_n826_, new_n747_ );
not g690 ( new_n828_, new_n822_ );
not g691 ( new_n829_, new_n825_ );
or g692 ( new_n830_, new_n828_, keyIn_0_37, new_n829_ );
and g693 ( new_n831_, new_n827_, new_n830_ );
or g694 ( new_n832_, new_n831_, new_n701_ );
and g695 ( new_n833_, new_n832_, new_n746_ );
not g696 ( new_n834_, new_n831_ );
and g697 ( new_n835_, new_n834_, keyIn_0_40, new_n612_ );
or g698 ( new_n836_, new_n833_, new_n835_ );
and g699 ( new_n837_, new_n836_, N65 );
not g700 ( new_n838_, new_n837_ );
not g701 ( new_n839_, new_n833_ );
not g702 ( new_n840_, new_n835_ );
and g703 ( new_n841_, new_n839_, new_n145_, new_n840_ );
not g704 ( new_n842_, new_n841_ );
and g705 ( new_n843_, new_n838_, new_n745_, new_n842_ );
or g706 ( new_n844_, new_n837_, new_n841_ );
and g707 ( new_n845_, new_n844_, keyIn_0_52 );
or g708 ( N740, new_n845_, new_n843_ );
not g709 ( new_n847_, keyIn_0_53 );
not g710 ( new_n848_, keyIn_0_41 );
or g711 ( new_n849_, new_n831_, new_n638_ );
and g712 ( new_n850_, new_n849_, new_n848_ );
and g713 ( new_n851_, new_n834_, keyIn_0_41, new_n637_ );
or g714 ( new_n852_, new_n850_, new_n851_ );
and g715 ( new_n853_, new_n852_, N69 );
not g716 ( new_n854_, new_n853_ );
not g717 ( new_n855_, new_n850_ );
not g718 ( new_n856_, new_n851_ );
and g719 ( new_n857_, new_n855_, new_n146_, new_n856_ );
not g720 ( new_n858_, new_n857_ );
and g721 ( new_n859_, new_n854_, new_n847_, new_n858_ );
or g722 ( new_n860_, new_n853_, new_n857_ );
and g723 ( new_n861_, new_n860_, keyIn_0_53 );
or g724 ( N741, new_n861_, new_n859_ );
not g725 ( new_n863_, keyIn_0_54 );
not g726 ( new_n864_, keyIn_0_42 );
or g727 ( new_n865_, new_n831_, new_n664_ );
and g728 ( new_n866_, new_n865_, new_n864_ );
and g729 ( new_n867_, new_n834_, keyIn_0_42, new_n350_ );
or g730 ( new_n868_, new_n866_, new_n867_ );
and g731 ( new_n869_, new_n868_, N73 );
not g732 ( new_n870_, new_n869_ );
not g733 ( new_n871_, new_n866_ );
not g734 ( new_n872_, new_n867_ );
and g735 ( new_n873_, new_n871_, new_n139_, new_n872_ );
not g736 ( new_n874_, new_n873_ );
and g737 ( new_n875_, new_n870_, new_n863_, new_n874_ );
or g738 ( new_n876_, new_n869_, new_n873_ );
and g739 ( new_n877_, new_n876_, keyIn_0_54 );
or g740 ( N742, new_n877_, new_n875_ );
not g741 ( new_n879_, keyIn_0_55 );
not g742 ( new_n880_, keyIn_0_43 );
or g743 ( new_n881_, new_n831_, new_n435_ );
and g744 ( new_n882_, new_n881_, new_n880_ );
and g745 ( new_n883_, new_n834_, keyIn_0_43, new_n434_ );
or g746 ( new_n884_, new_n882_, new_n883_ );
and g747 ( new_n885_, new_n884_, N77 );
not g748 ( new_n886_, new_n885_ );
not g749 ( new_n887_, new_n882_ );
not g750 ( new_n888_, new_n883_ );
and g751 ( new_n889_, new_n887_, new_n140_, new_n888_ );
not g752 ( new_n890_, new_n889_ );
and g753 ( new_n891_, new_n886_, new_n879_, new_n890_ );
or g754 ( new_n892_, new_n885_, new_n889_ );
and g755 ( new_n893_, new_n892_, keyIn_0_55 );
or g756 ( N743, new_n893_, new_n891_ );
not g757 ( new_n895_, keyIn_0_44 );
and g758 ( new_n896_, new_n552_, new_n823_ );
and g759 ( new_n897_, new_n822_, new_n896_ );
or g760 ( new_n898_, new_n897_, keyIn_0_38 );
not g761 ( new_n899_, keyIn_0_38 );
not g762 ( new_n900_, new_n896_ );
or g763 ( new_n901_, new_n828_, new_n899_, new_n900_ );
and g764 ( new_n902_, new_n898_, new_n901_ );
or g765 ( new_n903_, new_n902_, new_n701_ );
and g766 ( new_n904_, new_n903_, new_n895_ );
not g767 ( new_n905_, new_n902_ );
and g768 ( new_n906_, new_n905_, keyIn_0_44, new_n612_ );
or g769 ( new_n907_, new_n904_, new_n906_ );
and g770 ( new_n908_, new_n907_, N81 );
not g771 ( new_n909_, new_n908_ );
not g772 ( new_n910_, new_n904_ );
not g773 ( new_n911_, new_n906_ );
and g774 ( new_n912_, new_n910_, new_n160_, new_n911_ );
not g775 ( new_n913_, new_n912_ );
and g776 ( new_n914_, new_n909_, keyIn_0_56, new_n913_ );
not g777 ( new_n915_, keyIn_0_56 );
or g778 ( new_n916_, new_n908_, new_n912_ );
and g779 ( new_n917_, new_n916_, new_n915_ );
or g780 ( N744, new_n917_, new_n914_ );
not g781 ( new_n919_, keyIn_0_57 );
not g782 ( new_n920_, keyIn_0_45 );
or g783 ( new_n921_, new_n902_, new_n638_ );
and g784 ( new_n922_, new_n921_, new_n920_ );
and g785 ( new_n923_, new_n905_, keyIn_0_45, new_n637_ );
or g786 ( new_n924_, new_n922_, new_n923_ );
and g787 ( new_n925_, new_n924_, N85 );
not g788 ( new_n926_, new_n925_ );
not g789 ( new_n927_, new_n922_ );
not g790 ( new_n928_, new_n923_ );
and g791 ( new_n929_, new_n927_, new_n161_, new_n928_ );
not g792 ( new_n930_, new_n929_ );
and g793 ( new_n931_, new_n926_, new_n919_, new_n930_ );
or g794 ( new_n932_, new_n925_, new_n929_ );
and g795 ( new_n933_, new_n932_, keyIn_0_57 );
or g796 ( N745, new_n933_, new_n931_ );
not g797 ( new_n935_, keyIn_0_46 );
or g798 ( new_n936_, new_n902_, new_n664_ );
and g799 ( new_n937_, new_n936_, new_n935_ );
and g800 ( new_n938_, new_n905_, keyIn_0_46, new_n350_ );
or g801 ( new_n939_, new_n937_, new_n938_ );
and g802 ( new_n940_, new_n939_, N89 );
not g803 ( new_n941_, new_n940_ );
not g804 ( new_n942_, new_n937_ );
not g805 ( new_n943_, new_n938_ );
and g806 ( new_n944_, new_n942_, new_n154_, new_n943_ );
not g807 ( new_n945_, new_n944_ );
and g808 ( new_n946_, new_n941_, keyIn_0_58, new_n945_ );
not g809 ( new_n947_, keyIn_0_58 );
or g810 ( new_n948_, new_n940_, new_n944_ );
and g811 ( new_n949_, new_n948_, new_n947_ );
or g812 ( N746, new_n949_, new_n946_ );
not g813 ( new_n951_, keyIn_0_59 );
not g814 ( new_n952_, keyIn_0_47 );
or g815 ( new_n953_, new_n902_, new_n435_ );
and g816 ( new_n954_, new_n953_, new_n952_ );
and g817 ( new_n955_, new_n905_, keyIn_0_47, new_n434_ );
or g818 ( new_n956_, new_n954_, new_n955_ );
and g819 ( new_n957_, new_n956_, N93 );
not g820 ( new_n958_, new_n957_ );
not g821 ( new_n959_, new_n954_ );
not g822 ( new_n960_, new_n955_ );
and g823 ( new_n961_, new_n959_, new_n155_, new_n960_ );
not g824 ( new_n962_, new_n961_ );
and g825 ( new_n963_, new_n958_, new_n951_, new_n962_ );
or g826 ( new_n964_, new_n957_, new_n961_ );
and g827 ( new_n965_, new_n964_, keyIn_0_59 );
or g828 ( N747, new_n965_, new_n963_ );
not g829 ( new_n967_, keyIn_0_48 );
not g830 ( new_n968_, keyIn_0_39 );
and g831 ( new_n969_, new_n520_, new_n824_ );
and g832 ( new_n970_, new_n822_, new_n969_ );
or g833 ( new_n971_, new_n970_, new_n968_ );
not g834 ( new_n972_, new_n969_ );
or g835 ( new_n973_, new_n828_, keyIn_0_39, new_n972_ );
and g836 ( new_n974_, new_n971_, new_n973_ );
or g837 ( new_n975_, new_n974_, new_n701_ );
and g838 ( new_n976_, new_n975_, new_n967_ );
not g839 ( new_n977_, new_n974_ );
and g840 ( new_n978_, new_n977_, keyIn_0_48, new_n612_ );
or g841 ( new_n979_, new_n976_, new_n978_ );
and g842 ( new_n980_, new_n979_, N97 );
not g843 ( new_n981_, new_n980_ );
not g844 ( new_n982_, new_n976_ );
not g845 ( new_n983_, new_n978_ );
and g846 ( new_n984_, new_n982_, new_n442_, new_n983_ );
not g847 ( new_n985_, new_n984_ );
and g848 ( new_n986_, new_n981_, keyIn_0_60, new_n985_ );
not g849 ( new_n987_, keyIn_0_60 );
or g850 ( new_n988_, new_n980_, new_n984_ );
and g851 ( new_n989_, new_n988_, new_n987_ );
or g852 ( N748, new_n989_, new_n986_ );
not g853 ( new_n991_, keyIn_0_49 );
or g854 ( new_n992_, new_n974_, new_n638_ );
and g855 ( new_n993_, new_n992_, new_n991_ );
and g856 ( new_n994_, new_n977_, keyIn_0_49, new_n637_ );
or g857 ( new_n995_, new_n993_, new_n994_ );
and g858 ( new_n996_, new_n995_, N101 );
not g859 ( new_n997_, new_n996_ );
not g860 ( new_n998_, new_n993_ );
not g861 ( new_n999_, new_n994_ );
and g862 ( new_n1000_, new_n998_, new_n443_, new_n999_ );
not g863 ( new_n1001_, new_n1000_ );
and g864 ( new_n1002_, new_n997_, keyIn_0_61, new_n1001_ );
not g865 ( new_n1003_, keyIn_0_61 );
or g866 ( new_n1004_, new_n996_, new_n1000_ );
and g867 ( new_n1005_, new_n1004_, new_n1003_ );
or g868 ( N749, new_n1005_, new_n1002_ );
not g869 ( new_n1007_, keyIn_0_50 );
or g870 ( new_n1008_, new_n974_, new_n664_ );
and g871 ( new_n1009_, new_n1008_, new_n1007_ );
and g872 ( new_n1010_, new_n977_, keyIn_0_50, new_n350_ );
or g873 ( new_n1011_, new_n1009_, new_n1010_ );
and g874 ( new_n1012_, new_n1011_, N105 );
not g875 ( new_n1013_, new_n1012_ );
not g876 ( new_n1014_, new_n1009_ );
not g877 ( new_n1015_, new_n1010_ );
and g878 ( new_n1016_, new_n1014_, new_n295_, new_n1015_ );
not g879 ( new_n1017_, new_n1016_ );
and g880 ( new_n1018_, new_n1013_, keyIn_0_62, new_n1017_ );
not g881 ( new_n1019_, keyIn_0_62 );
or g882 ( new_n1020_, new_n1012_, new_n1016_ );
and g883 ( new_n1021_, new_n1020_, new_n1019_ );
or g884 ( N750, new_n1021_, new_n1018_ );
not g885 ( new_n1023_, keyIn_0_63 );
not g886 ( new_n1024_, keyIn_0_51 );
or g887 ( new_n1025_, new_n974_, new_n435_ );
and g888 ( new_n1026_, new_n1025_, new_n1024_ );
and g889 ( new_n1027_, new_n977_, keyIn_0_51, new_n434_ );
or g890 ( new_n1028_, new_n1026_, new_n1027_ );
and g891 ( new_n1029_, new_n1028_, new_n418_ );
not g892 ( new_n1030_, new_n1029_ );
not g893 ( new_n1031_, new_n1026_ );
not g894 ( new_n1032_, new_n1027_ );
and g895 ( new_n1033_, new_n1031_, N109, new_n1032_ );
not g896 ( new_n1034_, new_n1033_ );
and g897 ( new_n1035_, new_n1030_, new_n1023_, new_n1034_ );
or g898 ( new_n1036_, new_n1029_, new_n1033_ );
and g899 ( new_n1037_, new_n1036_, keyIn_0_63 );
or g900 ( N751, new_n1037_, new_n1035_ );
and g901 ( new_n1039_, new_n822_, new_n521_, new_n549_ );
and g902 ( new_n1040_, new_n1039_, new_n612_ );
not g903 ( new_n1041_, new_n1040_ );
and g904 ( new_n1042_, new_n1041_, N113 );
and g905 ( new_n1043_, new_n1040_, new_n484_ );
or g906 ( N752, new_n1042_, new_n1043_ );
and g907 ( new_n1045_, new_n1039_, new_n637_ );
not g908 ( new_n1046_, new_n1045_ );
and g909 ( new_n1047_, new_n1046_, N117 );
and g910 ( new_n1048_, new_n1045_, new_n485_ );
or g911 ( N753, new_n1047_, new_n1048_ );
and g912 ( new_n1050_, new_n1039_, new_n350_ );
not g913 ( new_n1051_, new_n1050_ );
and g914 ( new_n1052_, new_n1051_, N121 );
and g915 ( new_n1053_, new_n1050_, new_n296_ );
or g916 ( N754, new_n1052_, new_n1053_ );
and g917 ( new_n1055_, new_n1039_, new_n434_ );
not g918 ( new_n1056_, new_n1055_ );
and g919 ( new_n1057_, new_n1056_, N125 );
and g920 ( new_n1058_, new_n1055_, new_n419_ );
or g921 ( N755, new_n1057_, new_n1058_ );
endmodule