module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n170_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n1120_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n959_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1082_, new_n849_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n167_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n708_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n1028_, new_n508_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1113_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n140_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n1109_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n749_, new_n861_, new_n1095_, new_n310_, new_n144_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1118_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n1001_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1088_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n1122_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n138_, N1 );
nand g001 ( new_n139_, N81, N85 );
not g002 ( new_n140_, new_n139_ );
nor g003 ( new_n141_, N81, N85 );
nor g004 ( new_n142_, new_n140_, new_n141_ );
not g005 ( new_n143_, new_n142_ );
nand g006 ( new_n144_, N89, N93 );
not g007 ( new_n145_, new_n144_ );
nor g008 ( new_n146_, N89, N93 );
nor g009 ( new_n147_, new_n145_, new_n146_ );
not g010 ( new_n148_, new_n147_ );
nor g011 ( new_n149_, new_n143_, new_n148_ );
nor g012 ( new_n150_, new_n142_, new_n147_ );
nor g013 ( new_n151_, new_n149_, new_n150_ );
nand g014 ( new_n152_, N65, N69 );
not g015 ( new_n153_, new_n152_ );
nor g016 ( new_n154_, N65, N69 );
nor g017 ( new_n155_, new_n153_, new_n154_ );
not g018 ( new_n156_, new_n155_ );
nand g019 ( new_n157_, new_n156_, keyIn_0_5 );
not g020 ( new_n158_, keyIn_0_5 );
nand g021 ( new_n159_, new_n155_, new_n158_ );
nand g022 ( new_n160_, new_n157_, new_n159_ );
nand g023 ( new_n161_, N73, N77 );
not g024 ( new_n162_, new_n161_ );
nor g025 ( new_n163_, N73, N77 );
nor g026 ( new_n164_, new_n162_, new_n163_ );
not g027 ( new_n165_, new_n164_ );
nand g028 ( new_n166_, new_n165_, keyIn_0_6 );
not g029 ( new_n167_, keyIn_0_6 );
nand g030 ( new_n168_, new_n164_, new_n167_ );
nand g031 ( new_n169_, new_n166_, new_n168_ );
nand g032 ( new_n170_, new_n160_, new_n169_ );
not g033 ( new_n171_, new_n170_ );
nor g034 ( new_n172_, new_n160_, new_n169_ );
nor g035 ( new_n173_, new_n171_, new_n172_ );
not g036 ( new_n174_, new_n173_ );
nor g037 ( new_n175_, new_n174_, new_n151_ );
not g038 ( new_n176_, new_n151_ );
nor g039 ( new_n177_, new_n173_, new_n176_ );
nor g040 ( new_n178_, new_n175_, new_n177_ );
not g041 ( new_n179_, new_n178_ );
nand g042 ( new_n180_, N129, N137 );
not g043 ( new_n181_, new_n180_ );
nor g044 ( new_n182_, new_n179_, new_n181_ );
nor g045 ( new_n183_, new_n178_, new_n180_ );
nor g046 ( new_n184_, new_n182_, new_n183_ );
not g047 ( new_n185_, new_n184_ );
nand g048 ( new_n186_, N33, N49 );
not g049 ( new_n187_, new_n186_ );
nor g050 ( new_n188_, N33, N49 );
nor g051 ( new_n189_, new_n187_, new_n188_ );
nand g052 ( new_n190_, N1, N17 );
not g053 ( new_n191_, new_n190_ );
nor g054 ( new_n192_, N1, N17 );
nor g055 ( new_n193_, new_n191_, new_n192_ );
not g056 ( new_n194_, new_n193_ );
nor g057 ( new_n195_, new_n194_, new_n189_ );
nand g058 ( new_n196_, new_n194_, new_n189_ );
not g059 ( new_n197_, new_n196_ );
nor g060 ( new_n198_, new_n197_, new_n195_ );
nor g061 ( new_n199_, new_n185_, new_n198_ );
nand g062 ( new_n200_, new_n185_, new_n198_ );
not g063 ( new_n201_, new_n200_ );
nor g064 ( new_n202_, new_n201_, new_n199_ );
not g065 ( new_n203_, new_n202_ );
not g066 ( new_n204_, keyIn_0_23 );
nand g067 ( new_n205_, N132, N137 );
not g068 ( new_n206_, new_n205_ );
not g069 ( new_n207_, keyIn_0_19 );
nor g070 ( new_n208_, N121, N125 );
nand g071 ( new_n209_, N121, N125 );
not g072 ( new_n210_, new_n209_ );
nor g073 ( new_n211_, new_n210_, new_n208_ );
not g074 ( new_n212_, N113 );
nor g075 ( new_n213_, new_n212_, N117 );
not g076 ( new_n214_, new_n213_ );
not g077 ( new_n215_, N117 );
nor g078 ( new_n216_, new_n215_, N113 );
not g079 ( new_n217_, new_n216_ );
nand g080 ( new_n218_, new_n214_, new_n217_ );
nand g081 ( new_n219_, new_n218_, keyIn_0_7 );
not g082 ( new_n220_, new_n219_ );
nor g083 ( new_n221_, new_n218_, keyIn_0_7 );
nor g084 ( new_n222_, new_n220_, new_n221_ );
nand g085 ( new_n223_, new_n222_, new_n211_ );
not g086 ( new_n224_, new_n211_ );
not g087 ( new_n225_, keyIn_0_7 );
not g088 ( new_n226_, new_n218_ );
nand g089 ( new_n227_, new_n226_, new_n225_ );
nand g090 ( new_n228_, new_n227_, new_n219_ );
nand g091 ( new_n229_, new_n228_, new_n224_ );
nand g092 ( new_n230_, new_n223_, new_n229_ );
nand g093 ( new_n231_, new_n230_, new_n207_ );
nor g094 ( new_n232_, new_n228_, new_n224_ );
nor g095 ( new_n233_, new_n222_, new_n211_ );
nor g096 ( new_n234_, new_n233_, new_n232_ );
nand g097 ( new_n235_, new_n234_, keyIn_0_19 );
nand g098 ( new_n236_, new_n235_, new_n231_ );
nand g099 ( new_n237_, new_n236_, new_n151_ );
not g100 ( new_n238_, new_n231_ );
nor g101 ( new_n239_, new_n230_, new_n207_ );
nor g102 ( new_n240_, new_n238_, new_n239_ );
nand g103 ( new_n241_, new_n240_, new_n176_ );
nand g104 ( new_n242_, new_n241_, new_n237_ );
nand g105 ( new_n243_, new_n242_, keyIn_0_9 );
not g106 ( new_n244_, new_n243_ );
nor g107 ( new_n245_, new_n242_, keyIn_0_9 );
nor g108 ( new_n246_, new_n244_, new_n245_ );
nand g109 ( new_n247_, new_n246_, new_n206_ );
not g110 ( new_n248_, keyIn_0_9 );
not g111 ( new_n249_, new_n237_ );
nor g112 ( new_n250_, new_n236_, new_n151_ );
nor g113 ( new_n251_, new_n249_, new_n250_ );
nand g114 ( new_n252_, new_n251_, new_n248_ );
nand g115 ( new_n253_, new_n252_, new_n243_ );
nand g116 ( new_n254_, new_n253_, new_n205_ );
nand g117 ( new_n255_, new_n247_, new_n254_ );
nand g118 ( new_n256_, new_n255_, new_n204_ );
nor g119 ( new_n257_, new_n253_, new_n205_ );
not g120 ( new_n258_, new_n254_ );
nor g121 ( new_n259_, new_n258_, new_n257_ );
nand g122 ( new_n260_, new_n259_, keyIn_0_23 );
nand g123 ( new_n261_, new_n260_, new_n256_ );
nand g124 ( new_n262_, N13, N29 );
not g125 ( new_n263_, new_n262_ );
nor g126 ( new_n264_, N13, N29 );
nor g127 ( new_n265_, new_n263_, new_n264_ );
not g128 ( new_n266_, new_n265_ );
nor g129 ( new_n267_, new_n266_, keyIn_0_14 );
nand g130 ( new_n268_, new_n266_, keyIn_0_14 );
not g131 ( new_n269_, new_n268_ );
nor g132 ( new_n270_, new_n269_, new_n267_ );
not g133 ( new_n271_, new_n270_ );
not g134 ( new_n272_, N45 );
nor g135 ( new_n273_, new_n272_, N61 );
not g136 ( new_n274_, N61 );
nor g137 ( new_n275_, new_n274_, N45 );
nor g138 ( new_n276_, new_n273_, new_n275_ );
not g139 ( new_n277_, new_n276_ );
nor g140 ( new_n278_, new_n271_, new_n277_ );
nor g141 ( new_n279_, new_n270_, new_n276_ );
nor g142 ( new_n280_, new_n278_, new_n279_ );
nand g143 ( new_n281_, new_n261_, new_n280_ );
not g144 ( new_n282_, new_n281_ );
nor g145 ( new_n283_, new_n261_, new_n280_ );
nor g146 ( new_n284_, new_n282_, new_n283_ );
nand g147 ( new_n285_, N97, N101 );
not g148 ( new_n286_, new_n285_ );
nor g149 ( new_n287_, N97, N101 );
nor g150 ( new_n288_, new_n286_, new_n287_ );
nand g151 ( new_n289_, N105, N109 );
not g152 ( new_n290_, new_n289_ );
nor g153 ( new_n291_, N105, N109 );
nor g154 ( new_n292_, new_n290_, new_n291_ );
nand g155 ( new_n293_, new_n288_, new_n292_ );
not g156 ( new_n294_, new_n288_ );
not g157 ( new_n295_, new_n292_ );
nand g158 ( new_n296_, new_n294_, new_n295_ );
nand g159 ( new_n297_, new_n296_, new_n293_ );
nand g160 ( new_n298_, new_n297_, keyIn_0_18 );
not g161 ( new_n299_, new_n298_ );
nor g162 ( new_n300_, new_n297_, keyIn_0_18 );
nor g163 ( new_n301_, new_n299_, new_n300_ );
nand g164 ( new_n302_, new_n236_, new_n301_ );
not g165 ( new_n303_, new_n301_ );
nand g166 ( new_n304_, new_n240_, new_n303_ );
nand g167 ( new_n305_, new_n304_, new_n302_ );
nand g168 ( new_n306_, new_n305_, keyIn_0_22 );
not g169 ( new_n307_, keyIn_0_22 );
not g170 ( new_n308_, new_n302_ );
nor g171 ( new_n309_, new_n236_, new_n301_ );
nor g172 ( new_n310_, new_n308_, new_n309_ );
nand g173 ( new_n311_, new_n310_, new_n307_ );
nand g174 ( new_n312_, new_n311_, new_n306_ );
nand g175 ( new_n313_, new_n312_, keyIn_0_8 );
not g176 ( new_n314_, keyIn_0_8 );
nor g177 ( new_n315_, new_n310_, new_n307_ );
nor g178 ( new_n316_, new_n305_, keyIn_0_22 );
nor g179 ( new_n317_, new_n315_, new_n316_ );
nand g180 ( new_n318_, new_n317_, new_n314_ );
nand g181 ( new_n319_, new_n318_, new_n313_ );
nand g182 ( new_n320_, N130, N137 );
nand g183 ( new_n321_, new_n319_, new_n320_ );
nor g184 ( new_n322_, new_n317_, new_n314_ );
nor g185 ( new_n323_, new_n312_, keyIn_0_8 );
nor g186 ( new_n324_, new_n322_, new_n323_ );
not g187 ( new_n325_, new_n320_ );
nand g188 ( new_n326_, new_n324_, new_n325_ );
nand g189 ( new_n327_, new_n326_, new_n321_ );
nand g190 ( new_n328_, N37, N53 );
not g191 ( new_n329_, new_n328_ );
nor g192 ( new_n330_, N37, N53 );
nor g193 ( new_n331_, new_n329_, new_n330_ );
not g194 ( new_n332_, new_n331_ );
nor g195 ( new_n333_, new_n332_, keyIn_0_13 );
nand g196 ( new_n334_, new_n332_, keyIn_0_13 );
not g197 ( new_n335_, new_n334_ );
nor g198 ( new_n336_, new_n335_, new_n333_ );
nand g199 ( new_n337_, N5, N21 );
not g200 ( new_n338_, new_n337_ );
nor g201 ( new_n339_, N5, N21 );
nor g202 ( new_n340_, new_n338_, new_n339_ );
not g203 ( new_n341_, new_n340_ );
nor g204 ( new_n342_, new_n341_, keyIn_0_12 );
nand g205 ( new_n343_, new_n341_, keyIn_0_12 );
not g206 ( new_n344_, new_n343_ );
nor g207 ( new_n345_, new_n344_, new_n342_ );
not g208 ( new_n346_, new_n345_ );
nor g209 ( new_n347_, new_n346_, new_n336_ );
nand g210 ( new_n348_, new_n346_, new_n336_ );
not g211 ( new_n349_, new_n348_ );
nor g212 ( new_n350_, new_n349_, new_n347_ );
nand g213 ( new_n351_, new_n327_, new_n350_ );
nor g214 ( new_n352_, new_n324_, new_n325_ );
nor g215 ( new_n353_, new_n319_, new_n320_ );
nor g216 ( new_n354_, new_n352_, new_n353_ );
not g217 ( new_n355_, new_n350_ );
nand g218 ( new_n356_, new_n354_, new_n355_ );
nand g219 ( new_n357_, new_n356_, new_n351_ );
not g220 ( new_n358_, keyIn_0_24 );
nand g221 ( new_n359_, new_n174_, new_n301_ );
nand g222 ( new_n360_, new_n303_, new_n173_ );
nand g223 ( new_n361_, new_n359_, new_n360_ );
nand g224 ( new_n362_, N131, N137 );
not g225 ( new_n363_, new_n362_ );
nand g226 ( new_n364_, new_n361_, new_n363_ );
not g227 ( new_n365_, new_n364_ );
nor g228 ( new_n366_, new_n361_, new_n363_ );
nor g229 ( new_n367_, new_n365_, new_n366_ );
not g230 ( new_n368_, new_n367_ );
nand g231 ( new_n369_, N9, N25 );
not g232 ( new_n370_, new_n369_ );
nor g233 ( new_n371_, N9, N25 );
nor g234 ( new_n372_, new_n370_, new_n371_ );
not g235 ( new_n373_, new_n372_ );
nand g236 ( new_n374_, N41, N57 );
not g237 ( new_n375_, new_n374_ );
nor g238 ( new_n376_, N41, N57 );
nor g239 ( new_n377_, new_n375_, new_n376_ );
not g240 ( new_n378_, new_n377_ );
nor g241 ( new_n379_, new_n373_, new_n378_ );
nor g242 ( new_n380_, new_n372_, new_n377_ );
nor g243 ( new_n381_, new_n379_, new_n380_ );
nor g244 ( new_n382_, new_n368_, new_n381_ );
nand g245 ( new_n383_, new_n368_, new_n381_ );
not g246 ( new_n384_, new_n383_ );
nor g247 ( new_n385_, new_n384_, new_n382_ );
nand g248 ( new_n386_, new_n385_, new_n358_ );
not g249 ( new_n387_, new_n382_ );
nand g250 ( new_n388_, new_n387_, new_n383_ );
nand g251 ( new_n389_, new_n388_, keyIn_0_24 );
nand g252 ( new_n390_, new_n386_, new_n389_ );
nand g253 ( new_n391_, new_n357_, new_n390_ );
nor g254 ( new_n392_, new_n203_, keyIn_0_25 );
nand g255 ( new_n393_, new_n203_, keyIn_0_25 );
not g256 ( new_n394_, new_n393_ );
nor g257 ( new_n395_, new_n394_, new_n392_ );
not g258 ( new_n396_, new_n395_ );
nor g259 ( new_n397_, new_n391_, new_n396_ );
nor g260 ( new_n398_, new_n390_, new_n202_ );
not g261 ( new_n399_, new_n398_ );
nor g262 ( new_n400_, new_n357_, new_n399_ );
nor g263 ( new_n401_, new_n397_, new_n400_ );
nor g264 ( new_n402_, new_n401_, new_n284_ );
not g265 ( new_n403_, new_n256_ );
nor g266 ( new_n404_, new_n255_, new_n204_ );
nor g267 ( new_n405_, new_n403_, new_n404_ );
not g268 ( new_n406_, new_n280_ );
nand g269 ( new_n407_, new_n405_, new_n406_ );
nand g270 ( new_n408_, new_n407_, new_n281_ );
nand g271 ( new_n409_, new_n408_, new_n202_ );
nor g272 ( new_n410_, new_n390_, keyIn_0_26 );
not g273 ( new_n411_, new_n410_ );
nand g274 ( new_n412_, new_n390_, keyIn_0_26 );
nand g275 ( new_n413_, new_n411_, new_n412_ );
nand g276 ( new_n414_, new_n413_, new_n357_ );
nor g277 ( new_n415_, new_n414_, new_n409_ );
nand g278 ( new_n416_, new_n415_, keyIn_0_36 );
not g279 ( new_n417_, keyIn_0_36 );
nor g280 ( new_n418_, new_n284_, new_n203_ );
nor g281 ( new_n419_, new_n354_, new_n355_ );
nor g282 ( new_n420_, new_n327_, new_n350_ );
nor g283 ( new_n421_, new_n419_, new_n420_ );
not g284 ( new_n422_, new_n412_ );
nor g285 ( new_n423_, new_n422_, new_n410_ );
nor g286 ( new_n424_, new_n421_, new_n423_ );
nand g287 ( new_n425_, new_n418_, new_n424_ );
nand g288 ( new_n426_, new_n425_, new_n417_ );
nand g289 ( new_n427_, new_n426_, new_n416_ );
nor g290 ( new_n428_, new_n421_, new_n399_ );
nand g291 ( new_n429_, new_n428_, new_n284_ );
nand g292 ( new_n430_, new_n427_, new_n429_ );
nor g293 ( new_n431_, new_n430_, new_n402_ );
not g294 ( new_n432_, keyIn_0_21 );
not g295 ( new_n433_, keyIn_0_17 );
not g296 ( new_n434_, keyIn_0_2 );
not g297 ( new_n435_, N33 );
not g298 ( new_n436_, N37 );
nand g299 ( new_n437_, new_n435_, new_n436_ );
nand g300 ( new_n438_, N33, N37 );
nand g301 ( new_n439_, new_n437_, new_n438_ );
nand g302 ( new_n440_, new_n439_, new_n434_ );
nor g303 ( new_n441_, N33, N37 );
nor g304 ( new_n442_, new_n441_, new_n434_ );
nand g305 ( new_n443_, new_n442_, new_n438_ );
nand g306 ( new_n444_, new_n440_, new_n443_ );
not g307 ( new_n445_, new_n444_ );
not g308 ( new_n446_, keyIn_0_3 );
nor g309 ( new_n447_, N41, N45 );
nand g310 ( new_n448_, N41, N45 );
not g311 ( new_n449_, new_n448_ );
nor g312 ( new_n450_, new_n449_, new_n447_ );
nor g313 ( new_n451_, new_n450_, new_n446_ );
not g314 ( new_n452_, N41 );
nand g315 ( new_n453_, new_n452_, new_n272_ );
nand g316 ( new_n454_, new_n453_, new_n448_ );
nor g317 ( new_n455_, new_n454_, keyIn_0_3 );
nor g318 ( new_n456_, new_n451_, new_n455_ );
nand g319 ( new_n457_, new_n445_, new_n456_ );
nand g320 ( new_n458_, new_n454_, keyIn_0_3 );
nand g321 ( new_n459_, new_n450_, new_n446_ );
nand g322 ( new_n460_, new_n459_, new_n458_ );
nand g323 ( new_n461_, new_n460_, new_n444_ );
nand g324 ( new_n462_, new_n457_, new_n461_ );
nand g325 ( new_n463_, new_n462_, new_n433_ );
nor g326 ( new_n464_, new_n460_, new_n444_ );
not g327 ( new_n465_, new_n461_ );
nor g328 ( new_n466_, new_n465_, new_n464_ );
nand g329 ( new_n467_, new_n466_, keyIn_0_17 );
nand g330 ( new_n468_, new_n467_, new_n463_ );
nand g331 ( new_n469_, N1, N5 );
not g332 ( new_n470_, new_n469_ );
nor g333 ( new_n471_, N1, N5 );
nor g334 ( new_n472_, new_n470_, new_n471_ );
not g335 ( new_n473_, new_n472_ );
nand g336 ( new_n474_, N9, N13 );
not g337 ( new_n475_, new_n474_ );
nor g338 ( new_n476_, N9, N13 );
nor g339 ( new_n477_, new_n475_, new_n476_ );
not g340 ( new_n478_, new_n477_ );
nor g341 ( new_n479_, new_n473_, new_n478_ );
nor g342 ( new_n480_, new_n472_, new_n477_ );
nor g343 ( new_n481_, new_n479_, new_n480_ );
not g344 ( new_n482_, new_n481_ );
nand g345 ( new_n483_, new_n482_, keyIn_0_16 );
not g346 ( new_n484_, keyIn_0_16 );
nand g347 ( new_n485_, new_n481_, new_n484_ );
nand g348 ( new_n486_, new_n483_, new_n485_ );
nand g349 ( new_n487_, new_n468_, new_n486_ );
nor g350 ( new_n488_, new_n466_, keyIn_0_17 );
nor g351 ( new_n489_, new_n462_, new_n433_ );
nor g352 ( new_n490_, new_n488_, new_n489_ );
not g353 ( new_n491_, new_n486_ );
nand g354 ( new_n492_, new_n490_, new_n491_ );
nand g355 ( new_n493_, new_n492_, new_n487_ );
nand g356 ( new_n494_, new_n493_, new_n432_ );
nor g357 ( new_n495_, new_n490_, new_n491_ );
nor g358 ( new_n496_, new_n468_, new_n486_ );
nor g359 ( new_n497_, new_n495_, new_n496_ );
nand g360 ( new_n498_, new_n497_, keyIn_0_21 );
nand g361 ( new_n499_, new_n498_, new_n494_ );
nand g362 ( new_n500_, new_n499_, keyIn_0_10 );
not g363 ( new_n501_, keyIn_0_10 );
nor g364 ( new_n502_, new_n497_, keyIn_0_21 );
nor g365 ( new_n503_, new_n493_, new_n432_ );
nor g366 ( new_n504_, new_n502_, new_n503_ );
nand g367 ( new_n505_, new_n504_, new_n501_ );
nand g368 ( new_n506_, new_n505_, new_n500_ );
nand g369 ( new_n507_, N135, N137 );
nand g370 ( new_n508_, new_n506_, new_n507_ );
nor g371 ( new_n509_, new_n504_, new_n501_ );
nor g372 ( new_n510_, new_n499_, keyIn_0_10 );
nor g373 ( new_n511_, new_n509_, new_n510_ );
not g374 ( new_n512_, new_n507_ );
nand g375 ( new_n513_, new_n511_, new_n512_ );
nand g376 ( new_n514_, new_n513_, new_n508_ );
not g377 ( new_n515_, keyIn_0_20 );
nand g378 ( new_n516_, N73, N89 );
not g379 ( new_n517_, new_n516_ );
nor g380 ( new_n518_, N73, N89 );
nor g381 ( new_n519_, new_n517_, new_n518_ );
not g382 ( new_n520_, new_n519_ );
nand g383 ( new_n521_, N105, N121 );
not g384 ( new_n522_, new_n521_ );
nor g385 ( new_n523_, N105, N121 );
nor g386 ( new_n524_, new_n522_, new_n523_ );
not g387 ( new_n525_, new_n524_ );
nor g388 ( new_n526_, new_n520_, new_n525_ );
nor g389 ( new_n527_, new_n519_, new_n524_ );
nor g390 ( new_n528_, new_n526_, new_n527_ );
not g391 ( new_n529_, new_n528_ );
nand g392 ( new_n530_, new_n529_, new_n515_ );
not g393 ( new_n531_, new_n530_ );
nor g394 ( new_n532_, new_n529_, new_n515_ );
nor g395 ( new_n533_, new_n531_, new_n532_ );
not g396 ( new_n534_, new_n533_ );
nand g397 ( new_n535_, new_n514_, new_n534_ );
not g398 ( new_n536_, new_n535_ );
nor g399 ( new_n537_, new_n514_, new_n534_ );
nor g400 ( new_n538_, new_n536_, new_n537_ );
nor g401 ( new_n539_, new_n431_, new_n538_ );
not g402 ( new_n540_, new_n539_ );
nor g403 ( new_n541_, new_n540_, new_n203_ );
nor g404 ( new_n542_, N49, N53 );
nand g405 ( new_n543_, N49, N53 );
not g406 ( new_n544_, new_n543_ );
nor g407 ( new_n545_, new_n544_, new_n542_ );
not g408 ( new_n546_, new_n545_ );
not g409 ( new_n547_, N57 );
nor g410 ( new_n548_, new_n547_, N61 );
nor g411 ( new_n549_, new_n274_, N57 );
nor g412 ( new_n550_, new_n548_, new_n549_ );
not g413 ( new_n551_, new_n550_ );
nand g414 ( new_n552_, new_n551_, keyIn_0_4 );
nor g415 ( new_n553_, new_n551_, keyIn_0_4 );
not g416 ( new_n554_, new_n553_ );
nand g417 ( new_n555_, new_n554_, new_n552_ );
nor g418 ( new_n556_, new_n555_, new_n546_ );
not g419 ( new_n557_, new_n556_ );
nand g420 ( new_n558_, new_n555_, new_n546_ );
nand g421 ( new_n559_, new_n557_, new_n558_ );
nor g422 ( new_n560_, new_n490_, new_n559_ );
not g423 ( new_n561_, new_n558_ );
nor g424 ( new_n562_, new_n561_, new_n556_ );
nor g425 ( new_n563_, new_n562_, new_n468_ );
nor g426 ( new_n564_, new_n560_, new_n563_ );
not g427 ( new_n565_, new_n564_ );
nand g428 ( new_n566_, N134, N137 );
nor g429 ( new_n567_, new_n565_, new_n566_ );
not g430 ( new_n568_, new_n567_ );
nand g431 ( new_n569_, new_n565_, new_n566_ );
nand g432 ( new_n570_, new_n568_, new_n569_ );
nand g433 ( new_n571_, N101, N117 );
not g434 ( new_n572_, new_n571_ );
nor g435 ( new_n573_, N101, N117 );
nor g436 ( new_n574_, new_n572_, new_n573_ );
nand g437 ( new_n575_, N69, N85 );
not g438 ( new_n576_, new_n575_ );
nor g439 ( new_n577_, N69, N85 );
nor g440 ( new_n578_, new_n576_, new_n577_ );
not g441 ( new_n579_, new_n578_ );
nor g442 ( new_n580_, new_n579_, new_n574_ );
nand g443 ( new_n581_, new_n579_, new_n574_ );
not g444 ( new_n582_, new_n581_ );
nor g445 ( new_n583_, new_n582_, new_n580_ );
nand g446 ( new_n584_, new_n570_, new_n583_ );
not g447 ( new_n585_, new_n584_ );
nor g448 ( new_n586_, new_n570_, new_n583_ );
nor g449 ( new_n587_, new_n585_, new_n586_ );
nor g450 ( new_n588_, N25, N29 );
nand g451 ( new_n589_, N25, N29 );
not g452 ( new_n590_, new_n589_ );
nor g453 ( new_n591_, new_n590_, new_n588_ );
not g454 ( new_n592_, keyIn_0_1 );
not g455 ( new_n593_, N21 );
nand g456 ( new_n594_, new_n593_, N17 );
not g457 ( new_n595_, N17 );
nand g458 ( new_n596_, new_n595_, N21 );
nand g459 ( new_n597_, new_n594_, new_n596_ );
nand g460 ( new_n598_, new_n597_, keyIn_0_0 );
not g461 ( new_n599_, new_n598_ );
nor g462 ( new_n600_, new_n597_, keyIn_0_0 );
nor g463 ( new_n601_, new_n599_, new_n600_ );
nor g464 ( new_n602_, new_n601_, new_n592_ );
not g465 ( new_n603_, keyIn_0_0 );
not g466 ( new_n604_, new_n597_ );
nand g467 ( new_n605_, new_n604_, new_n603_ );
nand g468 ( new_n606_, new_n605_, new_n598_ );
nor g469 ( new_n607_, new_n606_, keyIn_0_1 );
nor g470 ( new_n608_, new_n602_, new_n607_ );
nand g471 ( new_n609_, new_n608_, new_n591_ );
not g472 ( new_n610_, new_n591_ );
nand g473 ( new_n611_, new_n606_, keyIn_0_1 );
nand g474 ( new_n612_, new_n601_, new_n592_ );
nand g475 ( new_n613_, new_n612_, new_n611_ );
nand g476 ( new_n614_, new_n613_, new_n610_ );
nand g477 ( new_n615_, new_n609_, new_n614_ );
nor g478 ( new_n616_, new_n615_, new_n486_ );
not g479 ( new_n617_, new_n616_ );
nand g480 ( new_n618_, new_n615_, new_n486_ );
nand g481 ( new_n619_, new_n617_, new_n618_ );
nand g482 ( new_n620_, N133, N137 );
nand g483 ( new_n621_, new_n619_, new_n620_ );
not g484 ( new_n622_, new_n618_ );
nor g485 ( new_n623_, new_n622_, new_n616_ );
not g486 ( new_n624_, new_n620_ );
nand g487 ( new_n625_, new_n623_, new_n624_ );
nand g488 ( new_n626_, new_n625_, new_n621_ );
not g489 ( new_n627_, N97 );
nor g490 ( new_n628_, new_n627_, N113 );
nor g491 ( new_n629_, new_n212_, N97 );
nor g492 ( new_n630_, new_n628_, new_n629_ );
not g493 ( new_n631_, new_n630_ );
nand g494 ( new_n632_, new_n631_, keyIn_0_15 );
not g495 ( new_n633_, new_n632_ );
nor g496 ( new_n634_, new_n631_, keyIn_0_15 );
nor g497 ( new_n635_, new_n633_, new_n634_ );
not g498 ( new_n636_, new_n635_ );
not g499 ( new_n637_, N65 );
nor g500 ( new_n638_, new_n637_, N81 );
not g501 ( new_n639_, N81 );
nor g502 ( new_n640_, new_n639_, N65 );
nor g503 ( new_n641_, new_n638_, new_n640_ );
nor g504 ( new_n642_, new_n636_, new_n641_ );
nand g505 ( new_n643_, new_n636_, new_n641_ );
not g506 ( new_n644_, new_n643_ );
nor g507 ( new_n645_, new_n644_, new_n642_ );
not g508 ( new_n646_, new_n645_ );
nor g509 ( new_n647_, new_n626_, new_n646_ );
nand g510 ( new_n648_, new_n626_, new_n646_ );
not g511 ( new_n649_, new_n648_ );
nor g512 ( new_n650_, new_n649_, new_n647_ );
nor g513 ( new_n651_, new_n587_, new_n650_ );
not g514 ( new_n652_, new_n651_ );
not g515 ( new_n653_, keyIn_0_11 );
nand g516 ( new_n654_, new_n615_, new_n562_ );
not g517 ( new_n655_, new_n654_ );
nor g518 ( new_n656_, new_n615_, new_n562_ );
nor g519 ( new_n657_, new_n655_, new_n656_ );
nand g520 ( new_n658_, new_n657_, new_n653_ );
nor g521 ( new_n659_, new_n613_, new_n610_ );
not g522 ( new_n660_, new_n614_ );
nor g523 ( new_n661_, new_n660_, new_n659_ );
nand g524 ( new_n662_, new_n661_, new_n559_ );
nand g525 ( new_n663_, new_n662_, new_n654_ );
nand g526 ( new_n664_, new_n663_, keyIn_0_11 );
nand g527 ( new_n665_, new_n658_, new_n664_ );
nand g528 ( new_n666_, N136, N137 );
nand g529 ( new_n667_, new_n665_, new_n666_ );
not g530 ( new_n668_, new_n667_ );
nor g531 ( new_n669_, new_n665_, new_n666_ );
nor g532 ( new_n670_, new_n668_, new_n669_ );
nand g533 ( new_n671_, N109, N125 );
not g534 ( new_n672_, new_n671_ );
nor g535 ( new_n673_, N109, N125 );
nor g536 ( new_n674_, new_n672_, new_n673_ );
nand g537 ( new_n675_, N77, N93 );
not g538 ( new_n676_, new_n675_ );
nor g539 ( new_n677_, N77, N93 );
nor g540 ( new_n678_, new_n676_, new_n677_ );
not g541 ( new_n679_, new_n678_ );
nor g542 ( new_n680_, new_n679_, new_n674_ );
nand g543 ( new_n681_, new_n679_, new_n674_ );
not g544 ( new_n682_, new_n681_ );
nor g545 ( new_n683_, new_n682_, new_n680_ );
nor g546 ( new_n684_, new_n670_, new_n683_ );
nor g547 ( new_n685_, new_n663_, keyIn_0_11 );
not g548 ( new_n686_, new_n664_ );
nor g549 ( new_n687_, new_n686_, new_n685_ );
not g550 ( new_n688_, new_n666_ );
nand g551 ( new_n689_, new_n687_, new_n688_ );
nand g552 ( new_n690_, new_n689_, new_n667_ );
not g553 ( new_n691_, new_n683_ );
nor g554 ( new_n692_, new_n690_, new_n691_ );
nor g555 ( new_n693_, new_n684_, new_n692_ );
nor g556 ( new_n694_, new_n652_, new_n693_ );
nand g557 ( new_n695_, new_n541_, new_n694_ );
nand g558 ( new_n696_, new_n695_, keyIn_0_41 );
nor g559 ( new_n697_, new_n695_, keyIn_0_41 );
not g560 ( new_n698_, new_n697_ );
nand g561 ( new_n699_, new_n698_, new_n696_ );
nand g562 ( new_n700_, new_n699_, new_n138_ );
not g563 ( new_n701_, new_n699_ );
nand g564 ( new_n702_, new_n701_, N1 );
nand g565 ( N724, new_n702_, new_n700_ );
nor g566 ( new_n704_, new_n540_, new_n357_ );
nand g567 ( new_n705_, new_n704_, new_n694_ );
nand g568 ( new_n706_, new_n705_, keyIn_0_42 );
nor g569 ( new_n707_, new_n705_, keyIn_0_42 );
not g570 ( new_n708_, new_n707_ );
nand g571 ( new_n709_, new_n708_, new_n706_ );
nand g572 ( new_n710_, new_n709_, N5 );
not g573 ( new_n711_, N5 );
not g574 ( new_n712_, new_n709_ );
nand g575 ( new_n713_, new_n712_, new_n711_ );
nand g576 ( N725, new_n713_, new_n710_ );
not g577 ( new_n715_, new_n390_ );
nand g578 ( new_n716_, new_n539_, new_n694_ );
nor g579 ( new_n717_, new_n716_, new_n715_ );
not g580 ( new_n718_, new_n717_ );
nand g581 ( new_n719_, new_n718_, N9 );
not g582 ( new_n720_, N9 );
nand g583 ( new_n721_, new_n717_, new_n720_ );
nand g584 ( N726, new_n719_, new_n721_ );
nor g585 ( new_n723_, new_n716_, new_n408_ );
not g586 ( new_n724_, new_n723_ );
nand g587 ( new_n725_, new_n724_, N13 );
not g588 ( new_n726_, N13 );
nand g589 ( new_n727_, new_n723_, new_n726_ );
nand g590 ( N727, new_n725_, new_n727_ );
nand g591 ( new_n729_, new_n690_, new_n691_ );
nand g592 ( new_n730_, new_n670_, new_n683_ );
nand g593 ( new_n731_, new_n730_, new_n729_ );
nor g594 ( new_n732_, new_n431_, new_n731_ );
nor g595 ( new_n733_, new_n511_, new_n512_ );
nor g596 ( new_n734_, new_n506_, new_n507_ );
nor g597 ( new_n735_, new_n733_, new_n734_ );
nand g598 ( new_n736_, new_n735_, new_n533_ );
nand g599 ( new_n737_, new_n736_, new_n535_ );
nor g600 ( new_n738_, new_n737_, new_n652_ );
not g601 ( new_n739_, new_n738_ );
nor g602 ( new_n740_, new_n739_, new_n203_ );
nand g603 ( new_n741_, new_n732_, new_n740_ );
not g604 ( new_n742_, new_n741_ );
nor g605 ( new_n743_, new_n742_, new_n595_ );
nor g606 ( new_n744_, new_n741_, N17 );
nor g607 ( new_n745_, new_n743_, new_n744_ );
not g608 ( new_n746_, new_n745_ );
nand g609 ( new_n747_, new_n746_, keyIn_0_54 );
not g610 ( new_n748_, keyIn_0_54 );
nand g611 ( new_n749_, new_n745_, new_n748_ );
nand g612 ( N728, new_n747_, new_n749_ );
nor g613 ( new_n751_, new_n739_, new_n357_ );
nand g614 ( new_n752_, new_n732_, new_n751_ );
not g615 ( new_n753_, new_n752_ );
nor g616 ( new_n754_, new_n753_, new_n593_ );
nor g617 ( new_n755_, new_n752_, N21 );
nor g618 ( new_n756_, new_n754_, new_n755_ );
not g619 ( new_n757_, new_n756_ );
nand g620 ( new_n758_, new_n757_, keyIn_0_55 );
not g621 ( new_n759_, keyIn_0_55 );
nand g622 ( new_n760_, new_n756_, new_n759_ );
nand g623 ( N729, new_n758_, new_n760_ );
not g624 ( new_n762_, N25 );
nor g625 ( new_n763_, new_n739_, new_n715_ );
nand g626 ( new_n764_, new_n732_, new_n763_ );
not g627 ( new_n765_, new_n764_ );
nand g628 ( new_n766_, new_n765_, new_n762_ );
nand g629 ( new_n767_, new_n764_, N25 );
nand g630 ( N730, new_n766_, new_n767_ );
not g631 ( new_n769_, keyIn_0_43 );
nor g632 ( new_n770_, new_n739_, new_n408_ );
nand g633 ( new_n771_, new_n732_, new_n770_ );
nor g634 ( new_n772_, new_n771_, new_n769_ );
nand g635 ( new_n773_, new_n771_, new_n769_ );
not g636 ( new_n774_, new_n773_ );
nor g637 ( new_n775_, new_n774_, new_n772_ );
not g638 ( new_n776_, new_n775_ );
nand g639 ( new_n777_, new_n776_, N29 );
not g640 ( new_n778_, N29 );
nand g641 ( new_n779_, new_n775_, new_n778_ );
nand g642 ( N731, new_n777_, new_n779_ );
nand g643 ( new_n781_, new_n587_, new_n650_ );
nor g644 ( new_n782_, new_n693_, new_n781_ );
nand g645 ( new_n783_, new_n541_, new_n782_ );
nand g646 ( new_n784_, new_n783_, N33 );
nor g647 ( new_n785_, new_n783_, N33 );
not g648 ( new_n786_, new_n785_ );
nand g649 ( new_n787_, new_n786_, new_n784_ );
nand g650 ( new_n788_, new_n787_, keyIn_0_56 );
not g651 ( new_n789_, keyIn_0_56 );
not g652 ( new_n790_, new_n787_ );
nand g653 ( new_n791_, new_n790_, new_n789_ );
nand g654 ( N732, new_n791_, new_n788_ );
nand g655 ( new_n793_, new_n704_, new_n782_ );
nand g656 ( new_n794_, new_n793_, new_n436_ );
nor g657 ( new_n795_, new_n793_, new_n436_ );
not g658 ( new_n796_, new_n795_ );
nand g659 ( new_n797_, new_n796_, new_n794_ );
nand g660 ( new_n798_, new_n797_, keyIn_0_57 );
not g661 ( new_n799_, keyIn_0_57 );
not g662 ( new_n800_, new_n797_ );
nand g663 ( new_n801_, new_n800_, new_n799_ );
nand g664 ( N733, new_n801_, new_n798_ );
not g665 ( new_n803_, keyIn_0_44 );
not g666 ( new_n804_, new_n782_ );
nor g667 ( new_n805_, new_n804_, new_n715_ );
nand g668 ( new_n806_, new_n539_, new_n805_ );
nor g669 ( new_n807_, new_n806_, new_n803_ );
nand g670 ( new_n808_, new_n806_, new_n803_ );
not g671 ( new_n809_, new_n808_ );
nor g672 ( new_n810_, new_n809_, new_n807_ );
not g673 ( new_n811_, new_n810_ );
nand g674 ( new_n812_, new_n811_, N41 );
nand g675 ( new_n813_, new_n810_, new_n452_ );
nand g676 ( N734, new_n812_, new_n813_ );
not g677 ( new_n815_, keyIn_0_58 );
nor g678 ( new_n816_, new_n408_, new_n804_ );
nand g679 ( new_n817_, new_n539_, new_n816_ );
nor g680 ( new_n818_, new_n817_, keyIn_0_45 );
nand g681 ( new_n819_, new_n817_, keyIn_0_45 );
not g682 ( new_n820_, new_n819_ );
nor g683 ( new_n821_, new_n820_, new_n818_ );
nor g684 ( new_n822_, new_n821_, N45 );
nand g685 ( new_n823_, new_n821_, N45 );
not g686 ( new_n824_, new_n823_ );
nor g687 ( new_n825_, new_n824_, new_n822_ );
nand g688 ( new_n826_, new_n825_, new_n815_ );
not g689 ( new_n827_, new_n822_ );
nand g690 ( new_n828_, new_n827_, new_n823_ );
nand g691 ( new_n829_, new_n828_, keyIn_0_58 );
nand g692 ( N735, new_n826_, new_n829_ );
not g693 ( new_n831_, N49 );
not g694 ( new_n832_, new_n402_ );
nor g695 ( new_n833_, new_n425_, new_n417_ );
nor g696 ( new_n834_, new_n415_, keyIn_0_36 );
nor g697 ( new_n835_, new_n833_, new_n834_ );
not g698 ( new_n836_, new_n429_ );
nor g699 ( new_n837_, new_n835_, new_n836_ );
nand g700 ( new_n838_, new_n837_, new_n832_ );
nand g701 ( new_n839_, new_n838_, new_n693_ );
nor g702 ( new_n840_, new_n538_, keyIn_0_27 );
nand g703 ( new_n841_, new_n538_, keyIn_0_27 );
not g704 ( new_n842_, new_n841_ );
nor g705 ( new_n843_, new_n842_, new_n781_ );
not g706 ( new_n844_, new_n843_ );
nor g707 ( new_n845_, new_n844_, new_n840_ );
not g708 ( new_n846_, new_n845_ );
nor g709 ( new_n847_, new_n839_, new_n846_ );
nand g710 ( new_n848_, new_n847_, keyIn_0_39 );
not g711 ( new_n849_, keyIn_0_39 );
nand g712 ( new_n850_, new_n732_, new_n845_ );
nand g713 ( new_n851_, new_n850_, new_n849_ );
nand g714 ( new_n852_, new_n848_, new_n851_ );
nand g715 ( new_n853_, new_n852_, new_n202_ );
nand g716 ( new_n854_, new_n853_, new_n831_ );
not g717 ( new_n855_, new_n854_ );
nor g718 ( new_n856_, new_n853_, new_n831_ );
nor g719 ( new_n857_, new_n855_, new_n856_ );
nand g720 ( new_n858_, new_n857_, keyIn_0_59 );
not g721 ( new_n859_, keyIn_0_59 );
not g722 ( new_n860_, new_n853_ );
nand g723 ( new_n861_, new_n860_, N49 );
nand g724 ( new_n862_, new_n861_, new_n854_ );
nand g725 ( new_n863_, new_n862_, new_n859_ );
nand g726 ( N736, new_n858_, new_n863_ );
not g727 ( new_n865_, keyIn_0_46 );
nand g728 ( new_n866_, new_n852_, new_n421_ );
nand g729 ( new_n867_, new_n866_, new_n865_ );
not g730 ( new_n868_, new_n867_ );
nor g731 ( new_n869_, new_n866_, new_n865_ );
nor g732 ( new_n870_, new_n868_, new_n869_ );
nand g733 ( new_n871_, new_n870_, N53 );
not g734 ( new_n872_, N53 );
not g735 ( new_n873_, new_n866_ );
nand g736 ( new_n874_, new_n873_, keyIn_0_46 );
nand g737 ( new_n875_, new_n874_, new_n867_ );
nand g738 ( new_n876_, new_n875_, new_n872_ );
nand g739 ( N737, new_n871_, new_n876_ );
nor g740 ( new_n878_, new_n850_, new_n849_ );
not g741 ( new_n879_, new_n851_ );
nor g742 ( new_n880_, new_n879_, new_n878_ );
nor g743 ( new_n881_, new_n880_, new_n715_ );
nand g744 ( new_n882_, new_n881_, new_n547_ );
not g745 ( new_n883_, new_n881_ );
nand g746 ( new_n884_, new_n883_, N57 );
nand g747 ( N738, new_n884_, new_n882_ );
nor g748 ( new_n886_, new_n880_, new_n408_ );
nand g749 ( new_n887_, new_n886_, new_n274_ );
not g750 ( new_n888_, new_n886_ );
nand g751 ( new_n889_, new_n888_, N61 );
nand g752 ( N739, new_n889_, new_n887_ );
not g753 ( new_n891_, keyIn_0_47 );
not g754 ( new_n892_, new_n647_ );
nand g755 ( new_n893_, new_n892_, new_n648_ );
not g756 ( new_n894_, keyIn_0_37 );
nor g757 ( new_n895_, new_n737_, keyIn_0_31 );
nand g758 ( new_n896_, new_n737_, keyIn_0_31 );
nand g759 ( new_n897_, new_n896_, new_n782_ );
nor g760 ( new_n898_, new_n897_, new_n895_ );
nand g761 ( new_n899_, new_n898_, new_n894_ );
nor g762 ( new_n900_, new_n898_, new_n894_ );
nand g763 ( new_n901_, new_n538_, keyIn_0_32 );
not g764 ( new_n902_, keyIn_0_32 );
nand g765 ( new_n903_, new_n737_, new_n902_ );
nand g766 ( new_n904_, new_n901_, new_n903_ );
nor g767 ( new_n905_, new_n731_, keyIn_0_33 );
nand g768 ( new_n906_, new_n731_, keyIn_0_33 );
nand g769 ( new_n907_, new_n906_, new_n651_ );
nor g770 ( new_n908_, new_n907_, new_n905_ );
nand g771 ( new_n909_, new_n904_, new_n908_ );
nor g772 ( new_n910_, new_n731_, keyIn_0_30 );
not g773 ( new_n911_, keyIn_0_30 );
nor g774 ( new_n912_, new_n693_, new_n911_ );
nor g775 ( new_n913_, new_n912_, new_n910_ );
nor g776 ( new_n914_, new_n650_, keyIn_0_29 );
not g777 ( new_n915_, keyIn_0_29 );
nor g778 ( new_n916_, new_n893_, new_n915_ );
nor g779 ( new_n917_, new_n914_, new_n916_ );
nor g780 ( new_n918_, new_n917_, new_n587_ );
nand g781 ( new_n919_, new_n737_, new_n918_ );
nor g782 ( new_n920_, new_n919_, new_n913_ );
nand g783 ( new_n921_, new_n587_, keyIn_0_28 );
not g784 ( new_n922_, keyIn_0_28 );
not g785 ( new_n923_, new_n586_ );
nand g786 ( new_n924_, new_n923_, new_n584_ );
nand g787 ( new_n925_, new_n924_, new_n922_ );
nand g788 ( new_n926_, new_n921_, new_n925_ );
nor g789 ( new_n927_, new_n731_, new_n893_ );
nand g790 ( new_n928_, new_n926_, new_n927_ );
nor g791 ( new_n929_, new_n928_, new_n737_ );
nor g792 ( new_n930_, new_n920_, new_n929_ );
nand g793 ( new_n931_, new_n909_, new_n930_ );
nor g794 ( new_n932_, new_n931_, new_n900_ );
nand g795 ( new_n933_, new_n932_, new_n899_ );
nand g796 ( new_n934_, new_n933_, keyIn_0_38 );
not g797 ( new_n935_, new_n934_ );
nor g798 ( new_n936_, new_n933_, keyIn_0_38 );
nor g799 ( new_n937_, new_n935_, new_n936_ );
nor g800 ( new_n938_, new_n409_, new_n391_ );
nand g801 ( new_n939_, new_n937_, new_n938_ );
nand g802 ( new_n940_, new_n939_, keyIn_0_40 );
not g803 ( new_n941_, keyIn_0_40 );
not g804 ( new_n942_, keyIn_0_38 );
not g805 ( new_n943_, new_n933_ );
nand g806 ( new_n944_, new_n943_, new_n942_ );
nand g807 ( new_n945_, new_n944_, new_n934_ );
not g808 ( new_n946_, new_n938_ );
nor g809 ( new_n947_, new_n945_, new_n946_ );
nand g810 ( new_n948_, new_n947_, new_n941_ );
nand g811 ( new_n949_, new_n940_, new_n948_ );
nand g812 ( new_n950_, new_n949_, new_n893_ );
nand g813 ( new_n951_, new_n950_, new_n891_ );
not g814 ( new_n952_, new_n951_ );
nor g815 ( new_n953_, new_n950_, new_n891_ );
nor g816 ( new_n954_, new_n952_, new_n953_ );
nand g817 ( new_n955_, new_n954_, new_n637_ );
not g818 ( new_n956_, new_n950_ );
nand g819 ( new_n957_, new_n956_, keyIn_0_47 );
nand g820 ( new_n958_, new_n957_, new_n951_ );
nand g821 ( new_n959_, new_n958_, N65 );
nand g822 ( N740, new_n955_, new_n959_ );
not g823 ( new_n961_, N69 );
not g824 ( new_n962_, keyIn_0_48 );
nand g825 ( new_n963_, new_n949_, new_n587_ );
nand g826 ( new_n964_, new_n963_, new_n962_ );
not g827 ( new_n965_, new_n964_ );
nor g828 ( new_n966_, new_n963_, new_n962_ );
nor g829 ( new_n967_, new_n965_, new_n966_ );
nand g830 ( new_n968_, new_n967_, new_n961_ );
not g831 ( new_n969_, new_n963_ );
nand g832 ( new_n970_, new_n969_, keyIn_0_48 );
nand g833 ( new_n971_, new_n970_, new_n964_ );
nand g834 ( new_n972_, new_n971_, N69 );
nand g835 ( N741, new_n968_, new_n972_ );
nand g836 ( new_n974_, new_n949_, new_n737_ );
nand g837 ( new_n975_, new_n974_, N73 );
not g838 ( new_n976_, N73 );
not g839 ( new_n977_, new_n974_ );
nand g840 ( new_n978_, new_n977_, new_n976_ );
nand g841 ( N742, new_n978_, new_n975_ );
not g842 ( new_n980_, N77 );
nand g843 ( new_n981_, new_n949_, new_n693_ );
nand g844 ( new_n982_, new_n981_, new_n980_ );
not g845 ( new_n983_, new_n982_ );
nor g846 ( new_n984_, new_n981_, new_n980_ );
nor g847 ( new_n985_, new_n983_, new_n984_ );
nand g848 ( new_n986_, new_n985_, keyIn_0_60 );
not g849 ( new_n987_, keyIn_0_60 );
not g850 ( new_n988_, new_n981_ );
nand g851 ( new_n989_, new_n988_, N77 );
nand g852 ( new_n990_, new_n989_, new_n982_ );
nand g853 ( new_n991_, new_n990_, new_n987_ );
nand g854 ( N743, new_n986_, new_n991_ );
not g855 ( new_n993_, keyIn_0_34 );
nor g856 ( new_n994_, new_n357_, new_n993_ );
nor g857 ( new_n995_, new_n421_, keyIn_0_34 );
nor g858 ( new_n996_, new_n390_, new_n203_ );
nand g859 ( new_n997_, new_n284_, new_n996_ );
nor g860 ( new_n998_, new_n995_, new_n997_ );
not g861 ( new_n999_, new_n998_ );
nor g862 ( new_n1000_, new_n999_, new_n994_ );
not g863 ( new_n1001_, new_n1000_ );
nor g864 ( new_n1002_, new_n945_, new_n1001_ );
not g865 ( new_n1003_, new_n1002_ );
nor g866 ( new_n1004_, new_n1003_, new_n650_ );
not g867 ( new_n1005_, new_n1004_ );
nand g868 ( new_n1006_, new_n1005_, N81 );
nand g869 ( new_n1007_, new_n1004_, new_n639_ );
nand g870 ( N744, new_n1006_, new_n1007_ );
not g871 ( new_n1009_, N85 );
nor g872 ( new_n1010_, new_n1003_, new_n924_ );
nor g873 ( new_n1011_, new_n1010_, keyIn_0_49 );
nand g874 ( new_n1012_, new_n1010_, keyIn_0_49 );
not g875 ( new_n1013_, new_n1012_ );
nor g876 ( new_n1014_, new_n1013_, new_n1011_ );
not g877 ( new_n1015_, new_n1014_ );
nand g878 ( new_n1016_, new_n1015_, new_n1009_ );
nand g879 ( new_n1017_, new_n1014_, N85 );
nand g880 ( N745, new_n1016_, new_n1017_ );
not g881 ( new_n1019_, keyIn_0_61 );
nand g882 ( new_n1020_, new_n937_, new_n737_ );
nor g883 ( new_n1021_, new_n1020_, new_n1001_ );
nor g884 ( new_n1022_, new_n1021_, N89 );
nand g885 ( new_n1023_, new_n1021_, N89 );
not g886 ( new_n1024_, new_n1023_ );
nor g887 ( new_n1025_, new_n1024_, new_n1022_ );
not g888 ( new_n1026_, new_n1025_ );
nand g889 ( new_n1027_, new_n1026_, new_n1019_ );
nand g890 ( new_n1028_, new_n1025_, keyIn_0_61 );
nand g891 ( N746, new_n1027_, new_n1028_ );
nor g892 ( new_n1030_, new_n1003_, new_n731_ );
not g893 ( new_n1031_, new_n1030_ );
nand g894 ( new_n1032_, new_n1031_, N93 );
not g895 ( new_n1033_, N93 );
nand g896 ( new_n1034_, new_n1030_, new_n1033_ );
nand g897 ( N747, new_n1032_, new_n1034_ );
not g898 ( new_n1036_, keyIn_0_35 );
nor g899 ( new_n1037_, new_n203_, new_n1036_ );
nor g900 ( new_n1038_, new_n202_, keyIn_0_35 );
nor g901 ( new_n1039_, new_n1037_, new_n1038_ );
nor g902 ( new_n1040_, new_n1039_, new_n715_ );
nand g903 ( new_n1041_, new_n421_, new_n1040_ );
nor g904 ( new_n1042_, new_n1041_, new_n284_ );
nand g905 ( new_n1043_, new_n937_, new_n1042_ );
nor g906 ( new_n1044_, new_n1043_, new_n650_ );
not g907 ( new_n1045_, new_n1044_ );
nand g908 ( new_n1046_, new_n1045_, N97 );
nand g909 ( new_n1047_, new_n1044_, new_n627_ );
nand g910 ( N748, new_n1046_, new_n1047_ );
not g911 ( new_n1049_, keyIn_0_50 );
nor g912 ( new_n1050_, new_n1043_, new_n924_ );
nor g913 ( new_n1051_, new_n1050_, new_n1049_ );
nand g914 ( new_n1052_, new_n1050_, new_n1049_ );
not g915 ( new_n1053_, new_n1052_ );
nor g916 ( new_n1054_, new_n1053_, new_n1051_ );
not g917 ( new_n1055_, new_n1054_ );
nand g918 ( new_n1056_, new_n1055_, N101 );
not g919 ( new_n1057_, N101 );
nand g920 ( new_n1058_, new_n1054_, new_n1057_ );
nand g921 ( N749, new_n1056_, new_n1058_ );
nor g922 ( new_n1060_, new_n1043_, new_n538_ );
not g923 ( new_n1061_, new_n1060_ );
nand g924 ( new_n1062_, new_n1061_, N105 );
not g925 ( new_n1063_, N105 );
nand g926 ( new_n1064_, new_n1060_, new_n1063_ );
nand g927 ( N750, new_n1062_, new_n1064_ );
nor g928 ( new_n1066_, new_n1043_, new_n731_ );
not g929 ( new_n1067_, new_n1066_ );
nand g930 ( new_n1068_, new_n1067_, N109 );
not g931 ( new_n1069_, N109 );
nand g932 ( new_n1070_, new_n1066_, new_n1069_ );
nand g933 ( N751, new_n1068_, new_n1070_ );
not g934 ( new_n1072_, new_n400_ );
nor g935 ( new_n1073_, new_n1072_, new_n408_ );
not g936 ( new_n1074_, new_n1073_ );
nor g937 ( new_n1075_, new_n1074_, new_n650_ );
nand g938 ( new_n1076_, new_n937_, new_n1075_ );
not g939 ( new_n1077_, new_n1076_ );
nand g940 ( new_n1078_, new_n1077_, new_n212_ );
nand g941 ( new_n1079_, new_n1076_, N113 );
nand g942 ( N752, new_n1078_, new_n1079_ );
nor g943 ( new_n1081_, new_n1074_, new_n924_ );
nand g944 ( new_n1082_, new_n937_, new_n1081_ );
not g945 ( new_n1083_, new_n1082_ );
nor g946 ( new_n1084_, new_n1083_, keyIn_0_51 );
nand g947 ( new_n1085_, new_n1083_, keyIn_0_51 );
not g948 ( new_n1086_, new_n1085_ );
nor g949 ( new_n1087_, new_n1086_, new_n1084_ );
not g950 ( new_n1088_, new_n1087_ );
nand g951 ( new_n1089_, new_n1088_, N117 );
nand g952 ( new_n1090_, new_n1087_, new_n215_ );
nand g953 ( N753, new_n1089_, new_n1090_ );
not g954 ( new_n1092_, keyIn_0_62 );
not g955 ( new_n1093_, N121 );
not g956 ( new_n1094_, keyIn_0_52 );
nor g957 ( new_n1095_, new_n1020_, new_n1074_ );
nor g958 ( new_n1096_, new_n1095_, new_n1094_ );
nor g959 ( new_n1097_, new_n945_, new_n538_ );
nand g960 ( new_n1098_, new_n1097_, new_n1073_ );
nor g961 ( new_n1099_, new_n1098_, keyIn_0_52 );
nor g962 ( new_n1100_, new_n1096_, new_n1099_ );
nor g963 ( new_n1101_, new_n1100_, new_n1093_ );
nand g964 ( new_n1102_, new_n1098_, keyIn_0_52 );
nand g965 ( new_n1103_, new_n1095_, new_n1094_ );
nand g966 ( new_n1104_, new_n1103_, new_n1102_ );
nor g967 ( new_n1105_, new_n1104_, N121 );
nor g968 ( new_n1106_, new_n1101_, new_n1105_ );
nand g969 ( new_n1107_, new_n1106_, new_n1092_ );
nand g970 ( new_n1108_, new_n1104_, N121 );
nand g971 ( new_n1109_, new_n1100_, new_n1093_ );
nand g972 ( new_n1110_, new_n1109_, new_n1108_ );
nand g973 ( new_n1111_, new_n1110_, keyIn_0_62 );
nand g974 ( N754, new_n1107_, new_n1111_ );
not g975 ( new_n1113_, keyIn_0_63 );
not g976 ( new_n1114_, keyIn_0_53 );
nor g977 ( new_n1115_, new_n1074_, new_n731_ );
nand g978 ( new_n1116_, new_n937_, new_n1115_ );
nand g979 ( new_n1117_, new_n1116_, new_n1114_ );
nor g980 ( new_n1118_, new_n1116_, new_n1114_ );
not g981 ( new_n1119_, new_n1118_ );
nand g982 ( new_n1120_, new_n1119_, new_n1117_ );
nor g983 ( new_n1121_, new_n1120_, N125 );
nand g984 ( new_n1122_, new_n1120_, N125 );
not g985 ( new_n1123_, new_n1122_ );
nor g986 ( new_n1124_, new_n1123_, new_n1121_ );
nand g987 ( new_n1125_, new_n1124_, new_n1113_ );
not g988 ( new_n1126_, new_n1121_ );
nand g989 ( new_n1127_, new_n1126_, new_n1122_ );
nand g990 ( new_n1128_, new_n1127_, keyIn_0_63 );
nand g991 ( N755, new_n1125_, new_n1128_ );
endmodule