module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g18881, g23612, g23652, g73, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29219, g29220, g29221, g30327, g30331,
         g30332, g31656, g31665, g34435, g34839, g36, g44, g53, g54, g56, g57,
         g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6753,
         g84, g90, g91, g92, g99, test_so10, test_so26, test_so35, test_so39,
         test_so42, test_so44, test_so46, test_so80, test_so86, test_so92,
         test_so100, g34783, n4895, n4837, n4920, n2787, n5045, g559, n4959,
         g33046, g5057, n5615, g34441, g2771, n5544, g33982, g1882, g34007,
         g2299, g24276, g4040, n5530, g30381, g2547, n5782, g30405, g3243,
         g25604, g452, g30416, g3542, g30466, g5232, g25736, g5813, g34617,
         g33974, g1744, g30505, g5909, g33554, g1802, n5536, g30432, g3554,
         g33064, g6219, n5385, g34881, g807, n5479, g6031, g24216, g847, n5709,
         g24232, n9367, g34733, g4172, g34882, g4372, g33026, g3512, g31867,
         n5471, g25668, g3490, n5454, g24344, n5432, g4235, g33966, g1600,
         g33550, g1714, n5460, g30393, g3155, n5366, g29248, g2236, g4571,
         g4555, g24274, g3698, g33973, g1736, g30360, g1968, n5664, g34460,
         g30494, g5607, g30384, g2657, n5316, g24340, n5439, g29223, g490,
         n5708, g26881, g311, n5317, g34252, g772, n5334, g30489, g5587,
         g29301, g6177, n5874, g6377, g33022, g3167, n5652, g30496, g5615,
         g33043, g4567, g29263, g30533, g6287, g24256, n5302, g34015, g2563,
         g34031, g4776, n5707, g34452, g4593, n5303, g34646, g6199, g34001,
         g2295, g25633, g1384, g24259, g1339, g33049, g5180, n5384, g34609,
         g2844, g31869, g1024, g30490, g30427, g3598, g21894, g4264, n5823,
         g33965, g767, n5333, g34645, g5853, g33571, g2089, g34267, g4933,
         g26971, g4521, n5752, g34644, g5507, g30534, g6291, g33535, g294,
         n5680, g30498, g25728, g25743, g25684, g3813, g25613, g562, g34438,
         g608, n5475, g24244, g1205, n5547, g30439, g3909, g30541, g6259,
         g30519, g5905, g25621, g921, g34807, g2955, g25599, g203, g24235,
         g34036, g4878, n5283, g30476, g5204, g30429, g3606, g32997, g1926,
         n5510, g33063, g6215, n5651, g30424, g3586, g32977, g291, n5679,
         g34026, g4674, n5440, g30420, g3570, g33560, g29226, g676, n5751,
         g25619, g843, g34455, g4332, n5540, g30457, g4153, g33625, g6336,
         n5592, g34790, g622, n5672, g30414, g3506, n5576, g26966, g4558,
         g25656, g3111, g30390, g25688, g34727, g939, g25594, g278, n5627,
         g26963, g4492, g34034, g4864, n5318, g33541, g1036, g28093, g24236,
         g1178, g30404, g3239, g28051, g718, g29303, g6195, n5741, g26917,
         g1135, n5328, g33624, g6395, n5396, g24337, g34911, g554, g33963,
         g496, g34627, g3853, g29282, g5134, n5807, g25676, g33013, g2485,
         n5509, g32981, g925, n5725, g34976, n9357, g30483, g5555, g32994,
         g1798, g28070, g34806, g2941, g30453, g3905, g33539, g763, n5332,
         g30526, g6255, g26951, g4375, g34035, g4871, n5443, g34636, g4722,
         g32978, g590, n5472, g30348, g1632, n5836, g24336, n5438, g3100,
         g24250, g29236, g1437, g29298, g6154, n5747, g1579, g30499, g5567,
         g33976, g1752, g32996, g1917, g30335, g744, n5470, g34637, g4737,
         n5867, g25694, g30528, g6267, g24251, g1442, g30521, g26960, g4477,
         n5849, g24239, g34259, g4643, n5382, g30474, g5264, n5703, g33016,
         g2610, g34643, g5160, g30510, g5933, g29239, g1454, g26897, g753,
         g34729, g1296, g34625, g3151, g34800, g24353, g6727, n5531, g33029,
         g3530, n5569, g4104, g24253, g1532, g24281, g33997, n9352, g34971,
         n9351, g34263, g4754, g24237, g1189, n5642, g33584, g2287, n5353,
         g24280, g4273, n5764, g26920, g1389, g33548, g29296, g5835, n5663,
         g30338, g1171, n5363, g21895, g4269, n5763, g33588, g2399, n5762,
         g34041, g4983, n5367, g30495, g5611, g29279, g4572, g25655, g3143,
         n5882, g34795, g2898, g24269, g3343, g30403, g3235, g33042, g30419,
         g3566, g34023, n9348, g28090, g4961, g34642, g4927, n5879, g30370,
         g2259, n5419, g34448, g2819, n5609, g26946, g5802, g34610, g2852,
         g24209, g417, n5358, g28047, g681, g24206, g437, g26891, g30504,
         g5901, g34798, g2886, g25669, g3494, n5889, g30480, g5511, n5575,
         g33027, g3518, n5645, g33972, g1604, g25697, g5092, g28099, g4831,
         g26947, g4382, g24350, g6386, g24210, g479, g30455, g3965, g28084,
         g33993, g2008, g736, g30444, g3933, g33537, g222, g25650, g3050,
         g25625, g1052, g30366, g2122, n5784, g33593, g2465, n5523, g30502,
         g5889, g33036, g4495, g25595, g34462, g33024, g3179, n5390, g33552,
         g1728, n5352, g34014, g2433, g29273, g3835, n5662, g25748, g6187,
         n5453, g34638, g4917, g30341, g1070, g26899, g822, n5422, g30336,
         g914, n5560, g5339, g26940, g4164, g25622, g34447, g2807, n5379,
         g33613, g4054, n5395, g25749, g6191, n5888, g25704, g5077, n5455,
         g33053, g5523, n5647, g3680, g30555, g6637, g25601, g174, n5402,
         g33971, g1682, g26892, g355, g1087, g26915, g1105, n5478, g33008,
         g30538, g6307, g3802, g25750, g6159, g30369, g2255, n5414, g34446,
         g2815, n5404, g29230, g911, n5559, g43, g33975, g1748, g30497, g5551,
         g30418, g3558, g25721, g5499, n5885, g34622, g30438, g3901, g34266,
         g4888, g30540, g6251, g32986, g1373, g25648, g33960, g157, n5678,
         g34442, g2783, n5403, g4281, g30421, g3574, g33573, g2112, g34730,
         g1283, g24205, g10122_Tj, g4297, n5698, g32979, g758, n5331, g34025,
         g4639, n5727, g25763, g6537, n5884, g30481, g5543, g30517, g5961,
         g30539, g6243, g34880, n9340, g24242, n5654, g30436, g29265, g3476,
         n5786, g32990, g1664, g24245, g1246, n5756, g30553, g6629, g26907,
         g246, n6008, g24278, g4049, g26955, g24282, g2932, g29276, g4575,
         g31894, g4098, n5350, g33037, g4498, g26894, g528, n5327, g34977,
         n5477, g25654, g3139, n5447, g33962, g34451, g4584, n5539, g34250,
         g142, n5724, g29295, g5831, g26905, g239, g25629, g1216, n5442,
         g34792, g2848, g25703, g5022, g32983, g1030, g30402, g3231, g25757,
         g1430, n9336, g33999, g2241, g24262, g1564, g25729, g6148, g30558,
         g6649, g34781, g110, g26901, g225, n5597, g26961, g33039, g4504,
         g33059, g5873, n5388, g31899, g5037, n5611, g33007, g2319, n5375,
         g25720, g5495, n5446, g21891, g30462, g5208, g30487, g5579, g33058,
         g5869, n5649, g24261, g1589, n5755, g25730, g5752, g30531, g6279,
         g30506, g34804, g2975, n5750, g25747, g6167, n5430, n5701, g33601,
         g2599, n5524, g26922, g1448, n5343, g29250, g2370, g30459, g5164,
         n5570, g1333, n5616, g33534, g153, n5677, g30543, g6549, n5571,
         g29275, g4087, n5480, g34030, g34980, g2984, g30451, g3961, g25627,
         g962, n5630, g34657, g101, g30552, g6625, g34979, n9332, g30337,
         g1018, g24254, g24277, g4045, g29237, g1467, g30378, g2461, n5840,
         g33019, n5300, g33623, g5990, n5589, g29235, g1256, n5558, g31902,
         g5029, n5601, g29306, g6519, n5806, g25689, g4169, n5729, g33978,
         g1816, g26970, g4369, g29278, g4578, g34253, g4459, n5765, g29272,
         g3831, n5872, g33595, g2514, g33610, g3288, n5400, g33589, g34605,
         g2145, n5307, g30350, g1700, n5417, g25611, g513, n5548, g2841, n5963,
         g33619, g5297, n5588, g34022, g2763, g34033, g4793, n5368, g34726,
         g952, g31870, g1263, n5674, g33985, g1950, g29283, g5138, n5871,
         g34003, g2307, g25677, g34463, g4664, g33006, g2223, g29292, g5808,
         n5749, g30557, g6645, g33989, g2016, g33033, g3873, n5387, n5699,
         g34005, g2315, g26932, g2811, g30516, g5957, g33575, g2047, g33032,
         g30486, g5575, g34974, n9327, g25678, g3752, g30440, g3917,
         DFF_480_n1, g1585, n5757, g26949, g4388, g30530, g6275, g30542, g6311,
         g25624, g1041, g30383, g33597, g2537, g34598, g26957, g4430, g26967,
         n9325, g28102, g4826, g30524, g6239, g26903, g232, g30475, g5268,
         g34647, g6545, g30377, n9324, g33553, g1772, n5504, g31903, g5052,
         n5607, g25715, g33984, g1890, g33602, g2629, n5521, g28045, g572,
         n5337, g34603, g2130, g33035, g4108, n5715, g4308, g24208, g475, g990,
         n5622, g31, n5469, g34970, n9322, g24213, g33614, g3990, n5594,
         g33060, g30362, g1992, g33023, g3171, n5603, g26898, g812, n5733,
         g25618, g832, g30518, g5897, g4570, n5702, g26959, g4455, g34801,
         g2902, g26884, g333, g25600, g168, g26933, g28066, g3684, g33612,
         g3639, n5591, g24268, g3338, n5527, g25716, g5406, g26906, g269,
         g24203, g401, g24346, g6040, g24207, g441, g25701, n5690, g29269,
         g3808, n5745, g9, n5468, g34255, g30450, g3957, g30456, g4093, n5340,
         g32991, g1760, n5602, g24348, n5437, g34249, g160, n5843, g30371,
         g2279, n5778, g29268, g3498, n5740, g29224, g586, n5336, g33017,
         g2619, n5508, g30339, g1183, n5599, g33967, g1608, g33559, g1779,
         g29255, g2652, g30368, g2193, n5839, g30375, g2393, n5421, g28052,
         g661, g28089, g4950, g33055, g5535, n5566, g30392, g2834, g30343,
         g1361, g30523, g6235, g24233, g1146, n5851, g33018, g32976, g150,
         n5676, g30349, g1696, n5628, g33067, g6555, g26900, g33034, g3881,
         n5564, g30551, g6621, g25667, g3470, n5424, g30452, g3897, g34719,
         g518, g538, g33607, g2606, n5311, g26923, g1472, n5290, g24211,
         g33050, g5188, n5567, g24341, g5689, n5529, g24201, g405, g30463,
         g5216, g6494, g34464, g4669, g24243, g996, g24335, g4531, g34611,
         g2860, g34262, g4743, g30546, g6593, g25591, g4411, g30347, g1413,
         g30556, g6641, g6, g33562, g1936, n5534, g55, g25610, g504, n5519,
         g33015, g2587, n5372, g31896, g4480, g34004, n9314, g30428, g30485,
         g5571, g30422, g3578, g25714, g29294, g5827, n5809, g30423, g3582,
         g30529, g6271, g34028, g4688, n5656, g33587, g2380, g30460, g5196,
         g30401, g3227, g33990, n9312, g29309, g6541, n5739, g30411, g3203,
         g33546, g1668, n5598, g28085, g4760, g26904, g262, g33556, g1840,
         n5451, g25722, g5467, g25605, g460, g33062, g6209, g26893, n5704,
         g28050, g655, g34626, g33583, g2204, n5620, g30472, g5256, g34454,
         g4608, n5274, g34850, g794, n5291, g4423, g24272, g3689, n5532, g5685,
         g24214, g703, n5821, g26909, g862, n5682, g30406, g3247, g33569,
         g2040, n5505, g34628, g4146, n5981, g34458, g4633, n5844, g24240,
         n5304, g34634, g4732, g25700, n5689, g29293, g5817, g33009, g2351,
         n5511, g33603, g2648, g24355, g6736, g34268, g4944, g25691, g4072,
         g26890, g29264, g3466, g28072, g4116, g31900, g5041, n5605, g26956,
         g4434, g29271, g3827, n5808, g29304, g6500, n5748, g29261, g3133,
         n5661, g28063, g3333, g979, n5320, g34027, g4681, g33961, g298, n5675,
         g33604, g32995, g1894, n5374, g34624, g2988, g30415, g3538, g33536,
         g301, g26888, n9306, DFF_709_n1, g28055, g827, n5728, g24238, g33600,
         g2555, n5351, g28105, g5011, g34721, g199, g29307, g6523, n5870,
         g30345, g34453, g4601, n5365, g32980, g854, g29238, g1484, n5865,
         g34639, g4922, g25695, g5080, n5893, g33057, g5863, g26969, g4581,
         n5670, g29253, g2518, g34021, g2567, g26895, g568, n5335, g30413,
         g3263, g30549, g6613, g24347, g25758, g6444, g34808, g2965, g30501,
         g5857, n5573, g33969, n9303, g34440, g890, n5305, g30433, g3562,
         g21900, g26921, g1404, g29270, g3817, n9302, g33038, g4501, g31865,
         g26926, g2724, n5301, g28083, g4704, g34797, g22, g2878, g30478,
         g5220, g34724, g617, n5339, g24212, g26883, g316, g32985, g1277,
         g25761, g6513, n5426, g26886, g336, n5824, g34796, g2882, g32982,
         g33561, g1906, n5503, g26880, g305, n5282, g34975, g8, g26931, g2799,
         g34641, g4912, g34629, g4157, n5983, g33598, g2541, n5461, g33576,
         g2153, n5356, g34720, g550, g26902, g255, g29244, g30468, g5240,
         g26924, g1478, n5289, g33031, g3863, g29245, g1959, g29266, g3480,
         n5868, g30559, g6653, g34794, g2864, g28087, g4894, g30435, g3857,
         n5572, g25609, g28057, g1002, g34439, g776, n5330, g28, n5324, g1236,
         g34260, g4646, n5712, g33012, g2476, g32989, g1657, n5525, g34006,
         g2375, g63, g358, g26910, g896, n5431, g28043, g33021, g3161, g29251,
         g2384, n5700, g34456, g4616, n5608, g26968, g4561, g33991, g2024,
         g3451, g26930, g2795, g34599, g613, n5474, g28082, g4527, g33557,
         g1844, g30511, g5937, g33045, g30379, g2523, n5281, g24267, n5436,
         g34020, g2643, g24249, g1489, n5850, g25592, g30382, n9295, g29285,
         g5156, n5734, n5526, n9294, g25662, g21896, g33563, g1955, g33622,
         g33582, g2273, n5458, g28086, g4771, g25744, g6098, g29262, g3147,
         n5738, g24270, g3347, g33581, g2269, g191, g24266, g2712, g34849,
         g626, n5288, g33618, g2729, g5357, n5393, g34038, g34032, g4709,
         n5518, g34803, g2927, g34459, g4340, n5653, g30509, g5929, g34640,
         g4907, g28069, g4035, g21899, g2946, g31868, g918, n5673, g26938,
         g4082, g25756, g30363, g30334, g577, n5294, g33970, g1620, g30391,
         g2831, g25615, g667, g33540, g930, n5731, g30445, g3937, g25617, g817,
         n5822, g24247, g1249, g24215, g837, n5562, g33964, g599, n5550,
         g25719, g5475, n5425, g29228, g30514, g5949, g33627, g6682, n5590,
         g24231, g904, g34615, g2873, n5488, g30356, g1854, n5785, g25696,
         g5084, n5681, g30493, g5603, n5726, g33594, g2495, n5522, g34009,
         g2437, g30365, g2102, n5666, g33004, g2208, g34018, g25685, g4064,
         n5416, g34040, g4899, n5517, g25639, g2719, n5465, g34029, g4785,
         n5361, g30488, g5583, g34600, g781, n5551, g29300, g6173, n5810,
         g34802, g2917, g25614, g686, g28058, g1252, n5554, g29225, g671,
         g33580, g30532, g6283, DFF_909_n1, g33054, g5527, n5389, g26962,
         g4489, g33564, g1974, n5450, g32984, g1270, n5716, g34039, g4966,
         n5706, g33065, g6227, n5568, g30443, g3929, g29291, g5503, n5737,
         g24279, g30508, g5925, g29232, g1124, g34269, g4955, g30464, g5224,
         g33988, g2012, g30522, g6203, n5574, g25708, g5120, g30374, g2389,
         n5631, g26953, g4438, g34008, g2429, g34444, g2787, n5610, g34731,
         g33606, g2675, n5457, g24334, g34265, g4836, n5713, g30340, g1199,
         g24257, n5401, g30482, g5547, g34604, g2138, n5275, g33591, g2338,
         n5310, g30525, g6247, g26929, g2791, g30448, g34602, g1291, n2549,
         g30513, g5945, g30469, g5244, g33608, g2759, g33626, g6741, n5398,
         g34725, g785, n5293, g30342, g1259, n5553, g29267, g3484, n5668,
         g25593, g209, n5595, g30548, g6609, g33052, g5517, g34012, g2449,
         g34017, n9281, DFF_961_n1, g24263, g2715, n5299, g26912, g936, n5557,
         g30364, g2098, n5280, g34254, g4462, n5671, g34251, g604, n5473,
         g30560, g6589, g33983, n9280, g24204, g429, g33980, g1870, g34631,
         g29243, g1825, g25623, g1008, n5321, g26950, g4392, n5710, g30431,
         g3546, g30467, g5236, g30353, g1768, n5834, g34467, g4854, g30442,
         g3925, g29305, g6509, g25616, g732, g29252, g2504, g4519, g4520,
         g33003, g2185, n5376, g34613, g37, g4031, g33570, g2070, n5535,
         g34734, g4176, g24275, n5435, g4405, g872, g29302, g6181, n5667,
         g24349, g34264, g4765, g30484, g5563, g25634, g1395, g33567, g1913,
         g33585, g2331, n5513, g30527, g6263, g34978, n9276, g30447, g3945,
         g347, n5860, g34256, g4473, g25630, g1266, g29290, g5489, n5660,
         g29227, g31872, g2748, n5516, g29287, g5471, g31897, g4540, g6723,
         g30562, g6605, g34011, n9274, g33996, g2173, g21898, g33014, g2491,
         g34465, g4849, g33995, g2169, g30372, n9273, g30545, g30389, g33590,
         g2407, n5459, g34616, g2868, g26927, g2767, g32992, g1783, n5596,
         g25631, g1312, n5466, g30477, g5212, g34632, g4245, g28046, g645,
         g4291, g26896, n5657, g25602, g26916, g1129, n5329, g33578, g2227,
         n5538, g33579, g2246, g30354, g1830, n5413, g30425, g3590, g24200,
         g392, g33544, g1592, n5362, g25764, g6505, g24246, g1221, g30507,
         g5921, g26889, g30333, g218, g32998, g1932, g32987, g1624, n5370,
         g25702, g5062, g29286, g5462, n5744, g34606, g2689, g33070, g6573,
         n5563, g29240, g1677, g32999, g2028, n5371, g33605, g2671, g24255,
         g26945, g33558, g1848, n5464, g25699, n5669, g29289, g5485, n5869,
         g30388, g2741, n5349, n5482, g29254, g2638, g28074, g4122, g34450,
         g4322, n5506, g30512, g5941, g33572, g2108, n5452, g25, g33551,
         g33538, g595, n5476, g33005, g2217, n5512, g24248, n9267, g33002,
         g2066, g24234, g1152, n5618, g30471, g5252, g34000, g2165, g34016,
         g2571, g33048, g5176, n5650, g25628, g26934, g2827, g34468, g4859,
         g24202, g424, g33542, g1274, n5730, n9265, n6006, g34445, g2803,
         n5545, g33555, g1821, g34013, g2509, g28091, g5073, g26919, n5556,
         g30554, g6633, g29281, g5124, g30537, g6303, g28092, g5069, g34732,
         g2994, n5634, g28049, g650, g33545, g1636, n5549, g30441, g3921,
         g29247, g24354, g6732, g25636, g1306, n5796, g26914, g1061, g25670,
         g3462, g33998, g2181, g25626, g956, n5341, g33977, g1756, g29297,
         g5849, n5736, g28071, g4112, g30387, n9262, g33577, g2197, n5514,
         g33592, g26913, g1046, g28044, g482, n5820, g26948, g4401, g30344,
         g1514, n5364, g26885, g329, n5766, g33069, g6565, n5386, g34621,
         g2950, g28059, g1345, g25762, g6533, n5445, g34633, g4727, g24352,
         g26925, g1536, g30446, g3941, g25597, g370, g24342, g5694, g30357,
         g1858, g26908, g446, g30399, g3219, g29242, g1811, g30547, g6601,
         g34010, g2441, g33986, g1874, g34257, g30544, g6581, g30561, g6597,
         g5008, g30430, g3610, g34799, g2890, g33565, g1978, g33968, g1612,
         g34843, g112, g34793, g2856, g33566, g1982, n5462, g30465, g28073,
         g4119, g24351, g6390, g30346, g1542, g21893, g4258, g4818, g31904,
         g5033, g34635, g4717, g25637, g1554, n5768, g29274, g3849, n5735,
         g30396, g3199, g25735, g34037, g4975, n5360, g34791, g790, n5292,
         g30520, g5913, g30358, g1902, n5837, g29299, g6163, g25690, g4125,
         g28096, g4821, n5880, g28088, g4939, g24241, n5392, g30397, g3207,
         g4483, g30409, g29284, g5142, n5658, g30470, g5248, g30367, g2126,
         g24273, g3694, g29288, g5481, n5805, g30359, g1964, n5315, g25698,
         g5097, n5753, g30398, g3215, n9255, n6005, g26952, g4427, g26928,
         g2779, n5694, g26954, g30351, g1720, n5780, g31871, g1367, g5112, g19,
         g26939, g4145, g33994, g2161, g25596, g376, n5633, g33586, g2361,
         n5537, g21901, DFF_1234_n1, g31866, g582, n5552, g33000, g2051,
         g26918, g1193, g30373, g2327, n5841, g28056, g907, n5555, g34601,
         g947, n5286, g30355, g1834, n5665, g30426, g3594, g34805, g2999,
         g34002, g2303, g28053, g29229, g723, n5826, g33620, g5703, n5397,
         g34722, g546, g33599, g2472, n5619, g30515, g5953, g25649, g33979,
         g1740, g30417, g3550, g3845, n5886, g33574, g2116, n5463, g30410,
         g30454, g3913, g34024, g33547, g1687, g30386, g2681, n5777, g33596,
         g2533, n5761, g26887, g324, n5827, g34607, g2697, n5308, g31895,
         g4417, g33068, g6561, n5646, g29233, g1141, g24258, n5655, g30376,
         g33549, g1710, g29308, g6527, n5659, g30408, g3255, g29241, g1691,
         g34620, g2936, g33621, g5644, n5593, g5152, n5883, g24339, g5352,
         g34443, g2775, n5378, g34619, g2922, g29234, g30503, g5893, g30550,
         g6617, g33001, g2060, n5507, g33040, g4512, g30492, g5599, g25664,
         g3401, g26944, g4366, g34614, g29260, g3129, n5861, g33047, g5170,
         g24298, g25733, g5821, n5429, g30536, g6299, g29246, g2079, g34261,
         g4698, g33611, g3703, n5399, g25638, g1559, n5441, g34728, n9247,
         g29222, g411, g25742, g30449, g3953, g34608, g2704, n5377, g24345,
         g6035, n5528, n9245, g25635, g1300, n5483, g25686, g4057, n5711,
         g30461, g5200, g34466, g4843, g31901, g5046, n5578, g29249, g2250,
         g26882, n5456, g33041, g33011, g2453, n5373, g25734, g5841, n5449,
         n5705, g34618, g2912, g33010, g2357, g31864, g164, n5561, g34630,
         g4253, n5484, g31898, g5016, n5369, g25653, g3119, n5423, g25632,
         g1351, n5322, g32988, g33616, g29280, g5115, n5743, g33609, g3352,
         n5604, g30563, g6657, g33044, g4552, g30437, g3893, g30412, g3211,
         g30491, g5595, g30434, g3614, g34612, g29259, g3125, n5781, g25681,
         g3821, n5428, g25687, g4141, n5612, g33617, g30479, g5272, g29256,
         g2735, n5600, g28054, g728, g30535, g6295, g30385, g2661, n5418,
         g30361, g1988, n5783, g25705, g24260, g1548, n5546, g29257, g3106,
         n5742, g34461, g4659, g34258, g4358, n5348, g32993, g1792, n5359,
         g33992, g2084, g30394, g3187, g34449, g4311, n5323, g34019, g2583,
         g18597, n9240, g29231, g1094, g25682, g21897, g4284, g30395, g3191,
         g21892, g4239, g4180, n5380, g28048, g691, n5520, g34723, g534,
         g25598, g385, n5632, g33987, g2004, g30380, g2527, n5420, g5456,
         g26965, n6007, g25706, g30458, g4507, n5846, g24338, g5348, g30400,
         g3223, g34623, g2970, g24343, g5698, g30473, g5260, g24252, g1521,
         g33028, g3522, n5383, g29258, g3115, g30407, g3251, g26958, g34457,
         g33568, g1996, n5355, g25663, g26964, g4515, g34735, g4300, g30352,
         n9236, g33543, g1379, g24271, n5433, g33981, g1878, g30500, g5619,
         g34649, g71, g29277, g25612, n5287, g28060, n2505, n2499, n2396,
         n2668, n3122, g72, n5960, n4689, n5961, n4708, n3593, n3595, n3574,
         n3576, n3517, n3519, n3628, n3630, n3555, n3557, n3646, n3648, n3536,
         n3538, n3611, n3613, n3765, n3505, n3525, n3635, n4888, n2595, n2527,
         n3524, n3005, n3623, n3549, n3799, n3033, n3622, n3587, n3586, n3605,
         n3604, n3568, n3567, n3548, n3512, n3511, n3531, n3530, n3641, n3640,
         n3131, n3111, n4537, n4201, n3745, n3684, n3274, n2982, n2706, n2649,
         n2556, n2509, n2487, n2427, n2423, n4826, n2421, n4172, n4173, n4190,
         n4191, n4388, n3951, n3774, n3842, n3808, n3908, n3984, n3875, n4015,
         n3446, n3914, n3406, n3780, n3481, n3957, n3426, n3848, n3491, n3990,
         n3416, n3814, n3436, n3881, n3502, n4022, n3501, n4027, n3407, n3785,
         n3482, n3962, n3427, n3853, n3437, n3886, n3417, n3819, n3492, n3995,
         n3447, n3919, n3682, n3272, n2980, n2704, n2647, n2554, n2507, n2485,
         n2425, n2419, n3743, n2405, n2760, n2552, n4198, n2404, n3653, n4962,
         n4948, n3195, n3116, n4945, n4525, n4518, n3281, n3277, n3276, n2989,
         n2991, n3687, n3279, n2710, n2707, n3174, n3362, n3676, n2644, n3115,
         n3833, n3023, n3933, n3729, n2601, n3664, n3662, n3673, n3671, n2607,
         n3506, n2790, n4490, n4178, n4514, n4196, n3736, n3741, n2598, n4804,
         n4811, n4814, n4519, n2594, n3084, n2590, n4722, n3125, n3105, n3145,
         n3164, n2422, n5121, n4037, n4034, n4039, n3972, n3969, n3929, n3926,
         n3863, n3860, n4003, n4002, n4032, n4035, n3797, n3792, n3790, n3795,
         n3891, n3893, n3827, n3826, n3896, n4007, n3931, n3793, n3924, n3831,
         n3829, n3927, n3974, n3898, n3970, n4000, n3865, n3861, n3824, n3894,
         n3967, n3858, n4005, n3395, n4956, n5026, n3941, n3733, n4798, n4805,
         n4175, n4193, n3738, n4721, n4523, n4524, n4526, n2573, n2577, n2563,
         n2567, n4938, n4913, n4714, n4516, n4517, n5111, n3730, n4305, n4283,
         n2608, n4447, n4448, n4402, n4403, n4425, n4426, n4436, n4437, n4391,
         n4392, n4379, n4380, n4414, n4415, n4458, n4459, n5016, n5014, n3064,
         n3065, n4535, n5112, n3675, counter_31, counter_30, counter_29,
         counter_28, counter_27, counter_26, counter_25, counter_24,
         counter_23, counter_22, counter_21, counter_20, counter_19,
         counter_18, counter_17, counter_16, counter_15, counter_14,
         counter_13, counter_12, counter_11, counter_10, counter_9, counter_8,
         counter_7, counter_6, counter_5, counter_4, counter_3, counter_2,
         counter_1, counter_0, carry_31, carry_30, carry_29, carry_28,
         carry_27, carry_26, carry_25, carry_24, carry_23, carry_22, carry_21,
         carry_20, carry_19, carry_18, carry_17, carry_16, carry_15, carry_14,
         carry_13, carry_12, carry_11, carry_10, carry_9, carry_8, carry_7,
         carry_6, carry_5, carry_4, carry_3, carry_2, N31, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N23, N24, N25, N26, N2, N3, N4, N16,
         N17, N18, N19, N20, N21, N22, N27, N28, N29, N30, N1, N32, n37, n87,
         n73, n86, n85, n84, n83, n82, n81, n80, n79, n78, n77, n76, n75, n74,
         n58, n59, n60, n61, n62, n63, n64, Trigger_out, n65, n66, n67, n68,
         n69, n70, n71, n72, n43, n45, n50, n51, n94, n106, n128, g33959, n175,
         n180, n181, n184, n187, n189, n191, n195, n196, n201, g33533, n240,
         n297, n301, n310, n342, n357, n410, n412, n417, n418, n473, g34788,
         n495, n507, n508, n509, n510, n514, n524, n525, n645, n657, n666,
         n668, n671, n672, n699, n704, n724, n725, n727, n728, n729, n730,
         n756, n770, n772, n776, n777, n797, n872, n875, n876, n877, n878,
         n915, n917, n927, n928, n952, n967, n1011, n1069, n1166, n1169, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1302, n1324, n1326,
         n1330, n1331, n1338, n1574, n1633, n1635, n1697, n7946, n7948, n7949,
         n7950, n7952, n7957, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7973, n7974, n7975, n7980, n7983, n7984, n7986, n7987, n7988, n7989,
         n7990, n7991, n7994, n7995, n7996, n7997, n7999, n8000, n8002, n8003,
         n8004, n8005, n8006, n8010, n8013, n8014, n8015, n8016, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8027, n8029, n8031, n8032, n8033,
         n8034, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8047, n8048,
         n8051, n8052, n8055, n8084, n8085, n8086, n8087, n8088, n8089, n8134,
         n8135, n8179, n8180, n8184, n8185, n8186, n8187, n8192, n8193, n8194,
         n8195, n8196, n8197, n8208, n8211, n8212, n8213, n8214, n8215, n8216,
         n8218, n8219, n8222, n8223, n8224, n8226, n8243, n8244, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8359, n8360, n8361, n8363, n8364, n8365, n8366,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8403, n8404, n8405, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, g32975, n8476, n8477, n8478, n8479, n8480, n8481,
         g31860, n8483, g31862, n8485, g31863, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9237, n9238, n9239, n9241, n9242,
         n9243, n9244, n9246, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9256, n9257, n9258, n9259, n9260, n9261, n9263, n9264, n9266, n9268,
         n9269, n9270, n9271, n9272, n9275, n9277, n9278, n9279, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9296, n9297, n9298, n9299, n9300, n9301, n9304, n9305, n9307, n9308,
         n9309, n9310, n9311, n9313, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9323, n9326, n9328, n9329, n9330, n9331, n9333, n9334, n9335,
         n9337, n9338, n9339, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9349, n9350, n9353, n9354, n9355, n9356, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         U5353_n1, U5355_n1, U5961_n1, U5962_n1, U5963_n1, U5964_n1, U5965_n1,
         U5966_n1, U5967_n1, U5968_n1, U6100_n1, U6211_n1, U6212_n1, U6213_n1,
         U6214_n1, U6215_n1, U6216_n1, U6217_n1, U6218_n1, U6279_n1, U6280_n1,
         U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1, U6286_n1, U6287_n1,
         U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1, U6338_n1, U6341_n1,
         U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1,
         U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1,
         U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1,
         U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1,
         U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6417_n1,
         U6446_n1, U6465_n1, U6497_n1, U6523_n1, U6542_n1, U6552_n1, U6553_n1,
         U6554_n1, U6555_n1, U6556_n1, U6559_n1, U6560_n1, U6561_n1, U6570_n1,
         U6911_n1, U6912_n1, U6917_n1, U6926_n1, U6927_n1, U6929_n1, U6931_n1,
         U6932_n1, U6933_n1, U6934_n1, U6935_n1, U6936_n1, U6937_n1, U6938_n1,
         U6939_n1, U6940_n1, U6941_n1, U6944_n1, U6950_n1, U6954_n1, U6955_n1,
         U6956_n1, U6957_n1, U7174_n1, U7248_n1, U7249_n1, U7402_n1, U7405_n1,
         U7413_n1, U7416_n1, U7427_n1, U7438_n1, U7449_n1, U7455_n1, U7464_n1,
         U7467_n1, U7482_n1, U7492_n1, U7513_n1, U7516_n1, U7549_n1, U7561_n1,
         U7574_n1, U7577_n1, U7585_n1, U7595_n1, U7614_n1, U7621_n1, U7629_n1,
         U7636_n1, U7639_n1, U7649_n1, U7652_n1, U7668_n1, U7673_n1, U7690_n1,
         U7707_n1, U7712_n1, U7792_n1, U7794_n1, U7895_n1, U7897_n1, U7977_n1,
         U8034_n1, U8036_n1, U8050_n1, U8055_n1, U8060_n1, U8070_n1, U8074_n1,
         U8088_n1, U8112_n1, U8113_n1, U8147_n1, U8165_n1, U8185_n1, U8192_n1,
         U8210_n1, U8223_n1, U8224_n1, U8281_n1, U8307_n1, U8974_n1, U8975_n1,
         U9065_n1, U9070_n1, U9075_n1, U9076_n1, U9080_n1, U9084_n1, U9085_n1,
         U9086_n1, U9090_n1, U9098_n1, U9099_n1, U9101_n1, U9107_n1, U9111_n1,
         U9116_n1, U9120_n1, U9124_n1, U9128_n1, U9132_n1, U9136_n1, U9315_n1,
         U9453_n1, U9825_n1, U9886_n1, U9927_n1, U9953_n1, U9957_n1, U9958_n1,
         U9968_n1, U9972_n1, U9992_n1, U10314_n1, U10318_n1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g34597 = 1'b0;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g29218 = g18881;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g24167 = g73;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20557 = g29213;
  assign g20652 = g29214;
  assign g20901 = g29215;
  assign g21176 = g29216;
  assign g21270 = g29217;
  assign g20654 = g29219;
  assign g21245 = g29220;
  assign g21292 = g29221;
  assign g23002 = g30327;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g31521 = g34435;
  assign g34956 = g34839;
  assign g21698 = g36;
  assign g24185 = g44;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18101 = g6746;
  assign g18097 = g6747;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18100 = g6751;
  assign g18092 = g6753;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g31861 = test_so10;
  assign g25219 = test_so10;
  assign g13881 = test_so26;
  assign g9615 = test_so35;
  assign g8785 = test_so39;
  assign g8291 = test_so42;
  assign g17316 = test_so44;
  assign g8178 = test_so46;
  assign g12470 = test_so80;
  assign g11447 = test_so86;
  assign g9682 = test_so92;
  assign g29210 = test_so100;
  assign g20049 = test_so100;
  assign g24166 = g72;
  assign g28753 = g33959;
  assign g27831 = g33533;
  assign g33894 = g34788;
  assign g26801 = g32975;
  assign g25114 = g31860;
  assign g25259 = g31862;
  assign g25167 = g31863;

  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(n8537), .CLK(n8842), .Q(
        g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(n8583), .CLK(n8888), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(n8582), .CLK(n8887), .Q(
        g1882) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(n8629), .CLK(n8934), .Q(
        g2299) );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(n8633), .CLK(n8938), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(n8594), .CLK(n8899), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(n8595), .CLK(n8900), .Q(g559) );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(n8639), .CLK(n8944), .Q(
        g3243) );
  SDFFX1 DFF_10_Q_reg ( .D(g25604), .SI(g3243), .SE(n8565), .CLK(n8870), .Q(
        g452) );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(n8580), .CLK(n8885), .Q(
        g3542) );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(n8571), .CLK(n8876), .Q(
        g5232) );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(n8628), .CLK(n8933), .Q(
        g5813), .QN(n8364) );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(n8610), .CLK(n8915), .Q(
        test_so1), .QN(n8520) );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(n8628), .CLK(n8933), 
        .Q(g1744) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(n8593), .CLK(n8898), .Q(
        g5909) );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(n8627), .CLK(n8932), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(n8580), .CLK(n8885), .Q(
        g3554) );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(n8608), .CLK(n8913), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(n8579), .CLK(n8884), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(n8579), .CLK(n8884), .Q(
        g6031) );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(n8565), .CLK(n8870), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(n8588), .CLK(n8893), .Q(
        n9367) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(n8570), .CLK(n8875), .Q(
        g4172) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(n8562), .CLK(n8867), .Q(
        g4372) );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(n8562), .CLK(n8867), .Q(
        g3512), .QN(n8308) );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(n8578), .CLK(n8883), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(g25668), .SI(test_si3), .SE(n8562), .CLK(n8867), 
        .Q(g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(n8547), .CLK(n8852), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(n8629), .CLK(n8934), .Q(
        g4235), .QN(n8291) );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(n8631), .CLK(n8936), .Q(
        g1600) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(n8545), .CLK(n8850), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(n8602), .CLK(n8907), .Q(
        g14451), .QN(n8389) );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(n8605), .CLK(n8910), .Q(
        g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(n8559), .CLK(n8864), .Q(
        g2236), .QN(n8305) );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(n8591), .CLK(n8896), .Q(
        g4555) );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(n8544), .CLK(n8849), .Q(
        g3698), .QN(n8425) );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(n8618), .CLK(n8923), .Q(
        g1736) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(n8618), .CLK(n8923), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(n8618), .CLK(n8923), .Q(
        test_so3), .QN(n8510) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(n8540), .CLK(n8845), 
        .Q(g5607) );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(n8540), .CLK(n8845), .Q(
        g2657), .QN(n5316) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(n8548), .CLK(n8853), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(n8623), .CLK(n8928), .Q(
        g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(n8623), .CLK(n8928), .Q(
        g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(n8579), .CLK(n8884), .Q(
        g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(n8544), .CLK(n8849), .Q(
        g5587) );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(n8549), .CLK(n8854), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(n8605), .CLK(n8910), .Q(
        g6377) );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(n8605), .CLK(n8910), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(n8538), .CLK(n8843), .Q(
        g5615) );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(n8628), .CLK(n8933), .Q(
        g4567) );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(n8544), .CLK(n8849), .Q(
        test_so4), .QN(n8508) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(n8592), .CLK(n8897), 
        .Q(g6287) );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(n8560), .CLK(n8865), .Q(
        g7946), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g7946), .SE(n8569), .CLK(n8874), .Q(
        g2563) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(n8616), .CLK(n8921), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(n8616), .CLK(n8921), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(n8616), .CLK(n8921), .Q(
        g6199) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(n8629), .CLK(n8934), .Q(
        g2295) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(n8546), .CLK(n8851), .Q(
        g1384), .QN(n8434) );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(n8589), .CLK(n8894), .Q(
        g1339) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(n8611), .CLK(n8916), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(n8561), .CLK(n8866), .Q(
        g2844) );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(n8553), .CLK(n8858), .Q(
        g1024), .QN(n8465) );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(n8540), .CLK(n8845), .Q(
        test_so5) );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(n8580), .CLK(n8885), 
        .Q(g3598) );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(n8546), .CLK(n8851), .Q(
        g4264), .QN(n5823) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(n8578), .CLK(n8883), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(n8578), .CLK(n8883), .Q(
        g5853) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(n8608), .CLK(n8913), .Q(
        g13865) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(n8584), .CLK(n8889), .Q(
        g2089) );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(n8552), .CLK(n8857), .Q(
        g4933) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(n8541), .CLK(n8846), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(n8542), .CLK(n8847), .Q(
        g5507) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(n8601), .CLK(n8906), .Q(
        g16656), .QN(n8388) );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(n8639), .CLK(n8944), .Q(
        g6291) );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(n8568), .CLK(n8873), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(n8643), .CLK(n8948), .Q(
        test_so6) );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(n8603), .CLK(n8908), 
        .Q(g9617) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(n8556), .CLK(n8861), .Q(
        g9741), .QN(n7983) );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(n8556), .CLK(n8861), .Q(
        g3813), .QN(n8394) );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(n8556), .CLK(n8861), .Q(
        g562) );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(n8595), .CLK(n8900), .Q(
        g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(n8626), .CLK(n8931), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(n8565), .CLK(n8870), .Q(
        g3909) );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(n8593), .CLK(n8898), .Q(
        g6259) );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(n8593), .CLK(n8898), .Q(
        g5905) );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(n8593), .CLK(n8898), .Q(
        g921), .QN(n8041) );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(n8537), .CLK(n8842), .Q(
        g2955), .QN(n8040) );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(n8622), .CLK(n8927), .Q(
        g203) );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(n8634), .CLK(n8939), .Q(
        test_so7), .QN(n8518) );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(n8574), .CLK(n8879), 
        .Q(g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(n8612), .CLK(n8917), .Q(
        g5204) );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(n8599), .CLK(n8904), .Q(
        g17604), .QN(n8370) );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(n8580), .CLK(n8885), .Q(
        g3606) );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(n8607), .CLK(n8912), .Q(
        g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(n8607), .CLK(n8912), .Q(
        g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(n8580), .CLK(n8885), .Q(
        g3586) );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(n8568), .CLK(n8873), .Q(
        g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(n8619), .CLK(n8924), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(n8580), .CLK(n8885), .Q(
        g3570) );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(n8596), .CLK(n8901), .Q(
        g9048), .QN(n7946) );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(n8596), .CLK(n8901), .Q(
        g17607), .QN(n8433) );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(n8635), .CLK(n8940), .Q(
        test_so8), .QN(n8502) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(n8555), .CLK(n8860), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(n8565), .CLK(n8870), .Q(
        g843), .QN(n8029) );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(n8614), .CLK(n8919), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(n8570), .CLK(n8875), .Q(
        g4153) );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(n8570), .CLK(n8875), .Q(
        g17711), .QN(n8340) );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(n8548), .CLK(n8853), .Q(
        g6336), .QN(n5592) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(n8596), .CLK(n8901), .Q(
        g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(n8602), .CLK(n8907), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(n8591), .CLK(n8896), .Q(
        g4558) );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(n8617), .CLK(n8922), .Q(
        g17685), .QN(n8376) );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(n8617), .CLK(n8922), .Q(
        g3111), .QN(n8397) );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(n8558), .CLK(n8863), .Q(
        g29217) );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g29217), .SE(n8558), .CLK(n8863), .Q(
        test_so9) );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(n8567), .CLK(n8872), 
        .Q(g939) );
  SDFFX1 DFF_128_Q_reg ( .D(g25594), .SI(g939), .SE(n8567), .CLK(n8872), .Q(
        g278), .QN(n5627) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(n8636), .CLK(n8941), .Q(
        g4492) );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(n8574), .CLK(n8879), .Q(
        g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(n8553), .CLK(n8858), .Q(
        g1036), .QN(n8464) );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(n8571), .CLK(n8876), .Q(
        g29220) );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g29220), .SE(n8628), .CLK(n8933), .Q(
        g1178) );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(n8609), .CLK(n8914), .Q(
        g3239) );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(n8609), .CLK(n8914), .Q(
        g718), .QN(n8455) );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(n8637), .CLK(n8942), .Q(
        g6195), .QN(n5741) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(n8576), .CLK(n8881), .Q(
        g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(n8605), .CLK(n8910), .Q(
        g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(n8627), .CLK(n8932), .Q(
        test_so10), .QN(n8494) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(n8641), .CLK(n8946), 
        .Q(g554) );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(n8557), .CLK(n8862), .Q(
        g496) );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(n8557), .CLK(n8862), .Q(
        g3853) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(n8557), .CLK(n8862), .Q(
        g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(n8557), .CLK(n8862), .Q(
        g17404), .QN(n8403) );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(n8603), .CLK(n8908), .Q(
        g8344) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(n8594), .CLK(n8899), .Q(
        g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(n8567), .CLK(n8872), .Q(
        g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(n8538), .CLK(n8843), .Q(
        n9357) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(n8538), .CLK(n8843), .Q(
        g5555) );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(n8604), .CLK(n8909), .Q(
        g14096) );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(n8597), .CLK(n8902), .Q(
        g1798) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(n8597), .CLK(n8902), .Q(
        test_so11), .QN(n8491) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(n8564), .CLK(n8869), 
        .Q(g2941), .QN(n8197) );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(n8564), .CLK(n8869), .Q(
        g3905) );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(n8578), .CLK(n8883), .Q(
        g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(n8639), .CLK(n8944), .Q(
        g6255) );
  SDFFX1 DFF_159_Q_reg ( .D(g26951), .SI(g6255), .SE(n8555), .CLK(n8860), .Q(
        g4375), .QN(n7950) );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(n8574), .CLK(n8879), .Q(
        g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(n8615), .CLK(n8920), .Q(
        g4722) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(n8595), .CLK(n8900), .Q(
        g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(n8600), .CLK(n8905), .Q(
        g13099), .QN(n8386) );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(n8583), .CLK(n8888), .Q(
        g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(n8627), .CLK(n8932), .Q(
        g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(n8627), .CLK(n8932), .Q(
        g3100), .QN(n7997) );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(n8586), .CLK(n8891), .Q(
        test_so12), .QN(n8523) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(n8586), .CLK(n8891), 
        .Q(g1437) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(n8548), .CLK(n8853), .Q(
        g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(n8589), .CLK(n8894), .Q(
        g1579), .QN(n8033) );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(n8538), .CLK(n8843), .Q(
        g5567) );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(n8590), .CLK(n8895), .Q(
        g1752) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(n8614), .CLK(n8919), .Q(
        g1917), .QN(n8449) );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(n8578), .CLK(n8883), .Q(
        g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(n8615), .CLK(n8920), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(n8616), .CLK(n8921), .Q(
        g8132) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(n8592), .CLK(n8897), .Q(
        g6267) );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(n8592), .CLK(n8897), .Q(
        g16659), .QN(n8384) );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(n8586), .CLK(n8891), .Q(
        g1442), .QN(n8222) );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(n8573), .CLK(n8878), .Q(
        test_so13) );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(n8619), .CLK(n8924), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(n8619), .CLK(n8924), .Q(
        g10500) );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(n8618), .CLK(n8923), .Q(
        g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(n8571), .CLK(n8876), .Q(
        g5264) );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(n8617), .CLK(n8922), .Q(
        g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(n8618), .CLK(n8923), .Q(
        g2610), .QN(n8442) );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(n8618), .CLK(n8923), .Q(
        g5160) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(n8598), .CLK(n8903), .Q(
        g5933) );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(n8589), .CLK(n8894), .Q(
        g1454) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(n8578), .CLK(n8883), .Q(
        g753), .QN(n8453) );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(n8578), .CLK(n8883), .Q(
        g1296), .QN(n7948) );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(n8578), .CLK(n8883), .Q(
        g3151) );
  SDFFX1 DFF_197_Q_reg ( .D(g34800), .SI(g3151), .SE(n8610), .CLK(n8915), .Q(
        test_so14) );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(n8600), .CLK(n8905), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(n8602), .CLK(n8907), .Q(
        g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(n357), .SI(g3530), .SE(n8597), .CLK(n8902), .Q(
        g4104), .QN(n8363) );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(n8560), .CLK(n8865), .Q(
        g1532), .QN(n8244) );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(n8561), .CLK(n8866), .Q(
        g9251), .QN(n8184) );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(n8557), .CLK(n8862), .Q(
        n9352) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(n8556), .CLK(n8861), .Q(
        n9351) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(n8556), .CLK(n8861), .Q(
        g4754) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(n8629), .CLK(n8934), .Q(
        g1189), .QN(n5642) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(n8629), .CLK(n8934), .Q(
        g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(n8547), .CLK(n8852), .Q(
        g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(n8546), .CLK(n8851), .Q(
        g1389), .QN(n8326) );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(n8631), .CLK(n8936), .Q(
        test_so15), .QN(n8532) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(n8547), .CLK(n8852), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(n8620), .CLK(n8925), .Q(
        g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(n8620), .CLK(n8925), .Q(
        g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(g33588), .SI(g4269), .SE(n8629), .CLK(n8934), .Q(
        g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(n8612), .CLK(n8917), .Q(
        g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(n8538), .CLK(n8843), .Q(
        g5611) );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(n8601), .CLK(n8906), .Q(
        g16627), .QN(n8390) );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(n8563), .CLK(n8868), .Q(
        g4572) );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(n8552), .CLK(n8857), .Q(
        g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(n8552), .CLK(n8857), .Q(
        g2898) );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(n8609), .CLK(n8914), .Q(
        g3343), .QN(n8084) );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(n8609), .CLK(n8914), .Q(
        g3235) );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(n8627), .CLK(n8932), .Q(
        test_so16) );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(n8602), .CLK(n8907), 
        .Q(g3566) );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(n8572), .CLK(n8877), .Q(
        n9348) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(n8539), .CLK(n8844), .Q(
        g4961) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(n8637), .CLK(n8942), .Q(
        g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(n8559), .CLK(n8864), .Q(
        g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(n8558), .CLK(n8863), .Q(
        g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(n8556), .CLK(n8861), .Q(
        g7257) );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(n8556), .CLK(n8861), .Q(
        g5802), .QN(n7995) );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(n8561), .CLK(n8866), .Q(
        g2852) );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(n8621), .CLK(n8926), .Q(
        g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(n8621), .CLK(n8926), .Q(
        g681), .QN(n8349) );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(n8581), .CLK(n8886), .Q(
        g437) );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(n8625), .CLK(n8930), .Q(
        test_so17), .QN(n8513) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(n8593), .CLK(n8898), 
        .Q(g5901) );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(n8553), .CLK(n8858), .Q(
        g2886) );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(n8544), .CLK(n8849), .Q(
        g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(n8544), .CLK(n8849), .Q(
        g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(n8562), .CLK(n8867), .Q(
        g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(n8631), .CLK(n8936), .Q(
        g1604) );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(n8537), .CLK(n8842), .Q(
        g5092) );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(n8573), .CLK(n8878), .Q(
        g4831) );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(n8573), .CLK(n8878), .Q(
        g4382) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(n8637), .CLK(n8942), .Q(
        g6386), .QN(n8085) );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(n8566), .CLK(n8871), .Q(
        g479), .QN(n8031) );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(n8543), .CLK(n8848), .Q(
        g3965) );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(n8548), .CLK(n8853), .Q(
        test_so18) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(n8584), .CLK(n8889), 
        .Q(g2008) );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(n8597), .CLK(n8902), .Q(
        g736) );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(n8604), .CLK(n8909), .Q(
        g3933) );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(n8568), .CLK(n8873), .Q(
        g222) );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(n8598), .CLK(n8903), .Q(
        g3050) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(n8598), .CLK(n8903), .Q(
        g1052), .QN(n8135) );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(n8598), .CLK(n8903), .Q(
        g17580), .QN(n8372) );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(n8614), .CLK(n8919), .Q(
        g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(n8569), .CLK(n8874), .Q(
        g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(n8603), .CLK(n8908), .Q(
        g5889) );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(n8621), .CLK(n8926), .Q(
        g4495) );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(n8621), .CLK(n8926), .Q(
        g8719), .QN(n8361) );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(n8541), .CLK(n8846), .Q(
        test_so19), .QN(n8522) );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(n8606), .CLK(n8911), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(n8627), .CLK(n8932), .Q(
        g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(n8635), .CLK(n8940), .Q(
        g2433) );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(n8543), .CLK(n8848), .Q(
        g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(g25748), .SI(g3835), .SE(n8608), .CLK(n8913), .Q(
        g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(n8608), .CLK(n8913), .Q(
        g4917) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(n8553), .CLK(n8858), .Q(
        g1070), .QN(n8462) );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(n8630), .CLK(n8935), .Q(
        g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(n8640), .CLK(n8945), .Q(
        g17715) );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(n8567), .CLK(n8872), .Q(
        g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(n8627), .CLK(n8932), .Q(
        g5339) );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(n8570), .CLK(n8875), .Q(
        g4164), .QN(n8187) );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(n8588), .CLK(n8893), .Q(
        test_so20), .QN(n8527) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(n8558), .CLK(n8863), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(n8642), .CLK(n8947), .Q(
        g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(n8549), .CLK(n8854), .Q(
        g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(n8549), .CLK(n8854), .Q(
        g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(n8549), .CLK(n8854), .Q(
        g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(n8602), .CLK(n8907), .Q(
        g3680) );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(n8591), .CLK(n8896), .Q(
        g6637) );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(n8622), .CLK(n8927), .Q(
        g174), .QN(n5402) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(n8545), .CLK(n8850), .Q(
        g1682), .QN(n8025) );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(n8625), .CLK(n8930), .Q(
        g355) );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(n8626), .CLK(n8931), .Q(
        g1087), .QN(n8214) );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(n8577), .CLK(n8882), .Q(
        g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(n8634), .CLK(n8939), .Q(
        test_so21), .QN(n8498) );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(n8639), .CLK(n8944), 
        .Q(g6307) );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(n8639), .CLK(n8944), .Q(
        g3802), .QN(n7991) );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(n8639), .CLK(n8944), .Q(
        g6159), .QN(n8366) );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(n8559), .CLK(n8864), .Q(
        g2255), .QN(n5414) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(n8558), .CLK(n8863), .Q(
        g2815), .QN(n5404) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(n8567), .CLK(n8872), .Q(
        g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n8472), .SI(g911), .SE(n8549), .CLK(n8854), .Q(g43) );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(n8549), .CLK(n8854), .Q(
        g16775), .QN(n8337) );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(n8590), .CLK(n8895), .Q(
        g1748) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(n8545), .CLK(n8850), .Q(
        g5551) );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(n8581), .CLK(n8886), .Q(
        g3558) );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(n8642), .CLK(n8947), .Q(
        g5499), .QN(n5885) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(n8564), .CLK(n8869), .Q(
        test_so22), .QN(n8519) );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(n8564), .CLK(n8869), 
        .Q(g3901) );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(n8572), .CLK(n8877), .Q(
        g4888) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(n8592), .CLK(n8897), .Q(
        g6251) );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(n8617), .CLK(n8922), .Q(
        g17649), .QN(n8378) );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(n8546), .CLK(n8851), .Q(
        g1373), .QN(n8328) );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(n8606), .CLK(n8911), .Q(
        g8215) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(n8575), .CLK(n8880), .Q(
        g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(n8582), .CLK(n8887), .Q(
        g2783), .QN(n5403) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(n8594), .CLK(n8899), .Q(
        g4281), .QN(n8212) );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(n8580), .CLK(n8885), .Q(
        g3574) );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(n8641), .CLK(n8946), .Q(
        g2112) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(n8641), .CLK(n8946), .Q(
        g1283) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(n8581), .CLK(n8886), .Q(
        test_so23) );
  SDFFX1 DFF_325_Q_reg ( .D(g10122_Tj), .SI(test_si24), .SE(n8547), .CLK(n8852), .Q(g4297), .QN(n8420) );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(n8547), .CLK(n8852), .Q(
        g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(n8554), .CLK(n8859), .Q(
        g13272), .QN(n8411) );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(n8578), .CLK(n8883), .Q(
        g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(g34025), .SI(g758), .SE(n8628), .CLK(n8933), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(n8560), .CLK(n8865), .Q(
        g6537), .QN(n5884) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(n8560), .CLK(n8865), .Q(
        g5543) );
  SDFFX1 DFF_334_Q_reg ( .D(g7946), .SI(g5543), .SE(n8560), .CLK(n8865), .Q(
        g8475), .QN(n8410) );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(n8573), .CLK(n8878), .Q(
        g5961) );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(n8638), .CLK(n8943), .Q(
        g6243) );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(n8638), .CLK(n8943), .Q(
        n9340), .QN(n14833) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(n8566), .CLK(n8871), .Q(
        g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(n8603), .CLK(n8908), .Q(
        test_so24) );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(n8563), .CLK(n8868), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(n8563), .CLK(n8868), .Q(
        g1664) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(n8566), .CLK(n8871), .Q(
        g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(n8607), .CLK(n8912), .Q(
        g6629) );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(n8581), .CLK(n8886), .Q(
        g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(n8550), .CLK(n8855), .Q(
        g4049), .QN(n8416) );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(n8641), .CLK(n8946), .Q(
        g7260) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(n8561), .CLK(n8866), .Q(
        g2932) );
  SDFFX1 DFF_350_Q_reg ( .D(g29276), .SI(g2932), .SE(n8572), .CLK(n8877), .Q(
        g4575) );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(n8600), .CLK(n8905), .Q(
        g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(n8622), .CLK(n8927), .Q(
        g4498) );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(n8622), .CLK(n8927), .Q(
        g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(n8537), .CLK(n8842), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(g25654), .SI(test_si26), .SE(n8606), .CLK(n8911), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(n8566), .CLK(n8871), .Q(
        g29215) );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g29215), .SE(n8614), .CLK(n8919), .Q(
        g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(n8568), .CLK(n8873), .Q(
        g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(n8626), .CLK(n8931), .Q(
        g17639) );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(n8547), .CLK(n8852), .Q(
        g5831) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(n8604), .CLK(n8909), .Q(
        g239), .QN(n8330) );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(n8631), .CLK(n8936), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(n8539), .CLK(n8844), .Q(
        g2848) );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(n8633), .CLK(n8938), .Q(
        g5022), .QN(n8437) );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(n8633), .CLK(n8938), .Q(
        g16955) );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(n8553), .CLK(n8858), .Q(
        g1030), .QN(n8327) );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(n8602), .CLK(n8907), .Q(
        test_so26) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(n8606), .CLK(n8911), 
        .Q(g3231) );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(n8624), .CLK(n8929), .Q(
        g9817), .QN(n7986) );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(n8624), .CLK(n8929), .Q(
        g1430), .QN(n8215) );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(n8583), .CLK(n8888), .Q(
        n9336) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(n8583), .CLK(n8888), .Q(
        g2241), .QN(n8024) );
  SDFFX1 DFF_375_Q_reg ( .D(g24262), .SI(g2241), .SE(n8624), .CLK(n8929), .Q(
        g1564), .QN(n8399) );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(n8556), .CLK(n8861), .Q(
        g9680), .QN(n7994) );
  SDFFX1 DFF_377_Q_reg ( .D(test_so92), .SI(g9680), .SE(n8556), .CLK(n8861), 
        .Q(g6148), .QN(n7984) );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(n8637), .CLK(n8942), .Q(
        g6649) );
  SDFFX1 DFF_379_Q_reg ( .D(g34781), .SI(g6649), .SE(n8597), .CLK(n8902), .Q(
        g110), .QN(n8470) );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(n8604), .CLK(n8909), .Q(
        g14147) );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(n8577), .CLK(n8882), .Q(
        g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(n8636), .CLK(n8941), .Q(
        test_so27) );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(n8573), .CLK(n8878), 
        .Q(g4504) );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(n8573), .CLK(n8878), .Q(
        g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(n8634), .CLK(n8939), .Q(
        g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(n8634), .CLK(n8939), .Q(
        g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(g25720), .SI(g2319), .SE(n8642), .CLK(n8947), .Q(
        g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(n8570), .CLK(n8875), .Q(
        g11770) );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(n8571), .CLK(n8876), .Q(
        g5208) );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(n8538), .CLK(n8843), .Q(
        g5579) );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(n8602), .CLK(n8907), .Q(
        g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(n8602), .CLK(n8907), .Q(
        g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(n8556), .CLK(n8861), .Q(
        g5752) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(n8597), .CLK(n8902), .Q(
        g6279) );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(n8597), .CLK(n8902), .Q(
        test_so28) );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(n8576), .CLK(n8881), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(n8549), .CLK(n8854), .Q(
        g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(n8549), .CLK(n8854), .Q(
        g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(n8586), .CLK(n8891), .Q(
        g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(n8589), .CLK(n8894), .Q(
        g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(n8604), .CLK(n8909), .Q(
        g14125) );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(n8611), .CLK(n8916), .Q(
        g2370), .QN(n8301) );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(n8611), .CLK(n8916), .Q(
        g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(n8611), .CLK(n8916), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(n8575), .CLK(n8880), .Q(
        g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(n8600), .CLK(n8905), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(n8600), .CLK(n8905), .Q(
        g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(n8616), .CLK(n8921), .Q(
        test_so29), .QN(n8504) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(n8610), .CLK(n8915), 
        .Q(g2984) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(n8543), .CLK(n8848), .Q(
        g3961) );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(n8628), .CLK(n8933), .Q(
        g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(n8548), .CLK(n8853), .Q(
        g101), .QN(n8290) );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(n8548), .CLK(n8853), .Q(
        g8918) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(n8625), .CLK(n8930), .Q(
        g6625) );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(n8553), .CLK(n8858), .Q(
        n9332) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(n8553), .CLK(n8858), .Q(
        g1018), .QN(n8324) );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(n8557), .CLK(n8862), .Q(
        g17320), .QN(n8405) );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(n8550), .CLK(n8855), .Q(
        g4045), .QN(n8089) );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(n8550), .CLK(n8855), .Q(
        g1467) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(n8569), .CLK(n8874), .Q(
        g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(n8613), .CLK(n8918), .Q(
        test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(n8557), .CLK(n8862), 
        .Q(g5990), .QN(n5589) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(n8588), .CLK(n8893), .Q(
        g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(n8633), .CLK(n8938), .Q(
        g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(g29306), .SI(g5029), .SE(n8600), .CLK(n8905), .Q(
        g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(n8600), .CLK(n8905), .Q(
        g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(n8577), .CLK(n8882), .Q(
        g1816), .QN(n7973) );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(n8620), .CLK(n8925), .Q(
        g4369) );
  SDFFX1 DFF_439_Q_reg ( .D(g29278), .SI(g4369), .SE(n8620), .CLK(n8925), .Q(
        g4578), .QN(n8445) );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(n8620), .CLK(n8925), .Q(
        g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(n8543), .CLK(n8848), .Q(
        g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(n8550), .CLK(n8855), .Q(
        g2514), .QN(n8003) );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(n8552), .CLK(n8857), .Q(
        g3288), .QN(n5400) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(n8590), .CLK(n8895), .Q(
        test_so31) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(n8545), .CLK(n8850), 
        .Q(g2145), .QN(n5307) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(n8545), .CLK(n8850), .Q(
        g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(n8622), .CLK(n8927), .Q(
        g513), .QN(n5548) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(n8559), .CLK(n8864), .Q(
        g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(n8551), .CLK(n8856), .Q(
        g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(n8613), .CLK(n8918), .Q(
        g2763), .QN(n7957) );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(n8616), .CLK(n8921), .Q(
        g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(n8628), .CLK(n8933), .Q(
        g952), .QN(n7949) );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(n8588), .CLK(n8893), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(n8638), .CLK(n8943), .Q(
        g1950), .QN(n8023) );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(n8551), .CLK(n8856), .Q(
        g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(n8632), .CLK(n8937), .Q(
        g2307) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(n8632), .CLK(n8937), .Q(
        test_so32) );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(n8541), .CLK(n8846), 
        .Q(g8398), .QN(n7990) );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(n8541), .CLK(n8846), .Q(
        g4664) );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(n8559), .CLK(n8864), .Q(
        g2223) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(n8547), .CLK(n8852), .Q(
        g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(n8607), .CLK(n8912), .Q(
        g6645) );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(n8585), .CLK(n8890), .Q(
        g2016) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(n8601), .CLK(n8906), .Q(
        g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(n8601), .CLK(n8906), .Q(
        g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(n8632), .CLK(n8937), .Q(
        g2315) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(n8558), .CLK(n8863), .Q(
        g2811), .QN(n7968) );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(n8593), .CLK(n8898), .Q(
        g5957) );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(n8585), .CLK(n8890), .Q(
        g2047) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(n8601), .CLK(n8906), .Q(
        test_so33), .QN(n8493) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(n8617), .CLK(n8922), 
        .Q(g17760), .QN(n8336) );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(n8540), .CLK(n8845), .Q(
        g5575) );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(n8541), .CLK(n8846), .Q(
        n9327) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(n8541), .CLK(n8846), .Q(
        g3752) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(n8603), .CLK(n8908), .Q(
        g3917) );
  SDFFX1 DFF_480_Q_reg ( .D(test_so86), .SI(g3917), .SE(n8574), .CLK(n8879), 
        .Q(g8783), .QN(DFF_480_n1) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(n8574), .CLK(n8879), .Q(
        g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(n8623), .CLK(n8928), .Q(
        g4388), .QN(n8401) );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(n8639), .CLK(n8944), .Q(
        g6275) );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(n8639), .CLK(n8944), .Q(
        g6311) );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(n8639), .CLK(n8944), .Q(
        g8916) );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(n8553), .CLK(n8858), .Q(
        g1041), .QN(n8435) );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(n8575), .CLK(n8880), .Q(
        test_so34), .QN(n8525) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(n8550), .CLK(n8855), 
        .Q(g2537) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(n8555), .CLK(n8860), .Q(
        g29221), .QN(g23612) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g29221), .SE(n8555), .CLK(n8860), .Q(
        g4430), .QN(n8398) );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(n8592), .CLK(n8897), .Q(
        n9325) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(n8592), .CLK(n8897), .Q(
        g4826), .QN(n8010) );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(n8592), .CLK(n8897), .Q(
        g6239) );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(n8578), .CLK(n8883), .Q(
        g232), .QN(n8329) );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(n8571), .CLK(n8876), .Q(
        g5268) );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(n8571), .CLK(n8876), .Q(
        g6545) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(n8590), .CLK(n8895), .Q(
        n9324) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(n8590), .CLK(n8895), .Q(
        g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(n8634), .CLK(n8939), .Q(
        g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(n8641), .CLK(n8946), .Q(
        test_so35), .QN(n7988) );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(n8582), .CLK(n8887), 
        .Q(g1890) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(n8631), .CLK(n8936), .Q(
        g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(n8595), .CLK(n8900), .Q(
        g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(n8595), .CLK(n8900), .Q(
        g2130) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(n8605), .CLK(n8910), .Q(
        g4108), .QN(n5715) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(n8605), .CLK(n8910), .Q(
        g4308), .QN(n8213) );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(n8581), .CLK(n8886), .Q(
        g475) );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(n8620), .CLK(n8925), .Q(
        g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(n8620), .CLK(n8925), .Q(
        g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(n8539), .CLK(n8844), .Q(
        n9322) );
  SDFFX1 DFF_515_Q_reg ( .D(g24213), .SI(n9322), .SE(n8539), .CLK(n8844), .Q(
        g12184) );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(n8539), .CLK(n8844), .Q(
        g3990), .QN(n5594) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(n8603), .CLK(n8908), .Q(
        test_so36), .QN(n8500) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(n8587), .CLK(n8892), 
        .Q(g1992) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(n8587), .CLK(n8892), .Q(
        g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(n8565), .CLK(n8870), .Q(
        g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(n8630), .CLK(n8935), .Q(
        g832), .QN(n8216) );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(n8598), .CLK(n8903), .Q(
        g5897) );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(n8598), .CLK(n8903), .Q(
        g25689) );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(n8591), .CLK(n8896), .Q(
        g4571) );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(n8635), .CLK(n8940), .Q(
        g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(n8635), .CLK(n8940), .Q(
        g4455) );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(n8564), .CLK(n8869), .Q(
        g2902), .QN(n8038) );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(n8625), .CLK(n8930), .Q(
        g333) );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(n8625), .CLK(n8930), .Q(
        g168) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(n8558), .CLK(n8863), .Q(
        test_so37) );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(n8563), .CLK(n8868), 
        .Q(g3684) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(n8540), .CLK(n8845), .Q(
        g3639), .QN(n5591) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(n8626), .CLK(n8931), .Q(
        g14597) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(n8608), .CLK(n8913), .Q(
        g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(n8581), .CLK(n8886), .Q(
        g5406) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(n8581), .CLK(n8886), .Q(
        g269), .QN(n8331) );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(n8641), .CLK(n8946), .Q(
        g401) );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(n8641), .CLK(n8946), .Q(
        g6040), .QN(n8086) );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(n8581), .CLK(n8886), .Q(
        g441) );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(n8632), .CLK(n8937), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(n8543), .CLK(n8848), .Q(
        g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(n8543), .CLK(n8848), .Q(
        g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(n8618), .CLK(n8923), .Q(
        test_so38), .QN(n8506) );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(n8564), .CLK(n8869), 
        .Q(g3957) );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(n8600), .CLK(n8905), .Q(
        g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(n8590), .CLK(n8895), .Q(
        g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(n8617), .CLK(n8922), .Q(
        g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(n8576), .CLK(n8881), .Q(
        g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(n8614), .CLK(n8919), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(n8614), .CLK(n8919), .Q(
        g3498), .QN(n5740) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(n8595), .CLK(n8900), .Q(
        g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(n8604), .CLK(n8909), .Q(
        g14201) );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(n8618), .CLK(n8923), .Q(
        g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(n8618), .CLK(n8923), .Q(
        g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(n8632), .CLK(n8937), .Q(
        g1608) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(n8632), .CLK(n8937), .Q(
        test_so39), .QN(n8320) );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(n8626), .CLK(n8931), 
        .Q(g17577), .QN(n8373) );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(n8628), .CLK(n8933), .Q(
        g1779) );
  SDFFX1 DFF_568_Q_reg ( .D(g29255), .SI(g1779), .SE(n8642), .CLK(n8947), .Q(
        g2652), .QN(n8293) );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(n8558), .CLK(n8863), .Q(
        g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(n8590), .CLK(n8895), .Q(
        g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(n8609), .CLK(n8914), .Q(
        g661) );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(n8540), .CLK(n8845), .Q(
        g4950) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(n8540), .CLK(n8845), .Q(
        g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(n8558), .CLK(n8863), .Q(
        g2834), .QN(g23652) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(n8546), .CLK(n8851), .Q(
        g1361), .QN(n8325) );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(n8608), .CLK(n8913), .Q(
        g6235) );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(n8634), .CLK(n8939), .Q(
        g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(n8618), .CLK(n8923), .Q(
        test_so40) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(n8575), .CLK(n8880), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(n8545), .CLK(n8850), .Q(
        g1696), .QN(n5628) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(n8603), .CLK(n8908), .Q(
        g6555), .QN(n8314) );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(n8603), .CLK(n8908), .Q(
        g14189) );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(n8603), .CLK(n8908), .Q(
        g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(n8591), .CLK(n8896), .Q(
        g6621) );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(n8544), .CLK(n8849), .Q(
        g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(n8604), .CLK(n8909), .Q(
        g3897) );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(n8568), .CLK(n8873), .Q(
        g538) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(n8586), .CLK(n8891), .Q(
        g2606), .QN(n5311) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(n8550), .CLK(n8855), .Q(
        g1472), .QN(n5290) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(n8555), .CLK(n8860), .Q(
        test_so41) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(n8611), .CLK(n8916), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(n8599), .CLK(n8904), .Q(
        g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(n8599), .CLK(n8904), .Q(
        g13259), .QN(n8418) );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(n8621), .CLK(n8926), .Q(
        g405), .QN(n8345) );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(n8571), .CLK(n8876), .Q(
        g5216) );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(n8624), .CLK(n8929), .Q(
        g6494), .QN(n7987) );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(n8541), .CLK(n8846), .Q(
        g4669) );
  SDFFX1 DFF_606_Q_reg ( .D(g24243), .SI(g4669), .SE(n8619), .CLK(n8924), .Q(
        g996) );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(n8541), .CLK(n8846), .Q(
        g4531), .QN(n8412) );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(n8561), .CLK(n8866), .Q(
        g2860) );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(n8548), .CLK(n8853), .Q(
        g4743) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(n8607), .CLK(n8912), .Q(
        g6593) );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(n8607), .CLK(n8912), .Q(
        test_so42), .QN(n8218) );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(n8556), .CLK(n8861), 
        .Q(g4411) );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(n8546), .CLK(n8851), .Q(
        g1413), .QN(n8461) );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(n8619), .CLK(n8924), 
        .Q(g26960) );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(n8626), .CLK(n8931), .Q(
        g13039), .QN(n8374) );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(n8627), .CLK(n8932), .Q(
        g6641) );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(n8627), .CLK(n8932), .Q(
        g6) );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(n8610), .CLK(n8915), .Q(
        g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n8471), .SI(g1936), .SE(n8610), .CLK(n8915), .Q(
        g55) );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(n8609), .CLK(n8914), .Q(
        g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(n8575), .CLK(n8880), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(n8620), .CLK(n8925), .Q(
        g4480) );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(n8632), .CLK(n8937), .Q(
        n9314) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(n8580), .CLK(n8885), .Q(
        test_so43) );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(n8544), .CLK(n8849), 
        .Q(g5571) );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(n8581), .CLK(n8886), .Q(
        g3578) );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(n8581), .CLK(n8886), .Q(
        g9555) );
  SDFFX1 DFF_632_Q_reg ( .D(g29294), .SI(g9555), .SE(n8579), .CLK(n8884), .Q(
        g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(n8580), .CLK(n8885), .Q(
        g3582) );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(n8592), .CLK(n8897), .Q(
        g6271) );
  SDFFX1 DFF_635_Q_reg ( .D(g34028), .SI(g6271), .SE(n8619), .CLK(n8924), .Q(
        g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(n8590), .CLK(n8895), .Q(
        g2380), .QN(n8002) );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(n8612), .CLK(n8917), .Q(
        g5196) );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(n8636), .CLK(n8941), .Q(
        g3227) );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(n8584), .CLK(n8889), .Q(
        n9312) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(n8601), .CLK(n8906), .Q(
        g14518), .QN(n8383) );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(n8601), .CLK(n8906), .Q(
        test_so44), .QN(n8509) );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(n8625), .CLK(n8930), 
        .Q(g6541), .QN(n5739) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(n8609), .CLK(n8914), .Q(
        g3203) );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(n8631), .CLK(n8936), .Q(
        g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(n8557), .CLK(n8862), .Q(
        g4760) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(n8557), .CLK(n8862), .Q(
        g262), .QN(n8333) );
  SDFFX1 DFF_649_Q_reg ( .D(g33556), .SI(g262), .SE(n8627), .CLK(n8932), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(n8565), .CLK(n8870), .Q(
        g5467), .QN(n8395) );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(n8565), .CLK(n8870), .Q(
        g460) );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(n8608), .CLK(n8913), .Q(
        g6209), .QN(n8312) );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(n8626), .CLK(n8931), .Q(
        g29211), .QN(n8359) );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g29211), .SE(n8626), .CLK(n8931), .Q(
        g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(n8632), .CLK(n8937), .Q(
        g655), .QN(n8454) );
  SDFFX1 DFF_657_Q_reg ( .D(g34626), .SI(g655), .SE(n8632), .CLK(n8937), .Q(
        test_so45) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(n8557), .CLK(n8862), 
        .Q(g2204), .QN(n5620) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(n8612), .CLK(n8917), .Q(
        g5256) );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(n8616), .CLK(n8921), .Q(
        g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(n8579), .CLK(n8884), .Q(
        g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(n8633), .CLK(n8938), .Q(
        g13906) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(n8563), .CLK(n8868), .Q(
        g4423) );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(n8563), .CLK(n8868), .Q(
        g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(n8599), .CLK(n8904), .Q(
        g5685) );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(n8566), .CLK(n8871), .Q(
        g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(n8577), .CLK(n8882), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(n8606), .CLK(n8911), .Q(
        g3247) );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(n8586), .CLK(n8891), .Q(
        g2040), .QN(n5505) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(n8586), .CLK(n8891), .Q(
        test_so46) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(n8570), .CLK(n8875), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(n8618), .CLK(n8923), .Q(
        g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(n8619), .CLK(n8924), .Q(
        g7916), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g7916), .SE(n8615), .CLK(n8920), .Q(
        g4732) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(n8615), .CLK(n8920), .Q(
        g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(n8547), .CLK(n8852), .Q(
        g5817), .QN(n8452) );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(n8610), .CLK(n8915), .Q(
        g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(n8640), .CLK(n8945), .Q(
        g2648), .QN(n8006) );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(n8640), .CLK(n8945), .Q(
        g6736), .QN(n8423) );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(n8540), .CLK(n8845), .Q(
        g4944) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(n8623), .CLK(n8928), .Q(
        g4072) );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(n8625), .CLK(n8930), .Q(
        g7540) );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(n8641), .CLK(n8946), .Q(
        test_so47) );
  SDFFX1 DFF_688_Q_reg ( .D(g29264), .SI(test_si48), .SE(n8544), .CLK(n8849), 
        .Q(g3466), .QN(n8430) );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(n8605), .CLK(n8910), .Q(
        g4116) );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(n8634), .CLK(n8939), .Q(
        g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(n8555), .CLK(n8860), .Q(
        g4434), .QN(n8016) );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(n8642), .CLK(n8947), .Q(
        g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(n8560), .CLK(n8865), .Q(
        g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(n8599), .CLK(n8904), .Q(
        g17813) );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(n8552), .CLK(n8857), .Q(
        g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(n8587), .CLK(n8892), .Q(
        g3333), .QN(n8013) );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(n8587), .CLK(n8892), .Q(
        g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(n8619), .CLK(n8924), .Q(
        g4681), .QN(n8224) );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(n8568), .CLK(n8873), .Q(
        g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(n8631), .CLK(n8936), .Q(
        test_so48), .QN(n8530) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(n8587), .CLK(n8892), 
        .Q(g8789), .QN(n8323) );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(n8587), .CLK(n8892), .Q(
        g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(n8561), .CLK(n8866), .Q(
        g2988) );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(n8602), .CLK(n8907), .Q(
        g3538) );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(n8576), .CLK(n8881), .Q(
        g301) );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(n8576), .CLK(n8881), .Q(
        n9306), .QN(DFF_709_n1) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(n8576), .CLK(n8881), .Q(
        g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(n8576), .CLK(n8881), .Q(
        g17291), .QN(n8369) );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(n8586), .CLK(n8891), .Q(
        g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(n8639), .CLK(n8944), .Q(
        g5011) );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(n8642), .CLK(n8947), .Q(
        g199) );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(n8560), .CLK(n8865), .Q(
        g6523), .QN(n5870) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(n8622), .CLK(n8927), .Q(
        test_so49), .QN(n8490) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(n8616), .CLK(n8921), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(n8565), .CLK(n8870), .Q(
        g854) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(n8622), .CLK(n8927), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(n8608), .CLK(n8913), .Q(
        g4922) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(n8537), .CLK(n8842), .Q(
        g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(n8603), .CLK(n8908), .Q(
        g5863), .QN(n8309) );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(n8620), .CLK(n8925), .Q(
        g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(g29253), .SI(g4581), .SE(n8569), .CLK(n8874), .Q(
        g2518), .QN(n8295) );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(n8569), .CLK(n8874), .Q(
        g2567) );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(n8595), .CLK(n8900), .Q(
        g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(n8607), .CLK(n8912), .Q(
        g3263) );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(n8607), .CLK(n8912), .Q(
        g6613) );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(n8641), .CLK(n8946), .Q(
        test_so50), .QN(n8512) );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(n8624), .CLK(n8929), 
        .Q(g6444) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(n8576), .CLK(n8881), .Q(
        g2965), .QN(n8039) );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(n8603), .CLK(n8908), .Q(
        g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(n8632), .CLK(n8937), .Q(
        n9303) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(n8577), .CLK(n8882), .Q(
        g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(n8596), .CLK(n8901), .Q(
        g17646), .QN(n8431) );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(n8581), .CLK(n8886), .Q(
        g3562) );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(n8547), .CLK(n8852), .Q(
        g10122_Tj), .QN(n8419) );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122_Tj), .SE(n8611), .CLK(n8916), 
        .Q(g1404), .QN(n8427) );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(n8543), .CLK(n8848), .Q(
        g3817), .QN(n8429) );
  SDFFX1 DFF_743_Q_reg ( .D(n8476), .SI(g3817), .SE(n8572), .CLK(n8877), .Q(
        n9302) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(n8572), .CLK(n8877), .Q(
        g4501) );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(n8567), .CLK(n8872), .Q(
        test_so51), .QN(n8524) );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(n8613), .CLK(n8918), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(n8551), .CLK(n8856), .Q(
        g4704) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(n8553), .CLK(n8858), .Q(
        g2878) );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(n8571), .CLK(n8876), .Q(
        g5220) );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(n8596), .CLK(n8901), .Q(
        g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(n8596), .CLK(n8901), .Q(
        g12368) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(n8596), .CLK(n8901), .Q(
        g316) );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(n8639), .CLK(n8944), .Q(
        g1277) );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(n8560), .CLK(n8865), .Q(
        g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(n8625), .CLK(n8930), .Q(
        g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(n8553), .CLK(n8858), .Q(
        g2882) );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(n8567), .CLK(n8872), .Q(
        test_so52) );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(n8610), .CLK(n8915), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(n8610), .CLK(n8915), .Q(
        g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(g34975), .SI(g305), .SE(n8643), .CLK(n8948), .Q(g8) );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(n8558), .CLK(n8863), .Q(
        g2799), .QN(n7965) );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(n8604), .CLK(n8909), .Q(
        g14167) );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(n8626), .CLK(n8931), .Q(
        g17787) );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(n8637), .CLK(n8942), .Q(
        g4912) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(n8570), .CLK(n8875), .Q(
        g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(n8550), .CLK(n8855), .Q(
        g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(n8640), .CLK(n8945), .Q(
        g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(n8555), .CLK(n8860), .Q(
        g550), .QN(n8208) );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(n8578), .CLK(n8883), .Q(
        g255), .QN(n8332) );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(n8640), .CLK(n8945), .Q(
        test_so53), .QN(n8517) );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(n8612), .CLK(n8917), 
        .Q(g5240) );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(n8587), .CLK(n8892), .Q(
        g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(n8601), .CLK(n8906), .Q(
        g3863), .QN(n8310) );
  SDFFX1 DFF_777_Q_reg ( .D(g29245), .SI(g3863), .SE(n8640), .CLK(n8945), .Q(
        g1959), .QN(n8296) );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(n8544), .CLK(n8849), .Q(
        g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(n8591), .CLK(n8896), .Q(
        g6653) );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(n8617), .CLK(n8922), .Q(
        g17764) );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(n8572), .CLK(n8877), .Q(
        g2864) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(n8572), .CLK(n8877), .Q(
        g4894) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(n8599), .CLK(n8904), .Q(
        g17678) );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(n8601), .CLK(n8906), .Q(
        g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(n8601), .CLK(n8906), .Q(
        g16693), .QN(n8382) );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(n8622), .CLK(n8927), .Q(
        test_so54) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(n8553), .CLK(n8858), 
        .Q(g1002), .QN(n8466) );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(n8579), .CLK(n8884), .Q(
        g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(n8579), .CLK(n8884), .Q(
        g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(n8619), .CLK(n8924), .Q(
        g1236), .QN(n8032) );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(n8619), .CLK(n8924), .Q(
        g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(n8619), .CLK(n8924), .Q(
        g2476), .QN(n8443) );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(n8563), .CLK(n8868), .Q(
        g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(n8589), .CLK(n8894), .Q(
        g2375), .QN(n8022) );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(n8541), .CLK(n8846), .Q(
        g63), .QN(n8346) );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(n8547), .CLK(n8852), .Q(
        g17739), .QN(n8338) );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(n8621), .CLK(n8926), .Q(
        g358), .QN(n8458) );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(n8621), .CLK(n8926), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(g28043), .SI(g896), .SE(n8567), .CLK(n8872), .Q(
        test_so55), .QN(n8515) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(n8606), .CLK(n8911), 
        .Q(g3161), .QN(n8315) );
  SDFFX1 DFF_804_Q_reg ( .D(g29251), .SI(g3161), .SE(n8635), .CLK(n8940), .Q(
        g2384), .QN(n8300) );
  SDFFX1 DFF_806_Q_reg ( .D(test_so80), .SI(g2384), .SE(n8600), .CLK(n8905), 
        .Q(g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(n8573), .CLK(n8878), .Q(
        g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(n8591), .CLK(n8896), .Q(
        g4561) );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(n8584), .CLK(n8889), .Q(
        g2024) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(n8562), .CLK(n8867), .Q(
        g3451), .QN(n7975) );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(n8582), .CLK(n8887), .Q(
        g2795), .QN(n7966) );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(n8596), .CLK(n8901), .Q(
        g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(n8542), .CLK(n8847), .Q(
        g4527), .QN(n8185) );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(n8577), .CLK(n8882), .Q(
        g1844) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(n8598), .CLK(n8903), .Q(
        g5937) );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(n8628), .CLK(n8933), .Q(
        test_so56) );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(n8550), .CLK(n8855), 
        .Q(g2523), .QN(n5281) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(n8635), .CLK(n8940), .Q(
        g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(n8586), .CLK(n8891), .Q(
        g2643), .QN(n8021) );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(n8586), .CLK(n8891), .Q(
        g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(n8568), .CLK(n8873), .Q(
        g8358), .QN(n8047) );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(n8550), .CLK(n8855), .Q(
        n9295) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(n8550), .CLK(n8855), .Q(
        g5156), .QN(n5734) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(n8566), .CLK(n8871), .Q(
        g30332), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(g34975), .SI(g30332), .SE(n8561), .CLK(n8866), .Q(
        n9294) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(n8562), .CLK(n8867), .Q(
        g8279) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(n8594), .CLK(n8899), .Q(
        g8839) );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(n8638), .CLK(n8943), .Q(
        g1955), .QN(n7999) );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(n8641), .CLK(n8946), .Q(
        test_so57), .QN(n8503) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(n8559), .CLK(n8864), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(n8617), .CLK(n8922), .Q(
        g14749) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(n8640), .CLK(n8945), .Q(
        g4771) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(n8556), .CLK(n8861), .Q(
        g6098) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(n8606), .CLK(n8911), .Q(
        g3147), .QN(n5738) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(n8637), .CLK(n8942), .Q(
        g3347), .QN(n8413) );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(n8559), .CLK(n8864), .Q(
        g2269) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(n8568), .CLK(n8873), .Q(
        g191), .QN(n8048) );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(n8568), .CLK(n8873), .Q(
        g2712), .QN(n8421) );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(n8596), .CLK(n8901), .Q(
        g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(n8551), .CLK(n8856), .Q(
        g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(n8613), .CLK(n8918), .Q(
        test_so58), .QN(n8505) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(n8585), .CLK(n8890), 
        .Q(g17819) );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(n8640), .CLK(n8945), .Q(
        g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(n8564), .CLK(n8869), .Q(
        g2927), .QN(n8036) );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(n8573), .CLK(n8878), .Q(
        g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(n8593), .CLK(n8898), .Q(
        g5929) );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(n8608), .CLK(n8913), .Q(
        g4907) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(n8608), .CLK(n8913), .Q(
        g16874) );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(n8574), .CLK(n8879), .Q(
        g4035), .QN(n8014) );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(n8574), .CLK(n8879), .Q(
        g2946) );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(n8567), .CLK(n8872), .Q(
        g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(n8623), .CLK(n8928), .Q(
        g4082), .QN(n8348) );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(n8624), .CLK(n8929), .Q(
        g9743) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(n8585), .CLK(n8890), .Q(
        test_so59), .QN(n8526) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(n8595), .CLK(n8900), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(n8632), .CLK(n8937), .Q(
        g1620) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(n8554), .CLK(n8859), .Q(
        g2831), .QN(g30331) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(n8554), .CLK(n8859), .Q(
        g667) );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(n8567), .CLK(n8872), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(n8630), .CLK(n8935), .Q(
        g3937) );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(n8630), .CLK(n8935), .Q(
        g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(n8630), .CLK(n8935), .Q(
        g1249), .QN(n8440) );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(n8565), .CLK(n8870), .Q(
        g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(n8602), .CLK(n8907), .Q(
        g16924) );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(n8595), .CLK(n8900), .Q(
        g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(n8539), .CLK(n8844), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(n8597), .CLK(n8902), .Q(
        test_so60) );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(n8598), .CLK(n8903), 
        .Q(g5949) );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(n8572), .CLK(n8877), .Q(
        g6682), .QN(n5590) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(n8572), .CLK(n8877), .Q(
        g904), .QN(n8441) );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(n8561), .CLK(n8866), .Q(
        g2873), .QN(n5488) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(n8638), .CLK(n8943), .Q(
        g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(n8537), .CLK(n8842), .Q(
        g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(n8544), .CLK(n8849), .Q(
        g5603) );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(n8542), .CLK(n8847), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(n8635), .CLK(n8940), .Q(
        g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(n8635), .CLK(n8940), .Q(
        g2437) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(n8585), .CLK(n8890), .Q(
        g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(n8614), .CLK(n8919), .Q(
        g2208), .QN(n8391) );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(n8570), .CLK(n8875), .Q(
        test_so61) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(n8605), .CLK(n8910), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(n8613), .CLK(n8918), .Q(
        g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(n8613), .CLK(n8918), .Q(
        g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(n8616), .CLK(n8921), .Q(
        g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(n8538), .CLK(n8843), .Q(
        g5583) );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(n8579), .CLK(n8884), .Q(
        g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(n8605), .CLK(n8910), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(n8605), .CLK(n8910), .Q(
        g17743) );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(n8564), .CLK(n8869), .Q(
        g2917), .QN(n8037) );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(n8609), .CLK(n8914), .Q(
        g686) );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(n8588), .CLK(n8893), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(n8554), .CLK(n8859), .Q(
        g671), .QN(n7980) );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(n8640), .CLK(n8945), .Q(
        test_so62), .QN(n8531) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(n8592), .CLK(n8897), 
        .Q(g6283) );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(n8617), .CLK(n8922), .Q(
        g14705) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(n8626), .CLK(n8931), .Q(
        g17519), .QN(n8375) );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(n8626), .CLK(n8931), .Q(
        g8784), .QN(DFF_909_n1) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(n8549), .CLK(n8854), .Q(
        g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(n8636), .CLK(n8941), .Q(
        g4489) );
  SDFFX1 DFF_912_Q_reg ( .D(g33564), .SI(g4489), .SE(n8636), .CLK(n8941), .Q(
        g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(n8589), .CLK(n8894), .Q(
        g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(n8613), .CLK(n8918), .Q(
        g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(n8597), .CLK(n8902), .Q(
        g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(n8565), .CLK(n8870), .Q(
        g3929) );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(n8565), .CLK(n8870), .Q(
        g5503), .QN(n5737) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(n8542), .CLK(n8847), .Q(
        test_so63) );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(n8593), .CLK(n8898), 
        .Q(g5925) );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(n8599), .CLK(n8904), .Q(
        g1124) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(n8539), .CLK(n8844), .Q(
        g4955) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(n8612), .CLK(n8917), .Q(
        g5224) );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(n8584), .CLK(n8889), .Q(
        g2012) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(n8607), .CLK(n8912), .Q(
        g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(n8551), .CLK(n8856), .Q(
        g5120), .QN(n8396) );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(n8626), .CLK(n8931), .Q(
        g17674), .QN(n8341) );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(n8590), .CLK(n8895), .Q(
        g2389), .QN(n5631) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(n8590), .CLK(n8895), .Q(
        g4438) );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(n8635), .CLK(n8940), .Q(
        g2429) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(n8582), .CLK(n8887), .Q(
        g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(n8641), .CLK(n8946), .Q(
        test_so64) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(n8540), .CLK(n8845), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(n8574), .CLK(n8879), .Q(
        g18881) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g18881), .SE(n8574), .CLK(n8879), .Q(
        g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(n8554), .CLK(n8859), .Q(
        g1199), .QN(n8052) );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(n8554), .CLK(n8859), .Q(
        g19357), .QN(n5401) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(n8545), .CLK(n8850), .Q(
        g5547) );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(n8545), .CLK(n8850), .Q(
        g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(n8601), .CLK(n8906), .Q(
        g16744), .QN(n8334) );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(n8629), .CLK(n8934), .Q(
        g2338), .QN(n5310) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(n8629), .CLK(n8934), .Q(
        g8919) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(n8592), .CLK(n8897), .Q(
        g6247) );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(n8582), .CLK(n8887), .Q(
        g2791), .QN(n7967) );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(n8604), .CLK(n8909), .Q(
        test_so65) );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(n8537), .CLK(n8842), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(n8593), .CLK(n8898), .Q(
        g5945) );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(n8593), .CLK(n8898), .Q(
        g5244) );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(n8613), .CLK(n8918), .Q(
        g2759), .QN(n8463) );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(n8572), .CLK(n8877), .Q(
        g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(n8579), .CLK(n8884), .Q(
        g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(n8588), .CLK(n8893), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(n8544), .CLK(n8849), .Q(
        g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(n8568), .CLK(n8873), .Q(
        g209), .QN(n5595) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(n8625), .CLK(n8930), .Q(
        g6609) );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(n8625), .CLK(n8930), .Q(
        g5517), .QN(n8311) );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(n8636), .CLK(n8941), .Q(
        g2449) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(n8574), .CLK(n8879), .Q(
        test_so66) );
  SDFFX1 DFF_961_Q_reg ( .D(g18881), .SI(test_si67), .SE(n8574), .CLK(n8879), 
        .Q(n9281), .QN(DFF_961_n1) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(n8559), .CLK(n8864), .Q(
        g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(n8566), .CLK(n8871), .Q(
        g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(n8585), .CLK(n8890), .Q(
        g2098), .QN(n5280) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(n8618), .CLK(n8923), .Q(
        g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(n8595), .CLK(n8900), .Q(
        g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(n8627), .CLK(n8932), .Q(
        g6589) );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(n8582), .CLK(n8887), .Q(
        n9280) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(n8617), .CLK(n8922), .Q(
        g17845) );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(n8617), .CLK(n8922), .Q(
        g17871) );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(n8582), .CLK(n8887), .Q(
        g429) );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(n8582), .CLK(n8887), .Q(
        g1870) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(n8582), .CLK(n8887), .Q(
        test_so67) );
  SDFFX1 DFF_977_Q_reg ( .D(g29243), .SI(test_si68), .SE(n8639), .CLK(n8944), 
        .Q(g1825), .QN(n8302) );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(n8587), .CLK(n8892), .Q(
        g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(n8588), .CLK(n8893), .Q(
        g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(test_so46), .SI(g4392), .SE(n8588), .CLK(n8893), 
        .Q(g8283), .QN(n8354) );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(n8580), .CLK(n8885), .Q(
        g3546) );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(n8571), .CLK(n8876), .Q(
        g5236) );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(n8590), .CLK(n8895), .Q(
        g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(n8612), .CLK(n8917), .Q(
        g4854) );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(n8564), .CLK(n8869), .Q(
        g3925) );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(n8560), .CLK(n8865), .Q(
        g6509), .QN(n8407) );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(n8578), .CLK(n8883), .Q(
        g732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(n8569), .CLK(n8874), .Q(
        g2504), .QN(n8294) );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(n8569), .CLK(n8874), .Q(
        test_so68), .QN(n8496) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(n8542), .CLK(n8847), 
        .Q(g4520) );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(n8542), .CLK(n8847), .Q(
        g8917) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(n8613), .CLK(n8918), .Q(
        g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(n8613), .CLK(n8918), .Q(
        g37), .QN(g30327) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(n8633), .CLK(n8938), .Q(
        g4031) );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(n8586), .CLK(n8891), .Q(
        g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(n8616), .CLK(n8921), .Q(
        g8235), .QN(n8352) );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(n8570), .CLK(n8875), .Q(
        g4176) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(n8549), .CLK(n8854), .Q(
        g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(n8589), .CLK(n8894), .Q(
        g4405) );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(n8604), .CLK(n8909), .Q(
        g872) );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(n8549), .CLK(n8854), .Q(
        g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(n8637), .CLK(n8942), .Q(
        test_so69), .QN(n8495) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(n8548), .CLK(n8853), 
        .Q(g4765) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(n8538), .CLK(n8843), .Q(
        g5563) );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(n8611), .CLK(n8916), .Q(
        g1395), .QN(n8134) );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(n8609), .CLK(n8914), .Q(
        g1913) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(n8629), .CLK(n8934), .Q(
        g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(n8597), .CLK(n8902), .Q(
        g6263) );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(n8542), .CLK(n8847), .Q(
        n9276) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(n8542), .CLK(n8847), .Q(
        g3945) );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(n8625), .CLK(n8930), .Q(
        g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(n8620), .CLK(n8925), .Q(
        g4473), .QN(n8422) );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(n8630), .CLK(n8935), .Q(
        g1266), .QN(n8042) );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(n8642), .CLK(n8947), .Q(
        g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(n8555), .CLK(n8860), .Q(
        test_so70), .QN(n8521) );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(n8613), .CLK(n8918), 
        .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(n8539), .CLK(n8844), .Q(
        g5471), .QN(n8450) );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(n8620), .CLK(n8925), .Q(
        g4540) );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(n8621), .CLK(n8926), .Q(
        g6723) );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(n8637), .CLK(n8942), .Q(
        g6605) );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(n8569), .CLK(n8874), .Q(
        n9274) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(n8557), .CLK(n8862), .Q(
        g2173) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(n8594), .CLK(n8899), .Q(
        g9019) );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(n8594), .CLK(n8899), .Q(
        g2491) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(n8612), .CLK(n8917), .Q(
        g4849), .QN(n8436) );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(n8584), .CLK(n8889), .Q(
        g2169) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(n8559), .CLK(n8864), .Q(
        n9273) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(n8559), .CLK(n8864), .Q(
        test_so71) );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(n8554), .CLK(n8859), 
        .Q(g29219) );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g29219), .SE(n8590), .CLK(n8895), 
        .Q(g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(n8561), .CLK(n8866), .Q(
        g2868), .QN(n8351) );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(n8583), .CLK(n8888), .Q(
        g2767), .QN(n7970) );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(n8615), .CLK(n8920), .Q(
        g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(n8615), .CLK(n8920), .Q(
        g16718), .QN(n8335) );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(n8589), .CLK(n8894), 
        .Q(g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(n8594), .CLK(n8899), .Q(
        g5212) );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(n8594), .CLK(n8899), .Q(
        g4245) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(n8594), .CLK(n8899), .Q(
        g645), .QN(n8316) );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(n8594), .CLK(n8899), .Q(
        g4291), .QN(n8211) );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(n8566), .CLK(n8871), .Q(
        g29212), .QN(n5657) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g29212), .SE(n8566), .CLK(n8871), 
        .Q(test_so72) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(n8599), .CLK(n8904), 
        .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(n8587), .CLK(n8892), .Q(
        g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(n8587), .CLK(n8892), .Q(
        g8788), .QN(n8322) );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(n8583), .CLK(n8888), .Q(
        g2246), .QN(n8005) );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(n8577), .CLK(n8882), .Q(
        g1830), .QN(n5413) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(n8580), .CLK(n8885), .Q(
        g3590) );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(n8566), .CLK(n8871), .Q(
        g392), .QN(n8344) );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(n8631), .CLK(n8936), .Q(
        g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(n8631), .CLK(n8936), .Q(
        g6505), .QN(n8365) );
  SDFFX1 DFF_1057_Q_reg ( .D(g24246), .SI(g6505), .SE(n8631), .CLK(n8936), .Q(
        g1221), .QN(n8400) );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(n8598), .CLK(n8903), .Q(
        g5921) );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(n8575), .CLK(n8880), .Q(
        g29216) );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g29216), .SE(n8575), .CLK(n8880), 
        .Q(test_so73) );
  SDFFX1 DFF_1061_Q_reg ( .D(test_so42), .SI(test_si74), .SE(n8607), .CLK(
        n8912), .Q(g218), .QN(n8219) );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(n8607), .CLK(n8912), .Q(
        g1932) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(n8614), .CLK(n8919), .Q(
        g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(n8632), .CLK(n8937), .Q(
        g5062), .QN(n8438) );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(n8538), .CLK(n8843), .Q(
        g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(n8539), .CLK(n8844), .Q(
        g2689) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(n8623), .CLK(n8928), .Q(
        g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(n8563), .CLK(n8868), .Q(
        g1677), .QN(n8299) );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(n8585), .CLK(n8890), .Q(
        g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(n8540), .CLK(n8845), .Q(
        g2671) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(n8589), .CLK(n8894), .Q(
        g10527) );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(n8589), .CLK(n8894), 
        .Q(g7243) );
  SDFFX1 DFF_1074_Q_reg ( .D(n8471), .SI(g7243), .SE(n8610), .CLK(n8915), .Q(
        test_so74) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(n8577), .CLK(n8882), 
        .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(n8537), .CLK(n8842), .Q(
        g29213), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g29213), .SE(n8537), .CLK(n8842), 
        .Q(g5485), .QN(n5869) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(n8596), .CLK(n8901), .Q(
        g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(n8597), .CLK(n8902), .Q(
        g11678), .QN(n5482) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(n8570), .CLK(n8875), 
        .Q(g2638), .QN(n8292) );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(n8570), .CLK(n8875), .Q(
        g4122) );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(n8614), .CLK(n8919), .Q(
        g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(n8593), .CLK(n8898), .Q(
        g5941) );
  SDFFX1 DFF_1086_Q_reg ( .D(g33572), .SI(g5941), .SE(n8585), .CLK(n8890), .Q(
        g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(n8585), .CLK(n8890), .Q(
        g13068), .QN(n8432) );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(n8585), .CLK(n8890), .Q(
        g25), .QN(n8350) );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(n8576), .CLK(n8881), .Q(
        test_so75) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(n8595), .CLK(n8900), 
        .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(n8559), .CLK(n8864), .Q(
        g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(n8554), .CLK(n8859), .Q(
        n9267) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(n8554), .CLK(n8859), .Q(
        g2066) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(n8634), .CLK(n8939), .Q(
        g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(n8571), .CLK(n8876), .Q(
        g5252) );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(n8584), .CLK(n8889), .Q(
        g2165) );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(n8569), .CLK(n8874), .Q(
        g2571) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(n8611), .CLK(n8916), .Q(
        g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(n8611), .CLK(n8916), .Q(
        g8403), .QN(n8355) );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(n8585), .CLK(n8890), .Q(
        g14673) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(n8585), .CLK(n8890), 
        .Q(test_so76), .QN(n8507) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(n8558), .CLK(n8863), 
        .Q(g2827), .QN(n7969) );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(n8604), .CLK(n8909), .Q(
        g14217) );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(n8612), .CLK(n8917), 
        .Q(g4859) );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(n8621), .CLK(n8926), .Q(
        g424) );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(n8589), .CLK(n8894), .Q(
        g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(n8589), .CLK(n8894), .Q(
        g17423), .QN(n8404) );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(n8638), .CLK(n8943), 
        .Q(n9265), .QN(n6006) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(n8558), .CLK(n8863), .Q(
        g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(n8577), .CLK(n8882), .Q(
        g1821), .QN(n8000) );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(n8550), .CLK(n8855), .Q(
        g2509), .QN(n8020) );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(n8537), .CLK(n8842), .Q(
        g5073), .QN(n8392) );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(n8588), .CLK(n8893), .Q(
        test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(n8616), .CLK(n8921), 
        .Q(g8353), .QN(n8353) );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(n8617), .CLK(n8922), .Q(
        g13085), .QN(n8377) );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(n8637), .CLK(n8942), 
        .Q(g6633) );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(n8551), .CLK(n8856), .Q(
        g5124), .QN(n8457) );
  SDFFX1 DFF_1122_Q_reg ( .D(test_so44), .SI(g5124), .SE(n8601), .CLK(n8906), 
        .Q(g17400), .QN(n8368) );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(n8592), .CLK(n8897), 
        .Q(g6303) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(n8537), .CLK(n8842), .Q(
        g5069) );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(n8561), .CLK(n8866), .Q(
        g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(n8630), .CLK(n8935), .Q(
        g650), .QN(n8317) );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(n8630), .CLK(n8935), .Q(
        g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(n8630), .CLK(n8935), .Q(
        g3921) );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(n8630), .CLK(n8935), .Q(
        test_so78), .QN(n8514) );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(n8640), .CLK(n8945), 
        .Q(g6732), .QN(n8179) );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(n8560), .CLK(n8865), .Q(
        g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(n8638), .CLK(n8943), .Q(
        g1061), .QN(n8426) );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(n8638), .CLK(n8943), .Q(
        g3462), .QN(n8393) );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(n8584), .CLK(n8889), .Q(
        g2181) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(n8584), .CLK(n8889), .Q(
        g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(n8628), .CLK(n8933), .Q(
        g1756) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(n8628), .CLK(n8933), .Q(
        g5849), .QN(n5736) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(n8633), .CLK(n8938), .Q(
        g4112) );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(n8540), .CLK(n8845), .Q(
        n9262) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(n8557), .CLK(n8862), .Q(
        g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(n8635), .CLK(n8940), .Q(
        test_so79), .QN(n8501) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(n8553), .CLK(n8858), 
        .Q(g1046), .QN(n8243) );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(n8622), .CLK(n8927), .Q(
        g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(n8622), .CLK(n8927), .Q(
        g4401), .QN(n8015) );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(n8622), .CLK(n8927), .Q(
        g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(n8623), .CLK(n8928), .Q(
        g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(n8623), .CLK(n8928), .Q(
        g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(n8564), .CLK(n8869), .Q(
        g2950), .QN(n8195) );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(n8546), .CLK(n8851), .Q(
        g1345), .QN(n8469) );
  SDFFX1 DFF_1154_Q_reg ( .D(g25762), .SI(g1345), .SE(n8625), .CLK(n8930), .Q(
        g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(n8615), .CLK(n8920), .Q(
        g14421), .QN(n8380) );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(n8615), .CLK(n8920), 
        .Q(g4727) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(n8600), .CLK(n8905), .Q(
        test_so80), .QN(n8497) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(n8546), .CLK(n8851), 
        .Q(g1536), .QN(n7952) );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(n8564), .CLK(n8869), .Q(
        g3941) );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(n8621), .CLK(n8926), .Q(
        g370), .QN(n8307) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(n8548), .CLK(n8853), .Q(
        g5694), .QN(n8088) );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(n8577), .CLK(n8882), .Q(
        g1858) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(n8577), .CLK(n8882), .Q(
        g446) );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(n8606), .CLK(n8911), .Q(
        g3219) );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(n8591), .CLK(n8896), .Q(
        g1811), .QN(n8303) );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(n8591), .CLK(n8896), .Q(
        g6601) );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(n8569), .CLK(n8874), .Q(
        g2441) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(n8638), .CLK(n8943), .Q(
        g1874) );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(n8573), .CLK(n8878), .Q(
        test_so81), .QN(n8492) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(n8624), .CLK(n8929), 
        .Q(g6581) );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(n8607), .CLK(n8912), .Q(
        g6597) );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(n8611), .CLK(n8916), .Q(
        g5008) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(n8562), .CLK(n8867), .Q(
        g3610) );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(n8561), .CLK(n8866), .Q(
        g2890) );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(n8636), .CLK(n8941), .Q(
        g1978) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(n8636), .CLK(n8941), .Q(
        g1612) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(n8586), .CLK(n8891), .Q(
        g112), .QN(n8342) );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(n8541), .CLK(n8846), .Q(
        g2856) );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(n8599), .CLK(n8904), .Q(
        g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(n8599), .CLK(n8904), .Q(
        g17722), .QN(n8385) );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(n8635), .CLK(n8940), 
        .Q(test_so82) );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(n8605), .CLK(n8910), 
        .Q(g4119) );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(n8605), .CLK(n8910), .Q(
        g6390), .QN(n8414) );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(n8546), .CLK(n8851), .Q(
        g1542), .QN(n8051) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(n8546), .CLK(n8851), .Q(
        g4258), .QN(n8428) );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(n8616), .CLK(n8921), .Q(
        g4818) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(n8633), .CLK(n8938), .Q(
        g5033), .QN(n8409) );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(n8615), .CLK(n8920), .Q(
        g4717) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(n8624), .CLK(n8929), .Q(
        g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(n8624), .CLK(n8929), .Q(
        g3849), .QN(n5735) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(n8624), .CLK(n8929), .Q(
        g17778), .QN(n8339) );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(n8609), .CLK(n8914), 
        .Q(g3199) );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(n8643), .CLK(n8948), .Q(
        test_so83) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(n8613), .CLK(n8918), 
        .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(n8579), .CLK(n8884), .Q(
        g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(n8593), .CLK(n8898), .Q(
        g5913) );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(n8582), .CLK(n8887), .Q(
        g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(n8549), .CLK(n8854), .Q(
        g6163), .QN(n8451) );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(n8600), .CLK(n8905), .Q(
        g4125), .QN(n8226) );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(n8640), .CLK(n8945), .Q(
        g4821), .QN(n5880) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(n8552), .CLK(n8857), .Q(
        g4939) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(n8588), .CLK(n8893), .Q(
        g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(n8636), .CLK(n8941), 
        .Q(g3207) );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(n8636), .CLK(n8941), .Q(
        g4483) );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(n8587), .CLK(n8892), .Q(
        test_so84) );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(n8551), .CLK(n8856), 
        .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(n8571), .CLK(n8876), .Q(
        g5248) );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(n8543), .CLK(n8848), .Q(
        g2126) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(n8543), .CLK(n8848), .Q(
        g3694), .QN(n8087) );
  SDFFX1 DFF_1215_Q_reg ( .D(g29288), .SI(g3694), .SE(n8539), .CLK(n8844), .Q(
        g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(n8539), .CLK(n8844), .Q(
        g1964), .QN(n5315) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(n8537), .CLK(n8842), .Q(
        g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(n8606), .CLK(n8911), .Q(
        g3215) );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(n8633), .CLK(n8938), .Q(
        g16748) );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(n8638), .CLK(n8943), 
        .Q(n9255), .QN(n6005) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(n8555), .CLK(n8860), .Q(
        g4427), .QN(n8318) );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(n8555), .CLK(n8860), .Q(
        test_so85) );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(n8583), .CLK(n8888), 
        .Q(g2779), .QN(n7964) );
  SDFFX1 DFF_1224_Q_reg ( .D(test_so39), .SI(g2779), .SE(n8583), .CLK(n8888), 
        .Q(g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(n8583), .CLK(n8888), .Q(
        g7245) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(n8614), .CLK(n8919), .Q(
        g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(n8546), .CLK(n8851), .Q(
        g1367), .QN(n8468) );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(n8633), .CLK(n8938), .Q(
        g5112) );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(n8633), .CLK(n8938), .Q(
        g19), .QN(n8447) );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(n8633), .CLK(n8938), .Q(
        g4145), .QN(n8186) );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(n8584), .CLK(n8889), .Q(
        g2161) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(n8621), .CLK(n8926), .Q(
        g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(n8629), .CLK(n8934), .Q(
        g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(n8574), .CLK(n8879), .Q(
        test_so86), .QN(DFF_1234_n1) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(n8595), .CLK(n8900), 
        .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(n8615), .CLK(n8920), .Q(
        g2051), .QN(n8448) );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(n8554), .CLK(n8859), .Q(
        g1193) );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(n8634), .CLK(n8939), .Q(
        g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(n8567), .CLK(n8872), .Q(
        g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(n8567), .CLK(n8872), .Q(
        g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(n8577), .CLK(n8882), .Q(
        g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(n8641), .CLK(n8946), .Q(
        g3594) );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(n8561), .CLK(n8866), .Q(
        g2999) );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(n8629), .CLK(n8934), .Q(
        g2303) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(n8630), .CLK(n8935), .Q(
        g17688), .QN(n8387) );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(n8630), .CLK(n8935), 
        .Q(test_so87) );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(n8642), .CLK(n8947), 
        .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(n8642), .CLK(n8947), .Q(
        g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(n8568), .CLK(n8873), .Q(
        g546) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(n8568), .CLK(n8873), .Q(
        g2472), .QN(n5619) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(n8598), .CLK(n8903), .Q(
        g5953) );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(n8598), .CLK(n8903), .Q(
        g8277), .QN(n7996) );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(n8627), .CLK(n8932), .Q(
        g1740) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(n8580), .CLK(n8885), .Q(
        g3550) );
  SDFFX1 DFF_1260_Q_reg ( .D(n514), .SI(g3550), .SE(n8543), .CLK(n8848), .Q(
        g3845), .QN(n5886) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(n8543), .CLK(n8848), .Q(
        g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(n8599), .CLK(n8904), .Q(
        g14635) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(n8606), .CLK(n8911), 
        .Q(test_so88) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(n8565), .CLK(n8870), 
        .Q(g3913) );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(n8563), .CLK(n8868), .Q(
        g10306) );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(n8545), .CLK(n8850), 
        .Q(g1687), .QN(n8004) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(n8575), .CLK(n8880), .Q(
        g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(g33596), .SI(g2681), .SE(n8575), .CLK(n8880), .Q(
        g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(n8575), .CLK(n8880), .Q(
        g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(n8575), .CLK(n8880), .Q(
        g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(g31895), .SI(g2697), .SE(n8573), .CLK(n8878), .Q(
        g4417), .QN(n8460) );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(n8600), .CLK(n8905), .Q(
        g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(n8588), .CLK(n8893), .Q(
        g1141) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(n8588), .CLK(n8893), .Q(
        g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(n8634), .CLK(n8939), 
        .Q(test_so89), .QN(n8533) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(n8545), .CLK(n8850), 
        .Q(g1710) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(n8560), .CLK(n8865), .Q(
        g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(n8636), .CLK(n8941), .Q(
        g3255) );
  SDFFX1 DFF_1281_Q_reg ( .D(g29241), .SI(g3255), .SE(n8563), .CLK(n8868), .Q(
        g1691), .QN(n8298) );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(n8563), .CLK(n8868), .Q(
        g2936), .QN(n8196) );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(n8642), .CLK(n8947), .Q(
        g5644), .QN(n5593) );
  SDFFX1 DFF_1284_Q_reg ( .D(n191), .SI(g5644), .SE(n8551), .CLK(n8856), .Q(
        g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(n8551), .CLK(n8856), .Q(
        g5352), .QN(n8444) );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(n8570), .CLK(n8875), .Q(
        g8915) );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(n8583), .CLK(n8888), .Q(
        g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(n8635), .CLK(n8940), .Q(
        g2922), .QN(n8194) );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(n8576), .CLK(n8881), .Q(
        test_so90) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(n8598), .CLK(n8903), 
        .Q(g5893) );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(n8615), .CLK(n8920), .Q(
        g16603), .QN(n8381) );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(n8637), .CLK(n8942), 
        .Q(g6617) );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(n8554), .CLK(n8859), .Q(
        g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(n8563), .CLK(n8868), .Q(
        g4512) );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(n8538), .CLK(n8843), .Q(
        g5599) );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(n8562), .CLK(n8867), .Q(
        g3401) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(n8562), .CLK(n8867), .Q(
        g4366) );
  SDFFX1 DFF_1300_Q_reg ( .D(test_so26), .SI(g4366), .SE(n8602), .CLK(n8907), 
        .Q(g16722) );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(n8614), .CLK(n8919), 
        .Q(g29214) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g29214), .SE(n8552), .CLK(n8857), 
        .Q(g3129), .QN(n5861) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(n8608), .CLK(n8913), .Q(
        test_so91) );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(n8611), .CLK(n8916), 
        .Q(g5170), .QN(n8313) );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(n8611), .CLK(n8916), .Q(
        g26959) );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(n8547), .CLK(n8852), 
        .Q(g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(n8592), .CLK(n8897), .Q(
        g6299) );
  SDFFX1 DFF_1308_Q_reg ( .D(g7916), .SI(g6299), .SE(n8619), .CLK(n8924), .Q(
        g8416), .QN(n8417) );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(n8554), .CLK(n8859), .Q(
        g2079), .QN(n8297) );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(n8551), .CLK(n8856), .Q(
        g4698) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(n8544), .CLK(n8849), .Q(
        g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(n8624), .CLK(n8929), .Q(
        g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(n8642), .CLK(n8947), .Q(
        n9247) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(n8566), .CLK(n8871), .Q(
        g411) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(n8597), .CLK(n8902), .Q(
        test_so92) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(n8631), .CLK(n8936), 
        .Q(g3953) );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(n8631), .CLK(n8936), .Q(
        g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(n8579), .CLK(n8884), .Q(
        g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(n8579), .CLK(n8884), .Q(
        n9245) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(n8623), .CLK(n8928), .Q(
        g1300), .QN(n5483) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(n8623), .CLK(n8928), .Q(
        g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(n8612), .CLK(n8917), .Q(
        g5200) );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(n8612), .CLK(n8917), .Q(
        g4843), .QN(n8360) );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(n8634), .CLK(n8939), .Q(
        g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(g29249), .SI(g5046), .SE(n8559), .CLK(n8864), .Q(
        g2250), .QN(n8304) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(n8623), .CLK(n8928), .Q(
        g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(n8628), .CLK(n8933), 
        .Q(test_so93) );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(n8569), .CLK(n8874), 
        .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(g25734), .SI(g2453), .SE(n8548), .CLK(n8853), .Q(
        g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(n8548), .CLK(n8853), .Q(
        g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(n8610), .CLK(n8915), 
        .Q(g2912), .QN(n8193) );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(n8610), .CLK(n8915), .Q(
        g2357) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(n8629), .CLK(n8934), .Q(
        g8920) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(n8575), .CLK(n8880), .Q(
        g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(n8542), .CLK(n8847), .Q(
        g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(n8634), .CLK(n8939), .Q(
        g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(n8552), .CLK(n8857), .Q(
        g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(n8546), .CLK(n8851), .Q(
        g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(n8583), .CLK(n8888), .Q(
        test_so94), .QN(n8499) );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(n8542), .CLK(n8847), 
        .Q(g4519) );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(n8552), .CLK(n8857), .Q(
        g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(n8552), .CLK(n8857), .Q(
        g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(n8591), .CLK(n8896), .Q(
        g6657) );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(n8591), .CLK(n8896), .Q(
        g4552) );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(n8604), .CLK(n8909), .Q(
        g3893) );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(n8636), .CLK(n8941), .Q(
        g3211) );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(n8599), .CLK(n8904), .Q(
        g13049), .QN(n8371) );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(n8615), .CLK(n8920), 
        .Q(g16624), .QN(n8379) );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(n8538), .CLK(n8843), 
        .Q(g5595) );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(n8562), .CLK(n8867), .Q(
        g3614) );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(n8562), .CLK(n8867), .Q(
        test_so95) );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(n8637), .CLK(n8942), 
        .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(n8608), .CLK(n8913), .Q(
        g16686) );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(n8543), .CLK(n8848), 
        .Q(g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(n8623), .CLK(n8928), .Q(
        g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(n8591), .CLK(n8896), .Q(
        g4570) );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(n8571), .CLK(n8876), .Q(
        g5272) );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(n8596), .CLK(n8901), .Q(
        g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(n8566), .CLK(n8871), .Q(
        g728), .QN(n8055) );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(n8638), .CLK(n8943), .Q(
        g6295) );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(n8540), .CLK(n8845), .Q(
        g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(n8637), .CLK(n8942), .Q(
        g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(n8551), .CLK(n8856), .Q(
        test_so96), .QN(n8516) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(n8624), .CLK(n8929), 
        .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(n8552), .CLK(n8857), .Q(
        g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(n8541), .CLK(n8846), .Q(
        g4659), .QN(n8439) );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(n8541), .CLK(n8846), .Q(
        g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(n8638), .CLK(n8943), .Q(
        g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(n8584), .CLK(n8889), .Q(
        g2084), .QN(n8019) );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(n8606), .CLK(n8911), .Q(
        g3187) );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(n8614), .CLK(n8919), .Q(
        g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(n8569), .CLK(n8874), .Q(
        g2583) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(n8576), .CLK(n8881), .Q(
        n9240) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(n8576), .CLK(n8881), .Q(
        g1094) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(n8603), .CLK(n8908), .Q(
        test_so97), .QN(n8528) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(n8594), .CLK(n8899), 
        .Q(g4284), .QN(n8034) );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(n8606), .CLK(n8911), .Q(
        g3191) );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(n8547), .CLK(n8852), .Q(
        g4239), .QN(n8027) );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(n8587), .CLK(n8892), .Q(
        g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(n8555), .CLK(n8860), .Q(
        g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(n8555), .CLK(n8860), .Q(
        g534) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(n8621), .CLK(n8926), .Q(
        g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(n8584), .CLK(n8889), .Q(
        g2004) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(n8550), .CLK(n8855), .Q(
        g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(n8581), .CLK(n8886), .Q(
        g5456), .QN(n7989) );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(n8572), .CLK(n8877), .Q(
        n6007), .QN(n8319) );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(n8612), .CLK(n8917), .Q(
        test_so98), .QN(n8529) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(n8620), .CLK(n8925), 
        .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(n8551), .CLK(n8856), .Q(
        g5348), .QN(n8180) );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(n8609), .CLK(n8914), .Q(
        g3223) );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(n8564), .CLK(n8869), .Q(
        g2970), .QN(n8192) );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(n8548), .CLK(n8853), .Q(
        g5698), .QN(n8424) );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(n8594), .CLK(n8899), .Q(
        g5260) );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(n8560), .CLK(n8865), .Q(
        g1521) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(n8562), .CLK(n8867), .Q(
        g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(n8552), .CLK(n8857), .Q(
        g3115), .QN(n8408) );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(n8609), .CLK(n8914), .Q(
        g3251) );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(n8573), .CLK(n8878), .Q(
        g12832) );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(n8573), .CLK(n8878), 
        .Q(test_so99), .QN(n8511) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(n8640), .CLK(n8945), 
        .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(n8642), .CLK(n8947), .Q(
        g8342), .QN(n7974) );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(n8542), .CLK(n8847), .Q(
        g4515), .QN(n8223) );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(n8583), .CLK(n8888), .Q(
        g8787), .QN(n8321) );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(n8542), .CLK(n8847), .Q(
        g4300) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(n8545), .CLK(n8850), .Q(
        n9236) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(n8545), .CLK(n8850), .Q(
        g1379), .QN(n8467) );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(n8602), .CLK(n8907), .Q(
        g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(n8582), .CLK(n8887), 
        .Q(g1878) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(n8538), .CLK(n8843), .Q(
        g5619) );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(n8539), .CLK(n8844), .Q(
        g71), .QN(n8289) );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(n8572), .CLK(n8877), .Q(
        test_so100) );
  SDFFX1 DFF_748_Q_reg ( .D(n1338), .SI(g4704), .SE(n8610), .CLK(n8915), .Q(
        g22), .QN(n8459) );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(n8622), .CLK(n8927), .Q(
        g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(n8596), .CLK(n8901), .Q(
        g2729), .QN(n8347) );
  HADDX1 Trojan_U1_1_30 ( .A0(counter_30), .B0(carry_30), .C1(carry_31), .SO(
        N31) );
  HADDX1 Trojan_U1_1_4 ( .A0(counter_4), .B0(carry_4), .C1(carry_5), .SO(N5)
         );
  HADDX1 Trojan_U1_1_5 ( .A0(counter_5), .B0(carry_5), .C1(carry_6), .SO(N6)
         );
  HADDX1 Trojan_U1_1_6 ( .A0(counter_6), .B0(carry_6), .C1(carry_7), .SO(N7)
         );
  HADDX1 Trojan_U1_1_7 ( .A0(counter_7), .B0(carry_7), .C1(carry_8), .SO(N8)
         );
  HADDX1 Trojan_U1_1_8 ( .A0(counter_8), .B0(carry_8), .C1(carry_9), .SO(N9)
         );
  HADDX1 Trojan_U1_1_9 ( .A0(counter_9), .B0(carry_9), .C1(carry_10), .SO(N10)
         );
  HADDX1 Trojan_U1_1_10 ( .A0(counter_10), .B0(carry_10), .C1(carry_11), .SO(
        N11) );
  HADDX1 Trojan_U1_1_11 ( .A0(counter_11), .B0(carry_11), .C1(carry_12), .SO(
        N12) );
  HADDX1 Trojan_U1_1_12 ( .A0(counter_12), .B0(carry_12), .C1(carry_13), .SO(
        N13) );
  HADDX1 Trojan_U1_1_13 ( .A0(counter_13), .B0(carry_13), .C1(carry_14), .SO(
        N14) );
  HADDX1 Trojan_U1_1_14 ( .A0(counter_14), .B0(carry_14), .C1(carry_15), .SO(
        N15) );
  HADDX1 Trojan_U1_1_22 ( .A0(counter_22), .B0(carry_22), .C1(carry_23), .SO(
        N23) );
  HADDX1 Trojan_U1_1_23 ( .A0(counter_23), .B0(carry_23), .C1(carry_24), .SO(
        N24) );
  HADDX1 Trojan_U1_1_24 ( .A0(counter_24), .B0(carry_24), .C1(carry_25), .SO(
        N25) );
  HADDX1 Trojan_U1_1_25 ( .A0(counter_25), .B0(carry_25), .C1(carry_26), .SO(
        N26) );
  HADDX1 Trojan_U1_1_1 ( .A0(counter_1), .B0(counter_0), .C1(carry_2), .SO(N2)
         );
  HADDX1 Trojan_U1_1_2 ( .A0(counter_2), .B0(carry_2), .C1(carry_3), .SO(N3)
         );
  HADDX1 Trojan_U1_1_3 ( .A0(counter_3), .B0(carry_3), .C1(carry_4), .SO(N4)
         );
  HADDX1 Trojan_U1_1_15 ( .A0(counter_15), .B0(carry_15), .C1(carry_16), .SO(
        N16) );
  HADDX1 Trojan_U1_1_16 ( .A0(counter_16), .B0(carry_16), .C1(carry_17), .SO(
        N17) );
  HADDX1 Trojan_U1_1_17 ( .A0(counter_17), .B0(carry_17), .C1(carry_18), .SO(
        N18) );
  HADDX1 Trojan_U1_1_18 ( .A0(counter_18), .B0(carry_18), .C1(carry_19), .SO(
        N19) );
  HADDX1 Trojan_U1_1_19 ( .A0(counter_19), .B0(carry_19), .C1(carry_20), .SO(
        N20) );
  HADDX1 Trojan_U1_1_20 ( .A0(counter_20), .B0(carry_20), .C1(carry_21), .SO(
        N21) );
  HADDX1 Trojan_U1_1_21 ( .A0(counter_21), .B0(carry_21), .C1(carry_22), .SO(
        N22) );
  HADDX1 Trojan_U1_1_26 ( .A0(counter_26), .B0(carry_26), .C1(carry_27), .SO(
        N27) );
  HADDX1 Trojan_U1_1_27 ( .A0(counter_27), .B0(carry_27), .C1(carry_28), .SO(
        N28) );
  HADDX1 Trojan_U1_1_28 ( .A0(counter_28), .B0(carry_28), .C1(carry_29), .SO(
        N29) );
  HADDX1 Trojan_U1_1_29 ( .A0(counter_29), .B0(carry_29), .C1(carry_30), .SO(
        N30) );
  INVX0 Trojan_U1 ( .INP(counter_0), .ZN(N1) );
  XOR2X1 Trojan_U2 ( .IN1(carry_31), .IN2(counter_31), .Q(N32) );
  DFFARX1 Trojan_counter_reg_31_ ( .D(N32), .CLK(n37), .RSTB(n8536), .Q(
        counter_31), .QN(n73) );
  DFFARX1 Trojan_counter_reg_1_ ( .D(N2), .CLK(n37), .RSTB(n8535), .Q(
        counter_1) );
  DFFARX1 Trojan_counter_reg_2_ ( .D(N3), .CLK(n37), .RSTB(n87), .Q(counter_2)
         );
  DFFARX1 Trojan_counter_reg_3_ ( .D(N4), .CLK(n37), .RSTB(n8536), .Q(
        counter_3), .QN(n86) );
  DFFARX1 Trojan_counter_reg_15_ ( .D(N16), .CLK(n37), .RSTB(n8535), .Q(
        counter_15), .QN(n85) );
  DFFARX1 Trojan_counter_reg_16_ ( .D(N17), .CLK(n37), .RSTB(n87), .Q(
        counter_16), .QN(n84) );
  DFFARX1 Trojan_counter_reg_17_ ( .D(N18), .CLK(n37), .RSTB(n8536), .Q(
        counter_17), .QN(n83) );
  DFFARX1 Trojan_counter_reg_18_ ( .D(N19), .CLK(n37), .RSTB(n8535), .Q(
        counter_18), .QN(n82) );
  DFFARX1 Trojan_counter_reg_19_ ( .D(N20), .CLK(n37), .RSTB(n87), .Q(
        counter_19), .QN(n81) );
  DFFARX1 Trojan_counter_reg_20_ ( .D(N21), .CLK(n37), .RSTB(n8536), .Q(
        counter_20), .QN(n80) );
  DFFARX1 Trojan_counter_reg_21_ ( .D(N22), .CLK(n37), .RSTB(n8535), .Q(
        counter_21), .QN(n79) );
  DFFARX1 Trojan_counter_reg_26_ ( .D(N27), .CLK(n37), .RSTB(n87), .Q(
        counter_26), .QN(n78) );
  DFFARX1 Trojan_counter_reg_27_ ( .D(N28), .CLK(n37), .RSTB(n8536), .Q(
        counter_27), .QN(n77) );
  DFFARX1 Trojan_counter_reg_28_ ( .D(N29), .CLK(n37), .RSTB(n8535), .Q(
        counter_28), .QN(n76) );
  DFFARX1 Trojan_counter_reg_29_ ( .D(N30), .CLK(n37), .RSTB(n87), .Q(
        counter_29), .QN(n75) );
  DFFARX1 Trojan_counter_reg_30_ ( .D(N31), .CLK(n37), .RSTB(n8536), .Q(
        counter_30), .QN(n74) );
  DFFARX1 Trojan_counter_reg_7_ ( .D(N8), .CLK(n37), .RSTB(n8535), .Q(
        counter_7) );
  DFFARX1 Trojan_counter_reg_11_ ( .D(N12), .CLK(n37), .RSTB(n87), .Q(
        counter_11) );
  DFFARX1 Trojan_counter_reg_25_ ( .D(N26), .CLK(n37), .RSTB(n8536), .Q(
        counter_25) );
  DFFARX1 Trojan_counter_reg_6_ ( .D(N7), .CLK(n37), .RSTB(n8535), .Q(
        counter_6) );
  DFFARX1 Trojan_counter_reg_10_ ( .D(N11), .CLK(n37), .RSTB(n87), .Q(
        counter_10) );
  DFFARX1 Trojan_counter_reg_12_ ( .D(N13), .CLK(n37), .RSTB(n8536), .Q(
        counter_12) );
  DFFARX1 Trojan_counter_reg_24_ ( .D(N25), .CLK(n37), .RSTB(n8535), .Q(
        counter_24) );
  DFFARX1 Trojan_counter_reg_4_ ( .D(N5), .CLK(n37), .RSTB(n87), .Q(counter_4)
         );
  DFFARX1 Trojan_counter_reg_5_ ( .D(N6), .CLK(n37), .RSTB(n8536), .Q(
        counter_5) );
  DFFARX1 Trojan_counter_reg_9_ ( .D(N10), .CLK(n37), .RSTB(n8535), .Q(
        counter_9) );
  DFFARX1 Trojan_counter_reg_14_ ( .D(N15), .CLK(n37), .RSTB(n87), .Q(
        counter_14) );
  DFFARX1 Trojan_counter_reg_23_ ( .D(N24), .CLK(n37), .RSTB(n8536), .Q(
        counter_23) );
  DFFARX1 Trojan_counter_reg_8_ ( .D(N9), .CLK(n37), .RSTB(n8535), .Q(
        counter_8) );
  DFFARX1 Trojan_counter_reg_13_ ( .D(N14), .CLK(n37), .RSTB(n87), .Q(
        counter_13) );
  DFFARX1 Trojan_counter_reg_22_ ( .D(N23), .CLK(n37), .RSTB(n8536), .Q(
        counter_22) );
  DFFARX1 Trojan_counter_reg_0_ ( .D(N1), .CLK(n37), .RSTB(n8535), .Q(
        counter_0) );
  NAND4X0 Trojan_U14 ( .IN1(n240), .IN2(n495), .IN3(n310), .IN4(n58), .QN(n87)
         );
  INVX0 Trojan_U15 ( .INP(n59), .ZN(n58) );
  NOR4X0 Trojan_U16 ( .IN1(n240), .IN2(n495), .IN3(n310), .IN4(n59), .QN(n37)
         );
  NAND3X0 Trojan_U17 ( .IN1(n2601), .IN2(n5111), .IN3(n60), .QN(n59) );
  AND3X1 Trojan_U18 ( .IN1(n2396), .IN2(n3279), .IN3(n8473), .Q(n60) );
  NOR4X0 Trojan_U19 ( .IN1(n61), .IN2(n62), .IN3(n63), .IN4(n64), .QN(
        Trigger_out) );
  NAND4X0 Trojan_U20 ( .IN1(n78), .IN2(n77), .IN3(n76), .IN4(n75), .QN(n64) );
  NAND4X0 Trojan_U21 ( .IN1(n74), .IN2(n73), .IN3(counter_6), .IN4(counter_5), 
        .QN(n63) );
  NAND4X0 Trojan_U22 ( .IN1(n80), .IN2(n79), .IN3(n81), .IN4(n65), .QN(n62) );
  NOR4X0 Trojan_U23 ( .IN1(counter_25), .IN2(counter_24), .IN3(counter_23), 
        .IN4(counter_22), .QN(n65) );
  NAND4X0 Trojan_U24 ( .IN1(n66), .IN2(n67), .IN3(n68), .IN4(n69), .QN(n61) );
  NOR4X0 Trojan_U25 ( .IN1(n70), .IN2(counter_12), .IN3(counter_14), .IN4(
        counter_13), .QN(n69) );
  NAND4X0 Trojan_U26 ( .IN1(n85), .IN2(n84), .IN3(n83), .IN4(n82), .QN(n70) );
  NOR4X0 Trojan_U27 ( .IN1(counter_11), .IN2(counter_10), .IN3(counter_9), 
        .IN4(counter_8), .QN(n68) );
  MUX21X1 Trojan_U28 ( .IN1(n71), .IN2(n72), .S(n86), .Q(n67) );
  OA21X1 Trojan_U29 ( .IN1(counter_1), .IN2(counter_0), .IN3(counter_2), .Q(
        n72) );
  NAND2X0 Trojan_U30 ( .IN1(counter_2), .IN2(counter_1), .QN(n71) );
  NOR2X0 Trojan_U31 ( .IN1(counter_7), .IN2(counter_4), .QN(n66) );
  MUX21X1 Trojan_Paylod ( .IN1(g10122_Tj), .IN2(g25715), .S(Trigger_out), .Q(
        g10122) );
  INVX0 U8468 ( .INP(n87), .ZN(n8534) );
  INVX0 U8469 ( .INP(n8534), .ZN(n8535) );
  INVX0 U8470 ( .INP(n8534), .ZN(n8536) );
  NBUFFX2 U8471 ( .INP(n8665), .Z(n8538) );
  NBUFFX2 U8472 ( .INP(n8665), .Z(n8537) );
  NBUFFX2 U8473 ( .INP(n8655), .Z(n8587) );
  NBUFFX2 U8474 ( .INP(n8655), .Z(n8585) );
  NBUFFX2 U8475 ( .INP(n8646), .Z(n8632) );
  NBUFFX2 U8476 ( .INP(n8662), .Z(n8551) );
  NBUFFX2 U8477 ( .INP(n8650), .Z(n8613) );
  NBUFFX2 U8478 ( .INP(n8647), .Z(n8624) );
  NBUFFX2 U8479 ( .INP(n8662), .Z(n8550) );
  NBUFFX2 U8480 ( .INP(n8645), .Z(n8638) );
  NBUFFX2 U8481 ( .INP(n8661), .Z(n8554) );
  NBUFFX2 U8482 ( .INP(n8657), .Z(n8575) );
  NBUFFX2 U8483 ( .INP(n8657), .Z(n8577) );
  NBUFFX2 U8484 ( .INP(n8646), .Z(n8630) );
  NBUFFX2 U8485 ( .INP(n8651), .Z(n8606) );
  NBUFFX2 U8486 ( .INP(n8664), .Z(n8543) );
  NBUFFX2 U8487 ( .INP(n8659), .Z(n8566) );
  NBUFFX2 U8488 ( .INP(n8647), .Z(n8625) );
  NBUFFX2 U8489 ( .INP(n8656), .Z(n8581) );
  NBUFFX2 U8490 ( .INP(n8648), .Z(n8621) );
  NBUFFX2 U8491 ( .INP(n8664), .Z(n8539) );
  NBUFFX2 U8492 ( .INP(n8658), .Z(n8572) );
  NBUFFX2 U8493 ( .INP(n8660), .Z(n8563) );
  NBUFFX2 U8494 ( .INP(n8648), .Z(n8620) );
  NBUFFX2 U8495 ( .INP(n8653), .Z(n8598) );
  NBUFFX2 U8496 ( .INP(n8658), .Z(n8573) );
  NBUFFX2 U8497 ( .INP(n8654), .Z(n8590) );
  NBUFFX2 U8498 ( .INP(n8655), .Z(n8586) );
  NBUFFX2 U8499 ( .INP(n8652), .Z(n8600) );
  NBUFFX2 U8500 ( .INP(n8649), .Z(n8615) );
  NBUFFX2 U8501 ( .INP(n8659), .Z(n8564) );
  NBUFFX2 U8502 ( .INP(n8653), .Z(n8597) );
  NBUFFX2 U8503 ( .INP(n8651), .Z(n8604) );
  NBUFFX2 U8504 ( .INP(n8661), .Z(n8557) );
  NBUFFX2 U8505 ( .INP(n8657), .Z(n8576) );
  NBUFFX2 U8506 ( .INP(n8645), .Z(n8637) );
  NBUFFX2 U8507 ( .INP(n8650), .Z(n8609) );
  NBUFFX2 U8508 ( .INP(n8645), .Z(n8636) );
  NBUFFX2 U8509 ( .INP(n8659), .Z(n8567) );
  NBUFFX2 U8510 ( .INP(n8661), .Z(n8558) );
  NBUFFX2 U8511 ( .INP(n8649), .Z(n8617) );
  NBUFFX2 U8512 ( .INP(n8649), .Z(n8614) );
  NBUFFX2 U8513 ( .INP(n8661), .Z(n8555) );
  NBUFFX2 U8514 ( .INP(n8645), .Z(n8635) );
  NBUFFX2 U8515 ( .INP(n8653), .Z(n8596) );
  NBUFFX2 U8516 ( .INP(n8648), .Z(n8619) );
  NBUFFX2 U8517 ( .INP(n8651), .Z(n8607) );
  NBUFFX2 U8518 ( .INP(n8652), .Z(n8599) );
  NBUFFX2 U8519 ( .INP(n8650), .Z(n8612) );
  NBUFFX2 U8520 ( .INP(n8657), .Z(n8574) );
  NBUFFX2 U8521 ( .INP(n8645), .Z(n8634) );
  NBUFFX2 U8522 ( .INP(n8648), .Z(n8622) );
  NBUFFX2 U8523 ( .INP(n8647), .Z(n8626) );
  NBUFFX2 U8524 ( .INP(n8661), .Z(n8556) );
  NBUFFX2 U8525 ( .INP(n8652), .Z(n8603) );
  NBUFFX2 U8526 ( .INP(n8659), .Z(n8568) );
  NBUFFX2 U8527 ( .INP(n8652), .Z(n8601) );
  NBUFFX2 U8528 ( .INP(n8664), .Z(n8542) );
  NBUFFX2 U8529 ( .INP(n8664), .Z(n8541) );
  NBUFFX2 U8530 ( .INP(n8662), .Z(n8552) );
  NBUFFX2 U8531 ( .INP(n8655), .Z(n8584) );
  NBUFFX2 U8532 ( .INP(n8662), .Z(n8553) );
  NBUFFX2 U8533 ( .INP(n8660), .Z(n8561) );
  NBUFFX2 U8534 ( .INP(n8650), .Z(n8611) );
  NBUFFX2 U8535 ( .INP(n8654), .Z(n8589) );
  NBUFFX2 U8536 ( .INP(n8663), .Z(n8546) );
  NBUFFX2 U8537 ( .INP(n8649), .Z(n8616) );
  NBUFFX2 U8538 ( .INP(n8658), .Z(n8569) );
  NBUFFX2 U8539 ( .INP(n8660), .Z(n8560) );
  NBUFFX2 U8540 ( .INP(n8654), .Z(n8592) );
  NBUFFX2 U8541 ( .INP(n8662), .Z(n8549) );
  NBUFFX2 U8542 ( .INP(n8648), .Z(n8623) );
  NBUFFX2 U8543 ( .INP(n8663), .Z(n8548) );
  NBUFFX2 U8544 ( .INP(n8664), .Z(n8540) );
  NBUFFX2 U8545 ( .INP(n8649), .Z(n8618) );
  NBUFFX2 U8546 ( .INP(n8663), .Z(n8544) );
  NBUFFX2 U8547 ( .INP(n8654), .Z(n8591) );
  NBUFFX2 U8548 ( .INP(n8660), .Z(n8559) );
  NBUFFX2 U8549 ( .INP(n8651), .Z(n8605) );
  NBUFFX2 U8550 ( .INP(n8652), .Z(n8602) );
  NBUFFX2 U8551 ( .INP(n8663), .Z(n8545) );
  NBUFFX2 U8552 ( .INP(n8646), .Z(n8631) );
  NBUFFX2 U8553 ( .INP(n8663), .Z(n8547) );
  NBUFFX2 U8554 ( .INP(n8657), .Z(n8578) );
  NBUFFX2 U8555 ( .INP(n8660), .Z(n8562) );
  NBUFFX2 U8556 ( .INP(n8658), .Z(n8570) );
  NBUFFX2 U8557 ( .INP(n8655), .Z(n8588) );
  NBUFFX2 U8558 ( .INP(n8656), .Z(n8579) );
  NBUFFX2 U8559 ( .INP(n8651), .Z(n8608) );
  NBUFFX2 U8560 ( .INP(n8647), .Z(n8627) );
  NBUFFX2 U8561 ( .INP(n8654), .Z(n8593) );
  NBUFFX2 U8562 ( .INP(n8650), .Z(n8610) );
  NBUFFX2 U8563 ( .INP(n8647), .Z(n8628) );
  NBUFFX2 U8564 ( .INP(n8658), .Z(n8571) );
  NBUFFX2 U8565 ( .INP(n8656), .Z(n8580) );
  NBUFFX2 U8566 ( .INP(n8659), .Z(n8565) );
  NBUFFX2 U8567 ( .INP(n8653), .Z(n8595) );
  NBUFFX2 U8568 ( .INP(n8653), .Z(n8594) );
  NBUFFX2 U8569 ( .INP(n8646), .Z(n8633) );
  NBUFFX2 U8570 ( .INP(n8646), .Z(n8629) );
  NBUFFX2 U8571 ( .INP(n8656), .Z(n8582) );
  NBUFFX2 U8572 ( .INP(n8656), .Z(n8583) );
  NBUFFX2 U8573 ( .INP(n8970), .Z(n8843) );
  NBUFFX2 U8574 ( .INP(n8970), .Z(n8842) );
  NBUFFX2 U8575 ( .INP(n8960), .Z(n8892) );
  NBUFFX2 U8576 ( .INP(n8960), .Z(n8890) );
  NBUFFX2 U8577 ( .INP(n8951), .Z(n8937) );
  NBUFFX2 U8578 ( .INP(n8967), .Z(n8856) );
  NBUFFX2 U8579 ( .INP(n8955), .Z(n8918) );
  NBUFFX2 U8580 ( .INP(n8952), .Z(n8929) );
  NBUFFX2 U8581 ( .INP(n8967), .Z(n8855) );
  NBUFFX2 U8582 ( .INP(n8950), .Z(n8943) );
  NBUFFX2 U8583 ( .INP(n8966), .Z(n8859) );
  NBUFFX2 U8584 ( .INP(n8962), .Z(n8880) );
  NBUFFX2 U8585 ( .INP(n8962), .Z(n8882) );
  NBUFFX2 U8586 ( .INP(n8951), .Z(n8935) );
  NBUFFX2 U8587 ( .INP(n8956), .Z(n8911) );
  NBUFFX2 U8588 ( .INP(n8969), .Z(n8848) );
  NBUFFX2 U8589 ( .INP(n8964), .Z(n8871) );
  NBUFFX2 U8590 ( .INP(n8952), .Z(n8930) );
  NBUFFX2 U8591 ( .INP(n8961), .Z(n8886) );
  NBUFFX2 U8592 ( .INP(n8953), .Z(n8926) );
  NBUFFX2 U8593 ( .INP(n8969), .Z(n8844) );
  NBUFFX2 U8594 ( .INP(n8963), .Z(n8877) );
  NBUFFX2 U8595 ( .INP(n8965), .Z(n8868) );
  NBUFFX2 U8596 ( .INP(n8953), .Z(n8925) );
  NBUFFX2 U8597 ( .INP(n8958), .Z(n8903) );
  NBUFFX2 U8598 ( .INP(n8963), .Z(n8878) );
  NBUFFX2 U8599 ( .INP(n8959), .Z(n8895) );
  NBUFFX2 U8600 ( .INP(n8960), .Z(n8891) );
  NBUFFX2 U8601 ( .INP(n8957), .Z(n8905) );
  NBUFFX2 U8602 ( .INP(n8954), .Z(n8920) );
  NBUFFX2 U8603 ( .INP(n8964), .Z(n8869) );
  NBUFFX2 U8604 ( .INP(n8958), .Z(n8902) );
  NBUFFX2 U8605 ( .INP(n8956), .Z(n8909) );
  NBUFFX2 U8606 ( .INP(n8966), .Z(n8862) );
  NBUFFX2 U8607 ( .INP(n8962), .Z(n8881) );
  NBUFFX2 U8608 ( .INP(n8950), .Z(n8942) );
  NBUFFX2 U8609 ( .INP(n8955), .Z(n8914) );
  NBUFFX2 U8610 ( .INP(n8950), .Z(n8941) );
  NBUFFX2 U8611 ( .INP(n8964), .Z(n8872) );
  NBUFFX2 U8612 ( .INP(n8966), .Z(n8863) );
  NBUFFX2 U8613 ( .INP(n8954), .Z(n8922) );
  NBUFFX2 U8614 ( .INP(n8954), .Z(n8919) );
  NBUFFX2 U8615 ( .INP(n8966), .Z(n8860) );
  NBUFFX2 U8616 ( .INP(n8950), .Z(n8940) );
  NBUFFX2 U8617 ( .INP(n8958), .Z(n8901) );
  NBUFFX2 U8618 ( .INP(n8953), .Z(n8924) );
  NBUFFX2 U8619 ( .INP(n8956), .Z(n8912) );
  NBUFFX2 U8620 ( .INP(n8957), .Z(n8904) );
  NBUFFX2 U8621 ( .INP(n8955), .Z(n8917) );
  NBUFFX2 U8622 ( .INP(n8962), .Z(n8879) );
  NBUFFX2 U8623 ( .INP(n8950), .Z(n8939) );
  NBUFFX2 U8624 ( .INP(n8953), .Z(n8927) );
  NBUFFX2 U8625 ( .INP(n8952), .Z(n8931) );
  NBUFFX2 U8626 ( .INP(n8966), .Z(n8861) );
  NBUFFX2 U8627 ( .INP(n8957), .Z(n8908) );
  NBUFFX2 U8628 ( .INP(n8964), .Z(n8873) );
  NBUFFX2 U8629 ( .INP(n8957), .Z(n8906) );
  NBUFFX2 U8630 ( .INP(n8969), .Z(n8847) );
  NBUFFX2 U8631 ( .INP(n8969), .Z(n8846) );
  NBUFFX2 U8632 ( .INP(n8967), .Z(n8857) );
  NBUFFX2 U8633 ( .INP(n8960), .Z(n8889) );
  NBUFFX2 U8634 ( .INP(n8967), .Z(n8858) );
  NBUFFX2 U8635 ( .INP(n8965), .Z(n8866) );
  NBUFFX2 U8636 ( .INP(n8955), .Z(n8916) );
  NBUFFX2 U8637 ( .INP(n8959), .Z(n8894) );
  NBUFFX2 U8638 ( .INP(n8968), .Z(n8851) );
  NBUFFX2 U8639 ( .INP(n8954), .Z(n8921) );
  NBUFFX2 U8640 ( .INP(n8963), .Z(n8874) );
  NBUFFX2 U8641 ( .INP(n8965), .Z(n8865) );
  NBUFFX2 U8642 ( .INP(n8959), .Z(n8897) );
  NBUFFX2 U8643 ( .INP(n8967), .Z(n8854) );
  NBUFFX2 U8644 ( .INP(n8953), .Z(n8928) );
  NBUFFX2 U8645 ( .INP(n8968), .Z(n8853) );
  NBUFFX2 U8646 ( .INP(n8969), .Z(n8845) );
  NBUFFX2 U8647 ( .INP(n8954), .Z(n8923) );
  NBUFFX2 U8648 ( .INP(n8968), .Z(n8849) );
  NBUFFX2 U8649 ( .INP(n8959), .Z(n8896) );
  NBUFFX2 U8650 ( .INP(n8965), .Z(n8864) );
  NBUFFX2 U8651 ( .INP(n8956), .Z(n8910) );
  NBUFFX2 U8652 ( .INP(n8957), .Z(n8907) );
  NBUFFX2 U8653 ( .INP(n8968), .Z(n8850) );
  NBUFFX2 U8654 ( .INP(n8951), .Z(n8936) );
  NBUFFX2 U8655 ( .INP(n8968), .Z(n8852) );
  NBUFFX2 U8656 ( .INP(n8962), .Z(n8883) );
  NBUFFX2 U8657 ( .INP(n8965), .Z(n8867) );
  NBUFFX2 U8658 ( .INP(n8963), .Z(n8875) );
  NBUFFX2 U8659 ( .INP(n8960), .Z(n8893) );
  NBUFFX2 U8660 ( .INP(n8961), .Z(n8884) );
  NBUFFX2 U8661 ( .INP(n8956), .Z(n8913) );
  NBUFFX2 U8662 ( .INP(n8952), .Z(n8932) );
  NBUFFX2 U8663 ( .INP(n8959), .Z(n8898) );
  NBUFFX2 U8664 ( .INP(n8955), .Z(n8915) );
  NBUFFX2 U8665 ( .INP(n8952), .Z(n8933) );
  NBUFFX2 U8666 ( .INP(n8963), .Z(n8876) );
  NBUFFX2 U8667 ( .INP(n8961), .Z(n8885) );
  NBUFFX2 U8668 ( .INP(n8964), .Z(n8870) );
  NBUFFX2 U8669 ( .INP(n8958), .Z(n8900) );
  NBUFFX2 U8670 ( .INP(n8958), .Z(n8899) );
  NBUFFX2 U8671 ( .INP(n8951), .Z(n8938) );
  NBUFFX2 U8672 ( .INP(n8951), .Z(n8934) );
  NBUFFX2 U8673 ( .INP(n8961), .Z(n8887) );
  NBUFFX2 U8674 ( .INP(n8961), .Z(n8888) );
  NBUFFX2 U8675 ( .INP(n8644), .Z(n8642) );
  NBUFFX2 U8676 ( .INP(n8644), .Z(n8640) );
  NBUFFX2 U8677 ( .INP(n8644), .Z(n8641) );
  NBUFFX2 U8678 ( .INP(n8644), .Z(n8639) );
  NBUFFX2 U8679 ( .INP(n8949), .Z(n8947) );
  NBUFFX2 U8680 ( .INP(n8949), .Z(n8945) );
  NBUFFX2 U8681 ( .INP(n8949), .Z(n8946) );
  NBUFFX2 U8682 ( .INP(n8949), .Z(n8944) );
  NBUFFX2 U8683 ( .INP(n8644), .Z(n8643) );
  NBUFFX2 U8684 ( .INP(n8949), .Z(n8948) );
  NBUFFX2 U8685 ( .INP(n8673), .Z(n8644) );
  NBUFFX2 U8686 ( .INP(n8672), .Z(n8645) );
  NBUFFX2 U8687 ( .INP(n8672), .Z(n8646) );
  NBUFFX2 U8688 ( .INP(n8672), .Z(n8647) );
  NBUFFX2 U8689 ( .INP(n8671), .Z(n8648) );
  NBUFFX2 U8690 ( .INP(n8671), .Z(n8649) );
  NBUFFX2 U8691 ( .INP(n8671), .Z(n8650) );
  NBUFFX2 U8692 ( .INP(n8670), .Z(n8651) );
  NBUFFX2 U8693 ( .INP(n8670), .Z(n8652) );
  NBUFFX2 U8694 ( .INP(n8670), .Z(n8653) );
  NBUFFX2 U8695 ( .INP(n8669), .Z(n8654) );
  NBUFFX2 U8696 ( .INP(n8669), .Z(n8655) );
  NBUFFX2 U8697 ( .INP(n8669), .Z(n8656) );
  NBUFFX2 U8698 ( .INP(n8668), .Z(n8657) );
  NBUFFX2 U8699 ( .INP(n8668), .Z(n8658) );
  NBUFFX2 U8700 ( .INP(n8668), .Z(n8659) );
  NBUFFX2 U8701 ( .INP(n8667), .Z(n8660) );
  NBUFFX2 U8702 ( .INP(n8667), .Z(n8661) );
  NBUFFX2 U8703 ( .INP(n8667), .Z(n8662) );
  NBUFFX2 U8704 ( .INP(n8666), .Z(n8663) );
  NBUFFX2 U8705 ( .INP(n8666), .Z(n8664) );
  NBUFFX2 U8706 ( .INP(n8666), .Z(n8665) );
  NBUFFX2 U8707 ( .INP(n8676), .Z(n8666) );
  NBUFFX2 U8708 ( .INP(n8676), .Z(n8667) );
  NBUFFX2 U8709 ( .INP(n8675), .Z(n8668) );
  NBUFFX2 U8710 ( .INP(n8675), .Z(n8669) );
  NBUFFX2 U8711 ( .INP(n8675), .Z(n8670) );
  NBUFFX2 U8712 ( .INP(n8674), .Z(n8671) );
  NBUFFX2 U8713 ( .INP(n8674), .Z(n8672) );
  NBUFFX2 U8714 ( .INP(n8674), .Z(n8673) );
  NBUFFX2 U8715 ( .INP(test_se), .Z(n8674) );
  NBUFFX2 U8716 ( .INP(test_se), .Z(n8675) );
  NBUFFX2 U8717 ( .INP(test_se), .Z(n8676) );
  NBUFFX2 U8718 ( .INP(n8779), .Z(n8677) );
  NBUFFX2 U8719 ( .INP(n8779), .Z(n8678) );
  NBUFFX2 U8720 ( .INP(n8778), .Z(n8679) );
  NBUFFX2 U8721 ( .INP(n8778), .Z(n8680) );
  NBUFFX2 U8722 ( .INP(n8778), .Z(n8681) );
  NBUFFX2 U8723 ( .INP(n8777), .Z(n8682) );
  NBUFFX2 U8724 ( .INP(n8777), .Z(n8683) );
  NBUFFX2 U8725 ( .INP(n8777), .Z(n8684) );
  NBUFFX2 U8726 ( .INP(n8776), .Z(n8685) );
  NBUFFX2 U8727 ( .INP(n8776), .Z(n8686) );
  NBUFFX2 U8728 ( .INP(n8776), .Z(n8687) );
  NBUFFX2 U8729 ( .INP(n8775), .Z(n8688) );
  NBUFFX2 U8730 ( .INP(n8775), .Z(n8689) );
  NBUFFX2 U8731 ( .INP(n8775), .Z(n8690) );
  NBUFFX2 U8732 ( .INP(n8774), .Z(n8691) );
  NBUFFX2 U8733 ( .INP(n8774), .Z(n8692) );
  NBUFFX2 U8734 ( .INP(n8774), .Z(n8693) );
  NBUFFX2 U8735 ( .INP(n8773), .Z(n8694) );
  NBUFFX2 U8736 ( .INP(n8773), .Z(n8695) );
  NBUFFX2 U8737 ( .INP(n8773), .Z(n8696) );
  NBUFFX2 U8738 ( .INP(n8772), .Z(n8697) );
  NBUFFX2 U8739 ( .INP(n8772), .Z(n8698) );
  NBUFFX2 U8740 ( .INP(n8772), .Z(n8699) );
  NBUFFX2 U8741 ( .INP(n8771), .Z(n8700) );
  NBUFFX2 U8742 ( .INP(n8771), .Z(n8701) );
  NBUFFX2 U8743 ( .INP(n8771), .Z(n8702) );
  NBUFFX2 U8744 ( .INP(n8770), .Z(n8703) );
  NBUFFX2 U8745 ( .INP(n8770), .Z(n8704) );
  NBUFFX2 U8746 ( .INP(n8770), .Z(n8705) );
  NBUFFX2 U8747 ( .INP(n8769), .Z(n8706) );
  NBUFFX2 U8748 ( .INP(n8769), .Z(n8707) );
  NBUFFX2 U8749 ( .INP(n8769), .Z(n8708) );
  NBUFFX2 U8750 ( .INP(n8768), .Z(n8709) );
  NBUFFX2 U8751 ( .INP(n8768), .Z(n8710) );
  NBUFFX2 U8752 ( .INP(n8768), .Z(n8711) );
  NBUFFX2 U8753 ( .INP(n8767), .Z(n8712) );
  NBUFFX2 U8754 ( .INP(n8767), .Z(n8713) );
  NBUFFX2 U8755 ( .INP(n8767), .Z(n8714) );
  NBUFFX2 U8756 ( .INP(n8766), .Z(n8715) );
  NBUFFX2 U8757 ( .INP(n8766), .Z(n8716) );
  NBUFFX2 U8758 ( .INP(n8766), .Z(n8717) );
  NBUFFX2 U8759 ( .INP(n8765), .Z(n8718) );
  NBUFFX2 U8760 ( .INP(n8765), .Z(n8719) );
  NBUFFX2 U8761 ( .INP(n8765), .Z(n8720) );
  NBUFFX2 U8762 ( .INP(n8764), .Z(n8721) );
  NBUFFX2 U8763 ( .INP(n8764), .Z(n8722) );
  NBUFFX2 U8764 ( .INP(n8764), .Z(n8723) );
  NBUFFX2 U8765 ( .INP(n8763), .Z(n8724) );
  NBUFFX2 U8766 ( .INP(n8763), .Z(n8725) );
  NBUFFX2 U8767 ( .INP(n8763), .Z(n8726) );
  NBUFFX2 U8768 ( .INP(n8762), .Z(n8727) );
  NBUFFX2 U8769 ( .INP(n8762), .Z(n8728) );
  NBUFFX2 U8770 ( .INP(n8762), .Z(n8729) );
  NBUFFX2 U8771 ( .INP(n8761), .Z(n8730) );
  NBUFFX2 U8772 ( .INP(n8761), .Z(n8731) );
  NBUFFX2 U8773 ( .INP(n8761), .Z(n8732) );
  NBUFFX2 U8774 ( .INP(n8760), .Z(n8733) );
  NBUFFX2 U8775 ( .INP(n8760), .Z(n8734) );
  NBUFFX2 U8776 ( .INP(n8760), .Z(n8735) );
  NBUFFX2 U8777 ( .INP(n8759), .Z(n8736) );
  NBUFFX2 U8778 ( .INP(n8759), .Z(n8737) );
  NBUFFX2 U8779 ( .INP(n8759), .Z(n8738) );
  NBUFFX2 U8780 ( .INP(n8758), .Z(n8739) );
  NBUFFX2 U8781 ( .INP(n8758), .Z(n8740) );
  NBUFFX2 U8782 ( .INP(n8758), .Z(n8741) );
  NBUFFX2 U8783 ( .INP(n8757), .Z(n8742) );
  NBUFFX2 U8784 ( .INP(n8757), .Z(n8743) );
  NBUFFX2 U8785 ( .INP(n8757), .Z(n8744) );
  NBUFFX2 U8786 ( .INP(n8756), .Z(n8745) );
  NBUFFX2 U8787 ( .INP(n8756), .Z(n8746) );
  NBUFFX2 U8788 ( .INP(n8756), .Z(n8747) );
  NBUFFX2 U8789 ( .INP(n8755), .Z(n8748) );
  NBUFFX2 U8790 ( .INP(n8755), .Z(n8749) );
  NBUFFX2 U8791 ( .INP(n8755), .Z(n8750) );
  NBUFFX2 U8792 ( .INP(n8754), .Z(n8751) );
  NBUFFX2 U8793 ( .INP(n8754), .Z(n8752) );
  NBUFFX2 U8794 ( .INP(n8754), .Z(n8753) );
  NBUFFX2 U8795 ( .INP(n8788), .Z(n8754) );
  NBUFFX2 U8796 ( .INP(n8788), .Z(n8755) );
  NBUFFX2 U8797 ( .INP(n8787), .Z(n8756) );
  NBUFFX2 U8798 ( .INP(n8787), .Z(n8757) );
  NBUFFX2 U8799 ( .INP(n8787), .Z(n8758) );
  NBUFFX2 U8800 ( .INP(n8786), .Z(n8759) );
  NBUFFX2 U8801 ( .INP(n8786), .Z(n8760) );
  NBUFFX2 U8802 ( .INP(n8786), .Z(n8761) );
  NBUFFX2 U8803 ( .INP(n8785), .Z(n8762) );
  NBUFFX2 U8804 ( .INP(n8785), .Z(n8763) );
  NBUFFX2 U8805 ( .INP(n8785), .Z(n8764) );
  NBUFFX2 U8806 ( .INP(n8784), .Z(n8765) );
  NBUFFX2 U8807 ( .INP(n8784), .Z(n8766) );
  NBUFFX2 U8808 ( .INP(n8784), .Z(n8767) );
  NBUFFX2 U8809 ( .INP(n8783), .Z(n8768) );
  NBUFFX2 U8810 ( .INP(n8783), .Z(n8769) );
  NBUFFX2 U8811 ( .INP(n8783), .Z(n8770) );
  NBUFFX2 U8812 ( .INP(n8782), .Z(n8771) );
  NBUFFX2 U8813 ( .INP(n8782), .Z(n8772) );
  NBUFFX2 U8814 ( .INP(n8782), .Z(n8773) );
  NBUFFX2 U8815 ( .INP(n8781), .Z(n8774) );
  NBUFFX2 U8816 ( .INP(n8781), .Z(n8775) );
  NBUFFX2 U8817 ( .INP(n8781), .Z(n8776) );
  NBUFFX2 U8818 ( .INP(n8780), .Z(n8777) );
  NBUFFX2 U8819 ( .INP(n8780), .Z(n8778) );
  NBUFFX2 U8820 ( .INP(n8780), .Z(n8779) );
  NBUFFX2 U8821 ( .INP(n8791), .Z(n8780) );
  NBUFFX2 U8822 ( .INP(n8791), .Z(n8781) );
  NBUFFX2 U8823 ( .INP(n8791), .Z(n8782) );
  NBUFFX2 U8824 ( .INP(n8790), .Z(n8783) );
  NBUFFX2 U8825 ( .INP(n8790), .Z(n8784) );
  NBUFFX2 U8826 ( .INP(n8790), .Z(n8785) );
  NBUFFX2 U8827 ( .INP(n8789), .Z(n8786) );
  NBUFFX2 U8828 ( .INP(n8789), .Z(n8787) );
  NBUFFX2 U8829 ( .INP(n8789), .Z(n8788) );
  NBUFFX2 U8830 ( .INP(g35), .Z(n8789) );
  NBUFFX2 U8831 ( .INP(g35), .Z(n8790) );
  NBUFFX2 U8832 ( .INP(g35), .Z(n8791) );
  INVX0 U8833 ( .INP(n8684), .ZN(n8792) );
  INVX0 U8834 ( .INP(n8683), .ZN(n8793) );
  INVX0 U8835 ( .INP(n8685), .ZN(n8794) );
  INVX0 U8836 ( .INP(n8684), .ZN(n8795) );
  INVX0 U8837 ( .INP(n8685), .ZN(n8796) );
  INVX0 U8838 ( .INP(n8685), .ZN(n8797) );
  INVX0 U8839 ( .INP(n8684), .ZN(n8798) );
  INVX0 U8840 ( .INP(n8683), .ZN(n8799) );
  INVX0 U8841 ( .INP(n8684), .ZN(n8800) );
  INVX0 U8842 ( .INP(n8684), .ZN(n8801) );
  INVX0 U8843 ( .INP(n8680), .ZN(n8802) );
  INVX0 U8844 ( .INP(n8684), .ZN(n8803) );
  INVX0 U8845 ( .INP(n8684), .ZN(n8804) );
  INVX0 U8846 ( .INP(n8684), .ZN(n8805) );
  INVX0 U8847 ( .INP(n8684), .ZN(n8806) );
  INVX0 U8848 ( .INP(n8683), .ZN(n8807) );
  INVX0 U8849 ( .INP(n8683), .ZN(n8808) );
  INVX0 U8850 ( .INP(n8683), .ZN(n8809) );
  INVX0 U8851 ( .INP(n8683), .ZN(n8810) );
  INVX0 U8852 ( .INP(n8683), .ZN(n8811) );
  INVX0 U8853 ( .INP(n8682), .ZN(n8812) );
  INVX0 U8854 ( .INP(n8683), .ZN(n8813) );
  INVX0 U8855 ( .INP(n8682), .ZN(n8814) );
  INVX0 U8856 ( .INP(n8682), .ZN(n8815) );
  INVX0 U8857 ( .INP(n8681), .ZN(n8816) );
  INVX0 U8858 ( .INP(n8682), .ZN(n8817) );
  INVX0 U8859 ( .INP(n8683), .ZN(n8818) );
  INVX0 U8860 ( .INP(n8682), .ZN(n8819) );
  INVX0 U8861 ( .INP(n8681), .ZN(n8820) );
  INVX0 U8862 ( .INP(n8682), .ZN(n8821) );
  INVX0 U8863 ( .INP(n8682), .ZN(n8822) );
  INVX0 U8864 ( .INP(n8682), .ZN(n8823) );
  INVX0 U8865 ( .INP(n8681), .ZN(n8824) );
  INVX0 U8866 ( .INP(n8681), .ZN(n8825) );
  INVX0 U8867 ( .INP(n8681), .ZN(n8826) );
  INVX0 U8868 ( .INP(n8681), .ZN(n8827) );
  INVX0 U8869 ( .INP(n8681), .ZN(n8828) );
  INVX0 U8870 ( .INP(n8680), .ZN(n8829) );
  INVX0 U8871 ( .INP(n8680), .ZN(n8830) );
  INVX0 U8872 ( .INP(n8680), .ZN(n8831) );
  INVX0 U8873 ( .INP(n8681), .ZN(n8832) );
  INVX0 U8874 ( .INP(n8680), .ZN(n8833) );
  INVX0 U8875 ( .INP(n8678), .ZN(n8834) );
  INVX0 U8876 ( .INP(n8680), .ZN(n8835) );
  INVX0 U8877 ( .INP(n8680), .ZN(n8836) );
  INVX0 U8878 ( .INP(n8680), .ZN(n8837) );
  INVX0 U8879 ( .INP(n8681), .ZN(n8838) );
  INVX0 U8880 ( .INP(n8682), .ZN(n8839) );
  INVX0 U8881 ( .INP(n8680), .ZN(n8840) );
  INVX0 U8882 ( .INP(n8679), .ZN(n8841) );
  NBUFFX2 U8883 ( .INP(n8978), .Z(n8949) );
  NBUFFX2 U8884 ( .INP(n8977), .Z(n8950) );
  NBUFFX2 U8885 ( .INP(n8977), .Z(n8951) );
  NBUFFX2 U8886 ( .INP(n8977), .Z(n8952) );
  NBUFFX2 U8887 ( .INP(n8976), .Z(n8953) );
  NBUFFX2 U8888 ( .INP(n8976), .Z(n8954) );
  NBUFFX2 U8889 ( .INP(n8976), .Z(n8955) );
  NBUFFX2 U8890 ( .INP(n8975), .Z(n8956) );
  NBUFFX2 U8891 ( .INP(n8975), .Z(n8957) );
  NBUFFX2 U8892 ( .INP(n8975), .Z(n8958) );
  NBUFFX2 U8893 ( .INP(n8974), .Z(n8959) );
  NBUFFX2 U8894 ( .INP(n8974), .Z(n8960) );
  NBUFFX2 U8895 ( .INP(n8974), .Z(n8961) );
  NBUFFX2 U8896 ( .INP(n8973), .Z(n8962) );
  NBUFFX2 U8897 ( .INP(n8973), .Z(n8963) );
  NBUFFX2 U8898 ( .INP(n8973), .Z(n8964) );
  NBUFFX2 U8899 ( .INP(n8972), .Z(n8965) );
  NBUFFX2 U8900 ( .INP(n8972), .Z(n8966) );
  NBUFFX2 U8901 ( .INP(n8972), .Z(n8967) );
  NBUFFX2 U8902 ( .INP(n8971), .Z(n8968) );
  NBUFFX2 U8903 ( .INP(n8971), .Z(n8969) );
  NBUFFX2 U8904 ( .INP(n8971), .Z(n8970) );
  NBUFFX2 U8905 ( .INP(n8981), .Z(n8971) );
  NBUFFX2 U8906 ( .INP(n8981), .Z(n8972) );
  NBUFFX2 U8907 ( .INP(n8980), .Z(n8973) );
  NBUFFX2 U8908 ( .INP(n8980), .Z(n8974) );
  NBUFFX2 U8909 ( .INP(n8980), .Z(n8975) );
  NBUFFX2 U8910 ( .INP(n8979), .Z(n8976) );
  NBUFFX2 U8911 ( .INP(n8979), .Z(n8977) );
  NBUFFX2 U8912 ( .INP(n8979), .Z(n8978) );
  NBUFFX2 U8913 ( .INP(CK), .Z(n8979) );
  NBUFFX2 U8914 ( .INP(CK), .Z(n8980) );
  NBUFFX2 U8915 ( .INP(CK), .Z(n8981) );
  INVX0 U8916 ( .INP(n8982), .ZN(n967) );
  INVX0 U8917 ( .INP(n8983), .ZN(n872) );
  AND3X1 U8918 ( .IN1(n8984), .IN2(n8985), .IN3(n8986), .Q(n8472) );
  INVX0 U8919 ( .INP(n8987), .ZN(n797) );
  INVX0 U8920 ( .INP(n8988), .ZN(n730) );
  INVX0 U8921 ( .INP(n8989), .ZN(n728) );
  INVX0 U8922 ( .INP(n8990), .ZN(n725) );
  OR4X1 U8923 ( .IN1(n8991), .IN2(n8992), .IN3(n8993), .IN4(n8994), .Q(n5961)
         );
  AND2X1 U8924 ( .IN1(n8180), .IN2(n8995), .Q(n8994) );
  AND2X1 U8925 ( .IN1(n8996), .IN2(g5348), .Q(n8993) );
  AND2X1 U8926 ( .IN1(n8444), .IN2(n8997), .Q(n8992) );
  AND2X1 U8927 ( .IN1(g31860), .IN2(g5352), .Q(n8991) );
  OR4X1 U8928 ( .IN1(n8998), .IN2(n8999), .IN3(n9000), .IN4(n9001), .Q(n5960)
         );
  AND2X1 U8929 ( .IN1(n8423), .IN2(n9002), .Q(n9001) );
  AND2X1 U8930 ( .IN1(n9003), .IN2(g6736), .Q(n9000) );
  AND2X1 U8931 ( .IN1(n8179), .IN2(n9004), .Q(n8999) );
  AND2X1 U8932 ( .IN1(n9005), .IN2(g6732), .Q(n8998) );
  INVX0 U8933 ( .INP(n9006), .ZN(n525) );
  INVX0 U8934 ( .INP(n9007), .ZN(n524) );
  OR3X1 U8935 ( .IN1(n9008), .IN2(n9009), .IN3(n9010), .Q(n514) );
  AND2X1 U8936 ( .IN1(n9011), .IN2(g3845), .Q(n9010) );
  AND4X1 U8937 ( .IN1(n9012), .IN2(n8752), .IN3(n5662), .IN4(n8528), .Q(n9009)
         );
  AND2X1 U8938 ( .IN1(test_so97), .IN2(n9013), .Q(n9008) );
  OR2X1 U8939 ( .IN1(n8801), .IN2(n9014), .Q(n9013) );
  AND2X1 U8940 ( .IN1(n9012), .IN2(g3835), .Q(n9014) );
  OR2X1 U8941 ( .IN1(n8299), .IN2(n9015), .Q(n4459) );
  OR2X1 U8942 ( .IN1(n8303), .IN2(n9016), .Q(n4448) );
  OR2X1 U8943 ( .IN1(n9017), .IN2(n8517), .Q(n4437) );
  OR2X1 U8944 ( .IN1(n8297), .IN2(n9018), .Q(n4426) );
  OR2X1 U8945 ( .IN1(n8305), .IN2(n9019), .Q(n4415) );
  OR2X1 U8946 ( .IN1(n8301), .IN2(n9020), .Q(n4403) );
  OR2X1 U8947 ( .IN1(n8294), .IN2(n9021), .Q(n4392) );
  OR2X1 U8948 ( .IN1(n8292), .IN2(n9022), .Q(n4380) );
  OR4X1 U8949 ( .IN1(n9023), .IN2(n9024), .IN3(n9025), .IN4(n9026), .Q(n4305)
         );
  OR2X1 U8950 ( .IN1(n9027), .IN2(n9028), .Q(n9026) );
  AND2X1 U8951 ( .IN1(g4646), .IN2(g29220), .Q(n9028) );
  AND2X1 U8952 ( .IN1(n5880), .IN2(g4674), .Q(n9027) );
  AND2X1 U8953 ( .IN1(g4831), .IN2(g4681), .Q(n9025) );
  AND3X1 U8954 ( .IN1(n9029), .IN2(n9030), .IN3(n5656), .Q(n9024) );
  OR3X1 U8955 ( .IN1(n9031), .IN2(n9032), .IN3(n9033), .Q(n9030) );
  AND3X1 U8956 ( .IN1(n9034), .IN2(n9035), .IN3(n5707), .Q(n9033) );
  OR2X1 U8957 ( .IN1(n5368), .IN2(g34657), .Q(n9035) );
  OR2X1 U8958 ( .IN1(n9036), .IN2(g4793), .Q(n9034) );
  AND2X1 U8959 ( .IN1(n9037), .IN2(n8504), .Q(n9036) );
  OR3X1 U8960 ( .IN1(n9038), .IN2(n9039), .IN3(n9040), .Q(n9037) );
  AND2X1 U8961 ( .IN1(n9041), .IN2(n5867), .Q(n9040) );
  AND2X1 U8962 ( .IN1(n9042), .IN2(n9043), .Q(n9032) );
  XOR2X1 U8963 ( .IN1(g34657), .IN2(n9044), .Q(n9043) );
  OR4X1 U8964 ( .IN1(n9045), .IN2(n9046), .IN3(n9047), .IN4(n9048), .Q(n9044)
         );
  AND2X1 U8965 ( .IN1(n9041), .IN2(g4727), .Q(n9048) );
  AND3X1 U8966 ( .IN1(n5361), .IN2(g4722), .IN3(n5518), .Q(n9047) );
  AND2X1 U8967 ( .IN1(n9038), .IN2(g4717), .Q(n9046) );
  AND2X1 U8968 ( .IN1(n9039), .IN2(g4732), .Q(n9045) );
  AND2X1 U8969 ( .IN1(n8010), .IN2(g4688), .Q(n9023) );
  OR4X1 U8970 ( .IN1(n9049), .IN2(n9050), .IN3(n9051), .IN4(n9052), .Q(n4283)
         );
  OR2X1 U8971 ( .IN1(n9053), .IN2(n9054), .Q(n9052) );
  AND2X1 U8972 ( .IN1(g4871), .IN2(g3684), .Q(n9054) );
  AND2X1 U8973 ( .IN1(n8013), .IN2(g4864), .Q(n9053) );
  AND2X1 U8976 ( .IN1(g4836), .IN2(g5011), .Q(n9051) );
  AND3X1 U8977 ( .IN1(n9055), .IN2(n9056), .IN3(n5283), .Q(n9050) );
  OR3X1 U8978 ( .IN1(n9057), .IN2(n9058), .IN3(n9059), .Q(n9056) );
  AND3X1 U8979 ( .IN1(n9060), .IN2(n9061), .IN3(n5706), .Q(n9059) );
  OR2X1 U8980 ( .IN1(n5367), .IN2(g34649), .Q(n9061) );
  OR2X1 U8981 ( .IN1(n9062), .IN2(g4983), .Q(n9060) );
  AND2X1 U8982 ( .IN1(n9063), .IN2(n8505), .Q(n9062) );
  OR3X1 U8983 ( .IN1(n9064), .IN2(n9065), .IN3(n9066), .Q(n9063) );
  AND2X1 U8984 ( .IN1(n9067), .IN2(n5879), .Q(n9066) );
  AND2X1 U8985 ( .IN1(n9068), .IN2(n9069), .Q(n9058) );
  XOR2X1 U8986 ( .IN1(g34649), .IN2(n9070), .Q(n9069) );
  OR4X1 U8987 ( .IN1(n9071), .IN2(n9072), .IN3(n9073), .IN4(n9074), .Q(n9070)
         );
  AND2X1 U8988 ( .IN1(n9067), .IN2(g4917), .Q(n9074) );
  AND3X1 U8989 ( .IN1(n5360), .IN2(g4912), .IN3(n5517), .Q(n9073) );
  AND2X1 U8990 ( .IN1(n9064), .IN2(g4907), .Q(n9072) );
  AND2X1 U8991 ( .IN1(n9065), .IN2(g4922), .Q(n9071) );
  AND2X1 U8992 ( .IN1(n8014), .IN2(g4878), .Q(n9049) );
  AND3X1 U8993 ( .IN1(n5652), .IN2(n5366), .IN3(n8315), .Q(n4034) );
  AND3X1 U8994 ( .IN1(n5645), .IN2(n5576), .IN3(n8308), .Q(n4002) );
  AND3X1 U8995 ( .IN1(n5572), .IN2(n8493), .IN3(n8310), .Q(n3969) );
  AND4X1 U8996 ( .IN1(n8984), .IN2(n8985), .IN3(n2760), .IN4(g43), .Q(n3933)
         );
  AND3X1 U8997 ( .IN1(n5650), .IN2(n5570), .IN3(n8313), .Q(n3926) );
  AND3X1 U8998 ( .IN1(n5647), .IN2(n5575), .IN3(n8311), .Q(n3893) );
  AND3X1 U8999 ( .IN1(n5649), .IN2(n5573), .IN3(n8309), .Q(n3860) );
  AND3X1 U9000 ( .IN1(n5651), .IN2(n5574), .IN3(n8312), .Q(n3826) );
  AND3X1 U9001 ( .IN1(n5646), .IN2(n5571), .IN3(n8314), .Q(n3792) );
  OR4X1 U9002 ( .IN1(g691), .IN2(g417), .IN3(n9075), .IN4(n9076), .Q(n3675) );
  AND2X1 U9003 ( .IN1(n9077), .IN2(g392), .Q(n9076) );
  OR2X1 U9004 ( .IN1(g441), .IN2(n9078), .Q(n9077) );
  XNOR2X1 U9005 ( .IN1(test_so72), .IN2(g452), .Q(n9078) );
  AND2X1 U9006 ( .IN1(n8344), .IN2(n9079), .Q(n9075) );
  OR2X1 U9007 ( .IN1(g411), .IN2(n9080), .Q(n9079) );
  XOR2X1 U9008 ( .IN1(test_so72), .IN2(n5402), .Q(n9080) );
  OR2X1 U9009 ( .IN1(n5349), .IN2(n9081), .Q(n3635) );
  INVX0 U9010 ( .INP(n9082), .ZN(n357) );
  AND2X1 U9011 ( .IN1(n3064), .IN2(n9083), .Q(n9082) );
  OR2X1 U9012 ( .IN1(n5715), .IN2(n9084), .Q(n9083) );
  AND2X1 U9013 ( .IN1(n9085), .IN2(n8699), .Q(n9084) );
  OR2X1 U9014 ( .IN1(g4104), .IN2(n9086), .Q(n9085) );
  AND2X1 U9015 ( .IN1(n9087), .IN2(n9088), .Q(n3174) );
  XOR2X1 U9016 ( .IN1(n5708), .IN2(g73), .Q(n9088) );
  XOR2X1 U9017 ( .IN1(g72), .IN2(n5820), .Q(n9087) );
  INVX0 U9018 ( .INP(n9089), .ZN(n310) );
  AND2X1 U9019 ( .IN1(g34979), .IN2(n9090), .Q(n9089) );
  AND2X1 U9020 ( .IN1(n2760), .IN2(n9302), .Q(n3084) );
  OR3X1 U9021 ( .IN1(n8363), .IN2(n8792), .IN3(n9091), .Q(n3065) );
  AND2X1 U9022 ( .IN1(n9092), .IN2(g4108), .Q(n9091) );
  INVX0 U9023 ( .INP(n9093), .ZN(n301) );
  INVX0 U9024 ( .INP(n9094), .ZN(n297) );
  XOR2X1 U9025 ( .IN1(n5323), .IN2(n2607), .Q(n2608) );
  AND2X1 U9026 ( .IN1(n9090), .IN2(g34971), .Q(n2396) );
  INVX0 U9027 ( .INP(n9095), .ZN(n201) );
  OR3X1 U9028 ( .IN1(n9096), .IN2(n9097), .IN3(n9098), .Q(n191) );
  AND2X1 U9029 ( .IN1(n9099), .IN2(g5152), .Q(n9098) );
  AND4X1 U9030 ( .IN1(g32975), .IN2(n8752), .IN3(n5658), .IN4(n8529), .Q(n9097) );
  AND2X1 U9031 ( .IN1(test_so98), .IN2(n9100), .Q(n9096) );
  OR2X1 U9032 ( .IN1(n8801), .IN2(n9101), .Q(n9100) );
  AND2X1 U9033 ( .IN1(g32975), .IN2(g5142), .Q(n9101) );
  INVX0 U9034 ( .INP(n9102), .ZN(n184) );
  INVX0 U9035 ( .INP(n9103), .ZN(n181) );
  INVX0 U9036 ( .INP(n9104), .ZN(n180) );
  INVX0 U9037 ( .INP(n9105), .ZN(n175) );
  INVX0 U9038 ( .INP(n9106), .ZN(n1633) );
  INVX0 U9039 ( .INP(n9107), .ZN(n1574) );
  INVX0 U9040 ( .INP(n9108), .ZN(n1285) );
  INVX0 U9041 ( .INP(n9109), .ZN(n1283) );
  INVX0 U9042 ( .INP(n9110), .ZN(n1281) );
  INVX0 U9043 ( .INP(n9111), .ZN(n1279) );
  OR2X1 U9044 ( .IN1(n9112), .IN2(n9113), .Q(g34980) );
  AND2X1 U9045 ( .IN1(n9114), .IN2(n8699), .Q(n9113) );
  OR2X1 U9046 ( .IN1(n9115), .IN2(g2984), .Q(n9114) );
  AND4X1 U9047 ( .IN1(n8471), .IN2(n9116), .IN3(n9117), .IN4(n9118), .Q(n9115)
         );
  INVX0 U9048 ( .INP(g56), .ZN(n9118) );
  AND2X1 U9049 ( .IN1(test_so14), .IN2(n8808), .Q(n9112) );
  OR2X1 U9050 ( .IN1(n8459), .IN2(n8471), .Q(g34972) );
  XOR3X1 U9051 ( .IN1(g34975), .IN2(g34974), .IN3(n9119), .Q(n8471) );
  XNOR3X1 U9052 ( .IN1(n9120), .IN2(g34978), .IN3(n9121), .Q(n9119) );
  XOR3X1 U9053 ( .IN1(g34977), .IN2(g34976), .IN3(g34979), .Q(n9121) );
  XOR3X1 U9054 ( .IN1(n9122), .IN2(g34971), .IN3(g34970), .Q(n9120) );
  AND2X1 U9055 ( .IN1(n9123), .IN2(g55), .Q(n9122) );
  OR2X1 U9056 ( .IN1(n8459), .IN2(g34979), .Q(g34927) );
  OR4X1 U9057 ( .IN1(n9124), .IN2(n9125), .IN3(n9126), .IN4(n9127), .Q(g34979)
         );
  OR4X1 U9058 ( .IN1(n9128), .IN2(n9129), .IN3(n9130), .IN4(n9131), .Q(n9127)
         );
  AND2X1 U9059 ( .IN1(n9132), .IN2(n9332), .Q(n9131) );
  AND2X1 U9060 ( .IN1(n9133), .IN2(g1283), .Q(n9130) );
  AND2X1 U9061 ( .IN1(n9134), .IN2(g2138), .Q(n9129) );
  AND2X1 U9062 ( .IN1(n9135), .IN2(g2697), .Q(n9128) );
  OR2X1 U9063 ( .IN1(n9136), .IN2(n9137), .Q(n9126) );
  AND2X1 U9064 ( .IN1(test_so67), .IN2(n9138), .Q(n9137) );
  AND2X1 U9066 ( .IN1(n9139), .IN2(g4146), .Q(n9136) );
  AND2X1 U9067 ( .IN1(n9140), .IN2(g939), .Q(n9125) );
  AND2X1 U9068 ( .IN1(n1338), .IN2(n9141), .Q(n9124) );
  OR4X1 U9069 ( .IN1(n9142), .IN2(n9143), .IN3(n9144), .IN4(n9145), .Q(n9141)
         );
  OR4X1 U9071 ( .IN1(n9146), .IN2(n9147), .IN3(n9148), .IN4(n9149), .Q(n9145)
         );
  OR3X1 U9072 ( .IN1(n9150), .IN2(n9151), .IN3(n9152), .Q(n9149) );
  AND2X1 U9073 ( .IN1(test_so14), .IN2(n9090), .Q(n9152) );
  AND2X1 U9074 ( .IN1(g92), .IN2(n9153), .Q(n9151) );
  AND2X1 U9077 ( .IN1(g127), .IN2(n9154), .Q(n9150) );
  AND2X1 U9078 ( .IN1(n9155), .IN2(g744), .Q(n9148) );
  AND2X1 U9079 ( .IN1(n9156), .IN2(g2886), .Q(n9147) );
  AND2X1 U9081 ( .IN1(n9157), .IN2(g785), .Q(n9146) );
  OR3X1 U9082 ( .IN1(n9158), .IN2(n9159), .IN3(n9160), .Q(n9144) );
  AND2X1 U9083 ( .IN1(n9161), .IN2(g2975), .Q(n9160) );
  AND2X1 U9087 ( .IN1(n9162), .IN2(g2970), .Q(n9159) );
  AND2X1 U9088 ( .IN1(n9163), .IN2(g604), .Q(n9158) );
  OR2X1 U9089 ( .IN1(n9164), .IN2(n9165), .Q(n9143) );
  AND2X1 U9091 ( .IN1(n9166), .IN2(g568), .Q(n9165) );
  AND2X1 U9092 ( .IN1(g29221), .IN2(n9167), .Q(n9164) );
  OR2X1 U9093 ( .IN1(n8459), .IN2(g34978), .Q(g34925) );
  OR4X1 U9094 ( .IN1(n9168), .IN2(n9169), .IN3(n9170), .IN4(n9171), .Q(g34978)
         );
  OR4X1 U9095 ( .IN1(n9172), .IN2(n9173), .IN3(n9174), .IN4(n9175), .Q(n9171)
         );
  AND2X1 U9096 ( .IN1(n9132), .IN2(n9276), .Q(n9175) );
  AND2X1 U9097 ( .IN1(n7948), .IN2(n9133), .Q(n9174) );
  AND2X1 U9100 ( .IN1(n9134), .IN2(g2130), .Q(n9173) );
  AND2X1 U9102 ( .IN1(n9135), .IN2(g2689), .Q(n9172) );
  OR2X1 U9103 ( .IN1(n9176), .IN2(n9177), .Q(n9170) );
  AND2X1 U9104 ( .IN1(n9138), .IN2(g4253), .Q(n9177) );
  AND2X1 U9105 ( .IN1(n9139), .IN2(g4176), .Q(n9176) );
  AND2X1 U9106 ( .IN1(n7949), .IN2(n9140), .Q(n9169) );
  AND2X1 U9108 ( .IN1(n1338), .IN2(n9178), .Q(n9168) );
  OR4X1 U9109 ( .IN1(n9179), .IN2(n9142), .IN3(n9180), .IN4(n9181), .Q(n9178)
         );
  OR4X1 U9110 ( .IN1(n9182), .IN2(n9183), .IN3(n9184), .IN4(n9185), .Q(n9181)
         );
  OR3X1 U9112 ( .IN1(n9186), .IN2(n9187), .IN3(n9188), .Q(n9185) );
  AND2X1 U9113 ( .IN1(n9157), .IN2(g790), .Q(n9188) );
  AND2X1 U9114 ( .IN1(n9153), .IN2(g29214), .Q(n9187) );
  AND2X1 U9115 ( .IN1(n9154), .IN2(g2873), .Q(n9186) );
  AND2X1 U9117 ( .IN1(n9163), .IN2(g608), .Q(n9184) );
  AND2X1 U9118 ( .IN1(test_so2), .IN2(n9155), .Q(n9183) );
  AND2X1 U9119 ( .IN1(n9156), .IN2(g2878), .Q(n9182) );
  OR3X1 U9121 ( .IN1(n9189), .IN2(n9190), .IN3(n9191), .Q(n9180) );
  AND2X1 U9122 ( .IN1(n8208), .IN2(n9167), .Q(n9191) );
  AND2X1 U9123 ( .IN1(n9161), .IN2(g2965), .Q(n9190) );
  AND2X1 U9125 ( .IN1(test_so22), .IN2(n9162), .Q(n9189) );
  AND2X1 U9126 ( .IN1(n9166), .IN2(g572), .Q(n9179) );
  OR2X1 U9127 ( .IN1(n8459), .IN2(g34977), .Q(g34923) );
  OR4X1 U9129 ( .IN1(n9192), .IN2(n9193), .IN3(n9194), .IN4(n9195), .Q(g34977)
         );
  OR4X1 U9130 ( .IN1(n9196), .IN2(n9142), .IN3(n9197), .IN4(n9198), .Q(n9195)
         );
  AND2X1 U9131 ( .IN1(n5867), .IN2(n9199), .Q(n9198) );
  AND2X1 U9133 ( .IN1(n9132), .IN2(n9245), .Q(n9197) );
  AND2X1 U9134 ( .IN1(n5879), .IN2(n9200), .Q(n9196) );
  OR3X1 U9135 ( .IN1(n9201), .IN2(n9202), .IN3(n9203), .Q(n9194) );
  AND2X1 U9137 ( .IN1(n1338), .IN2(n9204), .Q(n9203) );
  OR4X1 U9138 ( .IN1(n9205), .IN2(n9206), .IN3(n9207), .IN4(n9208), .Q(n9204)
         );
  OR4X1 U9139 ( .IN1(n9209), .IN2(n9210), .IN3(n9211), .IN4(n9212), .Q(n9208)
         );
  OR3X1 U9140 ( .IN1(n9213), .IN2(n9214), .IN3(n9215), .Q(n9212) );
  AND2X1 U9141 ( .IN1(g37), .IN2(n9153), .Q(n9215) );
  AND2X1 U9142 ( .IN1(n9154), .IN2(g2868), .Q(n9214) );
  AND2X1 U9143 ( .IN1(n9155), .IN2(g758), .Q(n9211) );
  AND2X1 U9144 ( .IN1(n9156), .IN2(g2882), .Q(n9210) );
  AND2X1 U9145 ( .IN1(n9157), .IN2(g794), .Q(n9209) );
  OR3X1 U9146 ( .IN1(n9216), .IN2(n9217), .IN3(n9218), .Q(n9207) );
  AND2X1 U9147 ( .IN1(n9161), .IN2(g2955), .Q(n9218) );
  AND2X1 U9148 ( .IN1(n9162), .IN2(g2950), .Q(n9217) );
  AND2X1 U9149 ( .IN1(n9163), .IN2(g613), .Q(n9216) );
  AND2X1 U9150 ( .IN1(n9166), .IN2(g586), .Q(n9206) );
  AND2X1 U9151 ( .IN1(n9167), .IN2(g534), .Q(n9205) );
  AND2X1 U9152 ( .IN1(n9138), .IN2(g4300), .Q(n9202) );
  AND2X1 U9153 ( .IN1(n9139), .IN2(g4172), .Q(n9201) );
  AND2X1 U9154 ( .IN1(n9133), .IN2(g1291), .Q(n9193) );
  AND2X1 U9155 ( .IN1(n9140), .IN2(g947), .Q(n9192) );
  OR2X1 U9156 ( .IN1(n8459), .IN2(g34976), .Q(g34921) );
  OR4X1 U9157 ( .IN1(n9219), .IN2(n9220), .IN3(n9221), .IN4(n9222), .Q(g34976)
         );
  OR4X1 U9158 ( .IN1(n9223), .IN2(n9142), .IN3(n9224), .IN4(n9225), .Q(n9222)
         );
  AND2X1 U9159 ( .IN1(n9199), .IN2(g4722), .Q(n9225) );
  AND2X1 U9160 ( .IN1(n9134), .IN2(g5160), .Q(n9224) );
  AND2X1 U9161 ( .IN1(n9200), .IN2(g4912), .Q(n9223) );
  OR3X1 U9162 ( .IN1(n9226), .IN2(n9227), .IN3(n9228), .Q(n9221) );
  AND2X1 U9163 ( .IN1(n1338), .IN2(n9229), .Q(n9228) );
  OR4X1 U9164 ( .IN1(n9230), .IN2(n9231), .IN3(n9232), .IN4(n9233), .Q(n9229)
         );
  OR4X1 U9165 ( .IN1(n9234), .IN2(n9235), .IN3(n9237), .IN4(n9238), .Q(n9233)
         );
  OR3X1 U9166 ( .IN1(n9213), .IN2(n9239), .IN3(n9241), .Q(n9238) );
  AND2X1 U9167 ( .IN1(n9157), .IN2(g807), .Q(n9241) );
  AND2X1 U9168 ( .IN1(n9154), .IN2(g2988), .Q(n9239) );
  AND2X1 U9169 ( .IN1(n9163), .IN2(g617), .Q(n9237) );
  AND2X1 U9170 ( .IN1(n9155), .IN2(g763), .Q(n9235) );
  AND2X1 U9171 ( .IN1(n9156), .IN2(g2898), .Q(n9234) );
  OR3X1 U9172 ( .IN1(n9242), .IN2(n9243), .IN3(n9244), .Q(n9232) );
  AND2X1 U9173 ( .IN1(n9161), .IN2(g2941), .Q(n9244) );
  AND2X1 U9174 ( .IN1(test_so95), .IN2(n9246), .Q(n9243) );
  AND2X1 U9175 ( .IN1(n9162), .IN2(g2936), .Q(n9242) );
  AND2X1 U9176 ( .IN1(n9166), .IN2(g577), .Q(n9231) );
  AND2X1 U9177 ( .IN1(test_so41), .IN2(n9167), .Q(n9230) );
  AND2X1 U9178 ( .IN1(n9248), .IN2(g1135), .Q(n9227) );
  AND2X1 U9179 ( .IN1(n9249), .IN2(g1478), .Q(n9226) );
  AND2X1 U9180 ( .IN1(n9135), .IN2(g6545), .Q(n9220) );
  AND2X1 U9181 ( .IN1(n9132), .IN2(n9357), .Q(n9219) );
  OR2X1 U9182 ( .IN1(n8459), .IN2(g34975), .Q(g34919) );
  OR4X1 U9183 ( .IN1(n9250), .IN2(n9251), .IN3(n9252), .IN4(n9253), .Q(g34975)
         );
  OR4X1 U9184 ( .IN1(n9254), .IN2(n9142), .IN3(n9256), .IN4(n9257), .Q(n9253)
         );
  AND2X1 U9185 ( .IN1(n9199), .IN2(g4717), .Q(n9257) );
  AND2X1 U9186 ( .IN1(n9134), .IN2(g5507), .Q(n9256) );
  AND2X1 U9187 ( .IN1(n9200), .IN2(g4907), .Q(n9254) );
  OR3X1 U9188 ( .IN1(n9258), .IN2(n9259), .IN3(n9260), .Q(n9252) );
  AND2X1 U9189 ( .IN1(n1338), .IN2(n9261), .Q(n9260) );
  OR4X1 U9190 ( .IN1(n9263), .IN2(n9264), .IN3(n9266), .IN4(n9268), .Q(n9261)
         );
  OR4X1 U9191 ( .IN1(n9269), .IN2(n9270), .IN3(n9271), .IN4(n9272), .Q(n9268)
         );
  OR2X1 U9192 ( .IN1(n9275), .IN2(n9277), .Q(n9272) );
  AND2X1 U9193 ( .IN1(n9166), .IN2(g582), .Q(n9277) );
  AND2X1 U9194 ( .IN1(n9167), .IN2(g546), .Q(n9275) );
  AND2X1 U9195 ( .IN1(n9161), .IN2(g2927), .Q(n9271) );
  AND2X1 U9196 ( .IN1(n9246), .IN2(g2860), .Q(n9270) );
  AND2X1 U9197 ( .IN1(n9162), .IN2(g2922), .Q(n9269) );
  OR3X1 U9198 ( .IN1(n9278), .IN2(n9279), .IN3(n9282), .Q(n9266) );
  AND2X1 U9199 ( .IN1(n9156), .IN2(g2864), .Q(n9282) );
  AND2X1 U9200 ( .IN1(n9157), .IN2(g554), .Q(n9279) );
  AND2X1 U9201 ( .IN1(n5634), .IN2(n9154), .Q(n9278) );
  AND2X1 U9202 ( .IN1(n9163), .IN2(g622), .Q(n9264) );
  AND2X1 U9203 ( .IN1(n9155), .IN2(g767), .Q(n9263) );
  AND2X1 U9204 ( .IN1(n9248), .IN2(g1105), .Q(n9259) );
  AND2X1 U9205 ( .IN1(n9249), .IN2(g1448), .Q(n9258) );
  AND2X1 U9206 ( .IN1(n9135), .IN2(g3151), .Q(n9251) );
  AND2X1 U9207 ( .IN1(n9132), .IN2(n9294), .Q(n9250) );
  OR2X1 U9208 ( .IN1(n8459), .IN2(g34974), .Q(g34917) );
  OR4X1 U9209 ( .IN1(n9283), .IN2(n9284), .IN3(n9285), .IN4(n9286), .Q(g34974)
         );
  OR4X1 U9210 ( .IN1(n9287), .IN2(n9288), .IN3(n9289), .IN4(n9290), .Q(n9286)
         );
  AND2X1 U9211 ( .IN1(n9134), .IN2(g5853), .Q(n9290) );
  AND2X1 U9212 ( .IN1(test_so45), .IN2(n9135), .Q(n9289) );
  AND2X1 U9213 ( .IN1(n9200), .IN2(g4922), .Q(n9288) );
  AND2X1 U9214 ( .IN1(n9199), .IN2(g4732), .Q(n9287) );
  OR3X1 U9215 ( .IN1(n9291), .IN2(n9292), .IN3(n9293), .Q(n9285) );
  AND2X1 U9216 ( .IN1(n9248), .IN2(g1129), .Q(n9293) );
  AND2X1 U9217 ( .IN1(n9249), .IN2(g1472), .Q(n9292) );
  AND2X1 U9218 ( .IN1(n9132), .IN2(n9327), .Q(n9284) );
  AND2X1 U9219 ( .IN1(n1338), .IN2(n9296), .Q(n9283) );
  OR2X1 U9220 ( .IN1(n9297), .IN2(n9298), .Q(n9296) );
  OR4X1 U9221 ( .IN1(n9299), .IN2(n9300), .IN3(n9301), .IN4(n9304), .Q(n9298)
         );
  AND2X1 U9222 ( .IN1(n9246), .IN2(g2852), .Q(n9304) );
  AND2X1 U9223 ( .IN1(n9162), .IN2(g2912), .Q(n9301) );
  AND2X1 U9224 ( .IN1(n9166), .IN2(g590), .Q(n9300) );
  AND2X1 U9225 ( .IN1(n9161), .IN2(g2917), .Q(n9299) );
  OR4X1 U9226 ( .IN1(n9305), .IN2(n9307), .IN3(n9308), .IN4(n9309), .Q(n9297)
         );
  AND2X1 U9227 ( .IN1(n9156), .IN2(g2856), .Q(n9309) );
  AND2X1 U9228 ( .IN1(n9154), .IN2(g2999), .Q(n9308) );
  AND2X1 U9229 ( .IN1(n9163), .IN2(g626), .Q(n9307) );
  AND2X1 U9230 ( .IN1(n9155), .IN2(g772), .Q(n9305) );
  OR2X1 U9231 ( .IN1(n8459), .IN2(g34971), .Q(g34915) );
  OR4X1 U9232 ( .IN1(n9310), .IN2(n9311), .IN3(n9313), .IN4(n9315), .Q(g34971)
         );
  OR4X1 U9233 ( .IN1(n9316), .IN2(n9317), .IN3(n9318), .IN4(n9319), .Q(n9315)
         );
  AND2X1 U9234 ( .IN1(n9132), .IN2(n9351), .Q(n9319) );
  AND2X1 U9235 ( .IN1(test_so64), .IN2(n9133), .Q(n9318) );
  AND2X1 U9236 ( .IN1(n9134), .IN2(g2145), .Q(n9317) );
  AND2X1 U9237 ( .IN1(n9135), .IN2(g2704), .Q(n9316) );
  OR2X1 U9238 ( .IN1(n9320), .IN2(n9321), .Q(n9313) );
  AND2X1 U9239 ( .IN1(n9138), .IN2(g4245), .Q(n9321) );
  AND2X1 U9240 ( .IN1(n9323), .IN2(n9326), .Q(n9138) );
  AND2X1 U9241 ( .IN1(n9139), .IN2(g4157), .Q(n9320) );
  AND2X1 U9242 ( .IN1(n1338), .IN2(n9246), .Q(n9139) );
  AND2X1 U9243 ( .IN1(n9140), .IN2(n9247), .Q(n9311) );
  AND2X1 U9244 ( .IN1(n1338), .IN2(n9328), .Q(n9310) );
  OR4X1 U9245 ( .IN1(n9329), .IN2(n9142), .IN3(n9330), .IN4(n9331), .Q(n9328)
         );
  OR4X1 U9246 ( .IN1(n9333), .IN2(n9334), .IN3(n9335), .IN4(n9337), .Q(n9331)
         );
  OR2X1 U9247 ( .IN1(n9213), .IN2(n9338), .Q(n9337) );
  AND2X1 U9248 ( .IN1(n9154), .IN2(g2890), .Q(n9338) );
  AND2X1 U9249 ( .IN1(n9326), .IN2(n9339), .Q(n9154) );
  AND4X1 U9250 ( .IN1(g28), .IN2(n9341), .IN3(n5477), .IN4(g19), .Q(n9213) );
  AND2X1 U9251 ( .IN1(g100), .IN2(n9153), .Q(n9335) );
  AND3X1 U9252 ( .IN1(g28), .IN2(n9342), .IN3(n9339), .Q(n9153) );
  AND2X1 U9253 ( .IN1(n9157), .IN2(g781), .Q(n9334) );
  AND2X1 U9254 ( .IN1(n9090), .IN2(g2984), .Q(n9333) );
  AND4X1 U9255 ( .IN1(test_so25), .IN2(n9341), .IN3(n5324), .IN4(n8447), .Q(
        n9090) );
  OR3X1 U9256 ( .IN1(n9343), .IN2(n9344), .IN3(n9345), .Q(n9330) );
  AND2X1 U9257 ( .IN1(n9167), .IN2(g199), .Q(n9345) );
  AND2X1 U9258 ( .IN1(n9163), .IN2(g599), .Q(n9344) );
  AND2X1 U9259 ( .IN1(test_so60), .IN2(n9155), .Q(n9343) );
  OR2X1 U9260 ( .IN1(n9346), .IN2(n9291), .Q(n9142) );
  AND3X1 U9261 ( .IN1(n1338), .IN2(n8841), .IN3(n9157), .Q(n9346) );
  AND2X1 U9262 ( .IN1(n9326), .IN2(n9347), .Q(n9157) );
  AND2X1 U9263 ( .IN1(n9166), .IN2(g562), .Q(n9329) );
  OR2X1 U9264 ( .IN1(n8459), .IN2(g34970), .Q(g34913) );
  OR4X1 U9265 ( .IN1(n9349), .IN2(n9350), .IN3(n9353), .IN4(n9354), .Q(g34970)
         );
  OR4X1 U9266 ( .IN1(n9355), .IN2(n9356), .IN3(n9358), .IN4(n9359), .Q(n9354)
         );
  AND2X1 U9267 ( .IN1(n1338), .IN2(n9360), .Q(n9359) );
  OR2X1 U9268 ( .IN1(n9361), .IN2(n9362), .Q(n9360) );
  OR4X1 U9269 ( .IN1(n9363), .IN2(n9364), .IN3(n9365), .IN4(n9366), .Q(n9362)
         );
  AND2X1 U9270 ( .IN1(n9161), .IN2(g2902), .Q(n9366) );
  AND3X1 U9271 ( .IN1(n5324), .IN2(n9368), .IN3(n9341), .Q(n9161) );
  AND2X1 U9272 ( .IN1(n9246), .IN2(g2844), .Q(n9365) );
  AND3X1 U9273 ( .IN1(g9), .IN2(n9368), .IN3(n9369), .Q(n9246) );
  AND2X1 U9274 ( .IN1(n9166), .IN2(g595), .Q(n9364) );
  AND2X1 U9275 ( .IN1(n9167), .IN2(g538), .Q(n9363) );
  AND2X1 U9276 ( .IN1(n9369), .IN2(n9347), .Q(n9167) );
  OR4X1 U9277 ( .IN1(n9370), .IN2(n9371), .IN3(n9372), .IN4(n9373), .Q(n9361)
         );
  AND2X1 U9278 ( .IN1(n9155), .IN2(g776), .Q(n9373) );
  AND2X1 U9279 ( .IN1(n9156), .IN2(g2848), .Q(n9372) );
  AND3X1 U9280 ( .IN1(g9), .IN2(n9368), .IN3(n9326), .Q(n9156) );
  AND2X1 U9281 ( .IN1(test_so1), .IN2(n9162), .Q(n9371) );
  AND3X1 U9282 ( .IN1(g28), .IN2(n9368), .IN3(n9341), .Q(n9162) );
  AND4X1 U9283 ( .IN1(n3395), .IN2(test_so85), .IN3(g8), .IN4(g9), .Q(n9341)
         );
  AND2X1 U9284 ( .IN1(n9163), .IN2(n9340), .Q(n9370) );
  AND2X1 U9285 ( .IN1(n9134), .IN2(g6199), .Q(n9358) );
  AND2X1 U9286 ( .IN1(n9369), .IN2(n9323), .Q(n9134) );
  AND2X1 U9287 ( .IN1(n9200), .IN2(g4917), .Q(n9356) );
  AND3X1 U9288 ( .IN1(n1338), .IN2(n9326), .IN3(n2527), .Q(n9200) );
  AND2X1 U9289 ( .IN1(n9199), .IN2(g4727), .Q(n9355) );
  AND3X1 U9290 ( .IN1(n9369), .IN2(n1338), .IN3(n2527), .Q(n9199) );
  OR3X1 U9291 ( .IN1(n9291), .IN2(n9374), .IN3(n9375), .Q(n9353) );
  AND2X1 U9292 ( .IN1(n9248), .IN2(g956), .Q(n9375) );
  AND2X1 U9293 ( .IN1(n9140), .IN2(n5286), .Q(n9248) );
  AND3X1 U9294 ( .IN1(n1338), .IN2(n9326), .IN3(n2552), .Q(n9140) );
  AND3X1 U9295 ( .IN1(g28), .IN2(n9376), .IN3(n5469), .Q(n9326) );
  AND2X1 U9296 ( .IN1(n9249), .IN2(g1300), .Q(n9374) );
  AND2X1 U9297 ( .IN1(n9133), .IN2(n2549), .Q(n9249) );
  AND3X1 U9298 ( .IN1(n9369), .IN2(n1338), .IN3(n9339), .Q(n9133) );
  AND3X1 U9299 ( .IN1(n8447), .IN2(n5468), .IN3(test_so25), .Q(n9339) );
  AND3X1 U9300 ( .IN1(n8841), .IN2(n9377), .IN3(n1338), .Q(n9291) );
  OR3X1 U9301 ( .IN1(n9163), .IN2(n9166), .IN3(n9155), .Q(n9377) );
  AND3X1 U9302 ( .IN1(g28), .IN2(n9347), .IN3(n9342), .Q(n9155) );
  AND2X1 U9303 ( .IN1(n9368), .IN2(n5468), .Q(n9347) );
  AND2X1 U9304 ( .IN1(n5477), .IN2(n8447), .Q(n9368) );
  AND3X1 U9305 ( .IN1(n5324), .IN2(n9342), .IN3(n2552), .Q(n9166) );
  AND2X1 U9306 ( .IN1(n9369), .IN2(n2552), .Q(n9163) );
  AND3X1 U9307 ( .IN1(n9376), .IN2(n5324), .IN3(n5469), .Q(n9369) );
  AND2X1 U9308 ( .IN1(n9135), .IN2(g3853), .Q(n9350) );
  AND3X1 U9309 ( .IN1(n5324), .IN2(n9323), .IN3(n9342), .Q(n9135) );
  AND2X1 U9310 ( .IN1(g31), .IN2(n9376), .Q(n9342) );
  INVX0 U9311 ( .INP(n9378), .ZN(n9376) );
  OR3X1 U9312 ( .IN1(test_so85), .IN2(g8), .IN3(g6), .Q(n9378) );
  AND4X1 U9313 ( .IN1(g9), .IN2(n1338), .IN3(n5477), .IN4(g19), .Q(n9323) );
  INVX0 U9314 ( .INP(n9379), .ZN(n1338) );
  AND2X1 U9316 ( .IN1(n9132), .IN2(n9322), .Q(n9349) );
  AND2X1 U9317 ( .IN1(n9116), .IN2(n9379), .Q(n9132) );
  OR4X1 U9318 ( .IN1(g53), .IN2(n9123), .IN3(test_so74), .IN4(g57), .Q(n9379)
         );
  OR2X1 U9319 ( .IN1(g56), .IN2(n9117), .Q(n9123) );
  INVX0 U9320 ( .INP(g54), .ZN(n9117) );
  INVX0 U9321 ( .INP(g53), .ZN(n9116) );
  OR2X1 U9322 ( .IN1(n9380), .IN2(n9381), .Q(g34911) );
  AND2X1 U9323 ( .IN1(n2404), .IN2(g554), .Q(n9381) );
  AND2X1 U9324 ( .IN1(n9382), .IN2(g807), .Q(n9380) );
  OR2X1 U9325 ( .IN1(n2405), .IN2(n8794), .Q(n9382) );
  OR2X1 U9326 ( .IN1(n9383), .IN2(n9384), .Q(g34882) );
  AND2X1 U9327 ( .IN1(n9385), .IN2(n8700), .Q(n9384) );
  OR3X1 U9328 ( .IN1(n9386), .IN2(n9387), .IN3(n9388), .Q(n9385) );
  AND3X1 U9329 ( .IN1(n5653), .IN2(n9389), .IN3(n9390), .Q(n9388) );
  OR2X1 U9330 ( .IN1(g4358), .IN2(n9391), .Q(n9389) );
  AND3X1 U9331 ( .IN1(n9391), .IN2(n8492), .IN3(n5348), .Q(n9387) );
  OR4X1 U9332 ( .IN1(test_so81), .IN2(g4340), .IN3(n9392), .IN4(n9393), .Q(
        n9391) );
  AND3X1 U9333 ( .IN1(n5506), .IN2(g4311), .IN3(g4332), .Q(n9393) );
  AND2X1 U9334 ( .IN1(n5540), .IN2(n9394), .Q(n9392) );
  OR3X1 U9335 ( .IN1(n9395), .IN2(n9396), .IN3(n9397), .Q(n9394) );
  AND3X1 U9336 ( .IN1(g90), .IN2(n5634), .IN3(n5506), .Q(n9396) );
  AND2X1 U9337 ( .IN1(n8223), .IN2(g4322), .Q(n9395) );
  AND3X1 U9338 ( .IN1(test_so81), .IN2(g4340), .IN3(g4358), .Q(n9386) );
  AND2X1 U9339 ( .IN1(n8829), .IN2(g4366), .Q(n9383) );
  OR3X1 U9340 ( .IN1(n9398), .IN2(n9399), .IN3(n9400), .Q(g34881) );
  AND2X1 U9341 ( .IN1(n8827), .IN2(g794), .Q(n9400) );
  AND2X1 U9342 ( .IN1(n2405), .IN2(n5479), .Q(n9399) );
  AND3X1 U9343 ( .IN1(n2404), .IN2(n9401), .IN3(g807), .Q(n9398) );
  INVX0 U9344 ( .INP(n2405), .ZN(n9401) );
  OR3X1 U9345 ( .IN1(n9402), .IN2(n9403), .IN3(n9404), .Q(g34880) );
  AND2X1 U9346 ( .IN1(n8827), .IN2(g626), .Q(n9404) );
  AND2X1 U9347 ( .IN1(n2422), .IN2(n14833), .Q(n9403) );
  AND3X1 U9348 ( .IN1(n2421), .IN2(n9405), .IN3(n9340), .Q(n9402) );
  INVX0 U9349 ( .INP(n2422), .ZN(n9405) );
  OR3X1 U9350 ( .IN1(n9406), .IN2(n9407), .IN3(n9408), .Q(g34850) );
  AND2X1 U9351 ( .IN1(n8827), .IN2(g790), .Q(n9408) );
  AND2X1 U9352 ( .IN1(n2419), .IN2(n5291), .Q(n9407) );
  AND3X1 U9353 ( .IN1(n2404), .IN2(n9409), .IN3(g794), .Q(n9406) );
  INVX0 U9354 ( .INP(n2419), .ZN(n9409) );
  OR3X1 U9355 ( .IN1(n9410), .IN2(n9411), .IN3(n9412), .Q(g34849) );
  AND2X1 U9356 ( .IN1(n8827), .IN2(g622), .Q(n9412) );
  AND2X1 U9357 ( .IN1(n2423), .IN2(n5288), .Q(n9411) );
  AND3X1 U9358 ( .IN1(n2421), .IN2(n9413), .IN3(g626), .Q(n9410) );
  INVX0 U9359 ( .INP(n2423), .ZN(n9413) );
  AND2X1 U9360 ( .IN1(n9414), .IN2(g4369), .Q(g34839) );
  OR3X1 U9361 ( .IN1(n9415), .IN2(n9416), .IN3(g4366), .Q(n9414) );
  AND2X1 U9362 ( .IN1(n9417), .IN2(g4332), .Q(n9416) );
  OR3X1 U9363 ( .IN1(n9418), .IN2(g4311), .IN3(n9419), .Q(n9417) );
  AND2X1 U9364 ( .IN1(n5540), .IN2(n9420), .Q(n9415) );
  OR3X1 U9365 ( .IN1(g73), .IN2(n9418), .IN3(g4311), .Q(n9420) );
  OR2X1 U9366 ( .IN1(n9421), .IN2(n9422), .Q(g34808) );
  AND2X1 U9367 ( .IN1(n9423), .IN2(n8700), .Q(n9422) );
  OR3X1 U9368 ( .IN1(n9424), .IN2(n9425), .IN3(g2965), .Q(n9423) );
  AND2X1 U9369 ( .IN1(n8827), .IN2(g2955), .Q(n9421) );
  OR2X1 U9370 ( .IN1(n9426), .IN2(n9427), .Q(g34807) );
  AND2X1 U9371 ( .IN1(n9428), .IN2(n8700), .Q(n9427) );
  OR4X1 U9372 ( .IN1(n9429), .IN2(n9430), .IN3(n9431), .IN4(n9432), .Q(n9428)
         );
  OR3X1 U9373 ( .IN1(n9433), .IN2(g2955), .IN3(g2946), .Q(n9432) );
  AND2X1 U9374 ( .IN1(n8827), .IN2(g2941), .Q(n9426) );
  OR2X1 U9375 ( .IN1(n9434), .IN2(n9435), .Q(g34806) );
  AND2X1 U9376 ( .IN1(n9436), .IN2(n8700), .Q(n9435) );
  OR3X1 U9377 ( .IN1(g2941), .IN2(g4072), .IN3(g4153), .Q(n9436) );
  AND2X1 U9378 ( .IN1(n8827), .IN2(g2927), .Q(n9434) );
  AND2X1 U9379 ( .IN1(n9437), .IN2(n8700), .Q(g34805) );
  OR2X1 U9380 ( .IN1(g2932), .IN2(g2999), .Q(n9437) );
  OR2X1 U9381 ( .IN1(n9438), .IN2(n9439), .Q(g34804) );
  AND2X1 U9382 ( .IN1(n9440), .IN2(n8701), .Q(n9439) );
  OR3X1 U9383 ( .IN1(n5796), .IN2(n5630), .IN3(g2975), .Q(n9440) );
  AND2X1 U9384 ( .IN1(n8827), .IN2(g2965), .Q(n9438) );
  OR2X1 U9385 ( .IN1(n9441), .IN2(n9442), .Q(g34803) );
  AND2X1 U9386 ( .IN1(n9443), .IN2(n8701), .Q(n9442) );
  OR3X1 U9387 ( .IN1(g2932), .IN2(n9444), .IN3(g2927), .Q(n9443) );
  AND2X1 U9388 ( .IN1(n8827), .IN2(g2917), .Q(n9441) );
  OR2X1 U9389 ( .IN1(n9445), .IN2(n9446), .Q(g34802) );
  AND2X1 U9390 ( .IN1(n9447), .IN2(n8701), .Q(n9446) );
  OR3X1 U9391 ( .IN1(n9448), .IN2(n9449), .IN3(g2917), .Q(n9447) );
  AND2X1 U9392 ( .IN1(n8827), .IN2(g2902), .Q(n9445) );
  OR2X1 U9393 ( .IN1(n9450), .IN2(n9451), .Q(g34801) );
  AND2X1 U9394 ( .IN1(n9452), .IN2(n8701), .Q(n9451) );
  OR4X1 U9395 ( .IN1(g2902), .IN2(g301), .IN3(n5520), .IN4(g209), .Q(n9452) );
  AND2X1 U9396 ( .IN1(n8827), .IN2(g2970), .Q(n9450) );
  OR2X1 U9397 ( .IN1(n9453), .IN2(n9454), .Q(g34800) );
  AND2X1 U9398 ( .IN1(n9455), .IN2(n8701), .Q(n9454) );
  OR2X1 U9399 ( .IN1(test_so14), .IN2(test_so74), .Q(n9455) );
  AND2X1 U9400 ( .IN1(n8827), .IN2(g2886), .Q(n9453) );
  OR2X1 U9401 ( .IN1(n9456), .IN2(n9457), .Q(g34799) );
  AND2X1 U9402 ( .IN1(n9458), .IN2(n8701), .Q(n9457) );
  OR2X1 U9403 ( .IN1(n9444), .IN2(g2890), .Q(n9458) );
  INVX0 U9404 ( .INP(g44), .ZN(n9444) );
  AND2X1 U9405 ( .IN1(n8827), .IN2(g2873), .Q(n9456) );
  OR2X1 U9406 ( .IN1(n9459), .IN2(n9460), .Q(g34798) );
  AND2X1 U9407 ( .IN1(n9461), .IN2(n8701), .Q(n9460) );
  OR2X1 U9408 ( .IN1(g2946), .IN2(g2886), .Q(n9461) );
  AND2X1 U9409 ( .IN1(n8827), .IN2(g2878), .Q(n9459) );
  OR2X1 U9410 ( .IN1(n9462), .IN2(n9463), .Q(g34797) );
  AND2X1 U9411 ( .IN1(n9464), .IN2(n8701), .Q(n9463) );
  OR2X1 U9412 ( .IN1(n9425), .IN2(g2878), .Q(n9464) );
  INVX0 U9413 ( .INP(g91), .ZN(n9425) );
  AND2X1 U9414 ( .IN1(n8827), .IN2(g2882), .Q(n9462) );
  OR2X1 U9415 ( .IN1(n9465), .IN2(n9466), .Q(g34796) );
  AND2X1 U9416 ( .IN1(n9467), .IN2(n8702), .Q(n9466) );
  OR2X1 U9417 ( .IN1(n9424), .IN2(g2882), .Q(n9467) );
  OR2X1 U9418 ( .IN1(n9468), .IN2(n9469), .Q(n9424) );
  AND2X1 U9419 ( .IN1(n8827), .IN2(g2898), .Q(n9465) );
  OR2X1 U9420 ( .IN1(n9470), .IN2(n9471), .Q(g34795) );
  AND2X1 U9421 ( .IN1(n9472), .IN2(n8702), .Q(n9471) );
  OR2X1 U9422 ( .IN1(n9430), .IN2(g2898), .Q(n9472) );
  INVX0 U9423 ( .INP(n9473), .ZN(n9430) );
  AND4X1 U9424 ( .IN1(n9474), .IN2(n9475), .IN3(n9476), .IN4(n9477), .Q(n9473)
         );
  AND2X1 U9425 ( .IN1(n5861), .IN2(n5882), .Q(n9477) );
  AND2X1 U9426 ( .IN1(n8828), .IN2(g2864), .Q(n9470) );
  OR2X1 U9427 ( .IN1(n9478), .IN2(n9479), .Q(g34794) );
  AND2X1 U9428 ( .IN1(n9480), .IN2(n8702), .Q(n9479) );
  OR2X1 U9429 ( .IN1(n9431), .IN2(g2864), .Q(n9480) );
  INVX0 U9430 ( .INP(n9481), .ZN(n9431) );
  AND3X1 U9431 ( .IN1(n9482), .IN2(n9483), .IN3(n9484), .Q(n9481) );
  AND2X1 U9432 ( .IN1(n8828), .IN2(g2856), .Q(n9478) );
  OR2X1 U9433 ( .IN1(n9485), .IN2(n9486), .Q(g34793) );
  AND2X1 U9434 ( .IN1(n9487), .IN2(n8702), .Q(n9486) );
  OR2X1 U9435 ( .IN1(n9429), .IN2(g2856), .Q(n9487) );
  OR2X1 U9436 ( .IN1(n9488), .IN2(n9489), .Q(n9429) );
  AND2X1 U9437 ( .IN1(n8828), .IN2(g2848), .Q(n9485) );
  OR2X1 U9438 ( .IN1(n9490), .IN2(n9491), .Q(g34792) );
  AND2X1 U9439 ( .IN1(n9492), .IN2(n8702), .Q(n9491) );
  OR2X1 U9440 ( .IN1(n9433), .IN2(g2848), .Q(n9492) );
  INVX0 U9441 ( .INP(n9493), .ZN(n9433) );
  AND2X1 U9442 ( .IN1(n9494), .IN2(n9495), .Q(n9493) );
  AND2X1 U9443 ( .IN1(n8828), .IN2(g29214), .Q(n9490) );
  OR3X1 U9444 ( .IN1(n9496), .IN2(n9497), .IN3(n9498), .Q(g34791) );
  AND2X1 U9445 ( .IN1(n8828), .IN2(g785), .Q(n9498) );
  AND2X1 U9446 ( .IN1(n2425), .IN2(n5292), .Q(n9497) );
  AND3X1 U9447 ( .IN1(n2404), .IN2(n9499), .IN3(g790), .Q(n9496) );
  INVX0 U9448 ( .INP(n2425), .ZN(n9499) );
  OR3X1 U9449 ( .IN1(n9500), .IN2(n9501), .IN3(n9502), .Q(g34790) );
  AND2X1 U9450 ( .IN1(n8828), .IN2(g617), .Q(n9502) );
  AND2X1 U9451 ( .IN1(n2427), .IN2(n5672), .Q(n9501) );
  AND3X1 U9452 ( .IN1(n2421), .IN2(n9503), .IN3(g622), .Q(n9500) );
  INVX0 U9454 ( .INP(n2427), .ZN(n9503) );
  AND2X1 U9455 ( .IN1(n9504), .IN2(g890), .Q(g34788) );
  OR2X1 U9456 ( .IN1(n8031), .IN2(n9505), .Q(n9504) );
  INVX0 U9457 ( .INP(n3195), .ZN(n9505) );
  OR2X1 U9458 ( .IN1(n9506), .IN2(n9507), .Q(g34783) );
  AND3X1 U9459 ( .IN1(n9508), .IN2(n9509), .IN3(n9510), .Q(n9507) );
  AND3X1 U9460 ( .IN1(n9511), .IN2(n9512), .IN3(n9513), .Q(n9506) );
  OR2X1 U9461 ( .IN1(n9514), .IN2(n9515), .Q(g34735) );
  AND2X1 U9462 ( .IN1(n9516), .IN2(n8703), .Q(n9515) );
  OR2X1 U9463 ( .IN1(test_so63), .IN2(g4300), .Q(n9516) );
  AND2X1 U9464 ( .IN1(n8828), .IN2(g4297), .Q(n9514) );
  OR2X1 U9465 ( .IN1(n9517), .IN2(n9518), .Q(g34734) );
  AND2X1 U9466 ( .IN1(n9519), .IN2(n8703), .Q(n9518) );
  OR2X1 U9467 ( .IN1(g4072), .IN2(g4176), .Q(n9519) );
  AND2X1 U9468 ( .IN1(n8828), .IN2(g4172), .Q(n9517) );
  AND2X1 U9469 ( .IN1(n9520), .IN2(n8702), .Q(g34733) );
  OR2X1 U9470 ( .IN1(g4153), .IN2(g4172), .Q(n9520) );
  OR2X1 U9471 ( .IN1(n9521), .IN2(n9522), .Q(g34732) );
  AND2X1 U9472 ( .IN1(n8828), .IN2(g2999), .Q(n9522) );
  AND2X1 U9473 ( .IN1(n8705), .IN2(g2994), .Q(n9521) );
  OR2X1 U9474 ( .IN1(n9523), .IN2(n9524), .Q(g34731) );
  AND2X1 U9475 ( .IN1(n9525), .IN2(n8703), .Q(n9524) );
  OR2X1 U9476 ( .IN1(test_so64), .IN2(n9448), .Q(n9525) );
  AND2X1 U9477 ( .IN1(n8828), .IN2(g1283), .Q(n9523) );
  OR2X1 U9478 ( .IN1(n9526), .IN2(n9527), .Q(g34730) );
  AND2X1 U9479 ( .IN1(n9528), .IN2(n8704), .Q(n9527) );
  OR2X1 U9480 ( .IN1(g1283), .IN2(g1277), .Q(n9528) );
  AND2X1 U9481 ( .IN1(n8828), .IN2(g1296), .Q(n9526) );
  OR3X1 U9482 ( .IN1(n9529), .IN2(n9530), .IN3(n2499), .Q(g34729) );
  AND2X1 U9483 ( .IN1(n8828), .IN2(g1291), .Q(n9530) );
  AND2X1 U9484 ( .IN1(n5796), .IN2(n8703), .Q(n9529) );
  OR2X1 U9485 ( .IN1(n9531), .IN2(n9532), .Q(g34728) );
  AND2X1 U9486 ( .IN1(n9533), .IN2(n8703), .Q(n9532) );
  OR2X1 U9487 ( .IN1(n9449), .IN2(n9247), .Q(n9533) );
  AND2X1 U9488 ( .IN1(n8828), .IN2(g939), .Q(n9531) );
  OR2X1 U9489 ( .IN1(n9534), .IN2(n9535), .Q(g34727) );
  AND2X1 U9490 ( .IN1(n9536), .IN2(n8704), .Q(n9535) );
  OR2X1 U9491 ( .IN1(test_so52), .IN2(g939), .Q(n9536) );
  AND2X1 U9492 ( .IN1(n8828), .IN2(g952), .Q(n9534) );
  OR3X1 U9493 ( .IN1(n9537), .IN2(n9538), .IN3(n2505), .Q(g34726) );
  AND2X1 U9494 ( .IN1(n8828), .IN2(g947), .Q(n9538) );
  AND2X1 U9495 ( .IN1(n5630), .IN2(n8703), .Q(n9537) );
  OR3X1 U9496 ( .IN1(n9539), .IN2(n9540), .IN3(n9541), .Q(g34725) );
  AND2X1 U9497 ( .IN1(n8828), .IN2(g781), .Q(n9541) );
  AND2X1 U9498 ( .IN1(n2485), .IN2(n5293), .Q(n9540) );
  AND3X1 U9499 ( .IN1(n2404), .IN2(n9542), .IN3(g785), .Q(n9539) );
  INVX0 U9500 ( .INP(n2485), .ZN(n9542) );
  OR3X1 U9501 ( .IN1(n9543), .IN2(n9544), .IN3(n9545), .Q(g34724) );
  AND2X1 U9502 ( .IN1(n8828), .IN2(g613), .Q(n9545) );
  AND2X1 U9503 ( .IN1(n2487), .IN2(n5339), .Q(n9544) );
  AND3X1 U9504 ( .IN1(n2421), .IN2(n9546), .IN3(g617), .Q(n9543) );
  INVX0 U9505 ( .INP(n2487), .ZN(n9546) );
  OR2X1 U9506 ( .IN1(n9547), .IN2(n9548), .Q(g34723) );
  AND2X1 U9507 ( .IN1(n9549), .IN2(n8703), .Q(n9548) );
  OR2X1 U9508 ( .IN1(g301), .IN2(g534), .Q(n9549) );
  AND2X1 U9509 ( .IN1(test_so41), .IN2(n8810), .Q(n9547) );
  OR2X1 U9510 ( .IN1(n9550), .IN2(n9551), .Q(g34722) );
  AND2X1 U9511 ( .IN1(n9552), .IN2(n8704), .Q(n9551) );
  OR2X1 U9512 ( .IN1(n5520), .IN2(g546), .Q(n9552) );
  AND2X1 U9513 ( .IN1(n8828), .IN2(g538), .Q(n9550) );
  OR2X1 U9514 ( .IN1(n9553), .IN2(n9554), .Q(g34721) );
  AND2X1 U9515 ( .IN1(n9555), .IN2(n8704), .Q(n9554) );
  OR2X1 U9516 ( .IN1(g199), .IN2(g222), .Q(n9555) );
  AND2X1 U9517 ( .IN1(g29221), .IN2(n8810), .Q(n9553) );
  OR2X1 U9518 ( .IN1(n9556), .IN2(n9557), .Q(g34720) );
  AND2X1 U9519 ( .IN1(n9558), .IN2(n8704), .Q(n9557) );
  OR2X1 U9520 ( .IN1(n5657), .IN2(g550), .Q(n9558) );
  AND2X1 U9521 ( .IN1(n8828), .IN2(g534), .Q(n9556) );
  AND2X1 U9522 ( .IN1(n9559), .IN2(n8702), .Q(g34719) );
  OR2X1 U9523 ( .IN1(g209), .IN2(g538), .Q(n9559) );
  AND2X1 U9524 ( .IN1(n8709), .IN2(g6545), .Q(g34647) );
  AND2X1 U9525 ( .IN1(n8708), .IN2(g6199), .Q(g34646) );
  AND2X1 U9526 ( .IN1(n8709), .IN2(g5853), .Q(g34645) );
  AND2X1 U9527 ( .IN1(n8709), .IN2(g5507), .Q(g34644) );
  AND2X1 U9528 ( .IN1(n8709), .IN2(g5160), .Q(g34643) );
  OR2X1 U9529 ( .IN1(n9560), .IN2(n9561), .Q(g34642) );
  AND2X1 U9530 ( .IN1(n8828), .IN2(g4912), .Q(n9561) );
  AND2X1 U9531 ( .IN1(n8710), .IN2(g4927), .Q(n9560) );
  OR2X1 U9532 ( .IN1(n9562), .IN2(n9563), .Q(g34641) );
  AND2X1 U9533 ( .IN1(n8828), .IN2(g4907), .Q(n9563) );
  AND2X1 U9534 ( .IN1(n8710), .IN2(g4912), .Q(n9562) );
  OR2X1 U9535 ( .IN1(n9564), .IN2(n9565), .Q(g34640) );
  AND2X1 U9536 ( .IN1(n8828), .IN2(g4922), .Q(n9565) );
  AND2X1 U9537 ( .IN1(n8710), .IN2(g4907), .Q(n9564) );
  OR2X1 U9538 ( .IN1(n9566), .IN2(n9567), .Q(g34639) );
  AND2X1 U9539 ( .IN1(n8829), .IN2(g4917), .Q(n9567) );
  AND2X1 U9540 ( .IN1(n8710), .IN2(g4922), .Q(n9566) );
  AND2X1 U9541 ( .IN1(n8711), .IN2(g4917), .Q(g34638) );
  OR2X1 U9542 ( .IN1(n9568), .IN2(n9569), .Q(g34637) );
  AND2X1 U9543 ( .IN1(n8829), .IN2(g4722), .Q(n9569) );
  AND2X1 U9544 ( .IN1(n8711), .IN2(g4737), .Q(n9568) );
  OR2X1 U9545 ( .IN1(n9570), .IN2(n9571), .Q(g34636) );
  AND2X1 U9546 ( .IN1(n8829), .IN2(g4717), .Q(n9571) );
  AND2X1 U9547 ( .IN1(n8711), .IN2(g4722), .Q(n9570) );
  OR2X1 U9548 ( .IN1(n9572), .IN2(n9573), .Q(g34635) );
  AND2X1 U9549 ( .IN1(n8829), .IN2(g4732), .Q(n9573) );
  AND2X1 U9550 ( .IN1(n8712), .IN2(g4717), .Q(n9572) );
  OR2X1 U9551 ( .IN1(n9574), .IN2(n9575), .Q(g34634) );
  AND2X1 U9552 ( .IN1(n8829), .IN2(g4727), .Q(n9575) );
  AND2X1 U9553 ( .IN1(n8712), .IN2(g4732), .Q(n9574) );
  AND2X1 U9554 ( .IN1(n8712), .IN2(g4727), .Q(g34633) );
  OR2X1 U9555 ( .IN1(n9576), .IN2(n9577), .Q(g34632) );
  AND2X1 U9556 ( .IN1(test_so67), .IN2(n8810), .Q(n9577) );
  AND2X1 U9557 ( .IN1(n8712), .IN2(g4245), .Q(n9576) );
  OR2X1 U9558 ( .IN1(n9578), .IN2(n9579), .Q(g34631) );
  AND2X1 U9559 ( .IN1(n8829), .IN2(g4253), .Q(n9579) );
  AND2X1 U9560 ( .IN1(test_so67), .IN2(n8689), .Q(n9578) );
  OR2X1 U9561 ( .IN1(n9580), .IN2(n9581), .Q(g34630) );
  AND2X1 U9562 ( .IN1(n8829), .IN2(g4300), .Q(n9581) );
  AND2X1 U9563 ( .IN1(n8712), .IN2(g4253), .Q(n9580) );
  OR2X1 U9564 ( .IN1(n9582), .IN2(n9583), .Q(g34629) );
  AND2X1 U9565 ( .IN1(n8829), .IN2(g4146), .Q(n9583) );
  AND2X1 U9566 ( .IN1(n8711), .IN2(g4157), .Q(n9582) );
  OR2X1 U9567 ( .IN1(n9584), .IN2(n9585), .Q(g34628) );
  AND2X1 U9568 ( .IN1(n8829), .IN2(g4176), .Q(n9585) );
  AND2X1 U9569 ( .IN1(n8711), .IN2(g4146), .Q(n9584) );
  AND2X1 U9570 ( .IN1(n8711), .IN2(g3853), .Q(g34627) );
  AND2X1 U9571 ( .IN1(test_so45), .IN2(n8689), .Q(g34626) );
  AND2X1 U9572 ( .IN1(n8711), .IN2(g3151), .Q(g34625) );
  OR2X1 U9573 ( .IN1(n9586), .IN2(n9587), .Q(g34624) );
  AND2X1 U9574 ( .IN1(n8829), .IN2(g2994), .Q(n9587) );
  AND2X1 U9575 ( .IN1(n8711), .IN2(g2988), .Q(n9586) );
  OR2X1 U9576 ( .IN1(n9588), .IN2(n9589), .Q(g34623) );
  AND2X1 U9577 ( .IN1(test_so22), .IN2(n8811), .Q(n9589) );
  AND2X1 U9578 ( .IN1(n8710), .IN2(g2970), .Q(n9588) );
  OR2X1 U9579 ( .IN1(n9590), .IN2(n9591), .Q(g34622) );
  AND2X1 U9580 ( .IN1(n8829), .IN2(g2950), .Q(n9591) );
  AND2X1 U9581 ( .IN1(test_so22), .IN2(n8689), .Q(n9590) );
  OR2X1 U9582 ( .IN1(n9592), .IN2(n9593), .Q(g34621) );
  AND2X1 U9583 ( .IN1(n8829), .IN2(g2936), .Q(n9593) );
  AND2X1 U9584 ( .IN1(n8710), .IN2(g2950), .Q(n9592) );
  OR2X1 U9585 ( .IN1(n9594), .IN2(n9595), .Q(g34620) );
  AND2X1 U9586 ( .IN1(n8829), .IN2(g2922), .Q(n9595) );
  AND2X1 U9587 ( .IN1(n8710), .IN2(g2936), .Q(n9594) );
  OR2X1 U9588 ( .IN1(n9596), .IN2(n9597), .Q(g34619) );
  AND2X1 U9589 ( .IN1(n8829), .IN2(g2912), .Q(n9597) );
  AND2X1 U9590 ( .IN1(n8709), .IN2(g2922), .Q(n9596) );
  OR2X1 U9591 ( .IN1(n9598), .IN2(n9599), .Q(g34618) );
  AND2X1 U9592 ( .IN1(test_so1), .IN2(n8810), .Q(n9599) );
  AND2X1 U9593 ( .IN1(n8708), .IN2(g2912), .Q(n9598) );
  OR2X1 U9594 ( .IN1(n9600), .IN2(n9601), .Q(g34617) );
  AND2X1 U9595 ( .IN1(n8829), .IN2(g2984), .Q(n9601) );
  AND2X1 U9596 ( .IN1(test_so1), .IN2(n8687), .Q(n9600) );
  OR2X1 U9597 ( .IN1(n9602), .IN2(n9603), .Q(g34616) );
  AND2X1 U9598 ( .IN1(n8829), .IN2(g2988), .Q(n9603) );
  AND2X1 U9599 ( .IN1(n8708), .IN2(g2868), .Q(n9602) );
  OR2X1 U9600 ( .IN1(n9604), .IN2(n9605), .Q(g34615) );
  AND2X1 U9601 ( .IN1(n8829), .IN2(g2868), .Q(n9605) );
  AND2X1 U9602 ( .IN1(n8708), .IN2(g2873), .Q(n9604) );
  OR2X1 U9603 ( .IN1(n9606), .IN2(n9607), .Q(g34614) );
  AND2X1 U9604 ( .IN1(g37), .IN2(n8810), .Q(n9607) );
  AND2X1 U9605 ( .IN1(n8708), .IN2(g29214), .Q(n9606) );
  OR2X1 U9606 ( .IN1(n9608), .IN2(n9609), .Q(g34613) );
  AND2X1 U9607 ( .IN1(g37), .IN2(n8687), .Q(n9609) );
  AND2X1 U9608 ( .IN1(test_so95), .IN2(n8810), .Q(n9608) );
  OR2X1 U9609 ( .IN1(n9610), .IN2(n9611), .Q(g34612) );
  AND2X1 U9610 ( .IN1(n8829), .IN2(g2860), .Q(n9611) );
  AND2X1 U9611 ( .IN1(test_so95), .IN2(n8687), .Q(n9610) );
  OR2X1 U9612 ( .IN1(n9612), .IN2(n9613), .Q(g34611) );
  AND2X1 U9613 ( .IN1(n8829), .IN2(g2852), .Q(n9613) );
  AND2X1 U9614 ( .IN1(n8707), .IN2(g2860), .Q(n9612) );
  OR2X1 U9615 ( .IN1(n9614), .IN2(n9615), .Q(g34610) );
  AND2X1 U9616 ( .IN1(n8829), .IN2(g2844), .Q(n9615) );
  AND2X1 U9617 ( .IN1(n8707), .IN2(g2852), .Q(n9614) );
  OR2X1 U9618 ( .IN1(n9616), .IN2(n9617), .Q(g34609) );
  AND2X1 U9619 ( .IN1(n8829), .IN2(g2890), .Q(n9617) );
  AND2X1 U9620 ( .IN1(n8707), .IN2(g2844), .Q(n9616) );
  OR2X1 U9621 ( .IN1(n9618), .IN2(n9619), .Q(g34608) );
  AND2X1 U9622 ( .IN1(n8830), .IN2(g2697), .Q(n9619) );
  AND2X1 U9623 ( .IN1(n8708), .IN2(g2704), .Q(n9618) );
  OR2X1 U9624 ( .IN1(n9620), .IN2(n9621), .Q(g34607) );
  AND2X1 U9625 ( .IN1(n8830), .IN2(g2689), .Q(n9621) );
  AND2X1 U9626 ( .IN1(n8706), .IN2(g2697), .Q(n9620) );
  AND2X1 U9627 ( .IN1(n8706), .IN2(g2689), .Q(g34606) );
  OR2X1 U9628 ( .IN1(n9622), .IN2(n9623), .Q(g34605) );
  AND2X1 U9629 ( .IN1(n8830), .IN2(g2138), .Q(n9623) );
  AND2X1 U9630 ( .IN1(n8706), .IN2(g2145), .Q(n9622) );
  OR2X1 U9631 ( .IN1(n9624), .IN2(n9625), .Q(g34604) );
  AND2X1 U9632 ( .IN1(n8830), .IN2(g2130), .Q(n9625) );
  AND2X1 U9633 ( .IN1(n8707), .IN2(g2138), .Q(n9624) );
  AND2X1 U9634 ( .IN1(n8706), .IN2(g2130), .Q(g34603) );
  AND2X1 U9635 ( .IN1(n8706), .IN2(g1291), .Q(g34602) );
  AND2X1 U9636 ( .IN1(n8706), .IN2(g947), .Q(g34601) );
  OR3X1 U9637 ( .IN1(n9626), .IN2(n9627), .IN3(n9628), .Q(g34600) );
  AND2X1 U9638 ( .IN1(n8830), .IN2(g776), .Q(n9628) );
  AND2X1 U9639 ( .IN1(n2507), .IN2(n5551), .Q(n9627) );
  AND3X1 U9640 ( .IN1(n2404), .IN2(n9629), .IN3(g781), .Q(n9626) );
  INVX0 U9641 ( .INP(n2507), .ZN(n9629) );
  OR3X1 U9642 ( .IN1(n9630), .IN2(n9631), .IN3(n9632), .Q(g34599) );
  AND2X1 U9643 ( .IN1(n8830), .IN2(g608), .Q(n9632) );
  AND2X1 U9644 ( .IN1(n2509), .IN2(n5474), .Q(n9631) );
  AND3X1 U9645 ( .IN1(n2421), .IN2(n9633), .IN3(g613), .Q(n9630) );
  INVX0 U9646 ( .INP(n2509), .ZN(n9633) );
  OR2X1 U9647 ( .IN1(n9634), .IN2(n9635), .Q(g34598) );
  AND2X1 U9648 ( .IN1(g29221), .IN2(n8687), .Q(n9635) );
  AND2X1 U9649 ( .IN1(n8830), .IN2(g550), .Q(n9634) );
  OR2X1 U9650 ( .IN1(n9636), .IN2(n9637), .Q(g34468) );
  AND2X1 U9651 ( .IN1(n9638), .IN2(g4859), .Q(n9637) );
  AND2X1 U9652 ( .IN1(n9639), .IN2(g4854), .Q(n9636) );
  OR2X1 U9653 ( .IN1(n8805), .IN2(n9640), .Q(n9639) );
  AND2X1 U9654 ( .IN1(n9641), .IN2(n9642), .Q(n9640) );
  OR2X1 U9655 ( .IN1(n9643), .IN2(n9644), .Q(g34467) );
  AND2X1 U9656 ( .IN1(n8830), .IN2(g4849), .Q(n9644) );
  AND2X1 U9657 ( .IN1(n9645), .IN2(n9638), .Q(n9643) );
  XOR2X1 U9658 ( .IN1(n9642), .IN2(g4854), .Q(n9645) );
  AND2X1 U9659 ( .IN1(g4849), .IN2(n2563), .Q(n9642) );
  OR2X1 U9660 ( .IN1(n9646), .IN2(n9647), .Q(g34466) );
  AND3X1 U9661 ( .IN1(n9638), .IN2(g4843), .IN3(n5283), .Q(n9647) );
  AND2X1 U9662 ( .IN1(n9648), .IN2(g4878), .Q(n9646) );
  OR2X1 U9663 ( .IN1(n8805), .IN2(n9649), .Q(n9648) );
  AND2X1 U9664 ( .IN1(n8360), .IN2(n9641), .Q(n9649) );
  OR3X1 U9665 ( .IN1(n9650), .IN2(n9651), .IN3(n9652), .Q(g34465) );
  AND2X1 U9666 ( .IN1(n8830), .IN2(g4843), .Q(n9652) );
  AND2X1 U9667 ( .IN1(n2567), .IN2(n9638), .Q(n9651) );
  AND3X1 U9668 ( .IN1(n9641), .IN2(n2563), .IN3(n8436), .Q(n9650) );
  OR2X1 U9669 ( .IN1(n9653), .IN2(n9654), .Q(g34464) );
  AND2X1 U9670 ( .IN1(n9655), .IN2(g4669), .Q(n9654) );
  AND2X1 U9671 ( .IN1(n9656), .IN2(g4664), .Q(n9653) );
  OR2X1 U9672 ( .IN1(n8805), .IN2(n9657), .Q(n9656) );
  AND2X1 U9673 ( .IN1(n9658), .IN2(n9659), .Q(n9657) );
  OR2X1 U9674 ( .IN1(n9660), .IN2(n9661), .Q(g34463) );
  AND2X1 U9675 ( .IN1(n8830), .IN2(g4659), .Q(n9661) );
  AND2X1 U9676 ( .IN1(n9662), .IN2(n9655), .Q(n9660) );
  XOR2X1 U9677 ( .IN1(n9659), .IN2(g4664), .Q(n9662) );
  AND2X1 U9678 ( .IN1(g4659), .IN2(n2573), .Q(n9659) );
  OR2X1 U9679 ( .IN1(n9663), .IN2(n9664), .Q(g34462) );
  AND3X1 U9680 ( .IN1(n9655), .IN2(test_so19), .IN3(n5656), .Q(n9664) );
  AND2X1 U9681 ( .IN1(n9665), .IN2(g4688), .Q(n9663) );
  OR2X1 U9682 ( .IN1(n8805), .IN2(n9666), .Q(n9665) );
  AND2X1 U9683 ( .IN1(n9658), .IN2(n8522), .Q(n9666) );
  OR3X1 U9684 ( .IN1(n9667), .IN2(n9668), .IN3(n9669), .Q(g34461) );
  AND2X1 U9685 ( .IN1(test_so19), .IN2(n8810), .Q(n9669) );
  AND2X1 U9686 ( .IN1(n2577), .IN2(n9655), .Q(n9668) );
  AND3X1 U9687 ( .IN1(n9658), .IN2(n2573), .IN3(n8439), .Q(n9667) );
  OR2X1 U9688 ( .IN1(n9670), .IN2(n9671), .Q(g34460) );
  AND2X1 U9689 ( .IN1(g34025), .IN2(test_so3), .Q(n9671) );
  AND2X1 U9690 ( .IN1(n9672), .IN2(g4639), .Q(n9670) );
  OR2X1 U9691 ( .IN1(n8805), .IN2(n9673), .Q(n9672) );
  AND3X1 U9692 ( .IN1(n9674), .IN2(n8510), .IN3(n5382), .Q(n9673) );
  OR2X1 U9693 ( .IN1(n9675), .IN2(n9676), .Q(g34459) );
  AND2X1 U9694 ( .IN1(n9677), .IN2(n8687), .Q(n9676) );
  OR2X1 U9695 ( .IN1(n9678), .IN2(n9679), .Q(n9677) );
  INVX0 U9696 ( .INP(n9674), .ZN(n9679) );
  AND2X1 U9697 ( .IN1(n9680), .IN2(n9681), .Q(n9678) );
  OR2X1 U9698 ( .IN1(n9682), .IN2(g4340), .Q(n9680) );
  AND2X1 U9699 ( .IN1(n8830), .IN2(g4643), .Q(n9675) );
  OR2X1 U9700 ( .IN1(n9683), .IN2(n9684), .Q(g34458) );
  AND2X1 U9701 ( .IN1(test_so99), .IN2(n9685), .Q(n9684) );
  OR2X1 U9702 ( .IN1(n8805), .IN2(n9686), .Q(n9685) );
  AND3X1 U9703 ( .IN1(n9687), .IN2(g4639), .IN3(n5844), .Q(n9686) );
  AND2X1 U9704 ( .IN1(n9688), .IN2(g4633), .Q(n9683) );
  OR2X1 U9705 ( .IN1(n9689), .IN2(n9690), .Q(n9688) );
  AND2X1 U9706 ( .IN1(n9691), .IN2(n8511), .Q(n9689) );
  OR3X1 U9707 ( .IN1(n9692), .IN2(n9693), .IN3(n9694), .Q(g34457) );
  AND2X1 U9708 ( .IN1(test_so3), .IN2(n8810), .Q(n9694) );
  AND3X1 U9709 ( .IN1(n9687), .IN2(g4639), .IN3(n8511), .Q(n9693) );
  AND2X1 U9710 ( .IN1(test_so99), .IN2(n9690), .Q(n9692) );
  OR2X1 U9711 ( .IN1(n9695), .IN2(g34025), .Q(n9690) );
  AND2X1 U9712 ( .IN1(n9691), .IN2(n8510), .Q(n9695) );
  OR2X1 U9713 ( .IN1(n9696), .IN2(n9697), .Q(g34456) );
  AND2X1 U9714 ( .IN1(n9698), .IN2(g4616), .Q(n9697) );
  AND2X1 U9715 ( .IN1(n9699), .IN2(g4608), .Q(n9696) );
  OR2X1 U9716 ( .IN1(n8805), .IN2(n9700), .Q(n9699) );
  AND2X1 U9717 ( .IN1(n2590), .IN2(n9701), .Q(n9700) );
  OR2X1 U9718 ( .IN1(n9702), .IN2(n9703), .Q(g34455) );
  AND2X1 U9719 ( .IN1(n2595), .IN2(g4332), .Q(n9703) );
  AND2X1 U9720 ( .IN1(n9704), .IN2(g4322), .Q(n9702) );
  OR2X1 U9721 ( .IN1(n8805), .IN2(n9705), .Q(n9704) );
  AND3X1 U9722 ( .IN1(n9674), .IN2(n9706), .IN3(n2594), .Q(n9705) );
  OR2X1 U9723 ( .IN1(n9707), .IN2(n9708), .Q(g34454) );
  AND2X1 U9724 ( .IN1(n8830), .IN2(g4601), .Q(n9708) );
  AND2X1 U9725 ( .IN1(n9709), .IN2(n9698), .Q(n9707) );
  XOR2X1 U9726 ( .IN1(n2590), .IN2(g4608), .Q(n9709) );
  OR3X1 U9727 ( .IN1(n9710), .IN2(n9711), .IN3(n9712), .Q(g34453) );
  AND2X1 U9728 ( .IN1(n8830), .IN2(g4593), .Q(n9712) );
  AND3X1 U9729 ( .IN1(n2598), .IN2(n9701), .IN3(n5365), .Q(n9711) );
  AND3X1 U9730 ( .IN1(n9698), .IN2(n9713), .IN3(g4601), .Q(n9710) );
  INVX0 U9731 ( .INP(n2598), .ZN(n9713) );
  OR2X1 U9732 ( .IN1(n9714), .IN2(n9715), .Q(g34452) );
  AND2X1 U9733 ( .IN1(n8830), .IN2(g4584), .Q(n9715) );
  AND2X1 U9734 ( .IN1(n9716), .IN2(n9698), .Q(n9714) );
  XOR2X1 U9735 ( .IN1(g4593), .IN2(n2601), .Q(n9716) );
  OR2X1 U9736 ( .IN1(n9717), .IN2(n9718), .Q(g34451) );
  AND2X1 U9737 ( .IN1(n8830), .IN2(g4332), .Q(n9718) );
  AND2X1 U9738 ( .IN1(n9719), .IN2(n9698), .Q(n9717) );
  AND2X1 U9739 ( .IN1(n8706), .IN2(n9701), .Q(n9698) );
  AND2X1 U9740 ( .IN1(n9674), .IN2(n9720), .Q(n9701) );
  INVX0 U9741 ( .INP(n9721), .ZN(n9720) );
  AND2X1 U9742 ( .IN1(n2601), .IN2(g4616), .Q(n9721) );
  AND2X1 U9743 ( .IN1(g4584), .IN2(n9722), .Q(n2601) );
  XOR2X1 U9744 ( .IN1(g4584), .IN2(n9722), .Q(n9719) );
  OR3X1 U9745 ( .IN1(n9723), .IN2(n9724), .IN3(n9725), .Q(g34450) );
  AND2X1 U9746 ( .IN1(n8830), .IN2(g4311), .Q(n9725) );
  AND3X1 U9747 ( .IN1(n2594), .IN2(n9674), .IN3(n5506), .Q(n9724) );
  AND3X1 U9748 ( .IN1(n2595), .IN2(n9726), .IN3(g4322), .Q(n9723) );
  INVX0 U9749 ( .INP(n2594), .ZN(n9726) );
  AND2X1 U9750 ( .IN1(n9706), .IN2(n9727), .Q(n2595) );
  INVX0 U9751 ( .INP(n9722), .ZN(n9706) );
  AND3X1 U9752 ( .IN1(g4332), .IN2(g4322), .IN3(n2607), .Q(n9722) );
  AND2X1 U9753 ( .IN1(g4358), .IN2(n9728), .Q(n2607) );
  OR3X1 U9754 ( .IN1(n9729), .IN2(n9730), .IN3(n9731), .Q(g34448) );
  AND3X1 U9755 ( .IN1(n9732), .IN2(n9733), .IN3(n9734), .Q(n9731) );
  OR2X1 U9756 ( .IN1(n9735), .IN2(n9736), .Q(n9732) );
  AND2X1 U9757 ( .IN1(n7969), .IN2(n8686), .Q(n9735) );
  AND2X1 U9758 ( .IN1(n8830), .IN2(g2827), .Q(n9730) );
  AND3X1 U9759 ( .IN1(n9737), .IN2(g2819), .IN3(n8731), .Q(n9729) );
  OR3X1 U9760 ( .IN1(n9738), .IN2(n9739), .IN3(n9740), .Q(g34447) );
  AND3X1 U9761 ( .IN1(n9741), .IN2(n9733), .IN3(n9742), .Q(n9740) );
  OR2X1 U9762 ( .IN1(n9743), .IN2(n9736), .Q(n9741) );
  AND2X1 U9763 ( .IN1(n7968), .IN2(n8686), .Q(n9743) );
  AND2X1 U9764 ( .IN1(n8830), .IN2(g2815), .Q(n9739) );
  AND3X1 U9765 ( .IN1(n9744), .IN2(g2807), .IN3(n8732), .Q(n9738) );
  OR3X1 U9766 ( .IN1(n9745), .IN2(n9746), .IN3(n9747), .Q(g34446) );
  AND3X1 U9767 ( .IN1(n9748), .IN2(n9733), .IN3(n9749), .Q(n9747) );
  INVX0 U9768 ( .INP(n9750), .ZN(n9748) );
  AND2X1 U9769 ( .IN1(n9751), .IN2(n9752), .Q(n9750) );
  OR2X1 U9770 ( .IN1(n8806), .IN2(test_so37), .Q(n9751) );
  AND2X1 U9771 ( .IN1(n8830), .IN2(g2819), .Q(n9746) );
  AND3X1 U9772 ( .IN1(n9753), .IN2(g2815), .IN3(n8731), .Q(n9745) );
  OR3X1 U9773 ( .IN1(n9754), .IN2(n9755), .IN3(n9756), .Q(g34445) );
  AND3X1 U9774 ( .IN1(n9757), .IN2(n9733), .IN3(n9758), .Q(n9756) );
  OR2X1 U9775 ( .IN1(n1697), .IN2(n6005), .Q(n9733) );
  OR2X1 U9776 ( .IN1(n9759), .IN2(n9736), .Q(n9757) );
  AND2X1 U9777 ( .IN1(n7965), .IN2(n8687), .Q(n9759) );
  AND2X1 U9778 ( .IN1(n8830), .IN2(g2807), .Q(n9755) );
  AND3X1 U9779 ( .IN1(n9760), .IN2(g2803), .IN3(n8731), .Q(n9754) );
  OR3X1 U9780 ( .IN1(n9761), .IN2(n9762), .IN3(n9763), .Q(g34444) );
  AND3X1 U9781 ( .IN1(n9764), .IN2(n9765), .IN3(n9734), .Q(n9763) );
  INVX0 U9782 ( .INP(n9737), .ZN(n9734) );
  OR2X1 U9783 ( .IN1(n9766), .IN2(n9736), .Q(n9764) );
  AND2X1 U9784 ( .IN1(n7966), .IN2(n8686), .Q(n9766) );
  AND2X1 U9785 ( .IN1(n8830), .IN2(g2795), .Q(n9762) );
  AND3X1 U9786 ( .IN1(n9737), .IN2(g2787), .IN3(n8731), .Q(n9761) );
  OR2X1 U9787 ( .IN1(n9767), .IN2(n9768), .Q(n9737) );
  OR3X1 U9788 ( .IN1(n9769), .IN2(n9770), .IN3(n9771), .Q(g34443) );
  AND3X1 U9789 ( .IN1(n9772), .IN2(n9765), .IN3(n9742), .Q(n9771) );
  OR2X1 U9790 ( .IN1(n9773), .IN2(n9736), .Q(n9772) );
  AND2X1 U9791 ( .IN1(n7964), .IN2(n8686), .Q(n9773) );
  AND2X1 U9792 ( .IN1(n8830), .IN2(g2783), .Q(n9770) );
  AND3X1 U9793 ( .IN1(n9744), .IN2(g2775), .IN3(n8731), .Q(n9769) );
  INVX0 U9794 ( .INP(n9742), .ZN(n9744) );
  AND3X1 U9795 ( .IN1(g2724), .IN2(n8347), .IN3(n9774), .Q(n9742) );
  OR3X1 U9796 ( .IN1(n9775), .IN2(n9776), .IN3(n9777), .Q(g34442) );
  AND3X1 U9797 ( .IN1(n9778), .IN2(n9765), .IN3(n9749), .Q(n9777) );
  INVX0 U9798 ( .INP(n9753), .ZN(n9749) );
  OR2X1 U9799 ( .IN1(n9779), .IN2(n9736), .Q(n9778) );
  AND2X1 U9800 ( .IN1(n7967), .IN2(n8686), .Q(n9779) );
  AND2X1 U9801 ( .IN1(n8831), .IN2(g2787), .Q(n9776) );
  AND3X1 U9802 ( .IN1(n9753), .IN2(g2783), .IN3(n8732), .Q(n9775) );
  OR2X1 U9803 ( .IN1(n9768), .IN2(n9780), .Q(n9753) );
  OR3X1 U9804 ( .IN1(n9781), .IN2(n9782), .IN3(n9783), .Q(g34441) );
  AND3X1 U9805 ( .IN1(n9784), .IN2(n9765), .IN3(n9758), .Q(n9783) );
  OR2X1 U9806 ( .IN1(n1697), .IN2(n6006), .Q(n9765) );
  OR2X1 U9807 ( .IN1(n9785), .IN2(n9736), .Q(n9784) );
  AND2X1 U9808 ( .IN1(n7970), .IN2(n8686), .Q(n9785) );
  AND2X1 U9809 ( .IN1(n8831), .IN2(g2775), .Q(n9782) );
  AND3X1 U9810 ( .IN1(n9760), .IN2(g2771), .IN3(n8731), .Q(n9781) );
  INVX0 U9811 ( .INP(n9758), .ZN(n9760) );
  AND2X1 U9812 ( .IN1(n9786), .IN2(n9774), .Q(n9758) );
  OR2X1 U9813 ( .IN1(n9787), .IN2(n9788), .Q(g34440) );
  AND2X1 U9814 ( .IN1(n9789), .IN2(n8686), .Q(n9788) );
  OR2X1 U9815 ( .IN1(n9790), .IN2(n9791), .Q(n9789) );
  AND2X1 U9816 ( .IN1(g890), .IN2(g896), .Q(n9791) );
  AND2X1 U9817 ( .IN1(n9792), .IN2(g862), .Q(n9790) );
  OR2X1 U9818 ( .IN1(n9793), .IN2(n5431), .Q(n9792) );
  AND2X1 U9819 ( .IN1(n9794), .IN2(n9795), .Q(n9793) );
  OR3X1 U9820 ( .IN1(n2644), .IN2(n9796), .IN3(g703), .Q(n9794) );
  AND2X1 U9821 ( .IN1(n8831), .IN2(g446), .Q(n9787) );
  OR3X1 U9822 ( .IN1(n9797), .IN2(n9798), .IN3(n9799), .Q(g34439) );
  AND2X1 U9823 ( .IN1(n8831), .IN2(g772), .Q(n9799) );
  AND2X1 U9824 ( .IN1(n2554), .IN2(n5330), .Q(n9798) );
  AND3X1 U9826 ( .IN1(n2404), .IN2(n9800), .IN3(g776), .Q(n9797) );
  INVX0 U9827 ( .INP(n2554), .ZN(n9800) );
  OR3X1 U9828 ( .IN1(n9801), .IN2(n9802), .IN3(n9803), .Q(g34438) );
  AND2X1 U9829 ( .IN1(n8831), .IN2(g604), .Q(n9803) );
  AND2X1 U9830 ( .IN1(n2556), .IN2(n5475), .Q(n9802) );
  AND3X1 U9831 ( .IN1(n2421), .IN2(n9804), .IN3(g608), .Q(n9801) );
  INVX0 U9832 ( .INP(n2556), .ZN(n9804) );
  AND4X1 U9833 ( .IN1(n8226), .IN2(n5711), .IN3(n5416), .IN4(n9805), .Q(g34435) );
  OR3X1 U9834 ( .IN1(n9806), .IN2(g4141), .IN3(g4082), .Q(n9805) );
  AND4X1 U9835 ( .IN1(test_so11), .IN2(n5350), .IN3(n9807), .IN4(g4112), .Q(
        n9806) );
  OR2X1 U9836 ( .IN1(n8476), .IN2(n9094), .Q(g34425) );
  OR2X1 U9837 ( .IN1(n9808), .IN2(n9809), .Q(n9094) );
  AND2X1 U9838 ( .IN1(n9810), .IN2(n9811), .Q(n9808) );
  OR2X1 U9839 ( .IN1(n9812), .IN2(n9813), .Q(n8476) );
  AND2X1 U9840 ( .IN1(n9814), .IN2(test_so81), .Q(n9813) );
  OR2X1 U9841 ( .IN1(n9815), .IN2(n9816), .Q(n9814) );
  AND2X1 U9842 ( .IN1(n9817), .IN2(g4358), .Q(n9816) );
  OR2X1 U9843 ( .IN1(n9818), .IN2(n9819), .Q(n9817) );
  AND2X1 U9844 ( .IN1(n9820), .IN2(n9509), .Q(n9819) );
  AND2X1 U9845 ( .IN1(n9821), .IN2(n9512), .Q(n9818) );
  AND2X1 U9846 ( .IN1(n5348), .IN2(n9822), .Q(n9815) );
  OR2X1 U9847 ( .IN1(n9823), .IN2(n9824), .Q(n9822) );
  AND2X1 U9848 ( .IN1(n9825), .IN2(n9509), .Q(n9824) );
  AND2X1 U9849 ( .IN1(n9826), .IN2(n9512), .Q(n9823) );
  AND2X1 U9850 ( .IN1(n9827), .IN2(n8492), .Q(n9812) );
  OR2X1 U9851 ( .IN1(n9828), .IN2(n9829), .Q(n9827) );
  AND2X1 U9852 ( .IN1(n9830), .IN2(g4358), .Q(n9829) );
  OR2X1 U9853 ( .IN1(n9831), .IN2(n9832), .Q(n9830) );
  AND2X1 U9854 ( .IN1(n9833), .IN2(n9509), .Q(n9832) );
  AND2X1 U9855 ( .IN1(n9834), .IN2(n9512), .Q(n9831) );
  AND2X1 U9856 ( .IN1(n5348), .IN2(n9835), .Q(n9828) );
  OR2X1 U9857 ( .IN1(n9836), .IN2(n9837), .Q(n9835) );
  AND2X1 U9858 ( .IN1(n9003), .IN2(n9509), .Q(n9837) );
  INVX0 U9859 ( .INP(n9810), .ZN(n9509) );
  AND2X1 U9860 ( .IN1(g31860), .IN2(n9512), .Q(n9836) );
  INVX0 U9861 ( .INP(n9811), .ZN(n9512) );
  OR3X1 U9862 ( .IN1(g34843), .IN2(n9838), .IN3(n9809), .Q(g34383) );
  AND2X1 U9863 ( .IN1(n9839), .IN2(n9840), .Q(n9838) );
  AND4X1 U9864 ( .IN1(n9841), .IN2(n9842), .IN3(n9843), .IN4(n9844), .Q(n9840)
         );
  AND4X1 U9865 ( .IN1(n915), .IN2(n928), .IN3(n927), .IN4(n917), .Q(n9839) );
  OR2X1 U9866 ( .IN1(n9845), .IN2(n9846), .Q(g34843) );
  OR4X1 U9867 ( .IN1(n9847), .IN2(n9848), .IN3(n9849), .IN4(n9850), .Q(n9846)
         );
  AND3X1 U9868 ( .IN1(n9851), .IN2(g2495), .IN3(n5523), .Q(n9850) );
  AND3X1 U9869 ( .IN1(n9852), .IN2(g2629), .IN3(n5524), .Q(n9849) );
  AND2X1 U9870 ( .IN1(g31862), .IN2(n9853), .Q(n9848) );
  AND3X1 U9871 ( .IN1(n5505), .IN2(g2070), .IN3(n9854), .Q(n9847) );
  OR4X1 U9872 ( .IN1(n9855), .IN2(n9856), .IN3(n9857), .IN4(n9858), .Q(n9845)
         );
  INVX0 U9873 ( .INP(n9859), .ZN(n9858) );
  INVX0 U9874 ( .INP(n9860), .ZN(n9857) );
  OR3X1 U9875 ( .IN1(n9861), .IN2(n9862), .IN3(n9863), .Q(g34269) );
  AND3X1 U9876 ( .IN1(n9864), .IN2(n9865), .IN3(n9866), .Q(n9863) );
  OR2X1 U9877 ( .IN1(n9867), .IN2(g4961), .Q(n9865) );
  AND2X1 U9878 ( .IN1(n8831), .IN2(g4961), .Q(n9862) );
  AND3X1 U9879 ( .IN1(n9868), .IN2(g4955), .IN3(n8731), .Q(n9861) );
  INVX0 U9880 ( .INP(n9864), .ZN(n9868) );
  OR2X1 U9881 ( .IN1(n9869), .IN2(n9870), .Q(n9864) );
  OR3X1 U9882 ( .IN1(n9871), .IN2(n9872), .IN3(n9873), .Q(g34268) );
  AND3X1 U9883 ( .IN1(n9874), .IN2(n9875), .IN3(n9866), .Q(n9873) );
  OR2X1 U9884 ( .IN1(n9867), .IN2(g4950), .Q(n9875) );
  AND2X1 U9885 ( .IN1(n8831), .IN2(g4950), .Q(n9872) );
  AND3X1 U9887 ( .IN1(n9876), .IN2(g4944), .IN3(n8731), .Q(n9871) );
  INVX0 U9888 ( .INP(n9874), .ZN(n9876) );
  OR2X1 U9889 ( .IN1(n9877), .IN2(n9870), .Q(n9874) );
  OR3X1 U9890 ( .IN1(n9878), .IN2(n9879), .IN3(n9880), .Q(g34267) );
  AND3X1 U9891 ( .IN1(n9881), .IN2(n9882), .IN3(n9866), .Q(n9880) );
  OR2X1 U9892 ( .IN1(n9867), .IN2(g4939), .Q(n9882) );
  AND2X1 U9893 ( .IN1(n8831), .IN2(g4939), .Q(n9879) );
  AND3X1 U9894 ( .IN1(n9883), .IN2(g4933), .IN3(n8731), .Q(n9878) );
  INVX0 U9895 ( .INP(n9881), .ZN(n9883) );
  OR2X1 U9896 ( .IN1(n9884), .IN2(n9870), .Q(n9881) );
  OR3X1 U9897 ( .IN1(n9885), .IN2(n9886), .IN3(n9887), .Q(g34266) );
  AND3X1 U9898 ( .IN1(n9888), .IN2(n9889), .IN3(n9866), .Q(n9887) );
  AND2X1 U9899 ( .IN1(n8705), .IN2(n9890), .Q(n9866) );
  OR2X1 U9900 ( .IN1(n9891), .IN2(n9867), .Q(n9890) );
  OR2X1 U9901 ( .IN1(n9867), .IN2(g4894), .Q(n9889) );
  INVX0 U9902 ( .INP(n9892), .ZN(n9867) );
  OR2X1 U9903 ( .IN1(n8289), .IN2(n9891), .Q(n9892) );
  AND2X1 U9904 ( .IN1(n8831), .IN2(g4894), .Q(n9886) );
  AND3X1 U9905 ( .IN1(n9893), .IN2(g4888), .IN3(n8730), .Q(n9885) );
  INVX0 U9906 ( .INP(n9888), .ZN(n9893) );
  OR2X1 U9907 ( .IN1(n9508), .IN2(n9870), .Q(n9888) );
  INVX0 U9908 ( .INP(n9891), .ZN(n9870) );
  OR3X1 U9909 ( .IN1(test_so46), .IN2(n9894), .IN3(g5008), .Q(n9891) );
  AND2X1 U9910 ( .IN1(n9638), .IN2(n9055), .Q(g34265) );
  AND3X1 U9911 ( .IN1(n5318), .IN2(n5443), .IN3(n5713), .Q(n9055) );
  AND2X1 U9912 ( .IN1(n8705), .IN2(n9641), .Q(n9638) );
  AND2X1 U9913 ( .IN1(n9895), .IN2(n9896), .Q(n9641) );
  INVX0 U9914 ( .INP(n9510), .ZN(n9895) );
  OR3X1 U9915 ( .IN1(n9897), .IN2(n9898), .IN3(n9899), .Q(g34264) );
  AND3X1 U9916 ( .IN1(n9900), .IN2(n9901), .IN3(n9902), .Q(n9899) );
  OR2X1 U9917 ( .IN1(n9903), .IN2(g4771), .Q(n9901) );
  AND2X1 U9918 ( .IN1(n8831), .IN2(g4771), .Q(n9898) );
  AND3X1 U9919 ( .IN1(n9904), .IN2(g4765), .IN3(n8730), .Q(n9897) );
  INVX0 U9920 ( .INP(n9900), .ZN(n9904) );
  OR2X1 U9921 ( .IN1(n9905), .IN2(n9906), .Q(n9900) );
  OR3X1 U9922 ( .IN1(n9907), .IN2(n9908), .IN3(n9909), .Q(g34263) );
  AND3X1 U9923 ( .IN1(n9910), .IN2(n9911), .IN3(n9902), .Q(n9909) );
  OR2X1 U9924 ( .IN1(n9903), .IN2(g4760), .Q(n9911) );
  AND2X1 U9925 ( .IN1(n8831), .IN2(g4760), .Q(n9908) );
  AND3X1 U9926 ( .IN1(n9912), .IN2(g4754), .IN3(n8732), .Q(n9907) );
  INVX0 U9928 ( .INP(n9910), .ZN(n9912) );
  OR2X1 U9929 ( .IN1(n9913), .IN2(n9906), .Q(n9910) );
  OR3X1 U9930 ( .IN1(n9914), .IN2(n9915), .IN3(n9916), .Q(g34262) );
  AND3X1 U9931 ( .IN1(n9917), .IN2(n9918), .IN3(n9902), .Q(n9916) );
  OR2X1 U9932 ( .IN1(n9903), .IN2(test_so18), .Q(n9918) );
  AND2X1 U9933 ( .IN1(test_so18), .IN2(n8810), .Q(n9915) );
  AND3X1 U9934 ( .IN1(n9919), .IN2(g4743), .IN3(n8730), .Q(n9914) );
  INVX0 U9935 ( .INP(n9917), .ZN(n9919) );
  OR2X1 U9936 ( .IN1(n9920), .IN2(n9906), .Q(n9917) );
  OR3X1 U9937 ( .IN1(n9921), .IN2(n9922), .IN3(n9923), .Q(g34261) );
  AND3X1 U9938 ( .IN1(n9924), .IN2(n9925), .IN3(n9902), .Q(n9923) );
  AND2X1 U9939 ( .IN1(n8705), .IN2(n9926), .Q(n9902) );
  OR2X1 U9940 ( .IN1(n9927), .IN2(n9903), .Q(n9926) );
  OR2X1 U9941 ( .IN1(n9903), .IN2(g4704), .Q(n9925) );
  INVX0 U9942 ( .INP(n9928), .ZN(n9903) );
  OR2X1 U9943 ( .IN1(n8290), .IN2(n9927), .Q(n9928) );
  AND2X1 U9944 ( .IN1(n8831), .IN2(g4704), .Q(n9922) );
  AND3X1 U9945 ( .IN1(n9929), .IN2(g4698), .IN3(n8748), .Q(n9921) );
  INVX0 U9946 ( .INP(n9924), .ZN(n9929) );
  OR2X1 U9947 ( .IN1(n9511), .IN2(n9906), .Q(n9924) );
  INVX0 U9948 ( .INP(n9927), .ZN(n9906) );
  OR3X1 U9949 ( .IN1(n9894), .IN2(g4818), .IN3(g8132), .Q(n9927) );
  AND2X1 U9950 ( .IN1(n9655), .IN2(n9029), .Q(g34260) );
  AND3X1 U9951 ( .IN1(n5440), .IN2(n5712), .IN3(n8224), .Q(n9029) );
  AND2X1 U9952 ( .IN1(n8706), .IN2(n9658), .Q(n9655) );
  AND2X1 U9954 ( .IN1(n9930), .IN2(n9931), .Q(n9658) );
  AND2X1 U9955 ( .IN1(n9932), .IN2(g4633), .Q(g34259) );
  OR2X1 U9956 ( .IN1(n8794), .IN2(n9933), .Q(n9932) );
  AND2X1 U9959 ( .IN1(n9687), .IN2(n5727), .Q(n9933) );
  AND3X1 U9960 ( .IN1(n9674), .IN2(test_so3), .IN3(n5382), .Q(n9687) );
  OR3X1 U9961 ( .IN1(n9934), .IN2(n9935), .IN3(n9936), .Q(g34258) );
  AND2X1 U9962 ( .IN1(test_so81), .IN2(n8810), .Q(n9936) );
  AND3X1 U9963 ( .IN1(n9728), .IN2(n9674), .IN3(n5348), .Q(n9935) );
  INVX0 U9964 ( .INP(n9937), .ZN(n9728) );
  AND3X1 U9965 ( .IN1(n9727), .IN2(n9937), .IN3(g4358), .Q(n9934) );
  OR2X1 U9966 ( .IN1(n8492), .IN2(n9681), .Q(n9937) );
  OR3X1 U9967 ( .IN1(n9938), .IN2(n9939), .IN3(n9940), .Q(g34257) );
  AND2X1 U9969 ( .IN1(n8831), .IN2(g4340), .Q(n9940) );
  AND3X1 U9970 ( .IN1(n9674), .IN2(n8492), .IN3(n9941), .Q(n9939) );
  AND3X1 U9971 ( .IN1(n9727), .IN2(test_so81), .IN3(n9681), .Q(n9938) );
  INVX0 U9973 ( .INP(n9941), .ZN(n9681) );
  AND2X1 U9974 ( .IN1(g4340), .IN2(n9682), .Q(n9941) );
  AND3X1 U9975 ( .IN1(n5727), .IN2(test_so3), .IN3(test_so99), .Q(n9682) );
  OR2X1 U9976 ( .IN1(n9942), .IN2(n9943), .Q(g34256) );
  AND2X1 U9977 ( .IN1(n9944), .IN2(n8685), .Q(n9943) );
  OR3X1 U9978 ( .IN1(n9945), .IN2(n9946), .IN3(g4459), .Q(n9944) );
  AND2X1 U9979 ( .IN1(n5671), .IN2(g4473), .Q(n9946) );
  AND2X1 U9980 ( .IN1(n8831), .IN2(g4369), .Q(n9942) );
  OR4X1 U9981 ( .IN1(n9947), .IN2(g4462), .IN3(n8792), .IN4(n9945), .Q(g34255)
         );
  AND2X1 U9982 ( .IN1(test_so38), .IN2(g4473), .Q(n9947) );
  OR2X1 U9983 ( .IN1(n9948), .IN2(n9949), .Q(g34254) );
  AND2X1 U9984 ( .IN1(n9945), .IN2(n8685), .Q(n9949) );
  AND2X1 U9985 ( .IN1(n9950), .IN2(g4473), .Q(n9948) );
  OR4X1 U9986 ( .IN1(n5382), .IN2(n8792), .IN3(test_so38), .IN4(n5671), .Q(
        n9950) );
  AND2X1 U9987 ( .IN1(n9951), .IN2(n8685), .Q(g34253) );
  OR3X1 U9988 ( .IN1(n5671), .IN2(n9945), .IN3(n8506), .Q(n9951) );
  AND3X1 U9989 ( .IN1(g26960), .IN2(n9952), .IN3(n5849), .Q(n9945) );
  OR2X1 U9990 ( .IN1(n9397), .IN2(n9953), .Q(n9952) );
  AND2X1 U9991 ( .IN1(n2668), .IN2(n5846), .Q(n9953) );
  OR3X1 U9993 ( .IN1(n9954), .IN2(n9955), .IN3(n9956), .Q(g34252) );
  AND2X1 U9994 ( .IN1(n8831), .IN2(g767), .Q(n9956) );
  AND2X1 U9995 ( .IN1(n2647), .IN2(n5334), .Q(n9955) );
  AND3X1 U9996 ( .IN1(n2404), .IN2(n9957), .IN3(g772), .Q(n9954) );
  INVX0 U9997 ( .INP(n2647), .ZN(n9957) );
  OR3X1 U9998 ( .IN1(n9958), .IN2(n9959), .IN3(n9960), .Q(g34251) );
  AND2X1 U9999 ( .IN1(n8831), .IN2(g599), .Q(n9960) );
  AND2X1 U10000 ( .IN1(n2649), .IN2(n5473), .Q(n9959) );
  AND3X1 U10001 ( .IN1(n2421), .IN2(n9961), .IN3(g604), .Q(n9958) );
  INVX0 U10002 ( .INP(n2649), .ZN(n9961) );
  OR3X1 U10003 ( .IN1(n9962), .IN2(n9963), .IN3(n9964), .Q(g34250) );
  AND2X1 U10004 ( .IN1(n8831), .IN2(g298), .Q(n9964) );
  AND2X1 U10005 ( .IN1(n5724), .IN2(n2707), .Q(n9963) );
  AND3X1 U10006 ( .IN1(n8473), .IN2(n9965), .IN3(g142), .Q(n9962) );
  INVX0 U10007 ( .INP(n2707), .ZN(n9965) );
  OR3X1 U10008 ( .IN1(n9966), .IN2(n9967), .IN3(n9968), .Q(g34249) );
  AND2X1 U10009 ( .IN1(n8831), .IN2(g157), .Q(n9968) );
  AND2X1 U10010 ( .IN1(n2710), .IN2(n5843), .Q(n9967) );
  AND3X1 U10011 ( .IN1(n9969), .IN2(n9970), .IN3(g160), .Q(n9966) );
  INVX0 U10012 ( .INP(n2710), .ZN(n9970) );
  OR3X1 U10013 ( .IN1(g34781), .IN2(n9971), .IN3(n9809), .Q(g34201) );
  AND4X1 U10014 ( .IN1(n724), .IN2(n1635), .IN3(n9972), .IN4(n9973), .Q(n9971)
         );
  AND4X1 U10015 ( .IN1(n1282), .IN2(n1284), .IN3(n1278), .IN4(n1280), .Q(n9973) );
  AND2X1 U10016 ( .IN1(n729), .IN2(n727), .Q(n9972) );
  OR4X1 U10017 ( .IN1(n9974), .IN2(n9975), .IN3(n9976), .IN4(n9977), .Q(g34781) );
  OR4X1 U10018 ( .IN1(n9978), .IN2(n9979), .IN3(n9980), .IN4(n9981), .Q(n9977)
         );
  AND2X1 U10019 ( .IN1(n9982), .IN2(n9983), .Q(n9981) );
  AND2X1 U10020 ( .IN1(n9984), .IN2(n3005), .Q(n9980) );
  AND2X1 U10021 ( .IN1(n9985), .IN2(n9986), .Q(n9979) );
  AND2X1 U10022 ( .IN1(n9987), .IN2(n9988), .Q(n9978) );
  OR2X1 U10023 ( .IN1(n9989), .IN2(n9990), .Q(n9976) );
  AND2X1 U10024 ( .IN1(n9991), .IN2(n9992), .Q(n9990) );
  AND2X1 U10025 ( .IN1(n9993), .IN2(n9994), .Q(n9989) );
  AND2X1 U10026 ( .IN1(g31863), .IN2(n9995), .Q(n9975) );
  AND2X1 U10027 ( .IN1(n9996), .IN2(n9997), .Q(n9974) );
  OR2X1 U10028 ( .IN1(n9998), .IN2(n9999), .Q(g34041) );
  AND2X1 U10029 ( .IN1(n8831), .IN2(g5008), .Q(n9999) );
  AND2X1 U10030 ( .IN1(n10000), .IN2(n10001), .Q(n9998) );
  XOR2X1 U10031 ( .IN1(n9510), .IN2(g4983), .Q(n10000) );
  OR4X1 U10032 ( .IN1(n10002), .IN2(n10003), .IN3(n10004), .IN4(n10005), .Q(
        g34040) );
  AND3X1 U10033 ( .IN1(n9065), .IN2(n9896), .IN3(n8752), .Q(n10005) );
  AND2X1 U10034 ( .IN1(n8831), .IN2(g4975), .Q(n10004) );
  AND2X1 U10035 ( .IN1(n10001), .IN2(g4899), .Q(n10003) );
  AND2X1 U10036 ( .IN1(n10006), .IN2(n9064), .Q(n10002) );
  OR2X1 U10037 ( .IN1(n10007), .IN2(n10008), .Q(g34039) );
  AND2X1 U10038 ( .IN1(n10001), .IN2(g4966), .Q(n10008) );
  AND2X1 U10039 ( .IN1(test_so58), .IN2(n10009), .Q(n10007) );
  OR2X1 U10040 ( .IN1(n8795), .IN2(n10010), .Q(n10009) );
  AND2X1 U10041 ( .IN1(n10011), .IN2(n10012), .Q(n10010) );
  OR3X1 U10042 ( .IN1(n10013), .IN2(n10014), .IN3(n10015), .Q(g34038) );
  AND2X1 U10043 ( .IN1(n8831), .IN2(g4983), .Q(n10015) );
  AND3X1 U10044 ( .IN1(n10011), .IN2(n8505), .IN3(n10012), .Q(n10014) );
  AND3X1 U10045 ( .IN1(test_so58), .IN2(n10001), .IN3(n10016), .Q(n10013) );
  OR3X1 U10046 ( .IN1(n10017), .IN2(n10018), .IN3(n10019), .Q(g34037) );
  AND2X1 U10047 ( .IN1(n8824), .IN2(g4966), .Q(n10019) );
  AND2X1 U10048 ( .IN1(n10006), .IN2(n5360), .Q(n10018) );
  AND3X1 U10049 ( .IN1(g4966), .IN2(n9896), .IN3(n10012), .Q(n10006) );
  AND2X1 U10050 ( .IN1(n10001), .IN2(g4975), .Q(n10017) );
  AND2X1 U10051 ( .IN1(n8705), .IN2(n10011), .Q(n10001) );
  AND2X1 U10052 ( .IN1(n9896), .IN2(n10020), .Q(n10011) );
  OR2X1 U10053 ( .IN1(n10016), .IN2(n5706), .Q(n10020) );
  INVX0 U10054 ( .INP(n10012), .ZN(n10016) );
  AND2X1 U10055 ( .IN1(g4983), .IN2(n9510), .Q(n10012) );
  AND2X1 U10056 ( .IN1(g4878), .IN2(n10021), .Q(n9510) );
  AND2X1 U10057 ( .IN1(n10022), .IN2(g4871), .Q(g34036) );
  AND2X1 U10058 ( .IN1(n10022), .IN2(g4864), .Q(g34035) );
  AND2X1 U10059 ( .IN1(n10022), .IN2(g4836), .Q(g34034) );
  OR2X1 U10060 ( .IN1(n8796), .IN2(n9896), .Q(n10022) );
  OR3X1 U10061 ( .IN1(n8346), .IN2(n1697), .IN3(n9810), .Q(n9896) );
  OR2X1 U10062 ( .IN1(n10023), .IN2(n10024), .Q(g34033) );
  AND2X1 U10063 ( .IN1(n8822), .IN2(g4818), .Q(n10024) );
  AND2X1 U10064 ( .IN1(n10025), .IN2(n10026), .Q(n10023) );
  XOR2X1 U10065 ( .IN1(g4793), .IN2(n9513), .Q(n10025) );
  OR4X1 U10066 ( .IN1(n10027), .IN2(n10028), .IN3(n10029), .IN4(n10030), .Q(
        g34032) );
  AND3X1 U10067 ( .IN1(n9039), .IN2(n9931), .IN3(n8751), .Q(n10030) );
  AND2X1 U10068 ( .IN1(n8822), .IN2(g4785), .Q(n10029) );
  AND2X1 U10069 ( .IN1(n10026), .IN2(g4709), .Q(n10028) );
  AND2X1 U10070 ( .IN1(n10031), .IN2(n9038), .Q(n10027) );
  OR2X1 U10071 ( .IN1(n10032), .IN2(n10033), .Q(g34031) );
  AND2X1 U10072 ( .IN1(n10026), .IN2(g4776), .Q(n10033) );
  AND2X1 U10073 ( .IN1(test_so29), .IN2(n10034), .Q(n10032) );
  OR2X1 U10074 ( .IN1(n8796), .IN2(n10035), .Q(n10034) );
  AND2X1 U10075 ( .IN1(n10036), .IN2(n10037), .Q(n10035) );
  OR3X1 U10076 ( .IN1(n10038), .IN2(n10039), .IN3(n10040), .Q(g34030) );
  AND2X1 U10077 ( .IN1(n8822), .IN2(g4793), .Q(n10040) );
  AND3X1 U10078 ( .IN1(n10036), .IN2(n8504), .IN3(n10037), .Q(n10039) );
  AND3X1 U10079 ( .IN1(test_so29), .IN2(n10026), .IN3(n10041), .Q(n10038) );
  OR3X1 U10080 ( .IN1(n10042), .IN2(n10043), .IN3(n10044), .Q(g34029) );
  AND2X1 U10081 ( .IN1(n8822), .IN2(g4776), .Q(n10044) );
  AND2X1 U10082 ( .IN1(n10031), .IN2(n5361), .Q(n10043) );
  AND3X1 U10083 ( .IN1(g4776), .IN2(n9931), .IN3(n10037), .Q(n10031) );
  INVX0 U10084 ( .INP(n10041), .ZN(n10037) );
  AND2X1 U10085 ( .IN1(n10026), .IN2(g4785), .Q(n10042) );
  AND2X1 U10086 ( .IN1(n8705), .IN2(n10036), .Q(n10026) );
  AND2X1 U10087 ( .IN1(n9931), .IN2(n10045), .Q(n10036) );
  OR2X1 U10088 ( .IN1(n10041), .IN2(n5707), .Q(n10045) );
  OR2X1 U10089 ( .IN1(n5368), .IN2(n9930), .Q(n10041) );
  INVX0 U10090 ( .INP(n9513), .ZN(n9930) );
  AND2X1 U10091 ( .IN1(g4688), .IN2(n10046), .Q(n9513) );
  AND2X1 U10092 ( .IN1(n9093), .IN2(g4674), .Q(g34027) );
  AND2X1 U10093 ( .IN1(n9093), .IN2(g4646), .Q(g34026) );
  OR2X1 U10094 ( .IN1(n8796), .IN2(n9931), .Q(n9093) );
  OR3X1 U10095 ( .IN1(n8346), .IN2(n1697), .IN3(n9811), .Q(n9931) );
  AND2X1 U10096 ( .IN1(n5727), .IN2(n9691), .Q(g34025) );
  AND2X1 U10097 ( .IN1(n9727), .IN2(n5382), .Q(n9691) );
  AND2X1 U10098 ( .IN1(n8706), .IN2(n9674), .Q(n9727) );
  OR2X1 U10099 ( .IN1(n10047), .IN2(DFF_961_n1), .Q(n9674) );
  AND2X1 U10100 ( .IN1(n10048), .IN2(n1697), .Q(n10047) );
  OR2X1 U10101 ( .IN1(n10049), .IN2(n10050), .Q(g34024) );
  AND3X1 U10102 ( .IN1(n10051), .IN2(n10052), .IN3(n8751), .Q(n10050) );
  OR2X1 U10103 ( .IN1(n10053), .IN2(n10054), .Q(n10052) );
  OR2X1 U10104 ( .IN1(n10048), .IN2(n10055), .Q(n10051) );
  AND2X1 U10105 ( .IN1(n8822), .IN2(g4492), .Q(n10049) );
  OR2X1 U10106 ( .IN1(n10056), .IN2(n10057), .Q(g34023) );
  AND2X1 U10107 ( .IN1(n10058), .IN2(n9325), .Q(n10057) );
  OR2X1 U10108 ( .IN1(n8797), .IN2(n10059), .Q(n10058) );
  AND4X1 U10109 ( .IN1(n10060), .IN2(g4555), .IN3(g4558), .IN4(g4561), .Q(
        n10059) );
  AND3X1 U10110 ( .IN1(n10054), .IN2(n8724), .IN3(n10060), .Q(n10056) );
  OR2X1 U10111 ( .IN1(n10048), .IN2(n10061), .Q(n10060) );
  INVX0 U10112 ( .INP(n9397), .ZN(n10048) );
  OR2X1 U10113 ( .IN1(n9397), .IN2(g2988), .Q(n10054) );
  OR4X1 U10114 ( .IN1(n2787), .IN2(n10062), .IN3(n10063), .IN4(n10064), .Q(
        g34022) );
  AND2X1 U10115 ( .IN1(n8822), .IN2(g2759), .Q(n10064) );
  AND3X1 U10116 ( .IN1(n10065), .IN2(g2763), .IN3(n8750), .Q(n10063) );
  INVX0 U10117 ( .INP(n10066), .ZN(n10065) );
  AND2X1 U10118 ( .IN1(n10066), .IN2(n7957), .Q(n10062) );
  AND2X1 U10119 ( .IN1(g2759), .IN2(n10067), .Q(n10066) );
  OR3X1 U10120 ( .IN1(n10068), .IN2(n10069), .IN3(n10070), .Q(g34021) );
  AND2X1 U10121 ( .IN1(n8822), .IN2(g2648), .Q(n10070) );
  AND2X1 U10122 ( .IN1(n10071), .IN2(g2567), .Q(n10069) );
  AND2X1 U10123 ( .IN1(n10072), .IN2(n10073), .Q(n10068) );
  OR2X1 U10124 ( .IN1(n10074), .IN2(n10075), .Q(g34020) );
  AND2X1 U10125 ( .IN1(n10076), .IN2(n8686), .Q(n10075) );
  OR2X1 U10126 ( .IN1(n10077), .IN2(n10078), .Q(n10076) );
  AND2X1 U10127 ( .IN1(n10079), .IN2(g2643), .Q(n10078) );
  OR2X1 U10128 ( .IN1(n10080), .IN2(n10081), .Q(n10079) );
  AND2X1 U10129 ( .IN1(n10082), .IN2(g2555), .Q(n10080) );
  AND2X1 U10130 ( .IN1(n10083), .IN2(n10084), .Q(n10077) );
  INVX0 U10131 ( .INP(n10082), .ZN(n10084) );
  OR2X1 U10132 ( .IN1(n10085), .IN2(n10072), .Q(n10083) );
  AND2X1 U10133 ( .IN1(n8021), .IN2(n10086), .Q(n10085) );
  AND2X1 U10134 ( .IN1(n10087), .IN2(g2629), .Q(n10074) );
  OR2X1 U10135 ( .IN1(n8796), .IN2(n10088), .Q(n10087) );
  AND2X1 U10136 ( .IN1(n10082), .IN2(g2643), .Q(n10088) );
  AND2X1 U10137 ( .IN1(n10089), .IN2(n10090), .Q(n10082) );
  OR2X1 U10138 ( .IN1(g1589), .IN2(n10091), .Q(n10090) );
  OR3X1 U10139 ( .IN1(n10092), .IN2(n10093), .IN3(n10094), .Q(g34019) );
  AND2X1 U10140 ( .IN1(n10095), .IN2(n10073), .Q(n10094) );
  AND2X1 U10141 ( .IN1(n8822), .IN2(g2571), .Q(n10093) );
  AND3X1 U10142 ( .IN1(n10096), .IN2(g2583), .IN3(n8751), .Q(n10092) );
  INVX0 U10143 ( .INP(n10095), .ZN(n10096) );
  AND2X1 U10144 ( .IN1(g2629), .IN2(n10097), .Q(n10095) );
  OR3X1 U10145 ( .IN1(n10098), .IN2(n10099), .IN3(n10100), .Q(g34018) );
  AND2X1 U10146 ( .IN1(n10101), .IN2(n10073), .Q(n10100) );
  INVX0 U10147 ( .INP(n10102), .ZN(n10101) );
  AND2X1 U10148 ( .IN1(n8823), .IN2(g2583), .Q(n10099) );
  AND3X1 U10149 ( .IN1(test_so61), .IN2(n10102), .IN3(n8750), .Q(n10098) );
  OR2X1 U10150 ( .IN1(n10081), .IN2(n10103), .Q(n10102) );
  OR3X1 U10151 ( .IN1(n10104), .IN2(n10105), .IN3(n10106), .Q(g34017) );
  AND2X1 U10152 ( .IN1(n10107), .IN2(n10073), .Q(n10106) );
  AND2X1 U10153 ( .IN1(test_so61), .IN2(n8810), .Q(n10105) );
  AND3X1 U10154 ( .IN1(test_so66), .IN2(n10108), .IN3(n8749), .Q(n10104) );
  INVX0 U10155 ( .INP(n10107), .ZN(n10108) );
  AND3X1 U10156 ( .IN1(g2629), .IN2(g2555), .IN3(n10086), .Q(n10107) );
  OR3X1 U10157 ( .IN1(n10109), .IN2(n10110), .IN3(n10111), .Q(g34016) );
  AND2X1 U10158 ( .IN1(n10112), .IN2(n10073), .Q(n10111) );
  AND2X1 U10159 ( .IN1(n8823), .IN2(g2563), .Q(n10110) );
  AND3X1 U10160 ( .IN1(n10113), .IN2(g2571), .IN3(n8751), .Q(n10109) );
  INVX0 U10161 ( .INP(n10112), .ZN(n10113) );
  AND3X1 U10162 ( .IN1(g2599), .IN2(n10086), .IN3(n5521), .Q(n10112) );
  OR3X1 U10163 ( .IN1(n10114), .IN2(n10115), .IN3(n10116), .Q(g34015) );
  AND2X1 U10164 ( .IN1(n10117), .IN2(n10073), .Q(n10116) );
  AND2X1 U10165 ( .IN1(n8707), .IN2(n10118), .Q(n10073) );
  INVX0 U10166 ( .INP(n10119), .ZN(n10118) );
  AND2X1 U10167 ( .IN1(n10089), .IN2(n10120), .Q(n10119) );
  OR2X1 U10168 ( .IN1(n10091), .IN2(g1585), .Q(n10120) );
  OR3X1 U10169 ( .IN1(n10121), .IN2(n10122), .IN3(n10123), .Q(n10089) );
  AND2X1 U10170 ( .IN1(n5483), .IN2(n10124), .Q(n10123) );
  INVX0 U10171 ( .INP(n10091), .ZN(n10122) );
  AND2X1 U10172 ( .IN1(n8823), .IN2(g2567), .Q(n10115) );
  AND3X1 U10173 ( .IN1(n10125), .IN2(g2563), .IN3(n8751), .Q(n10114) );
  INVX0 U10174 ( .INP(n10117), .ZN(n10125) );
  AND2X1 U10175 ( .IN1(g2555), .IN2(n10097), .Q(n10117) );
  OR3X1 U10176 ( .IN1(n10126), .IN2(n10127), .IN3(n10128), .Q(g34014) );
  AND2X1 U10177 ( .IN1(n8823), .IN2(g2514), .Q(n10128) );
  AND2X1 U10178 ( .IN1(n10129), .IN2(g2433), .Q(n10127) );
  AND2X1 U10179 ( .IN1(n10130), .IN2(n10131), .Q(n10126) );
  OR2X1 U10180 ( .IN1(n10132), .IN2(n10133), .Q(g34013) );
  AND2X1 U10181 ( .IN1(n10134), .IN2(n8685), .Q(n10133) );
  OR2X1 U10182 ( .IN1(n10135), .IN2(n10136), .Q(n10134) );
  AND2X1 U10183 ( .IN1(n10137), .IN2(g2509), .Q(n10136) );
  OR2X1 U10184 ( .IN1(n10138), .IN2(n10139), .Q(n10137) );
  AND2X1 U10185 ( .IN1(test_so79), .IN2(n10140), .Q(n10138) );
  AND2X1 U10186 ( .IN1(n10141), .IN2(n10142), .Q(n10135) );
  INVX0 U10187 ( .INP(n10140), .ZN(n10142) );
  OR2X1 U10188 ( .IN1(n10143), .IN2(n10130), .Q(n10141) );
  AND2X1 U10189 ( .IN1(n8020), .IN2(n10144), .Q(n10143) );
  AND2X1 U10190 ( .IN1(n10145), .IN2(g2495), .Q(n10132) );
  OR2X1 U10191 ( .IN1(n8797), .IN2(n10146), .Q(n10145) );
  AND2X1 U10192 ( .IN1(n10140), .IN2(g2509), .Q(n10146) );
  AND2X1 U10193 ( .IN1(n10147), .IN2(n10148), .Q(n10140) );
  OR2X1 U10194 ( .IN1(n10149), .IN2(n5755), .Q(n10148) );
  OR3X1 U10195 ( .IN1(n10150), .IN2(n10151), .IN3(n10152), .Q(g34012) );
  AND2X1 U10196 ( .IN1(n10153), .IN2(n10131), .Q(n10152) );
  AND2X1 U10197 ( .IN1(n8823), .IN2(g2437), .Q(n10151) );
  AND3X1 U10198 ( .IN1(n10154), .IN2(g2449), .IN3(n8750), .Q(n10150) );
  INVX0 U10199 ( .INP(n10153), .ZN(n10154) );
  AND2X1 U10200 ( .IN1(g2495), .IN2(n10155), .Q(n10153) );
  OR3X1 U10201 ( .IN1(n10156), .IN2(n10157), .IN3(n10158), .Q(g34011) );
  AND2X1 U10202 ( .IN1(n10159), .IN2(n10131), .Q(n10158) );
  INVX0 U10203 ( .INP(n10160), .ZN(n10159) );
  AND2X1 U10204 ( .IN1(n8823), .IN2(g2449), .Q(n10157) );
  AND3X1 U10205 ( .IN1(n10160), .IN2(n9274), .IN3(n8751), .Q(n10156) );
  OR2X1 U10206 ( .IN1(n10139), .IN2(n10161), .Q(n10160) );
  OR3X1 U10207 ( .IN1(n10162), .IN2(n10163), .IN3(n10164), .Q(g34010) );
  AND2X1 U10208 ( .IN1(n10165), .IN2(n10131), .Q(n10164) );
  AND2X1 U10209 ( .IN1(n8823), .IN2(n9274), .Q(n10163) );
  AND3X1 U10210 ( .IN1(n10166), .IN2(g2441), .IN3(n8751), .Q(n10162) );
  INVX0 U10211 ( .INP(n10165), .ZN(n10166) );
  AND3X1 U10212 ( .IN1(g2495), .IN2(n10144), .IN3(test_so79), .Q(n10165) );
  OR3X1 U10213 ( .IN1(n10167), .IN2(n10168), .IN3(n10169), .Q(g34009) );
  AND2X1 U10214 ( .IN1(n10170), .IN2(n10131), .Q(n10169) );
  AND2X1 U10215 ( .IN1(n8823), .IN2(g2429), .Q(n10168) );
  AND3X1 U10216 ( .IN1(n10171), .IN2(g2437), .IN3(n8749), .Q(n10167) );
  INVX0 U10217 ( .INP(n10170), .ZN(n10171) );
  AND3X1 U10218 ( .IN1(g2465), .IN2(n10144), .IN3(n5522), .Q(n10170) );
  OR3X1 U10219 ( .IN1(n10172), .IN2(n10173), .IN3(n10174), .Q(g34008) );
  AND2X1 U10220 ( .IN1(n10175), .IN2(n10131), .Q(n10174) );
  AND2X1 U10221 ( .IN1(n8708), .IN2(n10176), .Q(n10131) );
  INVX0 U10222 ( .INP(n10177), .ZN(n10176) );
  AND2X1 U10223 ( .IN1(n10147), .IN2(n10178), .Q(n10177) );
  OR2X1 U10224 ( .IN1(n5757), .IN2(n10149), .Q(n10178) );
  OR3X1 U10225 ( .IN1(n10121), .IN2(n10179), .IN3(n10180), .Q(n10147) );
  AND2X1 U10226 ( .IN1(n5290), .IN2(n10124), .Q(n10180) );
  INVX0 U10227 ( .INP(n10149), .ZN(n10179) );
  AND2X1 U10228 ( .IN1(n8823), .IN2(g2433), .Q(n10173) );
  AND3X1 U10229 ( .IN1(n10181), .IN2(g2429), .IN3(n8750), .Q(n10172) );
  INVX0 U10230 ( .INP(n10175), .ZN(n10181) );
  AND2X1 U10231 ( .IN1(test_so79), .IN2(n10155), .Q(n10175) );
  OR3X1 U10232 ( .IN1(n10182), .IN2(n10183), .IN3(n10184), .Q(g34007) );
  AND2X1 U10233 ( .IN1(n8823), .IN2(g2380), .Q(n10184) );
  AND2X1 U10234 ( .IN1(n10185), .IN2(g2299), .Q(n10183) );
  AND2X1 U10235 ( .IN1(n10186), .IN2(n10187), .Q(n10182) );
  OR2X1 U10236 ( .IN1(n10188), .IN2(n10189), .Q(g34006) );
  AND2X1 U10237 ( .IN1(n10190), .IN2(n8685), .Q(n10189) );
  OR2X1 U10238 ( .IN1(n10191), .IN2(n10192), .Q(n10190) );
  AND2X1 U10239 ( .IN1(n10193), .IN2(g2375), .Q(n10192) );
  OR2X1 U10240 ( .IN1(n10194), .IN2(n10195), .Q(n10193) );
  AND2X1 U10241 ( .IN1(n10196), .IN2(g2287), .Q(n10194) );
  AND2X1 U10242 ( .IN1(n10197), .IN2(n10198), .Q(n10191) );
  INVX0 U10243 ( .INP(n10196), .ZN(n10198) );
  OR2X1 U10244 ( .IN1(n10199), .IN2(n10186), .Q(n10197) );
  AND2X1 U10245 ( .IN1(n8022), .IN2(n10200), .Q(n10199) );
  AND2X1 U10246 ( .IN1(n10201), .IN2(g2361), .Q(n10188) );
  OR2X1 U10247 ( .IN1(n8797), .IN2(n10202), .Q(n10201) );
  AND2X1 U10248 ( .IN1(n10196), .IN2(g2375), .Q(n10202) );
  AND2X1 U10249 ( .IN1(n10203), .IN2(n10204), .Q(n10196) );
  OR2X1 U10250 ( .IN1(n10205), .IN2(g1589), .Q(n10204) );
  OR3X1 U10251 ( .IN1(n10206), .IN2(n10207), .IN3(n10208), .Q(g34005) );
  AND2X1 U10252 ( .IN1(n10209), .IN2(n10187), .Q(n10208) );
  INVX0 U10253 ( .INP(n10210), .ZN(n10209) );
  AND2X1 U10254 ( .IN1(n8823), .IN2(g2303), .Q(n10207) );
  AND3X1 U10255 ( .IN1(n10210), .IN2(g2315), .IN3(n8750), .Q(n10206) );
  OR2X1 U10256 ( .IN1(g2331), .IN2(n10211), .Q(n10210) );
  OR3X1 U10257 ( .IN1(n10212), .IN2(n10213), .IN3(n10214), .Q(g34004) );
  AND2X1 U10258 ( .IN1(n10215), .IN2(n10187), .Q(n10214) );
  INVX0 U10259 ( .INP(n10216), .ZN(n10215) );
  AND2X1 U10260 ( .IN1(n8823), .IN2(g2315), .Q(n10213) );
  AND3X1 U10261 ( .IN1(n10216), .IN2(n9314), .IN3(n8750), .Q(n10212) );
  OR2X1 U10262 ( .IN1(n10195), .IN2(n10217), .Q(n10216) );
  OR3X1 U10263 ( .IN1(n10218), .IN2(n10219), .IN3(n10220), .Q(g34003) );
  AND2X1 U10264 ( .IN1(n10221), .IN2(n10187), .Q(n10220) );
  INVX0 U10265 ( .INP(n10222), .ZN(n10221) );
  AND2X1 U10266 ( .IN1(n8823), .IN2(n9314), .Q(n10219) );
  AND3X1 U10267 ( .IN1(n10222), .IN2(g2307), .IN3(n8748), .Q(n10218) );
  OR2X1 U10268 ( .IN1(n5353), .IN2(n10211), .Q(n10222) );
  OR2X1 U10269 ( .IN1(n10195), .IN2(n5537), .Q(n10211) );
  OR3X1 U10270 ( .IN1(n10223), .IN2(n10224), .IN3(n10225), .Q(g34002) );
  AND2X1 U10271 ( .IN1(n10226), .IN2(n10187), .Q(n10225) );
  AND2X1 U10272 ( .IN1(n8823), .IN2(g2295), .Q(n10224) );
  AND3X1 U10273 ( .IN1(n10227), .IN2(g2303), .IN3(n8749), .Q(n10223) );
  INVX0 U10274 ( .INP(n10226), .ZN(n10227) );
  AND3X1 U10275 ( .IN1(g2331), .IN2(n10200), .IN3(n5537), .Q(n10226) );
  OR3X1 U10276 ( .IN1(n10228), .IN2(n10229), .IN3(n10230), .Q(g34001) );
  AND2X1 U10277 ( .IN1(n10231), .IN2(n10187), .Q(n10230) );
  AND2X1 U10278 ( .IN1(n8705), .IN2(n10232), .Q(n10187) );
  INVX0 U10279 ( .INP(n10233), .ZN(n10232) );
  AND2X1 U10280 ( .IN1(n10203), .IN2(n10234), .Q(n10233) );
  OR2X1 U10281 ( .IN1(g1585), .IN2(n10205), .Q(n10234) );
  OR3X1 U10282 ( .IN1(n10121), .IN2(n10235), .IN3(n10236), .Q(n10203) );
  AND2X1 U10283 ( .IN1(n5343), .IN2(n10124), .Q(n10236) );
  INVX0 U10284 ( .INP(n10205), .ZN(n10235) );
  AND2X1 U10285 ( .IN1(n8823), .IN2(g2299), .Q(n10229) );
  AND3X1 U10286 ( .IN1(n10237), .IN2(g2295), .IN3(n8749), .Q(n10228) );
  INVX0 U10287 ( .INP(n10231), .ZN(n10237) );
  AND3X1 U10288 ( .IN1(g2287), .IN2(n10200), .IN3(n5513), .Q(n10231) );
  OR3X1 U10289 ( .IN1(n10238), .IN2(n10239), .IN3(n10240), .Q(g34000) );
  AND2X1 U10290 ( .IN1(n8823), .IN2(g2246), .Q(n10240) );
  AND2X1 U10291 ( .IN1(n10241), .IN2(g2165), .Q(n10239) );
  AND2X1 U10292 ( .IN1(n10242), .IN2(n10243), .Q(n10238) );
  OR2X1 U10293 ( .IN1(n10244), .IN2(n10245), .Q(g33999) );
  AND2X1 U10294 ( .IN1(n10246), .IN2(n8685), .Q(n10245) );
  OR2X1 U10295 ( .IN1(n10247), .IN2(n10248), .Q(n10246) );
  AND2X1 U10296 ( .IN1(n10249), .IN2(g2241), .Q(n10248) );
  OR2X1 U10297 ( .IN1(n10250), .IN2(n10251), .Q(n10249) );
  AND2X1 U10298 ( .IN1(n10252), .IN2(g2153), .Q(n10250) );
  AND2X1 U10299 ( .IN1(n10253), .IN2(n10254), .Q(n10247) );
  INVX0 U10300 ( .INP(n10252), .ZN(n10254) );
  OR2X1 U10301 ( .IN1(n10255), .IN2(n10242), .Q(n10253) );
  AND2X1 U10302 ( .IN1(n8024), .IN2(n10256), .Q(n10255) );
  AND2X1 U10303 ( .IN1(n10257), .IN2(g2227), .Q(n10244) );
  OR2X1 U10304 ( .IN1(n8798), .IN2(n10258), .Q(n10257) );
  AND2X1 U10305 ( .IN1(n10252), .IN2(g2241), .Q(n10258) );
  AND2X1 U10306 ( .IN1(n10259), .IN2(n10260), .Q(n10252) );
  OR2X1 U10307 ( .IN1(n10261), .IN2(n5755), .Q(n10260) );
  OR3X1 U10308 ( .IN1(n10262), .IN2(n10263), .IN3(n10264), .Q(g33998) );
  AND2X1 U10309 ( .IN1(n10265), .IN2(n10243), .Q(n10264) );
  INVX0 U10310 ( .INP(n10266), .ZN(n10265) );
  AND2X1 U10311 ( .IN1(n8823), .IN2(g2169), .Q(n10263) );
  AND3X1 U10312 ( .IN1(n10266), .IN2(g2181), .IN3(n8750), .Q(n10262) );
  OR2X1 U10313 ( .IN1(g2197), .IN2(n10267), .Q(n10266) );
  OR3X1 U10315 ( .IN1(n10268), .IN2(n10269), .IN3(n10270), .Q(g33997) );
  AND2X1 U10316 ( .IN1(n10271), .IN2(n10243), .Q(n10270) );
  INVX0 U10317 ( .INP(n10272), .ZN(n10271) );
  AND2X1 U10319 ( .IN1(n8823), .IN2(g2181), .Q(n10269) );
  AND3X1 U10320 ( .IN1(n10272), .IN2(n9352), .IN3(n8749), .Q(n10268) );
  OR2X1 U10321 ( .IN1(n10251), .IN2(n10273), .Q(n10272) );
  OR3X1 U10322 ( .IN1(n10274), .IN2(n10275), .IN3(n10276), .Q(g33996) );
  AND2X1 U10323 ( .IN1(n10277), .IN2(n10243), .Q(n10276) );
  INVX0 U10324 ( .INP(n10278), .ZN(n10277) );
  AND2X1 U10325 ( .IN1(n8823), .IN2(n9352), .Q(n10275) );
  AND3X1 U10326 ( .IN1(n10278), .IN2(g2173), .IN3(n8746), .Q(n10274) );
  OR2X1 U10327 ( .IN1(n5356), .IN2(n10267), .Q(n10278) );
  OR2X1 U10328 ( .IN1(n10251), .IN2(n5538), .Q(n10267) );
  OR3X1 U10329 ( .IN1(n10279), .IN2(n10280), .IN3(n10281), .Q(g33995) );
  AND2X1 U10330 ( .IN1(n10282), .IN2(n10243), .Q(n10281) );
  AND2X1 U10331 ( .IN1(n8823), .IN2(g2161), .Q(n10280) );
  AND3X1 U10332 ( .IN1(n10283), .IN2(g2169), .IN3(n8749), .Q(n10279) );
  INVX0 U10333 ( .INP(n10282), .ZN(n10283) );
  AND3X1 U10334 ( .IN1(g2197), .IN2(n10256), .IN3(n5538), .Q(n10282) );
  OR3X1 U10335 ( .IN1(n10284), .IN2(n10285), .IN3(n10286), .Q(g33994) );
  AND2X1 U10336 ( .IN1(n10287), .IN2(n10243), .Q(n10286) );
  AND2X1 U10337 ( .IN1(n8705), .IN2(n10288), .Q(n10243) );
  INVX0 U10338 ( .INP(n10289), .ZN(n10288) );
  AND2X1 U10339 ( .IN1(n10259), .IN2(n10290), .Q(n10289) );
  OR2X1 U10340 ( .IN1(n5757), .IN2(n10261), .Q(n10290) );
  OR3X1 U10341 ( .IN1(n10121), .IN2(n10291), .IN3(n10292), .Q(n10259) );
  AND2X1 U10342 ( .IN1(n5289), .IN2(n10124), .Q(n10292) );
  INVX0 U10343 ( .INP(n10261), .ZN(n10291) );
  AND2X1 U10344 ( .IN1(g1291), .IN2(n10124), .Q(n10121) );
  AND2X1 U10345 ( .IN1(g4180), .IN2(n10293), .Q(n10124) );
  AND2X1 U10346 ( .IN1(n8823), .IN2(g2165), .Q(n10285) );
  AND3X1 U10347 ( .IN1(n10294), .IN2(g2161), .IN3(n8749), .Q(n10284) );
  INVX0 U10348 ( .INP(n10287), .ZN(n10294) );
  AND3X1 U10349 ( .IN1(g2153), .IN2(n10256), .IN3(n5514), .Q(n10287) );
  OR3X1 U10350 ( .IN1(n10295), .IN2(n10296), .IN3(n10297), .Q(g33993) );
  AND2X1 U10351 ( .IN1(n8823), .IN2(g2089), .Q(n10297) );
  AND2X1 U10352 ( .IN1(n10298), .IN2(g2008), .Q(n10296) );
  AND2X1 U10353 ( .IN1(n10299), .IN2(n10300), .Q(n10295) );
  OR2X1 U10354 ( .IN1(n10301), .IN2(n10302), .Q(g33992) );
  AND2X1 U10355 ( .IN1(n10303), .IN2(n8686), .Q(n10302) );
  OR2X1 U10356 ( .IN1(n10304), .IN2(n10305), .Q(n10303) );
  AND2X1 U10357 ( .IN1(n10306), .IN2(g2084), .Q(n10305) );
  OR2X1 U10358 ( .IN1(n10307), .IN2(n10308), .Q(n10306) );
  AND2X1 U10359 ( .IN1(n10309), .IN2(g1996), .Q(n10307) );
  AND2X1 U10360 ( .IN1(n10310), .IN2(n10311), .Q(n10304) );
  INVX0 U10361 ( .INP(n10309), .ZN(n10311) );
  OR2X1 U10362 ( .IN1(n10312), .IN2(n10299), .Q(n10310) );
  AND2X1 U10363 ( .IN1(n8019), .IN2(n10313), .Q(n10312) );
  AND2X1 U10364 ( .IN1(n10314), .IN2(g2070), .Q(n10301) );
  OR2X1 U10365 ( .IN1(n8798), .IN2(n10315), .Q(n10314) );
  AND2X1 U10366 ( .IN1(n10309), .IN2(g2084), .Q(n10315) );
  AND2X1 U10367 ( .IN1(n10316), .IN2(n10317), .Q(n10309) );
  OR2X1 U10368 ( .IN1(g1246), .IN2(n10318), .Q(n10317) );
  OR3X1 U10369 ( .IN1(n10319), .IN2(n10320), .IN3(n10321), .Q(g33991) );
  AND2X1 U10370 ( .IN1(n10322), .IN2(n10300), .Q(n10321) );
  INVX0 U10371 ( .INP(n10323), .ZN(n10322) );
  AND2X1 U10372 ( .IN1(n8824), .IN2(g2012), .Q(n10320) );
  AND3X1 U10373 ( .IN1(n10323), .IN2(g2024), .IN3(n8749), .Q(n10319) );
  OR2X1 U10374 ( .IN1(g2040), .IN2(n10324), .Q(n10323) );
  OR3X1 U10375 ( .IN1(n10325), .IN2(n10326), .IN3(n10327), .Q(g33990) );
  AND2X1 U10376 ( .IN1(n10328), .IN2(n10300), .Q(n10327) );
  INVX0 U10377 ( .INP(n10329), .ZN(n10328) );
  AND2X1 U10378 ( .IN1(n8824), .IN2(g2024), .Q(n10326) );
  AND3X1 U10379 ( .IN1(n10329), .IN2(n9312), .IN3(n8749), .Q(n10325) );
  OR2X1 U10380 ( .IN1(n10308), .IN2(n10330), .Q(n10329) );
  OR3X1 U10381 ( .IN1(n10331), .IN2(n10332), .IN3(n10333), .Q(g33989) );
  AND2X1 U10382 ( .IN1(n10334), .IN2(n10300), .Q(n10333) );
  INVX0 U10383 ( .INP(n10335), .ZN(n10334) );
  AND2X1 U10384 ( .IN1(n8824), .IN2(n9312), .Q(n10332) );
  AND3X1 U10385 ( .IN1(n10335), .IN2(g2016), .IN3(n8749), .Q(n10331) );
  OR2X1 U10386 ( .IN1(n5355), .IN2(n10324), .Q(n10335) );
  OR2X1 U10387 ( .IN1(n10308), .IN2(n5535), .Q(n10324) );
  OR3X1 U10388 ( .IN1(n10336), .IN2(n10337), .IN3(n10338), .Q(g33988) );
  AND2X1 U10389 ( .IN1(n10339), .IN2(n10300), .Q(n10338) );
  AND2X1 U10390 ( .IN1(n8824), .IN2(g2004), .Q(n10337) );
  AND3X1 U10391 ( .IN1(n10340), .IN2(g2012), .IN3(n8748), .Q(n10336) );
  INVX0 U10392 ( .INP(n10339), .ZN(n10340) );
  AND3X1 U10393 ( .IN1(g2040), .IN2(n10313), .IN3(n5535), .Q(n10339) );
  OR3X1 U10394 ( .IN1(n10341), .IN2(n10342), .IN3(n10343), .Q(g33987) );
  AND2X1 U10395 ( .IN1(n10344), .IN2(n10300), .Q(n10343) );
  AND2X1 U10396 ( .IN1(n8707), .IN2(n10345), .Q(n10300) );
  INVX0 U10397 ( .INP(n10346), .ZN(n10345) );
  AND2X1 U10398 ( .IN1(n10316), .IN2(n10347), .Q(n10346) );
  OR2X1 U10399 ( .IN1(n10318), .IN2(g30332), .Q(n10347) );
  OR3X1 U10400 ( .IN1(n10348), .IN2(n10349), .IN3(n10350), .Q(n10316) );
  AND2X1 U10401 ( .IN1(n5341), .IN2(n10351), .Q(n10350) );
  AND2X1 U10402 ( .IN1(n8824), .IN2(g2008), .Q(n10342) );
  AND3X1 U10403 ( .IN1(n10352), .IN2(g2004), .IN3(n8748), .Q(n10341) );
  INVX0 U10404 ( .INP(n10344), .ZN(n10352) );
  AND3X1 U10405 ( .IN1(g1996), .IN2(n10313), .IN3(n5505), .Q(n10344) );
  OR3X1 U10406 ( .IN1(n10353), .IN2(n10354), .IN3(n10355), .Q(g33986) );
  AND2X1 U10407 ( .IN1(n8824), .IN2(g1955), .Q(n10355) );
  AND2X1 U10408 ( .IN1(n10356), .IN2(g1874), .Q(n10354) );
  AND2X1 U10409 ( .IN1(n10357), .IN2(n10358), .Q(n10353) );
  OR2X1 U10410 ( .IN1(n10359), .IN2(n10360), .Q(g33985) );
  AND2X1 U10411 ( .IN1(n10361), .IN2(n8690), .Q(n10360) );
  OR2X1 U10412 ( .IN1(n10362), .IN2(n10363), .Q(n10361) );
  AND2X1 U10413 ( .IN1(n10364), .IN2(g1950), .Q(n10363) );
  OR2X1 U10414 ( .IN1(n10365), .IN2(n10366), .Q(n10364) );
  AND2X1 U10415 ( .IN1(test_so8), .IN2(n10367), .Q(n10365) );
  AND2X1 U10416 ( .IN1(n10368), .IN2(n10369), .Q(n10362) );
  INVX0 U10417 ( .INP(n10367), .ZN(n10369) );
  OR2X1 U10418 ( .IN1(n10370), .IN2(n10357), .Q(n10368) );
  AND2X1 U10419 ( .IN1(n8023), .IN2(n10371), .Q(n10370) );
  AND2X1 U10420 ( .IN1(n10372), .IN2(g1936), .Q(n10359) );
  OR2X1 U10421 ( .IN1(n8799), .IN2(n10373), .Q(n10372) );
  AND2X1 U10422 ( .IN1(n10367), .IN2(g1950), .Q(n10373) );
  AND2X1 U10423 ( .IN1(n10374), .IN2(n10375), .Q(n10367) );
  OR2X1 U10424 ( .IN1(n10376), .IN2(n5756), .Q(n10375) );
  OR3X1 U10425 ( .IN1(n10377), .IN2(n10378), .IN3(n10379), .Q(g33984) );
  AND2X1 U10426 ( .IN1(n10380), .IN2(n10358), .Q(n10379) );
  INVX0 U10427 ( .INP(n10381), .ZN(n10380) );
  AND2X1 U10428 ( .IN1(n8824), .IN2(g1878), .Q(n10378) );
  AND3X1 U10429 ( .IN1(n10381), .IN2(g1890), .IN3(n8748), .Q(n10377) );
  OR2X1 U10430 ( .IN1(g1906), .IN2(n10382), .Q(n10381) );
  OR3X1 U10431 ( .IN1(n10383), .IN2(n10384), .IN3(n10385), .Q(g33983) );
  AND2X1 U10432 ( .IN1(n10386), .IN2(n10358), .Q(n10385) );
  INVX0 U10433 ( .INP(n10387), .ZN(n10386) );
  AND2X1 U10434 ( .IN1(n8824), .IN2(g1890), .Q(n10384) );
  AND3X1 U10435 ( .IN1(n10387), .IN2(n9280), .IN3(n8748), .Q(n10383) );
  OR2X1 U10436 ( .IN1(n10366), .IN2(n10388), .Q(n10387) );
  OR3X1 U10437 ( .IN1(n10389), .IN2(n10390), .IN3(n10391), .Q(g33982) );
  AND2X1 U10438 ( .IN1(n10392), .IN2(n10358), .Q(n10391) );
  INVX0 U10439 ( .INP(n10393), .ZN(n10392) );
  AND2X1 U10440 ( .IN1(n8824), .IN2(n9280), .Q(n10390) );
  AND3X1 U10441 ( .IN1(n10393), .IN2(g1882), .IN3(n8748), .Q(n10389) );
  OR2X1 U10442 ( .IN1(n8502), .IN2(n10382), .Q(n10393) );
  OR2X1 U10443 ( .IN1(n10366), .IN2(n5534), .Q(n10382) );
  OR3X1 U10444 ( .IN1(n10394), .IN2(n10395), .IN3(n10396), .Q(g33981) );
  AND2X1 U10445 ( .IN1(n10397), .IN2(n10358), .Q(n10396) );
  AND2X1 U10446 ( .IN1(n8824), .IN2(g1870), .Q(n10395) );
  AND3X1 U10447 ( .IN1(n10398), .IN2(g1878), .IN3(n8748), .Q(n10394) );
  INVX0 U10448 ( .INP(n10397), .ZN(n10398) );
  AND3X1 U10449 ( .IN1(g1906), .IN2(n10371), .IN3(n5534), .Q(n10397) );
  OR3X1 U10450 ( .IN1(n10399), .IN2(n10400), .IN3(n10401), .Q(g33980) );
  AND2X1 U10451 ( .IN1(n10402), .IN2(n10358), .Q(n10401) );
  AND2X1 U10452 ( .IN1(n8706), .IN2(n10403), .Q(n10358) );
  INVX0 U10453 ( .INP(n10404), .ZN(n10403) );
  AND2X1 U10454 ( .IN1(n10374), .IN2(n10405), .Q(n10404) );
  OR2X1 U10455 ( .IN1(n5526), .IN2(n10376), .Q(n10405) );
  OR3X1 U10456 ( .IN1(n10348), .IN2(n10406), .IN3(n10407), .Q(n10374) );
  AND2X1 U10457 ( .IN1(n5329), .IN2(n10351), .Q(n10407) );
  INVX0 U10458 ( .INP(n10376), .ZN(n10406) );
  AND2X1 U10459 ( .IN1(n8824), .IN2(g1874), .Q(n10400) );
  AND3X1 U10460 ( .IN1(n10408), .IN2(g1870), .IN3(n8748), .Q(n10399) );
  INVX0 U10461 ( .INP(n10402), .ZN(n10408) );
  AND3X1 U10462 ( .IN1(n10371), .IN2(n5503), .IN3(test_so8), .Q(n10402) );
  OR3X1 U10463 ( .IN1(n10409), .IN2(n10410), .IN3(n10411), .Q(g33979) );
  AND2X1 U10464 ( .IN1(n8824), .IN2(g1821), .Q(n10411) );
  AND2X1 U10465 ( .IN1(n10412), .IN2(g1740), .Q(n10410) );
  AND2X1 U10466 ( .IN1(n10413), .IN2(n10414), .Q(n10409) );
  OR2X1 U10467 ( .IN1(n10415), .IN2(n10416), .Q(g33978) );
  AND2X1 U10468 ( .IN1(n10417), .IN2(n8690), .Q(n10416) );
  OR2X1 U10469 ( .IN1(n10418), .IN2(n10419), .Q(n10417) );
  AND2X1 U10470 ( .IN1(n10420), .IN2(g1816), .Q(n10419) );
  OR2X1 U10471 ( .IN1(n10421), .IN2(n10422), .Q(n10420) );
  AND2X1 U10472 ( .IN1(n10423), .IN2(g1728), .Q(n10421) );
  AND2X1 U10473 ( .IN1(n10424), .IN2(n10425), .Q(n10418) );
  INVX0 U10474 ( .INP(n10423), .ZN(n10425) );
  OR2X1 U10475 ( .IN1(n10426), .IN2(n10413), .Q(n10424) );
  AND2X1 U10476 ( .IN1(n7973), .IN2(n10427), .Q(n10426) );
  AND2X1 U10477 ( .IN1(n10428), .IN2(g1802), .Q(n10415) );
  OR2X1 U10478 ( .IN1(n8799), .IN2(n10429), .Q(n10428) );
  AND2X1 U10479 ( .IN1(n10423), .IN2(g1816), .Q(n10429) );
  AND2X1 U10480 ( .IN1(n10430), .IN2(n10431), .Q(n10423) );
  OR2X1 U10481 ( .IN1(n10432), .IN2(g1246), .Q(n10431) );
  OR3X1 U10482 ( .IN1(n10433), .IN2(n10434), .IN3(n10435), .Q(g33977) );
  AND2X1 U10483 ( .IN1(n10436), .IN2(n10414), .Q(n10435) );
  INVX0 U10484 ( .INP(n10437), .ZN(n10436) );
  AND2X1 U10485 ( .IN1(n8824), .IN2(g1744), .Q(n10434) );
  AND3X1 U10486 ( .IN1(n10437), .IN2(g1756), .IN3(n8748), .Q(n10433) );
  OR2X1 U10487 ( .IN1(g1772), .IN2(n10438), .Q(n10437) );
  OR3X1 U10488 ( .IN1(n10439), .IN2(n10440), .IN3(n10441), .Q(g33976) );
  AND2X1 U10489 ( .IN1(n10442), .IN2(n10414), .Q(n10441) );
  INVX0 U10490 ( .INP(n10443), .ZN(n10442) );
  AND2X1 U10491 ( .IN1(n8824), .IN2(g1756), .Q(n10440) );
  AND3X1 U10492 ( .IN1(n10443), .IN2(g1752), .IN3(n8748), .Q(n10439) );
  OR2X1 U10493 ( .IN1(n10422), .IN2(n10444), .Q(n10443) );
  OR3X1 U10494 ( .IN1(n10445), .IN2(n10446), .IN3(n10447), .Q(g33975) );
  AND2X1 U10495 ( .IN1(n10448), .IN2(n10414), .Q(n10447) );
  INVX0 U10496 ( .INP(n10449), .ZN(n10448) );
  AND2X1 U10497 ( .IN1(n8824), .IN2(g1752), .Q(n10446) );
  AND3X1 U10498 ( .IN1(n10449), .IN2(g1748), .IN3(n8747), .Q(n10445) );
  OR2X1 U10499 ( .IN1(n5352), .IN2(n10438), .Q(n10449) );
  OR2X1 U10500 ( .IN1(n10422), .IN2(n5536), .Q(n10438) );
  OR3X1 U10501 ( .IN1(n10450), .IN2(n10451), .IN3(n10452), .Q(g33974) );
  AND2X1 U10502 ( .IN1(n10453), .IN2(n10414), .Q(n10452) );
  AND2X1 U10503 ( .IN1(n8824), .IN2(g1736), .Q(n10451) );
  AND3X1 U10504 ( .IN1(n10454), .IN2(g1744), .IN3(n8747), .Q(n10450) );
  INVX0 U10505 ( .INP(n10453), .ZN(n10454) );
  AND3X1 U10506 ( .IN1(g1772), .IN2(n10427), .IN3(n5536), .Q(n10453) );
  OR3X1 U10507 ( .IN1(n10455), .IN2(n10456), .IN3(n10457), .Q(g33973) );
  AND2X1 U10508 ( .IN1(n10458), .IN2(n10414), .Q(n10457) );
  AND2X1 U10509 ( .IN1(n8707), .IN2(n10459), .Q(n10414) );
  INVX0 U10510 ( .INP(n10460), .ZN(n10459) );
  AND2X1 U10511 ( .IN1(n10430), .IN2(n10461), .Q(n10460) );
  OR2X1 U10512 ( .IN1(g30332), .IN2(n10432), .Q(n10461) );
  OR3X1 U10513 ( .IN1(n10348), .IN2(n10462), .IN3(n10463), .Q(n10430) );
  AND2X1 U10514 ( .IN1(n5478), .IN2(n10351), .Q(n10463) );
  INVX0 U10515 ( .INP(n10432), .ZN(n10462) );
  AND2X1 U10516 ( .IN1(n8824), .IN2(g1740), .Q(n10456) );
  AND3X1 U10517 ( .IN1(n10464), .IN2(g1736), .IN3(n8747), .Q(n10455) );
  INVX0 U10518 ( .INP(n10458), .ZN(n10464) );
  AND3X1 U10519 ( .IN1(g1728), .IN2(n10427), .IN3(n5504), .Q(n10458) );
  OR3X1 U10520 ( .IN1(n10465), .IN2(n10466), .IN3(n10467), .Q(g33972) );
  AND2X1 U10521 ( .IN1(n8824), .IN2(g1687), .Q(n10467) );
  AND2X1 U10522 ( .IN1(n10468), .IN2(g1604), .Q(n10466) );
  AND2X1 U10523 ( .IN1(n10469), .IN2(n10470), .Q(n10465) );
  OR2X1 U10524 ( .IN1(n10471), .IN2(n10472), .Q(g33971) );
  AND2X1 U10525 ( .IN1(n10473), .IN2(n8690), .Q(n10472) );
  OR2X1 U10526 ( .IN1(n10474), .IN2(n10475), .Q(n10473) );
  AND2X1 U10527 ( .IN1(n10476), .IN2(g1682), .Q(n10475) );
  OR2X1 U10528 ( .IN1(n10477), .IN2(n10478), .Q(n10476) );
  AND2X1 U10529 ( .IN1(n10479), .IN2(g1592), .Q(n10477) );
  AND2X1 U10530 ( .IN1(n10480), .IN2(n10481), .Q(n10474) );
  INVX0 U10531 ( .INP(n10479), .ZN(n10481) );
  OR2X1 U10532 ( .IN1(n10482), .IN2(n10469), .Q(n10480) );
  AND2X1 U10533 ( .IN1(n8025), .IN2(n10483), .Q(n10482) );
  AND2X1 U10534 ( .IN1(n10484), .IN2(g1668), .Q(n10471) );
  OR2X1 U10535 ( .IN1(n8800), .IN2(n10485), .Q(n10484) );
  AND2X1 U10536 ( .IN1(n10479), .IN2(g1682), .Q(n10485) );
  AND2X1 U10537 ( .IN1(n10486), .IN2(n10487), .Q(n10479) );
  OR2X1 U10538 ( .IN1(n10488), .IN2(n5756), .Q(n10487) );
  OR3X1 U10539 ( .IN1(n10489), .IN2(n10490), .IN3(n10491), .Q(g33970) );
  AND2X1 U10540 ( .IN1(n10492), .IN2(n10470), .Q(n10491) );
  AND2X1 U10541 ( .IN1(n8824), .IN2(g1608), .Q(n10490) );
  AND3X1 U10542 ( .IN1(n10493), .IN2(g1620), .IN3(n8747), .Q(n10489) );
  INVX0 U10543 ( .INP(n10492), .ZN(n10493) );
  AND2X1 U10544 ( .IN1(n10483), .IN2(g31862), .Q(n10492) );
  OR3X1 U10545 ( .IN1(n10494), .IN2(n10495), .IN3(n10496), .Q(g33969) );
  AND2X1 U10546 ( .IN1(n10497), .IN2(n10470), .Q(n10496) );
  AND2X1 U10547 ( .IN1(n8824), .IN2(g1620), .Q(n10495) );
  AND3X1 U10548 ( .IN1(n10498), .IN2(n9303), .IN3(n8747), .Q(n10494) );
  INVX0 U10549 ( .INP(n10497), .ZN(n10498) );
  AND2X1 U10550 ( .IN1(n5362), .IN2(n10499), .Q(n10497) );
  OR3X1 U10551 ( .IN1(n10500), .IN2(n10501), .IN3(n10502), .Q(g33968) );
  AND2X1 U10552 ( .IN1(n10503), .IN2(n10470), .Q(n10502) );
  AND2X1 U10553 ( .IN1(n8824), .IN2(n9303), .Q(n10501) );
  AND3X1 U10554 ( .IN1(n10504), .IN2(g1612), .IN3(n8747), .Q(n10500) );
  INVX0 U10555 ( .INP(n10503), .ZN(n10504) );
  AND2X1 U10556 ( .IN1(g1668), .IN2(n10505), .Q(n10503) );
  OR3X1 U10557 ( .IN1(n10506), .IN2(n10507), .IN3(n10508), .Q(g33967) );
  AND2X1 U10558 ( .IN1(n10509), .IN2(n10470), .Q(n10508) );
  AND2X1 U10559 ( .IN1(n8825), .IN2(g1600), .Q(n10507) );
  AND3X1 U10560 ( .IN1(n10510), .IN2(g1608), .IN3(n8747), .Q(n10506) );
  INVX0 U10561 ( .INP(n10509), .ZN(n10510) );
  AND2X1 U10562 ( .IN1(n5598), .IN2(n10499), .Q(n10509) );
  OR3X1 U10563 ( .IN1(n10511), .IN2(n10512), .IN3(n10513), .Q(g33966) );
  AND2X1 U10564 ( .IN1(n10514), .IN2(n10470), .Q(n10513) );
  INVX0 U10565 ( .INP(n10515), .ZN(n10470) );
  OR2X1 U10566 ( .IN1(n8800), .IN2(n10516), .Q(n10515) );
  AND2X1 U10567 ( .IN1(n10486), .IN2(n10517), .Q(n10516) );
  OR2X1 U10568 ( .IN1(n5526), .IN2(n10488), .Q(n10517) );
  OR3X1 U10569 ( .IN1(n10348), .IN2(n10518), .IN3(n10519), .Q(n10486) );
  AND2X1 U10570 ( .IN1(n5328), .IN2(n10351), .Q(n10519) );
  INVX0 U10571 ( .INP(n10488), .ZN(n10518) );
  AND2X1 U10572 ( .IN1(g947), .IN2(n10351), .Q(n10348) );
  AND2X1 U10573 ( .IN1(g4180), .IN2(n10520), .Q(n10351) );
  AND2X1 U10574 ( .IN1(n8825), .IN2(g1604), .Q(n10512) );
  AND3X1 U10575 ( .IN1(n10521), .IN2(g1600), .IN3(n8747), .Q(n10511) );
  INVX0 U10576 ( .INP(n10514), .ZN(n10521) );
  AND2X1 U10577 ( .IN1(n5549), .IN2(n10505), .Q(n10514) );
  OR3X1 U10578 ( .IN1(n10522), .IN2(n10523), .IN3(n10524), .Q(g33965) );
  AND2X1 U10579 ( .IN1(n8825), .IN2(g763), .Q(n10524) );
  AND2X1 U10580 ( .IN1(n2704), .IN2(n5333), .Q(n10523) );
  AND3X1 U10581 ( .IN1(n2404), .IN2(n10525), .IN3(g767), .Q(n10522) );
  INVX0 U10582 ( .INP(n2704), .ZN(n10525) );
  OR3X1 U10583 ( .IN1(n10526), .IN2(n10527), .IN3(n10528), .Q(g33964) );
  AND2X1 U10584 ( .IN1(n8825), .IN2(g595), .Q(n10528) );
  AND2X1 U10585 ( .IN1(n2706), .IN2(n5550), .Q(n10527) );
  AND3X1 U10586 ( .IN1(n2421), .IN2(n10529), .IN3(g599), .Q(n10526) );
  INVX0 U10587 ( .INP(n2706), .ZN(n10529) );
  OR2X1 U10588 ( .IN1(n10530), .IN2(n10531), .Q(g33963) );
  AND3X1 U10589 ( .IN1(n10532), .IN2(n10533), .IN3(n8747), .Q(n10531) );
  OR3X1 U10590 ( .IN1(g73), .IN2(n10534), .IN3(n10535), .Q(n10533) );
  AND2X1 U10591 ( .IN1(g72), .IN2(g262), .Q(n10535) );
  AND2X1 U10592 ( .IN1(n10536), .IN2(g269), .Q(n10534) );
  OR2X1 U10593 ( .IN1(n10537), .IN2(n9419), .Q(n10532) );
  AND2X1 U10594 ( .IN1(n10536), .IN2(g255), .Q(n10537) );
  AND2X1 U10595 ( .IN1(n8825), .IN2(g29215), .Q(n10530) );
  OR2X1 U10596 ( .IN1(n10538), .IN2(n10539), .Q(g33962) );
  AND3X1 U10597 ( .IN1(n10540), .IN2(n10541), .IN3(n8747), .Q(n10539) );
  OR2X1 U10598 ( .IN1(n10542), .IN2(n9419), .Q(n10541) );
  INVX0 U10599 ( .INP(g73), .ZN(n9419) );
  AND2X1 U10600 ( .IN1(n10543), .IN2(n10544), .Q(n10542) );
  OR2X1 U10601 ( .IN1(g72), .IN2(g232), .Q(n10544) );
  OR2X1 U10602 ( .IN1(n10536), .IN2(g225), .Q(n10543) );
  OR3X1 U10603 ( .IN1(g73), .IN2(n10545), .IN3(n10546), .Q(n10540) );
  AND2X1 U10604 ( .IN1(g72), .IN2(g239), .Q(n10546) );
  AND2X1 U10605 ( .IN1(n10536), .IN2(g246), .Q(n10545) );
  AND2X1 U10606 ( .IN1(n8825), .IN2(g479), .Q(n10538) );
  OR3X1 U10607 ( .IN1(n10547), .IN2(n10548), .IN3(n10549), .Q(g33961) );
  AND2X1 U10608 ( .IN1(n8825), .IN2(g294), .Q(n10549) );
  AND2X1 U10609 ( .IN1(n2989), .IN2(n5675), .Q(n10548) );
  AND3X1 U10610 ( .IN1(n8473), .IN2(n10550), .IN3(g298), .Q(n10547) );
  INVX0 U10611 ( .INP(n2989), .ZN(n10550) );
  OR3X1 U10612 ( .IN1(n10551), .IN2(n10552), .IN3(n10553), .Q(g33960) );
  AND2X1 U10613 ( .IN1(n8825), .IN2(g153), .Q(n10553) );
  AND2X1 U10614 ( .IN1(n2991), .IN2(n5678), .Q(n10552) );
  AND3X1 U10615 ( .IN1(n9969), .IN2(n10554), .IN3(g157), .Q(n10551) );
  INVX0 U10616 ( .INP(n2991), .ZN(n10554) );
  OR4X1 U10617 ( .IN1(g34649), .IN2(n9894), .IN3(n8355), .IN4(n8354), .Q(
        g33935) );
  OR4X1 U10618 ( .IN1(n10555), .IN2(n10556), .IN3(n10557), .IN4(n10558), .Q(
        g34649) );
  AND2X1 U10619 ( .IN1(n9067), .IN2(g4955), .Q(n10558) );
  AND2X1 U10620 ( .IN1(n9064), .IN2(g4933), .Q(n10556) );
  AND2X1 U10621 ( .IN1(n9065), .IN2(g4944), .Q(n10555) );
  OR3X1 U10622 ( .IN1(n5846), .IN2(n9894), .IN3(g18881), .Q(g33874) );
  OR4X1 U10623 ( .IN1(n9809), .IN2(n8986), .IN3(n10559), .IN4(n10560), .Q(
        g33659) );
  INVX0 U10624 ( .INP(n8984), .ZN(n10560) );
  XNOR2X1 U10625 ( .IN1(g4108), .IN2(g72), .Q(n8984) );
  INVX0 U10626 ( .INP(n8985), .ZN(n10559) );
  XNOR2X1 U10627 ( .IN1(g4104), .IN2(g73), .Q(n8985) );
  OR2X1 U10628 ( .IN1(n10561), .IN2(n10562), .Q(n8986) );
  AND2X1 U10629 ( .IN1(n10563), .IN2(g4098), .Q(n10562) );
  OR3X1 U10630 ( .IN1(n10564), .IN2(n10565), .IN3(n10566), .Q(n10563) );
  AND2X1 U10631 ( .IN1(n10567), .IN2(n10568), .Q(n10566) );
  AND2X1 U10632 ( .IN1(n10569), .IN2(n9807), .Q(n10565) );
  AND3X1 U10633 ( .IN1(n10570), .IN2(n10571), .IN3(g4093), .Q(n10564) );
  OR2X1 U10634 ( .IN1(n10572), .IN2(g4087), .Q(n10571) );
  OR2X1 U10635 ( .IN1(n5480), .IN2(n9012), .Q(n10570) );
  AND2X1 U10636 ( .IN1(n5350), .IN2(n10573), .Q(n10561) );
  OR3X1 U10637 ( .IN1(n10574), .IN2(n10575), .IN3(n10576), .Q(n10573) );
  AND2X1 U10638 ( .IN1(n10577), .IN2(n10568), .Q(n10576) );
  AND2X1 U10639 ( .IN1(g32975), .IN2(n9807), .Q(n10575) );
  AND3X1 U10640 ( .IN1(n10578), .IN2(n10579), .IN3(g4093), .Q(n10574) );
  OR2X1 U10641 ( .IN1(n10580), .IN2(g4087), .Q(n10579) );
  OR2X1 U10642 ( .IN1(n5480), .IN2(n10581), .Q(n10578) );
  OR2X1 U10643 ( .IN1(n9894), .IN2(n10582), .Q(n9809) );
  OR4X1 U10644 ( .IN1(g34657), .IN2(n9894), .IN3(n8353), .IN4(n8352), .Q(
        g33636) );
  INVX0 U10645 ( .INP(n2668), .ZN(n9894) );
  OR2X1 U10646 ( .IN1(n10583), .IN2(g134), .Q(n2668) );
  AND2X1 U10647 ( .IN1(g99), .IN2(g37), .Q(n10583) );
  OR4X1 U10648 ( .IN1(n10584), .IN2(n10585), .IN3(n10586), .IN4(n10587), .Q(
        g34657) );
  AND2X1 U10649 ( .IN1(n9041), .IN2(g4765), .Q(n10587) );
  AND2X1 U10650 ( .IN1(n9038), .IN2(g4743), .Q(n10585) );
  AND2X1 U10651 ( .IN1(n9039), .IN2(g4754), .Q(n10584) );
  OR2X1 U10652 ( .IN1(n10588), .IN2(n10589), .Q(g33627) );
  AND2X1 U10653 ( .IN1(n8825), .IN2(g6741), .Q(n10589) );
  AND2X1 U10654 ( .IN1(n10590), .IN2(n10591), .Q(n10588) );
  OR2X1 U10655 ( .IN1(n10592), .IN2(n10593), .Q(n10590) );
  AND2X1 U10656 ( .IN1(n9002), .IN2(n10594), .Q(n10593) );
  AND2X1 U10657 ( .IN1(n10595), .IN2(n8690), .Q(n10592) );
  OR2X1 U10658 ( .IN1(n10596), .IN2(n9005), .Q(n10595) );
  AND2X1 U10659 ( .IN1(n8479), .IN2(g6682), .Q(n10596) );
  OR3X1 U10660 ( .IN1(n10597), .IN2(n10598), .IN3(n10599), .Q(g33626) );
  AND2X1 U10661 ( .IN1(n10600), .IN2(g6741), .Q(n10599) );
  AND2X1 U10662 ( .IN1(n8825), .IN2(g6736), .Q(n10598) );
  AND4X1 U10663 ( .IN1(n10591), .IN2(n10594), .IN3(n5398), .IN4(n8721), .Q(
        n10597) );
  OR4X1 U10664 ( .IN1(n9810), .IN2(n10601), .IN3(test_so81), .IN4(n8479), .Q(
        n10591) );
  OR2X1 U10665 ( .IN1(n10602), .IN2(n10603), .Q(g33625) );
  AND2X1 U10666 ( .IN1(n8825), .IN2(g6395), .Q(n10603) );
  AND2X1 U10667 ( .IN1(n10604), .IN2(n10605), .Q(n10602) );
  OR2X1 U10668 ( .IN1(n10606), .IN2(n10607), .Q(n10604) );
  AND2X1 U10669 ( .IN1(n10608), .IN2(n10609), .Q(n10607) );
  AND2X1 U10670 ( .IN1(n10610), .IN2(n8690), .Q(n10606) );
  OR2X1 U10671 ( .IN1(n10611), .IN2(n10612), .Q(n10610) );
  AND2X1 U10672 ( .IN1(n10613), .IN2(g6336), .Q(n10611) );
  OR3X1 U10673 ( .IN1(n10614), .IN2(n10615), .IN3(n10616), .Q(g33624) );
  AND2X1 U10674 ( .IN1(n10617), .IN2(g6395), .Q(n10616) );
  AND2X1 U10675 ( .IN1(n8825), .IN2(g6390), .Q(n10615) );
  AND4X1 U10676 ( .IN1(n10609), .IN2(n10605), .IN3(n5396), .IN4(n8721), .Q(
        n10614) );
  OR4X1 U10677 ( .IN1(n10613), .IN2(n10618), .IN3(n9811), .IN4(n8492), .Q(
        n10605) );
  OR2X1 U10678 ( .IN1(n10619), .IN2(n10620), .Q(g33623) );
  AND2X1 U10679 ( .IN1(test_so57), .IN2(n8809), .Q(n10620) );
  AND2X1 U10680 ( .IN1(n10621), .IN2(n10622), .Q(n10619) );
  OR2X1 U10681 ( .IN1(n10623), .IN2(n10624), .Q(n10621) );
  AND2X1 U10682 ( .IN1(n10625), .IN2(n10626), .Q(n10624) );
  AND2X1 U10683 ( .IN1(n10627), .IN2(n8690), .Q(n10623) );
  OR2X1 U10684 ( .IN1(n10628), .IN2(n10629), .Q(n10627) );
  AND2X1 U10685 ( .IN1(n10630), .IN2(g5990), .Q(n10628) );
  OR3X1 U10686 ( .IN1(n10631), .IN2(n10632), .IN3(n10633), .Q(g33622) );
  AND2X1 U10687 ( .IN1(n10634), .IN2(test_so57), .Q(n10633) );
  AND2X1 U10688 ( .IN1(test_so50), .IN2(n8809), .Q(n10632) );
  AND4X1 U10689 ( .IN1(n10622), .IN2(n8503), .IN3(n10626), .IN4(n8721), .Q(
        n10631) );
  OR4X1 U10690 ( .IN1(n10618), .IN2(n10630), .IN3(test_so81), .IN4(n9811), .Q(
        n10622) );
  OR2X1 U10691 ( .IN1(n10635), .IN2(n10636), .Q(g33621) );
  AND2X1 U10692 ( .IN1(n8825), .IN2(g5703), .Q(n10636) );
  AND2X1 U10693 ( .IN1(n10637), .IN2(n10638), .Q(n10635) );
  OR2X1 U10694 ( .IN1(n10639), .IN2(n10640), .Q(n10637) );
  AND2X1 U10695 ( .IN1(n10641), .IN2(n10642), .Q(n10640) );
  AND2X1 U10696 ( .IN1(n10643), .IN2(n8691), .Q(n10639) );
  OR2X1 U10697 ( .IN1(n10644), .IN2(n10645), .Q(n10643) );
  AND2X1 U10698 ( .IN1(n10646), .IN2(g5644), .Q(n10644) );
  OR3X1 U10699 ( .IN1(n10647), .IN2(n10648), .IN3(n10649), .Q(g33620) );
  AND2X1 U10700 ( .IN1(n10650), .IN2(g5703), .Q(n10649) );
  AND2X1 U10701 ( .IN1(n8825), .IN2(g5698), .Q(n10648) );
  AND4X1 U10702 ( .IN1(n10642), .IN2(n10638), .IN3(n5397), .IN4(n8721), .Q(
        n10647) );
  OR4X1 U10703 ( .IN1(n10601), .IN2(n10646), .IN3(n9811), .IN4(n8492), .Q(
        n10638) );
  OR2X1 U10704 ( .IN1(n10651), .IN2(n10652), .Q(g33619) );
  AND2X1 U10705 ( .IN1(n8825), .IN2(g5357), .Q(n10652) );
  AND2X1 U10706 ( .IN1(n10653), .IN2(n10654), .Q(n10651) );
  OR2X1 U10707 ( .IN1(n10655), .IN2(n10656), .Q(n10653) );
  AND2X1 U10708 ( .IN1(n8997), .IN2(g33959), .Q(n10656) );
  AND2X1 U10709 ( .IN1(n10657), .IN2(n8691), .Q(n10655) );
  OR2X1 U10710 ( .IN1(n10658), .IN2(n8996), .Q(n10657) );
  AND2X1 U10711 ( .IN1(n8474), .IN2(g5297), .Q(n10658) );
  OR3X1 U10712 ( .IN1(n10659), .IN2(n10660), .IN3(n10661), .Q(g33618) );
  AND2X1 U10713 ( .IN1(n10662), .IN2(g5357), .Q(n10661) );
  AND2X1 U10714 ( .IN1(n8825), .IN2(g5352), .Q(n10660) );
  AND4X1 U10715 ( .IN1(n10654), .IN2(g33959), .IN3(n5393), .IN4(n8722), .Q(
        n10659) );
  OR4X1 U10716 ( .IN1(n9811), .IN2(n10601), .IN3(test_so81), .IN4(n8474), .Q(
        n10654) );
  OR2X1 U10717 ( .IN1(n10663), .IN2(g4311), .Q(n9811) );
  OR2X1 U10718 ( .IN1(n10664), .IN2(n10665), .Q(g33617) );
  AND2X1 U10719 ( .IN1(n10061), .IN2(n8691), .Q(n10665) );
  OR2X1 U10720 ( .IN1(n10666), .IN2(n10667), .Q(n10061) );
  AND2X1 U10721 ( .IN1(n10668), .IN2(g4581), .Q(n10667) );
  OR2X1 U10722 ( .IN1(n9397), .IN2(g4575), .Q(n10668) );
  AND2X1 U10723 ( .IN1(n5670), .IN2(g4552), .Q(n10666) );
  AND2X1 U10724 ( .IN1(n8825), .IN2(g4552), .Q(n10664) );
  OR2X1 U10725 ( .IN1(n10669), .IN2(n10670), .Q(g33616) );
  AND2X1 U10726 ( .IN1(n10055), .IN2(n8691), .Q(n10670) );
  OR2X1 U10727 ( .IN1(n10671), .IN2(n10672), .Q(n10055) );
  AND2X1 U10728 ( .IN1(n10673), .IN2(g4581), .Q(n10672) );
  OR2X1 U10729 ( .IN1(test_so100), .IN2(n9397), .Q(n10673) );
  AND2X1 U10730 ( .IN1(n5670), .IN2(g4512), .Q(n10671) );
  AND2X1 U10731 ( .IN1(n8825), .IN2(g4515), .Q(n10669) );
  OR2X1 U10732 ( .IN1(n10674), .IN2(n10675), .Q(g33614) );
  AND2X1 U10733 ( .IN1(n8825), .IN2(g4054), .Q(n10675) );
  AND2X1 U10734 ( .IN1(n10676), .IN2(n10677), .Q(n10674) );
  OR2X1 U10735 ( .IN1(n10678), .IN2(n10679), .Q(n10676) );
  AND2X1 U10736 ( .IN1(n10680), .IN2(n10681), .Q(n10679) );
  AND2X1 U10737 ( .IN1(n10682), .IN2(n8691), .Q(n10678) );
  OR2X1 U10738 ( .IN1(n10683), .IN2(n10684), .Q(n10682) );
  AND2X1 U10739 ( .IN1(n10685), .IN2(g3990), .Q(n10683) );
  OR3X1 U10740 ( .IN1(n10686), .IN2(n10687), .IN3(n10688), .Q(g33613) );
  AND2X1 U10741 ( .IN1(n10689), .IN2(g4054), .Q(n10688) );
  AND2X1 U10742 ( .IN1(n8825), .IN2(g4049), .Q(n10687) );
  AND4X1 U10743 ( .IN1(n10681), .IN2(n10677), .IN3(n5395), .IN4(n8722), .Q(
        n10686) );
  OR4X1 U10744 ( .IN1(n10618), .IN2(n10685), .IN3(n9810), .IN4(n8492), .Q(
        n10677) );
  OR2X1 U10745 ( .IN1(n10690), .IN2(n10691), .Q(g33612) );
  AND2X1 U10746 ( .IN1(n8825), .IN2(g3703), .Q(n10691) );
  AND2X1 U10747 ( .IN1(n10692), .IN2(n10693), .Q(n10690) );
  OR2X1 U10748 ( .IN1(n10694), .IN2(n10695), .Q(n10692) );
  AND2X1 U10749 ( .IN1(n10696), .IN2(n10697), .Q(n10695) );
  AND2X1 U10750 ( .IN1(n10698), .IN2(n8691), .Q(n10694) );
  OR2X1 U10751 ( .IN1(n10699), .IN2(n10700), .Q(n10698) );
  AND2X1 U10752 ( .IN1(n10701), .IN2(g3639), .Q(n10699) );
  OR3X1 U10753 ( .IN1(n10702), .IN2(n10703), .IN3(n10704), .Q(g33611) );
  AND2X1 U10754 ( .IN1(n10705), .IN2(g3703), .Q(n10704) );
  AND2X1 U10755 ( .IN1(n8825), .IN2(g3698), .Q(n10703) );
  AND4X1 U10756 ( .IN1(n10697), .IN2(n10693), .IN3(n5399), .IN4(n8721), .Q(
        n10702) );
  OR4X1 U10757 ( .IN1(n10618), .IN2(n10701), .IN3(test_so81), .IN4(n9810), .Q(
        n10693) );
  INVX0 U10758 ( .INP(n3033), .ZN(n10618) );
  OR2X1 U10759 ( .IN1(n10706), .IN2(n10707), .Q(g33610) );
  AND3X1 U10760 ( .IN1(n10708), .IN2(n10709), .IN3(n8745), .Q(n10707) );
  OR3X1 U10761 ( .IN1(n10710), .IN2(n10711), .IN3(n10712), .Q(n10708) );
  AND2X1 U10762 ( .IN1(n10713), .IN2(g3288), .Q(n10711) );
  AND2X1 U10763 ( .IN1(n10714), .IN2(n10715), .Q(n10710) );
  AND2X1 U10764 ( .IN1(n8826), .IN2(g3352), .Q(n10706) );
  OR3X1 U10765 ( .IN1(n10716), .IN2(n10717), .IN3(n10718), .Q(g33609) );
  AND2X1 U10766 ( .IN1(n10719), .IN2(g3352), .Q(n10718) );
  AND2X1 U10767 ( .IN1(n8826), .IN2(g3347), .Q(n10717) );
  AND4X1 U10768 ( .IN1(n10715), .IN2(n10709), .IN3(n5604), .IN4(n8722), .Q(
        n10716) );
  OR4X1 U10769 ( .IN1(n10601), .IN2(n10713), .IN3(n9810), .IN4(n8492), .Q(
        n10709) );
  OR2X1 U10770 ( .IN1(n5323), .IN2(n10663), .Q(n9810) );
  OR2X1 U10771 ( .IN1(n9418), .IN2(n10720), .Q(n10663) );
  XOR2X1 U10772 ( .IN1(n10721), .IN2(n5540), .Q(n10720) );
  XOR2X1 U10773 ( .IN1(n10536), .IN2(n5506), .Q(n9418) );
  INVX0 U10774 ( .INP(g72), .ZN(n10536) );
  INVX0 U10775 ( .INP(n3023), .ZN(n10601) );
  OR4X1 U10776 ( .IN1(n2787), .IN2(n10722), .IN3(n10723), .IN4(n10724), .Q(
        g33608) );
  AND2X1 U10777 ( .IN1(test_so30), .IN2(n8809), .Q(n10724) );
  AND3X1 U10778 ( .IN1(n10725), .IN2(g2759), .IN3(n8745), .Q(n10723) );
  INVX0 U10779 ( .INP(n10067), .ZN(n10725) );
  AND2X1 U10780 ( .IN1(n10067), .IN2(n8463), .Q(n10722) );
  AND2X1 U10781 ( .IN1(test_so30), .IN2(n2790), .Q(n10067) );
  INVX0 U10782 ( .INP(n10726), .ZN(g33607) );
  AND3X1 U10783 ( .IN1(n10727), .IN2(n10728), .IN3(n10729), .Q(n10726) );
  OR2X1 U10784 ( .IN1(n5351), .IN2(n8677), .Q(n10729) );
  OR3X1 U10785 ( .IN1(n10730), .IN2(n10731), .IN3(n10732), .Q(n10728) );
  AND2X1 U10786 ( .IN1(n10733), .IN2(n10734), .Q(n10731) );
  OR4X1 U10787 ( .IN1(n9752), .IN2(g2599), .IN3(n5521), .IN4(n915), .Q(n10734)
         );
  INVX0 U10788 ( .INP(n9852), .ZN(n915) );
  AND3X1 U10789 ( .IN1(g518), .IN2(n3116), .IN3(n5519), .Q(n9852) );
  OR2X1 U10790 ( .IN1(n8797), .IN2(n10735), .Q(n10733) );
  AND3X1 U10791 ( .IN1(g2629), .IN2(g112), .IN3(n5524), .Q(n10730) );
  OR2X1 U10792 ( .IN1(n5311), .IN2(n10736), .Q(n10727) );
  AND2X1 U10793 ( .IN1(n10737), .IN2(n10738), .Q(n10736) );
  OR2X1 U10794 ( .IN1(n3105), .IN2(n8794), .Q(n10738) );
  OR3X1 U10795 ( .IN1(n10739), .IN2(n10740), .IN3(n10741), .Q(g33606) );
  AND2X1 U10796 ( .IN1(n10071), .IN2(g2675), .Q(n10741) );
  AND2X1 U10797 ( .IN1(n8826), .IN2(g2671), .Q(n10740) );
  AND3X1 U10798 ( .IN1(n5457), .IN2(n10072), .IN3(n8745), .Q(n10739) );
  OR3X1 U10799 ( .IN1(n10742), .IN2(n10743), .IN3(n10744), .Q(g33605) );
  AND2X1 U10800 ( .IN1(n10071), .IN2(g2671), .Q(n10744) );
  AND4X1 U10801 ( .IN1(n10072), .IN2(n8752), .IN3(n5418), .IN4(n8530), .Q(
        n10743) );
  AND2X1 U10802 ( .IN1(test_so48), .IN2(n10745), .Q(n10742) );
  OR2X1 U10803 ( .IN1(n8796), .IN2(n10746), .Q(n10745) );
  AND2X1 U10804 ( .IN1(n10072), .IN2(g2661), .Q(n10746) );
  OR2X1 U10805 ( .IN1(n10747), .IN2(n10748), .Q(g33604) );
  AND2X1 U10806 ( .IN1(n10749), .IN2(g2661), .Q(n10748) );
  AND2X1 U10807 ( .IN1(test_so48), .IN2(n10071), .Q(n10747) );
  OR2X1 U10808 ( .IN1(n10750), .IN2(n10751), .Q(g33603) );
  AND2X1 U10809 ( .IN1(n10749), .IN2(g2643), .Q(n10751) );
  AND2X1 U10810 ( .IN1(n10071), .IN2(g2648), .Q(n10750) );
  INVX0 U10811 ( .INP(n10749), .ZN(n10071) );
  OR2X1 U10812 ( .IN1(n8796), .IN2(n10072), .Q(n10749) );
  AND3X1 U10813 ( .IN1(n10086), .IN2(n5351), .IN3(n5521), .Q(n10072) );
  OR2X1 U10814 ( .IN1(n10752), .IN2(n10753), .Q(g33602) );
  AND2X1 U10815 ( .IN1(n10754), .IN2(g2629), .Q(n10753) );
  AND2X1 U10816 ( .IN1(n10755), .IN2(g2599), .Q(n10752) );
  OR2X1 U10817 ( .IN1(n8797), .IN2(n10756), .Q(n10755) );
  AND2X1 U10818 ( .IN1(n10086), .IN2(n10735), .Q(n10756) );
  OR3X1 U10819 ( .IN1(n10757), .IN2(n10758), .IN3(n10759), .Q(g33601) );
  AND2X1 U10820 ( .IN1(n10754), .IN2(g2599), .Q(n10759) );
  AND4X1 U10821 ( .IN1(n10735), .IN2(g2555), .IN3(n10086), .IN4(n8722), .Q(
        n10758) );
  AND2X1 U10822 ( .IN1(n8826), .IN2(g2606), .Q(n10757) );
  OR2X1 U10823 ( .IN1(n10760), .IN2(n10761), .Q(g33600) );
  AND2X1 U10824 ( .IN1(n10754), .IN2(g2555), .Q(n10761) );
  AND2X1 U10825 ( .IN1(n8707), .IN2(n10081), .Q(n10754) );
  INVX0 U10826 ( .INP(n10086), .ZN(n10081) );
  AND4X1 U10827 ( .IN1(n5521), .IN2(n10762), .IN3(n8721), .IN4(n10735), .Q(
        n10760) );
  INVX0 U10828 ( .INP(n3111), .ZN(n10735) );
  OR2X1 U10829 ( .IN1(n10097), .IN2(g2555), .Q(n10762) );
  AND2X1 U10830 ( .IN1(n10086), .IN2(n5524), .Q(n10097) );
  OR2X1 U10831 ( .IN1(n645), .IN2(n10091), .Q(n10086) );
  OR3X1 U10832 ( .IN1(n10763), .IN2(n10764), .IN3(n10765), .Q(n10091) );
  AND2X1 U10833 ( .IN1(n2549), .IN2(g1300), .Q(n10765) );
  AND3X1 U10834 ( .IN1(g2689), .IN2(g2704), .IN3(g2697), .Q(n10764) );
  INVX0 U10835 ( .INP(n10732), .ZN(n645) );
  OR2X1 U10836 ( .IN1(n10766), .IN2(n8215), .Q(n10732) );
  AND3X1 U10837 ( .IN1(n10767), .IN2(n8490), .IN3(n5364), .Q(n10766) );
  INVX0 U10838 ( .INP(n10768), .ZN(g33599) );
  AND4X1 U10839 ( .IN1(n495), .IN2(n10769), .IN3(n10770), .IN4(n10771), .Q(
        n10768) );
  OR4X1 U10840 ( .IN1(n10772), .IN2(n10773), .IN3(n10774), .IN4(n8792), .Q(
        n10771) );
  OR2X1 U10841 ( .IN1(n8501), .IN2(n8677), .Q(n10770) );
  OR2X1 U10842 ( .IN1(n10775), .IN2(n5619), .Q(n10769) );
  AND2X1 U10843 ( .IN1(n10776), .IN2(n10737), .Q(n10775) );
  OR2X1 U10844 ( .IN1(n8795), .IN2(n3125), .Q(n10776) );
  OR4X1 U10845 ( .IN1(g2465), .IN2(n9752), .IN3(n10772), .IN4(n10777), .Q(n495) );
  OR3X1 U10846 ( .IN1(n5522), .IN2(n928), .IN3(n10773), .Q(n10777) );
  AND3X1 U10847 ( .IN1(g112), .IN2(g2495), .IN3(n5523), .Q(n10773) );
  INVX0 U10848 ( .INP(n9851), .ZN(n928) );
  AND3X1 U10849 ( .IN1(g504), .IN2(g518), .IN3(n3116), .Q(n9851) );
  OR3X1 U10850 ( .IN1(n10778), .IN2(n10779), .IN3(n10780), .Q(g33598) );
  AND2X1 U10851 ( .IN1(n10129), .IN2(g2541), .Q(n10780) );
  AND2X1 U10852 ( .IN1(n8826), .IN2(g2537), .Q(n10779) );
  AND3X1 U10853 ( .IN1(n5461), .IN2(n10130), .IN3(n8745), .Q(n10778) );
  OR3X1 U10854 ( .IN1(n10781), .IN2(n10782), .IN3(n10783), .Q(g33597) );
  AND2X1 U10855 ( .IN1(n10129), .IN2(g2537), .Q(n10783) );
  AND4X1 U10856 ( .IN1(n10130), .IN2(n8752), .IN3(n5420), .IN4(n5761), .Q(
        n10782) );
  AND2X1 U10857 ( .IN1(n10784), .IN2(g2533), .Q(n10781) );
  OR2X1 U10858 ( .IN1(n8795), .IN2(n10785), .Q(n10784) );
  AND2X1 U10859 ( .IN1(n10130), .IN2(g2527), .Q(n10785) );
  OR2X1 U10860 ( .IN1(n10786), .IN2(n10787), .Q(g33596) );
  AND2X1 U10861 ( .IN1(n10788), .IN2(g2527), .Q(n10787) );
  AND2X1 U10862 ( .IN1(n10129), .IN2(g2533), .Q(n10786) );
  OR2X1 U10863 ( .IN1(n10789), .IN2(n10790), .Q(g33595) );
  AND2X1 U10864 ( .IN1(n10788), .IN2(g2509), .Q(n10790) );
  AND2X1 U10865 ( .IN1(n10129), .IN2(g2514), .Q(n10789) );
  INVX0 U10866 ( .INP(n10788), .ZN(n10129) );
  OR2X1 U10867 ( .IN1(n8795), .IN2(n10130), .Q(n10788) );
  AND3X1 U10868 ( .IN1(n8501), .IN2(n10144), .IN3(n5522), .Q(n10130) );
  OR2X1 U10869 ( .IN1(n10791), .IN2(n10792), .Q(g33594) );
  AND2X1 U10870 ( .IN1(n10793), .IN2(g2495), .Q(n10792) );
  AND2X1 U10871 ( .IN1(n10794), .IN2(g2465), .Q(n10791) );
  OR2X1 U10872 ( .IN1(n8795), .IN2(n10795), .Q(n10794) );
  AND2X1 U10873 ( .IN1(n10144), .IN2(n10774), .Q(n10795) );
  OR3X1 U10874 ( .IN1(n10796), .IN2(n10797), .IN3(n10798), .Q(g33593) );
  AND2X1 U10875 ( .IN1(n10793), .IN2(g2465), .Q(n10798) );
  AND4X1 U10876 ( .IN1(n10144), .IN2(n10774), .IN3(test_so79), .IN4(n8722), 
        .Q(n10797) );
  AND2X1 U10877 ( .IN1(n8826), .IN2(g2472), .Q(n10796) );
  OR2X1 U10878 ( .IN1(n10799), .IN2(n10800), .Q(g33592) );
  AND2X1 U10879 ( .IN1(n10793), .IN2(test_so79), .Q(n10800) );
  AND2X1 U10880 ( .IN1(n8707), .IN2(n10139), .Q(n10793) );
  INVX0 U10881 ( .INP(n10144), .ZN(n10139) );
  AND4X1 U10882 ( .IN1(n5522), .IN2(n10801), .IN3(n8721), .IN4(n10774), .Q(
        n10799) );
  INVX0 U10883 ( .INP(n3131), .ZN(n10774) );
  OR2X1 U10884 ( .IN1(n10155), .IN2(test_so79), .Q(n10801) );
  AND2X1 U10885 ( .IN1(n10144), .IN2(n5523), .Q(n10155) );
  OR2X1 U10886 ( .IN1(n3122), .IN2(n10149), .Q(n10144) );
  OR3X1 U10887 ( .IN1(n10763), .IN2(n10802), .IN3(n10803), .Q(n10149) );
  AND2X1 U10888 ( .IN1(n2549), .IN2(g1472), .Q(n10803) );
  AND3X1 U10889 ( .IN1(g2697), .IN2(g2689), .IN3(n5377), .Q(n10802) );
  INVX0 U10890 ( .INP(n10772), .ZN(n3122) );
  OR2X1 U10891 ( .IN1(n8404), .IN2(n10804), .Q(n10772) );
  AND2X1 U10892 ( .IN1(n10805), .IN2(n10767), .Q(n10804) );
  INVX0 U10893 ( .INP(n10806), .ZN(g33591) );
  AND3X1 U10894 ( .IN1(n10807), .IN2(n10808), .IN3(n10809), .Q(n10806) );
  OR2X1 U10895 ( .IN1(n5353), .IN2(n8677), .Q(n10809) );
  OR3X1 U10896 ( .IN1(n10810), .IN2(n10811), .IN3(n10812), .Q(n10808) );
  AND2X1 U10897 ( .IN1(n10813), .IN2(n10814), .Q(n10811) );
  OR2X1 U10898 ( .IN1(n9752), .IN2(n9859), .Q(n10814) );
  OR3X1 U10899 ( .IN1(n5537), .IN2(n927), .IN3(g2331), .Q(n9859) );
  OR2X1 U10900 ( .IN1(n8798), .IN2(n10815), .Q(n10813) );
  AND3X1 U10901 ( .IN1(g2361), .IN2(g112), .IN3(n5513), .Q(n10810) );
  OR2X1 U10902 ( .IN1(n5310), .IN2(n10816), .Q(n10807) );
  AND2X1 U10903 ( .IN1(n10737), .IN2(n10817), .Q(n10816) );
  OR2X1 U10904 ( .IN1(n3145), .IN2(n8793), .Q(n10817) );
  OR3X1 U10905 ( .IN1(n10818), .IN2(n10819), .IN3(n10820), .Q(g33590) );
  AND2X1 U10906 ( .IN1(n10185), .IN2(g2407), .Q(n10820) );
  AND2X1 U10907 ( .IN1(test_so31), .IN2(n8809), .Q(n10819) );
  AND3X1 U10908 ( .IN1(n5459), .IN2(n10186), .IN3(n8744), .Q(n10818) );
  OR3X1 U10909 ( .IN1(n10821), .IN2(n10822), .IN3(n10823), .Q(g33589) );
  AND2X1 U10910 ( .IN1(test_so31), .IN2(n10185), .Q(n10823) );
  AND4X1 U10911 ( .IN1(n10186), .IN2(n8753), .IN3(n5421), .IN4(n5762), .Q(
        n10822) );
  AND2X1 U10912 ( .IN1(n10824), .IN2(g2399), .Q(n10821) );
  OR2X1 U10913 ( .IN1(n8796), .IN2(n10825), .Q(n10824) );
  AND2X1 U10914 ( .IN1(n10186), .IN2(g2393), .Q(n10825) );
  OR2X1 U10915 ( .IN1(n10826), .IN2(n10827), .Q(g33588) );
  AND2X1 U10916 ( .IN1(n10828), .IN2(g2393), .Q(n10827) );
  AND2X1 U10917 ( .IN1(n10185), .IN2(g2399), .Q(n10826) );
  OR2X1 U10918 ( .IN1(n10829), .IN2(n10830), .Q(g33587) );
  AND2X1 U10919 ( .IN1(n10828), .IN2(g2375), .Q(n10830) );
  AND2X1 U10920 ( .IN1(n10185), .IN2(g2380), .Q(n10829) );
  INVX0 U10921 ( .INP(n10828), .ZN(n10185) );
  OR2X1 U10922 ( .IN1(n8795), .IN2(n10186), .Q(n10828) );
  AND3X1 U10923 ( .IN1(n10200), .IN2(n5353), .IN3(n5537), .Q(n10186) );
  OR2X1 U10924 ( .IN1(n10831), .IN2(n10832), .Q(g33586) );
  AND2X1 U10925 ( .IN1(n10833), .IN2(g2361), .Q(n10832) );
  AND2X1 U10926 ( .IN1(n10834), .IN2(g2331), .Q(n10831) );
  OR2X1 U10927 ( .IN1(n8797), .IN2(n10835), .Q(n10834) );
  AND2X1 U10928 ( .IN1(n10815), .IN2(n10200), .Q(n10835) );
  OR3X1 U10929 ( .IN1(n10836), .IN2(n10837), .IN3(n10838), .Q(g33585) );
  AND2X1 U10930 ( .IN1(n10833), .IN2(g2331), .Q(n10838) );
  AND4X1 U10931 ( .IN1(n10200), .IN2(g2287), .IN3(n10815), .IN4(n8722), .Q(
        n10837) );
  AND2X1 U10932 ( .IN1(n8826), .IN2(g2338), .Q(n10836) );
  OR2X1 U10933 ( .IN1(n10839), .IN2(n10840), .Q(g33584) );
  AND2X1 U10934 ( .IN1(n10833), .IN2(g2287), .Q(n10840) );
  AND2X1 U10935 ( .IN1(n8707), .IN2(n10195), .Q(n10833) );
  INVX0 U10936 ( .INP(n10200), .ZN(n10195) );
  AND4X1 U10937 ( .IN1(n5537), .IN2(n10841), .IN3(n10815), .IN4(n8723), .Q(
        n10839) );
  OR2X1 U10938 ( .IN1(n927), .IN2(n10842), .Q(n10815) );
  OR3X1 U10939 ( .IN1(n5519), .IN2(n10843), .IN3(g518), .Q(n927) );
  OR2X1 U10940 ( .IN1(n10844), .IN2(g2287), .Q(n10841) );
  AND2X1 U10941 ( .IN1(n5513), .IN2(n10200), .Q(n10844) );
  OR2X1 U10942 ( .IN1(n342), .IN2(n10205), .Q(n10200) );
  OR3X1 U10943 ( .IN1(n10763), .IN2(n10845), .IN3(n10846), .Q(n10205) );
  AND2X1 U10944 ( .IN1(n2549), .IN2(g1448), .Q(n10846) );
  AND3X1 U10945 ( .IN1(g2689), .IN2(g2704), .IN3(n5308), .Q(n10845) );
  INVX0 U10946 ( .INP(n10812), .ZN(n342) );
  OR2X1 U10947 ( .IN1(n10847), .IN2(n8403), .Q(n10812) );
  AND2X1 U10948 ( .IN1(n10848), .IN2(n10767), .Q(n10847) );
  INVX0 U10949 ( .INP(n10849), .ZN(g33583) );
  AND3X1 U10950 ( .IN1(n10850), .IN2(n10851), .IN3(n10852), .Q(n10849) );
  OR2X1 U10951 ( .IN1(n5356), .IN2(n8677), .Q(n10852) );
  OR3X1 U10952 ( .IN1(n10853), .IN2(n10854), .IN3(n10855), .Q(n10851) );
  AND2X1 U10953 ( .IN1(n10856), .IN2(n10857), .Q(n10854) );
  OR2X1 U10954 ( .IN1(n9752), .IN2(n9860), .Q(n10857) );
  OR3X1 U10955 ( .IN1(n5538), .IN2(n917), .IN3(g2197), .Q(n9860) );
  OR2X1 U10956 ( .IN1(n8798), .IN2(n10858), .Q(n10856) );
  AND3X1 U10957 ( .IN1(g2227), .IN2(g112), .IN3(n5514), .Q(n10853) );
  OR2X1 U10958 ( .IN1(n5620), .IN2(n10859), .Q(n10850) );
  AND2X1 U10959 ( .IN1(n10737), .IN2(n10860), .Q(n10859) );
  OR2X1 U10960 ( .IN1(n3164), .IN2(n8794), .Q(n10860) );
  OR3X1 U10961 ( .IN1(n10861), .IN2(n10862), .IN3(n10863), .Q(g33582) );
  AND2X1 U10962 ( .IN1(n10241), .IN2(g2273), .Q(n10863) );
  AND2X1 U10963 ( .IN1(n8826), .IN2(g2269), .Q(n10862) );
  AND3X1 U10964 ( .IN1(n5458), .IN2(n10242), .IN3(n8744), .Q(n10861) );
  OR3X1 U10965 ( .IN1(n10864), .IN2(n10865), .IN3(n10866), .Q(g33581) );
  AND2X1 U10966 ( .IN1(n10241), .IN2(g2269), .Q(n10866) );
  AND4X1 U10967 ( .IN1(n10242), .IN2(n8752), .IN3(n5419), .IN4(n8531), .Q(
        n10865) );
  AND2X1 U10968 ( .IN1(test_so62), .IN2(n10867), .Q(n10864) );
  OR2X1 U10969 ( .IN1(n8799), .IN2(n10868), .Q(n10867) );
  AND2X1 U10970 ( .IN1(n10242), .IN2(g2259), .Q(n10868) );
  OR2X1 U10971 ( .IN1(n10869), .IN2(n10870), .Q(g33580) );
  AND2X1 U10972 ( .IN1(n10871), .IN2(g2259), .Q(n10870) );
  AND2X1 U10973 ( .IN1(test_so62), .IN2(n10241), .Q(n10869) );
  OR2X1 U10974 ( .IN1(n10872), .IN2(n10873), .Q(g33579) );
  AND2X1 U10975 ( .IN1(n10871), .IN2(g2241), .Q(n10873) );
  AND2X1 U10976 ( .IN1(n10241), .IN2(g2246), .Q(n10872) );
  INVX0 U10977 ( .INP(n10871), .ZN(n10241) );
  OR2X1 U10978 ( .IN1(n8800), .IN2(n10242), .Q(n10871) );
  AND3X1 U10979 ( .IN1(n10256), .IN2(n5356), .IN3(n5538), .Q(n10242) );
  OR2X1 U10980 ( .IN1(n10874), .IN2(n10875), .Q(g33578) );
  AND2X1 U10981 ( .IN1(n10876), .IN2(g2227), .Q(n10875) );
  AND2X1 U10982 ( .IN1(n10877), .IN2(g2197), .Q(n10874) );
  OR2X1 U10983 ( .IN1(n8801), .IN2(n10878), .Q(n10877) );
  AND2X1 U10984 ( .IN1(n10858), .IN2(n10256), .Q(n10878) );
  OR3X1 U10985 ( .IN1(n10879), .IN2(n10880), .IN3(n10881), .Q(g33577) );
  AND2X1 U10986 ( .IN1(n10876), .IN2(g2197), .Q(n10881) );
  AND4X1 U10987 ( .IN1(n10256), .IN2(g2153), .IN3(n10858), .IN4(n8723), .Q(
        n10880) );
  AND2X1 U10988 ( .IN1(n8826), .IN2(g2204), .Q(n10879) );
  OR2X1 U10989 ( .IN1(n10882), .IN2(n10883), .Q(g33576) );
  AND2X1 U10990 ( .IN1(n10876), .IN2(g2153), .Q(n10883) );
  AND2X1 U10991 ( .IN1(n8708), .IN2(n10251), .Q(n10876) );
  INVX0 U10992 ( .INP(n10256), .ZN(n10251) );
  AND4X1 U10993 ( .IN1(n5538), .IN2(n10884), .IN3(n10858), .IN4(n8722), .Q(
        n10882) );
  OR2X1 U10994 ( .IN1(n917), .IN2(n10842), .Q(n10858) );
  OR3X1 U10995 ( .IN1(n10843), .IN2(g518), .IN3(g504), .Q(n917) );
  INVX0 U10996 ( .INP(n3116), .ZN(n10843) );
  OR2X1 U10997 ( .IN1(n10885), .IN2(g2153), .Q(n10884) );
  AND2X1 U10998 ( .IN1(n5514), .IN2(n10256), .Q(n10885) );
  OR2X1 U10999 ( .IN1(n657), .IN2(n10261), .Q(n10256) );
  OR3X1 U11000 ( .IN1(n10763), .IN2(n10886), .IN3(n10887), .Q(n10261) );
  AND2X1 U11001 ( .IN1(n2549), .IN2(g1478), .Q(n10887) );
  AND3X1 U11002 ( .IN1(n5377), .IN2(g2689), .IN3(n5308), .Q(n10886) );
  INVX0 U11003 ( .INP(n10293), .ZN(n10763) );
  OR2X1 U11004 ( .IN1(n10888), .IN2(g134), .Q(n10293) );
  AND3X1 U11005 ( .IN1(n10889), .IN2(g691), .IN3(n5595), .Q(n10888) );
  INVX0 U11006 ( .INP(n10855), .ZN(n657) );
  OR2X1 U11007 ( .IN1(n10890), .IN2(n8405), .Q(n10855) );
  AND3X1 U11008 ( .IN1(g1514), .IN2(n8490), .IN3(n10767), .Q(n10890) );
  AND4X1 U11009 ( .IN1(n5768), .IN2(n8399), .IN3(test_so68), .IN4(n10891), .Q(
        n10767) );
  AND3X1 U11010 ( .IN1(g1404), .IN2(n5441), .IN3(n5546), .Q(n10891) );
  OR4X1 U11011 ( .IN1(n10892), .IN2(n10893), .IN3(n10894), .IN4(n10895), .Q(
        g33575) );
  INVX0 U11012 ( .INP(n10896), .ZN(n10895) );
  OR4X1 U11013 ( .IN1(n10897), .IN2(n10898), .IN3(n10899), .IN4(n8792), .Q(
        n10896) );
  AND2X1 U11014 ( .IN1(n8826), .IN2(g1996), .Q(n10894) );
  AND2X1 U11015 ( .IN1(n10900), .IN2(g2047), .Q(n10893) );
  OR2X1 U11016 ( .IN1(n10901), .IN2(n10902), .Q(n10900) );
  AND2X1 U11017 ( .IN1(n10903), .IN2(n8692), .Q(n10901) );
  INVX0 U11018 ( .INP(n240), .ZN(n10892) );
  OR4X1 U11019 ( .IN1(g2040), .IN2(n10903), .IN3(n9752), .IN4(n10904), .Q(n240) );
  OR2X1 U11020 ( .IN1(n5535), .IN2(n10898), .Q(n10904) );
  AND3X1 U11021 ( .IN1(g112), .IN2(g2070), .IN3(n5505), .Q(n10898) );
  OR2X1 U11022 ( .IN1(n10897), .IN2(n9841), .Q(n10903) );
  OR3X1 U11023 ( .IN1(n10905), .IN2(n10906), .IN3(n10907), .Q(g33574) );
  AND2X1 U11024 ( .IN1(n10298), .IN2(g2116), .Q(n10907) );
  AND2X1 U11025 ( .IN1(n8826), .IN2(g2112), .Q(n10906) );
  AND3X1 U11026 ( .IN1(n5463), .IN2(n10299), .IN3(n8744), .Q(n10905) );
  OR3X1 U11027 ( .IN1(n10908), .IN2(n10909), .IN3(n10910), .Q(g33573) );
  AND2X1 U11028 ( .IN1(n10298), .IN2(g2112), .Q(n10910) );
  AND4X1 U11029 ( .IN1(n10299), .IN2(n8753), .IN3(n5666), .IN4(n5452), .Q(
        n10909) );
  AND2X1 U11030 ( .IN1(n10911), .IN2(g2108), .Q(n10908) );
  OR2X1 U11031 ( .IN1(n8800), .IN2(n10912), .Q(n10911) );
  AND2X1 U11032 ( .IN1(n10299), .IN2(g2102), .Q(n10912) );
  OR2X1 U11033 ( .IN1(n10913), .IN2(n10914), .Q(g33572) );
  AND2X1 U11034 ( .IN1(n10915), .IN2(g2102), .Q(n10914) );
  AND2X1 U11035 ( .IN1(n10298), .IN2(g2108), .Q(n10913) );
  OR2X1 U11036 ( .IN1(n10916), .IN2(n10917), .Q(g33571) );
  AND2X1 U11037 ( .IN1(n10915), .IN2(g2084), .Q(n10917) );
  AND2X1 U11038 ( .IN1(n10298), .IN2(g2089), .Q(n10916) );
  INVX0 U11039 ( .INP(n10915), .ZN(n10298) );
  OR2X1 U11040 ( .IN1(n8800), .IN2(n10299), .Q(n10915) );
  AND3X1 U11041 ( .IN1(n10313), .IN2(n5355), .IN3(n5535), .Q(n10299) );
  OR2X1 U11042 ( .IN1(n10918), .IN2(n10919), .Q(g33570) );
  AND2X1 U11043 ( .IN1(n10920), .IN2(g2070), .Q(n10919) );
  AND2X1 U11044 ( .IN1(n10921), .IN2(g2040), .Q(n10918) );
  OR2X1 U11045 ( .IN1(n8800), .IN2(n10922), .Q(n10921) );
  AND2X1 U11046 ( .IN1(n10899), .IN2(n10313), .Q(n10922) );
  OR3X1 U11047 ( .IN1(n10923), .IN2(n10924), .IN3(n10925), .Q(g33569) );
  AND2X1 U11048 ( .IN1(n10920), .IN2(g2040), .Q(n10925) );
  AND4X1 U11049 ( .IN1(n10313), .IN2(g1996), .IN3(n10899), .IN4(n8723), .Q(
        n10924) );
  AND2X1 U11050 ( .IN1(n8826), .IN2(g2047), .Q(n10923) );
  OR2X1 U11051 ( .IN1(n10926), .IN2(n10927), .Q(g33568) );
  AND2X1 U11052 ( .IN1(n10920), .IN2(g1996), .Q(n10927) );
  AND2X1 U11053 ( .IN1(n8708), .IN2(n10308), .Q(n10920) );
  AND4X1 U11054 ( .IN1(n5535), .IN2(n10928), .IN3(n10899), .IN4(n8722), .Q(
        n10926) );
  OR2X1 U11055 ( .IN1(n9841), .IN2(n10842), .Q(n10899) );
  INVX0 U11056 ( .INP(n9854), .ZN(n9841) );
  AND3X1 U11057 ( .IN1(g518), .IN2(n5519), .IN3(n3195), .Q(n9854) );
  OR2X1 U11058 ( .IN1(n10929), .IN2(g1996), .Q(n10928) );
  AND2X1 U11059 ( .IN1(n5505), .IN2(n10313), .Q(n10929) );
  INVX0 U11060 ( .INP(n10308), .ZN(n10313) );
  AND2X1 U11061 ( .IN1(n10897), .IN2(n10349), .Q(n10308) );
  INVX0 U11062 ( .INP(n10318), .ZN(n10349) );
  OR3X1 U11063 ( .IN1(n10930), .IN2(n10931), .IN3(n10932), .Q(n10318) );
  AND2X1 U11064 ( .IN1(n5286), .IN2(g956), .Q(n10932) );
  AND3X1 U11065 ( .IN1(g2145), .IN2(g2130), .IN3(g2138), .Q(n10931) );
  OR2X1 U11066 ( .IN1(n10933), .IN2(n8214), .Q(n10897) );
  AND3X1 U11067 ( .IN1(n5363), .IN2(n10934), .IN3(n5599), .Q(n10933) );
  OR3X1 U11068 ( .IN1(n10935), .IN2(n10936), .IN3(n10937), .Q(g33567) );
  AND2X1 U11069 ( .IN1(test_so8), .IN2(n8808), .Q(n10937) );
  AND2X1 U11070 ( .IN1(n10938), .IN2(g1913), .Q(n10936) );
  OR2X1 U11071 ( .IN1(n10939), .IN2(n10902), .Q(n10938) );
  AND2X1 U11072 ( .IN1(n10940), .IN2(n8692), .Q(n10939) );
  OR2X1 U11073 ( .IN1(n9842), .IN2(n10941), .Q(n10940) );
  INVX0 U11074 ( .INP(n10942), .ZN(n9842) );
  AND3X1 U11075 ( .IN1(n10943), .IN2(n10944), .IN3(n10945), .Q(n10935) );
  OR3X1 U11076 ( .IN1(n8342), .IN2(n5534), .IN3(g1906), .Q(n10944) );
  OR2X1 U11077 ( .IN1(n10946), .IN2(n10947), .Q(n10943) );
  AND2X1 U11078 ( .IN1(n10948), .IN2(n8692), .Q(n10947) );
  AND2X1 U11079 ( .IN1(n9856), .IN2(n9736), .Q(n10946) );
  AND3X1 U11080 ( .IN1(g1936), .IN2(n10942), .IN3(n5503), .Q(n9856) );
  OR3X1 U11081 ( .IN1(n10949), .IN2(n10950), .IN3(n10951), .Q(g33566) );
  AND2X1 U11082 ( .IN1(n10356), .IN2(g1982), .Q(n10951) );
  AND2X1 U11083 ( .IN1(n8826), .IN2(g1978), .Q(n10950) );
  AND3X1 U11084 ( .IN1(n5462), .IN2(n10357), .IN3(n8744), .Q(n10949) );
  OR3X1 U11085 ( .IN1(n10952), .IN2(n10953), .IN3(n10954), .Q(g33565) );
  AND2X1 U11086 ( .IN1(n10356), .IN2(g1978), .Q(n10954) );
  AND4X1 U11087 ( .IN1(n10357), .IN2(n8752), .IN3(n5664), .IN4(n5450), .Q(
        n10953) );
  AND2X1 U11088 ( .IN1(n10955), .IN2(g1974), .Q(n10952) );
  OR2X1 U11089 ( .IN1(n8800), .IN2(n10956), .Q(n10955) );
  AND2X1 U11090 ( .IN1(n10357), .IN2(g1968), .Q(n10956) );
  OR2X1 U11091 ( .IN1(n10957), .IN2(n10958), .Q(g33564) );
  AND2X1 U11092 ( .IN1(n10959), .IN2(g1968), .Q(n10958) );
  AND2X1 U11093 ( .IN1(n10356), .IN2(g1974), .Q(n10957) );
  OR2X1 U11094 ( .IN1(n10960), .IN2(n10961), .Q(g33563) );
  AND2X1 U11095 ( .IN1(n10959), .IN2(g1950), .Q(n10961) );
  AND2X1 U11096 ( .IN1(n10356), .IN2(g1955), .Q(n10960) );
  INVX0 U11097 ( .INP(n10959), .ZN(n10356) );
  OR2X1 U11098 ( .IN1(n8799), .IN2(n10357), .Q(n10959) );
  AND3X1 U11099 ( .IN1(n8502), .IN2(n10371), .IN3(n5534), .Q(n10357) );
  OR2X1 U11100 ( .IN1(n10962), .IN2(n10963), .Q(g33562) );
  AND2X1 U11101 ( .IN1(n10964), .IN2(g1936), .Q(n10963) );
  AND2X1 U11102 ( .IN1(n10965), .IN2(g1906), .Q(n10962) );
  OR2X1 U11103 ( .IN1(n8799), .IN2(n10966), .Q(n10965) );
  AND2X1 U11104 ( .IN1(n10967), .IN2(n10371), .Q(n10966) );
  OR3X1 U11105 ( .IN1(n10968), .IN2(n10969), .IN3(n10970), .Q(g33561) );
  AND2X1 U11106 ( .IN1(n10964), .IN2(g1906), .Q(n10970) );
  AND4X1 U11107 ( .IN1(n10967), .IN2(n10371), .IN3(test_so8), .IN4(n8722), .Q(
        n10969) );
  AND2X1 U11108 ( .IN1(n8826), .IN2(g1913), .Q(n10968) );
  OR2X1 U11109 ( .IN1(n10971), .IN2(n10972), .Q(g33560) );
  AND2X1 U11110 ( .IN1(n10964), .IN2(test_so8), .Q(n10972) );
  AND2X1 U11111 ( .IN1(n8709), .IN2(n10366), .Q(n10964) );
  INVX0 U11112 ( .INP(n10371), .ZN(n10366) );
  AND4X1 U11113 ( .IN1(n5534), .IN2(n10973), .IN3(n10967), .IN4(n8722), .Q(
        n10971) );
  INVX0 U11114 ( .INP(n10948), .ZN(n10967) );
  AND2X1 U11115 ( .IN1(n10942), .IN2(n3115), .Q(n10948) );
  AND3X1 U11116 ( .IN1(g504), .IN2(g518), .IN3(n3195), .Q(n10942) );
  OR2X1 U11117 ( .IN1(n10974), .IN2(test_so8), .Q(n10973) );
  AND2X1 U11118 ( .IN1(n5503), .IN2(n10371), .Q(n10974) );
  OR2X1 U11119 ( .IN1(n10945), .IN2(n10376), .Q(n10371) );
  OR3X1 U11120 ( .IN1(n10930), .IN2(n10975), .IN3(n10976), .Q(n10376) );
  AND2X1 U11121 ( .IN1(n5286), .IN2(g1129), .Q(n10976) );
  AND3X1 U11122 ( .IN1(g2138), .IN2(g2130), .IN3(n5307), .Q(n10975) );
  INVX0 U11123 ( .INP(n10941), .ZN(n10945) );
  OR2X1 U11124 ( .IN1(n10977), .IN2(n8368), .Q(n10941) );
  AND3X1 U11125 ( .IN1(g1171), .IN2(g1183), .IN3(n10934), .Q(n10977) );
  OR3X1 U11126 ( .IN1(n10978), .IN2(n10979), .IN3(n10980), .Q(g33559) );
  AND2X1 U11127 ( .IN1(n8826), .IN2(g1728), .Q(n10980) );
  AND2X1 U11128 ( .IN1(n10981), .IN2(g1779), .Q(n10979) );
  OR2X1 U11129 ( .IN1(n10982), .IN2(n10902), .Q(n10981) );
  AND2X1 U11130 ( .IN1(n10983), .IN2(n8692), .Q(n10982) );
  OR2X1 U11131 ( .IN1(n9843), .IN2(n10984), .Q(n10983) );
  INVX0 U11132 ( .INP(n10985), .ZN(n9843) );
  AND3X1 U11133 ( .IN1(n10986), .IN2(n10987), .IN3(n10988), .Q(n10978) );
  OR3X1 U11134 ( .IN1(n8342), .IN2(n5536), .IN3(g1772), .Q(n10987) );
  OR2X1 U11135 ( .IN1(n10989), .IN2(n10990), .Q(n10986) );
  AND2X1 U11136 ( .IN1(n10991), .IN2(n8692), .Q(n10990) );
  AND2X1 U11137 ( .IN1(n9855), .IN2(n9736), .Q(n10989) );
  AND3X1 U11138 ( .IN1(g1802), .IN2(n10985), .IN3(n5504), .Q(n9855) );
  OR3X1 U11139 ( .IN1(n10992), .IN2(n10993), .IN3(n10994), .Q(g33558) );
  AND2X1 U11140 ( .IN1(n10412), .IN2(g1848), .Q(n10994) );
  AND2X1 U11141 ( .IN1(n8826), .IN2(g1844), .Q(n10993) );
  AND3X1 U11142 ( .IN1(n5464), .IN2(n10413), .IN3(n8743), .Q(n10992) );
  OR3X1 U11143 ( .IN1(n10995), .IN2(n10996), .IN3(n10997), .Q(g33557) );
  AND2X1 U11144 ( .IN1(n10412), .IN2(g1844), .Q(n10997) );
  AND4X1 U11145 ( .IN1(n10413), .IN2(n8752), .IN3(n5665), .IN4(n5451), .Q(
        n10996) );
  AND2X1 U11146 ( .IN1(n10998), .IN2(g1840), .Q(n10995) );
  OR2X1 U11147 ( .IN1(n8799), .IN2(n10999), .Q(n10998) );
  AND2X1 U11148 ( .IN1(n10413), .IN2(g1834), .Q(n10999) );
  OR2X1 U11149 ( .IN1(n11000), .IN2(n11001), .Q(g33556) );
  AND2X1 U11150 ( .IN1(n11002), .IN2(g1834), .Q(n11001) );
  AND2X1 U11151 ( .IN1(n10412), .IN2(g1840), .Q(n11000) );
  OR2X1 U11152 ( .IN1(n11003), .IN2(n11004), .Q(g33555) );
  AND2X1 U11153 ( .IN1(n11002), .IN2(g1816), .Q(n11004) );
  AND2X1 U11154 ( .IN1(n10412), .IN2(g1821), .Q(n11003) );
  INVX0 U11155 ( .INP(n11002), .ZN(n10412) );
  OR2X1 U11156 ( .IN1(n8799), .IN2(n10413), .Q(n11002) );
  AND3X1 U11157 ( .IN1(n10427), .IN2(n5352), .IN3(n5536), .Q(n10413) );
  OR2X1 U11158 ( .IN1(n11005), .IN2(n11006), .Q(g33554) );
  AND2X1 U11159 ( .IN1(n11007), .IN2(g1802), .Q(n11006) );
  AND2X1 U11160 ( .IN1(n11008), .IN2(g1772), .Q(n11005) );
  OR2X1 U11161 ( .IN1(n8798), .IN2(n11009), .Q(n11008) );
  AND2X1 U11162 ( .IN1(n11010), .IN2(n10427), .Q(n11009) );
  OR3X1 U11163 ( .IN1(n11011), .IN2(n11012), .IN3(n11013), .Q(g33553) );
  AND2X1 U11164 ( .IN1(n11007), .IN2(g1772), .Q(n11013) );
  AND4X1 U11165 ( .IN1(n10427), .IN2(g1728), .IN3(n11010), .IN4(n8722), .Q(
        n11012) );
  AND2X1 U11166 ( .IN1(n8826), .IN2(g1779), .Q(n11011) );
  OR2X1 U11167 ( .IN1(n11014), .IN2(n11015), .Q(g33552) );
  AND2X1 U11168 ( .IN1(n11007), .IN2(g1728), .Q(n11015) );
  AND2X1 U11169 ( .IN1(n8708), .IN2(n10422), .Q(n11007) );
  INVX0 U11170 ( .INP(n10427), .ZN(n10422) );
  AND4X1 U11171 ( .IN1(n5536), .IN2(n11016), .IN3(n11010), .IN4(n8723), .Q(
        n11014) );
  INVX0 U11172 ( .INP(n10991), .ZN(n11010) );
  AND2X1 U11173 ( .IN1(n10985), .IN2(n3115), .Q(n10991) );
  AND3X1 U11174 ( .IN1(g504), .IN2(n5287), .IN3(n3195), .Q(n10985) );
  OR2X1 U11175 ( .IN1(n11017), .IN2(g1728), .Q(n11016) );
  AND2X1 U11176 ( .IN1(n5504), .IN2(n10427), .Q(n11017) );
  OR2X1 U11177 ( .IN1(n10988), .IN2(n10432), .Q(n10427) );
  OR3X1 U11178 ( .IN1(n10930), .IN2(n11018), .IN3(n11019), .Q(n10432) );
  AND2X1 U11179 ( .IN1(n5286), .IN2(g1105), .Q(n11019) );
  AND3X1 U11180 ( .IN1(g2145), .IN2(g2130), .IN3(n5275), .Q(n11018) );
  INVX0 U11181 ( .INP(n10984), .ZN(n10988) );
  OR2X1 U11182 ( .IN1(n11020), .IN2(n8509), .Q(n10984) );
  AND2X1 U11183 ( .IN1(n11021), .IN2(n10934), .Q(n11020) );
  OR4X1 U11184 ( .IN1(n11022), .IN2(n11023), .IN3(n11024), .IN4(n11025), .Q(
        g33551) );
  AND2X1 U11185 ( .IN1(n11026), .IN2(n8692), .Q(n11025) );
  OR2X1 U11186 ( .IN1(n11027), .IN2(n11028), .Q(n11026) );
  AND2X1 U11187 ( .IN1(test_so75), .IN2(n11029), .Q(n11028) );
  OR2X1 U11188 ( .IN1(n9844), .IN2(n11030), .Q(n11029) );
  INVX0 U11189 ( .INP(n11031), .ZN(n11027) );
  OR3X1 U11190 ( .IN1(n11030), .IN2(n11032), .IN3(n11033), .Q(n11031) );
  AND2X1 U11191 ( .IN1(g112), .IN2(g31862), .Q(n11032) );
  AND2X1 U11192 ( .IN1(n8826), .IN2(g1592), .Q(n11024) );
  AND2X1 U11193 ( .IN1(test_so75), .IN2(n10902), .Q(n11023) );
  AND3X1 U11194 ( .IN1(n8342), .IN2(g33533), .IN3(n11034), .Q(n11022) );
  AND3X1 U11195 ( .IN1(n9853), .IN2(n9736), .IN3(g31862), .Q(n11034) );
  OR3X1 U11196 ( .IN1(n11035), .IN2(n11036), .IN3(n11037), .Q(g33550) );
  AND2X1 U11197 ( .IN1(n10468), .IN2(g1714), .Q(n11037) );
  AND2X1 U11198 ( .IN1(n8826), .IN2(g1710), .Q(n11036) );
  AND3X1 U11199 ( .IN1(n5460), .IN2(n10469), .IN3(n8743), .Q(n11035) );
  OR3X1 U11200 ( .IN1(n11038), .IN2(n11039), .IN3(n11040), .Q(g33549) );
  AND2X1 U11201 ( .IN1(n10468), .IN2(g1710), .Q(n11040) );
  AND4X1 U11202 ( .IN1(n10469), .IN2(n8752), .IN3(n5417), .IN4(n8532), .Q(
        n11039) );
  AND2X1 U11203 ( .IN1(test_so15), .IN2(n11041), .Q(n11038) );
  OR2X1 U11204 ( .IN1(n8797), .IN2(n11042), .Q(n11041) );
  AND2X1 U11205 ( .IN1(n10469), .IN2(g1700), .Q(n11042) );
  OR2X1 U11206 ( .IN1(n11043), .IN2(n11044), .Q(g33548) );
  AND2X1 U11207 ( .IN1(n11045), .IN2(g1700), .Q(n11044) );
  AND2X1 U11208 ( .IN1(test_so15), .IN2(n10468), .Q(n11043) );
  OR2X1 U11209 ( .IN1(n11046), .IN2(n11047), .Q(g33547) );
  AND2X1 U11210 ( .IN1(n11045), .IN2(g1682), .Q(n11047) );
  AND2X1 U11211 ( .IN1(n10468), .IN2(g1687), .Q(n11046) );
  INVX0 U11212 ( .INP(n11045), .ZN(n10468) );
  OR2X1 U11213 ( .IN1(n8797), .IN2(n10469), .Q(n11045) );
  AND3X1 U11214 ( .IN1(n10483), .IN2(n5362), .IN3(n5598), .Q(n10469) );
  OR3X1 U11215 ( .IN1(n11048), .IN2(n11049), .IN3(n11050), .Q(g33546) );
  AND2X1 U11216 ( .IN1(n8826), .IN2(g1636), .Q(n11050) );
  AND2X1 U11217 ( .IN1(n10499), .IN2(n11033), .Q(n11049) );
  AND2X1 U11218 ( .IN1(n10483), .IN2(g1636), .Q(n10499) );
  AND2X1 U11219 ( .IN1(n11051), .IN2(g1668), .Q(n11048) );
  OR3X1 U11220 ( .IN1(n11052), .IN2(n11053), .IN3(n11054), .Q(g33545) );
  AND2X1 U11221 ( .IN1(n11051), .IN2(g1636), .Q(n11054) );
  AND3X1 U11222 ( .IN1(n10505), .IN2(n11033), .IN3(n8743), .Q(n11053) );
  AND2X1 U11223 ( .IN1(n10483), .IN2(g1592), .Q(n10505) );
  AND2X1 U11224 ( .IN1(test_so75), .IN2(n8808), .Q(n11052) );
  OR2X1 U11225 ( .IN1(n11055), .IN2(n11056), .Q(g33544) );
  AND2X1 U11226 ( .IN1(n11051), .IN2(g1592), .Q(n11056) );
  AND2X1 U11227 ( .IN1(n8709), .IN2(n10478), .Q(n11051) );
  INVX0 U11228 ( .INP(n10483), .ZN(n10478) );
  AND4X1 U11229 ( .IN1(n5598), .IN2(n11057), .IN3(n11033), .IN4(n8723), .Q(
        n11055) );
  OR2X1 U11230 ( .IN1(n9844), .IN2(n10842), .Q(n11033) );
  INVX0 U11231 ( .INP(n3115), .ZN(n10842) );
  INVX0 U11232 ( .INP(n9853), .ZN(n9844) );
  AND3X1 U11233 ( .IN1(n5287), .IN2(n5519), .IN3(n3195), .Q(n9853) );
  OR2X1 U11234 ( .IN1(n11058), .IN2(g1592), .Q(n11057) );
  AND2X1 U11235 ( .IN1(n5549), .IN2(n10483), .Q(n11058) );
  OR2X1 U11236 ( .IN1(g33533), .IN2(n10488), .Q(n10483) );
  OR3X1 U11237 ( .IN1(n10930), .IN2(n11059), .IN3(n11060), .Q(n10488) );
  AND2X1 U11238 ( .IN1(n5286), .IN2(g1135), .Q(n11060) );
  AND3X1 U11239 ( .IN1(n5307), .IN2(g2130), .IN3(n5275), .Q(n11059) );
  INVX0 U11240 ( .INP(n10520), .ZN(n10930) );
  OR2X1 U11241 ( .IN1(n11061), .IN2(g134), .Q(n10520) );
  AND3X1 U11242 ( .IN1(n11062), .IN2(g691), .IN3(n5595), .Q(n11061) );
  OR2X1 U11243 ( .IN1(n11063), .IN2(n11064), .Q(g33543) );
  AND2X1 U11244 ( .IN1(n11065), .IN2(g1373), .Q(n11064) );
  OR2X1 U11245 ( .IN1(n8796), .IN2(n11066), .Q(n11065) );
  AND3X1 U11246 ( .IN1(n11067), .IN2(n11068), .IN3(n8467), .Q(n11066) );
  AND3X1 U11247 ( .IN1(n8727), .IN2(g1379), .IN3(n11069), .Q(n11063) );
  OR2X1 U11248 ( .IN1(n11070), .IN2(n11071), .Q(n11069) );
  AND2X1 U11249 ( .IN1(n8328), .IN2(n11068), .Q(n11070) );
  OR3X1 U11250 ( .IN1(n11072), .IN2(n11073), .IN3(n11074), .Q(g33542) );
  AND2X1 U11251 ( .IN1(n8826), .IN2(g1270), .Q(n11074) );
  AND2X1 U11252 ( .IN1(n5730), .IN2(n11075), .Q(n11073) );
  AND3X1 U11253 ( .IN1(n11076), .IN2(n11077), .IN3(g1274), .Q(n11072) );
  OR2X1 U11254 ( .IN1(n11078), .IN2(n11079), .Q(g33541) );
  AND2X1 U11255 ( .IN1(n11080), .IN2(g1030), .Q(n11079) );
  OR2X1 U11256 ( .IN1(n8796), .IN2(n11081), .Q(n11080) );
  AND3X1 U11257 ( .IN1(n11082), .IN2(n11083), .IN3(n8464), .Q(n11081) );
  AND3X1 U11258 ( .IN1(n8726), .IN2(g1036), .IN3(n11084), .Q(n11078) );
  OR2X1 U11259 ( .IN1(n11085), .IN2(n11086), .Q(n11084) );
  AND2X1 U11260 ( .IN1(n8327), .IN2(n11083), .Q(n11085) );
  OR3X1 U11261 ( .IN1(n11087), .IN2(n11088), .IN3(n11089), .Q(g33540) );
  AND2X1 U11262 ( .IN1(n8826), .IN2(g925), .Q(n11089) );
  AND2X1 U11263 ( .IN1(n5731), .IN2(n11090), .Q(n11088) );
  AND3X1 U11264 ( .IN1(n11091), .IN2(n11092), .IN3(g930), .Q(n11087) );
  OR3X1 U11265 ( .IN1(n11093), .IN2(n11094), .IN3(n11095), .Q(g33539) );
  AND2X1 U11266 ( .IN1(n8827), .IN2(g758), .Q(n11095) );
  AND2X1 U11267 ( .IN1(n2980), .IN2(n5332), .Q(n11094) );
  AND3X1 U11268 ( .IN1(n2404), .IN2(n11096), .IN3(g763), .Q(n11093) );
  INVX0 U11269 ( .INP(n2980), .ZN(n11096) );
  OR3X1 U11270 ( .IN1(n11097), .IN2(n11098), .IN3(n11099), .Q(g33538) );
  AND2X1 U11271 ( .IN1(n8827), .IN2(g590), .Q(n11099) );
  AND2X1 U11272 ( .IN1(n2982), .IN2(n5476), .Q(n11098) );
  AND3X1 U11273 ( .IN1(n2421), .IN2(n11100), .IN3(g595), .Q(n11097) );
  INVX0 U11274 ( .INP(n2982), .ZN(n11100) );
  OR2X1 U11275 ( .IN1(n11101), .IN2(n11102), .Q(g33537) );
  AND3X1 U11276 ( .IN1(n2707), .IN2(g142), .IN3(n8743), .Q(n11102) );
  AND2X1 U11277 ( .IN1(n8827), .IN2(g301), .Q(n11101) );
  AND2X1 U11278 ( .IN1(n11103), .IN2(g160), .Q(g33536) );
  OR2X1 U11279 ( .IN1(n2710), .IN2(n8793), .Q(n11103) );
  OR3X1 U11280 ( .IN1(n11104), .IN2(n11105), .IN3(n11106), .Q(g33535) );
  AND2X1 U11281 ( .IN1(n8827), .IN2(g291), .Q(n11106) );
  AND2X1 U11282 ( .IN1(n3276), .IN2(n5680), .Q(n11105) );
  AND3X1 U11283 ( .IN1(n8473), .IN2(n11107), .IN3(g294), .Q(n11104) );
  INVX0 U11284 ( .INP(n3276), .ZN(n11107) );
  OR3X1 U11285 ( .IN1(n11108), .IN2(n11109), .IN3(n11110), .Q(g33534) );
  AND2X1 U11286 ( .IN1(n8827), .IN2(g150), .Q(n11110) );
  AND2X1 U11287 ( .IN1(n3277), .IN2(n5677), .Q(n11109) );
  AND3X1 U11288 ( .IN1(n9969), .IN2(n11111), .IN3(g153), .Q(n11108) );
  INVX0 U11289 ( .INP(n3277), .ZN(n11111) );
  INVX0 U11290 ( .INP(n11030), .ZN(g33533) );
  OR2X1 U11291 ( .IN1(n11112), .IN2(n8369), .Q(n11030) );
  AND3X1 U11292 ( .IN1(n10934), .IN2(g1171), .IN3(n5599), .Q(n11112) );
  AND4X1 U11293 ( .IN1(n5442), .IN2(n5547), .IN3(n8400), .IN4(n11113), .Q(
        n10934) );
  AND3X1 U11294 ( .IN1(n8507), .IN2(g1061), .IN3(g979), .Q(n11113) );
  AND3X1 U11295 ( .IN1(n11114), .IN2(n11115), .IN3(n11116), .Q(g33435) );
  OR2X1 U11296 ( .IN1(n5610), .IN2(n9767), .Q(n11116) );
  OR3X1 U11297 ( .IN1(n11117), .IN2(n11118), .IN3(g2729), .Q(n11115) );
  AND2X1 U11298 ( .IN1(n5544), .IN2(n5301), .Q(n11118) );
  AND2X1 U11299 ( .IN1(n5378), .IN2(g2724), .Q(n11117) );
  OR2X1 U11300 ( .IN1(n5403), .IN2(n9780), .Q(n11114) );
  AND3X1 U11301 ( .IN1(n11119), .IN2(n11120), .IN3(n11121), .Q(g33079) );
  OR2X1 U11302 ( .IN1(n5609), .IN2(n9767), .Q(n11121) );
  OR3X1 U11303 ( .IN1(n11122), .IN2(n11123), .IN3(g2729), .Q(n11120) );
  AND2X1 U11304 ( .IN1(n5545), .IN2(n5301), .Q(n11123) );
  AND2X1 U11305 ( .IN1(n5379), .IN2(g2724), .Q(n11122) );
  OR2X1 U11306 ( .IN1(n5404), .IN2(n9780), .Q(n11119) );
  OR2X1 U11307 ( .IN1(n8347), .IN2(g2724), .Q(n9780) );
  OR2X1 U11308 ( .IN1(n11124), .IN2(n11125), .Q(g33070) );
  AND2X1 U11309 ( .IN1(n8827), .IN2(g6565), .Q(n11125) );
  AND2X1 U11310 ( .IN1(n11126), .IN2(n11127), .Q(n11124) );
  OR3X1 U11311 ( .IN1(n11128), .IN2(n11129), .IN3(n11130), .Q(n11126) );
  AND2X1 U11312 ( .IN1(g25756), .IN2(n5646), .Q(n11130) );
  AND2X1 U11313 ( .IN1(n11131), .IN2(n8693), .Q(n11129) );
  OR2X1 U11314 ( .IN1(n11132), .IN2(n11133), .Q(g33069) );
  AND2X1 U11315 ( .IN1(n11134), .IN2(g6565), .Q(n11133) );
  AND2X1 U11316 ( .IN1(n11135), .IN2(g6561), .Q(n11132) );
  OR2X1 U11317 ( .IN1(n8807), .IN2(n11136), .Q(n11135) );
  AND2X1 U11318 ( .IN1(n5386), .IN2(n11127), .Q(n11136) );
  OR2X1 U11319 ( .IN1(n11137), .IN2(n11138), .Q(g33068) );
  AND2X1 U11320 ( .IN1(n8838), .IN2(g6555), .Q(n11138) );
  AND3X1 U11321 ( .IN1(n11127), .IN2(n11139), .IN3(n5646), .Q(n11137) );
  INVX0 U11322 ( .INP(n704), .ZN(n11139) );
  OR2X1 U11323 ( .IN1(n11140), .IN2(n11141), .Q(g33067) );
  AND2X1 U11324 ( .IN1(n8836), .IN2(g6549), .Q(n11141) );
  AND2X1 U11325 ( .IN1(n11142), .IN2(n11127), .Q(n11140) );
  INVX0 U11326 ( .INP(n11143), .ZN(n11142) );
  AND2X1 U11327 ( .IN1(n11144), .IN2(n3407), .Q(n11143) );
  OR2X1 U11328 ( .IN1(n8806), .IN2(n3406), .Q(n11144) );
  OR2X1 U11329 ( .IN1(n11145), .IN2(n11146), .Q(g33065) );
  AND2X1 U11330 ( .IN1(n8836), .IN2(g6219), .Q(n11146) );
  AND2X1 U11331 ( .IN1(n11147), .IN2(n11148), .Q(n11145) );
  OR3X1 U11332 ( .IN1(n11149), .IN2(n11150), .IN3(n11151), .Q(n11147) );
  AND2X1 U11333 ( .IN1(g25742), .IN2(n5651), .Q(n11151) );
  AND2X1 U11334 ( .IN1(n8709), .IN2(n11152), .Q(n11150) );
  OR2X1 U11335 ( .IN1(n11153), .IN2(n11154), .Q(g33064) );
  AND2X1 U11336 ( .IN1(n11155), .IN2(g6219), .Q(n11154) );
  AND2X1 U11337 ( .IN1(n11156), .IN2(g6215), .Q(n11153) );
  OR2X1 U11338 ( .IN1(n8805), .IN2(n11157), .Q(n11156) );
  AND2X1 U11339 ( .IN1(n5385), .IN2(n11148), .Q(n11157) );
  OR2X1 U11340 ( .IN1(n11158), .IN2(n11159), .Q(g33063) );
  AND2X1 U11341 ( .IN1(n8836), .IN2(g6209), .Q(n11159) );
  AND3X1 U11342 ( .IN1(n11148), .IN2(n11160), .IN3(n5651), .Q(n11158) );
  INVX0 U11343 ( .INP(n952), .ZN(n11160) );
  OR2X1 U11344 ( .IN1(n11161), .IN2(n11162), .Q(g33062) );
  AND2X1 U11345 ( .IN1(n8836), .IN2(g6203), .Q(n11162) );
  AND2X1 U11346 ( .IN1(n11163), .IN2(n11148), .Q(n11161) );
  INVX0 U11347 ( .INP(n11164), .ZN(n11163) );
  AND2X1 U11348 ( .IN1(n11165), .IN2(n3417), .Q(n11164) );
  OR2X1 U11349 ( .IN1(n8805), .IN2(n3416), .Q(n11165) );
  OR2X1 U11350 ( .IN1(n11166), .IN2(n11167), .Q(g33060) );
  AND2X1 U11351 ( .IN1(n8836), .IN2(g5873), .Q(n11167) );
  AND2X1 U11352 ( .IN1(n11168), .IN2(n11169), .Q(n11166) );
  OR3X1 U11353 ( .IN1(n11170), .IN2(n11171), .IN3(n11172), .Q(n11168) );
  AND2X1 U11354 ( .IN1(g25728), .IN2(n5649), .Q(n11172) );
  AND2X1 U11355 ( .IN1(n8709), .IN2(n11173), .Q(n11171) );
  OR2X1 U11356 ( .IN1(n11174), .IN2(n11175), .Q(g33059) );
  AND2X1 U11357 ( .IN1(n11176), .IN2(g5873), .Q(n11175) );
  AND2X1 U11358 ( .IN1(n11177), .IN2(g5869), .Q(n11174) );
  OR2X1 U11359 ( .IN1(n8805), .IN2(n11178), .Q(n11177) );
  AND2X1 U11360 ( .IN1(n5388), .IN2(n11169), .Q(n11178) );
  OR2X1 U11361 ( .IN1(n11179), .IN2(n11180), .Q(g33058) );
  AND2X1 U11362 ( .IN1(n8836), .IN2(g5863), .Q(n11180) );
  AND3X1 U11363 ( .IN1(n11169), .IN2(n11181), .IN3(n5649), .Q(n11179) );
  INVX0 U11364 ( .INP(n1011), .ZN(n11181) );
  OR2X1 U11365 ( .IN1(n11182), .IN2(n11183), .Q(g33057) );
  AND2X1 U11366 ( .IN1(n8836), .IN2(g5857), .Q(n11183) );
  AND2X1 U11367 ( .IN1(n11184), .IN2(n11169), .Q(n11182) );
  INVX0 U11368 ( .INP(n11185), .ZN(n11184) );
  AND2X1 U11369 ( .IN1(n11186), .IN2(n3427), .Q(n11185) );
  OR2X1 U11370 ( .IN1(n8804), .IN2(n3426), .Q(n11186) );
  OR2X1 U11371 ( .IN1(n11187), .IN2(n11188), .Q(g33055) );
  AND2X1 U11372 ( .IN1(n8836), .IN2(g5527), .Q(n11188) );
  AND2X1 U11373 ( .IN1(n11189), .IN2(n11190), .Q(n11187) );
  OR3X1 U11374 ( .IN1(n11191), .IN2(n11192), .IN3(n11193), .Q(n11189) );
  AND2X1 U11375 ( .IN1(g25714), .IN2(n5647), .Q(n11193) );
  AND2X1 U11376 ( .IN1(n8709), .IN2(n11194), .Q(n11192) );
  OR2X1 U11377 ( .IN1(n11195), .IN2(n11196), .Q(g33054) );
  AND2X1 U11378 ( .IN1(n11197), .IN2(g5527), .Q(n11196) );
  AND2X1 U11379 ( .IN1(n11198), .IN2(g5523), .Q(n11195) );
  OR2X1 U11380 ( .IN1(n8804), .IN2(n11199), .Q(n11198) );
  AND2X1 U11381 ( .IN1(n5389), .IN2(n11190), .Q(n11199) );
  OR2X1 U11382 ( .IN1(n11200), .IN2(n11201), .Q(g33053) );
  AND2X1 U11383 ( .IN1(n8837), .IN2(g5517), .Q(n11201) );
  AND3X1 U11384 ( .IN1(n11190), .IN2(n11202), .IN3(n5647), .Q(n11200) );
  INVX0 U11385 ( .INP(n473), .ZN(n11202) );
  OR2X1 U11386 ( .IN1(n11203), .IN2(n11204), .Q(g33052) );
  AND2X1 U11387 ( .IN1(n8837), .IN2(g5511), .Q(n11204) );
  AND2X1 U11388 ( .IN1(n11205), .IN2(n11190), .Q(n11203) );
  INVX0 U11389 ( .INP(n11206), .ZN(n11205) );
  AND2X1 U11390 ( .IN1(n11207), .IN2(n3437), .Q(n11206) );
  OR2X1 U11391 ( .IN1(n8803), .IN2(n3436), .Q(n11207) );
  OR2X1 U11392 ( .IN1(n11208), .IN2(n11209), .Q(g33050) );
  AND2X1 U11393 ( .IN1(n8837), .IN2(g5180), .Q(n11209) );
  AND2X1 U11394 ( .IN1(n11210), .IN2(n11211), .Q(n11208) );
  OR3X1 U11395 ( .IN1(n11212), .IN2(n11213), .IN3(n11214), .Q(n11210) );
  AND2X1 U11396 ( .IN1(g25700), .IN2(n5650), .Q(n11214) );
  AND2X1 U11397 ( .IN1(n8710), .IN2(n11215), .Q(n11213) );
  OR2X1 U11398 ( .IN1(n11216), .IN2(n11217), .Q(g33049) );
  AND2X1 U11399 ( .IN1(n11218), .IN2(g5180), .Q(n11217) );
  AND2X1 U11400 ( .IN1(n11219), .IN2(g5176), .Q(n11216) );
  OR2X1 U11401 ( .IN1(n8803), .IN2(n11220), .Q(n11219) );
  AND2X1 U11402 ( .IN1(n5384), .IN2(n11211), .Q(n11220) );
  OR2X1 U11403 ( .IN1(n11221), .IN2(n11222), .Q(g33048) );
  AND2X1 U11404 ( .IN1(n8837), .IN2(g5170), .Q(n11222) );
  AND3X1 U11405 ( .IN1(n11211), .IN2(n11223), .IN3(n5650), .Q(n11221) );
  INVX0 U11406 ( .INP(n699), .ZN(n11223) );
  OR2X1 U11407 ( .IN1(n11224), .IN2(n11225), .Q(g33047) );
  AND2X1 U11408 ( .IN1(n8837), .IN2(g5164), .Q(n11225) );
  AND2X1 U11409 ( .IN1(n11226), .IN2(n11211), .Q(n11224) );
  INVX0 U11410 ( .INP(n11227), .ZN(n11226) );
  AND2X1 U11411 ( .IN1(n11228), .IN2(n3447), .Q(n11227) );
  OR2X1 U11412 ( .IN1(n8803), .IN2(n3446), .Q(n11228) );
  OR3X1 U11413 ( .IN1(n11229), .IN2(n11230), .IN3(n11231), .Q(g33046) );
  AND2X1 U11414 ( .IN1(n8837), .IN2(g5052), .Q(n11231) );
  AND3X1 U11415 ( .IN1(n11232), .IN2(n11233), .IN3(g5057), .Q(n11230) );
  INVX0 U11416 ( .INP(n11234), .ZN(n11233) );
  AND2X1 U11417 ( .IN1(n5615), .IN2(n11235), .Q(n11229) );
  OR2X1 U11418 ( .IN1(n11234), .IN2(n11236), .Q(n11235) );
  AND2X1 U11419 ( .IN1(g5052), .IN2(n11237), .Q(n11234) );
  OR3X1 U11420 ( .IN1(n11238), .IN2(n11239), .IN3(n11240), .Q(g33045) );
  AND2X1 U11421 ( .IN1(n11241), .IN2(g4567), .Q(n11240) );
  OR3X1 U11422 ( .IN1(n11242), .IN2(n11243), .IN3(n11239), .Q(g33044) );
  AND2X1 U11423 ( .IN1(test_so93), .IN2(n11241), .Q(n11242) );
  OR3X1 U11424 ( .IN1(n11244), .IN2(n11245), .IN3(n11246), .Q(g33043) );
  AND2X1 U11425 ( .IN1(test_so16), .IN2(n11241), .Q(n11246) );
  OR3X1 U11426 ( .IN1(n11244), .IN2(n11239), .IN3(n11247), .Q(g33042) );
  AND2X1 U11427 ( .IN1(n11241), .IN2(g4540), .Q(n11247) );
  INVX0 U11428 ( .INP(n11248), .ZN(n11239) );
  OR2X1 U11429 ( .IN1(n8445), .IN2(n11241), .Q(n11248) );
  OR3X1 U11430 ( .IN1(n11238), .IN2(n11245), .IN3(n11249), .Q(g33041) );
  AND2X1 U11431 ( .IN1(test_so56), .IN2(n11241), .Q(n11249) );
  OR3X1 U11432 ( .IN1(n11250), .IN2(n11243), .IN3(n11251), .Q(g33040) );
  AND2X1 U11433 ( .IN1(n11252), .IN2(n9397), .Q(n11243) );
  OR2X1 U11434 ( .IN1(g72), .IN2(g73), .Q(n9397) );
  AND2X1 U11435 ( .IN1(n11241), .IN2(g4504), .Q(n11250) );
  OR3X1 U11436 ( .IN1(n11238), .IN2(n11253), .IN3(n11254), .Q(g33039) );
  AND2X1 U11437 ( .IN1(n11241), .IN2(g4501), .Q(n11254) );
  OR3X1 U11438 ( .IN1(n11238), .IN2(n11251), .IN3(n11255), .Q(g33038) );
  AND2X1 U11439 ( .IN1(n11241), .IN2(g4498), .Q(n11255) );
  AND2X1 U11440 ( .IN1(n11256), .IN2(n11252), .Q(n11238) );
  OR2X1 U11441 ( .IN1(n11257), .IN2(g73), .Q(n11256) );
  OR3X1 U11442 ( .IN1(n11244), .IN2(n11253), .IN3(n11258), .Q(g33037) );
  AND2X1 U11443 ( .IN1(n11241), .IN2(g4495), .Q(n11258) );
  OR3X1 U11444 ( .IN1(n11244), .IN2(n11251), .IN3(n11259), .Q(g33036) );
  AND2X1 U11445 ( .IN1(n11241), .IN2(g4480), .Q(n11259) );
  AND2X1 U11446 ( .IN1(g4572), .IN2(n11252), .Q(n11251) );
  AND2X1 U11447 ( .IN1(n11260), .IN2(n11252), .Q(n11244) );
  OR2X1 U11448 ( .IN1(n10721), .IN2(g72), .Q(n11260) );
  OR4X1 U11449 ( .IN1(n8481), .IN2(n11261), .IN3(n11262), .IN4(n11263), .Q(
        g33035) );
  AND2X1 U11450 ( .IN1(n8837), .IN2(g4098), .Q(n11263) );
  AND3X1 U11451 ( .IN1(n9086), .IN2(g4108), .IN3(n8742), .Q(n11262) );
  AND2X1 U11452 ( .IN1(n9092), .IN2(n5715), .Q(n11261) );
  INVX0 U11453 ( .INP(n9086), .ZN(n9092) );
  OR2X1 U11454 ( .IN1(n5350), .IN2(n11264), .Q(n9086) );
  OR2X1 U11455 ( .IN1(n11265), .IN2(n11266), .Q(g33034) );
  AND2X1 U11456 ( .IN1(n8837), .IN2(g3873), .Q(n11266) );
  AND2X1 U11457 ( .IN1(n11267), .IN2(n11268), .Q(n11265) );
  OR3X1 U11458 ( .IN1(n11269), .IN2(n11270), .IN3(n11271), .Q(n11267) );
  AND2X1 U11459 ( .IN1(g25676), .IN2(n8493), .Q(n11271) );
  AND2X1 U11460 ( .IN1(n8710), .IN2(n11272), .Q(n11270) );
  OR2X1 U11461 ( .IN1(n11273), .IN2(n11274), .Q(g33033) );
  AND2X1 U11462 ( .IN1(n11275), .IN2(g3873), .Q(n11274) );
  AND2X1 U11463 ( .IN1(test_so33), .IN2(n11276), .Q(n11273) );
  OR2X1 U11464 ( .IN1(n8803), .IN2(n11277), .Q(n11276) );
  AND2X1 U11465 ( .IN1(n5387), .IN2(n11268), .Q(n11277) );
  OR2X1 U11466 ( .IN1(n11278), .IN2(n11279), .Q(g33032) );
  AND2X1 U11467 ( .IN1(n8837), .IN2(g3863), .Q(n11279) );
  AND3X1 U11468 ( .IN1(n11280), .IN2(n8493), .IN3(n11268), .Q(n11278) );
  INVX0 U11469 ( .INP(n1069), .ZN(n11280) );
  OR2X1 U11470 ( .IN1(n11281), .IN2(n11282), .Q(g33031) );
  AND2X1 U11471 ( .IN1(n8837), .IN2(g3857), .Q(n11282) );
  AND2X1 U11472 ( .IN1(n11283), .IN2(n11268), .Q(n11281) );
  INVX0 U11473 ( .INP(n11284), .ZN(n11283) );
  AND2X1 U11474 ( .IN1(n11285), .IN2(n3482), .Q(n11284) );
  OR2X1 U11475 ( .IN1(n8803), .IN2(n3481), .Q(n11285) );
  OR2X1 U11476 ( .IN1(n11286), .IN2(n11287), .Q(g33029) );
  AND2X1 U11477 ( .IN1(n8837), .IN2(g3522), .Q(n11287) );
  AND2X1 U11478 ( .IN1(n11288), .IN2(n11289), .Q(n11286) );
  OR3X1 U11479 ( .IN1(n11290), .IN2(n11291), .IN3(n11292), .Q(n11288) );
  AND2X1 U11480 ( .IN1(g25662), .IN2(n5645), .Q(n11292) );
  AND2X1 U11481 ( .IN1(n8710), .IN2(n11293), .Q(n11291) );
  OR2X1 U11482 ( .IN1(n11294), .IN2(n11295), .Q(g33028) );
  AND2X1 U11483 ( .IN1(n11296), .IN2(g3522), .Q(n11295) );
  AND2X1 U11484 ( .IN1(n11297), .IN2(g3518), .Q(n11294) );
  OR2X1 U11485 ( .IN1(n8802), .IN2(n11298), .Q(n11297) );
  AND2X1 U11486 ( .IN1(n5383), .IN2(n11289), .Q(n11298) );
  OR2X1 U11487 ( .IN1(n11299), .IN2(n11300), .Q(g33027) );
  AND2X1 U11488 ( .IN1(n8837), .IN2(g3512), .Q(n11300) );
  AND3X1 U11489 ( .IN1(n11289), .IN2(n11301), .IN3(n5645), .Q(n11299) );
  INVX0 U11490 ( .INP(n94), .ZN(n11301) );
  OR2X1 U11491 ( .IN1(n11302), .IN2(n11303), .Q(g33026) );
  AND2X1 U11492 ( .IN1(n8837), .IN2(g3506), .Q(n11303) );
  AND2X1 U11493 ( .IN1(n11304), .IN2(n11289), .Q(n11302) );
  INVX0 U11494 ( .INP(n11305), .ZN(n11304) );
  AND2X1 U11495 ( .IN1(n11306), .IN2(n3492), .Q(n11305) );
  OR2X1 U11496 ( .IN1(n8802), .IN2(n3491), .Q(n11306) );
  OR3X1 U11497 ( .IN1(n11307), .IN2(n11308), .IN3(n11309), .Q(g33024) );
  AND2X1 U11498 ( .IN1(g25648), .IN2(n11310), .Q(n11309) );
  AND3X1 U11499 ( .IN1(n11311), .IN2(n11312), .IN3(n8742), .Q(n11308) );
  OR2X1 U11500 ( .IN1(n11313), .IN2(n11314), .Q(n11311) );
  AND2X1 U11501 ( .IN1(n8837), .IN2(g3171), .Q(n11307) );
  OR2X1 U11502 ( .IN1(n11315), .IN2(n11316), .Q(g33023) );
  AND2X1 U11503 ( .IN1(n11317), .IN2(g3167), .Q(n11316) );
  OR2X1 U11504 ( .IN1(n8802), .IN2(n11318), .Q(n11317) );
  AND2X1 U11505 ( .IN1(n5603), .IN2(n11312), .Q(n11318) );
  AND3X1 U11506 ( .IN1(n8726), .IN2(g3171), .IN3(n11310), .Q(n11315) );
  OR2X1 U11507 ( .IN1(n11319), .IN2(n11320), .Q(g33022) );
  AND2X1 U11508 ( .IN1(n8837), .IN2(g3161), .Q(n11320) );
  AND2X1 U11509 ( .IN1(n11310), .IN2(n11321), .Q(n11319) );
  INVX0 U11510 ( .INP(n106), .ZN(n11321) );
  OR2X1 U11511 ( .IN1(n11322), .IN2(n11323), .Q(g33021) );
  AND2X1 U11512 ( .IN1(n8837), .IN2(g3155), .Q(n11323) );
  AND2X1 U11513 ( .IN1(n11324), .IN2(n11312), .Q(n11322) );
  INVX0 U11514 ( .INP(n11325), .ZN(n11324) );
  AND2X1 U11515 ( .IN1(n11326), .IN2(n3501), .Q(n11325) );
  OR2X1 U11516 ( .IN1(n8802), .IN2(n3502), .Q(n11326) );
  OR3X1 U11517 ( .IN1(n11327), .IN2(n11328), .IN3(n2787), .Q(g33019) );
  AND2X1 U11518 ( .IN1(n11329), .IN2(n8693), .Q(n11328) );
  XOR2X1 U11519 ( .IN1(test_so30), .IN2(n2790), .Q(n11329) );
  AND2X1 U11520 ( .IN1(n8837), .IN2(g2748), .Q(n11327) );
  OR4X1 U11521 ( .IN1(n11330), .IN2(n11331), .IN3(n11332), .IN4(n11333), .Q(
        g33018) );
  AND4X1 U11522 ( .IN1(n3511), .IN2(n11334), .IN3(n11335), .IN4(n8442), .Q(
        n11333) );
  AND2X1 U11523 ( .IN1(n9736), .IN2(g2619), .Q(n11335) );
  AND2X1 U11524 ( .IN1(n8837), .IN2(g2610), .Q(n11332) );
  AND2X1 U11525 ( .IN1(test_so40), .IN2(n11336), .Q(n11331) );
  OR3X1 U11526 ( .IN1(n10902), .IN2(n11337), .IN3(n11338), .Q(n11336) );
  AND2X1 U11527 ( .IN1(n1282), .IN2(n8694), .Q(n11338) );
  INVX0 U11528 ( .INP(n9988), .ZN(n1282) );
  AND3X1 U11529 ( .IN1(n3512), .IN2(n9109), .IN3(n3517), .Q(n11330) );
  AND2X1 U11530 ( .IN1(n9988), .IN2(n3524), .Q(n9109) );
  AND2X1 U11531 ( .IN1(n3505), .IN2(n3525), .Q(n9988) );
  OR3X1 U11532 ( .IN1(n8470), .IN2(n5508), .IN3(g2610), .Q(n3512) );
  OR4X1 U11533 ( .IN1(n11339), .IN2(n11340), .IN3(n3519), .IN4(n11341), .Q(
        g33017) );
  AND2X1 U11534 ( .IN1(n11337), .IN2(g2619), .Q(n11341) );
  AND2X1 U11535 ( .IN1(test_so40), .IN2(n8808), .Q(n11340) );
  AND2X1 U11536 ( .IN1(n3517), .IN2(g2610), .Q(n11339) );
  OR3X1 U11537 ( .IN1(n11342), .IN2(n11343), .IN3(n3519), .Q(g33016) );
  INVX0 U11538 ( .INP(n11344), .ZN(n11343) );
  OR2X1 U11539 ( .IN1(n11337), .IN2(n5372), .Q(n11344) );
  AND2X1 U11540 ( .IN1(n11337), .IN2(g2610), .Q(n11342) );
  OR4X1 U11541 ( .IN1(n11345), .IN2(n11346), .IN3(n3519), .IN4(n11347), .Q(
        g33015) );
  AND3X1 U11542 ( .IN1(n5508), .IN2(n11348), .IN3(n3517), .Q(n11347) );
  AND2X1 U11543 ( .IN1(test_so34), .IN2(n8809), .Q(n11346) );
  AND2X1 U11544 ( .IN1(n11337), .IN2(g2587), .Q(n11345) );
  OR4X1 U11545 ( .IN1(n11349), .IN2(n11350), .IN3(n11351), .IN4(n11352), .Q(
        g33014) );
  AND4X1 U11546 ( .IN1(n3530), .IN2(n11353), .IN3(n11354), .IN4(n8443), .Q(
        n11352) );
  AND2X1 U11547 ( .IN1(n9736), .IN2(g2485), .Q(n11354) );
  AND2X1 U11548 ( .IN1(n8837), .IN2(g2476), .Q(n11351) );
  AND2X1 U11549 ( .IN1(n11355), .IN2(g2491), .Q(n11350) );
  OR3X1 U11550 ( .IN1(n10902), .IN2(n11356), .IN3(n11357), .Q(n11355) );
  AND2X1 U11551 ( .IN1(n1284), .IN2(n8694), .Q(n11357) );
  INVX0 U11552 ( .INP(n9986), .ZN(n1284) );
  AND3X1 U11553 ( .IN1(n3531), .IN2(n9108), .IN3(n3536), .Q(n11349) );
  AND2X1 U11554 ( .IN1(n9986), .IN2(n3524), .Q(n9108) );
  AND3X1 U11555 ( .IN1(g2748), .IN2(n5349), .IN3(n3525), .Q(n9986) );
  OR3X1 U11556 ( .IN1(n8470), .IN2(n5509), .IN3(g2476), .Q(n3531) );
  OR4X1 U11557 ( .IN1(n11358), .IN2(n11359), .IN3(n3538), .IN4(n11360), .Q(
        g33013) );
  AND2X1 U11558 ( .IN1(n11356), .IN2(g2485), .Q(n11360) );
  AND2X1 U11559 ( .IN1(n8837), .IN2(g2491), .Q(n11359) );
  AND2X1 U11560 ( .IN1(n3536), .IN2(g2476), .Q(n11358) );
  OR3X1 U11561 ( .IN1(n11361), .IN2(n11362), .IN3(n3538), .Q(g33012) );
  INVX0 U11562 ( .INP(n11363), .ZN(n11362) );
  OR2X1 U11563 ( .IN1(n11356), .IN2(n5373), .Q(n11363) );
  AND2X1 U11564 ( .IN1(n11356), .IN2(g2476), .Q(n11361) );
  OR4X1 U11565 ( .IN1(n11364), .IN2(n11365), .IN3(n3538), .IN4(n11366), .Q(
        g33011) );
  AND3X1 U11566 ( .IN1(n5509), .IN2(n11367), .IN3(n3536), .Q(n11366) );
  AND2X1 U11567 ( .IN1(n8837), .IN2(g2461), .Q(n11365) );
  AND2X1 U11568 ( .IN1(n11356), .IN2(g2453), .Q(n11364) );
  OR4X1 U11569 ( .IN1(n11368), .IN2(n11369), .IN3(n11370), .IN4(n11371), .Q(
        g33010) );
  AND4X1 U11570 ( .IN1(n3548), .IN2(n11372), .IN3(n11373), .IN4(n8498), .Q(
        n11371) );
  AND2X1 U11571 ( .IN1(n9736), .IN2(g2351), .Q(n11373) );
  AND2X1 U11572 ( .IN1(test_so21), .IN2(n8808), .Q(n11370) );
  AND2X1 U11573 ( .IN1(n11374), .IN2(g2357), .Q(n11369) );
  OR3X1 U11574 ( .IN1(n10902), .IN2(n11375), .IN3(n11376), .Q(n11374) );
  AND2X1 U11575 ( .IN1(n1278), .IN2(n8694), .Q(n11376) );
  INVX0 U11576 ( .INP(n9997), .ZN(n1278) );
  AND3X1 U11577 ( .IN1(n3549), .IN2(n9111), .IN3(n3555), .Q(n11368) );
  AND2X1 U11578 ( .IN1(n9997), .IN2(n3524), .Q(n9111) );
  AND3X1 U11579 ( .IN1(g2741), .IN2(n5516), .IN3(n3525), .Q(n9997) );
  OR3X1 U11580 ( .IN1(test_so21), .IN2(n8470), .IN3(n5511), .Q(n3549) );
  OR4X1 U11581 ( .IN1(n11377), .IN2(n11378), .IN3(n3557), .IN4(n11379), .Q(
        g33009) );
  AND2X1 U11582 ( .IN1(n11375), .IN2(g2351), .Q(n11379) );
  AND2X1 U11583 ( .IN1(n8837), .IN2(g2357), .Q(n11378) );
  AND2X1 U11584 ( .IN1(n3555), .IN2(test_so21), .Q(n11377) );
  OR3X1 U11585 ( .IN1(n11380), .IN2(n11381), .IN3(n3557), .Q(g33008) );
  INVX0 U11586 ( .INP(n11382), .ZN(n11381) );
  OR2X1 U11587 ( .IN1(n11375), .IN2(n5375), .Q(n11382) );
  AND2X1 U11588 ( .IN1(n11375), .IN2(test_so21), .Q(n11380) );
  OR4X1 U11589 ( .IN1(n11383), .IN2(n11384), .IN3(n3557), .IN4(n11385), .Q(
        g33007) );
  AND3X1 U11590 ( .IN1(n5511), .IN2(n11386), .IN3(n3555), .Q(n11385) );
  AND2X1 U11591 ( .IN1(n8838), .IN2(g2327), .Q(n11384) );
  AND2X1 U11592 ( .IN1(n11375), .IN2(g2319), .Q(n11383) );
  OR4X1 U11593 ( .IN1(n11387), .IN2(n11388), .IN3(n11389), .IN4(n11390), .Q(
        g33006) );
  AND4X1 U11594 ( .IN1(n3567), .IN2(n11391), .IN3(n11392), .IN4(n8391), .Q(
        n11390) );
  AND2X1 U11595 ( .IN1(n9736), .IN2(g2217), .Q(n11392) );
  AND2X1 U11596 ( .IN1(n8838), .IN2(g2208), .Q(n11389) );
  AND2X1 U11597 ( .IN1(n11393), .IN2(g2223), .Q(n11388) );
  OR3X1 U11598 ( .IN1(n10902), .IN2(n11394), .IN3(n11395), .Q(n11393) );
  AND2X1 U11599 ( .IN1(n1280), .IN2(n8694), .Q(n11395) );
  INVX0 U11600 ( .INP(n9983), .ZN(n1280) );
  AND3X1 U11601 ( .IN1(n3568), .IN2(n9110), .IN3(n3574), .Q(n11387) );
  AND2X1 U11602 ( .IN1(n9983), .IN2(n3524), .Q(n9110) );
  AND3X1 U11603 ( .IN1(n5349), .IN2(n5516), .IN3(n3525), .Q(n9983) );
  OR3X1 U11604 ( .IN1(n8470), .IN2(n5512), .IN3(g2208), .Q(n3568) );
  OR4X1 U11605 ( .IN1(n11396), .IN2(n11397), .IN3(n3576), .IN4(n11398), .Q(
        g33005) );
  AND2X1 U11606 ( .IN1(n11394), .IN2(g2217), .Q(n11398) );
  AND2X1 U11607 ( .IN1(n8838), .IN2(g2223), .Q(n11397) );
  AND2X1 U11608 ( .IN1(n3574), .IN2(g2208), .Q(n11396) );
  OR3X1 U11609 ( .IN1(n11399), .IN2(n11400), .IN3(n3576), .Q(g33004) );
  INVX0 U11610 ( .INP(n11401), .ZN(n11400) );
  OR2X1 U11611 ( .IN1(n11394), .IN2(n5376), .Q(n11401) );
  AND2X1 U11612 ( .IN1(n11394), .IN2(g2208), .Q(n11399) );
  OR4X1 U11613 ( .IN1(n11402), .IN2(n11403), .IN3(n3576), .IN4(n11404), .Q(
        g33003) );
  AND3X1 U11614 ( .IN1(n5512), .IN2(n11405), .IN3(n3574), .Q(n11404) );
  AND2X1 U11615 ( .IN1(n8838), .IN2(g2193), .Q(n11403) );
  AND2X1 U11616 ( .IN1(n11394), .IN2(g2185), .Q(n11402) );
  OR4X1 U11617 ( .IN1(n11406), .IN2(n11407), .IN3(n11408), .IN4(n11409), .Q(
        g33002) );
  AND4X1 U11618 ( .IN1(n3586), .IN2(n11410), .IN3(n11411), .IN4(n8448), .Q(
        n11409) );
  AND2X1 U11619 ( .IN1(n9736), .IN2(g2060), .Q(n11411) );
  AND2X1 U11620 ( .IN1(n8838), .IN2(g2051), .Q(n11408) );
  AND2X1 U11621 ( .IN1(n11412), .IN2(g2066), .Q(n11407) );
  OR3X1 U11622 ( .IN1(n10902), .IN2(n11413), .IN3(n11414), .Q(n11412) );
  AND2X1 U11623 ( .IN1(n729), .IN2(n8694), .Q(n11414) );
  INVX0 U11624 ( .INP(n9994), .ZN(n729) );
  AND3X1 U11625 ( .IN1(n3587), .IN2(n8988), .IN3(n3593), .Q(n11406) );
  AND2X1 U11626 ( .IN1(n9994), .IN2(n3524), .Q(n8988) );
  AND3X1 U11627 ( .IN1(n5300), .IN2(n756), .IN3(n3505), .Q(n9994) );
  OR3X1 U11628 ( .IN1(n8470), .IN2(n5507), .IN3(g2051), .Q(n3587) );
  OR4X1 U11629 ( .IN1(n11415), .IN2(n11416), .IN3(n3595), .IN4(n11417), .Q(
        g33001) );
  AND2X1 U11630 ( .IN1(n11413), .IN2(g2060), .Q(n11417) );
  AND2X1 U11631 ( .IN1(n8838), .IN2(g2066), .Q(n11416) );
  AND2X1 U11632 ( .IN1(n3593), .IN2(g2051), .Q(n11415) );
  OR3X1 U11633 ( .IN1(n11418), .IN2(n11419), .IN3(n3595), .Q(g33000) );
  INVX0 U11634 ( .INP(n11420), .ZN(n11419) );
  OR2X1 U11635 ( .IN1(n11413), .IN2(n5371), .Q(n11420) );
  AND2X1 U11636 ( .IN1(n11413), .IN2(g2051), .Q(n11418) );
  OR4X1 U11637 ( .IN1(n11421), .IN2(n11422), .IN3(n3595), .IN4(n11423), .Q(
        g32999) );
  AND3X1 U11638 ( .IN1(n5507), .IN2(n11424), .IN3(n3593), .Q(n11423) );
  AND2X1 U11639 ( .IN1(test_so59), .IN2(n8809), .Q(n11422) );
  AND2X1 U11640 ( .IN1(n11413), .IN2(g2028), .Q(n11421) );
  OR4X1 U11641 ( .IN1(n11425), .IN2(n11426), .IN3(n11427), .IN4(n11428), .Q(
        g32998) );
  AND4X1 U11642 ( .IN1(n3604), .IN2(n11429), .IN3(n11430), .IN4(n8449), .Q(
        n11428) );
  AND2X1 U11643 ( .IN1(n9736), .IN2(g1926), .Q(n11430) );
  AND2X1 U11644 ( .IN1(n8838), .IN2(g1917), .Q(n11427) );
  AND2X1 U11645 ( .IN1(n11431), .IN2(g1932), .Q(n11426) );
  OR3X1 U11646 ( .IN1(n10902), .IN2(n11432), .IN3(n11433), .Q(n11431) );
  AND2X1 U11647 ( .IN1(n727), .IN2(n8694), .Q(n11433) );
  AND3X1 U11648 ( .IN1(n3605), .IN2(n8989), .IN3(n3611), .Q(n11425) );
  AND2X1 U11649 ( .IN1(n9992), .IN2(n3524), .Q(n8989) );
  INVX0 U11650 ( .INP(n727), .ZN(n9992) );
  OR4X1 U11651 ( .IN1(n11434), .IN2(g2741), .IN3(test_so30), .IN4(n5516), .Q(
        n727) );
  OR3X1 U11652 ( .IN1(n8470), .IN2(n5510), .IN3(g1917), .Q(n3605) );
  OR4X1 U11653 ( .IN1(n11435), .IN2(n11436), .IN3(n3613), .IN4(n11437), .Q(
        g32997) );
  AND2X1 U11654 ( .IN1(n11432), .IN2(g1926), .Q(n11437) );
  AND2X1 U11655 ( .IN1(n8838), .IN2(g1932), .Q(n11436) );
  AND2X1 U11656 ( .IN1(n3611), .IN2(g1917), .Q(n11435) );
  OR3X1 U11657 ( .IN1(n11438), .IN2(n11439), .IN3(n3613), .Q(g32996) );
  INVX0 U11658 ( .INP(n11440), .ZN(n11439) );
  OR2X1 U11659 ( .IN1(n11432), .IN2(n5374), .Q(n11440) );
  AND2X1 U11660 ( .IN1(n11432), .IN2(g1917), .Q(n11438) );
  OR4X1 U11661 ( .IN1(n11441), .IN2(n11442), .IN3(n3613), .IN4(n11443), .Q(
        g32995) );
  AND3X1 U11662 ( .IN1(n5510), .IN2(n11444), .IN3(n3611), .Q(n11443) );
  AND2X1 U11663 ( .IN1(n8838), .IN2(g1902), .Q(n11442) );
  AND2X1 U11664 ( .IN1(n11432), .IN2(g1894), .Q(n11441) );
  OR4X1 U11665 ( .IN1(n11445), .IN2(n11446), .IN3(n11447), .IN4(n11448), .Q(
        g32994) );
  AND4X1 U11666 ( .IN1(n3622), .IN2(n11449), .IN3(n11450), .IN4(n5596), .Q(
        n11448) );
  AND2X1 U11667 ( .IN1(n9736), .IN2(g1792), .Q(n11450) );
  AND2X1 U11668 ( .IN1(n8838), .IN2(g1783), .Q(n11447) );
  AND2X1 U11669 ( .IN1(n11451), .IN2(g1798), .Q(n11446) );
  OR3X1 U11670 ( .IN1(n10902), .IN2(n11452), .IN3(n11453), .Q(n11451) );
  AND2X1 U11671 ( .IN1(n8711), .IN2(n1635), .Q(n11453) );
  INVX0 U11672 ( .INP(n3005), .ZN(n1635) );
  AND3X1 U11673 ( .IN1(n3623), .IN2(n9106), .IN3(n3628), .Q(n11445) );
  AND2X1 U11674 ( .IN1(n3005), .IN2(n3524), .Q(n9106) );
  OR3X1 U11675 ( .IN1(n8470), .IN2(n5359), .IN3(g1783), .Q(n3623) );
  OR4X1 U11676 ( .IN1(n11454), .IN2(n11455), .IN3(n3630), .IN4(n11456), .Q(
        g32993) );
  AND2X1 U11677 ( .IN1(n11452), .IN2(g1792), .Q(n11456) );
  AND2X1 U11678 ( .IN1(n8838), .IN2(g1798), .Q(n11455) );
  AND2X1 U11679 ( .IN1(n3628), .IN2(g1783), .Q(n11454) );
  OR3X1 U11680 ( .IN1(n11457), .IN2(n11458), .IN3(n3630), .Q(g32992) );
  INVX0 U11681 ( .INP(n11459), .ZN(n11458) );
  OR2X1 U11682 ( .IN1(n11452), .IN2(n5602), .Q(n11459) );
  AND2X1 U11683 ( .IN1(n11452), .IN2(g1783), .Q(n11457) );
  OR4X1 U11684 ( .IN1(n11460), .IN2(n11461), .IN3(n3630), .IN4(n11462), .Q(
        g32991) );
  AND3X1 U11685 ( .IN1(n5359), .IN2(n11463), .IN3(n3628), .Q(n11462) );
  AND2X1 U11686 ( .IN1(n8838), .IN2(g1768), .Q(n11461) );
  AND2X1 U11687 ( .IN1(n11452), .IN2(g1760), .Q(n11460) );
  OR4X1 U11688 ( .IN1(n11464), .IN2(n11465), .IN3(n11466), .IN4(n11467), .Q(
        g32990) );
  AND4X1 U11689 ( .IN1(n3640), .IN2(n11468), .IN3(n11469), .IN4(n8499), .Q(
        n11467) );
  AND2X1 U11690 ( .IN1(n9736), .IN2(g1657), .Q(n11469) );
  AND2X1 U11691 ( .IN1(test_so94), .IN2(n8808), .Q(n11466) );
  AND2X1 U11692 ( .IN1(n11470), .IN2(g1664), .Q(n11465) );
  OR3X1 U11693 ( .IN1(n11471), .IN2(n10902), .IN3(n11472), .Q(n11470) );
  AND2X1 U11694 ( .IN1(n724), .IN2(n8694), .Q(n11472) );
  INVX0 U11695 ( .INP(n9995), .ZN(n724) );
  INVX0 U11696 ( .INP(n10737), .ZN(n10902) );
  OR2X1 U11697 ( .IN1(n2760), .IN2(n8794), .Q(n10737) );
  AND3X1 U11698 ( .IN1(n3641), .IN2(n8990), .IN3(n3646), .Q(n11464) );
  AND2X1 U11699 ( .IN1(n9995), .IN2(n3524), .Q(n8990) );
  AND2X1 U11700 ( .IN1(n756), .IN2(n3653), .Q(n9995) );
  INVX0 U11701 ( .INP(n11434), .ZN(n756) );
  OR2X1 U11702 ( .IN1(n11473), .IN2(n11474), .Q(n11434) );
  XOR2X1 U11703 ( .IN1(g2759), .IN2(g72), .Q(n11474) );
  XOR2X1 U11704 ( .IN1(g2763), .IN2(g73), .Q(n11473) );
  OR3X1 U11705 ( .IN1(test_so94), .IN2(n8470), .IN3(n5525), .Q(n3641) );
  OR4X1 U11706 ( .IN1(n11475), .IN2(n11476), .IN3(n3648), .IN4(n11477), .Q(
        g32989) );
  AND2X1 U11707 ( .IN1(n11471), .IN2(g1657), .Q(n11477) );
  AND2X1 U11708 ( .IN1(n8838), .IN2(g1664), .Q(n11476) );
  AND2X1 U11709 ( .IN1(n3646), .IN2(test_so94), .Q(n11475) );
  OR3X1 U11710 ( .IN1(n11478), .IN2(n11479), .IN3(n3648), .Q(g32988) );
  INVX0 U11711 ( .INP(n11480), .ZN(n11479) );
  OR2X1 U11712 ( .IN1(n11471), .IN2(n5370), .Q(n11480) );
  AND2X1 U11713 ( .IN1(n11471), .IN2(test_so94), .Q(n11478) );
  OR4X1 U11714 ( .IN1(n11481), .IN2(n11482), .IN3(n3648), .IN4(n11483), .Q(
        g32987) );
  AND3X1 U11715 ( .IN1(n5525), .IN2(n11484), .IN3(n3646), .Q(n11483) );
  AND2X1 U11716 ( .IN1(n8838), .IN2(g1632), .Q(n11482) );
  AND2X1 U11717 ( .IN1(n11471), .IN2(g1624), .Q(n11481) );
  OR3X1 U11718 ( .IN1(n11485), .IN2(n11486), .IN3(n11487), .Q(g32986) );
  AND3X1 U11719 ( .IN1(n11067), .IN2(n8328), .IN3(n11488), .Q(n11487) );
  INVX0 U11720 ( .INP(n11071), .ZN(n11067) );
  AND2X1 U11721 ( .IN1(n8838), .IN2(g1367), .Q(n11486) );
  AND3X1 U11722 ( .IN1(n11071), .IN2(g1373), .IN3(n8741), .Q(n11485) );
  OR2X1 U11723 ( .IN1(n11489), .IN2(n9104), .Q(n11071) );
  AND2X1 U11724 ( .IN1(n8468), .IN2(n11068), .Q(n11489) );
  AND2X1 U11725 ( .IN1(n11490), .IN2(g1274), .Q(g32985) );
  OR2X1 U11726 ( .IN1(n8801), .IN2(n11491), .Q(n11490) );
  AND2X1 U11727 ( .IN1(n11075), .IN2(n9448), .Q(n11491) );
  INVX0 U11728 ( .INP(n11077), .ZN(n11075) );
  OR2X1 U11729 ( .IN1(n5716), .IN2(n11492), .Q(n11077) );
  OR3X1 U11730 ( .IN1(n11493), .IN2(n11494), .IN3(n11495), .Q(g32984) );
  AND2X1 U11731 ( .IN1(n8838), .IN2(g1263), .Q(n11495) );
  AND2X1 U11732 ( .IN1(n5716), .IN2(n3662), .Q(n11494) );
  AND3X1 U11733 ( .IN1(n11076), .IN2(n11492), .IN3(g1270), .Q(n11493) );
  INVX0 U11734 ( .INP(n3662), .ZN(n11492) );
  OR3X1 U11735 ( .IN1(n11496), .IN2(n11497), .IN3(n11498), .Q(g32983) );
  AND3X1 U11736 ( .IN1(n11082), .IN2(n8327), .IN3(n11499), .Q(n11498) );
  INVX0 U11737 ( .INP(n11086), .ZN(n11082) );
  AND2X1 U11738 ( .IN1(n8838), .IN2(g1024), .Q(n11497) );
  AND3X1 U11739 ( .IN1(n11086), .IN2(g1030), .IN3(n8741), .Q(n11496) );
  OR2X1 U11740 ( .IN1(n11500), .IN2(n9007), .Q(n11086) );
  AND2X1 U11741 ( .IN1(n8465), .IN2(n11083), .Q(n11500) );
  AND2X1 U11742 ( .IN1(n11501), .IN2(g930), .Q(g32982) );
  OR2X1 U11743 ( .IN1(n8801), .IN2(n11502), .Q(n11501) );
  AND2X1 U11744 ( .IN1(n11090), .IN2(n9449), .Q(n11502) );
  INVX0 U11745 ( .INP(n11092), .ZN(n11090) );
  OR2X1 U11746 ( .IN1(n5725), .IN2(n11503), .Q(n11092) );
  OR3X1 U11747 ( .IN1(n11504), .IN2(n11505), .IN3(n11506), .Q(g32981) );
  AND2X1 U11748 ( .IN1(n8838), .IN2(g918), .Q(n11506) );
  AND2X1 U11749 ( .IN1(n5725), .IN2(n3671), .Q(n11505) );
  AND3X1 U11750 ( .IN1(n11091), .IN2(n11503), .IN3(g925), .Q(n11504) );
  INVX0 U11751 ( .INP(n3671), .ZN(n11503) );
  AND3X1 U11752 ( .IN1(n11507), .IN2(n11508), .IN3(n8741), .Q(g32980) );
  OR2X1 U11753 ( .IN1(n11509), .IN2(g854), .Q(n11508) );
  INVX0 U11754 ( .INP(n11510), .ZN(n11507) );
  AND2X1 U11755 ( .IN1(n11509), .IN2(n2644), .Q(n11510) );
  INVX0 U11756 ( .INP(n9796), .ZN(n11509) );
  OR4X1 U11757 ( .IN1(n5633), .IN2(g385), .IN3(n8361), .IN4(n8307), .Q(n9796)
         );
  OR3X1 U11758 ( .IN1(n11511), .IN2(n11512), .IN3(n11513), .Q(g32979) );
  AND2X1 U11759 ( .IN1(test_so2), .IN2(n8808), .Q(n11513) );
  AND2X1 U11760 ( .IN1(n3272), .IN2(n5331), .Q(n11512) );
  AND3X1 U11761 ( .IN1(n2404), .IN2(n11514), .IN3(g758), .Q(n11511) );
  INVX0 U11762 ( .INP(n3272), .ZN(n11514) );
  OR3X1 U11763 ( .IN1(n11515), .IN2(n11516), .IN3(n11517), .Q(g32978) );
  AND2X1 U11764 ( .IN1(n8838), .IN2(g582), .Q(n11517) );
  AND2X1 U11765 ( .IN1(n3274), .IN2(n5472), .Q(n11516) );
  AND3X1 U11766 ( .IN1(n2421), .IN2(n11518), .IN3(g590), .Q(n11515) );
  INVX0 U11767 ( .INP(n3274), .ZN(n11518) );
  OR3X1 U11768 ( .IN1(n11519), .IN2(n11520), .IN3(n11521), .Q(g32977) );
  AND2X1 U11769 ( .IN1(test_so51), .IN2(n8809), .Q(n11521) );
  AND2X1 U11770 ( .IN1(n3279), .IN2(n5679), .Q(n11520) );
  AND3X1 U11771 ( .IN1(n8473), .IN2(n11522), .IN3(g291), .Q(n11519) );
  INVX0 U11772 ( .INP(n3279), .ZN(n11522) );
  AND3X1 U11773 ( .IN1(n11523), .IN2(test_so51), .IN3(test_so55), .Q(n3279) );
  OR3X1 U11774 ( .IN1(n11524), .IN2(n11525), .IN3(n11526), .Q(g32976) );
  AND2X1 U11775 ( .IN1(n8838), .IN2(g164), .Q(n11526) );
  AND2X1 U11776 ( .IN1(n3281), .IN2(n5676), .Q(n11525) );
  AND3X1 U11777 ( .IN1(n9969), .IN2(n11527), .IN3(g150), .Q(n11524) );
  INVX0 U11778 ( .INP(n3281), .ZN(n11527) );
  AND4X1 U11779 ( .IN1(n11528), .IN2(n11529), .IN3(n11530), .IN4(n11531), .Q(
        g32185) );
  AND4X1 U11780 ( .IN1(n11532), .IN2(n11533), .IN3(n11534), .IN4(n11535), .Q(
        n11531) );
  OR2X1 U11781 ( .IN1(n8039), .IN2(n8519), .Q(n11535) );
  OR2X1 U11782 ( .IN1(n5750), .IN2(n8192), .Q(n11534) );
  OR2X1 U11783 ( .IN1(n8037), .IN2(n8193), .Q(n11533) );
  OR2X1 U11784 ( .IN1(n8036), .IN2(n8194), .Q(n11532) );
  OR2X1 U11785 ( .IN1(n8038), .IN2(n8520), .Q(n11530) );
  OR2X1 U11786 ( .IN1(n8196), .IN2(n8197), .Q(n11529) );
  OR2X1 U11787 ( .IN1(n8040), .IN2(n8195), .Q(n11528) );
  OR4X1 U11788 ( .IN1(n11536), .IN2(n11537), .IN3(n11538), .IN4(n11539), .Q(
        g31904) );
  AND2X1 U11789 ( .IN1(n8409), .IN2(n11540), .Q(n11539) );
  INVX0 U11790 ( .INP(n11541), .ZN(n11538) );
  OR4X1 U11791 ( .IN1(n11542), .IN2(n11540), .IN3(n11543), .IN4(n8409), .Q(
        n11541) );
  AND2X1 U11792 ( .IN1(n11544), .IN2(n8695), .Q(n11537) );
  AND2X1 U11793 ( .IN1(n8838), .IN2(g5029), .Q(n11536) );
  OR4X1 U11794 ( .IN1(n11236), .IN2(n11545), .IN3(n11546), .IN4(n11547), .Q(
        g31903) );
  AND2X1 U11795 ( .IN1(n11237), .IN2(n5607), .Q(n11547) );
  INVX0 U11796 ( .INP(n11548), .ZN(n11546) );
  OR4X1 U11797 ( .IN1(n11237), .IN2(n11549), .IN3(n11543), .IN4(n5607), .Q(
        n11548) );
  AND2X1 U11798 ( .IN1(g5046), .IN2(n11550), .Q(n11237) );
  AND2X1 U11799 ( .IN1(n8839), .IN2(g5046), .Q(n11545) );
  AND3X1 U11800 ( .IN1(n8727), .IN2(n5607), .IN3(n11549), .Q(n11236) );
  OR3X1 U11801 ( .IN1(n11551), .IN2(n11552), .IN3(n11553), .Q(g31902) );
  AND2X1 U11802 ( .IN1(n11542), .IN2(n8695), .Q(n11553) );
  AND2X1 U11803 ( .IN1(n11554), .IN2(g5016), .Q(n11552) );
  OR2X1 U11804 ( .IN1(n8801), .IN2(n11555), .Q(n11554) );
  AND2X1 U11805 ( .IN1(n5601), .IN2(g5062), .Q(n11555) );
  AND4X1 U11806 ( .IN1(n11232), .IN2(g5029), .IN3(n11556), .IN4(n11557), .Q(
        n11551) );
  OR2X1 U11807 ( .IN1(n8437), .IN2(g5016), .Q(n11557) );
  OR2X1 U11808 ( .IN1(n8438), .IN2(n5369), .Q(n11556) );
  OR4X1 U11809 ( .IN1(n11558), .IN2(n11559), .IN3(n11560), .IN4(n11561), .Q(
        g31901) );
  AND2X1 U11810 ( .IN1(n11550), .IN2(n5578), .Q(n11561) );
  INVX0 U11811 ( .INP(n11562), .ZN(n11560) );
  OR4X1 U11812 ( .IN1(n11563), .IN2(n11550), .IN3(n11543), .IN4(n5578), .Q(
        n11562) );
  INVX0 U11813 ( .INP(n11232), .ZN(n11543) );
  AND3X1 U11814 ( .IN1(g5037), .IN2(g5041), .IN3(n11564), .Q(n11550) );
  AND2X1 U11815 ( .IN1(n11549), .IN2(n8695), .Q(n11559) );
  AND2X1 U11816 ( .IN1(n5578), .IN2(n11563), .Q(n11549) );
  AND3X1 U11817 ( .IN1(n5605), .IN2(n11544), .IN3(n5611), .Q(n11563) );
  AND2X1 U11818 ( .IN1(n8839), .IN2(g5041), .Q(n11558) );
  OR3X1 U11819 ( .IN1(n11565), .IN2(n11566), .IN3(n11567), .Q(g31900) );
  AND2X1 U11820 ( .IN1(n11568), .IN2(n5605), .Q(n11567) );
  AND2X1 U11821 ( .IN1(n11569), .IN2(g5037), .Q(n11566) );
  OR3X1 U11822 ( .IN1(n11570), .IN2(n11571), .IN3(n8792), .Q(n11569) );
  AND2X1 U11823 ( .IN1(n11564), .IN2(n5605), .Q(n11571) );
  AND3X1 U11824 ( .IN1(n11232), .IN2(n11572), .IN3(g5041), .Q(n11570) );
  AND4X1 U11825 ( .IN1(n11573), .IN2(g5041), .IN3(n11232), .IN4(n5611), .Q(
        n11565) );
  OR4X1 U11826 ( .IN1(n11568), .IN2(n11574), .IN3(n11575), .IN4(n11576), .Q(
        g31899) );
  AND2X1 U11827 ( .IN1(n5611), .IN2(n11564), .Q(n11576) );
  AND4X1 U11828 ( .IN1(n11572), .IN2(n11573), .IN3(n11232), .IN4(g5037), .Q(
        n11575) );
  INVX0 U11829 ( .INP(n11544), .ZN(n11573) );
  INVX0 U11830 ( .INP(n11564), .ZN(n11572) );
  AND2X1 U11831 ( .IN1(g5033), .IN2(n11540), .Q(n11564) );
  AND3X1 U11832 ( .IN1(g5062), .IN2(g5029), .IN3(g5016), .Q(n11540) );
  AND2X1 U11833 ( .IN1(n8839), .IN2(g5033), .Q(n11574) );
  AND3X1 U11834 ( .IN1(n8727), .IN2(n11544), .IN3(n5611), .Q(n11568) );
  AND2X1 U11835 ( .IN1(n11542), .IN2(n8409), .Q(n11544) );
  AND3X1 U11836 ( .IN1(g5022), .IN2(n5369), .IN3(n5601), .Q(n11542) );
  OR3X1 U11837 ( .IN1(n11577), .IN2(n11578), .IN3(n11579), .Q(g31898) );
  AND3X1 U11838 ( .IN1(n11232), .IN2(n11580), .IN3(n5369), .Q(n11579) );
  AND4X1 U11839 ( .IN1(n11581), .IN2(n11582), .IN3(n11583), .IN4(n11584), .Q(
        n11232) );
  AND2X1 U11840 ( .IN1(n8711), .IN2(n11585), .Q(n11584) );
  AND2X1 U11841 ( .IN1(n8839), .IN2(g5022), .Q(n11578) );
  AND3X1 U11842 ( .IN1(n11586), .IN2(g5016), .IN3(n8730), .Q(n11577) );
  INVX0 U11843 ( .INP(n11580), .ZN(n11586) );
  OR2X1 U11844 ( .IN1(g5022), .IN2(g5062), .Q(n11580) );
  OR3X1 U11845 ( .IN1(n11245), .IN2(n11587), .IN3(n11588), .Q(g31897) );
  AND2X1 U11846 ( .IN1(n8839), .IN2(g4423), .Q(n11587) );
  AND2X1 U11847 ( .IN1(g4575), .IN2(n11252), .Q(n11245) );
  OR3X1 U11848 ( .IN1(n11253), .IN2(n11589), .IN3(n11588), .Q(g31896) );
  OR2X1 U11849 ( .IN1(n11590), .IN2(n11591), .Q(n11588) );
  AND2X1 U11850 ( .IN1(n11252), .IN2(n11592), .Q(n11591) );
  OR2X1 U11851 ( .IN1(n10721), .IN2(n11257), .Q(n11592) );
  INVX0 U11852 ( .INP(g72), .ZN(n11257) );
  INVX0 U11853 ( .INP(g73), .ZN(n10721) );
  AND3X1 U11854 ( .IN1(n8727), .IN2(g4372), .IN3(n5670), .Q(n11590) );
  INVX0 U11855 ( .INP(n11593), .ZN(n11589) );
  OR2X1 U11856 ( .IN1(n8677), .IN2(n5849), .Q(n11593) );
  AND2X1 U11857 ( .IN1(n11252), .IN2(test_so100), .Q(n11253) );
  INVX0 U11858 ( .INP(n11241), .ZN(n11252) );
  OR2X1 U11859 ( .IN1(n5670), .IN2(n8794), .Q(n11241) );
  OR2X1 U11860 ( .IN1(n11594), .IN2(n9736), .Q(g31895) );
  INVX0 U11861 ( .INP(n9752), .ZN(n9736) );
  OR2X1 U11862 ( .IN1(n8802), .IN2(n1697), .Q(n9752) );
  INVX0 U11863 ( .INP(n2760), .ZN(n1697) );
  AND2X1 U11864 ( .IN1(n8839), .IN2(g4382), .Q(n11594) );
  OR3X1 U11865 ( .IN1(n11595), .IN2(n11596), .IN3(n8481), .Q(g31894) );
  AND2X1 U11866 ( .IN1(n11597), .IN2(n8695), .Q(n11596) );
  XOR2X1 U11867 ( .IN1(n11264), .IN2(n5350), .Q(n11597) );
  OR2X1 U11868 ( .IN1(n5340), .IN2(n3729), .Q(n11264) );
  OR2X1 U11869 ( .IN1(n5480), .IN2(n11598), .Q(n3729) );
  AND2X1 U11870 ( .IN1(n8839), .IN2(g4093), .Q(n11595) );
  OR2X1 U11871 ( .IN1(n11599), .IN2(n11600), .Q(g31872) );
  AND2X1 U11872 ( .IN1(n8839), .IN2(g2741), .Q(n11600) );
  AND2X1 U11873 ( .IN1(n11601), .IN2(n3730), .Q(n11599) );
  XOR2X1 U11874 ( .IN1(n11602), .IN2(n5516), .Q(n11601) );
  OR2X1 U11875 ( .IN1(n5349), .IN2(n3506), .Q(n11602) );
  OR3X1 U11876 ( .IN1(n11603), .IN2(n11604), .IN3(n11605), .Q(g31871) );
  AND2X1 U11877 ( .IN1(n3733), .IN2(n11488), .Q(n11605) );
  AND3X1 U11878 ( .IN1(n9104), .IN2(g1367), .IN3(n8746), .Q(n11604) );
  OR2X1 U11879 ( .IN1(n11606), .IN2(n9103), .Q(n9104) );
  AND2X1 U11880 ( .IN1(n8325), .IN2(n11068), .Q(n11606) );
  AND2X1 U11881 ( .IN1(n8839), .IN2(g1361), .Q(n11603) );
  OR3X1 U11882 ( .IN1(n11607), .IN2(n11608), .IN3(n11609), .Q(g31870) );
  AND2X1 U11883 ( .IN1(n8839), .IN2(g1259), .Q(n11609) );
  AND2X1 U11884 ( .IN1(n3664), .IN2(n5674), .Q(n11608) );
  AND3X1 U11885 ( .IN1(n11076), .IN2(n11610), .IN3(g1263), .Q(n11607) );
  INVX0 U11886 ( .INP(n3664), .ZN(n11610) );
  OR3X1 U11887 ( .IN1(n11611), .IN2(n11612), .IN3(n11613), .Q(g31869) );
  AND2X1 U11888 ( .IN1(n3738), .IN2(n11499), .Q(n11613) );
  AND3X1 U11889 ( .IN1(n9007), .IN2(g1024), .IN3(n8741), .Q(n11612) );
  OR2X1 U11890 ( .IN1(n11614), .IN2(n9006), .Q(n9007) );
  AND2X1 U11891 ( .IN1(n8324), .IN2(n11083), .Q(n11614) );
  AND2X1 U11892 ( .IN1(n8839), .IN2(g1018), .Q(n11611) );
  OR3X1 U11893 ( .IN1(n11615), .IN2(n11616), .IN3(n11617), .Q(g31868) );
  AND2X1 U11894 ( .IN1(n8839), .IN2(g914), .Q(n11617) );
  AND2X1 U11895 ( .IN1(n3673), .IN2(n5673), .Q(n11616) );
  AND3X1 U11896 ( .IN1(n11091), .IN2(n11618), .IN3(g918), .Q(n11615) );
  INVX0 U11897 ( .INP(n3673), .ZN(n11618) );
  OR3X1 U11898 ( .IN1(n11619), .IN2(n11620), .IN3(n11621), .Q(g31867) );
  AND2X1 U11899 ( .IN1(n8839), .IN2(g744), .Q(n11621) );
  AND2X1 U11900 ( .IN1(n3682), .IN2(n5471), .Q(n11620) );
  AND3X1 U11901 ( .IN1(n2404), .IN2(test_so2), .IN3(n11622), .Q(n11619) );
  INVX0 U11902 ( .INP(n3682), .ZN(n11622) );
  OR3X1 U11903 ( .IN1(n11623), .IN2(n11624), .IN3(n11625), .Q(g31866) );
  AND2X1 U11904 ( .IN1(n8839), .IN2(g577), .Q(n11625) );
  AND2X1 U11905 ( .IN1(n3684), .IN2(n5552), .Q(n11624) );
  AND3X1 U11906 ( .IN1(n2421), .IN2(n11626), .IN3(g582), .Q(n11623) );
  INVX0 U11907 ( .INP(n3684), .ZN(n11626) );
  OR2X1 U11908 ( .IN1(n11627), .IN2(n11628), .Q(g31865) );
  AND3X1 U11909 ( .IN1(n8473), .IN2(test_so51), .IN3(n8515), .Q(n11628) );
  AND2X1 U11910 ( .IN1(test_so55), .IN2(n11629), .Q(n11627) );
  OR2X1 U11911 ( .IN1(n8802), .IN2(n11630), .Q(n11629) );
  AND2X1 U11912 ( .IN1(n11523), .IN2(n8524), .Q(n11630) );
  OR3X1 U11913 ( .IN1(n11631), .IN2(n11632), .IN3(n11633), .Q(g31864) );
  AND2X1 U11914 ( .IN1(test_so73), .IN2(n8808), .Q(n11633) );
  AND2X1 U11915 ( .IN1(n3687), .IN2(n5561), .Q(n11632) );
  AND3X1 U11916 ( .IN1(n9969), .IN2(n11634), .IN3(g164), .Q(n11631) );
  INVX0 U11917 ( .INP(n3687), .ZN(n11634) );
  AND3X1 U11918 ( .IN1(n11635), .IN2(n11636), .IN3(test_so73), .Q(n3687) );
  AND2X1 U11919 ( .IN1(g1668), .IN2(n5549), .Q(g31862) );
  OR2X1 U11920 ( .IN1(n11637), .IN2(n11638), .Q(g31793) );
  AND3X1 U11921 ( .IN1(n11639), .IN2(n9482), .IN3(n9484), .Q(n11638) );
  OR2X1 U11922 ( .IN1(n11640), .IN2(n11641), .Q(n11639) );
  AND2X1 U11923 ( .IN1(n11642), .IN2(n11643), .Q(n11641) );
  AND3X1 U11924 ( .IN1(n8318), .IN2(n11644), .IN3(n8319), .Q(n11640) );
  OR2X1 U11925 ( .IN1(n11645), .IN2(n11642), .Q(n11644) );
  AND2X1 U11926 ( .IN1(n11646), .IN2(n11643), .Q(n11645) );
  OR2X1 U11927 ( .IN1(n11647), .IN2(n11648), .Q(n11646) );
  AND3X1 U11928 ( .IN1(n11649), .IN2(n11650), .IN3(n11651), .Q(n11647) );
  OR2X1 U11929 ( .IN1(n11652), .IN2(n11653), .Q(n11651) );
  AND2X1 U11930 ( .IN1(n11654), .IN2(n11655), .Q(n11652) );
  OR2X1 U11931 ( .IN1(n11654), .IN2(n11655), .Q(n11649) );
  AND2X1 U11932 ( .IN1(n9483), .IN2(n11656), .Q(n11637) );
  OR2X1 U11933 ( .IN1(n11657), .IN2(n9484), .Q(n11656) );
  AND2X1 U11934 ( .IN1(n11658), .IN2(n11659), .Q(n9484) );
  AND2X1 U11935 ( .IN1(n11660), .IN2(n9482), .Q(n11657) );
  OR2X1 U11936 ( .IN1(n11659), .IN2(n11658), .Q(n11660) );
  AND4X1 U11937 ( .IN1(n8318), .IN2(n8319), .IN3(n11643), .IN4(n11642), .Q(
        n9483) );
  AND2X1 U11938 ( .IN1(n11650), .IN2(n11648), .Q(n11642) );
  AND3X1 U11939 ( .IN1(n11653), .IN2(n11655), .IN3(n11654), .Q(n11648) );
  OR2X1 U11940 ( .IN1(n8351), .IN2(n10582), .Q(g31665) );
  OR2X1 U11941 ( .IN1(n5488), .IN2(n10582), .Q(g31656) );
  INVX0 U11942 ( .INP(g113), .ZN(n10582) );
  OR3X1 U11943 ( .IN1(n11661), .IN2(n11662), .IN3(n11663), .Q(g30563) );
  AND2X1 U11944 ( .IN1(n8839), .IN2(g6653), .Q(n11663) );
  AND2X1 U11945 ( .IN1(n3765), .IN2(n10569), .Q(n11662) );
  AND2X1 U11946 ( .IN1(n11664), .IN2(g6657), .Q(n11661) );
  OR3X1 U11947 ( .IN1(n11665), .IN2(n11666), .IN3(n11667), .Q(g30562) );
  AND2X1 U11948 ( .IN1(n11668), .IN2(n3765), .Q(n11667) );
  INVX0 U11949 ( .INP(n11669), .ZN(n11668) );
  AND2X1 U11950 ( .IN1(n8839), .IN2(g6649), .Q(n11666) );
  AND3X1 U11951 ( .IN1(n11669), .IN2(g6605), .IN3(n8741), .Q(n11665) );
  OR2X1 U11952 ( .IN1(n5646), .IN2(n1331), .Q(n11669) );
  OR3X1 U11953 ( .IN1(n11670), .IN2(n11671), .IN3(n11672), .Q(g30561) );
  AND2X1 U11954 ( .IN1(n11128), .IN2(n3765), .Q(n11672) );
  INVX0 U11955 ( .INP(n11673), .ZN(n11128) );
  AND2X1 U11956 ( .IN1(n8839), .IN2(g6645), .Q(n11671) );
  AND3X1 U11957 ( .IN1(n11673), .IN2(g6597), .IN3(n8741), .Q(n11670) );
  OR2X1 U11958 ( .IN1(n5646), .IN2(n1324), .Q(n11673) );
  OR3X1 U11959 ( .IN1(n11674), .IN2(n11675), .IN3(n11676), .Q(g30560) );
  AND2X1 U11960 ( .IN1(n11677), .IN2(n3765), .Q(n11676) );
  INVX0 U11961 ( .INP(n11678), .ZN(n11677) );
  AND2X1 U11962 ( .IN1(n8839), .IN2(g6641), .Q(n11675) );
  AND3X1 U11963 ( .IN1(n11678), .IN2(g6589), .IN3(n8741), .Q(n11674) );
  OR2X1 U11964 ( .IN1(n5646), .IN2(n1326), .Q(n11678) );
  OR3X1 U11965 ( .IN1(n11679), .IN2(n11680), .IN3(n11681), .Q(g30559) );
  AND2X1 U11966 ( .IN1(n3774), .IN2(n11682), .Q(n11681) );
  AND3X1 U11967 ( .IN1(n11683), .IN2(g6653), .IN3(n8741), .Q(n11680) );
  OR2X1 U11968 ( .IN1(n704), .IN2(n1330), .Q(n11683) );
  AND2X1 U11969 ( .IN1(n8839), .IN2(g6637), .Q(n11679) );
  OR3X1 U11970 ( .IN1(n11684), .IN2(n11685), .IN3(n11686), .Q(g30558) );
  AND2X1 U11971 ( .IN1(n3774), .IN2(n11131), .Q(n11686) );
  AND3X1 U11972 ( .IN1(n11687), .IN2(g6649), .IN3(n8741), .Q(n11685) );
  OR2X1 U11973 ( .IN1(n704), .IN2(n1331), .Q(n11687) );
  AND2X1 U11974 ( .IN1(n8839), .IN2(g6633), .Q(n11684) );
  OR3X1 U11975 ( .IN1(n11688), .IN2(n11689), .IN3(n11690), .Q(g30557) );
  AND2X1 U11976 ( .IN1(n3774), .IN2(n11691), .Q(n11690) );
  AND3X1 U11977 ( .IN1(n11692), .IN2(g6645), .IN3(n8742), .Q(n11689) );
  OR2X1 U11978 ( .IN1(n704), .IN2(n1324), .Q(n11692) );
  AND2X1 U11979 ( .IN1(n8839), .IN2(g6629), .Q(n11688) );
  OR3X1 U11980 ( .IN1(n11693), .IN2(n11694), .IN3(n11695), .Q(g30556) );
  AND2X1 U11981 ( .IN1(n3774), .IN2(n11696), .Q(n11695) );
  AND3X1 U11982 ( .IN1(n11697), .IN2(g6641), .IN3(n8742), .Q(n11694) );
  OR2X1 U11983 ( .IN1(n704), .IN2(n1326), .Q(n11697) );
  OR2X1 U11984 ( .IN1(n8314), .IN2(n5571), .Q(n704) );
  AND2X1 U11985 ( .IN1(n8839), .IN2(g6625), .Q(n11693) );
  OR3X1 U11986 ( .IN1(n11698), .IN2(n11699), .IN3(n11700), .Q(g30555) );
  AND2X1 U11987 ( .IN1(n3780), .IN2(n11682), .Q(n11700) );
  AND3X1 U11988 ( .IN1(n11701), .IN2(g6637), .IN3(n8742), .Q(n11699) );
  OR2X1 U11989 ( .IN1(n3406), .IN2(n1330), .Q(n11701) );
  AND2X1 U11990 ( .IN1(n8840), .IN2(g6621), .Q(n11698) );
  OR3X1 U11991 ( .IN1(n11702), .IN2(n11703), .IN3(n11704), .Q(g30554) );
  AND2X1 U11992 ( .IN1(n3780), .IN2(n11131), .Q(n11704) );
  AND3X1 U11993 ( .IN1(n11705), .IN2(g6633), .IN3(n8742), .Q(n11703) );
  OR2X1 U11994 ( .IN1(n3406), .IN2(n1331), .Q(n11705) );
  AND2X1 U11995 ( .IN1(n8840), .IN2(g6617), .Q(n11702) );
  OR3X1 U11996 ( .IN1(n11706), .IN2(n11707), .IN3(n11708), .Q(g30553) );
  AND2X1 U11997 ( .IN1(n3780), .IN2(n11691), .Q(n11708) );
  AND3X1 U11998 ( .IN1(n11709), .IN2(g6629), .IN3(n8742), .Q(n11707) );
  OR2X1 U11999 ( .IN1(n3406), .IN2(n1324), .Q(n11709) );
  AND2X1 U12000 ( .IN1(n8840), .IN2(g6613), .Q(n11706) );
  OR3X1 U12001 ( .IN1(n11710), .IN2(n11711), .IN3(n11712), .Q(g30552) );
  AND2X1 U12002 ( .IN1(n3780), .IN2(n11696), .Q(n11712) );
  AND3X1 U12003 ( .IN1(n11713), .IN2(g6625), .IN3(n8742), .Q(n11711) );
  OR2X1 U12004 ( .IN1(n3406), .IN2(n1326), .Q(n11713) );
  OR2X1 U12005 ( .IN1(n8314), .IN2(g6549), .Q(n3406) );
  AND2X1 U12006 ( .IN1(n8840), .IN2(g6609), .Q(n11710) );
  OR3X1 U12007 ( .IN1(n11714), .IN2(n11715), .IN3(n11716), .Q(g30551) );
  AND2X1 U12008 ( .IN1(n3785), .IN2(n11682), .Q(n11716) );
  AND3X1 U12009 ( .IN1(n11717), .IN2(g6621), .IN3(n8742), .Q(n11715) );
  OR2X1 U12010 ( .IN1(n3407), .IN2(n1330), .Q(n11717) );
  AND2X1 U12011 ( .IN1(n8840), .IN2(g6601), .Q(n11714) );
  OR3X1 U12012 ( .IN1(n11718), .IN2(n11719), .IN3(n11720), .Q(g30550) );
  AND2X1 U12013 ( .IN1(n3785), .IN2(n11131), .Q(n11720) );
  INVX0 U12014 ( .INP(n1331), .ZN(n11131) );
  AND3X1 U12015 ( .IN1(n11721), .IN2(g6617), .IN3(n8742), .Q(n11719) );
  OR2X1 U12016 ( .IN1(n3407), .IN2(n1331), .Q(n11721) );
  OR2X1 U12017 ( .IN1(n5563), .IN2(g6565), .Q(n1331) );
  AND2X1 U12018 ( .IN1(n8840), .IN2(g6593), .Q(n11718) );
  OR3X1 U12019 ( .IN1(n11722), .IN2(n11723), .IN3(n11724), .Q(g30549) );
  AND2X1 U12020 ( .IN1(n3785), .IN2(n11691), .Q(n11724) );
  INVX0 U12021 ( .INP(n1324), .ZN(n11691) );
  AND3X1 U12022 ( .IN1(n11725), .IN2(g6613), .IN3(n8742), .Q(n11723) );
  OR2X1 U12023 ( .IN1(n3407), .IN2(n1324), .Q(n11725) );
  OR2X1 U12024 ( .IN1(n5386), .IN2(g6573), .Q(n1324) );
  AND2X1 U12025 ( .IN1(test_so71), .IN2(n8808), .Q(n11722) );
  OR3X1 U12026 ( .IN1(n11726), .IN2(n11727), .IN3(n11728), .Q(g30548) );
  AND2X1 U12027 ( .IN1(n3785), .IN2(n11696), .Q(n11728) );
  INVX0 U12028 ( .INP(n1326), .ZN(n11696) );
  AND3X1 U12029 ( .IN1(n11729), .IN2(g6609), .IN3(n8743), .Q(n11727) );
  OR2X1 U12030 ( .IN1(n3407), .IN2(n1326), .Q(n11729) );
  OR2X1 U12031 ( .IN1(g6565), .IN2(g6573), .Q(n1326) );
  OR2X1 U12032 ( .IN1(n5571), .IN2(g6555), .Q(n3407) );
  AND2X1 U12033 ( .IN1(n8840), .IN2(g6581), .Q(n11726) );
  OR3X1 U12034 ( .IN1(n11730), .IN2(n11731), .IN3(n11732), .Q(g30547) );
  AND2X1 U12035 ( .IN1(n8840), .IN2(g6605), .Q(n11732) );
  AND2X1 U12036 ( .IN1(n3790), .IN2(n3765), .Q(n11731) );
  AND3X1 U12037 ( .IN1(n8728), .IN2(g6601), .IN3(n11733), .Q(n11730) );
  INVX0 U12038 ( .INP(n3790), .ZN(n11733) );
  OR3X1 U12039 ( .IN1(n11734), .IN2(n11735), .IN3(n11736), .Q(g30546) );
  AND2X1 U12040 ( .IN1(n8840), .IN2(g6597), .Q(n11736) );
  AND2X1 U12041 ( .IN1(n3793), .IN2(n3765), .Q(n11735) );
  AND3X1 U12042 ( .IN1(n8728), .IN2(g6593), .IN3(n11737), .Q(n11734) );
  INVX0 U12043 ( .INP(n3793), .ZN(n11737) );
  OR3X1 U12044 ( .IN1(n11738), .IN2(n11739), .IN3(n11740), .Q(g30545) );
  AND2X1 U12045 ( .IN1(n8840), .IN2(g6589), .Q(n11740) );
  AND2X1 U12046 ( .IN1(n3795), .IN2(n3765), .Q(n11739) );
  AND3X1 U12047 ( .IN1(test_so71), .IN2(n8725), .IN3(n11741), .Q(n11738) );
  INVX0 U12048 ( .INP(n3795), .ZN(n11741) );
  OR3X1 U12049 ( .IN1(n11742), .IN2(n11743), .IN3(n11744), .Q(g30544) );
  AND2X1 U12050 ( .IN1(n8840), .IN2(g6573), .Q(n11744) );
  AND2X1 U12051 ( .IN1(n3797), .IN2(n3765), .Q(n11743) );
  AND3X1 U12052 ( .IN1(n8729), .IN2(g6581), .IN3(n11745), .Q(n11742) );
  INVX0 U12053 ( .INP(n3797), .ZN(n11745) );
  AND2X1 U12054 ( .IN1(n11134), .IN2(n5571), .Q(g30543) );
  AND3X1 U12055 ( .IN1(n8729), .IN2(n11127), .IN3(n5646), .Q(n11134) );
  OR2X1 U12056 ( .IN1(n11746), .IN2(n11747), .Q(n11127) );
  OR3X1 U12057 ( .IN1(n11748), .IN2(n11749), .IN3(n11750), .Q(g30542) );
  AND2X1 U12058 ( .IN1(n8840), .IN2(g6307), .Q(n11750) );
  AND2X1 U12059 ( .IN1(n10581), .IN2(n3765), .Q(n11749) );
  AND2X1 U12060 ( .IN1(n11751), .IN2(g6311), .Q(n11748) );
  OR3X1 U12061 ( .IN1(n11752), .IN2(n11753), .IN3(n11754), .Q(g30541) );
  AND2X1 U12062 ( .IN1(n11755), .IN2(n3765), .Q(n11754) );
  INVX0 U12063 ( .INP(n11756), .ZN(n11755) );
  AND2X1 U12064 ( .IN1(n8840), .IN2(g6303), .Q(n11753) );
  AND3X1 U12065 ( .IN1(n11756), .IN2(g6259), .IN3(n8743), .Q(n11752) );
  OR2X1 U12066 ( .IN1(n5651), .IN2(n43), .Q(n11756) );
  OR3X1 U12067 ( .IN1(n11757), .IN2(n11758), .IN3(n11759), .Q(g30540) );
  AND2X1 U12068 ( .IN1(n11149), .IN2(n3765), .Q(n11759) );
  INVX0 U12069 ( .INP(n11760), .ZN(n11149) );
  AND2X1 U12070 ( .IN1(n8840), .IN2(g6299), .Q(n11758) );
  AND3X1 U12071 ( .IN1(n11760), .IN2(g6251), .IN3(n8743), .Q(n11757) );
  OR2X1 U12072 ( .IN1(n5651), .IN2(n51), .Q(n11760) );
  OR3X1 U12073 ( .IN1(n11761), .IN2(n11762), .IN3(n11763), .Q(g30539) );
  AND2X1 U12074 ( .IN1(n11764), .IN2(n3765), .Q(n11763) );
  INVX0 U12075 ( .INP(n11765), .ZN(n11764) );
  AND2X1 U12076 ( .IN1(n8840), .IN2(g6295), .Q(n11762) );
  AND3X1 U12077 ( .IN1(n11765), .IN2(g6243), .IN3(n8743), .Q(n11761) );
  OR2X1 U12078 ( .IN1(n5651), .IN2(n45), .Q(n11765) );
  OR3X1 U12079 ( .IN1(n11766), .IN2(n11767), .IN3(n11768), .Q(g30538) );
  AND2X1 U12080 ( .IN1(n3808), .IN2(n11769), .Q(n11768) );
  AND3X1 U12081 ( .IN1(n11770), .IN2(g6307), .IN3(n8743), .Q(n11767) );
  OR2X1 U12082 ( .IN1(n952), .IN2(n50), .Q(n11770) );
  AND2X1 U12083 ( .IN1(n8840), .IN2(g6291), .Q(n11766) );
  OR3X1 U12084 ( .IN1(n11771), .IN2(n11772), .IN3(n11773), .Q(g30537) );
  AND2X1 U12085 ( .IN1(n3808), .IN2(n11152), .Q(n11773) );
  AND3X1 U12086 ( .IN1(n11774), .IN2(g6303), .IN3(n8743), .Q(n11772) );
  OR2X1 U12087 ( .IN1(n952), .IN2(n43), .Q(n11774) );
  AND2X1 U12088 ( .IN1(n8840), .IN2(g6287), .Q(n11771) );
  OR3X1 U12089 ( .IN1(n11775), .IN2(n11776), .IN3(n11777), .Q(g30536) );
  AND2X1 U12090 ( .IN1(n3808), .IN2(n11778), .Q(n11777) );
  AND3X1 U12091 ( .IN1(n11779), .IN2(g6299), .IN3(n8743), .Q(n11776) );
  OR2X1 U12092 ( .IN1(n952), .IN2(n51), .Q(n11779) );
  AND2X1 U12093 ( .IN1(n8840), .IN2(g6283), .Q(n11775) );
  OR3X1 U12094 ( .IN1(n11780), .IN2(n11781), .IN3(n11782), .Q(g30535) );
  AND2X1 U12095 ( .IN1(n3808), .IN2(n11783), .Q(n11782) );
  AND3X1 U12096 ( .IN1(n11784), .IN2(g6295), .IN3(n8743), .Q(n11781) );
  OR2X1 U12097 ( .IN1(n952), .IN2(n45), .Q(n11784) );
  OR2X1 U12098 ( .IN1(n8312), .IN2(n5574), .Q(n952) );
  AND2X1 U12099 ( .IN1(n8840), .IN2(g6279), .Q(n11780) );
  OR3X1 U12100 ( .IN1(n11785), .IN2(n11786), .IN3(n11787), .Q(g30534) );
  AND2X1 U12101 ( .IN1(n3814), .IN2(n11769), .Q(n11787) );
  AND3X1 U12102 ( .IN1(n11788), .IN2(g6291), .IN3(n8744), .Q(n11786) );
  OR2X1 U12103 ( .IN1(n50), .IN2(n3416), .Q(n11788) );
  AND2X1 U12104 ( .IN1(n8840), .IN2(g6275), .Q(n11785) );
  OR3X1 U12105 ( .IN1(n11789), .IN2(n11790), .IN3(n11791), .Q(g30533) );
  AND2X1 U12106 ( .IN1(n3814), .IN2(n11152), .Q(n11791) );
  AND3X1 U12107 ( .IN1(n11792), .IN2(g6287), .IN3(n8744), .Q(n11790) );
  OR2X1 U12108 ( .IN1(n43), .IN2(n3416), .Q(n11792) );
  AND2X1 U12109 ( .IN1(n8840), .IN2(g6271), .Q(n11789) );
  OR3X1 U12110 ( .IN1(n11793), .IN2(n11794), .IN3(n11795), .Q(g30532) );
  AND2X1 U12111 ( .IN1(n3814), .IN2(n11778), .Q(n11795) );
  AND3X1 U12112 ( .IN1(n11796), .IN2(g6283), .IN3(n8744), .Q(n11794) );
  OR2X1 U12113 ( .IN1(n51), .IN2(n3416), .Q(n11796) );
  AND2X1 U12114 ( .IN1(n8840), .IN2(g6267), .Q(n11793) );
  OR3X1 U12115 ( .IN1(n11797), .IN2(n11798), .IN3(n11799), .Q(g30531) );
  AND2X1 U12116 ( .IN1(n3814), .IN2(n11783), .Q(n11799) );
  AND3X1 U12117 ( .IN1(n11800), .IN2(g6279), .IN3(n8744), .Q(n11798) );
  OR2X1 U12118 ( .IN1(n45), .IN2(n3416), .Q(n11800) );
  OR2X1 U12119 ( .IN1(n8312), .IN2(g6203), .Q(n3416) );
  AND2X1 U12120 ( .IN1(n8841), .IN2(g6263), .Q(n11797) );
  OR3X1 U12121 ( .IN1(n11801), .IN2(n11802), .IN3(n11803), .Q(g30530) );
  AND2X1 U12122 ( .IN1(n3819), .IN2(n11769), .Q(n11803) );
  AND3X1 U12123 ( .IN1(n11804), .IN2(g6275), .IN3(n8744), .Q(n11802) );
  OR2X1 U12124 ( .IN1(n50), .IN2(n3417), .Q(n11804) );
  AND2X1 U12125 ( .IN1(n8841), .IN2(g6255), .Q(n11801) );
  OR3X1 U12126 ( .IN1(n11805), .IN2(n11806), .IN3(n11807), .Q(g30529) );
  AND2X1 U12127 ( .IN1(n3819), .IN2(n11152), .Q(n11807) );
  INVX0 U12128 ( .INP(n43), .ZN(n11152) );
  AND3X1 U12129 ( .IN1(n11808), .IN2(g6271), .IN3(n8744), .Q(n11806) );
  OR2X1 U12130 ( .IN1(n43), .IN2(n3417), .Q(n11808) );
  OR2X1 U12131 ( .IN1(n5568), .IN2(g6219), .Q(n43) );
  AND2X1 U12132 ( .IN1(n8841), .IN2(g6247), .Q(n11805) );
  OR3X1 U12133 ( .IN1(n11809), .IN2(n11810), .IN3(n11811), .Q(g30528) );
  AND2X1 U12134 ( .IN1(n3819), .IN2(n11778), .Q(n11811) );
  INVX0 U12135 ( .INP(n51), .ZN(n11778) );
  AND3X1 U12136 ( .IN1(n11812), .IN2(g6267), .IN3(n8744), .Q(n11810) );
  OR2X1 U12137 ( .IN1(n51), .IN2(n3417), .Q(n11812) );
  OR2X1 U12138 ( .IN1(n5385), .IN2(g6227), .Q(n51) );
  AND2X1 U12139 ( .IN1(n8841), .IN2(g6239), .Q(n11809) );
  OR3X1 U12140 ( .IN1(n11813), .IN2(n11814), .IN3(n11815), .Q(g30527) );
  AND2X1 U12141 ( .IN1(n3819), .IN2(n11783), .Q(n11815) );
  INVX0 U12142 ( .INP(n45), .ZN(n11783) );
  AND3X1 U12143 ( .IN1(n11816), .IN2(g6263), .IN3(n8744), .Q(n11814) );
  OR2X1 U12144 ( .IN1(n45), .IN2(n3417), .Q(n11816) );
  OR2X1 U12145 ( .IN1(n5574), .IN2(g6209), .Q(n3417) );
  OR2X1 U12146 ( .IN1(g6227), .IN2(g6219), .Q(n45) );
  AND2X1 U12147 ( .IN1(n8841), .IN2(g6235), .Q(n11813) );
  OR3X1 U12148 ( .IN1(n11817), .IN2(n11818), .IN3(n11819), .Q(g30526) );
  AND2X1 U12149 ( .IN1(n8841), .IN2(g6259), .Q(n11819) );
  AND2X1 U12150 ( .IN1(n3824), .IN2(n3765), .Q(n11818) );
  AND3X1 U12151 ( .IN1(n8729), .IN2(g6255), .IN3(n11820), .Q(n11817) );
  INVX0 U12152 ( .INP(n3824), .ZN(n11820) );
  OR3X1 U12153 ( .IN1(n11821), .IN2(n11822), .IN3(n11823), .Q(g30525) );
  AND2X1 U12154 ( .IN1(n8834), .IN2(g6251), .Q(n11823) );
  AND2X1 U12155 ( .IN1(n3827), .IN2(n3765), .Q(n11822) );
  AND3X1 U12156 ( .IN1(n8729), .IN2(g6247), .IN3(n11824), .Q(n11821) );
  INVX0 U12157 ( .INP(n3827), .ZN(n11824) );
  OR3X1 U12158 ( .IN1(n11825), .IN2(n11826), .IN3(n11827), .Q(g30524) );
  AND2X1 U12159 ( .IN1(n8831), .IN2(g6243), .Q(n11827) );
  AND2X1 U12160 ( .IN1(n3829), .IN2(n3765), .Q(n11826) );
  AND3X1 U12161 ( .IN1(n8730), .IN2(g6239), .IN3(n11828), .Q(n11825) );
  INVX0 U12162 ( .INP(n3829), .ZN(n11828) );
  OR3X1 U12163 ( .IN1(n11829), .IN2(n11830), .IN3(n11831), .Q(g30523) );
  AND2X1 U12164 ( .IN1(n8832), .IN2(g6227), .Q(n11831) );
  AND2X1 U12165 ( .IN1(n3831), .IN2(n3765), .Q(n11830) );
  AND3X1 U12166 ( .IN1(n8730), .IN2(g6235), .IN3(n11832), .Q(n11829) );
  INVX0 U12167 ( .INP(n3831), .ZN(n11832) );
  AND2X1 U12168 ( .IN1(n11155), .IN2(n5574), .Q(g30522) );
  AND3X1 U12169 ( .IN1(n8729), .IN2(n11148), .IN3(n5651), .Q(n11155) );
  OR3X1 U12170 ( .IN1(n5480), .IN2(n5340), .IN3(n11833), .Q(n11148) );
  OR3X1 U12171 ( .IN1(n11834), .IN2(n11835), .IN3(n11836), .Q(g30521) );
  AND2X1 U12172 ( .IN1(n8832), .IN2(g5961), .Q(n11836) );
  AND2X1 U12173 ( .IN1(n10580), .IN2(n3765), .Q(n11835) );
  AND2X1 U12174 ( .IN1(test_so13), .IN2(n11837), .Q(n11834) );
  OR3X1 U12175 ( .IN1(n11838), .IN2(n11839), .IN3(n11840), .Q(g30520) );
  AND2X1 U12176 ( .IN1(n11841), .IN2(n3765), .Q(n11840) );
  INVX0 U12177 ( .INP(n11842), .ZN(n11841) );
  AND2X1 U12178 ( .IN1(n8832), .IN2(g5957), .Q(n11839) );
  AND3X1 U12179 ( .IN1(n11842), .IN2(g5913), .IN3(n8744), .Q(n11838) );
  OR2X1 U12180 ( .IN1(n5649), .IN2(n666), .Q(n11842) );
  OR3X1 U12181 ( .IN1(n11843), .IN2(n11844), .IN3(n11845), .Q(g30519) );
  AND2X1 U12182 ( .IN1(n11170), .IN2(n3765), .Q(n11845) );
  INVX0 U12183 ( .INP(n11846), .ZN(n11170) );
  AND2X1 U12184 ( .IN1(n8832), .IN2(g5953), .Q(n11844) );
  AND3X1 U12185 ( .IN1(n11846), .IN2(g5905), .IN3(n8745), .Q(n11843) );
  OR2X1 U12186 ( .IN1(n5649), .IN2(n672), .Q(n11846) );
  OR3X1 U12187 ( .IN1(n11847), .IN2(n11848), .IN3(n11849), .Q(g30518) );
  AND2X1 U12188 ( .IN1(n11850), .IN2(n3765), .Q(n11849) );
  INVX0 U12189 ( .INP(n11851), .ZN(n11850) );
  AND2X1 U12190 ( .IN1(n8832), .IN2(g5949), .Q(n11848) );
  AND3X1 U12191 ( .IN1(n11851), .IN2(g5897), .IN3(n8745), .Q(n11847) );
  OR2X1 U12192 ( .IN1(n5649), .IN2(n668), .Q(n11851) );
  OR3X1 U12193 ( .IN1(n11852), .IN2(n11853), .IN3(n11854), .Q(g30517) );
  AND2X1 U12194 ( .IN1(n3842), .IN2(n11855), .Q(n11854) );
  AND3X1 U12195 ( .IN1(n11856), .IN2(g5961), .IN3(n8745), .Q(n11853) );
  OR2X1 U12196 ( .IN1(n671), .IN2(n1011), .Q(n11856) );
  AND2X1 U12197 ( .IN1(n8832), .IN2(g5945), .Q(n11852) );
  OR3X1 U12198 ( .IN1(n11857), .IN2(n11858), .IN3(n11859), .Q(g30516) );
  AND2X1 U12199 ( .IN1(n3842), .IN2(n11173), .Q(n11859) );
  AND3X1 U12200 ( .IN1(n11860), .IN2(g5957), .IN3(n8745), .Q(n11858) );
  OR2X1 U12201 ( .IN1(n666), .IN2(n1011), .Q(n11860) );
  AND2X1 U12202 ( .IN1(n8832), .IN2(g5941), .Q(n11857) );
  OR3X1 U12203 ( .IN1(n11861), .IN2(n11862), .IN3(n11863), .Q(g30515) );
  AND2X1 U12204 ( .IN1(n3842), .IN2(n11864), .Q(n11863) );
  AND3X1 U12205 ( .IN1(n11865), .IN2(g5953), .IN3(n8745), .Q(n11862) );
  OR2X1 U12206 ( .IN1(n672), .IN2(n1011), .Q(n11865) );
  AND2X1 U12207 ( .IN1(n8832), .IN2(g5937), .Q(n11861) );
  OR3X1 U12208 ( .IN1(n11866), .IN2(n11867), .IN3(n11868), .Q(g30514) );
  AND2X1 U12209 ( .IN1(n3842), .IN2(n11869), .Q(n11868) );
  AND3X1 U12210 ( .IN1(n11870), .IN2(g5949), .IN3(n8745), .Q(n11867) );
  OR2X1 U12211 ( .IN1(n668), .IN2(n1011), .Q(n11870) );
  OR2X1 U12212 ( .IN1(n8309), .IN2(n5573), .Q(n1011) );
  AND2X1 U12213 ( .IN1(n8832), .IN2(g5933), .Q(n11866) );
  OR3X1 U12214 ( .IN1(n11871), .IN2(n11872), .IN3(n11873), .Q(g30513) );
  AND2X1 U12215 ( .IN1(n3848), .IN2(n11855), .Q(n11873) );
  AND3X1 U12216 ( .IN1(n11874), .IN2(g5945), .IN3(n8745), .Q(n11872) );
  OR2X1 U12217 ( .IN1(n671), .IN2(n3426), .Q(n11874) );
  AND2X1 U12218 ( .IN1(n8832), .IN2(g5929), .Q(n11871) );
  OR3X1 U12219 ( .IN1(n11875), .IN2(n11876), .IN3(n11877), .Q(g30512) );
  AND2X1 U12220 ( .IN1(n3848), .IN2(n11173), .Q(n11877) );
  AND3X1 U12221 ( .IN1(n11878), .IN2(g5941), .IN3(n8745), .Q(n11876) );
  OR2X1 U12222 ( .IN1(n666), .IN2(n3426), .Q(n11878) );
  AND2X1 U12223 ( .IN1(n8832), .IN2(g5925), .Q(n11875) );
  OR3X1 U12224 ( .IN1(n11879), .IN2(n11880), .IN3(n11881), .Q(g30511) );
  AND2X1 U12225 ( .IN1(n3848), .IN2(n11864), .Q(n11881) );
  AND3X1 U12226 ( .IN1(n11882), .IN2(g5937), .IN3(n8745), .Q(n11880) );
  OR2X1 U12227 ( .IN1(n672), .IN2(n3426), .Q(n11882) );
  AND2X1 U12228 ( .IN1(n8832), .IN2(g5921), .Q(n11879) );
  OR3X1 U12229 ( .IN1(n11883), .IN2(n11884), .IN3(n11885), .Q(g30510) );
  AND2X1 U12230 ( .IN1(n3848), .IN2(n11869), .Q(n11885) );
  AND3X1 U12231 ( .IN1(n11886), .IN2(g5933), .IN3(n8746), .Q(n11884) );
  OR2X1 U12232 ( .IN1(n668), .IN2(n3426), .Q(n11886) );
  OR2X1 U12233 ( .IN1(n8309), .IN2(g5857), .Q(n3426) );
  AND2X1 U12234 ( .IN1(test_so28), .IN2(n8809), .Q(n11883) );
  OR3X1 U12235 ( .IN1(n11887), .IN2(n11888), .IN3(n11889), .Q(g30509) );
  AND2X1 U12236 ( .IN1(n3853), .IN2(n11855), .Q(n11889) );
  AND3X1 U12237 ( .IN1(n11890), .IN2(g5929), .IN3(n8746), .Q(n11888) );
  OR2X1 U12238 ( .IN1(n671), .IN2(n3427), .Q(n11890) );
  AND2X1 U12239 ( .IN1(n8832), .IN2(g5909), .Q(n11887) );
  OR3X1 U12240 ( .IN1(n11891), .IN2(n11892), .IN3(n11893), .Q(g30508) );
  AND2X1 U12241 ( .IN1(n3853), .IN2(n11173), .Q(n11893) );
  INVX0 U12242 ( .INP(n666), .ZN(n11173) );
  AND3X1 U12243 ( .IN1(n11894), .IN2(g5925), .IN3(n8746), .Q(n11892) );
  OR2X1 U12244 ( .IN1(n666), .IN2(n3427), .Q(n11894) );
  OR2X1 U12245 ( .IN1(n8500), .IN2(g5873), .Q(n666) );
  AND2X1 U12246 ( .IN1(n8832), .IN2(g5901), .Q(n11891) );
  OR3X1 U12247 ( .IN1(n11895), .IN2(n11896), .IN3(n11897), .Q(g30507) );
  AND2X1 U12248 ( .IN1(n3853), .IN2(n11864), .Q(n11897) );
  INVX0 U12249 ( .INP(n672), .ZN(n11864) );
  AND3X1 U12250 ( .IN1(n11898), .IN2(g5921), .IN3(n8746), .Q(n11896) );
  OR2X1 U12251 ( .IN1(n672), .IN2(n3427), .Q(n11898) );
  OR2X1 U12252 ( .IN1(test_so36), .IN2(n5388), .Q(n672) );
  AND2X1 U12253 ( .IN1(n8832), .IN2(g5893), .Q(n11895) );
  OR3X1 U12254 ( .IN1(n11899), .IN2(n11900), .IN3(n11901), .Q(g30506) );
  AND2X1 U12255 ( .IN1(n3853), .IN2(n11869), .Q(n11901) );
  INVX0 U12256 ( .INP(n668), .ZN(n11869) );
  AND3X1 U12257 ( .IN1(test_so28), .IN2(n11902), .IN3(n8746), .Q(n11900) );
  OR2X1 U12258 ( .IN1(n668), .IN2(n3427), .Q(n11902) );
  OR2X1 U12259 ( .IN1(n5573), .IN2(g5863), .Q(n3427) );
  OR2X1 U12260 ( .IN1(test_so36), .IN2(g5873), .Q(n668) );
  AND2X1 U12261 ( .IN1(n8832), .IN2(g5889), .Q(n11899) );
  OR3X1 U12262 ( .IN1(n11903), .IN2(n11904), .IN3(n11905), .Q(g30505) );
  AND2X1 U12263 ( .IN1(n8832), .IN2(g5913), .Q(n11905) );
  AND2X1 U12264 ( .IN1(n3858), .IN2(n3765), .Q(n11904) );
  AND3X1 U12265 ( .IN1(n8729), .IN2(g5909), .IN3(n11906), .Q(n11903) );
  INVX0 U12266 ( .INP(n3858), .ZN(n11906) );
  OR3X1 U12267 ( .IN1(n11907), .IN2(n11908), .IN3(n11909), .Q(g30504) );
  AND2X1 U12268 ( .IN1(n8832), .IN2(g5905), .Q(n11909) );
  AND2X1 U12269 ( .IN1(n3861), .IN2(n3765), .Q(n11908) );
  AND3X1 U12270 ( .IN1(n8730), .IN2(g5901), .IN3(n11910), .Q(n11907) );
  INVX0 U12271 ( .INP(n3861), .ZN(n11910) );
  OR3X1 U12272 ( .IN1(n11911), .IN2(n11912), .IN3(n11913), .Q(g30503) );
  AND2X1 U12273 ( .IN1(n8832), .IN2(g5897), .Q(n11913) );
  AND2X1 U12274 ( .IN1(n3863), .IN2(n3765), .Q(n11912) );
  AND3X1 U12275 ( .IN1(n8730), .IN2(g5893), .IN3(n11914), .Q(n11911) );
  INVX0 U12276 ( .INP(n3863), .ZN(n11914) );
  OR3X1 U12277 ( .IN1(n11915), .IN2(n11916), .IN3(n11917), .Q(g30502) );
  AND2X1 U12278 ( .IN1(test_so36), .IN2(n8810), .Q(n11917) );
  AND2X1 U12279 ( .IN1(n3865), .IN2(n3765), .Q(n11916) );
  AND3X1 U12280 ( .IN1(n8730), .IN2(g5889), .IN3(n11918), .Q(n11915) );
  INVX0 U12281 ( .INP(n3865), .ZN(n11918) );
  AND2X1 U12282 ( .IN1(n11176), .IN2(n5573), .Q(g30501) );
  AND3X1 U12283 ( .IN1(n8729), .IN2(n11169), .IN3(n5649), .Q(n11176) );
  OR3X1 U12284 ( .IN1(n5340), .IN2(g4087), .IN3(n11833), .Q(n11169) );
  OR3X1 U12285 ( .IN1(n11919), .IN2(n11920), .IN3(n11921), .Q(g30500) );
  AND2X1 U12286 ( .IN1(n8832), .IN2(g5615), .Q(n11921) );
  AND2X1 U12287 ( .IN1(n3765), .IN2(n10577), .Q(n11920) );
  AND2X1 U12288 ( .IN1(n11922), .IN2(g5619), .Q(n11919) );
  OR3X1 U12289 ( .IN1(n11923), .IN2(n11924), .IN3(n11925), .Q(g30499) );
  AND2X1 U12290 ( .IN1(n11926), .IN2(n3765), .Q(n11925) );
  INVX0 U12291 ( .INP(n11927), .ZN(n11926) );
  AND2X1 U12292 ( .IN1(n8832), .IN2(g5611), .Q(n11924) );
  AND3X1 U12293 ( .IN1(n11927), .IN2(g5567), .IN3(n8746), .Q(n11923) );
  OR2X1 U12294 ( .IN1(n5647), .IN2(n878), .Q(n11927) );
  OR3X1 U12295 ( .IN1(n11928), .IN2(n11929), .IN3(n11930), .Q(g30498) );
  AND2X1 U12296 ( .IN1(n11191), .IN2(n3765), .Q(n11930) );
  INVX0 U12297 ( .INP(n11931), .ZN(n11191) );
  AND2X1 U12298 ( .IN1(n8832), .IN2(g5607), .Q(n11929) );
  AND3X1 U12299 ( .IN1(test_so6), .IN2(n11931), .IN3(n8746), .Q(n11928) );
  OR2X1 U12300 ( .IN1(n5647), .IN2(n875), .Q(n11931) );
  OR3X1 U12301 ( .IN1(n11932), .IN2(n11933), .IN3(n11934), .Q(g30497) );
  AND2X1 U12302 ( .IN1(n11935), .IN2(n3765), .Q(n11934) );
  INVX0 U12303 ( .INP(n11936), .ZN(n11935) );
  AND2X1 U12304 ( .IN1(n8833), .IN2(g5603), .Q(n11933) );
  AND3X1 U12305 ( .IN1(n11936), .IN2(g5551), .IN3(n8746), .Q(n11932) );
  OR2X1 U12306 ( .IN1(n5647), .IN2(n876), .Q(n11936) );
  OR3X1 U12307 ( .IN1(n11937), .IN2(n11938), .IN3(n11939), .Q(g30496) );
  AND2X1 U12308 ( .IN1(n3875), .IN2(n11940), .Q(n11939) );
  AND3X1 U12309 ( .IN1(n11941), .IN2(g5615), .IN3(n8746), .Q(n11938) );
  OR2X1 U12310 ( .IN1(n877), .IN2(n473), .Q(n11941) );
  AND2X1 U12311 ( .IN1(n8833), .IN2(g5599), .Q(n11937) );
  OR3X1 U12312 ( .IN1(n11942), .IN2(n11943), .IN3(n11944), .Q(g30495) );
  AND2X1 U12313 ( .IN1(n3875), .IN2(n11194), .Q(n11944) );
  AND3X1 U12314 ( .IN1(n11945), .IN2(g5611), .IN3(n8746), .Q(n11943) );
  OR2X1 U12315 ( .IN1(n878), .IN2(n473), .Q(n11945) );
  AND2X1 U12316 ( .IN1(n8833), .IN2(g5595), .Q(n11942) );
  OR3X1 U12317 ( .IN1(n11946), .IN2(n11947), .IN3(n11948), .Q(g30494) );
  AND2X1 U12318 ( .IN1(n3875), .IN2(n11949), .Q(n11948) );
  AND3X1 U12319 ( .IN1(n11950), .IN2(g5607), .IN3(n8746), .Q(n11947) );
  OR2X1 U12320 ( .IN1(n875), .IN2(n473), .Q(n11950) );
  AND2X1 U12321 ( .IN1(test_so5), .IN2(n8809), .Q(n11946) );
  OR3X1 U12322 ( .IN1(n11951), .IN2(n11952), .IN3(n11953), .Q(g30493) );
  AND2X1 U12323 ( .IN1(n3875), .IN2(n11954), .Q(n11953) );
  AND3X1 U12324 ( .IN1(n11955), .IN2(g5603), .IN3(n8748), .Q(n11952) );
  OR2X1 U12325 ( .IN1(n876), .IN2(n473), .Q(n11955) );
  OR2X1 U12326 ( .IN1(n8311), .IN2(n5575), .Q(n473) );
  AND2X1 U12327 ( .IN1(n8833), .IN2(g5587), .Q(n11951) );
  OR3X1 U12328 ( .IN1(n11956), .IN2(n11957), .IN3(n11958), .Q(g30492) );
  AND2X1 U12329 ( .IN1(n3881), .IN2(n11940), .Q(n11958) );
  AND3X1 U12330 ( .IN1(n11959), .IN2(g5599), .IN3(n8749), .Q(n11957) );
  OR2X1 U12331 ( .IN1(n877), .IN2(n3436), .Q(n11959) );
  AND2X1 U12332 ( .IN1(n8833), .IN2(g5583), .Q(n11956) );
  OR3X1 U12333 ( .IN1(n11960), .IN2(n11961), .IN3(n11962), .Q(g30491) );
  AND2X1 U12334 ( .IN1(n3881), .IN2(n11194), .Q(n11962) );
  AND3X1 U12335 ( .IN1(n11963), .IN2(g5595), .IN3(n8750), .Q(n11961) );
  OR2X1 U12336 ( .IN1(n878), .IN2(n3436), .Q(n11963) );
  AND2X1 U12337 ( .IN1(n8833), .IN2(g5579), .Q(n11960) );
  OR3X1 U12338 ( .IN1(n11964), .IN2(n11965), .IN3(n11966), .Q(g30490) );
  AND2X1 U12339 ( .IN1(n3881), .IN2(n11949), .Q(n11966) );
  AND3X1 U12340 ( .IN1(test_so5), .IN2(n11967), .IN3(n8751), .Q(n11965) );
  OR2X1 U12341 ( .IN1(n875), .IN2(n3436), .Q(n11967) );
  AND2X1 U12342 ( .IN1(n8833), .IN2(g5575), .Q(n11964) );
  OR3X1 U12343 ( .IN1(n11968), .IN2(n11969), .IN3(n11970), .Q(g30489) );
  AND2X1 U12344 ( .IN1(n3881), .IN2(n11954), .Q(n11970) );
  AND3X1 U12345 ( .IN1(n11971), .IN2(g5587), .IN3(n8751), .Q(n11969) );
  OR2X1 U12346 ( .IN1(n876), .IN2(n3436), .Q(n11971) );
  OR2X1 U12347 ( .IN1(n8311), .IN2(g5511), .Q(n3436) );
  AND2X1 U12348 ( .IN1(n8833), .IN2(g5571), .Q(n11968) );
  OR3X1 U12349 ( .IN1(n11972), .IN2(n11973), .IN3(n11974), .Q(g30488) );
  AND2X1 U12350 ( .IN1(n3886), .IN2(n11940), .Q(n11974) );
  AND3X1 U12351 ( .IN1(n11975), .IN2(g5583), .IN3(n8751), .Q(n11973) );
  OR2X1 U12352 ( .IN1(n877), .IN2(n3437), .Q(n11975) );
  AND2X1 U12353 ( .IN1(n8833), .IN2(g5563), .Q(n11972) );
  OR3X1 U12354 ( .IN1(n11976), .IN2(n11977), .IN3(n11978), .Q(g30487) );
  AND2X1 U12355 ( .IN1(n3886), .IN2(n11194), .Q(n11978) );
  INVX0 U12356 ( .INP(n878), .ZN(n11194) );
  AND3X1 U12357 ( .IN1(n11979), .IN2(g5579), .IN3(n8751), .Q(n11977) );
  OR2X1 U12358 ( .IN1(n878), .IN2(n3437), .Q(n11979) );
  OR2X1 U12359 ( .IN1(n5566), .IN2(g5527), .Q(n878) );
  AND2X1 U12360 ( .IN1(n8833), .IN2(g5555), .Q(n11976) );
  OR3X1 U12361 ( .IN1(n11980), .IN2(n11981), .IN3(n11982), .Q(g30486) );
  AND2X1 U12362 ( .IN1(n3886), .IN2(n11949), .Q(n11982) );
  INVX0 U12363 ( .INP(n875), .ZN(n11949) );
  AND3X1 U12364 ( .IN1(n11983), .IN2(g5575), .IN3(n8752), .Q(n11981) );
  OR2X1 U12365 ( .IN1(n875), .IN2(n3437), .Q(n11983) );
  OR2X1 U12366 ( .IN1(n5389), .IN2(g5535), .Q(n875) );
  AND2X1 U12367 ( .IN1(n8833), .IN2(g5547), .Q(n11980) );
  OR3X1 U12368 ( .IN1(n11984), .IN2(n11985), .IN3(n11986), .Q(g30485) );
  AND2X1 U12369 ( .IN1(n3886), .IN2(n11954), .Q(n11986) );
  INVX0 U12370 ( .INP(n876), .ZN(n11954) );
  AND3X1 U12371 ( .IN1(n11987), .IN2(g5571), .IN3(n8752), .Q(n11985) );
  OR2X1 U12372 ( .IN1(n876), .IN2(n3437), .Q(n11987) );
  OR2X1 U12373 ( .IN1(n5575), .IN2(g5517), .Q(n3437) );
  OR2X1 U12374 ( .IN1(g5527), .IN2(g5535), .Q(n876) );
  AND2X1 U12375 ( .IN1(n8833), .IN2(g5543), .Q(n11984) );
  OR3X1 U12376 ( .IN1(n11988), .IN2(n11989), .IN3(n11990), .Q(g30484) );
  AND2X1 U12377 ( .IN1(n8833), .IN2(g5567), .Q(n11990) );
  AND2X1 U12378 ( .IN1(n3891), .IN2(n3765), .Q(n11989) );
  AND3X1 U12379 ( .IN1(n8727), .IN2(g5563), .IN3(n11991), .Q(n11988) );
  INVX0 U12380 ( .INP(n3891), .ZN(n11991) );
  OR3X1 U12381 ( .IN1(n11992), .IN2(n11993), .IN3(n11994), .Q(g30483) );
  AND2X1 U12382 ( .IN1(test_so6), .IN2(n8809), .Q(n11994) );
  AND2X1 U12383 ( .IN1(n3894), .IN2(n3765), .Q(n11993) );
  AND3X1 U12384 ( .IN1(n8728), .IN2(g5555), .IN3(n11995), .Q(n11992) );
  INVX0 U12385 ( .INP(n3894), .ZN(n11995) );
  OR3X1 U12386 ( .IN1(n11996), .IN2(n11997), .IN3(n11998), .Q(g30482) );
  AND2X1 U12387 ( .IN1(n8833), .IN2(g5551), .Q(n11998) );
  AND2X1 U12388 ( .IN1(n3896), .IN2(n3765), .Q(n11997) );
  AND3X1 U12389 ( .IN1(n8728), .IN2(g5547), .IN3(n11999), .Q(n11996) );
  INVX0 U12390 ( .INP(n3896), .ZN(n11999) );
  OR3X1 U12391 ( .IN1(n12000), .IN2(n12001), .IN3(n12002), .Q(g30481) );
  AND2X1 U12392 ( .IN1(n8833), .IN2(g5535), .Q(n12002) );
  AND2X1 U12393 ( .IN1(n3898), .IN2(n3765), .Q(n12001) );
  AND3X1 U12394 ( .IN1(n8728), .IN2(g5543), .IN3(n12003), .Q(n12000) );
  INVX0 U12395 ( .INP(n3898), .ZN(n12003) );
  AND2X1 U12396 ( .IN1(n11197), .IN2(n5575), .Q(g30480) );
  AND3X1 U12397 ( .IN1(n8728), .IN2(n11190), .IN3(n5647), .Q(n11197) );
  OR2X1 U12398 ( .IN1(n12004), .IN2(n11833), .Q(n11190) );
  OR3X1 U12399 ( .IN1(n12005), .IN2(n12006), .IN3(n12007), .Q(g30479) );
  AND2X1 U12400 ( .IN1(n8833), .IN2(g5268), .Q(n12007) );
  AND2X1 U12401 ( .IN1(n3765), .IN2(g32975), .Q(n12006) );
  AND2X1 U12402 ( .IN1(n9099), .IN2(g5272), .Q(n12005) );
  OR3X1 U12403 ( .IN1(n12008), .IN2(n12009), .IN3(n12010), .Q(g30478) );
  AND2X1 U12404 ( .IN1(n12011), .IN2(n3765), .Q(n12010) );
  INVX0 U12405 ( .INP(n12012), .ZN(n12011) );
  AND2X1 U12406 ( .IN1(n8833), .IN2(g5264), .Q(n12009) );
  AND3X1 U12407 ( .IN1(n12012), .IN2(g5220), .IN3(n8731), .Q(n12008) );
  OR2X1 U12408 ( .IN1(n5650), .IN2(n187), .Q(n12012) );
  OR3X1 U12409 ( .IN1(n12013), .IN2(n12014), .IN3(n12015), .Q(g30477) );
  AND2X1 U12410 ( .IN1(n11212), .IN2(n3765), .Q(n12015) );
  INVX0 U12411 ( .INP(n12016), .ZN(n11212) );
  AND2X1 U12412 ( .IN1(n8833), .IN2(g5260), .Q(n12014) );
  AND3X1 U12413 ( .IN1(n12016), .IN2(g5212), .IN3(n8733), .Q(n12013) );
  OR2X1 U12414 ( .IN1(n5650), .IN2(n196), .Q(n12016) );
  OR3X1 U12415 ( .IN1(n12017), .IN2(n12018), .IN3(n12019), .Q(g30476) );
  AND2X1 U12416 ( .IN1(n12020), .IN2(n3765), .Q(n12019) );
  INVX0 U12417 ( .INP(n12021), .ZN(n12020) );
  AND2X1 U12418 ( .IN1(n8833), .IN2(g5256), .Q(n12018) );
  AND3X1 U12419 ( .IN1(n12021), .IN2(g5204), .IN3(n8731), .Q(n12017) );
  OR2X1 U12420 ( .IN1(n5650), .IN2(n189), .Q(n12021) );
  OR3X1 U12421 ( .IN1(n12022), .IN2(n12023), .IN3(n12024), .Q(g30475) );
  AND2X1 U12422 ( .IN1(n3908), .IN2(n12025), .Q(n12024) );
  AND3X1 U12423 ( .IN1(n12026), .IN2(g5268), .IN3(n8732), .Q(n12023) );
  OR2X1 U12424 ( .IN1(n699), .IN2(n195), .Q(n12026) );
  AND2X1 U12425 ( .IN1(n8833), .IN2(g5252), .Q(n12022) );
  OR3X1 U12426 ( .IN1(n12027), .IN2(n12028), .IN3(n12029), .Q(g30474) );
  AND2X1 U12427 ( .IN1(n3908), .IN2(n11215), .Q(n12029) );
  AND3X1 U12428 ( .IN1(n12030), .IN2(g5264), .IN3(n8731), .Q(n12028) );
  OR2X1 U12429 ( .IN1(n699), .IN2(n187), .Q(n12030) );
  AND2X1 U12430 ( .IN1(n8833), .IN2(g5248), .Q(n12027) );
  OR3X1 U12431 ( .IN1(n12031), .IN2(n12032), .IN3(n12033), .Q(g30473) );
  AND2X1 U12432 ( .IN1(n3908), .IN2(n12034), .Q(n12033) );
  AND3X1 U12433 ( .IN1(n12035), .IN2(g5260), .IN3(n8734), .Q(n12032) );
  OR2X1 U12434 ( .IN1(n699), .IN2(n196), .Q(n12035) );
  AND2X1 U12435 ( .IN1(n8833), .IN2(g5244), .Q(n12031) );
  OR3X1 U12436 ( .IN1(n12036), .IN2(n12037), .IN3(n12038), .Q(g30472) );
  AND2X1 U12437 ( .IN1(n3908), .IN2(n12039), .Q(n12038) );
  AND3X1 U12438 ( .IN1(n12040), .IN2(g5256), .IN3(n8732), .Q(n12037) );
  OR2X1 U12439 ( .IN1(n699), .IN2(n189), .Q(n12040) );
  OR2X1 U12440 ( .IN1(n8313), .IN2(n5570), .Q(n699) );
  AND2X1 U12441 ( .IN1(n8834), .IN2(g5240), .Q(n12036) );
  OR3X1 U12442 ( .IN1(n12041), .IN2(n12042), .IN3(n12043), .Q(g30471) );
  AND2X1 U12443 ( .IN1(n3914), .IN2(n12025), .Q(n12043) );
  AND3X1 U12444 ( .IN1(n12044), .IN2(g5252), .IN3(n8732), .Q(n12042) );
  OR2X1 U12445 ( .IN1(n3446), .IN2(n195), .Q(n12044) );
  AND2X1 U12446 ( .IN1(n8834), .IN2(g5236), .Q(n12041) );
  OR3X1 U12447 ( .IN1(n12045), .IN2(n12046), .IN3(n12047), .Q(g30470) );
  AND2X1 U12448 ( .IN1(n3914), .IN2(n11215), .Q(n12047) );
  AND3X1 U12449 ( .IN1(n12048), .IN2(g5248), .IN3(n8732), .Q(n12046) );
  OR2X1 U12450 ( .IN1(n3446), .IN2(n187), .Q(n12048) );
  AND2X1 U12451 ( .IN1(n8834), .IN2(g5232), .Q(n12045) );
  OR3X1 U12452 ( .IN1(n12049), .IN2(n12050), .IN3(n12051), .Q(g30469) );
  AND2X1 U12453 ( .IN1(n3914), .IN2(n12034), .Q(n12051) );
  AND3X1 U12454 ( .IN1(n12052), .IN2(g5244), .IN3(n8732), .Q(n12050) );
  OR2X1 U12455 ( .IN1(n3446), .IN2(n196), .Q(n12052) );
  AND2X1 U12456 ( .IN1(test_so82), .IN2(n8810), .Q(n12049) );
  OR3X1 U12457 ( .IN1(n12053), .IN2(n12054), .IN3(n12055), .Q(g30468) );
  AND2X1 U12458 ( .IN1(n3914), .IN2(n12039), .Q(n12055) );
  AND3X1 U12459 ( .IN1(n12056), .IN2(g5240), .IN3(n8732), .Q(n12054) );
  OR2X1 U12460 ( .IN1(n3446), .IN2(n189), .Q(n12056) );
  OR2X1 U12461 ( .IN1(n8313), .IN2(g5164), .Q(n3446) );
  AND2X1 U12462 ( .IN1(n8834), .IN2(g5224), .Q(n12053) );
  OR3X1 U12463 ( .IN1(n12057), .IN2(n12058), .IN3(n12059), .Q(g30467) );
  AND2X1 U12464 ( .IN1(n3919), .IN2(n12025), .Q(n12059) );
  AND3X1 U12465 ( .IN1(n12060), .IN2(g5236), .IN3(n8732), .Q(n12058) );
  OR2X1 U12466 ( .IN1(n3447), .IN2(n195), .Q(n12060) );
  AND2X1 U12467 ( .IN1(n8834), .IN2(g5216), .Q(n12057) );
  OR3X1 U12468 ( .IN1(n12061), .IN2(n12062), .IN3(n12063), .Q(g30466) );
  AND2X1 U12469 ( .IN1(n3919), .IN2(n11215), .Q(n12063) );
  INVX0 U12470 ( .INP(n187), .ZN(n11215) );
  AND3X1 U12471 ( .IN1(n12064), .IN2(g5232), .IN3(n8732), .Q(n12062) );
  OR2X1 U12472 ( .IN1(n3447), .IN2(n187), .Q(n12064) );
  OR2X1 U12473 ( .IN1(n5567), .IN2(g5180), .Q(n187) );
  AND2X1 U12474 ( .IN1(n8834), .IN2(g5208), .Q(n12061) );
  OR3X1 U12475 ( .IN1(n12065), .IN2(n12066), .IN3(n12067), .Q(g30465) );
  AND2X1 U12476 ( .IN1(n3919), .IN2(n12034), .Q(n12067) );
  INVX0 U12477 ( .INP(n196), .ZN(n12034) );
  AND3X1 U12478 ( .IN1(test_so82), .IN2(n12068), .IN3(n8734), .Q(n12066) );
  OR2X1 U12479 ( .IN1(n3447), .IN2(n196), .Q(n12068) );
  OR2X1 U12480 ( .IN1(n5384), .IN2(g5188), .Q(n196) );
  AND2X1 U12481 ( .IN1(n8834), .IN2(g5200), .Q(n12065) );
  OR3X1 U12482 ( .IN1(n12069), .IN2(n12070), .IN3(n12071), .Q(g30464) );
  AND2X1 U12483 ( .IN1(n3919), .IN2(n12039), .Q(n12071) );
  INVX0 U12484 ( .INP(n189), .ZN(n12039) );
  AND3X1 U12485 ( .IN1(n12072), .IN2(g5224), .IN3(n8735), .Q(n12070) );
  OR2X1 U12486 ( .IN1(n3447), .IN2(n189), .Q(n12072) );
  OR2X1 U12487 ( .IN1(g5188), .IN2(g5180), .Q(n189) );
  OR2X1 U12488 ( .IN1(n5570), .IN2(g5170), .Q(n3447) );
  AND2X1 U12489 ( .IN1(n8834), .IN2(g5196), .Q(n12069) );
  OR3X1 U12490 ( .IN1(n12073), .IN2(n12074), .IN3(n12075), .Q(g30463) );
  AND2X1 U12491 ( .IN1(n8834), .IN2(g5220), .Q(n12075) );
  AND2X1 U12492 ( .IN1(n3924), .IN2(n3765), .Q(n12074) );
  AND3X1 U12493 ( .IN1(n8729), .IN2(g5216), .IN3(n12076), .Q(n12073) );
  INVX0 U12494 ( .INP(n3924), .ZN(n12076) );
  OR3X1 U12495 ( .IN1(n12077), .IN2(n12078), .IN3(n12079), .Q(g30462) );
  AND2X1 U12496 ( .IN1(n8834), .IN2(g5212), .Q(n12079) );
  AND2X1 U12497 ( .IN1(n3927), .IN2(n3765), .Q(n12078) );
  AND3X1 U12498 ( .IN1(n8727), .IN2(g5208), .IN3(n12080), .Q(n12077) );
  INVX0 U12499 ( .INP(n3927), .ZN(n12080) );
  OR3X1 U12500 ( .IN1(n12081), .IN2(n12082), .IN3(n12083), .Q(g30461) );
  AND2X1 U12501 ( .IN1(n8834), .IN2(g5204), .Q(n12083) );
  AND2X1 U12502 ( .IN1(n3929), .IN2(n3765), .Q(n12082) );
  AND3X1 U12503 ( .IN1(n8729), .IN2(g5200), .IN3(n12084), .Q(n12081) );
  INVX0 U12504 ( .INP(n3929), .ZN(n12084) );
  OR3X1 U12505 ( .IN1(n12085), .IN2(n12086), .IN3(n12087), .Q(g30460) );
  AND2X1 U12506 ( .IN1(n8834), .IN2(g5188), .Q(n12087) );
  AND2X1 U12507 ( .IN1(n3931), .IN2(n3765), .Q(n12086) );
  AND3X1 U12508 ( .IN1(n8728), .IN2(g5196), .IN3(n12088), .Q(n12085) );
  INVX0 U12509 ( .INP(n3931), .ZN(n12088) );
  AND2X1 U12510 ( .IN1(n11218), .IN2(n5570), .Q(g30459) );
  AND3X1 U12511 ( .IN1(n8729), .IN2(n11211), .IN3(n5650), .Q(n11218) );
  OR2X1 U12512 ( .IN1(n11746), .IN2(n11833), .Q(n11211) );
  INVX0 U12513 ( .INP(n3833), .ZN(n11833) );
  OR3X1 U12514 ( .IN1(n12089), .IN2(n12090), .IN3(n8792), .Q(g30458) );
  INVX0 U12515 ( .INP(n12091), .ZN(n12090) );
  OR2X1 U12516 ( .IN1(n12092), .IN2(n5846), .Q(n12091) );
  AND2X1 U12517 ( .IN1(n12092), .IN2(g113), .Q(n12089) );
  AND2X1 U12518 ( .IN1(g4473), .IN2(n5765), .Q(n12092) );
  OR2X1 U12519 ( .IN1(n12093), .IN2(n12094), .Q(g30457) );
  AND2X1 U12520 ( .IN1(n12095), .IN2(n8695), .Q(n12094) );
  OR2X1 U12521 ( .IN1(n12096), .IN2(n12097), .Q(n12095) );
  AND2X1 U12522 ( .IN1(n12098), .IN2(n5983), .Q(n12097) );
  XNOR2X1 U12523 ( .IN1(g115), .IN2(n12099), .Q(n12098) );
  AND2X1 U12524 ( .IN1(n12100), .IN2(n5981), .Q(n12096) );
  XNOR2X1 U12525 ( .IN1(g126), .IN2(n12101), .Q(n12100) );
  AND2X1 U12526 ( .IN1(n8834), .IN2(g4122), .Q(n12093) );
  OR3X1 U12527 ( .IN1(n12102), .IN2(n12103), .IN3(n12104), .Q(g30456) );
  AND2X1 U12528 ( .IN1(n8834), .IN2(g4087), .Q(n12104) );
  AND2X1 U12529 ( .IN1(n3941), .IN2(n12105), .Q(n12103) );
  AND3X1 U12530 ( .IN1(n10568), .IN2(g4169), .IN3(n12106), .Q(n12102) );
  OR3X1 U12531 ( .IN1(n12107), .IN2(n12108), .IN3(n12109), .Q(g30455) );
  AND2X1 U12532 ( .IN1(n8834), .IN2(g3961), .Q(n12109) );
  AND2X1 U12533 ( .IN1(n3765), .IN2(n9012), .Q(n12108) );
  AND2X1 U12534 ( .IN1(n9011), .IN2(g3965), .Q(n12107) );
  OR3X1 U12535 ( .IN1(n12110), .IN2(n12111), .IN3(n12112), .Q(g30454) );
  AND2X1 U12536 ( .IN1(n12113), .IN2(n3765), .Q(n12112) );
  INVX0 U12537 ( .INP(n12114), .ZN(n12113) );
  AND2X1 U12538 ( .IN1(n8834), .IN2(g3957), .Q(n12111) );
  AND3X1 U12539 ( .IN1(n12114), .IN2(g3913), .IN3(n8734), .Q(n12110) );
  OR2X1 U12540 ( .IN1(n770), .IN2(n8493), .Q(n12114) );
  OR3X1 U12541 ( .IN1(n12115), .IN2(n12116), .IN3(n12117), .Q(g30453) );
  AND2X1 U12542 ( .IN1(n11269), .IN2(n3765), .Q(n12117) );
  INVX0 U12543 ( .INP(n12118), .ZN(n11269) );
  AND2X1 U12544 ( .IN1(n8834), .IN2(g3953), .Q(n12116) );
  AND3X1 U12545 ( .IN1(n12118), .IN2(g3905), .IN3(n8734), .Q(n12115) );
  OR2X1 U12546 ( .IN1(n777), .IN2(n8493), .Q(n12118) );
  OR3X1 U12547 ( .IN1(n12119), .IN2(n12120), .IN3(n12121), .Q(g30452) );
  AND2X1 U12548 ( .IN1(n12122), .IN2(n3765), .Q(n12121) );
  INVX0 U12549 ( .INP(n12123), .ZN(n12122) );
  AND2X1 U12550 ( .IN1(test_so65), .IN2(n8810), .Q(n12120) );
  AND3X1 U12551 ( .IN1(n12123), .IN2(g3897), .IN3(n8735), .Q(n12119) );
  OR2X1 U12552 ( .IN1(n772), .IN2(n8493), .Q(n12123) );
  OR3X1 U12553 ( .IN1(n12124), .IN2(n12125), .IN3(n12126), .Q(g30451) );
  AND2X1 U12554 ( .IN1(n3951), .IN2(n12127), .Q(n12126) );
  AND3X1 U12555 ( .IN1(n12128), .IN2(g3961), .IN3(n8734), .Q(n12125) );
  OR2X1 U12556 ( .IN1(n776), .IN2(n1069), .Q(n12128) );
  AND2X1 U12557 ( .IN1(n8834), .IN2(g3945), .Q(n12124) );
  OR3X1 U12558 ( .IN1(n12129), .IN2(n12130), .IN3(n12131), .Q(g30450) );
  AND2X1 U12559 ( .IN1(n3951), .IN2(n11272), .Q(n12131) );
  AND3X1 U12560 ( .IN1(n12132), .IN2(g3957), .IN3(n8734), .Q(n12130) );
  OR2X1 U12561 ( .IN1(n770), .IN2(n1069), .Q(n12132) );
  AND2X1 U12562 ( .IN1(n8834), .IN2(g3941), .Q(n12129) );
  OR3X1 U12563 ( .IN1(n12133), .IN2(n12134), .IN3(n12135), .Q(g30449) );
  AND2X1 U12564 ( .IN1(n3951), .IN2(n12136), .Q(n12135) );
  AND3X1 U12565 ( .IN1(n12137), .IN2(g3953), .IN3(n8734), .Q(n12134) );
  OR2X1 U12566 ( .IN1(n777), .IN2(n1069), .Q(n12137) );
  AND2X1 U12567 ( .IN1(n8834), .IN2(g3937), .Q(n12133) );
  OR3X1 U12568 ( .IN1(n12138), .IN2(n12139), .IN3(n12140), .Q(g30448) );
  AND2X1 U12569 ( .IN1(n3951), .IN2(n12141), .Q(n12140) );
  AND3X1 U12570 ( .IN1(test_so65), .IN2(n12142), .IN3(n8735), .Q(n12139) );
  OR2X1 U12571 ( .IN1(n772), .IN2(n1069), .Q(n12142) );
  OR2X1 U12572 ( .IN1(n8310), .IN2(n5572), .Q(n1069) );
  AND2X1 U12573 ( .IN1(n8834), .IN2(g3933), .Q(n12138) );
  OR3X1 U12574 ( .IN1(n12143), .IN2(n12144), .IN3(n12145), .Q(g30447) );
  AND2X1 U12575 ( .IN1(n3957), .IN2(n12127), .Q(n12145) );
  AND3X1 U12576 ( .IN1(n12146), .IN2(g3945), .IN3(n8735), .Q(n12144) );
  OR2X1 U12577 ( .IN1(n776), .IN2(n3481), .Q(n12146) );
  AND2X1 U12578 ( .IN1(n8835), .IN2(g3929), .Q(n12143) );
  OR3X1 U12579 ( .IN1(n12147), .IN2(n12148), .IN3(n12149), .Q(g30446) );
  AND2X1 U12580 ( .IN1(n3957), .IN2(n11272), .Q(n12149) );
  AND3X1 U12581 ( .IN1(n12150), .IN2(g3941), .IN3(n8735), .Q(n12148) );
  OR2X1 U12582 ( .IN1(n770), .IN2(n3481), .Q(n12150) );
  AND2X1 U12583 ( .IN1(n8835), .IN2(g3925), .Q(n12147) );
  OR3X1 U12584 ( .IN1(n12151), .IN2(n12152), .IN3(n12153), .Q(g30445) );
  AND2X1 U12585 ( .IN1(n3957), .IN2(n12136), .Q(n12153) );
  AND3X1 U12586 ( .IN1(n12154), .IN2(g3937), .IN3(n8735), .Q(n12152) );
  OR2X1 U12587 ( .IN1(n777), .IN2(n3481), .Q(n12154) );
  AND2X1 U12588 ( .IN1(n8835), .IN2(g3921), .Q(n12151) );
  OR3X1 U12589 ( .IN1(n12155), .IN2(n12156), .IN3(n12157), .Q(g30444) );
  AND2X1 U12590 ( .IN1(n3957), .IN2(n12141), .Q(n12157) );
  AND3X1 U12591 ( .IN1(n12158), .IN2(g3933), .IN3(n8741), .Q(n12156) );
  OR2X1 U12592 ( .IN1(n772), .IN2(n3481), .Q(n12158) );
  OR2X1 U12593 ( .IN1(n8310), .IN2(g3857), .Q(n3481) );
  AND2X1 U12594 ( .IN1(n8835), .IN2(g3917), .Q(n12155) );
  OR3X1 U12595 ( .IN1(n12159), .IN2(n12160), .IN3(n12161), .Q(g30443) );
  AND2X1 U12596 ( .IN1(n3962), .IN2(n12127), .Q(n12161) );
  AND3X1 U12597 ( .IN1(n12162), .IN2(g3929), .IN3(n8736), .Q(n12160) );
  OR2X1 U12598 ( .IN1(n776), .IN2(n3482), .Q(n12162) );
  AND2X1 U12599 ( .IN1(n8835), .IN2(g3909), .Q(n12159) );
  OR3X1 U12600 ( .IN1(n12163), .IN2(n12164), .IN3(n12165), .Q(g30442) );
  AND2X1 U12601 ( .IN1(n3962), .IN2(n11272), .Q(n12165) );
  INVX0 U12602 ( .INP(n770), .ZN(n11272) );
  AND3X1 U12603 ( .IN1(n12166), .IN2(g3925), .IN3(n8736), .Q(n12164) );
  OR2X1 U12604 ( .IN1(n770), .IN2(n3482), .Q(n12166) );
  OR2X1 U12605 ( .IN1(n5564), .IN2(g3873), .Q(n770) );
  AND2X1 U12606 ( .IN1(n8835), .IN2(g3901), .Q(n12163) );
  OR3X1 U12607 ( .IN1(n12167), .IN2(n12168), .IN3(n12169), .Q(g30441) );
  AND2X1 U12608 ( .IN1(n3962), .IN2(n12136), .Q(n12169) );
  INVX0 U12609 ( .INP(n777), .ZN(n12136) );
  AND3X1 U12610 ( .IN1(n12170), .IN2(g3921), .IN3(n8736), .Q(n12168) );
  OR2X1 U12611 ( .IN1(n777), .IN2(n3482), .Q(n12170) );
  OR2X1 U12612 ( .IN1(n5387), .IN2(g3881), .Q(n777) );
  AND2X1 U12613 ( .IN1(n8835), .IN2(g3893), .Q(n12167) );
  OR3X1 U12614 ( .IN1(n12171), .IN2(n12172), .IN3(n12173), .Q(g30440) );
  AND2X1 U12615 ( .IN1(n3962), .IN2(n12141), .Q(n12173) );
  INVX0 U12616 ( .INP(n772), .ZN(n12141) );
  AND3X1 U12617 ( .IN1(n12174), .IN2(g3917), .IN3(n8736), .Q(n12172) );
  OR2X1 U12618 ( .IN1(n772), .IN2(n3482), .Q(n12174) );
  OR2X1 U12619 ( .IN1(n5572), .IN2(g3863), .Q(n3482) );
  OR2X1 U12620 ( .IN1(g3881), .IN2(g3873), .Q(n772) );
  AND2X1 U12621 ( .IN1(test_so24), .IN2(n8810), .Q(n12171) );
  OR3X1 U12622 ( .IN1(n12175), .IN2(n12176), .IN3(n12177), .Q(g30439) );
  AND2X1 U12623 ( .IN1(n8835), .IN2(g3913), .Q(n12177) );
  AND2X1 U12624 ( .IN1(n3967), .IN2(n3765), .Q(n12176) );
  AND3X1 U12625 ( .IN1(n8728), .IN2(g3909), .IN3(n12178), .Q(n12175) );
  INVX0 U12626 ( .INP(n3967), .ZN(n12178) );
  OR3X1 U12627 ( .IN1(n12179), .IN2(n12180), .IN3(n12181), .Q(g30438) );
  AND2X1 U12628 ( .IN1(n8835), .IN2(g3905), .Q(n12181) );
  AND2X1 U12629 ( .IN1(n3970), .IN2(n3765), .Q(n12180) );
  AND3X1 U12630 ( .IN1(n8730), .IN2(g3901), .IN3(n12182), .Q(n12179) );
  INVX0 U12631 ( .INP(n3970), .ZN(n12182) );
  OR3X1 U12632 ( .IN1(n12183), .IN2(n12184), .IN3(n12185), .Q(g30437) );
  AND2X1 U12633 ( .IN1(n8835), .IN2(g3897), .Q(n12185) );
  AND2X1 U12634 ( .IN1(n3972), .IN2(n3765), .Q(n12184) );
  AND3X1 U12635 ( .IN1(n8730), .IN2(g3893), .IN3(n12186), .Q(n12183) );
  INVX0 U12636 ( .INP(n3972), .ZN(n12186) );
  OR3X1 U12637 ( .IN1(n12187), .IN2(n12188), .IN3(n12189), .Q(g30436) );
  AND2X1 U12638 ( .IN1(n8835), .IN2(g3881), .Q(n12189) );
  AND2X1 U12639 ( .IN1(n3974), .IN2(n3765), .Q(n12188) );
  AND3X1 U12640 ( .IN1(test_so24), .IN2(n8724), .IN3(n12190), .Q(n12187) );
  INVX0 U12641 ( .INP(n3974), .ZN(n12190) );
  AND2X1 U12642 ( .IN1(n11275), .IN2(n5572), .Q(g30435) );
  AND3X1 U12643 ( .IN1(n8493), .IN2(n8724), .IN3(n11268), .Q(n11275) );
  OR3X1 U12644 ( .IN1(n5480), .IN2(n5340), .IN3(n11747), .Q(n11268) );
  OR3X1 U12645 ( .IN1(n12191), .IN2(n12192), .IN3(n12193), .Q(g30434) );
  AND2X1 U12646 ( .IN1(n8835), .IN2(g3610), .Q(n12193) );
  AND2X1 U12647 ( .IN1(n10572), .IN2(n3765), .Q(n12192) );
  AND2X1 U12648 ( .IN1(n12194), .IN2(g3614), .Q(n12191) );
  OR3X1 U12649 ( .IN1(n12195), .IN2(n12196), .IN3(n12197), .Q(g30433) );
  AND2X1 U12650 ( .IN1(n12198), .IN2(n3765), .Q(n12197) );
  INVX0 U12651 ( .INP(n12199), .ZN(n12198) );
  AND2X1 U12652 ( .IN1(n8835), .IN2(g3606), .Q(n12196) );
  AND3X1 U12653 ( .IN1(n12199), .IN2(g3562), .IN3(n8736), .Q(n12195) );
  OR2X1 U12654 ( .IN1(n5645), .IN2(n418), .Q(n12199) );
  OR3X1 U12655 ( .IN1(n12200), .IN2(n12201), .IN3(n12202), .Q(g30432) );
  AND2X1 U12656 ( .IN1(n11290), .IN2(n3765), .Q(n12202) );
  INVX0 U12657 ( .INP(n12203), .ZN(n11290) );
  AND2X1 U12658 ( .IN1(test_so43), .IN2(n8810), .Q(n12201) );
  AND3X1 U12659 ( .IN1(n12203), .IN2(g3554), .IN3(n8737), .Q(n12200) );
  OR2X1 U12660 ( .IN1(n5645), .IN2(n410), .Q(n12203) );
  OR3X1 U12661 ( .IN1(n12204), .IN2(n12205), .IN3(n12206), .Q(g30431) );
  AND2X1 U12662 ( .IN1(n12207), .IN2(n3765), .Q(n12206) );
  INVX0 U12663 ( .INP(n12208), .ZN(n12207) );
  AND2X1 U12664 ( .IN1(n8835), .IN2(g3598), .Q(n12205) );
  AND3X1 U12665 ( .IN1(n12208), .IN2(g3546), .IN3(n8737), .Q(n12204) );
  OR2X1 U12666 ( .IN1(n5645), .IN2(n412), .Q(n12208) );
  OR3X1 U12667 ( .IN1(n12209), .IN2(n12210), .IN3(n12211), .Q(g30430) );
  AND2X1 U12668 ( .IN1(n3984), .IN2(n12212), .Q(n12211) );
  AND3X1 U12669 ( .IN1(n12213), .IN2(g3610), .IN3(n8737), .Q(n12210) );
  OR2X1 U12670 ( .IN1(n94), .IN2(n417), .Q(n12213) );
  AND2X1 U12671 ( .IN1(n8835), .IN2(g3594), .Q(n12209) );
  OR3X1 U12672 ( .IN1(n12214), .IN2(n12215), .IN3(n12216), .Q(g30429) );
  AND2X1 U12673 ( .IN1(n3984), .IN2(n11293), .Q(n12216) );
  AND3X1 U12674 ( .IN1(n12217), .IN2(g3606), .IN3(n8737), .Q(n12215) );
  OR2X1 U12675 ( .IN1(n94), .IN2(n418), .Q(n12217) );
  AND2X1 U12676 ( .IN1(n8835), .IN2(g3590), .Q(n12214) );
  OR3X1 U12677 ( .IN1(n12218), .IN2(n12219), .IN3(n12220), .Q(g30428) );
  AND2X1 U12678 ( .IN1(n3984), .IN2(n12221), .Q(n12220) );
  AND3X1 U12679 ( .IN1(test_so43), .IN2(n12222), .IN3(n8737), .Q(n12219) );
  OR2X1 U12680 ( .IN1(n94), .IN2(n410), .Q(n12222) );
  AND2X1 U12681 ( .IN1(n8835), .IN2(g3586), .Q(n12218) );
  OR3X1 U12682 ( .IN1(n12223), .IN2(n12224), .IN3(n12225), .Q(g30427) );
  AND2X1 U12683 ( .IN1(n3984), .IN2(n12226), .Q(n12225) );
  AND3X1 U12684 ( .IN1(n12227), .IN2(g3598), .IN3(n8737), .Q(n12224) );
  OR2X1 U12685 ( .IN1(n94), .IN2(n412), .Q(n12227) );
  OR2X1 U12686 ( .IN1(n8308), .IN2(n5576), .Q(n94) );
  AND2X1 U12687 ( .IN1(n8835), .IN2(g3582), .Q(n12223) );
  OR3X1 U12688 ( .IN1(n12228), .IN2(n12229), .IN3(n12230), .Q(g30426) );
  AND2X1 U12689 ( .IN1(n3990), .IN2(n12212), .Q(n12230) );
  AND3X1 U12690 ( .IN1(n12231), .IN2(g3594), .IN3(n8738), .Q(n12229) );
  OR2X1 U12691 ( .IN1(n417), .IN2(n3491), .Q(n12231) );
  AND2X1 U12692 ( .IN1(n8835), .IN2(g3578), .Q(n12228) );
  OR3X1 U12693 ( .IN1(n12232), .IN2(n12233), .IN3(n12234), .Q(g30425) );
  AND2X1 U12694 ( .IN1(n3990), .IN2(n11293), .Q(n12234) );
  AND3X1 U12695 ( .IN1(n12235), .IN2(g3590), .IN3(n8738), .Q(n12233) );
  OR2X1 U12696 ( .IN1(n418), .IN2(n3491), .Q(n12235) );
  AND2X1 U12697 ( .IN1(n8835), .IN2(g3574), .Q(n12232) );
  OR3X1 U12698 ( .IN1(n12236), .IN2(n12237), .IN3(n12238), .Q(g30424) );
  AND2X1 U12699 ( .IN1(n3990), .IN2(n12221), .Q(n12238) );
  AND3X1 U12700 ( .IN1(n12239), .IN2(g3586), .IN3(n8738), .Q(n12237) );
  OR2X1 U12701 ( .IN1(n410), .IN2(n3491), .Q(n12239) );
  AND2X1 U12702 ( .IN1(n8835), .IN2(g3570), .Q(n12236) );
  OR3X1 U12703 ( .IN1(n12240), .IN2(n12241), .IN3(n12242), .Q(g30423) );
  AND2X1 U12704 ( .IN1(n3990), .IN2(n12226), .Q(n12242) );
  AND3X1 U12705 ( .IN1(n12243), .IN2(g3582), .IN3(n8738), .Q(n12241) );
  OR2X1 U12706 ( .IN1(n412), .IN2(n3491), .Q(n12243) );
  OR2X1 U12707 ( .IN1(n8308), .IN2(g3506), .Q(n3491) );
  AND2X1 U12708 ( .IN1(n8835), .IN2(g3566), .Q(n12240) );
  OR3X1 U12709 ( .IN1(n12244), .IN2(n12245), .IN3(n12246), .Q(g30422) );
  AND2X1 U12710 ( .IN1(n3995), .IN2(n12212), .Q(n12246) );
  AND3X1 U12711 ( .IN1(n12247), .IN2(g3578), .IN3(n8738), .Q(n12245) );
  OR2X1 U12712 ( .IN1(n417), .IN2(n3492), .Q(n12247) );
  AND2X1 U12713 ( .IN1(n8836), .IN2(g3558), .Q(n12244) );
  OR3X1 U12714 ( .IN1(n12248), .IN2(n12249), .IN3(n12250), .Q(g30421) );
  AND2X1 U12715 ( .IN1(n3995), .IN2(n11293), .Q(n12250) );
  INVX0 U12716 ( .INP(n418), .ZN(n11293) );
  AND3X1 U12717 ( .IN1(n12251), .IN2(g3574), .IN3(n8738), .Q(n12249) );
  OR2X1 U12718 ( .IN1(n418), .IN2(n3492), .Q(n12251) );
  OR2X1 U12719 ( .IN1(n5569), .IN2(g3522), .Q(n418) );
  AND2X1 U12720 ( .IN1(n8836), .IN2(g3550), .Q(n12248) );
  OR3X1 U12721 ( .IN1(n12252), .IN2(n12253), .IN3(n12254), .Q(g30420) );
  AND2X1 U12722 ( .IN1(n3995), .IN2(n12221), .Q(n12254) );
  INVX0 U12723 ( .INP(n410), .ZN(n12221) );
  AND3X1 U12724 ( .IN1(n12255), .IN2(g3570), .IN3(n8738), .Q(n12253) );
  OR2X1 U12725 ( .IN1(n410), .IN2(n3492), .Q(n12255) );
  OR2X1 U12726 ( .IN1(n5383), .IN2(g3530), .Q(n410) );
  AND2X1 U12727 ( .IN1(n8836), .IN2(g3542), .Q(n12252) );
  OR3X1 U12728 ( .IN1(n12256), .IN2(n12257), .IN3(n12258), .Q(g30419) );
  AND2X1 U12729 ( .IN1(n3995), .IN2(n12226), .Q(n12258) );
  INVX0 U12730 ( .INP(n412), .ZN(n12226) );
  AND3X1 U12731 ( .IN1(n12259), .IN2(g3566), .IN3(n8738), .Q(n12257) );
  OR2X1 U12732 ( .IN1(n412), .IN2(n3492), .Q(n12259) );
  OR2X1 U12733 ( .IN1(n5576), .IN2(g3512), .Q(n3492) );
  OR2X1 U12734 ( .IN1(g3522), .IN2(g3530), .Q(n412) );
  AND2X1 U12735 ( .IN1(n8836), .IN2(g3538), .Q(n12256) );
  OR3X1 U12736 ( .IN1(n12260), .IN2(n12261), .IN3(n12262), .Q(g30418) );
  AND2X1 U12737 ( .IN1(n8836), .IN2(g3562), .Q(n12262) );
  AND2X1 U12738 ( .IN1(n4000), .IN2(n3765), .Q(n12261) );
  AND3X1 U12739 ( .IN1(n8729), .IN2(g3558), .IN3(n12263), .Q(n12260) );
  INVX0 U12740 ( .INP(n4000), .ZN(n12263) );
  OR3X1 U12741 ( .IN1(n12264), .IN2(n12265), .IN3(n12266), .Q(g30417) );
  AND2X1 U12742 ( .IN1(n8836), .IN2(g3554), .Q(n12266) );
  AND2X1 U12743 ( .IN1(n4003), .IN2(n3765), .Q(n12265) );
  AND3X1 U12744 ( .IN1(n8729), .IN2(g3550), .IN3(n12267), .Q(n12264) );
  INVX0 U12745 ( .INP(n4003), .ZN(n12267) );
  OR3X1 U12746 ( .IN1(n12268), .IN2(n12269), .IN3(n12270), .Q(g30416) );
  AND2X1 U12747 ( .IN1(n8836), .IN2(g3546), .Q(n12270) );
  AND2X1 U12748 ( .IN1(n4005), .IN2(n3765), .Q(n12269) );
  AND3X1 U12749 ( .IN1(n8728), .IN2(g3542), .IN3(n12271), .Q(n12268) );
  INVX0 U12750 ( .INP(n4005), .ZN(n12271) );
  OR3X1 U12751 ( .IN1(n12272), .IN2(n12273), .IN3(n12274), .Q(g30415) );
  AND2X1 U12752 ( .IN1(n8836), .IN2(g3530), .Q(n12274) );
  AND2X1 U12753 ( .IN1(n4007), .IN2(n3765), .Q(n12273) );
  AND3X1 U12754 ( .IN1(n8728), .IN2(g3538), .IN3(n12275), .Q(n12272) );
  INVX0 U12755 ( .INP(n4007), .ZN(n12275) );
  AND2X1 U12756 ( .IN1(n11296), .IN2(n5576), .Q(g30414) );
  AND3X1 U12757 ( .IN1(n8728), .IN2(n11289), .IN3(n5645), .Q(n11296) );
  OR3X1 U12758 ( .IN1(n5340), .IN2(g4087), .IN3(n11747), .Q(n11289) );
  OR3X1 U12759 ( .IN1(n12276), .IN2(n12277), .IN3(n12278), .Q(g30413) );
  AND2X1 U12760 ( .IN1(test_so84), .IN2(n8809), .Q(n12278) );
  AND2X1 U12761 ( .IN1(n3765), .IN2(n10567), .Q(n12277) );
  AND2X1 U12762 ( .IN1(n12279), .IN2(g3263), .Q(n12276) );
  OR3X1 U12763 ( .IN1(n12280), .IN2(n12281), .IN3(n12282), .Q(g30412) );
  AND2X1 U12764 ( .IN1(n12283), .IN2(n3765), .Q(n12282) );
  INVX0 U12765 ( .INP(n12284), .ZN(n12283) );
  AND2X1 U12766 ( .IN1(n8836), .IN2(g3255), .Q(n12281) );
  AND3X1 U12767 ( .IN1(n12284), .IN2(g3211), .IN3(n8739), .Q(n12280) );
  OR2X1 U12768 ( .IN1(n5652), .IN2(n510), .Q(n12284) );
  OR3X1 U12769 ( .IN1(n12285), .IN2(n12286), .IN3(n12287), .Q(g30411) );
  AND2X1 U12770 ( .IN1(n11313), .IN2(n3765), .Q(n12287) );
  INVX0 U12771 ( .INP(n12288), .ZN(n11313) );
  AND2X1 U12772 ( .IN1(n8836), .IN2(g3251), .Q(n12286) );
  AND3X1 U12773 ( .IN1(n12288), .IN2(g3203), .IN3(n8739), .Q(n12285) );
  OR2X1 U12774 ( .IN1(n5652), .IN2(n507), .Q(n12288) );
  OR3X1 U12775 ( .IN1(n12289), .IN2(n12290), .IN3(n12291), .Q(g30410) );
  AND2X1 U12776 ( .IN1(n12292), .IN2(n3765), .Q(n12291) );
  INVX0 U12777 ( .INP(n12293), .ZN(n12292) );
  AND2X1 U12778 ( .IN1(n8836), .IN2(g3247), .Q(n12290) );
  AND3X1 U12779 ( .IN1(test_so88), .IN2(n12293), .IN3(n8739), .Q(n12289) );
  OR2X1 U12780 ( .IN1(n5652), .IN2(n508), .Q(n12293) );
  OR3X1 U12781 ( .IN1(n12294), .IN2(n12295), .IN3(n12296), .Q(g30409) );
  AND2X1 U12782 ( .IN1(n4015), .IN2(n12297), .Q(n12296) );
  AND3X1 U12783 ( .IN1(test_so84), .IN2(n12298), .IN3(n8739), .Q(n12295) );
  OR2X1 U12784 ( .IN1(n509), .IN2(n106), .Q(n12298) );
  AND2X1 U12785 ( .IN1(n8836), .IN2(g3243), .Q(n12294) );
  OR3X1 U12786 ( .IN1(n12299), .IN2(n12300), .IN3(n12301), .Q(g30408) );
  AND2X1 U12787 ( .IN1(n4015), .IN2(n11314), .Q(n12301) );
  AND3X1 U12788 ( .IN1(n12302), .IN2(g3255), .IN3(n8739), .Q(n12300) );
  OR2X1 U12789 ( .IN1(n510), .IN2(n106), .Q(n12302) );
  AND2X1 U12790 ( .IN1(n8836), .IN2(g3239), .Q(n12299) );
  OR3X1 U12791 ( .IN1(n12303), .IN2(n12304), .IN3(n12305), .Q(g30407) );
  AND2X1 U12792 ( .IN1(n4015), .IN2(n12306), .Q(n12305) );
  AND3X1 U12793 ( .IN1(n12307), .IN2(g3251), .IN3(n8740), .Q(n12304) );
  OR2X1 U12794 ( .IN1(n507), .IN2(n106), .Q(n12307) );
  AND2X1 U12795 ( .IN1(n8836), .IN2(g3235), .Q(n12303) );
  OR3X1 U12796 ( .IN1(n12308), .IN2(n12309), .IN3(n12310), .Q(g30406) );
  AND2X1 U12797 ( .IN1(n4015), .IN2(n12311), .Q(n12310) );
  AND3X1 U12798 ( .IN1(n12312), .IN2(g3247), .IN3(n8740), .Q(n12309) );
  OR2X1 U12799 ( .IN1(n508), .IN2(n106), .Q(n12312) );
  OR2X1 U12800 ( .IN1(n8315), .IN2(n5366), .Q(n106) );
  AND2X1 U12801 ( .IN1(n8814), .IN2(g3231), .Q(n12308) );
  OR3X1 U12802 ( .IN1(n12313), .IN2(n12314), .IN3(n12315), .Q(g30405) );
  AND2X1 U12803 ( .IN1(n4022), .IN2(n12297), .Q(n12315) );
  AND3X1 U12804 ( .IN1(n12316), .IN2(g3243), .IN3(n8740), .Q(n12314) );
  OR2X1 U12805 ( .IN1(n509), .IN2(n3502), .Q(n12316) );
  AND2X1 U12806 ( .IN1(n8811), .IN2(g3227), .Q(n12313) );
  OR3X1 U12807 ( .IN1(n12317), .IN2(n12318), .IN3(n12319), .Q(g30404) );
  AND2X1 U12808 ( .IN1(n4022), .IN2(n11314), .Q(n12319) );
  AND3X1 U12809 ( .IN1(n12320), .IN2(g3239), .IN3(n8740), .Q(n12318) );
  OR2X1 U12810 ( .IN1(n510), .IN2(n3502), .Q(n12320) );
  AND2X1 U12811 ( .IN1(n8811), .IN2(g3223), .Q(n12317) );
  OR3X1 U12812 ( .IN1(n12321), .IN2(n12322), .IN3(n12323), .Q(g30403) );
  AND2X1 U12813 ( .IN1(n4022), .IN2(n12306), .Q(n12323) );
  AND3X1 U12814 ( .IN1(n12324), .IN2(g3235), .IN3(n8740), .Q(n12322) );
  OR2X1 U12815 ( .IN1(n507), .IN2(n3502), .Q(n12324) );
  AND2X1 U12816 ( .IN1(n8811), .IN2(g3219), .Q(n12321) );
  OR3X1 U12817 ( .IN1(n12325), .IN2(n12326), .IN3(n12327), .Q(g30402) );
  AND2X1 U12818 ( .IN1(n4022), .IN2(n12311), .Q(n12327) );
  AND3X1 U12819 ( .IN1(n12328), .IN2(g3231), .IN3(n8740), .Q(n12326) );
  OR2X1 U12820 ( .IN1(n508), .IN2(n3502), .Q(n12328) );
  OR2X1 U12821 ( .IN1(n8315), .IN2(g3155), .Q(n3502) );
  AND2X1 U12822 ( .IN1(n8811), .IN2(g3215), .Q(n12325) );
  OR3X1 U12823 ( .IN1(n12329), .IN2(n12330), .IN3(n12331), .Q(g30401) );
  AND2X1 U12824 ( .IN1(n4027), .IN2(n12297), .Q(n12331) );
  AND3X1 U12825 ( .IN1(n12332), .IN2(g3227), .IN3(n8740), .Q(n12330) );
  OR2X1 U12826 ( .IN1(n509), .IN2(n3501), .Q(n12332) );
  AND2X1 U12827 ( .IN1(n8811), .IN2(g3207), .Q(n12329) );
  OR3X1 U12828 ( .IN1(n12333), .IN2(n12334), .IN3(n12335), .Q(g30400) );
  AND2X1 U12829 ( .IN1(n4027), .IN2(n11314), .Q(n12335) );
  INVX0 U12830 ( .INP(n510), .ZN(n11314) );
  AND3X1 U12831 ( .IN1(n12336), .IN2(g3223), .IN3(n8740), .Q(n12334) );
  OR2X1 U12832 ( .IN1(n510), .IN2(n3501), .Q(n12336) );
  OR2X1 U12833 ( .IN1(n5390), .IN2(g3171), .Q(n510) );
  AND2X1 U12834 ( .IN1(n8812), .IN2(g3199), .Q(n12333) );
  OR3X1 U12835 ( .IN1(n12337), .IN2(n12338), .IN3(n12339), .Q(g30399) );
  AND2X1 U12836 ( .IN1(n4027), .IN2(n12306), .Q(n12339) );
  INVX0 U12837 ( .INP(n507), .ZN(n12306) );
  AND3X1 U12838 ( .IN1(n12340), .IN2(g3219), .IN3(n8740), .Q(n12338) );
  OR2X1 U12839 ( .IN1(n507), .IN2(n3501), .Q(n12340) );
  OR2X1 U12840 ( .IN1(n5603), .IN2(g3179), .Q(n507) );
  AND2X1 U12841 ( .IN1(n8811), .IN2(g3191), .Q(n12337) );
  OR3X1 U12842 ( .IN1(n12341), .IN2(n12342), .IN3(n12343), .Q(g30398) );
  AND2X1 U12843 ( .IN1(n4027), .IN2(n12311), .Q(n12343) );
  INVX0 U12844 ( .INP(n508), .ZN(n12311) );
  AND3X1 U12845 ( .IN1(n12344), .IN2(g3215), .IN3(n8741), .Q(n12342) );
  OR2X1 U12846 ( .IN1(n508), .IN2(n3501), .Q(n12344) );
  OR2X1 U12847 ( .IN1(n5366), .IN2(g3161), .Q(n3501) );
  OR2X1 U12848 ( .IN1(g3171), .IN2(g3179), .Q(n508) );
  AND2X1 U12849 ( .IN1(n8811), .IN2(g3187), .Q(n12341) );
  OR3X1 U12850 ( .IN1(n12345), .IN2(n12346), .IN3(n12347), .Q(g30397) );
  AND2X1 U12851 ( .IN1(n8811), .IN2(g3211), .Q(n12347) );
  AND2X1 U12852 ( .IN1(n4032), .IN2(n3765), .Q(n12346) );
  AND3X1 U12853 ( .IN1(n8730), .IN2(g3207), .IN3(n12348), .Q(n12345) );
  INVX0 U12854 ( .INP(n4032), .ZN(n12348) );
  OR3X1 U12855 ( .IN1(n12349), .IN2(n12350), .IN3(n12351), .Q(g30396) );
  AND2X1 U12856 ( .IN1(n8811), .IN2(g3203), .Q(n12351) );
  AND2X1 U12857 ( .IN1(n4035), .IN2(n3765), .Q(n12350) );
  AND3X1 U12858 ( .IN1(n8726), .IN2(g3199), .IN3(n12352), .Q(n12349) );
  INVX0 U12859 ( .INP(n4035), .ZN(n12352) );
  OR3X1 U12860 ( .IN1(n12353), .IN2(n12354), .IN3(n12355), .Q(g30395) );
  AND2X1 U12861 ( .IN1(test_so88), .IN2(n8810), .Q(n12355) );
  AND2X1 U12862 ( .IN1(n4037), .IN2(n3765), .Q(n12354) );
  AND3X1 U12863 ( .IN1(n8728), .IN2(g3191), .IN3(n12356), .Q(n12353) );
  INVX0 U12864 ( .INP(n4037), .ZN(n12356) );
  OR3X1 U12865 ( .IN1(n12357), .IN2(n12358), .IN3(n12359), .Q(g30394) );
  AND2X1 U12866 ( .IN1(n8811), .IN2(g3179), .Q(n12359) );
  AND2X1 U12867 ( .IN1(n4039), .IN2(n3765), .Q(n12358) );
  AND3X1 U12868 ( .IN1(n8727), .IN2(g3187), .IN3(n12360), .Q(n12357) );
  INVX0 U12869 ( .INP(n4039), .ZN(n12360) );
  AND3X1 U12870 ( .IN1(n5366), .IN2(n8726), .IN3(n11310), .Q(g30393) );
  AND2X1 U12871 ( .IN1(n11312), .IN2(n5652), .Q(n11310) );
  OR2X1 U12872 ( .IN1(n12004), .IN2(n11747), .Q(n11312) );
  INVX0 U12873 ( .INP(n3799), .ZN(n11747) );
  OR2X1 U12874 ( .IN1(n12361), .IN2(n12362), .Q(g30392) );
  AND2X1 U12875 ( .IN1(n8811), .IN2(g2803), .Q(n12361) );
  OR2X1 U12876 ( .IN1(n12363), .IN2(n12364), .Q(g30391) );
  AND2X1 U12877 ( .IN1(n8812), .IN2(g2771), .Q(n12363) );
  OR2X1 U12878 ( .IN1(n12365), .IN2(n12362), .Q(g30390) );
  AND2X1 U12879 ( .IN1(n12366), .IN2(n8695), .Q(n12362) );
  OR2X1 U12880 ( .IN1(n12367), .IN2(n12368), .Q(n12366) );
  AND2X1 U12881 ( .IN1(n12369), .IN2(n12370), .Q(n12368) );
  AND4X1 U12882 ( .IN1(n12371), .IN2(n12372), .IN3(n12373), .IN4(n12374), .Q(
        n12369) );
  OR2X1 U12883 ( .IN1(n5545), .IN2(n12375), .Q(n12374) );
  OR2X1 U12884 ( .IN1(n5379), .IN2(n1169), .Q(n12373) );
  OR2X1 U12885 ( .IN1(n5609), .IN2(n12376), .Q(n12372) );
  OR2X1 U12886 ( .IN1(n5404), .IN2(n12377), .Q(n12371) );
  AND2X1 U12887 ( .IN1(n12378), .IN2(n12379), .Q(n12367) );
  AND4X1 U12888 ( .IN1(n12380), .IN2(n12381), .IN3(n12382), .IN4(n12383), .Q(
        n12378) );
  OR2X1 U12889 ( .IN1(n12375), .IN2(g2236), .Q(n12383) );
  OR2X1 U12890 ( .IN1(n1169), .IN2(g2370), .Q(n12382) );
  OR2X1 U12891 ( .IN1(n12376), .IN2(g2638), .Q(n12381) );
  OR2X1 U12892 ( .IN1(n12377), .IN2(g2504), .Q(n12380) );
  AND2X1 U12893 ( .IN1(g2834), .IN2(n8810), .Q(n12365) );
  OR2X1 U12894 ( .IN1(n12384), .IN2(n12364), .Q(g30389) );
  AND2X1 U12895 ( .IN1(n12385), .IN2(n8695), .Q(n12364) );
  OR2X1 U12896 ( .IN1(n12386), .IN2(n12387), .Q(n12385) );
  AND2X1 U12897 ( .IN1(n12388), .IN2(n12370), .Q(n12387) );
  AND4X1 U12898 ( .IN1(n12389), .IN2(n12390), .IN3(n12391), .IN4(n12392), .Q(
        n12388) );
  OR2X1 U12899 ( .IN1(n5544), .IN2(n12375), .Q(n12392) );
  OR2X1 U12900 ( .IN1(n5378), .IN2(n1169), .Q(n12391) );
  OR2X1 U12901 ( .IN1(n5610), .IN2(n12376), .Q(n12390) );
  OR2X1 U12902 ( .IN1(n5403), .IN2(n12377), .Q(n12389) );
  AND2X1 U12903 ( .IN1(n12393), .IN2(n12379), .Q(n12386) );
  INVX0 U12904 ( .INP(n12370), .ZN(n12379) );
  AND3X1 U12905 ( .IN1(n3653), .IN2(n9786), .IN3(n5600), .Q(n12370) );
  AND2X1 U12906 ( .IN1(n5349), .IN2(n12394), .Q(n3653) );
  INVX0 U12907 ( .INP(n9081), .ZN(n12394) );
  AND4X1 U12908 ( .IN1(n12395), .IN2(n12396), .IN3(n12397), .IN4(n12398), .Q(
        n12393) );
  OR2X1 U12909 ( .IN1(n12375), .IN2(g1677), .Q(n12398) );
  OR2X1 U12910 ( .IN1(n1169), .IN2(g1811), .Q(n12397) );
  OR2X1 U12911 ( .IN1(n12376), .IN2(g2079), .Q(n12396) );
  OR2X1 U12912 ( .IN1(test_so53), .IN2(n12377), .Q(n12395) );
  AND2X1 U12913 ( .IN1(g2831), .IN2(n8810), .Q(n12384) );
  OR2X1 U12914 ( .IN1(n12399), .IN2(n12400), .Q(g30388) );
  AND2X1 U12915 ( .IN1(n8811), .IN2(g2735), .Q(n12400) );
  AND2X1 U12916 ( .IN1(n12401), .IN2(n3730), .Q(n12399) );
  XOR2X1 U12917 ( .IN1(n3506), .IN2(n5349), .Q(n12401) );
  OR2X1 U12918 ( .IN1(n5600), .IN2(n12402), .Q(n3506) );
  OR3X1 U12919 ( .IN1(n12403), .IN2(n12404), .IN3(n12405), .Q(g30387) );
  AND2X1 U12920 ( .IN1(n12406), .IN2(n9262), .Q(n12405) );
  AND3X1 U12921 ( .IN1(n12407), .IN2(n5457), .IN3(n5777), .Q(n12404) );
  AND2X1 U12922 ( .IN1(n12408), .IN2(g2681), .Q(n12403) );
  OR2X1 U12923 ( .IN1(n8802), .IN2(n12409), .Q(n12408) );
  AND2X1 U12924 ( .IN1(n12410), .IN2(g2675), .Q(n12409) );
  OR2X1 U12925 ( .IN1(n12411), .IN2(n12412), .Q(g30386) );
  AND2X1 U12926 ( .IN1(n12413), .IN2(g2675), .Q(n12412) );
  AND2X1 U12927 ( .IN1(n12406), .IN2(g2681), .Q(n12411) );
  OR3X1 U12928 ( .IN1(n12414), .IN2(n12415), .IN3(n12416), .Q(g30385) );
  AND2X1 U12929 ( .IN1(n8811), .IN2(g2657), .Q(n12416) );
  AND2X1 U12930 ( .IN1(n12407), .IN2(n5418), .Q(n12415) );
  AND2X1 U12931 ( .IN1(n12406), .IN2(g2661), .Q(n12414) );
  INVX0 U12932 ( .INP(n12413), .ZN(n12406) );
  OR2X1 U12933 ( .IN1(n8802), .IN2(n12410), .Q(n12413) );
  OR3X1 U12934 ( .IN1(n12417), .IN2(n12418), .IN3(n12419), .Q(g30384) );
  AND2X1 U12935 ( .IN1(n8811), .IN2(g2652), .Q(n12419) );
  AND2X1 U12936 ( .IN1(n12420), .IN2(g2657), .Q(n12418) );
  OR2X1 U12937 ( .IN1(n12421), .IN2(n11337), .Q(n12420) );
  AND2X1 U12938 ( .IN1(n8718), .IN2(n11348), .Q(n12421) );
  AND3X1 U12939 ( .IN1(n3517), .IN2(n12422), .IN3(n8478), .Q(n12417) );
  XOR2X1 U12940 ( .IN1(n8293), .IN2(n8006), .Q(n12422) );
  OR3X1 U12941 ( .IN1(n12423), .IN2(n12424), .IN3(n12425), .Q(g30383) );
  AND2X1 U12942 ( .IN1(test_so66), .IN2(n8809), .Q(n12425) );
  AND2X1 U12943 ( .IN1(test_so34), .IN2(n12426), .Q(n12424) );
  OR2X1 U12944 ( .IN1(n12427), .IN2(n11337), .Q(n12426) );
  INVX0 U12945 ( .INP(n12428), .ZN(n12427) );
  OR2X1 U12946 ( .IN1(n9987), .IN2(n8793), .Q(n12428) );
  AND3X1 U12947 ( .IN1(n9987), .IN2(n10103), .IN3(n3517), .Q(n12423) );
  OR2X1 U12948 ( .IN1(n5524), .IN2(g2555), .Q(n10103) );
  OR3X1 U12949 ( .IN1(n12429), .IN2(n12430), .IN3(n12431), .Q(g30382) );
  AND2X1 U12950 ( .IN1(n12432), .IN2(n9295), .Q(n12431) );
  AND3X1 U12951 ( .IN1(n12433), .IN2(n5461), .IN3(n5782), .Q(n12430) );
  AND2X1 U12952 ( .IN1(n12434), .IN2(g2547), .Q(n12429) );
  OR2X1 U12953 ( .IN1(n8802), .IN2(n12435), .Q(n12434) );
  AND2X1 U12954 ( .IN1(n12436), .IN2(g2541), .Q(n12435) );
  OR2X1 U12955 ( .IN1(n12437), .IN2(n12438), .Q(g30381) );
  AND2X1 U12956 ( .IN1(n12439), .IN2(g2541), .Q(n12438) );
  AND2X1 U12957 ( .IN1(n12432), .IN2(g2547), .Q(n12437) );
  OR3X1 U12958 ( .IN1(n12440), .IN2(n12441), .IN3(n12442), .Q(g30380) );
  AND2X1 U12959 ( .IN1(n8812), .IN2(g2523), .Q(n12442) );
  AND2X1 U12960 ( .IN1(n12433), .IN2(n5420), .Q(n12441) );
  AND2X1 U12961 ( .IN1(n12432), .IN2(g2527), .Q(n12440) );
  INVX0 U12962 ( .INP(n12439), .ZN(n12432) );
  OR2X1 U12963 ( .IN1(n8803), .IN2(n12436), .Q(n12439) );
  OR3X1 U12964 ( .IN1(n12443), .IN2(n12444), .IN3(n12445), .Q(g30379) );
  AND2X1 U12965 ( .IN1(n8812), .IN2(g2518), .Q(n12445) );
  AND2X1 U12966 ( .IN1(n12446), .IN2(g2523), .Q(n12444) );
  OR2X1 U12967 ( .IN1(n12447), .IN2(n11356), .Q(n12446) );
  AND2X1 U12968 ( .IN1(n8712), .IN2(n11367), .Q(n12447) );
  AND3X1 U12969 ( .IN1(n3536), .IN2(n12448), .IN3(n8485), .Q(n12443) );
  XOR2X1 U12970 ( .IN1(n8295), .IN2(n8003), .Q(n12448) );
  OR3X1 U12971 ( .IN1(n12449), .IN2(n12450), .IN3(n12451), .Q(g30378) );
  AND2X1 U12972 ( .IN1(n8812), .IN2(g2441), .Q(n12451) );
  AND2X1 U12973 ( .IN1(n12452), .IN2(g2461), .Q(n12450) );
  OR2X1 U12974 ( .IN1(n12453), .IN2(n11356), .Q(n12452) );
  INVX0 U12975 ( .INP(n12454), .ZN(n12453) );
  OR2X1 U12976 ( .IN1(n9985), .IN2(n8793), .Q(n12454) );
  AND3X1 U12977 ( .IN1(n9985), .IN2(n10161), .IN3(n3536), .Q(n12449) );
  OR2X1 U12978 ( .IN1(n5523), .IN2(test_so79), .Q(n10161) );
  OR3X1 U12979 ( .IN1(n12455), .IN2(n12456), .IN3(n12457), .Q(g30377) );
  AND2X1 U12980 ( .IN1(n12458), .IN2(n9324), .Q(n12457) );
  AND3X1 U12981 ( .IN1(n12459), .IN2(n5459), .IN3(n8533), .Q(n12456) );
  AND2X1 U12982 ( .IN1(test_so89), .IN2(n12460), .Q(n12455) );
  OR2X1 U12983 ( .IN1(n8803), .IN2(n12461), .Q(n12460) );
  AND2X1 U12984 ( .IN1(n12462), .IN2(g2407), .Q(n12461) );
  OR2X1 U12985 ( .IN1(n12463), .IN2(n12464), .Q(g30376) );
  AND2X1 U12986 ( .IN1(n12465), .IN2(g2407), .Q(n12464) );
  AND2X1 U12987 ( .IN1(test_so89), .IN2(n12458), .Q(n12463) );
  OR3X1 U12988 ( .IN1(n12466), .IN2(n12467), .IN3(n12468), .Q(g30375) );
  AND2X1 U12989 ( .IN1(n8812), .IN2(g2389), .Q(n12468) );
  AND2X1 U12990 ( .IN1(n12459), .IN2(n5421), .Q(n12467) );
  AND2X1 U12991 ( .IN1(n12458), .IN2(g2393), .Q(n12466) );
  INVX0 U12992 ( .INP(n12465), .ZN(n12458) );
  OR2X1 U12993 ( .IN1(n8803), .IN2(n12462), .Q(n12465) );
  OR3X1 U12994 ( .IN1(n12469), .IN2(n12470), .IN3(n12471), .Q(g30374) );
  AND2X1 U12995 ( .IN1(n8812), .IN2(g2384), .Q(n12471) );
  AND2X1 U12996 ( .IN1(n12472), .IN2(g2389), .Q(n12470) );
  OR2X1 U12997 ( .IN1(n12473), .IN2(n11375), .Q(n12472) );
  AND2X1 U12998 ( .IN1(n8712), .IN2(n11386), .Q(n12473) );
  AND3X1 U12999 ( .IN1(n3555), .IN2(n12474), .IN3(n8480), .Q(n12469) );
  XOR2X1 U13000 ( .IN1(n8300), .IN2(n8002), .Q(n12474) );
  OR3X1 U13001 ( .IN1(n12475), .IN2(n12476), .IN3(n12477), .Q(g30373) );
  AND2X1 U13002 ( .IN1(n8812), .IN2(g2307), .Q(n12477) );
  AND2X1 U13003 ( .IN1(n12478), .IN2(g2327), .Q(n12476) );
  OR2X1 U13004 ( .IN1(n12479), .IN2(n11375), .Q(n12478) );
  INVX0 U13005 ( .INP(n12480), .ZN(n12479) );
  OR2X1 U13006 ( .IN1(n9996), .IN2(n8793), .Q(n12480) );
  AND3X1 U13007 ( .IN1(n9996), .IN2(n10217), .IN3(n3555), .Q(n12475) );
  OR2X1 U13008 ( .IN1(n5513), .IN2(g2287), .Q(n10217) );
  OR3X1 U13009 ( .IN1(n12481), .IN2(n12482), .IN3(n12483), .Q(g30372) );
  AND2X1 U13010 ( .IN1(n12484), .IN2(n9273), .Q(n12483) );
  AND3X1 U13011 ( .IN1(n12485), .IN2(n5458), .IN3(n5778), .Q(n12482) );
  AND2X1 U13012 ( .IN1(n12486), .IN2(g2279), .Q(n12481) );
  OR2X1 U13013 ( .IN1(n8804), .IN2(n12487), .Q(n12486) );
  AND2X1 U13014 ( .IN1(n12488), .IN2(g2273), .Q(n12487) );
  OR2X1 U13015 ( .IN1(n12489), .IN2(n12490), .Q(g30371) );
  AND2X1 U13016 ( .IN1(n12491), .IN2(g2273), .Q(n12490) );
  AND2X1 U13017 ( .IN1(n12484), .IN2(g2279), .Q(n12489) );
  OR3X1 U13018 ( .IN1(n12492), .IN2(n12493), .IN3(n12494), .Q(g30370) );
  AND2X1 U13019 ( .IN1(n8812), .IN2(g2255), .Q(n12494) );
  AND2X1 U13020 ( .IN1(n12485), .IN2(n5419), .Q(n12493) );
  AND2X1 U13021 ( .IN1(n12484), .IN2(g2259), .Q(n12492) );
  INVX0 U13022 ( .INP(n12491), .ZN(n12484) );
  OR2X1 U13023 ( .IN1(n8804), .IN2(n12488), .Q(n12491) );
  OR3X1 U13024 ( .IN1(n12495), .IN2(n12496), .IN3(n12497), .Q(g30369) );
  AND2X1 U13025 ( .IN1(n8812), .IN2(g2250), .Q(n12497) );
  AND2X1 U13026 ( .IN1(n12498), .IN2(g2255), .Q(n12496) );
  OR2X1 U13027 ( .IN1(n12499), .IN2(n11394), .Q(n12498) );
  AND2X1 U13028 ( .IN1(n8712), .IN2(n11405), .Q(n12499) );
  AND3X1 U13029 ( .IN1(n3574), .IN2(n12500), .IN3(n8487), .Q(n12495) );
  XOR2X1 U13030 ( .IN1(n8304), .IN2(n8005), .Q(n12500) );
  OR3X1 U13031 ( .IN1(n12501), .IN2(n12502), .IN3(n12503), .Q(g30368) );
  AND2X1 U13032 ( .IN1(n8812), .IN2(g2173), .Q(n12503) );
  AND2X1 U13033 ( .IN1(n12504), .IN2(g2193), .Q(n12502) );
  OR2X1 U13034 ( .IN1(n12505), .IN2(n11394), .Q(n12504) );
  INVX0 U13035 ( .INP(n12506), .ZN(n12505) );
  OR2X1 U13036 ( .IN1(n9982), .IN2(n8793), .Q(n12506) );
  AND3X1 U13037 ( .IN1(n9982), .IN2(n10273), .IN3(n3574), .Q(n12501) );
  OR2X1 U13038 ( .IN1(n5514), .IN2(g2153), .Q(n10273) );
  OR3X1 U13039 ( .IN1(n12507), .IN2(n12508), .IN3(n12509), .Q(g30367) );
  AND2X1 U13040 ( .IN1(n12510), .IN2(g2126), .Q(n12509) );
  AND3X1 U13041 ( .IN1(n12511), .IN2(n5463), .IN3(n5784), .Q(n12508) );
  AND2X1 U13042 ( .IN1(n12512), .IN2(g2122), .Q(n12507) );
  OR2X1 U13043 ( .IN1(n8805), .IN2(n12513), .Q(n12512) );
  AND2X1 U13044 ( .IN1(n12514), .IN2(g2116), .Q(n12513) );
  OR2X1 U13045 ( .IN1(n12515), .IN2(n12516), .Q(g30366) );
  AND2X1 U13046 ( .IN1(n12517), .IN2(g2116), .Q(n12516) );
  AND2X1 U13047 ( .IN1(n12510), .IN2(g2122), .Q(n12515) );
  OR3X1 U13048 ( .IN1(n12518), .IN2(n12519), .IN3(n12520), .Q(g30365) );
  AND2X1 U13049 ( .IN1(n8813), .IN2(g2098), .Q(n12520) );
  AND2X1 U13050 ( .IN1(n12511), .IN2(n5666), .Q(n12519) );
  AND2X1 U13051 ( .IN1(n12510), .IN2(g2102), .Q(n12518) );
  INVX0 U13052 ( .INP(n12517), .ZN(n12510) );
  OR2X1 U13053 ( .IN1(n8805), .IN2(n12514), .Q(n12517) );
  OR3X1 U13054 ( .IN1(n12521), .IN2(n12522), .IN3(n12523), .Q(g30364) );
  AND2X1 U13055 ( .IN1(test_so78), .IN2(n8809), .Q(n12523) );
  AND2X1 U13056 ( .IN1(n12524), .IN2(g2098), .Q(n12522) );
  OR2X1 U13057 ( .IN1(n12525), .IN2(n11413), .Q(n12524) );
  AND2X1 U13058 ( .IN1(n8712), .IN2(n11424), .Q(n12525) );
  AND3X1 U13059 ( .IN1(n8489), .IN2(n3593), .IN3(n12526), .Q(n12521) );
  XOR2X1 U13060 ( .IN1(g2089), .IN2(test_so78), .Q(n12526) );
  OR3X1 U13061 ( .IN1(n12527), .IN2(n12528), .IN3(n12529), .Q(g30363) );
  AND2X1 U13062 ( .IN1(n8813), .IN2(g2016), .Q(n12529) );
  AND2X1 U13063 ( .IN1(test_so59), .IN2(n12530), .Q(n12528) );
  OR2X1 U13064 ( .IN1(n12531), .IN2(n11413), .Q(n12530) );
  INVX0 U13065 ( .INP(n12532), .ZN(n12531) );
  OR2X1 U13066 ( .IN1(n9993), .IN2(n8793), .Q(n12532) );
  AND3X1 U13067 ( .IN1(n9993), .IN2(n10330), .IN3(n3593), .Q(n12527) );
  OR2X1 U13068 ( .IN1(n5505), .IN2(g1996), .Q(n10330) );
  OR3X1 U13069 ( .IN1(n12533), .IN2(n12534), .IN3(n12535), .Q(g30362) );
  AND2X1 U13070 ( .IN1(n12536), .IN2(g1992), .Q(n12535) );
  AND3X1 U13071 ( .IN1(n12537), .IN2(n5462), .IN3(n5783), .Q(n12534) );
  AND2X1 U13072 ( .IN1(n12538), .IN2(g1988), .Q(n12533) );
  OR2X1 U13073 ( .IN1(n8806), .IN2(n12539), .Q(n12538) );
  AND2X1 U13074 ( .IN1(n12540), .IN2(g1982), .Q(n12539) );
  OR2X1 U13075 ( .IN1(n12541), .IN2(n12542), .Q(g30361) );
  AND2X1 U13076 ( .IN1(n12543), .IN2(g1982), .Q(n12542) );
  AND2X1 U13077 ( .IN1(n12536), .IN2(g1988), .Q(n12541) );
  OR3X1 U13078 ( .IN1(n12544), .IN2(n12545), .IN3(n12546), .Q(g30360) );
  AND2X1 U13079 ( .IN1(n8813), .IN2(g1964), .Q(n12546) );
  AND2X1 U13080 ( .IN1(n12537), .IN2(n5664), .Q(n12545) );
  AND2X1 U13081 ( .IN1(n12536), .IN2(g1968), .Q(n12544) );
  INVX0 U13082 ( .INP(n12543), .ZN(n12536) );
  OR2X1 U13083 ( .IN1(n8806), .IN2(n12540), .Q(n12543) );
  OR3X1 U13084 ( .IN1(n12547), .IN2(n12548), .IN3(n12549), .Q(g30359) );
  AND2X1 U13085 ( .IN1(n8813), .IN2(g1959), .Q(n12549) );
  AND2X1 U13086 ( .IN1(n12550), .IN2(g1964), .Q(n12548) );
  OR2X1 U13087 ( .IN1(n12551), .IN2(n11432), .Q(n12550) );
  AND2X1 U13088 ( .IN1(n8713), .IN2(n11444), .Q(n12551) );
  AND3X1 U13089 ( .IN1(n3611), .IN2(n12552), .IN3(n8477), .Q(n12547) );
  XOR2X1 U13090 ( .IN1(n8296), .IN2(n7999), .Q(n12552) );
  OR3X1 U13091 ( .IN1(n12553), .IN2(n12554), .IN3(n12555), .Q(g30358) );
  AND2X1 U13092 ( .IN1(n8813), .IN2(g1882), .Q(n12555) );
  AND2X1 U13093 ( .IN1(n12556), .IN2(g1902), .Q(n12554) );
  OR2X1 U13094 ( .IN1(n12557), .IN2(n11432), .Q(n12556) );
  INVX0 U13095 ( .INP(n12558), .ZN(n12557) );
  OR2X1 U13096 ( .IN1(n9991), .IN2(n8792), .Q(n12558) );
  AND3X1 U13097 ( .IN1(n9991), .IN2(n10388), .IN3(n3611), .Q(n12553) );
  OR2X1 U13098 ( .IN1(n5503), .IN2(test_so8), .Q(n10388) );
  OR3X1 U13099 ( .IN1(n12559), .IN2(n12560), .IN3(n12561), .Q(g30357) );
  AND2X1 U13100 ( .IN1(n12562), .IN2(g1858), .Q(n12561) );
  AND3X1 U13101 ( .IN1(n12563), .IN2(n5464), .IN3(n5785), .Q(n12560) );
  AND2X1 U13102 ( .IN1(n12564), .IN2(g1854), .Q(n12559) );
  OR2X1 U13103 ( .IN1(n8795), .IN2(n12565), .Q(n12564) );
  AND2X1 U13104 ( .IN1(n12566), .IN2(g1848), .Q(n12565) );
  OR2X1 U13105 ( .IN1(n12567), .IN2(n12568), .Q(g30356) );
  AND2X1 U13106 ( .IN1(n12569), .IN2(g1848), .Q(n12568) );
  AND2X1 U13107 ( .IN1(n12562), .IN2(g1854), .Q(n12567) );
  OR3X1 U13108 ( .IN1(n12570), .IN2(n12571), .IN3(n12572), .Q(g30355) );
  AND2X1 U13109 ( .IN1(n8813), .IN2(g1830), .Q(n12572) );
  AND2X1 U13110 ( .IN1(n12563), .IN2(n5665), .Q(n12571) );
  AND2X1 U13111 ( .IN1(n12562), .IN2(g1834), .Q(n12570) );
  INVX0 U13112 ( .INP(n12569), .ZN(n12562) );
  OR2X1 U13113 ( .IN1(n8795), .IN2(n12566), .Q(n12569) );
  OR3X1 U13114 ( .IN1(n12573), .IN2(n12574), .IN3(n12575), .Q(g30354) );
  AND2X1 U13115 ( .IN1(n8813), .IN2(g1825), .Q(n12575) );
  AND2X1 U13116 ( .IN1(n12576), .IN2(g1830), .Q(n12574) );
  OR2X1 U13117 ( .IN1(n12577), .IN2(n11452), .Q(n12576) );
  AND2X1 U13118 ( .IN1(n8713), .IN2(n11463), .Q(n12577) );
  AND3X1 U13119 ( .IN1(n3628), .IN2(n12578), .IN3(n8483), .Q(n12573) );
  XOR2X1 U13120 ( .IN1(n8302), .IN2(n8000), .Q(n12578) );
  OR3X1 U13121 ( .IN1(n12579), .IN2(n12580), .IN3(n12581), .Q(g30353) );
  AND2X1 U13122 ( .IN1(n8813), .IN2(g1748), .Q(n12581) );
  AND2X1 U13123 ( .IN1(n12582), .IN2(g1768), .Q(n12580) );
  OR2X1 U13124 ( .IN1(n12583), .IN2(n11452), .Q(n12582) );
  INVX0 U13125 ( .INP(n12584), .ZN(n12583) );
  OR2X1 U13126 ( .IN1(n9984), .IN2(n8794), .Q(n12584) );
  AND3X1 U13127 ( .IN1(n9984), .IN2(n10444), .IN3(n3628), .Q(n12579) );
  OR2X1 U13128 ( .IN1(n5504), .IN2(g1728), .Q(n10444) );
  OR3X1 U13129 ( .IN1(n12585), .IN2(n12586), .IN3(n12587), .Q(g30352) );
  AND2X1 U13130 ( .IN1(n12588), .IN2(n9236), .Q(n12587) );
  AND4X1 U13131 ( .IN1(n5460), .IN2(n8753), .IN3(n12589), .IN4(n5780), .Q(
        n12586) );
  AND2X1 U13132 ( .IN1(n12590), .IN2(g1720), .Q(n12585) );
  OR2X1 U13133 ( .IN1(n8797), .IN2(n12591), .Q(n12590) );
  AND2X1 U13134 ( .IN1(n12589), .IN2(g1714), .Q(n12591) );
  OR2X1 U13135 ( .IN1(n12592), .IN2(n12593), .Q(g30351) );
  AND2X1 U13136 ( .IN1(n12594), .IN2(g1714), .Q(n12593) );
  AND2X1 U13137 ( .IN1(n12588), .IN2(g1720), .Q(n12592) );
  OR3X1 U13138 ( .IN1(n12595), .IN2(n12596), .IN3(n12597), .Q(g30350) );
  AND2X1 U13139 ( .IN1(n12588), .IN2(g1700), .Q(n12597) );
  INVX0 U13140 ( .INP(n12594), .ZN(n12588) );
  OR2X1 U13141 ( .IN1(n8796), .IN2(n12589), .Q(n12594) );
  AND2X1 U13142 ( .IN1(n8813), .IN2(g1696), .Q(n12596) );
  AND3X1 U13143 ( .IN1(n12589), .IN2(n5417), .IN3(n8741), .Q(n12595) );
  OR3X1 U13144 ( .IN1(n12598), .IN2(n12599), .IN3(n12600), .Q(g30349) );
  AND2X1 U13145 ( .IN1(n8813), .IN2(g1691), .Q(n12600) );
  AND2X1 U13146 ( .IN1(n12601), .IN2(g1696), .Q(n12599) );
  OR2X1 U13147 ( .IN1(n12602), .IN2(n11471), .Q(n12601) );
  AND2X1 U13148 ( .IN1(n8713), .IN2(n11484), .Q(n12602) );
  AND3X1 U13149 ( .IN1(n3646), .IN2(n12603), .IN3(n8488), .Q(n12598) );
  XOR2X1 U13150 ( .IN1(n8298), .IN2(n8004), .Q(n12603) );
  OR3X1 U13151 ( .IN1(n12604), .IN2(n12605), .IN3(n12606), .Q(g30348) );
  AND2X1 U13152 ( .IN1(n8813), .IN2(g1612), .Q(n12606) );
  AND2X1 U13153 ( .IN1(n12607), .IN2(g1632), .Q(n12605) );
  OR2X1 U13154 ( .IN1(n12608), .IN2(n11471), .Q(n12607) );
  INVX0 U13155 ( .INP(n12609), .ZN(n12608) );
  OR2X1 U13156 ( .IN1(g31863), .IN2(n8793), .Q(n12609) );
  AND3X1 U13157 ( .IN1(g31863), .IN2(n12610), .IN3(n3646), .Q(n12604) );
  OR2X1 U13158 ( .IN1(n5549), .IN2(g1592), .Q(n12610) );
  OR2X1 U13159 ( .IN1(n12611), .IN2(n12612), .Q(g30347) );
  INVX0 U13160 ( .INP(n12613), .ZN(n12612) );
  OR2X1 U13161 ( .IN1(n8678), .IN2(n8051), .Q(n12613) );
  AND3X1 U13162 ( .IN1(n12614), .IN2(n12615), .IN3(n12616), .Q(n12611) );
  INVX0 U13163 ( .INP(n12617), .ZN(n12614) );
  AND2X1 U13164 ( .IN1(n12618), .IN2(n12619), .Q(n12617) );
  OR2X1 U13165 ( .IN1(n8797), .IN2(n8461), .Q(n12619) );
  OR2X1 U13166 ( .IN1(n12620), .IN2(n12621), .Q(g30346) );
  AND4X1 U13167 ( .IN1(n12622), .IN2(n12618), .IN3(n12616), .IN4(n8723), .Q(
        n12621) );
  INVX0 U13168 ( .INP(n12623), .ZN(n12616) );
  INVX0 U13169 ( .INP(n12624), .ZN(n12622) );
  AND2X1 U13170 ( .IN1(n12625), .IN2(n8051), .Q(n12624) );
  AND2X1 U13171 ( .IN1(n8813), .IN2(g1536), .Q(n12620) );
  OR2X1 U13172 ( .IN1(n12626), .IN2(n12627), .Q(g30345) );
  AND2X1 U13173 ( .IN1(n12628), .IN2(g1514), .Q(n12627) );
  OR2X1 U13174 ( .IN1(n8797), .IN2(n12629), .Q(n12628) );
  XOR2X1 U13175 ( .IN1(n8490), .IN2(n5302), .Q(n12629) );
  AND2X1 U13176 ( .IN1(n12630), .IN2(n8694), .Q(n12626) );
  OR2X1 U13177 ( .IN1(n10848), .IN2(n12623), .Q(n12630) );
  AND2X1 U13178 ( .IN1(n12631), .IN2(n8694), .Q(g30344) );
  OR2X1 U13179 ( .IN1(n12623), .IN2(n12632), .Q(n12631) );
  XOR2X1 U13180 ( .IN1(n5364), .IN2(n5302), .Q(n12632) );
  OR2X1 U13181 ( .IN1(n12633), .IN2(n4173), .Q(n12623) );
  AND2X1 U13182 ( .IN1(n4172), .IN2(n10848), .Q(n12633) );
  INVX0 U13183 ( .INP(n12634), .ZN(n10848) );
  AND3X1 U13184 ( .IN1(n12635), .IN2(g7946), .IN3(n4895), .Q(n4172) );
  OR3X1 U13185 ( .IN1(n12636), .IN2(n12637), .IN3(n12638), .Q(g30343) );
  AND2X1 U13186 ( .IN1(n4175), .IN2(n11488), .Q(n12638) );
  AND3X1 U13187 ( .IN1(n9103), .IN2(g1361), .IN3(n8742), .Q(n12637) );
  OR2X1 U13188 ( .IN1(n12639), .IN2(n12640), .Q(n9103) );
  AND2X1 U13189 ( .IN1(n8469), .IN2(n11068), .Q(n12639) );
  AND2X1 U13190 ( .IN1(n8813), .IN2(g1345), .Q(n12636) );
  OR3X1 U13191 ( .IN1(n12641), .IN2(n12642), .IN3(n12643), .Q(g30342) );
  AND2X1 U13192 ( .IN1(n8813), .IN2(g1256), .Q(n12643) );
  AND2X1 U13193 ( .IN1(n3736), .IN2(n5553), .Q(n12642) );
  AND3X1 U13194 ( .IN1(n11076), .IN2(n12644), .IN3(g1259), .Q(n12641) );
  INVX0 U13195 ( .INP(n3736), .ZN(n12644) );
  OR2X1 U13196 ( .IN1(n12645), .IN2(n12646), .Q(g30341) );
  INVX0 U13197 ( .INP(n12647), .ZN(n12646) );
  OR2X1 U13198 ( .IN1(n8678), .IN2(n8052), .Q(n12647) );
  AND3X1 U13199 ( .IN1(n12648), .IN2(n12649), .IN3(n12650), .Q(n12645) );
  INVX0 U13200 ( .INP(n12651), .ZN(n12648) );
  AND2X1 U13201 ( .IN1(n12652), .IN2(n12653), .Q(n12651) );
  OR2X1 U13202 ( .IN1(n8798), .IN2(n8462), .Q(n12653) );
  OR2X1 U13203 ( .IN1(n12654), .IN2(n12655), .Q(g30340) );
  AND4X1 U13204 ( .IN1(n12656), .IN2(n12652), .IN3(n12650), .IN4(n8722), .Q(
        n12655) );
  INVX0 U13205 ( .INP(n12657), .ZN(n12650) );
  INVX0 U13206 ( .INP(n12658), .ZN(n12656) );
  AND2X1 U13207 ( .IN1(n12659), .IN2(n8052), .Q(n12658) );
  AND2X1 U13208 ( .IN1(n8813), .IN2(g1193), .Q(n12654) );
  OR2X1 U13209 ( .IN1(n12660), .IN2(n12661), .Q(g30339) );
  AND2X1 U13210 ( .IN1(n12662), .IN2(g1171), .Q(n12661) );
  OR2X1 U13211 ( .IN1(n8798), .IN2(n12663), .Q(n12662) );
  XOR2X1 U13212 ( .IN1(n5599), .IN2(n5304), .Q(n12663) );
  AND2X1 U13213 ( .IN1(n12664), .IN2(n8694), .Q(n12660) );
  OR2X1 U13214 ( .IN1(n11021), .IN2(n12657), .Q(n12664) );
  AND2X1 U13215 ( .IN1(n12665), .IN2(n8693), .Q(g30338) );
  OR2X1 U13216 ( .IN1(n12657), .IN2(n12666), .Q(n12665) );
  XOR2X1 U13217 ( .IN1(n5363), .IN2(n5304), .Q(n12666) );
  OR2X1 U13218 ( .IN1(n12667), .IN2(n4191), .Q(n12657) );
  AND2X1 U13219 ( .IN1(n4190), .IN2(n11021), .Q(n12667) );
  INVX0 U13220 ( .INP(n12668), .ZN(n11021) );
  AND3X1 U13221 ( .IN1(n12669), .IN2(g7916), .IN3(n4920), .Q(n4190) );
  OR3X1 U13222 ( .IN1(n12670), .IN2(n12671), .IN3(n12672), .Q(g30337) );
  AND2X1 U13223 ( .IN1(n4193), .IN2(n11499), .Q(n12672) );
  AND3X1 U13224 ( .IN1(n9006), .IN2(g1018), .IN3(n8742), .Q(n12671) );
  OR2X1 U13225 ( .IN1(n12673), .IN2(n12674), .Q(n9006) );
  AND2X1 U13226 ( .IN1(n8466), .IN2(n11083), .Q(n12673) );
  AND2X1 U13227 ( .IN1(n8813), .IN2(g1002), .Q(n12670) );
  OR3X1 U13228 ( .IN1(n12675), .IN2(n12676), .IN3(n12677), .Q(g30336) );
  AND2X1 U13229 ( .IN1(n8813), .IN2(g911), .Q(n12677) );
  AND2X1 U13230 ( .IN1(n3741), .IN2(n5560), .Q(n12676) );
  AND3X1 U13231 ( .IN1(n11091), .IN2(n12678), .IN3(g914), .Q(n12675) );
  INVX0 U13232 ( .INP(n3741), .ZN(n12678) );
  OR3X1 U13233 ( .IN1(n12679), .IN2(n12680), .IN3(n12681), .Q(g30335) );
  AND2X1 U13234 ( .IN1(test_so60), .IN2(n8810), .Q(n12681) );
  AND2X1 U13235 ( .IN1(n3743), .IN2(n5470), .Q(n12680) );
  AND3X1 U13236 ( .IN1(n2404), .IN2(n12682), .IN3(g744), .Q(n12679) );
  INVX0 U13237 ( .INP(n3743), .ZN(n12682) );
  AND3X1 U13238 ( .IN1(n4198), .IN2(test_so60), .IN3(n12683), .Q(n3743) );
  INVX0 U13239 ( .INP(n12684), .ZN(n12683) );
  OR2X1 U13240 ( .IN1(n5482), .IN2(g736), .Q(n4198) );
  OR3X1 U13241 ( .IN1(n12685), .IN2(n12686), .IN3(n12687), .Q(g30334) );
  AND2X1 U13242 ( .IN1(n8814), .IN2(g586), .Q(n12687) );
  AND2X1 U13243 ( .IN1(n3745), .IN2(n5294), .Q(n12686) );
  AND3X1 U13244 ( .IN1(n2421), .IN2(n12688), .IN3(g577), .Q(n12685) );
  INVX0 U13245 ( .INP(n3745), .ZN(n12688) );
  OR2X1 U13246 ( .IN1(n12689), .IN2(n12690), .Q(g30333) );
  AND2X1 U13247 ( .IN1(n8814), .IN2(g142), .Q(n12690) );
  AND2X1 U13248 ( .IN1(n9969), .IN2(n12691), .Q(n12689) );
  XOR2X1 U13249 ( .IN1(test_so73), .IN2(n11635), .Q(n12691) );
  AND2X1 U13250 ( .IN1(n8713), .IN2(n11636), .Q(n9969) );
  AND3X1 U13251 ( .IN1(g691), .IN2(n12692), .IN3(n12693), .Q(n11636) );
  INVX0 U13252 ( .INP(n12694), .ZN(n12693) );
  AND2X1 U13253 ( .IN1(n11635), .IN2(n12695), .Q(n12694) );
  OR3X1 U13254 ( .IN1(test_so72), .IN2(g174), .IN3(g168), .Q(n12695) );
  OR3X1 U13255 ( .IN1(n12696), .IN2(n12697), .IN3(n12698), .Q(g29309) );
  AND2X1 U13256 ( .IN1(n3765), .IN2(n12699), .Q(n12698) );
  OR2X1 U13257 ( .IN1(n10569), .IN2(n5739), .Q(n12699) );
  AND3X1 U13258 ( .IN1(n9107), .IN2(g6541), .IN3(n11664), .Q(n12697) );
  OR3X1 U13259 ( .IN1(n12700), .IN2(n12701), .IN3(n12702), .Q(g29308) );
  AND2X1 U13260 ( .IN1(n8814), .IN2(g6523), .Q(n12702) );
  AND2X1 U13261 ( .IN1(n5659), .IN2(n12703), .Q(n12701) );
  AND2X1 U13262 ( .IN1(n12704), .IN2(g6527), .Q(n12700) );
  OR3X1 U13263 ( .IN1(n12705), .IN2(n12706), .IN3(n12707), .Q(g29307) );
  AND2X1 U13264 ( .IN1(n12704), .IN2(g6523), .Q(n12707) );
  AND3X1 U13265 ( .IN1(n5426), .IN2(n12703), .IN3(n5806), .Q(n12706) );
  AND2X1 U13266 ( .IN1(n12708), .IN2(g6519), .Q(n12705) );
  OR2X1 U13267 ( .IN1(n8799), .IN2(n12709), .Q(n12708) );
  AND2X1 U13268 ( .IN1(n12710), .IN2(g6513), .Q(n12709) );
  OR2X1 U13269 ( .IN1(n12711), .IN2(n12712), .Q(g29306) );
  AND2X1 U13270 ( .IN1(n12713), .IN2(g6513), .Q(n12712) );
  AND2X1 U13271 ( .IN1(n12704), .IN2(g6519), .Q(n12711) );
  INVX0 U13272 ( .INP(n12713), .ZN(n12704) );
  OR2X1 U13273 ( .IN1(n8799), .IN2(n12710), .Q(n12713) );
  OR3X1 U13274 ( .IN1(n12714), .IN2(n12715), .IN3(n12716), .Q(g29305) );
  INVX0 U13275 ( .INP(n12717), .ZN(n12716) );
  OR2X1 U13276 ( .IN1(n11643), .IN2(n12710), .Q(n12717) );
  OR2X1 U13277 ( .IN1(n8407), .IN2(n8793), .Q(n11643) );
  AND3X1 U13278 ( .IN1(n12703), .IN2(g6505), .IN3(n5748), .Q(n12715) );
  AND2X1 U13279 ( .IN1(n8713), .IN2(n12710), .Q(n12703) );
  AND2X1 U13280 ( .IN1(n12718), .IN2(g6500), .Q(n12714) );
  OR2X1 U13281 ( .IN1(n8800), .IN2(n12719), .Q(n12718) );
  AND2X1 U13282 ( .IN1(n8365), .IN2(n12710), .Q(n12719) );
  AND2X1 U13283 ( .IN1(n10594), .IN2(n12720), .Q(n12710) );
  OR2X1 U13284 ( .IN1(n12721), .IN2(n12722), .Q(g29304) );
  AND2X1 U13285 ( .IN1(n12723), .IN2(n8693), .Q(n12722) );
  OR2X1 U13286 ( .IN1(n12724), .IN2(n12725), .Q(n12723) );
  AND2X1 U13287 ( .IN1(n12726), .IN2(n10594), .Q(n12725) );
  XNOR2X1 U13288 ( .IN1(n12727), .IN2(n12728), .Q(n12726) );
  OR2X1 U13289 ( .IN1(n5748), .IN2(n12720), .Q(n12728) );
  AND3X1 U13290 ( .IN1(g17722), .IN2(g6727), .IN3(n9003), .Q(n12720) );
  AND2X1 U13291 ( .IN1(n8479), .IN2(g6500), .Q(n12724) );
  AND2X1 U13292 ( .IN1(n8814), .IN2(g6505), .Q(n12721) );
  OR3X1 U13293 ( .IN1(n12696), .IN2(n12729), .IN3(n12730), .Q(g29303) );
  AND2X1 U13294 ( .IN1(n3765), .IN2(n12731), .Q(n12730) );
  OR2X1 U13295 ( .IN1(n10581), .IN2(n5741), .Q(n12731) );
  AND3X1 U13296 ( .IN1(n9107), .IN2(g6195), .IN3(n11751), .Q(n12729) );
  OR3X1 U13297 ( .IN1(n12732), .IN2(n12733), .IN3(n12734), .Q(g29302) );
  AND2X1 U13298 ( .IN1(n8814), .IN2(g6177), .Q(n12734) );
  AND2X1 U13299 ( .IN1(n5667), .IN2(n12735), .Q(n12733) );
  AND2X1 U13300 ( .IN1(n12736), .IN2(g6181), .Q(n12732) );
  OR3X1 U13301 ( .IN1(n12737), .IN2(n12738), .IN3(n12739), .Q(g29301) );
  AND2X1 U13302 ( .IN1(n12736), .IN2(g6177), .Q(n12739) );
  AND3X1 U13303 ( .IN1(n5430), .IN2(n12735), .IN3(n5810), .Q(n12738) );
  AND2X1 U13304 ( .IN1(n12740), .IN2(g6173), .Q(n12737) );
  OR2X1 U13305 ( .IN1(n8800), .IN2(n12741), .Q(n12740) );
  AND2X1 U13306 ( .IN1(n12742), .IN2(g6167), .Q(n12741) );
  OR2X1 U13307 ( .IN1(n12743), .IN2(n12744), .Q(g29300) );
  AND2X1 U13308 ( .IN1(n12745), .IN2(g6167), .Q(n12744) );
  AND2X1 U13309 ( .IN1(n12736), .IN2(g6173), .Q(n12743) );
  INVX0 U13310 ( .INP(n12745), .ZN(n12736) );
  OR2X1 U13311 ( .IN1(n8800), .IN2(n12742), .Q(n12745) );
  OR3X1 U13312 ( .IN1(n12746), .IN2(n12747), .IN3(n12748), .Q(g29299) );
  INVX0 U13313 ( .INP(n12749), .ZN(n12748) );
  OR2X1 U13314 ( .IN1(n11654), .IN2(n12742), .Q(n12749) );
  OR2X1 U13315 ( .IN1(n8451), .IN2(n8794), .Q(n11654) );
  AND3X1 U13316 ( .IN1(n12735), .IN2(g6159), .IN3(n5747), .Q(n12747) );
  AND2X1 U13317 ( .IN1(n8713), .IN2(n12742), .Q(n12735) );
  AND2X1 U13318 ( .IN1(n12750), .IN2(g6154), .Q(n12746) );
  OR2X1 U13319 ( .IN1(n8800), .IN2(n12751), .Q(n12750) );
  AND2X1 U13320 ( .IN1(n8366), .IN2(n12742), .Q(n12751) );
  AND2X1 U13321 ( .IN1(n10609), .IN2(n12752), .Q(n12742) );
  OR2X1 U13322 ( .IN1(n12753), .IN2(n12754), .Q(g29298) );
  AND2X1 U13323 ( .IN1(n12755), .IN2(n8693), .Q(n12754) );
  OR2X1 U13324 ( .IN1(n12756), .IN2(n12757), .Q(n12755) );
  AND2X1 U13325 ( .IN1(n12758), .IN2(n10609), .Q(n12757) );
  XNOR2X1 U13326 ( .IN1(n12759), .IN2(n12760), .Q(n12758) );
  OR2X1 U13327 ( .IN1(n5747), .IN2(n12752), .Q(n12760) );
  AND3X1 U13328 ( .IN1(g17685), .IN2(n9821), .IN3(test_so69), .Q(n12752) );
  AND2X1 U13329 ( .IN1(n10613), .IN2(g6154), .Q(n12756) );
  AND2X1 U13330 ( .IN1(n8814), .IN2(g6159), .Q(n12753) );
  OR3X1 U13331 ( .IN1(n12696), .IN2(n12761), .IN3(n12762), .Q(g29297) );
  AND2X1 U13332 ( .IN1(n3765), .IN2(n12763), .Q(n12762) );
  OR2X1 U13333 ( .IN1(n10580), .IN2(n5736), .Q(n12763) );
  AND3X1 U13334 ( .IN1(n9107), .IN2(g5849), .IN3(n11837), .Q(n12761) );
  OR3X1 U13335 ( .IN1(n12764), .IN2(n12765), .IN3(n12766), .Q(g29296) );
  AND2X1 U13336 ( .IN1(n8814), .IN2(g5831), .Q(n12766) );
  AND2X1 U13337 ( .IN1(n5663), .IN2(n12767), .Q(n12765) );
  AND2X1 U13338 ( .IN1(n12768), .IN2(g5835), .Q(n12764) );
  OR3X1 U13339 ( .IN1(n12769), .IN2(n12770), .IN3(n12771), .Q(g29295) );
  AND2X1 U13340 ( .IN1(n12768), .IN2(g5831), .Q(n12771) );
  AND3X1 U13341 ( .IN1(n5429), .IN2(n12767), .IN3(n5809), .Q(n12770) );
  AND2X1 U13342 ( .IN1(n12772), .IN2(g5827), .Q(n12769) );
  OR2X1 U13343 ( .IN1(n8801), .IN2(n12773), .Q(n12772) );
  AND2X1 U13344 ( .IN1(n12774), .IN2(g5821), .Q(n12773) );
  OR2X1 U13345 ( .IN1(n12775), .IN2(n12776), .Q(g29294) );
  AND2X1 U13346 ( .IN1(n12777), .IN2(g5821), .Q(n12776) );
  AND2X1 U13347 ( .IN1(n12768), .IN2(g5827), .Q(n12775) );
  INVX0 U13348 ( .INP(n12777), .ZN(n12768) );
  OR2X1 U13349 ( .IN1(n8801), .IN2(n12774), .Q(n12777) );
  OR3X1 U13350 ( .IN1(n12778), .IN2(n12779), .IN3(n12780), .Q(g29293) );
  INVX0 U13351 ( .INP(n12781), .ZN(n12780) );
  OR2X1 U13352 ( .IN1(n11655), .IN2(n12774), .Q(n12781) );
  OR2X1 U13353 ( .IN1(n8452), .IN2(n8794), .Q(n11655) );
  AND3X1 U13354 ( .IN1(n12767), .IN2(g5813), .IN3(n5749), .Q(n12779) );
  AND2X1 U13355 ( .IN1(n8713), .IN2(n12774), .Q(n12767) );
  AND2X1 U13356 ( .IN1(n12782), .IN2(g5808), .Q(n12778) );
  OR2X1 U13357 ( .IN1(n8801), .IN2(n12783), .Q(n12782) );
  AND2X1 U13358 ( .IN1(n8364), .IN2(n12774), .Q(n12783) );
  AND2X1 U13359 ( .IN1(n10626), .IN2(n12784), .Q(n12774) );
  OR2X1 U13360 ( .IN1(n12785), .IN2(n12786), .Q(g29292) );
  AND2X1 U13361 ( .IN1(n12787), .IN2(n8693), .Q(n12786) );
  OR2X1 U13362 ( .IN1(n12788), .IN2(n12789), .Q(n12787) );
  AND2X1 U13363 ( .IN1(n12790), .IN2(n10626), .Q(n12789) );
  XNOR2X1 U13364 ( .IN1(n12791), .IN2(n12792), .Q(n12790) );
  OR2X1 U13365 ( .IN1(n5749), .IN2(n12784), .Q(n12792) );
  AND3X1 U13366 ( .IN1(g17646), .IN2(g6035), .IN3(n9834), .Q(n12784) );
  AND2X1 U13367 ( .IN1(n10630), .IN2(g5808), .Q(n12788) );
  AND2X1 U13368 ( .IN1(n8814), .IN2(g5813), .Q(n12785) );
  OR3X1 U13369 ( .IN1(n12696), .IN2(n12793), .IN3(n12794), .Q(g29291) );
  AND2X1 U13370 ( .IN1(n3765), .IN2(n12795), .Q(n12794) );
  OR2X1 U13371 ( .IN1(n10577), .IN2(n5737), .Q(n12795) );
  AND3X1 U13372 ( .IN1(n9107), .IN2(g5503), .IN3(n11922), .Q(n12793) );
  OR3X1 U13373 ( .IN1(n12796), .IN2(n12797), .IN3(n12798), .Q(g29290) );
  AND2X1 U13374 ( .IN1(n8814), .IN2(g5485), .Q(n12798) );
  AND2X1 U13375 ( .IN1(n5660), .IN2(n12799), .Q(n12797) );
  AND2X1 U13376 ( .IN1(n12800), .IN2(g5489), .Q(n12796) );
  OR3X1 U13377 ( .IN1(n12801), .IN2(n12802), .IN3(n12803), .Q(g29289) );
  AND2X1 U13378 ( .IN1(n12800), .IN2(g5485), .Q(n12803) );
  AND3X1 U13379 ( .IN1(n5425), .IN2(n12799), .IN3(n5805), .Q(n12802) );
  AND2X1 U13380 ( .IN1(n12804), .IN2(g5481), .Q(n12801) );
  OR2X1 U13381 ( .IN1(n8801), .IN2(n12805), .Q(n12804) );
  AND2X1 U13382 ( .IN1(n12806), .IN2(g5475), .Q(n12805) );
  OR2X1 U13383 ( .IN1(n12807), .IN2(n12808), .Q(g29288) );
  AND2X1 U13384 ( .IN1(n12809), .IN2(g5475), .Q(n12808) );
  AND2X1 U13385 ( .IN1(n12800), .IN2(g5481), .Q(n12807) );
  INVX0 U13386 ( .INP(n12809), .ZN(n12800) );
  OR2X1 U13387 ( .IN1(n8801), .IN2(n12806), .Q(n12809) );
  OR3X1 U13388 ( .IN1(n12810), .IN2(n12811), .IN3(n12812), .Q(g29287) );
  INVX0 U13389 ( .INP(n12813), .ZN(n12812) );
  OR2X1 U13390 ( .IN1(n11653), .IN2(n12806), .Q(n12813) );
  OR2X1 U13391 ( .IN1(n8450), .IN2(n8794), .Q(n11653) );
  AND3X1 U13392 ( .IN1(n12799), .IN2(g5467), .IN3(n5744), .Q(n12811) );
  AND2X1 U13393 ( .IN1(n8713), .IN2(n12806), .Q(n12799) );
  AND2X1 U13394 ( .IN1(n12814), .IN2(g5462), .Q(n12810) );
  OR2X1 U13395 ( .IN1(n8800), .IN2(n12815), .Q(n12814) );
  AND2X1 U13396 ( .IN1(n8395), .IN2(n12806), .Q(n12815) );
  AND2X1 U13397 ( .IN1(n10642), .IN2(n12816), .Q(n12806) );
  OR2X1 U13398 ( .IN1(n12817), .IN2(n12818), .Q(g29286) );
  AND2X1 U13399 ( .IN1(n12819), .IN2(n8693), .Q(n12818) );
  OR2X1 U13400 ( .IN1(n12820), .IN2(n12821), .Q(n12819) );
  AND2X1 U13401 ( .IN1(n12822), .IN2(n10642), .Q(n12821) );
  XNOR2X1 U13402 ( .IN1(n12823), .IN2(n12824), .Q(n12822) );
  OR2X1 U13403 ( .IN1(n5744), .IN2(n12816), .Q(n12824) );
  AND3X1 U13404 ( .IN1(g17604), .IN2(g5689), .IN3(n9826), .Q(n12816) );
  AND2X1 U13405 ( .IN1(n10646), .IN2(g5462), .Q(n12820) );
  AND2X1 U13406 ( .IN1(n8814), .IN2(g5467), .Q(n12817) );
  OR3X1 U13407 ( .IN1(n12696), .IN2(n12825), .IN3(n12826), .Q(g29285) );
  AND2X1 U13408 ( .IN1(n3765), .IN2(n12827), .Q(n12826) );
  OR2X1 U13409 ( .IN1(g32975), .IN2(n5734), .Q(n12827) );
  AND3X1 U13410 ( .IN1(n9107), .IN2(g5156), .IN3(n9099), .Q(n12825) );
  OR3X1 U13411 ( .IN1(n12828), .IN2(n12829), .IN3(n12830), .Q(g29284) );
  AND2X1 U13412 ( .IN1(n8814), .IN2(g5138), .Q(n12830) );
  AND2X1 U13413 ( .IN1(n12831), .IN2(n5658), .Q(n12829) );
  AND2X1 U13414 ( .IN1(n12832), .IN2(g5142), .Q(n12828) );
  OR3X1 U13415 ( .IN1(n12833), .IN2(n12834), .IN3(n12835), .Q(g29283) );
  AND2X1 U13416 ( .IN1(n12832), .IN2(g5138), .Q(n12835) );
  AND3X1 U13417 ( .IN1(n12831), .IN2(n8516), .IN3(n5807), .Q(n12834) );
  AND2X1 U13418 ( .IN1(n12836), .IN2(g5134), .Q(n12833) );
  OR2X1 U13419 ( .IN1(n8799), .IN2(n12837), .Q(n12836) );
  AND2X1 U13420 ( .IN1(test_so96), .IN2(n12838), .Q(n12837) );
  OR2X1 U13421 ( .IN1(n12839), .IN2(n12840), .Q(g29282) );
  AND2X1 U13422 ( .IN1(test_so96), .IN2(n12841), .Q(n12840) );
  AND2X1 U13423 ( .IN1(n12832), .IN2(g5134), .Q(n12839) );
  INVX0 U13424 ( .INP(n12841), .ZN(n12832) );
  OR2X1 U13425 ( .IN1(n8799), .IN2(n12838), .Q(n12841) );
  OR3X1 U13426 ( .IN1(n12842), .IN2(n12843), .IN3(n12844), .Q(g29281) );
  INVX0 U13427 ( .INP(n12845), .ZN(n12844) );
  OR2X1 U13428 ( .IN1(n11650), .IN2(n12838), .Q(n12845) );
  OR2X1 U13429 ( .IN1(n8457), .IN2(n8794), .Q(n11650) );
  AND3X1 U13430 ( .IN1(n12831), .IN2(g5120), .IN3(n5743), .Q(n12843) );
  AND2X1 U13431 ( .IN1(n8713), .IN2(n12838), .Q(n12831) );
  AND2X1 U13432 ( .IN1(n12846), .IN2(g5115), .Q(n12842) );
  OR2X1 U13433 ( .IN1(n8798), .IN2(n12847), .Q(n12846) );
  AND2X1 U13434 ( .IN1(n8396), .IN2(n12838), .Q(n12847) );
  AND2X1 U13435 ( .IN1(g33959), .IN2(n12848), .Q(n12838) );
  OR2X1 U13436 ( .IN1(n12849), .IN2(n12850), .Q(g29280) );
  AND2X1 U13437 ( .IN1(n12851), .IN2(n8693), .Q(n12850) );
  OR2X1 U13438 ( .IN1(n12852), .IN2(n12853), .Q(n12851) );
  AND2X1 U13439 ( .IN1(n12854), .IN2(g33959), .Q(n12853) );
  XNOR2X1 U13440 ( .IN1(n12855), .IN2(n12856), .Q(n12854) );
  OR2X1 U13441 ( .IN1(n5743), .IN2(n12848), .Q(n12856) );
  AND3X1 U13442 ( .IN1(g17577), .IN2(g31860), .IN3(test_so10), .Q(n12848) );
  AND2X1 U13443 ( .IN1(n8474), .IN2(g5115), .Q(n12852) );
  AND2X1 U13444 ( .IN1(n8814), .IN2(g5120), .Q(n12849) );
  OR2X1 U13445 ( .IN1(n12857), .IN2(g29279), .Q(g29278) );
  AND2X1 U13446 ( .IN1(n8814), .IN2(g4572), .Q(n12857) );
  OR2X1 U13447 ( .IN1(n12858), .IN2(g29277), .Q(g29276) );
  AND2X1 U13448 ( .IN1(test_so100), .IN2(n8809), .Q(n12858) );
  OR2X1 U13449 ( .IN1(n12859), .IN2(n12860), .Q(g29275) );
  AND2X1 U13450 ( .IN1(test_so11), .IN2(n8809), .Q(n12860) );
  AND2X1 U13451 ( .IN1(n12861), .IN2(n12105), .Q(n12859) );
  XOR2X1 U13452 ( .IN1(n12106), .IN2(g4087), .Q(n12861) );
  INVX0 U13453 ( .INP(n11598), .ZN(n12106) );
  OR2X1 U13454 ( .IN1(n12862), .IN2(n8491), .Q(n11598) );
  OR3X1 U13455 ( .IN1(n12696), .IN2(n12863), .IN3(n12864), .Q(g29274) );
  AND2X1 U13456 ( .IN1(n3765), .IN2(n12865), .Q(n12864) );
  OR2X1 U13457 ( .IN1(n9012), .IN2(n5735), .Q(n12865) );
  AND3X1 U13458 ( .IN1(n9107), .IN2(g3849), .IN3(n9011), .Q(n12863) );
  OR3X1 U13459 ( .IN1(n12866), .IN2(n12867), .IN3(n12868), .Q(g29273) );
  AND2X1 U13460 ( .IN1(n8812), .IN2(g3831), .Q(n12868) );
  AND2X1 U13461 ( .IN1(n12869), .IN2(n5662), .Q(n12867) );
  AND2X1 U13462 ( .IN1(n12870), .IN2(g3835), .Q(n12866) );
  OR3X1 U13463 ( .IN1(n12871), .IN2(n12872), .IN3(n12873), .Q(g29272) );
  AND2X1 U13464 ( .IN1(n12870), .IN2(g3831), .Q(n12873) );
  AND3X1 U13465 ( .IN1(n5428), .IN2(n12869), .IN3(n5808), .Q(n12872) );
  AND2X1 U13466 ( .IN1(n12874), .IN2(g3827), .Q(n12871) );
  OR2X1 U13467 ( .IN1(n8795), .IN2(n12875), .Q(n12874) );
  AND2X1 U13468 ( .IN1(n12876), .IN2(g3821), .Q(n12875) );
  OR2X1 U13469 ( .IN1(n12877), .IN2(n12878), .Q(g29271) );
  AND2X1 U13470 ( .IN1(n12879), .IN2(g3821), .Q(n12878) );
  AND2X1 U13471 ( .IN1(n12870), .IN2(g3827), .Q(n12877) );
  INVX0 U13472 ( .INP(n12879), .ZN(n12870) );
  OR2X1 U13473 ( .IN1(n8797), .IN2(n12876), .Q(n12879) );
  OR3X1 U13474 ( .IN1(n12880), .IN2(n12881), .IN3(n12882), .Q(g29270) );
  INVX0 U13475 ( .INP(n12883), .ZN(n12882) );
  OR2X1 U13476 ( .IN1(n9482), .IN2(n12876), .Q(n12883) );
  OR2X1 U13477 ( .IN1(n8429), .IN2(n8794), .Q(n9482) );
  AND3X1 U13478 ( .IN1(n12869), .IN2(g3813), .IN3(n5745), .Q(n12881) );
  AND2X1 U13479 ( .IN1(n8713), .IN2(n12876), .Q(n12869) );
  AND2X1 U13480 ( .IN1(n12884), .IN2(g3808), .Q(n12880) );
  OR2X1 U13481 ( .IN1(n8795), .IN2(n12885), .Q(n12884) );
  AND2X1 U13482 ( .IN1(n8394), .IN2(n12876), .Q(n12885) );
  AND2X1 U13483 ( .IN1(n10681), .IN2(n12886), .Q(n12876) );
  OR2X1 U13484 ( .IN1(n12887), .IN2(n12888), .Q(g29269) );
  AND2X1 U13485 ( .IN1(n12889), .IN2(n8693), .Q(n12888) );
  OR2X1 U13486 ( .IN1(n12890), .IN2(n12891), .Q(n12889) );
  AND2X1 U13487 ( .IN1(n12892), .IN2(n10681), .Q(n12891) );
  XNOR2X1 U13488 ( .IN1(n12893), .IN2(n12894), .Q(n12892) );
  OR2X1 U13489 ( .IN1(n5745), .IN2(n12886), .Q(n12894) );
  AND3X1 U13490 ( .IN1(g16693), .IN2(g4040), .IN3(n9820), .Q(n12886) );
  AND2X1 U13491 ( .IN1(n10685), .IN2(g3808), .Q(n12890) );
  AND2X1 U13492 ( .IN1(n8814), .IN2(g3813), .Q(n12887) );
  OR3X1 U13493 ( .IN1(n12696), .IN2(n12895), .IN3(n12896), .Q(g29268) );
  AND2X1 U13494 ( .IN1(n3765), .IN2(n12897), .Q(n12896) );
  OR2X1 U13495 ( .IN1(n10572), .IN2(n5740), .Q(n12897) );
  AND3X1 U13496 ( .IN1(n9107), .IN2(g3498), .IN3(n12194), .Q(n12895) );
  OR3X1 U13497 ( .IN1(n12898), .IN2(n12899), .IN3(n12900), .Q(g29267) );
  AND2X1 U13498 ( .IN1(n8814), .IN2(g3480), .Q(n12900) );
  AND2X1 U13499 ( .IN1(n5668), .IN2(n12901), .Q(n12899) );
  AND2X1 U13500 ( .IN1(n12902), .IN2(g3484), .Q(n12898) );
  OR3X1 U13501 ( .IN1(n12903), .IN2(n12904), .IN3(n12905), .Q(g29266) );
  AND2X1 U13502 ( .IN1(n12902), .IN2(g3480), .Q(n12905) );
  AND3X1 U13503 ( .IN1(n5424), .IN2(n12901), .IN3(n5786), .Q(n12904) );
  AND2X1 U13504 ( .IN1(n12906), .IN2(g3476), .Q(n12903) );
  OR2X1 U13505 ( .IN1(n8800), .IN2(n12907), .Q(n12906) );
  AND2X1 U13506 ( .IN1(n12908), .IN2(g3470), .Q(n12907) );
  OR2X1 U13507 ( .IN1(n12909), .IN2(n12910), .Q(g29265) );
  AND2X1 U13508 ( .IN1(n12911), .IN2(g3470), .Q(n12910) );
  AND2X1 U13509 ( .IN1(n12902), .IN2(g3476), .Q(n12909) );
  INVX0 U13510 ( .INP(n12911), .ZN(n12902) );
  OR2X1 U13511 ( .IN1(n8799), .IN2(n12908), .Q(n12911) );
  OR3X1 U13512 ( .IN1(n12912), .IN2(n12913), .IN3(n12914), .Q(g29264) );
  INVX0 U13513 ( .INP(n12915), .ZN(n12914) );
  OR2X1 U13514 ( .IN1(n11658), .IN2(n12908), .Q(n12915) );
  OR2X1 U13515 ( .IN1(n8430), .IN2(n8793), .Q(n11658) );
  AND3X1 U13516 ( .IN1(n12901), .IN2(g3462), .IN3(n8508), .Q(n12913) );
  AND2X1 U13517 ( .IN1(n8714), .IN2(n12908), .Q(n12901) );
  AND2X1 U13518 ( .IN1(test_so4), .IN2(n12916), .Q(n12912) );
  OR2X1 U13519 ( .IN1(n8798), .IN2(n12917), .Q(n12916) );
  AND2X1 U13520 ( .IN1(n8393), .IN2(n12908), .Q(n12917) );
  AND2X1 U13521 ( .IN1(n10697), .IN2(n12918), .Q(n12908) );
  OR2X1 U13522 ( .IN1(n12919), .IN2(n12920), .Q(g29263) );
  AND2X1 U13523 ( .IN1(n12921), .IN2(n8693), .Q(n12920) );
  OR2X1 U13524 ( .IN1(n12922), .IN2(n12923), .Q(n12921) );
  AND2X1 U13525 ( .IN1(n12924), .IN2(n10697), .Q(n12923) );
  XNOR2X1 U13526 ( .IN1(n12925), .IN2(n12926), .Q(n12924) );
  OR2X1 U13527 ( .IN1(n8508), .IN2(n12918), .Q(n12926) );
  AND3X1 U13528 ( .IN1(g16656), .IN2(g3689), .IN3(n9833), .Q(n12918) );
  AND2X1 U13529 ( .IN1(test_so4), .IN2(n10701), .Q(n12922) );
  AND2X1 U13530 ( .IN1(n8813), .IN2(g3462), .Q(n12919) );
  OR3X1 U13531 ( .IN1(n12696), .IN2(n12927), .IN3(n12928), .Q(g29262) );
  AND2X1 U13532 ( .IN1(n3765), .IN2(n12929), .Q(n12928) );
  OR2X1 U13533 ( .IN1(n10567), .IN2(n5738), .Q(n12929) );
  AND3X1 U13534 ( .IN1(n9107), .IN2(g3147), .IN3(n12279), .Q(n12927) );
  AND2X1 U13535 ( .IN1(n9107), .IN2(n3765), .Q(n12696) );
  AND2X1 U13536 ( .IN1(g4180), .IN2(n8034), .Q(n9107) );
  OR3X1 U13537 ( .IN1(n12930), .IN2(n12931), .IN3(n12932), .Q(g29261) );
  AND2X1 U13538 ( .IN1(n8813), .IN2(g3129), .Q(n12932) );
  AND2X1 U13539 ( .IN1(n5661), .IN2(n12933), .Q(n12931) );
  AND2X1 U13540 ( .IN1(n12934), .IN2(g3133), .Q(n12930) );
  OR3X1 U13541 ( .IN1(n12935), .IN2(n12936), .IN3(n12937), .Q(g29260) );
  AND2X1 U13542 ( .IN1(n12934), .IN2(g3129), .Q(n12937) );
  AND3X1 U13543 ( .IN1(n5423), .IN2(n12933), .IN3(n5781), .Q(n12936) );
  AND2X1 U13544 ( .IN1(n12938), .IN2(g3125), .Q(n12935) );
  OR2X1 U13545 ( .IN1(n8795), .IN2(n12939), .Q(n12938) );
  AND2X1 U13546 ( .IN1(n12940), .IN2(g3119), .Q(n12939) );
  OR2X1 U13547 ( .IN1(n12941), .IN2(n12942), .Q(g29259) );
  AND2X1 U13548 ( .IN1(n12943), .IN2(g3119), .Q(n12942) );
  AND2X1 U13549 ( .IN1(n12934), .IN2(g3125), .Q(n12941) );
  INVX0 U13550 ( .INP(n12943), .ZN(n12934) );
  OR2X1 U13551 ( .IN1(n8796), .IN2(n12940), .Q(n12943) );
  OR3X1 U13552 ( .IN1(n12944), .IN2(n12945), .IN3(n12946), .Q(g29258) );
  INVX0 U13553 ( .INP(n12947), .ZN(n12946) );
  OR2X1 U13554 ( .IN1(n11659), .IN2(n12940), .Q(n12947) );
  OR2X1 U13555 ( .IN1(n8408), .IN2(n8793), .Q(n11659) );
  AND3X1 U13556 ( .IN1(n12933), .IN2(g3111), .IN3(n5742), .Q(n12945) );
  AND2X1 U13557 ( .IN1(n8714), .IN2(n12940), .Q(n12933) );
  AND2X1 U13558 ( .IN1(n12948), .IN2(g3106), .Q(n12944) );
  OR2X1 U13559 ( .IN1(n8806), .IN2(n12949), .Q(n12948) );
  AND2X1 U13560 ( .IN1(n8397), .IN2(n12940), .Q(n12949) );
  AND2X1 U13561 ( .IN1(n10715), .IN2(n12950), .Q(n12940) );
  OR2X1 U13562 ( .IN1(n12951), .IN2(n12952), .Q(g29257) );
  AND2X1 U13563 ( .IN1(n12953), .IN2(n8692), .Q(n12952) );
  OR2X1 U13564 ( .IN1(n12954), .IN2(n12955), .Q(n12953) );
  AND2X1 U13565 ( .IN1(n12956), .IN2(n10715), .Q(n12955) );
  XNOR2X1 U13566 ( .IN1(n12957), .IN2(n12958), .Q(n12956) );
  OR2X1 U13567 ( .IN1(n5742), .IN2(n12950), .Q(n12958) );
  AND3X1 U13568 ( .IN1(g16624), .IN2(g3338), .IN3(n9825), .Q(n12950) );
  AND2X1 U13569 ( .IN1(n10713), .IN2(g3106), .Q(n12954) );
  AND2X1 U13570 ( .IN1(n8813), .IN2(g3111), .Q(n12951) );
  OR4X1 U13571 ( .IN1(n2787), .IN2(n12959), .IN3(n12960), .IN4(n12961), .Q(
        g29256) );
  AND2X1 U13572 ( .IN1(n8813), .IN2(g2729), .Q(n12961) );
  AND3X1 U13573 ( .IN1(n12402), .IN2(g2735), .IN3(n8743), .Q(n12960) );
  AND2X1 U13574 ( .IN1(n5600), .IN2(n12962), .Q(n12959) );
  INVX0 U13575 ( .INP(n12402), .ZN(n12962) );
  OR2X1 U13576 ( .IN1(n12376), .IN2(n9767), .Q(n12402) );
  OR2X1 U13577 ( .IN1(n5301), .IN2(n8347), .Q(n9767) );
  OR2X1 U13578 ( .IN1(n12963), .IN2(n12964), .Q(g29255) );
  AND2X1 U13579 ( .IN1(n12965), .IN2(g2652), .Q(n12964) );
  OR2X1 U13580 ( .IN1(n12966), .IN2(n11337), .Q(n12965) );
  AND2X1 U13581 ( .IN1(n4379), .IN2(n8692), .Q(n12966) );
  AND2X1 U13582 ( .IN1(n12967), .IN2(g2638), .Q(n12963) );
  OR2X1 U13583 ( .IN1(n8805), .IN2(n12968), .Q(n12967) );
  AND2X1 U13584 ( .IN1(n11334), .IN2(n9022), .Q(n12968) );
  OR2X1 U13585 ( .IN1(n8478), .IN2(n8293), .Q(n9022) );
  OR4X1 U13586 ( .IN1(n12969), .IN2(n12970), .IN3(n12971), .IN4(n12972), .Q(
        g29254) );
  AND2X1 U13587 ( .IN1(n3517), .IN2(n12973), .Q(n12972) );
  OR4X1 U13588 ( .IN1(n12974), .IN2(n12975), .IN3(n12976), .IN4(n12977), .Q(
        n12973) );
  AND2X1 U13589 ( .IN1(n8442), .IN2(n12978), .Q(n12977) );
  OR2X1 U13590 ( .IN1(n12979), .IN2(n12980), .Q(n12978) );
  AND2X1 U13591 ( .IN1(g2619), .IN2(g2571), .Q(n12980) );
  AND2X1 U13592 ( .IN1(test_so61), .IN2(g2587), .Q(n12979) );
  AND3X1 U13593 ( .IN1(n5508), .IN2(n5372), .IN3(test_so66), .Q(n12976) );
  AND2X1 U13594 ( .IN1(n8478), .IN2(g2563), .Q(n12975) );
  INVX0 U13595 ( .INP(n11348), .ZN(n8478) );
  OR2X1 U13596 ( .IN1(n8442), .IN2(g2587), .Q(n11348) );
  AND2X1 U13597 ( .IN1(n9987), .IN2(g2583), .Q(n12974) );
  AND2X1 U13598 ( .IN1(g2610), .IN2(n5508), .Q(n9987) );
  AND2X1 U13599 ( .IN1(n8714), .IN2(n11334), .Q(n3517) );
  AND2X1 U13600 ( .IN1(n12407), .IN2(g2567), .Q(n12971) );
  AND2X1 U13601 ( .IN1(n8714), .IN2(n12410), .Q(n12407) );
  AND3X1 U13602 ( .IN1(g2619), .IN2(g2587), .IN3(n11334), .Q(n12410) );
  INVX0 U13603 ( .INP(n12981), .ZN(n11334) );
  AND2X1 U13604 ( .IN1(n8813), .IN2(g2619), .Q(n12970) );
  AND2X1 U13605 ( .IN1(n11337), .IN2(g2638), .Q(n12969) );
  AND2X1 U13606 ( .IN1(n8714), .IN2(n12981), .Q(n11337) );
  OR3X1 U13607 ( .IN1(n12982), .IN2(n12983), .IN3(n12376), .Q(n12981) );
  AND2X1 U13608 ( .IN1(n9786), .IN2(g2819), .Q(n12983) );
  OR2X1 U13609 ( .IN1(n12984), .IN2(n12985), .Q(g29253) );
  AND2X1 U13610 ( .IN1(n12986), .IN2(g2518), .Q(n12985) );
  OR2X1 U13611 ( .IN1(n12987), .IN2(n11356), .Q(n12986) );
  AND2X1 U13612 ( .IN1(n4391), .IN2(n8692), .Q(n12987) );
  AND2X1 U13613 ( .IN1(n12988), .IN2(g2504), .Q(n12984) );
  OR2X1 U13614 ( .IN1(n8803), .IN2(n12989), .Q(n12988) );
  AND2X1 U13615 ( .IN1(n11353), .IN2(n9021), .Q(n12989) );
  OR2X1 U13616 ( .IN1(n8485), .IN2(n8295), .Q(n9021) );
  OR4X1 U13617 ( .IN1(n12990), .IN2(n12991), .IN3(n12992), .IN4(n12993), .Q(
        g29252) );
  AND2X1 U13618 ( .IN1(n3536), .IN2(n12994), .Q(n12993) );
  OR4X1 U13619 ( .IN1(n12995), .IN2(n12996), .IN3(n12997), .IN4(n12998), .Q(
        n12994) );
  AND2X1 U13620 ( .IN1(n8443), .IN2(n12999), .Q(n12998) );
  OR2X1 U13621 ( .IN1(n13000), .IN2(n13001), .Q(n12999) );
  AND2X1 U13622 ( .IN1(g2485), .IN2(g2437), .Q(n13001) );
  AND2X1 U13623 ( .IN1(g2453), .IN2(n9274), .Q(n13000) );
  AND3X1 U13624 ( .IN1(n5373), .IN2(g2441), .IN3(n5509), .Q(n12997) );
  AND2X1 U13625 ( .IN1(n8485), .IN2(g2429), .Q(n12996) );
  INVX0 U13626 ( .INP(n11367), .ZN(n8485) );
  OR2X1 U13627 ( .IN1(n8443), .IN2(g2453), .Q(n11367) );
  AND2X1 U13628 ( .IN1(n9985), .IN2(g2449), .Q(n12995) );
  AND2X1 U13629 ( .IN1(g2476), .IN2(n5509), .Q(n9985) );
  AND2X1 U13630 ( .IN1(n8714), .IN2(n11353), .Q(n3536) );
  AND2X1 U13631 ( .IN1(n12433), .IN2(g2433), .Q(n12992) );
  AND2X1 U13632 ( .IN1(n8714), .IN2(n12436), .Q(n12433) );
  AND3X1 U13633 ( .IN1(g2485), .IN2(g2453), .IN3(n11353), .Q(n12436) );
  INVX0 U13634 ( .INP(n13002), .ZN(n11353) );
  AND2X1 U13635 ( .IN1(n8812), .IN2(g2485), .Q(n12991) );
  AND2X1 U13636 ( .IN1(n11356), .IN2(g2504), .Q(n12990) );
  AND2X1 U13637 ( .IN1(n8714), .IN2(n13002), .Q(n11356) );
  OR3X1 U13638 ( .IN1(n12982), .IN2(n13003), .IN3(n12377), .Q(n13002) );
  AND2X1 U13639 ( .IN1(n9786), .IN2(g2815), .Q(n13003) );
  OR2X1 U13640 ( .IN1(n13004), .IN2(n13005), .Q(g29251) );
  AND2X1 U13641 ( .IN1(n13006), .IN2(g2370), .Q(n13005) );
  OR2X1 U13642 ( .IN1(n8803), .IN2(n13007), .Q(n13006) );
  AND2X1 U13643 ( .IN1(n11372), .IN2(n9020), .Q(n13007) );
  OR2X1 U13644 ( .IN1(n8480), .IN2(n8300), .Q(n9020) );
  AND2X1 U13645 ( .IN1(n13008), .IN2(g2384), .Q(n13004) );
  OR2X1 U13646 ( .IN1(n13009), .IN2(n11375), .Q(n13008) );
  AND2X1 U13647 ( .IN1(n4402), .IN2(n8692), .Q(n13009) );
  OR4X1 U13648 ( .IN1(n13010), .IN2(n13011), .IN3(n13012), .IN4(n13013), .Q(
        g29250) );
  AND2X1 U13649 ( .IN1(n3555), .IN2(n13014), .Q(n13013) );
  OR4X1 U13650 ( .IN1(n13015), .IN2(n13016), .IN3(n13017), .IN4(n13018), .Q(
        n13014) );
  AND2X1 U13651 ( .IN1(n13019), .IN2(n8498), .Q(n13018) );
  OR2X1 U13652 ( .IN1(n13020), .IN2(n13021), .Q(n13019) );
  AND2X1 U13653 ( .IN1(g2351), .IN2(g2303), .Q(n13021) );
  AND2X1 U13654 ( .IN1(g2319), .IN2(n9314), .Q(n13020) );
  AND3X1 U13655 ( .IN1(n5375), .IN2(g2307), .IN3(n5511), .Q(n13017) );
  AND2X1 U13656 ( .IN1(n8480), .IN2(g2295), .Q(n13016) );
  INVX0 U13657 ( .INP(n11386), .ZN(n8480) );
  OR2X1 U13658 ( .IN1(g2319), .IN2(n8498), .Q(n11386) );
  AND2X1 U13659 ( .IN1(n9996), .IN2(g2315), .Q(n13015) );
  AND2X1 U13660 ( .IN1(test_so21), .IN2(n5511), .Q(n9996) );
  AND2X1 U13661 ( .IN1(n8714), .IN2(n11372), .Q(n3555) );
  AND2X1 U13662 ( .IN1(n12459), .IN2(g2299), .Q(n13012) );
  AND2X1 U13663 ( .IN1(n8714), .IN2(n12462), .Q(n12459) );
  AND3X1 U13664 ( .IN1(g2351), .IN2(g2319), .IN3(n11372), .Q(n12462) );
  INVX0 U13665 ( .INP(n13022), .ZN(n11372) );
  AND2X1 U13666 ( .IN1(n8812), .IN2(g2351), .Q(n13011) );
  AND2X1 U13667 ( .IN1(n11375), .IN2(g2370), .Q(n13010) );
  AND2X1 U13668 ( .IN1(n8715), .IN2(n13022), .Q(n11375) );
  OR3X1 U13669 ( .IN1(n1169), .IN2(n12982), .IN3(n13023), .Q(n13022) );
  AND2X1 U13670 ( .IN1(n9786), .IN2(g2807), .Q(n13023) );
  OR2X1 U13671 ( .IN1(n13024), .IN2(n13025), .Q(g29249) );
  AND2X1 U13672 ( .IN1(n13026), .IN2(g2236), .Q(n13025) );
  OR2X1 U13673 ( .IN1(n8803), .IN2(n13027), .Q(n13026) );
  AND2X1 U13674 ( .IN1(n11391), .IN2(n9019), .Q(n13027) );
  OR2X1 U13675 ( .IN1(n8487), .IN2(n8304), .Q(n9019) );
  AND2X1 U13676 ( .IN1(n13028), .IN2(g2250), .Q(n13024) );
  OR2X1 U13677 ( .IN1(n13029), .IN2(n11394), .Q(n13028) );
  AND2X1 U13678 ( .IN1(n4414), .IN2(n8691), .Q(n13029) );
  OR4X1 U13679 ( .IN1(n13030), .IN2(n13031), .IN3(n13032), .IN4(n13033), .Q(
        g29248) );
  AND2X1 U13680 ( .IN1(n3574), .IN2(n13034), .Q(n13033) );
  OR4X1 U13681 ( .IN1(n13035), .IN2(n13036), .IN3(n13037), .IN4(n13038), .Q(
        n13034) );
  AND2X1 U13682 ( .IN1(n8391), .IN2(n13039), .Q(n13038) );
  OR2X1 U13683 ( .IN1(n13040), .IN2(n13041), .Q(n13039) );
  AND2X1 U13684 ( .IN1(g2217), .IN2(g2169), .Q(n13041) );
  AND2X1 U13685 ( .IN1(g2185), .IN2(n9352), .Q(n13040) );
  AND3X1 U13686 ( .IN1(n5376), .IN2(g2173), .IN3(n5512), .Q(n13037) );
  AND2X1 U13687 ( .IN1(n8487), .IN2(g2161), .Q(n13036) );
  INVX0 U13688 ( .INP(n11405), .ZN(n8487) );
  OR2X1 U13689 ( .IN1(n8391), .IN2(g2185), .Q(n11405) );
  AND2X1 U13690 ( .IN1(n9982), .IN2(g2181), .Q(n13035) );
  AND2X1 U13691 ( .IN1(g2208), .IN2(n5512), .Q(n9982) );
  AND2X1 U13692 ( .IN1(n8715), .IN2(n11391), .Q(n3574) );
  AND2X1 U13693 ( .IN1(n12485), .IN2(g2165), .Q(n13032) );
  AND2X1 U13694 ( .IN1(n8715), .IN2(n12488), .Q(n12485) );
  AND3X1 U13695 ( .IN1(g2217), .IN2(g2185), .IN3(n11391), .Q(n12488) );
  INVX0 U13696 ( .INP(n13042), .ZN(n11391) );
  AND2X1 U13697 ( .IN1(n8812), .IN2(g2217), .Q(n13031) );
  AND2X1 U13698 ( .IN1(n11394), .IN2(g2236), .Q(n13030) );
  AND2X1 U13699 ( .IN1(n8715), .IN2(n13042), .Q(n11394) );
  OR2X1 U13700 ( .IN1(n13043), .IN2(n13044), .Q(n13042) );
  AND2X1 U13701 ( .IN1(n9786), .IN2(g2803), .Q(n13043) );
  OR2X1 U13702 ( .IN1(n13045), .IN2(n13046), .Q(g29247) );
  AND2X1 U13703 ( .IN1(test_so78), .IN2(n13047), .Q(n13046) );
  OR2X1 U13704 ( .IN1(n13048), .IN2(n11413), .Q(n13047) );
  AND2X1 U13705 ( .IN1(n4425), .IN2(n8691), .Q(n13048) );
  AND2X1 U13706 ( .IN1(n13049), .IN2(g2079), .Q(n13045) );
  OR2X1 U13707 ( .IN1(n8802), .IN2(n13050), .Q(n13049) );
  AND2X1 U13708 ( .IN1(n11410), .IN2(n9018), .Q(n13050) );
  OR2X1 U13709 ( .IN1(n8489), .IN2(n8514), .Q(n9018) );
  OR4X1 U13710 ( .IN1(n13051), .IN2(n13052), .IN3(n13053), .IN4(n13054), .Q(
        g29246) );
  AND2X1 U13711 ( .IN1(n3593), .IN2(n13055), .Q(n13054) );
  OR4X1 U13712 ( .IN1(n13056), .IN2(n13057), .IN3(n13058), .IN4(n13059), .Q(
        n13055) );
  AND2X1 U13713 ( .IN1(n8448), .IN2(n13060), .Q(n13059) );
  OR2X1 U13714 ( .IN1(n13061), .IN2(n13062), .Q(n13060) );
  AND2X1 U13715 ( .IN1(g2060), .IN2(g2012), .Q(n13062) );
  AND2X1 U13716 ( .IN1(g2028), .IN2(n9312), .Q(n13061) );
  AND3X1 U13717 ( .IN1(n5371), .IN2(g2016), .IN3(n5507), .Q(n13058) );
  AND2X1 U13718 ( .IN1(n8489), .IN2(g2004), .Q(n13057) );
  INVX0 U13719 ( .INP(n11424), .ZN(n8489) );
  OR2X1 U13720 ( .IN1(n8448), .IN2(g2028), .Q(n11424) );
  AND2X1 U13721 ( .IN1(n9993), .IN2(g2024), .Q(n13056) );
  AND2X1 U13722 ( .IN1(g2051), .IN2(n5507), .Q(n9993) );
  AND2X1 U13723 ( .IN1(n8715), .IN2(n11410), .Q(n3593) );
  AND2X1 U13724 ( .IN1(n12511), .IN2(g2008), .Q(n13053) );
  AND2X1 U13725 ( .IN1(n8715), .IN2(n12514), .Q(n12511) );
  AND3X1 U13726 ( .IN1(g2060), .IN2(g2028), .IN3(n11410), .Q(n12514) );
  INVX0 U13727 ( .INP(n13063), .ZN(n11410) );
  AND2X1 U13728 ( .IN1(n8812), .IN2(g2060), .Q(n13052) );
  AND2X1 U13729 ( .IN1(n11413), .IN2(g2079), .Q(n13051) );
  AND2X1 U13730 ( .IN1(n8715), .IN2(n13063), .Q(n11413) );
  OR3X1 U13731 ( .IN1(n12982), .IN2(n13064), .IN3(n12376), .Q(n13063) );
  AND2X1 U13732 ( .IN1(n9786), .IN2(g2787), .Q(n13064) );
  OR2X1 U13733 ( .IN1(n13065), .IN2(n13066), .Q(g29245) );
  AND2X1 U13734 ( .IN1(test_so53), .IN2(n13067), .Q(n13066) );
  OR2X1 U13735 ( .IN1(n8802), .IN2(n13068), .Q(n13067) );
  AND2X1 U13736 ( .IN1(n11429), .IN2(n9017), .Q(n13068) );
  OR2X1 U13737 ( .IN1(n8477), .IN2(n8296), .Q(n9017) );
  AND2X1 U13738 ( .IN1(n13069), .IN2(g1959), .Q(n13065) );
  OR2X1 U13739 ( .IN1(n13070), .IN2(n11432), .Q(n13069) );
  AND2X1 U13740 ( .IN1(n4436), .IN2(n8691), .Q(n13070) );
  OR4X1 U13741 ( .IN1(n13071), .IN2(n13072), .IN3(n13073), .IN4(n13074), .Q(
        g29244) );
  AND2X1 U13742 ( .IN1(n3611), .IN2(n13075), .Q(n13074) );
  OR4X1 U13743 ( .IN1(n13076), .IN2(n13077), .IN3(n13078), .IN4(n13079), .Q(
        n13075) );
  AND2X1 U13744 ( .IN1(n8449), .IN2(n13080), .Q(n13079) );
  OR2X1 U13745 ( .IN1(n13081), .IN2(n13082), .Q(n13080) );
  AND2X1 U13746 ( .IN1(g1926), .IN2(g1878), .Q(n13082) );
  AND2X1 U13747 ( .IN1(g1894), .IN2(n9280), .Q(n13081) );
  AND3X1 U13748 ( .IN1(n5374), .IN2(g1882), .IN3(n5510), .Q(n13078) );
  AND2X1 U13749 ( .IN1(n8477), .IN2(g1870), .Q(n13077) );
  INVX0 U13750 ( .INP(n11444), .ZN(n8477) );
  OR2X1 U13751 ( .IN1(n8449), .IN2(g1894), .Q(n11444) );
  AND2X1 U13752 ( .IN1(n9991), .IN2(g1890), .Q(n13076) );
  AND2X1 U13753 ( .IN1(g1917), .IN2(n5510), .Q(n9991) );
  AND2X1 U13754 ( .IN1(n8715), .IN2(n11429), .Q(n3611) );
  AND2X1 U13755 ( .IN1(n12537), .IN2(g1874), .Q(n13073) );
  AND2X1 U13756 ( .IN1(n8715), .IN2(n12540), .Q(n12537) );
  AND3X1 U13757 ( .IN1(g1926), .IN2(g1894), .IN3(n11429), .Q(n12540) );
  INVX0 U13758 ( .INP(n13083), .ZN(n11429) );
  AND2X1 U13759 ( .IN1(n8811), .IN2(g1926), .Q(n13072) );
  AND2X1 U13760 ( .IN1(n11432), .IN2(test_so53), .Q(n13071) );
  AND2X1 U13761 ( .IN1(n8715), .IN2(n13083), .Q(n11432) );
  OR3X1 U13762 ( .IN1(n12982), .IN2(n13084), .IN3(n12377), .Q(n13083) );
  INVX0 U13763 ( .INP(n13085), .ZN(n12377) );
  AND2X1 U13764 ( .IN1(n9786), .IN2(g2783), .Q(n13084) );
  OR2X1 U13765 ( .IN1(n13086), .IN2(n13087), .Q(g29243) );
  AND2X1 U13766 ( .IN1(n13088), .IN2(g1811), .Q(n13087) );
  OR2X1 U13767 ( .IN1(n8802), .IN2(n13089), .Q(n13088) );
  AND2X1 U13768 ( .IN1(n11449), .IN2(n9016), .Q(n13089) );
  OR2X1 U13769 ( .IN1(n8483), .IN2(n8302), .Q(n9016) );
  AND2X1 U13770 ( .IN1(n13090), .IN2(g1825), .Q(n13086) );
  OR2X1 U13771 ( .IN1(n13091), .IN2(n11452), .Q(n13090) );
  AND2X1 U13772 ( .IN1(n4447), .IN2(n8691), .Q(n13091) );
  OR4X1 U13773 ( .IN1(n13092), .IN2(n13093), .IN3(n13094), .IN4(n13095), .Q(
        g29242) );
  AND2X1 U13774 ( .IN1(n3628), .IN2(n13096), .Q(n13095) );
  OR4X1 U13775 ( .IN1(n13097), .IN2(n13098), .IN3(n13099), .IN4(n13100), .Q(
        n13096) );
  AND2X1 U13776 ( .IN1(n5596), .IN2(n13101), .Q(n13100) );
  OR2X1 U13777 ( .IN1(n13102), .IN2(n13103), .Q(n13101) );
  AND2X1 U13778 ( .IN1(g1760), .IN2(g1752), .Q(n13103) );
  AND2X1 U13779 ( .IN1(g1792), .IN2(g1744), .Q(n13102) );
  AND3X1 U13780 ( .IN1(n5602), .IN2(g1748), .IN3(n5359), .Q(n13099) );
  AND2X1 U13781 ( .IN1(n8483), .IN2(g1736), .Q(n13098) );
  INVX0 U13782 ( .INP(n11463), .ZN(n8483) );
  OR2X1 U13783 ( .IN1(n5596), .IN2(g1760), .Q(n11463) );
  AND2X1 U13784 ( .IN1(n9984), .IN2(g1756), .Q(n13097) );
  AND2X1 U13785 ( .IN1(g1783), .IN2(n5359), .Q(n9984) );
  AND2X1 U13786 ( .IN1(n8716), .IN2(n11449), .Q(n3628) );
  AND2X1 U13787 ( .IN1(n12563), .IN2(g1740), .Q(n13094) );
  AND2X1 U13788 ( .IN1(n8716), .IN2(n12566), .Q(n12563) );
  AND3X1 U13789 ( .IN1(g1760), .IN2(g1792), .IN3(n11449), .Q(n12566) );
  INVX0 U13790 ( .INP(n13104), .ZN(n11449) );
  AND2X1 U13791 ( .IN1(n8812), .IN2(g1792), .Q(n13093) );
  AND2X1 U13792 ( .IN1(n11452), .IN2(g1811), .Q(n13092) );
  AND2X1 U13793 ( .IN1(n8716), .IN2(n13104), .Q(n11452) );
  OR3X1 U13794 ( .IN1(n1169), .IN2(n12982), .IN3(n13105), .Q(n13104) );
  AND2X1 U13795 ( .IN1(n9786), .IN2(g2775), .Q(n13105) );
  OR2X1 U13796 ( .IN1(n5299), .IN2(g2719), .Q(n1169) );
  OR2X1 U13797 ( .IN1(n13106), .IN2(n13107), .Q(g29241) );
  AND2X1 U13798 ( .IN1(n13108), .IN2(g1677), .Q(n13107) );
  OR2X1 U13799 ( .IN1(n8802), .IN2(n13109), .Q(n13108) );
  AND2X1 U13800 ( .IN1(n11468), .IN2(n9015), .Q(n13109) );
  OR2X1 U13801 ( .IN1(n8488), .IN2(n8298), .Q(n9015) );
  AND2X1 U13802 ( .IN1(n13110), .IN2(g1691), .Q(n13106) );
  OR2X1 U13803 ( .IN1(n13111), .IN2(n11471), .Q(n13110) );
  AND2X1 U13804 ( .IN1(n4458), .IN2(n8690), .Q(n13111) );
  OR4X1 U13805 ( .IN1(n13112), .IN2(n13113), .IN3(n13114), .IN4(n13115), .Q(
        g29240) );
  AND2X1 U13806 ( .IN1(n11471), .IN2(g1677), .Q(n13115) );
  AND2X1 U13807 ( .IN1(n8716), .IN2(n13116), .Q(n11471) );
  AND2X1 U13808 ( .IN1(n3646), .IN2(n13117), .Q(n13114) );
  OR4X1 U13809 ( .IN1(n13118), .IN2(n13119), .IN3(n13120), .IN4(n13121), .Q(
        n13117) );
  AND2X1 U13810 ( .IN1(n13122), .IN2(n8499), .Q(n13121) );
  OR2X1 U13811 ( .IN1(n13123), .IN2(n13124), .Q(n13122) );
  AND2X1 U13812 ( .IN1(g1657), .IN2(g1608), .Q(n13124) );
  AND2X1 U13813 ( .IN1(g1624), .IN2(n9303), .Q(n13123) );
  AND3X1 U13814 ( .IN1(n5370), .IN2(g1612), .IN3(n5525), .Q(n13120) );
  AND2X1 U13815 ( .IN1(n8488), .IN2(g1600), .Q(n13119) );
  INVX0 U13816 ( .INP(n11484), .ZN(n8488) );
  OR2X1 U13817 ( .IN1(g1624), .IN2(n8499), .Q(n11484) );
  AND2X1 U13818 ( .IN1(g31863), .IN2(g1620), .Q(n13118) );
  AND2X1 U13819 ( .IN1(test_so94), .IN2(n5525), .Q(g31863) );
  AND2X1 U13820 ( .IN1(n8716), .IN2(n11468), .Q(n3646) );
  AND2X1 U13821 ( .IN1(n8811), .IN2(g1657), .Q(n13113) );
  AND2X1 U13822 ( .IN1(n12589), .IN2(g1604), .Q(n13112) );
  AND3X1 U13823 ( .IN1(g1657), .IN2(g1624), .IN3(n11468), .Q(n12589) );
  INVX0 U13824 ( .INP(n13116), .ZN(n11468) );
  OR2X1 U13825 ( .IN1(n13125), .IN2(n13044), .Q(n13116) );
  OR2X1 U13826 ( .IN1(n12982), .IN2(n12375), .Q(n13044) );
  OR2X1 U13827 ( .IN1(g2715), .IN2(g2719), .Q(n12375) );
  AND2X1 U13828 ( .IN1(n13126), .IN2(n9786), .Q(n12982) );
  INVX0 U13829 ( .INP(n4388), .ZN(n13126) );
  AND2X1 U13830 ( .IN1(n9786), .IN2(g2771), .Q(n13125) );
  AND2X1 U13831 ( .IN1(n5301), .IN2(n8347), .Q(n9786) );
  OR3X1 U13832 ( .IN1(n13127), .IN2(n13128), .IN3(n13129), .Q(g29239) );
  AND3X1 U13833 ( .IN1(n13130), .IN2(n13131), .IN3(n13132), .Q(n13129) );
  AND3X1 U13834 ( .IN1(n13133), .IN2(g1454), .IN3(n8747), .Q(n13128) );
  OR2X1 U13835 ( .IN1(n13130), .IN2(n13134), .Q(n13133) );
  XOR2X1 U13836 ( .IN1(n13135), .IN2(n5343), .Q(n13130) );
  AND2X1 U13837 ( .IN1(n8812), .IN2(g1478), .Q(n13127) );
  OR3X1 U13838 ( .IN1(n13136), .IN2(n13137), .IN3(n13138), .Q(g29238) );
  AND2X1 U13839 ( .IN1(n8811), .IN2(g1472), .Q(n13138) );
  AND2X1 U13840 ( .IN1(n13139), .IN2(g1484), .Q(n13137) );
  OR2X1 U13841 ( .IN1(n13140), .IN2(n13141), .Q(n13139) );
  AND2X1 U13842 ( .IN1(n13142), .IN2(n8690), .Q(n13140) );
  AND3X1 U13843 ( .IN1(n13142), .IN2(n13132), .IN3(n13143), .Q(n13136) );
  XOR2X1 U13844 ( .IN1(n13135), .IN2(n5483), .Q(n13142) );
  OR3X1 U13845 ( .IN1(n13144), .IN2(n13145), .IN3(n13146), .Q(g29237) );
  AND3X1 U13846 ( .IN1(n13147), .IN2(n13132), .IN3(n13148), .Q(n13146) );
  AND3X1 U13847 ( .IN1(n13149), .IN2(g1467), .IN3(n8747), .Q(n13145) );
  OR2X1 U13848 ( .IN1(n13147), .IN2(n13150), .Q(n13149) );
  INVX0 U13849 ( .INP(n13148), .ZN(n13150) );
  XOR2X1 U13850 ( .IN1(n13135), .IN2(n5290), .Q(n13147) );
  AND2X1 U13851 ( .IN1(n8812), .IN2(g1448), .Q(n13144) );
  OR3X1 U13852 ( .IN1(n13151), .IN2(n13152), .IN3(n13153), .Q(g29236) );
  AND3X1 U13853 ( .IN1(n13154), .IN2(n13132), .IN3(n13155), .Q(n13153) );
  AND3X1 U13854 ( .IN1(n8726), .IN2(n5850), .IN3(n8222), .Q(n13132) );
  AND3X1 U13855 ( .IN1(n13156), .IN2(g1437), .IN3(n8748), .Q(n13152) );
  OR2X1 U13856 ( .IN1(n13154), .IN2(n13157), .Q(n13156) );
  INVX0 U13857 ( .INP(n13155), .ZN(n13157) );
  XOR2X1 U13858 ( .IN1(n13135), .IN2(n5289), .Q(n13154) );
  OR2X1 U13859 ( .IN1(n9448), .IN2(n9267), .Q(n13135) );
  AND2X1 U13860 ( .IN1(n8811), .IN2(g1442), .Q(n13151) );
  OR3X1 U13861 ( .IN1(n13158), .IN2(n13159), .IN3(n13160), .Q(g29235) );
  AND2X1 U13862 ( .IN1(n8811), .IN2(g1252), .Q(n13160) );
  AND2X1 U13863 ( .IN1(n4178), .IN2(n5558), .Q(n13159) );
  AND3X1 U13864 ( .IN1(n11076), .IN2(n13161), .IN3(g1256), .Q(n13158) );
  INVX0 U13865 ( .INP(n4178), .ZN(n13161) );
  OR3X1 U13866 ( .IN1(n13162), .IN2(n13163), .IN3(n13164), .Q(g29234) );
  AND3X1 U13867 ( .IN1(n13165), .IN2(n13166), .IN3(n13167), .Q(n13164) );
  AND3X1 U13868 ( .IN1(test_so90), .IN2(n13168), .IN3(n8747), .Q(n13163) );
  OR2X1 U13869 ( .IN1(n13165), .IN2(n13169), .Q(n13168) );
  XOR2X1 U13870 ( .IN1(n13170), .IN2(n5478), .Q(n13165) );
  AND2X1 U13871 ( .IN1(n8811), .IN2(g1135), .Q(n13162) );
  OR3X1 U13872 ( .IN1(n13171), .IN2(n13172), .IN3(n13173), .Q(g29233) );
  AND2X1 U13873 ( .IN1(n8812), .IN2(g1129), .Q(n13173) );
  AND2X1 U13874 ( .IN1(n13174), .IN2(g1141), .Q(n13172) );
  OR2X1 U13875 ( .IN1(n13175), .IN2(n13176), .Q(n13174) );
  AND2X1 U13876 ( .IN1(n13177), .IN2(n8690), .Q(n13175) );
  AND3X1 U13877 ( .IN1(n13177), .IN2(n13167), .IN3(n13178), .Q(n13171) );
  XOR2X1 U13878 ( .IN1(n13170), .IN2(n5341), .Q(n13177) );
  OR3X1 U13879 ( .IN1(n13179), .IN2(n13180), .IN3(n13181), .Q(g29232) );
  AND3X1 U13880 ( .IN1(n13182), .IN2(n13167), .IN3(n13183), .Q(n13181) );
  AND3X1 U13881 ( .IN1(n13184), .IN2(g1124), .IN3(n8749), .Q(n13180) );
  OR2X1 U13882 ( .IN1(n13182), .IN2(n13185), .Q(n13184) );
  INVX0 U13883 ( .INP(n13183), .ZN(n13185) );
  XOR2X1 U13884 ( .IN1(n13170), .IN2(n5329), .Q(n13182) );
  AND2X1 U13885 ( .IN1(n8812), .IN2(g1105), .Q(n13179) );
  OR3X1 U13886 ( .IN1(n13186), .IN2(n13187), .IN3(n13188), .Q(g29231) );
  AND3X1 U13887 ( .IN1(n13189), .IN2(n13167), .IN3(n13190), .Q(n13188) );
  AND3X1 U13888 ( .IN1(n8518), .IN2(n8723), .IN3(n5851), .Q(n13167) );
  AND3X1 U13889 ( .IN1(n13191), .IN2(g1094), .IN3(n8749), .Q(n13187) );
  OR2X1 U13890 ( .IN1(n13189), .IN2(n13192), .Q(n13191) );
  INVX0 U13891 ( .INP(n13190), .ZN(n13192) );
  XOR2X1 U13892 ( .IN1(n13170), .IN2(n5328), .Q(n13189) );
  OR2X1 U13893 ( .IN1(n9449), .IN2(n9367), .Q(n13170) );
  INVX0 U13894 ( .INP(n11062), .ZN(n9449) );
  AND2X1 U13895 ( .IN1(test_so7), .IN2(n8809), .Q(n13186) );
  OR3X1 U13896 ( .IN1(n13193), .IN2(n13194), .IN3(n13195), .Q(g29230) );
  AND2X1 U13897 ( .IN1(n8822), .IN2(g907), .Q(n13195) );
  AND2X1 U13898 ( .IN1(n4196), .IN2(n5559), .Q(n13194) );
  AND3X1 U13899 ( .IN1(n11091), .IN2(n13196), .IN3(g911), .Q(n13193) );
  INVX0 U13900 ( .INP(n4196), .ZN(n13196) );
  OR3X1 U13901 ( .IN1(n13197), .IN2(n13198), .IN3(n13199), .Q(g29229) );
  AND2X1 U13902 ( .IN1(n8822), .IN2(g827), .Q(n13199) );
  AND3X1 U13903 ( .IN1(n4516), .IN2(n13200), .IN3(n5826), .Q(n13198) );
  AND2X1 U13904 ( .IN1(n4517), .IN2(g723), .Q(n13197) );
  OR2X1 U13905 ( .IN1(n13201), .IN2(n13202), .Q(g29228) );
  AND2X1 U13906 ( .IN1(n8822), .IN2(g736), .Q(n13202) );
  AND2X1 U13907 ( .IN1(n2404), .IN2(n13203), .Q(n13201) );
  XNOR2X1 U13908 ( .IN1(test_so60), .IN2(n12684), .Q(n13203) );
  OR2X1 U13909 ( .IN1(n13204), .IN2(n12692), .Q(n12684) );
  AND2X1 U13910 ( .IN1(n5482), .IN2(g12184), .Q(n13204) );
  OR3X1 U13911 ( .IN1(n13205), .IN2(n13206), .IN3(n13207), .Q(g29227) );
  AND2X1 U13912 ( .IN1(n8822), .IN2(g676), .Q(n13207) );
  AND2X1 U13913 ( .IN1(n4524), .IN2(test_so70), .Q(n13206) );
  AND3X1 U13914 ( .IN1(n4523), .IN2(n13208), .IN3(n8521), .Q(n13205) );
  OR3X1 U13915 ( .IN1(n13209), .IN2(n13210), .IN3(n13211), .Q(g29226) );
  AND2X1 U13916 ( .IN1(n8822), .IN2(g671), .Q(n13211) );
  AND3X1 U13917 ( .IN1(n4526), .IN2(n13208), .IN3(n5751), .Q(n13210) );
  AND3X1 U13918 ( .IN1(n4525), .IN2(n13212), .IN3(g676), .Q(n13209) );
  INVX0 U13919 ( .INP(n4526), .ZN(n13212) );
  OR2X1 U13920 ( .IN1(n13213), .IN2(n13214), .Q(g29225) );
  AND2X1 U13921 ( .IN1(n8822), .IN2(g667), .Q(n13214) );
  AND2X1 U13922 ( .IN1(n13215), .IN2(n4525), .Q(n13213) );
  AND2X1 U13923 ( .IN1(n8716), .IN2(n13208), .Q(n4525) );
  AND2X1 U13924 ( .IN1(g703), .IN2(n13216), .Q(n13208) );
  OR4X1 U13925 ( .IN1(n4535), .IN2(n13217), .IN3(n128), .IN4(n8349), .Q(n13216) );
  INVX0 U13926 ( .INP(n13218), .ZN(n13217) );
  XOR2X1 U13927 ( .IN1(g655), .IN2(g718), .Q(n4535) );
  XOR2X1 U13928 ( .IN1(n128), .IN2(n7980), .Q(n13215) );
  INVX0 U13929 ( .INP(n13219), .ZN(n128) );
  OR3X1 U13930 ( .IN1(n13220), .IN2(n13221), .IN3(n13222), .Q(g29224) );
  AND2X1 U13931 ( .IN1(n8822), .IN2(g572), .Q(n13222) );
  AND2X1 U13932 ( .IN1(n4201), .IN2(n5336), .Q(n13221) );
  AND3X1 U13933 ( .IN1(n2421), .IN2(n13223), .IN3(g586), .Q(n13220) );
  INVX0 U13934 ( .INP(n4201), .ZN(n13223) );
  OR3X1 U13935 ( .IN1(n13224), .IN2(n13225), .IN3(n13226), .Q(g29223) );
  AND2X1 U13936 ( .IN1(n13227), .IN2(n5708), .Q(n13226) );
  AND2X1 U13937 ( .IN1(n13228), .IN2(n8686), .Q(n13225) );
  INVX0 U13938 ( .INP(n13229), .ZN(n13228) );
  AND2X1 U13939 ( .IN1(n13230), .IN2(n13231), .Q(n13229) );
  OR2X1 U13940 ( .IN1(n13227), .IN2(n5708), .Q(n13230) );
  AND2X1 U13941 ( .IN1(g482), .IN2(n13232), .Q(n13227) );
  AND2X1 U13942 ( .IN1(n8822), .IN2(g482), .Q(n13224) );
  OR3X1 U13943 ( .IN1(n13233), .IN2(n13234), .IN3(n13235), .Q(g29222) );
  AND2X1 U13944 ( .IN1(n13236), .IN2(g411), .Q(n13235) );
  AND3X1 U13945 ( .IN1(n13237), .IN2(n3676), .IN3(n5358), .Q(n13234) );
  AND2X1 U13946 ( .IN1(n13238), .IN2(g417), .Q(n13233) );
  OR2X1 U13947 ( .IN1(n8801), .IN2(n13239), .Q(n13238) );
  AND2X1 U13948 ( .IN1(n4948), .IN2(n13240), .Q(n13239) );
  INVX0 U13949 ( .INP(n3676), .ZN(n13240) );
  XOR2X1 U13950 ( .IN1(n13241), .IN2(n5358), .Q(n3676) );
  OR2X1 U13951 ( .IN1(n13242), .IN2(n13243), .Q(n13241) );
  AND2X1 U13952 ( .IN1(n13244), .IN2(n8345), .Q(n13243) );
  OR2X1 U13953 ( .IN1(n13245), .IN2(n13246), .Q(n13244) );
  AND2X1 U13954 ( .IN1(n8344), .IN2(g424), .Q(n13246) );
  AND2X1 U13955 ( .IN1(g437), .IN2(g392), .Q(n13245) );
  AND2X1 U13956 ( .IN1(n13247), .IN2(g405), .Q(n13242) );
  OR2X1 U13957 ( .IN1(n13248), .IN2(n13249), .Q(n13247) );
  AND2X1 U13958 ( .IN1(g401), .IN2(g392), .Q(n13249) );
  AND2X1 U13959 ( .IN1(n8344), .IN2(g437), .Q(n13248) );
  OR3X1 U13960 ( .IN1(n13250), .IN2(n13251), .IN3(n13252), .Q(g28105) );
  AND2X1 U13961 ( .IN1(n10600), .IN2(g5011), .Q(n13252) );
  AND3X1 U13962 ( .IN1(n12727), .IN2(n10594), .IN3(n8750), .Q(n13251) );
  INVX0 U13963 ( .INP(n8479), .ZN(n10594) );
  OR2X1 U13964 ( .IN1(n13253), .IN2(n13254), .Q(n12727) );
  AND2X1 U13965 ( .IN1(n13255), .IN2(g6727), .Q(n13254) );
  OR4X1 U13966 ( .IN1(n13256), .IN2(n13257), .IN3(n13258), .IN4(n13259), .Q(
        n13255) );
  OR3X1 U13967 ( .IN1(n13260), .IN2(n13261), .IN3(n13262), .Q(n13259) );
  AND2X1 U13968 ( .IN1(n9003), .IN2(n13263), .Q(n13262) );
  OR2X1 U13969 ( .IN1(n13264), .IN2(n13265), .Q(n13263) );
  AND2X1 U13970 ( .IN1(g6641), .IN2(g17764), .Q(n13265) );
  AND2X1 U13971 ( .IN1(g6657), .IN2(g17722), .Q(n13264) );
  AND3X1 U13972 ( .IN1(g6609), .IN2(g17871), .IN3(n9002), .Q(n13261) );
  AND3X1 U13973 ( .IN1(g14749), .IN2(g6625), .IN3(n9005), .Q(n13260) );
  AND2X1 U13974 ( .IN1(n9004), .IN2(n13266), .Q(n13258) );
  OR2X1 U13975 ( .IN1(n13267), .IN2(n13268), .Q(n13266) );
  AND2X1 U13976 ( .IN1(g6581), .IN2(g13099), .Q(n13268) );
  AND2X1 U13977 ( .IN1(g6589), .IN2(g6723), .Q(n13267) );
  AND2X1 U13978 ( .IN1(test_so80), .IN2(n13269), .Q(n13257) );
  OR2X1 U13979 ( .IN1(n13270), .IN2(n13271), .Q(n13269) );
  AND2X1 U13980 ( .IN1(test_so71), .IN2(n9002), .Q(n13270) );
  AND2X1 U13981 ( .IN1(n13272), .IN2(n8497), .Q(n13256) );
  AND2X1 U13982 ( .IN1(n5531), .IN2(n13273), .Q(n13253) );
  OR4X1 U13983 ( .IN1(n13274), .IN2(n13275), .IN3(n13276), .IN4(n13277), .Q(
        n13273) );
  OR3X1 U13984 ( .IN1(n13278), .IN2(n13279), .IN3(n13280), .Q(n13277) );
  AND2X1 U13985 ( .IN1(n9005), .IN2(n13281), .Q(n13280) );
  OR2X1 U13986 ( .IN1(n13282), .IN2(n13283), .Q(n13281) );
  AND2X1 U13987 ( .IN1(g6593), .IN2(g13099), .Q(n13283) );
  AND2X1 U13988 ( .IN1(g6723), .IN2(g6605), .Q(n13282) );
  AND3X1 U13989 ( .IN1(g14749), .IN2(g6633), .IN3(n9004), .Q(n13279) );
  AND3X1 U13990 ( .IN1(g17871), .IN2(g6617), .IN3(n9003), .Q(n13278) );
  AND2X1 U13991 ( .IN1(n9002), .IN2(n13284), .Q(n13276) );
  OR2X1 U13992 ( .IN1(n13285), .IN2(n13286), .Q(n13284) );
  AND2X1 U13993 ( .IN1(g6597), .IN2(g17722), .Q(n13286) );
  AND2X1 U13994 ( .IN1(g17764), .IN2(g6649), .Q(n13285) );
  AND2X1 U13995 ( .IN1(test_so80), .IN2(n13287), .Q(n13275) );
  OR2X1 U13996 ( .IN1(n13288), .IN2(n13272), .Q(n13287) );
  OR3X1 U13997 ( .IN1(n13289), .IN2(n13290), .IN3(n13291), .Q(n13272) );
  AND3X1 U13998 ( .IN1(g14828), .IN2(g6621), .IN3(n9004), .Q(n13291) );
  AND3X1 U13999 ( .IN1(g6637), .IN2(g17778), .IN3(n9002), .Q(n13290) );
  AND2X1 U14000 ( .IN1(g6741), .IN2(n5590), .Q(n9002) );
  AND3X1 U14001 ( .IN1(g6653), .IN2(g17688), .IN3(n9005), .Q(n13289) );
  AND2X1 U14002 ( .IN1(n9003), .IN2(g6601), .Q(n13288) );
  AND2X1 U14003 ( .IN1(n13271), .IN2(n8497), .Q(n13274) );
  OR3X1 U14004 ( .IN1(n13292), .IN2(n13293), .IN3(n13294), .Q(n13271) );
  AND3X1 U14005 ( .IN1(g6645), .IN2(g17688), .IN3(n9004), .Q(n13294) );
  AND2X1 U14006 ( .IN1(n5590), .IN2(n5398), .Q(n9004) );
  AND3X1 U14007 ( .IN1(g14828), .IN2(g6613), .IN3(n9005), .Q(n13293) );
  AND2X1 U14008 ( .IN1(g6682), .IN2(n5398), .Q(n9005) );
  AND3X1 U14009 ( .IN1(g6629), .IN2(g17778), .IN3(n9003), .Q(n13292) );
  AND2X1 U14010 ( .IN1(g6682), .IN2(g6741), .Q(n9003) );
  AND2X1 U14011 ( .IN1(n8822), .IN2(g6657), .Q(n13250) );
  OR3X1 U14012 ( .IN1(n13295), .IN2(n13296), .IN3(n13297), .Q(g28102) );
  AND2X1 U14013 ( .IN1(n10617), .IN2(g4826), .Q(n13297) );
  AND3X1 U14014 ( .IN1(n10609), .IN2(n12759), .IN3(n8750), .Q(n13296) );
  OR2X1 U14015 ( .IN1(n13298), .IN2(n13299), .Q(n12759) );
  AND2X1 U14016 ( .IN1(n13300), .IN2(n8495), .Q(n13299) );
  OR4X1 U14017 ( .IN1(n13301), .IN2(n13302), .IN3(n13303), .IN4(n13304), .Q(
        n13300) );
  OR3X1 U14018 ( .IN1(n13305), .IN2(n13306), .IN3(n13307), .Q(n13304) );
  AND2X1 U14019 ( .IN1(n10608), .IN2(n13308), .Q(n13307) );
  OR2X1 U14020 ( .IN1(n13309), .IN2(n13310), .Q(n13308) );
  AND2X1 U14021 ( .IN1(g6251), .IN2(g17685), .Q(n13310) );
  AND2X1 U14022 ( .IN1(g17743), .IN2(g6303), .Q(n13309) );
  AND3X1 U14023 ( .IN1(g17845), .IN2(g6271), .IN3(n9821), .Q(n13306) );
  AND3X1 U14024 ( .IN1(g14705), .IN2(g6287), .IN3(n13311), .Q(n13305) );
  AND2X1 U14025 ( .IN1(n10612), .IN2(n13312), .Q(n13303) );
  OR2X1 U14026 ( .IN1(n13313), .IN2(n13314), .Q(n13312) );
  AND2X1 U14027 ( .IN1(g6247), .IN2(g13085), .Q(n13314) );
  AND2X1 U14028 ( .IN1(g6377), .IN2(g6259), .Q(n13313) );
  AND2X1 U14029 ( .IN1(n13315), .IN2(g12422), .Q(n13302) );
  OR2X1 U14030 ( .IN1(n13316), .IN2(n13317), .Q(n13315) );
  AND2X1 U14031 ( .IN1(n9821), .IN2(g6255), .Q(n13316) );
  AND2X1 U14032 ( .IN1(n5437), .IN2(n13318), .Q(n13301) );
  AND2X1 U14033 ( .IN1(test_so69), .IN2(n13319), .Q(n13298) );
  OR4X1 U14034 ( .IN1(n13320), .IN2(n13321), .IN3(n13322), .IN4(n13323), .Q(
        n13319) );
  OR3X1 U14035 ( .IN1(n13324), .IN2(n13325), .IN3(n13326), .Q(n13323) );
  AND2X1 U14036 ( .IN1(n13311), .IN2(n13327), .Q(n13326) );
  OR2X1 U14037 ( .IN1(n13328), .IN2(n13329), .Q(n13327) );
  AND2X1 U14038 ( .IN1(g6235), .IN2(g13085), .Q(n13329) );
  AND2X1 U14039 ( .IN1(g6243), .IN2(g6377), .Q(n13328) );
  AND3X1 U14040 ( .IN1(g14705), .IN2(g6279), .IN3(n10612), .Q(n13325) );
  AND3X1 U14041 ( .IN1(g6263), .IN2(g17845), .IN3(n10608), .Q(n13324) );
  AND2X1 U14042 ( .IN1(n9821), .IN2(n13330), .Q(n13322) );
  OR2X1 U14043 ( .IN1(n13331), .IN2(n13332), .Q(n13330) );
  AND2X1 U14044 ( .IN1(g6295), .IN2(g17743), .Q(n13332) );
  AND2X1 U14045 ( .IN1(g6311), .IN2(g17685), .Q(n13331) );
  AND2X1 U14046 ( .IN1(n13333), .IN2(g12422), .Q(n13321) );
  OR2X1 U14047 ( .IN1(n13334), .IN2(n13318), .Q(n13333) );
  OR3X1 U14048 ( .IN1(n13335), .IN2(n13336), .IN3(n13337), .Q(n13318) );
  AND3X1 U14049 ( .IN1(g14779), .IN2(g6267), .IN3(n10612), .Q(n13337) );
  AND3X1 U14050 ( .IN1(g6283), .IN2(g17760), .IN3(n9821), .Q(n13336) );
  AND3X1 U14051 ( .IN1(g6299), .IN2(g17649), .IN3(n13311), .Q(n13335) );
  AND2X1 U14052 ( .IN1(n10608), .IN2(g6239), .Q(n13334) );
  AND2X1 U14053 ( .IN1(n5437), .IN2(n13317), .Q(n13320) );
  OR3X1 U14054 ( .IN1(n13338), .IN2(n13339), .IN3(n13340), .Q(n13317) );
  AND3X1 U14055 ( .IN1(g6307), .IN2(g17649), .IN3(n10612), .Q(n13340) );
  AND3X1 U14056 ( .IN1(g6291), .IN2(g17760), .IN3(n10608), .Q(n13339) );
  AND3X1 U14057 ( .IN1(g14779), .IN2(g6275), .IN3(n13311), .Q(n13338) );
  AND2X1 U14058 ( .IN1(n8822), .IN2(g6311), .Q(n13295) );
  OR3X1 U14059 ( .IN1(n13341), .IN2(n13342), .IN3(n13343), .Q(g28099) );
  AND2X1 U14060 ( .IN1(n10634), .IN2(g4831), .Q(n13343) );
  AND3X1 U14061 ( .IN1(n10626), .IN2(n12791), .IN3(n8750), .Q(n13342) );
  OR2X1 U14062 ( .IN1(n13344), .IN2(n13345), .Q(n12791) );
  AND2X1 U14063 ( .IN1(n13346), .IN2(g6035), .Q(n13345) );
  OR4X1 U14064 ( .IN1(n13347), .IN2(n13348), .IN3(n13349), .IN4(n13350), .Q(
        n13346) );
  OR3X1 U14065 ( .IN1(n13351), .IN2(n13352), .IN3(n13353), .Q(n13350) );
  AND2X1 U14066 ( .IN1(n13354), .IN2(n13355), .Q(n13353) );
  OR2X1 U14067 ( .IN1(n13356), .IN2(n13357), .Q(n13355) );
  AND2X1 U14068 ( .IN1(g5889), .IN2(g13068), .Q(n13357) );
  AND2X1 U14069 ( .IN1(g5897), .IN2(g6031), .Q(n13356) );
  AND3X1 U14070 ( .IN1(g14673), .IN2(g5933), .IN3(n10629), .Q(n13352) );
  AND3X1 U14071 ( .IN1(n10625), .IN2(g17819), .IN3(test_so28), .Q(n13351) );
  AND2X1 U14072 ( .IN1(n9834), .IN2(n13358), .Q(n13349) );
  OR2X1 U14073 ( .IN1(n13359), .IN2(n13360), .Q(n13358) );
  AND2X1 U14074 ( .IN1(test_so13), .IN2(g17646), .Q(n13360) );
  AND2X1 U14075 ( .IN1(g5949), .IN2(g17715), .Q(n13359) );
  AND2X1 U14076 ( .IN1(n13361), .IN2(g12350), .Q(n13348) );
  OR2X1 U14077 ( .IN1(n13362), .IN2(n13363), .Q(n13361) );
  AND2X1 U14078 ( .IN1(n10625), .IN2(g5893), .Q(n13362) );
  AND2X1 U14079 ( .IN1(n5432), .IN2(n13364), .Q(n13347) );
  AND2X1 U14080 ( .IN1(n5528), .IN2(n13365), .Q(n13344) );
  OR4X1 U14081 ( .IN1(n13366), .IN2(n13367), .IN3(n13368), .IN4(n13369), .Q(
        n13365) );
  OR3X1 U14082 ( .IN1(n13370), .IN2(n13371), .IN3(n13372), .Q(n13369) );
  AND2X1 U14083 ( .IN1(n10625), .IN2(n13373), .Q(n13372) );
  OR2X1 U14084 ( .IN1(n13374), .IN2(n13375), .Q(n13373) );
  AND2X1 U14085 ( .IN1(g5905), .IN2(g17646), .Q(n13375) );
  AND2X1 U14086 ( .IN1(g17715), .IN2(g5957), .Q(n13374) );
  AND3X1 U14087 ( .IN1(g17819), .IN2(g5925), .IN3(n9834), .Q(n13371) );
  AND3X1 U14088 ( .IN1(g14673), .IN2(g5941), .IN3(n13354), .Q(n13370) );
  AND2X1 U14089 ( .IN1(n10629), .IN2(n13376), .Q(n13368) );
  OR2X1 U14090 ( .IN1(n13377), .IN2(n13378), .Q(n13376) );
  AND2X1 U14091 ( .IN1(g5901), .IN2(g13068), .Q(n13378) );
  AND2X1 U14092 ( .IN1(g6031), .IN2(g5913), .Q(n13377) );
  AND2X1 U14093 ( .IN1(n13379), .IN2(g12350), .Q(n13367) );
  OR2X1 U14094 ( .IN1(n13380), .IN2(n13364), .Q(n13379) );
  OR3X1 U14095 ( .IN1(n13381), .IN2(n13382), .IN3(n13383), .Q(n13364) );
  AND3X1 U14096 ( .IN1(g5961), .IN2(g17607), .IN3(n10629), .Q(n13383) );
  AND3X1 U14097 ( .IN1(g5945), .IN2(g17739), .IN3(n10625), .Q(n13382) );
  AND3X1 U14098 ( .IN1(g14738), .IN2(g5929), .IN3(n13354), .Q(n13381) );
  AND2X1 U14099 ( .IN1(n9834), .IN2(g5909), .Q(n13380) );
  AND2X1 U14100 ( .IN1(n5432), .IN2(n13363), .Q(n13366) );
  OR3X1 U14101 ( .IN1(n13384), .IN2(n13385), .IN3(n13386), .Q(n13363) );
  AND3X1 U14102 ( .IN1(g14738), .IN2(g5921), .IN3(n10629), .Q(n13386) );
  AND3X1 U14103 ( .IN1(g5937), .IN2(g17739), .IN3(n9834), .Q(n13385) );
  AND3X1 U14104 ( .IN1(g5953), .IN2(g17607), .IN3(n13354), .Q(n13384) );
  AND2X1 U14105 ( .IN1(test_so13), .IN2(n8808), .Q(n13341) );
  OR3X1 U14106 ( .IN1(n13387), .IN2(n13388), .IN3(n13389), .Q(g28096) );
  AND2X1 U14107 ( .IN1(n10650), .IN2(g4821), .Q(n13389) );
  AND3X1 U14108 ( .IN1(n10642), .IN2(n12823), .IN3(n8751), .Q(n13388) );
  OR2X1 U14109 ( .IN1(n13390), .IN2(n13391), .Q(n12823) );
  AND2X1 U14110 ( .IN1(n13392), .IN2(g5689), .Q(n13391) );
  OR4X1 U14111 ( .IN1(n13393), .IN2(n13394), .IN3(n13395), .IN4(n13396), .Q(
        n13392) );
  OR3X1 U14112 ( .IN1(n13397), .IN2(n13398), .IN3(n13399), .Q(n13396) );
  AND2X1 U14113 ( .IN1(n13400), .IN2(n13401), .Q(n13399) );
  OR2X1 U14114 ( .IN1(n13402), .IN2(n13403), .Q(n13401) );
  AND2X1 U14115 ( .IN1(g5543), .IN2(g13049), .Q(n13403) );
  AND2X1 U14116 ( .IN1(g5551), .IN2(g5685), .Q(n13402) );
  AND3X1 U14117 ( .IN1(g14635), .IN2(g5587), .IN3(n10645), .Q(n13398) );
  AND3X1 U14118 ( .IN1(g5571), .IN2(g17813), .IN3(n10641), .Q(n13397) );
  AND2X1 U14119 ( .IN1(n9826), .IN2(n13404), .Q(n13395) );
  OR2X1 U14120 ( .IN1(n13405), .IN2(n13406), .Q(n13404) );
  AND2X1 U14121 ( .IN1(g5603), .IN2(g17678), .Q(n13406) );
  AND2X1 U14122 ( .IN1(g5619), .IN2(g17604), .Q(n13405) );
  AND2X1 U14123 ( .IN1(n13407), .IN2(g12300), .Q(n13394) );
  OR2X1 U14124 ( .IN1(n13408), .IN2(n13409), .Q(n13407) );
  AND2X1 U14125 ( .IN1(n10641), .IN2(g5547), .Q(n13408) );
  AND2X1 U14126 ( .IN1(n5439), .IN2(n13410), .Q(n13393) );
  AND2X1 U14127 ( .IN1(n5529), .IN2(n13411), .Q(n13390) );
  OR4X1 U14128 ( .IN1(n13412), .IN2(n13413), .IN3(n13414), .IN4(n13415), .Q(
        n13411) );
  OR3X1 U14129 ( .IN1(n13416), .IN2(n13417), .IN3(n13418), .Q(n13415) );
  AND2X1 U14130 ( .IN1(n10641), .IN2(n13419), .Q(n13418) );
  OR2X1 U14131 ( .IN1(n13420), .IN2(n13421), .Q(n13419) );
  AND2X1 U14132 ( .IN1(test_so6), .IN2(g17604), .Q(n13421) );
  AND2X1 U14133 ( .IN1(g17678), .IN2(g5611), .Q(n13420) );
  AND3X1 U14134 ( .IN1(g17813), .IN2(g5579), .IN3(n9826), .Q(n13417) );
  AND3X1 U14135 ( .IN1(g14635), .IN2(g5595), .IN3(n13400), .Q(n13416) );
  AND2X1 U14136 ( .IN1(n10645), .IN2(n13422), .Q(n13414) );
  OR2X1 U14137 ( .IN1(n13423), .IN2(n13424), .Q(n13422) );
  AND2X1 U14138 ( .IN1(g5555), .IN2(g13049), .Q(n13424) );
  AND2X1 U14139 ( .IN1(g5685), .IN2(g5567), .Q(n13423) );
  AND2X1 U14140 ( .IN1(n13425), .IN2(g12300), .Q(n13413) );
  OR2X1 U14141 ( .IN1(n13426), .IN2(n13410), .Q(n13425) );
  OR3X1 U14142 ( .IN1(n13427), .IN2(n13428), .IN3(n13429), .Q(n13410) );
  AND3X1 U14143 ( .IN1(g5615), .IN2(g17580), .IN3(n10645), .Q(n13429) );
  AND3X1 U14144 ( .IN1(g5599), .IN2(g17711), .IN3(n10641), .Q(n13428) );
  AND3X1 U14145 ( .IN1(g14694), .IN2(g5583), .IN3(n13400), .Q(n13427) );
  AND2X1 U14146 ( .IN1(n9826), .IN2(g5563), .Q(n13426) );
  AND2X1 U14147 ( .IN1(n5439), .IN2(n13409), .Q(n13412) );
  OR3X1 U14148 ( .IN1(n13430), .IN2(n13431), .IN3(n13432), .Q(n13409) );
  AND3X1 U14149 ( .IN1(g14694), .IN2(g5575), .IN3(n10645), .Q(n13432) );
  AND3X1 U14150 ( .IN1(n9826), .IN2(g17711), .IN3(test_so5), .Q(n13431) );
  AND3X1 U14151 ( .IN1(g5607), .IN2(g17580), .IN3(n13400), .Q(n13430) );
  AND2X1 U14152 ( .IN1(n8822), .IN2(g5619), .Q(n13387) );
  OR3X1 U14153 ( .IN1(n13433), .IN2(n13434), .IN3(n13435), .Q(g28093) );
  AND2X1 U14154 ( .IN1(n10662), .IN2(g29220), .Q(n13435) );
  AND3X1 U14155 ( .IN1(n12855), .IN2(g33959), .IN3(n8750), .Q(n13434) );
  INVX0 U14156 ( .INP(n8474), .ZN(g33959) );
  OR2X1 U14157 ( .IN1(n13436), .IN2(n13437), .Q(n12855) );
  AND2X1 U14158 ( .IN1(n13438), .IN2(n8494), .Q(n13437) );
  OR4X1 U14159 ( .IN1(n13439), .IN2(n13440), .IN3(n13441), .IN4(n13442), .Q(
        n13438) );
  OR3X1 U14160 ( .IN1(n13443), .IN2(n13444), .IN3(n13445), .Q(n13442) );
  AND2X1 U14161 ( .IN1(n8996), .IN2(n13446), .Q(n13445) );
  OR2X1 U14162 ( .IN1(n13447), .IN2(n13448), .Q(n13446) );
  AND2X1 U14163 ( .IN1(g5208), .IN2(g13039), .Q(n13448) );
  AND2X1 U14164 ( .IN1(g5220), .IN2(g5339), .Q(n13447) );
  AND3X1 U14165 ( .IN1(g17787), .IN2(g5232), .IN3(g31860), .Q(n13444) );
  AND3X1 U14166 ( .IN1(g14597), .IN2(g5248), .IN3(n8995), .Q(n13443) );
  AND2X1 U14167 ( .IN1(n8997), .IN2(n13449), .Q(n13441) );
  OR2X1 U14168 ( .IN1(n13450), .IN2(n13451), .Q(n13449) );
  AND2X1 U14169 ( .IN1(g5212), .IN2(g17577), .Q(n13451) );
  AND2X1 U14170 ( .IN1(g17639), .IN2(g5264), .Q(n13450) );
  AND2X1 U14171 ( .IN1(n13452), .IN2(g12238), .Q(n13440) );
  OR2X1 U14172 ( .IN1(n13453), .IN2(n13454), .Q(n13452) );
  AND2X1 U14173 ( .IN1(g31860), .IN2(g5216), .Q(n13453) );
  AND2X1 U14174 ( .IN1(n5438), .IN2(n13455), .Q(n13439) );
  AND2X1 U14175 ( .IN1(test_so10), .IN2(n13456), .Q(n13436) );
  OR4X1 U14176 ( .IN1(n13457), .IN2(n13458), .IN3(n13459), .IN4(n13460), .Q(
        n13456) );
  OR3X1 U14177 ( .IN1(n13461), .IN2(n13462), .IN3(n13463), .Q(n13460) );
  AND2X1 U14178 ( .IN1(n8995), .IN2(n13464), .Q(n13463) );
  OR2X1 U14179 ( .IN1(n13465), .IN2(n13466), .Q(n13464) );
  AND2X1 U14180 ( .IN1(g5196), .IN2(g13039), .Q(n13466) );
  AND2X1 U14181 ( .IN1(g5339), .IN2(g5204), .Q(n13465) );
  AND3X1 U14182 ( .IN1(g5224), .IN2(g17787), .IN3(n8997), .Q(n13462) );
  AND3X1 U14183 ( .IN1(g14597), .IN2(g5240), .IN3(n8996), .Q(n13461) );
  AND2X1 U14184 ( .IN1(g31860), .IN2(n13467), .Q(n13459) );
  OR2X1 U14185 ( .IN1(n13468), .IN2(n13469), .Q(n13467) );
  AND2X1 U14186 ( .IN1(g5256), .IN2(g17639), .Q(n13469) );
  AND2X1 U14187 ( .IN1(g5272), .IN2(g17577), .Q(n13468) );
  AND2X1 U14188 ( .IN1(n13470), .IN2(g12238), .Q(n13458) );
  OR2X1 U14189 ( .IN1(n13471), .IN2(n13455), .Q(n13470) );
  OR3X1 U14190 ( .IN1(n13472), .IN2(n13473), .IN3(n13474), .Q(n13455) );
  AND3X1 U14191 ( .IN1(g5244), .IN2(g17674), .IN3(g31860), .Q(n13474) );
  AND2X1 U14192 ( .IN1(g5297), .IN2(g5357), .Q(g31860) );
  AND3X1 U14193 ( .IN1(g5260), .IN2(g17519), .IN3(n8995), .Q(n13473) );
  AND3X1 U14194 ( .IN1(n8996), .IN2(g14662), .IN3(test_so82), .Q(n13472) );
  AND2X1 U14195 ( .IN1(n8997), .IN2(g5200), .Q(n13471) );
  AND2X1 U14196 ( .IN1(n5438), .IN2(n13454), .Q(n13457) );
  OR3X1 U14197 ( .IN1(n13475), .IN2(n13476), .IN3(n13477), .Q(n13454) );
  AND3X1 U14198 ( .IN1(g5252), .IN2(g17674), .IN3(n8997), .Q(n13477) );
  AND2X1 U14199 ( .IN1(g5357), .IN2(n5588), .Q(n8997) );
  AND3X1 U14200 ( .IN1(g14662), .IN2(g5236), .IN3(n8995), .Q(n13476) );
  AND2X1 U14201 ( .IN1(n5393), .IN2(n5588), .Q(n8995) );
  AND3X1 U14202 ( .IN1(g5268), .IN2(g17519), .IN3(n8996), .Q(n13475) );
  AND2X1 U14203 ( .IN1(g5297), .IN2(n5393), .Q(n8996) );
  AND2X1 U14204 ( .IN1(n8822), .IN2(g5272), .Q(n13433) );
  OR2X1 U14205 ( .IN1(n13478), .IN2(n13479), .Q(g28092) );
  AND3X1 U14206 ( .IN1(n11582), .IN2(n11581), .IN3(n8751), .Q(n13479) );
  OR3X1 U14207 ( .IN1(g84), .IN2(n13480), .IN3(g5052), .Q(n11581) );
  OR3X1 U14208 ( .IN1(n13481), .IN2(n13480), .IN3(g5041), .Q(n11582) );
  OR3X1 U14209 ( .IN1(n8437), .IN2(n5615), .IN3(g5046), .Q(n13480) );
  AND2X1 U14210 ( .IN1(n8822), .IN2(g5057), .Q(n13478) );
  OR2X1 U14211 ( .IN1(n13482), .IN2(n13483), .Q(g28091) );
  AND3X1 U14212 ( .IN1(n11583), .IN2(n11585), .IN3(n8750), .Q(n13483) );
  OR3X1 U14213 ( .IN1(n5607), .IN2(g84), .IN3(n13484), .Q(n11585) );
  OR3X1 U14214 ( .IN1(n5605), .IN2(n13484), .IN3(n13481), .Q(n11583) );
  INVX0 U14215 ( .INP(g84), .ZN(n13481) );
  OR3X1 U14216 ( .IN1(n8438), .IN2(n5578), .IN3(g5057), .Q(n13484) );
  AND2X1 U14217 ( .IN1(n8821), .IN2(g5069), .Q(n13482) );
  OR2X1 U14218 ( .IN1(n13485), .IN2(n13486), .Q(g28090) );
  AND2X1 U14219 ( .IN1(n10689), .IN2(g4961), .Q(n13486) );
  AND3X1 U14220 ( .IN1(n13487), .IN2(n8723), .IN3(n9869), .Q(n13485) );
  AND2X1 U14221 ( .IN1(n9065), .IN2(n9057), .Q(n9869) );
  OR2X1 U14222 ( .IN1(n13488), .IN2(g4961), .Q(n13487) );
  AND2X1 U14223 ( .IN1(n10681), .IN2(n13489), .Q(n13488) );
  OR4X1 U14224 ( .IN1(n13490), .IN2(n13491), .IN3(n13492), .IN4(n13493), .Q(
        n13489) );
  AND2X1 U14225 ( .IN1(n8416), .IN2(n10680), .Q(n13493) );
  AND2X1 U14226 ( .IN1(n9820), .IN2(g4049), .Q(n13492) );
  AND2X1 U14227 ( .IN1(n8089), .IN2(n13494), .Q(n13491) );
  AND2X1 U14228 ( .IN1(n10684), .IN2(g4045), .Q(n13490) );
  OR2X1 U14229 ( .IN1(n13495), .IN2(n13496), .Q(g28089) );
  AND2X1 U14230 ( .IN1(n10705), .IN2(g4950), .Q(n13496) );
  AND3X1 U14231 ( .IN1(n13497), .IN2(n8725), .IN3(n9877), .Q(n13495) );
  AND2X1 U14232 ( .IN1(n9064), .IN2(n9057), .Q(n9877) );
  OR2X1 U14233 ( .IN1(n13498), .IN2(g4950), .Q(n13497) );
  AND2X1 U14234 ( .IN1(n10697), .IN2(n13499), .Q(n13498) );
  OR4X1 U14235 ( .IN1(n13500), .IN2(n13501), .IN3(n13502), .IN4(n13503), .Q(
        n13499) );
  AND2X1 U14236 ( .IN1(n8425), .IN2(n10696), .Q(n13503) );
  AND2X1 U14237 ( .IN1(n9833), .IN2(g3698), .Q(n13502) );
  AND2X1 U14238 ( .IN1(n8087), .IN2(n13504), .Q(n13501) );
  AND2X1 U14239 ( .IN1(n10700), .IN2(g3694), .Q(n13500) );
  OR2X1 U14240 ( .IN1(n13505), .IN2(n13506), .Q(g28088) );
  AND2X1 U14241 ( .IN1(n10719), .IN2(g4939), .Q(n13506) );
  AND3X1 U14242 ( .IN1(n13507), .IN2(n8724), .IN3(n9884), .Q(n13505) );
  AND3X1 U14243 ( .IN1(n5360), .IN2(n5517), .IN3(n9057), .Q(n9884) );
  OR2X1 U14244 ( .IN1(n13508), .IN2(g4939), .Q(n13507) );
  AND2X1 U14245 ( .IN1(n10715), .IN2(n13509), .Q(n13508) );
  OR4X1 U14246 ( .IN1(n13510), .IN2(n13511), .IN3(n13512), .IN4(n13513), .Q(
        n13509) );
  AND2X1 U14247 ( .IN1(n8413), .IN2(n10714), .Q(n13513) );
  AND2X1 U14248 ( .IN1(n9825), .IN2(g3347), .Q(n13512) );
  AND2X1 U14249 ( .IN1(n8084), .IN2(n13514), .Q(n13511) );
  AND2X1 U14250 ( .IN1(n10712), .IN2(g3343), .Q(n13510) );
  OR2X1 U14251 ( .IN1(n13515), .IN2(n13516), .Q(g28087) );
  AND2X1 U14252 ( .IN1(n10600), .IN2(g4894), .Q(n13516) );
  AND2X1 U14253 ( .IN1(n8716), .IN2(n8479), .Q(n10600) );
  OR2X1 U14254 ( .IN1(n13517), .IN2(n5713), .Q(n8479) );
  AND2X1 U14255 ( .IN1(n13518), .IN2(n10557), .Q(n13517) );
  AND3X1 U14256 ( .IN1(g4888), .IN2(n5360), .IN3(n5517), .Q(n10557) );
  AND3X1 U14257 ( .IN1(n13519), .IN2(n8724), .IN3(n9508), .Q(n13515) );
  AND2X1 U14258 ( .IN1(n9067), .IN2(n9057), .Q(n9508) );
  AND2X1 U14259 ( .IN1(g4983), .IN2(n9068), .Q(n9057) );
  OR2X1 U14260 ( .IN1(n4689), .IN2(g4894), .Q(n13519) );
  OR2X1 U14261 ( .IN1(n13520), .IN2(n13521), .Q(g28086) );
  AND2X1 U14262 ( .IN1(n10617), .IN2(g4771), .Q(n13521) );
  AND2X1 U14263 ( .IN1(n8716), .IN2(n10613), .Q(n10617) );
  AND3X1 U14264 ( .IN1(n13522), .IN2(n8723), .IN3(n9905), .Q(n13520) );
  AND2X1 U14265 ( .IN1(n9039), .IN2(n9031), .Q(n9905) );
  OR2X1 U14266 ( .IN1(n13523), .IN2(g4771), .Q(n13522) );
  AND2X1 U14267 ( .IN1(n10609), .IN2(n13524), .Q(n13523) );
  OR4X1 U14268 ( .IN1(n13525), .IN2(n13526), .IN3(n13527), .IN4(n13528), .Q(
        n13524) );
  AND2X1 U14269 ( .IN1(n8085), .IN2(n13311), .Q(n13528) );
  AND2X1 U14270 ( .IN1(n5396), .IN2(n5592), .Q(n13311) );
  AND2X1 U14271 ( .IN1(n10612), .IN2(g6386), .Q(n13527) );
  AND2X1 U14272 ( .IN1(g6336), .IN2(n5396), .Q(n10612) );
  AND2X1 U14273 ( .IN1(n8414), .IN2(n10608), .Q(n13526) );
  AND2X1 U14274 ( .IN1(g6395), .IN2(n5592), .Q(n10608) );
  AND2X1 U14275 ( .IN1(n9821), .IN2(g6390), .Q(n13525) );
  AND2X1 U14276 ( .IN1(g6336), .IN2(g6395), .Q(n9821) );
  INVX0 U14277 ( .INP(n10613), .ZN(n10609) );
  OR2X1 U14278 ( .IN1(n13529), .IN2(n5656), .Q(n10613) );
  AND3X1 U14279 ( .IN1(n13530), .IN2(g4765), .IN3(n9041), .Q(n13529) );
  OR2X1 U14280 ( .IN1(n13531), .IN2(n13532), .Q(g28085) );
  AND2X1 U14281 ( .IN1(n10634), .IN2(g4760), .Q(n13532) );
  AND2X1 U14282 ( .IN1(n8716), .IN2(n10630), .Q(n10634) );
  AND3X1 U14283 ( .IN1(n13533), .IN2(n8723), .IN3(n9913), .Q(n13531) );
  AND2X1 U14284 ( .IN1(n9038), .IN2(n9031), .Q(n9913) );
  OR2X1 U14285 ( .IN1(n13534), .IN2(g4760), .Q(n13533) );
  AND2X1 U14286 ( .IN1(n10626), .IN2(n13535), .Q(n13534) );
  OR4X1 U14287 ( .IN1(n13536), .IN2(n13537), .IN3(n13538), .IN4(n13539), .Q(
        n13535) );
  AND2X1 U14288 ( .IN1(n8086), .IN2(n13354), .Q(n13539) );
  AND2X1 U14289 ( .IN1(n8503), .IN2(n5589), .Q(n13354) );
  AND2X1 U14290 ( .IN1(n10629), .IN2(g6040), .Q(n13538) );
  AND2X1 U14291 ( .IN1(n8503), .IN2(g5990), .Q(n10629) );
  AND2X1 U14292 ( .IN1(test_so50), .IN2(n9834), .Q(n13537) );
  AND2X1 U14293 ( .IN1(g5990), .IN2(test_so57), .Q(n9834) );
  AND2X1 U14294 ( .IN1(n10625), .IN2(n8512), .Q(n13536) );
  AND2X1 U14295 ( .IN1(test_so57), .IN2(n5589), .Q(n10625) );
  INVX0 U14296 ( .INP(n10630), .ZN(n10626) );
  OR2X1 U14297 ( .IN1(n13540), .IN2(n8224), .Q(n10630) );
  AND3X1 U14298 ( .IN1(n13530), .IN2(g4754), .IN3(n9039), .Q(n13540) );
  AND2X1 U14299 ( .IN1(g4709), .IN2(n5361), .Q(n9039) );
  OR2X1 U14300 ( .IN1(n13541), .IN2(n13542), .Q(g28084) );
  AND2X1 U14301 ( .IN1(n10650), .IN2(test_so18), .Q(n13542) );
  AND2X1 U14302 ( .IN1(n8716), .IN2(n10646), .Q(n10650) );
  AND3X1 U14303 ( .IN1(n13543), .IN2(n8724), .IN3(n9920), .Q(n13541) );
  AND3X1 U14304 ( .IN1(n5361), .IN2(n5518), .IN3(n9031), .Q(n9920) );
  OR2X1 U14305 ( .IN1(n13544), .IN2(test_so18), .Q(n13543) );
  AND2X1 U14306 ( .IN1(n10642), .IN2(n13545), .Q(n13544) );
  OR4X1 U14307 ( .IN1(n13546), .IN2(n13547), .IN3(n13548), .IN4(n13549), .Q(
        n13545) );
  AND2X1 U14308 ( .IN1(n8088), .IN2(n13400), .Q(n13549) );
  AND2X1 U14309 ( .IN1(n5397), .IN2(n5593), .Q(n13400) );
  AND2X1 U14310 ( .IN1(n10645), .IN2(g5694), .Q(n13548) );
  AND2X1 U14311 ( .IN1(g5644), .IN2(n5397), .Q(n10645) );
  AND2X1 U14312 ( .IN1(n8424), .IN2(n10641), .Q(n13547) );
  AND2X1 U14313 ( .IN1(g5703), .IN2(n5593), .Q(n10641) );
  AND2X1 U14314 ( .IN1(n9826), .IN2(g5698), .Q(n13546) );
  AND2X1 U14315 ( .IN1(g5644), .IN2(g5703), .Q(n9826) );
  INVX0 U14316 ( .INP(n10646), .ZN(n10642) );
  OR2X1 U14317 ( .IN1(n13550), .IN2(n5440), .Q(n10646) );
  AND3X1 U14318 ( .IN1(n13530), .IN2(g4743), .IN3(n9038), .Q(n13550) );
  AND2X1 U14319 ( .IN1(g4785), .IN2(n5518), .Q(n9038) );
  OR2X1 U14320 ( .IN1(n13551), .IN2(n13552), .Q(g28083) );
  AND2X1 U14321 ( .IN1(n10662), .IN2(g4704), .Q(n13552) );
  AND2X1 U14322 ( .IN1(n8717), .IN2(n8474), .Q(n10662) );
  OR2X1 U14323 ( .IN1(n13553), .IN2(n5712), .Q(n8474) );
  AND2X1 U14324 ( .IN1(n13530), .IN2(n10586), .Q(n13553) );
  AND3X1 U14325 ( .IN1(g4698), .IN2(n5361), .IN3(n5518), .Q(n10586) );
  AND3X1 U14326 ( .IN1(n10046), .IN2(n9042), .IN3(n5368), .Q(n13530) );
  AND3X1 U14327 ( .IN1(g4659), .IN2(g4669), .IN3(test_so19), .Q(n10046) );
  AND3X1 U14328 ( .IN1(n13554), .IN2(n8724), .IN3(n9511), .Q(n13551) );
  AND2X1 U14329 ( .IN1(n9041), .IN2(n9031), .Q(n9511) );
  AND2X1 U14330 ( .IN1(g4793), .IN2(n9042), .Q(n9031) );
  AND2X1 U14331 ( .IN1(n8504), .IN2(g4776), .Q(n9042) );
  AND2X1 U14332 ( .IN1(g4709), .IN2(g4785), .Q(n9041) );
  OR2X1 U14333 ( .IN1(n4708), .IN2(g4704), .Q(n13554) );
  OR2X1 U14334 ( .IN1(n13555), .IN2(n13556), .Q(g28082) );
  AND3X1 U14335 ( .IN1(n9390), .IN2(n8724), .IN3(n5752), .Q(n13556) );
  AND2X1 U14336 ( .IN1(n13557), .IN2(g4521), .Q(n13555) );
  OR2X1 U14337 ( .IN1(n8802), .IN2(n13558), .Q(n13557) );
  XNOR2X1 U14338 ( .IN1(n10053), .IN2(n8185), .Q(n13558) );
  OR3X1 U14339 ( .IN1(n13559), .IN2(n13560), .IN3(n13561), .Q(g28074) );
  AND2X1 U14340 ( .IN1(n8821), .IN2(g4119), .Q(n13561) );
  AND2X1 U14341 ( .IN1(n4714), .IN2(n4721), .Q(n13560) );
  AND3X1 U14342 ( .IN1(n8727), .IN2(g4122), .IN3(n13562), .Q(n13559) );
  INVX0 U14343 ( .INP(n4714), .ZN(n13562) );
  OR3X1 U14344 ( .IN1(n13563), .IN2(n13564), .IN3(n13565), .Q(g28073) );
  AND2X1 U14345 ( .IN1(n13566), .IN2(n4721), .Q(n13565) );
  AND2X1 U14346 ( .IN1(n8821), .IN2(g4116), .Q(n13564) );
  AND3X1 U14347 ( .IN1(n13567), .IN2(g4119), .IN3(n8731), .Q(n13563) );
  INVX0 U14348 ( .INP(n13566), .ZN(n13567) );
  AND2X1 U14349 ( .IN1(g4057), .IN2(n13568), .Q(n13566) );
  OR3X1 U14350 ( .IN1(n13569), .IN2(n13570), .IN3(n13571), .Q(g28072) );
  AND2X1 U14351 ( .IN1(n13572), .IN2(n4721), .Q(n13571) );
  AND2X1 U14352 ( .IN1(n8821), .IN2(g4112), .Q(n13570) );
  AND3X1 U14353 ( .IN1(n13573), .IN2(g4116), .IN3(n8733), .Q(n13569) );
  INVX0 U14354 ( .INP(n13572), .ZN(n13573) );
  AND3X1 U14355 ( .IN1(g4064), .IN2(n5711), .IN3(n4722), .Q(n13572) );
  OR2X1 U14356 ( .IN1(n13574), .IN2(n13575), .Q(g28071) );
  INVX0 U14357 ( .INP(n13576), .ZN(n13575) );
  OR2X1 U14358 ( .IN1(n13577), .IN2(n8186), .Q(n13576) );
  AND2X1 U14359 ( .IN1(n13577), .IN2(g4112), .Q(n13574) );
  AND2X1 U14360 ( .IN1(n8717), .IN2(n13578), .Q(n13577) );
  INVX0 U14361 ( .INP(n13579), .ZN(n13578) );
  AND2X1 U14362 ( .IN1(n13568), .IN2(n5711), .Q(n13579) );
  AND2X1 U14363 ( .IN1(n5416), .IN2(n4722), .Q(n13568) );
  AND4X1 U14364 ( .IN1(n8491), .IN2(n9807), .IN3(n5350), .IN4(n13580), .Q(
        n4722) );
  AND2X1 U14365 ( .IN1(n5612), .IN2(n8348), .Q(n13580) );
  INVX0 U14366 ( .INP(n11746), .ZN(n9807) );
  OR2X1 U14367 ( .IN1(g4087), .IN2(g4093), .Q(n11746) );
  OR4X1 U14368 ( .IN1(n8481), .IN2(n13581), .IN3(n13582), .IN4(n13583), .Q(
        g28070) );
  AND2X1 U14369 ( .IN1(n8821), .IN2(g4082), .Q(n13583) );
  AND3X1 U14370 ( .IN1(test_so11), .IN2(n12862), .IN3(n8732), .Q(n13582) );
  AND2X1 U14371 ( .IN1(n13584), .IN2(n8491), .Q(n13581) );
  INVX0 U14372 ( .INP(n12862), .ZN(n13584) );
  OR2X1 U14373 ( .IN1(n8348), .IN2(n13585), .Q(n12862) );
  OR3X1 U14374 ( .IN1(n13586), .IN2(n13587), .IN3(n13588), .Q(g28069) );
  AND2X1 U14375 ( .IN1(n10689), .IN2(g4035), .Q(n13588) );
  AND2X1 U14376 ( .IN1(n8717), .IN2(n10685), .Q(n10689) );
  AND3X1 U14377 ( .IN1(n10681), .IN2(n12893), .IN3(n8733), .Q(n13587) );
  OR2X1 U14378 ( .IN1(n13589), .IN2(n13590), .Q(n12893) );
  AND2X1 U14379 ( .IN1(n13591), .IN2(g4040), .Q(n13590) );
  OR4X1 U14380 ( .IN1(n13592), .IN2(n13593), .IN3(n13594), .IN4(n13595), .Q(
        n13591) );
  OR3X1 U14381 ( .IN1(n13596), .IN2(n13597), .IN3(n13598), .Q(n13595) );
  AND2X1 U14382 ( .IN1(n9820), .IN2(n13599), .Q(n13598) );
  OR2X1 U14383 ( .IN1(n13600), .IN2(n13601), .Q(n13599) );
  AND2X1 U14384 ( .IN1(test_so65), .IN2(g16748), .Q(n13601) );
  AND2X1 U14385 ( .IN1(g3965), .IN2(g16693), .Q(n13600) );
  AND3X1 U14386 ( .IN1(g3917), .IN2(g16955), .IN3(n10680), .Q(n13597) );
  AND3X1 U14387 ( .IN1(g13906), .IN2(g3933), .IN3(n10684), .Q(n13596) );
  AND2X1 U14388 ( .IN1(n13494), .IN2(n13602), .Q(n13594) );
  OR2X1 U14389 ( .IN1(n13603), .IN2(n13604), .Q(n13602) );
  AND2X1 U14390 ( .IN1(test_so24), .IN2(g14518), .Q(n13604) );
  AND2X1 U14391 ( .IN1(g3897), .IN2(g4031), .Q(n13603) );
  AND2X1 U14392 ( .IN1(n13605), .IN2(g11418), .Q(n13593) );
  OR2X1 U14393 ( .IN1(n13606), .IN2(n13607), .Q(n13605) );
  AND2X1 U14394 ( .IN1(n10680), .IN2(g3893), .Q(n13606) );
  AND2X1 U14395 ( .IN1(n5435), .IN2(n13608), .Q(n13592) );
  AND2X1 U14396 ( .IN1(n5530), .IN2(n13609), .Q(n13589) );
  OR4X1 U14397 ( .IN1(n13610), .IN2(n13611), .IN3(n13612), .IN4(n13613), .Q(
        n13609) );
  OR3X1 U14398 ( .IN1(n13614), .IN2(n13615), .IN3(n13616), .Q(n13613) );
  AND2X1 U14399 ( .IN1(n10684), .IN2(n13617), .Q(n13616) );
  OR2X1 U14400 ( .IN1(n13618), .IN2(n13619), .Q(n13617) );
  AND2X1 U14401 ( .IN1(g3901), .IN2(g14518), .Q(n13619) );
  AND2X1 U14402 ( .IN1(g4031), .IN2(g3913), .Q(n13618) );
  AND3X1 U14403 ( .IN1(g13906), .IN2(g3941), .IN3(n13494), .Q(n13615) );
  AND3X1 U14404 ( .IN1(g16955), .IN2(g3925), .IN3(n9820), .Q(n13614) );
  AND2X1 U14405 ( .IN1(n10680), .IN2(n13620), .Q(n13612) );
  OR2X1 U14406 ( .IN1(n13621), .IN2(n13622), .Q(n13620) );
  AND2X1 U14407 ( .IN1(g3905), .IN2(g16693), .Q(n13622) );
  AND2X1 U14408 ( .IN1(g16748), .IN2(g3957), .Q(n13621) );
  AND2X1 U14409 ( .IN1(n13623), .IN2(g11418), .Q(n13611) );
  OR2X1 U14410 ( .IN1(n13624), .IN2(n13608), .Q(n13623) );
  OR3X1 U14411 ( .IN1(n13625), .IN2(n13626), .IN3(n13627), .Q(n13608) );
  AND3X1 U14412 ( .IN1(g13966), .IN2(g3929), .IN3(n13494), .Q(n13627) );
  AND3X1 U14413 ( .IN1(g3945), .IN2(g16775), .IN3(n10680), .Q(n13626) );
  AND2X1 U14414 ( .IN1(g4054), .IN2(n5594), .Q(n10680) );
  AND3X1 U14415 ( .IN1(g3961), .IN2(g16659), .IN3(n10684), .Q(n13625) );
  AND2X1 U14416 ( .IN1(n9820), .IN2(g3909), .Q(n13624) );
  AND2X1 U14417 ( .IN1(n5435), .IN2(n13607), .Q(n13610) );
  OR3X1 U14418 ( .IN1(n13628), .IN2(n13629), .IN3(n13630), .Q(n13607) );
  AND3X1 U14419 ( .IN1(g3953), .IN2(g16659), .IN3(n13494), .Q(n13630) );
  AND2X1 U14420 ( .IN1(n5395), .IN2(n5594), .Q(n13494) );
  AND3X1 U14421 ( .IN1(g13966), .IN2(g3921), .IN3(n10684), .Q(n13629) );
  AND2X1 U14422 ( .IN1(g3990), .IN2(n5395), .Q(n10684) );
  AND3X1 U14423 ( .IN1(g3937), .IN2(g16775), .IN3(n9820), .Q(n13628) );
  AND2X1 U14424 ( .IN1(g3990), .IN2(g4054), .Q(n9820) );
  INVX0 U14425 ( .INP(n10685), .ZN(n10681) );
  OR2X1 U14426 ( .IN1(n13631), .IN2(n5283), .Q(n10685) );
  AND3X1 U14427 ( .IN1(n13518), .IN2(g4955), .IN3(n9067), .Q(n13631) );
  AND2X1 U14428 ( .IN1(g4899), .IN2(g4975), .Q(n9067) );
  AND2X1 U14429 ( .IN1(n8821), .IN2(g3965), .Q(n13586) );
  OR3X1 U14430 ( .IN1(n13632), .IN2(n13633), .IN3(n13634), .Q(g28066) );
  AND2X1 U14431 ( .IN1(n10705), .IN2(g3684), .Q(n13634) );
  AND2X1 U14432 ( .IN1(n8717), .IN2(n10701), .Q(n10705) );
  AND3X1 U14433 ( .IN1(n10697), .IN2(n12925), .IN3(n8733), .Q(n13633) );
  OR2X1 U14434 ( .IN1(n13635), .IN2(n13636), .Q(n12925) );
  AND2X1 U14435 ( .IN1(n13637), .IN2(g3689), .Q(n13636) );
  OR4X1 U14436 ( .IN1(n13638), .IN2(n13639), .IN3(n13640), .IN4(n13641), .Q(
        n13637) );
  OR3X1 U14437 ( .IN1(n13642), .IN2(n13643), .IN3(n13644), .Q(n13641) );
  AND2X1 U14438 ( .IN1(n9833), .IN2(n13645), .Q(n13644) );
  OR2X1 U14439 ( .IN1(n13646), .IN2(n13647), .Q(n13645) );
  AND2X1 U14440 ( .IN1(g3598), .IN2(g16722), .Q(n13647) );
  AND2X1 U14441 ( .IN1(g3614), .IN2(g16656), .Q(n13646) );
  AND3X1 U14442 ( .IN1(g3566), .IN2(g16924), .IN3(n10696), .Q(n13643) );
  AND3X1 U14443 ( .IN1(n10700), .IN2(g3582), .IN3(test_so26), .Q(n13642) );
  AND2X1 U14444 ( .IN1(n13504), .IN2(n13648), .Q(n13640) );
  OR2X1 U14445 ( .IN1(n13649), .IN2(n13650), .Q(n13648) );
  AND2X1 U14446 ( .IN1(g3538), .IN2(g14451), .Q(n13650) );
  AND2X1 U14447 ( .IN1(g3546), .IN2(g3680), .Q(n13649) );
  AND2X1 U14448 ( .IN1(n13651), .IN2(g11388), .Q(n13639) );
  OR2X1 U14449 ( .IN1(n13652), .IN2(n13653), .Q(n13651) );
  AND2X1 U14450 ( .IN1(n10696), .IN2(g3542), .Q(n13652) );
  AND2X1 U14451 ( .IN1(n5433), .IN2(n13654), .Q(n13638) );
  AND2X1 U14452 ( .IN1(n5532), .IN2(n13655), .Q(n13635) );
  OR4X1 U14453 ( .IN1(n13656), .IN2(n13657), .IN3(n13658), .IN4(n13659), .Q(
        n13655) );
  OR3X1 U14454 ( .IN1(n13660), .IN2(n13661), .IN3(n13662), .Q(n13659) );
  AND2X1 U14455 ( .IN1(n10700), .IN2(n13663), .Q(n13662) );
  OR2X1 U14456 ( .IN1(n13664), .IN2(n13665), .Q(n13663) );
  AND2X1 U14457 ( .IN1(g3550), .IN2(g14451), .Q(n13665) );
  AND2X1 U14458 ( .IN1(g3680), .IN2(g3562), .Q(n13664) );
  AND3X1 U14459 ( .IN1(test_so26), .IN2(g3590), .IN3(n13504), .Q(n13661) );
  AND3X1 U14460 ( .IN1(g16924), .IN2(g3574), .IN3(n9833), .Q(n13660) );
  AND2X1 U14461 ( .IN1(n10696), .IN2(n13666), .Q(n13658) );
  OR2X1 U14462 ( .IN1(n13667), .IN2(n13668), .Q(n13666) );
  AND2X1 U14463 ( .IN1(g3554), .IN2(g16656), .Q(n13668) );
  AND2X1 U14464 ( .IN1(g16722), .IN2(g3606), .Q(n13667) );
  AND2X1 U14465 ( .IN1(n13669), .IN2(g11388), .Q(n13657) );
  OR2X1 U14466 ( .IN1(n13670), .IN2(n13654), .Q(n13669) );
  OR3X1 U14467 ( .IN1(n13671), .IN2(n13672), .IN3(n13673), .Q(n13654) );
  AND3X1 U14468 ( .IN1(g13926), .IN2(g3578), .IN3(n13504), .Q(n13673) );
  AND3X1 U14469 ( .IN1(g3594), .IN2(g16744), .IN3(n10696), .Q(n13672) );
  AND2X1 U14470 ( .IN1(g3703), .IN2(n5591), .Q(n10696) );
  AND3X1 U14471 ( .IN1(g3610), .IN2(g16627), .IN3(n10700), .Q(n13671) );
  AND2X1 U14472 ( .IN1(n9833), .IN2(g3558), .Q(n13670) );
  AND2X1 U14473 ( .IN1(n5433), .IN2(n13653), .Q(n13656) );
  OR3X1 U14474 ( .IN1(n13674), .IN2(n13675), .IN3(n13676), .Q(n13653) );
  AND3X1 U14475 ( .IN1(test_so43), .IN2(g16627), .IN3(n13504), .Q(n13676) );
  AND2X1 U14476 ( .IN1(n5399), .IN2(n5591), .Q(n13504) );
  AND3X1 U14477 ( .IN1(g13926), .IN2(g3570), .IN3(n10700), .Q(n13675) );
  AND2X1 U14478 ( .IN1(g3639), .IN2(n5399), .Q(n10700) );
  AND3X1 U14479 ( .IN1(g3586), .IN2(g16744), .IN3(n9833), .Q(n13674) );
  AND2X1 U14480 ( .IN1(g3639), .IN2(g3703), .Q(n9833) );
  INVX0 U14481 ( .INP(n10701), .ZN(n10697) );
  OR2X1 U14482 ( .IN1(n13677), .IN2(n5443), .Q(n10701) );
  AND3X1 U14483 ( .IN1(n13518), .IN2(g4944), .IN3(n9065), .Q(n13677) );
  AND2X1 U14484 ( .IN1(g4899), .IN2(n5360), .Q(n9065) );
  AND2X1 U14485 ( .IN1(n8821), .IN2(g3614), .Q(n13632) );
  OR3X1 U14486 ( .IN1(n13678), .IN2(n13679), .IN3(n13680), .Q(g28063) );
  AND2X1 U14487 ( .IN1(n10719), .IN2(g3333), .Q(n13680) );
  AND2X1 U14488 ( .IN1(n8717), .IN2(n10713), .Q(n10719) );
  AND3X1 U14489 ( .IN1(n10715), .IN2(n12957), .IN3(n8733), .Q(n13679) );
  OR2X1 U14490 ( .IN1(n13681), .IN2(n13682), .Q(n12957) );
  AND2X1 U14491 ( .IN1(n13683), .IN2(g3338), .Q(n13682) );
  OR4X1 U14492 ( .IN1(n13684), .IN2(n13685), .IN3(n13686), .IN4(n13687), .Q(
        n13683) );
  OR3X1 U14493 ( .IN1(n13688), .IN2(n13689), .IN3(n13690), .Q(n13687) );
  AND2X1 U14494 ( .IN1(n9825), .IN2(n13691), .Q(n13690) );
  OR2X1 U14495 ( .IN1(n13692), .IN2(n13693), .Q(n13691) );
  AND2X1 U14496 ( .IN1(g3247), .IN2(g16686), .Q(n13693) );
  AND2X1 U14497 ( .IN1(g3263), .IN2(g16624), .Q(n13692) );
  AND3X1 U14498 ( .IN1(g3215), .IN2(g16874), .IN3(n10714), .Q(n13689) );
  AND3X1 U14499 ( .IN1(g13865), .IN2(g3231), .IN3(n10712), .Q(n13688) );
  AND2X1 U14500 ( .IN1(n13514), .IN2(n13694), .Q(n13686) );
  OR2X1 U14501 ( .IN1(n13695), .IN2(n13696), .Q(n13694) );
  AND2X1 U14502 ( .IN1(test_so91), .IN2(test_so88), .Q(n13696) );
  AND2X1 U14503 ( .IN1(g3187), .IN2(g14421), .Q(n13695) );
  AND2X1 U14504 ( .IN1(n13697), .IN2(g11349), .Q(n13685) );
  OR2X1 U14505 ( .IN1(n13698), .IN2(n13699), .Q(n13697) );
  AND2X1 U14506 ( .IN1(n10714), .IN2(g3191), .Q(n13698) );
  AND2X1 U14507 ( .IN1(n5436), .IN2(n13700), .Q(n13684) );
  AND2X1 U14508 ( .IN1(n5527), .IN2(n13701), .Q(n13681) );
  OR4X1 U14509 ( .IN1(n13702), .IN2(n13703), .IN3(n13704), .IN4(n13705), .Q(
        n13701) );
  OR3X1 U14510 ( .IN1(n13706), .IN2(n13707), .IN3(n13708), .Q(n13705) );
  AND2X1 U14511 ( .IN1(n10712), .IN2(n13709), .Q(n13708) );
  OR2X1 U14512 ( .IN1(n13710), .IN2(n13711), .Q(n13709) );
  AND2X1 U14513 ( .IN1(g3199), .IN2(g14421), .Q(n13711) );
  AND2X1 U14514 ( .IN1(test_so91), .IN2(g3211), .Q(n13710) );
  AND3X1 U14515 ( .IN1(g13865), .IN2(g3239), .IN3(n13514), .Q(n13707) );
  AND3X1 U14516 ( .IN1(g16874), .IN2(g3223), .IN3(n9825), .Q(n13706) );
  AND2X1 U14517 ( .IN1(n10714), .IN2(n13712), .Q(n13704) );
  OR2X1 U14518 ( .IN1(n13713), .IN2(n13714), .Q(n13712) );
  AND2X1 U14519 ( .IN1(g3203), .IN2(g16624), .Q(n13714) );
  AND2X1 U14520 ( .IN1(g16686), .IN2(g3255), .Q(n13713) );
  AND2X1 U14521 ( .IN1(n13715), .IN2(g11349), .Q(n13703) );
  OR2X1 U14522 ( .IN1(n13716), .IN2(n13700), .Q(n13715) );
  OR3X1 U14523 ( .IN1(n13717), .IN2(n13718), .IN3(n13719), .Q(n13700) );
  AND3X1 U14524 ( .IN1(g13895), .IN2(g3227), .IN3(n13514), .Q(n13719) );
  AND3X1 U14525 ( .IN1(g3243), .IN2(g16718), .IN3(n10714), .Q(n13718) );
  AND2X1 U14526 ( .IN1(g3352), .IN2(n5400), .Q(n10714) );
  AND3X1 U14527 ( .IN1(test_so84), .IN2(g16603), .IN3(n10712), .Q(n13717) );
  AND2X1 U14528 ( .IN1(n9825), .IN2(g3207), .Q(n13716) );
  AND2X1 U14529 ( .IN1(n5436), .IN2(n13699), .Q(n13702) );
  OR3X1 U14530 ( .IN1(n13720), .IN2(n13721), .IN3(n13722), .Q(n13699) );
  AND3X1 U14531 ( .IN1(g3251), .IN2(g16603), .IN3(n13514), .Q(n13722) );
  AND2X1 U14532 ( .IN1(n5604), .IN2(n5400), .Q(n13514) );
  AND3X1 U14533 ( .IN1(g13895), .IN2(g3219), .IN3(n10712), .Q(n13721) );
  AND2X1 U14534 ( .IN1(g3288), .IN2(n5604), .Q(n10712) );
  AND3X1 U14535 ( .IN1(g3235), .IN2(g16718), .IN3(n9825), .Q(n13720) );
  AND2X1 U14536 ( .IN1(g3352), .IN2(g3288), .Q(n9825) );
  INVX0 U14537 ( .INP(n10713), .ZN(n10715) );
  OR2X1 U14538 ( .IN1(n13723), .IN2(n5318), .Q(n10713) );
  AND3X1 U14539 ( .IN1(n13518), .IN2(g4933), .IN3(n9064), .Q(n13723) );
  AND2X1 U14540 ( .IN1(g4975), .IN2(n5517), .Q(n9064) );
  AND3X1 U14541 ( .IN1(n10021), .IN2(n9068), .IN3(n5367), .Q(n13518) );
  AND2X1 U14542 ( .IN1(n8505), .IN2(g4966), .Q(n9068) );
  AND3X1 U14543 ( .IN1(g4849), .IN2(g4843), .IN3(g4859), .Q(n10021) );
  AND2X1 U14544 ( .IN1(n8821), .IN2(g3263), .Q(n13678) );
  OR4X1 U14545 ( .IN1(n2787), .IN2(n13724), .IN3(n13725), .IN4(n13726), .Q(
        g28060) );
  AND2X1 U14546 ( .IN1(n8821), .IN2(g2724), .Q(n13726) );
  AND3X1 U14547 ( .IN1(n13727), .IN2(g2729), .IN3(n8732), .Q(n13725) );
  AND2X1 U14548 ( .IN1(n13728), .IN2(n8347), .Q(n13724) );
  INVX0 U14549 ( .INP(n13727), .ZN(n13728) );
  OR2X1 U14550 ( .IN1(n5301), .IN2(n12376), .Q(n13727) );
  OR3X1 U14551 ( .IN1(n13729), .IN2(n13730), .IN3(n13731), .Q(g28059) );
  AND2X1 U14552 ( .IN1(n8821), .IN2(g1351), .Q(n13731) );
  AND2X1 U14553 ( .IN1(n4798), .IN2(n12640), .Q(n13730) );
  AND3X1 U14554 ( .IN1(n11488), .IN2(n8469), .IN3(n13732), .Q(n13729) );
  AND2X1 U14555 ( .IN1(n8717), .IN2(n11068), .Q(n11488) );
  AND4X1 U14556 ( .IN1(n13733), .IN2(n5466), .IN3(n13734), .IN4(n13735), .Q(
        n11068) );
  INVX0 U14557 ( .INP(n13736), .ZN(n13735) );
  AND3X1 U14558 ( .IN1(n13737), .IN2(g1351), .IN3(n13738), .Q(n13736) );
  OR2X1 U14559 ( .IN1(n13738), .IN2(g1351), .Q(n13734) );
  OR3X1 U14560 ( .IN1(n13739), .IN2(n13740), .IN3(n13741), .Q(g28058) );
  AND2X1 U14561 ( .IN1(test_so77), .IN2(n8808), .Q(n13741) );
  AND2X1 U14562 ( .IN1(n4490), .IN2(n5554), .Q(n13740) );
  AND3X1 U14563 ( .IN1(n11076), .IN2(n13742), .IN3(g1252), .Q(n13739) );
  INVX0 U14564 ( .INP(n4490), .ZN(n13742) );
  OR3X1 U14565 ( .IN1(n13743), .IN2(n13744), .IN3(n13745), .Q(g28057) );
  AND2X1 U14566 ( .IN1(n8821), .IN2(g1008), .Q(n13745) );
  AND2X1 U14567 ( .IN1(n4805), .IN2(n12674), .Q(n13744) );
  AND3X1 U14568 ( .IN1(n11499), .IN2(n8466), .IN3(n13746), .Q(n13743) );
  AND2X1 U14569 ( .IN1(n8717), .IN2(n11083), .Q(n11499) );
  AND4X1 U14570 ( .IN1(n8527), .IN2(n13747), .IN3(n13748), .IN4(n13749), .Q(
        n11083) );
  OR2X1 U14571 ( .IN1(g1008), .IN2(n13750), .Q(n13749) );
  INVX0 U14572 ( .INP(n13751), .ZN(n13748) );
  AND3X1 U14573 ( .IN1(n13752), .IN2(n13750), .IN3(g1008), .Q(n13751) );
  OR3X1 U14574 ( .IN1(n13753), .IN2(n13754), .IN3(n13755), .Q(g28056) );
  AND2X1 U14575 ( .IN1(n8821), .IN2(g936), .Q(n13755) );
  AND2X1 U14576 ( .IN1(n4514), .IN2(n5555), .Q(n13754) );
  AND3X1 U14577 ( .IN1(n11091), .IN2(n13756), .IN3(g907), .Q(n13753) );
  INVX0 U14578 ( .INP(n4514), .ZN(n13756) );
  OR3X1 U14579 ( .IN1(n13757), .IN2(n13758), .IN3(n13759), .Q(g28055) );
  AND2X1 U14580 ( .IN1(n8821), .IN2(g822), .Q(n13759) );
  AND3X1 U14581 ( .IN1(n4519), .IN2(n13200), .IN3(n5728), .Q(n13758) );
  AND3X1 U14582 ( .IN1(n4518), .IN2(n13760), .IN3(g827), .Q(n13757) );
  INVX0 U14583 ( .INP(n4519), .ZN(n13760) );
  OR2X1 U14584 ( .IN1(n13761), .IN2(n13762), .Q(g28054) );
  AND2X1 U14585 ( .IN1(n13763), .IN2(g661), .Q(n13762) );
  AND2X1 U14586 ( .IN1(n13764), .IN2(g728), .Q(n13761) );
  OR3X1 U14587 ( .IN1(n13765), .IN2(n13766), .IN3(n13767), .Q(g28053) );
  AND2X1 U14588 ( .IN1(n8821), .IN2(g681), .Q(n13767) );
  AND2X1 U14589 ( .IN1(n13236), .IN2(test_so87), .Q(n13766) );
  OR2X1 U14590 ( .IN1(n13768), .IN2(n13769), .Q(g28052) );
  AND2X1 U14591 ( .IN1(n13763), .IN2(g718), .Q(n13769) );
  AND2X1 U14592 ( .IN1(n13764), .IN2(g661), .Q(n13768) );
  OR2X1 U14593 ( .IN1(n13770), .IN2(n13771), .Q(g28051) );
  AND2X1 U14594 ( .IN1(n13763), .IN2(g655), .Q(n13771) );
  AND2X1 U14595 ( .IN1(n13764), .IN2(g718), .Q(n13770) );
  OR2X1 U14596 ( .IN1(n13772), .IN2(n13773), .Q(g28050) );
  AND2X1 U14597 ( .IN1(n13763), .IN2(g650), .Q(n13773) );
  AND2X1 U14598 ( .IN1(n13764), .IN2(g655), .Q(n13772) );
  OR3X1 U14599 ( .IN1(n13774), .IN2(n13775), .IN3(n13776), .Q(g28049) );
  AND2X1 U14600 ( .IN1(test_so87), .IN2(n8808), .Q(n13776) );
  AND2X1 U14601 ( .IN1(n13764), .IN2(g650), .Q(n13775) );
  AND2X1 U14602 ( .IN1(n13765), .IN2(g681), .Q(n13774) );
  OR3X1 U14603 ( .IN1(n13777), .IN2(n13778), .IN3(n13779), .Q(g28048) );
  INVX0 U14604 ( .INP(n13780), .ZN(n13779) );
  OR2X1 U14605 ( .IN1(n8679), .IN2(n5657), .Q(n13780) );
  AND2X1 U14606 ( .IN1(n13781), .IN2(n8983), .Q(n13778) );
  AND4X1 U14607 ( .IN1(n5112), .IN2(n5520), .IN3(g703), .IN4(n13218), .Q(n8983) );
  AND4X1 U14608 ( .IN1(test_so87), .IN2(n13782), .IN3(n8316), .IN4(n8317), .Q(
        n13218) );
  XOR2X1 U14609 ( .IN1(n8055), .IN2(g661), .Q(n13782) );
  AND2X1 U14610 ( .IN1(n13783), .IN2(g691), .Q(n13777) );
  OR2X1 U14611 ( .IN1(n13784), .IN2(n13785), .Q(n13783) );
  AND3X1 U14612 ( .IN1(g703), .IN2(n8521), .IN3(n8733), .Q(n13784) );
  OR2X1 U14613 ( .IN1(n13786), .IN2(n13787), .Q(g28047) );
  AND2X1 U14614 ( .IN1(n13763), .IN2(g645), .Q(n13787) );
  INVX0 U14615 ( .INP(n13764), .ZN(n13763) );
  AND2X1 U14616 ( .IN1(n13764), .IN2(g681), .Q(n13786) );
  OR2X1 U14617 ( .IN1(n13788), .IN2(n13789), .Q(g28046) );
  AND2X1 U14618 ( .IN1(n13764), .IN2(g645), .Q(n13789) );
  AND2X1 U14619 ( .IN1(n8717), .IN2(n13790), .Q(n13764) );
  AND2X1 U14620 ( .IN1(n13765), .IN2(g446), .Q(n13788) );
  AND2X1 U14621 ( .IN1(n8717), .IN2(n13791), .Q(n13765) );
  INVX0 U14622 ( .INP(n13790), .ZN(n13791) );
  OR3X1 U14623 ( .IN1(n13792), .IN2(n13793), .IN3(n13794), .Q(n13790) );
  AND2X1 U14624 ( .IN1(n5520), .IN2(n13795), .Q(n13793) );
  OR3X1 U14625 ( .IN1(n5358), .IN2(g411), .IN3(g424), .Q(n13795) );
  AND2X1 U14626 ( .IN1(n13796), .IN2(g691), .Q(n13792) );
  OR3X1 U14627 ( .IN1(n13797), .IN2(n13798), .IN3(n13799), .Q(g28045) );
  AND2X1 U14628 ( .IN1(n8821), .IN2(g568), .Q(n13799) );
  AND2X1 U14629 ( .IN1(n4537), .IN2(n5337), .Q(n13798) );
  AND3X1 U14630 ( .IN1(n2421), .IN2(n13800), .IN3(g572), .Q(n13797) );
  INVX0 U14631 ( .INP(n4537), .ZN(n13800) );
  OR2X1 U14632 ( .IN1(n13801), .IN2(n13802), .Q(g28044) );
  AND2X1 U14633 ( .IN1(n13803), .IN2(n8687), .Q(n13802) );
  OR2X1 U14634 ( .IN1(n4962), .IN2(n13804), .Q(n13803) );
  XOR2X1 U14635 ( .IN1(g482), .IN2(n13232), .Q(n13804) );
  AND2X1 U14636 ( .IN1(n13805), .IN2(n13806), .Q(n13232) );
  OR2X1 U14637 ( .IN1(g528), .IN2(n13807), .Q(n13805) );
  AND2X1 U14638 ( .IN1(n8821), .IN2(g528), .Q(n13801) );
  OR2X1 U14639 ( .IN1(n13808), .IN2(n13809), .Q(g28043) );
  AND2X1 U14640 ( .IN1(n8821), .IN2(g278), .Q(n13809) );
  AND2X1 U14641 ( .IN1(n8473), .IN2(n8515), .Q(n13808) );
  AND2X1 U14642 ( .IN1(n8717), .IN2(n11523), .Q(n8473) );
  AND4X1 U14643 ( .IN1(g691), .IN2(n12692), .IN3(n13810), .IN4(n13811), .Q(
        n11523) );
  OR2X1 U14644 ( .IN1(n13812), .IN2(n5627), .Q(n13810) );
  INVX0 U14645 ( .INP(n13813), .ZN(n13812) );
  OR4X1 U14646 ( .IN1(n13814), .IN2(n13815), .IN3(n13816), .IN4(n13817), .Q(
        n12692) );
  AND3X1 U14647 ( .IN1(n8454), .IN2(n8453), .IN3(n8455), .Q(n13817) );
  AND3X1 U14648 ( .IN1(g753), .IN2(g655), .IN3(g718), .Q(n13816) );
  AND2X1 U14649 ( .IN1(g807), .IN2(g554), .Q(n13814) );
  OR3X1 U14650 ( .IN1(n8792), .IN2(g1306), .IN3(g962), .Q(g28042) );
  OR3X1 U14651 ( .IN1(n8792), .IN2(n11062), .IN3(n10889), .Q(g28041) );
  INVX0 U14652 ( .INP(n9448), .ZN(n10889) );
  OR2X1 U14653 ( .IN1(n7952), .IN2(n13818), .Q(n9448) );
  AND2X1 U14654 ( .IN1(g1193), .IN2(n4837), .Q(n11062) );
  OR2X1 U14655 ( .IN1(n13819), .IN2(n13820), .Q(g28030) );
  AND3X1 U14656 ( .IN1(n9475), .IN2(n9474), .IN3(n9476), .Q(n13820) );
  AND3X1 U14657 ( .IN1(n5861), .IN2(n13821), .IN3(n5882), .Q(n13819) );
  OR2X1 U14658 ( .IN1(n13822), .IN2(n13823), .Q(n13821) );
  AND2X1 U14659 ( .IN1(n9476), .IN2(n9475), .Q(n13823) );
  AND2X1 U14660 ( .IN1(n13824), .IN2(n9474), .Q(n13822) );
  OR2X1 U14661 ( .IN1(n8804), .IN2(n13825), .Q(n9474) );
  AND2X1 U14662 ( .IN1(n5889), .IN2(n5868), .Q(n13825) );
  OR2X1 U14663 ( .IN1(n13826), .IN2(n13827), .Q(n13824) );
  AND2X1 U14664 ( .IN1(n9476), .IN2(n13828), .Q(n13827) );
  OR2X1 U14665 ( .IN1(n13829), .IN2(n13830), .Q(n13828) );
  AND4X1 U14666 ( .IN1(n5885), .IN2(n5869), .IN3(n13831), .IN4(n13832), .Q(
        n13829) );
  OR2X1 U14667 ( .IN1(n13833), .IN2(n13834), .Q(n13832) );
  OR2X1 U14668 ( .IN1(n13835), .IN2(n13836), .Q(n13831) );
  AND2X1 U14669 ( .IN1(n13837), .IN2(n13838), .Q(n9476) );
  AND2X1 U14670 ( .IN1(n9475), .IN2(n13839), .Q(n13826) );
  OR2X1 U14671 ( .IN1(n13838), .IN2(n13837), .Q(n13839) );
  OR2X1 U14672 ( .IN1(n8804), .IN2(n13840), .Q(n13837) );
  AND2X1 U14673 ( .IN1(n5883), .IN2(n5871), .Q(n13840) );
  OR2X1 U14674 ( .IN1(n8804), .IN2(n13841), .Q(n13838) );
  AND2X1 U14675 ( .IN1(n5886), .IN2(n5872), .Q(n13841) );
  AND2X1 U14676 ( .IN1(n13842), .IN2(n13830), .Q(n9475) );
  AND2X1 U14677 ( .IN1(n13834), .IN2(n13833), .Q(n13830) );
  AND2X1 U14678 ( .IN1(n13836), .IN2(n13835), .Q(n13833) );
  INVX0 U14679 ( .INP(n13843), .ZN(n13835) );
  AND2X1 U14680 ( .IN1(n8718), .IN2(n13844), .Q(n13843) );
  OR2X1 U14681 ( .IN1(g5831), .IN2(test_so83), .Q(n13844) );
  OR2X1 U14682 ( .IN1(n8804), .IN2(n13845), .Q(n13836) );
  AND2X1 U14683 ( .IN1(n5888), .IN2(n5874), .Q(n13845) );
  OR2X1 U14684 ( .IN1(n8804), .IN2(n13846), .Q(n13834) );
  AND2X1 U14685 ( .IN1(n5884), .IN2(n5870), .Q(n13846) );
  OR2X1 U14686 ( .IN1(n13847), .IN2(n8793), .Q(n13842) );
  AND2X1 U14687 ( .IN1(n5869), .IN2(n5885), .Q(n13847) );
  OR2X1 U14688 ( .IN1(n13848), .IN2(n13849), .Q(g26971) );
  AND2X1 U14689 ( .IN1(n13850), .IN2(n8687), .Q(n13849) );
  OR2X1 U14690 ( .IN1(n5670), .IN2(n8412), .Q(n13850) );
  AND2X1 U14691 ( .IN1(n8821), .IN2(g4512), .Q(n13848) );
  OR2X1 U14692 ( .IN1(n13851), .IN2(n13852), .Q(g26970) );
  AND2X1 U14693 ( .IN1(n8821), .IN2(g4459), .Q(n13852) );
  AND2X1 U14694 ( .IN1(n8718), .IN2(g4473), .Q(n13851) );
  OR2X1 U14695 ( .IN1(n13853), .IN2(n13854), .Q(g26969) );
  AND3X1 U14696 ( .IN1(n8422), .IN2(n8506), .IN3(n8733), .Q(n13854) );
  AND2X1 U14697 ( .IN1(n8821), .IN2(g4462), .Q(n13853) );
  OR2X1 U14698 ( .IN1(n13855), .IN2(n13856), .Q(g26968) );
  AND2X1 U14699 ( .IN1(n8821), .IN2(g4558), .Q(n13856) );
  OR2X1 U14700 ( .IN1(n13857), .IN2(n13858), .Q(g26967) );
  AND2X1 U14701 ( .IN1(n8821), .IN2(g4561), .Q(n13858) );
  OR2X1 U14702 ( .IN1(n13859), .IN2(n13860), .Q(g26966) );
  AND2X1 U14703 ( .IN1(n8820), .IN2(g4555), .Q(n13860) );
  XOR2X1 U14704 ( .IN1(n9348), .IN2(n13861), .Q(g26965) );
  AND2X1 U14705 ( .IN1(n8718), .IN2(g10306), .Q(n13861) );
  OR2X1 U14706 ( .IN1(n13862), .IN2(n13863), .Q(g26964) );
  INVX0 U14707 ( .INP(n13864), .ZN(n13863) );
  OR2X1 U14708 ( .IN1(n13865), .IN2(n8185), .Q(n13864) );
  AND2X1 U14709 ( .IN1(n8720), .IN2(n13866), .Q(n13865) );
  OR2X1 U14710 ( .IN1(g4521), .IN2(n10053), .Q(n13866) );
  AND3X1 U14711 ( .IN1(n13867), .IN2(n13868), .IN3(n8733), .Q(n13862) );
  OR2X1 U14712 ( .IN1(n5752), .IN2(g4515), .Q(n13868) );
  OR2X1 U14713 ( .IN1(n13869), .IN2(g4521), .Q(n13867) );
  AND2X1 U14714 ( .IN1(n10053), .IN2(n8185), .Q(n13869) );
  AND4X1 U14715 ( .IN1(g4483), .IN2(test_so27), .IN3(g4492), .IN4(g4489), .Q(
        n10053) );
  OR2X1 U14716 ( .IN1(n13857), .IN2(n13870), .Q(g26963) );
  AND2X1 U14717 ( .IN1(n8820), .IN2(g4489), .Q(n13870) );
  AND2X1 U14718 ( .IN1(g6750), .IN2(n8687), .Q(n13857) );
  OR2X1 U14719 ( .IN1(n13871), .IN2(n13855), .Q(g26962) );
  AND2X1 U14720 ( .IN1(g6749), .IN2(n8687), .Q(n13855) );
  AND2X1 U14721 ( .IN1(test_so27), .IN2(n8809), .Q(n13871) );
  OR2X1 U14722 ( .IN1(n13859), .IN2(n13872), .Q(g26961) );
  AND2X1 U14723 ( .IN1(n8820), .IN2(g4483), .Q(n13872) );
  AND2X1 U14724 ( .IN1(g6748), .IN2(n8688), .Q(n13859) );
  OR2X1 U14725 ( .IN1(n13873), .IN2(n13874), .Q(g26958) );
  AND2X1 U14726 ( .IN1(n8820), .IN2(g4455), .Q(n13873) );
  OR2X1 U14727 ( .IN1(n13875), .IN2(n13876), .Q(g26957) );
  AND2X1 U14728 ( .IN1(test_so47), .IN2(n8688), .Q(n13876) );
  AND2X1 U14729 ( .IN1(n13877), .IN2(g4434), .Q(n13875) );
  OR2X1 U14730 ( .IN1(n8795), .IN2(n13878), .Q(n13877) );
  AND2X1 U14731 ( .IN1(n13879), .IN2(g4392), .Q(n13878) );
  OR2X1 U14732 ( .IN1(n13880), .IN2(n9336), .Q(g26956) );
  AND3X1 U14733 ( .IN1(n13879), .IN2(g4430), .IN3(n13881), .Q(n13880) );
  OR2X1 U14734 ( .IN1(n13882), .IN2(n13883), .Q(g26955) );
  AND2X1 U14735 ( .IN1(n13884), .IN2(g4438), .Q(n13883) );
  AND2X1 U14736 ( .IN1(n13879), .IN2(n13885), .Q(n13882) );
  OR3X1 U14737 ( .IN1(n13886), .IN2(n13887), .IN3(n13888), .Q(g26954) );
  AND2X1 U14738 ( .IN1(test_so47), .IN2(n8808), .Q(n13888) );
  AND2X1 U14739 ( .IN1(n13889), .IN2(g4438), .Q(n13887) );
  AND2X1 U14740 ( .IN1(n13881), .IN2(n13879), .Q(n13886) );
  INVX0 U14741 ( .INP(n13890), .ZN(n13879) );
  OR4X1 U14742 ( .IN1(test_so47), .IN2(g4438), .IN3(n9336), .IN4(n13891), .Q(
        n13890) );
  OR2X1 U14743 ( .IN1(g7245), .IN2(g7260), .Q(n13891) );
  OR2X1 U14744 ( .IN1(n13892), .IN2(n13893), .Q(g26952) );
  AND2X1 U14745 ( .IN1(n13894), .IN2(n8688), .Q(n13893) );
  OR2X1 U14746 ( .IN1(n13895), .IN2(n13896), .Q(n13894) );
  XOR2X1 U14747 ( .IN1(n8016), .IN2(n8015), .Q(n13896) );
  AND2X1 U14748 ( .IN1(n8398), .IN2(g4388), .Q(n13895) );
  AND2X1 U14749 ( .IN1(n13897), .IN2(g4430), .Q(n13892) );
  OR2X1 U14750 ( .IN1(n8401), .IN2(n8793), .Q(n13897) );
  OR2X1 U14751 ( .IN1(n13898), .IN2(g26953), .Q(g26951) );
  AND2X1 U14752 ( .IN1(n8820), .IN2(g4427), .Q(n13898) );
  OR2X1 U14753 ( .IN1(n13899), .IN2(n13874), .Q(g26950) );
  OR2X1 U14754 ( .IN1(n13900), .IN2(n13901), .Q(n13874) );
  AND2X1 U14755 ( .IN1(n13902), .IN2(n8688), .Q(n13901) );
  AND2X1 U14756 ( .IN1(n13885), .IN2(n13903), .Q(n13900) );
  AND2X1 U14757 ( .IN1(n8820), .IN2(g4417), .Q(n13899) );
  OR2X1 U14758 ( .IN1(n13904), .IN2(n13905), .Q(g26949) );
  AND2X1 U14759 ( .IN1(n8720), .IN2(g4411), .Q(n13905) );
  AND2X1 U14760 ( .IN1(n13906), .IN2(g4401), .Q(n13904) );
  OR2X1 U14761 ( .IN1(n8797), .IN2(n13907), .Q(n13906) );
  AND2X1 U14762 ( .IN1(n13908), .IN2(g4392), .Q(n13907) );
  OR2X1 U14763 ( .IN1(n13909), .IN2(g4405), .Q(g26948) );
  AND3X1 U14764 ( .IN1(n13908), .IN2(g4388), .IN3(n13881), .Q(n13909) );
  OR3X1 U14765 ( .IN1(n13910), .IN2(n13911), .IN3(n13912), .Q(g26947) );
  AND2X1 U14766 ( .IN1(n13913), .IN2(n8688), .Q(n13911) );
  OR2X1 U14767 ( .IN1(n13914), .IN2(n13902), .Q(n13913) );
  AND3X1 U14768 ( .IN1(n13908), .IN2(n5710), .IN3(n8460), .Q(n13902) );
  AND3X1 U14769 ( .IN1(n13903), .IN2(g4382), .IN3(n7950), .Q(n13914) );
  AND2X1 U14770 ( .IN1(n8820), .IN2(g4388), .Q(n13910) );
  OR2X1 U14771 ( .IN1(n13915), .IN2(n13916), .Q(g26946) );
  AND2X1 U14772 ( .IN1(n13884), .IN2(g4375), .Q(n13916) );
  AND2X1 U14773 ( .IN1(n13908), .IN2(n13885), .Q(n13915) );
  AND2X1 U14774 ( .IN1(g4392), .IN2(n8688), .Q(n13885) );
  OR3X1 U14775 ( .IN1(n13917), .IN2(n13912), .IN3(n13918), .Q(g26945) );
  AND2X1 U14776 ( .IN1(n8820), .IN2(g4411), .Q(n13918) );
  AND2X1 U14777 ( .IN1(n13889), .IN2(g4375), .Q(n13912) );
  INVX0 U14778 ( .INP(n13884), .ZN(n13889) );
  OR2X1 U14779 ( .IN1(n8799), .IN2(g4382), .Q(n13884) );
  AND2X1 U14780 ( .IN1(n13881), .IN2(n13908), .Q(n13917) );
  INVX0 U14781 ( .INP(n13903), .ZN(n13908) );
  OR4X1 U14782 ( .IN1(g4405), .IN2(g4375), .IN3(g4411), .IN4(n13919), .Q(
        n13903) );
  OR2X1 U14783 ( .IN1(g7257), .IN2(g7243), .Q(n13919) );
  AND2X1 U14784 ( .IN1(n8721), .IN2(n5710), .Q(n13881) );
  AND2X1 U14785 ( .IN1(n13920), .IN2(n8688), .Q(g26944) );
  INVX0 U14786 ( .INP(n13921), .ZN(n13920) );
  AND4X1 U14787 ( .IN1(n9390), .IN2(n13922), .IN3(g4358), .IN4(test_so81), .Q(
        n13921) );
  INVX0 U14788 ( .INP(n13923), .ZN(n9390) );
  OR2X1 U14789 ( .IN1(n13924), .IN2(g135), .Q(n13923) );
  AND3X1 U14790 ( .IN1(n13925), .IN2(n13926), .IN3(n13927), .Q(n13924) );
  OR3X1 U14791 ( .IN1(g4616), .IN2(n13928), .IN3(n13929), .Q(n13927) );
  XOR2X1 U14792 ( .IN1(n5539), .IN2(n5274), .Q(n13929) );
  XOR2X1 U14793 ( .IN1(n5365), .IN2(n5303), .Q(n13928) );
  OR4X1 U14794 ( .IN1(n5303), .IN2(g4601), .IN3(g4608), .IN4(n5539), .Q(n13926) );
  OR3X1 U14795 ( .IN1(n5274), .IN2(g4593), .IN3(g4584), .Q(n13925) );
  OR2X1 U14796 ( .IN1(n13930), .IN2(n13931), .Q(g26940) );
  AND2X1 U14797 ( .IN1(n12099), .IN2(n8688), .Q(n13931) );
  OR2X1 U14798 ( .IN1(n13932), .IN2(n13933), .Q(n12099) );
  AND2X1 U14799 ( .IN1(g114), .IN2(n5983), .Q(n13933) );
  AND2X1 U14800 ( .IN1(g116), .IN2(g4157), .Q(n13932) );
  AND2X1 U14801 ( .IN1(n8820), .IN2(g4153), .Q(n13930) );
  OR2X1 U14802 ( .IN1(n13934), .IN2(n13935), .Q(g26939) );
  AND2X1 U14803 ( .IN1(n12101), .IN2(n8688), .Q(n13935) );
  OR2X1 U14804 ( .IN1(n13936), .IN2(n13937), .Q(n12101) );
  AND2X1 U14805 ( .IN1(g120), .IN2(n5981), .Q(n13937) );
  AND2X1 U14806 ( .IN1(g124), .IN2(g4146), .Q(n13936) );
  AND2X1 U14807 ( .IN1(n8820), .IN2(g4104), .Q(n13934) );
  OR3X1 U14808 ( .IN1(n13938), .IN2(n13939), .IN3(n8481), .Q(g26938) );
  AND2X1 U14809 ( .IN1(n13940), .IN2(n8688), .Q(n13939) );
  XOR2X1 U14810 ( .IN1(n13585), .IN2(n8348), .Q(n13940) );
  OR2X1 U14811 ( .IN1(n5612), .IN2(n1166), .Q(n13585) );
  AND2X1 U14812 ( .IN1(n8820), .IN2(g4141), .Q(n13938) );
  OR3X1 U14813 ( .IN1(n13941), .IN2(n13942), .IN3(n13943), .Q(g26934) );
  AND2X1 U14814 ( .IN1(n4888), .IN2(g2827), .Q(n13943) );
  AND2X1 U14815 ( .IN1(test_so37), .IN2(n8808), .Q(n13942) );
  AND2X1 U14816 ( .IN1(n13944), .IN2(n8525), .Q(n13941) );
  OR3X1 U14817 ( .IN1(n13945), .IN2(n13946), .IN3(n13947), .Q(g26933) );
  AND2X1 U14818 ( .IN1(test_so37), .IN2(n4888), .Q(n13947) );
  AND2X1 U14819 ( .IN1(n8820), .IN2(g2811), .Q(n13946) );
  AND2X1 U14820 ( .IN1(n5840), .IN2(n13944), .Q(n13945) );
  OR3X1 U14821 ( .IN1(n13948), .IN2(n13949), .IN3(n13950), .Q(g26932) );
  AND2X1 U14822 ( .IN1(n4888), .IN2(g2811), .Q(n13950) );
  AND2X1 U14823 ( .IN1(n8820), .IN2(g2799), .Q(n13949) );
  AND2X1 U14824 ( .IN1(n5841), .IN2(n13944), .Q(n13948) );
  OR3X1 U14825 ( .IN1(n13951), .IN2(n13952), .IN3(n13953), .Q(g26931) );
  AND2X1 U14826 ( .IN1(n4888), .IN2(g2799), .Q(n13953) );
  AND2X1 U14827 ( .IN1(n8820), .IN2(g29219), .Q(n13952) );
  AND2X1 U14828 ( .IN1(n5839), .IN2(n13944), .Q(n13951) );
  OR3X1 U14829 ( .IN1(n13954), .IN2(n13955), .IN3(n13956), .Q(g26930) );
  AND2X1 U14830 ( .IN1(n4888), .IN2(g2795), .Q(n13956) );
  AND2X1 U14831 ( .IN1(n8820), .IN2(g2791), .Q(n13955) );
  AND2X1 U14832 ( .IN1(n13944), .IN2(n8526), .Q(n13954) );
  OR3X1 U14833 ( .IN1(n13957), .IN2(n13958), .IN3(n13959), .Q(g26929) );
  AND2X1 U14834 ( .IN1(n4888), .IN2(g2791), .Q(n13959) );
  AND2X1 U14835 ( .IN1(n8820), .IN2(g2779), .Q(n13958) );
  AND2X1 U14836 ( .IN1(n5837), .IN2(n13944), .Q(n13957) );
  OR3X1 U14837 ( .IN1(n13960), .IN2(n13961), .IN3(n13962), .Q(g26928) );
  AND2X1 U14838 ( .IN1(n4888), .IN2(g2779), .Q(n13962) );
  AND2X1 U14839 ( .IN1(n8820), .IN2(g2767), .Q(n13961) );
  AND2X1 U14840 ( .IN1(n5834), .IN2(n13944), .Q(n13960) );
  OR3X1 U14841 ( .IN1(n13963), .IN2(n13964), .IN3(n13965), .Q(g26927) );
  AND2X1 U14842 ( .IN1(n4888), .IN2(g2767), .Q(n13965) );
  AND2X1 U14843 ( .IN1(n8820), .IN2(g2763), .Q(n13964) );
  AND2X1 U14844 ( .IN1(n5836), .IN2(n13944), .Q(n13963) );
  AND3X1 U14845 ( .IN1(n9768), .IN2(n9081), .IN3(n4888), .Q(n13944) );
  OR2X1 U14846 ( .IN1(test_so30), .IN2(g2748), .Q(n9081) );
  INVX0 U14847 ( .INP(n9774), .ZN(n9768) );
  AND3X1 U14848 ( .IN1(g2735), .IN2(n3505), .IN3(test_so30), .Q(n9774) );
  AND2X1 U14849 ( .IN1(g2748), .IN2(g2741), .Q(n3505) );
  OR2X1 U14850 ( .IN1(n13966), .IN2(n13967), .Q(g26926) );
  AND2X1 U14851 ( .IN1(n8820), .IN2(g2719), .Q(n13967) );
  AND2X1 U14852 ( .IN1(n13968), .IN2(n3730), .Q(n13966) );
  XOR2X1 U14853 ( .IN1(n12376), .IN2(n5301), .Q(n13968) );
  OR2X1 U14854 ( .IN1(n5465), .IN2(n5299), .Q(n12376) );
  OR2X1 U14855 ( .IN1(n13969), .IN2(n13970), .Q(g26925) );
  AND2X1 U14856 ( .IN1(n13971), .IN2(n8689), .Q(n13970) );
  OR2X1 U14857 ( .IN1(n13972), .IN2(n4173), .Q(n13971) );
  AND2X1 U14858 ( .IN1(n12615), .IN2(g1536), .Q(n13972) );
  OR2X1 U14859 ( .IN1(n8461), .IN2(n12618), .Q(n12615) );
  OR2X1 U14860 ( .IN1(n8051), .IN2(n12625), .Q(n12618) );
  OR3X1 U14861 ( .IN1(n5302), .IN2(n12635), .IN3(n12634), .Q(n12625) );
  AND3X1 U14862 ( .IN1(g1521), .IN2(g1339), .IN3(n8244), .Q(n12635) );
  AND2X1 U14863 ( .IN1(n8820), .IN2(g1532), .Q(n13969) );
  OR3X1 U14864 ( .IN1(n13973), .IN2(n13974), .IN3(n13975), .Q(g26924) );
  AND2X1 U14865 ( .IN1(n13976), .IN2(n5289), .Q(n13975) );
  AND2X1 U14866 ( .IN1(n8820), .IN2(g1437), .Q(n13974) );
  AND3X1 U14867 ( .IN1(n13977), .IN2(g1478), .IN3(n8733), .Q(n13973) );
  INVX0 U14868 ( .INP(n13976), .ZN(n13977) );
  AND3X1 U14869 ( .IN1(g1437), .IN2(n13155), .IN3(n13978), .Q(n13976) );
  AND3X1 U14870 ( .IN1(n8490), .IN2(g13272), .IN3(g1514), .Q(n13155) );
  OR3X1 U14871 ( .IN1(n13979), .IN2(n13980), .IN3(n13981), .Q(g26923) );
  AND2X1 U14872 ( .IN1(n13982), .IN2(n5290), .Q(n13981) );
  AND2X1 U14873 ( .IN1(n8820), .IN2(g1467), .Q(n13980) );
  AND3X1 U14874 ( .IN1(n13983), .IN2(g1472), .IN3(n8733), .Q(n13979) );
  INVX0 U14875 ( .INP(n13982), .ZN(n13983) );
  AND3X1 U14876 ( .IN1(g1467), .IN2(n13148), .IN3(n13978), .Q(n13982) );
  AND2X1 U14877 ( .IN1(g13272), .IN2(n10805), .Q(n13148) );
  OR3X1 U14878 ( .IN1(n13984), .IN2(n13985), .IN3(n13986), .Q(g26922) );
  AND2X1 U14879 ( .IN1(n13987), .IN2(n5343), .Q(n13986) );
  AND2X1 U14880 ( .IN1(n8819), .IN2(g1454), .Q(n13985) );
  AND3X1 U14881 ( .IN1(n13988), .IN2(g1448), .IN3(n8733), .Q(n13984) );
  INVX0 U14882 ( .INP(n13987), .ZN(n13988) );
  AND3X1 U14883 ( .IN1(g1454), .IN2(n13131), .IN3(n13978), .Q(n13987) );
  INVX0 U14884 ( .INP(n13134), .ZN(n13131) );
  OR2X1 U14885 ( .IN1(n8411), .IN2(n12634), .Q(n13134) );
  OR2X1 U14886 ( .IN1(g1514), .IN2(n8490), .Q(n12634) );
  OR2X1 U14887 ( .IN1(n13989), .IN2(n13990), .Q(g26921) );
  AND3X1 U14888 ( .IN1(n13991), .IN2(n8496), .IN3(n8734), .Q(n13990) );
  XOR2X1 U14889 ( .IN1(n13992), .IN2(n8427), .Q(n13991) );
  AND2X1 U14890 ( .IN1(n8819), .IN2(g1395), .Q(n13989) );
  OR3X1 U14891 ( .IN1(n13993), .IN2(n13994), .IN3(n13995), .Q(g26920) );
  AND2X1 U14892 ( .IN1(n4913), .IN2(n13996), .Q(n13995) );
  AND3X1 U14893 ( .IN1(n9105), .IN2(g1389), .IN3(n8733), .Q(n13994) );
  OR2X1 U14894 ( .IN1(n13997), .IN2(n13998), .Q(n9105) );
  AND2X1 U14895 ( .IN1(n8434), .IN2(g1351), .Q(n13997) );
  AND2X1 U14896 ( .IN1(n8819), .IN2(g1384), .Q(n13993) );
  OR3X1 U14897 ( .IN1(n13999), .IN2(n14000), .IN3(n14001), .Q(g26919) );
  AND2X1 U14898 ( .IN1(n8819), .IN2(g1266), .Q(n14001) );
  AND2X1 U14899 ( .IN1(n4804), .IN2(n5556), .Q(n14000) );
  AND3X1 U14900 ( .IN1(test_so77), .IN2(n11076), .IN3(n14002), .Q(n13999) );
  INVX0 U14901 ( .INP(n4804), .ZN(n14002) );
  AND3X1 U14902 ( .IN1(g1249), .IN2(g1266), .IN3(g12923), .Q(n4804) );
  OR2X1 U14903 ( .IN1(n14003), .IN2(n14004), .Q(g26918) );
  AND2X1 U14904 ( .IN1(n14005), .IN2(n8689), .Q(n14004) );
  OR2X1 U14905 ( .IN1(n14006), .IN2(n4191), .Q(n14005) );
  AND2X1 U14906 ( .IN1(n12649), .IN2(g1193), .Q(n14006) );
  OR2X1 U14907 ( .IN1(n8462), .IN2(n12652), .Q(n12649) );
  OR2X1 U14908 ( .IN1(n8052), .IN2(n12659), .Q(n12652) );
  OR3X1 U14909 ( .IN1(n5304), .IN2(n12669), .IN3(n12668), .Q(n12659) );
  AND3X1 U14910 ( .IN1(g996), .IN2(g1178), .IN3(n5642), .Q(n12669) );
  AND2X1 U14911 ( .IN1(n8819), .IN2(g1189), .Q(n14003) );
  OR3X1 U14912 ( .IN1(n14007), .IN2(n14008), .IN3(n14009), .Q(g26917) );
  AND2X1 U14913 ( .IN1(n14010), .IN2(n5328), .Q(n14009) );
  AND2X1 U14914 ( .IN1(n8819), .IN2(g1094), .Q(n14008) );
  AND3X1 U14915 ( .IN1(n14011), .IN2(g1135), .IN3(n8733), .Q(n14007) );
  INVX0 U14916 ( .INP(n14010), .ZN(n14011) );
  AND3X1 U14917 ( .IN1(g1094), .IN2(n13190), .IN3(n14012), .Q(n14010) );
  AND3X1 U14918 ( .IN1(g13259), .IN2(g1171), .IN3(n5599), .Q(n13190) );
  OR3X1 U14919 ( .IN1(n14013), .IN2(n14014), .IN3(n14015), .Q(g26916) );
  AND2X1 U14920 ( .IN1(n14016), .IN2(n5329), .Q(n14015) );
  AND2X1 U14921 ( .IN1(n8819), .IN2(g1124), .Q(n14014) );
  AND3X1 U14922 ( .IN1(n14017), .IN2(g1129), .IN3(n8734), .Q(n14013) );
  INVX0 U14923 ( .INP(n14016), .ZN(n14017) );
  AND3X1 U14924 ( .IN1(g1124), .IN2(n13183), .IN3(n14012), .Q(n14016) );
  AND3X1 U14925 ( .IN1(g13259), .IN2(g1183), .IN3(g1171), .Q(n13183) );
  OR3X1 U14926 ( .IN1(n14018), .IN2(n14019), .IN3(n14020), .Q(g26915) );
  AND2X1 U14927 ( .IN1(n14021), .IN2(n5478), .Q(n14020) );
  AND2X1 U14928 ( .IN1(test_so90), .IN2(n8809), .Q(n14019) );
  AND3X1 U14929 ( .IN1(n14022), .IN2(g1105), .IN3(n8734), .Q(n14018) );
  INVX0 U14930 ( .INP(n14021), .ZN(n14022) );
  AND3X1 U14931 ( .IN1(n13166), .IN2(test_so90), .IN3(n14012), .Q(n14021) );
  INVX0 U14932 ( .INP(n13169), .ZN(n13166) );
  OR2X1 U14933 ( .IN1(n8418), .IN2(n12668), .Q(n13169) );
  OR2X1 U14934 ( .IN1(n5599), .IN2(g1171), .Q(n12668) );
  OR2X1 U14935 ( .IN1(n14023), .IN2(n14024), .Q(g26914) );
  AND3X1 U14936 ( .IN1(n5320), .IN2(n14025), .IN3(n8734), .Q(n14024) );
  XOR2X1 U14937 ( .IN1(n14026), .IN2(n8426), .Q(n14025) );
  AND2X1 U14938 ( .IN1(n8819), .IN2(g1052), .Q(n14023) );
  OR3X1 U14939 ( .IN1(n14027), .IN2(n14028), .IN3(n14029), .Q(g26913) );
  AND2X1 U14940 ( .IN1(n4938), .IN2(n14030), .Q(n14029) );
  AND3X1 U14941 ( .IN1(n8987), .IN2(g1046), .IN3(n8734), .Q(n14028) );
  OR2X1 U14942 ( .IN1(n14031), .IN2(n14032), .Q(n8987) );
  AND2X1 U14943 ( .IN1(n8435), .IN2(g1008), .Q(n14031) );
  AND2X1 U14944 ( .IN1(n8819), .IN2(g1041), .Q(n14027) );
  OR3X1 U14945 ( .IN1(n14033), .IN2(n14034), .IN3(n14035), .Q(g26912) );
  AND2X1 U14946 ( .IN1(n8819), .IN2(g921), .Q(n14035) );
  AND2X1 U14947 ( .IN1(n4811), .IN2(n5557), .Q(n14034) );
  AND3X1 U14948 ( .IN1(n11091), .IN2(n14036), .IN3(g936), .Q(n14033) );
  INVX0 U14949 ( .INP(n4811), .ZN(n14036) );
  AND3X1 U14950 ( .IN1(g904), .IN2(g921), .IN3(g12919), .Q(n4811) );
  XOR2X1 U14951 ( .IN1(g862), .IN2(n14037), .Q(g26910) );
  AND2X1 U14952 ( .IN1(n5305), .IN2(n8689), .Q(n14037) );
  OR2X1 U14953 ( .IN1(n14038), .IN2(n14039), .Q(g26909) );
  AND2X1 U14954 ( .IN1(n14040), .IN2(n8689), .Q(n14039) );
  OR2X1 U14955 ( .IN1(n14041), .IN2(n14042), .Q(n14040) );
  AND2X1 U14956 ( .IN1(n5305), .IN2(g896), .Q(n14042) );
  AND2X1 U14957 ( .IN1(n5431), .IN2(g862), .Q(n14041) );
  AND2X1 U14958 ( .IN1(n8819), .IN2(g890), .Q(n14038) );
  OR3X1 U14959 ( .IN1(n14043), .IN2(n14044), .IN3(n14045), .Q(g26908) );
  AND2X1 U14960 ( .IN1(n4945), .IN2(g446), .Q(n14045) );
  AND2X1 U14961 ( .IN1(n8819), .IN2(g246), .Q(n14044) );
  AND2X1 U14962 ( .IN1(n14046), .IN2(g872), .Q(n14043) );
  OR3X1 U14963 ( .IN1(n14047), .IN2(n14048), .IN3(n14049), .Q(g26907) );
  AND2X1 U14964 ( .IN1(n4945), .IN2(g246), .Q(n14049) );
  AND2X1 U14965 ( .IN1(n8819), .IN2(g269), .Q(n14048) );
  AND2X1 U14966 ( .IN1(n14046), .IN2(g14167), .Q(n14047) );
  OR3X1 U14967 ( .IN1(n14050), .IN2(n14051), .IN3(n14052), .Q(g26906) );
  AND2X1 U14968 ( .IN1(n4945), .IN2(g269), .Q(n14052) );
  AND2X1 U14969 ( .IN1(n8819), .IN2(g239), .Q(n14051) );
  AND2X1 U14970 ( .IN1(n14046), .IN2(g14147), .Q(n14050) );
  OR3X1 U14971 ( .IN1(n14053), .IN2(n14054), .IN3(n14055), .Q(g26905) );
  AND2X1 U14972 ( .IN1(n4945), .IN2(g239), .Q(n14055) );
  AND2X1 U14973 ( .IN1(n8819), .IN2(g262), .Q(n14054) );
  AND2X1 U14974 ( .IN1(n14046), .IN2(g14125), .Q(n14053) );
  OR3X1 U14975 ( .IN1(n14056), .IN2(n14057), .IN3(n14058), .Q(g26904) );
  AND2X1 U14976 ( .IN1(n4945), .IN2(g262), .Q(n14058) );
  AND2X1 U14977 ( .IN1(n8819), .IN2(g232), .Q(n14057) );
  AND2X1 U14978 ( .IN1(n14046), .IN2(g14096), .Q(n14056) );
  OR3X1 U14979 ( .IN1(n14059), .IN2(n14060), .IN3(n14061), .Q(g26903) );
  AND2X1 U14980 ( .IN1(n4945), .IN2(g232), .Q(n14061) );
  AND2X1 U14981 ( .IN1(n8819), .IN2(g255), .Q(n14060) );
  AND2X1 U14982 ( .IN1(n14046), .IN2(g14217), .Q(n14059) );
  OR3X1 U14983 ( .IN1(n14062), .IN2(n14063), .IN3(n14064), .Q(g26902) );
  AND2X1 U14984 ( .IN1(n4945), .IN2(g255), .Q(n14064) );
  AND2X1 U14985 ( .IN1(n8819), .IN2(g225), .Q(n14063) );
  AND2X1 U14986 ( .IN1(n14046), .IN2(g14201), .Q(n14062) );
  OR3X1 U14987 ( .IN1(n14065), .IN2(n14066), .IN3(n14067), .Q(g26901) );
  AND2X1 U14988 ( .IN1(n4945), .IN2(g225), .Q(n14067) );
  AND2X1 U14989 ( .IN1(n8819), .IN2(g872), .Q(n14066) );
  AND2X1 U14990 ( .IN1(n14046), .IN2(g14189), .Q(n14065) );
  AND2X1 U14991 ( .IN1(n8982), .IN2(n8689), .Q(n14046) );
  AND3X1 U14992 ( .IN1(g890), .IN2(n5431), .IN3(n5682), .Q(n8982) );
  OR2X1 U14993 ( .IN1(n14068), .IN2(n14069), .Q(g26899) );
  AND2X1 U14994 ( .IN1(n8819), .IN2(g832), .Q(n14069) );
  AND2X1 U14995 ( .IN1(n14070), .IN2(n4518), .Q(n14068) );
  XOR2X1 U14996 ( .IN1(g822), .IN2(n4814), .Q(n14070) );
  AND3X1 U14997 ( .IN1(g832), .IN2(g817), .IN3(n4948), .Q(n4814) );
  OR2X1 U14998 ( .IN1(n14071), .IN2(n14072), .Q(g26898) );
  AND2X1 U14999 ( .IN1(n14073), .IN2(g843), .Q(n14072) );
  OR2X1 U15000 ( .IN1(n8800), .IN2(n14074), .Q(n14073) );
  AND3X1 U15001 ( .IN1(n5733), .IN2(g837), .IN3(n14075), .Q(n14074) );
  AND3X1 U15002 ( .IN1(g837), .IN2(g812), .IN3(n14076), .Q(n14071) );
  OR2X1 U15003 ( .IN1(n14077), .IN2(n13236), .Q(n14076) );
  AND2X1 U15004 ( .IN1(n14078), .IN2(n8689), .Q(n14077) );
  OR2X1 U15005 ( .IN1(n5709), .IN2(n8029), .Q(n14078) );
  OR2X1 U15006 ( .IN1(n14079), .IN2(n14080), .Q(g26897) );
  AND2X1 U15007 ( .IN1(n14081), .IN2(g732), .Q(n14080) );
  INVX0 U15008 ( .INP(n14082), .ZN(n14081) );
  AND2X1 U15009 ( .IN1(n14082), .IN2(g753), .Q(n14079) );
  AND2X1 U15010 ( .IN1(n8721), .IN2(n13815), .Q(n14082) );
  OR3X1 U15011 ( .IN1(n14083), .IN2(n14084), .IN3(n14085), .Q(g26896) );
  AND2X1 U15012 ( .IN1(n4956), .IN2(n13219), .Q(n14085) );
  AND2X1 U15013 ( .IN1(n14086), .IN2(g728), .Q(n14084) );
  INVX0 U15014 ( .INP(n14087), .ZN(n14083) );
  OR2X1 U15015 ( .IN1(n14086), .IN2(n5657), .Q(n14087) );
  OR2X1 U15016 ( .IN1(n8800), .IN2(n13219), .Q(n14086) );
  AND4X1 U15017 ( .IN1(n13807), .IN2(test_so54), .IN3(n5519), .IN4(n4948), .Q(
        n13219) );
  OR3X1 U15018 ( .IN1(n14088), .IN2(n14089), .IN3(n14090), .Q(g26895) );
  AND2X1 U15019 ( .IN1(n8819), .IN2(g562), .Q(n14090) );
  AND2X1 U15020 ( .IN1(n4826), .IN2(n5335), .Q(n14089) );
  AND3X1 U15021 ( .IN1(n2421), .IN2(n14091), .IN3(g568), .Q(n14088) );
  INVX0 U15022 ( .INP(n4826), .ZN(n14091) );
  AND3X1 U15023 ( .IN1(n14092), .IN2(g562), .IN3(n4959), .Q(n4826) );
  OR2X1 U15024 ( .IN1(n14093), .IN2(n14094), .Q(g26894) );
  AND4X1 U15025 ( .IN1(n14095), .IN2(n14096), .IN3(n13231), .IN4(n8723), .Q(
        n14094) );
  INVX0 U15026 ( .INP(n14097), .ZN(n14096) );
  AND2X1 U15027 ( .IN1(g528), .IN2(n13806), .Q(n14097) );
  OR2X1 U15028 ( .IN1(n14098), .IN2(g528), .Q(n14095) );
  AND2X1 U15029 ( .IN1(n13806), .IN2(n14099), .Q(n14098) );
  INVX0 U15030 ( .INP(n13807), .ZN(n14099) );
  AND3X1 U15031 ( .IN1(g482), .IN2(g490), .IN3(n5327), .Q(n13807) );
  AND3X1 U15032 ( .IN1(g518), .IN2(n5548), .IN3(n14100), .Q(n13806) );
  AND2X1 U15033 ( .IN1(n8819), .IN2(g518), .Q(n14093) );
  OR2X1 U15034 ( .IN1(n14101), .IN2(n14102), .Q(g26893) );
  AND2X1 U15035 ( .IN1(n14103), .IN2(n8689), .Q(n14102) );
  OR2X1 U15036 ( .IN1(n14104), .IN2(n14105), .Q(n14103) );
  AND2X1 U15037 ( .IN1(test_so17), .IN2(n14106), .Q(n14105) );
  AND2X1 U15038 ( .IN1(g29211), .IN2(n8513), .Q(n14104) );
  AND2X1 U15039 ( .IN1(n8818), .IN2(g355), .Q(n14101) );
  OR2X1 U15040 ( .IN1(n14107), .IN2(n14108), .Q(g26892) );
  AND2X1 U15041 ( .IN1(test_so17), .IN2(n8809), .Q(n14108) );
  AND3X1 U15042 ( .IN1(n8726), .IN2(n14106), .IN3(n8513), .Q(n14107) );
  OR2X1 U15043 ( .IN1(g333), .IN2(g355), .Q(n14106) );
  OR2X1 U15044 ( .IN1(n14109), .IN2(n14110), .Q(g26891) );
  AND3X1 U15045 ( .IN1(n8727), .IN2(g7540), .IN3(n5860), .Q(n14110) );
  AND2X1 U15046 ( .IN1(n8818), .IN2(g347), .Q(n14109) );
  OR2X1 U15047 ( .IN1(n14111), .IN2(n14112), .Q(g26890) );
  AND2X1 U15048 ( .IN1(n8818), .IN2(g333), .Q(n14112) );
  AND2X1 U15049 ( .IN1(n5860), .IN2(n8690), .Q(n14111) );
  OR2X1 U15050 ( .IN1(n14113), .IN2(n14114), .Q(g26889) );
  AND4X1 U15051 ( .IN1(g329), .IN2(DFF_709_n1), .IN3(n14115), .IN4(n8723), .Q(
        n14114) );
  AND2X1 U15052 ( .IN1(n8818), .IN2(g29211), .Q(n14113) );
  OR2X1 U15053 ( .IN1(n14116), .IN2(n14117), .Q(g26888) );
  AND2X1 U15054 ( .IN1(n8818), .IN2(g29216), .Q(n14117) );
  AND2X1 U15055 ( .IN1(n8720), .IN2(g316), .Q(n14116) );
  OR3X1 U15056 ( .IN1(n14118), .IN2(n14119), .IN3(n14120), .Q(g26887) );
  AND3X1 U15057 ( .IN1(n5317), .IN2(g324), .IN3(n8735), .Q(n14119) );
  AND2X1 U15058 ( .IN1(n8818), .IN2(g336), .Q(n14118) );
  OR3X1 U15059 ( .IN1(n14121), .IN2(n14122), .IN3(n14123), .Q(g26886) );
  AND2X1 U15060 ( .IN1(n14120), .IN2(n14124), .Q(n14123) );
  AND2X1 U15061 ( .IN1(n8818), .IN2(g311), .Q(n14122) );
  AND3X1 U15062 ( .IN1(n14115), .IN2(g336), .IN3(n8734), .Q(n14121) );
  OR2X1 U15063 ( .IN1(n14125), .IN2(n14126), .Q(g26884) );
  AND2X1 U15064 ( .IN1(n14127), .IN2(n8704), .Q(n14126) );
  OR2X1 U15065 ( .IN1(n14128), .IN2(n14129), .Q(n14127) );
  AND2X1 U15066 ( .IN1(n14124), .IN2(n14130), .Q(n14129) );
  OR3X1 U15067 ( .IN1(n14131), .IN2(n14132), .IN3(g26885), .Q(n14130) );
  AND2X1 U15068 ( .IN1(g305), .IN2(g336), .Q(n14132) );
  AND2X1 U15069 ( .IN1(n5824), .IN2(g311), .Q(n14131) );
  AND4X1 U15070 ( .IN1(n5766), .IN2(n5456), .IN3(n5282), .IN4(n5317), .Q(
        n14128) );
  AND2X1 U15071 ( .IN1(n8818), .IN2(g329), .Q(n14125) );
  OR2X1 U15072 ( .IN1(n14133), .IN2(n14134), .Q(g26883) );
  AND2X1 U15073 ( .IN1(n14124), .IN2(n8703), .Q(n14134) );
  INVX0 U15074 ( .INP(n14115), .ZN(n14124) );
  OR2X1 U15075 ( .IN1(n14135), .IN2(n14136), .Q(n14115) );
  AND2X1 U15076 ( .IN1(n5827), .IN2(n5317), .Q(n14136) );
  AND2X1 U15077 ( .IN1(n5282), .IN2(g324), .Q(n14135) );
  AND2X1 U15078 ( .IN1(n8818), .IN2(g324), .Q(n14133) );
  OR3X1 U15079 ( .IN1(n14137), .IN2(n14138), .IN3(n14120), .Q(g26882) );
  AND2X1 U15080 ( .IN1(g305), .IN2(n8705), .Q(n14120) );
  AND2X1 U15081 ( .IN1(n8818), .IN2(g316), .Q(n14138) );
  AND2X1 U15082 ( .IN1(n8721), .IN2(g311), .Q(n14137) );
  OR2X1 U15083 ( .IN1(n14139), .IN2(n14140), .Q(g26881) );
  AND2X1 U15084 ( .IN1(n8818), .IN2(g305), .Q(n14140) );
  AND2X1 U15085 ( .IN1(g6744), .IN2(n8705), .Q(n14139) );
  INVX0 U15086 ( .INP(n14141), .ZN(g26877) );
  AND3X1 U15087 ( .IN1(n8726), .IN2(n9469), .IN3(n9468), .Q(n14141) );
  OR2X1 U15088 ( .IN1(n14142), .IN2(n14143), .Q(n9468) );
  OR4X1 U15089 ( .IN1(g2472), .IN2(g2204), .IN3(g2491), .IN4(g2223), .Q(n14143) );
  OR4X1 U15090 ( .IN1(g2338), .IN2(g2606), .IN3(test_so40), .IN4(g2357), .Q(
        n14142) );
  OR2X1 U15091 ( .IN1(n14144), .IN2(n14145), .Q(n9469) );
  OR4X1 U15092 ( .IN1(g2066), .IN2(g1798), .IN3(g1779), .IN4(g2047), .Q(n14145) );
  OR4X1 U15093 ( .IN1(g1913), .IN2(g1932), .IN3(test_so75), .IN4(g1664), .Q(
        n14144) );
  INVX0 U15094 ( .INP(n14146), .ZN(g26876) );
  AND3X1 U15095 ( .IN1(n8726), .IN2(n9489), .IN3(n9488), .Q(n14146) );
  OR2X1 U15096 ( .IN1(n14147), .IN2(n14148), .Q(n9488) );
  OR4X1 U15097 ( .IN1(n9324), .IN2(n9262), .IN3(n9295), .IN4(n9273), .Q(n14148) );
  OR4X1 U15098 ( .IN1(g2269), .IN2(g2537), .IN3(test_so31), .IN4(g2671), .Q(
        n14147) );
  OR2X1 U15099 ( .IN1(n14149), .IN2(n14150), .Q(n9489) );
  OR4X1 U15100 ( .IN1(g1858), .IN2(n9236), .IN3(g1992), .IN4(g2126), .Q(n14150) );
  OR4X1 U15101 ( .IN1(g1844), .IN2(g2112), .IN3(g1710), .IN4(g1978), .Q(n14149) );
  OR3X1 U15102 ( .IN1(n8792), .IN2(n9495), .IN3(n9494), .Q(g26875) );
  AND4X1 U15103 ( .IN1(n5414), .IN2(n5631), .IN3(n5281), .IN4(n5316), .Q(n9494) );
  AND4X1 U15104 ( .IN1(n5413), .IN2(n5628), .IN3(n5280), .IN4(n5315), .Q(n9495) );
  OR2X1 U15105 ( .IN1(n14151), .IN2(n14152), .Q(g25764) );
  AND2X1 U15106 ( .IN1(n14153), .IN2(g6541), .Q(n14152) );
  AND2X1 U15107 ( .IN1(n11664), .IN2(g6505), .Q(n14151) );
  OR3X1 U15108 ( .IN1(n14154), .IN2(n14155), .IN3(n14156), .Q(g25763) );
  AND2X1 U15109 ( .IN1(n11664), .IN2(g6537), .Q(n14156) );
  AND4X1 U15110 ( .IN1(n10569), .IN2(n8752), .IN3(n5659), .IN4(n5445), .Q(
        n14155) );
  AND2X1 U15111 ( .IN1(n14157), .IN2(g6533), .Q(n14154) );
  OR2X1 U15112 ( .IN1(n8799), .IN2(n14158), .Q(n14157) );
  AND2X1 U15113 ( .IN1(n10569), .IN2(g6527), .Q(n14158) );
  OR2X1 U15114 ( .IN1(n14159), .IN2(n14160), .Q(g25762) );
  AND2X1 U15115 ( .IN1(n14153), .IN2(g6527), .Q(n14160) );
  AND2X1 U15116 ( .IN1(n11664), .IN2(g6533), .Q(n14159) );
  OR3X1 U15117 ( .IN1(n14161), .IN2(n14162), .IN3(n14163), .Q(g25761) );
  AND2X1 U15118 ( .IN1(n11664), .IN2(g6513), .Q(n14163) );
  INVX0 U15119 ( .INP(n14153), .ZN(n11664) );
  OR2X1 U15120 ( .IN1(n8799), .IN2(n10569), .Q(n14153) );
  INVX0 U15121 ( .INP(n14164), .ZN(n14162) );
  OR2X1 U15122 ( .IN1(n8679), .IN2(n8407), .Q(n14164) );
  AND3X1 U15123 ( .IN1(n5426), .IN2(n10569), .IN3(n8735), .Q(n14161) );
  AND2X1 U15124 ( .IN1(g6561), .IN2(n11682), .Q(n10569) );
  INVX0 U15125 ( .INP(n1330), .ZN(n11682) );
  OR2X1 U15126 ( .IN1(n5563), .IN2(n5386), .Q(n1330) );
  OR2X1 U15127 ( .IN1(n14165), .IN2(n14166), .Q(g25758) );
  AND3X1 U15128 ( .IN1(n7986), .IN2(n14167), .IN3(n8735), .Q(n14166) );
  OR2X1 U15129 ( .IN1(n14168), .IN2(g6444), .Q(n14167) );
  AND2X1 U15130 ( .IN1(n7987), .IN2(g9743), .Q(n14168) );
  AND2X1 U15131 ( .IN1(n8818), .IN2(g6494), .Q(n14165) );
  OR2X1 U15132 ( .IN1(n14169), .IN2(n14170), .Q(g25757) );
  AND2X1 U15133 ( .IN1(n8818), .IN2(g6444), .Q(n14170) );
  AND2X1 U15134 ( .IN1(n8720), .IN2(g6727), .Q(n14169) );
  AND2X1 U15135 ( .IN1(g6573), .IN2(n8704), .Q(g25756) );
  OR2X1 U15136 ( .IN1(n14171), .IN2(n14172), .Q(g25750) );
  AND2X1 U15137 ( .IN1(n14173), .IN2(g6195), .Q(n14172) );
  AND2X1 U15138 ( .IN1(n11751), .IN2(g6159), .Q(n14171) );
  OR3X1 U15139 ( .IN1(n14174), .IN2(n14175), .IN3(n14176), .Q(g25749) );
  AND2X1 U15140 ( .IN1(n11751), .IN2(g6191), .Q(n14176) );
  AND4X1 U15141 ( .IN1(n10581), .IN2(n8753), .IN3(n5667), .IN4(n5453), .Q(
        n14175) );
  AND2X1 U15142 ( .IN1(n14177), .IN2(g6187), .Q(n14174) );
  OR2X1 U15143 ( .IN1(n8798), .IN2(n14178), .Q(n14177) );
  AND2X1 U15144 ( .IN1(n10581), .IN2(g6181), .Q(n14178) );
  OR2X1 U15145 ( .IN1(n14179), .IN2(n14180), .Q(g25748) );
  AND2X1 U15146 ( .IN1(n14173), .IN2(g6181), .Q(n14180) );
  AND2X1 U15147 ( .IN1(n11751), .IN2(g6187), .Q(n14179) );
  OR3X1 U15148 ( .IN1(n14181), .IN2(n14182), .IN3(n14183), .Q(g25747) );
  AND2X1 U15149 ( .IN1(n11751), .IN2(g6167), .Q(n14183) );
  INVX0 U15150 ( .INP(n14173), .ZN(n11751) );
  OR2X1 U15151 ( .IN1(n8798), .IN2(n10581), .Q(n14173) );
  INVX0 U15152 ( .INP(n14184), .ZN(n14182) );
  OR2X1 U15153 ( .IN1(n8679), .IN2(n8451), .Q(n14184) );
  AND3X1 U15154 ( .IN1(n5430), .IN2(n10581), .IN3(n8735), .Q(n14181) );
  AND2X1 U15155 ( .IN1(g6215), .IN2(n11769), .Q(n10581) );
  INVX0 U15156 ( .INP(n50), .ZN(n11769) );
  OR2X1 U15157 ( .IN1(n5568), .IN2(n5385), .Q(n50) );
  OR2X1 U15158 ( .IN1(n14185), .IN2(n14186), .Q(g25744) );
  AND3X1 U15159 ( .IN1(n7983), .IN2(n14187), .IN3(n8735), .Q(n14186) );
  OR2X1 U15160 ( .IN1(n14188), .IN2(g6098), .Q(n14187) );
  AND2X1 U15161 ( .IN1(test_so92), .IN2(n7984), .Q(n14188) );
  AND2X1 U15162 ( .IN1(n8818), .IN2(g6148), .Q(n14185) );
  OR2X1 U15163 ( .IN1(n14189), .IN2(n14190), .Q(g25743) );
  AND2X1 U15164 ( .IN1(n8818), .IN2(g6098), .Q(n14190) );
  AND2X1 U15165 ( .IN1(test_so69), .IN2(n8704), .Q(n14189) );
  AND2X1 U15166 ( .IN1(g6227), .IN2(n8704), .Q(g25742) );
  OR2X1 U15167 ( .IN1(n14191), .IN2(n14192), .Q(g25736) );
  AND2X1 U15168 ( .IN1(n14193), .IN2(g5849), .Q(n14192) );
  AND2X1 U15169 ( .IN1(n11837), .IN2(g5813), .Q(n14191) );
  OR3X1 U15170 ( .IN1(n14194), .IN2(n14195), .IN3(n14196), .Q(g25735) );
  AND2X1 U15171 ( .IN1(test_so83), .IN2(n11837), .Q(n14196) );
  AND4X1 U15172 ( .IN1(n10580), .IN2(n8752), .IN3(n5663), .IN4(n5449), .Q(
        n14195) );
  AND2X1 U15173 ( .IN1(n14197), .IN2(g5841), .Q(n14194) );
  OR2X1 U15174 ( .IN1(n8798), .IN2(n14198), .Q(n14197) );
  AND2X1 U15175 ( .IN1(n10580), .IN2(g5835), .Q(n14198) );
  OR2X1 U15176 ( .IN1(n14199), .IN2(n14200), .Q(g25734) );
  AND2X1 U15177 ( .IN1(n14193), .IN2(g5835), .Q(n14200) );
  AND2X1 U15178 ( .IN1(n11837), .IN2(g5841), .Q(n14199) );
  OR3X1 U15179 ( .IN1(n14201), .IN2(n14202), .IN3(n14203), .Q(g25733) );
  AND2X1 U15180 ( .IN1(n11837), .IN2(g5821), .Q(n14203) );
  INVX0 U15181 ( .INP(n14193), .ZN(n11837) );
  OR2X1 U15182 ( .IN1(n8798), .IN2(n10580), .Q(n14193) );
  INVX0 U15183 ( .INP(n14204), .ZN(n14202) );
  OR2X1 U15184 ( .IN1(n8679), .IN2(n8452), .Q(n14204) );
  AND3X1 U15185 ( .IN1(n5429), .IN2(n10580), .IN3(n8735), .Q(n14201) );
  AND2X1 U15186 ( .IN1(g5869), .IN2(n11855), .Q(n10580) );
  INVX0 U15187 ( .INP(n671), .ZN(n11855) );
  OR2X1 U15188 ( .IN1(n5388), .IN2(n8500), .Q(n671) );
  OR2X1 U15189 ( .IN1(n14205), .IN2(n14206), .Q(g25730) );
  AND3X1 U15190 ( .IN1(n7994), .IN2(n14207), .IN3(n8735), .Q(n14206) );
  OR2X1 U15191 ( .IN1(n14208), .IN2(g5752), .Q(n14207) );
  AND2X1 U15192 ( .IN1(n7995), .IN2(g9617), .Q(n14208) );
  AND2X1 U15193 ( .IN1(n8818), .IN2(g5802), .Q(n14205) );
  OR2X1 U15194 ( .IN1(n14209), .IN2(n14210), .Q(g25729) );
  AND2X1 U15195 ( .IN1(n8818), .IN2(g5752), .Q(n14210) );
  AND2X1 U15196 ( .IN1(n8720), .IN2(g6035), .Q(n14209) );
  AND2X1 U15197 ( .IN1(n8721), .IN2(test_so36), .Q(g25728) );
  OR2X1 U15198 ( .IN1(n14211), .IN2(n14212), .Q(g25722) );
  AND2X1 U15199 ( .IN1(n14213), .IN2(g5503), .Q(n14212) );
  AND2X1 U15200 ( .IN1(n11922), .IN2(g5467), .Q(n14211) );
  OR3X1 U15201 ( .IN1(n14214), .IN2(n14215), .IN3(n14216), .Q(g25721) );
  AND2X1 U15202 ( .IN1(n11922), .IN2(g5499), .Q(n14216) );
  AND4X1 U15203 ( .IN1(n10577), .IN2(n8753), .IN3(n5660), .IN4(n5446), .Q(
        n14215) );
  AND2X1 U15204 ( .IN1(n14217), .IN2(g5495), .Q(n14214) );
  OR2X1 U15205 ( .IN1(n8798), .IN2(n14218), .Q(n14217) );
  AND2X1 U15206 ( .IN1(n10577), .IN2(g5489), .Q(n14218) );
  OR2X1 U15207 ( .IN1(n14219), .IN2(n14220), .Q(g25720) );
  AND2X1 U15208 ( .IN1(n14213), .IN2(g5489), .Q(n14220) );
  AND2X1 U15209 ( .IN1(n11922), .IN2(g5495), .Q(n14219) );
  OR3X1 U15210 ( .IN1(n14221), .IN2(n14222), .IN3(n14223), .Q(g25719) );
  AND2X1 U15211 ( .IN1(n11922), .IN2(g5475), .Q(n14223) );
  INVX0 U15212 ( .INP(n14213), .ZN(n11922) );
  OR2X1 U15213 ( .IN1(n8798), .IN2(n10577), .Q(n14213) );
  INVX0 U15214 ( .INP(n14224), .ZN(n14222) );
  OR2X1 U15215 ( .IN1(n8679), .IN2(n8450), .Q(n14224) );
  AND3X1 U15216 ( .IN1(n5425), .IN2(n10577), .IN3(n8736), .Q(n14221) );
  AND2X1 U15217 ( .IN1(g5523), .IN2(n11940), .Q(n10577) );
  INVX0 U15218 ( .INP(n877), .ZN(n11940) );
  OR2X1 U15219 ( .IN1(n5566), .IN2(n5389), .Q(n877) );
  OR2X1 U15220 ( .IN1(n14225), .IN2(n14226), .Q(g25716) );
  AND3X1 U15221 ( .IN1(n14227), .IN2(n7988), .IN3(n8736), .Q(n14226) );
  OR2X1 U15222 ( .IN1(n14228), .IN2(g5406), .Q(n14227) );
  AND2X1 U15223 ( .IN1(n7989), .IN2(g9555), .Q(n14228) );
  AND2X1 U15224 ( .IN1(n8818), .IN2(g5456), .Q(n14225) );
  OR2X1 U15225 ( .IN1(n14229), .IN2(n14230), .Q(g25715) );
  AND2X1 U15226 ( .IN1(n8818), .IN2(g5406), .Q(n14230) );
  AND2X1 U15227 ( .IN1(n8720), .IN2(g5689), .Q(n14229) );
  AND2X1 U15228 ( .IN1(g5535), .IN2(n8704), .Q(g25714) );
  OR2X1 U15229 ( .IN1(n14231), .IN2(n14232), .Q(g25708) );
  AND2X1 U15230 ( .IN1(n14233), .IN2(g5156), .Q(n14232) );
  AND2X1 U15231 ( .IN1(n9099), .IN2(g5120), .Q(n14231) );
  OR2X1 U15232 ( .IN1(n14234), .IN2(n14235), .Q(g25706) );
  AND2X1 U15233 ( .IN1(n14233), .IN2(g5142), .Q(n14235) );
  AND2X1 U15234 ( .IN1(test_so98), .IN2(n9099), .Q(n14234) );
  OR3X1 U15235 ( .IN1(n14236), .IN2(n14237), .IN3(n14238), .Q(g25705) );
  AND2X1 U15236 ( .IN1(test_so96), .IN2(n9099), .Q(n14238) );
  INVX0 U15237 ( .INP(n14233), .ZN(n9099) );
  OR2X1 U15238 ( .IN1(n8797), .IN2(g32975), .Q(n14233) );
  INVX0 U15239 ( .INP(n14239), .ZN(n14237) );
  OR2X1 U15240 ( .IN1(n8678), .IN2(n8457), .Q(n14239) );
  AND3X1 U15241 ( .IN1(g32975), .IN2(n8516), .IN3(n8736), .Q(n14236) );
  AND2X1 U15242 ( .IN1(g5176), .IN2(n12025), .Q(g32975) );
  INVX0 U15243 ( .INP(n195), .ZN(n12025) );
  OR2X1 U15244 ( .IN1(n5567), .IN2(n5384), .Q(n195) );
  AND2X1 U15245 ( .IN1(n14240), .IN2(g5073), .Q(g25704) );
  OR2X1 U15246 ( .IN1(n8797), .IN2(g5069), .Q(n14240) );
  OR2X1 U15247 ( .IN1(n14241), .IN2(n14242), .Q(g25703) );
  AND3X1 U15248 ( .IN1(n5689), .IN2(n14243), .IN3(n8736), .Q(n14242) );
  INVX0 U15249 ( .INP(n14244), .ZN(n14243) );
  AND2X1 U15250 ( .IN1(n14245), .IN2(n8437), .Q(n14244) );
  OR2X1 U15251 ( .IN1(g5112), .IN2(n5690), .Q(n14245) );
  AND2X1 U15252 ( .IN1(n8818), .IN2(g5112), .Q(n14241) );
  OR2X1 U15253 ( .IN1(n14246), .IN2(n14247), .Q(g25702) );
  AND3X1 U15254 ( .IN1(n5690), .IN2(n14248), .IN3(n8736), .Q(n14247) );
  OR2X1 U15255 ( .IN1(n14249), .IN2(g5062), .Q(n14248) );
  INVX0 U15256 ( .INP(n14250), .ZN(n14249) );
  OR2X1 U15257 ( .IN1(n5689), .IN2(test_so32), .Q(n14250) );
  AND2X1 U15258 ( .IN1(test_so32), .IN2(n8810), .Q(n14246) );
  OR2X1 U15259 ( .IN1(n14251), .IN2(n14252), .Q(g25701) );
  AND2X1 U15260 ( .IN1(n8818), .IN2(g5062), .Q(n14252) );
  AND2X1 U15261 ( .IN1(test_so10), .IN2(n8703), .Q(n14251) );
  AND2X1 U15262 ( .IN1(g5188), .IN2(n8703), .Q(g25700) );
  OR3X1 U15263 ( .IN1(n14253), .IN2(n14254), .IN3(n14255), .Q(g25699) );
  AND2X1 U15264 ( .IN1(n8817), .IN2(g5097), .Q(n14255) );
  AND2X1 U15265 ( .IN1(n5014), .IN2(n5669), .Q(n14254) );
  INVX0 U15266 ( .INP(n14256), .ZN(n14253) );
  OR3X1 U15267 ( .IN1(n8792), .IN2(n5014), .IN3(n5669), .Q(n14256) );
  OR3X1 U15268 ( .IN1(n14257), .IN2(n14258), .IN3(n14259), .Q(g25698) );
  AND2X1 U15269 ( .IN1(n8817), .IN2(g5092), .Q(n14259) );
  AND2X1 U15270 ( .IN1(n5016), .IN2(n5753), .Q(n14258) );
  AND3X1 U15271 ( .IN1(n8726), .IN2(n14260), .IN3(g5097), .Q(n14257) );
  INVX0 U15272 ( .INP(n5016), .ZN(n14260) );
  XNOR2X1 U15273 ( .IN1(n5681), .IN2(n14261), .Q(g25697) );
  AND2X1 U15274 ( .IN1(n8720), .IN2(g5092), .Q(n14261) );
  OR3X1 U15275 ( .IN1(n14262), .IN2(n14263), .IN3(n14264), .Q(g25696) );
  AND3X1 U15276 ( .IN1(n8727), .IN2(g5077), .IN3(n8392), .Q(n14264) );
  AND3X1 U15277 ( .IN1(n14265), .IN2(n14266), .IN3(n5893), .Q(n14263) );
  OR2X1 U15278 ( .IN1(n5455), .IN2(g5069), .Q(n14266) );
  INVX0 U15279 ( .INP(n14267), .ZN(n14262) );
  OR2X1 U15280 ( .IN1(n14265), .IN2(n5893), .Q(n14267) );
  AND2X1 U15281 ( .IN1(n8720), .IN2(n5681), .Q(n14265) );
  AND2X1 U15282 ( .IN1(n14268), .IN2(g5077), .Q(g25695) );
  OR3X1 U15283 ( .IN1(n14269), .IN2(n14270), .IN3(n8792), .Q(n14268) );
  AND2X1 U15284 ( .IN1(n8392), .IN2(n5681), .Q(n14270) );
  INVX0 U15285 ( .INP(n14271), .ZN(n14269) );
  OR2X1 U15286 ( .IN1(g5069), .IN2(n5681), .Q(n14271) );
  OR2X1 U15287 ( .IN1(n14272), .IN2(n14273), .Q(g25691) );
  AND2X1 U15288 ( .IN1(n8817), .IN2(g4125), .Q(n14273) );
  AND2X1 U15289 ( .IN1(n8481), .IN2(n14274), .Q(n14272) );
  OR4X1 U15290 ( .IN1(n8491), .IN2(g4064), .IN3(g4057), .IN4(n14275), .Q(
        n14274) );
  OR4X1 U15291 ( .IN1(g4141), .IN2(g4082), .IN3(n5350), .IN4(n12004), .Q(
        n14275) );
  INVX0 U15292 ( .INP(n10568), .ZN(n12004) );
  AND2X1 U15293 ( .IN1(g4087), .IN2(n5340), .Q(n10568) );
  OR2X1 U15294 ( .IN1(n14276), .IN2(n14277), .Q(g25690) );
  AND3X1 U15295 ( .IN1(n8226), .IN2(g25689), .IN3(n8736), .Q(n14277) );
  AND2X1 U15296 ( .IN1(n8817), .IN2(g4169), .Q(n14276) );
  OR3X1 U15297 ( .IN1(n14278), .IN2(n14279), .IN3(n14280), .Q(g25687) );
  AND2X1 U15298 ( .IN1(n8817), .IN2(g4057), .Q(n14280) );
  AND2X1 U15299 ( .IN1(n5026), .IN2(n12105), .Q(n14279) );
  AND3X1 U15300 ( .IN1(n14281), .IN2(g4169), .IN3(n5612), .Q(n14278) );
  INVX0 U15301 ( .INP(n1166), .ZN(n14281) );
  OR2X1 U15302 ( .IN1(n5416), .IN2(n5711), .Q(n1166) );
  OR2X1 U15303 ( .IN1(n14282), .IN2(n14283), .Q(g25686) );
  AND3X1 U15304 ( .IN1(n12105), .IN2(g4057), .IN3(n5416), .Q(n14283) );
  AND2X1 U15305 ( .IN1(g4169), .IN2(n8702), .Q(n12105) );
  AND2X1 U15306 ( .IN1(n14284), .IN2(g4064), .Q(n14282) );
  OR2X1 U15307 ( .IN1(n8796), .IN2(n14285), .Q(n14284) );
  AND2X1 U15308 ( .IN1(n5711), .IN2(g4169), .Q(n14285) );
  OR3X1 U15309 ( .IN1(n14286), .IN2(n14287), .IN3(n8481), .Q(g25685) );
  AND2X1 U15310 ( .IN1(n8720), .IN2(n5729), .Q(n8481) );
  AND2X1 U15311 ( .IN1(n8817), .IN2(g4072), .Q(n14287) );
  AND2X1 U15312 ( .IN1(n5416), .IN2(n8702), .Q(n14286) );
  OR2X1 U15313 ( .IN1(n14288), .IN2(n14289), .Q(g25684) );
  AND2X1 U15314 ( .IN1(n14290), .IN2(g3849), .Q(n14289) );
  AND2X1 U15315 ( .IN1(n9011), .IN2(g3813), .Q(n14288) );
  OR2X1 U15316 ( .IN1(n14291), .IN2(n14292), .Q(g25682) );
  AND2X1 U15317 ( .IN1(n14290), .IN2(g3835), .Q(n14292) );
  AND2X1 U15318 ( .IN1(test_so97), .IN2(n9011), .Q(n14291) );
  OR3X1 U15319 ( .IN1(n14293), .IN2(n14294), .IN3(n14295), .Q(g25681) );
  AND2X1 U15320 ( .IN1(n9011), .IN2(g3821), .Q(n14295) );
  INVX0 U15321 ( .INP(n14290), .ZN(n9011) );
  OR2X1 U15322 ( .IN1(n8796), .IN2(n9012), .Q(n14290) );
  INVX0 U15323 ( .INP(n14296), .ZN(n14294) );
  OR2X1 U15324 ( .IN1(n8678), .IN2(n8429), .Q(n14296) );
  AND3X1 U15325 ( .IN1(n5428), .IN2(n9012), .IN3(n8736), .Q(n14293) );
  AND2X1 U15326 ( .IN1(n12127), .IN2(test_so33), .Q(n9012) );
  INVX0 U15327 ( .INP(n776), .ZN(n12127) );
  OR2X1 U15328 ( .IN1(n5564), .IN2(n5387), .Q(n776) );
  OR2X1 U15329 ( .IN1(n14297), .IN2(n14298), .Q(g25678) );
  AND3X1 U15330 ( .IN1(n7990), .IN2(n14299), .IN3(n8736), .Q(n14298) );
  OR2X1 U15331 ( .IN1(n14300), .IN2(g3752), .Q(n14299) );
  AND2X1 U15332 ( .IN1(n7991), .IN2(g8344), .Q(n14300) );
  AND2X1 U15333 ( .IN1(n8817), .IN2(g3802), .Q(n14297) );
  OR2X1 U15334 ( .IN1(n14301), .IN2(n14302), .Q(g25677) );
  AND2X1 U15335 ( .IN1(n8817), .IN2(g3752), .Q(n14302) );
  AND2X1 U15336 ( .IN1(n8720), .IN2(g4040), .Q(n14301) );
  AND2X1 U15337 ( .IN1(g3881), .IN2(n8701), .Q(g25676) );
  OR2X1 U15338 ( .IN1(n14303), .IN2(n14304), .Q(g25670) );
  AND2X1 U15339 ( .IN1(n14305), .IN2(g3498), .Q(n14304) );
  AND2X1 U15340 ( .IN1(n12194), .IN2(g3462), .Q(n14303) );
  OR3X1 U15341 ( .IN1(n14306), .IN2(n14307), .IN3(n14308), .Q(g25669) );
  AND2X1 U15342 ( .IN1(n12194), .IN2(g3494), .Q(n14308) );
  AND4X1 U15343 ( .IN1(n10572), .IN2(n8753), .IN3(n5668), .IN4(n5454), .Q(
        n14307) );
  AND2X1 U15344 ( .IN1(n14309), .IN2(g3490), .Q(n14306) );
  OR2X1 U15345 ( .IN1(n8796), .IN2(n14310), .Q(n14309) );
  AND2X1 U15346 ( .IN1(n10572), .IN2(g3484), .Q(n14310) );
  OR2X1 U15347 ( .IN1(n14311), .IN2(n14312), .Q(g25668) );
  AND2X1 U15348 ( .IN1(n14305), .IN2(g3484), .Q(n14312) );
  AND2X1 U15349 ( .IN1(n12194), .IN2(g3490), .Q(n14311) );
  OR3X1 U15350 ( .IN1(n14313), .IN2(n14314), .IN3(n14315), .Q(g25667) );
  AND2X1 U15351 ( .IN1(n12194), .IN2(g3470), .Q(n14315) );
  INVX0 U15352 ( .INP(n14305), .ZN(n12194) );
  OR2X1 U15353 ( .IN1(n8795), .IN2(n10572), .Q(n14305) );
  INVX0 U15354 ( .INP(n14316), .ZN(n14314) );
  OR2X1 U15355 ( .IN1(n8678), .IN2(n8430), .Q(n14316) );
  AND3X1 U15356 ( .IN1(n5424), .IN2(n10572), .IN3(n8737), .Q(n14313) );
  AND2X1 U15357 ( .IN1(g3518), .IN2(n12212), .Q(n10572) );
  INVX0 U15358 ( .INP(n417), .ZN(n12212) );
  OR2X1 U15359 ( .IN1(n5569), .IN2(n5383), .Q(n417) );
  OR2X1 U15360 ( .IN1(n14317), .IN2(n14318), .Q(g25664) );
  AND3X1 U15361 ( .IN1(n7974), .IN2(n14319), .IN3(n8737), .Q(n14318) );
  OR2X1 U15362 ( .IN1(n14320), .IN2(g3401), .Q(n14319) );
  AND2X1 U15363 ( .IN1(n7975), .IN2(g8279), .Q(n14320) );
  AND2X1 U15364 ( .IN1(n8817), .IN2(g3451), .Q(n14317) );
  OR2X1 U15365 ( .IN1(n14321), .IN2(n14322), .Q(g25663) );
  AND2X1 U15366 ( .IN1(n8817), .IN2(g3401), .Q(n14322) );
  AND2X1 U15367 ( .IN1(n8719), .IN2(g3689), .Q(n14321) );
  AND2X1 U15368 ( .IN1(g3530), .IN2(n8701), .Q(g25662) );
  OR2X1 U15369 ( .IN1(n14323), .IN2(n14324), .Q(g25656) );
  AND2X1 U15370 ( .IN1(n14325), .IN2(g3147), .Q(n14324) );
  AND2X1 U15371 ( .IN1(n12279), .IN2(g3111), .Q(n14323) );
  OR3X1 U15372 ( .IN1(n14326), .IN2(n14327), .IN3(n14328), .Q(g25655) );
  INVX0 U15373 ( .INP(n14329), .ZN(n14328) );
  OR2X1 U15374 ( .IN1(n14325), .IN2(n5882), .Q(n14329) );
  AND4X1 U15375 ( .IN1(n10567), .IN2(n8753), .IN3(n5661), .IN4(n5447), .Q(
        n14327) );
  AND2X1 U15376 ( .IN1(n14330), .IN2(g3139), .Q(n14326) );
  OR2X1 U15377 ( .IN1(n8795), .IN2(n14331), .Q(n14330) );
  AND2X1 U15378 ( .IN1(n10567), .IN2(g3133), .Q(n14331) );
  OR2X1 U15379 ( .IN1(n14332), .IN2(n14333), .Q(g25654) );
  AND2X1 U15380 ( .IN1(n14325), .IN2(g3133), .Q(n14333) );
  AND2X1 U15381 ( .IN1(n12279), .IN2(g3139), .Q(n14332) );
  OR3X1 U15382 ( .IN1(n14334), .IN2(n14335), .IN3(n14336), .Q(g25653) );
  AND2X1 U15383 ( .IN1(n12279), .IN2(g3119), .Q(n14336) );
  INVX0 U15384 ( .INP(n14325), .ZN(n12279) );
  OR2X1 U15385 ( .IN1(n8796), .IN2(n10567), .Q(n14325) );
  INVX0 U15386 ( .INP(n14337), .ZN(n14335) );
  OR2X1 U15387 ( .IN1(n8678), .IN2(n8408), .Q(n14337) );
  AND3X1 U15388 ( .IN1(n5423), .IN2(n10567), .IN3(n8737), .Q(n14334) );
  AND2X1 U15389 ( .IN1(g3167), .IN2(n12297), .Q(n10567) );
  INVX0 U15390 ( .INP(n509), .ZN(n12297) );
  OR2X1 U15391 ( .IN1(n5603), .IN2(n5390), .Q(n509) );
  OR2X1 U15392 ( .IN1(n14338), .IN2(n14339), .Q(g25650) );
  AND3X1 U15393 ( .IN1(n7996), .IN2(n14340), .IN3(n8737), .Q(n14339) );
  OR2X1 U15394 ( .IN1(n14341), .IN2(g3050), .Q(n14340) );
  AND2X1 U15395 ( .IN1(n7997), .IN2(g8215), .Q(n14341) );
  AND2X1 U15396 ( .IN1(n8817), .IN2(g3100), .Q(n14338) );
  OR2X1 U15397 ( .IN1(n14342), .IN2(n14343), .Q(g25649) );
  AND2X1 U15398 ( .IN1(n8817), .IN2(g3050), .Q(n14343) );
  AND2X1 U15399 ( .IN1(n8719), .IN2(g3338), .Q(n14342) );
  AND2X1 U15400 ( .IN1(g3179), .IN2(n8700), .Q(g25648) );
  OR3X1 U15401 ( .IN1(n14344), .IN2(n14345), .IN3(n5045), .Q(g25639) );
  AND2X1 U15402 ( .IN1(n13085), .IN2(n8700), .Q(n14345) );
  AND2X1 U15403 ( .IN1(g2719), .IN2(n5299), .Q(n13085) );
  AND2X1 U15404 ( .IN1(n8817), .IN2(g2715), .Q(n14344) );
  OR2X1 U15405 ( .IN1(n14346), .IN2(n14347), .Q(g25638) );
  AND2X1 U15406 ( .IN1(n14348), .IN2(n8700), .Q(n14347) );
  OR2X1 U15407 ( .IN1(n14349), .IN2(n14350), .Q(n14348) );
  AND3X1 U15408 ( .IN1(n14351), .IN2(n5768), .IN3(n5441), .Q(n14350) );
  AND2X1 U15409 ( .IN1(n14352), .IN2(g1559), .Q(n14349) );
  AND2X1 U15410 ( .IN1(n8817), .IN2(g1564), .Q(n14346) );
  OR2X1 U15411 ( .IN1(n14353), .IN2(n14354), .Q(g25637) );
  AND2X1 U15412 ( .IN1(n14355), .IN2(g1559), .Q(n14354) );
  OR2X1 U15413 ( .IN1(n8795), .IN2(n14356), .Q(n14355) );
  AND2X1 U15414 ( .IN1(n14351), .IN2(n5768), .Q(n14356) );
  AND3X1 U15415 ( .IN1(n8726), .IN2(g1554), .IN3(n14352), .Q(n14353) );
  OR3X1 U15416 ( .IN1(n14357), .IN2(n14358), .IN3(n14359), .Q(g25636) );
  AND2X1 U15417 ( .IN1(n14360), .IN2(n10805), .Q(n14359) );
  AND3X1 U15418 ( .IN1(n14361), .IN2(g1306), .IN3(n8737), .Q(n14358) );
  INVX0 U15419 ( .INP(n14362), .ZN(n14361) );
  AND2X1 U15420 ( .IN1(g7946), .IN2(n10805), .Q(n14362) );
  AND2X1 U15421 ( .IN1(g1514), .IN2(test_so49), .Q(n10805) );
  AND2X1 U15422 ( .IN1(n8817), .IN2(g1521), .Q(n14357) );
  OR2X1 U15423 ( .IN1(n14363), .IN2(n14364), .Q(g25635) );
  AND2X1 U15424 ( .IN1(n14365), .IN2(g1300), .Q(n14364) );
  OR2X1 U15425 ( .IN1(n14366), .IN2(n13141), .Q(n14365) );
  AND2X1 U15426 ( .IN1(n14367), .IN2(n8700), .Q(n14366) );
  OR2X1 U15427 ( .IN1(n5865), .IN2(n14368), .Q(n14367) );
  AND2X1 U15428 ( .IN1(n14369), .IN2(g1484), .Q(n14363) );
  OR2X1 U15429 ( .IN1(n8807), .IN2(n14370), .Q(n14369) );
  AND3X1 U15430 ( .IN1(n13143), .IN2(n5483), .IN3(n13978), .Q(n14370) );
  INVX0 U15431 ( .INP(n14368), .ZN(n13978) );
  OR2X1 U15432 ( .IN1(n8222), .IN2(test_so12), .Q(n14368) );
  AND3X1 U15433 ( .IN1(n13992), .IN2(n8496), .IN3(n14371), .Q(g25634) );
  OR2X1 U15434 ( .IN1(n14372), .IN2(n14373), .Q(n14371) );
  AND2X1 U15435 ( .IN1(n8719), .IN2(g1395), .Q(n14373) );
  AND2X1 U15436 ( .IN1(n11076), .IN2(n14374), .Q(n14372) );
  INVX0 U15437 ( .INP(n14375), .ZN(n14374) );
  OR3X1 U15438 ( .IN1(n8134), .IN2(n5655), .IN3(n14375), .Q(n13992) );
  OR3X1 U15439 ( .IN1(n14376), .IN2(n14377), .IN3(n14378), .Q(g25633) );
  AND3X1 U15440 ( .IN1(n14379), .IN2(n8434), .IN3(n13996), .Q(n14378) );
  AND2X1 U15441 ( .IN1(n8817), .IN2(g1379), .Q(n14377) );
  AND3X1 U15442 ( .IN1(n13998), .IN2(g1384), .IN3(n8737), .Q(n14376) );
  OR2X1 U15443 ( .IN1(n14380), .IN2(n14381), .Q(g25632) );
  AND3X1 U15444 ( .IN1(n14382), .IN2(n14383), .IN3(n13996), .Q(n14381) );
  AND2X1 U15445 ( .IN1(g1351), .IN2(n8700), .Q(n13996) );
  OR2X1 U15446 ( .IN1(n12640), .IN2(n14384), .Q(n14383) );
  OR2X1 U15447 ( .IN1(n8326), .IN2(n13998), .Q(n14382) );
  AND2X1 U15448 ( .IN1(n14385), .IN2(g1312), .Q(n14380) );
  OR2X1 U15449 ( .IN1(n8806), .IN2(n14379), .Q(n14385) );
  AND2X1 U15450 ( .IN1(n14386), .IN2(n8699), .Q(g25631) );
  OR2X1 U15451 ( .IN1(n14387), .IN2(n14388), .Q(n14386) );
  AND2X1 U15452 ( .IN1(n13998), .IN2(g1312), .Q(n14388) );
  AND3X1 U15453 ( .IN1(n14389), .IN2(n14390), .IN3(n13732), .Q(n14387) );
  INVX0 U15454 ( .INP(n12640), .ZN(n13732) );
  OR2X1 U15455 ( .IN1(n9102), .IN2(g1351), .Q(n14390) );
  AND4X1 U15456 ( .IN1(g1379), .IN2(n13738), .IN3(g1345), .IN4(g1367), .Q(
        n9102) );
  OR2X1 U15457 ( .IN1(n5322), .IN2(n14391), .Q(n14389) );
  AND2X1 U15458 ( .IN1(n13737), .IN2(n13733), .Q(n14391) );
  OR2X1 U15459 ( .IN1(n8326), .IN2(n13738), .Q(n13733) );
  INVX0 U15460 ( .INP(n14384), .ZN(n13737) );
  OR2X1 U15461 ( .IN1(n8328), .IN2(n8325), .Q(n14384) );
  OR2X1 U15462 ( .IN1(n14392), .IN2(n14393), .Q(g25630) );
  AND2X1 U15463 ( .IN1(g24247), .IN2(g1266), .Q(n14393) );
  AND2X1 U15464 ( .IN1(n14394), .IN2(g1249), .Q(n14392) );
  OR2X1 U15465 ( .IN1(n8806), .IN2(n14395), .Q(n14394) );
  AND2X1 U15466 ( .IN1(n8042), .IN2(g12923), .Q(n14395) );
  OR2X1 U15467 ( .IN1(n14396), .IN2(n14397), .Q(g25629) );
  AND2X1 U15468 ( .IN1(n14398), .IN2(n8699), .Q(n14397) );
  OR2X1 U15469 ( .IN1(n14399), .IN2(n14400), .Q(n14398) );
  AND3X1 U15470 ( .IN1(n14401), .IN2(n8507), .IN3(n5442), .Q(n14400) );
  AND2X1 U15471 ( .IN1(n14402), .IN2(g1216), .Q(n14399) );
  AND2X1 U15472 ( .IN1(n8817), .IN2(g1221), .Q(n14396) );
  OR2X1 U15473 ( .IN1(n14403), .IN2(n14404), .Q(g25628) );
  AND2X1 U15474 ( .IN1(n14405), .IN2(g1216), .Q(n14404) );
  OR2X1 U15475 ( .IN1(n8806), .IN2(n14406), .Q(n14405) );
  AND2X1 U15476 ( .IN1(n14401), .IN2(n8507), .Q(n14406) );
  AND3X1 U15477 ( .IN1(n14402), .IN2(n8724), .IN3(test_so76), .Q(n14403) );
  INVX0 U15478 ( .INP(n14401), .ZN(n14402) );
  OR2X1 U15479 ( .IN1(n14407), .IN2(n14408), .Q(g25627) );
  AND2X1 U15480 ( .IN1(n14409), .IN2(n8699), .Q(n14408) );
  OR2X1 U15481 ( .IN1(n14410), .IN2(n14411), .Q(n14409) );
  AND2X1 U15482 ( .IN1(n14412), .IN2(g962), .Q(n14411) );
  INVX0 U15483 ( .INP(n14413), .ZN(n14412) );
  AND2X1 U15484 ( .IN1(n14413), .IN2(g996), .Q(n14410) );
  AND3X1 U15485 ( .IN1(g1183), .IN2(g1171), .IN3(g7916), .Q(n14413) );
  AND2X1 U15486 ( .IN1(n8817), .IN2(g1178), .Q(n14407) );
  OR2X1 U15487 ( .IN1(n14414), .IN2(n14415), .Q(g25626) );
  AND2X1 U15488 ( .IN1(n14416), .IN2(g956), .Q(n14415) );
  OR2X1 U15489 ( .IN1(n14417), .IN2(n13176), .Q(n14416) );
  AND2X1 U15490 ( .IN1(n14418), .IN2(n8699), .Q(n14417) );
  INVX0 U15491 ( .INP(n14419), .ZN(n14418) );
  AND2X1 U15492 ( .IN1(g1141), .IN2(n14012), .Q(n14419) );
  AND2X1 U15493 ( .IN1(n14420), .IN2(g1141), .Q(n14414) );
  OR2X1 U15494 ( .IN1(n8804), .IN2(n14421), .Q(n14420) );
  AND3X1 U15495 ( .IN1(n13178), .IN2(n5341), .IN3(n14012), .Q(n14421) );
  AND2X1 U15496 ( .IN1(test_so7), .IN2(n5618), .Q(n14012) );
  AND3X1 U15497 ( .IN1(n14422), .IN2(n14026), .IN3(n5320), .Q(g25625) );
  OR3X1 U15498 ( .IN1(n8135), .IN2(n5654), .IN3(n14423), .Q(n14026) );
  OR2X1 U15499 ( .IN1(n14424), .IN2(n14425), .Q(n14422) );
  AND2X1 U15500 ( .IN1(n8719), .IN2(g1052), .Q(n14425) );
  AND2X1 U15501 ( .IN1(n11091), .IN2(n14426), .Q(n14424) );
  INVX0 U15502 ( .INP(n14423), .ZN(n14426) );
  OR3X1 U15503 ( .IN1(n14427), .IN2(n14428), .IN3(n14429), .Q(g25624) );
  AND3X1 U15504 ( .IN1(n14430), .IN2(n8435), .IN3(n14030), .Q(n14429) );
  AND2X1 U15505 ( .IN1(n8817), .IN2(g1036), .Q(n14428) );
  AND3X1 U15506 ( .IN1(n14032), .IN2(g1041), .IN3(n8737), .Q(n14427) );
  OR2X1 U15507 ( .IN1(n14431), .IN2(n14432), .Q(g25623) );
  AND3X1 U15508 ( .IN1(n14433), .IN2(n14434), .IN3(n14030), .Q(n14432) );
  AND2X1 U15509 ( .IN1(g1008), .IN2(n8699), .Q(n14030) );
  INVX0 U15510 ( .INP(n14435), .ZN(n14434) );
  AND2X1 U15511 ( .IN1(n13746), .IN2(n13752), .Q(n14435) );
  OR2X1 U15512 ( .IN1(n8243), .IN2(n14032), .Q(n14433) );
  AND2X1 U15513 ( .IN1(test_so20), .IN2(n14436), .Q(n14431) );
  OR2X1 U15514 ( .IN1(n8806), .IN2(n14430), .Q(n14436) );
  INVX0 U15515 ( .INP(n14032), .ZN(n14430) );
  AND2X1 U15516 ( .IN1(n14437), .IN2(n8699), .Q(g25622) );
  OR2X1 U15517 ( .IN1(n14438), .IN2(n14439), .Q(n14437) );
  AND2X1 U15518 ( .IN1(test_so20), .IN2(n14032), .Q(n14439) );
  AND3X1 U15519 ( .IN1(n14440), .IN2(n14441), .IN3(n13746), .Q(n14438) );
  INVX0 U15520 ( .INP(n12674), .ZN(n13746) );
  OR2X1 U15521 ( .IN1(n9095), .IN2(g1008), .Q(n14441) );
  AND4X1 U15522 ( .IN1(g1036), .IN2(n13750), .IN3(g1002), .IN4(g1024), .Q(
        n9095) );
  OR2X1 U15523 ( .IN1(n5321), .IN2(n14442), .Q(n14440) );
  AND2X1 U15524 ( .IN1(n13752), .IN2(n13747), .Q(n14442) );
  OR2X1 U15525 ( .IN1(n8243), .IN2(n13750), .Q(n13747) );
  AND2X1 U15526 ( .IN1(g1030), .IN2(g1018), .Q(n13752) );
  OR2X1 U15527 ( .IN1(n14443), .IN2(n14444), .Q(g25621) );
  AND2X1 U15528 ( .IN1(g24231), .IN2(g921), .Q(n14444) );
  AND2X1 U15529 ( .IN1(n14445), .IN2(g904), .Q(n14443) );
  OR2X1 U15530 ( .IN1(n8806), .IN2(n14446), .Q(n14445) );
  AND2X1 U15531 ( .IN1(n8041), .IN2(g12919), .Q(n14446) );
  AND2X1 U15532 ( .IN1(n14447), .IN2(g837), .Q(g25619) );
  OR2X1 U15533 ( .IN1(n8806), .IN2(n14448), .Q(n14447) );
  XOR2X1 U15534 ( .IN1(n14075), .IN2(g843), .Q(n14448) );
  OR2X1 U15535 ( .IN1(n14449), .IN2(n14450), .Q(g25618) );
  AND2X1 U15536 ( .IN1(n14451), .IN2(g832), .Q(n14450) );
  OR2X1 U15537 ( .IN1(n14452), .IN2(n14453), .Q(n14451) );
  AND2X1 U15538 ( .IN1(n5822), .IN2(n4518), .Q(n14453) );
  AND2X1 U15539 ( .IN1(n8719), .IN2(n13200), .Q(n4518) );
  AND2X1 U15540 ( .IN1(n13236), .IN2(n13200), .Q(n14452) );
  AND2X1 U15541 ( .IN1(n14454), .IN2(g817), .Q(n14449) );
  OR2X1 U15542 ( .IN1(n8806), .IN2(n14455), .Q(n14454) );
  AND3X1 U15543 ( .IN1(n4948), .IN2(n13200), .IN3(n8216), .Q(n14455) );
  OR2X1 U15544 ( .IN1(n14456), .IN2(n14457), .Q(g25617) );
  AND2X1 U15545 ( .IN1(n8817), .IN2(g812), .Q(n14457) );
  AND3X1 U15546 ( .IN1(n14458), .IN2(n14459), .IN3(n13200), .Q(n14456) );
  OR2X1 U15547 ( .IN1(n14460), .IN2(n5709), .Q(n13200) );
  AND2X1 U15548 ( .IN1(n5733), .IN2(g837), .Q(n14460) );
  OR2X1 U15549 ( .IN1(n13237), .IN2(g817), .Q(n14459) );
  OR2X1 U15550 ( .IN1(n5822), .IN2(n13236), .Q(n14458) );
  AND2X1 U15551 ( .IN1(n14461), .IN2(n8699), .Q(g25616) );
  XOR3X1 U15552 ( .IN1(n14462), .IN2(n14463), .IN3(n14464), .Q(n14461) );
  XOR2X1 U15553 ( .IN1(g225), .IN2(n14465), .Q(n14464) );
  AND2X1 U15554 ( .IN1(g732), .IN2(n13815), .Q(n14465) );
  OR4X1 U15555 ( .IN1(n13796), .IN2(n13794), .IN3(g528), .IN4(n14466), .Q(
        n13815) );
  OR2X1 U15556 ( .IN1(g490), .IN2(g482), .Q(n14466) );
  OR2X1 U15557 ( .IN1(test_so54), .IN2(g518), .Q(n13796) );
  XOR3X1 U15558 ( .IN1(n8331), .IN2(n8330), .IN3(n14467), .Q(n14463) );
  XOR2X1 U15559 ( .IN1(n8333), .IN2(n8332), .Q(n14467) );
  XOR2X1 U15560 ( .IN1(n8329), .IN2(n6008), .Q(n14462) );
  OR2X1 U15561 ( .IN1(n14468), .IN2(n14469), .Q(g25615) );
  AND2X1 U15562 ( .IN1(n14470), .IN2(g686), .Q(n14469) );
  AND2X1 U15563 ( .IN1(n13785), .IN2(g667), .Q(n14468) );
  OR3X1 U15564 ( .IN1(n14471), .IN2(n14472), .IN3(n14473), .Q(g25614) );
  AND2X1 U15565 ( .IN1(n8817), .IN2(g691), .Q(n14473) );
  AND2X1 U15566 ( .IN1(n5111), .IN2(n14100), .Q(n14472) );
  AND2X1 U15567 ( .IN1(n13785), .IN2(g686), .Q(n14471) );
  OR2X1 U15568 ( .IN1(n14474), .IN2(n14475), .Q(g25613) );
  AND2X1 U15569 ( .IN1(n8817), .IN2(g559), .Q(n14475) );
  AND3X1 U15570 ( .IN1(n2421), .IN2(n14476), .IN3(n14477), .Q(n14474) );
  XOR2X1 U15571 ( .IN1(n14092), .IN2(g562), .Q(n14477) );
  INVX0 U15572 ( .INP(n14478), .ZN(n14092) );
  OR2X1 U15573 ( .IN1(n14479), .IN2(n8359), .Q(n14478) );
  AND2X1 U15574 ( .IN1(n7946), .IN2(g12368), .Q(n14479) );
  OR2X1 U15575 ( .IN1(n5288), .IN2(n14833), .Q(n14476) );
  OR2X1 U15576 ( .IN1(n14480), .IN2(n14481), .Q(g25612) );
  AND2X1 U15577 ( .IN1(n13785), .IN2(g518), .Q(n14481) );
  AND2X1 U15578 ( .IN1(n14482), .IN2(g513), .Q(n14480) );
  OR2X1 U15579 ( .IN1(n14483), .IN2(n14484), .Q(g25611) );
  AND2X1 U15580 ( .IN1(n13785), .IN2(g513), .Q(n14484) );
  AND2X1 U15581 ( .IN1(n14482), .IN2(g504), .Q(n14483) );
  OR2X1 U15582 ( .IN1(n8806), .IN2(n14485), .Q(n14482) );
  AND2X1 U15583 ( .IN1(n14100), .IN2(n13231), .Q(n14485) );
  INVX0 U15584 ( .INP(n4962), .ZN(n13231) );
  OR3X1 U15585 ( .IN1(n14486), .IN2(n14487), .IN3(n14488), .Q(g25610) );
  AND2X1 U15586 ( .IN1(test_so54), .IN2(n14470), .Q(n14487) );
  AND2X1 U15587 ( .IN1(n13785), .IN2(g504), .Q(n14486) );
  OR3X1 U15588 ( .IN1(n14488), .IN2(n14489), .IN3(n14490), .Q(g25609) );
  AND2X1 U15589 ( .IN1(n13781), .IN2(n5287), .Q(n14490) );
  AND2X1 U15590 ( .IN1(test_so54), .IN2(n14491), .Q(n14489) );
  OR2X1 U15591 ( .IN1(n14492), .IN2(n13785), .Q(n14491) );
  INVX0 U15592 ( .INP(n14470), .ZN(n13785) );
  OR2X1 U15593 ( .IN1(n8806), .IN2(n14100), .Q(n14470) );
  AND2X1 U15594 ( .IN1(n5548), .IN2(n8699), .Q(n14492) );
  AND2X1 U15595 ( .IN1(n13781), .IN2(n4962), .Q(n14488) );
  AND2X1 U15596 ( .IN1(n8719), .IN2(n14100), .Q(n13781) );
  AND3X1 U15597 ( .IN1(g358), .IN2(g385), .IN3(n5633), .Q(n14100) );
  OR3X1 U15598 ( .IN1(n14493), .IN2(n14494), .IN3(n14495), .Q(g25605) );
  AND2X1 U15599 ( .IN1(n14496), .IN2(g460), .Q(n14495) );
  AND3X1 U15600 ( .IN1(n14497), .IN2(g246), .IN3(n8738), .Q(n14494) );
  AND2X1 U15601 ( .IN1(n8816), .IN2(g168), .Q(n14493) );
  OR2X1 U15602 ( .IN1(n14498), .IN2(n14499), .Q(g25604) );
  AND2X1 U15603 ( .IN1(n14500), .IN2(g460), .Q(n14499) );
  AND2X1 U15604 ( .IN1(n14496), .IN2(g452), .Q(n14498) );
  OR3X1 U15605 ( .IN1(n14501), .IN2(n14502), .IN3(n14503), .Q(g25602) );
  AND2X1 U15606 ( .IN1(n14496), .IN2(test_so72), .Q(n14503) );
  AND3X1 U15607 ( .IN1(n14497), .IN2(g446), .IN3(n8738), .Q(n14502) );
  AND2X1 U15608 ( .IN1(n8816), .IN2(g405), .Q(n14501) );
  OR2X1 U15609 ( .IN1(n14504), .IN2(n14505), .Q(g25601) );
  AND2X1 U15610 ( .IN1(test_so72), .IN2(n14500), .Q(n14505) );
  AND2X1 U15611 ( .IN1(n14496), .IN2(g174), .Q(n14504) );
  OR2X1 U15612 ( .IN1(n14506), .IN2(n14507), .Q(g25600) );
  AND2X1 U15613 ( .IN1(n14500), .IN2(g174), .Q(n14507) );
  AND2X1 U15614 ( .IN1(n14496), .IN2(g168), .Q(n14506) );
  INVX0 U15615 ( .INP(n14500), .ZN(n14496) );
  OR2X1 U15616 ( .IN1(n8806), .IN2(n14497), .Q(n14500) );
  INVX0 U15617 ( .INP(n13794), .ZN(n14497) );
  OR2X1 U15618 ( .IN1(n5121), .IN2(g370), .Q(n13794) );
  OR2X1 U15619 ( .IN1(n14508), .IN2(n14509), .Q(g25599) );
  INVX0 U15620 ( .INP(n9795), .ZN(n14509) );
  AND2X1 U15621 ( .IN1(n8816), .IN2(g385), .Q(n14508) );
  OR2X1 U15622 ( .IN1(n14510), .IN2(n14511), .Q(g25598) );
  AND2X1 U15623 ( .IN1(n14512), .IN2(g376), .Q(n14511) );
  OR2X1 U15624 ( .IN1(n8805), .IN2(n14513), .Q(n14512) );
  AND2X1 U15625 ( .IN1(n5121), .IN2(g358), .Q(n14513) );
  AND3X1 U15626 ( .IN1(n8726), .IN2(g385), .IN3(n5121), .Q(n14510) );
  OR3X1 U15627 ( .IN1(n8458), .IN2(n5633), .IN3(n5632), .Q(n5121) );
  OR2X1 U15628 ( .IN1(n14514), .IN2(n14515), .Q(g25597) );
  AND2X1 U15629 ( .IN1(n14516), .IN2(n8698), .Q(n14515) );
  XOR2X1 U15630 ( .IN1(n9795), .IN2(n8307), .Q(n14516) );
  OR3X1 U15631 ( .IN1(n8361), .IN2(n5633), .IN3(n5632), .Q(n9795) );
  AND2X1 U15632 ( .IN1(n8816), .IN2(g358), .Q(n14514) );
  OR2X1 U15633 ( .IN1(n14517), .IN2(n14518), .Q(g25596) );
  AND2X1 U15634 ( .IN1(n14519), .IN2(n8698), .Q(n14518) );
  XOR2X1 U15635 ( .IN1(n8458), .IN2(n5633), .Q(n14519) );
  AND2X1 U15636 ( .IN1(n8816), .IN2(g370), .Q(n14517) );
  AND3X1 U15637 ( .IN1(n8458), .IN2(n8724), .IN3(n8361), .Q(g25595) );
  AND3X1 U15638 ( .IN1(n13813), .IN2(n8725), .IN3(n13811), .Q(g25594) );
  OR2X1 U15639 ( .IN1(n14520), .IN2(g278), .Q(n13811) );
  AND4X1 U15640 ( .IN1(n6008), .IN2(n8329), .IN3(n8330), .IN4(n14521), .Q(
        n14520) );
  AND4X1 U15641 ( .IN1(g269), .IN2(n5597), .IN3(g262), .IN4(g255), .Q(n14521)
         );
  OR4X1 U15642 ( .IN1(g269), .IN2(g255), .IN3(g262), .IN4(n14522), .Q(n13813)
         );
  OR4X1 U15643 ( .IN1(n6008), .IN2(n5597), .IN3(n8330), .IN4(n8329), .Q(n14522) );
  OR2X1 U15644 ( .IN1(n14523), .IN2(n14524), .Q(g25593) );
  AND2X1 U15645 ( .IN1(n14525), .IN2(n8698), .Q(n14524) );
  OR2X1 U15646 ( .IN1(n14526), .IN2(n14527), .Q(n14525) );
  AND2X1 U15647 ( .IN1(n14528), .IN2(n14529), .Q(n14527) );
  INVX0 U15648 ( .INP(n14530), .ZN(n14529) );
  AND2X1 U15649 ( .IN1(n14530), .IN2(g209), .Q(n14526) );
  INVX0 U15650 ( .INP(n14531), .ZN(n14523) );
  OR2X1 U15651 ( .IN1(n8679), .IN2(n8048), .Q(n14531) );
  OR2X1 U15652 ( .IN1(n14532), .IN2(n14533), .Q(g25592) );
  AND2X1 U15653 ( .IN1(n14534), .IN2(n8698), .Q(n14533) );
  XOR2X1 U15654 ( .IN1(n14535), .IN2(n8047), .Q(n14534) );
  OR2X1 U15655 ( .IN1(n14530), .IN2(n14528), .Q(n14535) );
  XOR2X1 U15656 ( .IN1(n8047), .IN2(n8048), .Q(n14528) );
  OR2X1 U15657 ( .IN1(n8219), .IN2(n8218), .Q(n14530) );
  AND2X1 U15658 ( .IN1(n8816), .IN2(g222), .Q(n14532) );
  OR2X1 U15659 ( .IN1(n14536), .IN2(n14537), .Q(g25591) );
  AND2X1 U15660 ( .IN1(n8816), .IN2(g209), .Q(n14537) );
  AND2X1 U15661 ( .IN1(n8219), .IN2(n8698), .Q(n14536) );
  AND2X1 U15662 ( .IN1(n14538), .IN2(g6732), .Q(g24355) );
  OR2X1 U15663 ( .IN1(n8804), .IN2(n14539), .Q(n14538) );
  OR2X1 U15664 ( .IN1(n14540), .IN2(n14541), .Q(g24354) );
  AND3X1 U15665 ( .IN1(n8423), .IN2(n14539), .IN3(n8738), .Q(n14541) );
  OR2X1 U15666 ( .IN1(n5531), .IN2(n14542), .Q(n14539) );
  AND2X1 U15667 ( .IN1(n8816), .IN2(g6727), .Q(n14540) );
  OR2X1 U15668 ( .IN1(n14543), .IN2(n14544), .Q(g24353) );
  AND2X1 U15669 ( .IN1(n14545), .IN2(n8698), .Q(n14544) );
  XOR2X1 U15670 ( .IN1(n14542), .IN2(n5531), .Q(n14545) );
  OR4X1 U15671 ( .IN1(n5700), .IN2(n8497), .IN3(n8387), .IN4(n8339), .Q(n14542) );
  AND2X1 U15672 ( .IN1(n8816), .IN2(g6723), .Q(n14543) );
  AND4X1 U15673 ( .IN1(n14546), .IN2(n14547), .IN3(n8387), .IN4(n14548), .Q(
        g24352) );
  AND3X1 U15674 ( .IN1(n8385), .IN2(n8724), .IN3(n8386), .Q(n14548) );
  OR2X1 U15675 ( .IN1(n8339), .IN2(g14828), .Q(n14547) );
  OR2X1 U15676 ( .IN1(test_so80), .IN2(n5700), .Q(n14546) );
  AND2X1 U15677 ( .IN1(n14549), .IN2(g6386), .Q(g24351) );
  OR2X1 U15678 ( .IN1(n8804), .IN2(n14550), .Q(n14549) );
  OR2X1 U15679 ( .IN1(n14551), .IN2(n14552), .Q(g24350) );
  AND3X1 U15680 ( .IN1(n8414), .IN2(n14550), .IN3(n8738), .Q(n14552) );
  OR2X1 U15681 ( .IN1(n8495), .IN2(n14553), .Q(n14550) );
  AND2X1 U15682 ( .IN1(test_so69), .IN2(n8809), .Q(n14551) );
  OR2X1 U15683 ( .IN1(n14554), .IN2(n14555), .Q(g24349) );
  AND2X1 U15684 ( .IN1(n14556), .IN2(n8698), .Q(n14555) );
  XOR2X1 U15685 ( .IN1(n8495), .IN2(n14553), .Q(n14556) );
  OR4X1 U15686 ( .IN1(n5703), .IN2(n5437), .IN3(n8378), .IN4(n8336), .Q(n14553) );
  AND2X1 U15687 ( .IN1(n8816), .IN2(g6377), .Q(n14554) );
  AND4X1 U15688 ( .IN1(n14557), .IN2(n14558), .IN3(n8378), .IN4(n14559), .Q(
        g24348) );
  AND3X1 U15689 ( .IN1(n8376), .IN2(n8724), .IN3(n8377), .Q(n14559) );
  OR2X1 U15690 ( .IN1(n8336), .IN2(g14779), .Q(n14558) );
  OR2X1 U15691 ( .IN1(n5703), .IN2(g12422), .Q(n14557) );
  AND2X1 U15692 ( .IN1(n14560), .IN2(g6040), .Q(g24347) );
  OR2X1 U15693 ( .IN1(n8804), .IN2(n14561), .Q(n14560) );
  OR2X1 U15694 ( .IN1(n14562), .IN2(n14563), .Q(g24346) );
  AND3X1 U15695 ( .IN1(n14561), .IN2(n8512), .IN3(n8738), .Q(n14563) );
  OR2X1 U15696 ( .IN1(n5528), .IN2(n14564), .Q(n14561) );
  AND2X1 U15697 ( .IN1(n8816), .IN2(g6035), .Q(n14562) );
  OR2X1 U15698 ( .IN1(n14565), .IN2(n14566), .Q(g24345) );
  AND2X1 U15699 ( .IN1(n14567), .IN2(n8698), .Q(n14566) );
  XOR2X1 U15700 ( .IN1(n14564), .IN2(n5528), .Q(n14567) );
  OR4X1 U15701 ( .IN1(n5698), .IN2(n5432), .IN3(n8433), .IN4(n8338), .Q(n14564) );
  AND2X1 U15702 ( .IN1(n8816), .IN2(g6031), .Q(n14565) );
  AND4X1 U15703 ( .IN1(n14568), .IN2(n14569), .IN3(n8433), .IN4(n14570), .Q(
        g24344) );
  AND3X1 U15704 ( .IN1(n8431), .IN2(n8725), .IN3(n8432), .Q(n14570) );
  OR2X1 U15705 ( .IN1(n8338), .IN2(g14738), .Q(n14569) );
  OR2X1 U15706 ( .IN1(n5698), .IN2(g12350), .Q(n14568) );
  AND2X1 U15707 ( .IN1(n14571), .IN2(g5694), .Q(g24343) );
  OR2X1 U15708 ( .IN1(n8804), .IN2(n14572), .Q(n14571) );
  OR2X1 U15709 ( .IN1(n14573), .IN2(n14574), .Q(g24342) );
  AND3X1 U15710 ( .IN1(n8424), .IN2(n14572), .IN3(n8739), .Q(n14574) );
  OR2X1 U15711 ( .IN1(n5529), .IN2(n14575), .Q(n14572) );
  AND2X1 U15712 ( .IN1(n8816), .IN2(g5689), .Q(n14573) );
  OR2X1 U15713 ( .IN1(n14576), .IN2(n14577), .Q(g24341) );
  AND2X1 U15714 ( .IN1(n14578), .IN2(n8698), .Q(n14577) );
  XOR2X1 U15715 ( .IN1(n14575), .IN2(n5529), .Q(n14578) );
  OR4X1 U15716 ( .IN1(n5705), .IN2(n5439), .IN3(n8372), .IN4(n8340), .Q(n14575) );
  AND2X1 U15717 ( .IN1(n8816), .IN2(g5685), .Q(n14576) );
  AND4X1 U15718 ( .IN1(n14579), .IN2(n14580), .IN3(n8372), .IN4(n14581), .Q(
        g24340) );
  AND3X1 U15719 ( .IN1(n8370), .IN2(n8725), .IN3(n8371), .Q(n14581) );
  OR2X1 U15720 ( .IN1(n8340), .IN2(g14694), .Q(n14580) );
  OR2X1 U15721 ( .IN1(n5705), .IN2(g12300), .Q(n14579) );
  AND2X1 U15722 ( .IN1(n14582), .IN2(g5348), .Q(g24339) );
  OR2X1 U15723 ( .IN1(n8804), .IN2(n14583), .Q(n14582) );
  OR2X1 U15724 ( .IN1(n14584), .IN2(n14585), .Q(g24338) );
  AND3X1 U15725 ( .IN1(n8444), .IN2(n14583), .IN3(n8739), .Q(n14585) );
  OR2X1 U15726 ( .IN1(n8494), .IN2(n14586), .Q(n14583) );
  AND2X1 U15727 ( .IN1(test_so10), .IN2(n8810), .Q(n14584) );
  OR2X1 U15728 ( .IN1(n14587), .IN2(n14588), .Q(g24337) );
  AND2X1 U15729 ( .IN1(n14589), .IN2(n8698), .Q(n14588) );
  XOR2X1 U15730 ( .IN1(n8494), .IN2(n14586), .Q(n14589) );
  OR4X1 U15731 ( .IN1(n5704), .IN2(n5438), .IN3(n8375), .IN4(n8341), .Q(n14586) );
  AND2X1 U15732 ( .IN1(n8816), .IN2(g5339), .Q(n14587) );
  AND4X1 U15733 ( .IN1(n14590), .IN2(n14591), .IN3(n8375), .IN4(n14592), .Q(
        g24336) );
  AND3X1 U15734 ( .IN1(n8373), .IN2(n8725), .IN3(n8374), .Q(n14592) );
  OR2X1 U15735 ( .IN1(n8341), .IN2(g14662), .Q(n14591) );
  OR2X1 U15736 ( .IN1(n5704), .IN2(g12238), .Q(n14590) );
  OR2X1 U15737 ( .IN1(n14593), .IN2(n14594), .Q(g24335) );
  AND2X1 U15738 ( .IN1(n8816), .IN2(g18881), .Q(n14594) );
  AND3X1 U15739 ( .IN1(n5653), .IN2(g4643), .IN3(n14595), .Q(n14593) );
  OR2X1 U15740 ( .IN1(n14596), .IN2(n14597), .Q(g24334) );
  AND2X1 U15741 ( .IN1(n8816), .IN2(g4358), .Q(n14597) );
  AND4X1 U15742 ( .IN1(n13922), .IN2(n5608), .IN3(n14595), .IN4(n14598), .Q(
        n14596) );
  AND4X1 U15743 ( .IN1(n5274), .IN2(n5539), .IN3(n5303), .IN4(n5365), .Q(
        n14598) );
  AND4X1 U15744 ( .IN1(n8492), .IN2(n8753), .IN3(n5506), .IN4(n14599), .Q(
        n14595) );
  AND3X1 U15745 ( .IN1(n5540), .IN2(n5323), .IN3(n5348), .Q(n14599) );
  AND4X1 U15746 ( .IN1(n5727), .IN2(test_so3), .IN3(g4633), .IN4(g4340), .Q(
        n13922) );
  AND2X1 U15747 ( .IN1(n8816), .IN2(g4392), .Q(g24298) );
  OR2X1 U15748 ( .IN1(n14600), .IN2(n14601), .Q(g24282) );
  AND2X1 U15749 ( .IN1(g24281), .IN2(g9251), .Q(n14601) );
  AND2X1 U15750 ( .IN1(n14602), .IN2(g4308), .Q(n14600) );
  OR2X1 U15751 ( .IN1(n8184), .IN2(n8793), .Q(n14602) );
  AND2X1 U15752 ( .IN1(n8719), .IN2(n8213), .Q(g24281) );
  OR2X1 U15753 ( .IN1(n14603), .IN2(n14604), .Q(g24280) );
  AND2X1 U15754 ( .IN1(n14605), .IN2(g4273), .Q(n14604) );
  OR2X1 U15755 ( .IN1(n14606), .IN2(n14607), .Q(n14605) );
  AND2X1 U15756 ( .IN1(n5763), .IN2(n8697), .Q(n14606) );
  AND2X1 U15757 ( .IN1(n14608), .IN2(g4269), .Q(n14603) );
  OR2X1 U15758 ( .IN1(n8803), .IN2(n14609), .Q(n14608) );
  AND3X1 U15759 ( .IN1(g4264), .IN2(g4258), .IN3(n5764), .Q(n14609) );
  OR2X1 U15760 ( .IN1(n14610), .IN2(n14611), .Q(g24279) );
  AND2X1 U15761 ( .IN1(n14612), .IN2(n8697), .Q(n14611) );
  XNOR2X1 U15762 ( .IN1(n14613), .IN2(n14614), .Q(n14612) );
  OR2X1 U15763 ( .IN1(n14615), .IN2(n14616), .Q(n14613) );
  AND3X1 U15764 ( .IN1(n5726), .IN2(n14617), .IN3(n8291), .Q(n14616) );
  OR4X1 U15765 ( .IN1(g11770), .IN2(g8916), .IN3(g8915), .IN4(n14618), .Q(
        n14617) );
  OR4X1 U15766 ( .IN1(g8920), .IN2(g8919), .IN3(g8918), .IN4(g8917), .Q(n14618) );
  INVX0 U15767 ( .INP(n14619), .ZN(n14615) );
  OR2X1 U15768 ( .IN1(n5726), .IN2(n8291), .Q(n14619) );
  AND2X1 U15769 ( .IN1(n8816), .IN2(g4235), .Q(n14610) );
  AND2X1 U15770 ( .IN1(n14620), .IN2(g4045), .Q(g24278) );
  OR2X1 U15771 ( .IN1(n8803), .IN2(n14621), .Q(n14620) );
  OR2X1 U15772 ( .IN1(n14622), .IN2(n14623), .Q(g24277) );
  AND3X1 U15773 ( .IN1(n8416), .IN2(n14621), .IN3(n8739), .Q(n14623) );
  OR2X1 U15774 ( .IN1(n5530), .IN2(n14624), .Q(n14621) );
  AND2X1 U15775 ( .IN1(n8816), .IN2(g4040), .Q(n14622) );
  OR2X1 U15776 ( .IN1(n14625), .IN2(n14626), .Q(g24276) );
  AND2X1 U15777 ( .IN1(n14627), .IN2(n8697), .Q(n14626) );
  XOR2X1 U15778 ( .IN1(n14624), .IN2(n5530), .Q(n14627) );
  OR4X1 U15779 ( .IN1(n5701), .IN2(n5435), .IN3(n8384), .IN4(n8337), .Q(n14624) );
  AND2X1 U15780 ( .IN1(n8816), .IN2(g4031), .Q(n14625) );
  AND4X1 U15781 ( .IN1(n14628), .IN2(n14629), .IN3(n8384), .IN4(n14630), .Q(
        g24275) );
  AND3X1 U15782 ( .IN1(n8382), .IN2(n8725), .IN3(n8383), .Q(n14630) );
  OR2X1 U15783 ( .IN1(n8337), .IN2(g13966), .Q(n14629) );
  OR2X1 U15784 ( .IN1(n5701), .IN2(g11418), .Q(n14628) );
  AND2X1 U15785 ( .IN1(n14631), .IN2(g3694), .Q(g24274) );
  OR2X1 U15786 ( .IN1(n8803), .IN2(n14632), .Q(n14631) );
  OR2X1 U15787 ( .IN1(n14633), .IN2(n14634), .Q(g24273) );
  AND3X1 U15788 ( .IN1(n8425), .IN2(n14632), .IN3(n8739), .Q(n14634) );
  OR2X1 U15789 ( .IN1(n5532), .IN2(n14635), .Q(n14632) );
  AND2X1 U15790 ( .IN1(n8816), .IN2(g3689), .Q(n14633) );
  OR2X1 U15791 ( .IN1(n14636), .IN2(n14637), .Q(g24272) );
  AND2X1 U15792 ( .IN1(n14638), .IN2(n8697), .Q(n14637) );
  XOR2X1 U15793 ( .IN1(n14635), .IN2(n5532), .Q(n14638) );
  OR4X1 U15794 ( .IN1(n5699), .IN2(n5433), .IN3(n8390), .IN4(n8334), .Q(n14635) );
  AND2X1 U15795 ( .IN1(n8815), .IN2(g3680), .Q(n14636) );
  AND4X1 U15796 ( .IN1(n14639), .IN2(n14640), .IN3(n8390), .IN4(n14641), .Q(
        g24271) );
  AND3X1 U15797 ( .IN1(n8388), .IN2(n8725), .IN3(n8389), .Q(n14641) );
  OR2X1 U15798 ( .IN1(n8334), .IN2(g13926), .Q(n14640) );
  OR2X1 U15799 ( .IN1(n5699), .IN2(g11388), .Q(n14639) );
  AND2X1 U15800 ( .IN1(n14642), .IN2(g3343), .Q(g24270) );
  OR2X1 U15801 ( .IN1(n8803), .IN2(n14643), .Q(n14642) );
  OR2X1 U15802 ( .IN1(n14644), .IN2(n14645), .Q(g24269) );
  AND3X1 U15803 ( .IN1(n8413), .IN2(n14643), .IN3(n8739), .Q(n14645) );
  OR2X1 U15804 ( .IN1(n5527), .IN2(n14646), .Q(n14643) );
  AND2X1 U15805 ( .IN1(n8815), .IN2(g3338), .Q(n14644) );
  OR2X1 U15806 ( .IN1(n14647), .IN2(n14648), .Q(g24268) );
  AND2X1 U15807 ( .IN1(n14649), .IN2(n8697), .Q(n14648) );
  XOR2X1 U15808 ( .IN1(n14646), .IN2(n5527), .Q(n14649) );
  OR4X1 U15809 ( .IN1(n5702), .IN2(n5436), .IN3(n8381), .IN4(n8335), .Q(n14646) );
  AND2X1 U15810 ( .IN1(test_so91), .IN2(n8811), .Q(n14647) );
  AND4X1 U15811 ( .IN1(n14650), .IN2(n14651), .IN3(n8381), .IN4(n14652), .Q(
        g24267) );
  AND3X1 U15812 ( .IN1(n8379), .IN2(n8725), .IN3(n8380), .Q(n14652) );
  OR2X1 U15813 ( .IN1(n8335), .IN2(g13895), .Q(n14651) );
  OR2X1 U15814 ( .IN1(n5702), .IN2(g11349), .Q(n14650) );
  OR2X1 U15815 ( .IN1(n14653), .IN2(n14654), .Q(g24266) );
  AND3X1 U15816 ( .IN1(test_so9), .IN2(n8421), .IN3(n8739), .Q(n14654) );
  AND2X1 U15817 ( .IN1(n8815), .IN2(g2841), .Q(n14653) );
  OR3X1 U15818 ( .IN1(n14655), .IN2(n14656), .IN3(n2787), .Q(g24263) );
  AND2X1 U15819 ( .IN1(n8719), .IN2(n5963), .Q(n2787) );
  AND2X1 U15820 ( .IN1(n8815), .IN2(g2712), .Q(n14656) );
  AND2X1 U15821 ( .IN1(n5299), .IN2(n8697), .Q(n14655) );
  OR3X1 U15822 ( .IN1(n14657), .IN2(n14658), .IN3(n14659), .Q(g24262) );
  AND2X1 U15823 ( .IN1(n14660), .IN2(n8399), .Q(n14659) );
  AND2X1 U15824 ( .IN1(n8815), .IN2(g1548), .Q(n14658) );
  AND3X1 U15825 ( .IN1(n14661), .IN2(g1564), .IN3(n8739), .Q(n14657) );
  OR2X1 U15826 ( .IN1(n14662), .IN2(n11076), .Q(g24261) );
  AND2X1 U15827 ( .IN1(n8815), .IN2(g1585), .Q(n14662) );
  XNOR2X1 U15828 ( .IN1(n8215), .IN2(n14663), .Q(g24260) );
  AND2X1 U15829 ( .IN1(n8719), .IN2(g1548), .Q(n14663) );
  OR2X1 U15830 ( .IN1(n14664), .IN2(n11076), .Q(g24259) );
  AND2X1 U15831 ( .IN1(n8815), .IN2(g1579), .Q(n14664) );
  OR2X1 U15832 ( .IN1(n14665), .IN2(n14666), .Q(g24258) );
  AND2X1 U15833 ( .IN1(n8815), .IN2(g1554), .Q(n14666) );
  AND2X1 U15834 ( .IN1(n8719), .IN2(g496), .Q(n14665) );
  XOR2X1 U15835 ( .IN1(n5616), .IN2(n14667), .Q(g24257) );
  OR2X1 U15836 ( .IN1(n14668), .IN2(n8793), .Q(n14667) );
  OR2X1 U15837 ( .IN1(n14669), .IN2(n14670), .Q(g24256) );
  AND2X1 U15838 ( .IN1(n14671), .IN2(n8697), .Q(n14670) );
  OR2X1 U15839 ( .IN1(n14672), .IN2(n14673), .Q(n14671) );
  AND4X1 U15840 ( .IN1(n8410), .IN2(n14375), .IN3(n8411), .IN4(n14668), .Q(
        n14673) );
  INVX0 U15841 ( .INP(n14674), .ZN(n14672) );
  OR2X1 U15842 ( .IN1(n14668), .IN2(n14675), .Q(n14674) );
  AND3X1 U15843 ( .IN1(n14375), .IN2(n8410), .IN3(n8411), .Q(n14675) );
  AND3X1 U15844 ( .IN1(n5616), .IN2(n5302), .IN3(n5401), .Q(n14375) );
  OR3X1 U15845 ( .IN1(n1302), .IN2(n13998), .IN3(n14676), .Q(n14668) );
  XOR2X1 U15846 ( .IN1(test_so68), .IN2(n8033), .Q(n14676) );
  AND2X1 U15847 ( .IN1(n8815), .IN2(g1339), .Q(n14669) );
  OR3X1 U15848 ( .IN1(n14677), .IN2(n14678), .IN3(n14679), .Q(g24255) );
  AND2X1 U15849 ( .IN1(n11076), .IN2(g17423), .Q(n14679) );
  AND2X1 U15850 ( .IN1(n8815), .IN2(g1589), .Q(n14678) );
  AND3X1 U15851 ( .IN1(n8404), .IN2(g10527), .IN3(n8739), .Q(n14677) );
  AND3X1 U15852 ( .IN1(n8405), .IN2(n8403), .IN3(n14680), .Q(g24254) );
  AND3X1 U15853 ( .IN1(n14681), .IN2(n8725), .IN3(n8404), .Q(n14680) );
  OR3X1 U15854 ( .IN1(n5768), .IN2(n14682), .IN3(n14352), .Q(n14681) );
  INVX0 U15855 ( .INP(n14351), .ZN(n14352) );
  AND2X1 U15856 ( .IN1(g1564), .IN2(n14660), .Q(n14351) );
  INVX0 U15857 ( .INP(n14661), .ZN(n14660) );
  OR2X1 U15858 ( .IN1(n5546), .IN2(n8215), .Q(n14661) );
  AND2X1 U15859 ( .IN1(n14379), .IN2(n13818), .Q(n14682) );
  INVX0 U15860 ( .INP(n1302), .ZN(n13818) );
  OR2X1 U15861 ( .IN1(g1351), .IN2(g1312), .Q(n1302) );
  INVX0 U15862 ( .INP(n13998), .ZN(n14379) );
  OR2X1 U15863 ( .IN1(n12640), .IN2(n13738), .Q(n13998) );
  XOR2X1 U15864 ( .IN1(g1339), .IN2(n8496), .Q(n13738) );
  AND2X1 U15865 ( .IN1(n8496), .IN2(n5616), .Q(n12640) );
  OR2X1 U15866 ( .IN1(n14683), .IN2(n14684), .Q(g24253) );
  AND2X1 U15867 ( .IN1(n14685), .IN2(n8697), .Q(n14684) );
  OR2X1 U15868 ( .IN1(n14686), .IN2(n14687), .Q(n14685) );
  AND2X1 U15869 ( .IN1(g7946), .IN2(g1521), .Q(n14687) );
  AND2X1 U15870 ( .IN1(n5302), .IN2(g1532), .Q(n14686) );
  AND2X1 U15871 ( .IN1(n8815), .IN2(g1306), .Q(n14683) );
  OR3X1 U15872 ( .IN1(n14688), .IN2(n14689), .IN3(n14360), .Q(g24252) );
  AND3X1 U15873 ( .IN1(g1339), .IN2(g7946), .IN3(n8740), .Q(n14360) );
  AND3X1 U15874 ( .IN1(n5302), .IN2(g1521), .IN3(n8740), .Q(n14689) );
  AND2X1 U15875 ( .IN1(test_so49), .IN2(n8809), .Q(n14688) );
  OR2X1 U15876 ( .IN1(n14690), .IN2(n14691), .Q(g24251) );
  AND2X1 U15877 ( .IN1(test_so12), .IN2(n14692), .Q(n14691) );
  AND2X1 U15878 ( .IN1(n13141), .IN2(g1442), .Q(n14690) );
  OR2X1 U15879 ( .IN1(n14693), .IN2(n14694), .Q(g24250) );
  AND2X1 U15880 ( .IN1(n14692), .IN2(g1489), .Q(n14694) );
  AND2X1 U15881 ( .IN1(test_so12), .IN2(n13141), .Q(n14693) );
  OR2X1 U15882 ( .IN1(n14695), .IN2(n14696), .Q(g24249) );
  AND2X1 U15883 ( .IN1(n14697), .IN2(g1489), .Q(n14696) );
  OR2X1 U15884 ( .IN1(n14698), .IN2(n13141), .Q(n14697) );
  INVX0 U15885 ( .INP(n14692), .ZN(n13141) );
  OR2X1 U15886 ( .IN1(n8802), .IN2(n13143), .Q(n14692) );
  AND2X1 U15887 ( .IN1(n8718), .IN2(n8523), .Q(n14698) );
  AND3X1 U15888 ( .IN1(n8222), .IN2(n8725), .IN3(n13143), .Q(n14695) );
  AND3X1 U15889 ( .IN1(n8490), .IN2(g13272), .IN3(n5364), .Q(n13143) );
  OR3X1 U15890 ( .IN1(n14699), .IN2(n14700), .IN3(n14701), .Q(g24248) );
  XOR2X1 U15891 ( .IN1(g1404), .IN2(n14702), .Q(n14701) );
  AND2X1 U15892 ( .IN1(n5655), .IN2(n8697), .Q(n14702) );
  AND2X1 U15893 ( .IN1(n5401), .IN2(n8697), .Q(n14700) );
  AND2X1 U15894 ( .IN1(n11076), .IN2(g1395), .Q(n14699) );
  AND2X1 U15895 ( .IN1(n11076), .IN2(n8440), .Q(g24247) );
  AND2X1 U15896 ( .IN1(g12923), .IN2(n8696), .Q(n11076) );
  OR3X1 U15897 ( .IN1(n14703), .IN2(n14704), .IN3(n14705), .Q(g24246) );
  AND2X1 U15898 ( .IN1(n14706), .IN2(n8400), .Q(n14705) );
  AND2X1 U15899 ( .IN1(n8815), .IN2(g1205), .Q(n14704) );
  AND3X1 U15900 ( .IN1(n14707), .IN2(g1221), .IN3(n8740), .Q(n14703) );
  OR2X1 U15901 ( .IN1(n14708), .IN2(n11091), .Q(g24245) );
  AND2X1 U15902 ( .IN1(n8815), .IN2(g30332), .Q(n14708) );
  XNOR2X1 U15903 ( .IN1(n8214), .IN2(n14709), .Q(g24244) );
  AND2X1 U15904 ( .IN1(n8718), .IN2(g1205), .Q(n14709) );
  OR2X1 U15905 ( .IN1(n14710), .IN2(n11091), .Q(g24243) );
  AND2X1 U15906 ( .IN1(n8815), .IN2(g1236), .Q(n14710) );
  OR2X1 U15907 ( .IN1(n14711), .IN2(n14712), .Q(g24242) );
  AND2X1 U15908 ( .IN1(test_so76), .IN2(n8809), .Q(n14712) );
  AND2X1 U15909 ( .IN1(n8718), .IN2(g29215), .Q(n14711) );
  XOR2X1 U15910 ( .IN1(n5622), .IN2(n14713), .Q(g24241) );
  OR2X1 U15911 ( .IN1(n14714), .IN2(n8794), .Q(n14713) );
  OR2X1 U15912 ( .IN1(n14715), .IN2(n14716), .Q(g24240) );
  AND2X1 U15913 ( .IN1(n14717), .IN2(n8696), .Q(n14716) );
  OR2X1 U15914 ( .IN1(n14718), .IN2(n14719), .Q(n14717) );
  AND4X1 U15915 ( .IN1(n8417), .IN2(n14423), .IN3(n8418), .IN4(n14714), .Q(
        n14719) );
  INVX0 U15916 ( .INP(n14720), .ZN(n14718) );
  OR2X1 U15917 ( .IN1(n14714), .IN2(n14721), .Q(n14720) );
  AND3X1 U15918 ( .IN1(n14423), .IN2(n8417), .IN3(n8418), .Q(n14721) );
  AND3X1 U15919 ( .IN1(n5622), .IN2(n5304), .IN3(n5392), .Q(n14423) );
  OR3X1 U15920 ( .IN1(n4837), .IN2(n14722), .IN3(n14032), .Q(n14714) );
  XOR2X1 U15921 ( .IN1(n8032), .IN2(g979), .Q(n14722) );
  AND2X1 U15922 ( .IN1(n8815), .IN2(g996), .Q(n14715) );
  OR3X1 U15923 ( .IN1(n14723), .IN2(n14724), .IN3(n14725), .Q(g24239) );
  AND2X1 U15924 ( .IN1(n11091), .IN2(g17400), .Q(n14725) );
  AND2X1 U15925 ( .IN1(n8815), .IN2(g1246), .Q(n14724) );
  AND3X1 U15926 ( .IN1(n8368), .IN2(g10500), .IN3(n8740), .Q(n14723) );
  AND3X1 U15927 ( .IN1(n8369), .IN2(n8368), .IN3(n14726), .Q(g24238) );
  AND3X1 U15928 ( .IN1(n8727), .IN2(n8509), .IN3(n14727), .Q(n14726) );
  INVX0 U15929 ( .INP(n14728), .ZN(n14727) );
  AND3X1 U15930 ( .IN1(n14729), .IN2(n14401), .IN3(test_so76), .Q(n14728) );
  AND2X1 U15931 ( .IN1(g1221), .IN2(n14706), .Q(n14401) );
  INVX0 U15932 ( .INP(n14707), .ZN(n14706) );
  OR2X1 U15933 ( .IN1(n5547), .IN2(n8214), .Q(n14707) );
  OR2X1 U15934 ( .IN1(n14032), .IN2(n4837), .Q(n14729) );
  OR2X1 U15935 ( .IN1(test_so20), .IN2(g1008), .Q(n4837) );
  OR2X1 U15936 ( .IN1(n12674), .IN2(n13750), .Q(n14032) );
  XOR2X1 U15937 ( .IN1(g996), .IN2(n5320), .Q(n13750) );
  AND2X1 U15938 ( .IN1(n5320), .IN2(n5622), .Q(n12674) );
  OR2X1 U15939 ( .IN1(n14730), .IN2(n14731), .Q(g24237) );
  AND2X1 U15940 ( .IN1(n14732), .IN2(n8696), .Q(n14731) );
  OR2X1 U15941 ( .IN1(n14733), .IN2(n14734), .Q(n14732) );
  AND2X1 U15942 ( .IN1(g7916), .IN2(g1178), .Q(n14734) );
  AND2X1 U15943 ( .IN1(n5304), .IN2(g1189), .Q(n14733) );
  AND2X1 U15944 ( .IN1(n8815), .IN2(g962), .Q(n14730) );
  OR2X1 U15945 ( .IN1(n14735), .IN2(n14736), .Q(g24236) );
  AND2X1 U15946 ( .IN1(n14737), .IN2(n8696), .Q(n14736) );
  OR2X1 U15947 ( .IN1(n14738), .IN2(n14739), .Q(n14737) );
  AND2X1 U15948 ( .IN1(g7916), .IN2(g996), .Q(n14739) );
  AND2X1 U15949 ( .IN1(n5304), .IN2(g1178), .Q(n14738) );
  AND2X1 U15950 ( .IN1(n8815), .IN2(g1183), .Q(n14735) );
  OR2X1 U15951 ( .IN1(n14740), .IN2(n14741), .Q(g24235) );
  AND2X1 U15952 ( .IN1(n14742), .IN2(g1152), .Q(n14741) );
  AND2X1 U15953 ( .IN1(n13176), .IN2(test_so7), .Q(n14740) );
  OR2X1 U15954 ( .IN1(n14743), .IN2(n14744), .Q(g24234) );
  AND2X1 U15955 ( .IN1(n14742), .IN2(g1146), .Q(n14744) );
  AND2X1 U15956 ( .IN1(n13176), .IN2(g1152), .Q(n14743) );
  OR2X1 U15957 ( .IN1(n14745), .IN2(n14746), .Q(g24233) );
  AND2X1 U15958 ( .IN1(n14747), .IN2(g1146), .Q(n14746) );
  OR2X1 U15959 ( .IN1(n14748), .IN2(n13176), .Q(n14747) );
  INVX0 U15960 ( .INP(n14742), .ZN(n13176) );
  OR2X1 U15961 ( .IN1(n8801), .IN2(n13178), .Q(n14742) );
  AND2X1 U15962 ( .IN1(n5618), .IN2(n8696), .Q(n14748) );
  AND3X1 U15963 ( .IN1(n8727), .IN2(n8518), .IN3(n13178), .Q(n14745) );
  AND3X1 U15964 ( .IN1(g13259), .IN2(n5363), .IN3(n5599), .Q(n13178) );
  OR3X1 U15965 ( .IN1(n14749), .IN2(n14750), .IN3(n14751), .Q(g24232) );
  XOR2X1 U15966 ( .IN1(g1061), .IN2(n14752), .Q(n14751) );
  AND2X1 U15967 ( .IN1(n5654), .IN2(n8696), .Q(n14752) );
  AND2X1 U15968 ( .IN1(n5392), .IN2(n8696), .Q(n14750) );
  AND2X1 U15969 ( .IN1(n11091), .IN2(g1052), .Q(n14749) );
  AND2X1 U15970 ( .IN1(n11091), .IN2(n8441), .Q(g24231) );
  AND2X1 U15971 ( .IN1(g12919), .IN2(n8696), .Q(n11091) );
  OR2X1 U15972 ( .IN1(n14753), .IN2(n14754), .Q(g24216) );
  AND2X1 U15973 ( .IN1(n14755), .IN2(g854), .Q(n14754) );
  AND2X1 U15974 ( .IN1(n13236), .IN2(g847), .Q(n14753) );
  OR2X1 U15975 ( .IN1(n14756), .IN2(n14757), .Q(g24215) );
  AND2X1 U15976 ( .IN1(n14758), .IN2(g703), .Q(n14757) );
  OR2X1 U15977 ( .IN1(n8801), .IN2(n14759), .Q(n14758) );
  AND2X1 U15978 ( .IN1(n5562), .IN2(n14075), .Q(n14759) );
  AND2X1 U15979 ( .IN1(g847), .IN2(n4948), .Q(n14075) );
  AND2X1 U15980 ( .IN1(n14760), .IN2(g837), .Q(n14756) );
  OR2X1 U15981 ( .IN1(n14761), .IN2(n13236), .Q(n14760) );
  AND3X1 U15982 ( .IN1(n14762), .IN2(n8726), .IN3(n14763), .Q(n14761) );
  OR2X1 U15983 ( .IN1(n5728), .IN2(n8216), .Q(n14763) );
  OR3X1 U15984 ( .IN1(n14764), .IN2(n14765), .IN3(n14766), .Q(g24214) );
  AND2X1 U15985 ( .IN1(n14767), .IN2(g703), .Q(n14766) );
  OR2X1 U15986 ( .IN1(n14768), .IN2(n13236), .Q(n14767) );
  AND2X1 U15987 ( .IN1(n14769), .IN2(n8696), .Q(n14768) );
  OR2X1 U15988 ( .IN1(n5562), .IN2(n14762), .Q(n14769) );
  OR2X1 U15989 ( .IN1(n5709), .IN2(n5733), .Q(n14762) );
  AND4X1 U15990 ( .IN1(n13237), .IN2(g822), .IN3(n14770), .IN4(n5709), .Q(
        n14765) );
  AND2X1 U15991 ( .IN1(g817), .IN2(g723), .Q(n14770) );
  AND2X1 U15992 ( .IN1(n8815), .IN2(g847), .Q(n14764) );
  OR2X1 U15993 ( .IN1(n14771), .IN2(g24212), .Q(g24213) );
  AND2X1 U15994 ( .IN1(n8815), .IN2(g753), .Q(n14771) );
  OR2X1 U15995 ( .IN1(n14772), .IN2(n14773), .Q(g24211) );
  AND2X1 U15996 ( .IN1(n8815), .IN2(g546), .Q(n14773) );
  AND2X1 U15997 ( .IN1(n2404), .IN2(n14774), .Q(n14772) );
  OR2X1 U15998 ( .IN1(n5520), .IN2(test_so41), .Q(n14774) );
  AND3X1 U15999 ( .IN1(n14775), .IN2(n8725), .IN3(n11635), .Q(g24210) );
  AND3X1 U16000 ( .IN1(g203), .IN2(g518), .IN3(n5548), .Q(n11635) );
  OR2X1 U16001 ( .IN1(n14776), .IN2(n14777), .Q(n14775) );
  AND2X1 U16002 ( .IN1(g174), .IN2(g168), .Q(n14777) );
  AND2X1 U16003 ( .IN1(test_so72), .IN2(n14778), .Q(n14776) );
  OR2X1 U16004 ( .IN1(g174), .IN2(g168), .Q(n14778) );
  OR2X1 U16005 ( .IN1(n14779), .IN2(n14780), .Q(g24209) );
  AND2X1 U16006 ( .IN1(n13237), .IN2(g446), .Q(n14780) );
  AND2X1 U16007 ( .IN1(n13236), .IN2(g417), .Q(n14779) );
  OR3X1 U16008 ( .IN1(n14781), .IN2(n14782), .IN3(n14783), .Q(g24208) );
  AND2X1 U16009 ( .IN1(n8815), .IN2(g424), .Q(n14783) );
  AND2X1 U16010 ( .IN1(n13237), .IN2(g246), .Q(n14782) );
  AND2X1 U16011 ( .IN1(n13236), .IN2(g475), .Q(n14781) );
  OR2X1 U16012 ( .IN1(n14784), .IN2(n14785), .Q(g24207) );
  AND2X1 U16013 ( .IN1(n14755), .IN2(g475), .Q(n14785) );
  AND2X1 U16014 ( .IN1(n13236), .IN2(g441), .Q(n14784) );
  OR2X1 U16015 ( .IN1(n14786), .IN2(n14787), .Q(g24206) );
  AND2X1 U16016 ( .IN1(n14755), .IN2(g441), .Q(n14787) );
  AND2X1 U16017 ( .IN1(n13236), .IN2(g437), .Q(n14786) );
  OR3X1 U16018 ( .IN1(n14788), .IN2(n14789), .IN3(n14790), .Q(g24205) );
  AND2X1 U16019 ( .IN1(n8814), .IN2(g437), .Q(n14790) );
  AND2X1 U16020 ( .IN1(n13237), .IN2(g269), .Q(n14789) );
  AND2X1 U16021 ( .IN1(test_so23), .IN2(n13236), .Q(n14788) );
  OR2X1 U16022 ( .IN1(n14791), .IN2(n14792), .Q(g24204) );
  AND2X1 U16023 ( .IN1(test_so23), .IN2(n14755), .Q(n14792) );
  AND2X1 U16024 ( .IN1(n13236), .IN2(g429), .Q(n14791) );
  OR2X1 U16025 ( .IN1(n14793), .IN2(n14794), .Q(g24203) );
  AND2X1 U16026 ( .IN1(n14755), .IN2(g429), .Q(n14794) );
  AND2X1 U16027 ( .IN1(n13236), .IN2(g401), .Q(n14793) );
  OR2X1 U16028 ( .IN1(n14795), .IN2(n14796), .Q(g24202) );
  AND2X1 U16029 ( .IN1(n14755), .IN2(g411), .Q(n14796) );
  AND2X1 U16030 ( .IN1(n13236), .IN2(g424), .Q(n14795) );
  OR2X1 U16031 ( .IN1(n14797), .IN2(n14798), .Q(g24201) );
  AND2X1 U16032 ( .IN1(n14755), .IN2(g392), .Q(n14798) );
  AND2X1 U16033 ( .IN1(n13236), .IN2(g405), .Q(n14797) );
  OR3X1 U16034 ( .IN1(n14799), .IN2(n14800), .IN3(n14801), .Q(g24200) );
  AND2X1 U16035 ( .IN1(n8814), .IN2(g401), .Q(n14801) );
  AND2X1 U16036 ( .IN1(n13236), .IN2(g392), .Q(n14800) );
  INVX0 U16037 ( .INP(n14755), .ZN(n13236) );
  OR2X1 U16038 ( .IN1(n4948), .IN2(n8794), .Q(n14755) );
  AND3X1 U16039 ( .IN1(n5821), .IN2(g854), .IN3(n13237), .Q(n14799) );
  AND2X1 U16040 ( .IN1(n8718), .IN2(n4948), .Q(n13237) );
  AND2X1 U16041 ( .IN1(n8459), .IN2(n8350), .Q(g23190) );
  OR2X1 U16042 ( .IN1(n14802), .IN2(n14803), .Q(g21901) );
  AND2X1 U16043 ( .IN1(n14804), .IN2(n8696), .Q(n14803) );
  OR2X1 U16044 ( .IN1(n14805), .IN2(n14806), .Q(n14804) );
  AND2X1 U16045 ( .IN1(n5380), .IN2(n14807), .Q(n14806) );
  OR2X1 U16046 ( .IN1(n14808), .IN2(g8786), .Q(n14807) );
  AND4X1 U16047 ( .IN1(n8322), .IN2(n8321), .IN3(n8323), .IN4(n14809), .Q(
        n14808) );
  AND4X1 U16048 ( .IN1(DFF_480_n1), .IN2(DFF_909_n1), .IN3(n8320), .IN4(
        DFF_1234_n1), .Q(n14809) );
  AND2X1 U16049 ( .IN1(n5694), .IN2(g4180), .Q(n14805) );
  AND2X1 U16050 ( .IN1(n8814), .IN2(g2946), .Q(n14802) );
  OR2X1 U16051 ( .IN1(n14810), .IN2(n14811), .Q(g21900) );
  AND3X1 U16052 ( .IN1(n8420), .IN2(n8419), .IN3(n8741), .Q(n14811) );
  AND2X1 U16053 ( .IN1(n8814), .IN2(g4239), .Q(n14810) );
  XNOR2X1 U16054 ( .IN1(n8211), .IN2(n14812), .Q(g21899) );
  AND2X1 U16055 ( .IN1(n8718), .IN2(g9019), .Q(n14812) );
  OR2X1 U16056 ( .IN1(n14813), .IN2(n14814), .Q(g21898) );
  INVX0 U16057 ( .INP(n14815), .ZN(n14814) );
  OR2X1 U16058 ( .IN1(n8677), .IN2(n8034), .Q(n14815) );
  AND2X1 U16059 ( .IN1(n8211), .IN2(n8695), .Q(n14813) );
  XNOR2X1 U16060 ( .IN1(n8212), .IN2(n14816), .Q(g21897) );
  AND2X1 U16061 ( .IN1(n8718), .IN2(g8839), .Q(n14816) );
  OR2X1 U16062 ( .IN1(n14817), .IN2(n14818), .Q(g21896) );
  AND2X1 U16063 ( .IN1(n8814), .IN2(g4245), .Q(n14818) );
  AND2X1 U16064 ( .IN1(n8212), .IN2(n8695), .Q(n14817) );
  OR2X1 U16065 ( .IN1(n14819), .IN2(n14820), .Q(g21895) );
  AND2X1 U16066 ( .IN1(n14607), .IN2(g4269), .Q(n14820) );
  OR2X1 U16067 ( .IN1(n14821), .IN2(g21893), .Q(n14607) );
  AND2X1 U16068 ( .IN1(n5823), .IN2(n8695), .Q(n14821) );
  AND2X1 U16069 ( .IN1(n14822), .IN2(g4264), .Q(n14819) );
  OR2X1 U16070 ( .IN1(n8801), .IN2(n14823), .Q(n14822) );
  AND2X1 U16071 ( .IN1(n5763), .IN2(g4258), .Q(n14823) );
  OR2X1 U16072 ( .IN1(n14824), .IN2(n14825), .Q(g21894) );
  AND2X1 U16073 ( .IN1(g21893), .IN2(g4264), .Q(n14825) );
  AND2X1 U16074 ( .IN1(n14826), .IN2(g4258), .Q(n14824) );
  OR2X1 U16075 ( .IN1(n5823), .IN2(n8794), .Q(n14826) );
  AND2X1 U16076 ( .IN1(n8712), .IN2(n8428), .Q(g21893) );
  OR2X1 U16077 ( .IN1(n14827), .IN2(n14828), .Q(g21892) );
  AND2X1 U16078 ( .IN1(n8814), .IN2(g4273), .Q(n14828) );
  AND2X1 U16079 ( .IN1(n8027), .IN2(n8702), .Q(n14827) );
  OR2X1 U16080 ( .IN1(n14829), .IN2(n14830), .Q(g21891) );
  AND2X1 U16081 ( .IN1(n14614), .IN2(n8677), .Q(n14830) );
  OR2X1 U16082 ( .IN1(n14831), .IN2(n14832), .Q(n14614) );
  AND2X1 U16083 ( .IN1(n8186), .IN2(n5484), .Q(n14832) );
  AND2X1 U16084 ( .IN1(n8187), .IN2(g4253), .Q(n14831) );
  AND2X1 U16085 ( .IN1(n8818), .IN2(g4180), .Q(n14829) );
  AND2X1 U16086 ( .IN1(n8812), .IN2(n9240), .Q(g21727) );
  AND2X1 U16087 ( .IN1(n8822), .IN2(g2975), .Q(g18597) );
  INVX0 U16088 ( .INP(g5), .ZN(g12833) );
  OR2X1 U5116_U1 ( .IN1(g34783), .IN2(n297), .Q(g34221) );
  OR2X1 U5126_U1 ( .IN1(n1302), .IN2(n184), .Q(n4895) );
  OR2X1 U5127_U1 ( .IN1(n4837), .IN2(n201), .Q(n4920) );
  OR2X1 U5128_U1 ( .IN1(n2787), .IN2(n1169), .Q(n5045) );
  OR2X1 U5129_U1 ( .IN1(g559), .IN2(g9048), .Q(n4959) );
  INVX0 U5353_U2 ( .INP(n8479), .ZN(U5353_n1) );
  AND2X1 U5353_U1 ( .IN1(n5960), .IN2(U5353_n1), .Q(n4689) );
  INVX0 U5355_U2 ( .INP(n8474), .ZN(U5355_n1) );
  AND2X1 U5355_U1 ( .IN1(n5961), .IN2(U5355_n1), .Q(n4708) );
  INVX0 U5961_U2 ( .INP(n730), .ZN(U5961_n1) );
  AND2X1 U5961_U1 ( .IN1(n3593), .IN2(U5961_n1), .Q(n3595) );
  INVX0 U5962_U2 ( .INP(n1281), .ZN(U5962_n1) );
  AND2X1 U5962_U1 ( .IN1(n3574), .IN2(U5962_n1), .Q(n3576) );
  INVX0 U5963_U2 ( .INP(n1283), .ZN(U5963_n1) );
  AND2X1 U5963_U1 ( .IN1(n3517), .IN2(U5963_n1), .Q(n3519) );
  INVX0 U5964_U2 ( .INP(n1633), .ZN(U5964_n1) );
  AND2X1 U5964_U1 ( .IN1(n3628), .IN2(U5964_n1), .Q(n3630) );
  INVX0 U5965_U2 ( .INP(n1279), .ZN(U5965_n1) );
  AND2X1 U5965_U1 ( .IN1(n3555), .IN2(U5965_n1), .Q(n3557) );
  INVX0 U5966_U2 ( .INP(n725), .ZN(U5966_n1) );
  AND2X1 U5966_U1 ( .IN1(n3646), .IN2(U5966_n1), .Q(n3648) );
  INVX0 U5967_U2 ( .INP(n1285), .ZN(U5967_n1) );
  AND2X1 U5967_U1 ( .IN1(n3536), .IN2(U5967_n1), .Q(n3538) );
  INVX0 U5968_U2 ( .INP(n728), .ZN(U5968_n1) );
  AND2X1 U5968_U1 ( .IN1(n3611), .IN2(U5968_n1), .Q(n3613) );
  AND2X1 U6100_U2 ( .IN1(n3635), .IN2(U6100_n1), .Q(n4888) );
  INVX0 U6100_U1 ( .INP(n8807), .ZN(U6100_n1) );
  INVX0 U6211_U2 ( .INP(n1635), .ZN(U6211_n1) );
  AND2X1 U6211_U1 ( .IN1(n3623), .IN2(U6211_n1), .Q(n3622) );
  INVX0 U6212_U2 ( .INP(n729), .ZN(U6212_n1) );
  AND2X1 U6212_U1 ( .IN1(n3587), .IN2(U6212_n1), .Q(n3586) );
  INVX0 U6213_U2 ( .INP(n727), .ZN(U6213_n1) );
  AND2X1 U6213_U1 ( .IN1(n3605), .IN2(U6213_n1), .Q(n3604) );
  INVX0 U6214_U2 ( .INP(n1280), .ZN(U6214_n1) );
  AND2X1 U6214_U1 ( .IN1(n3568), .IN2(U6214_n1), .Q(n3567) );
  INVX0 U6215_U2 ( .INP(n1278), .ZN(U6215_n1) );
  AND2X1 U6215_U1 ( .IN1(n3549), .IN2(U6215_n1), .Q(n3548) );
  INVX0 U6216_U2 ( .INP(n1282), .ZN(U6216_n1) );
  AND2X1 U6216_U1 ( .IN1(n3512), .IN2(U6216_n1), .Q(n3511) );
  INVX0 U6217_U2 ( .INP(n1284), .ZN(U6217_n1) );
  AND2X1 U6217_U1 ( .IN1(n3531), .IN2(U6217_n1), .Q(n3530) );
  INVX0 U6218_U2 ( .INP(n724), .ZN(U6218_n1) );
  AND2X1 U6218_U1 ( .IN1(n3641), .IN2(U6218_n1), .Q(n3640) );
  INVX0 U6279_U2 ( .INP(n5337), .ZN(U6279_n1) );
  AND2X1 U6279_U1 ( .IN1(n4537), .IN2(U6279_n1), .Q(n4201) );
  INVX0 U6280_U2 ( .INP(n5336), .ZN(U6280_n1) );
  AND2X1 U6280_U1 ( .IN1(n4201), .IN2(U6280_n1), .Q(n3745) );
  INVX0 U6281_U2 ( .INP(n5294), .ZN(U6281_n1) );
  AND2X1 U6281_U1 ( .IN1(n3745), .IN2(U6281_n1), .Q(n3684) );
  INVX0 U6282_U2 ( .INP(n5552), .ZN(U6282_n1) );
  AND2X1 U6282_U1 ( .IN1(n3684), .IN2(U6282_n1), .Q(n3274) );
  INVX0 U6283_U2 ( .INP(n5472), .ZN(U6283_n1) );
  AND2X1 U6283_U1 ( .IN1(n3274), .IN2(U6283_n1), .Q(n2982) );
  INVX0 U6284_U2 ( .INP(n5476), .ZN(U6284_n1) );
  AND2X1 U6284_U1 ( .IN1(n2982), .IN2(U6284_n1), .Q(n2706) );
  INVX0 U6285_U2 ( .INP(n5550), .ZN(U6285_n1) );
  AND2X1 U6285_U1 ( .IN1(n2706), .IN2(U6285_n1), .Q(n2649) );
  INVX0 U6286_U2 ( .INP(n5473), .ZN(U6286_n1) );
  AND2X1 U6286_U1 ( .IN1(n2649), .IN2(U6286_n1), .Q(n2556) );
  INVX0 U6287_U2 ( .INP(n5475), .ZN(U6287_n1) );
  AND2X1 U6287_U1 ( .IN1(n2556), .IN2(U6287_n1), .Q(n2509) );
  INVX0 U6288_U2 ( .INP(n5474), .ZN(U6288_n1) );
  AND2X1 U6288_U1 ( .IN1(n2509), .IN2(U6288_n1), .Q(n2487) );
  INVX0 U6289_U2 ( .INP(n5339), .ZN(U6289_n1) );
  AND2X1 U6289_U1 ( .IN1(n2487), .IN2(U6289_n1), .Q(n2427) );
  INVX0 U6290_U2 ( .INP(n5672), .ZN(U6290_n1) );
  AND2X1 U6290_U1 ( .IN1(n2427), .IN2(U6290_n1), .Q(n2423) );
  INVX0 U6291_U2 ( .INP(n5335), .ZN(U6291_n1) );
  AND2X1 U6291_U1 ( .IN1(n4826), .IN2(U6291_n1), .Q(n4537) );
  AND2X1 U6292_U2 ( .IN1(n4959), .IN2(U6292_n1), .Q(n2421) );
  INVX0 U6292_U1 ( .INP(n8808), .ZN(U6292_n1) );
  AND2X1 U6338_U2 ( .IN1(n1574), .IN2(U6338_n1), .Q(n3765) );
  INVX0 U6338_U1 ( .INP(n8807), .ZN(U6338_n1) );
  INVX0 U6341_U2 ( .INP(n1069), .ZN(U6341_n1) );
  AND2X1 U6341_U1 ( .IN1(n3765), .IN2(U6341_n1), .Q(n3951) );
  INVX0 U6342_U2 ( .INP(n704), .ZN(U6342_n1) );
  AND2X1 U6342_U1 ( .IN1(n3765), .IN2(U6342_n1), .Q(n3774) );
  INVX0 U6343_U2 ( .INP(n1011), .ZN(U6343_n1) );
  AND2X1 U6343_U1 ( .IN1(n3765), .IN2(U6343_n1), .Q(n3842) );
  INVX0 U6344_U2 ( .INP(n952), .ZN(U6344_n1) );
  AND2X1 U6344_U1 ( .IN1(n3765), .IN2(U6344_n1), .Q(n3808) );
  INVX0 U6345_U2 ( .INP(n699), .ZN(U6345_n1) );
  AND2X1 U6345_U1 ( .IN1(n3765), .IN2(U6345_n1), .Q(n3908) );
  INVX0 U6346_U2 ( .INP(n94), .ZN(U6346_n1) );
  AND2X1 U6346_U1 ( .IN1(n3765), .IN2(U6346_n1), .Q(n3984) );
  INVX0 U6347_U2 ( .INP(n473), .ZN(U6347_n1) );
  AND2X1 U6347_U1 ( .IN1(n3765), .IN2(U6347_n1), .Q(n3875) );
  INVX0 U6348_U2 ( .INP(n106), .ZN(U6348_n1) );
  AND2X1 U6348_U1 ( .IN1(n3765), .IN2(U6348_n1), .Q(n4015) );
  INVX0 U6349_U2 ( .INP(n3446), .ZN(U6349_n1) );
  AND2X1 U6349_U1 ( .IN1(n3765), .IN2(U6349_n1), .Q(n3914) );
  INVX0 U6350_U2 ( .INP(n3406), .ZN(U6350_n1) );
  AND2X1 U6350_U1 ( .IN1(n3765), .IN2(U6350_n1), .Q(n3780) );
  INVX0 U6351_U2 ( .INP(n3481), .ZN(U6351_n1) );
  AND2X1 U6351_U1 ( .IN1(n3765), .IN2(U6351_n1), .Q(n3957) );
  INVX0 U6352_U2 ( .INP(n3426), .ZN(U6352_n1) );
  AND2X1 U6352_U1 ( .IN1(n3765), .IN2(U6352_n1), .Q(n3848) );
  INVX0 U6353_U2 ( .INP(n3491), .ZN(U6353_n1) );
  AND2X1 U6353_U1 ( .IN1(n3765), .IN2(U6353_n1), .Q(n3990) );
  INVX0 U6354_U2 ( .INP(n3416), .ZN(U6354_n1) );
  AND2X1 U6354_U1 ( .IN1(n3765), .IN2(U6354_n1), .Q(n3814) );
  INVX0 U6355_U2 ( .INP(n3436), .ZN(U6355_n1) );
  AND2X1 U6355_U1 ( .IN1(n3765), .IN2(U6355_n1), .Q(n3881) );
  INVX0 U6356_U2 ( .INP(n3502), .ZN(U6356_n1) );
  AND2X1 U6356_U1 ( .IN1(n3765), .IN2(U6356_n1), .Q(n4022) );
  INVX0 U6357_U2 ( .INP(n3501), .ZN(U6357_n1) );
  AND2X1 U6357_U1 ( .IN1(n3765), .IN2(U6357_n1), .Q(n4027) );
  INVX0 U6358_U2 ( .INP(n3407), .ZN(U6358_n1) );
  AND2X1 U6358_U1 ( .IN1(n3765), .IN2(U6358_n1), .Q(n3785) );
  INVX0 U6359_U2 ( .INP(n3482), .ZN(U6359_n1) );
  AND2X1 U6359_U1 ( .IN1(n3765), .IN2(U6359_n1), .Q(n3962) );
  INVX0 U6360_U2 ( .INP(n3427), .ZN(U6360_n1) );
  AND2X1 U6360_U1 ( .IN1(n3765), .IN2(U6360_n1), .Q(n3853) );
  INVX0 U6361_U2 ( .INP(n3437), .ZN(U6361_n1) );
  AND2X1 U6361_U1 ( .IN1(n3765), .IN2(U6361_n1), .Q(n3886) );
  INVX0 U6362_U2 ( .INP(n3417), .ZN(U6362_n1) );
  AND2X1 U6362_U1 ( .IN1(n3765), .IN2(U6362_n1), .Q(n3819) );
  INVX0 U6363_U2 ( .INP(n3492), .ZN(U6363_n1) );
  AND2X1 U6363_U1 ( .IN1(n3765), .IN2(U6363_n1), .Q(n3995) );
  INVX0 U6364_U2 ( .INP(n3447), .ZN(U6364_n1) );
  AND2X1 U6364_U1 ( .IN1(n3765), .IN2(U6364_n1), .Q(n3919) );
  INVX0 U6365_U2 ( .INP(n5471), .ZN(U6365_n1) );
  AND2X1 U6365_U1 ( .IN1(n3682), .IN2(U6365_n1), .Q(n3272) );
  INVX0 U6366_U2 ( .INP(n5331), .ZN(U6366_n1) );
  AND2X1 U6366_U1 ( .IN1(n3272), .IN2(U6366_n1), .Q(n2980) );
  INVX0 U6367_U2 ( .INP(n5332), .ZN(U6367_n1) );
  AND2X1 U6367_U1 ( .IN1(n2980), .IN2(U6367_n1), .Q(n2704) );
  INVX0 U6368_U2 ( .INP(n5333), .ZN(U6368_n1) );
  AND2X1 U6368_U1 ( .IN1(n2704), .IN2(U6368_n1), .Q(n2647) );
  INVX0 U6369_U2 ( .INP(n5334), .ZN(U6369_n1) );
  AND2X1 U6369_U1 ( .IN1(n2647), .IN2(U6369_n1), .Q(n2554) );
  INVX0 U6370_U2 ( .INP(n5330), .ZN(U6370_n1) );
  AND2X1 U6370_U1 ( .IN1(n2554), .IN2(U6370_n1), .Q(n2507) );
  INVX0 U6371_U2 ( .INP(n5551), .ZN(U6371_n1) );
  AND2X1 U6371_U1 ( .IN1(n2507), .IN2(U6371_n1), .Q(n2485) );
  INVX0 U6372_U2 ( .INP(n5293), .ZN(U6372_n1) );
  AND2X1 U6372_U1 ( .IN1(n2485), .IN2(U6372_n1), .Q(n2425) );
  INVX0 U6373_U2 ( .INP(n5292), .ZN(U6373_n1) );
  AND2X1 U6373_U1 ( .IN1(n2425), .IN2(U6373_n1), .Q(n2419) );
  INVX0 U6374_U2 ( .INP(n5470), .ZN(U6374_n1) );
  AND2X1 U6374_U1 ( .IN1(n3743), .IN2(U6374_n1), .Q(n3682) );
  INVX0 U6375_U2 ( .INP(n5291), .ZN(U6375_n1) );
  AND2X1 U6375_U1 ( .IN1(n2419), .IN2(U6375_n1), .Q(n2405) );
  AND2X1 U6417_U2 ( .IN1(n4198), .IN2(U6417_n1), .Q(n2404) );
  INVX0 U6417_U1 ( .INP(n8808), .ZN(U6417_n1) );
  INVX0 U6446_U2 ( .INP(n1697), .ZN(U6446_n1) );
  AND2X1 U6446_U1 ( .IN1(g110), .IN2(U6446_n1), .Q(n3524) );
  INVX0 U6465_U2 ( .INP(n5600), .ZN(U6465_n1) );
  AND2X1 U6465_U1 ( .IN1(n3653), .IN2(U6465_n1), .Q(n4388) );
  INVX0 U6497_U2 ( .INP(n3635), .ZN(U6497_n1) );
  AND2X1 U6497_U1 ( .IN1(n756), .IN2(U6497_n1), .Q(n3005) );
  AND2X1 U6523_U2 ( .IN1(n967), .IN2(U6523_n1), .Q(n4945) );
  INVX0 U6523_U1 ( .INP(n8807), .ZN(U6523_n1) );
  INVX0 U6542_U2 ( .INP(n5300), .ZN(U6542_n1) );
  AND2X1 U6542_U1 ( .IN1(n756), .IN2(U6542_n1), .Q(n3525) );
  INVX0 U6552_U2 ( .INP(n5676), .ZN(U6552_n1) );
  AND2X1 U6552_U1 ( .IN1(n3281), .IN2(U6552_n1), .Q(n3277) );
  INVX0 U6553_U2 ( .INP(n5680), .ZN(U6553_n1) );
  AND2X1 U6553_U1 ( .IN1(n3276), .IN2(U6553_n1), .Q(n2989) );
  INVX0 U6554_U2 ( .INP(n5677), .ZN(U6554_n1) );
  AND2X1 U6554_U1 ( .IN1(n3277), .IN2(U6554_n1), .Q(n2991) );
  INVX0 U6555_U2 ( .INP(n5561), .ZN(U6555_n1) );
  AND2X1 U6555_U1 ( .IN1(n3687), .IN2(U6555_n1), .Q(n3281) );
  INVX0 U6556_U2 ( .INP(n5679), .ZN(U6556_n1) );
  AND2X1 U6556_U1 ( .IN1(n3279), .IN2(U6556_n1), .Q(n3276) );
  INVX0 U6559_U2 ( .INP(n5678), .ZN(U6559_n1) );
  AND2X1 U6559_U1 ( .IN1(n2991), .IN2(U6559_n1), .Q(n2710) );
  INVX0 U6560_U2 ( .INP(n5675), .ZN(U6560_n1) );
  AND2X1 U6560_U1 ( .IN1(n2989), .IN2(U6560_n1), .Q(n2707) );
  INVX0 U6561_U2 ( .INP(n5327), .ZN(U6561_n1) );
  AND2X1 U6561_U1 ( .IN1(n3174), .IN2(U6561_n1), .Q(n3116) );
  INVX0 U6570_U2 ( .INP(n5477), .ZN(U6570_n1) );
  AND2X1 U6570_U1 ( .IN1(n3362), .IN2(U6570_n1), .Q(n2527) );
  INVX0 U6911_U2 ( .INP(n915), .ZN(U6911_n1) );
  AND2X1 U6911_U1 ( .IN1(n3115), .IN2(U6911_n1), .Q(n3111) );
  INVX0 U6912_U2 ( .INP(n928), .ZN(U6912_n1) );
  AND2X1 U6912_U1 ( .IN1(n3115), .IN2(U6912_n1), .Q(n3131) );
  INVX0 U6917_U2 ( .INP(n5350), .ZN(U6917_n1) );
  AND2X1 U6917_U1 ( .IN1(n3933), .IN2(U6917_n1), .Q(n3799) );
  INVX0 U6926_U2 ( .INP(n5674), .ZN(U6926_n1) );
  AND2X1 U6926_U1 ( .IN1(n3664), .IN2(U6926_n1), .Q(n3662) );
  INVX0 U6927_U2 ( .INP(n5673), .ZN(U6927_n1) );
  AND2X1 U6927_U1 ( .IN1(n3673), .IN2(U6927_n1), .Q(n3671) );
  INVX0 U6929_U2 ( .INP(n3506), .ZN(U6929_n1) );
  AND2X1 U6929_U1 ( .IN1(n3505), .IN2(U6929_n1), .Q(n2790) );
  INVX0 U6931_U2 ( .INP(n5554), .ZN(U6931_n1) );
  AND2X1 U6931_U1 ( .IN1(n4490), .IN2(U6931_n1), .Q(n4178) );
  INVX0 U6932_U2 ( .INP(n5555), .ZN(U6932_n1) );
  AND2X1 U6932_U1 ( .IN1(n4514), .IN2(U6932_n1), .Q(n4196) );
  INVX0 U6933_U2 ( .INP(n5558), .ZN(U6933_n1) );
  AND2X1 U6933_U1 ( .IN1(n4178), .IN2(U6933_n1), .Q(n3736) );
  INVX0 U6934_U2 ( .INP(n5559), .ZN(U6934_n1) );
  AND2X1 U6934_U1 ( .IN1(n4196), .IN2(U6934_n1), .Q(n3741) );
  INVX0 U6935_U2 ( .INP(n5553), .ZN(U6935_n1) );
  AND2X1 U6935_U1 ( .IN1(n3736), .IN2(U6935_n1), .Q(n3664) );
  INVX0 U6936_U2 ( .INP(n5560), .ZN(U6936_n1) );
  AND2X1 U6936_U1 ( .IN1(n3741), .IN2(U6936_n1), .Q(n3673) );
  INVX0 U6937_U2 ( .INP(n5303), .ZN(U6937_n1) );
  AND2X1 U6937_U1 ( .IN1(n2601), .IN2(U6937_n1), .Q(n2598) );
  INVX0 U6938_U2 ( .INP(n5556), .ZN(U6938_n1) );
  AND2X1 U6938_U1 ( .IN1(n4804), .IN2(U6938_n1), .Q(n4490) );
  INVX0 U6939_U2 ( .INP(n5557), .ZN(U6939_n1) );
  AND2X1 U6939_U1 ( .IN1(n4811), .IN2(U6939_n1), .Q(n4514) );
  INVX0 U6940_U2 ( .INP(n5422), .ZN(U6940_n1) );
  AND2X1 U6940_U1 ( .IN1(n4814), .IN2(U6940_n1), .Q(n4519) );
  INVX0 U6941_U2 ( .INP(n5323), .ZN(U6941_n1) );
  AND2X1 U6941_U1 ( .IN1(n2607), .IN2(U6941_n1), .Q(n2594) );
  INVX0 U6944_U2 ( .INP(n5348), .ZN(U6944_n1) );
  AND2X1 U6944_U1 ( .IN1(n3084), .IN2(U6944_n1), .Q(n3033) );
  INVX0 U6950_U2 ( .INP(n5365), .ZN(U6950_n1) );
  AND2X1 U6950_U1 ( .IN1(n2598), .IN2(U6950_n1), .Q(n2590) );
  INVX0 U6954_U2 ( .INP(n928), .ZN(U6954_n1) );
  AND2X1 U6954_U1 ( .IN1(n3122), .IN2(U6954_n1), .Q(n3125) );
  INVX0 U6955_U2 ( .INP(n915), .ZN(U6955_n1) );
  AND2X1 U6955_U1 ( .IN1(n645), .IN2(U6955_n1), .Q(n3105) );
  INVX0 U6956_U2 ( .INP(n927), .ZN(U6956_n1) );
  AND2X1 U6956_U1 ( .IN1(n342), .IN2(U6956_n1), .Q(n3145) );
  INVX0 U6957_U2 ( .INP(n917), .ZN(U6957_n1) );
  AND2X1 U6957_U1 ( .IN1(n657), .IN2(U6957_n1), .Q(n3164) );
  INVX0 U7174_U2 ( .INP(n5288), .ZN(U7174_n1) );
  AND2X1 U7174_U1 ( .IN1(n2423), .IN2(U7174_n1), .Q(n2422) );
  INVX0 U7248_U2 ( .INP(g1536), .ZN(U7248_n1) );
  AND2X1 U7248_U1 ( .IN1(n4172), .IN2(U7248_n1), .Q(n4173) );
  INVX0 U7249_U2 ( .INP(g1193), .ZN(U7249_n1) );
  AND2X1 U7249_U1 ( .IN1(n4190), .IN2(U7249_n1), .Q(n4191) );
  INVX0 U7402_U2 ( .INP(n507), .ZN(U7402_n1) );
  AND2X1 U7402_U1 ( .IN1(n4034), .IN2(U7402_n1), .Q(n4037) );
  INVX0 U7405_U2 ( .INP(n508), .ZN(U7405_n1) );
  AND2X1 U7405_U1 ( .IN1(n4034), .IN2(U7405_n1), .Q(n4039) );
  INVX0 U7413_U2 ( .INP(n777), .ZN(U7413_n1) );
  AND2X1 U7413_U1 ( .IN1(n3969), .IN2(U7413_n1), .Q(n3972) );
  INVX0 U7416_U2 ( .INP(n196), .ZN(U7416_n1) );
  AND2X1 U7416_U1 ( .IN1(n3926), .IN2(U7416_n1), .Q(n3929) );
  INVX0 U7427_U2 ( .INP(n672), .ZN(U7427_n1) );
  AND2X1 U7427_U1 ( .IN1(n3860), .IN2(U7427_n1), .Q(n3863) );
  INVX0 U7438_U2 ( .INP(n418), .ZN(U7438_n1) );
  AND2X1 U7438_U1 ( .IN1(n4002), .IN2(U7438_n1), .Q(n4003) );
  INVX0 U7449_U2 ( .INP(n509), .ZN(U7449_n1) );
  AND2X1 U7449_U1 ( .IN1(n4034), .IN2(U7449_n1), .Q(n4032) );
  INVX0 U7455_U2 ( .INP(n510), .ZN(U7455_n1) );
  AND2X1 U7455_U1 ( .IN1(n4034), .IN2(U7455_n1), .Q(n4035) );
  INVX0 U7464_U2 ( .INP(n1326), .ZN(U7464_n1) );
  AND2X1 U7464_U1 ( .IN1(n3792), .IN2(U7464_n1), .Q(n3797) );
  INVX0 U7467_U2 ( .INP(n1330), .ZN(U7467_n1) );
  AND2X1 U7467_U1 ( .IN1(n3792), .IN2(U7467_n1), .Q(n3790) );
  INVX0 U7482_U2 ( .INP(n1324), .ZN(U7482_n1) );
  AND2X1 U7482_U1 ( .IN1(n3792), .IN2(U7482_n1), .Q(n3795) );
  INVX0 U7492_U2 ( .INP(n877), .ZN(U7492_n1) );
  AND2X1 U7492_U1 ( .IN1(n3893), .IN2(U7492_n1), .Q(n3891) );
  INVX0 U7513_U2 ( .INP(n43), .ZN(U7513_n1) );
  AND2X1 U7513_U1 ( .IN1(n3826), .IN2(U7513_n1), .Q(n3827) );
  INVX0 U7516_U2 ( .INP(n875), .ZN(U7516_n1) );
  AND2X1 U7516_U1 ( .IN1(n3893), .IN2(U7516_n1), .Q(n3896) );
  INVX0 U7549_U2 ( .INP(n412), .ZN(U7549_n1) );
  AND2X1 U7549_U1 ( .IN1(n4002), .IN2(U7549_n1), .Q(n4007) );
  INVX0 U7561_U2 ( .INP(n189), .ZN(U7561_n1) );
  AND2X1 U7561_U1 ( .IN1(n3926), .IN2(U7561_n1), .Q(n3931) );
  INVX0 U7574_U2 ( .INP(n1331), .ZN(U7574_n1) );
  AND2X1 U7574_U1 ( .IN1(n3792), .IN2(U7574_n1), .Q(n3793) );
  INVX0 U7577_U2 ( .INP(n195), .ZN(U7577_n1) );
  AND2X1 U7577_U1 ( .IN1(n3926), .IN2(U7577_n1), .Q(n3924) );
  INVX0 U7585_U2 ( .INP(n45), .ZN(U7585_n1) );
  AND2X1 U7585_U1 ( .IN1(n3826), .IN2(U7585_n1), .Q(n3831) );
  INVX0 U7595_U2 ( .INP(n51), .ZN(U7595_n1) );
  AND2X1 U7595_U1 ( .IN1(n3826), .IN2(U7595_n1), .Q(n3829) );
  INVX0 U7614_U2 ( .INP(n187), .ZN(U7614_n1) );
  AND2X1 U7614_U1 ( .IN1(n3926), .IN2(U7614_n1), .Q(n3927) );
  INVX0 U7621_U2 ( .INP(n772), .ZN(U7621_n1) );
  AND2X1 U7621_U1 ( .IN1(n3969), .IN2(U7621_n1), .Q(n3974) );
  INVX0 U7629_U2 ( .INP(n876), .ZN(U7629_n1) );
  AND2X1 U7629_U1 ( .IN1(n3893), .IN2(U7629_n1), .Q(n3898) );
  INVX0 U7636_U2 ( .INP(n770), .ZN(U7636_n1) );
  AND2X1 U7636_U1 ( .IN1(n3969), .IN2(U7636_n1), .Q(n3970) );
  INVX0 U7639_U2 ( .INP(n417), .ZN(U7639_n1) );
  AND2X1 U7639_U1 ( .IN1(n4002), .IN2(U7639_n1), .Q(n4000) );
  INVX0 U7649_U2 ( .INP(n668), .ZN(U7649_n1) );
  AND2X1 U7649_U1 ( .IN1(n3860), .IN2(U7649_n1), .Q(n3865) );
  INVX0 U7652_U2 ( .INP(n666), .ZN(U7652_n1) );
  AND2X1 U7652_U1 ( .IN1(n3860), .IN2(U7652_n1), .Q(n3861) );
  INVX0 U7668_U2 ( .INP(n50), .ZN(U7668_n1) );
  AND2X1 U7668_U1 ( .IN1(n3826), .IN2(U7668_n1), .Q(n3824) );
  INVX0 U7673_U2 ( .INP(n878), .ZN(U7673_n1) );
  AND2X1 U7673_U1 ( .IN1(n3893), .IN2(U7673_n1), .Q(n3894) );
  INVX0 U7690_U2 ( .INP(n776), .ZN(U7690_n1) );
  AND2X1 U7690_U1 ( .IN1(n3969), .IN2(U7690_n1), .Q(n3967) );
  INVX0 U7707_U2 ( .INP(n671), .ZN(U7707_n1) );
  AND2X1 U7707_U1 ( .IN1(n3860), .IN2(U7707_n1), .Q(n3858) );
  INVX0 U7712_U2 ( .INP(n410), .ZN(U7712_n1) );
  AND2X1 U7712_U1 ( .IN1(n4002), .IN2(U7712_n1), .Q(n4005) );
  AND2X1 U7792_U2 ( .IN1(g952), .IN2(U7792_n1), .Q(n2505) );
  INVX0 U7792_U1 ( .INP(n8808), .ZN(U7792_n1) );
  AND2X1 U7794_U2 ( .IN1(g1296), .IN2(U7794_n1), .Q(n2499) );
  INVX0 U7794_U1 ( .INP(n8807), .ZN(U7794_n1) );
  INVX0 U7895_U2 ( .INP(g113), .ZN(U7895_n1) );
  AND2X1 U7895_U1 ( .IN1(n2668), .IN2(U7895_n1), .Q(n2760) );
  INVX0 U7897_U2 ( .INP(g31), .ZN(U7897_n1) );
  AND2X1 U7897_U1 ( .IN1(g6), .IN2(U7897_n1), .Q(n3395) );
  AND2X1 U7977_U2 ( .IN1(g661), .IN2(U7977_n1), .Q(n4956) );
  INVX0 U7977_U1 ( .INP(n8808), .ZN(U7977_n1) );
  INVX0 U8034_U2 ( .INP(n5612), .ZN(U8034_n1) );
  AND2X1 U8034_U1 ( .IN1(n1166), .IN2(U8034_n1), .Q(n5026) );
  INVX0 U8036_U2 ( .INP(n5340), .ZN(U8036_n1) );
  AND2X1 U8036_U1 ( .IN1(n3729), .IN2(U8036_n1), .Q(n3941) );
  INVX0 U8050_U2 ( .INP(g1367), .ZN(U8050_n1) );
  AND2X1 U8050_U1 ( .IN1(n180), .IN2(U8050_n1), .Q(n3733) );
  AND2X1 U8055_U2 ( .IN1(g1345), .IN2(U8055_n1), .Q(n4798) );
  INVX0 U8055_U1 ( .INP(n8807), .ZN(U8055_n1) );
  AND2X1 U8060_U2 ( .IN1(g1002), .IN2(U8060_n1), .Q(n4805) );
  INVX0 U8060_U1 ( .INP(n8808), .ZN(U8060_n1) );
  INVX0 U8070_U2 ( .INP(g1361), .ZN(U8070_n1) );
  AND2X1 U8070_U1 ( .IN1(n181), .IN2(U8070_n1), .Q(n4175) );
  INVX0 U8074_U2 ( .INP(g1018), .ZN(U8074_n1) );
  AND2X1 U8074_U1 ( .IN1(n525), .IN2(U8074_n1), .Q(n4193) );
  INVX0 U8088_U2 ( .INP(g1024), .ZN(U8088_n1) );
  AND2X1 U8088_U1 ( .IN1(n524), .IN2(U8088_n1), .Q(n3738) );
  INVX0 U8112_U2 ( .INP(n4523), .ZN(U8112_n1) );
  AND2X1 U8112_U1 ( .IN1(n4525), .IN2(U8112_n1), .Q(n4524) );
  INVX0 U8113_U2 ( .INP(n5751), .ZN(U8113_n1) );
  AND2X1 U8113_U1 ( .IN1(n4526), .IN2(U8113_n1), .Q(n4523) );
  INVX0 U8147_U2 ( .INP(n2573), .ZN(U8147_n1) );
  AND2X1 U8147_U1 ( .IN1(g4659), .IN2(U8147_n1), .Q(n2577) );
  INVX0 U8165_U2 ( .INP(n2563), .ZN(U8165_n1) );
  AND2X1 U8165_U1 ( .IN1(g4849), .IN2(U8165_n1), .Q(n2567) );
  INVX0 U8185_U2 ( .INP(g1046), .ZN(U8185_n1) );
  AND2X1 U8185_U1 ( .IN1(n797), .IN2(U8185_n1), .Q(n4938) );
  INVX0 U8192_U2 ( .INP(g1389), .ZN(U8192_n1) );
  AND2X1 U8192_U1 ( .IN1(n175), .IN2(U8192_n1), .Q(n4913) );
  INVX0 U8210_U2 ( .INP(n1166), .ZN(U8210_n1) );
  AND2X1 U8210_U1 ( .IN1(n4722), .IN2(U8210_n1), .Q(n4714) );
  INVX0 U8223_U2 ( .INP(n4516), .ZN(U8223_n1) );
  AND2X1 U8223_U1 ( .IN1(n4518), .IN2(U8223_n1), .Q(n4517) );
  INVX0 U8224_U2 ( .INP(n5728), .ZN(U8224_n1) );
  AND2X1 U8224_U1 ( .IN1(n4519), .IN2(U8224_n1), .Q(n4516) );
  AND2X1 U8281_U2 ( .IN1(n872), .IN2(U8281_n1), .Q(n5111) );
  INVX0 U8281_U1 ( .INP(n8807), .ZN(U8281_n1) );
  AND2X1 U8307_U2 ( .IN1(g29216), .IN2(U8307_n1), .Q(g26900) );
  INVX0 U8307_U1 ( .INP(n8808), .ZN(U8307_n1) );
  INVX0 U8974_U2 ( .INP(test_so25), .ZN(U8974_n1) );
  AND2X1 U8974_U1 ( .IN1(n3362), .IN2(U8974_n1), .Q(n2552) );
  INVX0 U8975_U2 ( .INP(g528), .ZN(U8975_n1) );
  AND2X1 U8975_U1 ( .IN1(n3174), .IN2(U8975_n1), .Q(n3195) );
  AND2X1 U9065_U2 ( .IN1(g4145), .IN2(U9065_n1), .Q(n4721) );
  INVX0 U9065_U1 ( .INP(n8807), .ZN(U9065_n1) );
  AND2X1 U9070_U2 ( .IN1(g2841), .IN2(U9070_n1), .Q(n3730) );
  INVX0 U9070_U1 ( .INP(n8808), .ZN(U9070_n1) );
  INVX0 U9075_U2 ( .INP(g9), .ZN(U9075_n1) );
  AND2X1 U9075_U1 ( .IN1(g19), .IN2(U9075_n1), .Q(n3362) );
  AND2X1 U9076_U2 ( .IN1(g113), .IN2(U9076_n1), .Q(g25694) );
  INVX0 U9076_U1 ( .INP(n8807), .ZN(U9076_n1) );
  AND2X1 U9080_U2 ( .IN1(n4305), .IN2(U9080_n1), .Q(g29277) );
  INVX0 U9080_U1 ( .INP(n8807), .ZN(U9080_n1) );
  AND2X1 U9084_U2 ( .IN1(g4423), .IN2(U9084_n1), .Q(g26953) );
  INVX0 U9084_U1 ( .INP(n8807), .ZN(U9084_n1) );
  AND2X1 U9085_U2 ( .IN1(g64), .IN2(U9085_n1), .Q(g24212) );
  INVX0 U9085_U1 ( .INP(n8807), .ZN(U9085_n1) );
  AND2X1 U9086_U2 ( .IN1(n4283), .IN2(U9086_n1), .Q(g29279) );
  INVX0 U9086_U1 ( .INP(n8807), .ZN(U9086_n1) );
  AND2X1 U9090_U2 ( .IN1(g125), .IN2(U9090_n1), .Q(g25688) );
  INVX0 U9090_U1 ( .INP(n8807), .ZN(U9090_n1) );
  INVX0 U9098_U2 ( .INP(n301), .ZN(U9098_n1) );
  AND2X1 U9098_U1 ( .IN1(g4681), .IN2(U9098_n1), .Q(g34028) );
  INVX0 U9099_U2 ( .INP(n2608), .ZN(U9099_n1) );
  AND2X1 U9099_U1 ( .IN1(n2595), .IN2(U9099_n1), .Q(g34449) );
  AND2X1 U9101_U2 ( .IN1(g6745), .IN2(U9101_n1), .Q(g26880) );
  INVX0 U9101_U1 ( .INP(n8807), .ZN(U9101_n1) );
  INVX0 U9107_U2 ( .INP(n8483), .ZN(U9107_n1) );
  AND2X1 U9107_U1 ( .IN1(n4448), .IN2(U9107_n1), .Q(n4447) );
  INVX0 U9111_U2 ( .INP(n8480), .ZN(U9111_n1) );
  AND2X1 U9111_U1 ( .IN1(n4403), .IN2(U9111_n1), .Q(n4402) );
  INVX0 U9116_U2 ( .INP(n8489), .ZN(U9116_n1) );
  AND2X1 U9116_U1 ( .IN1(n4426), .IN2(U9116_n1), .Q(n4425) );
  INVX0 U9120_U2 ( .INP(n8477), .ZN(U9120_n1) );
  AND2X1 U9120_U1 ( .IN1(n4437), .IN2(U9120_n1), .Q(n4436) );
  INVX0 U9124_U2 ( .INP(n8485), .ZN(U9124_n1) );
  AND2X1 U9124_U1 ( .IN1(n4392), .IN2(U9124_n1), .Q(n4391) );
  INVX0 U9128_U2 ( .INP(n8478), .ZN(U9128_n1) );
  AND2X1 U9128_U1 ( .IN1(n4380), .IN2(U9128_n1), .Q(n4379) );
  INVX0 U9132_U2 ( .INP(n8487), .ZN(U9132_n1) );
  AND2X1 U9132_U1 ( .IN1(n4415), .IN2(U9132_n1), .Q(n4414) );
  INVX0 U9136_U2 ( .INP(n8488), .ZN(U9136_n1) );
  AND2X1 U9136_U1 ( .IN1(n4459), .IN2(U9136_n1), .Q(n4458) );
  INVX0 U9315_U2 ( .INP(n5753), .ZN(U9315_n1) );
  AND2X1 U9315_U1 ( .IN1(n5016), .IN2(U9315_n1), .Q(n5014) );
  INVX0 U9453_U2 ( .INP(n8481), .ZN(U9453_n1) );
  AND2X1 U9453_U1 ( .IN1(n3065), .IN2(U9453_n1), .Q(n3064) );
  INVX0 U9825_U2 ( .INP(n1697), .ZN(U9825_n1) );
  AND2X1 U9825_U1 ( .IN1(g112), .IN2(U9825_n1), .Q(n3115) );
  INVX0 U9886_U2 ( .INP(n5121), .ZN(U9886_n1) );
  AND2X1 U9886_U1 ( .IN1(g370), .IN2(U9886_n1), .Q(n4948) );
  INVX0 U9927_U2 ( .INP(g4098), .ZN(U9927_n1) );
  AND2X1 U9927_U1 ( .IN1(n3933), .IN2(U9927_n1), .Q(n3833) );
  INVX0 U9953_U2 ( .INP(n128), .ZN(U9953_n1) );
  AND2X1 U9953_U1 ( .IN1(g671), .IN2(U9953_n1), .Q(n4526) );
  INVX0 U9957_U2 ( .INP(n5283), .ZN(U9957_n1) );
  AND2X1 U9957_U1 ( .IN1(g4843), .IN2(U9957_n1), .Q(n2563) );
  INVX0 U9958_U2 ( .INP(n5656), .ZN(U9958_n1) );
  AND2X1 U9958_U1 ( .IN1(test_so19), .IN2(U9958_n1), .Q(n2573) );
  INVX0 U9968_U2 ( .INP(g4358), .ZN(U9968_n1) );
  AND2X1 U9968_U1 ( .IN1(n3084), .IN2(U9968_n1), .Q(n3023) );
  INVX0 U9972_U2 ( .INP(n4535), .ZN(U9972_n1) );
  AND2X1 U9972_U1 ( .IN1(g681), .IN2(U9972_n1), .Q(n5112) );
  INVX0 U9992_U2 ( .INP(n3676), .ZN(U9992_n1) );
  AND2X1 U9992_U1 ( .IN1(n3675), .IN2(U9992_n1), .Q(n2644) );
  INVX0 U10314_U2 ( .INP(g686), .ZN(U10314_n1) );
  AND2X1 U10314_U1 ( .IN1(g667), .IN2(U10314_n1), .Q(n4962) );
  INVX0 U10318_U2 ( .INP(n5681), .ZN(U10318_n1) );
  AND2X1 U10318_U1 ( .IN1(g5092), .IN2(U10318_n1), .Q(n5016) );
endmodule

