module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n462_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n449_, new_n364_, new_n580_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n530_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n139_, new_n314_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n227_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n570_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n182_, new_n407_, new_n480_, new_n513_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n522_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n131_, new_n255_, new_n533_, new_n459_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n440_, new_n531_, new_n252_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n134_, new_n433_, new_n435_, new_n265_, new_n370_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n412_, new_n327_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n545_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n284_, new_n119_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

nand g000 ( new_n119_, N29, N42, N75 );
not g001 ( N388, new_n119_ );
nand g002 ( new_n121_, N29, N36, N80 );
not g003 ( N389, new_n121_ );
nand g004 ( new_n123_, N29, N36, N42 );
not g005 ( N390, new_n123_ );
nand g006 ( new_n125_, N85, N86 );
not g007 ( N391, new_n125_ );
nand g008 ( new_n127_, N1, N8 );
not g009 ( new_n128_, new_n127_ );
nand g010 ( new_n129_, new_n128_, N13, N17 );
not g011 ( N418, new_n129_ );
not g012 ( new_n131_, N13 );
not g013 ( new_n132_, N17 );
nand g014 ( new_n133_, N1, N26 );
nor g015 ( new_n134_, new_n133_, new_n131_, new_n132_ );
nand g016 ( N419, new_n134_, new_n123_ );
nand g017 ( N420, N59, N75, N80 );
nand g018 ( N421, N36, N59, N80 );
nand g019 ( N422, N36, N42, N59 );
not g020 ( new_n139_, N90 );
nor g021 ( new_n140_, N87, N88 );
nor g022 ( N423, new_n140_, new_n139_ );
nand g023 ( N446, new_n134_, N390 );
nand g024 ( new_n143_, keyIn_0_0, N1, N26, N51 );
not g025 ( new_n144_, keyIn_0_0 );
nand g026 ( new_n145_, N1, N26, N51 );
nand g027 ( new_n146_, new_n145_, new_n144_ );
nand g028 ( new_n147_, new_n146_, new_n143_ );
not g029 ( N447, new_n147_ );
nand g030 ( new_n149_, new_n128_, N13, N55 );
nand g031 ( new_n150_, N29, N68 );
nor g032 ( N448, new_n149_, new_n150_ );
not g033 ( new_n152_, N74 );
nand g034 ( new_n153_, N59, N68 );
nor g035 ( N449, new_n149_, new_n152_, new_n153_ );
not g036 ( new_n155_, N89 );
nor g037 ( N450, new_n140_, new_n155_ );
nand g038 ( new_n157_, N111, N116 );
not g039 ( new_n158_, N111 );
not g040 ( new_n159_, N116 );
nand g041 ( new_n160_, new_n158_, new_n159_ );
nand g042 ( new_n161_, new_n160_, new_n157_ );
nand g043 ( new_n162_, N121, N126 );
not g044 ( new_n163_, N121 );
not g045 ( new_n164_, N126 );
nand g046 ( new_n165_, new_n163_, new_n164_ );
nand g047 ( new_n166_, new_n165_, new_n162_ );
nand g048 ( new_n167_, new_n161_, new_n166_ );
nand g049 ( new_n168_, new_n160_, new_n165_, new_n157_, new_n162_ );
nand g050 ( new_n169_, new_n167_, new_n168_ );
nand g051 ( new_n170_, new_n169_, N135 );
not g052 ( new_n171_, N135 );
nand g053 ( new_n172_, new_n167_, new_n171_, new_n168_ );
nand g054 ( new_n173_, new_n170_, new_n172_ );
not g055 ( new_n174_, N130 );
nand g056 ( new_n175_, N91, N96 );
not g057 ( new_n176_, N91 );
not g058 ( new_n177_, N96 );
nand g059 ( new_n178_, new_n176_, new_n177_ );
nand g060 ( new_n179_, new_n178_, new_n175_ );
nand g061 ( new_n180_, N101, N106 );
not g062 ( new_n181_, N101 );
not g063 ( new_n182_, N106 );
nand g064 ( new_n183_, new_n181_, new_n182_ );
nand g065 ( new_n184_, new_n183_, new_n180_ );
nand g066 ( new_n185_, new_n179_, new_n184_ );
nand g067 ( new_n186_, new_n178_, new_n183_, new_n175_, new_n180_ );
nand g068 ( new_n187_, new_n185_, new_n186_ );
nand g069 ( new_n188_, new_n187_, new_n174_ );
nand g070 ( new_n189_, new_n185_, N130, new_n186_ );
nand g071 ( new_n190_, new_n188_, new_n189_ );
nand g072 ( new_n191_, new_n173_, new_n190_ );
nand g073 ( new_n192_, new_n170_, new_n188_, new_n172_, new_n189_ );
nand g074 ( N767, new_n191_, new_n192_ );
nand g075 ( new_n194_, N183, N189 );
not g076 ( new_n195_, N183 );
not g077 ( new_n196_, N189 );
nand g078 ( new_n197_, new_n195_, new_n196_ );
nand g079 ( new_n198_, new_n197_, new_n194_ );
nand g080 ( new_n199_, N195, N201 );
not g081 ( new_n200_, N195 );
not g082 ( new_n201_, N201 );
nand g083 ( new_n202_, new_n200_, new_n201_ );
nand g084 ( new_n203_, new_n202_, new_n199_ );
nand g085 ( new_n204_, new_n198_, new_n203_ );
nand g086 ( new_n205_, new_n197_, new_n202_, new_n194_, new_n199_ );
nand g087 ( new_n206_, new_n204_, new_n205_ );
nand g088 ( new_n207_, new_n206_, N207 );
not g089 ( new_n208_, N207 );
nand g090 ( new_n209_, new_n204_, new_n208_, new_n205_ );
nand g091 ( new_n210_, new_n207_, new_n209_ );
nand g092 ( new_n211_, N159, N165 );
not g093 ( new_n212_, N159 );
not g094 ( new_n213_, N165 );
nand g095 ( new_n214_, new_n212_, new_n213_ );
nand g096 ( new_n215_, new_n214_, new_n211_ );
nand g097 ( new_n216_, N171, N177 );
not g098 ( new_n217_, N171 );
not g099 ( new_n218_, N177 );
nand g100 ( new_n219_, new_n217_, new_n218_ );
nand g101 ( new_n220_, new_n219_, new_n216_ );
nand g102 ( new_n221_, new_n215_, new_n220_ );
nand g103 ( new_n222_, new_n214_, new_n219_, new_n211_, new_n216_ );
nand g104 ( new_n223_, new_n221_, new_n222_ );
nand g105 ( new_n224_, new_n223_, new_n174_ );
nand g106 ( new_n225_, new_n221_, N130, new_n222_ );
nand g107 ( new_n226_, new_n224_, new_n225_ );
nand g108 ( new_n227_, new_n210_, new_n226_ );
nand g109 ( new_n228_, new_n207_, new_n224_, new_n209_, new_n225_ );
nand g110 ( N768, new_n227_, new_n228_ );
not g111 ( new_n230_, keyIn_0_27 );
not g112 ( new_n231_, keyIn_0_23 );
not g113 ( new_n232_, keyIn_0_21 );
not g114 ( new_n233_, keyIn_0_15 );
not g115 ( new_n234_, keyIn_0_10 );
nand g116 ( new_n235_, new_n147_, keyIn_0_6 );
not g117 ( new_n236_, keyIn_0_6 );
nand g118 ( new_n237_, new_n146_, new_n236_, new_n143_ );
nand g119 ( new_n238_, new_n235_, new_n237_ );
nand g120 ( new_n239_, new_n238_, new_n234_ );
nand g121 ( new_n240_, new_n235_, keyIn_0_10, new_n237_ );
nand g122 ( new_n241_, new_n239_, new_n240_ );
not g123 ( new_n242_, N42 );
nand g124 ( new_n243_, new_n132_, new_n242_ );
nand g125 ( new_n244_, new_n243_, keyIn_0_4 );
not g126 ( new_n245_, keyIn_0_4 );
nand g127 ( new_n246_, new_n245_, new_n132_, new_n242_ );
nand g128 ( new_n247_, new_n244_, new_n246_ );
not g129 ( new_n248_, keyIn_0_5 );
nand g130 ( new_n249_, new_n248_, N17, N42 );
nand g131 ( new_n250_, N17, N42 );
nand g132 ( new_n251_, new_n250_, keyIn_0_5 );
nand g133 ( new_n252_, new_n251_, new_n249_ );
nand g134 ( new_n253_, new_n247_, keyIn_0_9, new_n252_ );
nand g135 ( new_n254_, N59, N156 );
not g136 ( new_n255_, new_n254_ );
not g137 ( new_n256_, keyIn_0_9 );
nand g138 ( new_n257_, new_n247_, new_n252_ );
nand g139 ( new_n258_, new_n257_, new_n256_ );
nand g140 ( new_n259_, new_n258_, new_n253_, new_n255_ );
not g141 ( new_n260_, new_n259_ );
nand g142 ( new_n261_, new_n260_, new_n233_, new_n241_ );
nand g143 ( new_n262_, new_n260_, new_n241_ );
nand g144 ( new_n263_, new_n262_, keyIn_0_15 );
nand g145 ( new_n264_, new_n263_, new_n261_ );
not g146 ( new_n265_, keyIn_0_2 );
nand g147 ( new_n266_, new_n265_, N42, N59, N75 );
nand g148 ( new_n267_, N42, N59, N75 );
nand g149 ( new_n268_, new_n267_, keyIn_0_2 );
nand g150 ( new_n269_, new_n268_, new_n266_ );
nand g151 ( new_n270_, new_n269_, keyIn_0_8 );
not g152 ( new_n271_, keyIn_0_8 );
nand g153 ( new_n272_, new_n268_, new_n271_, new_n266_ );
nand g154 ( new_n273_, new_n270_, new_n272_ );
nand g155 ( new_n274_, new_n128_, keyIn_0_1, N17, N51 );
not g156 ( new_n275_, keyIn_0_1 );
nand g157 ( new_n276_, new_n128_, N17, N51 );
nand g158 ( new_n277_, new_n276_, new_n275_ );
nand g159 ( new_n278_, new_n277_, new_n274_ );
nand g160 ( new_n279_, new_n278_, keyIn_0_7 );
not g161 ( new_n280_, keyIn_0_7 );
nand g162 ( new_n281_, new_n277_, new_n280_, new_n274_ );
nand g163 ( new_n282_, new_n279_, new_n281_ );
nand g164 ( new_n283_, new_n282_, keyIn_0_11, new_n273_ );
not g165 ( new_n284_, keyIn_0_11 );
nand g166 ( new_n285_, new_n282_, new_n273_ );
nand g167 ( new_n286_, new_n285_, new_n284_ );
nand g168 ( new_n287_, new_n286_, new_n283_ );
nand g169 ( new_n288_, new_n264_, keyIn_0_17, new_n287_ );
not g170 ( new_n289_, keyIn_0_17 );
nand g171 ( new_n290_, new_n264_, new_n287_ );
nand g172 ( new_n291_, new_n290_, new_n289_ );
nand g173 ( new_n292_, new_n291_, new_n288_ );
nand g174 ( new_n293_, new_n292_, N126 );
nand g175 ( new_n294_, new_n255_, keyIn_0_3 );
not g176 ( new_n295_, keyIn_0_3 );
nand g177 ( new_n296_, new_n254_, new_n295_ );
nand g178 ( new_n297_, new_n241_, new_n294_, new_n296_ );
not g179 ( new_n298_, new_n297_ );
nand g180 ( new_n299_, new_n298_, N17 );
nand g181 ( new_n300_, new_n299_, keyIn_0_16 );
not g182 ( new_n301_, keyIn_0_16 );
nand g183 ( new_n302_, new_n298_, new_n301_, N17 );
nand g184 ( new_n303_, new_n300_, N1, new_n302_ );
nand g185 ( new_n304_, new_n303_, N153 );
nand g186 ( new_n305_, new_n293_, new_n232_, new_n304_ );
nand g187 ( new_n306_, new_n293_, new_n304_ );
nand g188 ( new_n307_, new_n306_, keyIn_0_21 );
not g189 ( new_n308_, N268 );
not g190 ( new_n309_, keyIn_0_14 );
nand g191 ( new_n310_, N29, N75, N80 );
not g192 ( new_n311_, new_n310_ );
nand g193 ( new_n312_, new_n241_, new_n309_, N55, new_n311_ );
nand g194 ( new_n313_, new_n241_, N55, new_n311_ );
nand g195 ( new_n314_, new_n313_, keyIn_0_14 );
nand g196 ( new_n315_, new_n314_, new_n308_, new_n312_ );
not g197 ( new_n316_, new_n315_ );
nand g198 ( new_n317_, new_n316_, keyIn_0_19 );
not g199 ( new_n318_, keyIn_0_19 );
nand g200 ( new_n319_, new_n315_, new_n318_ );
nand g201 ( new_n320_, new_n317_, new_n319_ );
not g202 ( new_n321_, new_n320_ );
nand g203 ( new_n322_, new_n307_, new_n305_, new_n321_ );
nand g204 ( new_n323_, new_n322_, new_n231_ );
nand g205 ( new_n324_, new_n307_, keyIn_0_23, new_n305_, new_n321_ );
nand g206 ( new_n325_, new_n323_, new_n324_ );
nand g207 ( new_n326_, new_n325_, N201 );
nand g208 ( new_n327_, new_n323_, new_n201_, new_n324_ );
nand g209 ( new_n328_, new_n326_, new_n327_ );
not g210 ( new_n329_, new_n328_ );
nand g211 ( new_n330_, new_n329_, N261 );
not g212 ( new_n331_, N261 );
nand g213 ( new_n332_, new_n328_, new_n331_ );
nand g214 ( new_n333_, new_n330_, N219, new_n332_ );
nand g215 ( new_n334_, new_n329_, N228 );
not g216 ( new_n335_, new_n334_ );
not g217 ( new_n336_, new_n326_ );
nand g218 ( new_n337_, new_n336_, N237 );
not g219 ( new_n338_, new_n337_ );
nand g220 ( new_n339_, new_n325_, N246 );
nand g221 ( new_n340_, N42, N72, N73 );
nor g222 ( new_n341_, new_n149_, new_n340_, new_n153_ );
nand g223 ( new_n342_, new_n341_, N201 );
nand g224 ( new_n343_, N255, N267 );
nand g225 ( new_n344_, N121, N210 );
nand g226 ( new_n345_, new_n339_, new_n342_, new_n343_, new_n344_ );
nor g227 ( new_n346_, new_n335_, new_n338_, new_n345_ );
nand g228 ( new_n347_, new_n346_, new_n333_ );
nand g229 ( new_n348_, new_n347_, new_n230_ );
nand g230 ( new_n349_, new_n346_, keyIn_0_27, new_n333_ );
nand g231 ( N850, new_n348_, new_n349_ );
nand g232 ( new_n351_, new_n292_, N116 );
nand g233 ( new_n352_, new_n303_, N146 );
nand g234 ( new_n353_, new_n352_, new_n315_ );
not g235 ( new_n354_, new_n353_ );
nand g236 ( new_n355_, new_n354_, new_n196_, new_n351_ );
not g237 ( new_n356_, keyIn_0_22 );
not g238 ( new_n357_, keyIn_0_20 );
nand g239 ( new_n358_, new_n292_, N121 );
nand g240 ( new_n359_, new_n303_, N149 );
nand g241 ( new_n360_, new_n358_, new_n357_, new_n359_ );
nand g242 ( new_n361_, new_n358_, new_n359_ );
nand g243 ( new_n362_, new_n361_, keyIn_0_20 );
not g244 ( new_n363_, keyIn_0_18 );
nand g245 ( new_n364_, new_n316_, new_n363_ );
nand g246 ( new_n365_, new_n315_, keyIn_0_18 );
nand g247 ( new_n366_, new_n364_, new_n365_ );
not g248 ( new_n367_, new_n366_ );
nand g249 ( new_n368_, new_n362_, new_n360_, new_n367_ );
nand g250 ( new_n369_, new_n368_, new_n356_ );
nand g251 ( new_n370_, new_n362_, keyIn_0_22, new_n360_, new_n367_ );
nand g252 ( new_n371_, new_n369_, new_n370_ );
nand g253 ( new_n372_, new_n371_, new_n200_ );
nand g254 ( new_n373_, new_n372_, N261, new_n327_, new_n355_ );
nand g255 ( new_n374_, new_n373_, keyIn_0_24 );
nand g256 ( new_n375_, new_n354_, new_n351_ );
nand g257 ( new_n376_, new_n375_, N189 );
nand g258 ( new_n377_, new_n369_, N195, new_n370_ );
not g259 ( new_n378_, new_n377_ );
nand g260 ( new_n379_, new_n378_, new_n355_ );
nand g261 ( new_n380_, new_n374_, new_n376_, new_n379_ );
not g262 ( new_n381_, new_n380_ );
not g263 ( new_n382_, keyIn_0_24 );
nand g264 ( new_n383_, new_n327_, N261 );
not g265 ( new_n384_, new_n383_ );
nand g266 ( new_n385_, new_n384_, new_n382_, new_n355_, new_n372_ );
not g267 ( new_n386_, keyIn_0_25 );
nand g268 ( new_n387_, new_n372_, N201, new_n325_, new_n355_ );
nand g269 ( new_n388_, new_n387_, new_n386_ );
nand g270 ( new_n389_, new_n336_, keyIn_0_25, new_n355_, new_n372_ );
nand g271 ( new_n390_, new_n385_, new_n388_, new_n389_ );
not g272 ( new_n391_, new_n390_ );
nand g273 ( new_n392_, new_n391_, new_n381_, keyIn_0_26 );
not g274 ( new_n393_, keyIn_0_26 );
nand g275 ( new_n394_, new_n391_, new_n381_ );
nand g276 ( new_n395_, new_n394_, new_n393_ );
nand g277 ( new_n396_, new_n395_, new_n392_ );
nand g278 ( new_n397_, new_n292_, N111 );
nand g279 ( new_n398_, new_n303_, N143 );
nand g280 ( new_n399_, new_n398_, new_n315_ );
not g281 ( new_n400_, new_n399_ );
nand g282 ( new_n401_, new_n400_, new_n397_ );
nand g283 ( new_n402_, new_n401_, N183 );
nand g284 ( new_n403_, new_n400_, new_n195_, new_n397_ );
nand g285 ( new_n404_, new_n402_, new_n403_ );
not g286 ( new_n405_, new_n404_ );
nand g287 ( new_n406_, new_n396_, new_n405_ );
nand g288 ( new_n407_, new_n395_, new_n392_, new_n404_ );
nand g289 ( new_n408_, new_n406_, N219, new_n407_ );
nand g290 ( new_n409_, new_n405_, N228 );
nand g291 ( new_n410_, new_n401_, N183, N237 );
nand g292 ( new_n411_, new_n401_, N246 );
nand g293 ( new_n412_, N106, N210 );
nand g294 ( new_n413_, new_n341_, N183 );
nand g295 ( new_n414_, new_n410_, new_n411_, new_n412_, new_n413_ );
not g296 ( new_n415_, new_n414_ );
nand g297 ( N863, new_n408_, new_n409_, new_n415_ );
nand g298 ( new_n417_, new_n383_, new_n326_ );
nand g299 ( new_n418_, new_n417_, new_n372_ );
nand g300 ( new_n419_, new_n418_, new_n377_ );
nand g301 ( new_n420_, new_n376_, new_n355_ );
not g302 ( new_n421_, new_n420_ );
nand g303 ( new_n422_, new_n419_, new_n421_ );
nand g304 ( new_n423_, new_n418_, new_n377_, new_n420_ );
nand g305 ( new_n424_, new_n422_, N219, new_n423_ );
nand g306 ( new_n425_, new_n421_, N228 );
not g307 ( new_n426_, new_n425_ );
nand g308 ( new_n427_, new_n375_, N189, N237 );
not g309 ( new_n428_, new_n427_ );
nand g310 ( new_n429_, new_n375_, N246 );
nand g311 ( new_n430_, new_n341_, N189 );
nand g312 ( new_n431_, N255, N259 );
nand g313 ( new_n432_, N111, N210 );
nand g314 ( new_n433_, new_n429_, new_n430_, new_n431_, new_n432_ );
nor g315 ( new_n434_, new_n426_, new_n428_, new_n433_ );
nand g316 ( new_n435_, new_n424_, new_n434_ );
nand g317 ( new_n436_, new_n435_, keyIn_0_30 );
not g318 ( new_n437_, keyIn_0_30 );
nand g319 ( new_n438_, new_n424_, new_n437_, new_n434_ );
nand g320 ( N864, new_n436_, new_n438_ );
not g321 ( new_n440_, keyIn_0_31 );
nand g322 ( new_n441_, new_n417_, new_n372_, new_n377_ );
nand g323 ( new_n442_, new_n372_, new_n377_ );
nand g324 ( new_n443_, new_n442_, new_n326_, new_n383_ );
nand g325 ( new_n444_, new_n441_, N219, new_n443_ );
nand g326 ( new_n445_, new_n372_, N228, new_n377_ );
not g327 ( new_n446_, new_n445_ );
nand g328 ( new_n447_, new_n378_, N237 );
not g329 ( new_n448_, new_n447_ );
nand g330 ( new_n449_, new_n369_, N246, new_n370_ );
nand g331 ( new_n450_, new_n341_, N195 );
nand g332 ( new_n451_, N255, N260 );
nand g333 ( new_n452_, N116, N210 );
nand g334 ( new_n453_, new_n449_, new_n450_, new_n451_, new_n452_ );
nor g335 ( new_n454_, new_n446_, new_n448_, new_n453_ );
nand g336 ( new_n455_, new_n454_, new_n444_ );
nand g337 ( new_n456_, new_n455_, new_n440_ );
nand g338 ( new_n457_, new_n454_, new_n444_, keyIn_0_31 );
nand g339 ( N865, new_n456_, new_n457_ );
nand g340 ( new_n459_, new_n396_, new_n403_ );
nand g341 ( new_n460_, new_n459_, new_n402_ );
nand g342 ( new_n461_, new_n292_, N96 );
not g343 ( new_n462_, keyIn_0_12 );
nand g344 ( new_n463_, new_n298_, new_n462_, N55 );
nand g345 ( new_n464_, new_n298_, N55 );
nand g346 ( new_n465_, new_n464_, keyIn_0_12 );
nand g347 ( new_n466_, new_n465_, new_n463_ );
nand g348 ( new_n467_, new_n466_, N146 );
not g349 ( new_n468_, new_n467_ );
nand g350 ( new_n469_, N51, N138 );
not g351 ( new_n470_, new_n469_ );
nand g352 ( new_n471_, new_n241_, keyIn_0_13, N17, new_n311_ );
not g353 ( new_n472_, keyIn_0_13 );
nand g354 ( new_n473_, new_n241_, N17, new_n311_ );
nand g355 ( new_n474_, new_n473_, new_n472_ );
nand g356 ( new_n475_, new_n474_, new_n308_, new_n471_ );
not g357 ( new_n476_, new_n475_ );
nor g358 ( new_n477_, new_n468_, new_n470_, new_n476_ );
nand g359 ( new_n478_, new_n477_, new_n213_, new_n461_ );
nand g360 ( new_n479_, new_n292_, N101 );
nand g361 ( new_n480_, new_n466_, N149 );
not g362 ( new_n481_, new_n480_ );
nand g363 ( new_n482_, N17, N138 );
not g364 ( new_n483_, new_n482_ );
nor g365 ( new_n484_, new_n481_, new_n476_, new_n483_ );
nand g366 ( new_n485_, new_n484_, new_n217_, new_n479_ );
nand g367 ( new_n486_, new_n478_, new_n485_ );
not g368 ( new_n487_, new_n486_ );
nand g369 ( new_n488_, new_n292_, N106 );
nand g370 ( new_n489_, new_n466_, N153 );
not g371 ( new_n490_, new_n489_ );
nand g372 ( new_n491_, N138, N152 );
not g373 ( new_n492_, new_n491_ );
nor g374 ( new_n493_, new_n490_, new_n476_, new_n492_ );
nand g375 ( new_n494_, new_n493_, new_n218_, new_n488_ );
nand g376 ( new_n495_, new_n487_, new_n494_ );
not g377 ( new_n496_, new_n495_ );
nand g378 ( new_n497_, new_n460_, new_n496_ );
nand g379 ( new_n498_, new_n497_, keyIn_0_28 );
not g380 ( new_n499_, keyIn_0_28 );
nand g381 ( new_n500_, new_n460_, new_n499_, new_n496_ );
nand g382 ( new_n501_, new_n477_, new_n461_ );
nand g383 ( new_n502_, new_n501_, N165 );
nand g384 ( new_n503_, new_n493_, new_n488_ );
nand g385 ( new_n504_, new_n503_, N177 );
nand g386 ( new_n505_, new_n484_, new_n479_ );
nand g387 ( new_n506_, new_n505_, N171 );
nand g388 ( new_n507_, new_n504_, new_n506_ );
nand g389 ( new_n508_, new_n487_, new_n507_ );
nand g390 ( new_n509_, new_n508_, new_n502_ );
not g391 ( new_n510_, new_n509_ );
nand g392 ( new_n511_, new_n498_, keyIn_0_29, new_n500_, new_n510_ );
not g393 ( new_n512_, keyIn_0_29 );
nand g394 ( new_n513_, new_n498_, new_n500_, new_n510_ );
nand g395 ( new_n514_, new_n513_, new_n512_ );
nand g396 ( new_n515_, new_n514_, new_n511_ );
nand g397 ( new_n516_, new_n292_, N91 );
nand g398 ( new_n517_, new_n466_, N143 );
not g399 ( new_n518_, new_n517_ );
nand g400 ( new_n519_, N8, N138 );
not g401 ( new_n520_, new_n519_ );
nor g402 ( new_n521_, new_n518_, new_n476_, new_n520_ );
nand g403 ( new_n522_, new_n521_, new_n212_, new_n516_ );
nand g404 ( new_n523_, new_n515_, new_n522_ );
nand g405 ( new_n524_, new_n521_, new_n516_ );
nand g406 ( new_n525_, new_n524_, N159 );
nand g407 ( N866, new_n523_, new_n525_ );
nand g408 ( new_n527_, new_n460_, new_n494_, new_n504_ );
nand g409 ( new_n528_, new_n504_, new_n494_ );
nand g410 ( new_n529_, new_n459_, new_n402_, new_n528_ );
nand g411 ( new_n530_, new_n527_, N219, new_n529_ );
nand g412 ( new_n531_, new_n504_, N228, new_n494_ );
nand g413 ( new_n532_, new_n503_, N177, N237 );
nand g414 ( new_n533_, new_n503_, N246 );
nand g415 ( new_n534_, N101, N210 );
nand g416 ( new_n535_, new_n341_, N177 );
nand g417 ( new_n536_, new_n532_, new_n533_, new_n534_, new_n535_ );
not g418 ( new_n537_, new_n536_ );
nand g419 ( N874, new_n530_, new_n531_, new_n537_ );
nand g420 ( new_n539_, new_n525_, new_n522_ );
not g421 ( new_n540_, new_n539_ );
nand g422 ( new_n541_, new_n515_, new_n540_ );
nand g423 ( new_n542_, new_n514_, new_n511_, new_n539_ );
nand g424 ( new_n543_, new_n541_, N219, new_n542_ );
nand g425 ( new_n544_, new_n540_, N228 );
not g426 ( new_n545_, new_n544_ );
nand g427 ( new_n546_, new_n524_, N159, N237 );
nand g428 ( new_n547_, new_n524_, N246 );
nand g429 ( new_n548_, new_n341_, N159 );
nand g430 ( new_n549_, N210, N268 );
nand g431 ( new_n550_, new_n546_, new_n547_, new_n548_, new_n549_ );
nor g432 ( new_n551_, new_n545_, new_n550_ );
nand g433 ( N878, new_n543_, new_n551_ );
nand g434 ( new_n553_, new_n460_, new_n494_ );
nand g435 ( new_n554_, new_n553_, new_n504_ );
nand g436 ( new_n555_, new_n554_, new_n485_ );
nand g437 ( new_n556_, new_n502_, new_n478_ );
nand g438 ( new_n557_, new_n555_, new_n506_, new_n556_ );
nand g439 ( new_n558_, new_n555_, new_n506_ );
not g440 ( new_n559_, new_n556_ );
nand g441 ( new_n560_, new_n558_, new_n559_ );
nand g442 ( new_n561_, new_n560_, N219, new_n557_ );
nand g443 ( new_n562_, new_n559_, N228 );
nand g444 ( new_n563_, new_n501_, N165, N237 );
nand g445 ( new_n564_, new_n501_, N246 );
nand g446 ( new_n565_, N91, N210 );
nand g447 ( new_n566_, new_n341_, N165 );
nand g448 ( new_n567_, new_n563_, new_n564_, new_n565_, new_n566_ );
not g449 ( new_n568_, new_n567_ );
nand g450 ( N879, new_n561_, new_n562_, new_n568_ );
nand g451 ( new_n570_, new_n554_, new_n485_, new_n506_ );
nand g452 ( new_n571_, new_n506_, new_n485_ );
nand g453 ( new_n572_, new_n553_, new_n504_, new_n571_ );
nand g454 ( new_n573_, new_n570_, N219, new_n572_ );
nand g455 ( new_n574_, new_n506_, N228, new_n485_ );
nand g456 ( new_n575_, new_n505_, N171, N237 );
nand g457 ( new_n576_, new_n505_, N246 );
nand g458 ( new_n577_, N96, N210 );
nand g459 ( new_n578_, new_n341_, N171 );
nand g460 ( new_n579_, new_n575_, new_n576_, new_n577_, new_n578_ );
not g461 ( new_n580_, new_n579_ );
nand g462 ( N880, new_n573_, new_n574_, new_n580_ );
endmodule