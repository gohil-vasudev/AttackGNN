module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n888_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n504_, new_n862_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n774_, new_n716_, new_n701_, new_n792_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n890_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n848_, new_n277_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n696_, new_n939_, new_n208_, new_n632_, new_n671_, new_n528_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n901_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n851_, new_n932_, new_n878_, new_n543_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n918_, new_n810_, new_n808_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n719_, new_n869_, new_n273_, new_n224_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n741_, new_n806_, new_n605_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n612_, new_n919_, new_n302_, new_n755_, new_n225_, new_n922_, new_n387_, new_n615_, new_n476_, new_n722_, new_n856_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n584_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n756_, new_n495_, new_n823_, new_n431_, new_n927_, new_n818_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n865_, new_n358_, new_n877_, new_n348_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n896_, new_n226_, new_n802_, new_n697_, new_n709_, new_n373_, new_n866_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n573_, new_n765_, new_n405_;

xnor g000 ( new_n202_, N81, N85 );
xnor g001 ( new_n203_, new_n202_, keyIn_0_10 );
xnor g002 ( new_n204_, N89, N93 );
xnor g003 ( new_n205_, new_n204_, keyIn_0_11 );
xnor g004 ( new_n206_, new_n203_, new_n205_ );
xnor g005 ( new_n207_, new_n206_, keyIn_0_33 );
xnor g006 ( new_n208_, N65, N69 );
xnor g007 ( new_n209_, new_n208_, keyIn_0_8 );
xor g008 ( new_n210_, N73, N77 );
xnor g009 ( new_n211_, new_n210_, keyIn_0_9 );
xnor g010 ( new_n212_, new_n211_, new_n209_ );
xnor g011 ( new_n213_, new_n212_, keyIn_0_32 );
xnor g012 ( new_n214_, new_n213_, new_n207_ );
xnor g013 ( new_n215_, new_n214_, keyIn_0_43 );
nand g014 ( new_n216_, N129, N137 );
xor g015 ( new_n217_, new_n215_, new_n216_ );
xnor g016 ( new_n218_, new_n217_, keyIn_0_47 );
xor g017 ( new_n219_, N1, N17 );
xnor g018 ( new_n220_, N33, N49 );
xnor g019 ( new_n221_, new_n219_, new_n220_ );
xnor g020 ( new_n222_, new_n218_, new_n221_ );
xor g021 ( new_n223_, new_n222_, keyIn_0_55 );
not g022 ( new_n224_, keyIn_0_35 );
xnor g023 ( new_n225_, N113, N117 );
xnor g024 ( new_n226_, new_n225_, keyIn_0_14 );
not g025 ( new_n227_, keyIn_0_15 );
xnor g026 ( new_n228_, N121, N125 );
xnor g027 ( new_n229_, new_n228_, new_n227_ );
xnor g028 ( new_n230_, new_n226_, new_n229_ );
xnor g029 ( new_n231_, new_n230_, new_n224_ );
xnor g030 ( new_n232_, new_n207_, new_n231_ );
xnor g031 ( new_n233_, new_n232_, keyIn_0_46 );
nand g032 ( new_n234_, N132, N137 );
xor g033 ( new_n235_, new_n233_, new_n234_ );
xnor g034 ( new_n236_, new_n235_, keyIn_0_50 );
xnor g035 ( new_n237_, N13, N29 );
xnor g036 ( new_n238_, new_n237_, keyIn_0_23 );
xor g037 ( new_n239_, N45, N61 );
xnor g038 ( new_n240_, new_n238_, new_n239_ );
xnor g039 ( new_n241_, new_n236_, new_n240_ );
xnor g040 ( new_n242_, new_n241_, keyIn_0_58 );
not g041 ( new_n243_, new_n242_ );
xnor g042 ( new_n244_, N97, N101 );
xnor g043 ( new_n245_, new_n244_, keyIn_0_12 );
xnor g044 ( new_n246_, N105, N109 );
xnor g045 ( new_n247_, new_n246_, keyIn_0_13 );
xnor g046 ( new_n248_, new_n245_, new_n247_ );
xnor g047 ( new_n249_, new_n248_, keyIn_0_34 );
xnor g048 ( new_n250_, new_n231_, new_n249_ );
xnor g049 ( new_n251_, new_n250_, keyIn_0_44 );
nand g050 ( new_n252_, N130, N137 );
xor g051 ( new_n253_, new_n251_, new_n252_ );
xnor g052 ( new_n254_, new_n253_, keyIn_0_48 );
xor g053 ( new_n255_, N5, N21 );
xnor g054 ( new_n256_, N37, N53 );
xnor g055 ( new_n257_, new_n255_, new_n256_ );
xnor g056 ( new_n258_, new_n254_, new_n257_ );
xnor g057 ( new_n259_, new_n258_, keyIn_0_56 );
nand g058 ( new_n260_, new_n243_, new_n259_ );
xnor g059 ( new_n261_, new_n213_, new_n249_ );
xnor g060 ( new_n262_, new_n261_, keyIn_0_45 );
nand g061 ( new_n263_, N131, N137 );
and g062 ( new_n264_, new_n263_, keyIn_0_16 );
not g063 ( new_n265_, N137 );
not g064 ( new_n266_, keyIn_0_16 );
nand g065 ( new_n267_, new_n266_, N131 );
nor g066 ( new_n268_, new_n267_, new_n265_ );
nor g067 ( new_n269_, new_n268_, new_n264_ );
xor g068 ( new_n270_, new_n262_, new_n269_ );
xnor g069 ( new_n271_, new_n270_, keyIn_0_49 );
xnor g070 ( new_n272_, N41, N57 );
xnor g071 ( new_n273_, new_n272_, keyIn_0_22 );
xor g072 ( new_n274_, N9, N25 );
xnor g073 ( new_n275_, new_n274_, keyIn_0_21 );
xnor g074 ( new_n276_, new_n275_, new_n273_ );
xnor g075 ( new_n277_, new_n276_, keyIn_0_36 );
xnor g076 ( new_n278_, new_n271_, new_n277_ );
xnor g077 ( new_n279_, new_n278_, keyIn_0_57 );
not g078 ( new_n280_, new_n279_ );
nand g079 ( new_n281_, new_n260_, new_n280_ );
nor g080 ( new_n282_, new_n260_, new_n280_ );
not g081 ( new_n283_, new_n259_ );
nand g082 ( new_n284_, new_n283_, new_n242_ );
nand g083 ( new_n285_, new_n284_, new_n223_ );
nor g084 ( new_n286_, new_n282_, new_n285_ );
nand g085 ( new_n287_, new_n286_, new_n281_ );
xnor g086 ( new_n288_, new_n279_, keyIn_0_63 );
nor g087 ( new_n289_, new_n260_, new_n223_ );
nand g088 ( new_n290_, new_n289_, new_n288_ );
nand g089 ( new_n291_, new_n287_, new_n290_ );
not g090 ( new_n292_, keyIn_0_61 );
not g091 ( new_n293_, keyIn_0_53 );
not g092 ( new_n294_, keyIn_0_28 );
xnor g093 ( new_n295_, N1, N5 );
nand g094 ( new_n296_, new_n295_, keyIn_0_0 );
nand g095 ( new_n297_, N1, N5 );
nor g096 ( new_n298_, N1, N5 );
nor g097 ( new_n299_, new_n298_, keyIn_0_0 );
nand g098 ( new_n300_, new_n299_, new_n297_ );
nand g099 ( new_n301_, new_n296_, new_n300_ );
xnor g100 ( new_n302_, N9, N13 );
nand g101 ( new_n303_, new_n302_, keyIn_0_1 );
nand g102 ( new_n304_, N9, N13 );
nor g103 ( new_n305_, N9, N13 );
nor g104 ( new_n306_, new_n305_, keyIn_0_1 );
nand g105 ( new_n307_, new_n306_, new_n304_ );
nand g106 ( new_n308_, new_n303_, new_n307_ );
nand g107 ( new_n309_, new_n301_, new_n308_ );
and g108 ( new_n310_, new_n296_, new_n300_ );
and g109 ( new_n311_, new_n303_, new_n307_ );
nand g110 ( new_n312_, new_n310_, new_n311_ );
nand g111 ( new_n313_, new_n312_, new_n309_ );
nand g112 ( new_n314_, new_n313_, new_n294_ );
and g113 ( new_n315_, new_n301_, new_n308_ );
nor g114 ( new_n316_, new_n301_, new_n308_ );
nor g115 ( new_n317_, new_n315_, new_n316_ );
nand g116 ( new_n318_, new_n317_, keyIn_0_28 );
nand g117 ( new_n319_, new_n318_, new_n314_ );
not g118 ( new_n320_, keyIn_0_4 );
xnor g119 ( new_n321_, N33, N37 );
nand g120 ( new_n322_, new_n321_, new_n320_ );
nand g121 ( new_n323_, N33, N37 );
nor g122 ( new_n324_, N33, N37 );
nor g123 ( new_n325_, new_n324_, new_n320_ );
nand g124 ( new_n326_, new_n325_, new_n323_ );
nand g125 ( new_n327_, new_n322_, new_n326_ );
xnor g126 ( new_n328_, N41, N45 );
nand g127 ( new_n329_, new_n328_, keyIn_0_5 );
nand g128 ( new_n330_, N41, N45 );
nor g129 ( new_n331_, N41, N45 );
nor g130 ( new_n332_, new_n331_, keyIn_0_5 );
nand g131 ( new_n333_, new_n332_, new_n330_ );
nand g132 ( new_n334_, new_n329_, new_n333_ );
xnor g133 ( new_n335_, new_n327_, new_n334_ );
xnor g134 ( new_n336_, new_n335_, keyIn_0_30 );
nand g135 ( new_n337_, new_n336_, new_n319_ );
xnor g136 ( new_n338_, new_n313_, keyIn_0_28 );
not g137 ( new_n339_, keyIn_0_30 );
nand g138 ( new_n340_, new_n335_, new_n339_ );
and g139 ( new_n341_, new_n327_, new_n334_ );
nor g140 ( new_n342_, new_n327_, new_n334_ );
nor g141 ( new_n343_, new_n341_, new_n342_ );
nand g142 ( new_n344_, new_n343_, keyIn_0_30 );
nand g143 ( new_n345_, new_n344_, new_n340_ );
nand g144 ( new_n346_, new_n338_, new_n345_ );
nand g145 ( new_n347_, new_n337_, new_n346_ );
nand g146 ( new_n348_, new_n347_, keyIn_0_41 );
not g147 ( new_n349_, keyIn_0_41 );
xnor g148 ( new_n350_, new_n345_, new_n319_ );
nand g149 ( new_n351_, new_n350_, new_n349_ );
nand g150 ( new_n352_, new_n351_, new_n348_ );
nand g151 ( new_n353_, N135, N137 );
nand g152 ( new_n354_, new_n353_, keyIn_0_19 );
not g153 ( new_n355_, N135 );
nor g154 ( new_n356_, new_n355_, keyIn_0_19 );
nand g155 ( new_n357_, new_n356_, N137 );
nand g156 ( new_n358_, new_n357_, new_n354_ );
nand g157 ( new_n359_, new_n352_, new_n358_ );
xnor g158 ( new_n360_, new_n347_, new_n349_ );
not g159 ( new_n361_, new_n358_ );
nand g160 ( new_n362_, new_n360_, new_n361_ );
nand g161 ( new_n363_, new_n362_, new_n359_ );
nand g162 ( new_n364_, new_n363_, new_n293_ );
xnor g163 ( new_n365_, new_n352_, new_n361_ );
nand g164 ( new_n366_, new_n365_, keyIn_0_53 );
nand g165 ( new_n367_, new_n366_, new_n364_ );
xnor g166 ( new_n368_, N73, N89 );
xnor g167 ( new_n369_, new_n368_, keyIn_0_26 );
xor g168 ( new_n370_, N105, N121 );
xnor g169 ( new_n371_, new_n370_, keyIn_0_27 );
xnor g170 ( new_n372_, new_n371_, new_n369_ );
xnor g171 ( new_n373_, new_n372_, keyIn_0_38 );
nand g172 ( new_n374_, new_n367_, new_n373_ );
xnor g173 ( new_n375_, new_n363_, keyIn_0_53 );
not g174 ( new_n376_, new_n373_ );
nand g175 ( new_n377_, new_n375_, new_n376_ );
nand g176 ( new_n378_, new_n377_, new_n374_ );
nand g177 ( new_n379_, new_n378_, new_n292_ );
xnor g178 ( new_n380_, new_n367_, new_n376_ );
nand g179 ( new_n381_, new_n380_, keyIn_0_61 );
nand g180 ( new_n382_, new_n381_, new_n379_ );
not g181 ( new_n383_, keyIn_0_29 );
not g182 ( new_n384_, keyIn_0_2 );
xnor g183 ( new_n385_, N17, N21 );
nand g184 ( new_n386_, new_n385_, new_n384_ );
nand g185 ( new_n387_, N17, N21 );
nor g186 ( new_n388_, N17, N21 );
nor g187 ( new_n389_, new_n388_, new_n384_ );
nand g188 ( new_n390_, new_n389_, new_n387_ );
nand g189 ( new_n391_, new_n386_, new_n390_ );
xnor g190 ( new_n392_, N25, N29 );
nand g191 ( new_n393_, new_n392_, keyIn_0_3 );
nand g192 ( new_n394_, N25, N29 );
nor g193 ( new_n395_, N25, N29 );
nor g194 ( new_n396_, new_n395_, keyIn_0_3 );
nand g195 ( new_n397_, new_n396_, new_n394_ );
nand g196 ( new_n398_, new_n393_, new_n397_ );
xnor g197 ( new_n399_, new_n391_, new_n398_ );
nand g198 ( new_n400_, new_n399_, new_n383_ );
and g199 ( new_n401_, new_n391_, new_n398_ );
nor g200 ( new_n402_, new_n391_, new_n398_ );
nor g201 ( new_n403_, new_n401_, new_n402_ );
nand g202 ( new_n404_, new_n403_, keyIn_0_29 );
nand g203 ( new_n405_, new_n404_, new_n400_ );
not g204 ( new_n406_, keyIn_0_31 );
xnor g205 ( new_n407_, N49, N53 );
nand g206 ( new_n408_, new_n407_, keyIn_0_6 );
nand g207 ( new_n409_, N49, N53 );
nor g208 ( new_n410_, N49, N53 );
nor g209 ( new_n411_, new_n410_, keyIn_0_6 );
nand g210 ( new_n412_, new_n411_, new_n409_ );
nand g211 ( new_n413_, new_n408_, new_n412_ );
xnor g212 ( new_n414_, N57, N61 );
nand g213 ( new_n415_, new_n414_, keyIn_0_7 );
nand g214 ( new_n416_, N57, N61 );
nor g215 ( new_n417_, N57, N61 );
nor g216 ( new_n418_, new_n417_, keyIn_0_7 );
nand g217 ( new_n419_, new_n418_, new_n416_ );
nand g218 ( new_n420_, new_n415_, new_n419_ );
nand g219 ( new_n421_, new_n413_, new_n420_ );
and g220 ( new_n422_, new_n408_, new_n412_ );
and g221 ( new_n423_, new_n415_, new_n419_ );
nand g222 ( new_n424_, new_n422_, new_n423_ );
nand g223 ( new_n425_, new_n424_, new_n421_ );
nand g224 ( new_n426_, new_n425_, new_n406_ );
and g225 ( new_n427_, new_n413_, new_n420_ );
nor g226 ( new_n428_, new_n413_, new_n420_ );
nor g227 ( new_n429_, new_n427_, new_n428_ );
nand g228 ( new_n430_, new_n429_, keyIn_0_31 );
nand g229 ( new_n431_, new_n430_, new_n426_ );
xnor g230 ( new_n432_, new_n405_, new_n431_ );
xnor g231 ( new_n433_, new_n432_, keyIn_0_42 );
nand g232 ( new_n434_, N136, N137 );
nand g233 ( new_n435_, new_n434_, keyIn_0_20 );
not g234 ( new_n436_, N136 );
nor g235 ( new_n437_, new_n436_, keyIn_0_20 );
nand g236 ( new_n438_, new_n437_, N137 );
nand g237 ( new_n439_, new_n438_, new_n435_ );
nand g238 ( new_n440_, new_n433_, new_n439_ );
not g239 ( new_n441_, keyIn_0_42 );
xnor g240 ( new_n442_, new_n432_, new_n441_ );
not g241 ( new_n443_, new_n439_ );
nand g242 ( new_n444_, new_n442_, new_n443_ );
nand g243 ( new_n445_, new_n444_, new_n440_ );
xnor g244 ( new_n446_, new_n445_, keyIn_0_54 );
xor g245 ( new_n447_, N77, N93 );
xnor g246 ( new_n448_, N109, N125 );
xnor g247 ( new_n449_, new_n447_, new_n448_ );
nand g248 ( new_n450_, new_n446_, new_n449_ );
not g249 ( new_n451_, keyIn_0_54 );
xnor g250 ( new_n452_, new_n445_, new_n451_ );
not g251 ( new_n453_, new_n449_ );
nand g252 ( new_n454_, new_n452_, new_n453_ );
nand g253 ( new_n455_, new_n454_, new_n450_ );
xnor g254 ( new_n456_, new_n455_, keyIn_0_62 );
not g255 ( new_n457_, keyIn_0_51 );
xnor g256 ( new_n458_, new_n405_, new_n319_ );
nand g257 ( new_n459_, new_n458_, keyIn_0_39 );
not g258 ( new_n460_, keyIn_0_39 );
xnor g259 ( new_n461_, new_n338_, new_n405_ );
nand g260 ( new_n462_, new_n461_, new_n460_ );
nand g261 ( new_n463_, new_n462_, new_n459_ );
and g262 ( new_n464_, N133, N137 );
or g263 ( new_n465_, new_n464_, keyIn_0_17 );
not g264 ( new_n466_, new_n465_ );
nand g265 ( new_n467_, keyIn_0_17, N133 );
nor g266 ( new_n468_, new_n467_, new_n265_ );
nor g267 ( new_n469_, new_n466_, new_n468_ );
nand g268 ( new_n470_, new_n463_, new_n469_ );
xnor g269 ( new_n471_, new_n458_, new_n460_ );
not g270 ( new_n472_, new_n469_ );
nand g271 ( new_n473_, new_n471_, new_n472_ );
nand g272 ( new_n474_, new_n473_, new_n470_ );
nand g273 ( new_n475_, new_n474_, new_n457_ );
xnor g274 ( new_n476_, new_n463_, new_n472_ );
nand g275 ( new_n477_, new_n476_, keyIn_0_51 );
nand g276 ( new_n478_, new_n477_, new_n475_ );
xnor g277 ( new_n479_, N65, N81 );
xnor g278 ( new_n480_, N97, N113 );
xnor g279 ( new_n481_, new_n479_, new_n480_ );
not g280 ( new_n482_, new_n481_ );
nand g281 ( new_n483_, new_n478_, new_n482_ );
xnor g282 ( new_n484_, new_n474_, keyIn_0_51 );
nand g283 ( new_n485_, new_n484_, new_n481_ );
nand g284 ( new_n486_, new_n485_, new_n483_ );
nand g285 ( new_n487_, new_n486_, keyIn_0_59 );
not g286 ( new_n488_, keyIn_0_59 );
xnor g287 ( new_n489_, new_n478_, new_n481_ );
nand g288 ( new_n490_, new_n489_, new_n488_ );
nand g289 ( new_n491_, new_n490_, new_n487_ );
not g290 ( new_n492_, keyIn_0_52 );
nand g291 ( new_n493_, new_n345_, new_n431_ );
xnor g292 ( new_n494_, new_n425_, keyIn_0_31 );
nand g293 ( new_n495_, new_n336_, new_n494_ );
nand g294 ( new_n496_, new_n495_, new_n493_ );
nand g295 ( new_n497_, new_n496_, keyIn_0_40 );
not g296 ( new_n498_, keyIn_0_40 );
and g297 ( new_n499_, new_n345_, new_n431_ );
nor g298 ( new_n500_, new_n345_, new_n431_ );
nor g299 ( new_n501_, new_n499_, new_n500_ );
nand g300 ( new_n502_, new_n501_, new_n498_ );
nand g301 ( new_n503_, new_n502_, new_n497_ );
and g302 ( new_n504_, N134, N137 );
or g303 ( new_n505_, new_n504_, keyIn_0_18 );
not g304 ( new_n506_, new_n505_ );
nand g305 ( new_n507_, keyIn_0_18, N134 );
nor g306 ( new_n508_, new_n507_, new_n265_ );
nor g307 ( new_n509_, new_n506_, new_n508_ );
nand g308 ( new_n510_, new_n503_, new_n509_ );
xnor g309 ( new_n511_, new_n496_, new_n498_ );
not g310 ( new_n512_, new_n509_ );
nand g311 ( new_n513_, new_n511_, new_n512_ );
nand g312 ( new_n514_, new_n513_, new_n510_ );
nand g313 ( new_n515_, new_n514_, new_n492_ );
xnor g314 ( new_n516_, new_n503_, new_n512_ );
nand g315 ( new_n517_, new_n516_, keyIn_0_52 );
nand g316 ( new_n518_, new_n517_, new_n515_ );
xnor g317 ( new_n519_, N101, N117 );
xnor g318 ( new_n520_, new_n519_, keyIn_0_25 );
xor g319 ( new_n521_, N69, N85 );
xnor g320 ( new_n522_, new_n521_, keyIn_0_24 );
xnor g321 ( new_n523_, new_n522_, new_n520_ );
xnor g322 ( new_n524_, new_n523_, keyIn_0_37 );
not g323 ( new_n525_, new_n524_ );
nand g324 ( new_n526_, new_n518_, new_n525_ );
xnor g325 ( new_n527_, new_n514_, keyIn_0_52 );
nand g326 ( new_n528_, new_n527_, new_n524_ );
nand g327 ( new_n529_, new_n528_, new_n526_ );
nand g328 ( new_n530_, new_n529_, keyIn_0_60 );
not g329 ( new_n531_, keyIn_0_60 );
xnor g330 ( new_n532_, new_n518_, new_n524_ );
nand g331 ( new_n533_, new_n532_, new_n531_ );
nand g332 ( new_n534_, new_n533_, new_n530_ );
nor g333 ( new_n535_, new_n491_, new_n534_ );
nand g334 ( new_n536_, new_n535_, new_n456_ );
nor g335 ( new_n537_, new_n536_, new_n382_ );
nand g336 ( new_n538_, new_n291_, new_n537_ );
nor g337 ( new_n539_, new_n538_, new_n223_ );
xor g338 ( N724, new_n539_, N1 );
nor g339 ( new_n541_, new_n538_, new_n259_ );
xor g340 ( N725, new_n541_, N5 );
nor g341 ( new_n543_, new_n538_, new_n279_ );
xor g342 ( N726, new_n543_, N9 );
nor g343 ( new_n545_, new_n538_, new_n243_ );
xor g344 ( N727, new_n545_, N13 );
not g345 ( new_n547_, new_n223_ );
not g346 ( new_n548_, keyIn_0_76 );
xnor g347 ( new_n549_, new_n486_, new_n488_ );
xnor g348 ( new_n550_, new_n529_, new_n531_ );
nand g349 ( new_n551_, new_n549_, new_n550_ );
xnor g350 ( new_n552_, new_n378_, keyIn_0_61 );
nor g351 ( new_n553_, new_n456_, new_n552_ );
not g352 ( new_n554_, new_n553_ );
nor g353 ( new_n555_, new_n554_, new_n551_ );
nand g354 ( new_n556_, new_n291_, new_n555_ );
xnor g355 ( new_n557_, new_n556_, new_n548_ );
nand g356 ( new_n558_, new_n557_, new_n547_ );
xnor g357 ( new_n559_, new_n558_, keyIn_0_82 );
xnor g358 ( new_n560_, new_n559_, N17 );
xnor g359 ( N728, new_n560_, keyIn_0_105 );
not g360 ( new_n562_, keyIn_0_106 );
nand g361 ( new_n563_, new_n557_, new_n283_ );
xnor g362 ( new_n564_, new_n563_, keyIn_0_83 );
xnor g363 ( new_n565_, new_n564_, N21 );
xnor g364 ( N729, new_n565_, new_n562_ );
nand g365 ( new_n567_, new_n557_, new_n280_ );
xnor g366 ( N730, new_n567_, N25 );
not g367 ( new_n569_, keyIn_0_107 );
not g368 ( new_n570_, keyIn_0_84 );
nand g369 ( new_n571_, new_n557_, new_n242_ );
xnor g370 ( new_n572_, new_n571_, new_n570_ );
xnor g371 ( new_n573_, new_n572_, N29 );
xnor g372 ( N731, new_n573_, new_n569_ );
not g373 ( new_n575_, keyIn_0_77 );
not g374 ( new_n576_, keyIn_0_62 );
xnor g375 ( new_n577_, new_n455_, new_n576_ );
nand g376 ( new_n578_, new_n491_, new_n534_ );
nor g377 ( new_n579_, new_n578_, new_n577_ );
and g378 ( new_n580_, new_n579_, new_n552_ );
nand g379 ( new_n581_, new_n291_, new_n580_ );
xnor g380 ( new_n582_, new_n581_, new_n575_ );
nand g381 ( new_n583_, new_n582_, new_n547_ );
xnor g382 ( new_n584_, new_n583_, keyIn_0_85 );
xnor g383 ( new_n585_, new_n584_, N33 );
xnor g384 ( N732, new_n585_, keyIn_0_108 );
not g385 ( new_n587_, keyIn_0_109 );
not g386 ( new_n588_, keyIn_0_86 );
nand g387 ( new_n589_, new_n582_, new_n283_ );
xnor g388 ( new_n590_, new_n589_, new_n588_ );
xnor g389 ( new_n591_, new_n590_, N37 );
xnor g390 ( N733, new_n591_, new_n587_ );
nand g391 ( new_n593_, new_n582_, new_n280_ );
xnor g392 ( new_n594_, new_n593_, keyIn_0_87 );
xnor g393 ( new_n595_, new_n594_, N41 );
xnor g394 ( N734, new_n595_, keyIn_0_110 );
nand g395 ( new_n597_, new_n582_, new_n242_ );
xnor g396 ( new_n598_, new_n597_, keyIn_0_88 );
xnor g397 ( new_n599_, new_n598_, N45 );
xnor g398 ( N735, new_n599_, keyIn_0_111 );
nor g399 ( new_n601_, new_n554_, new_n578_ );
nand g400 ( new_n602_, new_n291_, new_n601_ );
nor g401 ( new_n603_, new_n602_, new_n223_ );
xor g402 ( N736, new_n603_, N49 );
nor g403 ( new_n605_, new_n602_, new_n259_ );
xor g404 ( N737, new_n605_, N53 );
nor g405 ( new_n607_, new_n602_, new_n279_ );
xor g406 ( N738, new_n607_, N57 );
nor g407 ( new_n609_, new_n602_, new_n243_ );
xor g408 ( N739, new_n609_, N61 );
not g409 ( new_n611_, N65 );
not g410 ( new_n612_, keyIn_0_89 );
not g411 ( new_n613_, keyIn_0_78 );
nor g412 ( new_n614_, new_n549_, new_n534_ );
nor g413 ( new_n615_, new_n577_, new_n382_ );
nand g414 ( new_n616_, new_n615_, new_n614_ );
xnor g415 ( new_n617_, new_n616_, keyIn_0_72 );
nor g416 ( new_n618_, new_n551_, new_n577_ );
xnor g417 ( new_n619_, new_n382_, keyIn_0_66 );
nand g418 ( new_n620_, new_n618_, new_n619_ );
nand g419 ( new_n621_, new_n620_, keyIn_0_74 );
not g420 ( new_n622_, keyIn_0_74 );
not g421 ( new_n623_, keyIn_0_66 );
xnor g422 ( new_n624_, new_n382_, new_n623_ );
nor g423 ( new_n625_, new_n624_, new_n536_ );
nand g424 ( new_n626_, new_n625_, new_n622_ );
nand g425 ( new_n627_, new_n626_, new_n621_ );
nand g426 ( new_n628_, new_n627_, new_n617_ );
nand g427 ( new_n629_, new_n550_, new_n491_ );
nor g428 ( new_n630_, new_n629_, new_n456_ );
xnor g429 ( new_n631_, new_n382_, keyIn_0_64 );
nand g430 ( new_n632_, new_n631_, new_n630_ );
xnor g431 ( new_n633_, new_n632_, keyIn_0_71 );
not g432 ( new_n634_, keyIn_0_73 );
nand g433 ( new_n635_, new_n382_, keyIn_0_65 );
not g434 ( new_n636_, keyIn_0_65 );
nand g435 ( new_n637_, new_n552_, new_n636_ );
nand g436 ( new_n638_, new_n637_, new_n635_ );
nand g437 ( new_n639_, new_n579_, new_n638_ );
xnor g438 ( new_n640_, new_n639_, new_n634_ );
nand g439 ( new_n641_, new_n633_, new_n640_ );
nor g440 ( new_n642_, new_n641_, new_n628_ );
nand g441 ( new_n643_, new_n642_, keyIn_0_75 );
not g442 ( new_n644_, keyIn_0_75 );
and g443 ( new_n645_, new_n627_, new_n617_ );
not g444 ( new_n646_, keyIn_0_71 );
xnor g445 ( new_n647_, new_n632_, new_n646_ );
xnor g446 ( new_n648_, new_n639_, keyIn_0_73 );
nor g447 ( new_n649_, new_n647_, new_n648_ );
nand g448 ( new_n650_, new_n645_, new_n649_ );
nand g449 ( new_n651_, new_n650_, new_n644_ );
nand g450 ( new_n652_, new_n651_, new_n643_ );
nor g451 ( new_n653_, new_n279_, new_n242_ );
nand g452 ( new_n654_, new_n653_, new_n547_ );
xor g453 ( new_n655_, new_n259_, keyIn_0_67 );
nor g454 ( new_n656_, new_n655_, new_n654_ );
nand g455 ( new_n657_, new_n652_, new_n656_ );
xnor g456 ( new_n658_, new_n657_, new_n613_ );
nand g457 ( new_n659_, new_n658_, new_n549_ );
nand g458 ( new_n660_, new_n659_, new_n612_ );
xnor g459 ( new_n661_, new_n657_, keyIn_0_78 );
nor g460 ( new_n662_, new_n661_, new_n491_ );
nand g461 ( new_n663_, new_n662_, keyIn_0_89 );
nand g462 ( new_n664_, new_n663_, new_n660_ );
nand g463 ( new_n665_, new_n664_, new_n611_ );
xnor g464 ( new_n666_, new_n659_, keyIn_0_89 );
nand g465 ( new_n667_, new_n666_, N65 );
nand g466 ( new_n668_, new_n667_, new_n665_ );
nand g467 ( new_n669_, new_n668_, keyIn_0_112 );
not g468 ( new_n670_, keyIn_0_112 );
xnor g469 ( new_n671_, new_n664_, N65 );
nand g470 ( new_n672_, new_n671_, new_n670_ );
nand g471 ( N740, new_n672_, new_n669_ );
not g472 ( new_n674_, keyIn_0_113 );
not g473 ( new_n675_, N69 );
nand g474 ( new_n676_, new_n658_, new_n534_ );
nand g475 ( new_n677_, new_n676_, keyIn_0_90 );
not g476 ( new_n678_, keyIn_0_90 );
nor g477 ( new_n679_, new_n661_, new_n550_ );
nand g478 ( new_n680_, new_n679_, new_n678_ );
nand g479 ( new_n681_, new_n680_, new_n677_ );
nand g480 ( new_n682_, new_n681_, new_n675_ );
xnor g481 ( new_n683_, new_n676_, new_n678_ );
nand g482 ( new_n684_, new_n683_, N69 );
nand g483 ( new_n685_, new_n684_, new_n682_ );
nand g484 ( new_n686_, new_n685_, new_n674_ );
xnor g485 ( new_n687_, new_n681_, N69 );
nand g486 ( new_n688_, new_n687_, keyIn_0_113 );
nand g487 ( N741, new_n688_, new_n686_ );
not g488 ( new_n690_, keyIn_0_114 );
not g489 ( new_n691_, N73 );
nand g490 ( new_n692_, new_n658_, new_n552_ );
nand g491 ( new_n693_, new_n692_, keyIn_0_91 );
not g492 ( new_n694_, keyIn_0_91 );
nor g493 ( new_n695_, new_n661_, new_n382_ );
nand g494 ( new_n696_, new_n695_, new_n694_ );
nand g495 ( new_n697_, new_n696_, new_n693_ );
nand g496 ( new_n698_, new_n697_, new_n691_ );
xnor g497 ( new_n699_, new_n692_, new_n694_ );
nand g498 ( new_n700_, new_n699_, N73 );
nand g499 ( new_n701_, new_n700_, new_n698_ );
nand g500 ( new_n702_, new_n701_, new_n690_ );
xnor g501 ( new_n703_, new_n697_, N73 );
nand g502 ( new_n704_, new_n703_, keyIn_0_114 );
nand g503 ( N742, new_n704_, new_n702_ );
not g504 ( new_n706_, N77 );
nand g505 ( new_n707_, new_n658_, new_n577_ );
nand g506 ( new_n708_, new_n707_, keyIn_0_92 );
not g507 ( new_n709_, keyIn_0_92 );
nor g508 ( new_n710_, new_n661_, new_n456_ );
nand g509 ( new_n711_, new_n710_, new_n709_ );
nand g510 ( new_n712_, new_n711_, new_n708_ );
nand g511 ( new_n713_, new_n712_, new_n706_ );
xnor g512 ( new_n714_, new_n707_, new_n709_ );
nand g513 ( new_n715_, new_n714_, N77 );
nand g514 ( new_n716_, new_n715_, new_n713_ );
nand g515 ( new_n717_, new_n716_, keyIn_0_115 );
not g516 ( new_n718_, keyIn_0_115 );
xnor g517 ( new_n719_, new_n712_, N77 );
nand g518 ( new_n720_, new_n719_, new_n718_ );
nand g519 ( N743, new_n720_, new_n717_ );
not g520 ( new_n722_, keyIn_0_116 );
not g521 ( new_n723_, N81 );
nor g522 ( new_n724_, new_n243_, new_n223_ );
nand g523 ( new_n725_, new_n724_, new_n259_ );
xnor g524 ( new_n726_, new_n279_, keyIn_0_68 );
nor g525 ( new_n727_, new_n725_, new_n726_ );
nand g526 ( new_n728_, new_n652_, new_n727_ );
xnor g527 ( new_n729_, new_n728_, keyIn_0_79 );
nand g528 ( new_n730_, new_n729_, new_n549_ );
nand g529 ( new_n731_, new_n730_, keyIn_0_93 );
not g530 ( new_n732_, keyIn_0_93 );
not g531 ( new_n733_, keyIn_0_79 );
xnor g532 ( new_n734_, new_n728_, new_n733_ );
nor g533 ( new_n735_, new_n734_, new_n491_ );
nand g534 ( new_n736_, new_n735_, new_n732_ );
nand g535 ( new_n737_, new_n736_, new_n731_ );
nand g536 ( new_n738_, new_n737_, new_n723_ );
xnor g537 ( new_n739_, new_n730_, new_n732_ );
nand g538 ( new_n740_, new_n739_, N81 );
nand g539 ( new_n741_, new_n740_, new_n738_ );
nand g540 ( new_n742_, new_n741_, new_n722_ );
xnor g541 ( new_n743_, new_n737_, N81 );
nand g542 ( new_n744_, new_n743_, keyIn_0_116 );
nand g543 ( N744, new_n744_, new_n742_ );
not g544 ( new_n746_, N85 );
nand g545 ( new_n747_, new_n729_, new_n534_ );
nand g546 ( new_n748_, new_n747_, keyIn_0_94 );
not g547 ( new_n749_, keyIn_0_94 );
nor g548 ( new_n750_, new_n734_, new_n550_ );
nand g549 ( new_n751_, new_n750_, new_n749_ );
nand g550 ( new_n752_, new_n751_, new_n748_ );
nand g551 ( new_n753_, new_n752_, new_n746_ );
xnor g552 ( new_n754_, new_n747_, new_n749_ );
nand g553 ( new_n755_, new_n754_, N85 );
nand g554 ( new_n756_, new_n755_, new_n753_ );
nand g555 ( new_n757_, new_n756_, keyIn_0_117 );
not g556 ( new_n758_, keyIn_0_117 );
xnor g557 ( new_n759_, new_n752_, N85 );
nand g558 ( new_n760_, new_n759_, new_n758_ );
nand g559 ( N745, new_n760_, new_n757_ );
not g560 ( new_n762_, keyIn_0_118 );
not g561 ( new_n763_, N89 );
nand g562 ( new_n764_, new_n729_, new_n552_ );
nand g563 ( new_n765_, new_n764_, keyIn_0_95 );
not g564 ( new_n766_, keyIn_0_95 );
nor g565 ( new_n767_, new_n734_, new_n382_ );
nand g566 ( new_n768_, new_n767_, new_n766_ );
nand g567 ( new_n769_, new_n768_, new_n765_ );
nand g568 ( new_n770_, new_n769_, new_n763_ );
xnor g569 ( new_n771_, new_n764_, new_n766_ );
nand g570 ( new_n772_, new_n771_, N89 );
nand g571 ( new_n773_, new_n772_, new_n770_ );
nand g572 ( new_n774_, new_n773_, new_n762_ );
xnor g573 ( new_n775_, new_n769_, N89 );
nand g574 ( new_n776_, new_n775_, keyIn_0_118 );
nand g575 ( N746, new_n776_, new_n774_ );
not g576 ( new_n778_, keyIn_0_119 );
not g577 ( new_n779_, N93 );
nand g578 ( new_n780_, new_n729_, new_n577_ );
nand g579 ( new_n781_, new_n780_, keyIn_0_96 );
not g580 ( new_n782_, keyIn_0_96 );
nor g581 ( new_n783_, new_n734_, new_n456_ );
nand g582 ( new_n784_, new_n783_, new_n782_ );
nand g583 ( new_n785_, new_n784_, new_n781_ );
nand g584 ( new_n786_, new_n785_, new_n779_ );
xnor g585 ( new_n787_, new_n780_, new_n782_ );
nand g586 ( new_n788_, new_n787_, N93 );
nand g587 ( new_n789_, new_n788_, new_n786_ );
nand g588 ( new_n790_, new_n789_, new_n778_ );
xnor g589 ( new_n791_, new_n785_, N93 );
nand g590 ( new_n792_, new_n791_, keyIn_0_119 );
nand g591 ( N747, new_n792_, new_n790_ );
not g592 ( new_n794_, keyIn_0_120 );
not g593 ( new_n795_, keyIn_0_80 );
nor g594 ( new_n796_, new_n547_, new_n259_ );
and g595 ( new_n797_, new_n796_, new_n653_ );
nand g596 ( new_n798_, new_n652_, new_n797_ );
xnor g597 ( new_n799_, new_n798_, new_n795_ );
nand g598 ( new_n800_, new_n799_, new_n549_ );
nand g599 ( new_n801_, new_n800_, keyIn_0_97 );
not g600 ( new_n802_, keyIn_0_97 );
xnor g601 ( new_n803_, new_n798_, keyIn_0_80 );
nor g602 ( new_n804_, new_n803_, new_n491_ );
nand g603 ( new_n805_, new_n804_, new_n802_ );
nand g604 ( new_n806_, new_n805_, new_n801_ );
nand g605 ( new_n807_, new_n806_, N97 );
not g606 ( new_n808_, N97 );
xnor g607 ( new_n809_, new_n800_, new_n802_ );
nand g608 ( new_n810_, new_n809_, new_n808_ );
nand g609 ( new_n811_, new_n810_, new_n807_ );
nand g610 ( new_n812_, new_n811_, new_n794_ );
xnor g611 ( new_n813_, new_n806_, new_n808_ );
nand g612 ( new_n814_, new_n813_, keyIn_0_120 );
nand g613 ( N748, new_n814_, new_n812_ );
not g614 ( new_n816_, N101 );
nand g615 ( new_n817_, new_n799_, new_n534_ );
nand g616 ( new_n818_, new_n817_, keyIn_0_98 );
not g617 ( new_n819_, keyIn_0_98 );
nor g618 ( new_n820_, new_n803_, new_n550_ );
nand g619 ( new_n821_, new_n820_, new_n819_ );
nand g620 ( new_n822_, new_n821_, new_n818_ );
nand g621 ( new_n823_, new_n822_, new_n816_ );
xnor g622 ( new_n824_, new_n817_, new_n819_ );
nand g623 ( new_n825_, new_n824_, N101 );
nand g624 ( new_n826_, new_n825_, new_n823_ );
nand g625 ( new_n827_, new_n826_, keyIn_0_121 );
not g626 ( new_n828_, keyIn_0_121 );
xnor g627 ( new_n829_, new_n822_, N101 );
nand g628 ( new_n830_, new_n829_, new_n828_ );
nand g629 ( N749, new_n830_, new_n827_ );
nand g630 ( new_n832_, new_n799_, new_n552_ );
nand g631 ( new_n833_, new_n832_, keyIn_0_99 );
not g632 ( new_n834_, keyIn_0_99 );
nor g633 ( new_n835_, new_n803_, new_n382_ );
nand g634 ( new_n836_, new_n835_, new_n834_ );
nand g635 ( new_n837_, new_n836_, new_n833_ );
nand g636 ( new_n838_, new_n837_, N105 );
not g637 ( new_n839_, N105 );
xnor g638 ( new_n840_, new_n832_, new_n834_ );
nand g639 ( new_n841_, new_n840_, new_n839_ );
nand g640 ( new_n842_, new_n841_, new_n838_ );
nand g641 ( new_n843_, new_n842_, keyIn_0_122 );
not g642 ( new_n844_, keyIn_0_122 );
xnor g643 ( new_n845_, new_n837_, new_n839_ );
nand g644 ( new_n846_, new_n845_, new_n844_ );
nand g645 ( N750, new_n846_, new_n843_ );
not g646 ( new_n848_, keyIn_0_123 );
nand g647 ( new_n849_, new_n799_, new_n577_ );
nand g648 ( new_n850_, new_n849_, keyIn_0_100 );
not g649 ( new_n851_, keyIn_0_100 );
nor g650 ( new_n852_, new_n803_, new_n456_ );
nand g651 ( new_n853_, new_n852_, new_n851_ );
nand g652 ( new_n854_, new_n853_, new_n850_ );
nand g653 ( new_n855_, new_n854_, N109 );
not g654 ( new_n856_, N109 );
xnor g655 ( new_n857_, new_n849_, new_n851_ );
nand g656 ( new_n858_, new_n857_, new_n856_ );
nand g657 ( new_n859_, new_n858_, new_n855_ );
nand g658 ( new_n860_, new_n859_, new_n848_ );
xnor g659 ( new_n861_, new_n854_, new_n856_ );
nand g660 ( new_n862_, new_n861_, keyIn_0_123 );
nand g661 ( N751, new_n862_, new_n860_ );
not g662 ( new_n864_, N113 );
not g663 ( new_n865_, keyIn_0_81 );
and g664 ( new_n866_, new_n547_, keyIn_0_69 );
or g665 ( new_n867_, new_n866_, new_n284_ );
not g666 ( new_n868_, keyIn_0_70 );
nand g667 ( new_n869_, new_n280_, new_n868_ );
nor g668 ( new_n870_, new_n280_, new_n868_ );
nor g669 ( new_n871_, new_n547_, keyIn_0_69 );
nor g670 ( new_n872_, new_n871_, new_n870_ );
nand g671 ( new_n873_, new_n872_, new_n869_ );
nor g672 ( new_n874_, new_n873_, new_n867_ );
nand g673 ( new_n875_, new_n652_, new_n874_ );
xnor g674 ( new_n876_, new_n875_, new_n865_ );
nand g675 ( new_n877_, new_n876_, new_n549_ );
nand g676 ( new_n878_, new_n877_, keyIn_0_101 );
not g677 ( new_n879_, keyIn_0_101 );
xnor g678 ( new_n880_, new_n875_, keyIn_0_81 );
nor g679 ( new_n881_, new_n880_, new_n491_ );
nand g680 ( new_n882_, new_n881_, new_n879_ );
nand g681 ( new_n883_, new_n882_, new_n878_ );
nand g682 ( new_n884_, new_n883_, new_n864_ );
xnor g683 ( new_n885_, new_n877_, new_n879_ );
nand g684 ( new_n886_, new_n885_, N113 );
nand g685 ( new_n887_, new_n886_, new_n884_ );
nand g686 ( new_n888_, new_n887_, keyIn_0_124 );
not g687 ( new_n889_, keyIn_0_124 );
xnor g688 ( new_n890_, new_n883_, N113 );
nand g689 ( new_n891_, new_n890_, new_n889_ );
nand g690 ( N752, new_n891_, new_n888_ );
not g691 ( new_n893_, keyIn_0_125 );
not g692 ( new_n894_, N117 );
nand g693 ( new_n895_, new_n876_, new_n534_ );
nand g694 ( new_n896_, new_n895_, keyIn_0_102 );
not g695 ( new_n897_, keyIn_0_102 );
nor g696 ( new_n898_, new_n880_, new_n550_ );
nand g697 ( new_n899_, new_n898_, new_n897_ );
nand g698 ( new_n900_, new_n899_, new_n896_ );
nand g699 ( new_n901_, new_n900_, new_n894_ );
xnor g700 ( new_n902_, new_n895_, new_n897_ );
nand g701 ( new_n903_, new_n902_, N117 );
nand g702 ( new_n904_, new_n903_, new_n901_ );
nand g703 ( new_n905_, new_n904_, new_n893_ );
xnor g704 ( new_n906_, new_n900_, N117 );
nand g705 ( new_n907_, new_n906_, keyIn_0_125 );
nand g706 ( N753, new_n907_, new_n905_ );
not g707 ( new_n909_, N121 );
not g708 ( new_n910_, keyIn_0_103 );
nand g709 ( new_n911_, new_n876_, new_n552_ );
nand g710 ( new_n912_, new_n911_, new_n910_ );
nor g711 ( new_n913_, new_n880_, new_n382_ );
nand g712 ( new_n914_, new_n913_, keyIn_0_103 );
nand g713 ( new_n915_, new_n914_, new_n912_ );
nand g714 ( new_n916_, new_n915_, new_n909_ );
xnor g715 ( new_n917_, new_n911_, keyIn_0_103 );
nand g716 ( new_n918_, new_n917_, N121 );
nand g717 ( new_n919_, new_n918_, new_n916_ );
nand g718 ( new_n920_, new_n919_, keyIn_0_126 );
not g719 ( new_n921_, keyIn_0_126 );
xnor g720 ( new_n922_, new_n915_, N121 );
nand g721 ( new_n923_, new_n922_, new_n921_ );
nand g722 ( N754, new_n923_, new_n920_ );
not g723 ( new_n925_, keyIn_0_127 );
not g724 ( new_n926_, N125 );
nand g725 ( new_n927_, new_n876_, new_n577_ );
nand g726 ( new_n928_, new_n927_, keyIn_0_104 );
not g727 ( new_n929_, keyIn_0_104 );
nor g728 ( new_n930_, new_n880_, new_n456_ );
nand g729 ( new_n931_, new_n930_, new_n929_ );
nand g730 ( new_n932_, new_n931_, new_n928_ );
nand g731 ( new_n933_, new_n932_, new_n926_ );
xnor g732 ( new_n934_, new_n927_, new_n929_ );
nand g733 ( new_n935_, new_n934_, N125 );
nand g734 ( new_n936_, new_n935_, new_n933_ );
nand g735 ( new_n937_, new_n936_, new_n925_ );
xnor g736 ( new_n938_, new_n932_, N125 );
nand g737 ( new_n939_, new_n938_, keyIn_0_127 );
nand g738 ( N755, new_n939_, new_n937_ );
endmodule