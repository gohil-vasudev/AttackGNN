module add_mul_combine_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_mul_0_, Result_mul_1_, Result_mul_2_, 
        Result_mul_3_, Result_mul_4_, Result_mul_5_, Result_mul_6_, 
        Result_mul_7_, Result_mul_8_, Result_mul_9_, Result_mul_10_, 
        Result_mul_11_, Result_mul_12_, Result_mul_13_, Result_mul_14_, 
        Result_mul_15_, Result_mul_16_, Result_mul_17_, Result_mul_18_, 
        Result_mul_19_, Result_mul_20_, Result_mul_21_, Result_mul_22_, 
        Result_mul_23_, Result_mul_24_, Result_mul_25_, Result_mul_26_, 
        Result_mul_27_, Result_mul_28_, Result_mul_29_, Result_mul_30_, 
        Result_mul_31_, Result_add_0_, Result_add_1_, Result_add_2_, 
        Result_add_3_, Result_add_4_, Result_add_5_, Result_add_6_, 
        Result_add_7_, Result_add_8_, Result_add_9_, Result_add_10_, 
        Result_add_11_, Result_add_12_, Result_add_13_, Result_add_14_, 
        Result_add_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_;
  wire   n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687;

  XOR2_X1 U1882 ( .A(n1834), .B(n1835), .Z(Result_mul_9_) );
  AND2_X1 U1883 ( .A1(n1836), .A2(n1837), .ZN(n1835) );
  OR2_X1 U1884 ( .A1(n1838), .A2(n1839), .ZN(n1837) );
  AND2_X1 U1885 ( .A1(n1840), .A2(n1841), .ZN(n1839) );
  INV_X1 U1886 ( .A(n1842), .ZN(n1836) );
  XOR2_X1 U1887 ( .A(n1843), .B(n1844), .Z(Result_mul_8_) );
  XOR2_X1 U1888 ( .A(n1845), .B(n1846), .Z(Result_mul_7_) );
  AND2_X1 U1889 ( .A1(n1847), .A2(n1848), .ZN(n1846) );
  OR2_X1 U1890 ( .A1(n1849), .A2(n1850), .ZN(n1848) );
  AND2_X1 U1891 ( .A1(n1851), .A2(n1852), .ZN(n1850) );
  INV_X1 U1892 ( .A(n1853), .ZN(n1847) );
  XOR2_X1 U1893 ( .A(n1854), .B(n1855), .Z(Result_mul_6_) );
  XOR2_X1 U1894 ( .A(n1856), .B(n1857), .Z(Result_mul_5_) );
  AND2_X1 U1895 ( .A1(n1858), .A2(n1859), .ZN(n1857) );
  OR2_X1 U1896 ( .A1(n1860), .A2(n1861), .ZN(n1859) );
  AND2_X1 U1897 ( .A1(n1862), .A2(n1863), .ZN(n1861) );
  INV_X1 U1898 ( .A(n1864), .ZN(n1858) );
  XOR2_X1 U1899 ( .A(n1865), .B(n1866), .Z(Result_mul_4_) );
  XOR2_X1 U1900 ( .A(n1867), .B(n1868), .Z(Result_mul_3_) );
  AND2_X1 U1901 ( .A1(n1869), .A2(n1870), .ZN(n1868) );
  OR2_X1 U1902 ( .A1(n1871), .A2(n1872), .ZN(n1870) );
  AND2_X1 U1903 ( .A1(n1873), .A2(n1874), .ZN(n1872) );
  INV_X1 U1904 ( .A(n1875), .ZN(n1869) );
  OR2_X1 U1905 ( .A1(n1876), .A2(n1877), .ZN(Result_mul_30_) );
  AND2_X1 U1906 ( .A1(b_15_), .A2(n1878), .ZN(n1877) );
  OR2_X1 U1907 ( .A1(n1879), .A2(n1880), .ZN(n1878) );
  AND2_X1 U1908 ( .A1(a_14_), .A2(n1881), .ZN(n1879) );
  AND2_X1 U1909 ( .A1(b_14_), .A2(n1882), .ZN(n1876) );
  OR2_X1 U1910 ( .A1(n1883), .A2(n1884), .ZN(n1882) );
  AND2_X1 U1911 ( .A1(a_15_), .A2(n1885), .ZN(n1883) );
  XOR2_X1 U1912 ( .A(n1886), .B(n1887), .Z(Result_mul_2_) );
  XNOR2_X1 U1913 ( .A(n1888), .B(n1889), .ZN(Result_mul_29_) );
  XNOR2_X1 U1914 ( .A(n1890), .B(n1891), .ZN(n1888) );
  XOR2_X1 U1915 ( .A(n1892), .B(n1893), .Z(Result_mul_28_) );
  XNOR2_X1 U1916 ( .A(n1894), .B(n1895), .ZN(n1892) );
  XOR2_X1 U1917 ( .A(n1896), .B(n1897), .Z(Result_mul_27_) );
  XNOR2_X1 U1918 ( .A(n1898), .B(n1899), .ZN(n1896) );
  XOR2_X1 U1919 ( .A(n1900), .B(n1901), .Z(Result_mul_26_) );
  XNOR2_X1 U1920 ( .A(n1902), .B(n1903), .ZN(n1900) );
  XNOR2_X1 U1921 ( .A(n1904), .B(n1905), .ZN(Result_mul_25_) );
  XOR2_X1 U1922 ( .A(n1906), .B(n1907), .Z(n1905) );
  XNOR2_X1 U1923 ( .A(n1908), .B(n1909), .ZN(Result_mul_24_) );
  XOR2_X1 U1924 ( .A(n1910), .B(n1911), .Z(n1909) );
  XNOR2_X1 U1925 ( .A(n1912), .B(n1913), .ZN(Result_mul_23_) );
  XOR2_X1 U1926 ( .A(n1914), .B(n1915), .Z(n1913) );
  XNOR2_X1 U1927 ( .A(n1916), .B(n1917), .ZN(Result_mul_22_) );
  XOR2_X1 U1928 ( .A(n1918), .B(n1919), .Z(n1917) );
  XNOR2_X1 U1929 ( .A(n1920), .B(n1921), .ZN(Result_mul_21_) );
  XOR2_X1 U1930 ( .A(n1922), .B(n1923), .Z(n1921) );
  XNOR2_X1 U1931 ( .A(n1924), .B(n1925), .ZN(Result_mul_20_) );
  XOR2_X1 U1932 ( .A(n1926), .B(n1927), .Z(n1925) );
  XOR2_X1 U1933 ( .A(n1928), .B(n1929), .Z(Result_mul_1_) );
  AND2_X1 U1934 ( .A1(n1930), .A2(n1931), .ZN(n1929) );
  OR2_X1 U1935 ( .A1(n1932), .A2(n1933), .ZN(n1931) );
  AND2_X1 U1936 ( .A1(n1934), .A2(n1935), .ZN(n1932) );
  INV_X1 U1937 ( .A(n1936), .ZN(n1930) );
  XNOR2_X1 U1938 ( .A(n1937), .B(n1938), .ZN(Result_mul_19_) );
  XOR2_X1 U1939 ( .A(n1939), .B(n1940), .Z(n1938) );
  XNOR2_X1 U1940 ( .A(n1941), .B(n1942), .ZN(Result_mul_18_) );
  XOR2_X1 U1941 ( .A(n1943), .B(n1944), .Z(n1942) );
  XNOR2_X1 U1942 ( .A(n1945), .B(n1946), .ZN(Result_mul_17_) );
  XOR2_X1 U1943 ( .A(n1947), .B(n1948), .Z(n1946) );
  XNOR2_X1 U1944 ( .A(n1949), .B(n1950), .ZN(Result_mul_16_) );
  XOR2_X1 U1945 ( .A(n1951), .B(n1952), .Z(n1950) );
  XNOR2_X1 U1946 ( .A(n1953), .B(n1954), .ZN(Result_mul_15_) );
  AND2_X1 U1947 ( .A1(n1955), .A2(n1956), .ZN(Result_mul_14_) );
  OR2_X1 U1948 ( .A1(n1957), .A2(n1958), .ZN(n1955) );
  AND2_X1 U1949 ( .A1(n1959), .A2(n1954), .ZN(n1957) );
  XNOR2_X1 U1950 ( .A(n1960), .B(n1961), .ZN(Result_mul_13_) );
  OR2_X1 U1951 ( .A1(n1962), .A2(n1963), .ZN(n1961) );
  AND2_X1 U1952 ( .A1(n1964), .A2(n1965), .ZN(n1962) );
  OR2_X1 U1953 ( .A1(n1966), .A2(n1967), .ZN(n1964) );
  XOR2_X1 U1954 ( .A(n1968), .B(n1969), .Z(Result_mul_12_) );
  AND2_X1 U1955 ( .A1(n1970), .A2(n1971), .ZN(n1969) );
  OR2_X1 U1956 ( .A1(n1972), .A2(n1973), .ZN(n1971) );
  INV_X1 U1957 ( .A(n1974), .ZN(n1970) );
  XOR2_X1 U1958 ( .A(n1975), .B(n1976), .Z(Result_mul_11_) );
  AND2_X1 U1959 ( .A1(n1977), .A2(n1978), .ZN(n1976) );
  OR2_X1 U1960 ( .A1(n1979), .A2(n1980), .ZN(n1978) );
  AND2_X1 U1961 ( .A1(n1981), .A2(n1982), .ZN(n1979) );
  INV_X1 U1962 ( .A(n1983), .ZN(n1977) );
  XOR2_X1 U1963 ( .A(n1984), .B(n1985), .Z(Result_mul_10_) );
  AND2_X1 U1964 ( .A1(n1986), .A2(n1987), .ZN(n1985) );
  OR2_X1 U1965 ( .A1(n1988), .A2(n1989), .ZN(n1987) );
  AND2_X1 U1966 ( .A1(n1990), .A2(n1991), .ZN(n1988) );
  INV_X1 U1967 ( .A(n1992), .ZN(n1986) );
  OR3_X1 U1968 ( .A1(n1936), .A2(n1993), .A3(n1994), .ZN(Result_mul_0_) );
  INV_X1 U1969 ( .A(n1995), .ZN(n1994) );
  OR2_X1 U1970 ( .A1(n1996), .A2(n1997), .ZN(n1995) );
  AND2_X1 U1971 ( .A1(n1928), .A2(n1933), .ZN(n1993) );
  AND2_X1 U1972 ( .A1(n1886), .A2(n1887), .ZN(n1928) );
  XNOR2_X1 U1973 ( .A(n1935), .B(n1998), .ZN(n1887) );
  OR2_X1 U1974 ( .A1(n1999), .A2(n2000), .ZN(n1886) );
  OR2_X1 U1975 ( .A1(n2001), .A2(n1875), .ZN(n1999) );
  AND3_X1 U1976 ( .A1(n1874), .A2(n1873), .A3(n1871), .ZN(n1875) );
  INV_X1 U1977 ( .A(n2002), .ZN(n1873) );
  AND2_X1 U1978 ( .A1(n1867), .A2(n1871), .ZN(n2001) );
  INV_X1 U1979 ( .A(n2003), .ZN(n1871) );
  OR2_X1 U1980 ( .A1(n2004), .A2(n2000), .ZN(n2003) );
  INV_X1 U1981 ( .A(n2005), .ZN(n2000) );
  OR2_X1 U1982 ( .A1(n2006), .A2(n2007), .ZN(n2005) );
  AND2_X1 U1983 ( .A1(n2006), .A2(n2007), .ZN(n2004) );
  OR2_X1 U1984 ( .A1(n2008), .A2(n2009), .ZN(n2007) );
  AND2_X1 U1985 ( .A1(n2010), .A2(n2011), .ZN(n2009) );
  AND2_X1 U1986 ( .A1(n2012), .A2(n2013), .ZN(n2008) );
  OR2_X1 U1987 ( .A1(n2011), .A2(n2010), .ZN(n2013) );
  XOR2_X1 U1988 ( .A(n2014), .B(n2015), .Z(n2006) );
  XOR2_X1 U1989 ( .A(n2016), .B(n2017), .Z(n2015) );
  AND2_X1 U1990 ( .A1(n1865), .A2(n1866), .ZN(n1867) );
  XNOR2_X1 U1991 ( .A(n1874), .B(n2002), .ZN(n1866) );
  OR2_X1 U1992 ( .A1(n2018), .A2(n2019), .ZN(n2002) );
  AND2_X1 U1993 ( .A1(n2020), .A2(n2021), .ZN(n2019) );
  AND2_X1 U1994 ( .A1(n2022), .A2(n2023), .ZN(n2018) );
  OR2_X1 U1995 ( .A1(n2021), .A2(n2020), .ZN(n2023) );
  XNOR2_X1 U1996 ( .A(n2012), .B(n2024), .ZN(n1874) );
  XOR2_X1 U1997 ( .A(n2011), .B(n2010), .Z(n2024) );
  OR2_X1 U1998 ( .A1(n2025), .A2(n1997), .ZN(n2010) );
  OR2_X1 U1999 ( .A1(n2026), .A2(n2027), .ZN(n2011) );
  AND2_X1 U2000 ( .A1(n2028), .A2(n2029), .ZN(n2027) );
  AND2_X1 U2001 ( .A1(n2030), .A2(n2031), .ZN(n2026) );
  OR2_X1 U2002 ( .A1(n2029), .A2(n2028), .ZN(n2031) );
  XOR2_X1 U2003 ( .A(n2032), .B(n2033), .Z(n2012) );
  XOR2_X1 U2004 ( .A(n2034), .B(n2035), .Z(n2033) );
  OR2_X1 U2005 ( .A1(n2036), .A2(n2037), .ZN(n1865) );
  OR2_X1 U2006 ( .A1(n2038), .A2(n1864), .ZN(n2036) );
  AND3_X1 U2007 ( .A1(n1863), .A2(n1862), .A3(n1860), .ZN(n1864) );
  INV_X1 U2008 ( .A(n2039), .ZN(n1862) );
  AND2_X1 U2009 ( .A1(n1856), .A2(n1860), .ZN(n2038) );
  INV_X1 U2010 ( .A(n2040), .ZN(n1860) );
  OR2_X1 U2011 ( .A1(n2041), .A2(n2037), .ZN(n2040) );
  INV_X1 U2012 ( .A(n2042), .ZN(n2037) );
  OR2_X1 U2013 ( .A1(n2043), .A2(n2044), .ZN(n2042) );
  AND2_X1 U2014 ( .A1(n2043), .A2(n2044), .ZN(n2041) );
  OR2_X1 U2015 ( .A1(n2045), .A2(n2046), .ZN(n2044) );
  AND2_X1 U2016 ( .A1(n2047), .A2(n2048), .ZN(n2046) );
  AND2_X1 U2017 ( .A1(n2049), .A2(n2050), .ZN(n2045) );
  OR2_X1 U2018 ( .A1(n2048), .A2(n2047), .ZN(n2050) );
  XOR2_X1 U2019 ( .A(n2022), .B(n2051), .Z(n2043) );
  XOR2_X1 U2020 ( .A(n2021), .B(n2020), .Z(n2051) );
  OR2_X1 U2021 ( .A1(n2052), .A2(n1997), .ZN(n2020) );
  OR2_X1 U2022 ( .A1(n2053), .A2(n2054), .ZN(n2021) );
  AND2_X1 U2023 ( .A1(n2055), .A2(n2056), .ZN(n2054) );
  AND2_X1 U2024 ( .A1(n2057), .A2(n2058), .ZN(n2053) );
  OR2_X1 U2025 ( .A1(n2056), .A2(n2055), .ZN(n2058) );
  XOR2_X1 U2026 ( .A(n2030), .B(n2059), .Z(n2022) );
  XOR2_X1 U2027 ( .A(n2029), .B(n2028), .Z(n2059) );
  OR2_X1 U2028 ( .A1(n2025), .A2(n2060), .ZN(n2028) );
  OR2_X1 U2029 ( .A1(n2061), .A2(n2062), .ZN(n2029) );
  AND2_X1 U2030 ( .A1(n2063), .A2(n2064), .ZN(n2062) );
  AND2_X1 U2031 ( .A1(n2065), .A2(n2066), .ZN(n2061) );
  OR2_X1 U2032 ( .A1(n2064), .A2(n2063), .ZN(n2066) );
  XNOR2_X1 U2033 ( .A(n2067), .B(n2068), .ZN(n2030) );
  XNOR2_X1 U2034 ( .A(n2069), .B(n2070), .ZN(n2067) );
  AND2_X1 U2035 ( .A1(n1854), .A2(n1855), .ZN(n1856) );
  XNOR2_X1 U2036 ( .A(n1863), .B(n2039), .ZN(n1855) );
  OR2_X1 U2037 ( .A1(n2071), .A2(n2072), .ZN(n2039) );
  AND2_X1 U2038 ( .A1(n2073), .A2(n2074), .ZN(n2072) );
  AND2_X1 U2039 ( .A1(n2075), .A2(n2076), .ZN(n2071) );
  OR2_X1 U2040 ( .A1(n2074), .A2(n2073), .ZN(n2076) );
  XNOR2_X1 U2041 ( .A(n2049), .B(n2077), .ZN(n1863) );
  XOR2_X1 U2042 ( .A(n2048), .B(n2047), .Z(n2077) );
  OR2_X1 U2043 ( .A1(n2078), .A2(n1997), .ZN(n2047) );
  OR2_X1 U2044 ( .A1(n2079), .A2(n2080), .ZN(n2048) );
  AND2_X1 U2045 ( .A1(n2081), .A2(n2082), .ZN(n2080) );
  AND2_X1 U2046 ( .A1(n2083), .A2(n2084), .ZN(n2079) );
  OR2_X1 U2047 ( .A1(n2082), .A2(n2081), .ZN(n2084) );
  XOR2_X1 U2048 ( .A(n2057), .B(n2085), .Z(n2049) );
  XOR2_X1 U2049 ( .A(n2056), .B(n2055), .Z(n2085) );
  OR2_X1 U2050 ( .A1(n2052), .A2(n2060), .ZN(n2055) );
  OR2_X1 U2051 ( .A1(n2086), .A2(n2087), .ZN(n2056) );
  AND2_X1 U2052 ( .A1(n2088), .A2(n2089), .ZN(n2087) );
  AND2_X1 U2053 ( .A1(n2090), .A2(n2091), .ZN(n2086) );
  OR2_X1 U2054 ( .A1(n2089), .A2(n2088), .ZN(n2091) );
  XOR2_X1 U2055 ( .A(n2065), .B(n2092), .Z(n2057) );
  XOR2_X1 U2056 ( .A(n2064), .B(n2063), .Z(n2092) );
  OR2_X1 U2057 ( .A1(n2025), .A2(n2093), .ZN(n2063) );
  OR2_X1 U2058 ( .A1(n2094), .A2(n2095), .ZN(n2064) );
  AND2_X1 U2059 ( .A1(n2096), .A2(n2097), .ZN(n2095) );
  AND2_X1 U2060 ( .A1(n2098), .A2(n2099), .ZN(n2094) );
  OR2_X1 U2061 ( .A1(n2096), .A2(n2097), .ZN(n2098) );
  XOR2_X1 U2062 ( .A(n2100), .B(n2101), .Z(n2065) );
  XOR2_X1 U2063 ( .A(n2102), .B(n2103), .Z(n2101) );
  OR2_X1 U2064 ( .A1(n2104), .A2(n2105), .ZN(n1854) );
  OR2_X1 U2065 ( .A1(n2106), .A2(n1853), .ZN(n2104) );
  AND3_X1 U2066 ( .A1(n1852), .A2(n1851), .A3(n1849), .ZN(n1853) );
  INV_X1 U2067 ( .A(n2107), .ZN(n1851) );
  AND2_X1 U2068 ( .A1(n1845), .A2(n1849), .ZN(n2106) );
  INV_X1 U2069 ( .A(n2108), .ZN(n1849) );
  OR2_X1 U2070 ( .A1(n2109), .A2(n2105), .ZN(n2108) );
  INV_X1 U2071 ( .A(n2110), .ZN(n2105) );
  OR2_X1 U2072 ( .A1(n2111), .A2(n2112), .ZN(n2110) );
  AND2_X1 U2073 ( .A1(n2111), .A2(n2112), .ZN(n2109) );
  OR2_X1 U2074 ( .A1(n2113), .A2(n2114), .ZN(n2112) );
  AND2_X1 U2075 ( .A1(n2115), .A2(n2116), .ZN(n2114) );
  AND2_X1 U2076 ( .A1(n2117), .A2(n2118), .ZN(n2113) );
  OR2_X1 U2077 ( .A1(n2116), .A2(n2115), .ZN(n2118) );
  XOR2_X1 U2078 ( .A(n2075), .B(n2119), .Z(n2111) );
  XOR2_X1 U2079 ( .A(n2074), .B(n2073), .Z(n2119) );
  OR2_X1 U2080 ( .A1(n2120), .A2(n1997), .ZN(n2073) );
  OR2_X1 U2081 ( .A1(n2121), .A2(n2122), .ZN(n2074) );
  AND2_X1 U2082 ( .A1(n2123), .A2(n2124), .ZN(n2122) );
  AND2_X1 U2083 ( .A1(n2125), .A2(n2126), .ZN(n2121) );
  OR2_X1 U2084 ( .A1(n2124), .A2(n2123), .ZN(n2126) );
  XOR2_X1 U2085 ( .A(n2083), .B(n2127), .Z(n2075) );
  XOR2_X1 U2086 ( .A(n2082), .B(n2081), .Z(n2127) );
  OR2_X1 U2087 ( .A1(n2078), .A2(n2060), .ZN(n2081) );
  OR2_X1 U2088 ( .A1(n2128), .A2(n2129), .ZN(n2082) );
  AND2_X1 U2089 ( .A1(n2130), .A2(n2131), .ZN(n2129) );
  AND2_X1 U2090 ( .A1(n2132), .A2(n2133), .ZN(n2128) );
  OR2_X1 U2091 ( .A1(n2131), .A2(n2130), .ZN(n2133) );
  XOR2_X1 U2092 ( .A(n2090), .B(n2134), .Z(n2083) );
  XOR2_X1 U2093 ( .A(n2089), .B(n2088), .Z(n2134) );
  OR2_X1 U2094 ( .A1(n2052), .A2(n2093), .ZN(n2088) );
  OR2_X1 U2095 ( .A1(n2135), .A2(n2136), .ZN(n2089) );
  AND2_X1 U2096 ( .A1(n2137), .A2(n2138), .ZN(n2136) );
  AND2_X1 U2097 ( .A1(n2139), .A2(n2140), .ZN(n2135) );
  OR2_X1 U2098 ( .A1(n2138), .A2(n2137), .ZN(n2140) );
  XNOR2_X1 U2099 ( .A(n2141), .B(n2096), .ZN(n2090) );
  XOR2_X1 U2100 ( .A(n2142), .B(n2143), .Z(n2096) );
  XOR2_X1 U2101 ( .A(n2144), .B(n2145), .Z(n2143) );
  XNOR2_X1 U2102 ( .A(n2099), .B(n2097), .ZN(n2141) );
  OR2_X1 U2103 ( .A1(n2146), .A2(n2147), .ZN(n2097) );
  AND2_X1 U2104 ( .A1(n2148), .A2(n2149), .ZN(n2147) );
  AND2_X1 U2105 ( .A1(n2150), .A2(n2151), .ZN(n2146) );
  OR2_X1 U2106 ( .A1(n2149), .A2(n2148), .ZN(n2151) );
  AND2_X1 U2107 ( .A1(n1843), .A2(n1844), .ZN(n1845) );
  XNOR2_X1 U2108 ( .A(n1852), .B(n2107), .ZN(n1844) );
  OR2_X1 U2109 ( .A1(n2152), .A2(n2153), .ZN(n2107) );
  AND2_X1 U2110 ( .A1(n2154), .A2(n2155), .ZN(n2153) );
  AND2_X1 U2111 ( .A1(n2156), .A2(n2157), .ZN(n2152) );
  OR2_X1 U2112 ( .A1(n2155), .A2(n2154), .ZN(n2157) );
  XNOR2_X1 U2113 ( .A(n2117), .B(n2158), .ZN(n1852) );
  XOR2_X1 U2114 ( .A(n2116), .B(n2115), .Z(n2158) );
  OR2_X1 U2115 ( .A1(n2159), .A2(n1997), .ZN(n2115) );
  OR2_X1 U2116 ( .A1(n2160), .A2(n2161), .ZN(n2116) );
  AND2_X1 U2117 ( .A1(n2162), .A2(n2163), .ZN(n2161) );
  AND2_X1 U2118 ( .A1(n2164), .A2(n2165), .ZN(n2160) );
  OR2_X1 U2119 ( .A1(n2163), .A2(n2162), .ZN(n2165) );
  XOR2_X1 U2120 ( .A(n2125), .B(n2166), .Z(n2117) );
  XOR2_X1 U2121 ( .A(n2124), .B(n2123), .Z(n2166) );
  OR2_X1 U2122 ( .A1(n2120), .A2(n2060), .ZN(n2123) );
  OR2_X1 U2123 ( .A1(n2167), .A2(n2168), .ZN(n2124) );
  AND2_X1 U2124 ( .A1(n2169), .A2(n2170), .ZN(n2168) );
  AND2_X1 U2125 ( .A1(n2171), .A2(n2172), .ZN(n2167) );
  OR2_X1 U2126 ( .A1(n2170), .A2(n2169), .ZN(n2172) );
  XOR2_X1 U2127 ( .A(n2132), .B(n2173), .Z(n2125) );
  XOR2_X1 U2128 ( .A(n2131), .B(n2130), .Z(n2173) );
  OR2_X1 U2129 ( .A1(n2078), .A2(n2093), .ZN(n2130) );
  OR2_X1 U2130 ( .A1(n2174), .A2(n2175), .ZN(n2131) );
  AND2_X1 U2131 ( .A1(n2176), .A2(n2177), .ZN(n2175) );
  AND2_X1 U2132 ( .A1(n2178), .A2(n2179), .ZN(n2174) );
  OR2_X1 U2133 ( .A1(n2177), .A2(n2176), .ZN(n2179) );
  XOR2_X1 U2134 ( .A(n2139), .B(n2180), .Z(n2132) );
  XOR2_X1 U2135 ( .A(n2138), .B(n2137), .Z(n2180) );
  OR2_X1 U2136 ( .A1(n2052), .A2(n2181), .ZN(n2137) );
  OR2_X1 U2137 ( .A1(n2182), .A2(n2183), .ZN(n2138) );
  AND2_X1 U2138 ( .A1(n2184), .A2(n2185), .ZN(n2183) );
  AND2_X1 U2139 ( .A1(n2186), .A2(n2187), .ZN(n2182) );
  OR2_X1 U2140 ( .A1(n2184), .A2(n2185), .ZN(n2186) );
  XOR2_X1 U2141 ( .A(n2150), .B(n2188), .Z(n2139) );
  XOR2_X1 U2142 ( .A(n2149), .B(n2148), .Z(n2188) );
  OR2_X1 U2143 ( .A1(n2189), .A2(n2025), .ZN(n2148) );
  OR2_X1 U2144 ( .A1(n2190), .A2(n2191), .ZN(n2149) );
  AND2_X1 U2145 ( .A1(n2192), .A2(n2193), .ZN(n2191) );
  AND2_X1 U2146 ( .A1(n2194), .A2(n2195), .ZN(n2190) );
  OR2_X1 U2147 ( .A1(n2193), .A2(n2192), .ZN(n2195) );
  XOR2_X1 U2148 ( .A(n2196), .B(n2197), .Z(n2150) );
  XOR2_X1 U2149 ( .A(n2198), .B(n2199), .Z(n2197) );
  OR2_X1 U2150 ( .A1(n2200), .A2(n2201), .ZN(n1843) );
  OR2_X1 U2151 ( .A1(n2202), .A2(n1842), .ZN(n2200) );
  AND3_X1 U2152 ( .A1(n1841), .A2(n1840), .A3(n1838), .ZN(n1842) );
  INV_X1 U2153 ( .A(n2203), .ZN(n1840) );
  AND2_X1 U2154 ( .A1(n1838), .A2(n1834), .ZN(n2202) );
  OR2_X1 U2155 ( .A1(n2204), .A2(n1992), .ZN(n1834) );
  AND3_X1 U2156 ( .A1(n1991), .A2(n1989), .A3(n1990), .ZN(n1992) );
  INV_X1 U2157 ( .A(n2205), .ZN(n1990) );
  AND2_X1 U2158 ( .A1(n1989), .A2(n1984), .ZN(n2204) );
  OR2_X1 U2159 ( .A1(n2206), .A2(n1983), .ZN(n1984) );
  AND3_X1 U2160 ( .A1(n1982), .A2(n1980), .A3(n1981), .ZN(n1983) );
  INV_X1 U2161 ( .A(n2207), .ZN(n1981) );
  AND2_X1 U2162 ( .A1(n1980), .A2(n1975), .ZN(n2206) );
  OR2_X1 U2163 ( .A1(n2208), .A2(n1974), .ZN(n1975) );
  AND2_X1 U2164 ( .A1(n1973), .A2(n1972), .ZN(n1974) );
  AND2_X1 U2165 ( .A1(n1973), .A2(n1968), .ZN(n2208) );
  OR2_X1 U2166 ( .A1(n2209), .A2(n1963), .ZN(n1968) );
  INV_X1 U2167 ( .A(n2210), .ZN(n1963) );
  OR3_X1 U2168 ( .A1(n1967), .A2(n1966), .A3(n1965), .ZN(n2210) );
  INV_X1 U2169 ( .A(n2211), .ZN(n2209) );
  OR2_X1 U2170 ( .A1(n1956), .A2(n1965), .ZN(n2211) );
  OR2_X1 U2171 ( .A1(n2212), .A2(n1972), .ZN(n1965) );
  INV_X1 U2172 ( .A(n2213), .ZN(n1972) );
  OR2_X1 U2173 ( .A1(n2214), .A2(n2215), .ZN(n2213) );
  AND2_X1 U2174 ( .A1(n2214), .A2(n2215), .ZN(n2212) );
  OR2_X1 U2175 ( .A1(n2216), .A2(n2217), .ZN(n2215) );
  AND2_X1 U2176 ( .A1(n2218), .A2(n2219), .ZN(n2217) );
  AND2_X1 U2177 ( .A1(n2220), .A2(n2221), .ZN(n2216) );
  OR2_X1 U2178 ( .A1(n2219), .A2(n2218), .ZN(n2221) );
  XOR2_X1 U2179 ( .A(n2222), .B(n2223), .Z(n2214) );
  XOR2_X1 U2180 ( .A(n2224), .B(n2225), .Z(n2223) );
  INV_X1 U2181 ( .A(n1960), .ZN(n1956) );
  AND3_X1 U2182 ( .A1(n1954), .A2(n1958), .A3(n1959), .ZN(n1960) );
  INV_X1 U2183 ( .A(n1953), .ZN(n1959) );
  OR2_X1 U2184 ( .A1(n2226), .A2(n2227), .ZN(n1953) );
  AND2_X1 U2185 ( .A1(n1952), .A2(n1951), .ZN(n2227) );
  AND2_X1 U2186 ( .A1(n1949), .A2(n2228), .ZN(n2226) );
  OR2_X1 U2187 ( .A1(n1952), .A2(n1951), .ZN(n2228) );
  OR2_X1 U2188 ( .A1(n2229), .A2(n2230), .ZN(n1951) );
  AND2_X1 U2189 ( .A1(n1948), .A2(n1947), .ZN(n2230) );
  AND2_X1 U2190 ( .A1(n1945), .A2(n2231), .ZN(n2229) );
  OR2_X1 U2191 ( .A1(n1948), .A2(n1947), .ZN(n2231) );
  OR2_X1 U2192 ( .A1(n2232), .A2(n2233), .ZN(n1947) );
  AND2_X1 U2193 ( .A1(n1944), .A2(n1943), .ZN(n2233) );
  AND2_X1 U2194 ( .A1(n1941), .A2(n2234), .ZN(n2232) );
  OR2_X1 U2195 ( .A1(n1944), .A2(n1943), .ZN(n2234) );
  OR2_X1 U2196 ( .A1(n2235), .A2(n2236), .ZN(n1943) );
  AND2_X1 U2197 ( .A1(n1940), .A2(n1939), .ZN(n2236) );
  AND2_X1 U2198 ( .A1(n1937), .A2(n2237), .ZN(n2235) );
  OR2_X1 U2199 ( .A1(n1940), .A2(n1939), .ZN(n2237) );
  OR2_X1 U2200 ( .A1(n2238), .A2(n2239), .ZN(n1939) );
  AND2_X1 U2201 ( .A1(n1927), .A2(n1926), .ZN(n2239) );
  AND2_X1 U2202 ( .A1(n1924), .A2(n2240), .ZN(n2238) );
  OR2_X1 U2203 ( .A1(n1927), .A2(n1926), .ZN(n2240) );
  OR2_X1 U2204 ( .A1(n2241), .A2(n2242), .ZN(n1926) );
  AND2_X1 U2205 ( .A1(n1923), .A2(n1922), .ZN(n2242) );
  AND2_X1 U2206 ( .A1(n1920), .A2(n2243), .ZN(n2241) );
  OR2_X1 U2207 ( .A1(n1923), .A2(n1922), .ZN(n2243) );
  OR2_X1 U2208 ( .A1(n2244), .A2(n2245), .ZN(n1922) );
  AND2_X1 U2209 ( .A1(n1919), .A2(n1918), .ZN(n2245) );
  AND2_X1 U2210 ( .A1(n1916), .A2(n2246), .ZN(n2244) );
  OR2_X1 U2211 ( .A1(n1919), .A2(n1918), .ZN(n2246) );
  OR2_X1 U2212 ( .A1(n2247), .A2(n2248), .ZN(n1918) );
  AND2_X1 U2213 ( .A1(n1915), .A2(n1914), .ZN(n2248) );
  AND2_X1 U2214 ( .A1(n1912), .A2(n2249), .ZN(n2247) );
  OR2_X1 U2215 ( .A1(n1915), .A2(n1914), .ZN(n2249) );
  OR2_X1 U2216 ( .A1(n2250), .A2(n2251), .ZN(n1914) );
  AND2_X1 U2217 ( .A1(n1911), .A2(n1910), .ZN(n2251) );
  AND2_X1 U2218 ( .A1(n1908), .A2(n2252), .ZN(n2250) );
  OR2_X1 U2219 ( .A1(n1911), .A2(n1910), .ZN(n2252) );
  OR2_X1 U2220 ( .A1(n2253), .A2(n2254), .ZN(n1910) );
  AND2_X1 U2221 ( .A1(n1907), .A2(n1906), .ZN(n2254) );
  AND2_X1 U2222 ( .A1(n1904), .A2(n2255), .ZN(n2253) );
  OR2_X1 U2223 ( .A1(n1907), .A2(n1906), .ZN(n2255) );
  OR2_X1 U2224 ( .A1(n2256), .A2(n2257), .ZN(n1906) );
  AND2_X1 U2225 ( .A1(n1903), .A2(n1902), .ZN(n2257) );
  AND2_X1 U2226 ( .A1(n1901), .A2(n2258), .ZN(n2256) );
  OR2_X1 U2227 ( .A1(n1903), .A2(n1902), .ZN(n2258) );
  OR2_X1 U2228 ( .A1(n2259), .A2(n2260), .ZN(n1902) );
  AND2_X1 U2229 ( .A1(n1899), .A2(n1898), .ZN(n2260) );
  AND2_X1 U2230 ( .A1(n1897), .A2(n2261), .ZN(n2259) );
  OR2_X1 U2231 ( .A1(n1899), .A2(n1898), .ZN(n2261) );
  OR2_X1 U2232 ( .A1(n2262), .A2(n2263), .ZN(n1898) );
  AND2_X1 U2233 ( .A1(n1895), .A2(n1894), .ZN(n2263) );
  AND2_X1 U2234 ( .A1(n1893), .A2(n2264), .ZN(n2262) );
  OR2_X1 U2235 ( .A1(n1895), .A2(n1894), .ZN(n2264) );
  OR2_X1 U2236 ( .A1(n2265), .A2(n2266), .ZN(n1894) );
  AND2_X1 U2237 ( .A1(n1889), .A2(n2267), .ZN(n2266) );
  AND2_X1 U2238 ( .A1(n1891), .A2(n2268), .ZN(n2265) );
  OR2_X1 U2239 ( .A1(n1889), .A2(n2267), .ZN(n2268) );
  INV_X1 U2240 ( .A(n1890), .ZN(n2267) );
  OR2_X1 U2241 ( .A1(n1885), .A2(n2269), .ZN(n1889) );
  INV_X1 U2242 ( .A(n2270), .ZN(n1891) );
  OR3_X1 U2243 ( .A1(n2271), .A2(n2272), .A3(n2273), .ZN(n2270) );
  AND2_X1 U2244 ( .A1(b_14_), .A2(n1880), .ZN(n2273) );
  AND2_X1 U2245 ( .A1(b_13_), .A2(n2274), .ZN(n2272) );
  OR2_X1 U2246 ( .A1(n2275), .A2(n1884), .ZN(n2274) );
  AND2_X1 U2247 ( .A1(a_15_), .A2(n1881), .ZN(n2275) );
  AND2_X1 U2248 ( .A1(n2276), .A2(n2277), .ZN(n2271) );
  OR2_X1 U2249 ( .A1(n1885), .A2(n2278), .ZN(n1895) );
  XNOR2_X1 U2250 ( .A(n2279), .B(n2280), .ZN(n1893) );
  XNOR2_X1 U2251 ( .A(n2281), .B(n2282), .ZN(n2280) );
  OR2_X1 U2252 ( .A1(n1885), .A2(n2283), .ZN(n1899) );
  XOR2_X1 U2253 ( .A(n2284), .B(n2285), .Z(n1897) );
  XOR2_X1 U2254 ( .A(n2286), .B(n2287), .Z(n2285) );
  OR2_X1 U2255 ( .A1(n1885), .A2(n2288), .ZN(n1903) );
  XOR2_X1 U2256 ( .A(n2289), .B(n2290), .Z(n1901) );
  XOR2_X1 U2257 ( .A(n2291), .B(n2292), .Z(n2290) );
  OR2_X1 U2258 ( .A1(n1885), .A2(n2293), .ZN(n1907) );
  XOR2_X1 U2259 ( .A(n2294), .B(n2295), .Z(n1904) );
  XOR2_X1 U2260 ( .A(n2296), .B(n2297), .Z(n2295) );
  OR2_X1 U2261 ( .A1(n1885), .A2(n2298), .ZN(n1911) );
  XOR2_X1 U2262 ( .A(n2299), .B(n2300), .Z(n1908) );
  XOR2_X1 U2263 ( .A(n2301), .B(n2302), .Z(n2300) );
  OR2_X1 U2264 ( .A1(n1885), .A2(n2303), .ZN(n1915) );
  XOR2_X1 U2265 ( .A(n2304), .B(n2305), .Z(n1912) );
  XOR2_X1 U2266 ( .A(n2306), .B(n2307), .Z(n2305) );
  OR2_X1 U2267 ( .A1(n1885), .A2(n2308), .ZN(n1919) );
  XOR2_X1 U2268 ( .A(n2309), .B(n2310), .Z(n1916) );
  XOR2_X1 U2269 ( .A(n2311), .B(n2312), .Z(n2310) );
  OR2_X1 U2270 ( .A1(n1885), .A2(n2313), .ZN(n1923) );
  XOR2_X1 U2271 ( .A(n2314), .B(n2315), .Z(n1920) );
  XOR2_X1 U2272 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR2_X1 U2273 ( .A1(n1885), .A2(n2189), .ZN(n1927) );
  XOR2_X1 U2274 ( .A(n2318), .B(n2319), .Z(n1924) );
  XOR2_X1 U2275 ( .A(n2320), .B(n2321), .Z(n2319) );
  OR2_X1 U2276 ( .A1(n1885), .A2(n2181), .ZN(n1940) );
  XOR2_X1 U2277 ( .A(n2322), .B(n2323), .Z(n1937) );
  XOR2_X1 U2278 ( .A(n2324), .B(n2325), .Z(n2323) );
  OR2_X1 U2279 ( .A1(n1885), .A2(n2093), .ZN(n1944) );
  XOR2_X1 U2280 ( .A(n2326), .B(n2327), .Z(n1941) );
  XOR2_X1 U2281 ( .A(n2328), .B(n2329), .Z(n2327) );
  OR2_X1 U2282 ( .A1(n1885), .A2(n2060), .ZN(n1948) );
  XOR2_X1 U2283 ( .A(n2330), .B(n2331), .Z(n1945) );
  XOR2_X1 U2284 ( .A(n2332), .B(n2333), .Z(n2331) );
  OR2_X1 U2285 ( .A1(n1885), .A2(n1997), .ZN(n1952) );
  INV_X1 U2286 ( .A(b_15_), .ZN(n1885) );
  XOR2_X1 U2287 ( .A(n2334), .B(n2335), .Z(n1949) );
  XOR2_X1 U2288 ( .A(n2336), .B(n2337), .Z(n2335) );
  XOR2_X1 U2289 ( .A(n1966), .B(n1967), .Z(n1958) );
  OR2_X1 U2290 ( .A1(n2338), .A2(n2339), .ZN(n1967) );
  AND2_X1 U2291 ( .A1(n2340), .A2(n2341), .ZN(n2339) );
  AND2_X1 U2292 ( .A1(n2342), .A2(n2343), .ZN(n2338) );
  OR2_X1 U2293 ( .A1(n2340), .A2(n2341), .ZN(n2343) );
  XOR2_X1 U2294 ( .A(n2220), .B(n2344), .Z(n1966) );
  XOR2_X1 U2295 ( .A(n2219), .B(n2218), .Z(n2344) );
  OR2_X1 U2296 ( .A1(n2277), .A2(n1997), .ZN(n2218) );
  OR2_X1 U2297 ( .A1(n2345), .A2(n2346), .ZN(n2219) );
  AND2_X1 U2298 ( .A1(n2347), .A2(n2348), .ZN(n2346) );
  AND2_X1 U2299 ( .A1(n2349), .A2(n2350), .ZN(n2345) );
  OR2_X1 U2300 ( .A1(n2348), .A2(n2347), .ZN(n2350) );
  XOR2_X1 U2301 ( .A(n2351), .B(n2352), .Z(n2220) );
  XOR2_X1 U2302 ( .A(n2353), .B(n2354), .Z(n2352) );
  XNOR2_X1 U2303 ( .A(n2342), .B(n2355), .ZN(n1954) );
  XOR2_X1 U2304 ( .A(n2341), .B(n2340), .Z(n2355) );
  OR2_X1 U2305 ( .A1(n1881), .A2(n1997), .ZN(n2340) );
  OR2_X1 U2306 ( .A1(n2356), .A2(n2357), .ZN(n2341) );
  AND2_X1 U2307 ( .A1(n2337), .A2(n2336), .ZN(n2357) );
  AND2_X1 U2308 ( .A1(n2334), .A2(n2358), .ZN(n2356) );
  OR2_X1 U2309 ( .A1(n2336), .A2(n2337), .ZN(n2358) );
  OR2_X1 U2310 ( .A1(n1881), .A2(n2060), .ZN(n2337) );
  OR2_X1 U2311 ( .A1(n2359), .A2(n2360), .ZN(n2336) );
  AND2_X1 U2312 ( .A1(n2333), .A2(n2332), .ZN(n2360) );
  AND2_X1 U2313 ( .A1(n2330), .A2(n2361), .ZN(n2359) );
  OR2_X1 U2314 ( .A1(n2332), .A2(n2333), .ZN(n2361) );
  OR2_X1 U2315 ( .A1(n1881), .A2(n2093), .ZN(n2333) );
  OR2_X1 U2316 ( .A1(n2362), .A2(n2363), .ZN(n2332) );
  AND2_X1 U2317 ( .A1(n2329), .A2(n2328), .ZN(n2363) );
  AND2_X1 U2318 ( .A1(n2326), .A2(n2364), .ZN(n2362) );
  OR2_X1 U2319 ( .A1(n2328), .A2(n2329), .ZN(n2364) );
  OR2_X1 U2320 ( .A1(n1881), .A2(n2181), .ZN(n2329) );
  OR2_X1 U2321 ( .A1(n2365), .A2(n2366), .ZN(n2328) );
  AND2_X1 U2322 ( .A1(n2325), .A2(n2324), .ZN(n2366) );
  AND2_X1 U2323 ( .A1(n2322), .A2(n2367), .ZN(n2365) );
  OR2_X1 U2324 ( .A1(n2324), .A2(n2325), .ZN(n2367) );
  OR2_X1 U2325 ( .A1(n1881), .A2(n2189), .ZN(n2325) );
  OR2_X1 U2326 ( .A1(n2368), .A2(n2369), .ZN(n2324) );
  AND2_X1 U2327 ( .A1(n2321), .A2(n2320), .ZN(n2369) );
  AND2_X1 U2328 ( .A1(n2318), .A2(n2370), .ZN(n2368) );
  OR2_X1 U2329 ( .A1(n2320), .A2(n2321), .ZN(n2370) );
  OR2_X1 U2330 ( .A1(n1881), .A2(n2313), .ZN(n2321) );
  OR2_X1 U2331 ( .A1(n2371), .A2(n2372), .ZN(n2320) );
  AND2_X1 U2332 ( .A1(n2317), .A2(n2316), .ZN(n2372) );
  AND2_X1 U2333 ( .A1(n2314), .A2(n2373), .ZN(n2371) );
  OR2_X1 U2334 ( .A1(n2316), .A2(n2317), .ZN(n2373) );
  OR2_X1 U2335 ( .A1(n1881), .A2(n2308), .ZN(n2317) );
  OR2_X1 U2336 ( .A1(n2374), .A2(n2375), .ZN(n2316) );
  AND2_X1 U2337 ( .A1(n2312), .A2(n2311), .ZN(n2375) );
  AND2_X1 U2338 ( .A1(n2309), .A2(n2376), .ZN(n2374) );
  OR2_X1 U2339 ( .A1(n2311), .A2(n2312), .ZN(n2376) );
  OR2_X1 U2340 ( .A1(n1881), .A2(n2303), .ZN(n2312) );
  OR2_X1 U2341 ( .A1(n2377), .A2(n2378), .ZN(n2311) );
  AND2_X1 U2342 ( .A1(n2307), .A2(n2306), .ZN(n2378) );
  AND2_X1 U2343 ( .A1(n2304), .A2(n2379), .ZN(n2377) );
  OR2_X1 U2344 ( .A1(n2306), .A2(n2307), .ZN(n2379) );
  OR2_X1 U2345 ( .A1(n1881), .A2(n2298), .ZN(n2307) );
  OR2_X1 U2346 ( .A1(n2380), .A2(n2381), .ZN(n2306) );
  AND2_X1 U2347 ( .A1(n2302), .A2(n2301), .ZN(n2381) );
  AND2_X1 U2348 ( .A1(n2299), .A2(n2382), .ZN(n2380) );
  OR2_X1 U2349 ( .A1(n2301), .A2(n2302), .ZN(n2382) );
  OR2_X1 U2350 ( .A1(n1881), .A2(n2293), .ZN(n2302) );
  OR2_X1 U2351 ( .A1(n2383), .A2(n2384), .ZN(n2301) );
  AND2_X1 U2352 ( .A1(n2297), .A2(n2296), .ZN(n2384) );
  AND2_X1 U2353 ( .A1(n2294), .A2(n2385), .ZN(n2383) );
  OR2_X1 U2354 ( .A1(n2296), .A2(n2297), .ZN(n2385) );
  OR2_X1 U2355 ( .A1(n1881), .A2(n2288), .ZN(n2297) );
  OR2_X1 U2356 ( .A1(n2386), .A2(n2387), .ZN(n2296) );
  AND2_X1 U2357 ( .A1(n2292), .A2(n2291), .ZN(n2387) );
  AND2_X1 U2358 ( .A1(n2289), .A2(n2388), .ZN(n2386) );
  OR2_X1 U2359 ( .A1(n2291), .A2(n2292), .ZN(n2388) );
  OR2_X1 U2360 ( .A1(n1881), .A2(n2283), .ZN(n2292) );
  OR2_X1 U2361 ( .A1(n2389), .A2(n2390), .ZN(n2291) );
  AND2_X1 U2362 ( .A1(n2287), .A2(n2286), .ZN(n2390) );
  AND2_X1 U2363 ( .A1(n2284), .A2(n2391), .ZN(n2389) );
  OR2_X1 U2364 ( .A1(n2286), .A2(n2287), .ZN(n2391) );
  OR2_X1 U2365 ( .A1(n1881), .A2(n2278), .ZN(n2287) );
  OR2_X1 U2366 ( .A1(n2392), .A2(n2393), .ZN(n2286) );
  AND2_X1 U2367 ( .A1(n2279), .A2(n2282), .ZN(n2393) );
  AND2_X1 U2368 ( .A1(n2281), .A2(n2394), .ZN(n2392) );
  OR2_X1 U2369 ( .A1(n2282), .A2(n2279), .ZN(n2394) );
  OR2_X1 U2370 ( .A1(n1881), .A2(n2269), .ZN(n2279) );
  OR3_X1 U2371 ( .A1(n1881), .A2(n2277), .A3(n2395), .ZN(n2282) );
  INV_X1 U2372 ( .A(n2396), .ZN(n2281) );
  OR2_X1 U2373 ( .A1(n2397), .A2(n2398), .ZN(n2396) );
  AND2_X1 U2374 ( .A1(b_13_), .A2(n2399), .ZN(n2398) );
  OR2_X1 U2375 ( .A1(n2400), .A2(n1880), .ZN(n2399) );
  AND2_X1 U2376 ( .A1(a_14_), .A2(n2401), .ZN(n2400) );
  AND2_X1 U2377 ( .A1(b_12_), .A2(n2402), .ZN(n2397) );
  OR2_X1 U2378 ( .A1(n2403), .A2(n1884), .ZN(n2402) );
  AND2_X1 U2379 ( .A1(a_15_), .A2(n2277), .ZN(n2403) );
  XOR2_X1 U2380 ( .A(n2404), .B(n2405), .Z(n2284) );
  XNOR2_X1 U2381 ( .A(n2406), .B(n2407), .ZN(n2404) );
  XOR2_X1 U2382 ( .A(n2408), .B(n2409), .Z(n2289) );
  XOR2_X1 U2383 ( .A(n2410), .B(n2411), .Z(n2409) );
  XOR2_X1 U2384 ( .A(n2412), .B(n2413), .Z(n2294) );
  XOR2_X1 U2385 ( .A(n2414), .B(n2415), .Z(n2413) );
  XOR2_X1 U2386 ( .A(n2416), .B(n2417), .Z(n2299) );
  XOR2_X1 U2387 ( .A(n2418), .B(n2419), .Z(n2417) );
  XOR2_X1 U2388 ( .A(n2420), .B(n2421), .Z(n2304) );
  XOR2_X1 U2389 ( .A(n2422), .B(n2423), .Z(n2421) );
  XOR2_X1 U2390 ( .A(n2424), .B(n2425), .Z(n2309) );
  XOR2_X1 U2391 ( .A(n2426), .B(n2427), .Z(n2425) );
  XOR2_X1 U2392 ( .A(n2428), .B(n2429), .Z(n2314) );
  XOR2_X1 U2393 ( .A(n2430), .B(n2431), .Z(n2429) );
  XOR2_X1 U2394 ( .A(n2432), .B(n2433), .Z(n2318) );
  XOR2_X1 U2395 ( .A(n2434), .B(n2435), .Z(n2433) );
  XOR2_X1 U2396 ( .A(n2436), .B(n2437), .Z(n2322) );
  XOR2_X1 U2397 ( .A(n2438), .B(n2439), .Z(n2437) );
  XOR2_X1 U2398 ( .A(n2440), .B(n2441), .Z(n2326) );
  XOR2_X1 U2399 ( .A(n2442), .B(n2443), .Z(n2441) );
  XOR2_X1 U2400 ( .A(n2444), .B(n2445), .Z(n2330) );
  XOR2_X1 U2401 ( .A(n2446), .B(n2447), .Z(n2445) );
  XOR2_X1 U2402 ( .A(n2448), .B(n2449), .Z(n2334) );
  XOR2_X1 U2403 ( .A(n2450), .B(n2451), .Z(n2449) );
  XOR2_X1 U2404 ( .A(n2349), .B(n2452), .Z(n2342) );
  XOR2_X1 U2405 ( .A(n2348), .B(n2347), .Z(n2452) );
  OR2_X1 U2406 ( .A1(n2277), .A2(n2060), .ZN(n2347) );
  OR2_X1 U2407 ( .A1(n2453), .A2(n2454), .ZN(n2348) );
  AND2_X1 U2408 ( .A1(n2451), .A2(n2450), .ZN(n2454) );
  AND2_X1 U2409 ( .A1(n2448), .A2(n2455), .ZN(n2453) );
  OR2_X1 U2410 ( .A1(n2450), .A2(n2451), .ZN(n2455) );
  OR2_X1 U2411 ( .A1(n2277), .A2(n2093), .ZN(n2451) );
  OR2_X1 U2412 ( .A1(n2456), .A2(n2457), .ZN(n2450) );
  AND2_X1 U2413 ( .A1(n2447), .A2(n2446), .ZN(n2457) );
  AND2_X1 U2414 ( .A1(n2444), .A2(n2458), .ZN(n2456) );
  OR2_X1 U2415 ( .A1(n2446), .A2(n2447), .ZN(n2458) );
  OR2_X1 U2416 ( .A1(n2277), .A2(n2181), .ZN(n2447) );
  OR2_X1 U2417 ( .A1(n2459), .A2(n2460), .ZN(n2446) );
  AND2_X1 U2418 ( .A1(n2443), .A2(n2442), .ZN(n2460) );
  AND2_X1 U2419 ( .A1(n2440), .A2(n2461), .ZN(n2459) );
  OR2_X1 U2420 ( .A1(n2442), .A2(n2443), .ZN(n2461) );
  OR2_X1 U2421 ( .A1(n2277), .A2(n2189), .ZN(n2443) );
  OR2_X1 U2422 ( .A1(n2462), .A2(n2463), .ZN(n2442) );
  AND2_X1 U2423 ( .A1(n2439), .A2(n2438), .ZN(n2463) );
  AND2_X1 U2424 ( .A1(n2436), .A2(n2464), .ZN(n2462) );
  OR2_X1 U2425 ( .A1(n2438), .A2(n2439), .ZN(n2464) );
  OR2_X1 U2426 ( .A1(n2277), .A2(n2313), .ZN(n2439) );
  OR2_X1 U2427 ( .A1(n2465), .A2(n2466), .ZN(n2438) );
  AND2_X1 U2428 ( .A1(n2435), .A2(n2434), .ZN(n2466) );
  AND2_X1 U2429 ( .A1(n2432), .A2(n2467), .ZN(n2465) );
  OR2_X1 U2430 ( .A1(n2434), .A2(n2435), .ZN(n2467) );
  OR2_X1 U2431 ( .A1(n2277), .A2(n2308), .ZN(n2435) );
  OR2_X1 U2432 ( .A1(n2468), .A2(n2469), .ZN(n2434) );
  AND2_X1 U2433 ( .A1(n2431), .A2(n2430), .ZN(n2469) );
  AND2_X1 U2434 ( .A1(n2428), .A2(n2470), .ZN(n2468) );
  OR2_X1 U2435 ( .A1(n2430), .A2(n2431), .ZN(n2470) );
  OR2_X1 U2436 ( .A1(n2277), .A2(n2303), .ZN(n2431) );
  OR2_X1 U2437 ( .A1(n2471), .A2(n2472), .ZN(n2430) );
  AND2_X1 U2438 ( .A1(n2427), .A2(n2426), .ZN(n2472) );
  AND2_X1 U2439 ( .A1(n2424), .A2(n2473), .ZN(n2471) );
  OR2_X1 U2440 ( .A1(n2426), .A2(n2427), .ZN(n2473) );
  OR2_X1 U2441 ( .A1(n2277), .A2(n2298), .ZN(n2427) );
  OR2_X1 U2442 ( .A1(n2474), .A2(n2475), .ZN(n2426) );
  AND2_X1 U2443 ( .A1(n2423), .A2(n2422), .ZN(n2475) );
  AND2_X1 U2444 ( .A1(n2420), .A2(n2476), .ZN(n2474) );
  OR2_X1 U2445 ( .A1(n2422), .A2(n2423), .ZN(n2476) );
  OR2_X1 U2446 ( .A1(n2277), .A2(n2293), .ZN(n2423) );
  OR2_X1 U2447 ( .A1(n2477), .A2(n2478), .ZN(n2422) );
  AND2_X1 U2448 ( .A1(n2419), .A2(n2418), .ZN(n2478) );
  AND2_X1 U2449 ( .A1(n2416), .A2(n2479), .ZN(n2477) );
  OR2_X1 U2450 ( .A1(n2418), .A2(n2419), .ZN(n2479) );
  OR2_X1 U2451 ( .A1(n2277), .A2(n2288), .ZN(n2419) );
  OR2_X1 U2452 ( .A1(n2480), .A2(n2481), .ZN(n2418) );
  AND2_X1 U2453 ( .A1(n2415), .A2(n2414), .ZN(n2481) );
  AND2_X1 U2454 ( .A1(n2412), .A2(n2482), .ZN(n2480) );
  OR2_X1 U2455 ( .A1(n2414), .A2(n2415), .ZN(n2482) );
  OR2_X1 U2456 ( .A1(n2277), .A2(n2283), .ZN(n2415) );
  OR2_X1 U2457 ( .A1(n2483), .A2(n2484), .ZN(n2414) );
  AND2_X1 U2458 ( .A1(n2411), .A2(n2410), .ZN(n2484) );
  AND2_X1 U2459 ( .A1(n2408), .A2(n2485), .ZN(n2483) );
  OR2_X1 U2460 ( .A1(n2410), .A2(n2411), .ZN(n2485) );
  OR2_X1 U2461 ( .A1(n2277), .A2(n2278), .ZN(n2411) );
  OR2_X1 U2462 ( .A1(n2486), .A2(n2487), .ZN(n2410) );
  AND2_X1 U2463 ( .A1(n2407), .A2(n2405), .ZN(n2487) );
  AND2_X1 U2464 ( .A1(n2488), .A2(n2489), .ZN(n2486) );
  OR2_X1 U2465 ( .A1(n2407), .A2(n2405), .ZN(n2488) );
  OR3_X1 U2466 ( .A1(n2277), .A2(n2401), .A3(n2395), .ZN(n2405) );
  INV_X1 U2467 ( .A(n2490), .ZN(n2407) );
  OR2_X1 U2468 ( .A1(n2491), .A2(n2492), .ZN(n2490) );
  AND2_X1 U2469 ( .A1(b_12_), .A2(n2493), .ZN(n2492) );
  OR2_X1 U2470 ( .A1(n2494), .A2(n1880), .ZN(n2493) );
  AND2_X1 U2471 ( .A1(a_14_), .A2(n2495), .ZN(n2494) );
  AND2_X1 U2472 ( .A1(b_11_), .A2(n2496), .ZN(n2491) );
  OR2_X1 U2473 ( .A1(n2497), .A2(n1884), .ZN(n2496) );
  AND2_X1 U2474 ( .A1(a_15_), .A2(n2401), .ZN(n2497) );
  XNOR2_X1 U2475 ( .A(n2498), .B(n2499), .ZN(n2408) );
  XNOR2_X1 U2476 ( .A(n2500), .B(n2501), .ZN(n2499) );
  XNOR2_X1 U2477 ( .A(n2502), .B(n2503), .ZN(n2412) );
  XNOR2_X1 U2478 ( .A(n2504), .B(n2505), .ZN(n2502) );
  XOR2_X1 U2479 ( .A(n2506), .B(n2507), .Z(n2416) );
  XOR2_X1 U2480 ( .A(n2508), .B(n2509), .Z(n2507) );
  XOR2_X1 U2481 ( .A(n2510), .B(n2511), .Z(n2420) );
  XOR2_X1 U2482 ( .A(n2512), .B(n2513), .Z(n2511) );
  XOR2_X1 U2483 ( .A(n2514), .B(n2515), .Z(n2424) );
  XOR2_X1 U2484 ( .A(n2516), .B(n2517), .Z(n2515) );
  XOR2_X1 U2485 ( .A(n2518), .B(n2519), .Z(n2428) );
  XOR2_X1 U2486 ( .A(n2520), .B(n2521), .Z(n2519) );
  XOR2_X1 U2487 ( .A(n2522), .B(n2523), .Z(n2432) );
  XOR2_X1 U2488 ( .A(n2524), .B(n2525), .Z(n2523) );
  XOR2_X1 U2489 ( .A(n2526), .B(n2527), .Z(n2436) );
  XOR2_X1 U2490 ( .A(n2528), .B(n2529), .Z(n2527) );
  XOR2_X1 U2491 ( .A(n2530), .B(n2531), .Z(n2440) );
  XOR2_X1 U2492 ( .A(n2532), .B(n2533), .Z(n2531) );
  XOR2_X1 U2493 ( .A(n2534), .B(n2535), .Z(n2444) );
  XOR2_X1 U2494 ( .A(n2536), .B(n2537), .Z(n2535) );
  XOR2_X1 U2495 ( .A(n2538), .B(n2539), .Z(n2448) );
  XOR2_X1 U2496 ( .A(n2540), .B(n2541), .Z(n2539) );
  XOR2_X1 U2497 ( .A(n2542), .B(n2543), .Z(n2349) );
  XOR2_X1 U2498 ( .A(n2544), .B(n2545), .Z(n2543) );
  XNOR2_X1 U2499 ( .A(n1982), .B(n2207), .ZN(n1973) );
  OR2_X1 U2500 ( .A1(n2546), .A2(n2547), .ZN(n2207) );
  AND2_X1 U2501 ( .A1(n2225), .A2(n2224), .ZN(n2547) );
  AND2_X1 U2502 ( .A1(n2222), .A2(n2548), .ZN(n2546) );
  OR2_X1 U2503 ( .A1(n2224), .A2(n2225), .ZN(n2548) );
  OR2_X1 U2504 ( .A1(n2401), .A2(n1997), .ZN(n2225) );
  OR2_X1 U2505 ( .A1(n2549), .A2(n2550), .ZN(n2224) );
  AND2_X1 U2506 ( .A1(n2354), .A2(n2353), .ZN(n2550) );
  AND2_X1 U2507 ( .A1(n2351), .A2(n2551), .ZN(n2549) );
  OR2_X1 U2508 ( .A1(n2353), .A2(n2354), .ZN(n2551) );
  OR2_X1 U2509 ( .A1(n2401), .A2(n2060), .ZN(n2354) );
  OR2_X1 U2510 ( .A1(n2552), .A2(n2553), .ZN(n2353) );
  AND2_X1 U2511 ( .A1(n2545), .A2(n2544), .ZN(n2553) );
  AND2_X1 U2512 ( .A1(n2542), .A2(n2554), .ZN(n2552) );
  OR2_X1 U2513 ( .A1(n2544), .A2(n2545), .ZN(n2554) );
  OR2_X1 U2514 ( .A1(n2401), .A2(n2093), .ZN(n2545) );
  OR2_X1 U2515 ( .A1(n2555), .A2(n2556), .ZN(n2544) );
  AND2_X1 U2516 ( .A1(n2541), .A2(n2540), .ZN(n2556) );
  AND2_X1 U2517 ( .A1(n2538), .A2(n2557), .ZN(n2555) );
  OR2_X1 U2518 ( .A1(n2540), .A2(n2541), .ZN(n2557) );
  OR2_X1 U2519 ( .A1(n2401), .A2(n2181), .ZN(n2541) );
  OR2_X1 U2520 ( .A1(n2558), .A2(n2559), .ZN(n2540) );
  AND2_X1 U2521 ( .A1(n2537), .A2(n2536), .ZN(n2559) );
  AND2_X1 U2522 ( .A1(n2534), .A2(n2560), .ZN(n2558) );
  OR2_X1 U2523 ( .A1(n2536), .A2(n2537), .ZN(n2560) );
  OR2_X1 U2524 ( .A1(n2401), .A2(n2189), .ZN(n2537) );
  OR2_X1 U2525 ( .A1(n2561), .A2(n2562), .ZN(n2536) );
  AND2_X1 U2526 ( .A1(n2533), .A2(n2532), .ZN(n2562) );
  AND2_X1 U2527 ( .A1(n2530), .A2(n2563), .ZN(n2561) );
  OR2_X1 U2528 ( .A1(n2532), .A2(n2533), .ZN(n2563) );
  OR2_X1 U2529 ( .A1(n2401), .A2(n2313), .ZN(n2533) );
  OR2_X1 U2530 ( .A1(n2564), .A2(n2565), .ZN(n2532) );
  AND2_X1 U2531 ( .A1(n2529), .A2(n2528), .ZN(n2565) );
  AND2_X1 U2532 ( .A1(n2526), .A2(n2566), .ZN(n2564) );
  OR2_X1 U2533 ( .A1(n2528), .A2(n2529), .ZN(n2566) );
  OR2_X1 U2534 ( .A1(n2401), .A2(n2308), .ZN(n2529) );
  OR2_X1 U2535 ( .A1(n2567), .A2(n2568), .ZN(n2528) );
  AND2_X1 U2536 ( .A1(n2525), .A2(n2524), .ZN(n2568) );
  AND2_X1 U2537 ( .A1(n2522), .A2(n2569), .ZN(n2567) );
  OR2_X1 U2538 ( .A1(n2524), .A2(n2525), .ZN(n2569) );
  OR2_X1 U2539 ( .A1(n2401), .A2(n2303), .ZN(n2525) );
  OR2_X1 U2540 ( .A1(n2570), .A2(n2571), .ZN(n2524) );
  AND2_X1 U2541 ( .A1(n2521), .A2(n2520), .ZN(n2571) );
  AND2_X1 U2542 ( .A1(n2518), .A2(n2572), .ZN(n2570) );
  OR2_X1 U2543 ( .A1(n2520), .A2(n2521), .ZN(n2572) );
  OR2_X1 U2544 ( .A1(n2401), .A2(n2298), .ZN(n2521) );
  OR2_X1 U2545 ( .A1(n2573), .A2(n2574), .ZN(n2520) );
  AND2_X1 U2546 ( .A1(n2517), .A2(n2516), .ZN(n2574) );
  AND2_X1 U2547 ( .A1(n2514), .A2(n2575), .ZN(n2573) );
  OR2_X1 U2548 ( .A1(n2516), .A2(n2517), .ZN(n2575) );
  OR2_X1 U2549 ( .A1(n2401), .A2(n2293), .ZN(n2517) );
  OR2_X1 U2550 ( .A1(n2576), .A2(n2577), .ZN(n2516) );
  AND2_X1 U2551 ( .A1(n2513), .A2(n2512), .ZN(n2577) );
  AND2_X1 U2552 ( .A1(n2510), .A2(n2578), .ZN(n2576) );
  OR2_X1 U2553 ( .A1(n2512), .A2(n2513), .ZN(n2578) );
  OR2_X1 U2554 ( .A1(n2401), .A2(n2288), .ZN(n2513) );
  OR2_X1 U2555 ( .A1(n2579), .A2(n2580), .ZN(n2512) );
  AND2_X1 U2556 ( .A1(n2509), .A2(n2508), .ZN(n2580) );
  AND2_X1 U2557 ( .A1(n2506), .A2(n2581), .ZN(n2579) );
  OR2_X1 U2558 ( .A1(n2508), .A2(n2509), .ZN(n2581) );
  OR2_X1 U2559 ( .A1(n2401), .A2(n2283), .ZN(n2509) );
  OR2_X1 U2560 ( .A1(n2582), .A2(n2583), .ZN(n2508) );
  AND2_X1 U2561 ( .A1(n2503), .A2(n2505), .ZN(n2583) );
  AND2_X1 U2562 ( .A1(n2584), .A2(n2504), .ZN(n2582) );
  OR2_X1 U2563 ( .A1(n2505), .A2(n2503), .ZN(n2584) );
  XNOR2_X1 U2564 ( .A(n2585), .B(n2586), .ZN(n2503) );
  XNOR2_X1 U2565 ( .A(n2587), .B(n2588), .ZN(n2586) );
  OR2_X1 U2566 ( .A1(n2589), .A2(n2590), .ZN(n2505) );
  AND2_X1 U2567 ( .A1(n2498), .A2(n2501), .ZN(n2590) );
  AND2_X1 U2568 ( .A1(n2500), .A2(n2591), .ZN(n2589) );
  OR2_X1 U2569 ( .A1(n2501), .A2(n2498), .ZN(n2591) );
  OR2_X1 U2570 ( .A1(n2269), .A2(n2401), .ZN(n2498) );
  OR3_X1 U2571 ( .A1(n2401), .A2(n2395), .A3(n2495), .ZN(n2501) );
  INV_X1 U2572 ( .A(n2592), .ZN(n2500) );
  OR2_X1 U2573 ( .A1(n2593), .A2(n2594), .ZN(n2592) );
  AND2_X1 U2574 ( .A1(b_11_), .A2(n2595), .ZN(n2594) );
  OR2_X1 U2575 ( .A1(n2596), .A2(n1880), .ZN(n2595) );
  AND2_X1 U2576 ( .A1(a_14_), .A2(n2597), .ZN(n2596) );
  AND2_X1 U2577 ( .A1(b_10_), .A2(n2598), .ZN(n2593) );
  OR2_X1 U2578 ( .A1(n2599), .A2(n1884), .ZN(n2598) );
  AND2_X1 U2579 ( .A1(a_15_), .A2(n2495), .ZN(n2599) );
  XNOR2_X1 U2580 ( .A(n2600), .B(n2601), .ZN(n2506) );
  XNOR2_X1 U2581 ( .A(n2602), .B(n2603), .ZN(n2600) );
  XNOR2_X1 U2582 ( .A(n2604), .B(n2605), .ZN(n2510) );
  XNOR2_X1 U2583 ( .A(n2606), .B(n2607), .ZN(n2604) );
  XOR2_X1 U2584 ( .A(n2608), .B(n2609), .Z(n2514) );
  XOR2_X1 U2585 ( .A(n2610), .B(n2611), .Z(n2609) );
  XOR2_X1 U2586 ( .A(n2612), .B(n2613), .Z(n2518) );
  XOR2_X1 U2587 ( .A(n2614), .B(n2615), .Z(n2613) );
  XOR2_X1 U2588 ( .A(n2616), .B(n2617), .Z(n2522) );
  XOR2_X1 U2589 ( .A(n2618), .B(n2619), .Z(n2617) );
  XOR2_X1 U2590 ( .A(n2620), .B(n2621), .Z(n2526) );
  XOR2_X1 U2591 ( .A(n2622), .B(n2623), .Z(n2621) );
  XOR2_X1 U2592 ( .A(n2624), .B(n2625), .Z(n2530) );
  XOR2_X1 U2593 ( .A(n2626), .B(n2627), .Z(n2625) );
  XOR2_X1 U2594 ( .A(n2628), .B(n2629), .Z(n2534) );
  XOR2_X1 U2595 ( .A(n2630), .B(n2631), .Z(n2629) );
  XOR2_X1 U2596 ( .A(n2632), .B(n2633), .Z(n2538) );
  XOR2_X1 U2597 ( .A(n2634), .B(n2635), .Z(n2633) );
  XOR2_X1 U2598 ( .A(n2636), .B(n2637), .Z(n2542) );
  XOR2_X1 U2599 ( .A(n2638), .B(n2639), .Z(n2637) );
  XOR2_X1 U2600 ( .A(n2640), .B(n2641), .Z(n2351) );
  XOR2_X1 U2601 ( .A(n2642), .B(n2643), .Z(n2641) );
  XOR2_X1 U2602 ( .A(n2644), .B(n2645), .Z(n2222) );
  XOR2_X1 U2603 ( .A(n2646), .B(n2647), .Z(n2645) );
  XNOR2_X1 U2604 ( .A(n2648), .B(n2649), .ZN(n1982) );
  XOR2_X1 U2605 ( .A(n2650), .B(n2651), .Z(n2649) );
  XNOR2_X1 U2606 ( .A(n1991), .B(n2205), .ZN(n1980) );
  OR2_X1 U2607 ( .A1(n2652), .A2(n2653), .ZN(n2205) );
  AND2_X1 U2608 ( .A1(n2651), .A2(n2650), .ZN(n2653) );
  AND2_X1 U2609 ( .A1(n2648), .A2(n2654), .ZN(n2652) );
  OR2_X1 U2610 ( .A1(n2650), .A2(n2651), .ZN(n2654) );
  OR2_X1 U2611 ( .A1(n2495), .A2(n1997), .ZN(n2651) );
  OR2_X1 U2612 ( .A1(n2655), .A2(n2656), .ZN(n2650) );
  AND2_X1 U2613 ( .A1(n2647), .A2(n2646), .ZN(n2656) );
  AND2_X1 U2614 ( .A1(n2644), .A2(n2657), .ZN(n2655) );
  OR2_X1 U2615 ( .A1(n2646), .A2(n2647), .ZN(n2657) );
  OR2_X1 U2616 ( .A1(n2495), .A2(n2060), .ZN(n2647) );
  OR2_X1 U2617 ( .A1(n2658), .A2(n2659), .ZN(n2646) );
  AND2_X1 U2618 ( .A1(n2643), .A2(n2642), .ZN(n2659) );
  AND2_X1 U2619 ( .A1(n2640), .A2(n2660), .ZN(n2658) );
  OR2_X1 U2620 ( .A1(n2642), .A2(n2643), .ZN(n2660) );
  OR2_X1 U2621 ( .A1(n2495), .A2(n2093), .ZN(n2643) );
  OR2_X1 U2622 ( .A1(n2661), .A2(n2662), .ZN(n2642) );
  AND2_X1 U2623 ( .A1(n2639), .A2(n2638), .ZN(n2662) );
  AND2_X1 U2624 ( .A1(n2636), .A2(n2663), .ZN(n2661) );
  OR2_X1 U2625 ( .A1(n2638), .A2(n2639), .ZN(n2663) );
  OR2_X1 U2626 ( .A1(n2495), .A2(n2181), .ZN(n2639) );
  OR2_X1 U2627 ( .A1(n2664), .A2(n2665), .ZN(n2638) );
  AND2_X1 U2628 ( .A1(n2635), .A2(n2634), .ZN(n2665) );
  AND2_X1 U2629 ( .A1(n2632), .A2(n2666), .ZN(n2664) );
  OR2_X1 U2630 ( .A1(n2634), .A2(n2635), .ZN(n2666) );
  OR2_X1 U2631 ( .A1(n2495), .A2(n2189), .ZN(n2635) );
  OR2_X1 U2632 ( .A1(n2667), .A2(n2668), .ZN(n2634) );
  AND2_X1 U2633 ( .A1(n2631), .A2(n2630), .ZN(n2668) );
  AND2_X1 U2634 ( .A1(n2628), .A2(n2669), .ZN(n2667) );
  OR2_X1 U2635 ( .A1(n2630), .A2(n2631), .ZN(n2669) );
  OR2_X1 U2636 ( .A1(n2495), .A2(n2313), .ZN(n2631) );
  OR2_X1 U2637 ( .A1(n2670), .A2(n2671), .ZN(n2630) );
  AND2_X1 U2638 ( .A1(n2627), .A2(n2626), .ZN(n2671) );
  AND2_X1 U2639 ( .A1(n2624), .A2(n2672), .ZN(n2670) );
  OR2_X1 U2640 ( .A1(n2626), .A2(n2627), .ZN(n2672) );
  OR2_X1 U2641 ( .A1(n2495), .A2(n2308), .ZN(n2627) );
  OR2_X1 U2642 ( .A1(n2673), .A2(n2674), .ZN(n2626) );
  AND2_X1 U2643 ( .A1(n2623), .A2(n2622), .ZN(n2674) );
  AND2_X1 U2644 ( .A1(n2620), .A2(n2675), .ZN(n2673) );
  OR2_X1 U2645 ( .A1(n2622), .A2(n2623), .ZN(n2675) );
  OR2_X1 U2646 ( .A1(n2495), .A2(n2303), .ZN(n2623) );
  OR2_X1 U2647 ( .A1(n2676), .A2(n2677), .ZN(n2622) );
  AND2_X1 U2648 ( .A1(n2619), .A2(n2618), .ZN(n2677) );
  AND2_X1 U2649 ( .A1(n2616), .A2(n2678), .ZN(n2676) );
  OR2_X1 U2650 ( .A1(n2618), .A2(n2619), .ZN(n2678) );
  OR2_X1 U2651 ( .A1(n2495), .A2(n2298), .ZN(n2619) );
  OR2_X1 U2652 ( .A1(n2679), .A2(n2680), .ZN(n2618) );
  AND2_X1 U2653 ( .A1(n2615), .A2(n2614), .ZN(n2680) );
  AND2_X1 U2654 ( .A1(n2612), .A2(n2681), .ZN(n2679) );
  OR2_X1 U2655 ( .A1(n2614), .A2(n2615), .ZN(n2681) );
  OR2_X1 U2656 ( .A1(n2495), .A2(n2293), .ZN(n2615) );
  OR2_X1 U2657 ( .A1(n2682), .A2(n2683), .ZN(n2614) );
  AND2_X1 U2658 ( .A1(n2611), .A2(n2610), .ZN(n2683) );
  AND2_X1 U2659 ( .A1(n2608), .A2(n2684), .ZN(n2682) );
  OR2_X1 U2660 ( .A1(n2610), .A2(n2611), .ZN(n2684) );
  OR2_X1 U2661 ( .A1(n2495), .A2(n2288), .ZN(n2611) );
  OR2_X1 U2662 ( .A1(n2685), .A2(n2686), .ZN(n2610) );
  AND2_X1 U2663 ( .A1(n2605), .A2(n2607), .ZN(n2686) );
  AND2_X1 U2664 ( .A1(n2687), .A2(n2606), .ZN(n2685) );
  OR2_X1 U2665 ( .A1(n2607), .A2(n2605), .ZN(n2687) );
  XNOR2_X1 U2666 ( .A(n2688), .B(n2689), .ZN(n2605) );
  XNOR2_X1 U2667 ( .A(n2690), .B(n2691), .ZN(n2688) );
  OR2_X1 U2668 ( .A1(n2692), .A2(n2693), .ZN(n2607) );
  AND2_X1 U2669 ( .A1(n2603), .A2(n2602), .ZN(n2693) );
  AND2_X1 U2670 ( .A1(n2601), .A2(n2694), .ZN(n2692) );
  OR2_X1 U2671 ( .A1(n2602), .A2(n2603), .ZN(n2694) );
  OR2_X1 U2672 ( .A1(n2278), .A2(n2495), .ZN(n2603) );
  OR2_X1 U2673 ( .A1(n2695), .A2(n2696), .ZN(n2602) );
  AND2_X1 U2674 ( .A1(n2585), .A2(n2588), .ZN(n2696) );
  AND2_X1 U2675 ( .A1(n2587), .A2(n2697), .ZN(n2695) );
  OR2_X1 U2676 ( .A1(n2588), .A2(n2585), .ZN(n2697) );
  OR2_X1 U2677 ( .A1(n2269), .A2(n2495), .ZN(n2585) );
  OR3_X1 U2678 ( .A1(n2395), .A2(n2495), .A3(n2597), .ZN(n2588) );
  INV_X1 U2679 ( .A(n2698), .ZN(n2587) );
  OR2_X1 U2680 ( .A1(n2699), .A2(n2700), .ZN(n2698) );
  AND2_X1 U2681 ( .A1(b_9_), .A2(n2701), .ZN(n2700) );
  OR2_X1 U2682 ( .A1(n2702), .A2(n1884), .ZN(n2701) );
  AND2_X1 U2683 ( .A1(a_15_), .A2(n2597), .ZN(n2702) );
  AND2_X1 U2684 ( .A1(b_10_), .A2(n2703), .ZN(n2699) );
  OR2_X1 U2685 ( .A1(n2704), .A2(n1880), .ZN(n2703) );
  AND2_X1 U2686 ( .A1(a_14_), .A2(n2705), .ZN(n2704) );
  XNOR2_X1 U2687 ( .A(n2706), .B(n2707), .ZN(n2601) );
  XNOR2_X1 U2688 ( .A(n2708), .B(n2709), .ZN(n2707) );
  XOR2_X1 U2689 ( .A(n2710), .B(n2711), .Z(n2608) );
  XOR2_X1 U2690 ( .A(n2712), .B(n2713), .Z(n2711) );
  XNOR2_X1 U2691 ( .A(n2714), .B(n2715), .ZN(n2612) );
  XNOR2_X1 U2692 ( .A(n2716), .B(n2717), .ZN(n2714) );
  XOR2_X1 U2693 ( .A(n2718), .B(n2719), .Z(n2616) );
  XOR2_X1 U2694 ( .A(n2720), .B(n2721), .Z(n2719) );
  XOR2_X1 U2695 ( .A(n2722), .B(n2723), .Z(n2620) );
  XOR2_X1 U2696 ( .A(n2724), .B(n2725), .Z(n2723) );
  XOR2_X1 U2697 ( .A(n2726), .B(n2727), .Z(n2624) );
  XOR2_X1 U2698 ( .A(n2728), .B(n2729), .Z(n2727) );
  XOR2_X1 U2699 ( .A(n2730), .B(n2731), .Z(n2628) );
  XOR2_X1 U2700 ( .A(n2732), .B(n2733), .Z(n2731) );
  XOR2_X1 U2701 ( .A(n2734), .B(n2735), .Z(n2632) );
  XOR2_X1 U2702 ( .A(n2736), .B(n2737), .Z(n2735) );
  XOR2_X1 U2703 ( .A(n2738), .B(n2739), .Z(n2636) );
  XOR2_X1 U2704 ( .A(n2740), .B(n2741), .Z(n2739) );
  XOR2_X1 U2705 ( .A(n2742), .B(n2743), .Z(n2640) );
  XOR2_X1 U2706 ( .A(n2744), .B(n2745), .Z(n2743) );
  XOR2_X1 U2707 ( .A(n2746), .B(n2747), .Z(n2644) );
  XOR2_X1 U2708 ( .A(n2748), .B(n2749), .Z(n2747) );
  XOR2_X1 U2709 ( .A(n2750), .B(n2751), .Z(n2648) );
  XOR2_X1 U2710 ( .A(n2752), .B(n2753), .Z(n2751) );
  XNOR2_X1 U2711 ( .A(n2754), .B(n2755), .ZN(n1991) );
  XOR2_X1 U2712 ( .A(n2756), .B(n2757), .Z(n2755) );
  XNOR2_X1 U2713 ( .A(n1841), .B(n2203), .ZN(n1989) );
  OR2_X1 U2714 ( .A1(n2758), .A2(n2759), .ZN(n2203) );
  AND2_X1 U2715 ( .A1(n2757), .A2(n2756), .ZN(n2759) );
  AND2_X1 U2716 ( .A1(n2754), .A2(n2760), .ZN(n2758) );
  OR2_X1 U2717 ( .A1(n2756), .A2(n2757), .ZN(n2760) );
  OR2_X1 U2718 ( .A1(n2597), .A2(n1997), .ZN(n2757) );
  OR2_X1 U2719 ( .A1(n2761), .A2(n2762), .ZN(n2756) );
  AND2_X1 U2720 ( .A1(n2753), .A2(n2752), .ZN(n2762) );
  AND2_X1 U2721 ( .A1(n2750), .A2(n2763), .ZN(n2761) );
  OR2_X1 U2722 ( .A1(n2752), .A2(n2753), .ZN(n2763) );
  OR2_X1 U2723 ( .A1(n2597), .A2(n2060), .ZN(n2753) );
  OR2_X1 U2724 ( .A1(n2764), .A2(n2765), .ZN(n2752) );
  AND2_X1 U2725 ( .A1(n2749), .A2(n2748), .ZN(n2765) );
  AND2_X1 U2726 ( .A1(n2746), .A2(n2766), .ZN(n2764) );
  OR2_X1 U2727 ( .A1(n2748), .A2(n2749), .ZN(n2766) );
  OR2_X1 U2728 ( .A1(n2597), .A2(n2093), .ZN(n2749) );
  OR2_X1 U2729 ( .A1(n2767), .A2(n2768), .ZN(n2748) );
  AND2_X1 U2730 ( .A1(n2742), .A2(n2745), .ZN(n2768) );
  AND2_X1 U2731 ( .A1(n2769), .A2(n2744), .ZN(n2767) );
  OR2_X1 U2732 ( .A1(n2770), .A2(n2771), .ZN(n2744) );
  AND2_X1 U2733 ( .A1(n2741), .A2(n2740), .ZN(n2771) );
  AND2_X1 U2734 ( .A1(n2738), .A2(n2772), .ZN(n2770) );
  OR2_X1 U2735 ( .A1(n2740), .A2(n2741), .ZN(n2772) );
  OR2_X1 U2736 ( .A1(n2597), .A2(n2189), .ZN(n2741) );
  OR2_X1 U2737 ( .A1(n2773), .A2(n2774), .ZN(n2740) );
  AND2_X1 U2738 ( .A1(n2734), .A2(n2737), .ZN(n2774) );
  AND2_X1 U2739 ( .A1(n2775), .A2(n2736), .ZN(n2773) );
  OR2_X1 U2740 ( .A1(n2776), .A2(n2777), .ZN(n2736) );
  AND2_X1 U2741 ( .A1(n2730), .A2(n2733), .ZN(n2777) );
  AND2_X1 U2742 ( .A1(n2778), .A2(n2732), .ZN(n2776) );
  OR2_X1 U2743 ( .A1(n2779), .A2(n2780), .ZN(n2732) );
  AND2_X1 U2744 ( .A1(n2726), .A2(n2729), .ZN(n2780) );
  AND2_X1 U2745 ( .A1(n2781), .A2(n2728), .ZN(n2779) );
  OR2_X1 U2746 ( .A1(n2782), .A2(n2783), .ZN(n2728) );
  AND2_X1 U2747 ( .A1(n2722), .A2(n2725), .ZN(n2783) );
  AND2_X1 U2748 ( .A1(n2784), .A2(n2724), .ZN(n2782) );
  OR2_X1 U2749 ( .A1(n2785), .A2(n2786), .ZN(n2724) );
  AND2_X1 U2750 ( .A1(n2718), .A2(n2721), .ZN(n2786) );
  AND2_X1 U2751 ( .A1(n2787), .A2(n2720), .ZN(n2785) );
  OR2_X1 U2752 ( .A1(n2788), .A2(n2789), .ZN(n2720) );
  AND2_X1 U2753 ( .A1(n2715), .A2(n2717), .ZN(n2789) );
  AND2_X1 U2754 ( .A1(n2790), .A2(n2716), .ZN(n2788) );
  OR2_X1 U2755 ( .A1(n2717), .A2(n2715), .ZN(n2790) );
  XOR2_X1 U2756 ( .A(n2791), .B(n2792), .Z(n2715) );
  XOR2_X1 U2757 ( .A(n2793), .B(n2794), .Z(n2792) );
  OR2_X1 U2758 ( .A1(n2795), .A2(n2796), .ZN(n2717) );
  AND2_X1 U2759 ( .A1(n2710), .A2(n2713), .ZN(n2796) );
  AND2_X1 U2760 ( .A1(n2797), .A2(n2712), .ZN(n2795) );
  OR2_X1 U2761 ( .A1(n2798), .A2(n2799), .ZN(n2712) );
  AND2_X1 U2762 ( .A1(n2689), .A2(n2691), .ZN(n2799) );
  AND2_X1 U2763 ( .A1(n2800), .A2(n2690), .ZN(n2798) );
  OR2_X1 U2764 ( .A1(n2801), .A2(n2802), .ZN(n2690) );
  AND2_X1 U2765 ( .A1(n2706), .A2(n2709), .ZN(n2802) );
  AND2_X1 U2766 ( .A1(n2708), .A2(n2803), .ZN(n2801) );
  OR2_X1 U2767 ( .A1(n2709), .A2(n2706), .ZN(n2803) );
  OR2_X1 U2768 ( .A1(n2269), .A2(n2597), .ZN(n2706) );
  OR3_X1 U2769 ( .A1(n2395), .A2(n2597), .A3(n2705), .ZN(n2709) );
  INV_X1 U2770 ( .A(n2804), .ZN(n2708) );
  OR2_X1 U2771 ( .A1(n2805), .A2(n2806), .ZN(n2804) );
  AND2_X1 U2772 ( .A1(b_9_), .A2(n2807), .ZN(n2806) );
  OR2_X1 U2773 ( .A1(n2808), .A2(n1880), .ZN(n2807) );
  AND2_X1 U2774 ( .A1(a_14_), .A2(n2809), .ZN(n2808) );
  AND2_X1 U2775 ( .A1(b_8_), .A2(n2810), .ZN(n2805) );
  OR2_X1 U2776 ( .A1(n2811), .A2(n1884), .ZN(n2810) );
  AND2_X1 U2777 ( .A1(a_15_), .A2(n2705), .ZN(n2811) );
  OR2_X1 U2778 ( .A1(n2691), .A2(n2689), .ZN(n2800) );
  XNOR2_X1 U2779 ( .A(n2812), .B(n2813), .ZN(n2689) );
  XNOR2_X1 U2780 ( .A(n2814), .B(n2815), .ZN(n2813) );
  OR2_X1 U2781 ( .A1(n2278), .A2(n2597), .ZN(n2691) );
  OR2_X1 U2782 ( .A1(n2713), .A2(n2710), .ZN(n2797) );
  XNOR2_X1 U2783 ( .A(n2816), .B(n2817), .ZN(n2710) );
  XNOR2_X1 U2784 ( .A(n2818), .B(n2819), .ZN(n2816) );
  OR2_X1 U2785 ( .A1(n2283), .A2(n2597), .ZN(n2713) );
  OR2_X1 U2786 ( .A1(n2721), .A2(n2718), .ZN(n2787) );
  XOR2_X1 U2787 ( .A(n2820), .B(n2821), .Z(n2718) );
  XOR2_X1 U2788 ( .A(n2822), .B(n2823), .Z(n2821) );
  OR2_X1 U2789 ( .A1(n2597), .A2(n2293), .ZN(n2721) );
  OR2_X1 U2790 ( .A1(n2725), .A2(n2722), .ZN(n2784) );
  XNOR2_X1 U2791 ( .A(n2824), .B(n2825), .ZN(n2722) );
  XNOR2_X1 U2792 ( .A(n2826), .B(n2827), .ZN(n2824) );
  OR2_X1 U2793 ( .A1(n2597), .A2(n2298), .ZN(n2725) );
  OR2_X1 U2794 ( .A1(n2729), .A2(n2726), .ZN(n2781) );
  XOR2_X1 U2795 ( .A(n2828), .B(n2829), .Z(n2726) );
  XOR2_X1 U2796 ( .A(n2830), .B(n2831), .Z(n2829) );
  OR2_X1 U2797 ( .A1(n2597), .A2(n2303), .ZN(n2729) );
  OR2_X1 U2798 ( .A1(n2733), .A2(n2730), .ZN(n2778) );
  XOR2_X1 U2799 ( .A(n2832), .B(n2833), .Z(n2730) );
  XOR2_X1 U2800 ( .A(n2834), .B(n2835), .Z(n2833) );
  OR2_X1 U2801 ( .A1(n2597), .A2(n2308), .ZN(n2733) );
  OR2_X1 U2802 ( .A1(n2737), .A2(n2734), .ZN(n2775) );
  XOR2_X1 U2803 ( .A(n2836), .B(n2837), .Z(n2734) );
  XOR2_X1 U2804 ( .A(n2838), .B(n2839), .Z(n2837) );
  OR2_X1 U2805 ( .A1(n2597), .A2(n2313), .ZN(n2737) );
  XOR2_X1 U2806 ( .A(n2840), .B(n2841), .Z(n2738) );
  XOR2_X1 U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  OR2_X1 U2808 ( .A1(n2745), .A2(n2742), .ZN(n2769) );
  XOR2_X1 U2809 ( .A(n2844), .B(n2845), .Z(n2742) );
  XOR2_X1 U2810 ( .A(n2846), .B(n2847), .Z(n2845) );
  OR2_X1 U2811 ( .A1(n2597), .A2(n2181), .ZN(n2745) );
  XOR2_X1 U2812 ( .A(n2848), .B(n2849), .Z(n2746) );
  XOR2_X1 U2813 ( .A(n2850), .B(n2851), .Z(n2849) );
  XOR2_X1 U2814 ( .A(n2852), .B(n2853), .Z(n2750) );
  XOR2_X1 U2815 ( .A(n2854), .B(n2855), .Z(n2853) );
  XOR2_X1 U2816 ( .A(n2856), .B(n2857), .Z(n2754) );
  XOR2_X1 U2817 ( .A(n2858), .B(n2859), .Z(n2857) );
  XNOR2_X1 U2818 ( .A(n2860), .B(n2861), .ZN(n1841) );
  XOR2_X1 U2819 ( .A(n2862), .B(n2863), .Z(n2861) );
  INV_X1 U2820 ( .A(n2864), .ZN(n1838) );
  OR2_X1 U2821 ( .A1(n2865), .A2(n2201), .ZN(n2864) );
  INV_X1 U2822 ( .A(n2866), .ZN(n2201) );
  OR2_X1 U2823 ( .A1(n2867), .A2(n2868), .ZN(n2866) );
  AND2_X1 U2824 ( .A1(n2867), .A2(n2868), .ZN(n2865) );
  OR2_X1 U2825 ( .A1(n2869), .A2(n2870), .ZN(n2868) );
  AND2_X1 U2826 ( .A1(n2863), .A2(n2862), .ZN(n2870) );
  AND2_X1 U2827 ( .A1(n2860), .A2(n2871), .ZN(n2869) );
  OR2_X1 U2828 ( .A1(n2862), .A2(n2863), .ZN(n2871) );
  OR2_X1 U2829 ( .A1(n2705), .A2(n1997), .ZN(n2863) );
  OR2_X1 U2830 ( .A1(n2872), .A2(n2873), .ZN(n2862) );
  AND2_X1 U2831 ( .A1(n2859), .A2(n2858), .ZN(n2873) );
  AND2_X1 U2832 ( .A1(n2856), .A2(n2874), .ZN(n2872) );
  OR2_X1 U2833 ( .A1(n2858), .A2(n2859), .ZN(n2874) );
  OR2_X1 U2834 ( .A1(n2705), .A2(n2060), .ZN(n2859) );
  OR2_X1 U2835 ( .A1(n2875), .A2(n2876), .ZN(n2858) );
  AND2_X1 U2836 ( .A1(n2855), .A2(n2854), .ZN(n2876) );
  AND2_X1 U2837 ( .A1(n2852), .A2(n2877), .ZN(n2875) );
  OR2_X1 U2838 ( .A1(n2854), .A2(n2855), .ZN(n2877) );
  OR2_X1 U2839 ( .A1(n2705), .A2(n2093), .ZN(n2855) );
  OR2_X1 U2840 ( .A1(n2878), .A2(n2879), .ZN(n2854) );
  AND2_X1 U2841 ( .A1(n2851), .A2(n2850), .ZN(n2879) );
  AND2_X1 U2842 ( .A1(n2848), .A2(n2880), .ZN(n2878) );
  OR2_X1 U2843 ( .A1(n2850), .A2(n2851), .ZN(n2880) );
  OR2_X1 U2844 ( .A1(n2705), .A2(n2181), .ZN(n2851) );
  OR2_X1 U2845 ( .A1(n2881), .A2(n2882), .ZN(n2850) );
  AND2_X1 U2846 ( .A1(n2844), .A2(n2847), .ZN(n2882) );
  AND2_X1 U2847 ( .A1(n2883), .A2(n2846), .ZN(n2881) );
  OR2_X1 U2848 ( .A1(n2884), .A2(n2885), .ZN(n2846) );
  AND2_X1 U2849 ( .A1(n2843), .A2(n2842), .ZN(n2885) );
  AND2_X1 U2850 ( .A1(n2840), .A2(n2886), .ZN(n2884) );
  OR2_X1 U2851 ( .A1(n2842), .A2(n2843), .ZN(n2886) );
  OR2_X1 U2852 ( .A1(n2705), .A2(n2313), .ZN(n2843) );
  OR2_X1 U2853 ( .A1(n2887), .A2(n2888), .ZN(n2842) );
  AND2_X1 U2854 ( .A1(n2836), .A2(n2839), .ZN(n2888) );
  AND2_X1 U2855 ( .A1(n2889), .A2(n2838), .ZN(n2887) );
  OR2_X1 U2856 ( .A1(n2890), .A2(n2891), .ZN(n2838) );
  AND2_X1 U2857 ( .A1(n2832), .A2(n2835), .ZN(n2891) );
  AND2_X1 U2858 ( .A1(n2892), .A2(n2834), .ZN(n2890) );
  OR2_X1 U2859 ( .A1(n2893), .A2(n2894), .ZN(n2834) );
  AND2_X1 U2860 ( .A1(n2828), .A2(n2831), .ZN(n2894) );
  AND2_X1 U2861 ( .A1(n2895), .A2(n2830), .ZN(n2893) );
  OR2_X1 U2862 ( .A1(n2896), .A2(n2897), .ZN(n2830) );
  AND2_X1 U2863 ( .A1(n2825), .A2(n2827), .ZN(n2897) );
  AND2_X1 U2864 ( .A1(n2898), .A2(n2826), .ZN(n2896) );
  OR2_X1 U2865 ( .A1(n2827), .A2(n2825), .ZN(n2898) );
  XOR2_X1 U2866 ( .A(n2899), .B(n2900), .Z(n2825) );
  XOR2_X1 U2867 ( .A(n2901), .B(n2902), .Z(n2900) );
  OR2_X1 U2868 ( .A1(n2903), .A2(n2904), .ZN(n2827) );
  AND2_X1 U2869 ( .A1(n2820), .A2(n2823), .ZN(n2904) );
  AND2_X1 U2870 ( .A1(n2905), .A2(n2822), .ZN(n2903) );
  OR2_X1 U2871 ( .A1(n2906), .A2(n2907), .ZN(n2822) );
  AND2_X1 U2872 ( .A1(n2791), .A2(n2794), .ZN(n2907) );
  AND2_X1 U2873 ( .A1(n2908), .A2(n2793), .ZN(n2906) );
  OR2_X1 U2874 ( .A1(n2909), .A2(n2910), .ZN(n2793) );
  AND2_X1 U2875 ( .A1(n2817), .A2(n2819), .ZN(n2910) );
  AND2_X1 U2876 ( .A1(n2911), .A2(n2818), .ZN(n2909) );
  OR2_X1 U2877 ( .A1(n2912), .A2(n2913), .ZN(n2818) );
  AND2_X1 U2878 ( .A1(n2812), .A2(n2815), .ZN(n2913) );
  AND2_X1 U2879 ( .A1(n2814), .A2(n2914), .ZN(n2912) );
  OR2_X1 U2880 ( .A1(n2815), .A2(n2812), .ZN(n2914) );
  OR2_X1 U2881 ( .A1(n2269), .A2(n2705), .ZN(n2812) );
  OR3_X1 U2882 ( .A1(n2395), .A2(n2705), .A3(n2809), .ZN(n2815) );
  INV_X1 U2883 ( .A(n2915), .ZN(n2814) );
  OR2_X1 U2884 ( .A1(n2916), .A2(n2917), .ZN(n2915) );
  AND2_X1 U2885 ( .A1(b_8_), .A2(n2918), .ZN(n2917) );
  OR2_X1 U2886 ( .A1(n2919), .A2(n1880), .ZN(n2918) );
  AND2_X1 U2887 ( .A1(a_14_), .A2(n2159), .ZN(n2919) );
  AND2_X1 U2888 ( .A1(b_7_), .A2(n2920), .ZN(n2916) );
  OR2_X1 U2889 ( .A1(n2921), .A2(n1884), .ZN(n2920) );
  AND2_X1 U2890 ( .A1(a_15_), .A2(n2809), .ZN(n2921) );
  OR2_X1 U2891 ( .A1(n2819), .A2(n2817), .ZN(n2911) );
  XNOR2_X1 U2892 ( .A(n2922), .B(n2923), .ZN(n2817) );
  XNOR2_X1 U2893 ( .A(n2924), .B(n2925), .ZN(n2923) );
  OR2_X1 U2894 ( .A1(n2278), .A2(n2705), .ZN(n2819) );
  OR2_X1 U2895 ( .A1(n2794), .A2(n2791), .ZN(n2908) );
  XNOR2_X1 U2896 ( .A(n2926), .B(n2927), .ZN(n2791) );
  XNOR2_X1 U2897 ( .A(n2928), .B(n2929), .ZN(n2926) );
  OR2_X1 U2898 ( .A1(n2283), .A2(n2705), .ZN(n2794) );
  OR2_X1 U2899 ( .A1(n2823), .A2(n2820), .ZN(n2905) );
  XOR2_X1 U2900 ( .A(n2930), .B(n2931), .Z(n2820) );
  XOR2_X1 U2901 ( .A(n2932), .B(n2933), .Z(n2931) );
  OR2_X1 U2902 ( .A1(n2288), .A2(n2705), .ZN(n2823) );
  OR2_X1 U2903 ( .A1(n2831), .A2(n2828), .ZN(n2895) );
  XOR2_X1 U2904 ( .A(n2934), .B(n2935), .Z(n2828) );
  XOR2_X1 U2905 ( .A(n2936), .B(n2937), .Z(n2935) );
  OR2_X1 U2906 ( .A1(n2705), .A2(n2298), .ZN(n2831) );
  OR2_X1 U2907 ( .A1(n2835), .A2(n2832), .ZN(n2892) );
  XNOR2_X1 U2908 ( .A(n2938), .B(n2939), .ZN(n2832) );
  XNOR2_X1 U2909 ( .A(n2940), .B(n2941), .ZN(n2938) );
  OR2_X1 U2910 ( .A1(n2705), .A2(n2303), .ZN(n2835) );
  OR2_X1 U2911 ( .A1(n2839), .A2(n2836), .ZN(n2889) );
  XOR2_X1 U2912 ( .A(n2942), .B(n2943), .Z(n2836) );
  XOR2_X1 U2913 ( .A(n2944), .B(n2945), .Z(n2943) );
  OR2_X1 U2914 ( .A1(n2705), .A2(n2308), .ZN(n2839) );
  XOR2_X1 U2915 ( .A(n2946), .B(n2947), .Z(n2840) );
  XOR2_X1 U2916 ( .A(n2948), .B(n2949), .Z(n2947) );
  OR2_X1 U2917 ( .A1(n2847), .A2(n2844), .ZN(n2883) );
  XOR2_X1 U2918 ( .A(n2950), .B(n2951), .Z(n2844) );
  XOR2_X1 U2919 ( .A(n2952), .B(n2953), .Z(n2951) );
  OR2_X1 U2920 ( .A1(n2705), .A2(n2189), .ZN(n2847) );
  XOR2_X1 U2921 ( .A(n2954), .B(n2955), .Z(n2848) );
  XOR2_X1 U2922 ( .A(n2956), .B(n2957), .Z(n2955) );
  XOR2_X1 U2923 ( .A(n2958), .B(n2959), .Z(n2852) );
  XOR2_X1 U2924 ( .A(n2960), .B(n2961), .Z(n2959) );
  XOR2_X1 U2925 ( .A(n2962), .B(n2963), .Z(n2856) );
  XOR2_X1 U2926 ( .A(n2964), .B(n2965), .Z(n2963) );
  XOR2_X1 U2927 ( .A(n2966), .B(n2967), .Z(n2860) );
  XOR2_X1 U2928 ( .A(n2968), .B(n2969), .Z(n2967) );
  XOR2_X1 U2929 ( .A(n2156), .B(n2970), .Z(n2867) );
  XOR2_X1 U2930 ( .A(n2155), .B(n2154), .Z(n2970) );
  OR2_X1 U2931 ( .A1(n2809), .A2(n1997), .ZN(n2154) );
  OR2_X1 U2932 ( .A1(n2971), .A2(n2972), .ZN(n2155) );
  AND2_X1 U2933 ( .A1(n2969), .A2(n2968), .ZN(n2972) );
  AND2_X1 U2934 ( .A1(n2966), .A2(n2973), .ZN(n2971) );
  OR2_X1 U2935 ( .A1(n2968), .A2(n2969), .ZN(n2973) );
  OR2_X1 U2936 ( .A1(n2809), .A2(n2060), .ZN(n2969) );
  OR2_X1 U2937 ( .A1(n2974), .A2(n2975), .ZN(n2968) );
  AND2_X1 U2938 ( .A1(n2965), .A2(n2964), .ZN(n2975) );
  AND2_X1 U2939 ( .A1(n2962), .A2(n2976), .ZN(n2974) );
  OR2_X1 U2940 ( .A1(n2964), .A2(n2965), .ZN(n2976) );
  OR2_X1 U2941 ( .A1(n2809), .A2(n2093), .ZN(n2965) );
  OR2_X1 U2942 ( .A1(n2977), .A2(n2978), .ZN(n2964) );
  AND2_X1 U2943 ( .A1(n2961), .A2(n2960), .ZN(n2978) );
  AND2_X1 U2944 ( .A1(n2958), .A2(n2979), .ZN(n2977) );
  OR2_X1 U2945 ( .A1(n2960), .A2(n2961), .ZN(n2979) );
  OR2_X1 U2946 ( .A1(n2809), .A2(n2181), .ZN(n2961) );
  OR2_X1 U2947 ( .A1(n2980), .A2(n2981), .ZN(n2960) );
  AND2_X1 U2948 ( .A1(n2957), .A2(n2956), .ZN(n2981) );
  AND2_X1 U2949 ( .A1(n2954), .A2(n2982), .ZN(n2980) );
  OR2_X1 U2950 ( .A1(n2956), .A2(n2957), .ZN(n2982) );
  OR2_X1 U2951 ( .A1(n2809), .A2(n2189), .ZN(n2957) );
  OR2_X1 U2952 ( .A1(n2983), .A2(n2984), .ZN(n2956) );
  AND2_X1 U2953 ( .A1(n2950), .A2(n2953), .ZN(n2984) );
  AND2_X1 U2954 ( .A1(n2985), .A2(n2952), .ZN(n2983) );
  OR2_X1 U2955 ( .A1(n2986), .A2(n2987), .ZN(n2952) );
  AND2_X1 U2956 ( .A1(n2949), .A2(n2948), .ZN(n2987) );
  AND2_X1 U2957 ( .A1(n2946), .A2(n2988), .ZN(n2986) );
  OR2_X1 U2958 ( .A1(n2948), .A2(n2949), .ZN(n2988) );
  OR2_X1 U2959 ( .A1(n2809), .A2(n2308), .ZN(n2949) );
  OR2_X1 U2960 ( .A1(n2989), .A2(n2990), .ZN(n2948) );
  AND2_X1 U2961 ( .A1(n2942), .A2(n2945), .ZN(n2990) );
  AND2_X1 U2962 ( .A1(n2991), .A2(n2944), .ZN(n2989) );
  OR2_X1 U2963 ( .A1(n2992), .A2(n2993), .ZN(n2944) );
  AND2_X1 U2964 ( .A1(n2939), .A2(n2941), .ZN(n2993) );
  AND2_X1 U2965 ( .A1(n2994), .A2(n2940), .ZN(n2992) );
  OR2_X1 U2966 ( .A1(n2941), .A2(n2939), .ZN(n2994) );
  XOR2_X1 U2967 ( .A(n2995), .B(n2996), .Z(n2939) );
  XOR2_X1 U2968 ( .A(n2997), .B(n2998), .Z(n2996) );
  OR2_X1 U2969 ( .A1(n2999), .A2(n3000), .ZN(n2941) );
  AND2_X1 U2970 ( .A1(n2934), .A2(n2937), .ZN(n3000) );
  AND2_X1 U2971 ( .A1(n3001), .A2(n2936), .ZN(n2999) );
  OR2_X1 U2972 ( .A1(n3002), .A2(n3003), .ZN(n2936) );
  AND2_X1 U2973 ( .A1(n2899), .A2(n2902), .ZN(n3003) );
  AND2_X1 U2974 ( .A1(n3004), .A2(n2901), .ZN(n3002) );
  OR2_X1 U2975 ( .A1(n3005), .A2(n3006), .ZN(n2901) );
  AND2_X1 U2976 ( .A1(n2930), .A2(n2933), .ZN(n3006) );
  AND2_X1 U2977 ( .A1(n3007), .A2(n2932), .ZN(n3005) );
  OR2_X1 U2978 ( .A1(n3008), .A2(n3009), .ZN(n2932) );
  AND2_X1 U2979 ( .A1(n2927), .A2(n2929), .ZN(n3009) );
  AND2_X1 U2980 ( .A1(n3010), .A2(n2928), .ZN(n3008) );
  OR2_X1 U2981 ( .A1(n3011), .A2(n3012), .ZN(n2928) );
  AND2_X1 U2982 ( .A1(n2922), .A2(n2925), .ZN(n3012) );
  AND2_X1 U2983 ( .A1(n2924), .A2(n3013), .ZN(n3011) );
  OR2_X1 U2984 ( .A1(n2925), .A2(n2922), .ZN(n3013) );
  OR2_X1 U2985 ( .A1(n2269), .A2(n2809), .ZN(n2922) );
  OR3_X1 U2986 ( .A1(n2395), .A2(n2809), .A3(n2159), .ZN(n2925) );
  INV_X1 U2987 ( .A(n3014), .ZN(n2924) );
  OR2_X1 U2988 ( .A1(n3015), .A2(n3016), .ZN(n3014) );
  AND2_X1 U2989 ( .A1(b_7_), .A2(n3017), .ZN(n3016) );
  OR2_X1 U2990 ( .A1(n3018), .A2(n1880), .ZN(n3017) );
  AND2_X1 U2991 ( .A1(a_14_), .A2(n2120), .ZN(n3018) );
  AND2_X1 U2992 ( .A1(b_6_), .A2(n3019), .ZN(n3015) );
  OR2_X1 U2993 ( .A1(n3020), .A2(n1884), .ZN(n3019) );
  AND2_X1 U2994 ( .A1(a_15_), .A2(n2159), .ZN(n3020) );
  OR2_X1 U2995 ( .A1(n2929), .A2(n2927), .ZN(n3010) );
  XNOR2_X1 U2996 ( .A(n3021), .B(n3022), .ZN(n2927) );
  XNOR2_X1 U2997 ( .A(n3023), .B(n3024), .ZN(n3022) );
  OR2_X1 U2998 ( .A1(n2278), .A2(n2809), .ZN(n2929) );
  OR2_X1 U2999 ( .A1(n2933), .A2(n2930), .ZN(n3007) );
  XNOR2_X1 U3000 ( .A(n3025), .B(n3026), .ZN(n2930) );
  XNOR2_X1 U3001 ( .A(n3027), .B(n3028), .ZN(n3025) );
  OR2_X1 U3002 ( .A1(n2283), .A2(n2809), .ZN(n2933) );
  OR2_X1 U3003 ( .A1(n2902), .A2(n2899), .ZN(n3004) );
  XOR2_X1 U3004 ( .A(n3029), .B(n3030), .Z(n2899) );
  XOR2_X1 U3005 ( .A(n3031), .B(n3032), .Z(n3030) );
  OR2_X1 U3006 ( .A1(n2288), .A2(n2809), .ZN(n2902) );
  OR2_X1 U3007 ( .A1(n2937), .A2(n2934), .ZN(n3001) );
  XOR2_X1 U3008 ( .A(n3033), .B(n3034), .Z(n2934) );
  XOR2_X1 U3009 ( .A(n3035), .B(n3036), .Z(n3034) );
  OR2_X1 U3010 ( .A1(n2293), .A2(n2809), .ZN(n2937) );
  OR2_X1 U3011 ( .A1(n2945), .A2(n2942), .ZN(n2991) );
  XOR2_X1 U3012 ( .A(n3037), .B(n3038), .Z(n2942) );
  XOR2_X1 U3013 ( .A(n3039), .B(n3040), .Z(n3038) );
  OR2_X1 U3014 ( .A1(n2809), .A2(n2303), .ZN(n2945) );
  XNOR2_X1 U3015 ( .A(n3041), .B(n3042), .ZN(n2946) );
  XNOR2_X1 U3016 ( .A(n3043), .B(n3044), .ZN(n3041) );
  OR2_X1 U3017 ( .A1(n2953), .A2(n2950), .ZN(n2985) );
  XOR2_X1 U3018 ( .A(n3045), .B(n3046), .Z(n2950) );
  XOR2_X1 U3019 ( .A(n3047), .B(n3048), .Z(n3046) );
  OR2_X1 U3020 ( .A1(n2809), .A2(n2313), .ZN(n2953) );
  XOR2_X1 U3021 ( .A(n3049), .B(n3050), .Z(n2954) );
  XOR2_X1 U3022 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR2_X1 U3023 ( .A(n3053), .B(n3054), .Z(n2958) );
  XOR2_X1 U3024 ( .A(n3055), .B(n3056), .Z(n3054) );
  XOR2_X1 U3025 ( .A(n3057), .B(n3058), .Z(n2962) );
  XOR2_X1 U3026 ( .A(n3059), .B(n3060), .Z(n3058) );
  XOR2_X1 U3027 ( .A(n3061), .B(n3062), .Z(n2966) );
  XOR2_X1 U3028 ( .A(n3063), .B(n3064), .Z(n3062) );
  XOR2_X1 U3029 ( .A(n2164), .B(n3065), .Z(n2156) );
  XOR2_X1 U3030 ( .A(n2163), .B(n2162), .Z(n3065) );
  OR2_X1 U3031 ( .A1(n2159), .A2(n2060), .ZN(n2162) );
  OR2_X1 U3032 ( .A1(n3066), .A2(n3067), .ZN(n2163) );
  AND2_X1 U3033 ( .A1(n3064), .A2(n3063), .ZN(n3067) );
  AND2_X1 U3034 ( .A1(n3061), .A2(n3068), .ZN(n3066) );
  OR2_X1 U3035 ( .A1(n3063), .A2(n3064), .ZN(n3068) );
  OR2_X1 U3036 ( .A1(n2159), .A2(n2093), .ZN(n3064) );
  OR2_X1 U3037 ( .A1(n3069), .A2(n3070), .ZN(n3063) );
  AND2_X1 U3038 ( .A1(n3060), .A2(n3059), .ZN(n3070) );
  AND2_X1 U3039 ( .A1(n3057), .A2(n3071), .ZN(n3069) );
  OR2_X1 U3040 ( .A1(n3059), .A2(n3060), .ZN(n3071) );
  OR2_X1 U3041 ( .A1(n2159), .A2(n2181), .ZN(n3060) );
  OR2_X1 U3042 ( .A1(n3072), .A2(n3073), .ZN(n3059) );
  AND2_X1 U3043 ( .A1(n3056), .A2(n3055), .ZN(n3073) );
  AND2_X1 U3044 ( .A1(n3053), .A2(n3074), .ZN(n3072) );
  OR2_X1 U3045 ( .A1(n3055), .A2(n3056), .ZN(n3074) );
  OR2_X1 U3046 ( .A1(n2159), .A2(n2189), .ZN(n3056) );
  OR2_X1 U3047 ( .A1(n3075), .A2(n3076), .ZN(n3055) );
  AND2_X1 U3048 ( .A1(n3052), .A2(n3051), .ZN(n3076) );
  AND2_X1 U3049 ( .A1(n3049), .A2(n3077), .ZN(n3075) );
  OR2_X1 U3050 ( .A1(n3051), .A2(n3052), .ZN(n3077) );
  OR2_X1 U3051 ( .A1(n2159), .A2(n2313), .ZN(n3052) );
  OR2_X1 U3052 ( .A1(n3078), .A2(n3079), .ZN(n3051) );
  AND2_X1 U3053 ( .A1(n3045), .A2(n3048), .ZN(n3079) );
  AND2_X1 U3054 ( .A1(n3080), .A2(n3047), .ZN(n3078) );
  OR2_X1 U3055 ( .A1(n3081), .A2(n3082), .ZN(n3047) );
  AND2_X1 U3056 ( .A1(n3042), .A2(n3044), .ZN(n3082) );
  AND2_X1 U3057 ( .A1(n3083), .A2(n3043), .ZN(n3081) );
  OR2_X1 U3058 ( .A1(n3042), .A2(n3044), .ZN(n3083) );
  OR2_X1 U3059 ( .A1(n3084), .A2(n3085), .ZN(n3044) );
  AND2_X1 U3060 ( .A1(n3037), .A2(n3040), .ZN(n3085) );
  AND2_X1 U3061 ( .A1(n3086), .A2(n3039), .ZN(n3084) );
  OR2_X1 U3062 ( .A1(n3087), .A2(n3088), .ZN(n3039) );
  AND2_X1 U3063 ( .A1(n2995), .A2(n2998), .ZN(n3088) );
  AND2_X1 U3064 ( .A1(n3089), .A2(n2997), .ZN(n3087) );
  OR2_X1 U3065 ( .A1(n3090), .A2(n3091), .ZN(n2997) );
  AND2_X1 U3066 ( .A1(n3033), .A2(n3036), .ZN(n3091) );
  AND2_X1 U3067 ( .A1(n3092), .A2(n3035), .ZN(n3090) );
  OR2_X1 U3068 ( .A1(n3093), .A2(n3094), .ZN(n3035) );
  AND2_X1 U3069 ( .A1(n3029), .A2(n3032), .ZN(n3094) );
  AND2_X1 U3070 ( .A1(n3095), .A2(n3031), .ZN(n3093) );
  OR2_X1 U3071 ( .A1(n3096), .A2(n3097), .ZN(n3031) );
  AND2_X1 U3072 ( .A1(n3026), .A2(n3028), .ZN(n3097) );
  AND2_X1 U3073 ( .A1(n3098), .A2(n3027), .ZN(n3096) );
  OR2_X1 U3074 ( .A1(n3099), .A2(n3100), .ZN(n3027) );
  AND2_X1 U3075 ( .A1(n3021), .A2(n3024), .ZN(n3100) );
  AND2_X1 U3076 ( .A1(n3023), .A2(n3101), .ZN(n3099) );
  OR2_X1 U3077 ( .A1(n3024), .A2(n3021), .ZN(n3101) );
  OR2_X1 U3078 ( .A1(n2269), .A2(n2159), .ZN(n3021) );
  OR3_X1 U3079 ( .A1(n2395), .A2(n2159), .A3(n2120), .ZN(n3024) );
  INV_X1 U3080 ( .A(n3102), .ZN(n3023) );
  OR2_X1 U3081 ( .A1(n3103), .A2(n3104), .ZN(n3102) );
  AND2_X1 U3082 ( .A1(b_6_), .A2(n3105), .ZN(n3104) );
  OR2_X1 U3083 ( .A1(n3106), .A2(n1880), .ZN(n3105) );
  AND2_X1 U3084 ( .A1(a_14_), .A2(n2078), .ZN(n3106) );
  AND2_X1 U3085 ( .A1(b_5_), .A2(n3107), .ZN(n3103) );
  OR2_X1 U3086 ( .A1(n3108), .A2(n1884), .ZN(n3107) );
  AND2_X1 U3087 ( .A1(a_15_), .A2(n2120), .ZN(n3108) );
  OR2_X1 U3088 ( .A1(n3028), .A2(n3026), .ZN(n3098) );
  XNOR2_X1 U3089 ( .A(n3109), .B(n3110), .ZN(n3026) );
  XNOR2_X1 U3090 ( .A(n3111), .B(n3112), .ZN(n3110) );
  OR2_X1 U3091 ( .A1(n2278), .A2(n2159), .ZN(n3028) );
  OR2_X1 U3092 ( .A1(n3032), .A2(n3029), .ZN(n3095) );
  XNOR2_X1 U3093 ( .A(n3113), .B(n3114), .ZN(n3029) );
  XNOR2_X1 U3094 ( .A(n3115), .B(n3116), .ZN(n3113) );
  OR2_X1 U3095 ( .A1(n2283), .A2(n2159), .ZN(n3032) );
  OR2_X1 U3096 ( .A1(n3036), .A2(n3033), .ZN(n3092) );
  XOR2_X1 U3097 ( .A(n3117), .B(n3118), .Z(n3033) );
  XOR2_X1 U3098 ( .A(n3119), .B(n3120), .Z(n3118) );
  OR2_X1 U3099 ( .A1(n2288), .A2(n2159), .ZN(n3036) );
  OR2_X1 U3100 ( .A1(n2998), .A2(n2995), .ZN(n3089) );
  XOR2_X1 U3101 ( .A(n3121), .B(n3122), .Z(n2995) );
  XOR2_X1 U3102 ( .A(n3123), .B(n3124), .Z(n3122) );
  OR2_X1 U3103 ( .A1(n2293), .A2(n2159), .ZN(n2998) );
  OR2_X1 U3104 ( .A1(n3040), .A2(n3037), .ZN(n3086) );
  XOR2_X1 U3105 ( .A(n3125), .B(n3126), .Z(n3037) );
  XOR2_X1 U3106 ( .A(n3127), .B(n3128), .Z(n3126) );
  OR2_X1 U3107 ( .A1(n2298), .A2(n2159), .ZN(n3040) );
  XOR2_X1 U3108 ( .A(n3129), .B(n3130), .Z(n3042) );
  XOR2_X1 U3109 ( .A(n3131), .B(n3132), .Z(n3130) );
  OR2_X1 U3110 ( .A1(n3048), .A2(n3045), .ZN(n3080) );
  XOR2_X1 U3111 ( .A(n3133), .B(n3134), .Z(n3045) );
  XOR2_X1 U3112 ( .A(n3135), .B(n3136), .Z(n3134) );
  OR2_X1 U3113 ( .A1(n2159), .A2(n2308), .ZN(n3048) );
  XNOR2_X1 U3114 ( .A(n3137), .B(n3138), .ZN(n3049) );
  XNOR2_X1 U3115 ( .A(n3139), .B(n3140), .ZN(n3137) );
  XOR2_X1 U3116 ( .A(n3141), .B(n3142), .Z(n3053) );
  XOR2_X1 U3117 ( .A(n3143), .B(n3144), .Z(n3142) );
  XOR2_X1 U3118 ( .A(n3145), .B(n3146), .Z(n3057) );
  XOR2_X1 U3119 ( .A(n3147), .B(n3148), .Z(n3146) );
  XOR2_X1 U3120 ( .A(n3149), .B(n3150), .Z(n3061) );
  XOR2_X1 U3121 ( .A(n3151), .B(n3152), .Z(n3150) );
  XOR2_X1 U3122 ( .A(n2171), .B(n3153), .Z(n2164) );
  XOR2_X1 U3123 ( .A(n2170), .B(n2169), .Z(n3153) );
  OR2_X1 U3124 ( .A1(n2120), .A2(n2093), .ZN(n2169) );
  OR2_X1 U3125 ( .A1(n3154), .A2(n3155), .ZN(n2170) );
  AND2_X1 U3126 ( .A1(n3152), .A2(n3151), .ZN(n3155) );
  AND2_X1 U3127 ( .A1(n3149), .A2(n3156), .ZN(n3154) );
  OR2_X1 U3128 ( .A1(n3151), .A2(n3152), .ZN(n3156) );
  OR2_X1 U3129 ( .A1(n2120), .A2(n2181), .ZN(n3152) );
  OR2_X1 U3130 ( .A1(n3157), .A2(n3158), .ZN(n3151) );
  AND2_X1 U3131 ( .A1(n3148), .A2(n3147), .ZN(n3158) );
  AND2_X1 U3132 ( .A1(n3145), .A2(n3159), .ZN(n3157) );
  OR2_X1 U3133 ( .A1(n3147), .A2(n3148), .ZN(n3159) );
  OR2_X1 U3134 ( .A1(n2120), .A2(n2189), .ZN(n3148) );
  OR2_X1 U3135 ( .A1(n3160), .A2(n3161), .ZN(n3147) );
  AND2_X1 U3136 ( .A1(n3144), .A2(n3143), .ZN(n3161) );
  AND2_X1 U3137 ( .A1(n3141), .A2(n3162), .ZN(n3160) );
  OR2_X1 U3138 ( .A1(n3143), .A2(n3144), .ZN(n3162) );
  OR2_X1 U3139 ( .A1(n2120), .A2(n2313), .ZN(n3144) );
  OR2_X1 U3140 ( .A1(n3163), .A2(n3164), .ZN(n3143) );
  AND2_X1 U3141 ( .A1(n3138), .A2(n3140), .ZN(n3164) );
  AND2_X1 U3142 ( .A1(n3165), .A2(n3139), .ZN(n3163) );
  OR2_X1 U3143 ( .A1(n3138), .A2(n3140), .ZN(n3165) );
  OR2_X1 U3144 ( .A1(n3166), .A2(n3167), .ZN(n3140) );
  AND2_X1 U3145 ( .A1(n3133), .A2(n3136), .ZN(n3167) );
  AND2_X1 U3146 ( .A1(n3168), .A2(n3135), .ZN(n3166) );
  OR2_X1 U3147 ( .A1(n3169), .A2(n3170), .ZN(n3135) );
  AND2_X1 U3148 ( .A1(n3132), .A2(n3131), .ZN(n3170) );
  AND2_X1 U3149 ( .A1(n3129), .A2(n3171), .ZN(n3169) );
  OR2_X1 U3150 ( .A1(n3131), .A2(n3132), .ZN(n3171) );
  OR2_X1 U3151 ( .A1(n2298), .A2(n2120), .ZN(n3132) );
  OR2_X1 U3152 ( .A1(n3172), .A2(n3173), .ZN(n3131) );
  AND2_X1 U3153 ( .A1(n3125), .A2(n3128), .ZN(n3173) );
  AND2_X1 U3154 ( .A1(n3174), .A2(n3127), .ZN(n3172) );
  OR2_X1 U3155 ( .A1(n3175), .A2(n3176), .ZN(n3127) );
  AND2_X1 U3156 ( .A1(n3121), .A2(n3124), .ZN(n3176) );
  AND2_X1 U3157 ( .A1(n3177), .A2(n3123), .ZN(n3175) );
  OR2_X1 U3158 ( .A1(n3178), .A2(n3179), .ZN(n3123) );
  AND2_X1 U3159 ( .A1(n3117), .A2(n3120), .ZN(n3179) );
  AND2_X1 U3160 ( .A1(n3180), .A2(n3119), .ZN(n3178) );
  OR2_X1 U3161 ( .A1(n3181), .A2(n3182), .ZN(n3119) );
  AND2_X1 U3162 ( .A1(n3114), .A2(n3116), .ZN(n3182) );
  AND2_X1 U3163 ( .A1(n3183), .A2(n3115), .ZN(n3181) );
  OR2_X1 U3164 ( .A1(n3184), .A2(n3185), .ZN(n3115) );
  AND2_X1 U3165 ( .A1(n3109), .A2(n3112), .ZN(n3185) );
  AND2_X1 U3166 ( .A1(n3111), .A2(n3186), .ZN(n3184) );
  OR2_X1 U3167 ( .A1(n3112), .A2(n3109), .ZN(n3186) );
  OR2_X1 U3168 ( .A1(n2269), .A2(n2120), .ZN(n3109) );
  OR3_X1 U3169 ( .A1(n2395), .A2(n2120), .A3(n2078), .ZN(n3112) );
  INV_X1 U3170 ( .A(n3187), .ZN(n3111) );
  OR2_X1 U3171 ( .A1(n3188), .A2(n3189), .ZN(n3187) );
  AND2_X1 U3172 ( .A1(b_5_), .A2(n3190), .ZN(n3189) );
  OR2_X1 U3173 ( .A1(n3191), .A2(n1880), .ZN(n3190) );
  AND2_X1 U3174 ( .A1(a_14_), .A2(n2052), .ZN(n3191) );
  AND2_X1 U3175 ( .A1(b_4_), .A2(n3192), .ZN(n3188) );
  OR2_X1 U3176 ( .A1(n3193), .A2(n1884), .ZN(n3192) );
  AND2_X1 U3177 ( .A1(a_15_), .A2(n2078), .ZN(n3193) );
  OR2_X1 U3178 ( .A1(n3116), .A2(n3114), .ZN(n3183) );
  XNOR2_X1 U3179 ( .A(n3194), .B(n3195), .ZN(n3114) );
  XNOR2_X1 U3180 ( .A(n3196), .B(n3197), .ZN(n3195) );
  OR2_X1 U3181 ( .A1(n2278), .A2(n2120), .ZN(n3116) );
  OR2_X1 U3182 ( .A1(n3120), .A2(n3117), .ZN(n3180) );
  XNOR2_X1 U3183 ( .A(n3198), .B(n3199), .ZN(n3117) );
  XNOR2_X1 U3184 ( .A(n3200), .B(n3201), .ZN(n3198) );
  OR2_X1 U3185 ( .A1(n2283), .A2(n2120), .ZN(n3120) );
  OR2_X1 U3186 ( .A1(n3124), .A2(n3121), .ZN(n3177) );
  XOR2_X1 U3187 ( .A(n3202), .B(n3203), .Z(n3121) );
  XOR2_X1 U3188 ( .A(n3204), .B(n3205), .Z(n3203) );
  OR2_X1 U3189 ( .A1(n2288), .A2(n2120), .ZN(n3124) );
  OR2_X1 U3190 ( .A1(n3128), .A2(n3125), .ZN(n3174) );
  XOR2_X1 U3191 ( .A(n3206), .B(n3207), .Z(n3125) );
  XOR2_X1 U3192 ( .A(n3208), .B(n3209), .Z(n3207) );
  OR2_X1 U3193 ( .A1(n2293), .A2(n2120), .ZN(n3128) );
  XOR2_X1 U3194 ( .A(n3210), .B(n3211), .Z(n3129) );
  XOR2_X1 U3195 ( .A(n3212), .B(n3213), .Z(n3211) );
  OR2_X1 U3196 ( .A1(n3136), .A2(n3133), .ZN(n3168) );
  XOR2_X1 U3197 ( .A(n3214), .B(n3215), .Z(n3133) );
  XOR2_X1 U3198 ( .A(n3216), .B(n3217), .Z(n3215) );
  OR2_X1 U3199 ( .A1(n2303), .A2(n2120), .ZN(n3136) );
  XOR2_X1 U3200 ( .A(n3218), .B(n3219), .Z(n3138) );
  XOR2_X1 U3201 ( .A(n3220), .B(n3221), .Z(n3219) );
  XOR2_X1 U3202 ( .A(n3222), .B(n3223), .Z(n3141) );
  XOR2_X1 U3203 ( .A(n3224), .B(n3225), .Z(n3223) );
  XNOR2_X1 U3204 ( .A(n3226), .B(n3227), .ZN(n3145) );
  XNOR2_X1 U3205 ( .A(n3228), .B(n3229), .ZN(n3226) );
  XOR2_X1 U3206 ( .A(n3230), .B(n3231), .Z(n3149) );
  XOR2_X1 U3207 ( .A(n3232), .B(n3233), .Z(n3231) );
  XOR2_X1 U3208 ( .A(n2178), .B(n3234), .Z(n2171) );
  XOR2_X1 U3209 ( .A(n2177), .B(n2176), .Z(n3234) );
  OR2_X1 U3210 ( .A1(n2078), .A2(n2181), .ZN(n2176) );
  OR2_X1 U3211 ( .A1(n3235), .A2(n3236), .ZN(n2177) );
  AND2_X1 U3212 ( .A1(n3233), .A2(n3232), .ZN(n3236) );
  AND2_X1 U3213 ( .A1(n3230), .A2(n3237), .ZN(n3235) );
  OR2_X1 U3214 ( .A1(n3232), .A2(n3233), .ZN(n3237) );
  OR2_X1 U3215 ( .A1(n2078), .A2(n2189), .ZN(n3233) );
  OR2_X1 U3216 ( .A1(n3238), .A2(n3239), .ZN(n3232) );
  AND2_X1 U3217 ( .A1(n3227), .A2(n3229), .ZN(n3239) );
  AND2_X1 U3218 ( .A1(n3240), .A2(n3228), .ZN(n3238) );
  OR2_X1 U3219 ( .A1(n3227), .A2(n3229), .ZN(n3240) );
  OR2_X1 U3220 ( .A1(n3241), .A2(n3242), .ZN(n3229) );
  AND2_X1 U3221 ( .A1(n3225), .A2(n3224), .ZN(n3242) );
  AND2_X1 U3222 ( .A1(n3222), .A2(n3243), .ZN(n3241) );
  OR2_X1 U3223 ( .A1(n3224), .A2(n3225), .ZN(n3243) );
  OR2_X1 U3224 ( .A1(n2308), .A2(n2078), .ZN(n3225) );
  OR2_X1 U3225 ( .A1(n3244), .A2(n3245), .ZN(n3224) );
  AND2_X1 U3226 ( .A1(n3221), .A2(n3220), .ZN(n3245) );
  AND2_X1 U3227 ( .A1(n3218), .A2(n3246), .ZN(n3244) );
  OR2_X1 U3228 ( .A1(n3220), .A2(n3221), .ZN(n3246) );
  OR2_X1 U3229 ( .A1(n2303), .A2(n2078), .ZN(n3221) );
  OR2_X1 U3230 ( .A1(n3247), .A2(n3248), .ZN(n3220) );
  AND2_X1 U3231 ( .A1(n3214), .A2(n3217), .ZN(n3248) );
  AND2_X1 U3232 ( .A1(n3249), .A2(n3216), .ZN(n3247) );
  OR2_X1 U3233 ( .A1(n3250), .A2(n3251), .ZN(n3216) );
  AND2_X1 U3234 ( .A1(n3213), .A2(n3212), .ZN(n3251) );
  AND2_X1 U3235 ( .A1(n3210), .A2(n3252), .ZN(n3250) );
  OR2_X1 U3236 ( .A1(n3212), .A2(n3213), .ZN(n3252) );
  OR2_X1 U3237 ( .A1(n2293), .A2(n2078), .ZN(n3213) );
  OR2_X1 U3238 ( .A1(n3253), .A2(n3254), .ZN(n3212) );
  AND2_X1 U3239 ( .A1(n3206), .A2(n3209), .ZN(n3254) );
  AND2_X1 U3240 ( .A1(n3255), .A2(n3208), .ZN(n3253) );
  OR2_X1 U3241 ( .A1(n3256), .A2(n3257), .ZN(n3208) );
  AND2_X1 U3242 ( .A1(n3202), .A2(n3205), .ZN(n3257) );
  AND2_X1 U3243 ( .A1(n3258), .A2(n3204), .ZN(n3256) );
  OR2_X1 U3244 ( .A1(n3259), .A2(n3260), .ZN(n3204) );
  AND2_X1 U3245 ( .A1(n3199), .A2(n3201), .ZN(n3260) );
  AND2_X1 U3246 ( .A1(n3261), .A2(n3200), .ZN(n3259) );
  OR2_X1 U3247 ( .A1(n3262), .A2(n3263), .ZN(n3200) );
  AND2_X1 U3248 ( .A1(n3194), .A2(n3197), .ZN(n3263) );
  AND2_X1 U3249 ( .A1(n3196), .A2(n3264), .ZN(n3262) );
  OR2_X1 U3250 ( .A1(n3197), .A2(n3194), .ZN(n3264) );
  OR2_X1 U3251 ( .A1(n2269), .A2(n2078), .ZN(n3194) );
  OR3_X1 U3252 ( .A1(n2395), .A2(n2078), .A3(n2052), .ZN(n3197) );
  INV_X1 U3253 ( .A(n3265), .ZN(n3196) );
  OR2_X1 U3254 ( .A1(n3266), .A2(n3267), .ZN(n3265) );
  AND2_X1 U3255 ( .A1(b_4_), .A2(n3268), .ZN(n3267) );
  OR2_X1 U3256 ( .A1(n3269), .A2(n1880), .ZN(n3268) );
  AND2_X1 U3257 ( .A1(a_14_), .A2(n2025), .ZN(n3269) );
  AND2_X1 U3258 ( .A1(b_3_), .A2(n3270), .ZN(n3266) );
  OR2_X1 U3259 ( .A1(n3271), .A2(n1884), .ZN(n3270) );
  AND2_X1 U3260 ( .A1(a_15_), .A2(n2052), .ZN(n3271) );
  OR2_X1 U3261 ( .A1(n3201), .A2(n3199), .ZN(n3261) );
  XNOR2_X1 U3262 ( .A(n3272), .B(n3273), .ZN(n3199) );
  XNOR2_X1 U3263 ( .A(n3274), .B(n3275), .ZN(n3273) );
  OR2_X1 U3264 ( .A1(n2278), .A2(n2078), .ZN(n3201) );
  OR2_X1 U3265 ( .A1(n3205), .A2(n3202), .ZN(n3258) );
  XNOR2_X1 U3266 ( .A(n3276), .B(n3277), .ZN(n3202) );
  XNOR2_X1 U3267 ( .A(n3278), .B(n3279), .ZN(n3276) );
  OR2_X1 U3268 ( .A1(n2283), .A2(n2078), .ZN(n3205) );
  OR2_X1 U3269 ( .A1(n3209), .A2(n3206), .ZN(n3255) );
  XOR2_X1 U3270 ( .A(n3280), .B(n3281), .Z(n3206) );
  XOR2_X1 U3271 ( .A(n3282), .B(n3283), .Z(n3281) );
  OR2_X1 U3272 ( .A1(n2288), .A2(n2078), .ZN(n3209) );
  XOR2_X1 U3273 ( .A(n3284), .B(n3285), .Z(n3210) );
  XOR2_X1 U3274 ( .A(n3286), .B(n3287), .Z(n3285) );
  OR2_X1 U3275 ( .A1(n3217), .A2(n3214), .ZN(n3249) );
  XOR2_X1 U3276 ( .A(n3288), .B(n3289), .Z(n3214) );
  XOR2_X1 U3277 ( .A(n3290), .B(n3291), .Z(n3289) );
  OR2_X1 U3278 ( .A1(n2298), .A2(n2078), .ZN(n3217) );
  XOR2_X1 U3279 ( .A(n3292), .B(n3293), .Z(n3218) );
  XOR2_X1 U3280 ( .A(n3294), .B(n3295), .Z(n3293) );
  XOR2_X1 U3281 ( .A(n3296), .B(n3297), .Z(n3222) );
  XOR2_X1 U3282 ( .A(n3298), .B(n3299), .Z(n3297) );
  XOR2_X1 U3283 ( .A(n3300), .B(n3301), .Z(n3227) );
  XOR2_X1 U3284 ( .A(n3302), .B(n3303), .Z(n3301) );
  XOR2_X1 U3285 ( .A(n3304), .B(n3305), .Z(n3230) );
  XOR2_X1 U3286 ( .A(n3306), .B(n3307), .Z(n3305) );
  XNOR2_X1 U3287 ( .A(n3308), .B(n2184), .ZN(n2178) );
  XOR2_X1 U3288 ( .A(n2194), .B(n3309), .Z(n2184) );
  XOR2_X1 U3289 ( .A(n2193), .B(n2192), .Z(n3309) );
  OR2_X1 U3290 ( .A1(n2313), .A2(n2025), .ZN(n2192) );
  OR2_X1 U3291 ( .A1(n3310), .A2(n3311), .ZN(n2193) );
  AND2_X1 U3292 ( .A1(n3312), .A2(n3313), .ZN(n3311) );
  AND2_X1 U3293 ( .A1(n3314), .A2(n3315), .ZN(n3310) );
  OR2_X1 U3294 ( .A1(n3313), .A2(n3312), .ZN(n3315) );
  XOR2_X1 U3295 ( .A(n3316), .B(n3317), .Z(n2194) );
  XOR2_X1 U3296 ( .A(n3318), .B(n3319), .Z(n3317) );
  XNOR2_X1 U3297 ( .A(n2187), .B(n2185), .ZN(n3308) );
  OR2_X1 U3298 ( .A1(n3320), .A2(n3321), .ZN(n2185) );
  AND2_X1 U3299 ( .A1(n3307), .A2(n3306), .ZN(n3321) );
  AND2_X1 U3300 ( .A1(n3304), .A2(n3322), .ZN(n3320) );
  OR2_X1 U3301 ( .A1(n3306), .A2(n3307), .ZN(n3322) );
  OR2_X1 U3302 ( .A1(n2313), .A2(n2052), .ZN(n3307) );
  OR2_X1 U3303 ( .A1(n3323), .A2(n3324), .ZN(n3306) );
  AND2_X1 U3304 ( .A1(n3303), .A2(n3302), .ZN(n3324) );
  AND2_X1 U3305 ( .A1(n3300), .A2(n3325), .ZN(n3323) );
  OR2_X1 U3306 ( .A1(n3302), .A2(n3303), .ZN(n3325) );
  OR2_X1 U3307 ( .A1(n2308), .A2(n2052), .ZN(n3303) );
  OR2_X1 U3308 ( .A1(n3326), .A2(n3327), .ZN(n3302) );
  AND2_X1 U3309 ( .A1(n3299), .A2(n3298), .ZN(n3327) );
  AND2_X1 U3310 ( .A1(n3296), .A2(n3328), .ZN(n3326) );
  OR2_X1 U3311 ( .A1(n3298), .A2(n3299), .ZN(n3328) );
  OR2_X1 U3312 ( .A1(n2303), .A2(n2052), .ZN(n3299) );
  OR2_X1 U3313 ( .A1(n3329), .A2(n3330), .ZN(n3298) );
  AND2_X1 U3314 ( .A1(n3295), .A2(n3294), .ZN(n3330) );
  AND2_X1 U3315 ( .A1(n3292), .A2(n3331), .ZN(n3329) );
  OR2_X1 U3316 ( .A1(n3294), .A2(n3295), .ZN(n3331) );
  OR2_X1 U3317 ( .A1(n2298), .A2(n2052), .ZN(n3295) );
  OR2_X1 U3318 ( .A1(n3332), .A2(n3333), .ZN(n3294) );
  AND2_X1 U3319 ( .A1(n3288), .A2(n3291), .ZN(n3333) );
  AND2_X1 U3320 ( .A1(n3334), .A2(n3290), .ZN(n3332) );
  OR2_X1 U3321 ( .A1(n3335), .A2(n3336), .ZN(n3290) );
  AND2_X1 U3322 ( .A1(n3287), .A2(n3286), .ZN(n3336) );
  AND2_X1 U3323 ( .A1(n3284), .A2(n3337), .ZN(n3335) );
  OR2_X1 U3324 ( .A1(n3286), .A2(n3287), .ZN(n3337) );
  OR2_X1 U3325 ( .A1(n2288), .A2(n2052), .ZN(n3287) );
  OR2_X1 U3326 ( .A1(n3338), .A2(n3339), .ZN(n3286) );
  AND2_X1 U3327 ( .A1(n3280), .A2(n3283), .ZN(n3339) );
  AND2_X1 U3328 ( .A1(n3340), .A2(n3282), .ZN(n3338) );
  OR2_X1 U3329 ( .A1(n3341), .A2(n3342), .ZN(n3282) );
  AND2_X1 U3330 ( .A1(n3277), .A2(n3279), .ZN(n3342) );
  AND2_X1 U3331 ( .A1(n3343), .A2(n3278), .ZN(n3341) );
  OR2_X1 U3332 ( .A1(n3344), .A2(n3345), .ZN(n3278) );
  AND2_X1 U3333 ( .A1(n3272), .A2(n3275), .ZN(n3345) );
  AND2_X1 U3334 ( .A1(n3274), .A2(n3346), .ZN(n3344) );
  OR2_X1 U3335 ( .A1(n3275), .A2(n3272), .ZN(n3346) );
  OR2_X1 U3336 ( .A1(n2269), .A2(n2052), .ZN(n3272) );
  OR3_X1 U3337 ( .A1(n2395), .A2(n2052), .A3(n2025), .ZN(n3275) );
  INV_X1 U3338 ( .A(n3347), .ZN(n3274) );
  OR2_X1 U3339 ( .A1(n3348), .A2(n3349), .ZN(n3347) );
  AND2_X1 U3340 ( .A1(b_3_), .A2(n3350), .ZN(n3349) );
  OR2_X1 U3341 ( .A1(n3351), .A2(n1880), .ZN(n3350) );
  AND2_X1 U3342 ( .A1(a_14_), .A2(n3352), .ZN(n3351) );
  AND2_X1 U3343 ( .A1(b_2_), .A2(n3353), .ZN(n3348) );
  OR2_X1 U3344 ( .A1(n3354), .A2(n1884), .ZN(n3353) );
  AND2_X1 U3345 ( .A1(a_15_), .A2(n2025), .ZN(n3354) );
  OR2_X1 U3346 ( .A1(n3279), .A2(n3277), .ZN(n3343) );
  XNOR2_X1 U3347 ( .A(n3355), .B(n3356), .ZN(n3277) );
  XNOR2_X1 U3348 ( .A(n3357), .B(n3358), .ZN(n3356) );
  OR2_X1 U3349 ( .A1(n2278), .A2(n2052), .ZN(n3279) );
  OR2_X1 U3350 ( .A1(n3283), .A2(n3280), .ZN(n3340) );
  XNOR2_X1 U3351 ( .A(n3359), .B(n3360), .ZN(n3280) );
  XNOR2_X1 U3352 ( .A(n3361), .B(n3362), .ZN(n3359) );
  OR2_X1 U3353 ( .A1(n2283), .A2(n2052), .ZN(n3283) );
  XOR2_X1 U3354 ( .A(n3363), .B(n3364), .Z(n3284) );
  XOR2_X1 U3355 ( .A(n3365), .B(n3366), .Z(n3364) );
  OR2_X1 U3356 ( .A1(n3291), .A2(n3288), .ZN(n3334) );
  XOR2_X1 U3357 ( .A(n3367), .B(n3368), .Z(n3288) );
  XOR2_X1 U3358 ( .A(n3369), .B(n3370), .Z(n3368) );
  OR2_X1 U3359 ( .A1(n2293), .A2(n2052), .ZN(n3291) );
  XOR2_X1 U3360 ( .A(n3371), .B(n3372), .Z(n3292) );
  XOR2_X1 U3361 ( .A(n3373), .B(n3374), .Z(n3372) );
  XOR2_X1 U3362 ( .A(n3375), .B(n3376), .Z(n3296) );
  XOR2_X1 U3363 ( .A(n3377), .B(n3378), .Z(n3376) );
  XOR2_X1 U3364 ( .A(n3379), .B(n3380), .Z(n3300) );
  XOR2_X1 U3365 ( .A(n3381), .B(n3382), .Z(n3380) );
  XOR2_X1 U3366 ( .A(n3314), .B(n3383), .Z(n3304) );
  XOR2_X1 U3367 ( .A(n3313), .B(n3312), .Z(n3383) );
  OR2_X1 U3368 ( .A1(n2308), .A2(n2025), .ZN(n3312) );
  OR2_X1 U3369 ( .A1(n3384), .A2(n3385), .ZN(n3313) );
  AND2_X1 U3370 ( .A1(n3382), .A2(n3381), .ZN(n3385) );
  AND2_X1 U3371 ( .A1(n3379), .A2(n3386), .ZN(n3384) );
  OR2_X1 U3372 ( .A1(n3381), .A2(n3382), .ZN(n3386) );
  OR2_X1 U3373 ( .A1(n2303), .A2(n2025), .ZN(n3382) );
  OR2_X1 U3374 ( .A1(n3387), .A2(n3388), .ZN(n3381) );
  AND2_X1 U3375 ( .A1(n3378), .A2(n3377), .ZN(n3388) );
  AND2_X1 U3376 ( .A1(n3375), .A2(n3389), .ZN(n3387) );
  OR2_X1 U3377 ( .A1(n3377), .A2(n3378), .ZN(n3389) );
  OR2_X1 U3378 ( .A1(n2298), .A2(n2025), .ZN(n3378) );
  OR2_X1 U3379 ( .A1(n3390), .A2(n3391), .ZN(n3377) );
  AND2_X1 U3380 ( .A1(n3374), .A2(n3373), .ZN(n3391) );
  AND2_X1 U3381 ( .A1(n3371), .A2(n3392), .ZN(n3390) );
  OR2_X1 U3382 ( .A1(n3373), .A2(n3374), .ZN(n3392) );
  OR2_X1 U3383 ( .A1(n2293), .A2(n2025), .ZN(n3374) );
  OR2_X1 U3384 ( .A1(n3393), .A2(n3394), .ZN(n3373) );
  AND2_X1 U3385 ( .A1(n3367), .A2(n3370), .ZN(n3394) );
  AND2_X1 U3386 ( .A1(n3395), .A2(n3369), .ZN(n3393) );
  OR2_X1 U3387 ( .A1(n3396), .A2(n3397), .ZN(n3369) );
  AND2_X1 U3388 ( .A1(n3366), .A2(n3365), .ZN(n3397) );
  AND2_X1 U3389 ( .A1(n3363), .A2(n3398), .ZN(n3396) );
  OR2_X1 U3390 ( .A1(n3365), .A2(n3366), .ZN(n3398) );
  OR2_X1 U3391 ( .A1(n2283), .A2(n2025), .ZN(n3366) );
  OR2_X1 U3392 ( .A1(n3399), .A2(n3400), .ZN(n3365) );
  AND2_X1 U3393 ( .A1(n3360), .A2(n3362), .ZN(n3400) );
  AND2_X1 U3394 ( .A1(n3401), .A2(n3361), .ZN(n3399) );
  OR2_X1 U3395 ( .A1(n3402), .A2(n3403), .ZN(n3361) );
  AND2_X1 U3396 ( .A1(n3355), .A2(n3358), .ZN(n3403) );
  AND2_X1 U3397 ( .A1(n3357), .A2(n3404), .ZN(n3402) );
  OR2_X1 U3398 ( .A1(n3358), .A2(n3355), .ZN(n3404) );
  OR2_X1 U3399 ( .A1(n2269), .A2(n2025), .ZN(n3355) );
  OR3_X1 U3400 ( .A1(n2395), .A2(n2025), .A3(n3352), .ZN(n3358) );
  INV_X1 U3401 ( .A(n3405), .ZN(n3357) );
  OR2_X1 U3402 ( .A1(n3406), .A2(n3407), .ZN(n3405) );
  AND2_X1 U3403 ( .A1(b_2_), .A2(n3408), .ZN(n3407) );
  OR2_X1 U3404 ( .A1(n3409), .A2(n1880), .ZN(n3408) );
  AND2_X1 U3405 ( .A1(a_14_), .A2(n3410), .ZN(n3409) );
  AND2_X1 U3406 ( .A1(b_1_), .A2(n3411), .ZN(n3406) );
  OR2_X1 U3407 ( .A1(n3412), .A2(n1884), .ZN(n3411) );
  AND2_X1 U3408 ( .A1(a_15_), .A2(n3352), .ZN(n3412) );
  OR2_X1 U3409 ( .A1(n3362), .A2(n3360), .ZN(n3401) );
  XNOR2_X1 U3410 ( .A(n3413), .B(n3414), .ZN(n3360) );
  XNOR2_X1 U3411 ( .A(n3415), .B(n3416), .ZN(n3414) );
  OR2_X1 U3412 ( .A1(n2278), .A2(n2025), .ZN(n3362) );
  XNOR2_X1 U3413 ( .A(n3417), .B(n3418), .ZN(n3363) );
  XNOR2_X1 U3414 ( .A(n3419), .B(n3420), .ZN(n3417) );
  OR2_X1 U3415 ( .A1(n3370), .A2(n3367), .ZN(n3395) );
  XOR2_X1 U3416 ( .A(n3421), .B(n3422), .Z(n3367) );
  XOR2_X1 U3417 ( .A(n3423), .B(n3424), .Z(n3422) );
  OR2_X1 U3418 ( .A1(n2288), .A2(n2025), .ZN(n3370) );
  XOR2_X1 U3419 ( .A(n3425), .B(n3426), .Z(n3371) );
  XOR2_X1 U3420 ( .A(n3427), .B(n3428), .Z(n3426) );
  XOR2_X1 U3421 ( .A(n3429), .B(n3430), .Z(n3375) );
  XOR2_X1 U3422 ( .A(n3431), .B(n3432), .Z(n3430) );
  XOR2_X1 U3423 ( .A(n3433), .B(n3434), .Z(n3379) );
  XOR2_X1 U3424 ( .A(n3435), .B(n3436), .Z(n3434) );
  XOR2_X1 U3425 ( .A(n3437), .B(n3438), .Z(n3314) );
  XOR2_X1 U3426 ( .A(n3439), .B(n3440), .Z(n3438) );
  AND3_X1 U3427 ( .A1(n1935), .A2(n1933), .A3(n1934), .ZN(n1936) );
  INV_X1 U3428 ( .A(n1998), .ZN(n1934) );
  OR2_X1 U3429 ( .A1(n3441), .A2(n3442), .ZN(n1998) );
  AND2_X1 U3430 ( .A1(n2017), .A2(n2016), .ZN(n3442) );
  AND2_X1 U3431 ( .A1(n2014), .A2(n3443), .ZN(n3441) );
  OR2_X1 U3432 ( .A1(n2016), .A2(n2017), .ZN(n3443) );
  OR2_X1 U3433 ( .A1(n3352), .A2(n1997), .ZN(n2017) );
  OR2_X1 U3434 ( .A1(n3444), .A2(n3445), .ZN(n2016) );
  AND2_X1 U3435 ( .A1(n2035), .A2(n2034), .ZN(n3445) );
  AND2_X1 U3436 ( .A1(n2032), .A2(n3446), .ZN(n3444) );
  OR2_X1 U3437 ( .A1(n2034), .A2(n2035), .ZN(n3446) );
  OR2_X1 U3438 ( .A1(n3352), .A2(n2060), .ZN(n2035) );
  OR2_X1 U3439 ( .A1(n3447), .A2(n3448), .ZN(n2034) );
  AND2_X1 U3440 ( .A1(n2068), .A2(n2070), .ZN(n3448) );
  AND2_X1 U3441 ( .A1(n3449), .A2(n2069), .ZN(n3447) );
  OR2_X1 U3442 ( .A1(n2068), .A2(n2070), .ZN(n3449) );
  OR2_X1 U3443 ( .A1(n3450), .A2(n3451), .ZN(n2070) );
  AND2_X1 U3444 ( .A1(n2103), .A2(n2102), .ZN(n3451) );
  AND2_X1 U3445 ( .A1(n2100), .A2(n3452), .ZN(n3450) );
  OR2_X1 U3446 ( .A1(n2102), .A2(n2103), .ZN(n3452) );
  OR2_X1 U3447 ( .A1(n2181), .A2(n3352), .ZN(n2103) );
  OR2_X1 U3448 ( .A1(n3453), .A2(n3454), .ZN(n2102) );
  AND2_X1 U3449 ( .A1(n2145), .A2(n2144), .ZN(n3454) );
  AND2_X1 U3450 ( .A1(n2142), .A2(n3455), .ZN(n3453) );
  OR2_X1 U3451 ( .A1(n2144), .A2(n2145), .ZN(n3455) );
  OR2_X1 U3452 ( .A1(n2189), .A2(n3352), .ZN(n2145) );
  OR2_X1 U3453 ( .A1(n3456), .A2(n3457), .ZN(n2144) );
  AND2_X1 U3454 ( .A1(n2199), .A2(n2198), .ZN(n3457) );
  AND2_X1 U3455 ( .A1(n2196), .A2(n3458), .ZN(n3456) );
  OR2_X1 U3456 ( .A1(n2198), .A2(n2199), .ZN(n3458) );
  OR2_X1 U3457 ( .A1(n2313), .A2(n3352), .ZN(n2199) );
  OR2_X1 U3458 ( .A1(n3459), .A2(n3460), .ZN(n2198) );
  AND2_X1 U3459 ( .A1(n3319), .A2(n3318), .ZN(n3460) );
  AND2_X1 U3460 ( .A1(n3316), .A2(n3461), .ZN(n3459) );
  OR2_X1 U3461 ( .A1(n3318), .A2(n3319), .ZN(n3461) );
  OR2_X1 U3462 ( .A1(n2308), .A2(n3352), .ZN(n3319) );
  OR2_X1 U3463 ( .A1(n3462), .A2(n3463), .ZN(n3318) );
  AND2_X1 U3464 ( .A1(n3440), .A2(n3439), .ZN(n3463) );
  AND2_X1 U3465 ( .A1(n3437), .A2(n3464), .ZN(n3462) );
  OR2_X1 U3466 ( .A1(n3439), .A2(n3440), .ZN(n3464) );
  OR2_X1 U3467 ( .A1(n2303), .A2(n3352), .ZN(n3440) );
  OR2_X1 U3468 ( .A1(n3465), .A2(n3466), .ZN(n3439) );
  AND2_X1 U3469 ( .A1(n3436), .A2(n3435), .ZN(n3466) );
  AND2_X1 U3470 ( .A1(n3433), .A2(n3467), .ZN(n3465) );
  OR2_X1 U3471 ( .A1(n3435), .A2(n3436), .ZN(n3467) );
  OR2_X1 U3472 ( .A1(n2298), .A2(n3352), .ZN(n3436) );
  OR2_X1 U3473 ( .A1(n3468), .A2(n3469), .ZN(n3435) );
  AND2_X1 U3474 ( .A1(n3432), .A2(n3431), .ZN(n3469) );
  AND2_X1 U3475 ( .A1(n3429), .A2(n3470), .ZN(n3468) );
  OR2_X1 U3476 ( .A1(n3431), .A2(n3432), .ZN(n3470) );
  OR2_X1 U3477 ( .A1(n2293), .A2(n3352), .ZN(n3432) );
  OR2_X1 U3478 ( .A1(n3471), .A2(n3472), .ZN(n3431) );
  AND2_X1 U3479 ( .A1(n3428), .A2(n3427), .ZN(n3472) );
  AND2_X1 U3480 ( .A1(n3425), .A2(n3473), .ZN(n3471) );
  OR2_X1 U3481 ( .A1(n3427), .A2(n3428), .ZN(n3473) );
  OR2_X1 U3482 ( .A1(n2288), .A2(n3352), .ZN(n3428) );
  OR2_X1 U3483 ( .A1(n3474), .A2(n3475), .ZN(n3427) );
  AND2_X1 U3484 ( .A1(n3421), .A2(n3424), .ZN(n3475) );
  AND2_X1 U3485 ( .A1(n3476), .A2(n3423), .ZN(n3474) );
  OR2_X1 U3486 ( .A1(n3477), .A2(n3478), .ZN(n3423) );
  AND2_X1 U3487 ( .A1(n3420), .A2(n3419), .ZN(n3478) );
  AND2_X1 U3488 ( .A1(n3418), .A2(n3479), .ZN(n3477) );
  OR2_X1 U3489 ( .A1(n3419), .A2(n3420), .ZN(n3479) );
  OR2_X1 U3490 ( .A1(n2278), .A2(n3352), .ZN(n3420) );
  OR2_X1 U3491 ( .A1(n3480), .A2(n3481), .ZN(n3419) );
  AND2_X1 U3492 ( .A1(n3413), .A2(n3416), .ZN(n3481) );
  AND2_X1 U3493 ( .A1(n3415), .A2(n3482), .ZN(n3480) );
  OR2_X1 U3494 ( .A1(n3416), .A2(n3413), .ZN(n3482) );
  OR2_X1 U3495 ( .A1(n2269), .A2(n3352), .ZN(n3413) );
  OR3_X1 U3496 ( .A1(n2395), .A2(n3352), .A3(n3410), .ZN(n3416) );
  INV_X1 U3497 ( .A(n3483), .ZN(n3415) );
  OR2_X1 U3498 ( .A1(n3484), .A2(n3485), .ZN(n3483) );
  AND2_X1 U3499 ( .A1(b_1_), .A2(n3486), .ZN(n3485) );
  OR2_X1 U3500 ( .A1(n3487), .A2(n1880), .ZN(n3486) );
  AND2_X1 U3501 ( .A1(n3488), .A2(a_14_), .ZN(n1880) );
  AND2_X1 U3502 ( .A1(a_14_), .A2(n3489), .ZN(n3487) );
  AND2_X1 U3503 ( .A1(b_0_), .A2(n3490), .ZN(n3484) );
  OR2_X1 U3504 ( .A1(n3491), .A2(n1884), .ZN(n3490) );
  AND2_X1 U3505 ( .A1(n3492), .A2(a_15_), .ZN(n1884) );
  AND2_X1 U3506 ( .A1(a_15_), .A2(n3410), .ZN(n3491) );
  XNOR2_X1 U3507 ( .A(n3493), .B(n3494), .ZN(n3418) );
  OR2_X1 U3508 ( .A1(n3495), .A2(n3496), .ZN(n3493) );
  INV_X1 U3509 ( .A(n3497), .ZN(n3496) );
  AND2_X1 U3510 ( .A1(n3498), .A2(n3499), .ZN(n3495) );
  OR2_X1 U3511 ( .A1(n3492), .A2(n3489), .ZN(n3498) );
  OR2_X1 U3512 ( .A1(n3424), .A2(n3421), .ZN(n3476) );
  XOR2_X1 U3513 ( .A(n3500), .B(n3501), .Z(n3421) );
  XOR2_X1 U3514 ( .A(n3502), .B(n3503), .Z(n3500) );
  OR2_X1 U3515 ( .A1(n2283), .A2(n3352), .ZN(n3424) );
  XNOR2_X1 U3516 ( .A(n3504), .B(n3505), .ZN(n3425) );
  XNOR2_X1 U3517 ( .A(n3506), .B(n3507), .ZN(n3504) );
  XNOR2_X1 U3518 ( .A(n3508), .B(n3509), .ZN(n3429) );
  XNOR2_X1 U3519 ( .A(n3510), .B(n3511), .ZN(n3508) );
  XNOR2_X1 U3520 ( .A(n3512), .B(n3513), .ZN(n3433) );
  XNOR2_X1 U3521 ( .A(n3514), .B(n3515), .ZN(n3512) );
  XOR2_X1 U3522 ( .A(n3516), .B(n3517), .Z(n3437) );
  XOR2_X1 U3523 ( .A(n3518), .B(n3519), .Z(n3517) );
  XOR2_X1 U3524 ( .A(n3520), .B(n3521), .Z(n3316) );
  XOR2_X1 U3525 ( .A(n3522), .B(n3523), .Z(n3521) );
  XOR2_X1 U3526 ( .A(n3524), .B(n3525), .Z(n2196) );
  XOR2_X1 U3527 ( .A(n3526), .B(n3527), .Z(n3525) );
  XOR2_X1 U3528 ( .A(n3528), .B(n3529), .Z(n2142) );
  XOR2_X1 U3529 ( .A(n3530), .B(n3531), .Z(n3529) );
  XOR2_X1 U3530 ( .A(n3532), .B(n3533), .Z(n2100) );
  XOR2_X1 U3531 ( .A(n3534), .B(n3535), .Z(n3533) );
  XOR2_X1 U3532 ( .A(n3536), .B(n3537), .Z(n2068) );
  XOR2_X1 U3533 ( .A(n3538), .B(n3539), .Z(n3537) );
  XOR2_X1 U3534 ( .A(n3540), .B(n3541), .Z(n2032) );
  XOR2_X1 U3535 ( .A(n3542), .B(n3543), .Z(n3541) );
  XOR2_X1 U3536 ( .A(n3544), .B(n3545), .Z(n2014) );
  XOR2_X1 U3537 ( .A(n3546), .B(n3547), .Z(n3545) );
  XOR2_X1 U3538 ( .A(n3548), .B(n1996), .Z(n1933) );
  OR2_X1 U3539 ( .A1(n3549), .A2(n3550), .ZN(n1996) );
  AND2_X1 U3540 ( .A1(n3551), .A2(n3552), .ZN(n3550) );
  AND2_X1 U3541 ( .A1(n3553), .A2(n3554), .ZN(n3549) );
  OR2_X1 U3542 ( .A1(n3552), .A2(n3551), .ZN(n3553) );
  OR2_X1 U3543 ( .A1(n1997), .A2(n3489), .ZN(n3548) );
  XNOR2_X1 U3544 ( .A(n3551), .B(n3555), .ZN(n1935) );
  XOR2_X1 U3545 ( .A(n3552), .B(n3554), .Z(n3555) );
  OR2_X1 U3546 ( .A1(n3410), .A2(n1997), .ZN(n3554) );
  INV_X1 U3547 ( .A(a_0_), .ZN(n1997) );
  OR2_X1 U3548 ( .A1(n3556), .A2(n3557), .ZN(n3552) );
  AND2_X1 U3549 ( .A1(n3544), .A2(n3546), .ZN(n3557) );
  AND2_X1 U3550 ( .A1(n3558), .A2(n3547), .ZN(n3556) );
  OR2_X1 U3551 ( .A1(n3546), .A2(n3544), .ZN(n3558) );
  OR2_X1 U3552 ( .A1(n2093), .A2(n3489), .ZN(n3544) );
  OR2_X1 U3553 ( .A1(n3559), .A2(n3560), .ZN(n3546) );
  AND2_X1 U3554 ( .A1(n3540), .A2(n3542), .ZN(n3560) );
  AND2_X1 U3555 ( .A1(n3561), .A2(n3543), .ZN(n3559) );
  OR2_X1 U3556 ( .A1(n2181), .A2(n3489), .ZN(n3543) );
  OR2_X1 U3557 ( .A1(n3542), .A2(n3540), .ZN(n3561) );
  OR2_X1 U3558 ( .A1(n2093), .A2(n3410), .ZN(n3540) );
  OR2_X1 U3559 ( .A1(n3562), .A2(n3563), .ZN(n3542) );
  AND2_X1 U3560 ( .A1(n3536), .A2(n3538), .ZN(n3563) );
  AND2_X1 U3561 ( .A1(n3564), .A2(n3539), .ZN(n3562) );
  OR2_X1 U3562 ( .A1(n2189), .A2(n3489), .ZN(n3539) );
  OR2_X1 U3563 ( .A1(n3538), .A2(n3536), .ZN(n3564) );
  OR2_X1 U3564 ( .A1(n2181), .A2(n3410), .ZN(n3536) );
  OR2_X1 U3565 ( .A1(n3565), .A2(n3566), .ZN(n3538) );
  AND2_X1 U3566 ( .A1(n3532), .A2(n3534), .ZN(n3566) );
  AND2_X1 U3567 ( .A1(n3567), .A2(n3535), .ZN(n3565) );
  OR2_X1 U3568 ( .A1(n2313), .A2(n3489), .ZN(n3535) );
  OR2_X1 U3569 ( .A1(n3534), .A2(n3532), .ZN(n3567) );
  OR2_X1 U3570 ( .A1(n2189), .A2(n3410), .ZN(n3532) );
  OR2_X1 U3571 ( .A1(n3568), .A2(n3569), .ZN(n3534) );
  AND2_X1 U3572 ( .A1(n3528), .A2(n3530), .ZN(n3569) );
  AND2_X1 U3573 ( .A1(n3570), .A2(n3531), .ZN(n3568) );
  OR2_X1 U3574 ( .A1(n2308), .A2(n3489), .ZN(n3531) );
  OR2_X1 U3575 ( .A1(n3530), .A2(n3528), .ZN(n3570) );
  OR2_X1 U3576 ( .A1(n2313), .A2(n3410), .ZN(n3528) );
  OR2_X1 U3577 ( .A1(n3571), .A2(n3572), .ZN(n3530) );
  AND2_X1 U3578 ( .A1(n3524), .A2(n3526), .ZN(n3572) );
  AND2_X1 U3579 ( .A1(n3573), .A2(n3527), .ZN(n3571) );
  OR2_X1 U3580 ( .A1(n2303), .A2(n3489), .ZN(n3527) );
  OR2_X1 U3581 ( .A1(n3526), .A2(n3524), .ZN(n3573) );
  OR2_X1 U3582 ( .A1(n2308), .A2(n3410), .ZN(n3524) );
  OR2_X1 U3583 ( .A1(n3574), .A2(n3575), .ZN(n3526) );
  AND2_X1 U3584 ( .A1(n3520), .A2(n3522), .ZN(n3575) );
  AND2_X1 U3585 ( .A1(n3576), .A2(n3523), .ZN(n3574) );
  OR2_X1 U3586 ( .A1(n2298), .A2(n3489), .ZN(n3523) );
  OR2_X1 U3587 ( .A1(n3522), .A2(n3520), .ZN(n3576) );
  OR2_X1 U3588 ( .A1(n2303), .A2(n3410), .ZN(n3520) );
  OR2_X1 U3589 ( .A1(n3577), .A2(n3578), .ZN(n3522) );
  AND2_X1 U3590 ( .A1(n3516), .A2(n3518), .ZN(n3578) );
  AND2_X1 U3591 ( .A1(n3579), .A2(n3519), .ZN(n3577) );
  OR2_X1 U3592 ( .A1(n2293), .A2(n3489), .ZN(n3519) );
  OR2_X1 U3593 ( .A1(n3518), .A2(n3516), .ZN(n3579) );
  OR2_X1 U3594 ( .A1(n2298), .A2(n3410), .ZN(n3516) );
  OR2_X1 U3595 ( .A1(n3580), .A2(n3581), .ZN(n3518) );
  AND2_X1 U3596 ( .A1(n3513), .A2(n3515), .ZN(n3581) );
  AND2_X1 U3597 ( .A1(n3582), .A2(n3514), .ZN(n3580) );
  OR2_X1 U3598 ( .A1(n2288), .A2(n3489), .ZN(n3514) );
  OR2_X1 U3599 ( .A1(n3515), .A2(n3513), .ZN(n3582) );
  OR2_X1 U3600 ( .A1(n2293), .A2(n3410), .ZN(n3513) );
  OR2_X1 U3601 ( .A1(n3583), .A2(n3584), .ZN(n3515) );
  AND2_X1 U3602 ( .A1(n3509), .A2(n3511), .ZN(n3584) );
  AND2_X1 U3603 ( .A1(n3585), .A2(n3510), .ZN(n3583) );
  OR2_X1 U3604 ( .A1(n2283), .A2(n3489), .ZN(n3510) );
  OR2_X1 U3605 ( .A1(n3511), .A2(n3509), .ZN(n3585) );
  OR2_X1 U3606 ( .A1(n2288), .A2(n3410), .ZN(n3509) );
  OR2_X1 U3607 ( .A1(n3586), .A2(n3587), .ZN(n3511) );
  AND2_X1 U3608 ( .A1(n3505), .A2(n3507), .ZN(n3587) );
  AND2_X1 U3609 ( .A1(n3588), .A2(n3506), .ZN(n3586) );
  OR2_X1 U3610 ( .A1(n2278), .A2(n3489), .ZN(n3506) );
  OR2_X1 U3611 ( .A1(n3507), .A2(n3505), .ZN(n3588) );
  OR2_X1 U3612 ( .A1(n2283), .A2(n3410), .ZN(n3505) );
  OR2_X1 U3613 ( .A1(n3589), .A2(n3590), .ZN(n3507) );
  AND2_X1 U3614 ( .A1(n3501), .A2(n3503), .ZN(n3590) );
  AND2_X1 U3615 ( .A1(n3502), .A2(n3591), .ZN(n3589) );
  OR2_X1 U3616 ( .A1(n3503), .A2(n3501), .ZN(n3591) );
  OR2_X1 U3617 ( .A1(n2278), .A2(n3410), .ZN(n3501) );
  OR2_X1 U3618 ( .A1(n2269), .A2(n3489), .ZN(n3503) );
  AND2_X1 U3619 ( .A1(n3497), .A2(n3494), .ZN(n3502) );
  OR3_X1 U3620 ( .A1(n2395), .A2(n3410), .A3(n3489), .ZN(n3494) );
  OR2_X1 U3621 ( .A1(n3492), .A2(n3488), .ZN(n2395) );
  OR3_X1 U3622 ( .A1(n3492), .A2(n3489), .A3(n3499), .ZN(n3497) );
  OR2_X1 U3623 ( .A1(n2269), .A2(n3410), .ZN(n3499) );
  OR2_X1 U3624 ( .A1(n2060), .A2(n3489), .ZN(n3551) );
  INV_X1 U3625 ( .A(b_0_), .ZN(n3489) );
  OR3_X1 U3626 ( .A1(n3592), .A2(n3593), .A3(n3594), .ZN(Result_add_9_) );
  AND2_X1 U3627 ( .A1(n3595), .A2(n3596), .ZN(n3594) );
  AND2_X1 U3628 ( .A1(n3597), .A2(n2705), .ZN(n3593) );
  XNOR2_X1 U3629 ( .A(n2293), .B(n3595), .ZN(n3597) );
  INV_X1 U3630 ( .A(n3598), .ZN(n3595) );
  AND3_X1 U3631 ( .A1(n3598), .A2(n2293), .A3(b_9_), .ZN(n3592) );
  XNOR2_X1 U3632 ( .A(n3599), .B(n3600), .ZN(Result_add_8_) );
  AND2_X1 U3633 ( .A1(n2940), .A2(n3601), .ZN(n3600) );
  INV_X1 U3634 ( .A(n3602), .ZN(n3601) );
  OR3_X1 U3635 ( .A1(n3603), .A2(n3604), .A3(n3605), .ZN(Result_add_7_) );
  INV_X1 U3636 ( .A(n3606), .ZN(n3605) );
  OR2_X1 U3637 ( .A1(n3607), .A2(n3043), .ZN(n3606) );
  AND2_X1 U3638 ( .A1(n3608), .A2(n2159), .ZN(n3604) );
  XNOR2_X1 U3639 ( .A(a_7_), .B(n3607), .ZN(n3608) );
  AND3_X1 U3640 ( .A1(n3607), .A2(n2303), .A3(b_7_), .ZN(n3603) );
  XOR2_X1 U3641 ( .A(n3609), .B(n3610), .Z(Result_add_6_) );
  OR2_X1 U3642 ( .A1(n3611), .A2(n3612), .ZN(n3610) );
  OR3_X1 U3643 ( .A1(n3613), .A2(n3614), .A3(n3615), .ZN(Result_add_5_) );
  INV_X1 U3644 ( .A(n3616), .ZN(n3615) );
  OR2_X1 U3645 ( .A1(n3617), .A2(n3228), .ZN(n3616) );
  AND2_X1 U3646 ( .A1(n3618), .A2(n2078), .ZN(n3614) );
  XNOR2_X1 U3647 ( .A(a_5_), .B(n3617), .ZN(n3618) );
  AND3_X1 U3648 ( .A1(n3617), .A2(n2313), .A3(b_5_), .ZN(n3613) );
  XOR2_X1 U3649 ( .A(n3619), .B(n3620), .Z(Result_add_4_) );
  OR2_X1 U3650 ( .A1(n3621), .A2(n3622), .ZN(n3620) );
  OR3_X1 U3651 ( .A1(n3623), .A2(n3624), .A3(n3625), .ZN(Result_add_3_) );
  INV_X1 U3652 ( .A(n3626), .ZN(n3625) );
  OR2_X1 U3653 ( .A1(n3627), .A2(n2099), .ZN(n3626) );
  AND2_X1 U3654 ( .A1(n3628), .A2(n2025), .ZN(n3624) );
  XNOR2_X1 U3655 ( .A(a_3_), .B(n3627), .ZN(n3628) );
  AND3_X1 U3656 ( .A1(n3627), .A2(n2181), .A3(b_3_), .ZN(n3623) );
  XOR2_X1 U3657 ( .A(n3629), .B(n3630), .Z(Result_add_2_) );
  OR2_X1 U3658 ( .A1(n3631), .A2(n3632), .ZN(n3630) );
  OR3_X1 U3659 ( .A1(n3633), .A2(n3634), .A3(n3635), .ZN(Result_add_1_) );
  INV_X1 U3660 ( .A(n3636), .ZN(n3635) );
  OR2_X1 U3661 ( .A1(n3637), .A2(n3547), .ZN(n3636) );
  AND2_X1 U3662 ( .A1(n3638), .A2(n3410), .ZN(n3634) );
  XNOR2_X1 U3663 ( .A(a_1_), .B(n3637), .ZN(n3638) );
  AND3_X1 U3664 ( .A1(n3637), .A2(n2060), .A3(b_1_), .ZN(n3633) );
  XNOR2_X1 U3665 ( .A(b_15_), .B(n3488), .ZN(Result_add_15_) );
  INV_X1 U3666 ( .A(a_15_), .ZN(n3488) );
  OR3_X1 U3667 ( .A1(n3639), .A2(n3640), .A3(n1890), .ZN(Result_add_14_) );
  AND2_X1 U3668 ( .A1(n2276), .A2(Result_mul_31_), .ZN(n1890) );
  INV_X1 U3669 ( .A(n3641), .ZN(n3640) );
  OR3_X1 U3670 ( .A1(Result_mul_31_), .A2(a_14_), .A3(n1881), .ZN(n3641) );
  AND2_X1 U3671 ( .A1(n3642), .A2(n1881), .ZN(n3639) );
  INV_X1 U3672 ( .A(b_14_), .ZN(n1881) );
  XNOR2_X1 U3673 ( .A(n3492), .B(Result_mul_31_), .ZN(n3642) );
  INV_X1 U3674 ( .A(a_14_), .ZN(n3492) );
  OR3_X1 U3675 ( .A1(n3643), .A2(n3644), .A3(n3645), .ZN(Result_add_13_) );
  AND2_X1 U3676 ( .A1(n2406), .A2(n3646), .ZN(n3645) );
  AND2_X1 U3677 ( .A1(n3647), .A2(n2277), .ZN(n3644) );
  XNOR2_X1 U3678 ( .A(n3648), .B(a_13_), .ZN(n3647) );
  AND3_X1 U3679 ( .A1(n3648), .A2(n2269), .A3(b_13_), .ZN(n3643) );
  XNOR2_X1 U3680 ( .A(n3649), .B(n3650), .ZN(Result_add_12_) );
  AND2_X1 U3681 ( .A1(n2504), .A2(n3651), .ZN(n3650) );
  INV_X1 U3682 ( .A(n3652), .ZN(n3651) );
  OR3_X1 U3683 ( .A1(n3653), .A2(n3654), .A3(n3655), .ZN(Result_add_11_) );
  AND2_X1 U3684 ( .A1(n3656), .A2(n3657), .ZN(n3655) );
  AND2_X1 U3685 ( .A1(n3658), .A2(n2495), .ZN(n3654) );
  XNOR2_X1 U3686 ( .A(n2283), .B(n3656), .ZN(n3658) );
  INV_X1 U3687 ( .A(n3659), .ZN(n3656) );
  AND3_X1 U3688 ( .A1(n3659), .A2(n2283), .A3(b_11_), .ZN(n3653) );
  XNOR2_X1 U3689 ( .A(n3660), .B(n3661), .ZN(Result_add_10_) );
  AND2_X1 U3690 ( .A1(n2716), .A2(n3662), .ZN(n3661) );
  INV_X1 U3691 ( .A(n3663), .ZN(n3662) );
  XOR2_X1 U3692 ( .A(n3664), .B(n3665), .Z(Result_add_0_) );
  XNOR2_X1 U3693 ( .A(a_0_), .B(b_0_), .ZN(n3665) );
  OR2_X1 U3694 ( .A1(n3666), .A2(n3667), .ZN(n3664) );
  AND2_X1 U3695 ( .A1(n2060), .A2(n3410), .ZN(n3667) );
  AND2_X1 U3696 ( .A1(n3637), .A2(n3547), .ZN(n3666) );
  OR2_X1 U3697 ( .A1(n2060), .A2(n3410), .ZN(n3547) );
  INV_X1 U3698 ( .A(b_1_), .ZN(n3410) );
  INV_X1 U3699 ( .A(a_1_), .ZN(n2060) );
  OR2_X1 U3700 ( .A1(n3668), .A2(n3631), .ZN(n3637) );
  AND2_X1 U3701 ( .A1(n2093), .A2(n3352), .ZN(n3631) );
  INV_X1 U3702 ( .A(b_2_), .ZN(n3352) );
  INV_X1 U3703 ( .A(a_2_), .ZN(n2093) );
  AND2_X1 U3704 ( .A1(n3629), .A2(n2069), .ZN(n3668) );
  INV_X1 U3705 ( .A(n3632), .ZN(n2069) );
  AND2_X1 U3706 ( .A1(a_2_), .A2(b_2_), .ZN(n3632) );
  OR2_X1 U3707 ( .A1(n3669), .A2(n3670), .ZN(n3629) );
  AND2_X1 U3708 ( .A1(n2181), .A2(n2025), .ZN(n3670) );
  AND2_X1 U3709 ( .A1(n3627), .A2(n2099), .ZN(n3669) );
  OR2_X1 U3710 ( .A1(n2181), .A2(n2025), .ZN(n2099) );
  INV_X1 U3711 ( .A(b_3_), .ZN(n2025) );
  INV_X1 U3712 ( .A(a_3_), .ZN(n2181) );
  OR2_X1 U3713 ( .A1(n3671), .A2(n3621), .ZN(n3627) );
  AND2_X1 U3714 ( .A1(n2189), .A2(n2052), .ZN(n3621) );
  INV_X1 U3715 ( .A(b_4_), .ZN(n2052) );
  INV_X1 U3716 ( .A(a_4_), .ZN(n2189) );
  AND2_X1 U3717 ( .A1(n3619), .A2(n2187), .ZN(n3671) );
  INV_X1 U3718 ( .A(n3622), .ZN(n2187) );
  AND2_X1 U3719 ( .A1(a_4_), .A2(b_4_), .ZN(n3622) );
  OR2_X1 U3720 ( .A1(n3672), .A2(n3673), .ZN(n3619) );
  AND2_X1 U3721 ( .A1(n2313), .A2(n2078), .ZN(n3673) );
  AND2_X1 U3722 ( .A1(n3617), .A2(n3228), .ZN(n3672) );
  OR2_X1 U3723 ( .A1(n2313), .A2(n2078), .ZN(n3228) );
  INV_X1 U3724 ( .A(b_5_), .ZN(n2078) );
  INV_X1 U3725 ( .A(a_5_), .ZN(n2313) );
  OR2_X1 U3726 ( .A1(n3674), .A2(n3611), .ZN(n3617) );
  AND2_X1 U3727 ( .A1(n2308), .A2(n2120), .ZN(n3611) );
  INV_X1 U3728 ( .A(b_6_), .ZN(n2120) );
  INV_X1 U3729 ( .A(a_6_), .ZN(n2308) );
  AND2_X1 U3730 ( .A1(n3609), .A2(n3139), .ZN(n3674) );
  INV_X1 U3731 ( .A(n3612), .ZN(n3139) );
  AND2_X1 U3732 ( .A1(a_6_), .A2(b_6_), .ZN(n3612) );
  OR2_X1 U3733 ( .A1(n3675), .A2(n3676), .ZN(n3609) );
  AND2_X1 U3734 ( .A1(n2303), .A2(n2159), .ZN(n3676) );
  AND2_X1 U3735 ( .A1(n3607), .A2(n3043), .ZN(n3675) );
  OR2_X1 U3736 ( .A1(n2303), .A2(n2159), .ZN(n3043) );
  INV_X1 U3737 ( .A(b_7_), .ZN(n2159) );
  INV_X1 U3738 ( .A(a_7_), .ZN(n2303) );
  OR2_X1 U3739 ( .A1(n3677), .A2(n3602), .ZN(n3607) );
  AND2_X1 U3740 ( .A1(n2298), .A2(n2809), .ZN(n3602) );
  AND2_X1 U3741 ( .A1(n3599), .A2(n2940), .ZN(n3677) );
  OR2_X1 U3742 ( .A1(n2298), .A2(n2809), .ZN(n2940) );
  INV_X1 U3743 ( .A(b_8_), .ZN(n2809) );
  INV_X1 U3744 ( .A(a_8_), .ZN(n2298) );
  OR2_X1 U3745 ( .A1(n3678), .A2(n3679), .ZN(n3599) );
  AND2_X1 U3746 ( .A1(n2293), .A2(n2705), .ZN(n3679) );
  INV_X1 U3747 ( .A(b_9_), .ZN(n2705) );
  INV_X1 U3748 ( .A(a_9_), .ZN(n2293) );
  AND2_X1 U3749 ( .A1(n3598), .A2(n2826), .ZN(n3678) );
  INV_X1 U3750 ( .A(n3596), .ZN(n2826) );
  AND2_X1 U3751 ( .A1(a_9_), .A2(b_9_), .ZN(n3596) );
  OR2_X1 U3752 ( .A1(n3680), .A2(n3663), .ZN(n3598) );
  AND2_X1 U3753 ( .A1(n2288), .A2(n2597), .ZN(n3663) );
  AND2_X1 U3754 ( .A1(n3660), .A2(n2716), .ZN(n3680) );
  OR2_X1 U3755 ( .A1(n2288), .A2(n2597), .ZN(n2716) );
  INV_X1 U3756 ( .A(b_10_), .ZN(n2597) );
  INV_X1 U3757 ( .A(a_10_), .ZN(n2288) );
  OR2_X1 U3758 ( .A1(n3681), .A2(n3682), .ZN(n3660) );
  AND2_X1 U3759 ( .A1(n2283), .A2(n2495), .ZN(n3682) );
  INV_X1 U3760 ( .A(b_11_), .ZN(n2495) );
  INV_X1 U3761 ( .A(a_11_), .ZN(n2283) );
  AND2_X1 U3762 ( .A1(n3659), .A2(n2606), .ZN(n3681) );
  INV_X1 U3763 ( .A(n3657), .ZN(n2606) );
  AND2_X1 U3764 ( .A1(a_11_), .A2(b_11_), .ZN(n3657) );
  OR2_X1 U3765 ( .A1(n3683), .A2(n3652), .ZN(n3659) );
  AND2_X1 U3766 ( .A1(n2278), .A2(n2401), .ZN(n3652) );
  AND2_X1 U3767 ( .A1(n3649), .A2(n2504), .ZN(n3683) );
  OR2_X1 U3768 ( .A1(n2278), .A2(n2401), .ZN(n2504) );
  INV_X1 U3769 ( .A(b_12_), .ZN(n2401) );
  INV_X1 U3770 ( .A(a_12_), .ZN(n2278) );
  OR2_X1 U3771 ( .A1(n3684), .A2(n3685), .ZN(n3649) );
  AND2_X1 U3772 ( .A1(n2269), .A2(n2277), .ZN(n3685) );
  INV_X1 U3773 ( .A(b_13_), .ZN(n2277) );
  INV_X1 U3774 ( .A(a_13_), .ZN(n2269) );
  AND2_X1 U3775 ( .A1(n3648), .A2(n2489), .ZN(n3684) );
  INV_X1 U3776 ( .A(n2406), .ZN(n2489) );
  AND2_X1 U3777 ( .A1(b_13_), .A2(a_13_), .ZN(n2406) );
  INV_X1 U3778 ( .A(n3646), .ZN(n3648) );
  OR2_X1 U3779 ( .A1(n3686), .A2(n2276), .ZN(n3646) );
  AND2_X1 U3780 ( .A1(a_14_), .A2(b_14_), .ZN(n2276) );
  AND2_X1 U3781 ( .A1(Result_mul_31_), .A2(n3687), .ZN(n3686) );
  OR2_X1 U3782 ( .A1(a_14_), .A2(b_14_), .ZN(n3687) );
  AND2_X1 U3783 ( .A1(a_15_), .A2(b_15_), .ZN(Result_mul_31_) );
endmodule

