module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n317_, new_n344_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n701_, new_n792_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n785_, new_n477_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n939_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n918_, new_n810_, new_n808_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n302_, new_n191_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n856_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n865_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n573_, new_n405_;

not g000 ( new_n151_, N75 );
nand g001 ( new_n152_, N29, N42 );
nor g002 ( N388, new_n152_, new_n151_ );
not g003 ( new_n154_, N80 );
nand g004 ( new_n155_, N29, N36 );
nor g005 ( N389, new_n155_, new_n154_ );
not g006 ( new_n157_, N42 );
nor g007 ( N390, new_n155_, new_n157_ );
nand g008 ( new_n159_, N85, N86 );
not g009 ( N391, new_n159_ );
not g010 ( new_n161_, N17 );
nand g011 ( new_n162_, N1, N8 );
not g012 ( new_n163_, new_n162_ );
nand g013 ( new_n164_, new_n163_, N13 );
nor g014 ( N418, new_n164_, new_n161_ );
not g015 ( new_n166_, N390 );
nand g016 ( new_n167_, N1, N26 );
nand g017 ( new_n168_, N13, N17 );
nor g018 ( new_n169_, new_n167_, new_n168_ );
nand g019 ( N419, new_n166_, new_n169_ );
nand g020 ( new_n171_, N59, N75 );
not g021 ( new_n172_, new_n171_ );
nand g022 ( N420, new_n172_, N80 );
nand g023 ( new_n174_, N36, N59 );
not g024 ( new_n175_, new_n174_ );
nand g025 ( N421, new_n175_, N80 );
nand g026 ( N422, new_n175_, N42 );
not g027 ( new_n178_, N90 );
nor g028 ( new_n179_, N87, N88 );
nor g029 ( N423, new_n179_, new_n178_ );
nand g030 ( N446, new_n169_, N390 );
not g031 ( new_n182_, N51 );
nor g032 ( new_n183_, new_n167_, new_n182_ );
nor g033 ( new_n184_, new_n183_, keyIn_0_0 );
not g034 ( new_n185_, keyIn_0_0 );
not g035 ( new_n186_, new_n167_ );
nand g036 ( new_n187_, new_n186_, N51 );
nor g037 ( new_n188_, new_n187_, new_n185_ );
nor g038 ( N447, new_n188_, new_n184_ );
not g039 ( new_n190_, new_n164_ );
nand g040 ( new_n191_, new_n190_, N55 );
nand g041 ( new_n192_, N29, N68 );
nor g042 ( N448, new_n191_, new_n192_ );
nand g043 ( new_n194_, N59, N68 );
not g044 ( new_n195_, new_n194_ );
nand g045 ( new_n196_, new_n195_, N74 );
nor g046 ( N449, new_n191_, new_n196_ );
not g047 ( new_n198_, N89 );
nor g048 ( N450, new_n179_, new_n198_ );
not g049 ( new_n200_, N135 );
nand g050 ( new_n201_, N111, N116 );
not g051 ( new_n202_, new_n201_ );
nor g052 ( new_n203_, N111, N116 );
nor g053 ( new_n204_, new_n202_, new_n203_ );
nand g054 ( new_n205_, N121, N126 );
not g055 ( new_n206_, new_n205_ );
nor g056 ( new_n207_, N121, N126 );
nor g057 ( new_n208_, new_n206_, new_n207_ );
nor g058 ( new_n209_, new_n204_, new_n208_ );
nand g059 ( new_n210_, new_n204_, new_n208_ );
not g060 ( new_n211_, new_n210_ );
nor g061 ( new_n212_, new_n211_, new_n209_ );
not g062 ( new_n213_, new_n212_ );
nand g063 ( new_n214_, new_n213_, new_n200_ );
nand g064 ( new_n215_, new_n214_, keyIn_0_21 );
not g065 ( new_n216_, new_n215_ );
nor g066 ( new_n217_, new_n214_, keyIn_0_21 );
nor g067 ( new_n218_, new_n216_, new_n217_ );
nor g068 ( new_n219_, new_n213_, new_n200_ );
nor g069 ( new_n220_, new_n218_, new_n219_ );
not g070 ( new_n221_, new_n220_ );
nand g071 ( new_n222_, N91, N96 );
not g072 ( new_n223_, new_n222_ );
nor g073 ( new_n224_, N91, N96 );
nor g074 ( new_n225_, new_n223_, new_n224_ );
nand g075 ( new_n226_, N101, N106 );
not g076 ( new_n227_, new_n226_ );
nor g077 ( new_n228_, N101, N106 );
nor g078 ( new_n229_, new_n227_, new_n228_ );
nor g079 ( new_n230_, new_n225_, new_n229_ );
nand g080 ( new_n231_, new_n225_, new_n229_ );
not g081 ( new_n232_, new_n231_ );
nor g082 ( new_n233_, new_n232_, new_n230_ );
not g083 ( new_n234_, new_n233_ );
nand g084 ( new_n235_, new_n234_, N130 );
not g085 ( new_n236_, new_n235_ );
nor g086 ( new_n237_, new_n234_, N130 );
nor g087 ( new_n238_, new_n236_, new_n237_ );
not g088 ( new_n239_, new_n238_ );
nand g089 ( new_n240_, new_n221_, new_n239_ );
nand g090 ( new_n241_, new_n220_, new_n238_ );
nand g091 ( N767, new_n240_, new_n241_ );
not g092 ( new_n243_, N207 );
nand g093 ( new_n244_, N195, N201 );
not g094 ( new_n245_, new_n244_ );
nor g095 ( new_n246_, N195, N201 );
nor g096 ( new_n247_, new_n245_, new_n246_ );
nand g097 ( new_n248_, keyIn_0_6, N183 );
nor g098 ( new_n249_, new_n247_, new_n248_ );
nand g099 ( new_n250_, new_n247_, new_n248_ );
not g100 ( new_n251_, new_n250_ );
nor g101 ( new_n252_, new_n251_, new_n249_ );
not g102 ( new_n253_, N189 );
nor g103 ( new_n254_, keyIn_0_6, N183 );
nor g104 ( new_n255_, new_n254_, new_n253_ );
not g105 ( new_n256_, new_n255_ );
nor g106 ( new_n257_, new_n252_, new_n256_ );
nand g107 ( new_n258_, new_n252_, new_n256_ );
not g108 ( new_n259_, new_n258_ );
nor g109 ( new_n260_, new_n259_, new_n257_ );
nor g110 ( new_n261_, new_n260_, new_n243_ );
nand g111 ( new_n262_, new_n260_, new_n243_ );
not g112 ( new_n263_, new_n262_ );
nor g113 ( new_n264_, new_n263_, new_n261_ );
not g114 ( new_n265_, new_n264_ );
not g115 ( new_n266_, N130 );
not g116 ( new_n267_, N159 );
nor g117 ( new_n268_, new_n267_, N165 );
not g118 ( new_n269_, N165 );
nor g119 ( new_n270_, new_n269_, N159 );
nor g120 ( new_n271_, new_n268_, new_n270_ );
nand g121 ( new_n272_, N171, N177 );
not g122 ( new_n273_, new_n272_ );
nor g123 ( new_n274_, N171, N177 );
nor g124 ( new_n275_, new_n273_, new_n274_ );
nor g125 ( new_n276_, new_n271_, new_n275_ );
nand g126 ( new_n277_, new_n271_, new_n275_ );
not g127 ( new_n278_, new_n277_ );
nor g128 ( new_n279_, new_n278_, new_n276_ );
nor g129 ( new_n280_, new_n279_, new_n266_ );
nand g130 ( new_n281_, new_n279_, new_n266_ );
not g131 ( new_n282_, new_n281_ );
nor g132 ( new_n283_, new_n282_, new_n280_ );
not g133 ( new_n284_, new_n283_ );
nand g134 ( new_n285_, new_n265_, new_n284_ );
nand g135 ( new_n286_, new_n264_, new_n283_ );
nand g136 ( N768, new_n285_, new_n286_ );
not g137 ( new_n288_, N201 );
not g138 ( new_n289_, keyIn_0_16 );
not g139 ( new_n290_, keyIn_0_12 );
nand g140 ( new_n291_, new_n187_, new_n185_ );
nand g141 ( new_n292_, new_n183_, keyIn_0_0 );
nand g142 ( new_n293_, new_n291_, new_n292_ );
nand g143 ( new_n294_, new_n293_, keyIn_0_8 );
not g144 ( new_n295_, keyIn_0_8 );
nand g145 ( new_n296_, N447, new_n295_ );
nand g146 ( new_n297_, new_n296_, new_n294_ );
nand g147 ( new_n298_, new_n297_, new_n290_ );
nor g148 ( new_n299_, N447, new_n295_ );
nor g149 ( new_n300_, new_n293_, keyIn_0_8 );
nor g150 ( new_n301_, new_n299_, new_n300_ );
nand g151 ( new_n302_, new_n301_, keyIn_0_12 );
nand g152 ( new_n303_, new_n302_, new_n298_ );
not g153 ( new_n304_, keyIn_0_3 );
nand g154 ( new_n305_, N59, N156 );
nand g155 ( new_n306_, new_n305_, new_n304_ );
not g156 ( new_n307_, new_n306_ );
nor g157 ( new_n308_, new_n305_, new_n304_ );
nor g158 ( new_n309_, new_n307_, new_n308_ );
nor g159 ( new_n310_, new_n309_, new_n161_ );
nand g160 ( new_n311_, new_n303_, new_n310_ );
nor g161 ( new_n312_, new_n311_, new_n289_ );
not g162 ( new_n313_, new_n312_ );
nand g163 ( new_n314_, new_n311_, new_n289_ );
nand g164 ( new_n315_, new_n314_, N1 );
not g165 ( new_n316_, new_n315_ );
nand g166 ( new_n317_, new_n316_, new_n313_ );
nand g167 ( new_n318_, new_n317_, keyIn_0_18 );
not g168 ( new_n319_, keyIn_0_18 );
nor g169 ( new_n320_, new_n315_, new_n312_ );
nand g170 ( new_n321_, new_n320_, new_n319_ );
nand g171 ( new_n322_, new_n318_, new_n321_ );
nand g172 ( new_n323_, new_n322_, N153 );
nor g173 ( new_n324_, N17, N42 );
nor g174 ( new_n325_, new_n324_, keyIn_0_4 );
not g175 ( new_n326_, keyIn_0_5 );
nand g176 ( new_n327_, N17, N42 );
nand g177 ( new_n328_, new_n327_, new_n326_ );
not g178 ( new_n329_, new_n328_ );
nor g179 ( new_n330_, new_n329_, new_n325_ );
nand g180 ( new_n331_, keyIn_0_5, N17 );
nor g181 ( new_n332_, new_n331_, new_n157_ );
nand g182 ( new_n333_, new_n324_, keyIn_0_4 );
not g183 ( new_n334_, new_n333_ );
nor g184 ( new_n335_, new_n334_, new_n332_ );
nand g185 ( new_n336_, new_n335_, new_n330_ );
nor g186 ( new_n337_, new_n336_, keyIn_0_11 );
not g187 ( new_n338_, new_n305_ );
nand g188 ( new_n339_, new_n336_, keyIn_0_11 );
nand g189 ( new_n340_, new_n339_, new_n338_ );
nor g190 ( new_n341_, new_n340_, new_n337_ );
nand g191 ( new_n342_, new_n303_, new_n341_ );
nand g192 ( new_n343_, new_n342_, keyIn_0_15 );
nor g193 ( new_n344_, new_n342_, keyIn_0_15 );
not g194 ( new_n345_, new_n344_ );
nand g195 ( new_n346_, new_n345_, new_n343_ );
not g196 ( new_n347_, keyIn_0_13 );
not g197 ( new_n348_, keyIn_0_10 );
not g198 ( new_n349_, keyIn_0_2 );
nand g199 ( new_n350_, N42, N59 );
nor g200 ( new_n351_, new_n350_, new_n151_ );
nor g201 ( new_n352_, new_n351_, new_n349_ );
nand g202 ( new_n353_, new_n351_, new_n349_ );
not g203 ( new_n354_, new_n353_ );
nor g204 ( new_n355_, new_n354_, new_n352_ );
nor g205 ( new_n356_, new_n355_, new_n348_ );
nand g206 ( new_n357_, new_n355_, new_n348_ );
not g207 ( new_n358_, new_n357_ );
nor g208 ( new_n359_, new_n358_, new_n356_ );
not g209 ( new_n360_, new_n359_ );
not g210 ( new_n361_, keyIn_0_9 );
nand g211 ( new_n362_, N17, N51 );
nor g212 ( new_n363_, new_n162_, new_n362_ );
nor g213 ( new_n364_, new_n363_, keyIn_0_1 );
nand g214 ( new_n365_, new_n363_, keyIn_0_1 );
not g215 ( new_n366_, new_n365_ );
nor g216 ( new_n367_, new_n366_, new_n364_ );
nor g217 ( new_n368_, new_n367_, new_n361_ );
nand g218 ( new_n369_, new_n367_, new_n361_ );
not g219 ( new_n370_, new_n369_ );
nor g220 ( new_n371_, new_n370_, new_n368_ );
nand g221 ( new_n372_, new_n360_, new_n371_ );
nand g222 ( new_n373_, new_n372_, new_n347_ );
nor g223 ( new_n374_, new_n372_, new_n347_ );
not g224 ( new_n375_, new_n374_ );
nand g225 ( new_n376_, new_n375_, new_n373_ );
nand g226 ( new_n377_, new_n346_, new_n376_ );
nand g227 ( new_n378_, new_n377_, keyIn_0_17 );
not g228 ( new_n379_, keyIn_0_17 );
not g229 ( new_n380_, new_n343_ );
nor g230 ( new_n381_, new_n380_, new_n344_ );
not g231 ( new_n382_, new_n373_ );
nor g232 ( new_n383_, new_n382_, new_n374_ );
nor g233 ( new_n384_, new_n381_, new_n383_ );
nand g234 ( new_n385_, new_n384_, new_n379_ );
nand g235 ( new_n386_, new_n385_, new_n378_ );
nand g236 ( new_n387_, new_n386_, N126 );
nand g237 ( new_n388_, new_n387_, new_n323_ );
nand g238 ( new_n389_, new_n388_, keyIn_0_27 );
not g239 ( new_n390_, new_n389_ );
nor g240 ( new_n391_, new_n388_, keyIn_0_27 );
nor g241 ( new_n392_, new_n390_, new_n391_ );
not g242 ( new_n393_, N55 );
nand g243 ( new_n394_, N29, N75 );
nor g244 ( new_n395_, new_n394_, new_n154_ );
nand g245 ( new_n396_, new_n303_, new_n395_ );
nor g246 ( new_n397_, new_n396_, new_n393_ );
nor g247 ( new_n398_, new_n397_, keyIn_0_14 );
nand g248 ( new_n399_, new_n397_, keyIn_0_14 );
not g249 ( new_n400_, new_n399_ );
nor g250 ( new_n401_, new_n400_, new_n398_ );
nor g251 ( new_n402_, new_n401_, N268 );
nor g252 ( new_n403_, new_n392_, new_n402_ );
nor g253 ( new_n404_, new_n403_, keyIn_0_30 );
not g254 ( new_n405_, new_n404_ );
nand g255 ( new_n406_, new_n403_, keyIn_0_30 );
nand g256 ( new_n407_, new_n405_, new_n406_ );
nor g257 ( new_n408_, new_n407_, new_n288_ );
not g258 ( new_n409_, keyIn_0_35 );
nand g259 ( new_n410_, new_n407_, new_n288_ );
nand g260 ( new_n411_, new_n410_, new_n409_ );
not g261 ( new_n412_, new_n410_ );
nand g262 ( new_n413_, new_n412_, keyIn_0_35 );
nand g263 ( new_n414_, new_n413_, new_n411_ );
nor g264 ( new_n415_, new_n414_, new_n408_ );
nand g265 ( new_n416_, new_n415_, N261 );
not g266 ( new_n417_, N219 );
nor g267 ( new_n418_, new_n415_, N261 );
nor g268 ( new_n419_, new_n418_, new_n417_ );
nand g269 ( new_n420_, new_n419_, new_n416_ );
not g270 ( new_n421_, N228 );
not g271 ( new_n422_, new_n415_ );
nor g272 ( new_n423_, new_n422_, new_n421_ );
nand g273 ( new_n424_, new_n408_, N237 );
not g274 ( new_n425_, N246 );
nor g275 ( new_n426_, new_n407_, new_n425_ );
not g276 ( new_n427_, N73 );
nand g277 ( new_n428_, N42, N72 );
nor g278 ( new_n429_, new_n428_, new_n427_ );
nand g279 ( new_n430_, new_n429_, new_n195_ );
nor g280 ( new_n431_, new_n191_, new_n430_ );
nand g281 ( new_n432_, new_n431_, N201 );
not g282 ( new_n433_, keyIn_0_7 );
nand g283 ( new_n434_, N121, N210 );
nor g284 ( new_n435_, new_n434_, new_n433_ );
nand g285 ( new_n436_, N255, N267 );
nand g286 ( new_n437_, new_n434_, new_n433_ );
nand g287 ( new_n438_, new_n437_, new_n436_ );
nor g288 ( new_n439_, new_n438_, new_n435_ );
nand g289 ( new_n440_, new_n432_, new_n439_ );
nor g290 ( new_n441_, new_n426_, new_n440_ );
nand g291 ( new_n442_, new_n441_, new_n424_ );
nor g292 ( new_n443_, new_n423_, new_n442_ );
nand g293 ( N850, new_n420_, new_n443_ );
not g294 ( new_n445_, keyIn_0_38 );
not g295 ( new_n446_, keyIn_0_32 );
not g296 ( new_n447_, keyIn_0_25 );
nand g297 ( new_n448_, new_n322_, N146 );
nand g298 ( new_n449_, new_n448_, keyIn_0_22 );
nor g299 ( new_n450_, new_n448_, keyIn_0_22 );
not g300 ( new_n451_, new_n450_ );
nand g301 ( new_n452_, new_n451_, new_n449_ );
not g302 ( new_n453_, keyIn_0_23 );
nand g303 ( new_n454_, new_n386_, N116 );
nor g304 ( new_n455_, new_n454_, new_n453_ );
nand g305 ( new_n456_, new_n454_, new_n453_ );
not g306 ( new_n457_, new_n456_ );
nor g307 ( new_n458_, new_n457_, new_n455_ );
nand g308 ( new_n459_, new_n458_, new_n452_ );
nand g309 ( new_n460_, new_n459_, new_n447_ );
not g310 ( new_n461_, new_n449_ );
nor g311 ( new_n462_, new_n461_, new_n450_ );
not g312 ( new_n463_, new_n454_ );
nand g313 ( new_n464_, new_n463_, keyIn_0_23 );
nand g314 ( new_n465_, new_n464_, new_n456_ );
nor g315 ( new_n466_, new_n465_, new_n462_ );
nand g316 ( new_n467_, new_n466_, keyIn_0_25 );
nand g317 ( new_n468_, new_n460_, new_n467_ );
not g318 ( new_n469_, keyIn_0_20 );
not g319 ( new_n470_, new_n402_ );
nand g320 ( new_n471_, new_n470_, new_n469_ );
nand g321 ( new_n472_, new_n402_, keyIn_0_20 );
nand g322 ( new_n473_, new_n471_, new_n472_ );
nand g323 ( new_n474_, new_n468_, new_n473_ );
nand g324 ( new_n475_, new_n474_, keyIn_0_28 );
not g325 ( new_n476_, keyIn_0_28 );
not g326 ( new_n477_, new_n474_ );
nand g327 ( new_n478_, new_n477_, new_n476_ );
nand g328 ( new_n479_, new_n478_, new_n475_ );
nand g329 ( new_n480_, new_n479_, new_n253_ );
nand g330 ( new_n481_, new_n480_, new_n446_ );
not g331 ( new_n482_, new_n481_ );
nor g332 ( new_n483_, new_n480_, new_n446_ );
nor g333 ( new_n484_, new_n482_, new_n483_ );
not g334 ( new_n485_, keyIn_0_34 );
not g335 ( new_n486_, N195 );
not g336 ( new_n487_, keyIn_0_29 );
not g337 ( new_n488_, keyIn_0_26 );
not g338 ( new_n489_, keyIn_0_24 );
nand g339 ( new_n490_, new_n386_, N121 );
nor g340 ( new_n491_, new_n490_, new_n489_ );
nand g341 ( new_n492_, new_n322_, N149 );
nand g342 ( new_n493_, new_n490_, new_n489_ );
nand g343 ( new_n494_, new_n493_, new_n492_ );
nor g344 ( new_n495_, new_n494_, new_n491_ );
nand g345 ( new_n496_, new_n495_, new_n488_ );
nor g346 ( new_n497_, new_n495_, new_n488_ );
nor g347 ( new_n498_, new_n497_, new_n402_ );
nand g348 ( new_n499_, new_n498_, new_n496_ );
nand g349 ( new_n500_, new_n499_, new_n487_ );
not g350 ( new_n501_, new_n496_ );
not g351 ( new_n502_, new_n491_ );
not g352 ( new_n503_, new_n494_ );
nand g353 ( new_n504_, new_n503_, new_n502_ );
nand g354 ( new_n505_, new_n504_, keyIn_0_26 );
nand g355 ( new_n506_, new_n505_, new_n470_ );
nor g356 ( new_n507_, new_n506_, new_n501_ );
nand g357 ( new_n508_, new_n507_, keyIn_0_29 );
nand g358 ( new_n509_, new_n508_, new_n500_ );
nand g359 ( new_n510_, new_n509_, new_n486_ );
nand g360 ( new_n511_, new_n510_, new_n485_ );
nor g361 ( new_n512_, new_n507_, keyIn_0_29 );
nor g362 ( new_n513_, new_n499_, new_n487_ );
nor g363 ( new_n514_, new_n512_, new_n513_ );
nor g364 ( new_n515_, new_n514_, N195 );
nand g365 ( new_n516_, new_n515_, keyIn_0_34 );
nand g366 ( new_n517_, new_n516_, new_n511_ );
not g367 ( new_n518_, N261 );
nor g368 ( new_n519_, new_n414_, new_n518_ );
nand g369 ( new_n520_, new_n519_, new_n517_ );
nor g370 ( new_n521_, new_n520_, new_n484_ );
nor g371 ( new_n522_, new_n521_, new_n445_ );
not g372 ( new_n523_, new_n522_ );
nand g373 ( new_n524_, new_n521_, new_n445_ );
nand g374 ( new_n525_, new_n523_, new_n524_ );
not g375 ( new_n526_, keyIn_0_39 );
not g376 ( new_n527_, keyIn_0_36 );
not g377 ( new_n528_, new_n475_ );
nor g378 ( new_n529_, new_n474_, keyIn_0_28 );
nor g379 ( new_n530_, new_n528_, new_n529_ );
nand g380 ( new_n531_, new_n530_, N189 );
nand g381 ( new_n532_, new_n531_, keyIn_0_31 );
not g382 ( new_n533_, keyIn_0_31 );
nor g383 ( new_n534_, new_n479_, new_n253_ );
nand g384 ( new_n535_, new_n534_, new_n533_ );
nand g385 ( new_n536_, new_n532_, new_n535_ );
nand g386 ( new_n537_, new_n536_, new_n527_ );
not g387 ( new_n538_, new_n536_ );
nand g388 ( new_n539_, new_n538_, keyIn_0_36 );
nand g389 ( new_n540_, new_n539_, new_n537_ );
nand g390 ( new_n541_, new_n540_, new_n526_ );
not g391 ( new_n542_, new_n537_ );
nor g392 ( new_n543_, new_n536_, new_n527_ );
nor g393 ( new_n544_, new_n542_, new_n543_ );
nand g394 ( new_n545_, new_n544_, keyIn_0_39 );
nand g395 ( new_n546_, new_n545_, new_n541_ );
nor g396 ( new_n547_, new_n525_, new_n546_ );
not g397 ( new_n548_, keyIn_0_40 );
not g398 ( new_n549_, new_n483_ );
nand g399 ( new_n550_, new_n549_, new_n481_ );
not g400 ( new_n551_, keyIn_0_33 );
nand g401 ( new_n552_, new_n514_, N195 );
nand g402 ( new_n553_, new_n552_, new_n551_ );
nor g403 ( new_n554_, new_n509_, new_n486_ );
nand g404 ( new_n555_, new_n554_, keyIn_0_33 );
nand g405 ( new_n556_, new_n553_, new_n555_ );
nand g406 ( new_n557_, new_n556_, keyIn_0_37 );
not g407 ( new_n558_, new_n557_ );
nor g408 ( new_n559_, new_n556_, keyIn_0_37 );
nor g409 ( new_n560_, new_n558_, new_n559_ );
nand g410 ( new_n561_, new_n560_, new_n550_ );
nor g411 ( new_n562_, new_n561_, new_n548_ );
nand g412 ( new_n563_, new_n561_, new_n548_ );
nand g413 ( new_n564_, new_n517_, new_n408_ );
nor g414 ( new_n565_, new_n484_, new_n564_ );
nor g415 ( new_n566_, new_n565_, keyIn_0_41 );
not g416 ( new_n567_, keyIn_0_41 );
not g417 ( new_n568_, new_n408_ );
not g418 ( new_n569_, new_n511_ );
nor g419 ( new_n570_, new_n510_, new_n485_ );
nor g420 ( new_n571_, new_n569_, new_n570_ );
nor g421 ( new_n572_, new_n571_, new_n568_ );
nand g422 ( new_n573_, new_n572_, new_n550_ );
nor g423 ( new_n574_, new_n573_, new_n567_ );
nor g424 ( new_n575_, new_n574_, new_n566_ );
nand g425 ( new_n576_, new_n575_, new_n563_ );
nor g426 ( new_n577_, new_n576_, new_n562_ );
nand g427 ( new_n578_, new_n577_, new_n547_ );
nand g428 ( new_n579_, new_n578_, keyIn_0_42 );
not g429 ( new_n580_, keyIn_0_42 );
not g430 ( new_n581_, new_n524_ );
nor g431 ( new_n582_, new_n581_, new_n522_ );
nor g432 ( new_n583_, new_n544_, keyIn_0_39 );
nor g433 ( new_n584_, new_n540_, new_n526_ );
nor g434 ( new_n585_, new_n583_, new_n584_ );
nand g435 ( new_n586_, new_n585_, new_n582_ );
not g436 ( new_n587_, new_n562_ );
not g437 ( new_n588_, keyIn_0_37 );
nor g438 ( new_n589_, new_n554_, keyIn_0_33 );
nor g439 ( new_n590_, new_n552_, new_n551_ );
nor g440 ( new_n591_, new_n590_, new_n589_ );
nand g441 ( new_n592_, new_n591_, new_n588_ );
nand g442 ( new_n593_, new_n592_, new_n557_ );
nor g443 ( new_n594_, new_n593_, new_n484_ );
nor g444 ( new_n595_, new_n594_, keyIn_0_40 );
nand g445 ( new_n596_, new_n573_, new_n567_ );
nand g446 ( new_n597_, new_n565_, keyIn_0_41 );
nand g447 ( new_n598_, new_n596_, new_n597_ );
nor g448 ( new_n599_, new_n595_, new_n598_ );
nand g449 ( new_n600_, new_n599_, new_n587_ );
nor g450 ( new_n601_, new_n586_, new_n600_ );
nand g451 ( new_n602_, new_n601_, new_n580_ );
nand g452 ( new_n603_, new_n602_, new_n579_ );
not g453 ( new_n604_, N183 );
not g454 ( new_n605_, N143 );
not g455 ( new_n606_, new_n322_ );
nor g456 ( new_n607_, new_n606_, new_n605_ );
nand g457 ( new_n608_, new_n386_, N111 );
not g458 ( new_n609_, new_n608_ );
not g459 ( new_n610_, keyIn_0_19 );
nand g460 ( new_n611_, new_n470_, new_n610_ );
not g461 ( new_n612_, new_n611_ );
nor g462 ( new_n613_, new_n470_, new_n610_ );
nor g463 ( new_n614_, new_n612_, new_n613_ );
nor g464 ( new_n615_, new_n614_, new_n609_ );
not g465 ( new_n616_, new_n615_ );
nor g466 ( new_n617_, new_n616_, new_n607_ );
nor g467 ( new_n618_, new_n617_, new_n604_ );
not g468 ( new_n619_, new_n618_ );
nand g469 ( new_n620_, new_n617_, new_n604_ );
nand g470 ( new_n621_, new_n619_, new_n620_ );
not g471 ( new_n622_, new_n621_ );
nand g472 ( new_n623_, new_n603_, new_n622_ );
nor g473 ( new_n624_, new_n603_, new_n622_ );
nor g474 ( new_n625_, new_n624_, new_n417_ );
nand g475 ( new_n626_, new_n625_, new_n623_ );
nor g476 ( new_n627_, new_n621_, new_n421_ );
nand g477 ( new_n628_, new_n618_, N237 );
nor g478 ( new_n629_, new_n617_, new_n425_ );
nand g479 ( new_n630_, new_n431_, N183 );
nand g480 ( new_n631_, N106, N210 );
nand g481 ( new_n632_, new_n630_, new_n631_ );
nor g482 ( new_n633_, new_n629_, new_n632_ );
nand g483 ( new_n634_, new_n633_, new_n628_ );
nor g484 ( new_n635_, new_n627_, new_n634_ );
nand g485 ( N863, new_n626_, new_n635_ );
not g486 ( new_n637_, keyIn_0_50 );
nor g487 ( new_n638_, new_n484_, new_n536_ );
nor g488 ( new_n639_, new_n519_, new_n408_ );
nor g489 ( new_n640_, new_n639_, new_n571_ );
nor g490 ( new_n641_, new_n640_, new_n560_ );
not g491 ( new_n642_, new_n641_ );
nor g492 ( new_n643_, new_n642_, new_n638_ );
nand g493 ( new_n644_, new_n642_, new_n638_ );
nand g494 ( new_n645_, new_n644_, N219 );
nor g495 ( new_n646_, new_n645_, new_n643_ );
nand g496 ( new_n647_, N111, N210 );
not g497 ( new_n648_, new_n647_ );
nor g498 ( new_n649_, new_n646_, new_n648_ );
not g499 ( new_n650_, new_n649_ );
nand g500 ( new_n651_, new_n650_, new_n637_ );
nand g501 ( new_n652_, new_n649_, keyIn_0_50 );
nand g502 ( new_n653_, new_n651_, new_n652_ );
not g503 ( new_n654_, N237 );
nor g504 ( new_n655_, new_n540_, new_n654_ );
nand g505 ( new_n656_, new_n638_, N228 );
nor g506 ( new_n657_, new_n479_, new_n425_ );
nand g507 ( new_n658_, new_n431_, N189 );
nand g508 ( new_n659_, N255, N259 );
nand g509 ( new_n660_, new_n658_, new_n659_ );
nor g510 ( new_n661_, new_n657_, new_n660_ );
nand g511 ( new_n662_, new_n656_, new_n661_ );
nor g512 ( new_n663_, new_n655_, new_n662_ );
nand g513 ( N864, new_n653_, new_n663_ );
nor g514 ( new_n665_, new_n571_, new_n591_ );
not g515 ( new_n666_, new_n665_ );
nand g516 ( new_n667_, new_n666_, new_n639_ );
nor g517 ( new_n668_, new_n666_, new_n639_ );
nor g518 ( new_n669_, new_n668_, new_n417_ );
nand g519 ( new_n670_, new_n669_, new_n667_ );
nor g520 ( new_n671_, new_n593_, new_n654_ );
nand g521 ( new_n672_, new_n665_, N228 );
nor g522 ( new_n673_, new_n509_, new_n425_ );
nand g523 ( new_n674_, new_n431_, N195 );
nand g524 ( new_n675_, N255, N260 );
nand g525 ( new_n676_, N116, N210 );
nand g526 ( new_n677_, new_n675_, new_n676_ );
not g527 ( new_n678_, new_n677_ );
nand g528 ( new_n679_, new_n674_, new_n678_ );
nor g529 ( new_n680_, new_n673_, new_n679_ );
nand g530 ( new_n681_, new_n672_, new_n680_ );
nor g531 ( new_n682_, new_n681_, new_n671_ );
nand g532 ( N865, new_n670_, new_n682_ );
not g533 ( new_n684_, keyIn_0_48 );
nand g534 ( new_n685_, new_n603_, new_n620_ );
nand g535 ( new_n686_, new_n685_, keyIn_0_43 );
not g536 ( new_n687_, new_n686_ );
nor g537 ( new_n688_, new_n685_, keyIn_0_43 );
nor g538 ( new_n689_, new_n687_, new_n688_ );
nor g539 ( new_n690_, new_n689_, new_n618_ );
nor g540 ( new_n691_, new_n690_, keyIn_0_44 );
not g541 ( new_n692_, keyIn_0_44 );
not g542 ( new_n693_, new_n688_ );
nand g543 ( new_n694_, new_n693_, new_n686_ );
nand g544 ( new_n695_, new_n694_, new_n619_ );
nor g545 ( new_n696_, new_n695_, new_n692_ );
nor g546 ( new_n697_, new_n691_, new_n696_ );
nand g547 ( new_n698_, new_n386_, N96 );
not g548 ( new_n699_, N146 );
nor g549 ( new_n700_, new_n309_, new_n393_ );
nand g550 ( new_n701_, new_n303_, new_n700_ );
nor g551 ( new_n702_, new_n701_, new_n699_ );
nand g552 ( new_n703_, N51, N138 );
not g553 ( new_n704_, new_n396_ );
nor g554 ( new_n705_, new_n161_, N268 );
nand g555 ( new_n706_, new_n704_, new_n705_ );
nand g556 ( new_n707_, new_n706_, new_n703_ );
nor g557 ( new_n708_, new_n707_, new_n702_ );
nand g558 ( new_n709_, new_n698_, new_n708_ );
nor g559 ( new_n710_, new_n709_, N165 );
nand g560 ( new_n711_, new_n386_, N101 );
not g561 ( new_n712_, N149 );
nor g562 ( new_n713_, new_n701_, new_n712_ );
nand g563 ( new_n714_, N17, N138 );
nand g564 ( new_n715_, new_n706_, new_n714_ );
nor g565 ( new_n716_, new_n715_, new_n713_ );
nand g566 ( new_n717_, new_n711_, new_n716_ );
nor g567 ( new_n718_, new_n717_, N171 );
nor g568 ( new_n719_, new_n710_, new_n718_ );
nand g569 ( new_n720_, new_n386_, N106 );
not g570 ( new_n721_, N153 );
nor g571 ( new_n722_, new_n701_, new_n721_ );
nand g572 ( new_n723_, N138, N152 );
nand g573 ( new_n724_, new_n706_, new_n723_ );
nor g574 ( new_n725_, new_n724_, new_n722_ );
nand g575 ( new_n726_, new_n720_, new_n725_ );
nor g576 ( new_n727_, new_n726_, N177 );
not g577 ( new_n728_, new_n727_ );
nand g578 ( new_n729_, new_n719_, new_n728_ );
not g579 ( new_n730_, new_n729_ );
nand g580 ( new_n731_, new_n697_, new_n730_ );
nor g581 ( new_n732_, new_n731_, keyIn_0_47 );
not g582 ( new_n733_, new_n732_ );
not g583 ( new_n734_, keyIn_0_47 );
nand g584 ( new_n735_, new_n695_, new_n692_ );
nand g585 ( new_n736_, new_n690_, keyIn_0_44 );
nand g586 ( new_n737_, new_n736_, new_n735_ );
nor g587 ( new_n738_, new_n737_, new_n729_ );
nor g588 ( new_n739_, new_n738_, new_n734_ );
nand g589 ( new_n740_, new_n717_, N171 );
nand g590 ( new_n741_, new_n726_, N177 );
nand g591 ( new_n742_, new_n740_, new_n741_ );
nand g592 ( new_n743_, new_n719_, new_n742_ );
nand g593 ( new_n744_, new_n709_, N165 );
nand g594 ( new_n745_, new_n743_, new_n744_ );
nor g595 ( new_n746_, new_n739_, new_n745_ );
nand g596 ( new_n747_, new_n746_, new_n733_ );
nand g597 ( new_n748_, new_n747_, new_n684_ );
nand g598 ( new_n749_, new_n731_, keyIn_0_47 );
not g599 ( new_n750_, new_n745_ );
nand g600 ( new_n751_, new_n749_, new_n750_ );
nor g601 ( new_n752_, new_n751_, new_n732_ );
nand g602 ( new_n753_, new_n752_, keyIn_0_48 );
nand g603 ( new_n754_, new_n748_, new_n753_ );
nand g604 ( new_n755_, new_n386_, N91 );
nor g605 ( new_n756_, new_n701_, new_n605_ );
nand g606 ( new_n757_, N8, N138 );
nand g607 ( new_n758_, new_n706_, new_n757_ );
nor g608 ( new_n759_, new_n758_, new_n756_ );
nand g609 ( new_n760_, new_n755_, new_n759_ );
nor g610 ( new_n761_, new_n760_, N159 );
not g611 ( new_n762_, new_n761_ );
nand g612 ( new_n763_, new_n754_, new_n762_ );
nand g613 ( new_n764_, new_n760_, N159 );
nand g614 ( N866, new_n763_, new_n764_ );
not g615 ( new_n766_, keyIn_0_57 );
not g616 ( new_n767_, keyIn_0_53 );
not g617 ( new_n768_, keyIn_0_49 );
not g618 ( new_n769_, new_n741_ );
nor g619 ( new_n770_, new_n769_, new_n727_ );
not g620 ( new_n771_, new_n770_ );
nor g621 ( new_n772_, new_n737_, new_n771_ );
nor g622 ( new_n773_, new_n772_, keyIn_0_46 );
nand g623 ( new_n774_, new_n772_, keyIn_0_46 );
not g624 ( new_n775_, new_n774_ );
nor g625 ( new_n776_, new_n775_, new_n773_ );
not g626 ( new_n777_, keyIn_0_45 );
nor g627 ( new_n778_, new_n697_, new_n770_ );
not g628 ( new_n779_, new_n778_ );
nand g629 ( new_n780_, new_n779_, new_n777_ );
not g630 ( new_n781_, new_n780_ );
nor g631 ( new_n782_, new_n779_, new_n777_ );
nor g632 ( new_n783_, new_n781_, new_n782_ );
nor g633 ( new_n784_, new_n783_, new_n776_ );
not g634 ( new_n785_, new_n784_ );
nand g635 ( new_n786_, new_n785_, new_n768_ );
nor g636 ( new_n787_, new_n785_, new_n768_ );
nor g637 ( new_n788_, new_n787_, new_n417_ );
nand g638 ( new_n789_, new_n788_, new_n786_ );
not g639 ( new_n790_, new_n789_ );
nor g640 ( new_n791_, new_n790_, new_n767_ );
nor g641 ( new_n792_, new_n789_, keyIn_0_53 );
nor g642 ( new_n793_, new_n791_, new_n792_ );
not g643 ( new_n794_, new_n793_ );
nand g644 ( new_n795_, N101, N210 );
nand g645 ( new_n796_, new_n794_, new_n795_ );
nand g646 ( new_n797_, new_n796_, keyIn_0_55 );
not g647 ( new_n798_, new_n797_ );
nor g648 ( new_n799_, new_n796_, keyIn_0_55 );
nor g649 ( new_n800_, new_n798_, new_n799_ );
nor g650 ( new_n801_, new_n771_, new_n421_ );
nor g651 ( new_n802_, new_n741_, new_n654_ );
nand g652 ( new_n803_, new_n726_, N246 );
nand g653 ( new_n804_, new_n431_, N177 );
nand g654 ( new_n805_, new_n803_, new_n804_ );
nor g655 ( new_n806_, new_n802_, new_n805_ );
not g656 ( new_n807_, new_n806_ );
nor g657 ( new_n808_, new_n801_, new_n807_ );
not g658 ( new_n809_, new_n808_ );
nor g659 ( new_n810_, new_n800_, new_n809_ );
nor g660 ( new_n811_, new_n810_, new_n766_ );
nand g661 ( new_n812_, new_n810_, new_n766_ );
not g662 ( new_n813_, new_n812_ );
nor g663 ( new_n814_, new_n813_, new_n811_ );
not g664 ( new_n815_, new_n814_ );
nor g665 ( new_n816_, new_n815_, keyIn_0_59 );
not g666 ( new_n817_, new_n816_ );
nand g667 ( new_n818_, new_n815_, keyIn_0_59 );
nand g668 ( new_n819_, new_n817_, new_n818_ );
nand g669 ( new_n820_, new_n819_, keyIn_0_61 );
not g670 ( new_n821_, keyIn_0_61 );
not g671 ( new_n822_, new_n818_ );
nor g672 ( new_n823_, new_n822_, new_n816_ );
nand g673 ( new_n824_, new_n823_, new_n821_ );
nand g674 ( N874, new_n824_, new_n820_ );
not g675 ( new_n826_, keyIn_0_62 );
not g676 ( new_n827_, keyIn_0_54 );
not g677 ( new_n828_, keyIn_0_51 );
not g678 ( new_n829_, new_n764_ );
nor g679 ( new_n830_, new_n829_, new_n761_ );
nor g680 ( new_n831_, new_n754_, new_n830_ );
nor g681 ( new_n832_, new_n831_, new_n828_ );
nand g682 ( new_n833_, new_n754_, new_n830_ );
nand g683 ( new_n834_, new_n833_, keyIn_0_52 );
not g684 ( new_n835_, new_n834_ );
nor g685 ( new_n836_, new_n835_, new_n832_ );
nor g686 ( new_n837_, new_n833_, keyIn_0_52 );
nor g687 ( new_n838_, new_n752_, keyIn_0_48 );
nor g688 ( new_n839_, new_n747_, new_n684_ );
nor g689 ( new_n840_, new_n838_, new_n839_ );
not g690 ( new_n841_, new_n830_ );
nand g691 ( new_n842_, new_n840_, new_n841_ );
nor g692 ( new_n843_, new_n842_, keyIn_0_51 );
nor g693 ( new_n844_, new_n843_, new_n837_ );
nand g694 ( new_n845_, new_n844_, new_n836_ );
nand g695 ( new_n846_, new_n845_, new_n827_ );
nand g696 ( new_n847_, new_n842_, keyIn_0_51 );
nand g697 ( new_n848_, new_n847_, new_n834_ );
not g698 ( new_n849_, keyIn_0_52 );
not g699 ( new_n850_, new_n833_ );
nand g700 ( new_n851_, new_n850_, new_n849_ );
nand g701 ( new_n852_, new_n831_, new_n828_ );
nand g702 ( new_n853_, new_n851_, new_n852_ );
nor g703 ( new_n854_, new_n853_, new_n848_ );
nand g704 ( new_n855_, new_n854_, keyIn_0_54 );
nand g705 ( new_n856_, new_n846_, new_n855_ );
nand g706 ( new_n857_, new_n856_, N219 );
nand g707 ( new_n858_, new_n857_, keyIn_0_56 );
not g708 ( new_n859_, keyIn_0_56 );
not g709 ( new_n860_, new_n857_ );
nand g710 ( new_n861_, new_n860_, new_n859_ );
nand g711 ( new_n862_, new_n861_, new_n858_ );
nand g712 ( new_n863_, N210, N268 );
nand g713 ( new_n864_, new_n862_, new_n863_ );
nor g714 ( new_n865_, new_n864_, keyIn_0_58 );
not g715 ( new_n866_, new_n865_ );
nand g716 ( new_n867_, new_n864_, keyIn_0_58 );
nor g717 ( new_n868_, new_n841_, new_n421_ );
nand g718 ( new_n869_, new_n829_, N237 );
nand g719 ( new_n870_, new_n760_, N246 );
nand g720 ( new_n871_, new_n431_, N159 );
nand g721 ( new_n872_, new_n870_, new_n871_ );
not g722 ( new_n873_, new_n872_ );
nand g723 ( new_n874_, new_n869_, new_n873_ );
nor g724 ( new_n875_, new_n868_, new_n874_ );
nand g725 ( new_n876_, new_n867_, new_n875_ );
not g726 ( new_n877_, new_n876_ );
nand g727 ( new_n878_, new_n877_, new_n866_ );
nand g728 ( new_n879_, new_n878_, keyIn_0_60 );
not g729 ( new_n880_, keyIn_0_60 );
nor g730 ( new_n881_, new_n876_, new_n865_ );
nand g731 ( new_n882_, new_n881_, new_n880_ );
nand g732 ( new_n883_, new_n879_, new_n882_ );
nand g733 ( new_n884_, new_n883_, new_n826_ );
nor g734 ( new_n885_, new_n881_, new_n880_ );
nor g735 ( new_n886_, new_n878_, keyIn_0_60 );
nor g736 ( new_n887_, new_n886_, new_n885_ );
nand g737 ( new_n888_, new_n887_, keyIn_0_62 );
nand g738 ( new_n889_, new_n888_, new_n884_ );
nand g739 ( new_n890_, new_n889_, keyIn_0_63 );
not g740 ( new_n891_, keyIn_0_63 );
nor g741 ( new_n892_, new_n887_, keyIn_0_62 );
nor g742 ( new_n893_, new_n883_, new_n826_ );
nor g743 ( new_n894_, new_n892_, new_n893_ );
nand g744 ( new_n895_, new_n894_, new_n891_ );
nand g745 ( N878, new_n895_, new_n890_ );
nor g746 ( new_n897_, new_n737_, new_n727_ );
nor g747 ( new_n898_, new_n897_, new_n769_ );
nor g748 ( new_n899_, new_n898_, new_n718_ );
not g749 ( new_n900_, new_n899_ );
nand g750 ( new_n901_, new_n900_, new_n740_ );
not g751 ( new_n902_, new_n744_ );
nor g752 ( new_n903_, new_n902_, new_n710_ );
nand g753 ( new_n904_, new_n901_, new_n903_ );
nor g754 ( new_n905_, new_n901_, new_n903_ );
nor g755 ( new_n906_, new_n905_, new_n417_ );
nand g756 ( new_n907_, new_n906_, new_n904_ );
not g757 ( new_n908_, new_n903_ );
nor g758 ( new_n909_, new_n908_, new_n421_ );
nand g759 ( new_n910_, new_n902_, N237 );
nand g760 ( new_n911_, new_n709_, N246 );
nand g761 ( new_n912_, new_n431_, N165 );
nand g762 ( new_n913_, N91, N210 );
nand g763 ( new_n914_, new_n912_, new_n913_ );
not g764 ( new_n915_, new_n914_ );
nand g765 ( new_n916_, new_n911_, new_n915_ );
not g766 ( new_n917_, new_n916_ );
nand g767 ( new_n918_, new_n910_, new_n917_ );
nor g768 ( new_n919_, new_n909_, new_n918_ );
nand g769 ( N879, new_n907_, new_n919_ );
nand g770 ( new_n921_, new_n899_, new_n740_ );
not g771 ( new_n922_, new_n898_ );
not g772 ( new_n923_, new_n740_ );
nor g773 ( new_n924_, new_n923_, new_n718_ );
nor g774 ( new_n925_, new_n922_, new_n924_ );
nor g775 ( new_n926_, new_n925_, new_n417_ );
nand g776 ( new_n927_, new_n926_, new_n921_ );
not g777 ( new_n928_, new_n924_ );
nor g778 ( new_n929_, new_n928_, new_n421_ );
nand g779 ( new_n930_, new_n923_, N237 );
nand g780 ( new_n931_, new_n717_, N246 );
nand g781 ( new_n932_, new_n431_, N171 );
nand g782 ( new_n933_, N96, N210 );
nand g783 ( new_n934_, new_n932_, new_n933_ );
not g784 ( new_n935_, new_n934_ );
nand g785 ( new_n936_, new_n931_, new_n935_ );
not g786 ( new_n937_, new_n936_ );
nand g787 ( new_n938_, new_n930_, new_n937_ );
nor g788 ( new_n939_, new_n929_, new_n938_ );
nand g789 ( N880, new_n927_, new_n939_ );
endmodule