module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, WX660, WX661, n3513, WX662, WX663, n3511,
         WX664, WX665, n3509, WX666, WX667, WX668, WX669, n3505, WX670, WX671,
         n3503, WX672, WX673, n3501, WX674, WX675, WX676, WX677, n3497, WX678,
         WX679, n3495, WX680, WX681, n3493, WX682, WX683, n3491, WX684, WX685,
         n3489, WX686, WX688, WX689, n3485, WX690, WX691, n3483, WX692, WX693,
         n3481, WX694, WX695, n3479, WX696, WX697, n3477, WX698, WX699, n3475,
         WX700, WX701, n3473, WX702, WX703, n3471, WX704, WX705, n3469, WX706,
         WX707, n3467, WX708, WX709, WX710, WX711, WX712, WX713, WX714, WX715,
         WX716, WX717, WX718, WX719, WX720, WX721, WX722, WX724, WX725, WX726,
         WX727, WX728, WX729, WX730, WX731, WX732, WX733, WX734, WX735, WX736,
         WX737, WX738, WX739, WX740, WX741, WX742, WX743, WX744, WX745, WX746,
         WX747, WX748, WX749, WX750, WX751, WX752, WX753, WX754, WX755, WX756,
         WX757, WX758, WX760, WX761, WX762, WX763, WX764, WX765, WX766, WX767,
         WX768, WX769, WX770, WX771, WX772, WX773, WX774, WX775, WX776, WX777,
         WX778, WX779, WX780, WX781, WX782, WX783, WX784, WX785, WX786, WX787,
         WX788, WX789, WX790, WX791, WX792, WX793, WX794, WX796, WX797, WX798,
         WX799, WX800, WX801, WX802, WX803, WX804, WX805, WX806, WX807, WX808,
         WX809, WX810, WX811, WX812, WX813, WX814, WX815, WX816, WX817, WX818,
         WX819, WX820, WX821, WX822, WX823, WX824, WX825, WX826, WX827, WX828,
         WX829, WX830, WX832, WX833, WX834, WX835, WX836, WX837, WX838, WX839,
         WX840, WX841, WX842, WX843, WX844, WX845, WX846, WX847, WX848, WX849,
         WX850, WX851, WX852, WX853, WX854, WX855, WX856, WX857, WX858, WX859,
         WX860, WX861, WX862, WX863, WX864, WX865, WX866, WX868, WX869, WX870,
         WX871, WX872, WX873, WX874, WX875, WX876, WX877, WX878, WX879, WX880,
         WX881, WX882, WX883, WX884, WX885, WX886, WX887, WX888, WX889, WX890,
         WX891, WX892, WX893, WX894, WX895, WX896, WX897, WX898, WX899, WX1264,
         DFF_160_n1, WX1266, WX1268, DFF_162_n1, WX1270, WX1272, DFF_164_n1,
         WX1274, DFF_165_n1, WX1276, DFF_166_n1, WX1278, DFF_167_n1, WX1280,
         DFF_168_n1, WX1282, DFF_169_n1, WX1284, WX1286, DFF_171_n1, WX1288,
         DFF_172_n1, WX1290, DFF_173_n1, WX1292, DFF_174_n1, WX1294,
         DFF_175_n1, WX1296, DFF_176_n1, WX1298, DFF_177_n1, WX1300,
         DFF_178_n1, WX1302, WX1304, DFF_180_n1, WX1306, DFF_181_n1, WX1308,
         DFF_182_n1, WX1310, DFF_183_n1, WX1312, DFF_184_n1, WX1314,
         DFF_185_n1, WX1316, DFF_186_n1, WX1318, DFF_187_n1, WX1320,
         DFF_188_n1, WX1322, DFF_189_n1, WX1324, DFF_190_n1, WX1326,
         DFF_191_n1, WX1777, WX1778, WX1779, n8702, WX1781, n8701, WX1783,
         n8700, WX1785, n8699, WX1787, WX1789, n8696, WX1791, n8695, WX1793,
         n8694, WX1795, n8693, WX1797, n8692, WX1799, n8691, WX1801, n8690,
         WX1803, n8689, WX1805, n8688, WX1807, n8687, WX1809, n8686, WX1811,
         n8685, WX1813, n8684, WX1815, n8683, WX1817, n8682, WX1819, n8681,
         WX1821, n8680, WX1823, WX1825, n8677, WX1827, n8676, WX1829, n8675,
         WX1831, n8674, WX1833, n8673, WX1835, n8672, WX1837, n8671, WX1839,
         n8670, WX1937, n8669, WX1939, n8668, WX1941, n8667, WX1943, n8666,
         WX1945, n8665, WX1947, n8664, WX1949, n8663, WX1951, n8662, WX1953,
         n8661, WX1955, WX1957, n8658, WX1959, n8657, WX1961, n8656, WX1963,
         n8655, WX1965, n8654, WX1967, n8653, WX1969, WX1970, WX1971, WX1972,
         WX1973, WX1974, WX1975, WX1976, WX1977, WX1978, WX1979, WX1980,
         WX1981, WX1982, WX1983, WX1984, WX1985, WX1986, WX1987, WX1988,
         WX1989, WX1990, WX1991, WX1993, WX1994, WX1995, WX1996, WX1997,
         WX1998, WX1999, WX2000, WX2001, WX2002, WX2003, WX2004, WX2005,
         WX2006, WX2007, WX2008, WX2009, WX2010, WX2011, WX2012, WX2013,
         WX2014, WX2015, WX2016, WX2017, WX2018, WX2019, WX2020, WX2021,
         WX2022, WX2023, WX2024, WX2025, WX2026, WX2027, WX2029, WX2030,
         WX2031, WX2032, WX2033, WX2034, WX2035, WX2036, n3783, WX2037, WX2038,
         WX2039, WX2040, WX2041, WX2042, WX2043, WX2044, n3775, WX2045, WX2046,
         WX2047, WX2048, WX2049, WX2050, WX2051, WX2052, WX2053, WX2054,
         WX2055, WX2056, n3763, WX2057, WX2058, WX2059, WX2060, WX2061, WX2062,
         WX2063, WX2065, WX2066, WX2067, WX2068, WX2069, WX2070, WX2071,
         WX2072, WX2073, WX2074, WX2075, WX2076, WX2077, WX2078, WX2079,
         WX2080, WX2081, WX2082, WX2083, WX2084, WX2085, WX2086, WX2087,
         WX2088, WX2089, WX2090, WX2091, WX2092, WX2093, WX2094, WX2095,
         WX2096, WX2097, WX2098, WX2099, WX2101, WX2102, WX2103, WX2104,
         WX2105, WX2106, WX2107, WX2108, WX2109, WX2110, WX2111, WX2112,
         WX2113, WX2114, WX2115, WX2116, WX2117, WX2118, WX2119, WX2120,
         WX2121, WX2122, WX2123, WX2124, WX2125, WX2126, WX2127, WX2128,
         WX2129, WX2130, WX2131, WX2132, WX2133, WX2134, WX2135, WX2137,
         WX2138, WX2139, WX2140, WX2141, WX2142, WX2143, WX2144, WX2145,
         WX2146, WX2147, WX2148, WX2149, WX2150, WX2151, WX2152, WX2153,
         WX2154, WX2155, WX2156, WX2157, WX2158, WX2159, WX2160, WX2161,
         WX2162, WX2163, WX2164, WX2165, WX2166, WX2167, WX2168, WX2169,
         WX2170, WX2171, WX2173, WX2174, WX2175, WX2176, WX2177, WX2178,
         WX2179, WX2180, WX2181, WX2182, WX2183, WX2184, WX2185, WX2186,
         WX2187, WX2188, WX2189, WX2190, WX2191, WX2192, WX2557, DFF_352_n1,
         WX2559, DFF_353_n1, WX2561, DFF_354_n1, WX2563, WX2565, DFF_356_n1,
         WX2567, DFF_357_n1, WX2569, DFF_358_n1, WX2571, WX2573, DFF_360_n1,
         WX2575, WX2577, WX2579, DFF_363_n1, WX2581, DFF_364_n1, WX2583,
         DFF_365_n1, WX2585, DFF_366_n1, WX2587, WX2589, DFF_368_n1, WX2591,
         DFF_369_n1, WX2593, DFF_370_n1, WX2595, DFF_371_n1, WX2597,
         DFF_372_n1, WX2599, DFF_373_n1, WX2601, DFF_374_n1, WX2603,
         DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609, DFF_378_n1, WX2611,
         WX2613, DFF_380_n1, WX2615, DFF_381_n1, WX2617, DFF_382_n1, WX2619,
         DFF_383_n1, WX3070, WX3071, WX3072, n8644, WX3074, n8643, WX3076,
         n8642, WX3078, n8641, WX3080, n8640, WX3082, n8639, WX3084, n8638,
         WX3086, n8637, WX3088, n8636, WX3090, n8635, WX3092, WX3094, n8632,
         WX3096, n8631, WX3098, n8630, WX3100, n8629, WX3102, n8628, WX3104,
         n8627, WX3106, n8626, WX3108, n8625, WX3110, n8624, WX3112, n8623,
         WX3114, n8622, WX3116, n8621, WX3118, n8620, WX3120, n8619, WX3122,
         n8618, WX3124, n8617, WX3126, n8616, WX3128, WX3130, n8613, WX3132,
         n8612, WX3230, n8611, WX3232, n8610, WX3234, n8609, WX3236, n8608,
         WX3238, n8607, WX3240, n8606, WX3242, n8605, WX3244, n8604, WX3246,
         n8603, WX3248, n8602, WX3250, n8601, WX3252, n8600, WX3254, n8599,
         WX3256, n8598, WX3258, n8597, WX3260, WX3262, WX3263, WX3264, WX3265,
         WX3266, WX3267, WX3268, WX3269, WX3270, WX3271, WX3272, WX3273,
         WX3274, WX3275, WX3276, WX3277, WX3278, WX3279, WX3280, WX3281,
         WX3282, WX3283, WX3284, WX3285, WX3286, WX3287, WX3288, WX3289,
         WX3290, WX3291, WX3292, WX3293, WX3294, WX3295, WX3296, WX3298,
         WX3299, WX3300, WX3301, WX3302, WX3303, WX3304, WX3305, WX3306,
         WX3307, WX3308, WX3309, WX3310, WX3311, WX3312, WX3313, WX3314,
         WX3315, WX3316, WX3317, WX3318, WX3319, WX3320, WX3321, WX3322,
         WX3323, WX3324, WX3325, WX3326, WX3327, WX3328, WX3329, WX3330,
         WX3331, WX3332, WX3334, WX3335, WX3336, WX3337, WX3338, WX3339,
         WX3340, WX3341, n3739, WX3342, WX3343, WX3344, WX3345, n3735, WX3346,
         WX3347, WX3348, WX3349, WX3350, WX3351, WX3352, WX3353, WX3354,
         WX3355, WX3356, WX3357, WX3358, WX3359, WX3360, WX3361, WX3362,
         WX3363, WX3364, WX3365, WX3366, WX3367, WX3368, WX3370, WX3371,
         WX3372, WX3373, WX3374, WX3375, WX3376, WX3377, WX3378, WX3379,
         WX3380, WX3381, WX3382, WX3383, WX3384, WX3385, WX3386, WX3387,
         WX3388, WX3389, WX3390, WX3391, WX3392, WX3393, WX3394, WX3395,
         WX3396, WX3397, WX3398, WX3399, WX3400, WX3401, WX3402, WX3403,
         WX3404, WX3406, WX3407, WX3408, WX3409, WX3410, WX3411, WX3412,
         WX3413, WX3414, WX3415, WX3416, WX3417, WX3418, WX3419, WX3420,
         WX3421, WX3422, WX3423, WX3424, WX3425, WX3426, WX3427, WX3428,
         WX3429, WX3430, WX3431, WX3432, WX3433, WX3434, WX3435, WX3436,
         WX3437, WX3438, WX3440, WX3441, WX3442, WX3443, WX3444, WX3445,
         WX3446, WX3447, WX3448, WX3449, WX3450, WX3451, WX3452, WX3453,
         WX3454, WX3455, WX3456, WX3457, WX3458, WX3459, WX3460, WX3461,
         WX3462, WX3463, WX3464, WX3465, WX3466, WX3467, WX3468, WX3469,
         WX3470, WX3471, WX3472, WX3474, WX3475, WX3476, WX3477, WX3478,
         WX3479, WX3480, WX3481, WX3482, WX3483, WX3484, WX3485, WX3850,
         DFF_544_n1, WX3852, DFF_545_n1, WX3854, DFF_546_n1, WX3856, WX3858,
         DFF_548_n1, WX3860, WX3862, DFF_550_n1, WX3864, DFF_551_n1, WX3866,
         DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872, DFF_555_n1, WX3874,
         DFF_556_n1, WX3876, DFF_557_n1, WX3878, DFF_558_n1, WX3880, WX3882,
         DFF_560_n1, WX3884, DFF_561_n1, WX3886, DFF_562_n1, WX3888,
         DFF_563_n1, WX3890, DFF_564_n1, WX3892, DFF_565_n1, WX3894, WX3896,
         DFF_567_n1, WX3898, DFF_568_n1, WX3900, DFF_569_n1, WX3902,
         DFF_570_n1, WX3904, WX3906, DFF_572_n1, WX3908, DFF_573_n1, WX3910,
         DFF_574_n1, WX3912, DFF_575_n1, WX4363, WX4364, WX4365, n8586, WX4367,
         n8585, WX4369, n8584, WX4371, n8583, WX4373, n8582, WX4375, n8581,
         WX4377, n8580, WX4379, n8579, WX4381, n8578, WX4383, n8577, WX4385,
         n8576, WX4387, WX4389, n8573, WX4391, n8572, WX4393, n8571, WX4395,
         n8570, WX4397, n8569, WX4399, n8568, WX4401, n8567, WX4403, n8566,
         WX4405, n8565, WX4407, n8564, WX4409, n8563, WX4411, n8562, WX4413,
         n8561, WX4415, n8560, WX4417, n8559, WX4419, n8558, WX4421, WX4423,
         n8555, WX4425, n8554, WX4523, n8553, WX4525, n8552, WX4527, n8551,
         WX4529, n8550, WX4531, n8549, WX4533, n8548, WX4535, n8547, WX4537,
         n8546, WX4539, n8545, WX4541, n8544, WX4543, n8543, WX4545, n8542,
         WX4547, n8541, WX4549, n8540, WX4551, WX4553, n8537, WX4555, WX4556,
         WX4557, WX4558, WX4559, WX4560, WX4561, WX4562, WX4563, WX4564,
         WX4565, WX4566, WX4567, WX4568, WX4569, WX4570, WX4571, WX4572,
         WX4573, WX4574, WX4575, WX4576, WX4577, WX4578, WX4579, WX4580,
         WX4581, WX4582, WX4583, WX4584, WX4585, WX4587, WX4588, WX4589,
         WX4590, WX4591, WX4592, WX4593, WX4594, WX4595, WX4596, WX4597,
         WX4598, WX4599, WX4600, WX4601, WX4602, WX4603, WX4604, WX4605,
         WX4606, WX4607, WX4608, WX4609, WX4610, WX4611, WX4612, WX4613,
         WX4614, WX4615, WX4616, WX4617, WX4618, WX4619, WX4621, WX4622,
         WX4623, WX4624, n3717, WX4625, WX4626, WX4627, WX4628, n3713, WX4629,
         WX4630, WX4631, WX4632, WX4633, WX4634, WX4635, WX4636, WX4637,
         WX4638, WX4639, WX4640, WX4641, WX4642, WX4643, WX4644, WX4645,
         WX4646, WX4647, WX4648, WX4649, WX4650, n3691, WX4651, WX4652, WX4653,
         WX4655, WX4656, WX4657, WX4658, WX4659, WX4660, WX4661, WX4662,
         WX4663, WX4664, WX4665, WX4666, WX4667, WX4668, WX4669, WX4670,
         WX4671, WX4672, WX4673, WX4674, WX4675, WX4676, WX4677, WX4678,
         WX4679, WX4680, WX4681, WX4682, WX4683, WX4684, WX4685, WX4686,
         WX4687, WX4689, WX4690, WX4691, WX4692, WX4693, WX4694, WX4695,
         WX4696, WX4697, WX4698, WX4699, WX4700, WX4701, WX4702, WX4703,
         WX4704, WX4705, WX4706, WX4707, WX4708, WX4709, WX4710, WX4711,
         WX4712, WX4713, WX4714, WX4715, WX4716, WX4717, WX4718, WX4719,
         WX4720, WX4721, WX4723, WX4724, WX4725, WX4726, WX4727, WX4728,
         WX4729, WX4730, WX4731, WX4732, WX4733, WX4734, WX4735, WX4736,
         WX4737, WX4738, WX4739, WX4740, WX4741, WX4742, WX4743, WX4744,
         WX4745, WX4746, WX4747, WX4748, WX4749, WX4750, WX4751, WX4752,
         WX4753, WX4754, WX4755, WX4757, WX4758, WX4759, WX4760, WX4761,
         WX4762, WX4763, WX4764, WX4765, WX4766, WX4767, WX4768, WX4769,
         WX4770, WX4771, WX4772, WX4773, WX4774, WX4775, WX4776, WX4777,
         WX4778, WX5143, DFF_736_n1, WX5145, DFF_737_n1, WX5147, DFF_738_n1,
         WX5149, WX5151, DFF_740_n1, WX5153, WX5155, DFF_742_n1, WX5157,
         DFF_743_n1, WX5159, DFF_744_n1, WX5161, DFF_745_n1, WX5163,
         DFF_746_n1, WX5165, DFF_747_n1, WX5167, DFF_748_n1, WX5169,
         DFF_749_n1, WX5171, DFF_750_n1, WX5173, WX5175, DFF_752_n1, WX5177,
         DFF_753_n1, WX5179, DFF_754_n1, WX5181, DFF_755_n1, WX5183,
         DFF_756_n1, WX5185, DFF_757_n1, WX5187, WX5189, DFF_759_n1, WX5191,
         DFF_760_n1, WX5193, DFF_761_n1, WX5195, DFF_762_n1, WX5197, WX5199,
         DFF_764_n1, WX5201, DFF_765_n1, WX5203, DFF_766_n1, WX5205,
         DFF_767_n1, WX5656, WX5657, WX5658, n8528, WX5660, n8527, WX5662,
         n8526, WX5664, n8525, WX5666, n8524, WX5668, n8523, WX5670, WX5672,
         n8520, WX5674, n8519, WX5676, n8518, WX5678, n8517, WX5680, n8516,
         WX5682, n8515, WX5684, n8514, WX5686, n8513, WX5688, n8512, WX5690,
         n8511, WX5692, n8510, WX5694, n8509, WX5696, n8508, WX5698, n8507,
         WX5700, n8506, WX5702, n8505, WX5704, WX5706, n8502, WX5708, n8501,
         WX5710, n8500, WX5712, n8499, WX5714, n8498, WX5716, n8497, WX5718,
         n8496, WX5816, n8495, WX5818, n8494, WX5820, n8493, WX5822, n8492,
         WX5824, n8491, WX5826, n8490, WX5828, n8489, WX5830, n8488, WX5832,
         n8487, WX5834, WX5836, n8484, WX5838, n8483, WX5840, n8482, WX5842,
         n8481, WX5844, n8480, WX5846, n8479, WX5848, WX5849, WX5850, WX5851,
         WX5852, WX5853, WX5854, WX5855, WX5856, WX5857, WX5858, WX5859,
         WX5860, WX5861, WX5862, WX5863, WX5864, WX5865, WX5866, WX5867,
         WX5868, WX5870, WX5871, WX5872, WX5873, WX5874, WX5875, WX5876,
         WX5877, WX5878, WX5879, WX5880, WX5881, WX5882, WX5883, WX5884,
         WX5885, WX5886, WX5887, WX5888, WX5889, WX5890, WX5891, WX5892,
         WX5893, WX5894, WX5895, WX5896, WX5897, WX5898, WX5899, WX5900,
         WX5901, WX5902, WX5904, WX5905, WX5906, WX5907, WX5908, WX5909,
         WX5910, WX5911, WX5912, WX5913, WX5914, WX5915, WX5916, WX5917,
         WX5918, WX5919, WX5920, WX5921, WX5922, WX5923, WX5924, WX5925,
         WX5926, WX5927, WX5928, WX5929, WX5930, WX5931, WX5932, WX5933, n3669,
         WX5934, WX5935, WX5936, WX5938, WX5939, WX5940, WX5941, n3661, WX5942,
         WX5943, WX5944, WX5945, WX5946, WX5947, WX5948, WX5949, WX5950,
         WX5951, WX5952, WX5953, WX5954, WX5955, WX5956, WX5957, WX5958,
         WX5959, WX5960, WX5961, WX5962, WX5963, WX5964, WX5965, WX5966,
         WX5967, WX5968, WX5969, WX5970, WX5972, WX5973, WX5974, WX5975,
         WX5976, WX5977, WX5978, WX5979, WX5980, WX5981, WX5982, WX5983,
         WX5984, WX5985, WX5986, WX5987, WX5988, WX5989, WX5990, WX5991,
         WX5992, WX5993, WX5994, WX5995, WX5996, WX5997, WX5998, WX5999,
         WX6000, WX6001, WX6002, WX6003, WX6004, WX6006, WX6007, WX6008,
         WX6009, WX6010, WX6011, WX6012, WX6013, WX6014, WX6015, WX6016,
         WX6017, WX6018, WX6019, WX6020, WX6021, WX6022, WX6023, WX6024,
         WX6025, WX6026, WX6027, WX6028, WX6029, WX6030, WX6031, WX6032,
         WX6033, WX6034, WX6035, WX6036, WX6037, WX6038, WX6040, WX6041,
         WX6042, WX6043, WX6044, WX6045, WX6046, WX6047, WX6048, WX6049,
         WX6050, WX6051, WX6052, WX6053, WX6054, WX6055, WX6056, WX6057,
         WX6058, WX6059, WX6060, WX6061, WX6062, WX6063, WX6064, WX6065,
         WX6066, WX6067, WX6068, WX6069, WX6070, WX6071, WX6436, WX6438,
         DFF_929_n1, WX6440, DFF_930_n1, WX6442, WX6444, DFF_932_n1, WX6446,
         DFF_933_n1, WX6448, DFF_934_n1, WX6450, DFF_935_n1, WX6452,
         DFF_936_n1, WX6454, DFF_937_n1, WX6456, WX6458, DFF_939_n1, WX6460,
         DFF_940_n1, WX6462, DFF_941_n1, WX6464, DFF_942_n1, WX6466,
         DFF_943_n1, WX6468, DFF_944_n1, WX6470, WX6472, DFF_946_n1, WX6474,
         DFF_947_n1, WX6476, DFF_948_n1, WX6478, DFF_949_n1, WX6480,
         DFF_950_n1, WX6482, DFF_951_n1, WX6484, DFF_952_n1, WX6486,
         DFF_953_n1, WX6488, DFF_954_n1, WX6490, DFF_955_n1, WX6492,
         DFF_956_n1, WX6494, DFF_957_n1, WX6496, DFF_958_n1, WX6498,
         DFF_959_n1, WX6949, WX6950, WX6951, n8470, WX6953, WX6955, n8467,
         WX6957, n8466, WX6959, n8465, WX6961, n8464, WX6963, n8463, WX6965,
         n8462, WX6967, n8461, WX6969, n8460, WX6971, n8459, WX6973, n8458,
         WX6975, n8457, WX6977, n8456, WX6979, n8455, WX6981, n8454, WX6983,
         n8453, WX6985, n8452, WX6987, WX6989, n8449, WX6991, n8448, WX6993,
         n8447, WX6995, n8446, WX6997, n8445, WX6999, n8444, WX7001, n8443,
         WX7003, n8442, WX7005, n8441, WX7007, n8440, WX7009, n8439, WX7011,
         n8438, WX7109, n8437, WX7111, n8436, WX7113, n8435, WX7115, n8434,
         WX7117, WX7119, n8431, WX7121, n8430, WX7123, n8429, WX7125, n8428,
         WX7127, n8427, WX7129, n8426, WX7131, n8425, WX7133, n8424, WX7135,
         n8423, WX7137, n8422, WX7139, n8421, WX7141, WX7142, WX7143, WX7144,
         WX7145, WX7146, WX7147, WX7148, WX7149, WX7150, WX7151, WX7153,
         WX7154, WX7155, WX7156, WX7157, WX7158, WX7159, WX7160, WX7161,
         WX7162, WX7163, WX7164, WX7165, WX7166, WX7167, WX7168, WX7169,
         WX7170, WX7171, WX7172, WX7173, WX7174, WX7175, WX7176, WX7177,
         WX7178, WX7179, WX7180, WX7181, WX7182, WX7183, WX7184, WX7185,
         WX7187, WX7188, WX7189, WX7190, WX7191, WX7192, WX7193, WX7194,
         WX7195, WX7196, WX7197, WX7198, WX7199, WX7200, WX7201, WX7202,
         WX7203, WX7204, WX7205, WX7206, WX7207, WX7208, WX7209, WX7210,
         WX7211, WX7212, WX7213, WX7214, WX7215, WX7216, n3647, WX7217, WX7218,
         WX7219, WX7221, WX7222, WX7223, WX7224, n3639, WX7225, WX7226, WX7227,
         WX7228, n3635, WX7229, WX7230, WX7231, WX7232, WX7233, WX7234, WX7235,
         WX7236, WX7237, WX7238, WX7239, WX7240, WX7241, WX7242, WX7243,
         WX7244, WX7245, WX7246, WX7247, WX7248, WX7249, WX7250, WX7251,
         WX7252, WX7253, WX7255, WX7256, WX7257, WX7258, WX7259, WX7260,
         WX7261, WX7262, WX7263, WX7264, WX7265, WX7266, WX7267, WX7268,
         WX7269, WX7270, WX7271, WX7272, WX7273, WX7274, WX7275, WX7276,
         WX7277, WX7278, WX7279, WX7280, WX7281, WX7282, WX7283, WX7284,
         WX7285, WX7286, WX7287, WX7289, WX7290, WX7291, WX7292, WX7293,
         WX7294, WX7295, WX7296, WX7297, WX7298, WX7299, WX7300, WX7301,
         WX7302, WX7303, WX7304, WX7305, WX7306, WX7307, WX7308, WX7309,
         WX7310, WX7311, WX7312, WX7313, WX7314, WX7315, WX7316, WX7317,
         WX7318, WX7319, WX7320, WX7321, WX7323, WX7324, WX7325, WX7326,
         WX7327, WX7328, WX7329, WX7330, WX7331, WX7332, WX7333, WX7334,
         WX7335, WX7336, WX7337, WX7338, WX7339, WX7340, WX7341, WX7342,
         WX7343, WX7344, WX7345, WX7346, WX7347, WX7348, WX7349, WX7350,
         WX7351, WX7352, WX7353, WX7354, WX7355, WX7357, WX7358, WX7359,
         WX7360, WX7361, WX7362, WX7363, WX7364, WX7729, DFF_1120_n1, WX7731,
         DFF_1121_n1, WX7733, DFF_1122_n1, WX7735, DFF_1123_n1, WX7737,
         DFF_1124_n1, WX7739, DFF_1125_n1, WX7741, DFF_1126_n1, WX7743,
         DFF_1127_n1, WX7745, DFF_1128_n1, WX7747, DFF_1129_n1, WX7749, WX7751,
         DFF_1131_n1, WX7753, WX7755, DFF_1133_n1, WX7757, DFF_1134_n1, WX7759,
         WX7761, DFF_1136_n1, WX7763, DFF_1137_n1, WX7765, DFF_1138_n1, WX7767,
         DFF_1139_n1, WX7769, WX7771, DFF_1141_n1, WX7773, DFF_1142_n1, WX7775,
         DFF_1143_n1, WX7777, DFF_1144_n1, WX7779, DFF_1145_n1, WX7781,
         DFF_1146_n1, WX7783, DFF_1147_n1, WX7785, DFF_1148_n1, WX7787, WX7789,
         DFF_1150_n1, WX7791, DFF_1151_n1, WX8242, WX8243, WX8244, n8411,
         WX8246, n8410, WX8248, n8409, WX8250, n8408, WX8252, n8407, WX8254,
         n8406, WX8256, n8405, WX8258, n8404, WX8260, n8403, WX8262, n8402,
         WX8264, n8401, WX8266, n8400, WX8268, n8399, WX8270, WX8272, n8396,
         WX8274, n8395, WX8276, n8394, WX8278, n8393, WX8280, n8392, WX8282,
         n8391, WX8284, n8390, WX8286, n8389, WX8288, n8388, WX8290, n8387,
         WX8292, n8386, WX8294, n8385, WX8296, n8384, WX8298, n8383, WX8300,
         n8382, WX8302, n8381, WX8304, WX8402, n8378, WX8404, n8377, WX8406,
         n8376, WX8408, n8375, WX8410, n8374, WX8412, n8373, WX8414, n8372,
         WX8416, n8371, WX8418, n8370, WX8420, n8369, WX8422, n8368, WX8424,
         n8367, WX8426, n8366, WX8428, n8365, WX8430, n8364, WX8432, n8363,
         WX8434, WX8436, WX8437, WX8438, WX8439, WX8440, WX8441, WX8442,
         WX8443, WX8444, WX8445, WX8446, WX8447, WX8448, WX8449, WX8450,
         WX8451, WX8452, WX8453, WX8454, WX8455, WX8456, WX8457, WX8458,
         WX8459, WX8460, WX8461, WX8462, WX8463, WX8464, WX8465, WX8466,
         WX8467, WX8468, WX8470, WX8471, WX8472, WX8473, WX8474, WX8475,
         WX8476, WX8477, WX8478, WX8479, WX8480, WX8481, WX8482, WX8483,
         WX8484, WX8485, WX8486, WX8487, WX8488, WX8489, WX8490, WX8491,
         WX8492, WX8493, WX8494, WX8495, WX8496, WX8497, WX8498, WX8499, n3625,
         WX8500, WX8501, WX8502, WX8504, WX8505, WX8506, WX8507, n3617, WX8508,
         WX8509, WX8510, WX8511, n3613, WX8512, WX8513, WX8514, WX8515, WX8516,
         WX8517, WX8518, WX8519, WX8520, WX8521, WX8522, WX8523, WX8524,
         WX8525, WX8526, WX8527, WX8528, WX8529, WX8530, WX8531, WX8532,
         WX8533, WX8534, WX8535, WX8536, WX8538, WX8539, WX8540, WX8541,
         WX8542, WX8543, WX8544, WX8545, WX8546, WX8547, WX8548, WX8549,
         WX8550, WX8551, WX8552, WX8553, WX8554, WX8555, WX8556, WX8557,
         WX8558, WX8559, WX8560, WX8561, WX8562, WX8563, WX8564, WX8565,
         WX8566, WX8567, WX8568, WX8569, WX8570, WX8572, WX8573, WX8574,
         WX8575, WX8576, WX8577, WX8578, WX8579, WX8580, WX8581, WX8582,
         WX8583, WX8584, WX8585, WX8586, WX8587, WX8588, WX8589, WX8590,
         WX8591, WX8592, WX8593, WX8594, WX8595, WX8596, WX8597, WX8598,
         WX8599, WX8600, WX8601, WX8602, WX8603, WX8604, WX8606, WX8607,
         WX8608, WX8609, WX8610, WX8611, WX8612, WX8613, WX8614, WX8615,
         WX8616, WX8617, WX8618, WX8619, WX8620, WX8621, WX8622, WX8623,
         WX8624, WX8625, WX8626, WX8627, WX8628, WX8629, WX8630, WX8631,
         WX8632, WX8633, WX8634, WX8635, WX8636, WX8637, WX8638, WX8640,
         WX8641, WX8642, WX8643, WX8644, WX8645, WX8646, WX8647, WX8648,
         WX8649, WX8650, WX8651, WX8652, WX8653, WX8654, WX8655, WX8656,
         WX8657, WX9022, DFF_1312_n1, WX9024, DFF_1313_n1, WX9026, DFF_1314_n1,
         WX9028, WX9030, DFF_1316_n1, WX9032, DFF_1317_n1, WX9034, DFF_1318_n1,
         WX9036, WX9038, WX9040, DFF_1321_n1, WX9042, WX9044, DFF_1323_n1,
         WX9046, DFF_1324_n1, WX9048, DFF_1325_n1, WX9050, DFF_1326_n1, WX9052,
         WX9054, DFF_1328_n1, WX9056, DFF_1329_n1, WX9058, DFF_1330_n1, WX9060,
         DFF_1331_n1, WX9062, DFF_1332_n1, WX9064, DFF_1333_n1, WX9066,
         DFF_1334_n1, WX9068, DFF_1335_n1, WX9070, WX9072, WX9074, DFF_1338_n1,
         WX9076, DFF_1339_n1, WX9078, DFF_1340_n1, WX9080, DFF_1341_n1, WX9082,
         DFF_1342_n1, WX9084, DFF_1343_n1, WX9535, WX9536, WX9537, n8353,
         WX9539, n8352, WX9541, n8351, WX9543, n8350, WX9545, n8349, WX9547,
         n8348, WX9549, n8347, WX9551, n8346, WX9553, WX9555, n8343, WX9557,
         n8342, WX9559, n8341, WX9561, n8340, WX9563, n8339, WX9565, n8338,
         WX9567, n8337, WX9569, n8336, WX9571, n8335, WX9573, n8334, WX9575,
         n8333, WX9577, n8332, WX9579, n8331, WX9581, n8330, WX9583, n8329,
         WX9585, n8328, WX9587, WX9589, n8325, WX9591, n8324, WX9593, n8323,
         WX9595, n8322, WX9597, n8321, WX9695, n8320, WX9697, n8319, WX9699,
         n8318, WX9701, n8317, WX9703, n8316, WX9705, n8315, WX9707, n8314,
         WX9709, n8313, WX9711, n8312, WX9713, n8311, WX9715, n8310, WX9717,
         WX9719, n8307, WX9721, n8306, WX9723, n8305, WX9725, n8304, WX9727,
         WX9728, WX9729, WX9730, WX9731, WX9732, WX9733, WX9734, WX9735,
         WX9736, WX9737, WX9738, WX9739, WX9740, WX9741, WX9742, WX9743,
         WX9744, WX9745, WX9746, WX9747, WX9748, WX9749, WX9750, WX9751,
         WX9753, WX9754, WX9755, WX9756, WX9757, WX9758, WX9759, WX9760,
         WX9761, WX9762, WX9763, WX9764, WX9765, WX9766, WX9767, WX9768,
         WX9769, WX9770, WX9771, WX9772, WX9773, WX9774, WX9775, WX9776,
         WX9777, WX9778, WX9779, WX9780, WX9781, WX9782, WX9783, WX9784,
         WX9785, WX9787, WX9788, WX9789, WX9790, WX9791, WX9792, WX9793,
         WX9794, n3591, WX9795, WX9796, WX9797, WX9798, WX9799, WX9800, WX9801,
         WX9802, WX9803, WX9804, WX9805, WX9806, WX9807, WX9808, WX9809,
         WX9810, WX9811, WX9812, WX9813, WX9814, WX9815, WX9816, n3569, WX9817,
         WX9818, WX9819, WX9821, WX9822, WX9823, WX9824, WX9825, WX9826,
         WX9827, WX9828, WX9829, WX9830, WX9831, WX9832, WX9833, WX9834,
         WX9835, WX9836, WX9837, WX9838, WX9839, WX9840, WX9841, WX9842,
         WX9843, WX9844, WX9845, WX9846, WX9847, WX9848, WX9849, WX9850,
         WX9851, WX9852, WX9853, WX9855, WX9856, WX9857, WX9858, WX9859,
         WX9860, WX9861, WX9862, WX9863, WX9864, WX9865, WX9866, WX9867,
         WX9868, WX9869, WX9870, WX9871, WX9872, WX9873, WX9874, WX9875,
         WX9876, WX9877, WX9878, WX9879, WX9880, WX9881, WX9882, WX9883,
         WX9884, WX9885, WX9886, WX9887, WX9889, WX9890, WX9891, WX9892,
         WX9893, WX9894, WX9895, WX9896, WX9897, WX9898, WX9899, WX9900,
         WX9901, WX9902, WX9903, WX9904, WX9905, WX9906, WX9907, WX9908,
         WX9909, WX9910, WX9911, WX9912, WX9913, WX9914, WX9915, WX9916,
         WX9917, WX9918, WX9919, WX9920, WX9921, WX9923, WX9924, WX9925,
         WX9926, WX9927, WX9928, WX9929, WX9930, WX9931, WX9932, WX9933,
         WX9934, WX9935, WX9936, WX9937, WX9938, WX9939, WX9940, WX9941,
         WX9942, WX9943, WX9944, WX9945, WX9946, WX9947, WX9948, WX9949,
         WX9950, WX10315, DFF_1504_n1, WX10317, DFF_1505_n1, WX10319, WX10321,
         WX10323, DFF_1508_n1, WX10325, DFF_1509_n1, WX10327, DFF_1510_n1,
         WX10329, DFF_1511_n1, WX10331, DFF_1512_n1, WX10333, DFF_1513_n1,
         WX10335, WX10337, DFF_1515_n1, WX10339, DFF_1516_n1, WX10341, WX10343,
         DFF_1518_n1, WX10345, WX10347, DFF_1520_n1, WX10349, DFF_1521_n1,
         WX10351, DFF_1522_n1, WX10353, WX10355, DFF_1524_n1, WX10357,
         DFF_1525_n1, WX10359, DFF_1526_n1, WX10361, DFF_1527_n1, WX10363,
         DFF_1528_n1, WX10365, DFF_1529_n1, WX10367, DFF_1530_n1, WX10369,
         DFF_1531_n1, WX10371, DFF_1532_n1, WX10373, DFF_1533_n1, WX10375,
         WX10377, DFF_1535_n1, WX10828, WX10829, WX10830, n8295, WX10832,
         n8294, WX10834, n8293, WX10836, WX10838, n8290, WX10840, n8289,
         WX10842, n8288, WX10844, n8287, WX10846, n8286, WX10848, n8285,
         WX10850, n8284, WX10852, n8283, WX10854, n8282, WX10856, n8281,
         WX10858, n8280, WX10860, n8279, WX10862, n8278, WX10864, n8277,
         WX10866, n8276, WX10868, n8275, WX10870, WX10872, n8272, WX10874,
         n8271, WX10876, n8270, WX10878, n8269, WX10880, n8268, WX10882, n8267,
         WX10884, n8266, WX10886, n8265, WX10888, n8264, WX10890, n8263,
         WX10988, n8262, WX10990, n8261, WX10992, n8260, WX10994, n8259,
         WX10996, n8258, WX10998, n8257, WX11000, WX11002, n8254, WX11004,
         n8253, WX11006, n8252, WX11008, n8251, WX11010, n8250, WX11012, n8249,
         WX11014, n8248, WX11016, n8247, WX11018, n8246, WX11020, WX11021,
         WX11022, WX11023, WX11024, WX11025, WX11026, WX11027, WX11028,
         WX11029, WX11030, WX11031, WX11032, WX11033, WX11034, WX11036,
         WX11037, WX11038, WX11039, WX11040, WX11041, WX11042, WX11043,
         WX11044, WX11045, WX11046, WX11047, WX11048, WX11049, WX11050,
         WX11051, WX11052, WX11053, WX11054, WX11055, WX11056, WX11057,
         WX11058, WX11059, WX11060, WX11061, WX11062, WX11063, WX11064,
         WX11065, WX11066, WX11067, WX11068, WX11070, WX11071, WX11072,
         WX11073, WX11074, WX11075, WX11076, WX11077, WX11078, WX11079,
         WX11080, WX11081, WX11082, WX11083, WX11084, WX11085, WX11086,
         WX11087, WX11088, WX11089, WX11090, WX11091, WX11092, WX11093,
         WX11094, WX11095, WX11096, WX11097, WX11098, WX11099, n3547, WX11100,
         WX11101, WX11102, WX11104, WX11105, WX11106, WX11107, n3539, WX11108,
         WX11109, WX11110, WX11111, n3535, WX11112, WX11113, WX11114, WX11115,
         WX11116, WX11117, WX11118, WX11119, WX11120, WX11121, WX11122,
         WX11123, WX11124, WX11125, WX11126, WX11127, WX11128, WX11129,
         WX11130, WX11131, WX11132, WX11133, WX11134, WX11135, WX11136,
         WX11138, WX11139, WX11140, WX11141, WX11142, WX11143, WX11144,
         WX11145, WX11146, WX11147, WX11148, WX11149, WX11150, WX11151,
         WX11152, WX11153, WX11154, WX11155, WX11156, WX11155_Tj_Payload,
         test_se_Trojan, WX11157, WX11158, WX11159, WX11160, WX11161, WX11162,
         WX11163, WX11164, WX11165, WX11166, WX11167, WX11168, WX11169,
         WX11170, WX11172, WX11173, WX11174, WX11175, WX11176, WX11177,
         WX11178, WX11179, WX11180, WX11181, WX11182, WX11183, WX11184,
         WX11185, WX11186, WX11187, WX11188, WX11189, WX11190, WX11191,
         WX11192, WX11193, WX11194, WX11195, WX11196, WX11197, WX11198,
         WX11199, WX11200, WX11201, WX11202, WX11203, WX11204, WX11206,
         WX11207, WX11208, WX11209, WX11210, WX11211, WX11212, WX11213,
         WX11214, WX11215, WX11216, WX11217, WX11218, WX11219, WX11220,
         WX11221, WX11222, WX11223, WX11224, WX11225, WX11226, WX11227,
         WX11228, WX11229, WX11230, WX11231, WX11232, WX11233, WX11234,
         WX11235, WX11236, WX11237, WX11238, WX11240, WX11241, WX11242,
         WX11243, WX11608, DFF_1696_n1, WX11610, WX11612, DFF_1698_n1, WX11614,
         DFF_1699_n1, WX11616, DFF_1700_n1, WX11618, DFF_1701_n1, WX11620,
         DFF_1702_n1, WX11622, DFF_1703_n1, WX11624, DFF_1704_n1, WX11626,
         DFF_1705_n1, WX11628, DFF_1706_n1, WX11630, DFF_1707_n1, WX11632,
         DFF_1708_n1, WX11634, DFF_1709_n1, WX11636, WX11638, DFF_1711_n1,
         WX11640, DFF_1712_n1, WX11642, DFF_1713_n1, WX11644, WX11646,
         DFF_1715_n1, WX11648, DFF_1716_n1, WX11650, DFF_1717_n1, WX11652,
         DFF_1718_n1, WX11654, DFF_1719_n1, WX11656, DFF_1720_n1, WX11658,
         DFF_1721_n1, WX11660, DFF_1722_n1, WX11662, DFF_1723_n1, WX11664,
         DFF_1724_n1, WX11666, DFF_1725_n1, WX11668, DFF_1726_n1, WX11670,
         n2245, n2153, n3278, n2152, n2148, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4,
         Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         test_se_NOT, Tj_Trigger, Trojan_SE, n281, n2335, n2337, n2338, n2340,
         n2342, n2344, n2346, n2348, n2350, n2352, n2354, n2356, n2357, n2359,
         n2360, n2362, n2363, n2365, n2366, n2368, n2370, n2372, n2374, n2376,
         n2377, n2379, n2380, n2382, n2383, n2385, n2387, n2389, n2391, n2393,
         n2395, n2397, n2399, n2401, n2403, n2405, n2407, n2409, n2411, n2413,
         n2415, n2417, n2419, n2421, n2423, n2424, n2426, n2427, n2429, n2430,
         n2432, n2434, n2436, n2438, n2440, n2441, n2443, n2444, n2446, n2447,
         n2449, n2450, n2452, n2454, n2456, n2457, n2459, n2460, n2462, n2463,
         n2465, n2466, n2468, n2470, n2472, n2474, n2476, n2478, n2480, n2482,
         n2484, n2485, n2487, n2489, n2491, n2493, n2495, n2497, n2499, n2501,
         n2503, n2505, n2506, n2508, n2509, n2510, n2512, n2514, n2516, n2518,
         n2520, n2522, n2523, n2525, n2527, n2528, n2530, n2532, n2534, n2535,
         n2537, n2539, n2540, n2542, n2544, n2546, n2547, n2549, n2551, n2553,
         n2555, n2557, n2558, n2560, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2928, n2929, n2931, n2933, n2935, n2937, n2939, n2940, n2942, n2944,
         n2946, n2947, n2949, n2951, n2953, n2954, n2955, n2956, n2958, n2959,
         n2961, n2963, n2965, n2967, n2968, n2970, n2971, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2981, n2982, n2983, n2985, n2986, n2988,
         n2990, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3468, n3470, n3472, n3474, n3476, n3478,
         n3480, n3482, n3484, n3486, n3487, n3488, n3490, n3492, n3494, n3496,
         n3498, n3499, n3500, n3502, n3504, n3506, n3507, n3508, n3510, n3512,
         n3514, n3515, n3516, n3518, n3520, n3522, n3523, n3524, n3526, n3528,
         n3530, n3531, n3532, n3533, n3534, n3536, n3537, n3538, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3614, n3615,
         n3616, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3636, n3637, n3638,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3714,
         n3715, n3716, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3736,
         n3737, n3738, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, U3558_n1, U3871_n1, U3991_n1, U5716_n1, U5717_n1,
         U5718_n1, U5719_n1, U5720_n1, U5721_n1, U5722_n1, U5723_n1, U5724_n1,
         U5725_n1, U5726_n1, U5727_n1, U5728_n1, U5729_n1, U5730_n1, U5731_n1,
         U5732_n1, U5733_n1, U5734_n1, U5735_n1, U5736_n1, U5737_n1, U5738_n1,
         U5739_n1, U5740_n1, U5741_n1, U5742_n1, U5743_n1, U5744_n1, U5745_n1,
         U5746_n1, U5747_n1, U5748_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1,
         U5753_n1, U5754_n1, U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1,
         U5760_n1, U5761_n1, U5762_n1, U5763_n1, U5764_n1, U5765_n1, U5766_n1,
         U5767_n1, U5768_n1, U5769_n1, U5770_n1, U5771_n1, U5772_n1, U5773_n1,
         U5774_n1, U5775_n1, U5776_n1, U5777_n1, U5778_n1, U5779_n1, U5780_n1,
         U5781_n1, U5782_n1, U5783_n1, U5784_n1, U5785_n1, U5786_n1, U5787_n1,
         U5788_n1, U5789_n1, U5790_n1, U5791_n1, U5792_n1, U5793_n1, U5794_n1,
         U5795_n1, U5796_n1, U5797_n1, U5798_n1, U5799_n1, U5800_n1, U5801_n1,
         U5802_n1, U5803_n1, U5804_n1, U5805_n1, U5806_n1, U5807_n1, U5808_n1,
         U5809_n1, U5810_n1, U5811_n1, U5812_n1, U5813_n1, U5814_n1, U5815_n1,
         U5816_n1, U5817_n1, U5818_n1, U5819_n1, U5820_n1, U5821_n1, U5822_n1,
         U5823_n1, U5824_n1, U5825_n1, U5826_n1, U5827_n1, U5828_n1, U5829_n1,
         U5830_n1, U5831_n1, U5832_n1, U5833_n1, U5834_n1, U5835_n1, U5836_n1,
         U5837_n1, U5838_n1, U5839_n1, U5840_n1, U5841_n1, U5842_n1, U5843_n1,
         U5844_n1, U5845_n1, U5846_n1, U5847_n1, U5848_n1, U5849_n1, U5850_n1,
         U5851_n1, U5852_n1, U5853_n1, U5854_n1, U5855_n1, U5856_n1, U5857_n1,
         U5858_n1, U5859_n1, U5860_n1, U5861_n1, U5862_n1, U5863_n1, U5864_n1,
         U5865_n1, U5866_n1, U5867_n1, U5868_n1, U5869_n1, U5870_n1, U5871_n1,
         U5872_n1, U5873_n1, U5874_n1, U5875_n1, U5876_n1, U5877_n1, U5878_n1,
         U5879_n1, U5880_n1, U5881_n1, U5882_n1, U5883_n1, U5884_n1, U5885_n1,
         U5886_n1, U5887_n1, U5888_n1, U5889_n1, U5890_n1, U5891_n1, U5892_n1,
         U5893_n1, U5894_n1, U5895_n1, U5896_n1, U5897_n1, U5898_n1, U5899_n1,
         U5900_n1, U5901_n1, U5902_n1, U5903_n1, U5904_n1, U5905_n1, U5906_n1,
         U5907_n1, U5908_n1, U5909_n1, U5910_n1, U5911_n1, U5912_n1, U5913_n1,
         U5914_n1, U5915_n1, U5916_n1, U5917_n1, U5918_n1, U5919_n1, U5920_n1,
         U5921_n1, U5922_n1, U5923_n1, U5924_n1, U5925_n1, U5926_n1, U5927_n1,
         U5928_n1, U5929_n1, U5930_n1, U5931_n1, U5932_n1, U5933_n1, U5934_n1,
         U5935_n1, U5936_n1, U5937_n1, U5938_n1, U5939_n1, U5940_n1, U5941_n1,
         U5942_n1, U5943_n1, U5944_n1, U5945_n1, U5946_n1, U5947_n1, U5948_n1,
         U5949_n1, U5950_n1, U5951_n1, U5952_n1, U5953_n1, U5954_n1, U5955_n1,
         U5956_n1, U5957_n1, U5958_n1, U5959_n1, U5960_n1, U5961_n1, U5962_n1,
         U5963_n1, U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1, U5969_n1,
         U5970_n1, U5971_n1, U5972_n1, U5973_n1, U5974_n1, U5975_n1, U5976_n1,
         U5977_n1, U5978_n1, U5979_n1, U5980_n1, U5981_n1, U5982_n1, U5983_n1,
         U5984_n1, U5985_n1, U5986_n1, U5987_n1, U5988_n1, U5989_n1, U5990_n1,
         U5991_n1, U5992_n1, U5993_n1, U5994_n1, U5995_n1, U5996_n1, U5997_n1,
         U5998_n1, U5999_n1, U6000_n1, U6001_n1, U6002_n1, U6003_n1, U6004_n1,
         U6005_n1, U6006_n1, U6007_n1, U6008_n1, U6009_n1, U6010_n1, U6011_n1,
         U6012_n1, U6013_n1, U6014_n1, U6015_n1, U6016_n1, U6017_n1, U6018_n1,
         U6019_n1, U6020_n1, U6021_n1, U6022_n1, U6023_n1, U6024_n1, U6025_n1,
         U6026_n1, U6027_n1, U6028_n1, U6029_n1, U6030_n1, U6031_n1, U6032_n1,
         U6033_n1, U6034_n1, U6035_n1, U6036_n1, U6037_n1, U6038_n1, U6039_n1,
         U6040_n1, U6041_n1, U6042_n1, U6043_n1, U6044_n1, U6045_n1, U6046_n1,
         U6047_n1, U6048_n1, U6049_n1, U6050_n1, U6051_n1, U6052_n1, U6053_n1,
         U6054_n1, U6055_n1, U6056_n1, U6057_n1, U6058_n1, U6059_n1, U6060_n1,
         U6061_n1, U6062_n1, U6063_n1, U6064_n1, U6065_n1, U6066_n1, U6067_n1,
         U6068_n1, U6069_n1, U6070_n1, U6071_n1, U6072_n1, U6073_n1, U6074_n1,
         U6075_n1, U6076_n1, U6077_n1, U6078_n1, U6079_n1, U6080_n1, U6081_n1,
         U6082_n1, U6083_n1, U6084_n1, U6085_n1, U6086_n1, U6087_n1, U6088_n1,
         U6089_n1, U6090_n1, U6091_n1, U6092_n1, U6093_n1, U6094_n1, U6095_n1,
         U6096_n1, U6097_n1, U6098_n1, U6099_n1, U6100_n1, U6101_n1, U6102_n1,
         U6103_n1, U6104_n1, U6105_n1, U6106_n1, U6107_n1, U6108_n1, U6109_n1,
         U6110_n1, U6111_n1, U6112_n1, U6113_n1, U6114_n1, U6115_n1, U6116_n1,
         U6117_n1, U6118_n1, U6119_n1, U6120_n1, U6121_n1, U6122_n1, U6123_n1,
         U6124_n1, U6125_n1, U6126_n1, U6127_n1, U6128_n1, U6129_n1, U6130_n1,
         U6131_n1, U6132_n1, U6133_n1, U6134_n1, U6135_n1, U6136_n1, U6137_n1,
         U6138_n1, U6139_n1, U6140_n1, U6141_n1, U6142_n1, U6143_n1, U6144_n1,
         U6145_n1, U6146_n1, U6147_n1, U6148_n1, U6149_n1, U6150_n1, U6151_n1,
         U6152_n1, U6153_n1, U6154_n1, U6155_n1, U6156_n1, U6157_n1, U6158_n1,
         U6159_n1, U6160_n1, U6161_n1, U6162_n1, U6163_n1, U6164_n1, U6165_n1,
         U6166_n1, U6167_n1, U6168_n1, U6169_n1, U6170_n1, U6171_n1, U6172_n1,
         U6173_n1, U6174_n1, U6175_n1, U6176_n1, U6177_n1, U6178_n1, U6179_n1,
         U6180_n1, U6181_n1, U6182_n1, U6183_n1, U6184_n1, U6185_n1, U6186_n1,
         U6187_n1, U6188_n1, U6189_n1, U6190_n1, U6191_n1, U6192_n1, U6193_n1,
         U6194_n1, U6195_n1, U6196_n1, U6197_n1, U6198_n1, U6199_n1, U6200_n1,
         U6201_n1, U6202_n1, U6203_n1, U6204_n1, U6205_n1, U6206_n1, U6207_n1,
         U6208_n1, U6209_n1, U6210_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1,
         U6215_n1, U6216_n1, U6217_n1, U6218_n1, U6219_n1, U6220_n1, U6221_n1,
         U6222_n1, U6223_n1, U6224_n1, U6225_n1, U6226_n1, U6227_n1, U6228_n1,
         U6229_n1, U6230_n1, U6231_n1, U6232_n1, U6233_n1, U6234_n1, U6235_n1,
         U6236_n1, U6237_n1, U6238_n1, U6239_n1, U6240_n1, U6241_n1, U6242_n1,
         U6243_n1, U6244_n1, U6245_n1, U6246_n1, U6247_n1, U6248_n1, U6249_n1,
         U6250_n1, U6251_n1, U6252_n1, U6253_n1, U6254_n1, U6255_n1, U6256_n1,
         U6257_n1, U6258_n1, U6259_n1, U6260_n1, U6261_n1, U6262_n1, U6263_n1,
         U6264_n1, U6265_n1, U6266_n1, U6267_n1, U6268_n1, U6269_n1, U6270_n1,
         U6271_n1, U6272_n1, U6273_n1, U6274_n1, U6275_n1, U6276_n1, U6277_n1,
         U6278_n1, U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1,
         U6285_n1, U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1,
         U6292_n1, U6293_n1, U6294_n1, U6295_n1, U6296_n1, U6297_n1, U6298_n1,
         U6299_n1, U6300_n1, U6301_n1, U6302_n1, U6303_n1, U6304_n1, U6305_n1,
         U6306_n1, U6307_n1, U6308_n1, U6309_n1, U6310_n1, U6311_n1, U6312_n1,
         U6313_n1, U6314_n1, U6315_n1, U6316_n1, U6317_n1, U6318_n1, U6319_n1,
         U6320_n1, U6321_n1, U6322_n1, U6323_n1, U6324_n1, U6325_n1, U6326_n1,
         U6327_n1, U6328_n1, U6329_n1, U6330_n1, U6331_n1, U6332_n1, U6333_n1,
         U6334_n1, U6335_n1, U6336_n1, U6337_n1, U6338_n1, U6339_n1, U6340_n1,
         U6341_n1, U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1,
         U6348_n1, U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1,
         U6355_n1, U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1,
         U6362_n1, U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1,
         U6369_n1, U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1,
         U6376_n1, U6377_n1, U6378_n1, U6379_n1, U6380_n1, U6381_n1, U6382_n1,
         U6383_n1, U6384_n1, U6385_n1, U6386_n1, U6387_n1, U6388_n1, U6389_n1,
         U6390_n1, U6391_n1, U6392_n1, U6393_n1, U6394_n1, U6395_n1, U6396_n1,
         U6397_n1, U6398_n1, U6399_n1, U6400_n1, U6401_n1, U6402_n1, U6403_n1,
         U6404_n1, U6405_n1, U6406_n1, U6407_n1, U6408_n1, U6409_n1, U6410_n1,
         U6411_n1, U6412_n1, U6413_n1, U6414_n1, U6415_n1, U6416_n1, U6417_n1,
         U6418_n1, U6419_n1, U6420_n1, U6421_n1, U6422_n1, U6423_n1, U6424_n1,
         U6425_n1, U6426_n1, U6427_n1, U6428_n1, U6429_n1, U6430_n1, U6431_n1,
         U6432_n1, U6433_n1, U6434_n1, U6435_n1, U6436_n1, U6437_n1, U6438_n1,
         U6439_n1, U6440_n1, U6441_n1, U6442_n1, U6443_n1, U6444_n1, U6445_n1,
         U6446_n1, U6447_n1, U6448_n1, U6449_n1, U6450_n1, U6451_n1, U6452_n1,
         U6453_n1, U6454_n1, U6455_n1, U6456_n1, U6457_n1, U6458_n1, U6459_n1,
         U6460_n1, U6461_n1, U6462_n1, U6463_n1, U6464_n1, U6465_n1, U6466_n1,
         U6467_n1, U6468_n1, U6469_n1, U6470_n1, U6471_n1, U6472_n1, U6473_n1,
         U6474_n1, U6475_n1, U6476_n1, U6477_n1, U6478_n1, U6479_n1, U6480_n1,
         U6481_n1, U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n3393), .CLK(n3757), .Q(
        WX485) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n3388), .CLK(n3759), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n3388), .CLK(n3759), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n3388), .CLK(n3759), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n3388), .CLK(n3759), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n3389), .CLK(n3759), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n3389), .CLK(n3759), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n3389), .CLK(n3759), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n3389), .CLK(n3759), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n3389), .CLK(n3758), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n3389), .CLK(n3758), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n3390), .CLK(n3758), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n3390), .CLK(n3758), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n3390), .CLK(n3758), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(n3390), .CLK(n3758), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n3390), .CLK(n3758), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n3390), .CLK(n3758), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n3391), .CLK(n3758), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n3391), .CLK(n3758), .Q(
        WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n3391), .CLK(n3758), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n3391), .CLK(n3758), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(n3391), .CLK(n3757), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n3391), .CLK(n3757), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n3392), .CLK(n3757), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n3392), .CLK(n3757), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n3392), .CLK(n3757), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n3392), .CLK(n3757), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n3392), .CLK(n3757), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n3392), .CLK(n3757), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n3393), .CLK(n3757), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n3393), .CLK(n3757), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n3393), .CLK(n3757), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n3388), .CLK(n3759), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n3388), .CLK(n3759), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n3387), .CLK(n3759), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n3387), .CLK(n3759), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n3106), .CLK(n3903), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n3106), .CLK(n3903), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n3106), .CLK(n3903), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n3386), .CLK(n3760), .Q(
        WX659) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n3386), .CLK(n3760), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n3386), .CLK(n3760), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n3385), .CLK(n3760), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n3385), .CLK(n3761), .Q(
        WX667) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n3385), .CLK(n3761), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n3384), .CLK(n3761), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n3384), .CLK(n3761), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n3383), .CLK(n3761), .Q(
        WX675) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n3383), .CLK(n3762), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n3382), .CLK(n3762), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n3381), .CLK(n3762), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n3381), .CLK(n3764), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n3380), .CLK(n3764), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n3379), .CLK(n3764), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n3378), .CLK(n3765), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n3378), .CLK(n3765), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n3377), .CLK(n3765), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n3377), .CLK(n3766), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n3376), .CLK(n3766), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n3375), .CLK(n3766), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n3375), .CLK(n3767), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n3374), .CLK(n3767), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n3373), .CLK(n3767), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n3373), .CLK(n3768), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n3372), .CLK(n3768), .Q(
        WX709), .QN(n6223) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n3372), .CLK(n3768), .Q(
        WX711), .QN(n2926) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n3371), .CLK(n3769), .Q(
        WX713) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n3387), .CLK(n3760), .Q(
        WX715), .QN(n6226) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n3387), .CLK(n3760), .Q(
        WX717) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n3387), .CLK(n3760), .Q(
        WX719) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n3387), .CLK(n3760), .Q(
        WX721) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n3386), .CLK(n3760), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n3386), .CLK(n3760), .Q(
        WX725) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n3386), .CLK(n3760), .Q(
        WX727), .QN(n2965) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n3385), .CLK(n3760), .Q(
        WX729), .QN(n2971) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n3385), .CLK(n3761), .Q(
        WX731), .QN(n6232) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n3385), .CLK(n3761), .Q(
        WX733) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n3384), .CLK(n3761), .Q(
        WX735) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n3384), .CLK(n3761), .Q(
        WX737) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n3383), .CLK(n3762), .Q(
        WX739), .QN(n2958) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n3383), .CLK(n3762), .Q(
        WX741), .QN(n2968) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n3382), .CLK(n3762), .Q(
        WX743) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n3381), .CLK(n3762), .Q(
        WX745) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n3381), .CLK(n3764), .Q(
        WX747) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n3380), .CLK(n3764), .Q(
        WX749) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n3379), .CLK(n3764), .Q(
        WX751), .QN(n6241) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n3379), .CLK(n3765), .Q(
        WX753), .QN(n6219) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n3378), .CLK(n3765), .Q(
        WX755) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n3377), .CLK(n3765), .Q(
        WX757), .QN(n2983) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n3377), .CLK(n3766), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n3376), .CLK(n3766), .Q(
        WX761) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n3375), .CLK(n3766), .Q(
        WX763) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n3375), .CLK(n3767), .Q(
        WX765) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n3374), .CLK(n3767), .Q(
        WX767), .QN(n2981) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n3373), .CLK(n3767), .Q(
        WX769) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n3373), .CLK(n3768), .Q(
        WX771), .QN(n2988) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n3372), .CLK(n3768), .Q(
        WX773), .QN(n2977) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n3371), .CLK(n3768), .Q(
        WX775) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n3371), .CLK(n3769), .Q(
        WX777), .QN(n6225) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n3371), .CLK(n3769), .Q(
        WX779) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n3370), .CLK(n3769), .Q(
        WX781), .QN(n6227) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n3370), .CLK(n3769), .Q(
        WX783), .QN(n6228) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n3370), .CLK(n3769), .Q(
        WX785), .QN(n6229) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n3369), .CLK(n3769), .Q(
        WX787), .QN(n6230) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n3369), .CLK(n3770), .Q(
        WX789), .QN(n6231) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n3369), .CLK(n3770), .Q(
        WX791) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n3368), .CLK(n3770), .Q(
        WX793) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n3368), .CLK(n3770), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n3384), .CLK(n3761), 
        .Q(WX797), .QN(n6233) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n3384), .CLK(n3761), .Q(
        WX799), .QN(n6234) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n3383), .CLK(n3761), .Q(
        WX801), .QN(n6235) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n3383), .CLK(n3762), .Q(
        WX803), .QN(n6236) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n3382), .CLK(n3762), .Q(
        WX805) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n3382), .CLK(n3762), .Q(
        WX807), .QN(n6237) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n3381), .CLK(n3764), .Q(
        WX809), .QN(n6238) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n3380), .CLK(n3764), .Q(
        WX811), .QN(n6239) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n3380), .CLK(n3764), .Q(
        WX813), .QN(n6240) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n3379), .CLK(n3765), .Q(
        WX815) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n3379), .CLK(n3765), .Q(
        WX817), .QN(n2953) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n3378), .CLK(n3765), .Q(
        WX819), .QN(n6220) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n3377), .CLK(n3766), .Q(
        WX821) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n3376), .CLK(n3766), .Q(
        WX823), .QN(n2974) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n3376), .CLK(n3766), .Q(
        WX825), .QN(n6221) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n3375), .CLK(n3767), .Q(
        WX827), .QN(n6222) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n3374), .CLK(n3767), .Q(
        WX829), .QN(n6224) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n3374), .CLK(n3767), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n3373), .CLK(n3768), 
        .Q(WX833), .QN(n6242) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n3372), .CLK(n3768), .Q(
        WX835) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n3372), .CLK(n3768), .Q(
        WX837), .QN(n2978) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n3371), .CLK(n3768), .Q(
        WX839), .QN(n2928) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n3371), .CLK(n3769), .Q(
        WX841), .QN(n2933) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n3370), .CLK(n3769), .Q(
        WX843), .QN(n2939) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n3370), .CLK(n3769), .Q(
        WX845), .QN(n2942) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n3370), .CLK(n3769), .Q(
        WX847), .QN(n2944) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n3369), .CLK(n3769), .Q(
        WX849), .QN(n2949) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n3369), .CLK(n3770), .Q(
        WX851), .QN(n2955) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n3369), .CLK(n3770), .Q(
        WX853), .QN(n2956) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n3368), .CLK(n3770), .Q(
        WX855), .QN(n2967) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n3368), .CLK(n3770), .Q(
        WX857), .QN(n2973) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n3368), .CLK(n3770), .Q(
        WX859), .QN(n2976) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n3368), .CLK(n3770), .Q(
        WX861), .QN(n2931) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n3367), .CLK(n3770), .Q(
        WX863), .QN(n2940) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n3367), .CLK(n3770), .Q(
        WX865), .QN(n2947) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n3367), .CLK(n3771), .Q(
        test_so8) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n3382), .CLK(n3762), 
        .Q(WX869), .QN(n2970) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n3382), .CLK(n3762), .Q(
        WX871), .QN(n2979) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n3381), .CLK(n3764), .Q(
        WX873), .QN(n2935) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n3380), .CLK(n3764), .Q(
        WX875), .QN(n2951) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n3380), .CLK(n3764), .Q(
        WX877), .QN(n2986) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n3379), .CLK(n3765), .Q(
        WX879), .QN(n2946) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n3378), .CLK(n3765), .Q(
        WX881), .QN(n2954) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n3378), .CLK(n3765), .Q(
        WX883), .QN(n2959) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n3377), .CLK(n3766), .Q(
        WX885), .QN(n2985) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n3376), .CLK(n3766), .Q(
        WX887), .QN(n2975) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n3376), .CLK(n3766), .Q(
        WX889), .QN(n2961) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n3375), .CLK(n3767), .Q(
        WX891), .QN(n2963) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n3374), .CLK(n3767), .Q(
        WX893), .QN(n2929) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n3374), .CLK(n3767), .Q(
        WX895), .QN(n2982) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n3373), .CLK(n3768), .Q(
        WX897), .QN(n2937) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n3372), .CLK(n3768), .Q(
        WX899), .QN(n2990) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n3109), .CLK(n3902), .Q(
        CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n3109), .CLK(n3902), 
        .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n3109), .CLK(n3902), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n3109), .CLK(n3902), 
        .Q(CRC_OUT_9_3) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n3109), .CLK(n3902), 
        .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n3108), .CLK(n3902), 
        .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n3108), .CLK(n3902), 
        .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n3108), .CLK(n3902), 
        .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n3108), .CLK(n3902), 
        .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n3108), .CLK(n3902), 
        .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n3108), .CLK(n3902), 
        .Q(CRC_OUT_9_10) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n3107), .CLK(n3903), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n3107), .CLK(n3903), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n3107), .CLK(n3903), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n3107), .CLK(n3903), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n3107), .CLK(n3903), .Q(CRC_OUT_9_15), .QN(DFF_175_n1) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n3107), .CLK(n3903), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n3106), .CLK(n3903), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n3106), .CLK(n3903), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n3106), .CLK(n3903), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n3367), .CLK(n3771), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n3367), .CLK(n3771), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n3367), .CLK(n3771), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n3366), .CLK(n3771), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n3366), .CLK(n3771), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n3366), .CLK(n3771), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n3366), .CLK(n3771), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n3366), .CLK(n3771), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n3366), .CLK(n3771), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n3365), .CLK(n3771), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(n3365), .CLK(n3771), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n3365), .CLK(n3772), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(WX1777), .SI(CRC_OUT_9_31), .SE(n3365), .CLK(n3772), .Q(WX1778) );
  SDFFX1 DFF_193_Q_reg ( .D(WX1779), .SI(WX1778), .SE(n3360), .CLK(n3774), .Q(
        n8702) );
  SDFFX1 DFF_194_Q_reg ( .D(WX1781), .SI(n8702), .SE(n3360), .CLK(n3774), .Q(
        n8701) );
  SDFFX1 DFF_195_Q_reg ( .D(WX1783), .SI(n8701), .SE(n3360), .CLK(n3774), .Q(
        n8700) );
  SDFFX1 DFF_196_Q_reg ( .D(WX1785), .SI(n8700), .SE(n3360), .CLK(n3774), .Q(
        n8699) );
  SDFFX1 DFF_197_Q_reg ( .D(WX1787), .SI(n8699), .SE(n3360), .CLK(n3774), .Q(
        test_so11) );
  SDFFX1 DFF_198_Q_reg ( .D(WX1789), .SI(test_si12), .SE(n3361), .CLK(n3774), 
        .Q(n8696) );
  SDFFX1 DFF_199_Q_reg ( .D(WX1791), .SI(n8696), .SE(n3361), .CLK(n3774), .Q(
        n8695) );
  SDFFX1 DFF_200_Q_reg ( .D(WX1793), .SI(n8695), .SE(n3361), .CLK(n3774), .Q(
        n8694) );
  SDFFX1 DFF_201_Q_reg ( .D(WX1795), .SI(n8694), .SE(n3361), .CLK(n3774), .Q(
        n8693) );
  SDFFX1 DFF_202_Q_reg ( .D(WX1797), .SI(n8693), .SE(n3361), .CLK(n3773), .Q(
        n8692) );
  SDFFX1 DFF_203_Q_reg ( .D(WX1799), .SI(n8692), .SE(n3361), .CLK(n3773), .Q(
        n8691) );
  SDFFX1 DFF_204_Q_reg ( .D(WX1801), .SI(n8691), .SE(n3362), .CLK(n3773), .Q(
        n8690) );
  SDFFX1 DFF_205_Q_reg ( .D(WX1803), .SI(n8690), .SE(n3362), .CLK(n3773), .Q(
        n8689) );
  SDFFX1 DFF_206_Q_reg ( .D(WX1805), .SI(n8689), .SE(n3362), .CLK(n3773), .Q(
        n8688) );
  SDFFX1 DFF_207_Q_reg ( .D(WX1807), .SI(n8688), .SE(n3362), .CLK(n3773), .Q(
        n8687) );
  SDFFX1 DFF_208_Q_reg ( .D(WX1809), .SI(n8687), .SE(n3362), .CLK(n3773), .Q(
        n8686) );
  SDFFX1 DFF_209_Q_reg ( .D(WX1811), .SI(n8686), .SE(n3362), .CLK(n3773), .Q(
        n8685) );
  SDFFX1 DFF_210_Q_reg ( .D(WX1813), .SI(n8685), .SE(n3363), .CLK(n3773), .Q(
        n8684) );
  SDFFX1 DFF_211_Q_reg ( .D(WX1815), .SI(n8684), .SE(n3363), .CLK(n3773), .Q(
        n8683) );
  SDFFX1 DFF_212_Q_reg ( .D(WX1817), .SI(n8683), .SE(n3363), .CLK(n3773), .Q(
        n8682) );
  SDFFX1 DFF_213_Q_reg ( .D(WX1819), .SI(n8682), .SE(n3363), .CLK(n3773), .Q(
        n8681) );
  SDFFX1 DFF_214_Q_reg ( .D(WX1821), .SI(n8681), .SE(n3363), .CLK(n3772), .Q(
        n8680) );
  SDFFX1 DFF_215_Q_reg ( .D(WX1823), .SI(n8680), .SE(n3363), .CLK(n3772), .Q(
        test_so12) );
  SDFFX1 DFF_216_Q_reg ( .D(WX1825), .SI(test_si13), .SE(n3364), .CLK(n3772), 
        .Q(n8677) );
  SDFFX1 DFF_217_Q_reg ( .D(WX1827), .SI(n8677), .SE(n3364), .CLK(n3772), .Q(
        n8676) );
  SDFFX1 DFF_218_Q_reg ( .D(WX1829), .SI(n8676), .SE(n3364), .CLK(n3772), .Q(
        n8675) );
  SDFFX1 DFF_219_Q_reg ( .D(WX1831), .SI(n8675), .SE(n3364), .CLK(n3772), .Q(
        n8674) );
  SDFFX1 DFF_220_Q_reg ( .D(WX1833), .SI(n8674), .SE(n3364), .CLK(n3772), .Q(
        n8673) );
  SDFFX1 DFF_221_Q_reg ( .D(WX1835), .SI(n8673), .SE(n3364), .CLK(n3772), .Q(
        n8672) );
  SDFFX1 DFF_222_Q_reg ( .D(WX1837), .SI(n8672), .SE(n3365), .CLK(n3772), .Q(
        n8671) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n3365), .CLK(n3772), .Q(
        n8670) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n3360), .CLK(n3774), .Q(
        n8669), .QN(n6189) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n3359), .CLK(n3776), .Q(
        n8668), .QN(n6188) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n3359), .CLK(n3776), .Q(
        n8667), .QN(n6186) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n3358), .CLK(n3776), .Q(
        n8666), .QN(n6184) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n3358), .CLK(n3776), .Q(
        n8665), .QN(n6182) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n3356), .CLK(n3777), .Q(
        n8664), .QN(n6180) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n3356), .CLK(n3777), .Q(
        n8663), .QN(n6178) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n3355), .CLK(n3778), .Q(
        n8662), .QN(n6176) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n3355), .CLK(n3778), .Q(
        n8661), .QN(n6174) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n3109), .CLK(n3902), .Q(
        test_so13) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n3353), .CLK(n3778), 
        .Q(n8658), .QN(n6170) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n3353), .CLK(n3779), .Q(
        n8657), .QN(n6168) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n3352), .CLK(n3779), .Q(
        n8656), .QN(n6166) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n3352), .CLK(n3779), .Q(
        n8655), .QN(n6164) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n3117), .CLK(n3898), .Q(
        n8654), .QN(n6162) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n3117), .CLK(n3898), .Q(
        n8653), .QN(n6160) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n3350), .CLK(n3780), .Q(
        WX1970), .QN(n2675) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n3350), .CLK(n3780), .Q(
        WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n3350), .CLK(n3780), .Q(
        WX1974), .QN(n2674) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n3350), .CLK(n3780), .Q(
        WX1976), .QN(n2673) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n3349), .CLK(n3780), .Q(
        WX1978), .QN(n2672) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n3349), .CLK(n3780), .Q(
        WX1980) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n3349), .CLK(n3781), .Q(
        WX1982), .QN(n2670) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n3349), .CLK(n3781), .Q(
        WX1984), .QN(n2669) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n3349), .CLK(n3781), .Q(
        WX1986), .QN(n2668) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n3349), .CLK(n3781), .Q(
        WX1988), .QN(n2667) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n3348), .CLK(n3781), .Q(
        WX1990), .QN(n2666) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n3348), .CLK(n3781), .Q(
        test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n3110), .CLK(n3901), 
        .Q(WX1994), .QN(n2665) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n3110), .CLK(n3901), .Q(
        WX1996), .QN(n2664) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n3110), .CLK(n3901), .Q(
        WX1998), .QN(n2663) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n3110), .CLK(n3901), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n3359), .CLK(n3774), .Q(
        WX2002), .QN(n2348) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n3359), .CLK(n3776), .Q(
        WX2004), .QN(n2560) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n3358), .CLK(n3776), .Q(
        WX2006), .QN(n2558) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n3358), .CLK(n3776), .Q(
        WX2008), .QN(n2557) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n3357), .CLK(n3776), .Q(
        WX2010), .QN(n2555) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n3357), .CLK(n3777), .Q(
        WX2012), .QN(n2553) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n3356), .CLK(n3777), .Q(
        WX2014), .QN(n2551) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n3356), .CLK(n3777), .Q(
        WX2016), .QN(n2549) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n3355), .CLK(n3778), .Q(
        WX2018), .QN(n2547) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n3354), .CLK(n3778), .Q(
        WX2020), .QN(n2546) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n3354), .CLK(n3778), .Q(
        WX2022), .QN(n2544) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n3353), .CLK(n3779), .Q(
        WX2024), .QN(n2542) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n3352), .CLK(n3779), .Q(
        WX2026), .QN(n2540) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n3352), .CLK(n3779), .Q(
        test_so15) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n3117), .CLK(n3898), 
        .Q(WX2030), .QN(n2537) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n3117), .CLK(n3898), .Q(
        WX2032), .QN(n2535) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n3117), .CLK(n3898), .Q(
        WX2034) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n3117), .CLK(n3898), .Q(
        WX2036), .QN(n3783) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n3116), .CLK(n3898), .Q(
        WX2038) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n3116), .CLK(n3898), .Q(
        WX2040) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n3115), .CLK(n3899), .Q(
        WX2042) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n3115), .CLK(n3899), .Q(
        WX2044), .QN(n3775) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n3114), .CLK(n3899), .Q(
        WX2046) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n3114), .CLK(n3899), .Q(
        WX2048) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n3113), .CLK(n3900), .Q(
        WX2050) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n3113), .CLK(n3900), .Q(
        WX2052) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n3112), .CLK(n3900), .Q(
        WX2054) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n3348), .CLK(n3781), .Q(
        WX2056), .QN(n3763) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n3348), .CLK(n3781), .Q(
        WX2058) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n3348), .CLK(n3781), .Q(
        WX2060) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n3348), .CLK(n3781), .Q(
        WX2062) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n3347), .CLK(n3781), .Q(
        test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n3359), .CLK(n3774), 
        .Q(WX2066) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n3359), .CLK(n3776), .Q(
        WX2068) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n3358), .CLK(n3776), .Q(
        WX2070) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n3358), .CLK(n3776), .Q(
        WX2072) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n3357), .CLK(n3776), .Q(
        WX2074) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n3357), .CLK(n3777), .Q(
        WX2076) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n3356), .CLK(n3777), .Q(
        WX2078) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n3355), .CLK(n3777), .Q(
        WX2080) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n3355), .CLK(n3778), .Q(
        WX2082) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n3354), .CLK(n3778), .Q(
        WX2084), .QN(n6172) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n3354), .CLK(n3778), .Q(
        WX2086) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n3353), .CLK(n3779), .Q(
        WX2088) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n3352), .CLK(n3779), .Q(
        WX2090) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n3351), .CLK(n3779), .Q(
        WX2092), .QN(n2539) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n3351), .CLK(n3780), .Q(
        WX2094) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n3351), .CLK(n3780), .Q(
        WX2096) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n3350), .CLK(n3780), .Q(
        WX2098), .QN(n6158) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n3116), .CLK(n3898), .Q(
        test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n3116), .CLK(n3898), 
        .Q(WX2102), .QN(n6155) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n3115), .CLK(n3899), .Q(
        WX2104), .QN(n6153) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n3115), .CLK(n3899), .Q(
        WX2106), .QN(n6152) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n3114), .CLK(n3899), .Q(
        WX2108), .QN(n2671) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n3114), .CLK(n3899), .Q(
        WX2110), .QN(n6149) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n3113), .CLK(n3900), .Q(
        WX2112), .QN(n6147) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n3113), .CLK(n3900), .Q(
        WX2114), .QN(n6146) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n3112), .CLK(n3900), .Q(
        WX2116), .QN(n6144) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n3112), .CLK(n3900), .Q(
        WX2118), .QN(n6143) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n3112), .CLK(n3900), .Q(
        WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n3111), .CLK(n3901), .Q(
        WX2122), .QN(n6140) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n3111), .CLK(n3901), .Q(
        WX2124), .QN(n6138) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n3111), .CLK(n3901), .Q(
        WX2126), .QN(n6136) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n3347), .CLK(n3781), .Q(
        WX2128), .QN(n2662) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n3347), .CLK(n3782), .Q(
        WX2130), .QN(n2900) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n3347), .CLK(n3782), .Q(
        WX2132), .QN(n2901) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n3347), .CLK(n3782), .Q(
        WX2134), .QN(n2902) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n3347), .CLK(n3782), .Q(
        test_so18) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n3357), .CLK(n3777), 
        .Q(WX2138), .QN(n2903) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n3357), .CLK(n3777), .Q(
        WX2140), .QN(n2904) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n3356), .CLK(n3777), .Q(
        WX2142), .QN(n2905) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n3355), .CLK(n3777), .Q(
        WX2144), .QN(n2906) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n3354), .CLK(n3778), .Q(
        WX2146), .QN(n2907) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n3354), .CLK(n3778), .Q(
        WX2148), .QN(n2908) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n3353), .CLK(n3778), .Q(
        WX2150), .QN(n2909) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n3353), .CLK(n3779), .Q(
        WX2152), .QN(n2910) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n3352), .CLK(n3779), .Q(
        WX2154), .QN(n2911) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n3351), .CLK(n3779), .Q(
        WX2156), .QN(n2912) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n3351), .CLK(n3780), .Q(
        WX2158), .QN(n2913) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n3351), .CLK(n3780), .Q(
        WX2160), .QN(n2703) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n3350), .CLK(n3780), .Q(
        WX2162), .QN(n2914) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n3116), .CLK(n3898), .Q(
        WX2164), .QN(n2915) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n3116), .CLK(n3898), .Q(
        WX2166), .QN(n2916) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n3115), .CLK(n3899), .Q(
        WX2168), .QN(n2917) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n3115), .CLK(n3899), .Q(
        WX2170), .QN(n2704) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n3114), .CLK(n3899), .Q(
        test_so19) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n3114), .CLK(n3899), 
        .Q(WX2174), .QN(n2918) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n3113), .CLK(n3900), .Q(
        WX2176), .QN(n2919) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n3113), .CLK(n3900), .Q(
        WX2178), .QN(n2920) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n3112), .CLK(n3900), .Q(
        WX2180), .QN(n2921) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n3112), .CLK(n3900), .Q(
        WX2182), .QN(n2922) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n3111), .CLK(n3901), .Q(
        WX2184), .QN(n2705) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n3111), .CLK(n3901), .Q(
        WX2186), .QN(n2923) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n3111), .CLK(n3901), .Q(
        WX2188), .QN(n2924) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n3110), .CLK(n3901), .Q(
        WX2190), .QN(n2925) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n3110), .CLK(n3901), .Q(
        WX2192), .QN(n2713) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n3123), .CLK(n3895), .Q(
        CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n3122), .CLK(n3895), 
        .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n3122), .CLK(n3895), 
        .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n3122), .CLK(n3895), 
        .Q(CRC_OUT_8_3) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n3122), .CLK(n3895), 
        .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n3122), .CLK(n3895), 
        .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n3122), .CLK(n3895), 
        .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n3121), .CLK(n3896), 
        .Q(test_so20) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n3121), .CLK(n3896), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n3121), .CLK(n3896), 
        .Q(CRC_OUT_8_9) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n3121), .CLK(n3896), 
        .Q(CRC_OUT_8_10) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n3121), .CLK(n3896), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n3121), .CLK(n3896), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n3120), .CLK(n3896), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n3120), .CLK(n3896), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n3120), .CLK(n3896), .Q(CRC_OUT_8_15) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n3120), .CLK(n3896), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n3120), .CLK(n3896), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n3120), .CLK(n3896), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n3119), .CLK(n3897), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n3119), .CLK(n3897), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n3119), .CLK(n3897), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n3119), .CLK(n3897), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n3119), .CLK(n3897), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n3119), .CLK(n3897), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n3118), .CLK(n3897), .Q(test_so21) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n3118), .CLK(n3897), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n3118), .CLK(n3897), .Q(CRC_OUT_8_27) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n3118), .CLK(n3897), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n3118), .CLK(n3897), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n3118), .CLK(n3897), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n3346), .CLK(n3782), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(WX3070), .SI(CRC_OUT_8_31), .SE(n3346), .CLK(n3782), .Q(WX3071) );
  SDFFX1 DFF_385_Q_reg ( .D(WX3072), .SI(WX3071), .SE(n3341), .CLK(n3786), .Q(
        n8644) );
  SDFFX1 DFF_386_Q_reg ( .D(WX3074), .SI(n8644), .SE(n3341), .CLK(n3785), .Q(
        n8643) );
  SDFFX1 DFF_387_Q_reg ( .D(WX3076), .SI(n8643), .SE(n3341), .CLK(n3785), .Q(
        n8642) );
  SDFFX1 DFF_388_Q_reg ( .D(WX3078), .SI(n8642), .SE(n3342), .CLK(n3785), .Q(
        n8641) );
  SDFFX1 DFF_389_Q_reg ( .D(WX3080), .SI(n8641), .SE(n3342), .CLK(n3785), .Q(
        n8640) );
  SDFFX1 DFF_390_Q_reg ( .D(WX3082), .SI(n8640), .SE(n3342), .CLK(n3785), .Q(
        n8639) );
  SDFFX1 DFF_391_Q_reg ( .D(WX3084), .SI(n8639), .SE(n3342), .CLK(n3785), .Q(
        n8638) );
  SDFFX1 DFF_392_Q_reg ( .D(WX3086), .SI(n8638), .SE(n3342), .CLK(n3785), .Q(
        n8637) );
  SDFFX1 DFF_393_Q_reg ( .D(WX3088), .SI(n8637), .SE(n3342), .CLK(n3785), .Q(
        n8636) );
  SDFFX1 DFF_394_Q_reg ( .D(WX3090), .SI(n8636), .SE(n3343), .CLK(n3785), .Q(
        n8635) );
  SDFFX1 DFF_395_Q_reg ( .D(WX3092), .SI(n8635), .SE(n3343), .CLK(n3785), .Q(
        test_so22) );
  SDFFX1 DFF_396_Q_reg ( .D(WX3094), .SI(test_si23), .SE(n3343), .CLK(n3785), 
        .Q(n8632) );
  SDFFX1 DFF_397_Q_reg ( .D(WX3096), .SI(n8632), .SE(n3343), .CLK(n3785), .Q(
        n8631) );
  SDFFX1 DFF_398_Q_reg ( .D(WX3098), .SI(n8631), .SE(n3343), .CLK(n3784), .Q(
        n8630) );
  SDFFX1 DFF_399_Q_reg ( .D(WX3100), .SI(n8630), .SE(n3343), .CLK(n3784), .Q(
        n8629) );
  SDFFX1 DFF_400_Q_reg ( .D(WX3102), .SI(n8629), .SE(n3344), .CLK(n3784), .Q(
        n8628) );
  SDFFX1 DFF_401_Q_reg ( .D(WX3104), .SI(n8628), .SE(n3344), .CLK(n3784), .Q(
        n8627) );
  SDFFX1 DFF_402_Q_reg ( .D(WX3106), .SI(n8627), .SE(n3344), .CLK(n3784), .Q(
        n8626) );
  SDFFX1 DFF_403_Q_reg ( .D(WX3108), .SI(n8626), .SE(n3344), .CLK(n3784), .Q(
        n8625) );
  SDFFX1 DFF_404_Q_reg ( .D(WX3110), .SI(n8625), .SE(n3344), .CLK(n3784), .Q(
        n8624) );
  SDFFX1 DFF_405_Q_reg ( .D(WX3112), .SI(n8624), .SE(n3344), .CLK(n3784), .Q(
        n8623) );
  SDFFX1 DFF_406_Q_reg ( .D(WX3114), .SI(n8623), .SE(n3345), .CLK(n3784), .Q(
        n8622) );
  SDFFX1 DFF_407_Q_reg ( .D(WX3116), .SI(n8622), .SE(n3345), .CLK(n3784), .Q(
        n8621) );
  SDFFX1 DFF_408_Q_reg ( .D(WX3118), .SI(n8621), .SE(n3345), .CLK(n3784), .Q(
        n8620) );
  SDFFX1 DFF_409_Q_reg ( .D(WX3120), .SI(n8620), .SE(n3345), .CLK(n3784), .Q(
        n8619) );
  SDFFX1 DFF_410_Q_reg ( .D(WX3122), .SI(n8619), .SE(n3345), .CLK(n3782), .Q(
        n8618) );
  SDFFX1 DFF_411_Q_reg ( .D(WX3124), .SI(n8618), .SE(n3345), .CLK(n3782), .Q(
        n8617) );
  SDFFX1 DFF_412_Q_reg ( .D(WX3126), .SI(n8617), .SE(n3346), .CLK(n3782), .Q(
        n8616) );
  SDFFX1 DFF_413_Q_reg ( .D(WX3128), .SI(n8616), .SE(n3346), .CLK(n3782), .Q(
        test_so23) );
  SDFFX1 DFF_414_Q_reg ( .D(WX3130), .SI(test_si24), .SE(n3346), .CLK(n3782), 
        .Q(n8613) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n3346), .CLK(n3782), .Q(
        n8612) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n3341), .CLK(n3786), .Q(
        n8611), .QN(n6190) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n3340), .CLK(n3786), .Q(
        n8610), .QN(n6187) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n3340), .CLK(n3786), .Q(
        n8609), .QN(n6185) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n3340), .CLK(n3786), .Q(
        n8608), .QN(n6183) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n3340), .CLK(n3786), .Q(
        n8607), .QN(n6181) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n3339), .CLK(n3787), .Q(
        n8606), .QN(n6179) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n3339), .CLK(n3787), .Q(
        n8605), .QN(n6177) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n3338), .CLK(n3787), .Q(
        n8604), .QN(n6175) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n3338), .CLK(n3787), .Q(
        n8603), .QN(n6173) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n3337), .CLK(n3788), .Q(
        n8602), .QN(n6171) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n3337), .CLK(n3788), .Q(
        n8601), .QN(n6169) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n3336), .CLK(n3788), .Q(
        n8600), .QN(n6167) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n3335), .CLK(n3788), .Q(
        n8599), .QN(n6165) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n3334), .CLK(n3789), .Q(
        n8598), .QN(n6163) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n3334), .CLK(n3789), .Q(
        n8597), .QN(n6161) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n3123), .CLK(n3895), .Q(
        test_so24) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n3125), .CLK(n3894), 
        .Q(WX3263), .QN(n2661) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n3123), .CLK(n3895), .Q(
        WX3265), .QN(n2660) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n3123), .CLK(n3895), .Q(
        WX3267), .QN(n2659) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n3331), .CLK(n3791), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n3331), .CLK(n3791), .Q(
        WX3271), .QN(n2657) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n3330), .CLK(n3791), .Q(
        WX3273), .QN(n2656) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n3329), .CLK(n3791), .Q(
        WX3275), .QN(n2655) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n3329), .CLK(n3792), .Q(
        WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n3328), .CLK(n3792), .Q(
        WX3279), .QN(n2654) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n3327), .CLK(n3792), .Q(
        WX3281) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n3327), .CLK(n3793), .Q(
        WX3283), .QN(n2652) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n3326), .CLK(n3793), .Q(
        WX3285), .QN(n2651) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n3325), .CLK(n3793), .Q(
        WX3287), .QN(n2650) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n3325), .CLK(n3794), .Q(
        WX3289), .QN(n2649) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n3324), .CLK(n3794), .Q(
        WX3291), .QN(n2648) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n3323), .CLK(n3794), .Q(
        WX3293), .QN(n2647) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n3341), .CLK(n3786), .Q(
        WX3295), .QN(n2346) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n3341), .CLK(n3786), .Q(
        test_so25) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n3340), .CLK(n3786), 
        .Q(WX3299), .QN(n2532) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n3340), .CLK(n3786), .Q(
        WX3301), .QN(n2530) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n3339), .CLK(n3786), .Q(
        WX3303), .QN(n2528) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n3339), .CLK(n3786), .Q(
        WX3305), .QN(n2527) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n3339), .CLK(n3787), .Q(
        WX3307), .QN(n2525) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n3338), .CLK(n3787), .Q(
        WX3309), .QN(n2523) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n3338), .CLK(n3787), .Q(
        WX3311), .QN(n2522) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n3337), .CLK(n3787), .Q(
        WX3313), .QN(n2520) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n3337), .CLK(n3788), .Q(
        WX3315), .QN(n2518) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n3336), .CLK(n3788), .Q(
        WX3317), .QN(n2516) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n3335), .CLK(n3788), .Q(
        WX3319), .QN(n2514) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n3335), .CLK(n3789), .Q(
        WX3321), .QN(n2512) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n3334), .CLK(n3789), .Q(
        WX3323), .QN(n2510) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n3333), .CLK(n3789), .Q(
        WX3325), .QN(n2509) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n3333), .CLK(n3790), .Q(
        WX3327) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n3332), .CLK(n3790), .Q(
        WX3329) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n3332), .CLK(n3790), .Q(
        WX3331) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n3331), .CLK(n3790), .Q(
        test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n3331), .CLK(n3791), 
        .Q(WX3335) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n3330), .CLK(n3791), .Q(
        WX3337) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n3329), .CLK(n3791), .Q(
        WX3339) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n3329), .CLK(n3792), .Q(
        WX3341), .QN(n3739) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n3328), .CLK(n3792), .Q(
        WX3343) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n3327), .CLK(n3792), .Q(
        WX3345), .QN(n3735) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n3327), .CLK(n3793), .Q(
        WX3347) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n3326), .CLK(n3793), .Q(
        WX3349) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n3325), .CLK(n3793), .Q(
        WX3351) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n3325), .CLK(n3794), .Q(
        WX3353) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n3324), .CLK(n3794), .Q(
        WX3355) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n3323), .CLK(n3794), .Q(
        WX3357) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n3323), .CLK(n3795), .Q(
        WX3359) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n3322), .CLK(n3795), .Q(
        WX3361), .QN(n2534) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n3322), .CLK(n3795), .Q(
        WX3363) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n3322), .CLK(n3795), .Q(
        WX3365) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n3321), .CLK(n3795), .Q(
        WX3367) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n3321), .CLK(n3796), .Q(
        test_so27) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n3339), .CLK(n3787), 
        .Q(WX3371) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n3338), .CLK(n3787), .Q(
        WX3373) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n3338), .CLK(n3787), .Q(
        WX3375) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n3337), .CLK(n3787), .Q(
        WX3377) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n3336), .CLK(n3788), .Q(
        WX3379) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n3336), .CLK(n3788), .Q(
        WX3381) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n3335), .CLK(n3789), .Q(
        WX3383) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n3335), .CLK(n3789), .Q(
        WX3385) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n3334), .CLK(n3789), .Q(
        WX3387) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n3333), .CLK(n3789), .Q(
        WX3389), .QN(n6159) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n3333), .CLK(n3790), .Q(
        WX3391), .QN(n6157) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n3332), .CLK(n3790), .Q(
        WX3393), .QN(n6156) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n3332), .CLK(n3790), .Q(
        WX3395), .QN(n6154) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n3331), .CLK(n3790), .Q(
        WX3397), .QN(n2658) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n3330), .CLK(n3791), .Q(
        WX3399), .QN(n6151) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n3330), .CLK(n3791), .Q(
        WX3401), .QN(n6150) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n3329), .CLK(n3792), .Q(
        WX3403), .QN(n6148) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n3328), .CLK(n3792), .Q(
        test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n3328), .CLK(n3792), 
        .Q(WX3407), .QN(n6145) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n3327), .CLK(n3793), .Q(
        WX3409), .QN(n2653) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n3326), .CLK(n3793), .Q(
        WX3411), .QN(n6142) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n3326), .CLK(n3793), .Q(
        WX3413), .QN(n6141) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n3325), .CLK(n3794), .Q(
        WX3415), .QN(n6139) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n3324), .CLK(n3794), .Q(
        WX3417), .QN(n6137) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n3324), .CLK(n3794), .Q(
        WX3419), .QN(n6135) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n3323), .CLK(n3795), .Q(
        WX3421), .QN(n6134) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n3323), .CLK(n3795), .Q(
        WX3423), .QN(n2874) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n3322), .CLK(n3795), .Q(
        WX3425), .QN(n2875) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n3322), .CLK(n3795), .Q(
        WX3427), .QN(n2876) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n3322), .CLK(n3795), .Q(
        WX3429), .QN(n2877) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n3321), .CLK(n3795), .Q(
        WX3431), .QN(n2878) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n3321), .CLK(n3796), .Q(
        WX3433), .QN(n2879) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n3321), .CLK(n3796), .Q(
        WX3435), .QN(n2880) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n3321), .CLK(n3796), .Q(
        WX3437), .QN(n2881) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n3320), .CLK(n3796), .Q(
        test_so29) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n3337), .CLK(n3788), 
        .Q(WX3441), .QN(n2882) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n3336), .CLK(n3788), .Q(
        WX3443), .QN(n2883) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n3336), .CLK(n3788), .Q(
        WX3445), .QN(n2884) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n3335), .CLK(n3789), .Q(
        WX3447), .QN(n2885) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n3334), .CLK(n3789), .Q(
        WX3449), .QN(n2886) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n3334), .CLK(n3789), .Q(
        WX3451), .QN(n2887) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n3333), .CLK(n3790), .Q(
        WX3453), .QN(n2700) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n3333), .CLK(n3790), .Q(
        WX3455), .QN(n2888) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n3332), .CLK(n3790), .Q(
        WX3457), .QN(n2889) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n3332), .CLK(n3790), .Q(
        WX3459), .QN(n2890) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n3331), .CLK(n3791), .Q(
        WX3461), .QN(n2891) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n3330), .CLK(n3791), .Q(
        WX3463), .QN(n2701) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n3330), .CLK(n3791), .Q(
        WX3465), .QN(n2892) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n3329), .CLK(n3792), .Q(
        WX3467), .QN(n2893) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n3328), .CLK(n3792), .Q(
        WX3469), .QN(n2894) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n3328), .CLK(n3792), .Q(
        WX3471), .QN(n2895) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n3327), .CLK(n3793), .Q(
        test_so30) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n3326), .CLK(n3793), 
        .Q(WX3475), .QN(n2896) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n3326), .CLK(n3793), .Q(
        WX3477), .QN(n2702) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n3325), .CLK(n3794), .Q(
        WX3479), .QN(n2897) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n3324), .CLK(n3794), .Q(
        WX3481), .QN(n2898) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n3324), .CLK(n3794), .Q(
        WX3483), .QN(n2899) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n3323), .CLK(n3795), .Q(
        WX3485), .QN(n2712) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n3128), .CLK(n3892), .Q(
        CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n3127), .CLK(n3893), 
        .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n3127), .CLK(n3893), 
        .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n3127), .CLK(n3893), 
        .Q(CRC_OUT_7_3) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n3127), .CLK(n3893), 
        .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n3127), .CLK(n3893), 
        .Q(CRC_OUT_7_5) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n3127), .CLK(n3893), 
        .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n3126), .CLK(n3893), 
        .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n3126), .CLK(n3893), 
        .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n3126), .CLK(n3893), 
        .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n3126), .CLK(n3893), 
        .Q(test_so31) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n3126), .CLK(n3893), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n3126), .CLK(n3893), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n3125), .CLK(n3894), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n3125), .CLK(n3894), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n3125), .CLK(n3894), .Q(CRC_OUT_7_15) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n3125), .CLK(n3894), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n3125), .CLK(n3894), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n3124), .CLK(n3894), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n3124), .CLK(n3894), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n3124), .CLK(n3894), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n3124), .CLK(n3894), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n3124), .CLK(n3894), .Q(CRC_OUT_7_22) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n3124), .CLK(n3894), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n3123), .CLK(n3895), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n3123), .CLK(n3895), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n3320), .CLK(n3796), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n3320), .CLK(n3796), .Q(test_so32) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n3320), .CLK(n3796), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n3320), .CLK(n3796), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n3320), .CLK(n3796), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n3319), .CLK(n3796), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(WX4363), .SI(CRC_OUT_7_31), .SE(n3319), .CLK(n3796), .Q(WX4364) );
  SDFFX1 DFF_577_Q_reg ( .D(WX4365), .SI(WX4364), .SE(n3314), .CLK(n3799), .Q(
        n8586) );
  SDFFX1 DFF_578_Q_reg ( .D(WX4367), .SI(n8586), .SE(n3314), .CLK(n3799), .Q(
        n8585) );
  SDFFX1 DFF_579_Q_reg ( .D(WX4369), .SI(n8585), .SE(n3314), .CLK(n3799), .Q(
        n8584) );
  SDFFX1 DFF_580_Q_reg ( .D(WX4371), .SI(n8584), .SE(n3315), .CLK(n3799), .Q(
        n8583) );
  SDFFX1 DFF_581_Q_reg ( .D(WX4373), .SI(n8583), .SE(n3315), .CLK(n3799), .Q(
        n8582) );
  SDFFX1 DFF_582_Q_reg ( .D(WX4375), .SI(n8582), .SE(n3315), .CLK(n3799), .Q(
        n8581) );
  SDFFX1 DFF_583_Q_reg ( .D(WX4377), .SI(n8581), .SE(n3315), .CLK(n3799), .Q(
        n8580) );
  SDFFX1 DFF_584_Q_reg ( .D(WX4379), .SI(n8580), .SE(n3315), .CLK(n3798), .Q(
        n8579) );
  SDFFX1 DFF_585_Q_reg ( .D(WX4381), .SI(n8579), .SE(n3315), .CLK(n3798), .Q(
        n8578) );
  SDFFX1 DFF_586_Q_reg ( .D(WX4383), .SI(n8578), .SE(n3316), .CLK(n3798), .Q(
        n8577) );
  SDFFX1 DFF_587_Q_reg ( .D(WX4385), .SI(n8577), .SE(n3316), .CLK(n3798), .Q(
        n8576) );
  SDFFX1 DFF_588_Q_reg ( .D(WX4387), .SI(n8576), .SE(n3316), .CLK(n3798), .Q(
        test_so33) );
  SDFFX1 DFF_589_Q_reg ( .D(WX4389), .SI(test_si34), .SE(n3316), .CLK(n3798), 
        .Q(n8573) );
  SDFFX1 DFF_590_Q_reg ( .D(WX4391), .SI(n8573), .SE(n3316), .CLK(n3798), .Q(
        n8572) );
  SDFFX1 DFF_591_Q_reg ( .D(WX4393), .SI(n8572), .SE(n3316), .CLK(n3798), .Q(
        n8571) );
  SDFFX1 DFF_592_Q_reg ( .D(WX4395), .SI(n8571), .SE(n3317), .CLK(n3798), .Q(
        n8570) );
  SDFFX1 DFF_593_Q_reg ( .D(WX4397), .SI(n8570), .SE(n3317), .CLK(n3798), .Q(
        n8569) );
  SDFFX1 DFF_594_Q_reg ( .D(WX4399), .SI(n8569), .SE(n3317), .CLK(n3798), .Q(
        n8568) );
  SDFFX1 DFF_595_Q_reg ( .D(WX4401), .SI(n8568), .SE(n3317), .CLK(n3798), .Q(
        n8567) );
  SDFFX1 DFF_596_Q_reg ( .D(WX4403), .SI(n8567), .SE(n3317), .CLK(n3797), .Q(
        n8566) );
  SDFFX1 DFF_597_Q_reg ( .D(WX4405), .SI(n8566), .SE(n3317), .CLK(n3797), .Q(
        n8565) );
  SDFFX1 DFF_598_Q_reg ( .D(WX4407), .SI(n8565), .SE(n3318), .CLK(n3797), .Q(
        n8564) );
  SDFFX1 DFF_599_Q_reg ( .D(WX4409), .SI(n8564), .SE(n3318), .CLK(n3797), .Q(
        n8563) );
  SDFFX1 DFF_600_Q_reg ( .D(WX4411), .SI(n8563), .SE(n3318), .CLK(n3797), .Q(
        n8562) );
  SDFFX1 DFF_601_Q_reg ( .D(WX4413), .SI(n8562), .SE(n3318), .CLK(n3797), .Q(
        n8561) );
  SDFFX1 DFF_602_Q_reg ( .D(WX4415), .SI(n8561), .SE(n3318), .CLK(n3797), .Q(
        n8560) );
  SDFFX1 DFF_603_Q_reg ( .D(WX4417), .SI(n8560), .SE(n3318), .CLK(n3797), .Q(
        n8559) );
  SDFFX1 DFF_604_Q_reg ( .D(WX4419), .SI(n8559), .SE(n3319), .CLK(n3797), .Q(
        n8558) );
  SDFFX1 DFF_605_Q_reg ( .D(WX4421), .SI(n8558), .SE(n3319), .CLK(n3797), .Q(
        test_so34) );
  SDFFX1 DFF_606_Q_reg ( .D(WX4423), .SI(test_si35), .SE(n3319), .CLK(n3797), 
        .Q(n8555) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n3319), .CLK(n3797), .Q(
        n8554) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n3314), .CLK(n3799), .Q(
        n8553), .QN(n6133) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n3313), .CLK(n3799), .Q(
        n8552), .QN(n6132) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n3313), .CLK(n3799), .Q(
        n8551), .QN(n6131) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n3312), .CLK(n3800), .Q(
        n8550), .QN(n6130) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n3312), .CLK(n3800), .Q(
        n8549), .QN(n6129) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n3311), .CLK(n3801), .Q(
        n8548), .QN(n6128) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n3311), .CLK(n3801), .Q(
        n8547), .QN(n6127) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n3310), .CLK(n3801), .Q(
        n8546), .QN(n6126) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n3310), .CLK(n3801), .Q(
        n8545), .QN(n6125) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n3308), .CLK(n3802), .Q(
        n8544), .QN(n6124) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n3308), .CLK(n3802), .Q(
        n8543), .QN(n6123) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n3307), .CLK(n3803), .Q(
        n8542), .QN(n6122) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n3307), .CLK(n3803), .Q(
        n8541), .QN(n6121) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n3306), .CLK(n3803), .Q(
        n8540), .QN(n6120) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n3306), .CLK(n3803), .Q(
        test_so35) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n3304), .CLK(n3804), 
        .Q(n8537), .QN(n6118) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n3304), .CLK(n3804), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n3304), .CLK(n3804), .Q(
        WX4558), .QN(n2645) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n3303), .CLK(n3805), .Q(
        WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n3302), .CLK(n3805), .Q(
        WX4562), .QN(n2644) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n3302), .CLK(n3805), .Q(
        WX4564) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n3301), .CLK(n3806), .Q(
        WX4566), .QN(n2642) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n3300), .CLK(n3806), .Q(
        WX4568), .QN(n2641) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n3300), .CLK(n3806), .Q(
        WX4570), .QN(n2640) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n3299), .CLK(n3807), .Q(
        WX4572), .QN(n2639) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n3298), .CLK(n3807), .Q(
        WX4574), .QN(n2638) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n3298), .CLK(n3807), .Q(
        WX4576), .QN(n2637) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n3297), .CLK(n3808), .Q(
        WX4578), .QN(n2636) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n3296), .CLK(n3808), .Q(
        WX4580), .QN(n2635) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n3296), .CLK(n3808), .Q(
        WX4582), .QN(n2634) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n3295), .CLK(n3809), .Q(
        WX4584), .QN(n2633) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n3294), .CLK(n3809), .Q(
        test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n3314), .CLK(n3799), 
        .Q(WX4588), .QN(n2344) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n3314), .CLK(n3799), .Q(
        WX4590), .QN(n2508) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n3313), .CLK(n3800), .Q(
        WX4592), .QN(n2506) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n3313), .CLK(n3800), .Q(
        WX4594), .QN(n2505) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n3312), .CLK(n3800), .Q(
        WX4596), .QN(n2503) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n3312), .CLK(n3800), .Q(
        WX4598), .QN(n2501) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n3311), .CLK(n3801), .Q(
        WX4600), .QN(n2499) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n3310), .CLK(n3801), .Q(
        WX4602), .QN(n2497) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n3309), .CLK(n3801), .Q(
        WX4604), .QN(n2495) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n3309), .CLK(n3802), .Q(
        WX4606), .QN(n2493) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n3308), .CLK(n3802), .Q(
        WX4608), .QN(n2491) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n3308), .CLK(n3802), .Q(
        WX4610), .QN(n2489) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n3307), .CLK(n3803), .Q(
        WX4612), .QN(n2487) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n3306), .CLK(n3803), .Q(
        WX4614), .QN(n2485) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n3305), .CLK(n3803), .Q(
        WX4616), .QN(n2484) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n3305), .CLK(n3804), .Q(
        WX4618), .QN(n2482) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n3304), .CLK(n3804), .Q(
        test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n3303), .CLK(n3804), 
        .Q(WX4622) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n3303), .CLK(n3805), .Q(
        WX4624), .QN(n3717) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n3302), .CLK(n3805), .Q(
        WX4626) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n3301), .CLK(n3805), .Q(
        WX4628), .QN(n3713) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n3301), .CLK(n3806), .Q(
        WX4630) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n3300), .CLK(n3806), .Q(
        WX4632) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n3299), .CLK(n3806), .Q(
        WX4634) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n3299), .CLK(n3807), .Q(
        WX4636) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n3298), .CLK(n3807), .Q(
        WX4638) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n3297), .CLK(n3807), .Q(
        WX4640) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n3297), .CLK(n3808), .Q(
        WX4642) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n3296), .CLK(n3808), .Q(
        WX4644) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n3295), .CLK(n3808), .Q(
        WX4646) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n3295), .CLK(n3809), .Q(
        WX4648) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n3294), .CLK(n3809), .Q(
        WX4650), .QN(n3691) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n3294), .CLK(n3809), .Q(
        WX4652) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n3293), .CLK(n3809), .Q(
        test_so38) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n3313), .CLK(n3800), 
        .Q(WX4656) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n3313), .CLK(n3800), .Q(
        WX4658) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n3312), .CLK(n3800), .Q(
        WX4660) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n3311), .CLK(n3800), .Q(
        WX4662) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n3311), .CLK(n3801), .Q(
        WX4664) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n3310), .CLK(n3801), .Q(
        WX4666) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n3309), .CLK(n3801), .Q(
        WX4668) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n3309), .CLK(n3802), .Q(
        WX4670) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n3308), .CLK(n3802), .Q(
        WX4672) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n3307), .CLK(n3802), .Q(
        WX4674) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n3307), .CLK(n3803), .Q(
        WX4676) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n3306), .CLK(n3803), .Q(
        WX4678) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n3305), .CLK(n3803), .Q(
        WX4680), .QN(n6119) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n3305), .CLK(n3804), .Q(
        WX4682) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n3304), .CLK(n3804), .Q(
        WX4684), .QN(n2646) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n3303), .CLK(n3804), .Q(
        WX4686), .QN(n6117) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n3303), .CLK(n3805), .Q(
        test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n3302), .CLK(n3805), 
        .Q(WX4690), .QN(n6116) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n3301), .CLK(n3805), .Q(
        WX4692), .QN(n2643) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n3301), .CLK(n3806), .Q(
        WX4694), .QN(n6115) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n3300), .CLK(n3806), .Q(
        WX4696), .QN(n6114) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n3299), .CLK(n3806), .Q(
        WX4698), .QN(n6113) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n3299), .CLK(n3807), .Q(
        WX4700), .QN(n6112) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n3298), .CLK(n3807), .Q(
        WX4702), .QN(n6111) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n3297), .CLK(n3807), .Q(
        WX4704), .QN(n6110) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n3297), .CLK(n3808), .Q(
        WX4706), .QN(n6109) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n3296), .CLK(n3808), .Q(
        WX4708), .QN(n6108) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n3295), .CLK(n3808), .Q(
        WX4710), .QN(n6107) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n3295), .CLK(n3809), .Q(
        WX4712), .QN(n6106) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n3294), .CLK(n3809), .Q(
        WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n3293), .CLK(n3809), .Q(
        WX4716), .QN(n2847) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n3293), .CLK(n3810), .Q(
        WX4718), .QN(n2848) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n3293), .CLK(n3810), .Q(
        WX4720), .QN(n2849) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n3293), .CLK(n3810), .Q(
        test_so40) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n3312), .CLK(n3800), 
        .Q(WX4724), .QN(n2850) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n3311), .CLK(n3800), .Q(
        WX4726), .QN(n2851) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n3310), .CLK(n3801), .Q(
        WX4728), .QN(n2852) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n3310), .CLK(n3801), .Q(
        WX4730), .QN(n2853) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n3309), .CLK(n3802), .Q(
        WX4732), .QN(n2854) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n3309), .CLK(n3802), .Q(
        WX4734), .QN(n2855) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n3308), .CLK(n3802), .Q(
        WX4736), .QN(n2856) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n3307), .CLK(n3802), .Q(
        WX4738), .QN(n2857) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n3306), .CLK(n3803), .Q(
        WX4740), .QN(n2858) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n3306), .CLK(n3803), .Q(
        WX4742), .QN(n2859) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n3305), .CLK(n3804), .Q(
        WX4744), .QN(n2860) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n3305), .CLK(n3804), .Q(
        WX4746), .QN(n2698) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n3304), .CLK(n3804), .Q(
        WX4748), .QN(n2861) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n3303), .CLK(n3805), .Q(
        WX4750), .QN(n2862) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n3302), .CLK(n3805), .Q(
        WX4752), .QN(n2863) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n3302), .CLK(n3805), .Q(
        WX4754), .QN(n2864) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n3301), .CLK(n3806), .Q(
        test_so41) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n3300), .CLK(n3806), 
        .Q(WX4758), .QN(n2865) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n3300), .CLK(n3806), .Q(
        WX4760), .QN(n2866) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n3299), .CLK(n3807), .Q(
        WX4762), .QN(n2867) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n3298), .CLK(n3807), .Q(
        WX4764), .QN(n2868) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n3298), .CLK(n3807), .Q(
        WX4766), .QN(n2869) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n3297), .CLK(n3808), .Q(
        WX4768), .QN(n2870) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n3296), .CLK(n3808), .Q(
        WX4770), .QN(n2699) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n3296), .CLK(n3808), .Q(
        WX4772), .QN(n2871) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n3295), .CLK(n3809), .Q(
        WX4774), .QN(n2872) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n3294), .CLK(n3809), .Q(
        WX4776), .QN(n2873) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n3294), .CLK(n3809), .Q(
        WX4778), .QN(n2711) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n3133), .CLK(n3890), .Q(
        CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n3132), .CLK(n3890), 
        .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n3132), .CLK(n3890), 
        .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n3132), .CLK(n3890), 
        .Q(CRC_OUT_6_3) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n3132), .CLK(n3890), 
        .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n3132), .CLK(n3890), 
        .Q(test_so42) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n3132), .CLK(n3890), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n3131), .CLK(n3891), 
        .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n3131), .CLK(n3891), 
        .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n3131), .CLK(n3891), 
        .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n3131), .CLK(n3891), 
        .Q(CRC_OUT_6_10), .QN(DFF_746_n1) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n3131), .CLK(n3891), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n3131), .CLK(n3891), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n3130), .CLK(n3891), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n3130), .CLK(n3891), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n3130), .CLK(n3891), .Q(CRC_OUT_6_15) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n3130), .CLK(n3891), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n3130), .CLK(n3891), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n3130), .CLK(n3891), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n3129), .CLK(n3892), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n3129), .CLK(n3892), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n3129), .CLK(n3892), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n3129), .CLK(n3892), .Q(test_so43) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n3129), .CLK(n3892), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n3129), .CLK(n3892), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n3128), .CLK(n3892), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n3128), .CLK(n3892), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n3128), .CLK(n3892), .Q(CRC_OUT_6_27) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n3128), .CLK(n3892), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n3128), .CLK(n3892), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n3293), .CLK(n3810), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n3292), .CLK(n3810), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(WX5656), .SI(CRC_OUT_6_31), .SE(n3292), .CLK(n3810), .Q(WX5657) );
  SDFFX1 DFF_769_Q_reg ( .D(WX5658), .SI(WX5657), .SE(n3287), .CLK(n3813), .Q(
        n8528) );
  SDFFX1 DFF_770_Q_reg ( .D(WX5660), .SI(n8528), .SE(n3287), .CLK(n3812), .Q(
        n8527) );
  SDFFX1 DFF_771_Q_reg ( .D(WX5662), .SI(n8527), .SE(n3287), .CLK(n3812), .Q(
        n8526) );
  SDFFX1 DFF_772_Q_reg ( .D(WX5664), .SI(n8526), .SE(n3288), .CLK(n3812), .Q(
        n8525) );
  SDFFX1 DFF_773_Q_reg ( .D(WX5666), .SI(n8525), .SE(n3288), .CLK(n3812), .Q(
        n8524) );
  SDFFX1 DFF_774_Q_reg ( .D(WX5668), .SI(n8524), .SE(n3288), .CLK(n3812), .Q(
        n8523) );
  SDFFX1 DFF_775_Q_reg ( .D(WX5670), .SI(n8523), .SE(n3288), .CLK(n3812), .Q(
        test_so44) );
  SDFFX1 DFF_776_Q_reg ( .D(WX5672), .SI(test_si45), .SE(n3288), .CLK(n3812), 
        .Q(n8520) );
  SDFFX1 DFF_777_Q_reg ( .D(WX5674), .SI(n8520), .SE(n3288), .CLK(n3812), .Q(
        n8519) );
  SDFFX1 DFF_778_Q_reg ( .D(WX5676), .SI(n8519), .SE(n3289), .CLK(n3812), .Q(
        n8518) );
  SDFFX1 DFF_779_Q_reg ( .D(WX5678), .SI(n8518), .SE(n3289), .CLK(n3812), .Q(
        n8517) );
  SDFFX1 DFF_780_Q_reg ( .D(WX5680), .SI(n8517), .SE(n3289), .CLK(n3812), .Q(
        n8516) );
  SDFFX1 DFF_781_Q_reg ( .D(WX5682), .SI(n8516), .SE(n3289), .CLK(n3812), .Q(
        n8515) );
  SDFFX1 DFF_782_Q_reg ( .D(WX5684), .SI(n8515), .SE(n3289), .CLK(n3811), .Q(
        n8514) );
  SDFFX1 DFF_783_Q_reg ( .D(WX5686), .SI(n8514), .SE(n3289), .CLK(n3811), .Q(
        n8513) );
  SDFFX1 DFF_784_Q_reg ( .D(WX5688), .SI(n8513), .SE(n3290), .CLK(n3811), .Q(
        n8512) );
  SDFFX1 DFF_785_Q_reg ( .D(WX5690), .SI(n8512), .SE(n3290), .CLK(n3811), .Q(
        n8511) );
  SDFFX1 DFF_786_Q_reg ( .D(WX5692), .SI(n8511), .SE(n3290), .CLK(n3811), .Q(
        n8510) );
  SDFFX1 DFF_787_Q_reg ( .D(WX5694), .SI(n8510), .SE(n3290), .CLK(n3811), .Q(
        n8509) );
  SDFFX1 DFF_788_Q_reg ( .D(WX5696), .SI(n8509), .SE(n3290), .CLK(n3811), .Q(
        n8508) );
  SDFFX1 DFF_789_Q_reg ( .D(WX5698), .SI(n8508), .SE(n3290), .CLK(n3811), .Q(
        n8507) );
  SDFFX1 DFF_790_Q_reg ( .D(WX5700), .SI(n8507), .SE(n3291), .CLK(n3811), .Q(
        n8506) );
  SDFFX1 DFF_791_Q_reg ( .D(WX5702), .SI(n8506), .SE(n3291), .CLK(n3811), .Q(
        n8505) );
  SDFFX1 DFF_792_Q_reg ( .D(WX5704), .SI(n8505), .SE(n3291), .CLK(n3811), .Q(
        test_so45) );
  SDFFX1 DFF_793_Q_reg ( .D(WX5706), .SI(test_si46), .SE(n3291), .CLK(n3811), 
        .Q(n8502) );
  SDFFX1 DFF_794_Q_reg ( .D(WX5708), .SI(n8502), .SE(n3291), .CLK(n3810), .Q(
        n8501) );
  SDFFX1 DFF_795_Q_reg ( .D(WX5710), .SI(n8501), .SE(n3291), .CLK(n3810), .Q(
        n8500) );
  SDFFX1 DFF_796_Q_reg ( .D(WX5712), .SI(n8500), .SE(n3292), .CLK(n3810), .Q(
        n8499) );
  SDFFX1 DFF_797_Q_reg ( .D(WX5714), .SI(n8499), .SE(n3292), .CLK(n3810), .Q(
        n8498) );
  SDFFX1 DFF_798_Q_reg ( .D(WX5716), .SI(n8498), .SE(n3292), .CLK(n3810), .Q(
        n8497) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n3292), .CLK(n3810), .Q(
        n8496) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n3287), .CLK(n3813), .Q(
        n8495), .QN(n6105) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n3286), .CLK(n3813), .Q(
        n8494), .QN(n6104) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n3286), .CLK(n3813), .Q(
        n8493), .QN(n6103) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n3286), .CLK(n3813), .Q(
        n8492), .QN(n6102) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n3286), .CLK(n3813), .Q(
        n8491), .QN(n6101) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n3285), .CLK(n3814), .Q(
        n8490), .QN(n6100) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n3285), .CLK(n3814), .Q(
        n8489), .QN(n6099) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n3284), .CLK(n3814), .Q(
        n8488), .QN(n6098) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n3284), .CLK(n3814), .Q(
        n8487), .QN(n6097) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n3133), .CLK(n3890), .Q(
        test_so46) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n3284), .CLK(n3814), 
        .Q(n8484), .QN(n6095) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n3283), .CLK(n3814), .Q(
        n8483), .QN(n6094) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n3134), .CLK(n3889), .Q(
        n8482), .QN(n6093) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n3283), .CLK(n3815), .Q(
        n8481), .QN(n6092) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n3282), .CLK(n3815), .Q(
        n8480), .QN(n6091) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n3282), .CLK(n3815), .Q(
        n8479), .QN(n6090) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n3135), .CLK(n3889), .Q(
        WX5849), .QN(n2632) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n3135), .CLK(n3889), .Q(
        WX5851), .QN(n2631) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n3135), .CLK(n3889), .Q(
        WX5853), .QN(n2630) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n3134), .CLK(n3889), .Q(
        WX5855), .QN(n2629) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n3256), .CLK(n3827), .Q(
        WX5857), .QN(n2628) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n3256), .CLK(n3827), .Q(
        WX5859), .QN(n2627) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n3134), .CLK(n3889), .Q(
        WX5861), .QN(n2626) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n3134), .CLK(n3889), .Q(
        WX5863), .QN(n2625) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n3133), .CLK(n3890), .Q(
        WX5865), .QN(n2624) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n3133), .CLK(n3890), .Q(
        WX5867), .QN(n2623) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n3133), .CLK(n3890), .Q(
        test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n3133), .CLK(n3890), 
        .Q(WX5871), .QN(n2622) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n3274), .CLK(n3819), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n3274), .CLK(n3819), .Q(
        WX5875), .QN(n2620) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n3273), .CLK(n3819), .Q(
        WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n3272), .CLK(n3819), .Q(
        WX5879), .QN(n2619) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n3287), .CLK(n3813), .Q(
        WX5881), .QN(n2342) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n3287), .CLK(n3813), .Q(
        WX5883), .QN(n2480) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n3286), .CLK(n3813), .Q(
        WX5885), .QN(n2478) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n3286), .CLK(n3813), .Q(
        WX5887), .QN(n2476) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n3285), .CLK(n3813), .Q(
        WX5889), .QN(n2474) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n3285), .CLK(n3813), .Q(
        WX5891), .QN(n2472) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n3285), .CLK(n3814), .Q(
        WX5893), .QN(n2470) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n3285), .CLK(n3814), .Q(
        WX5895), .QN(n2468) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n3284), .CLK(n3814), .Q(
        WX5897), .QN(n2466) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n3284), .CLK(n3814), .Q(
        WX5899), .QN(n2465) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n3284), .CLK(n3814), .Q(
        WX5901), .QN(n2463) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n3283), .CLK(n3814), .Q(
        test_so48) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n3134), .CLK(n3889), 
        .Q(WX5905), .QN(n2460) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n3282), .CLK(n3815), .Q(
        WX5907), .QN(n2459) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n3282), .CLK(n3815), .Q(
        WX5909), .QN(n2457) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n3282), .CLK(n3815), .Q(
        WX5911), .QN(n2456) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n3281), .CLK(n3815), .Q(
        WX5913) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n3281), .CLK(n3816), .Q(
        WX5915) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n3280), .CLK(n3816), .Q(
        WX5917) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n3280), .CLK(n3816), .Q(
        WX5919) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n3279), .CLK(n3816), .Q(
        WX5921) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n3279), .CLK(n3817), .Q(
        WX5923) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n3277), .CLK(n3817), .Q(
        WX5925) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n3277), .CLK(n3817), .Q(
        WX5927) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n3276), .CLK(n3817), .Q(
        WX5929) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n3276), .CLK(n3818), .Q(
        WX5931) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n3275), .CLK(n3818), .Q(
        WX5933), .QN(n3669) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n3275), .CLK(n3818), .Q(
        WX5935) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n3274), .CLK(n3818), .Q(
        test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n3273), .CLK(n3819), 
        .Q(WX5939) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n3273), .CLK(n3819), .Q(
        WX5941), .QN(n3661) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n3272), .CLK(n3820), .Q(
        WX5943) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n3272), .CLK(n3820), .Q(
        WX5945) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n3271), .CLK(n3820), .Q(
        WX5947) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n3271), .CLK(n3820), .Q(
        WX5949) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n3271), .CLK(n3820), .Q(
        WX5951) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n3270), .CLK(n3820), .Q(
        WX5953) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n3270), .CLK(n3821), .Q(
        WX5955) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n3270), .CLK(n3821), .Q(
        WX5957) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n3269), .CLK(n3821), .Q(
        WX5959) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n3269), .CLK(n3821), .Q(
        WX5961) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n3269), .CLK(n3821), .Q(
        WX5963), .QN(n6096) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n3268), .CLK(n3821), .Q(
        WX5965) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n3283), .CLK(n3815), .Q(
        WX5967), .QN(n2462) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n3283), .CLK(n3815), .Q(
        WX5969) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n3283), .CLK(n3815), .Q(
        test_so50) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n3282), .CLK(n3815), 
        .Q(WX5973) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n3281), .CLK(n3815), .Q(
        WX5975) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n3281), .CLK(n3816), .Q(
        WX5977), .QN(n6089) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n3281), .CLK(n3816), .Q(
        WX5979), .QN(n6088) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n3280), .CLK(n3816), .Q(
        WX5981), .QN(n6087) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n3280), .CLK(n3816), .Q(
        WX5983), .QN(n6086) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n3279), .CLK(n3817), .Q(
        WX5985), .QN(n6085) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n3279), .CLK(n3817), .Q(
        WX5987), .QN(n6084) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n3277), .CLK(n3817), .Q(
        WX5989), .QN(n6083) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n3277), .CLK(n3817), .Q(
        WX5991), .QN(n6082) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n3276), .CLK(n3818), .Q(
        WX5993), .QN(n6081) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n3276), .CLK(n3818), .Q(
        WX5995), .QN(n6080) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n3275), .CLK(n3818), .Q(
        WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n3275), .CLK(n3818), .Q(
        WX5999), .QN(n6079) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n3274), .CLK(n3819), .Q(
        WX6001), .QN(n2621) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n3273), .CLK(n3819), .Q(
        WX6003), .QN(n6078) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n3273), .CLK(n3819), .Q(
        test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n3272), .CLK(n3820), 
        .Q(WX6007), .QN(n6077) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n3271), .CLK(n3820), .Q(
        WX6009), .QN(n2819) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n3271), .CLK(n3820), .Q(
        WX6011), .QN(n2820) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n3271), .CLK(n3820), .Q(
        WX6013), .QN(n2821) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n3270), .CLK(n3820), .Q(
        WX6015), .QN(n2822) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n3270), .CLK(n3821), .Q(
        WX6017), .QN(n2823) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n3270), .CLK(n3821), .Q(
        WX6019), .QN(n2824) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n3269), .CLK(n3821), .Q(
        WX6021), .QN(n2825) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n3269), .CLK(n3821), .Q(
        WX6023), .QN(n2826) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n3269), .CLK(n3821), .Q(
        WX6025), .QN(n2827) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n3268), .CLK(n3821), .Q(
        WX6027), .QN(n2828) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n3268), .CLK(n3822), .Q(
        WX6029), .QN(n2829) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n3268), .CLK(n3822), .Q(
        WX6031), .QN(n2830) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n3268), .CLK(n3822), .Q(
        WX6033), .QN(n2831) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n3268), .CLK(n3822), .Q(
        WX6035), .QN(n2832) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n3267), .CLK(n3822), .Q(
        WX6037), .QN(n2833) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n3267), .CLK(n3822), .Q(
        test_so52) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n3281), .CLK(n3816), 
        .Q(WX6041), .QN(n2834) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n3280), .CLK(n3816), .Q(
        WX6043), .QN(n2835) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n3280), .CLK(n3816), .Q(
        WX6045), .QN(n2836) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n3279), .CLK(n3816), .Q(
        WX6047), .QN(n2837) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n3279), .CLK(n3817), .Q(
        WX6049), .QN(n2696) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n3277), .CLK(n3817), .Q(
        WX6051), .QN(n2838) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n3277), .CLK(n3817), .Q(
        WX6053), .QN(n2839) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n3276), .CLK(n3817), .Q(
        WX6055), .QN(n2840) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n3276), .CLK(n3818), .Q(
        WX6057), .QN(n2841) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n3275), .CLK(n3818), .Q(
        WX6059), .QN(n2842) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n3275), .CLK(n3818), .Q(
        WX6061), .QN(n2843) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n3274), .CLK(n3818), .Q(
        WX6063), .QN(n2697) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n3274), .CLK(n3819), .Q(
        WX6065), .QN(n2844) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n3273), .CLK(n3819), .Q(
        WX6067), .QN(n2845) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n3272), .CLK(n3819), .Q(
        WX6069), .QN(n2846) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n3272), .CLK(n3820), .Q(
        WX6071), .QN(n2710) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n3260), .CLK(n3826), .Q(
        test_so53) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n3260), .CLK(n3826), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n3260), .CLK(n3826), 
        .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n3259), .CLK(n3826), 
        .Q(CRC_OUT_5_3) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n3259), .CLK(n3826), 
        .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n3259), .CLK(n3826), 
        .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n3259), .CLK(n3826), 
        .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n3259), .CLK(n3826), 
        .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n3259), .CLK(n3826), 
        .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n3258), .CLK(n3826), 
        .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n3258), .CLK(n3826), 
        .Q(CRC_OUT_5_10) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n3258), .CLK(n3827), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n3258), .CLK(n3827), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n3258), .CLK(n3827), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n3258), .CLK(n3827), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n3257), .CLK(n3827), .Q(CRC_OUT_5_15), .QN(DFF_943_n1) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n3257), .CLK(n3827), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n3257), .CLK(n3827), .Q(test_so54) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n3257), .CLK(n3827), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n3257), .CLK(n3827), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n3257), .CLK(n3827), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n3267), .CLK(n3822), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n3267), .CLK(n3822), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n3267), .CLK(n3822), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n3267), .CLK(n3822), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n3266), .CLK(n3822), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n3266), .CLK(n3822), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n3266), .CLK(n3823), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n3266), .CLK(n3823), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n3266), .CLK(n3823), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n3266), .CLK(n3823), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n3265), .CLK(n3823), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(WX6949), .SI(CRC_OUT_5_31), .SE(n3265), .CLK(n3823), .Q(WX6950) );
  SDFFX1 DFF_961_Q_reg ( .D(WX6951), .SI(WX6950), .SE(n3260), .CLK(n3826), .Q(
        n8470) );
  SDFFX1 DFF_962_Q_reg ( .D(WX6953), .SI(n8470), .SE(n3260), .CLK(n3825), .Q(
        test_so55) );
  SDFFX1 DFF_963_Q_reg ( .D(WX6955), .SI(test_si56), .SE(n3260), .CLK(n3825), 
        .Q(n8467) );
  SDFFX1 DFF_964_Q_reg ( .D(WX6957), .SI(n8467), .SE(n3261), .CLK(n3825), .Q(
        n8466) );
  SDFFX1 DFF_965_Q_reg ( .D(WX6959), .SI(n8466), .SE(n3261), .CLK(n3825), .Q(
        n8465) );
  SDFFX1 DFF_966_Q_reg ( .D(WX6961), .SI(n8465), .SE(n3261), .CLK(n3825), .Q(
        n8464) );
  SDFFX1 DFF_967_Q_reg ( .D(WX6963), .SI(n8464), .SE(n3261), .CLK(n3825), .Q(
        n8463) );
  SDFFX1 DFF_968_Q_reg ( .D(WX6965), .SI(n8463), .SE(n3261), .CLK(n3825), .Q(
        n8462) );
  SDFFX1 DFF_969_Q_reg ( .D(WX6967), .SI(n8462), .SE(n3261), .CLK(n3825), .Q(
        n8461) );
  SDFFX1 DFF_970_Q_reg ( .D(WX6969), .SI(n8461), .SE(n3262), .CLK(n3825), .Q(
        n8460) );
  SDFFX1 DFF_971_Q_reg ( .D(WX6971), .SI(n8460), .SE(n3262), .CLK(n3825), .Q(
        n8459) );
  SDFFX1 DFF_972_Q_reg ( .D(WX6973), .SI(n8459), .SE(n3262), .CLK(n3825), .Q(
        n8458) );
  SDFFX1 DFF_973_Q_reg ( .D(WX6975), .SI(n8458), .SE(n3262), .CLK(n3825), .Q(
        n8457) );
  SDFFX1 DFF_974_Q_reg ( .D(WX6977), .SI(n8457), .SE(n3262), .CLK(n3824), .Q(
        n8456) );
  SDFFX1 DFF_975_Q_reg ( .D(WX6979), .SI(n8456), .SE(n3262), .CLK(n3824), .Q(
        n8455) );
  SDFFX1 DFF_976_Q_reg ( .D(WX6981), .SI(n8455), .SE(n3263), .CLK(n3824), .Q(
        n8454) );
  SDFFX1 DFF_977_Q_reg ( .D(WX6983), .SI(n8454), .SE(n3263), .CLK(n3824), .Q(
        n8453) );
  SDFFX1 DFF_978_Q_reg ( .D(WX6985), .SI(n8453), .SE(n3263), .CLK(n3824), .Q(
        n8452) );
  SDFFX1 DFF_979_Q_reg ( .D(WX6987), .SI(n8452), .SE(n3263), .CLK(n3824), .Q(
        test_so56) );
  SDFFX1 DFF_980_Q_reg ( .D(WX6989), .SI(test_si57), .SE(n3263), .CLK(n3824), 
        .Q(n8449) );
  SDFFX1 DFF_981_Q_reg ( .D(WX6991), .SI(n8449), .SE(n3263), .CLK(n3824), .Q(
        n8448) );
  SDFFX1 DFF_982_Q_reg ( .D(WX6993), .SI(n8448), .SE(n3264), .CLK(n3824), .Q(
        n8447) );
  SDFFX1 DFF_983_Q_reg ( .D(WX6995), .SI(n8447), .SE(n3264), .CLK(n3824), .Q(
        n8446) );
  SDFFX1 DFF_984_Q_reg ( .D(WX6997), .SI(n8446), .SE(n3264), .CLK(n3824), .Q(
        n8445) );
  SDFFX1 DFF_985_Q_reg ( .D(WX6999), .SI(n8445), .SE(n3264), .CLK(n3824), .Q(
        n8444) );
  SDFFX1 DFF_986_Q_reg ( .D(WX7001), .SI(n8444), .SE(n3264), .CLK(n3823), .Q(
        n8443) );
  SDFFX1 DFF_987_Q_reg ( .D(WX7003), .SI(n8443), .SE(n3264), .CLK(n3823), .Q(
        n8442) );
  SDFFX1 DFF_988_Q_reg ( .D(WX7005), .SI(n8442), .SE(n3265), .CLK(n3823), .Q(
        n8441) );
  SDFFX1 DFF_989_Q_reg ( .D(WX7007), .SI(n8441), .SE(n3265), .CLK(n3823), .Q(
        n8440) );
  SDFFX1 DFF_990_Q_reg ( .D(WX7009), .SI(n8440), .SE(n3265), .CLK(n3823), .Q(
        n8439) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n3265), .CLK(n3823), .Q(
        n8438) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n3250), .CLK(n3831), .Q(
        n8437), .QN(n6076) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n3250), .CLK(n3831), .Q(
        n8436), .QN(n6075) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n3249), .CLK(n3831), .Q(
        n8435), .QN(n6074) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n3248), .CLK(n3831), .Q(
        n8434), .QN(n6073) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n3134), .CLK(n3889), .Q(
        test_so57) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n3247), .CLK(n3832), 
        .Q(n8431), .QN(n6071) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n3247), .CLK(n3832), .Q(
        n8430), .QN(n6070) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n3135), .CLK(n3889), .Q(
        n8429), .QN(n6069) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n3245), .CLK(n3833), .Q(
        n8428), .QN(n6068) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n3244), .CLK(n3833), .Q(
        n8427), .QN(n6067) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n3244), .CLK(n3834), .Q(
        n8426), .QN(n6066) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n3243), .CLK(n3834), .Q(
        n8425), .QN(n6065) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n3243), .CLK(n3834), .Q(
        n8424), .QN(n6064) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n3242), .CLK(n3835), .Q(
        n8423), .QN(n6063) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n3242), .CLK(n3835), .Q(
        n8422), .QN(n6062) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n3240), .CLK(n3835), .Q(
        n8421), .QN(n6061) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n3240), .CLK(n3836), .Q(
        WX7142), .QN(n2618) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n3240), .CLK(n3836), 
        .Q(WX7144), .QN(n2617) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n3239), .CLK(n3836), 
        .Q(WX7146), .QN(n2616) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n3238), .CLK(n3837), 
        .Q(WX7148), .QN(n2615) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n3238), .CLK(n3837), 
        .Q(WX7150), .QN(n2614) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n3256), .CLK(n3828), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n3135), .CLK(n3889), 
        .Q(WX7154), .QN(n2613) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n3255), .CLK(n3828), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n3255), .CLK(n3828), 
        .Q(WX7158), .QN(n2611) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n3254), .CLK(n3828), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n3254), .CLK(n3829), 
        .Q(WX7162), .QN(n2610) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n3254), .CLK(n3829), 
        .Q(WX7164) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n3253), .CLK(n3829), 
        .Q(WX7166), .QN(n2608) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n3252), .CLK(n3829), 
        .Q(WX7168), .QN(n2607) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n3252), .CLK(n3830), 
        .Q(WX7170), .QN(n2606) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n3251), .CLK(n3830), 
        .Q(WX7172), .QN(n2605) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n3250), .CLK(n3830), 
        .Q(WX7174), .QN(n2340) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n3250), .CLK(n3831), 
        .Q(WX7176), .QN(n2454) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n3249), .CLK(n3831), 
        .Q(WX7178), .QN(n2452) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n3248), .CLK(n3832), 
        .Q(WX7180), .QN(n2450) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n3248), .CLK(n3832), 
        .Q(WX7182), .QN(n2449) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n3247), .CLK(n3832), 
        .Q(WX7184), .QN(n2447) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n3246), .CLK(n3832), 
        .Q(test_so59) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n3135), .CLK(n3889), 
        .Q(WX7188), .QN(n2444) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n3245), .CLK(n3833), 
        .Q(WX7190), .QN(n2443) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n3245), .CLK(n3833), 
        .Q(WX7192), .QN(n2441) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n3244), .CLK(n3834), 
        .Q(WX7194), .QN(n2440) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n3244), .CLK(n3834), 
        .Q(WX7196), .QN(n2438) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n3243), .CLK(n3834), 
        .Q(WX7198), .QN(n2436) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n3242), .CLK(n3835), 
        .Q(WX7200), .QN(n2434) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n3241), .CLK(n3835), 
        .Q(WX7202), .QN(n2432) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n3241), .CLK(n3835), 
        .Q(WX7204), .QN(n2430) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n3240), .CLK(n3836), 
        .Q(WX7206) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n3239), .CLK(n3836), 
        .Q(WX7208) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n3239), .CLK(n3836), 
        .Q(WX7210) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n3238), .CLK(n3837), 
        .Q(WX7212) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n3237), .CLK(n3837), 
        .Q(WX7214) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n3255), .CLK(n3828), 
        .Q(WX7216), .QN(n3647) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n3255), .CLK(n3828), 
        .Q(WX7218) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n3255), .CLK(n3828), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n3255), .CLK(n3828), 
        .Q(WX7222) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n3254), .CLK(n3829), 
        .Q(WX7224), .QN(n3639) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n3254), .CLK(n3829), 
        .Q(WX7226) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n3253), .CLK(n3829), 
        .Q(WX7228), .QN(n3635) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n3253), .CLK(n3829), 
        .Q(WX7230) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n3252), .CLK(n3830), 
        .Q(WX7232) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n3252), .CLK(n3830), 
        .Q(WX7234) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n3251), .CLK(n3830), 
        .Q(WX7236) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n3250), .CLK(n3831), 
        .Q(WX7238) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n3249), .CLK(n3831), 
        .Q(WX7240) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n3249), .CLK(n3831), 
        .Q(WX7242) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n3248), .CLK(n3832), 
        .Q(WX7244) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n3248), .CLK(n3832), 
        .Q(WX7246), .QN(n6072) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n3247), .CLK(n3832), 
        .Q(WX7248) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n3246), .CLK(n3833), 
        .Q(WX7250), .QN(n2446) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n3246), .CLK(n3833), 
        .Q(WX7252) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n3246), .CLK(n3833), 
        .Q(test_so61) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n3245), .CLK(n3833), 
        .Q(WX7256) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n3244), .CLK(n3834), 
        .Q(WX7258) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n3243), .CLK(n3834), 
        .Q(WX7260) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n3243), .CLK(n3834), 
        .Q(WX7262) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n3242), .CLK(n3835), 
        .Q(WX7264) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n3241), .CLK(n3835), 
        .Q(WX7266) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n3241), .CLK(n3835), 
        .Q(WX7268) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n3240), .CLK(n3836), 
        .Q(WX7270), .QN(n6060) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n3239), .CLK(n3836), 
        .Q(WX7272), .QN(n6059) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n3239), .CLK(n3836), 
        .Q(WX7274), .QN(n6058) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n3238), .CLK(n3837), 
        .Q(WX7276), .QN(n6057) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n3237), .CLK(n3837), 
        .Q(WX7278), .QN(n6056) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n3237), .CLK(n3837), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n3237), .CLK(n3837), 
        .Q(WX7282), .QN(n6055) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n3236), .CLK(n3838), 
        .Q(WX7284), .QN(n2612) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n3236), .CLK(n3838), 
        .Q(WX7286), .QN(n6054) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n3236), .CLK(n3838), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n3254), .CLK(n3829), 
        .Q(WX7290), .QN(n6053) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n3253), .CLK(n3829), 
        .Q(WX7292), .QN(n2609) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n3253), .CLK(n3829), 
        .Q(WX7294), .QN(n6052) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n3252), .CLK(n3830), 
        .Q(WX7296), .QN(n6051) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n3251), .CLK(n3830), 
        .Q(WX7298), .QN(n6050) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n3251), .CLK(n3830), 
        .Q(WX7300), .QN(n6049) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n3250), .CLK(n3831), 
        .Q(WX7302), .QN(n2792) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n3249), .CLK(n3831), 
        .Q(WX7304), .QN(n2793) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n3249), .CLK(n3831), 
        .Q(WX7306), .QN(n2794) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n3248), .CLK(n3832), 
        .Q(WX7308), .QN(n2795) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n3247), .CLK(n3832), 
        .Q(WX7310), .QN(n2796) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n3247), .CLK(n3832), 
        .Q(WX7312), .QN(n2797) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n3246), .CLK(n3833), 
        .Q(WX7314), .QN(n2798) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n3246), .CLK(n3833), 
        .Q(WX7316), .QN(n2799) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n3245), .CLK(n3833), 
        .Q(WX7318), .QN(n2800) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n3245), .CLK(n3833), 
        .Q(WX7320), .QN(n2801) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n3244), .CLK(n3834), 
        .Q(test_so63) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n3243), .CLK(n3834), 
        .Q(WX7324), .QN(n2802) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n3242), .CLK(n3834), 
        .Q(WX7326), .QN(n2803) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n3242), .CLK(n3835), 
        .Q(WX7328), .QN(n2804) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n3241), .CLK(n3835), 
        .Q(WX7330), .QN(n2805) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n3241), .CLK(n3835), 
        .Q(WX7332), .QN(n2694) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n3240), .CLK(n3836), 
        .Q(WX7334), .QN(n2806) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n3239), .CLK(n3836), 
        .Q(WX7336), .QN(n2807) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n3238), .CLK(n3836), 
        .Q(WX7338), .QN(n2808) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n3238), .CLK(n3837), 
        .Q(WX7340), .QN(n2809) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n3237), .CLK(n3837), 
        .Q(WX7342), .QN(n2695) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n3237), .CLK(n3837), 
        .Q(WX7344), .QN(n2810) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n3236), .CLK(n3837), 
        .Q(WX7346), .QN(n2811) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n3236), .CLK(n3838), 
        .Q(WX7348), .QN(n2812) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n3236), .CLK(n3838), 
        .Q(WX7350), .QN(n2813) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n3235), .CLK(n3838), 
        .Q(WX7352), .QN(n2814) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n3235), .CLK(n3838), 
        .Q(WX7354), .QN(n2815) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n3235), .CLK(n3838), 
        .Q(test_so64) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n3253), .CLK(n3829), 
        .Q(WX7358), .QN(n2816) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n3252), .CLK(n3830), 
        .Q(WX7360), .QN(n2817) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n3251), .CLK(n3830), 
        .Q(WX7362), .QN(n2818) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n3251), .CLK(n3830), 
        .Q(WX7364), .QN(n2709) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n3136), .CLK(n3888), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n3136), .CLK(n3888), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n3136), .CLK(n3888), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n3136), .CLK(n3888), .Q(CRC_OUT_4_3), .QN(DFF_1123_n1) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n3136), .CLK(n3888), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n3136), .CLK(n3888), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n3235), .CLK(n3838), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n3235), .CLK(n3838), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n3235), .CLK(n3838), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n3234), .CLK(n3838), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n3234), .CLK(n3839), .Q(CRC_OUT_4_10) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n3234), .CLK(
        n3839), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n3234), .CLK(
        n3839), .Q(test_so65) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n3234), .CLK(n3839), 
        .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n3234), .CLK(
        n3839), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n3233), .CLK(
        n3839), .Q(CRC_OUT_4_15) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n3233), .CLK(
        n3839), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n3233), .CLK(
        n3839), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n3233), .CLK(
        n3839), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n3233), .CLK(
        n3839), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n3233), .CLK(
        n3839), .Q(CRC_OUT_4_20) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n3232), .CLK(
        n3839), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n3232), .CLK(
        n3840), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n3232), .CLK(
        n3840), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n3232), .CLK(
        n3840), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n3232), .CLK(
        n3840), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n3232), .CLK(
        n3840), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n3231), .CLK(
        n3840), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n3231), .CLK(
        n3840), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n3231), .CLK(
        n3840), .Q(test_so66) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n3231), .CLK(n3840), 
        .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n3231), .CLK(
        n3840), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(WX8242), .SI(CRC_OUT_4_31), .SE(n3231), .CLK(
        n3840), .Q(WX8243) );
  SDFFX1 DFF_1153_Q_reg ( .D(WX8244), .SI(WX8243), .SE(n3225), .CLK(n3843), 
        .Q(n8411) );
  SDFFX1 DFF_1154_Q_reg ( .D(WX8246), .SI(n8411), .SE(n3226), .CLK(n3843), .Q(
        n8410) );
  SDFFX1 DFF_1155_Q_reg ( .D(WX8248), .SI(n8410), .SE(n3226), .CLK(n3843), .Q(
        n8409) );
  SDFFX1 DFF_1156_Q_reg ( .D(WX8250), .SI(n8409), .SE(n3226), .CLK(n3843), .Q(
        n8408) );
  SDFFX1 DFF_1157_Q_reg ( .D(WX8252), .SI(n8408), .SE(n3226), .CLK(n3843), .Q(
        n8407) );
  SDFFX1 DFF_1158_Q_reg ( .D(WX8254), .SI(n8407), .SE(n3226), .CLK(n3843), .Q(
        n8406) );
  SDFFX1 DFF_1159_Q_reg ( .D(WX8256), .SI(n8406), .SE(n3226), .CLK(n3842), .Q(
        n8405) );
  SDFFX1 DFF_1160_Q_reg ( .D(WX8258), .SI(n8405), .SE(n3227), .CLK(n3842), .Q(
        n8404) );
  SDFFX1 DFF_1161_Q_reg ( .D(WX8260), .SI(n8404), .SE(n3227), .CLK(n3842), .Q(
        n8403) );
  SDFFX1 DFF_1162_Q_reg ( .D(WX8262), .SI(n8403), .SE(n3227), .CLK(n3842), .Q(
        n8402) );
  SDFFX1 DFF_1163_Q_reg ( .D(WX8264), .SI(n8402), .SE(n3227), .CLK(n3842), .Q(
        n8401) );
  SDFFX1 DFF_1164_Q_reg ( .D(WX8266), .SI(n8401), .SE(n3227), .CLK(n3842), .Q(
        n8400) );
  SDFFX1 DFF_1165_Q_reg ( .D(WX8268), .SI(n8400), .SE(n3227), .CLK(n3842), .Q(
        n8399) );
  SDFFX1 DFF_1166_Q_reg ( .D(WX8270), .SI(n8399), .SE(n3228), .CLK(n3842), .Q(
        test_so67) );
  SDFFX1 DFF_1167_Q_reg ( .D(WX8272), .SI(test_si68), .SE(n3228), .CLK(n3842), 
        .Q(n8396) );
  SDFFX1 DFF_1168_Q_reg ( .D(WX8274), .SI(n8396), .SE(n3228), .CLK(n3842), .Q(
        n8395) );
  SDFFX1 DFF_1169_Q_reg ( .D(WX8276), .SI(n8395), .SE(n3228), .CLK(n3842), .Q(
        n8394) );
  SDFFX1 DFF_1170_Q_reg ( .D(WX8278), .SI(n8394), .SE(n3228), .CLK(n3842), .Q(
        n8393) );
  SDFFX1 DFF_1171_Q_reg ( .D(WX8280), .SI(n8393), .SE(n3228), .CLK(n3841), .Q(
        n8392) );
  SDFFX1 DFF_1172_Q_reg ( .D(WX8282), .SI(n8392), .SE(n3229), .CLK(n3841), .Q(
        n8391) );
  SDFFX1 DFF_1173_Q_reg ( .D(WX8284), .SI(n8391), .SE(n3229), .CLK(n3841), .Q(
        n8390) );
  SDFFX1 DFF_1174_Q_reg ( .D(WX8286), .SI(n8390), .SE(n3229), .CLK(n3841), .Q(
        n8389) );
  SDFFX1 DFF_1175_Q_reg ( .D(WX8288), .SI(n8389), .SE(n3229), .CLK(n3841), .Q(
        n8388) );
  SDFFX1 DFF_1176_Q_reg ( .D(WX8290), .SI(n8388), .SE(n3229), .CLK(n3841), .Q(
        n8387) );
  SDFFX1 DFF_1177_Q_reg ( .D(WX8292), .SI(n8387), .SE(n3229), .CLK(n3841), .Q(
        n8386) );
  SDFFX1 DFF_1178_Q_reg ( .D(WX8294), .SI(n8386), .SE(n3230), .CLK(n3841), .Q(
        n8385) );
  SDFFX1 DFF_1179_Q_reg ( .D(WX8296), .SI(n8385), .SE(n3230), .CLK(n3841), .Q(
        n8384) );
  SDFFX1 DFF_1180_Q_reg ( .D(WX8298), .SI(n8384), .SE(n3230), .CLK(n3841), .Q(
        n8383) );
  SDFFX1 DFF_1181_Q_reg ( .D(WX8300), .SI(n8383), .SE(n3230), .CLK(n3841), .Q(
        n8382) );
  SDFFX1 DFF_1182_Q_reg ( .D(WX8302), .SI(n8382), .SE(n3230), .CLK(n3841), .Q(
        n8381) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n3230), .CLK(n3840), .Q(
        test_so68) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n3225), .CLK(n3843), 
        .Q(n8378), .QN(n6048) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n3225), .CLK(n3843), .Q(
        n8377), .QN(n6047) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n3225), .CLK(n3843), .Q(
        n8376), .QN(n6046) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n3224), .CLK(n3844), .Q(
        n8375), .QN(n6045) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n3224), .CLK(n3844), .Q(
        n8374), .QN(n6044) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n3223), .CLK(n3844), .Q(
        n8373), .QN(n6043) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n3223), .CLK(n3844), .Q(
        n8372), .QN(n6042) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n3222), .CLK(n3845), .Q(
        n8371), .QN(n6041) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n3222), .CLK(n3845), .Q(
        n8370), .QN(n6040) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n3220), .CLK(n3845), .Q(
        n8369), .QN(n6039) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n3220), .CLK(n3846), .Q(
        n8368), .QN(n6038) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n3219), .CLK(n3846), .Q(
        n8367), .QN(n6037) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n3219), .CLK(n3846), .Q(
        n8366), .QN(n6036) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n3218), .CLK(n3847), .Q(
        n8365), .QN(n6035) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n3218), .CLK(n3847), .Q(
        n8364), .QN(n6034) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n3216), .CLK(n3847), .Q(
        n8363), .QN(n6033) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n3216), .CLK(n3848), .Q(
        test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n3137), .CLK(n3888), 
        .Q(WX8437), .QN(n2604) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n3215), .CLK(n3848), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n3214), .CLK(n3848), 
        .Q(WX8441), .QN(n2602) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n3256), .CLK(n3828), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n3256), .CLK(n3828), 
        .Q(WX8445), .QN(n2601) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n3212), .CLK(n3850), 
        .Q(WX8447) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n3212), .CLK(n3850), 
        .Q(WX8449), .QN(n2599) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n3211), .CLK(n3850), 
        .Q(WX8451), .QN(n2598) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n3211), .CLK(n3850), 
        .Q(WX8453), .QN(n2597) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n3210), .CLK(n3851), 
        .Q(WX8455), .QN(n2596) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n3209), .CLK(n3851), 
        .Q(WX8457), .QN(n2595) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n3209), .CLK(n3851), 
        .Q(WX8459), .QN(n2594) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n3208), .CLK(n3852), 
        .Q(WX8461), .QN(n2593) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n3207), .CLK(n3852), 
        .Q(WX8463), .QN(n2592) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n3207), .CLK(n3852), 
        .Q(WX8465), .QN(n2591) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n3225), .CLK(n3843), 
        .Q(WX8467), .QN(n2338) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n3225), .CLK(n3843), 
        .Q(test_so70) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n3224), .CLK(n3843), 
        .Q(WX8471), .QN(n2427) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n3224), .CLK(n3844), 
        .Q(WX8473), .QN(n2426) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n3224), .CLK(n3844), 
        .Q(WX8475), .QN(n2424) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n3223), .CLK(n3844), 
        .Q(WX8477), .QN(n2423) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n3223), .CLK(n3844), 
        .Q(WX8479), .QN(n2421) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n3222), .CLK(n3845), 
        .Q(WX8481), .QN(n2419) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n3221), .CLK(n3845), 
        .Q(WX8483), .QN(n2417) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n3221), .CLK(n3845), 
        .Q(WX8485), .QN(n2415) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n3220), .CLK(n3846), 
        .Q(WX8487), .QN(n2413) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n3220), .CLK(n3846), 
        .Q(WX8489), .QN(n2411) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n3219), .CLK(n3846), 
        .Q(WX8491), .QN(n2409) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n3218), .CLK(n3847), 
        .Q(WX8493), .QN(n2407) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n3217), .CLK(n3847), 
        .Q(WX8495), .QN(n2405) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n3217), .CLK(n3847), 
        .Q(WX8497), .QN(n2403) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n3216), .CLK(n3848), 
        .Q(WX8499), .QN(n3625) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n3216), .CLK(n3848), 
        .Q(WX8501) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n3215), .CLK(n3848), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n3214), .CLK(n3849), 
        .Q(WX8505) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n3214), .CLK(n3849), 
        .Q(WX8507), .QN(n3617) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n3213), .CLK(n3849), 
        .Q(WX8509) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n3213), .CLK(n3849), 
        .Q(WX8511), .QN(n3613) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n3212), .CLK(n3850), 
        .Q(WX8513) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n3211), .CLK(n3850), 
        .Q(WX8515) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n3211), .CLK(n3850), 
        .Q(WX8517) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n3210), .CLK(n3851), 
        .Q(WX8519) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n3209), .CLK(n3851), 
        .Q(WX8521) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n3209), .CLK(n3851), 
        .Q(WX8523) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n3208), .CLK(n3852), 
        .Q(WX8525) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n3207), .CLK(n3852), 
        .Q(WX8527) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n3207), .CLK(n3852), 
        .Q(WX8529) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n3206), .CLK(n3853), 
        .Q(WX8531) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n3206), .CLK(n3853), 
        .Q(WX8533), .QN(n2429) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n3205), .CLK(n3853), 
        .Q(WX8535) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n3205), .CLK(n3853), 
        .Q(test_so72) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n3224), .CLK(n3844), 
        .Q(WX8539) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n3223), .CLK(n3844), 
        .Q(WX8541) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n3223), .CLK(n3844), 
        .Q(WX8543) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n3222), .CLK(n3845), 
        .Q(WX8545) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n3221), .CLK(n3845), 
        .Q(WX8547) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n3221), .CLK(n3845), 
        .Q(WX8549) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n3220), .CLK(n3846), 
        .Q(WX8551) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n3219), .CLK(n3846), 
        .Q(WX8553) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n3219), .CLK(n3846), 
        .Q(WX8555) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n3218), .CLK(n3847), 
        .Q(WX8557) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n3217), .CLK(n3847), 
        .Q(WX8559) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n3217), .CLK(n3847), 
        .Q(WX8561) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n3216), .CLK(n3848), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n3215), .CLK(n3848), 
        .Q(WX8565), .QN(n6032) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n3215), .CLK(n3848), 
        .Q(WX8567), .QN(n2603) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n3214), .CLK(n3849), 
        .Q(WX8569), .QN(n6031) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n3214), .CLK(n3849), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n3213), .CLK(n3849), 
        .Q(WX8573), .QN(n6030) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n3213), .CLK(n3849), 
        .Q(WX8575), .QN(n2600) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n3212), .CLK(n3850), 
        .Q(WX8577), .QN(n6029) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n3211), .CLK(n3850), 
        .Q(WX8579), .QN(n6028) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n3210), .CLK(n3850), 
        .Q(WX8581), .QN(n6027) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n3210), .CLK(n3851), 
        .Q(WX8583), .QN(n6026) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n3209), .CLK(n3851), 
        .Q(WX8585), .QN(n6025) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n3208), .CLK(n3851), 
        .Q(WX8587), .QN(n6024) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n3208), .CLK(n3852), 
        .Q(WX8589), .QN(n6023) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n3207), .CLK(n3852), 
        .Q(WX8591), .QN(n6022) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n3206), .CLK(n3852), 
        .Q(WX8593), .QN(n6021) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n3206), .CLK(n3853), 
        .Q(WX8595), .QN(n2766) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n3206), .CLK(n3853), 
        .Q(WX8597), .QN(n2767) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n3205), .CLK(n3853), 
        .Q(WX8599), .QN(n2768) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n3205), .CLK(n3853), 
        .Q(WX8601), .QN(n2769) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n3205), .CLK(n3853), 
        .Q(WX8603), .QN(n2770) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n3205), .CLK(n3853), 
        .Q(test_so74) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n3222), .CLK(n3844), 
        .Q(WX8607), .QN(n2771) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n3222), .CLK(n3845), 
        .Q(WX8609), .QN(n2772) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n3221), .CLK(n3845), 
        .Q(WX8611), .QN(n2773) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n3221), .CLK(n3845), 
        .Q(WX8613), .QN(n2774) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n3220), .CLK(n3846), 
        .Q(WX8615), .QN(n2775) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n3219), .CLK(n3846), 
        .Q(WX8617), .QN(n2776) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n3218), .CLK(n3846), 
        .Q(WX8619), .QN(n2777) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n3218), .CLK(n3847), 
        .Q(WX8621), .QN(n2778) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n3217), .CLK(n3847), 
        .Q(WX8623), .QN(n2779) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n3217), .CLK(n3847), 
        .Q(WX8625), .QN(n2691) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n3216), .CLK(n3848), 
        .Q(WX8627), .QN(n2780) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n3215), .CLK(n3848), 
        .Q(WX8629), .QN(n2781) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n3215), .CLK(n3848), 
        .Q(WX8631), .QN(n2782) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n3214), .CLK(n3849), 
        .Q(WX8633), .QN(n2783) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n3213), .CLK(n3849), 
        .Q(WX8635), .QN(n2692) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n3213), .CLK(n3849), 
        .Q(WX8637), .QN(n2784) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n3212), .CLK(n3849), 
        .Q(test_so75) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n3212), .CLK(n3850), 
        .Q(WX8641), .QN(n2785) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n3211), .CLK(n3850), 
        .Q(WX8643), .QN(n2786) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n3210), .CLK(n3851), 
        .Q(WX8645), .QN(n2787) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n3210), .CLK(n3851), 
        .Q(WX8647), .QN(n2788) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n3209), .CLK(n3851), 
        .Q(WX8649), .QN(n2693) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n3208), .CLK(n3852), 
        .Q(WX8651), .QN(n2789) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n3208), .CLK(n3852), 
        .Q(WX8653), .QN(n2790) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n3207), .CLK(n3852), 
        .Q(WX8655), .QN(n2791) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n3206), .CLK(n3853), 
        .Q(WX8657), .QN(n2708) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n3141), .CLK(n3886), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n3141), .CLK(n3886), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n3141), .CLK(n3886), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n3141), .CLK(n3886), .Q(CRC_OUT_3_3) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n3141), .CLK(n3886), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n3140), .CLK(n3886), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n3140), .CLK(n3886), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n3140), .CLK(n3886), .Q(test_so76) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n3140), .CLK(n3886), 
        .Q(CRC_OUT_3_8) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n3140), .CLK(n3886), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n3140), .CLK(n3886), .Q(CRC_OUT_3_10) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n3139), .CLK(
        n3887), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n3139), .CLK(
        n3887), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n3139), .CLK(
        n3887), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n3139), .CLK(
        n3887), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n3139), .CLK(
        n3887), .Q(CRC_OUT_3_15) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n3139), .CLK(
        n3887), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n3138), .CLK(
        n3887), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n3138), .CLK(
        n3887), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n3138), .CLK(
        n3887), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n3138), .CLK(
        n3887), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n3138), .CLK(
        n3887), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n3138), .CLK(
        n3887), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n3137), .CLK(
        n3888), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n3137), .CLK(
        n3888), .Q(test_so77) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n3137), .CLK(n3888), 
        .Q(CRC_OUT_3_25) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n3137), .CLK(
        n3888), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n3137), .CLK(
        n3888), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n3204), .CLK(
        n3853), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n3204), .CLK(
        n3854), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n3204), .CLK(
        n3854), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n3204), .CLK(
        n3854), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(WX9535), .SI(CRC_OUT_3_31), .SE(n3204), .CLK(
        n3854), .Q(WX9536) );
  SDFFX1 DFF_1345_Q_reg ( .D(WX9537), .SI(WX9536), .SE(n3199), .CLK(n3856), 
        .Q(n8353) );
  SDFFX1 DFF_1346_Q_reg ( .D(WX9539), .SI(n8353), .SE(n3199), .CLK(n3856), .Q(
        n8352) );
  SDFFX1 DFF_1347_Q_reg ( .D(WX9541), .SI(n8352), .SE(n3199), .CLK(n3856), .Q(
        n8351) );
  SDFFX1 DFF_1348_Q_reg ( .D(WX9543), .SI(n8351), .SE(n3199), .CLK(n3856), .Q(
        n8350) );
  SDFFX1 DFF_1349_Q_reg ( .D(WX9545), .SI(n8350), .SE(n3199), .CLK(n3856), .Q(
        n8349) );
  SDFFX1 DFF_1350_Q_reg ( .D(WX9547), .SI(n8349), .SE(n3199), .CLK(n3856), .Q(
        n8348) );
  SDFFX1 DFF_1351_Q_reg ( .D(WX9549), .SI(n8348), .SE(n3200), .CLK(n3856), .Q(
        n8347) );
  SDFFX1 DFF_1352_Q_reg ( .D(WX9551), .SI(n8347), .SE(n3200), .CLK(n3856), .Q(
        n8346) );
  SDFFX1 DFF_1353_Q_reg ( .D(WX9553), .SI(n8346), .SE(n3200), .CLK(n3856), .Q(
        test_so78) );
  SDFFX1 DFF_1354_Q_reg ( .D(WX9555), .SI(test_si79), .SE(n3200), .CLK(n3856), 
        .Q(n8343) );
  SDFFX1 DFF_1355_Q_reg ( .D(WX9557), .SI(n8343), .SE(n3200), .CLK(n3856), .Q(
        n8342) );
  SDFFX1 DFF_1356_Q_reg ( .D(WX9559), .SI(n8342), .SE(n3200), .CLK(n3855), .Q(
        n8341) );
  SDFFX1 DFF_1357_Q_reg ( .D(WX9561), .SI(n8341), .SE(n3201), .CLK(n3855), .Q(
        n8340) );
  SDFFX1 DFF_1358_Q_reg ( .D(WX9563), .SI(n8340), .SE(n3201), .CLK(n3855), .Q(
        n8339) );
  SDFFX1 DFF_1359_Q_reg ( .D(WX9565), .SI(n8339), .SE(n3201), .CLK(n3855), .Q(
        n8338) );
  SDFFX1 DFF_1360_Q_reg ( .D(WX9567), .SI(n8338), .SE(n3201), .CLK(n3855), .Q(
        n8337) );
  SDFFX1 DFF_1361_Q_reg ( .D(WX9569), .SI(n8337), .SE(n3201), .CLK(n3855), .Q(
        n8336) );
  SDFFX1 DFF_1362_Q_reg ( .D(WX9571), .SI(n8336), .SE(n3201), .CLK(n3855), .Q(
        n8335) );
  SDFFX1 DFF_1363_Q_reg ( .D(WX9573), .SI(n8335), .SE(n3202), .CLK(n3855), .Q(
        n8334) );
  SDFFX1 DFF_1364_Q_reg ( .D(WX9575), .SI(n8334), .SE(n3202), .CLK(n3855), .Q(
        n8333) );
  SDFFX1 DFF_1365_Q_reg ( .D(WX9577), .SI(n8333), .SE(n3202), .CLK(n3855), .Q(
        n8332) );
  SDFFX1 DFF_1366_Q_reg ( .D(WX9579), .SI(n8332), .SE(n3202), .CLK(n3855), .Q(
        n8331) );
  SDFFX1 DFF_1367_Q_reg ( .D(WX9581), .SI(n8331), .SE(n3202), .CLK(n3855), .Q(
        n8330) );
  SDFFX1 DFF_1368_Q_reg ( .D(WX9583), .SI(n8330), .SE(n3202), .CLK(n3854), .Q(
        n8329) );
  SDFFX1 DFF_1369_Q_reg ( .D(WX9585), .SI(n8329), .SE(n3203), .CLK(n3854), .Q(
        n8328) );
  SDFFX1 DFF_1370_Q_reg ( .D(WX9587), .SI(n8328), .SE(n3203), .CLK(n3854), .Q(
        test_so79) );
  SDFFX1 DFF_1371_Q_reg ( .D(WX9589), .SI(test_si80), .SE(n3203), .CLK(n3854), 
        .Q(n8325) );
  SDFFX1 DFF_1372_Q_reg ( .D(WX9591), .SI(n8325), .SE(n3203), .CLK(n3854), .Q(
        n8324) );
  SDFFX1 DFF_1373_Q_reg ( .D(WX9593), .SI(n8324), .SE(n3203), .CLK(n3854), .Q(
        n8323) );
  SDFFX1 DFF_1374_Q_reg ( .D(WX9595), .SI(n8323), .SE(n3203), .CLK(n3854), .Q(
        n8322) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n3204), .CLK(n3854), .Q(
        n8321) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n3198), .CLK(n3856), .Q(
        n8320), .QN(n6020) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n3198), .CLK(n3857), .Q(
        n8319), .QN(n6019) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n3198), .CLK(n3857), .Q(
        n8318), .QN(n6018) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n3197), .CLK(n3857), .Q(
        n8317), .QN(n6017) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n3197), .CLK(n3857), .Q(
        n8316), .QN(n6016) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n3197), .CLK(n3857), .Q(
        n8315), .QN(n6015) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n3196), .CLK(n3857), .Q(
        n8314), .QN(n6014) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n3196), .CLK(n3858), .Q(
        n8313), .QN(n6013) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n3196), .CLK(n3858), .Q(
        n8312), .QN(n6012) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n3195), .CLK(n3858), .Q(
        n8311), .QN(n6011) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n3195), .CLK(n3858), .Q(
        n8310), .QN(n6010) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n3141), .CLK(n3886), .Q(
        test_so80) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n3194), .CLK(n3858), 
        .Q(n8307), .QN(n6008) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n3194), .CLK(n3859), .Q(
        n8306), .QN(n6007) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n3143), .CLK(n3885), .Q(
        n8305), .QN(n6006) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n3193), .CLK(n3859), .Q(
        n8304), .QN(n6005) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n3143), .CLK(n3885), .Q(
        WX9728), .QN(n2590) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n3192), .CLK(n3859), 
        .Q(WX9730) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n3192), .CLK(n3860), 
        .Q(WX9732), .QN(n2588) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n3192), .CLK(n3860), 
        .Q(WX9734), .QN(n2587) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n3256), .CLK(n3828), 
        .Q(WX9736), .QN(n2586) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n3143), .CLK(n3885), 
        .Q(WX9738), .QN(n2585) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n3143), .CLK(n3885), 
        .Q(WX9740), .QN(n2584) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n3142), .CLK(n3885), 
        .Q(WX9742), .QN(n2583) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n3142), .CLK(n3885), 
        .Q(WX9744), .QN(n2582) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n3142), .CLK(n3885), 
        .Q(WX9746), .QN(n2581) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n3142), .CLK(n3885), 
        .Q(WX9748), .QN(n2580) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n3142), .CLK(n3885), 
        .Q(WX9750), .QN(n2579) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n3142), .CLK(n3885), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n3146), .CLK(n3883), 
        .Q(WX9754), .QN(n2578) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n3185), .CLK(n3863), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n3185), .CLK(n3863), 
        .Q(WX9758), .QN(n2576) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n3198), .CLK(n3857), 
        .Q(WX9760), .QN(n2337) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n3198), .CLK(n3857), 
        .Q(WX9762), .QN(n2401) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n3198), .CLK(n3857), 
        .Q(WX9764), .QN(n2399) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n3197), .CLK(n3857), 
        .Q(WX9766), .QN(n2397) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n3197), .CLK(n3857), 
        .Q(WX9768), .QN(n2395) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n3197), .CLK(n3857), 
        .Q(WX9770), .QN(n2393) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n3196), .CLK(n3858), 
        .Q(WX9772), .QN(n2391) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n3196), .CLK(n3858), 
        .Q(WX9774), .QN(n2389) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n3196), .CLK(n3858), 
        .Q(WX9776), .QN(n2387) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n3195), .CLK(n3858), 
        .Q(WX9778), .QN(n2385) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n3195), .CLK(n3858), 
        .Q(WX9780), .QN(n2383) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n3195), .CLK(n3858), 
        .Q(WX9782), .QN(n2382) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n3195), .CLK(n3858), 
        .Q(WX9784), .QN(n2380) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n3194), .CLK(n3859), 
        .Q(test_so82) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n3143), .CLK(n3885), 
        .Q(WX9788), .QN(n2377) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n3193), .CLK(n3859), 
        .Q(WX9790), .QN(n2376) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n3193), .CLK(n3859), 
        .Q(WX9792) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n3193), .CLK(n3859), 
        .Q(WX9794), .QN(n3591) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n3192), .CLK(n3860), 
        .Q(WX9796) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n3191), .CLK(n3860), 
        .Q(WX9798) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n3191), .CLK(n3860), 
        .Q(WX9800) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n3190), .CLK(n3860), 
        .Q(WX9802) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n3190), .CLK(n3861), 
        .Q(WX9804) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n3189), .CLK(n3861), 
        .Q(WX9806) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n3189), .CLK(n3861), 
        .Q(WX9808) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n3188), .CLK(n3861), 
        .Q(WX9810) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n3188), .CLK(n3862), 
        .Q(WX9812) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n3187), .CLK(n3862), 
        .Q(WX9814) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n3187), .CLK(n3862), 
        .Q(WX9816), .QN(n3569) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n3186), .CLK(n3862), 
        .Q(WX9818) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n3186), .CLK(n3863), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n3185), .CLK(n3863), 
        .Q(WX9822) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n3185), .CLK(n3863), 
        .Q(WX9824) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n3184), .CLK(n3864), 
        .Q(WX9826) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n3184), .CLK(n3864), 
        .Q(WX9828) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n3184), .CLK(n3864), 
        .Q(WX9830) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n3183), .CLK(n3864), 
        .Q(WX9832) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n3183), .CLK(n3864), 
        .Q(WX9834) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n3183), .CLK(n3864), 
        .Q(WX9836) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n3182), .CLK(n3865), 
        .Q(WX9838) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n3182), .CLK(n3865), 
        .Q(WX9840) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n3182), .CLK(n3865), 
        .Q(WX9842) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n3181), .CLK(n3865), 
        .Q(WX9844) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n3181), .CLK(n3865), 
        .Q(WX9846), .QN(n6009) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n3181), .CLK(n3865), 
        .Q(WX9848) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n3194), .CLK(n3859), 
        .Q(WX9850), .QN(n2379) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n3194), .CLK(n3859), 
        .Q(WX9852) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n3194), .CLK(n3859), 
        .Q(test_so84) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n3193), .CLK(n3859), 
        .Q(WX9856), .QN(n6004) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n3193), .CLK(n3859), 
        .Q(WX9858), .QN(n2589) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n3192), .CLK(n3860), 
        .Q(WX9860), .QN(n6003) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n3191), .CLK(n3860), 
        .Q(WX9862), .QN(n6002) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n3191), .CLK(n3860), 
        .Q(WX9864), .QN(n6001) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n3190), .CLK(n3861), 
        .Q(WX9866), .QN(n6000) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n3190), .CLK(n3861), 
        .Q(WX9868), .QN(n5999) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n3189), .CLK(n3861), 
        .Q(WX9870), .QN(n5998) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n3189), .CLK(n3861), 
        .Q(WX9872), .QN(n5997) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n3188), .CLK(n3862), 
        .Q(WX9874), .QN(n5996) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n3188), .CLK(n3862), 
        .Q(WX9876), .QN(n5995) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n3187), .CLK(n3862), 
        .Q(WX9878), .QN(n5994) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n3187), .CLK(n3862), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n3186), .CLK(n3863), 
        .Q(WX9882), .QN(n5993) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n3186), .CLK(n3863), 
        .Q(WX9884), .QN(n2577) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n3185), .CLK(n3863), 
        .Q(WX9886), .QN(n5992) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n3184), .CLK(n3863), 
        .Q(test_so85) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n3184), .CLK(n3864), 
        .Q(WX9890), .QN(n2740) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n3184), .CLK(n3864), 
        .Q(WX9892), .QN(n2741) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n3183), .CLK(n3864), 
        .Q(WX9894), .QN(n2742) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n3183), .CLK(n3864), 
        .Q(WX9896), .QN(n2743) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n3183), .CLK(n3864), 
        .Q(WX9898), .QN(n2744) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n3182), .CLK(n3864), 
        .Q(WX9900), .QN(n2745) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n3182), .CLK(n3865), 
        .Q(WX9902), .QN(n2746) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n3182), .CLK(n3865), 
        .Q(WX9904), .QN(n2747) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n3181), .CLK(n3865), 
        .Q(WX9906), .QN(n2748) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n3181), .CLK(n3865), 
        .Q(WX9908), .QN(n2749) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n3181), .CLK(n3865), 
        .Q(WX9910), .QN(n2750) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n3180), .CLK(n3865), 
        .Q(WX9912), .QN(n2751) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n3180), .CLK(n3866), 
        .Q(WX9914), .QN(n2752) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n3180), .CLK(n3866), 
        .Q(WX9916), .QN(n2753) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n3180), .CLK(n3866), 
        .Q(WX9918), .QN(n2688) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n3180), .CLK(n3866), 
        .Q(WX9920), .QN(n2754) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n3180), .CLK(n3866), 
        .Q(test_so86) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n3192), .CLK(n3860), 
        .Q(WX9924), .QN(n2755) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n3191), .CLK(n3860), 
        .Q(WX9926), .QN(n2756) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n3191), .CLK(n3860), 
        .Q(WX9928), .QN(n2689) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n3190), .CLK(n3861), 
        .Q(WX9930), .QN(n2757) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n3190), .CLK(n3861), 
        .Q(WX9932), .QN(n2758) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n3189), .CLK(n3861), 
        .Q(WX9934), .QN(n2759) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n3189), .CLK(n3861), 
        .Q(WX9936), .QN(n2760) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n3188), .CLK(n3862), 
        .Q(WX9938), .QN(n2761) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n3188), .CLK(n3862), 
        .Q(WX9940), .QN(n2762) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n3187), .CLK(n3862), 
        .Q(WX9942), .QN(n2690) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n3187), .CLK(n3862), 
        .Q(WX9944), .QN(n2763) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n3186), .CLK(n3863), 
        .Q(WX9946), .QN(n2764) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n3186), .CLK(n3863), 
        .Q(WX9948), .QN(n2765) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n3185), .CLK(n3863), 
        .Q(WX9950), .QN(n2707) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n3147), .CLK(n3883), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n3146), .CLK(
        n3883), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n3146), .CLK(
        n3883), .Q(test_so87) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n3146), .CLK(n3883), 
        .Q(CRC_OUT_2_3) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n3146), .CLK(
        n3883), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n3146), .CLK(
        n3883), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n3145), .CLK(
        n3884), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n3145), .CLK(
        n3884), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n3145), .CLK(
        n3884), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n3145), .CLK(
        n3884), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n3145), .CLK(
        n3884), .Q(CRC_OUT_2_10) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n3145), .CLK(
        n3884), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n3144), .CLK(
        n3884), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n3144), .CLK(
        n3884), .Q(CRC_OUT_2_13) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n3144), .CLK(
        n3884), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n3144), .CLK(
        n3884), .Q(CRC_OUT_2_15) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n3144), .CLK(
        n3884), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n3144), .CLK(
        n3884), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n3143), .CLK(
        n3885), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n3179), .CLK(
        n3866), .Q(test_so88) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n3179), .CLK(n3866), 
        .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n3179), .CLK(
        n3866), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n3179), .CLK(
        n3866), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n3179), .CLK(
        n3866), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n3179), .CLK(
        n3866), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n3178), .CLK(
        n3866), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n3178), .CLK(
        n3867), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n3178), .CLK(
        n3867), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n3178), .CLK(
        n3867), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n3178), .CLK(
        n3867), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n3178), .CLK(
        n3867), .Q(CRC_OUT_2_30) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n3177), .CLK(
        n3867), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(WX10828), .SI(CRC_OUT_2_31), .SE(n3177), .CLK(
        n3867), .Q(WX10829) );
  SDFFX1 DFF_1537_Q_reg ( .D(WX10830), .SI(WX10829), .SE(n3172), .CLK(n3870), 
        .Q(n8295) );
  SDFFX1 DFF_1538_Q_reg ( .D(WX10832), .SI(n8295), .SE(n3172), .CLK(n3870), 
        .Q(n8294) );
  SDFFX1 DFF_1539_Q_reg ( .D(WX10834), .SI(n8294), .SE(n3172), .CLK(n3869), 
        .Q(n8293) );
  SDFFX1 DFF_1540_Q_reg ( .D(WX10836), .SI(n8293), .SE(n3173), .CLK(n3869), 
        .Q(test_so89) );
  SDFFX1 DFF_1541_Q_reg ( .D(WX10838), .SI(test_si90), .SE(n3173), .CLK(n3869), 
        .Q(n8290) );
  SDFFX1 DFF_1542_Q_reg ( .D(WX10840), .SI(n8290), .SE(n3173), .CLK(n3869), 
        .Q(n8289) );
  SDFFX1 DFF_1543_Q_reg ( .D(WX10842), .SI(n8289), .SE(n3173), .CLK(n3869), 
        .Q(n8288) );
  SDFFX1 DFF_1544_Q_reg ( .D(WX10844), .SI(n8288), .SE(n3173), .CLK(n3869), 
        .Q(n8287) );
  SDFFX1 DFF_1545_Q_reg ( .D(WX10846), .SI(n8287), .SE(n3173), .CLK(n3869), 
        .Q(n8286) );
  SDFFX1 DFF_1546_Q_reg ( .D(WX10848), .SI(n8286), .SE(n3174), .CLK(n3869), 
        .Q(n8285) );
  SDFFX1 DFF_1547_Q_reg ( .D(WX10850), .SI(n8285), .SE(n3174), .CLK(n3869), 
        .Q(n8284) );
  SDFFX1 DFF_1548_Q_reg ( .D(WX10852), .SI(n8284), .SE(n3174), .CLK(n3869), 
        .Q(n8283) );
  SDFFX1 DFF_1549_Q_reg ( .D(WX10854), .SI(n8283), .SE(n3174), .CLK(n3869), 
        .Q(n8282) );
  SDFFX1 DFF_1550_Q_reg ( .D(WX10856), .SI(n8282), .SE(n3174), .CLK(n3869), 
        .Q(n8281) );
  SDFFX1 DFF_1551_Q_reg ( .D(WX10858), .SI(n8281), .SE(n3174), .CLK(n3868), 
        .Q(n8280) );
  SDFFX1 DFF_1552_Q_reg ( .D(WX10860), .SI(n8280), .SE(n3175), .CLK(n3868), 
        .Q(n8279) );
  SDFFX1 DFF_1553_Q_reg ( .D(WX10862), .SI(n8279), .SE(n3175), .CLK(n3868), 
        .Q(n8278) );
  SDFFX1 DFF_1554_Q_reg ( .D(WX10864), .SI(n8278), .SE(n3175), .CLK(n3868), 
        .Q(n8277) );
  SDFFX1 DFF_1555_Q_reg ( .D(WX10866), .SI(n8277), .SE(n3175), .CLK(n3868), 
        .Q(n8276) );
  SDFFX1 DFF_1556_Q_reg ( .D(WX10868), .SI(n8276), .SE(n3175), .CLK(n3868), 
        .Q(n8275) );
  SDFFX1 DFF_1557_Q_reg ( .D(WX10870), .SI(n8275), .SE(n3175), .CLK(n3868), 
        .Q(test_so90) );
  SDFFX1 DFF_1558_Q_reg ( .D(WX10872), .SI(test_si91), .SE(n3176), .CLK(n3868), 
        .Q(n8272) );
  SDFFX1 DFF_1559_Q_reg ( .D(WX10874), .SI(n8272), .SE(n3176), .CLK(n3868), 
        .Q(n8271) );
  SDFFX1 DFF_1560_Q_reg ( .D(WX10876), .SI(n8271), .SE(n3176), .CLK(n3868), 
        .Q(n8270) );
  SDFFX1 DFF_1561_Q_reg ( .D(WX10878), .SI(n8270), .SE(n3176), .CLK(n3868), 
        .Q(n8269) );
  SDFFX1 DFF_1562_Q_reg ( .D(WX10880), .SI(n8269), .SE(n3176), .CLK(n3868), 
        .Q(n8268) );
  SDFFX1 DFF_1563_Q_reg ( .D(WX10882), .SI(n8268), .SE(n3176), .CLK(n3867), 
        .Q(n8267) );
  SDFFX1 DFF_1564_Q_reg ( .D(WX10884), .SI(n8267), .SE(n3177), .CLK(n3867), 
        .Q(n8266) );
  SDFFX1 DFF_1565_Q_reg ( .D(WX10886), .SI(n8266), .SE(n3177), .CLK(n3867), 
        .Q(n8265) );
  SDFFX1 DFF_1566_Q_reg ( .D(WX10888), .SI(n8265), .SE(n3177), .CLK(n3867), 
        .Q(n8264) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n3177), .CLK(n3867), 
        .Q(n8263) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n3172), .CLK(n3870), 
        .Q(n8262), .QN(n6218) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n3171), .CLK(n3870), 
        .Q(n8261), .QN(n6217) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n3171), .CLK(n3870), 
        .Q(n8260), .QN(n6216) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n3171), .CLK(n3870), 
        .Q(n8259), .QN(n6215) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n3171), .CLK(n3870), 
        .Q(n8258), .QN(n6214) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n3170), .CLK(n3871), 
        .Q(n8257), .QN(n6213) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n3170), .CLK(n3871), 
        .Q(test_so91) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n3169), .CLK(n3871), 
        .Q(n8254), .QN(n6211) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n3169), .CLK(n3871), 
        .Q(n8253), .QN(n6210) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n3147), .CLK(n3883), 
        .Q(n8252), .QN(n6209) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n3168), .CLK(n3871), 
        .Q(n8251), .QN(n6208) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n3168), .CLK(n3872), 
        .Q(n8250), .QN(n6207) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n3168), .CLK(n3872), 
        .Q(n8249), .QN(n6206) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n3167), .CLK(n3872), 
        .Q(n8248), .QN(n6205) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n3166), .CLK(n3872), 
        .Q(n8247), .QN(n6204) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n3165), .CLK(n3873), 
        .Q(n8246), .QN(n6203) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n3165), .CLK(n3873), 
        .Q(WX11021), .QN(n2575) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n3164), .CLK(n3873), 
        .Q(WX11023), .QN(n2574) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n3164), .CLK(n3874), 
        .Q(WX11025), .QN(n2573) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n3163), .CLK(n3874), 
        .Q(WX11027), .QN(n2572) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n3162), .CLK(n3875), 
        .Q(WX11029), .QN(n2571) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n3162), .CLK(n3875), 
        .Q(WX11031), .QN(n2570) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n3161), .CLK(n3875), 
        .Q(WX11033), .QN(n2569) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n3161), .CLK(n3875), 
        .Q(test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n3147), .CLK(n3883), 
        .Q(WX11037), .QN(n2568) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n3160), .CLK(n3876), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n3160), .CLK(n3876), 
        .Q(WX11041), .QN(n2566) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n3159), .CLK(n3877), 
        .Q(WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n3159), .CLK(n3877), 
        .Q(WX11045), .QN(n2565) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n3158), .CLK(n3877), 
        .Q(WX11047) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n3157), .CLK(n3878), 
        .Q(WX11049), .QN(n2563) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n3157), .CLK(n3878), 
        .Q(WX11051), .QN(n2562) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n3172), .CLK(n3870), 
        .Q(WX11053), .QN(n2335) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n3172), .CLK(n3870), 
        .Q(WX11055), .QN(n2374) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n3171), .CLK(n3870), 
        .Q(WX11057), .QN(n2372) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n3171), .CLK(n3870), 
        .Q(WX11059), .QN(n2370) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n3170), .CLK(n3870), 
        .Q(WX11061), .QN(n2368) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n3170), .CLK(n3871), 
        .Q(WX11063), .QN(n2366) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n3170), .CLK(n3871), 
        .Q(WX11065), .QN(n2365) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n3170), .CLK(n3871), 
        .Q(WX11067), .QN(n2363) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n3169), .CLK(n3871), 
        .Q(test_so93) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n3147), .CLK(n3883), 
        .Q(WX11071), .QN(n2360) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n3168), .CLK(n3872), 
        .Q(WX11073), .QN(n2359) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n3168), .CLK(n3872), 
        .Q(WX11075), .QN(n2357) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n3167), .CLK(n3872), 
        .Q(WX11077), .QN(n2356) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n3167), .CLK(n3872), 
        .Q(WX11079), .QN(n2354) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n3166), .CLK(n3873), 
        .Q(WX11081), .QN(n2352) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n3166), .CLK(n3873), 
        .Q(WX11083), .QN(n2350) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n3165), .CLK(n3873), 
        .Q(WX11085) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n3164), .CLK(n3874), 
        .Q(WX11087) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n3164), .CLK(n3874), 
        .Q(WX11089) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n3163), .CLK(n3874), 
        .Q(WX11091) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n3162), .CLK(n3875), 
        .Q(WX11093) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n3162), .CLK(n3875), 
        .Q(WX11095) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n3161), .CLK(n3875), 
        .Q(WX11097) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n3161), .CLK(n3875), 
        .Q(WX11099), .QN(n3547) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n3160), .CLK(n3876), 
        .Q(WX11101) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n3160), .CLK(n3876), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n3159), .CLK(n3876), 
        .Q(WX11105) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n3159), .CLK(n3877), 
        .Q(WX11107), .QN(n3539) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n3158), .CLK(n3877), 
        .Q(WX11109) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n3158), .CLK(n3877), 
        .Q(WX11111), .QN(n3535) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n3157), .CLK(n3878), 
        .Q(WX11113) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n3156), .CLK(n3878), 
        .Q(WX11115) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n3156), .CLK(n3878), 
        .Q(WX11117) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n3156), .CLK(n3878), 
        .Q(WX11119) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n3155), .CLK(n3879), 
        .Q(WX11121) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n3155), .CLK(n3879), 
        .Q(WX11123) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n3155), .CLK(n3879), 
        .Q(WX11125) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n3154), .CLK(n3879), 
        .Q(WX11127) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n3154), .CLK(n3879), 
        .Q(WX11129), .QN(n6212) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n3154), .CLK(n3879), 
        .Q(WX11131) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n3169), .CLK(n3871), 
        .Q(WX11133), .QN(n2362) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n3169), .CLK(n3871), 
        .Q(WX11135) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n3169), .CLK(n3871), 
        .Q(test_so95) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n3168), .CLK(n3872), 
        .Q(WX11139) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n3167), .CLK(n3872), 
        .Q(WX11141) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n3167), .CLK(n3872), 
        .Q(WX11143) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n3166), .CLK(n3873), 
        .Q(WX11145) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n3166), .CLK(n3873), 
        .Q(WX11147) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n3165), .CLK(n3873), 
        .Q(WX11149), .QN(n6202) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n3164), .CLK(n3874), 
        .Q(WX11151), .QN(n6201) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n3163), .CLK(n3874), 
        .Q(WX11153), .QN(n6200) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n3163), .CLK(n3874), 
        .Q(WX11155), .QN(n6199) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155_Tj_Payload), .SE(
        test_se_Trojan), .CLK(n3828), .Q(WX11157), .QN(n6198) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(test_se_Trojan), 
        .CLK(n3875), .Q(WX11159), .QN(n6197) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(test_se_Trojan), 
        .CLK(n3875), .Q(WX11161), .QN(n6196) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(test_se_Trojan), 
        .CLK(n3876), .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(test_se_Trojan), 
        .CLK(n3876), .Q(WX11165), .QN(n6195) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(test_se_Trojan), 
        .CLK(n3876), .Q(WX11167), .QN(n2567) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(test_se_Trojan), 
        .CLK(n3876), .Q(WX11169), .QN(n6194) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(test_se_Trojan), 
        .CLK(n3877), .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n3158), .CLK(n3877), 
        .Q(WX11173), .QN(n6193) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n3158), .CLK(n3877), 
        .Q(WX11175), .QN(n2564) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n3157), .CLK(n3878), 
        .Q(WX11177), .QN(n6192) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n3156), .CLK(n3878), 
        .Q(WX11179), .QN(n6191) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n3156), .CLK(n3878), 
        .Q(WX11181), .QN(n2714) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n3155), .CLK(n3879), 
        .Q(WX11183), .QN(n2715) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n3155), .CLK(n3879), 
        .Q(WX11185), .QN(n2716) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n3155), .CLK(n3879), 
        .Q(WX11187), .QN(n2717) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n3154), .CLK(n3879), 
        .Q(WX11189), .QN(n2718) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n3154), .CLK(n3879), 
        .Q(WX11191), .QN(n2719) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n3154), .CLK(n3879), 
        .Q(WX11193), .QN(n2720) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n3153), .CLK(n3880), 
        .Q(WX11195), .QN(n2721) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n3153), .CLK(n3880), 
        .Q(WX11197), .QN(n2722) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n3153), .CLK(n3880), 
        .Q(WX11199), .QN(n2723) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n3153), .CLK(n3880), 
        .Q(WX11201), .QN(n2724) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n3153), .CLK(n3880), 
        .Q(WX11203), .QN(n2725) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n3153), .CLK(n3880), 
        .Q(test_so97) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n3167), .CLK(n3872), 
        .Q(WX11207), .QN(n2726) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n3166), .CLK(n3873), 
        .Q(WX11209), .QN(n2727) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n3165), .CLK(n3873), 
        .Q(WX11211), .QN(n2685) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n3165), .CLK(n3873), 
        .Q(WX11213), .QN(n2728) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n3164), .CLK(n3874), 
        .Q(WX11215), .QN(n2729) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n3163), .CLK(n3874), 
        .Q(WX11217), .QN(n2730) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n3163), .CLK(n3874), 
        .Q(WX11219), .QN(n2731) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n3162), .CLK(n3874), 
        .Q(WX11221), .QN(n2686) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n3162), .CLK(n3875), 
        .Q(WX11223), .QN(n2732) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n3161), .CLK(n3875), 
        .Q(WX11225), .QN(n2733) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n3161), .CLK(n3876), 
        .Q(WX11227), .QN(n2734) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n3160), .CLK(n3876), 
        .Q(WX11229), .QN(n2735) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n3160), .CLK(n3876), 
        .Q(WX11231), .QN(n2736) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n3159), .CLK(n3877), 
        .Q(WX11233), .QN(n2737) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n3159), .CLK(n3877), 
        .Q(WX11235), .QN(n2687) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n3158), .CLK(n3877), 
        .Q(WX11237), .QN(n2738) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n3157), .CLK(n3878), 
        .Q(test_so98) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n3157), .CLK(n3878), 
        .Q(WX11241), .QN(n2739) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n3156), .CLK(n3878), 
        .Q(WX11243), .QN(n2706) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n3151), .CLK(n3881), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n3151), .CLK(
        n3881), .Q(CRC_OUT_1_1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n3151), .CLK(
        n3881), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n3151), .CLK(
        n3881), .Q(CRC_OUT_1_3), .QN(DFF_1699_n1) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n3150), .CLK(
        n3881), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n3150), .CLK(
        n3881), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n3150), .CLK(
        n3881), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n3150), .CLK(
        n3881), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n3150), .CLK(
        n3881), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n3150), .CLK(
        n3881), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n3149), .CLK(
        n3882), .Q(CRC_OUT_1_10), .QN(DFF_1706_n1) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n3149), .CLK(
        n3882), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n3149), .CLK(
        n3882), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n3149), .CLK(
        n3882), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n3149), .CLK(
        n3882), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n3149), .CLK(n3882), .Q(CRC_OUT_1_15), .QN(DFF_1711_n1) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n3148), .CLK(
        n3882), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n3148), .CLK(
        n3882), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n3148), .CLK(
        n3882), .Q(CRC_OUT_1_18) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n3148), .CLK(
        n3882), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n3148), .CLK(
        n3882), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n3148), .CLK(
        n3882), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n3147), .CLK(
        n3883), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n3147), .CLK(
        n3883), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n3152), .CLK(
        n3880), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n3152), .CLK(
        n3880), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n3152), .CLK(
        n3880), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n3152), .CLK(
        n3880), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n3152), .CLK(
        n3880), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n3152), .CLK(
        n3880), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n3151), .CLK(
        n3881), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n3151), .CLK(
        n3881), .Q(test_so100) );
  AND2X1 Trojan1 ( .IN1(WX742), .IN2(WX7249), .Q(Tj_OUT1) );
  AND2X1 Trojan2 ( .IN1(WX5922), .IN2(WX5960), .Q(Tj_OUT2) );
  AND2X1 Trojan3 ( .IN1(WX4697), .IN2(WX9032), .Q(Tj_OUT3) );
  AND2X1 Trojan4 ( .IN1(WX8298), .IN2(WX10846), .Q(Tj_OUT4) );
  NOR4X0 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .QN(Tj_OUT1234) );
  AND2X1 Trojan5 ( .IN1(WX3340), .IN2(WX6476), .Q(Tj_OUT5) );
  AND2X1 Trojan6 ( .IN1(WX9819), .IN2(WX1813), .Q(Tj_OUT6) );
  AND2X1 Trojan7 ( .IN1(WX5710), .IN2(WX3458), .Q(Tj_OUT7) );
  AND2X1 Trojan8 ( .IN1(WX9060), .IN2(WX7749), .Q(Tj_OUT8) );
  NOR4X0 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .QN(Tj_OUT5678) );
  INVX0 TrojanINV_test_se ( .INP(n3393), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  DFFX2 TrojanScanEnable ( .D(1'b1), .CLK(Tj_Trigger), .Q(Trojan_SE) );
  MUX21X1 Trojan_Payload1 ( .IN1(n3393), .IN2(1'b1), .S(Trojan_SE), .Q(
        test_se_Trojan) );
  MUX21X1 Trojan_Payload2 ( .IN1(WX11155), .IN2(WX3442), .S(Trojan_SE), .Q(
        WX11155_Tj_Payload) );
  NBUFFX2 U3327 ( .INP(n3071), .Z(n3069) );
  NBUFFX2 U3328 ( .INP(n3075), .Z(n3047) );
  NBUFFX2 U3329 ( .INP(n3075), .Z(n3048) );
  NBUFFX2 U3330 ( .INP(n3075), .Z(n3049) );
  NBUFFX2 U3331 ( .INP(n3075), .Z(n3050) );
  NBUFFX2 U3332 ( .INP(n3073), .Z(n3057) );
  NBUFFX2 U3333 ( .INP(n3073), .Z(n3059) );
  NBUFFX2 U3334 ( .INP(n3073), .Z(n3060) );
  NBUFFX2 U3335 ( .INP(n3072), .Z(n3061) );
  NBUFFX2 U3336 ( .INP(n3072), .Z(n3062) );
  NBUFFX2 U3337 ( .INP(n3072), .Z(n3063) );
  NBUFFX2 U3338 ( .INP(n3074), .Z(n3051) );
  NBUFFX2 U3339 ( .INP(n3074), .Z(n3052) );
  NBUFFX2 U3340 ( .INP(n3073), .Z(n3058) );
  NBUFFX2 U3341 ( .INP(n3074), .Z(n3053) );
  NBUFFX2 U3342 ( .INP(n3074), .Z(n3054) );
  NBUFFX2 U3343 ( .INP(n3074), .Z(n3055) );
  NBUFFX2 U3344 ( .INP(n3073), .Z(n3056) );
  NBUFFX2 U3345 ( .INP(n3072), .Z(n3065) );
  NBUFFX2 U3346 ( .INP(n3072), .Z(n3064) );
  NBUFFX2 U3347 ( .INP(n3071), .Z(n3066) );
  NBUFFX2 U3348 ( .INP(n3071), .Z(n3067) );
  NBUFFX2 U3349 ( .INP(n3071), .Z(n3068) );
  NBUFFX2 U3350 ( .INP(n3071), .Z(n3070) );
  NBUFFX2 U3351 ( .INP(n3932), .Z(n3760) );
  NBUFFX2 U3352 ( .INP(n3932), .Z(n3758) );
  NBUFFX2 U3353 ( .INP(n3932), .Z(n3759) );
  NBUFFX2 U3354 ( .INP(n3932), .Z(n3757) );
  NBUFFX2 U3355 ( .INP(n3908), .Z(n3882) );
  NBUFFX2 U3356 ( .INP(n3908), .Z(n3881) );
  NBUFFX2 U3357 ( .INP(n3908), .Z(n3880) );
  NBUFFX2 U3358 ( .INP(n3908), .Z(n3879) );
  NBUFFX2 U3359 ( .INP(n3909), .Z(n3878) );
  NBUFFX2 U3360 ( .INP(n3909), .Z(n3877) );
  NBUFFX2 U3361 ( .INP(n3909), .Z(n3876) );
  NBUFFX2 U3362 ( .INP(n3909), .Z(n3875) );
  NBUFFX2 U3363 ( .INP(n3909), .Z(n3874) );
  NBUFFX2 U3364 ( .INP(n3910), .Z(n3873) );
  NBUFFX2 U3365 ( .INP(n3910), .Z(n3872) );
  NBUFFX2 U3366 ( .INP(n3910), .Z(n3871) );
  NBUFFX2 U3367 ( .INP(n3911), .Z(n3868) );
  NBUFFX2 U3368 ( .INP(n3910), .Z(n3869) );
  NBUFFX2 U3369 ( .INP(n3910), .Z(n3870) );
  NBUFFX2 U3370 ( .INP(n3911), .Z(n3867) );
  NBUFFX2 U3371 ( .INP(n3907), .Z(n3884) );
  NBUFFX2 U3372 ( .INP(n3911), .Z(n3866) );
  NBUFFX2 U3373 ( .INP(n3911), .Z(n3865) );
  NBUFFX2 U3374 ( .INP(n3911), .Z(n3864) );
  NBUFFX2 U3375 ( .INP(n3912), .Z(n3862) );
  NBUFFX2 U3376 ( .INP(n3912), .Z(n3861) );
  NBUFFX2 U3377 ( .INP(n3912), .Z(n3863) );
  NBUFFX2 U3378 ( .INP(n3908), .Z(n3883) );
  NBUFFX2 U3379 ( .INP(n3912), .Z(n3860) );
  NBUFFX2 U3380 ( .INP(n3907), .Z(n3885) );
  NBUFFX2 U3381 ( .INP(n3912), .Z(n3859) );
  NBUFFX2 U3382 ( .INP(n3913), .Z(n3858) );
  NBUFFX2 U3383 ( .INP(n3913), .Z(n3857) );
  NBUFFX2 U3384 ( .INP(n3913), .Z(n3855) );
  NBUFFX2 U3385 ( .INP(n3913), .Z(n3856) );
  NBUFFX2 U3386 ( .INP(n3913), .Z(n3854) );
  NBUFFX2 U3387 ( .INP(n3907), .Z(n3887) );
  NBUFFX2 U3388 ( .INP(n3907), .Z(n3886) );
  NBUFFX2 U3389 ( .INP(n3914), .Z(n3853) );
  NBUFFX2 U3390 ( .INP(n3914), .Z(n3849) );
  NBUFFX2 U3391 ( .INP(n3914), .Z(n3852) );
  NBUFFX2 U3392 ( .INP(n3914), .Z(n3851) );
  NBUFFX2 U3393 ( .INP(n3914), .Z(n3850) );
  NBUFFX2 U3394 ( .INP(n3915), .Z(n3848) );
  NBUFFX2 U3395 ( .INP(n3915), .Z(n3847) );
  NBUFFX2 U3396 ( .INP(n3915), .Z(n3846) );
  NBUFFX2 U3397 ( .INP(n3915), .Z(n3845) );
  NBUFFX2 U3398 ( .INP(n3915), .Z(n3844) );
  NBUFFX2 U3399 ( .INP(n3916), .Z(n3841) );
  NBUFFX2 U3400 ( .INP(n3916), .Z(n3842) );
  NBUFFX2 U3401 ( .INP(n3916), .Z(n3843) );
  NBUFFX2 U3402 ( .INP(n3916), .Z(n3840) );
  NBUFFX2 U3403 ( .INP(n3916), .Z(n3839) );
  NBUFFX2 U3404 ( .INP(n3907), .Z(n3888) );
  NBUFFX2 U3405 ( .INP(n3917), .Z(n3838) );
  NBUFFX2 U3406 ( .INP(n3918), .Z(n3830) );
  NBUFFX2 U3407 ( .INP(n3918), .Z(n3829) );
  NBUFFX2 U3408 ( .INP(n3919), .Z(n3828) );
  NBUFFX2 U3409 ( .INP(n3917), .Z(n3837) );
  NBUFFX2 U3410 ( .INP(n3917), .Z(n3836) );
  NBUFFX2 U3411 ( .INP(n3917), .Z(n3835) );
  NBUFFX2 U3412 ( .INP(n3917), .Z(n3834) );
  NBUFFX2 U3413 ( .INP(n3918), .Z(n3833) );
  NBUFFX2 U3414 ( .INP(n3918), .Z(n3832) );
  NBUFFX2 U3415 ( .INP(n3918), .Z(n3831) );
  NBUFFX2 U3416 ( .INP(n3919), .Z(n3824) );
  NBUFFX2 U3417 ( .INP(n3919), .Z(n3825) );
  NBUFFX2 U3418 ( .INP(n3920), .Z(n3823) );
  NBUFFX2 U3419 ( .INP(n3919), .Z(n3826) );
  NBUFFX2 U3420 ( .INP(n3920), .Z(n3822) );
  NBUFFX2 U3421 ( .INP(n3920), .Z(n3821) );
  NBUFFX2 U3422 ( .INP(n3920), .Z(n3820) );
  NBUFFX2 U3423 ( .INP(n3921), .Z(n3818) );
  NBUFFX2 U3424 ( .INP(n3921), .Z(n3817) );
  NBUFFX2 U3425 ( .INP(n3921), .Z(n3816) );
  NBUFFX2 U3426 ( .INP(n3920), .Z(n3819) );
  NBUFFX2 U3427 ( .INP(n3919), .Z(n3827) );
  NBUFFX2 U3428 ( .INP(n3921), .Z(n3815) );
  NBUFFX2 U3429 ( .INP(n3906), .Z(n3889) );
  NBUFFX2 U3430 ( .INP(n3921), .Z(n3814) );
  NBUFFX2 U3431 ( .INP(n3922), .Z(n3811) );
  NBUFFX2 U3432 ( .INP(n3922), .Z(n3812) );
  NBUFFX2 U3433 ( .INP(n3922), .Z(n3813) );
  NBUFFX2 U3434 ( .INP(n3906), .Z(n3891) );
  NBUFFX2 U3435 ( .INP(n3906), .Z(n3890) );
  NBUFFX2 U3436 ( .INP(n3922), .Z(n3810) );
  NBUFFX2 U3437 ( .INP(n3922), .Z(n3809) );
  NBUFFX2 U3438 ( .INP(n3923), .Z(n3808) );
  NBUFFX2 U3439 ( .INP(n3923), .Z(n3807) );
  NBUFFX2 U3440 ( .INP(n3923), .Z(n3806) );
  NBUFFX2 U3441 ( .INP(n3923), .Z(n3805) );
  NBUFFX2 U3442 ( .INP(n3923), .Z(n3804) );
  NBUFFX2 U3443 ( .INP(n3924), .Z(n3803) );
  NBUFFX2 U3444 ( .INP(n3924), .Z(n3802) );
  NBUFFX2 U3445 ( .INP(n3924), .Z(n3801) );
  NBUFFX2 U3446 ( .INP(n3924), .Z(n3800) );
  NBUFFX2 U3447 ( .INP(n3925), .Z(n3797) );
  NBUFFX2 U3448 ( .INP(n3925), .Z(n3798) );
  NBUFFX2 U3449 ( .INP(n3924), .Z(n3799) );
  NBUFFX2 U3450 ( .INP(n3906), .Z(n3893) );
  NBUFFX2 U3451 ( .INP(n3906), .Z(n3892) );
  NBUFFX2 U3452 ( .INP(n3925), .Z(n3796) );
  NBUFFX2 U3453 ( .INP(n3925), .Z(n3795) );
  NBUFFX2 U3454 ( .INP(n3926), .Z(n3790) );
  NBUFFX2 U3455 ( .INP(n3925), .Z(n3794) );
  NBUFFX2 U3456 ( .INP(n3926), .Z(n3793) );
  NBUFFX2 U3457 ( .INP(n3926), .Z(n3792) );
  NBUFFX2 U3458 ( .INP(n3926), .Z(n3791) );
  NBUFFX2 U3459 ( .INP(n3905), .Z(n3894) );
  NBUFFX2 U3460 ( .INP(n3926), .Z(n3789) );
  NBUFFX2 U3461 ( .INP(n3927), .Z(n3788) );
  NBUFFX2 U3462 ( .INP(n3927), .Z(n3787) );
  NBUFFX2 U3463 ( .INP(n3927), .Z(n3784) );
  NBUFFX2 U3464 ( .INP(n3927), .Z(n3785) );
  NBUFFX2 U3465 ( .INP(n3927), .Z(n3786) );
  NBUFFX2 U3466 ( .INP(n3905), .Z(n3897) );
  NBUFFX2 U3467 ( .INP(n3905), .Z(n3896) );
  NBUFFX2 U3468 ( .INP(n3905), .Z(n3895) );
  NBUFFX2 U3469 ( .INP(n3928), .Z(n3782) );
  NBUFFX2 U3470 ( .INP(n3904), .Z(n3900) );
  NBUFFX2 U3471 ( .INP(n3904), .Z(n3899) );
  NBUFFX2 U3472 ( .INP(n3904), .Z(n3901) );
  NBUFFX2 U3473 ( .INP(n3928), .Z(n3781) );
  NBUFFX2 U3474 ( .INP(n3928), .Z(n3780) );
  NBUFFX2 U3475 ( .INP(n3905), .Z(n3898) );
  NBUFFX2 U3476 ( .INP(n3928), .Z(n3779) );
  NBUFFX2 U3477 ( .INP(n3928), .Z(n3778) );
  NBUFFX2 U3478 ( .INP(n3929), .Z(n3777) );
  NBUFFX2 U3479 ( .INP(n3929), .Z(n3776) );
  NBUFFX2 U3480 ( .INP(n3929), .Z(n3773) );
  NBUFFX2 U3481 ( .INP(n3929), .Z(n3774) );
  NBUFFX2 U3482 ( .INP(n3929), .Z(n3772) );
  NBUFFX2 U3483 ( .INP(n3904), .Z(n3902) );
  NBUFFX2 U3484 ( .INP(n3930), .Z(n3771) );
  NBUFFX2 U3485 ( .INP(n3930), .Z(n3770) );
  NBUFFX2 U3486 ( .INP(n3930), .Z(n3769) );
  NBUFFX2 U3487 ( .INP(n3930), .Z(n3768) );
  NBUFFX2 U3488 ( .INP(n3930), .Z(n3767) );
  NBUFFX2 U3489 ( .INP(n3931), .Z(n3766) );
  NBUFFX2 U3490 ( .INP(n3931), .Z(n3765) );
  NBUFFX2 U3491 ( .INP(n3931), .Z(n3764) );
  NBUFFX2 U3492 ( .INP(n3931), .Z(n3762) );
  NBUFFX2 U3493 ( .INP(n3931), .Z(n3761) );
  NBUFFX2 U3494 ( .INP(n3904), .Z(n3903) );
  NBUFFX2 U3495 ( .INP(n2997), .Z(n3019) );
  NBUFFX2 U3496 ( .INP(n2997), .Z(n3020) );
  NBUFFX2 U3497 ( .INP(n2997), .Z(n3018) );
  NBUFFX2 U3498 ( .INP(n3102), .Z(n3095) );
  NBUFFX2 U3499 ( .INP(n3101), .Z(n3099) );
  NBUFFX2 U3500 ( .INP(n3101), .Z(n3098) );
  NBUFFX2 U3501 ( .INP(n3101), .Z(n3096) );
  NBUFFX2 U3502 ( .INP(n3101), .Z(n3097) );
  NBUFFX2 U3503 ( .INP(n2996), .Z(n3017) );
  NBUFFX2 U3504 ( .INP(n2996), .Z(n3016) );
  NBUFFX2 U3505 ( .INP(n3102), .Z(n3094) );
  NBUFFX2 U3506 ( .INP(n3101), .Z(n3100) );
  NBUFFX2 U3507 ( .INP(n3105), .Z(n3080) );
  NBUFFX2 U3508 ( .INP(n3105), .Z(n3078) );
  NBUFFX2 U3509 ( .INP(n3105), .Z(n3079) );
  NBUFFX2 U3510 ( .INP(n3103), .Z(n3088) );
  NBUFFX2 U3511 ( .INP(n3103), .Z(n3089) );
  NBUFFX2 U3512 ( .INP(n3103), .Z(n3090) );
  NBUFFX2 U3513 ( .INP(n3102), .Z(n3091) );
  NBUFFX2 U3514 ( .INP(n3104), .Z(n3081) );
  NBUFFX2 U3515 ( .INP(n3104), .Z(n3083) );
  NBUFFX2 U3516 ( .INP(n3104), .Z(n3084) );
  NBUFFX2 U3517 ( .INP(n3104), .Z(n3085) );
  NBUFFX2 U3518 ( .INP(n3103), .Z(n3086) );
  NBUFFX2 U3519 ( .INP(n3103), .Z(n3087) );
  NBUFFX2 U3520 ( .INP(n3102), .Z(n3093) );
  NBUFFX2 U3521 ( .INP(n3102), .Z(n3092) );
  NBUFFX2 U3522 ( .INP(n3104), .Z(n3082) );
  NBUFFX2 U3523 ( .INP(n2995), .Z(n3009) );
  NBUFFX2 U3524 ( .INP(n2994), .Z(n3007) );
  NBUFFX2 U3525 ( .INP(n2994), .Z(n3006) );
  NBUFFX2 U3526 ( .INP(n2995), .Z(n3008) );
  NBUFFX2 U3527 ( .INP(n2994), .Z(n3005) );
  NBUFFX2 U3528 ( .INP(n2994), .Z(n3004) );
  NBUFFX2 U3529 ( .INP(n2993), .Z(n2999) );
  NBUFFX2 U3530 ( .INP(n2993), .Z(n2998) );
  NBUFFX2 U3531 ( .INP(n2994), .Z(n3003) );
  NBUFFX2 U3532 ( .INP(n2996), .Z(n3014) );
  NBUFFX2 U3533 ( .INP(n2996), .Z(n3015) );
  NBUFFX2 U3534 ( .INP(n2996), .Z(n3013) );
  NBUFFX2 U3535 ( .INP(n2995), .Z(n3012) );
  NBUFFX2 U3536 ( .INP(n2995), .Z(n3011) );
  NBUFFX2 U3537 ( .INP(n2995), .Z(n3010) );
  NBUFFX2 U3538 ( .INP(n2993), .Z(n3002) );
  NBUFFX2 U3539 ( .INP(n2993), .Z(n3001) );
  NBUFFX2 U3540 ( .INP(n2993), .Z(n3000) );
  NBUFFX2 U3541 ( .INP(n2997), .Z(n3021) );
  NBUFFX2 U3542 ( .INP(n3022), .Z(n3028) );
  NBUFFX2 U3543 ( .INP(n3027), .Z(n3043) );
  NBUFFX2 U3544 ( .INP(n3022), .Z(n3029) );
  NBUFFX2 U3545 ( .INP(n3022), .Z(n3030) );
  NBUFFX2 U3546 ( .INP(n3023), .Z(n3031) );
  NBUFFX2 U3547 ( .INP(n3023), .Z(n3032) );
  NBUFFX2 U3548 ( .INP(n3024), .Z(n3036) );
  NBUFFX2 U3549 ( .INP(n3025), .Z(n3037) );
  NBUFFX2 U3550 ( .INP(n3025), .Z(n3038) );
  NBUFFX2 U3551 ( .INP(n3025), .Z(n3039) );
  NBUFFX2 U3552 ( .INP(n3026), .Z(n3040) );
  NBUFFX2 U3553 ( .INP(n3026), .Z(n3041) );
  NBUFFX2 U3554 ( .INP(n3026), .Z(n3042) );
  NBUFFX2 U3555 ( .INP(n3023), .Z(n3033) );
  NBUFFX2 U3556 ( .INP(n3024), .Z(n3034) );
  NBUFFX2 U3557 ( .INP(n3024), .Z(n3035) );
  NBUFFX2 U3559 ( .INP(n3027), .Z(n3044) );
  NBUFFX2 U3560 ( .INP(n3580), .Z(n3577) );
  NBUFFX2 U3561 ( .INP(n3580), .Z(n3578) );
  NBUFFX2 U3562 ( .INP(n3583), .Z(n3567) );
  NBUFFX2 U3563 ( .INP(n3583), .Z(n3568) );
  NBUFFX2 U3564 ( .INP(n3583), .Z(n3570) );
  NBUFFX2 U3565 ( .INP(n3582), .Z(n3571) );
  NBUFFX2 U3566 ( .INP(n3582), .Z(n3572) );
  NBUFFX2 U3567 ( .INP(n3582), .Z(n3573) );
  NBUFFX2 U3568 ( .INP(n3581), .Z(n3574) );
  NBUFFX2 U3569 ( .INP(n3581), .Z(n3575) );
  NBUFFX2 U3570 ( .INP(n3581), .Z(n3576) );
  NBUFFX2 U3571 ( .INP(n3580), .Z(n3579) );
  NBUFFX2 U3572 ( .INP(n2148), .Z(n3022) );
  NBUFFX2 U3573 ( .INP(n2148), .Z(n3025) );
  NBUFFX2 U3574 ( .INP(n2148), .Z(n3026) );
  NBUFFX2 U3575 ( .INP(n2148), .Z(n3023) );
  NBUFFX2 U3576 ( .INP(n2148), .Z(n3024) );
  NBUFFX2 U3577 ( .INP(n2148), .Z(n3027) );
  NBUFFX2 U3578 ( .INP(TM1), .Z(n3583) );
  NBUFFX2 U3579 ( .INP(TM1), .Z(n3582) );
  NBUFFX2 U3580 ( .INP(TM1), .Z(n3580) );
  NBUFFX2 U3581 ( .INP(TM1), .Z(n3581) );
  NBUFFX2 U3582 ( .INP(n3947), .Z(n2993) );
  NBUFFX2 U3583 ( .INP(n3947), .Z(n2994) );
  NBUFFX2 U3584 ( .INP(n3947), .Z(n2995) );
  NBUFFX2 U3585 ( .INP(n3947), .Z(n2996) );
  NBUFFX2 U3586 ( .INP(n3947), .Z(n2997) );
  NBUFFX2 U3587 ( .INP(n2152), .Z(n3045) );
  NBUFFX2 U3588 ( .INP(n2152), .Z(n3046) );
  NBUFFX2 U3589 ( .INP(n3045), .Z(n3071) );
  NBUFFX2 U3590 ( .INP(n3045), .Z(n3072) );
  NBUFFX2 U3591 ( .INP(n3045), .Z(n3073) );
  NBUFFX2 U3592 ( .INP(n3046), .Z(n3074) );
  NBUFFX2 U3593 ( .INP(n3046), .Z(n3075) );
  NBUFFX2 U3594 ( .INP(n2153), .Z(n3076) );
  NBUFFX2 U3595 ( .INP(n2153), .Z(n3077) );
  NBUFFX2 U3596 ( .INP(n3076), .Z(n3101) );
  NBUFFX2 U3597 ( .INP(n3076), .Z(n3102) );
  NBUFFX2 U3598 ( .INP(n3076), .Z(n3103) );
  NBUFFX2 U3599 ( .INP(n3077), .Z(n3104) );
  NBUFFX2 U3600 ( .INP(n3077), .Z(n3105) );
  NBUFFX2 U3601 ( .INP(n3507), .Z(n3106) );
  NBUFFX2 U3602 ( .INP(n3507), .Z(n3107) );
  NBUFFX2 U3603 ( .INP(n3506), .Z(n3108) );
  NBUFFX2 U3604 ( .INP(n3506), .Z(n3109) );
  NBUFFX2 U3605 ( .INP(n3506), .Z(n3110) );
  NBUFFX2 U3606 ( .INP(n3504), .Z(n3111) );
  NBUFFX2 U3607 ( .INP(n3504), .Z(n3112) );
  NBUFFX2 U3608 ( .INP(n3504), .Z(n3113) );
  NBUFFX2 U3609 ( .INP(n3502), .Z(n3114) );
  NBUFFX2 U3610 ( .INP(n3502), .Z(n3115) );
  NBUFFX2 U3611 ( .INP(n3502), .Z(n3116) );
  NBUFFX2 U3612 ( .INP(n3500), .Z(n3117) );
  NBUFFX2 U3613 ( .INP(n3500), .Z(n3118) );
  NBUFFX2 U3614 ( .INP(n3500), .Z(n3119) );
  NBUFFX2 U3615 ( .INP(n3499), .Z(n3120) );
  NBUFFX2 U3616 ( .INP(n3499), .Z(n3121) );
  NBUFFX2 U3617 ( .INP(n3499), .Z(n3122) );
  NBUFFX2 U3618 ( .INP(n3498), .Z(n3123) );
  NBUFFX2 U3619 ( .INP(n3498), .Z(n3124) );
  NBUFFX2 U3620 ( .INP(n3498), .Z(n3125) );
  NBUFFX2 U3621 ( .INP(n3496), .Z(n3126) );
  NBUFFX2 U3622 ( .INP(n3496), .Z(n3127) );
  NBUFFX2 U3623 ( .INP(n3496), .Z(n3128) );
  NBUFFX2 U3624 ( .INP(n3494), .Z(n3129) );
  NBUFFX2 U3625 ( .INP(n3494), .Z(n3130) );
  NBUFFX2 U3626 ( .INP(n3494), .Z(n3131) );
  NBUFFX2 U3627 ( .INP(n3492), .Z(n3132) );
  NBUFFX2 U3628 ( .INP(n3492), .Z(n3133) );
  NBUFFX2 U3629 ( .INP(n3492), .Z(n3134) );
  NBUFFX2 U3630 ( .INP(n3490), .Z(n3135) );
  NBUFFX2 U3631 ( .INP(n3490), .Z(n3136) );
  NBUFFX2 U3632 ( .INP(n3490), .Z(n3137) );
  NBUFFX2 U3633 ( .INP(n3488), .Z(n3138) );
  NBUFFX2 U3634 ( .INP(n3488), .Z(n3139) );
  NBUFFX2 U3635 ( .INP(n3488), .Z(n3140) );
  NBUFFX2 U3636 ( .INP(n3487), .Z(n3141) );
  NBUFFX2 U3637 ( .INP(n3487), .Z(n3142) );
  NBUFFX2 U3638 ( .INP(n3487), .Z(n3143) );
  NBUFFX2 U3639 ( .INP(n3486), .Z(n3144) );
  NBUFFX2 U3640 ( .INP(n3486), .Z(n3145) );
  NBUFFX2 U3641 ( .INP(n3486), .Z(n3146) );
  NBUFFX2 U3642 ( .INP(n3484), .Z(n3147) );
  NBUFFX2 U3643 ( .INP(n3484), .Z(n3148) );
  NBUFFX2 U3644 ( .INP(n3484), .Z(n3149) );
  NBUFFX2 U3645 ( .INP(n3482), .Z(n3150) );
  NBUFFX2 U3646 ( .INP(n3482), .Z(n3151) );
  NBUFFX2 U3647 ( .INP(n3482), .Z(n3152) );
  NBUFFX2 U3648 ( .INP(n3480), .Z(n3153) );
  NBUFFX2 U3649 ( .INP(n3480), .Z(n3154) );
  NBUFFX2 U3650 ( .INP(n3480), .Z(n3155) );
  NBUFFX2 U3651 ( .INP(n3478), .Z(n3156) );
  NBUFFX2 U3652 ( .INP(n3478), .Z(n3157) );
  NBUFFX2 U3653 ( .INP(n3478), .Z(n3158) );
  NBUFFX2 U3654 ( .INP(n3476), .Z(n3159) );
  NBUFFX2 U3655 ( .INP(n3476), .Z(n3160) );
  NBUFFX2 U3656 ( .INP(n3476), .Z(n3161) );
  NBUFFX2 U3657 ( .INP(n3474), .Z(n3162) );
  NBUFFX2 U3658 ( .INP(n3474), .Z(n3163) );
  NBUFFX2 U3659 ( .INP(n3474), .Z(n3164) );
  NBUFFX2 U3660 ( .INP(n3472), .Z(n3165) );
  NBUFFX2 U3661 ( .INP(n3472), .Z(n3166) );
  NBUFFX2 U3662 ( .INP(n3472), .Z(n3167) );
  NBUFFX2 U3663 ( .INP(n3470), .Z(n3168) );
  NBUFFX2 U3664 ( .INP(n3470), .Z(n3169) );
  NBUFFX2 U3665 ( .INP(n3470), .Z(n3170) );
  NBUFFX2 U3666 ( .INP(n3468), .Z(n3171) );
  NBUFFX2 U3667 ( .INP(n3468), .Z(n3172) );
  NBUFFX2 U3668 ( .INP(n3468), .Z(n3173) );
  NBUFFX2 U3669 ( .INP(n3466), .Z(n3174) );
  NBUFFX2 U3670 ( .INP(n3466), .Z(n3175) );
  NBUFFX2 U3671 ( .INP(n3466), .Z(n3176) );
  NBUFFX2 U3672 ( .INP(n3465), .Z(n3177) );
  NBUFFX2 U3673 ( .INP(n3465), .Z(n3178) );
  NBUFFX2 U3674 ( .INP(n3465), .Z(n3179) );
  NBUFFX2 U3675 ( .INP(n3464), .Z(n3180) );
  NBUFFX2 U3676 ( .INP(n3464), .Z(n3181) );
  NBUFFX2 U3677 ( .INP(n3464), .Z(n3182) );
  NBUFFX2 U3678 ( .INP(n3463), .Z(n3183) );
  NBUFFX2 U3679 ( .INP(n3463), .Z(n3184) );
  NBUFFX2 U3680 ( .INP(n3463), .Z(n3185) );
  NBUFFX2 U3681 ( .INP(n3462), .Z(n3186) );
  NBUFFX2 U3682 ( .INP(n3462), .Z(n3187) );
  NBUFFX2 U3683 ( .INP(n3462), .Z(n3188) );
  NBUFFX2 U3684 ( .INP(n3461), .Z(n3189) );
  NBUFFX2 U3685 ( .INP(n3461), .Z(n3190) );
  NBUFFX2 U3686 ( .INP(n3461), .Z(n3191) );
  NBUFFX2 U3687 ( .INP(n3460), .Z(n3192) );
  NBUFFX2 U3688 ( .INP(n3460), .Z(n3193) );
  NBUFFX2 U3689 ( .INP(n3460), .Z(n3194) );
  NBUFFX2 U3690 ( .INP(n3459), .Z(n3195) );
  NBUFFX2 U3691 ( .INP(n3459), .Z(n3196) );
  NBUFFX2 U3692 ( .INP(n3459), .Z(n3197) );
  NBUFFX2 U3693 ( .INP(n3458), .Z(n3198) );
  NBUFFX2 U3694 ( .INP(n3458), .Z(n3199) );
  NBUFFX2 U3695 ( .INP(n3458), .Z(n3200) );
  NBUFFX2 U3696 ( .INP(n3457), .Z(n3201) );
  NBUFFX2 U3697 ( .INP(n3457), .Z(n3202) );
  NBUFFX2 U3698 ( .INP(n3457), .Z(n3203) );
  NBUFFX2 U3699 ( .INP(n3456), .Z(n3204) );
  NBUFFX2 U3700 ( .INP(n3456), .Z(n3205) );
  NBUFFX2 U3701 ( .INP(n3456), .Z(n3206) );
  NBUFFX2 U3702 ( .INP(n3455), .Z(n3207) );
  NBUFFX2 U3703 ( .INP(n3455), .Z(n3208) );
  NBUFFX2 U3704 ( .INP(n3455), .Z(n3209) );
  NBUFFX2 U3705 ( .INP(n3454), .Z(n3210) );
  NBUFFX2 U3706 ( .INP(n3454), .Z(n3211) );
  NBUFFX2 U3707 ( .INP(n3454), .Z(n3212) );
  NBUFFX2 U3708 ( .INP(n3453), .Z(n3213) );
  NBUFFX2 U3709 ( .INP(n3453), .Z(n3214) );
  NBUFFX2 U3710 ( .INP(n3453), .Z(n3215) );
  NBUFFX2 U3711 ( .INP(n3452), .Z(n3216) );
  NBUFFX2 U3712 ( .INP(n3452), .Z(n3217) );
  NBUFFX2 U3713 ( .INP(n3452), .Z(n3218) );
  NBUFFX2 U3714 ( .INP(n3451), .Z(n3219) );
  NBUFFX2 U3715 ( .INP(n3451), .Z(n3220) );
  NBUFFX2 U3716 ( .INP(n3451), .Z(n3221) );
  NBUFFX2 U3717 ( .INP(n3450), .Z(n3222) );
  NBUFFX2 U3718 ( .INP(n3450), .Z(n3223) );
  NBUFFX2 U3719 ( .INP(n3450), .Z(n3224) );
  NBUFFX2 U3720 ( .INP(n3449), .Z(n3225) );
  NBUFFX2 U3721 ( .INP(n3449), .Z(n3226) );
  NBUFFX2 U3722 ( .INP(n3449), .Z(n3227) );
  NBUFFX2 U3723 ( .INP(n3448), .Z(n3228) );
  NBUFFX2 U3724 ( .INP(n3448), .Z(n3229) );
  NBUFFX2 U3725 ( .INP(n3448), .Z(n3230) );
  NBUFFX2 U3726 ( .INP(n3447), .Z(n3231) );
  NBUFFX2 U3727 ( .INP(n3447), .Z(n3232) );
  NBUFFX2 U3728 ( .INP(n3447), .Z(n3233) );
  NBUFFX2 U3729 ( .INP(n3446), .Z(n3234) );
  NBUFFX2 U3730 ( .INP(n3446), .Z(n3235) );
  NBUFFX2 U3731 ( .INP(n3446), .Z(n3236) );
  NBUFFX2 U3732 ( .INP(n3445), .Z(n3237) );
  NBUFFX2 U3733 ( .INP(n3445), .Z(n3238) );
  NBUFFX2 U3734 ( .INP(n3445), .Z(n3239) );
  NBUFFX2 U3735 ( .INP(n3444), .Z(n3240) );
  NBUFFX2 U3736 ( .INP(n3444), .Z(n3241) );
  NBUFFX2 U3737 ( .INP(n3444), .Z(n3242) );
  NBUFFX2 U3738 ( .INP(n3443), .Z(n3243) );
  NBUFFX2 U3739 ( .INP(n3443), .Z(n3244) );
  NBUFFX2 U3740 ( .INP(n3443), .Z(n3245) );
  NBUFFX2 U3741 ( .INP(n3442), .Z(n3246) );
  NBUFFX2 U3742 ( .INP(n3442), .Z(n3247) );
  NBUFFX2 U3743 ( .INP(n3442), .Z(n3248) );
  NBUFFX2 U3744 ( .INP(n3441), .Z(n3249) );
  NBUFFX2 U3745 ( .INP(n3441), .Z(n3250) );
  NBUFFX2 U3746 ( .INP(n3441), .Z(n3251) );
  NBUFFX2 U3747 ( .INP(n3440), .Z(n3252) );
  NBUFFX2 U3748 ( .INP(n3440), .Z(n3253) );
  NBUFFX2 U3749 ( .INP(n3440), .Z(n3254) );
  NBUFFX2 U3750 ( .INP(n3439), .Z(n3255) );
  NBUFFX2 U3751 ( .INP(n3439), .Z(n3256) );
  NBUFFX2 U3752 ( .INP(n3439), .Z(n3257) );
  NBUFFX2 U3753 ( .INP(n3438), .Z(n3258) );
  NBUFFX2 U3754 ( .INP(n3438), .Z(n3259) );
  NBUFFX2 U3755 ( .INP(n3438), .Z(n3260) );
  NBUFFX2 U3756 ( .INP(n3437), .Z(n3261) );
  NBUFFX2 U3757 ( .INP(n3437), .Z(n3262) );
  NBUFFX2 U3758 ( .INP(n3437), .Z(n3263) );
  NBUFFX2 U3759 ( .INP(n3436), .Z(n3264) );
  NBUFFX2 U3760 ( .INP(n3436), .Z(n3265) );
  NBUFFX2 U3761 ( .INP(n3436), .Z(n3266) );
  NBUFFX2 U3762 ( .INP(n3435), .Z(n3267) );
  NBUFFX2 U3763 ( .INP(n3435), .Z(n3268) );
  NBUFFX2 U3764 ( .INP(n3435), .Z(n3269) );
  NBUFFX2 U3765 ( .INP(n3434), .Z(n3270) );
  NBUFFX2 U3766 ( .INP(n3434), .Z(n3271) );
  NBUFFX2 U3767 ( .INP(n3434), .Z(n3272) );
  NBUFFX2 U3768 ( .INP(n3433), .Z(n3273) );
  NBUFFX2 U3769 ( .INP(n3433), .Z(n3274) );
  NBUFFX2 U3770 ( .INP(n3433), .Z(n3275) );
  NBUFFX2 U3771 ( .INP(n3432), .Z(n3276) );
  NBUFFX2 U3772 ( .INP(n3432), .Z(n3277) );
  NBUFFX2 U3773 ( .INP(n3432), .Z(n3279) );
  NBUFFX2 U3774 ( .INP(n3431), .Z(n3280) );
  NBUFFX2 U3775 ( .INP(n3431), .Z(n3281) );
  NBUFFX2 U3776 ( .INP(n3431), .Z(n3282) );
  NBUFFX2 U3777 ( .INP(n3430), .Z(n3283) );
  NBUFFX2 U3778 ( .INP(n3430), .Z(n3284) );
  NBUFFX2 U3779 ( .INP(n3430), .Z(n3285) );
  NBUFFX2 U3780 ( .INP(n3429), .Z(n3286) );
  NBUFFX2 U3781 ( .INP(n3429), .Z(n3287) );
  NBUFFX2 U3782 ( .INP(n3429), .Z(n3288) );
  NBUFFX2 U3783 ( .INP(n3428), .Z(n3289) );
  NBUFFX2 U3784 ( .INP(n3428), .Z(n3290) );
  NBUFFX2 U3785 ( .INP(n3428), .Z(n3291) );
  NBUFFX2 U3786 ( .INP(n3427), .Z(n3292) );
  NBUFFX2 U3787 ( .INP(n3427), .Z(n3293) );
  NBUFFX2 U3788 ( .INP(n3427), .Z(n3294) );
  NBUFFX2 U3789 ( .INP(n3426), .Z(n3295) );
  NBUFFX2 U3790 ( .INP(n3426), .Z(n3296) );
  NBUFFX2 U3791 ( .INP(n3426), .Z(n3297) );
  NBUFFX2 U3792 ( .INP(n3425), .Z(n3298) );
  NBUFFX2 U3793 ( .INP(n3425), .Z(n3299) );
  NBUFFX2 U3794 ( .INP(n3425), .Z(n3300) );
  NBUFFX2 U3795 ( .INP(n3424), .Z(n3301) );
  NBUFFX2 U3796 ( .INP(n3424), .Z(n3302) );
  NBUFFX2 U3797 ( .INP(n3424), .Z(n3303) );
  NBUFFX2 U3798 ( .INP(n3423), .Z(n3304) );
  NBUFFX2 U3799 ( .INP(n3423), .Z(n3305) );
  NBUFFX2 U3800 ( .INP(n3423), .Z(n3306) );
  NBUFFX2 U3801 ( .INP(n3422), .Z(n3307) );
  NBUFFX2 U3802 ( .INP(n3422), .Z(n3308) );
  NBUFFX2 U3803 ( .INP(n3422), .Z(n3309) );
  NBUFFX2 U3804 ( .INP(n3421), .Z(n3310) );
  NBUFFX2 U3805 ( .INP(n3421), .Z(n3311) );
  NBUFFX2 U3806 ( .INP(n3421), .Z(n3312) );
  NBUFFX2 U3807 ( .INP(n3420), .Z(n3313) );
  NBUFFX2 U3808 ( .INP(n3420), .Z(n3314) );
  NBUFFX2 U3809 ( .INP(n3420), .Z(n3315) );
  NBUFFX2 U3810 ( .INP(n3419), .Z(n3316) );
  NBUFFX2 U3811 ( .INP(n3419), .Z(n3317) );
  NBUFFX2 U3812 ( .INP(n3419), .Z(n3318) );
  NBUFFX2 U3813 ( .INP(n3418), .Z(n3319) );
  NBUFFX2 U3814 ( .INP(n3418), .Z(n3320) );
  NBUFFX2 U3815 ( .INP(n3418), .Z(n3321) );
  NBUFFX2 U3816 ( .INP(n3417), .Z(n3322) );
  NBUFFX2 U3817 ( .INP(n3417), .Z(n3323) );
  NBUFFX2 U3818 ( .INP(n3417), .Z(n3324) );
  NBUFFX2 U3819 ( .INP(n3416), .Z(n3325) );
  NBUFFX2 U3820 ( .INP(n3416), .Z(n3326) );
  NBUFFX2 U3821 ( .INP(n3416), .Z(n3327) );
  NBUFFX2 U3822 ( .INP(n3415), .Z(n3328) );
  NBUFFX2 U3823 ( .INP(n3415), .Z(n3329) );
  NBUFFX2 U3824 ( .INP(n3415), .Z(n3330) );
  NBUFFX2 U3825 ( .INP(n3414), .Z(n3331) );
  NBUFFX2 U3826 ( .INP(n3414), .Z(n3332) );
  NBUFFX2 U3827 ( .INP(n3414), .Z(n3333) );
  NBUFFX2 U3828 ( .INP(n3413), .Z(n3334) );
  NBUFFX2 U3829 ( .INP(n3413), .Z(n3335) );
  NBUFFX2 U3830 ( .INP(n3413), .Z(n3336) );
  NBUFFX2 U3831 ( .INP(n3412), .Z(n3337) );
  NBUFFX2 U3832 ( .INP(n3412), .Z(n3338) );
  NBUFFX2 U3833 ( .INP(n3412), .Z(n3339) );
  NBUFFX2 U3834 ( .INP(n3411), .Z(n3340) );
  NBUFFX2 U3835 ( .INP(n3411), .Z(n3341) );
  NBUFFX2 U3836 ( .INP(n3411), .Z(n3342) );
  NBUFFX2 U3837 ( .INP(n3410), .Z(n3343) );
  NBUFFX2 U3838 ( .INP(n3410), .Z(n3344) );
  NBUFFX2 U3839 ( .INP(n3410), .Z(n3345) );
  NBUFFX2 U3840 ( .INP(n3409), .Z(n3346) );
  NBUFFX2 U3841 ( .INP(n3409), .Z(n3347) );
  NBUFFX2 U3842 ( .INP(n3409), .Z(n3348) );
  NBUFFX2 U3843 ( .INP(n3408), .Z(n3349) );
  NBUFFX2 U3844 ( .INP(n3408), .Z(n3350) );
  NBUFFX2 U3845 ( .INP(n3408), .Z(n3351) );
  NBUFFX2 U3846 ( .INP(n3407), .Z(n3352) );
  NBUFFX2 U3847 ( .INP(n3407), .Z(n3353) );
  NBUFFX2 U3848 ( .INP(n3407), .Z(n3354) );
  NBUFFX2 U3849 ( .INP(n3406), .Z(n3355) );
  NBUFFX2 U3850 ( .INP(n3406), .Z(n3356) );
  NBUFFX2 U3851 ( .INP(n3406), .Z(n3357) );
  NBUFFX2 U3852 ( .INP(n3405), .Z(n3358) );
  NBUFFX2 U3853 ( .INP(n3405), .Z(n3359) );
  NBUFFX2 U3854 ( .INP(n3405), .Z(n3360) );
  NBUFFX2 U3855 ( .INP(n3404), .Z(n3361) );
  NBUFFX2 U3856 ( .INP(n3404), .Z(n3362) );
  NBUFFX2 U3857 ( .INP(n3404), .Z(n3363) );
  NBUFFX2 U3858 ( .INP(n3403), .Z(n3364) );
  NBUFFX2 U3859 ( .INP(n3403), .Z(n3365) );
  NBUFFX2 U3860 ( .INP(n3403), .Z(n3366) );
  NBUFFX2 U3861 ( .INP(n3402), .Z(n3367) );
  NBUFFX2 U3862 ( .INP(n3402), .Z(n3368) );
  NBUFFX2 U3863 ( .INP(n3402), .Z(n3369) );
  NBUFFX2 U3864 ( .INP(n3401), .Z(n3370) );
  NBUFFX2 U3865 ( .INP(n3401), .Z(n3371) );
  NBUFFX2 U3866 ( .INP(n3401), .Z(n3372) );
  NBUFFX2 U3867 ( .INP(n3400), .Z(n3373) );
  NBUFFX2 U3868 ( .INP(n3400), .Z(n3374) );
  NBUFFX2 U3869 ( .INP(n3400), .Z(n3375) );
  NBUFFX2 U3870 ( .INP(n3399), .Z(n3376) );
  NBUFFX2 U3872 ( .INP(n3399), .Z(n3377) );
  NBUFFX2 U3873 ( .INP(n3399), .Z(n3378) );
  NBUFFX2 U3874 ( .INP(n3398), .Z(n3379) );
  NBUFFX2 U3875 ( .INP(n3398), .Z(n3380) );
  NBUFFX2 U3876 ( .INP(n3398), .Z(n3381) );
  NBUFFX2 U3877 ( .INP(n3397), .Z(n3382) );
  NBUFFX2 U3878 ( .INP(n3397), .Z(n3383) );
  NBUFFX2 U3879 ( .INP(n3397), .Z(n3384) );
  NBUFFX2 U3880 ( .INP(n3396), .Z(n3385) );
  NBUFFX2 U3881 ( .INP(n3396), .Z(n3386) );
  NBUFFX2 U3882 ( .INP(n3396), .Z(n3387) );
  NBUFFX2 U3883 ( .INP(n3395), .Z(n3388) );
  NBUFFX2 U3884 ( .INP(n3395), .Z(n3389) );
  NBUFFX2 U3885 ( .INP(n3395), .Z(n3390) );
  NBUFFX2 U3886 ( .INP(n3394), .Z(n3391) );
  NBUFFX2 U3887 ( .INP(n3394), .Z(n3392) );
  NBUFFX2 U3888 ( .INP(n3394), .Z(n3393) );
  NBUFFX2 U3889 ( .INP(n3551), .Z(n3394) );
  NBUFFX2 U3890 ( .INP(n3551), .Z(n3395) );
  NBUFFX2 U3891 ( .INP(n3551), .Z(n3396) );
  NBUFFX2 U3892 ( .INP(n3550), .Z(n3397) );
  NBUFFX2 U3893 ( .INP(n3550), .Z(n3398) );
  NBUFFX2 U3894 ( .INP(n3550), .Z(n3399) );
  NBUFFX2 U3895 ( .INP(n3549), .Z(n3400) );
  NBUFFX2 U3896 ( .INP(n3549), .Z(n3401) );
  NBUFFX2 U3897 ( .INP(n3549), .Z(n3402) );
  NBUFFX2 U3898 ( .INP(n3548), .Z(n3403) );
  NBUFFX2 U3899 ( .INP(n3548), .Z(n3404) );
  NBUFFX2 U3900 ( .INP(n3548), .Z(n3405) );
  NBUFFX2 U3901 ( .INP(n3546), .Z(n3406) );
  NBUFFX2 U3902 ( .INP(n3546), .Z(n3407) );
  NBUFFX2 U3903 ( .INP(n3546), .Z(n3408) );
  NBUFFX2 U3904 ( .INP(n3545), .Z(n3409) );
  NBUFFX2 U3905 ( .INP(n3545), .Z(n3410) );
  NBUFFX2 U3906 ( .INP(n3545), .Z(n3411) );
  NBUFFX2 U3907 ( .INP(n3544), .Z(n3412) );
  NBUFFX2 U3908 ( .INP(n3544), .Z(n3413) );
  NBUFFX2 U3909 ( .INP(n3544), .Z(n3414) );
  NBUFFX2 U3910 ( .INP(n3543), .Z(n3415) );
  NBUFFX2 U3911 ( .INP(n3543), .Z(n3416) );
  NBUFFX2 U3912 ( .INP(n3543), .Z(n3417) );
  NBUFFX2 U3913 ( .INP(n3542), .Z(n3418) );
  NBUFFX2 U3914 ( .INP(n3542), .Z(n3419) );
  NBUFFX2 U3915 ( .INP(n3542), .Z(n3420) );
  NBUFFX2 U3916 ( .INP(n3541), .Z(n3421) );
  NBUFFX2 U3917 ( .INP(n3541), .Z(n3422) );
  NBUFFX2 U3918 ( .INP(n3541), .Z(n3423) );
  NBUFFX2 U3919 ( .INP(n3540), .Z(n3424) );
  NBUFFX2 U3920 ( .INP(n3540), .Z(n3425) );
  NBUFFX2 U3921 ( .INP(n3540), .Z(n3426) );
  NBUFFX2 U3922 ( .INP(n3538), .Z(n3427) );
  NBUFFX2 U3923 ( .INP(n3538), .Z(n3428) );
  NBUFFX2 U3924 ( .INP(n3538), .Z(n3429) );
  NBUFFX2 U3925 ( .INP(n3537), .Z(n3430) );
  NBUFFX2 U3926 ( .INP(n3537), .Z(n3431) );
  NBUFFX2 U3927 ( .INP(n3537), .Z(n3432) );
  NBUFFX2 U3928 ( .INP(n3536), .Z(n3433) );
  NBUFFX2 U3929 ( .INP(n3536), .Z(n3434) );
  NBUFFX2 U3930 ( .INP(n3536), .Z(n3435) );
  NBUFFX2 U3931 ( .INP(n3534), .Z(n3436) );
  NBUFFX2 U3932 ( .INP(n3534), .Z(n3437) );
  NBUFFX2 U3933 ( .INP(n3534), .Z(n3438) );
  NBUFFX2 U3934 ( .INP(n3533), .Z(n3439) );
  NBUFFX2 U3935 ( .INP(n3533), .Z(n3440) );
  NBUFFX2 U3936 ( .INP(n3533), .Z(n3441) );
  NBUFFX2 U3937 ( .INP(n3532), .Z(n3442) );
  NBUFFX2 U3938 ( .INP(n3532), .Z(n3443) );
  NBUFFX2 U3939 ( .INP(n3532), .Z(n3444) );
  NBUFFX2 U3940 ( .INP(n3531), .Z(n3445) );
  NBUFFX2 U3941 ( .INP(n3531), .Z(n3446) );
  NBUFFX2 U3942 ( .INP(n3531), .Z(n3447) );
  NBUFFX2 U3943 ( .INP(n3530), .Z(n3448) );
  NBUFFX2 U3944 ( .INP(n3530), .Z(n3449) );
  NBUFFX2 U3945 ( .INP(n3530), .Z(n3450) );
  NBUFFX2 U3946 ( .INP(n3528), .Z(n3451) );
  NBUFFX2 U3947 ( .INP(n3528), .Z(n3452) );
  NBUFFX2 U3948 ( .INP(n3528), .Z(n3453) );
  NBUFFX2 U3949 ( .INP(n3526), .Z(n3454) );
  NBUFFX2 U3950 ( .INP(n3526), .Z(n3455) );
  NBUFFX2 U3951 ( .INP(n3526), .Z(n3456) );
  NBUFFX2 U3952 ( .INP(n3524), .Z(n3457) );
  NBUFFX2 U3953 ( .INP(n3524), .Z(n3458) );
  NBUFFX2 U3954 ( .INP(n3524), .Z(n3459) );
  NBUFFX2 U3955 ( .INP(n3523), .Z(n3460) );
  NBUFFX2 U3956 ( .INP(n3523), .Z(n3461) );
  NBUFFX2 U3957 ( .INP(n3523), .Z(n3462) );
  NBUFFX2 U3958 ( .INP(n3522), .Z(n3463) );
  NBUFFX2 U3959 ( .INP(n3522), .Z(n3464) );
  NBUFFX2 U3960 ( .INP(n3522), .Z(n3465) );
  NBUFFX2 U3961 ( .INP(n3520), .Z(n3466) );
  NBUFFX2 U3962 ( .INP(n3520), .Z(n3468) );
  NBUFFX2 U3963 ( .INP(n3520), .Z(n3470) );
  NBUFFX2 U3964 ( .INP(n3518), .Z(n3472) );
  NBUFFX2 U3965 ( .INP(n3518), .Z(n3474) );
  NBUFFX2 U3966 ( .INP(n3518), .Z(n3476) );
  NBUFFX2 U3967 ( .INP(n3516), .Z(n3478) );
  NBUFFX2 U3968 ( .INP(n3516), .Z(n3480) );
  NBUFFX2 U3969 ( .INP(n3516), .Z(n3482) );
  NBUFFX2 U3970 ( .INP(n3515), .Z(n3484) );
  NBUFFX2 U3971 ( .INP(n3515), .Z(n3486) );
  NBUFFX2 U3972 ( .INP(n3515), .Z(n3487) );
  NBUFFX2 U3973 ( .INP(n3514), .Z(n3488) );
  NBUFFX2 U3974 ( .INP(n3514), .Z(n3490) );
  NBUFFX2 U3975 ( .INP(n3514), .Z(n3492) );
  NBUFFX2 U3976 ( .INP(n3512), .Z(n3494) );
  NBUFFX2 U3977 ( .INP(n3512), .Z(n3496) );
  NBUFFX2 U3978 ( .INP(n3512), .Z(n3498) );
  NBUFFX2 U3979 ( .INP(n3510), .Z(n3499) );
  NBUFFX2 U3980 ( .INP(n3510), .Z(n3500) );
  NBUFFX2 U3981 ( .INP(n3510), .Z(n3502) );
  NBUFFX2 U3982 ( .INP(n3508), .Z(n3504) );
  NBUFFX2 U3983 ( .INP(n3508), .Z(n3506) );
  NBUFFX2 U3984 ( .INP(n3508), .Z(n3507) );
  NBUFFX2 U3985 ( .INP(n3562), .Z(n3508) );
  NBUFFX2 U3986 ( .INP(n3562), .Z(n3510) );
  NBUFFX2 U3987 ( .INP(n3561), .Z(n3512) );
  NBUFFX2 U3988 ( .INP(n3561), .Z(n3514) );
  NBUFFX2 U3989 ( .INP(n3561), .Z(n3515) );
  NBUFFX2 U3990 ( .INP(n3560), .Z(n3516) );
  NBUFFX2 U3992 ( .INP(n3560), .Z(n3518) );
  NBUFFX2 U3993 ( .INP(n3560), .Z(n3520) );
  NBUFFX2 U3994 ( .INP(n3559), .Z(n3522) );
  NBUFFX2 U3995 ( .INP(n3559), .Z(n3523) );
  NBUFFX2 U3996 ( .INP(n3559), .Z(n3524) );
  NBUFFX2 U3997 ( .INP(n3558), .Z(n3526) );
  NBUFFX2 U3998 ( .INP(n3558), .Z(n3528) );
  NBUFFX2 U3999 ( .INP(n3558), .Z(n3530) );
  NBUFFX2 U4000 ( .INP(n3557), .Z(n3531) );
  NBUFFX2 U4001 ( .INP(n3557), .Z(n3532) );
  NBUFFX2 U4002 ( .INP(n3557), .Z(n3533) );
  NBUFFX2 U4003 ( .INP(n3556), .Z(n3534) );
  NBUFFX2 U4004 ( .INP(n3556), .Z(n3536) );
  NBUFFX2 U4005 ( .INP(n3556), .Z(n3537) );
  NBUFFX2 U4006 ( .INP(n3555), .Z(n3538) );
  NBUFFX2 U4007 ( .INP(n3555), .Z(n3540) );
  NBUFFX2 U4008 ( .INP(n3555), .Z(n3541) );
  NBUFFX2 U4009 ( .INP(n3554), .Z(n3542) );
  NBUFFX2 U4010 ( .INP(n3554), .Z(n3543) );
  NBUFFX2 U4011 ( .INP(n3554), .Z(n3544) );
  NBUFFX2 U4012 ( .INP(n3553), .Z(n3545) );
  NBUFFX2 U4013 ( .INP(n3553), .Z(n3546) );
  NBUFFX2 U4014 ( .INP(n3553), .Z(n3548) );
  NBUFFX2 U4015 ( .INP(n3552), .Z(n3549) );
  NBUFFX2 U4016 ( .INP(n3552), .Z(n3550) );
  NBUFFX2 U4017 ( .INP(n3552), .Z(n3551) );
  NBUFFX2 U4018 ( .INP(n3566), .Z(n3552) );
  NBUFFX2 U4019 ( .INP(n3566), .Z(n3553) );
  NBUFFX2 U4020 ( .INP(n3565), .Z(n3554) );
  NBUFFX2 U4021 ( .INP(n3565), .Z(n3555) );
  NBUFFX2 U4022 ( .INP(n3565), .Z(n3556) );
  NBUFFX2 U4023 ( .INP(n3564), .Z(n3557) );
  NBUFFX2 U4024 ( .INP(n3564), .Z(n3558) );
  NBUFFX2 U4025 ( .INP(n3564), .Z(n3559) );
  NBUFFX2 U4026 ( .INP(n3563), .Z(n3560) );
  NBUFFX2 U4027 ( .INP(n3563), .Z(n3561) );
  NBUFFX2 U4028 ( .INP(n3563), .Z(n3562) );
  NBUFFX2 U4029 ( .INP(test_se), .Z(n3563) );
  NBUFFX2 U4030 ( .INP(test_se), .Z(n3564) );
  NBUFFX2 U4031 ( .INP(test_se), .Z(n3565) );
  NBUFFX2 U4032 ( .INP(test_se), .Z(n3566) );
  NBUFFX2 U4033 ( .INP(n3645), .Z(n3584) );
  NBUFFX2 U4034 ( .INP(n3645), .Z(n3585) );
  NBUFFX2 U4035 ( .INP(n3645), .Z(n3586) );
  NBUFFX2 U4036 ( .INP(n3644), .Z(n3587) );
  NBUFFX2 U4037 ( .INP(n3644), .Z(n3588) );
  NBUFFX2 U4038 ( .INP(n3644), .Z(n3589) );
  NBUFFX2 U4039 ( .INP(n3643), .Z(n3590) );
  NBUFFX2 U4040 ( .INP(n3643), .Z(n3592) );
  NBUFFX2 U4041 ( .INP(n3643), .Z(n3593) );
  NBUFFX2 U4042 ( .INP(n3642), .Z(n3594) );
  NBUFFX2 U4043 ( .INP(n3642), .Z(n3595) );
  NBUFFX2 U4044 ( .INP(n3642), .Z(n3596) );
  NBUFFX2 U4045 ( .INP(n3641), .Z(n3597) );
  NBUFFX2 U4046 ( .INP(n3641), .Z(n3598) );
  NBUFFX2 U4047 ( .INP(n3641), .Z(n3599) );
  NBUFFX2 U4048 ( .INP(n3640), .Z(n3600) );
  NBUFFX2 U4049 ( .INP(n3640), .Z(n3601) );
  NBUFFX2 U4050 ( .INP(n3640), .Z(n3602) );
  NBUFFX2 U4051 ( .INP(n3638), .Z(n3603) );
  NBUFFX2 U4052 ( .INP(n3638), .Z(n3604) );
  NBUFFX2 U4053 ( .INP(n3638), .Z(n3605) );
  NBUFFX2 U4054 ( .INP(n3637), .Z(n3606) );
  NBUFFX2 U4055 ( .INP(n3637), .Z(n3607) );
  NBUFFX2 U4056 ( .INP(n3637), .Z(n3608) );
  NBUFFX2 U4057 ( .INP(n3636), .Z(n3609) );
  NBUFFX2 U4058 ( .INP(n3636), .Z(n3610) );
  NBUFFX2 U4059 ( .INP(n3636), .Z(n3611) );
  NBUFFX2 U4060 ( .INP(n3634), .Z(n3612) );
  NBUFFX2 U4061 ( .INP(n3634), .Z(n3614) );
  NBUFFX2 U4062 ( .INP(n3634), .Z(n3615) );
  NBUFFX2 U4063 ( .INP(n3633), .Z(n3616) );
  NBUFFX2 U4064 ( .INP(n3633), .Z(n3618) );
  NBUFFX2 U4065 ( .INP(n3633), .Z(n3619) );
  NBUFFX2 U4066 ( .INP(n3632), .Z(n3620) );
  NBUFFX2 U4067 ( .INP(n3632), .Z(n3621) );
  NBUFFX2 U4068 ( .INP(n3632), .Z(n3622) );
  NBUFFX2 U4069 ( .INP(n3631), .Z(n3623) );
  NBUFFX2 U4070 ( .INP(n3631), .Z(n3624) );
  NBUFFX2 U4071 ( .INP(n3631), .Z(n3626) );
  NBUFFX2 U4072 ( .INP(n3630), .Z(n3627) );
  NBUFFX2 U4073 ( .INP(n3630), .Z(n3628) );
  NBUFFX2 U4074 ( .INP(n3630), .Z(n3629) );
  NBUFFX2 U4075 ( .INP(n3651), .Z(n3630) );
  NBUFFX2 U4076 ( .INP(n3651), .Z(n3631) );
  NBUFFX2 U4077 ( .INP(n3650), .Z(n3632) );
  NBUFFX2 U4078 ( .INP(n3650), .Z(n3633) );
  NBUFFX2 U4079 ( .INP(n3650), .Z(n3634) );
  NBUFFX2 U4080 ( .INP(n3649), .Z(n3636) );
  NBUFFX2 U4081 ( .INP(n3649), .Z(n3637) );
  NBUFFX2 U4082 ( .INP(n3649), .Z(n3638) );
  NBUFFX2 U4083 ( .INP(n3648), .Z(n3640) );
  NBUFFX2 U4084 ( .INP(n3648), .Z(n3641) );
  NBUFFX2 U4085 ( .INP(n3648), .Z(n3642) );
  NBUFFX2 U4086 ( .INP(n3646), .Z(n3643) );
  NBUFFX2 U4087 ( .INP(n3646), .Z(n3644) );
  NBUFFX2 U4088 ( .INP(n3646), .Z(n3645) );
  NBUFFX2 U4089 ( .INP(RESET), .Z(n3646) );
  NBUFFX2 U4090 ( .INP(RESET), .Z(n3648) );
  NBUFFX2 U4091 ( .INP(RESET), .Z(n3649) );
  NBUFFX2 U4092 ( .INP(RESET), .Z(n3650) );
  NBUFFX2 U4093 ( .INP(RESET), .Z(n3651) );
  INVX0 U4094 ( .INP(n3584), .ZN(n3652) );
  INVX0 U4095 ( .INP(n3584), .ZN(n3653) );
  INVX0 U4096 ( .INP(n3584), .ZN(n3654) );
  INVX0 U4097 ( .INP(n3584), .ZN(n3655) );
  INVX0 U4098 ( .INP(n3584), .ZN(n3656) );
  INVX0 U4099 ( .INP(n3584), .ZN(n3657) );
  INVX0 U4100 ( .INP(n3585), .ZN(n3658) );
  INVX0 U4101 ( .INP(n3585), .ZN(n3659) );
  INVX0 U4102 ( .INP(n3585), .ZN(n3660) );
  INVX0 U4103 ( .INP(n3585), .ZN(n3662) );
  INVX0 U4104 ( .INP(n3586), .ZN(n3663) );
  INVX0 U4105 ( .INP(n3586), .ZN(n3664) );
  INVX0 U4106 ( .INP(n3586), .ZN(n3665) );
  INVX0 U4107 ( .INP(n3590), .ZN(n3666) );
  INVX0 U4108 ( .INP(n3586), .ZN(n3667) );
  INVX0 U4109 ( .INP(n3586), .ZN(n3668) );
  INVX0 U4110 ( .INP(n3586), .ZN(n3670) );
  INVX0 U4111 ( .INP(n3586), .ZN(n3671) );
  INVX0 U4112 ( .INP(n3586), .ZN(n3672) );
  INVX0 U4113 ( .INP(n3587), .ZN(n3673) );
  INVX0 U4114 ( .INP(n3587), .ZN(n3674) );
  INVX0 U4115 ( .INP(n3587), .ZN(n3675) );
  INVX0 U4116 ( .INP(n3587), .ZN(n3676) );
  INVX0 U4117 ( .INP(n3587), .ZN(n3677) );
  INVX0 U4118 ( .INP(n3587), .ZN(n3678) );
  INVX0 U4119 ( .INP(n3587), .ZN(n3679) );
  INVX0 U4120 ( .INP(n3587), .ZN(n3680) );
  INVX0 U4121 ( .INP(n3588), .ZN(n3681) );
  INVX0 U4122 ( .INP(n3588), .ZN(n3682) );
  INVX0 U4123 ( .INP(n3588), .ZN(n3683) );
  INVX0 U4124 ( .INP(n3588), .ZN(n3684) );
  INVX0 U4125 ( .INP(n3588), .ZN(n3685) );
  INVX0 U4126 ( .INP(n3588), .ZN(n3686) );
  INVX0 U4127 ( .INP(n3588), .ZN(n3687) );
  INVX0 U4128 ( .INP(n3588), .ZN(n3688) );
  INVX0 U4129 ( .INP(n3589), .ZN(n3689) );
  INVX0 U4130 ( .INP(n3589), .ZN(n3690) );
  INVX0 U4131 ( .INP(n3589), .ZN(n3692) );
  INVX0 U4132 ( .INP(n3589), .ZN(n3693) );
  INVX0 U4133 ( .INP(n3589), .ZN(n3694) );
  INVX0 U4134 ( .INP(n3589), .ZN(n3695) );
  INVX0 U4135 ( .INP(n3589), .ZN(n3696) );
  INVX0 U4136 ( .INP(n3589), .ZN(n3697) );
  INVX0 U4137 ( .INP(n3590), .ZN(n3698) );
  INVX0 U4138 ( .INP(n3590), .ZN(n3699) );
  INVX0 U4139 ( .INP(n3590), .ZN(n3700) );
  INVX0 U4140 ( .INP(n3590), .ZN(n3701) );
  INVX0 U4141 ( .INP(n3590), .ZN(n3702) );
  INVX0 U4142 ( .INP(n3590), .ZN(n3703) );
  INVX0 U4143 ( .INP(n3590), .ZN(n3704) );
  INVX0 U4144 ( .INP(n3592), .ZN(n3705) );
  INVX0 U4145 ( .INP(n3592), .ZN(n3706) );
  INVX0 U4146 ( .INP(n3592), .ZN(n3707) );
  INVX0 U4147 ( .INP(n3592), .ZN(n3708) );
  INVX0 U4148 ( .INP(n3592), .ZN(n3709) );
  INVX0 U4149 ( .INP(n3592), .ZN(n3710) );
  INVX0 U4150 ( .INP(n3592), .ZN(n3711) );
  INVX0 U4151 ( .INP(n3592), .ZN(n3712) );
  INVX0 U4152 ( .INP(n3593), .ZN(n3714) );
  INVX0 U4153 ( .INP(n3593), .ZN(n3715) );
  INVX0 U4154 ( .INP(n3593), .ZN(n3716) );
  INVX0 U4155 ( .INP(n3593), .ZN(n3718) );
  INVX0 U4156 ( .INP(n3593), .ZN(n3719) );
  INVX0 U4157 ( .INP(n3593), .ZN(n3720) );
  INVX0 U4158 ( .INP(n3593), .ZN(n3721) );
  INVX0 U4159 ( .INP(n3593), .ZN(n3722) );
  INVX0 U4160 ( .INP(n3594), .ZN(n3723) );
  INVX0 U4161 ( .INP(n3594), .ZN(n3724) );
  INVX0 U4162 ( .INP(n3594), .ZN(n3725) );
  INVX0 U4163 ( .INP(n3594), .ZN(n3726) );
  INVX0 U4164 ( .INP(n3594), .ZN(n3727) );
  INVX0 U4165 ( .INP(n3594), .ZN(n3728) );
  INVX0 U4166 ( .INP(n3594), .ZN(n3729) );
  INVX0 U4167 ( .INP(n3594), .ZN(n3730) );
  INVX0 U4168 ( .INP(n3595), .ZN(n3731) );
  INVX0 U4169 ( .INP(n3595), .ZN(n3732) );
  INVX0 U4170 ( .INP(n3595), .ZN(n3733) );
  INVX0 U4171 ( .INP(n3595), .ZN(n3734) );
  INVX0 U4172 ( .INP(n3595), .ZN(n3736) );
  INVX0 U4173 ( .INP(n3595), .ZN(n3737) );
  INVX0 U4174 ( .INP(n3595), .ZN(n3738) );
  INVX0 U4175 ( .INP(n3596), .ZN(n3740) );
  INVX0 U4176 ( .INP(n3596), .ZN(n3741) );
  INVX0 U4177 ( .INP(n3596), .ZN(n3742) );
  INVX0 U4178 ( .INP(n3596), .ZN(n3743) );
  INVX0 U4179 ( .INP(n3596), .ZN(n3744) );
  INVX0 U4180 ( .INP(n3596), .ZN(n3745) );
  INVX0 U4181 ( .INP(n3596), .ZN(n3746) );
  INVX0 U4182 ( .INP(n3596), .ZN(n3747) );
  INVX0 U4183 ( .INP(n3597), .ZN(n3748) );
  INVX0 U4184 ( .INP(n3597), .ZN(n3749) );
  INVX0 U4185 ( .INP(n3597), .ZN(n3750) );
  INVX0 U4186 ( .INP(n3597), .ZN(n3751) );
  INVX0 U4187 ( .INP(n3597), .ZN(n3752) );
  INVX0 U4188 ( .INP(n3597), .ZN(n3753) );
  INVX0 U4189 ( .INP(n3597), .ZN(n3754) );
  INVX0 U4190 ( .INP(n3595), .ZN(n3755) );
  INVX0 U4191 ( .INP(n3584), .ZN(n3756) );
  NBUFFX2 U4192 ( .INP(n3942), .Z(n3904) );
  NBUFFX2 U4193 ( .INP(n3942), .Z(n3905) );
  NBUFFX2 U4194 ( .INP(n3941), .Z(n3906) );
  NBUFFX2 U4195 ( .INP(n3941), .Z(n3907) );
  NBUFFX2 U4196 ( .INP(n3941), .Z(n3908) );
  NBUFFX2 U4197 ( .INP(n3940), .Z(n3909) );
  NBUFFX2 U4198 ( .INP(n3940), .Z(n3910) );
  NBUFFX2 U4199 ( .INP(n3940), .Z(n3911) );
  NBUFFX2 U4200 ( .INP(n3939), .Z(n3912) );
  NBUFFX2 U4201 ( .INP(n3939), .Z(n3913) );
  NBUFFX2 U4202 ( .INP(n3939), .Z(n3914) );
  NBUFFX2 U4203 ( .INP(n3938), .Z(n3915) );
  NBUFFX2 U4204 ( .INP(n3938), .Z(n3916) );
  NBUFFX2 U4205 ( .INP(n3938), .Z(n3917) );
  NBUFFX2 U4206 ( .INP(n3937), .Z(n3918) );
  NBUFFX2 U4207 ( .INP(n3937), .Z(n3919) );
  NBUFFX2 U4208 ( .INP(n3937), .Z(n3920) );
  NBUFFX2 U4209 ( .INP(n3936), .Z(n3921) );
  NBUFFX2 U4210 ( .INP(n3936), .Z(n3922) );
  NBUFFX2 U4211 ( .INP(n3936), .Z(n3923) );
  NBUFFX2 U4212 ( .INP(n3935), .Z(n3924) );
  NBUFFX2 U4213 ( .INP(n3935), .Z(n3925) );
  NBUFFX2 U4214 ( .INP(n3935), .Z(n3926) );
  NBUFFX2 U4215 ( .INP(n3934), .Z(n3927) );
  NBUFFX2 U4216 ( .INP(n3934), .Z(n3928) );
  NBUFFX2 U4217 ( .INP(n3934), .Z(n3929) );
  NBUFFX2 U4218 ( .INP(n3933), .Z(n3930) );
  NBUFFX2 U4219 ( .INP(n3933), .Z(n3931) );
  NBUFFX2 U4220 ( .INP(n3933), .Z(n3932) );
  NBUFFX2 U4221 ( .INP(CK), .Z(n3933) );
  NBUFFX2 U4222 ( .INP(CK), .Z(n3934) );
  NBUFFX2 U4223 ( .INP(n3942), .Z(n3935) );
  NBUFFX2 U4224 ( .INP(CK), .Z(n3936) );
  NBUFFX2 U4225 ( .INP(n3938), .Z(n3937) );
  NBUFFX2 U4226 ( .INP(CK), .Z(n3938) );
  NBUFFX2 U4227 ( .INP(n3933), .Z(n3939) );
  NBUFFX2 U4228 ( .INP(n3934), .Z(n3940) );
  NBUFFX2 U4229 ( .INP(n3936), .Z(n3941) );
  NBUFFX2 U4230 ( .INP(n3771), .Z(n3942) );
  NOR2X0 U4231 ( .IN1(n3579), .IN2(n3652), .QN(n3278) );
  NOR2X0 U4232 ( .IN1(n6005), .IN2(n3652), .QN(WX9789) );
  NOR2X0 U4233 ( .IN1(n6006), .IN2(n3652), .QN(WX9787) );
  NOR2X0 U4234 ( .IN1(n6007), .IN2(n3652), .QN(WX9785) );
  NOR2X0 U4235 ( .IN1(n6008), .IN2(n3652), .QN(WX9783) );
  AND2X1 U4236 ( .IN1(n3602), .IN2(test_so80), .Q(WX9781) );
  NOR2X0 U4237 ( .IN1(n6010), .IN2(n3652), .QN(WX9779) );
  NOR2X0 U4238 ( .IN1(n6011), .IN2(n3652), .QN(WX9777) );
  NOR2X0 U4239 ( .IN1(n6012), .IN2(n3652), .QN(WX9775) );
  NOR2X0 U4240 ( .IN1(n6013), .IN2(n3652), .QN(WX9773) );
  NOR2X0 U4241 ( .IN1(n6014), .IN2(n3652), .QN(WX9771) );
  NOR2X0 U4242 ( .IN1(n6015), .IN2(n3652), .QN(WX9769) );
  NOR2X0 U4243 ( .IN1(n6016), .IN2(n3652), .QN(WX9767) );
  NOR2X0 U4244 ( .IN1(n6017), .IN2(n3653), .QN(WX9765) );
  NOR2X0 U4245 ( .IN1(n6018), .IN2(n3653), .QN(WX9763) );
  NOR2X0 U4246 ( .IN1(n6019), .IN2(n3653), .QN(WX9761) );
  NOR2X0 U4247 ( .IN1(n6020), .IN2(n3653), .QN(WX9759) );
  NAND4X0 U4248 ( .IN1(n3943), .IN2(n3944), .IN3(n3945), .IN4(n3946), .QN(
        WX9757) );
  NAND2X0 U4249 ( .IN1(n3006), .IN2(n3948), .QN(n3946) );
  NAND2X0 U4250 ( .IN1(n3078), .IN2(n3949), .QN(n3945) );
  NAND2X0 U4251 ( .IN1(n3028), .IN2(WX9595), .QN(n3944) );
  NAND2X0 U4252 ( .IN1(n3047), .IN2(CRC_OUT_2_0), .QN(n3943) );
  NAND4X0 U4253 ( .IN1(n3950), .IN2(n3951), .IN3(n3952), .IN4(n3953), .QN(
        WX9755) );
  NAND2X0 U4254 ( .IN1(n3954), .IN2(n3021), .QN(n3953) );
  NAND2X0 U4255 ( .IN1(n3090), .IN2(n3955), .QN(n3952) );
  NAND2X0 U4256 ( .IN1(WX9593), .IN2(n3028), .QN(n3951) );
  NAND2X0 U4257 ( .IN1(n3064), .IN2(CRC_OUT_2_1), .QN(n3950) );
  NAND4X0 U4258 ( .IN1(n3956), .IN2(n3957), .IN3(n3958), .IN4(n3959), .QN(
        WX9753) );
  NAND2X0 U4259 ( .IN1(n3008), .IN2(n3960), .QN(n3959) );
  NAND2X0 U4260 ( .IN1(n3961), .IN2(n3096), .QN(n3958) );
  NAND2X0 U4261 ( .IN1(WX9591), .IN2(n3028), .QN(n3957) );
  NAND2X0 U4262 ( .IN1(test_so87), .IN2(n3070), .QN(n3956) );
  NAND4X0 U4263 ( .IN1(n3962), .IN2(n3963), .IN3(n3964), .IN4(n3965), .QN(
        WX9751) );
  NAND2X0 U4264 ( .IN1(n3966), .IN2(n3020), .QN(n3965) );
  NAND2X0 U4265 ( .IN1(n3087), .IN2(n3967), .QN(n3964) );
  NAND2X0 U4266 ( .IN1(WX9589), .IN2(n3028), .QN(n3963) );
  NAND2X0 U4267 ( .IN1(n3058), .IN2(CRC_OUT_2_3), .QN(n3962) );
  NAND4X0 U4268 ( .IN1(n3968), .IN2(n3969), .IN3(n3970), .IN4(n3971), .QN(
        WX9749) );
  NAND2X0 U4269 ( .IN1(n3008), .IN2(n3972), .QN(n3971) );
  NAND2X0 U4270 ( .IN1(n3973), .IN2(n3097), .QN(n3970) );
  NAND2X0 U4271 ( .IN1(WX9587), .IN2(n3028), .QN(n3969) );
  NAND2X0 U4272 ( .IN1(n3058), .IN2(CRC_OUT_2_4), .QN(n3968) );
  NAND4X0 U4273 ( .IN1(n3974), .IN2(n3975), .IN3(n3976), .IN4(n3977), .QN(
        WX9747) );
  NAND2X0 U4274 ( .IN1(n3008), .IN2(n3978), .QN(n3977) );
  NAND2X0 U4275 ( .IN1(n3087), .IN2(n3979), .QN(n3976) );
  NAND2X0 U4276 ( .IN1(WX9585), .IN2(n3028), .QN(n3975) );
  NAND2X0 U4277 ( .IN1(n3058), .IN2(CRC_OUT_2_5), .QN(n3974) );
  NAND4X0 U4278 ( .IN1(n3980), .IN2(n3981), .IN3(n3982), .IN4(n3983), .QN(
        WX9745) );
  NAND2X0 U4279 ( .IN1(n3008), .IN2(n3984), .QN(n3983) );
  NAND2X0 U4280 ( .IN1(n3985), .IN2(n3097), .QN(n3982) );
  NAND2X0 U4281 ( .IN1(WX9583), .IN2(n3028), .QN(n3981) );
  NAND2X0 U4282 ( .IN1(n3058), .IN2(CRC_OUT_2_6), .QN(n3980) );
  NAND4X0 U4283 ( .IN1(n3986), .IN2(n3987), .IN3(n3988), .IN4(n3989), .QN(
        WX9743) );
  NAND2X0 U4284 ( .IN1(n3008), .IN2(n3990), .QN(n3989) );
  NAND2X0 U4285 ( .IN1(n3087), .IN2(n3991), .QN(n3988) );
  NAND2X0 U4286 ( .IN1(WX9581), .IN2(n3028), .QN(n3987) );
  NAND2X0 U4287 ( .IN1(n3059), .IN2(CRC_OUT_2_7), .QN(n3986) );
  NAND4X0 U4288 ( .IN1(n3992), .IN2(n3993), .IN3(n3994), .IN4(n3995), .QN(
        WX9741) );
  NAND2X0 U4289 ( .IN1(n3007), .IN2(n3996), .QN(n3995) );
  NAND2X0 U4290 ( .IN1(n3997), .IN2(n3096), .QN(n3994) );
  NAND2X0 U4291 ( .IN1(WX9579), .IN2(n3028), .QN(n3993) );
  NAND2X0 U4292 ( .IN1(n3059), .IN2(CRC_OUT_2_8), .QN(n3992) );
  NAND4X0 U4293 ( .IN1(n3998), .IN2(n3999), .IN3(n4000), .IN4(n4001), .QN(
        WX9739) );
  NAND2X0 U4294 ( .IN1(n3007), .IN2(n4002), .QN(n4001) );
  NAND2X0 U4295 ( .IN1(n3087), .IN2(n4003), .QN(n4000) );
  NAND2X0 U4296 ( .IN1(WX9577), .IN2(n3028), .QN(n3999) );
  NAND2X0 U4297 ( .IN1(n3059), .IN2(CRC_OUT_2_9), .QN(n3998) );
  NAND4X0 U4298 ( .IN1(n4004), .IN2(n4005), .IN3(n4006), .IN4(n4007), .QN(
        WX9737) );
  NAND2X0 U4299 ( .IN1(n3007), .IN2(n4008), .QN(n4007) );
  NAND2X0 U4300 ( .IN1(n3087), .IN2(n4009), .QN(n4006) );
  NAND2X0 U4301 ( .IN1(WX9575), .IN2(n3028), .QN(n4005) );
  NAND2X0 U4302 ( .IN1(n3059), .IN2(CRC_OUT_2_10), .QN(n4004) );
  NAND4X0 U4303 ( .IN1(n4010), .IN2(n4011), .IN3(n4012), .IN4(n4013), .QN(
        WX9735) );
  NAND2X0 U4304 ( .IN1(n3007), .IN2(n4014), .QN(n4013) );
  NAND2X0 U4305 ( .IN1(n3087), .IN2(n4015), .QN(n4012) );
  NAND2X0 U4306 ( .IN1(WX9573), .IN2(n3028), .QN(n4011) );
  NAND2X0 U4307 ( .IN1(n3059), .IN2(CRC_OUT_2_11), .QN(n4010) );
  NAND4X0 U4308 ( .IN1(n4016), .IN2(n4017), .IN3(n4018), .IN4(n4019), .QN(
        WX9733) );
  NAND2X0 U4309 ( .IN1(n3007), .IN2(n4020), .QN(n4019) );
  NAND2X0 U4310 ( .IN1(n3087), .IN2(n4021), .QN(n4018) );
  NAND2X0 U4311 ( .IN1(WX9571), .IN2(n3028), .QN(n4017) );
  NAND2X0 U4312 ( .IN1(n3059), .IN2(CRC_OUT_2_12), .QN(n4016) );
  NAND4X0 U4313 ( .IN1(n4022), .IN2(n4023), .IN3(n4024), .IN4(n4025), .QN(
        WX9731) );
  NAND2X0 U4314 ( .IN1(n3007), .IN2(n4026), .QN(n4025) );
  NAND2X0 U4315 ( .IN1(n3088), .IN2(n4027), .QN(n4024) );
  NAND2X0 U4316 ( .IN1(WX9569), .IN2(n3028), .QN(n4023) );
  NAND2X0 U4317 ( .IN1(n3059), .IN2(CRC_OUT_2_13), .QN(n4022) );
  NAND4X0 U4318 ( .IN1(n4028), .IN2(n4029), .IN3(n4030), .IN4(n4031), .QN(
        WX9729) );
  NAND2X0 U4319 ( .IN1(n4032), .IN2(n3020), .QN(n4031) );
  NAND2X0 U4320 ( .IN1(n3088), .IN2(n4033), .QN(n4030) );
  NAND2X0 U4321 ( .IN1(WX9567), .IN2(n3028), .QN(n4029) );
  NAND2X0 U4322 ( .IN1(n3059), .IN2(CRC_OUT_2_14), .QN(n4028) );
  NAND4X0 U4323 ( .IN1(n4034), .IN2(n4035), .IN3(n4036), .IN4(n4037), .QN(
        WX9727) );
  NAND2X0 U4324 ( .IN1(n3007), .IN2(n4038), .QN(n4037) );
  NAND2X0 U4325 ( .IN1(n3088), .IN2(n4039), .QN(n4036) );
  NAND2X0 U4326 ( .IN1(WX9565), .IN2(n3028), .QN(n4035) );
  NAND2X0 U4327 ( .IN1(n3059), .IN2(CRC_OUT_2_15), .QN(n4034) );
  NAND4X0 U4328 ( .IN1(n4040), .IN2(n4041), .IN3(n4042), .IN4(n4043), .QN(
        WX9725) );
  NAND2X0 U4329 ( .IN1(n4044), .IN2(n3020), .QN(n4043) );
  NAND2X0 U4330 ( .IN1(n3088), .IN2(n4045), .QN(n4042) );
  NAND2X0 U4331 ( .IN1(WX9563), .IN2(n3029), .QN(n4041) );
  NAND2X0 U4332 ( .IN1(n3059), .IN2(CRC_OUT_2_16), .QN(n4040) );
  NAND4X0 U4333 ( .IN1(n4046), .IN2(n4047), .IN3(n4048), .IN4(n4049), .QN(
        WX9723) );
  NAND2X0 U4334 ( .IN1(n3007), .IN2(n4050), .QN(n4049) );
  NAND2X0 U4335 ( .IN1(n3088), .IN2(n4051), .QN(n4048) );
  NAND2X0 U4336 ( .IN1(WX9561), .IN2(n3029), .QN(n4047) );
  NAND2X0 U4337 ( .IN1(n3059), .IN2(CRC_OUT_2_17), .QN(n4046) );
  NAND4X0 U4338 ( .IN1(n4052), .IN2(n4053), .IN3(n4054), .IN4(n4055), .QN(
        WX9721) );
  NAND2X0 U4339 ( .IN1(n4056), .IN2(n3020), .QN(n4055) );
  NAND2X0 U4340 ( .IN1(n3088), .IN2(n4057), .QN(n4054) );
  NAND2X0 U4341 ( .IN1(WX9559), .IN2(n3029), .QN(n4053) );
  NAND2X0 U4342 ( .IN1(n3059), .IN2(CRC_OUT_2_18), .QN(n4052) );
  NAND4X0 U4343 ( .IN1(n4058), .IN2(n4059), .IN3(n4060), .IN4(n4061), .QN(
        WX9719) );
  NAND2X0 U4344 ( .IN1(n3007), .IN2(n4062), .QN(n4061) );
  NAND2X0 U4345 ( .IN1(n4063), .IN2(n3097), .QN(n4060) );
  NAND2X0 U4346 ( .IN1(WX9557), .IN2(n3029), .QN(n4059) );
  NAND2X0 U4347 ( .IN1(test_so88), .IN2(n3069), .QN(n4058) );
  NAND4X0 U4348 ( .IN1(n4064), .IN2(n4065), .IN3(n4066), .IN4(n4067), .QN(
        WX9717) );
  NAND2X0 U4349 ( .IN1(n4068), .IN2(n3020), .QN(n4067) );
  NAND2X0 U4350 ( .IN1(n3088), .IN2(n4069), .QN(n4066) );
  NAND2X0 U4351 ( .IN1(WX9555), .IN2(n3029), .QN(n4065) );
  NAND2X0 U4352 ( .IN1(n3060), .IN2(CRC_OUT_2_20), .QN(n4064) );
  NAND4X0 U4353 ( .IN1(n4070), .IN2(n4071), .IN3(n4072), .IN4(n4073), .QN(
        WX9715) );
  NAND2X0 U4354 ( .IN1(n3007), .IN2(n4074), .QN(n4073) );
  NAND2X0 U4355 ( .IN1(n4075), .IN2(n3098), .QN(n4072) );
  NAND2X0 U4356 ( .IN1(WX9553), .IN2(n3029), .QN(n4071) );
  NAND2X0 U4357 ( .IN1(n3060), .IN2(CRC_OUT_2_21), .QN(n4070) );
  NAND4X0 U4358 ( .IN1(n4076), .IN2(n4077), .IN3(n4078), .IN4(n4079), .QN(
        WX9713) );
  NAND2X0 U4359 ( .IN1(n3007), .IN2(n4080), .QN(n4079) );
  NAND2X0 U4360 ( .IN1(n3088), .IN2(n4081), .QN(n4078) );
  NAND2X0 U4361 ( .IN1(WX9551), .IN2(n3029), .QN(n4077) );
  NAND2X0 U4362 ( .IN1(n3060), .IN2(CRC_OUT_2_22), .QN(n4076) );
  NAND4X0 U4363 ( .IN1(n4082), .IN2(n4083), .IN3(n4084), .IN4(n4085), .QN(
        WX9711) );
  NAND2X0 U4364 ( .IN1(n3007), .IN2(n4086), .QN(n4085) );
  NAND2X0 U4365 ( .IN1(n4087), .IN2(n3098), .QN(n4084) );
  NAND2X0 U4366 ( .IN1(WX9549), .IN2(n3029), .QN(n4083) );
  NAND2X0 U4367 ( .IN1(n3060), .IN2(CRC_OUT_2_23), .QN(n4082) );
  NAND4X0 U4368 ( .IN1(n4088), .IN2(n4089), .IN3(n4090), .IN4(n4091), .QN(
        WX9709) );
  NAND2X0 U4369 ( .IN1(n3006), .IN2(n4092), .QN(n4091) );
  NAND2X0 U4370 ( .IN1(n3088), .IN2(n4093), .QN(n4090) );
  NAND2X0 U4371 ( .IN1(WX9547), .IN2(n3029), .QN(n4089) );
  NAND2X0 U4372 ( .IN1(n3060), .IN2(CRC_OUT_2_24), .QN(n4088) );
  NAND4X0 U4373 ( .IN1(n4094), .IN2(n4095), .IN3(n4096), .IN4(n4097), .QN(
        WX9707) );
  NAND2X0 U4374 ( .IN1(n3006), .IN2(n4098), .QN(n4097) );
  NAND2X0 U4375 ( .IN1(n4099), .IN2(n3098), .QN(n4096) );
  NAND2X0 U4376 ( .IN1(WX9545), .IN2(n3029), .QN(n4095) );
  NAND2X0 U4377 ( .IN1(n3060), .IN2(CRC_OUT_2_25), .QN(n4094) );
  NAND4X0 U4378 ( .IN1(n4100), .IN2(n4101), .IN3(n4102), .IN4(n4103), .QN(
        WX9705) );
  NAND2X0 U4379 ( .IN1(n3006), .IN2(n4104), .QN(n4103) );
  NAND2X0 U4380 ( .IN1(n3088), .IN2(n4105), .QN(n4102) );
  NAND2X0 U4381 ( .IN1(WX9543), .IN2(n3029), .QN(n4101) );
  NAND2X0 U4382 ( .IN1(n3060), .IN2(CRC_OUT_2_26), .QN(n4100) );
  NAND4X0 U4383 ( .IN1(n4106), .IN2(n4107), .IN3(n4108), .IN4(n4109), .QN(
        WX9703) );
  NAND2X0 U4384 ( .IN1(n3006), .IN2(n4110), .QN(n4109) );
  NAND2X0 U4385 ( .IN1(n3088), .IN2(n4111), .QN(n4108) );
  NAND2X0 U4386 ( .IN1(WX9541), .IN2(n3029), .QN(n4107) );
  NAND2X0 U4387 ( .IN1(n3060), .IN2(CRC_OUT_2_27), .QN(n4106) );
  NAND4X0 U4388 ( .IN1(n4112), .IN2(n4113), .IN3(n4114), .IN4(n4115), .QN(
        WX9701) );
  NAND2X0 U4389 ( .IN1(n3006), .IN2(n4116), .QN(n4115) );
  NAND2X0 U4390 ( .IN1(n3088), .IN2(n4117), .QN(n4114) );
  NAND2X0 U4391 ( .IN1(WX9539), .IN2(n3029), .QN(n4113) );
  NAND2X0 U4392 ( .IN1(n3060), .IN2(CRC_OUT_2_28), .QN(n4112) );
  NAND4X0 U4393 ( .IN1(n4118), .IN2(n4119), .IN3(n4120), .IN4(n4121), .QN(
        WX9699) );
  NAND2X0 U4394 ( .IN1(n3006), .IN2(n4122), .QN(n4121) );
  NAND2X0 U4395 ( .IN1(n3089), .IN2(n4123), .QN(n4120) );
  NAND2X0 U4396 ( .IN1(WX9537), .IN2(n3029), .QN(n4119) );
  NAND2X0 U4397 ( .IN1(n3060), .IN2(CRC_OUT_2_29), .QN(n4118) );
  NAND4X0 U4398 ( .IN1(n4124), .IN2(n4125), .IN3(n4126), .IN4(n4127), .QN(
        WX9697) );
  NAND2X0 U4399 ( .IN1(n3006), .IN2(n4128), .QN(n4127) );
  NAND2X0 U4400 ( .IN1(n3089), .IN2(n4129), .QN(n4126) );
  NAND2X0 U4401 ( .IN1(WX9535), .IN2(n3029), .QN(n4125) );
  NAND2X0 U4402 ( .IN1(n3060), .IN2(CRC_OUT_2_30), .QN(n4124) );
  NAND4X0 U4403 ( .IN1(n4130), .IN2(n4131), .IN3(n4132), .IN4(n4133), .QN(
        WX9695) );
  NAND2X0 U4404 ( .IN1(n4134), .IN2(n3019), .QN(n4133) );
  NAND2X0 U4405 ( .IN1(n3089), .IN2(n4135), .QN(n4132) );
  NAND2X0 U4406 ( .IN1(n3060), .IN2(CRC_OUT_2_31), .QN(n4131) );
  NAND2X0 U4407 ( .IN1(n2245), .IN2(WX9536), .QN(n4130) );
  NOR2X0 U4408 ( .IN1(n3736), .IN2(WX9536), .QN(WX9597) );
  AND2X1 U4409 ( .IN1(n3601), .IN2(n8321), .Q(WX9595) );
  AND2X1 U4410 ( .IN1(n3601), .IN2(n8322), .Q(WX9593) );
  AND2X1 U4411 ( .IN1(n3601), .IN2(n8323), .Q(WX9591) );
  AND2X1 U4412 ( .IN1(n3600), .IN2(n8324), .Q(WX9589) );
  AND2X1 U4413 ( .IN1(n3601), .IN2(n8325), .Q(WX9587) );
  AND2X1 U4414 ( .IN1(test_so79), .IN2(n3598), .Q(WX9585) );
  AND2X1 U4415 ( .IN1(n3601), .IN2(n8328), .Q(WX9583) );
  AND2X1 U4416 ( .IN1(n3600), .IN2(n8329), .Q(WX9581) );
  AND2X1 U4417 ( .IN1(n3601), .IN2(n8330), .Q(WX9579) );
  AND2X1 U4418 ( .IN1(n3600), .IN2(n8331), .Q(WX9577) );
  AND2X1 U4419 ( .IN1(n3601), .IN2(n8332), .Q(WX9575) );
  AND2X1 U4420 ( .IN1(n3600), .IN2(n8333), .Q(WX9573) );
  AND2X1 U4421 ( .IN1(n3600), .IN2(n8334), .Q(WX9571) );
  AND2X1 U4422 ( .IN1(n3600), .IN2(n8335), .Q(WX9569) );
  AND2X1 U4423 ( .IN1(n3600), .IN2(n8336), .Q(WX9567) );
  AND2X1 U4424 ( .IN1(n3599), .IN2(n8337), .Q(WX9565) );
  AND2X1 U4425 ( .IN1(n3599), .IN2(n8338), .Q(WX9563) );
  AND2X1 U4426 ( .IN1(n3600), .IN2(n8339), .Q(WX9561) );
  AND2X1 U4427 ( .IN1(n3606), .IN2(n8340), .Q(WX9559) );
  AND2X1 U4428 ( .IN1(n3629), .IN2(n8341), .Q(WX9557) );
  AND2X1 U4429 ( .IN1(n3629), .IN2(n8342), .Q(WX9555) );
  AND2X1 U4430 ( .IN1(n3628), .IN2(n8343), .Q(WX9553) );
  AND2X1 U4431 ( .IN1(test_so78), .IN2(n3597), .Q(WX9551) );
  AND2X1 U4432 ( .IN1(n3628), .IN2(n8346), .Q(WX9549) );
  AND2X1 U4433 ( .IN1(n3628), .IN2(n8347), .Q(WX9547) );
  AND2X1 U4434 ( .IN1(n3628), .IN2(n8348), .Q(WX9545) );
  AND2X1 U4435 ( .IN1(n3628), .IN2(n8349), .Q(WX9543) );
  AND2X1 U4436 ( .IN1(n3628), .IN2(n8350), .Q(WX9541) );
  AND2X1 U4437 ( .IN1(n3628), .IN2(n8351), .Q(WX9539) );
  AND2X1 U4438 ( .IN1(n3628), .IN2(n8352), .Q(WX9537) );
  AND2X1 U4439 ( .IN1(n3627), .IN2(n8353), .Q(WX9535) );
  NOR2X0 U4440 ( .IN1(n3751), .IN2(n4136), .QN(WX9084) );
  XOR2X1 U4441 ( .IN1(n2766), .IN2(DFF_1342_n1), .Q(n4136) );
  NOR2X0 U4442 ( .IN1(n3745), .IN2(n4137), .QN(WX9082) );
  XOR2X1 U4443 ( .IN1(n2767), .IN2(DFF_1341_n1), .Q(n4137) );
  NOR2X0 U4444 ( .IN1(n3745), .IN2(n4138), .QN(WX9080) );
  XOR2X1 U4445 ( .IN1(n2768), .IN2(DFF_1340_n1), .Q(n4138) );
  NOR2X0 U4446 ( .IN1(n3745), .IN2(n4139), .QN(WX9078) );
  XOR2X1 U4447 ( .IN1(n2769), .IN2(DFF_1339_n1), .Q(n4139) );
  NOR2X0 U4448 ( .IN1(n3745), .IN2(n4140), .QN(WX9076) );
  XOR2X1 U4449 ( .IN1(n2770), .IN2(DFF_1338_n1), .Q(n4140) );
  NOR2X0 U4450 ( .IN1(n3745), .IN2(n4141), .QN(WX9074) );
  XOR2X1 U4451 ( .IN1(CRC_OUT_3_25), .IN2(test_so74), .Q(n4141) );
  NOR2X0 U4452 ( .IN1(n3745), .IN2(n4142), .QN(WX9072) );
  XNOR2X1 U4453 ( .IN1(n2771), .IN2(test_so77), .Q(n4142) );
  NOR2X0 U4454 ( .IN1(n3745), .IN2(n4143), .QN(WX9070) );
  XOR2X1 U4455 ( .IN1(n2772), .IN2(DFF_1335_n1), .Q(n4143) );
  NOR2X0 U4456 ( .IN1(n3745), .IN2(n4144), .QN(WX9068) );
  XOR2X1 U4457 ( .IN1(n2773), .IN2(DFF_1334_n1), .Q(n4144) );
  NOR2X0 U4458 ( .IN1(n3745), .IN2(n4145), .QN(WX9066) );
  XOR2X1 U4459 ( .IN1(n2774), .IN2(DFF_1333_n1), .Q(n4145) );
  NOR2X0 U4460 ( .IN1(n3745), .IN2(n4146), .QN(WX9064) );
  XOR2X1 U4461 ( .IN1(n2775), .IN2(DFF_1332_n1), .Q(n4146) );
  NOR2X0 U4462 ( .IN1(n3745), .IN2(n4147), .QN(WX9062) );
  XOR2X1 U4463 ( .IN1(n2776), .IN2(DFF_1331_n1), .Q(n4147) );
  NOR2X0 U4464 ( .IN1(n3746), .IN2(n4148), .QN(WX9060) );
  XOR2X1 U4465 ( .IN1(n2777), .IN2(DFF_1330_n1), .Q(n4148) );
  NOR2X0 U4466 ( .IN1(n3746), .IN2(n4149), .QN(WX9058) );
  XOR2X1 U4467 ( .IN1(n2778), .IN2(DFF_1329_n1), .Q(n4149) );
  NOR2X0 U4468 ( .IN1(n3746), .IN2(n4150), .QN(WX9056) );
  XOR2X1 U4469 ( .IN1(n2779), .IN2(DFF_1328_n1), .Q(n4150) );
  NOR2X0 U4470 ( .IN1(n3746), .IN2(n4151), .QN(WX9054) );
  XOR3X1 U4471 ( .IN1(n2691), .IN2(DFF_1343_n1), .IN3(CRC_OUT_3_15), .Q(n4151)
         );
  NOR2X0 U4472 ( .IN1(n3746), .IN2(n4152), .QN(WX9052) );
  XOR2X1 U4473 ( .IN1(n2780), .IN2(DFF_1326_n1), .Q(n4152) );
  NOR2X0 U4474 ( .IN1(n3746), .IN2(n4153), .QN(WX9050) );
  XOR2X1 U4475 ( .IN1(n2781), .IN2(DFF_1325_n1), .Q(n4153) );
  NOR2X0 U4476 ( .IN1(n3746), .IN2(n4154), .QN(WX9048) );
  XOR2X1 U4477 ( .IN1(n2782), .IN2(DFF_1324_n1), .Q(n4154) );
  NOR2X0 U4478 ( .IN1(n3746), .IN2(n4155), .QN(WX9046) );
  XOR2X1 U4479 ( .IN1(n2783), .IN2(DFF_1323_n1), .Q(n4155) );
  NOR2X0 U4480 ( .IN1(n3746), .IN2(n4156), .QN(WX9044) );
  XOR3X1 U4481 ( .IN1(n2692), .IN2(DFF_1343_n1), .IN3(CRC_OUT_3_10), .Q(n4156)
         );
  NOR2X0 U4482 ( .IN1(n3746), .IN2(n4157), .QN(WX9042) );
  XOR2X1 U4483 ( .IN1(n2784), .IN2(DFF_1321_n1), .Q(n4157) );
  NOR2X0 U4484 ( .IN1(n3746), .IN2(n4158), .QN(WX9040) );
  XOR2X1 U4485 ( .IN1(CRC_OUT_3_8), .IN2(test_so75), .Q(n4158) );
  NOR2X0 U4486 ( .IN1(n3746), .IN2(n4159), .QN(WX9038) );
  XNOR2X1 U4487 ( .IN1(n2785), .IN2(test_so76), .Q(n4159) );
  NOR2X0 U4488 ( .IN1(n3746), .IN2(n4160), .QN(WX9036) );
  XOR2X1 U4489 ( .IN1(n2786), .IN2(DFF_1318_n1), .Q(n4160) );
  NOR2X0 U4490 ( .IN1(n3747), .IN2(n4161), .QN(WX9034) );
  XOR2X1 U4491 ( .IN1(n2787), .IN2(DFF_1317_n1), .Q(n4161) );
  NOR2X0 U4492 ( .IN1(n3747), .IN2(n4162), .QN(WX9032) );
  XOR2X1 U4493 ( .IN1(n2788), .IN2(DFF_1316_n1), .Q(n4162) );
  NOR2X0 U4494 ( .IN1(n3747), .IN2(n4163), .QN(WX9030) );
  XOR3X1 U4495 ( .IN1(n2693), .IN2(DFF_1343_n1), .IN3(CRC_OUT_3_3), .Q(n4163)
         );
  NOR2X0 U4496 ( .IN1(n3747), .IN2(n4164), .QN(WX9028) );
  XOR2X1 U4497 ( .IN1(n2789), .IN2(DFF_1314_n1), .Q(n4164) );
  NOR2X0 U4498 ( .IN1(n3747), .IN2(n4165), .QN(WX9026) );
  XOR2X1 U4499 ( .IN1(n2790), .IN2(DFF_1313_n1), .Q(n4165) );
  NOR2X0 U4500 ( .IN1(n3747), .IN2(n4166), .QN(WX9024) );
  XOR2X1 U4501 ( .IN1(n2791), .IN2(DFF_1312_n1), .Q(n4166) );
  NOR2X0 U4502 ( .IN1(n3747), .IN2(n4167), .QN(WX9022) );
  XOR2X1 U4503 ( .IN1(n2708), .IN2(DFF_1343_n1), .Q(n4167) );
  NOR2X0 U4504 ( .IN1(n6033), .IN2(n3653), .QN(WX8496) );
  NOR2X0 U4505 ( .IN1(n6034), .IN2(n3653), .QN(WX8494) );
  NOR2X0 U4506 ( .IN1(n6035), .IN2(n3653), .QN(WX8492) );
  NOR2X0 U4507 ( .IN1(n6036), .IN2(n3653), .QN(WX8490) );
  NOR2X0 U4508 ( .IN1(n6037), .IN2(n3653), .QN(WX8488) );
  NOR2X0 U4509 ( .IN1(n6038), .IN2(n3653), .QN(WX8486) );
  NOR2X0 U4510 ( .IN1(n6039), .IN2(n3653), .QN(WX8484) );
  NOR2X0 U4511 ( .IN1(n6040), .IN2(n3653), .QN(WX8482) );
  NOR2X0 U4512 ( .IN1(n6041), .IN2(n3654), .QN(WX8480) );
  NOR2X0 U4513 ( .IN1(n6042), .IN2(n3654), .QN(WX8478) );
  NOR2X0 U4514 ( .IN1(n6043), .IN2(n3654), .QN(WX8476) );
  NOR2X0 U4515 ( .IN1(n6044), .IN2(n3654), .QN(WX8474) );
  NOR2X0 U4516 ( .IN1(n6045), .IN2(n3654), .QN(WX8472) );
  NOR2X0 U4517 ( .IN1(n6046), .IN2(n3654), .QN(WX8470) );
  NOR2X0 U4518 ( .IN1(n6047), .IN2(n3654), .QN(WX8468) );
  NOR2X0 U4519 ( .IN1(n6048), .IN2(n3654), .QN(WX8466) );
  NAND4X0 U4520 ( .IN1(n4168), .IN2(n4169), .IN3(n4170), .IN4(n4171), .QN(
        WX8464) );
  NAND2X0 U4521 ( .IN1(n3089), .IN2(n3948), .QN(n4171) );
  XNOR3X1 U4522 ( .IN1(n2707), .IN2(n2576), .IN3(n4172), .Q(n3948) );
  XOR2X1 U4523 ( .IN1(WX9822), .IN2(n5992), .Q(n4172) );
  NAND2X0 U4524 ( .IN1(n3006), .IN2(n4173), .QN(n4170) );
  NAND2X0 U4525 ( .IN1(WX8302), .IN2(n3029), .QN(n4169) );
  NAND2X0 U4526 ( .IN1(n3061), .IN2(CRC_OUT_3_0), .QN(n4168) );
  NAND4X0 U4527 ( .IN1(n4174), .IN2(n4175), .IN3(n4176), .IN4(n4177), .QN(
        WX8462) );
  NAND2X0 U4528 ( .IN1(n3954), .IN2(n3098), .QN(n4177) );
  XOR3X1 U4529 ( .IN1(n2765), .IN2(n2577), .IN3(n4178), .Q(n3954) );
  XOR2X1 U4530 ( .IN1(WX9756), .IN2(test_so83), .Q(n4178) );
  NAND2X0 U4531 ( .IN1(n3006), .IN2(n4179), .QN(n4176) );
  NAND2X0 U4532 ( .IN1(WX8300), .IN2(n3029), .QN(n4175) );
  NAND2X0 U4533 ( .IN1(n3061), .IN2(CRC_OUT_3_1), .QN(n4174) );
  NAND4X0 U4534 ( .IN1(n4180), .IN2(n4181), .IN3(n4182), .IN4(n4183), .QN(
        WX8460) );
  NAND2X0 U4535 ( .IN1(n3089), .IN2(n3960), .QN(n4183) );
  XNOR3X1 U4536 ( .IN1(n2764), .IN2(n2578), .IN3(n4184), .Q(n3960) );
  XOR2X1 U4537 ( .IN1(WX9818), .IN2(n5993), .Q(n4184) );
  NAND2X0 U4538 ( .IN1(n3006), .IN2(n4185), .QN(n4182) );
  NAND2X0 U4539 ( .IN1(WX8298), .IN2(n3030), .QN(n4181) );
  NAND2X0 U4540 ( .IN1(n3061), .IN2(CRC_OUT_3_2), .QN(n4180) );
  NAND4X0 U4541 ( .IN1(n4186), .IN2(n4187), .IN3(n4188), .IN4(n4189), .QN(
        WX8458) );
  NAND2X0 U4542 ( .IN1(n3966), .IN2(n3098), .QN(n4189) );
  XOR3X1 U4543 ( .IN1(n3569), .IN2(n2763), .IN3(n4190), .Q(n3966) );
  XOR2X1 U4544 ( .IN1(WX9880), .IN2(test_so81), .Q(n4190) );
  NAND2X0 U4545 ( .IN1(n3006), .IN2(n4191), .QN(n4188) );
  NAND2X0 U4546 ( .IN1(WX8296), .IN2(n3030), .QN(n4187) );
  NAND2X0 U4547 ( .IN1(n3061), .IN2(CRC_OUT_3_3), .QN(n4186) );
  NAND4X0 U4548 ( .IN1(n4192), .IN2(n4193), .IN3(n4194), .IN4(n4195), .QN(
        WX8456) );
  NAND2X0 U4549 ( .IN1(n3089), .IN2(n3972), .QN(n4195) );
  XNOR3X1 U4550 ( .IN1(n2690), .IN2(n2579), .IN3(n4196), .Q(n3972) );
  XOR2X1 U4551 ( .IN1(WX9814), .IN2(n5994), .Q(n4196) );
  NAND2X0 U4552 ( .IN1(n3008), .IN2(n4197), .QN(n4194) );
  NAND2X0 U4553 ( .IN1(WX8294), .IN2(n3030), .QN(n4193) );
  NAND2X0 U4554 ( .IN1(n3061), .IN2(CRC_OUT_3_4), .QN(n4192) );
  NAND4X0 U4555 ( .IN1(n4198), .IN2(n4199), .IN3(n4200), .IN4(n4201), .QN(
        WX8454) );
  NAND2X0 U4556 ( .IN1(n3089), .IN2(n3978), .QN(n4201) );
  XNOR3X1 U4557 ( .IN1(n2762), .IN2(n2580), .IN3(n4202), .Q(n3978) );
  XOR2X1 U4558 ( .IN1(WX9812), .IN2(n5995), .Q(n4202) );
  NAND2X0 U4559 ( .IN1(n3005), .IN2(n4203), .QN(n4200) );
  NAND2X0 U4560 ( .IN1(WX8292), .IN2(n3030), .QN(n4199) );
  NAND2X0 U4561 ( .IN1(n3061), .IN2(CRC_OUT_3_5), .QN(n4198) );
  NAND4X0 U4562 ( .IN1(n4204), .IN2(n4205), .IN3(n4206), .IN4(n4207), .QN(
        WX8452) );
  NAND2X0 U4563 ( .IN1(n3089), .IN2(n3984), .QN(n4207) );
  XNOR3X1 U4564 ( .IN1(n2761), .IN2(n2581), .IN3(n4208), .Q(n3984) );
  XOR2X1 U4565 ( .IN1(WX9810), .IN2(n5996), .Q(n4208) );
  NAND2X0 U4566 ( .IN1(n3005), .IN2(n4209), .QN(n4206) );
  NAND2X0 U4567 ( .IN1(WX8290), .IN2(n3030), .QN(n4205) );
  NAND2X0 U4568 ( .IN1(n3061), .IN2(CRC_OUT_3_6), .QN(n4204) );
  NAND4X0 U4569 ( .IN1(n4210), .IN2(n4211), .IN3(n4212), .IN4(n4213), .QN(
        WX8450) );
  NAND2X0 U4570 ( .IN1(n3089), .IN2(n3990), .QN(n4213) );
  XNOR3X1 U4571 ( .IN1(n2760), .IN2(n2582), .IN3(n4214), .Q(n3990) );
  XOR2X1 U4572 ( .IN1(WX9808), .IN2(n5997), .Q(n4214) );
  NAND2X0 U4573 ( .IN1(n3005), .IN2(n4215), .QN(n4212) );
  NAND2X0 U4574 ( .IN1(WX8288), .IN2(n3030), .QN(n4211) );
  NAND2X0 U4575 ( .IN1(test_so76), .IN2(n3070), .QN(n4210) );
  NAND4X0 U4576 ( .IN1(n4216), .IN2(n4217), .IN3(n4218), .IN4(n4219), .QN(
        WX8448) );
  NAND2X0 U4577 ( .IN1(n3089), .IN2(n3996), .QN(n4219) );
  XNOR3X1 U4578 ( .IN1(n2759), .IN2(n2583), .IN3(n4220), .Q(n3996) );
  XOR2X1 U4579 ( .IN1(WX9806), .IN2(n5998), .Q(n4220) );
  NAND2X0 U4580 ( .IN1(n3005), .IN2(n4221), .QN(n4218) );
  NAND2X0 U4581 ( .IN1(WX8286), .IN2(n3030), .QN(n4217) );
  NAND2X0 U4582 ( .IN1(n3061), .IN2(CRC_OUT_3_8), .QN(n4216) );
  NAND4X0 U4583 ( .IN1(n4222), .IN2(n4223), .IN3(n4224), .IN4(n4225), .QN(
        WX8446) );
  NAND2X0 U4584 ( .IN1(n3089), .IN2(n4002), .QN(n4225) );
  XNOR3X1 U4585 ( .IN1(n2758), .IN2(n2584), .IN3(n4226), .Q(n4002) );
  XOR2X1 U4586 ( .IN1(WX9804), .IN2(n5999), .Q(n4226) );
  NAND2X0 U4587 ( .IN1(n4227), .IN2(n3018), .QN(n4224) );
  NAND2X0 U4588 ( .IN1(WX8284), .IN2(n3030), .QN(n4223) );
  NAND2X0 U4589 ( .IN1(n3061), .IN2(CRC_OUT_3_9), .QN(n4222) );
  NAND4X0 U4590 ( .IN1(n4228), .IN2(n4229), .IN3(n4230), .IN4(n4231), .QN(
        WX8444) );
  NAND2X0 U4591 ( .IN1(n3089), .IN2(n4008), .QN(n4231) );
  XNOR3X1 U4592 ( .IN1(n2757), .IN2(n2585), .IN3(n4232), .Q(n4008) );
  XOR2X1 U4593 ( .IN1(WX9802), .IN2(n6000), .Q(n4232) );
  NAND2X0 U4594 ( .IN1(n3005), .IN2(n4233), .QN(n4230) );
  NAND2X0 U4595 ( .IN1(WX8282), .IN2(n3030), .QN(n4229) );
  NAND2X0 U4596 ( .IN1(n3061), .IN2(CRC_OUT_3_10), .QN(n4228) );
  NAND4X0 U4597 ( .IN1(n4234), .IN2(n4235), .IN3(n4236), .IN4(n4237), .QN(
        WX8442) );
  NAND2X0 U4598 ( .IN1(n3090), .IN2(n4014), .QN(n4237) );
  XNOR3X1 U4599 ( .IN1(n2689), .IN2(n2586), .IN3(n4238), .Q(n4014) );
  XOR2X1 U4600 ( .IN1(WX9800), .IN2(n6001), .Q(n4238) );
  NAND2X0 U4601 ( .IN1(n4239), .IN2(n3018), .QN(n4236) );
  NAND2X0 U4602 ( .IN1(WX8280), .IN2(n3030), .QN(n4235) );
  NAND2X0 U4603 ( .IN1(n3061), .IN2(CRC_OUT_3_11), .QN(n4234) );
  NAND4X0 U4604 ( .IN1(n4240), .IN2(n4241), .IN3(n4242), .IN4(n4243), .QN(
        WX8440) );
  NAND2X0 U4605 ( .IN1(n3091), .IN2(n4020), .QN(n4243) );
  XNOR3X1 U4606 ( .IN1(n2756), .IN2(n2587), .IN3(n4244), .Q(n4020) );
  XOR2X1 U4607 ( .IN1(WX9798), .IN2(n6002), .Q(n4244) );
  NAND2X0 U4608 ( .IN1(n3005), .IN2(n4245), .QN(n4242) );
  NAND2X0 U4609 ( .IN1(WX8278), .IN2(n3030), .QN(n4241) );
  NAND2X0 U4610 ( .IN1(n3061), .IN2(CRC_OUT_3_12), .QN(n4240) );
  NAND4X0 U4611 ( .IN1(n4246), .IN2(n4247), .IN3(n4248), .IN4(n4249), .QN(
        WX8438) );
  NAND2X0 U4612 ( .IN1(n3090), .IN2(n4026), .QN(n4249) );
  XNOR3X1 U4613 ( .IN1(n2755), .IN2(n2588), .IN3(n4250), .Q(n4026) );
  XOR2X1 U4614 ( .IN1(WX9796), .IN2(n6003), .Q(n4250) );
  NAND2X0 U4615 ( .IN1(n4251), .IN2(n3018), .QN(n4248) );
  NAND2X0 U4616 ( .IN1(WX8276), .IN2(n3030), .QN(n4247) );
  NAND2X0 U4617 ( .IN1(n3062), .IN2(CRC_OUT_3_13), .QN(n4246) );
  NAND4X0 U4618 ( .IN1(n4252), .IN2(n4253), .IN3(n4254), .IN4(n4255), .QN(
        WX8436) );
  NAND2X0 U4619 ( .IN1(n4032), .IN2(n3099), .QN(n4255) );
  XOR3X1 U4620 ( .IN1(n3591), .IN2(n2589), .IN3(n4256), .Q(n4032) );
  XOR2X1 U4621 ( .IN1(WX9730), .IN2(test_so86), .Q(n4256) );
  NAND2X0 U4622 ( .IN1(n3005), .IN2(n4257), .QN(n4254) );
  NAND2X0 U4623 ( .IN1(WX8274), .IN2(n3030), .QN(n4253) );
  NAND2X0 U4624 ( .IN1(n3062), .IN2(CRC_OUT_3_14), .QN(n4252) );
  NAND4X0 U4625 ( .IN1(n4258), .IN2(n4259), .IN3(n4260), .IN4(n4261), .QN(
        WX8434) );
  NAND2X0 U4626 ( .IN1(n3090), .IN2(n4038), .QN(n4261) );
  XNOR3X1 U4627 ( .IN1(n2754), .IN2(n2590), .IN3(n4262), .Q(n4038) );
  XOR2X1 U4628 ( .IN1(WX9792), .IN2(n6004), .Q(n4262) );
  NAND2X0 U4629 ( .IN1(n4263), .IN2(n3017), .QN(n4260) );
  NAND2X0 U4630 ( .IN1(WX8272), .IN2(n3030), .QN(n4259) );
  NAND2X0 U4631 ( .IN1(n3062), .IN2(CRC_OUT_3_15), .QN(n4258) );
  NAND4X0 U4632 ( .IN1(n4264), .IN2(n4265), .IN3(n4266), .IN4(n4267), .QN(
        WX8432) );
  NAND2X0 U4633 ( .IN1(n4044), .IN2(n3099), .QN(n4267) );
  XOR3X1 U4634 ( .IN1(n2376), .IN2(n3579), .IN3(n4268), .Q(n4044) );
  XNOR3X1 U4635 ( .IN1(test_so84), .IN2(n6005), .IN3(n2688), .Q(n4268) );
  NAND2X0 U4636 ( .IN1(n3005), .IN2(n4269), .QN(n4266) );
  NAND2X0 U4637 ( .IN1(WX8270), .IN2(n3030), .QN(n4265) );
  NAND2X0 U4638 ( .IN1(n3062), .IN2(CRC_OUT_3_16), .QN(n4264) );
  NAND4X0 U4639 ( .IN1(n4270), .IN2(n4271), .IN3(n4272), .IN4(n4273), .QN(
        WX8430) );
  NAND2X0 U4640 ( .IN1(n3090), .IN2(n4050), .QN(n4273) );
  XNOR3X1 U4641 ( .IN1(n2377), .IN2(n3567), .IN3(n4274), .Q(n4050) );
  XOR3X1 U4642 ( .IN1(n6006), .IN2(n2753), .IN3(WX9852), .Q(n4274) );
  NAND2X0 U4643 ( .IN1(n3005), .IN2(n4275), .QN(n4272) );
  NAND2X0 U4644 ( .IN1(WX8268), .IN2(n3030), .QN(n4271) );
  NAND2X0 U4645 ( .IN1(n3062), .IN2(CRC_OUT_3_17), .QN(n4270) );
  NAND4X0 U4646 ( .IN1(n4276), .IN2(n4277), .IN3(n4278), .IN4(n4279), .QN(
        WX8428) );
  NAND2X0 U4647 ( .IN1(n4056), .IN2(n3099), .QN(n4279) );
  XOR3X1 U4648 ( .IN1(n2379), .IN2(n3579), .IN3(n4280), .Q(n4056) );
  XNOR3X1 U4649 ( .IN1(test_so82), .IN2(n6007), .IN3(n2752), .Q(n4280) );
  NAND2X0 U4650 ( .IN1(n3005), .IN2(n4281), .QN(n4278) );
  NAND2X0 U4651 ( .IN1(WX8266), .IN2(n3030), .QN(n4277) );
  NAND2X0 U4652 ( .IN1(n3062), .IN2(CRC_OUT_3_18), .QN(n4276) );
  NAND4X0 U4653 ( .IN1(n4282), .IN2(n4283), .IN3(n4284), .IN4(n4285), .QN(
        WX8426) );
  NAND2X0 U4654 ( .IN1(n3090), .IN2(n4062), .QN(n4285) );
  XNOR3X1 U4655 ( .IN1(n2380), .IN2(n3567), .IN3(n4286), .Q(n4062) );
  XOR3X1 U4656 ( .IN1(n6008), .IN2(n2751), .IN3(WX9848), .Q(n4286) );
  NAND2X0 U4657 ( .IN1(n3005), .IN2(n4287), .QN(n4284) );
  NAND2X0 U4658 ( .IN1(WX8264), .IN2(n3031), .QN(n4283) );
  NAND2X0 U4659 ( .IN1(n3062), .IN2(CRC_OUT_3_19), .QN(n4282) );
  NAND4X0 U4660 ( .IN1(n4288), .IN2(n4289), .IN3(n4290), .IN4(n4291), .QN(
        WX8424) );
  NAND2X0 U4661 ( .IN1(n4068), .IN2(n3099), .QN(n4291) );
  XOR3X1 U4662 ( .IN1(n2382), .IN2(n3579), .IN3(n4292), .Q(n4068) );
  XNOR3X1 U4663 ( .IN1(test_so80), .IN2(n6009), .IN3(n2750), .Q(n4292) );
  NAND2X0 U4664 ( .IN1(n3005), .IN2(n4293), .QN(n4290) );
  NAND2X0 U4665 ( .IN1(WX8262), .IN2(n3031), .QN(n4289) );
  NAND2X0 U4666 ( .IN1(n3062), .IN2(CRC_OUT_3_20), .QN(n4288) );
  NAND4X0 U4667 ( .IN1(n4294), .IN2(n4295), .IN3(n4296), .IN4(n4297), .QN(
        WX8422) );
  NAND2X0 U4668 ( .IN1(n3090), .IN2(n4074), .QN(n4297) );
  XNOR3X1 U4669 ( .IN1(n2383), .IN2(n3567), .IN3(n4298), .Q(n4074) );
  XOR3X1 U4670 ( .IN1(n6010), .IN2(n2749), .IN3(WX9844), .Q(n4298) );
  NAND2X0 U4671 ( .IN1(n3004), .IN2(n4299), .QN(n4296) );
  NAND2X0 U4672 ( .IN1(WX8260), .IN2(n3031), .QN(n4295) );
  NAND2X0 U4673 ( .IN1(n3062), .IN2(CRC_OUT_3_21), .QN(n4294) );
  NAND4X0 U4674 ( .IN1(n4300), .IN2(n4301), .IN3(n4302), .IN4(n4303), .QN(
        WX8420) );
  NAND2X0 U4675 ( .IN1(n3090), .IN2(n4080), .QN(n4303) );
  XNOR3X1 U4676 ( .IN1(n2385), .IN2(n3567), .IN3(n4304), .Q(n4080) );
  XOR3X1 U4677 ( .IN1(n6011), .IN2(n2748), .IN3(WX9842), .Q(n4304) );
  NAND2X0 U4678 ( .IN1(n3004), .IN2(n4305), .QN(n4302) );
  NAND2X0 U4679 ( .IN1(WX8258), .IN2(n3031), .QN(n4301) );
  NAND2X0 U4680 ( .IN1(n3062), .IN2(CRC_OUT_3_22), .QN(n4300) );
  NAND4X0 U4681 ( .IN1(n4306), .IN2(n4307), .IN3(n4308), .IN4(n4309), .QN(
        WX8418) );
  NAND2X0 U4682 ( .IN1(n3090), .IN2(n4086), .QN(n4309) );
  XNOR3X1 U4683 ( .IN1(n2387), .IN2(n3567), .IN3(n4310), .Q(n4086) );
  XOR3X1 U4684 ( .IN1(n6012), .IN2(n2747), .IN3(WX9840), .Q(n4310) );
  NAND2X0 U4685 ( .IN1(n3004), .IN2(n4311), .QN(n4308) );
  NAND2X0 U4686 ( .IN1(WX8256), .IN2(n3031), .QN(n4307) );
  NAND2X0 U4687 ( .IN1(n3062), .IN2(CRC_OUT_3_23), .QN(n4306) );
  NAND4X0 U4688 ( .IN1(n4312), .IN2(n4313), .IN3(n4314), .IN4(n4315), .QN(
        WX8416) );
  NAND2X0 U4689 ( .IN1(n3090), .IN2(n4092), .QN(n4315) );
  XNOR3X1 U4690 ( .IN1(n2389), .IN2(n3567), .IN3(n4316), .Q(n4092) );
  XOR3X1 U4691 ( .IN1(n6013), .IN2(n2746), .IN3(WX9838), .Q(n4316) );
  NAND2X0 U4692 ( .IN1(n3004), .IN2(n4317), .QN(n4314) );
  NAND2X0 U4693 ( .IN1(WX8254), .IN2(n3031), .QN(n4313) );
  NAND2X0 U4694 ( .IN1(test_so77), .IN2(n3069), .QN(n4312) );
  NAND4X0 U4695 ( .IN1(n4318), .IN2(n4319), .IN3(n4320), .IN4(n4321), .QN(
        WX8414) );
  NAND2X0 U4696 ( .IN1(n3090), .IN2(n4098), .QN(n4321) );
  XNOR3X1 U4697 ( .IN1(n2391), .IN2(n3567), .IN3(n4322), .Q(n4098) );
  XOR3X1 U4698 ( .IN1(n6014), .IN2(n2745), .IN3(WX9836), .Q(n4322) );
  NAND2X0 U4699 ( .IN1(n3004), .IN2(n4323), .QN(n4320) );
  NAND2X0 U4700 ( .IN1(WX8252), .IN2(n3031), .QN(n4319) );
  NAND2X0 U4701 ( .IN1(n3062), .IN2(CRC_OUT_3_25), .QN(n4318) );
  NAND4X0 U4702 ( .IN1(n4324), .IN2(n4325), .IN3(n4326), .IN4(n4327), .QN(
        WX8412) );
  NAND2X0 U4703 ( .IN1(n3090), .IN2(n4104), .QN(n4327) );
  XNOR3X1 U4704 ( .IN1(n2393), .IN2(n3567), .IN3(n4328), .Q(n4104) );
  XOR3X1 U4705 ( .IN1(n6015), .IN2(n2744), .IN3(WX9834), .Q(n4328) );
  NAND2X0 U4706 ( .IN1(n4329), .IN2(n3017), .QN(n4326) );
  NAND2X0 U4707 ( .IN1(WX8250), .IN2(n3031), .QN(n4325) );
  NAND2X0 U4708 ( .IN1(n3063), .IN2(CRC_OUT_3_26), .QN(n4324) );
  NAND4X0 U4709 ( .IN1(n4330), .IN2(n4331), .IN3(n4332), .IN4(n4333), .QN(
        WX8410) );
  NAND2X0 U4710 ( .IN1(n3091), .IN2(n4110), .QN(n4333) );
  XNOR3X1 U4711 ( .IN1(n2395), .IN2(n3567), .IN3(n4334), .Q(n4110) );
  XOR3X1 U4712 ( .IN1(n6016), .IN2(n2743), .IN3(WX9832), .Q(n4334) );
  NAND2X0 U4713 ( .IN1(n3004), .IN2(n4335), .QN(n4332) );
  NAND2X0 U4714 ( .IN1(WX8248), .IN2(n3031), .QN(n4331) );
  NAND2X0 U4715 ( .IN1(n3063), .IN2(CRC_OUT_3_27), .QN(n4330) );
  NAND4X0 U4716 ( .IN1(n4336), .IN2(n4337), .IN3(n4338), .IN4(n4339), .QN(
        WX8408) );
  NAND2X0 U4717 ( .IN1(n3091), .IN2(n4116), .QN(n4339) );
  XNOR3X1 U4718 ( .IN1(n2397), .IN2(n3567), .IN3(n4340), .Q(n4116) );
  XOR3X1 U4719 ( .IN1(n6017), .IN2(n2742), .IN3(WX9830), .Q(n4340) );
  NAND2X0 U4720 ( .IN1(n4341), .IN2(n3017), .QN(n4338) );
  NAND2X0 U4721 ( .IN1(WX8246), .IN2(n3031), .QN(n4337) );
  NAND2X0 U4722 ( .IN1(n3063), .IN2(CRC_OUT_3_28), .QN(n4336) );
  NAND4X0 U4723 ( .IN1(n4342), .IN2(n4343), .IN3(n4344), .IN4(n4345), .QN(
        WX8406) );
  NAND2X0 U4724 ( .IN1(n3091), .IN2(n4122), .QN(n4345) );
  XNOR3X1 U4725 ( .IN1(n2399), .IN2(n3567), .IN3(n4346), .Q(n4122) );
  XOR3X1 U4726 ( .IN1(n6018), .IN2(n2741), .IN3(WX9828), .Q(n4346) );
  NAND2X0 U4727 ( .IN1(n3004), .IN2(n4347), .QN(n4344) );
  NAND2X0 U4728 ( .IN1(WX8244), .IN2(n3031), .QN(n4343) );
  NAND2X0 U4729 ( .IN1(n3063), .IN2(CRC_OUT_3_29), .QN(n4342) );
  NAND4X0 U4730 ( .IN1(n4348), .IN2(n4349), .IN3(n4350), .IN4(n4351), .QN(
        WX8404) );
  NAND2X0 U4731 ( .IN1(n3091), .IN2(n4128), .QN(n4351) );
  XNOR3X1 U4732 ( .IN1(n2401), .IN2(n3567), .IN3(n4352), .Q(n4128) );
  XOR3X1 U4733 ( .IN1(n6019), .IN2(n2740), .IN3(WX9826), .Q(n4352) );
  NAND2X0 U4734 ( .IN1(n4353), .IN2(n3017), .QN(n4350) );
  NAND2X0 U4735 ( .IN1(WX8242), .IN2(n3031), .QN(n4349) );
  NAND2X0 U4736 ( .IN1(n3063), .IN2(CRC_OUT_3_30), .QN(n4348) );
  NAND4X0 U4737 ( .IN1(n4354), .IN2(n4355), .IN3(n4356), .IN4(n4357), .QN(
        WX8402) );
  NAND2X0 U4738 ( .IN1(n4134), .IN2(n3100), .QN(n4357) );
  XOR3X1 U4739 ( .IN1(n2337), .IN2(n3578), .IN3(n4358), .Q(n4134) );
  XOR3X1 U4740 ( .IN1(test_so85), .IN2(n6020), .IN3(WX9824), .Q(n4358) );
  NAND2X0 U4741 ( .IN1(n3004), .IN2(n4359), .QN(n4356) );
  NAND2X0 U4742 ( .IN1(n3063), .IN2(CRC_OUT_3_31), .QN(n4355) );
  NAND2X0 U4743 ( .IN1(n2245), .IN2(WX8243), .QN(n4354) );
  NOR2X0 U4744 ( .IN1(n3747), .IN2(WX8243), .QN(WX8304) );
  AND2X1 U4745 ( .IN1(test_so68), .IN2(n3598), .Q(WX8302) );
  AND2X1 U4746 ( .IN1(n3627), .IN2(n8381), .Q(WX8300) );
  AND2X1 U4747 ( .IN1(n3627), .IN2(n8382), .Q(WX8298) );
  AND2X1 U4748 ( .IN1(n3627), .IN2(n8383), .Q(WX8296) );
  AND2X1 U4749 ( .IN1(n3627), .IN2(n8384), .Q(WX8294) );
  AND2X1 U4750 ( .IN1(n3627), .IN2(n8385), .Q(WX8292) );
  AND2X1 U4751 ( .IN1(n3627), .IN2(n8386), .Q(WX8290) );
  AND2X1 U4752 ( .IN1(n3627), .IN2(n8387), .Q(WX8288) );
  AND2X1 U4753 ( .IN1(n3626), .IN2(n8388), .Q(WX8286) );
  AND2X1 U4754 ( .IN1(n3626), .IN2(n8389), .Q(WX8284) );
  AND2X1 U4755 ( .IN1(n3626), .IN2(n8390), .Q(WX8282) );
  AND2X1 U4756 ( .IN1(n3626), .IN2(n8391), .Q(WX8280) );
  AND2X1 U4757 ( .IN1(n3626), .IN2(n8392), .Q(WX8278) );
  AND2X1 U4758 ( .IN1(n3626), .IN2(n8393), .Q(WX8276) );
  AND2X1 U4759 ( .IN1(n3626), .IN2(n8394), .Q(WX8274) );
  AND2X1 U4760 ( .IN1(n3626), .IN2(n8395), .Q(WX8272) );
  AND2X1 U4761 ( .IN1(n3626), .IN2(n8396), .Q(WX8270) );
  AND2X1 U4762 ( .IN1(test_so67), .IN2(n3598), .Q(WX8268) );
  AND2X1 U4763 ( .IN1(n3624), .IN2(n8399), .Q(WX8266) );
  AND2X1 U4764 ( .IN1(n3624), .IN2(n8400), .Q(WX8264) );
  AND2X1 U4765 ( .IN1(n3624), .IN2(n8401), .Q(WX8262) );
  AND2X1 U4766 ( .IN1(n3624), .IN2(n8402), .Q(WX8260) );
  AND2X1 U4767 ( .IN1(n3624), .IN2(n8403), .Q(WX8258) );
  AND2X1 U4768 ( .IN1(n3624), .IN2(n8404), .Q(WX8256) );
  AND2X1 U4769 ( .IN1(n3624), .IN2(n8405), .Q(WX8254) );
  AND2X1 U4770 ( .IN1(n3624), .IN2(n8406), .Q(WX8252) );
  AND2X1 U4771 ( .IN1(n3623), .IN2(n8407), .Q(WX8250) );
  AND2X1 U4772 ( .IN1(n3623), .IN2(n8408), .Q(WX8248) );
  AND2X1 U4773 ( .IN1(n3623), .IN2(n8409), .Q(WX8246) );
  AND2X1 U4774 ( .IN1(n3623), .IN2(n8410), .Q(WX8244) );
  AND2X1 U4775 ( .IN1(n3623), .IN2(n8411), .Q(WX8242) );
  NOR2X0 U4776 ( .IN1(n3747), .IN2(n4360), .QN(WX7791) );
  XOR2X1 U4777 ( .IN1(n2792), .IN2(DFF_1150_n1), .Q(n4360) );
  NOR2X0 U4778 ( .IN1(n3747), .IN2(n4361), .QN(WX7789) );
  XNOR2X1 U4779 ( .IN1(n2793), .IN2(test_so66), .Q(n4361) );
  NOR2X0 U4780 ( .IN1(n3747), .IN2(n4362), .QN(WX7787) );
  XOR2X1 U4781 ( .IN1(n2794), .IN2(DFF_1148_n1), .Q(n4362) );
  NOR2X0 U4782 ( .IN1(n3747), .IN2(n4363), .QN(WX7785) );
  XOR2X1 U4783 ( .IN1(n2795), .IN2(DFF_1147_n1), .Q(n4363) );
  NOR2X0 U4784 ( .IN1(n3747), .IN2(n4364), .QN(WX7783) );
  XOR2X1 U4785 ( .IN1(n2796), .IN2(DFF_1146_n1), .Q(n4364) );
  NOR2X0 U4786 ( .IN1(n3748), .IN2(n4365), .QN(WX7781) );
  XOR2X1 U4787 ( .IN1(n2797), .IN2(DFF_1145_n1), .Q(n4365) );
  NOR2X0 U4788 ( .IN1(n3748), .IN2(n4366), .QN(WX7779) );
  XOR2X1 U4789 ( .IN1(n2798), .IN2(DFF_1144_n1), .Q(n4366) );
  NOR2X0 U4790 ( .IN1(n3748), .IN2(n4367), .QN(WX7777) );
  XOR2X1 U4791 ( .IN1(n2799), .IN2(DFF_1143_n1), .Q(n4367) );
  NOR2X0 U4792 ( .IN1(n3748), .IN2(n4368), .QN(WX7775) );
  XOR2X1 U4793 ( .IN1(n2800), .IN2(DFF_1142_n1), .Q(n4368) );
  NOR2X0 U4794 ( .IN1(n3748), .IN2(n4369), .QN(WX7773) );
  XOR2X1 U4795 ( .IN1(n2801), .IN2(DFF_1141_n1), .Q(n4369) );
  NOR2X0 U4796 ( .IN1(n3748), .IN2(n4370), .QN(WX7771) );
  XOR2X1 U4797 ( .IN1(CRC_OUT_4_20), .IN2(test_so63), .Q(n4370) );
  NOR2X0 U4798 ( .IN1(n3748), .IN2(n4371), .QN(WX7769) );
  XOR2X1 U4799 ( .IN1(n2802), .IN2(DFF_1139_n1), .Q(n4371) );
  NOR2X0 U4800 ( .IN1(n3748), .IN2(n4372), .QN(WX7767) );
  XOR2X1 U4801 ( .IN1(n2803), .IN2(DFF_1138_n1), .Q(n4372) );
  NOR2X0 U4802 ( .IN1(n3748), .IN2(n4373), .QN(WX7765) );
  XOR2X1 U4803 ( .IN1(n2804), .IN2(DFF_1137_n1), .Q(n4373) );
  NOR2X0 U4804 ( .IN1(n3748), .IN2(n4374), .QN(WX7763) );
  XOR2X1 U4805 ( .IN1(n2805), .IN2(DFF_1136_n1), .Q(n4374) );
  NOR2X0 U4806 ( .IN1(n3748), .IN2(n4375), .QN(WX7761) );
  XOR3X1 U4807 ( .IN1(n2694), .IN2(DFF_1151_n1), .IN3(CRC_OUT_4_15), .Q(n4375)
         );
  NOR2X0 U4808 ( .IN1(n3748), .IN2(n4376), .QN(WX7759) );
  XOR2X1 U4809 ( .IN1(n2806), .IN2(DFF_1134_n1), .Q(n4376) );
  NOR2X0 U4810 ( .IN1(n3748), .IN2(n4377), .QN(WX7757) );
  XOR2X1 U4811 ( .IN1(n2807), .IN2(DFF_1133_n1), .Q(n4377) );
  NOR2X0 U4812 ( .IN1(n3749), .IN2(n4378), .QN(WX7755) );
  XNOR2X1 U4813 ( .IN1(n2808), .IN2(test_so65), .Q(n4378) );
  NOR2X0 U4814 ( .IN1(n3749), .IN2(n4379), .QN(WX7753) );
  XOR2X1 U4815 ( .IN1(n2809), .IN2(DFF_1131_n1), .Q(n4379) );
  NOR2X0 U4816 ( .IN1(n3749), .IN2(n4380), .QN(WX7751) );
  XOR3X1 U4817 ( .IN1(n2695), .IN2(DFF_1151_n1), .IN3(CRC_OUT_4_10), .Q(n4380)
         );
  NOR2X0 U4818 ( .IN1(n3749), .IN2(n4381), .QN(WX7749) );
  XOR2X1 U4819 ( .IN1(n2810), .IN2(DFF_1129_n1), .Q(n4381) );
  NOR2X0 U4820 ( .IN1(n3749), .IN2(n4382), .QN(WX7747) );
  XOR2X1 U4821 ( .IN1(n2811), .IN2(DFF_1128_n1), .Q(n4382) );
  NOR2X0 U4822 ( .IN1(n3749), .IN2(n4383), .QN(WX7745) );
  XOR2X1 U4823 ( .IN1(n2812), .IN2(DFF_1127_n1), .Q(n4383) );
  NOR2X0 U4824 ( .IN1(n3749), .IN2(n4384), .QN(WX7743) );
  XOR2X1 U4825 ( .IN1(n2813), .IN2(DFF_1126_n1), .Q(n4384) );
  NOR2X0 U4826 ( .IN1(n3749), .IN2(n4385), .QN(WX7741) );
  XOR2X1 U4827 ( .IN1(n2814), .IN2(DFF_1125_n1), .Q(n4385) );
  NOR2X0 U4828 ( .IN1(n3749), .IN2(n4386), .QN(WX7739) );
  XOR2X1 U4829 ( .IN1(n2815), .IN2(DFF_1124_n1), .Q(n4386) );
  NOR2X0 U4830 ( .IN1(n3749), .IN2(n4387), .QN(WX7737) );
  XOR3X1 U4831 ( .IN1(test_so64), .IN2(DFF_1151_n1), .IN3(DFF_1123_n1), .Q(
        n4387) );
  NOR2X0 U4832 ( .IN1(n3749), .IN2(n4388), .QN(WX7735) );
  XOR2X1 U4833 ( .IN1(n2816), .IN2(DFF_1122_n1), .Q(n4388) );
  NOR2X0 U4834 ( .IN1(n3749), .IN2(n4389), .QN(WX7733) );
  XOR2X1 U4835 ( .IN1(n2817), .IN2(DFF_1121_n1), .Q(n4389) );
  NOR2X0 U4836 ( .IN1(n3749), .IN2(n4390), .QN(WX7731) );
  XOR2X1 U4837 ( .IN1(n2818), .IN2(DFF_1120_n1), .Q(n4390) );
  NOR2X0 U4838 ( .IN1(n3750), .IN2(n4391), .QN(WX7729) );
  XOR2X1 U4839 ( .IN1(n2709), .IN2(DFF_1151_n1), .Q(n4391) );
  NOR2X0 U4840 ( .IN1(n6061), .IN2(n3654), .QN(WX7203) );
  NOR2X0 U4841 ( .IN1(n6062), .IN2(n3654), .QN(WX7201) );
  NOR2X0 U4842 ( .IN1(n6063), .IN2(n3654), .QN(WX7199) );
  NOR2X0 U4843 ( .IN1(n6064), .IN2(n3654), .QN(WX7197) );
  NOR2X0 U4844 ( .IN1(n6065), .IN2(n3655), .QN(WX7195) );
  NOR2X0 U4845 ( .IN1(n6066), .IN2(n3655), .QN(WX7193) );
  NOR2X0 U4846 ( .IN1(n6067), .IN2(n3655), .QN(WX7191) );
  NOR2X0 U4847 ( .IN1(n6068), .IN2(n3655), .QN(WX7189) );
  NOR2X0 U4848 ( .IN1(n6069), .IN2(n3655), .QN(WX7187) );
  NOR2X0 U4849 ( .IN1(n6070), .IN2(n3655), .QN(WX7185) );
  NOR2X0 U4850 ( .IN1(n6071), .IN2(n3655), .QN(WX7183) );
  AND2X1 U4851 ( .IN1(n3623), .IN2(test_so57), .Q(WX7181) );
  NOR2X0 U4852 ( .IN1(n6073), .IN2(n3655), .QN(WX7179) );
  NOR2X0 U4853 ( .IN1(n6074), .IN2(n3655), .QN(WX7177) );
  NOR2X0 U4854 ( .IN1(n6075), .IN2(n3655), .QN(WX7175) );
  NOR2X0 U4855 ( .IN1(n6076), .IN2(n3655), .QN(WX7173) );
  NAND4X0 U4856 ( .IN1(n4392), .IN2(n4393), .IN3(n4394), .IN4(n4395), .QN(
        WX7171) );
  NAND2X0 U4857 ( .IN1(n3091), .IN2(n4173), .QN(n4395) );
  XNOR3X1 U4858 ( .IN1(n2708), .IN2(n2591), .IN3(n4396), .Q(n4173) );
  XOR2X1 U4859 ( .IN1(WX8529), .IN2(n6021), .Q(n4396) );
  NAND2X0 U4860 ( .IN1(n3004), .IN2(n4397), .QN(n4394) );
  NAND2X0 U4861 ( .IN1(WX7009), .IN2(n3031), .QN(n4393) );
  NAND2X0 U4862 ( .IN1(n3063), .IN2(CRC_OUT_4_0), .QN(n4392) );
  NAND4X0 U4863 ( .IN1(n4398), .IN2(n4399), .IN3(n4400), .IN4(n4401), .QN(
        WX7169) );
  NAND2X0 U4864 ( .IN1(n3091), .IN2(n4179), .QN(n4401) );
  XNOR3X1 U4865 ( .IN1(n2791), .IN2(n2592), .IN3(n4402), .Q(n4179) );
  XOR2X1 U4866 ( .IN1(WX8527), .IN2(n6022), .Q(n4402) );
  NAND2X0 U4867 ( .IN1(n3004), .IN2(n4403), .QN(n4400) );
  NAND2X0 U4868 ( .IN1(WX7007), .IN2(n3031), .QN(n4399) );
  NAND2X0 U4869 ( .IN1(n3063), .IN2(CRC_OUT_4_1), .QN(n4398) );
  NAND4X0 U4870 ( .IN1(n4404), .IN2(n4405), .IN3(n4406), .IN4(n4407), .QN(
        WX7167) );
  NAND2X0 U4871 ( .IN1(n3091), .IN2(n4185), .QN(n4407) );
  XNOR3X1 U4872 ( .IN1(n2790), .IN2(n2593), .IN3(n4408), .Q(n4185) );
  XOR2X1 U4873 ( .IN1(WX8525), .IN2(n6023), .Q(n4408) );
  NAND2X0 U4874 ( .IN1(n3004), .IN2(n4409), .QN(n4406) );
  NAND2X0 U4875 ( .IN1(WX7005), .IN2(n3031), .QN(n4405) );
  NAND2X0 U4876 ( .IN1(n3063), .IN2(CRC_OUT_4_2), .QN(n4404) );
  NAND4X0 U4877 ( .IN1(n4410), .IN2(n4411), .IN3(n4412), .IN4(n4413), .QN(
        WX7165) );
  NAND2X0 U4878 ( .IN1(n3091), .IN2(n4191), .QN(n4413) );
  XNOR3X1 U4879 ( .IN1(n2789), .IN2(n2594), .IN3(n4414), .Q(n4191) );
  XOR2X1 U4880 ( .IN1(WX8523), .IN2(n6024), .Q(n4414) );
  NAND2X0 U4881 ( .IN1(n3004), .IN2(n4415), .QN(n4412) );
  NAND2X0 U4882 ( .IN1(WX7003), .IN2(n3031), .QN(n4411) );
  NAND2X0 U4883 ( .IN1(n3063), .IN2(CRC_OUT_4_3), .QN(n4410) );
  NAND4X0 U4884 ( .IN1(n4416), .IN2(n4417), .IN3(n4418), .IN4(n4419), .QN(
        WX7163) );
  NAND2X0 U4885 ( .IN1(n3091), .IN2(n4197), .QN(n4419) );
  XNOR3X1 U4886 ( .IN1(n2693), .IN2(n2595), .IN3(n4420), .Q(n4197) );
  XOR2X1 U4887 ( .IN1(WX8521), .IN2(n6025), .Q(n4420) );
  NAND2X0 U4888 ( .IN1(n4421), .IN2(n3017), .QN(n4418) );
  NAND2X0 U4889 ( .IN1(WX7001), .IN2(n3031), .QN(n4417) );
  NAND2X0 U4890 ( .IN1(n3063), .IN2(CRC_OUT_4_4), .QN(n4416) );
  NAND4X0 U4891 ( .IN1(n4422), .IN2(n4423), .IN3(n4424), .IN4(n4425), .QN(
        WX7161) );
  NAND2X0 U4892 ( .IN1(n3091), .IN2(n4203), .QN(n4425) );
  XNOR3X1 U4893 ( .IN1(n2788), .IN2(n2596), .IN3(n4426), .Q(n4203) );
  XOR2X1 U4894 ( .IN1(WX8519), .IN2(n6026), .Q(n4426) );
  NAND2X0 U4895 ( .IN1(n3003), .IN2(n4427), .QN(n4424) );
  NAND2X0 U4896 ( .IN1(WX6999), .IN2(n3032), .QN(n4423) );
  NAND2X0 U4897 ( .IN1(n3063), .IN2(CRC_OUT_4_5), .QN(n4422) );
  NAND4X0 U4898 ( .IN1(n4428), .IN2(n4429), .IN3(n4430), .IN4(n4431), .QN(
        WX7159) );
  NAND2X0 U4899 ( .IN1(n3091), .IN2(n4209), .QN(n4431) );
  XNOR3X1 U4900 ( .IN1(n2787), .IN2(n2597), .IN3(n4432), .Q(n4209) );
  XOR2X1 U4901 ( .IN1(WX8517), .IN2(n6027), .Q(n4432) );
  NAND2X0 U4902 ( .IN1(n4433), .IN2(n3017), .QN(n4430) );
  NAND2X0 U4903 ( .IN1(WX6997), .IN2(n3032), .QN(n4429) );
  NAND2X0 U4904 ( .IN1(n3064), .IN2(CRC_OUT_4_6), .QN(n4428) );
  NAND4X0 U4905 ( .IN1(n4434), .IN2(n4435), .IN3(n4436), .IN4(n4437), .QN(
        WX7157) );
  NAND2X0 U4906 ( .IN1(n3092), .IN2(n4215), .QN(n4437) );
  XNOR3X1 U4907 ( .IN1(n2786), .IN2(n2598), .IN3(n4438), .Q(n4215) );
  XOR2X1 U4908 ( .IN1(WX8515), .IN2(n6028), .Q(n4438) );
  NAND2X0 U4909 ( .IN1(n3003), .IN2(n4439), .QN(n4436) );
  NAND2X0 U4910 ( .IN1(WX6995), .IN2(n3032), .QN(n4435) );
  NAND2X0 U4911 ( .IN1(n3064), .IN2(CRC_OUT_4_7), .QN(n4434) );
  NAND4X0 U4912 ( .IN1(n4440), .IN2(n4441), .IN3(n4442), .IN4(n4443), .QN(
        WX7155) );
  NAND2X0 U4913 ( .IN1(n3092), .IN2(n4221), .QN(n4443) );
  XNOR3X1 U4914 ( .IN1(n2785), .IN2(n2599), .IN3(n4444), .Q(n4221) );
  XOR2X1 U4915 ( .IN1(WX8513), .IN2(n6029), .Q(n4444) );
  NAND2X0 U4916 ( .IN1(n4445), .IN2(n3017), .QN(n4442) );
  NAND2X0 U4917 ( .IN1(WX6993), .IN2(n3032), .QN(n4441) );
  NAND2X0 U4918 ( .IN1(n3064), .IN2(CRC_OUT_4_8), .QN(n4440) );
  NAND4X0 U4919 ( .IN1(n4446), .IN2(n4447), .IN3(n4448), .IN4(n4449), .QN(
        WX7153) );
  NAND2X0 U4920 ( .IN1(n4227), .IN2(n3100), .QN(n4449) );
  XOR3X1 U4921 ( .IN1(n3613), .IN2(n2600), .IN3(n4450), .Q(n4227) );
  XOR2X1 U4922 ( .IN1(WX8447), .IN2(test_so75), .Q(n4450) );
  NAND2X0 U4923 ( .IN1(n3003), .IN2(n4451), .QN(n4448) );
  NAND2X0 U4924 ( .IN1(WX6991), .IN2(n3032), .QN(n4447) );
  NAND2X0 U4925 ( .IN1(n3064), .IN2(CRC_OUT_4_9), .QN(n4446) );
  NAND4X0 U4926 ( .IN1(n4452), .IN2(n4453), .IN3(n4454), .IN4(n4455), .QN(
        WX7151) );
  NAND2X0 U4927 ( .IN1(n3092), .IN2(n4233), .QN(n4455) );
  XNOR3X1 U4928 ( .IN1(n2784), .IN2(n2601), .IN3(n4456), .Q(n4233) );
  XOR2X1 U4929 ( .IN1(WX8509), .IN2(n6030), .Q(n4456) );
  NAND2X0 U4930 ( .IN1(n4457), .IN2(n3016), .QN(n4454) );
  NAND2X0 U4931 ( .IN1(WX6989), .IN2(n3032), .QN(n4453) );
  NAND2X0 U4932 ( .IN1(n3064), .IN2(CRC_OUT_4_10), .QN(n4452) );
  NAND4X0 U4933 ( .IN1(n4458), .IN2(n4459), .IN3(n4460), .IN4(n4461), .QN(
        WX7149) );
  NAND2X0 U4934 ( .IN1(n4239), .IN2(n3100), .QN(n4461) );
  XOR3X1 U4935 ( .IN1(n3617), .IN2(n2692), .IN3(n4462), .Q(n4239) );
  XOR2X1 U4936 ( .IN1(WX8443), .IN2(test_so73), .Q(n4462) );
  NAND2X0 U4937 ( .IN1(n3003), .IN2(n4463), .QN(n4460) );
  NAND2X0 U4938 ( .IN1(WX6987), .IN2(n3032), .QN(n4459) );
  NAND2X0 U4939 ( .IN1(n3064), .IN2(CRC_OUT_4_11), .QN(n4458) );
  NAND4X0 U4940 ( .IN1(n4464), .IN2(n4465), .IN3(n4466), .IN4(n4467), .QN(
        WX7147) );
  NAND2X0 U4941 ( .IN1(n3092), .IN2(n4245), .QN(n4467) );
  XNOR3X1 U4942 ( .IN1(n2783), .IN2(n2602), .IN3(n4468), .Q(n4245) );
  XOR2X1 U4943 ( .IN1(WX8505), .IN2(n6031), .Q(n4468) );
  NAND2X0 U4944 ( .IN1(n3003), .IN2(n4469), .QN(n4466) );
  NAND2X0 U4945 ( .IN1(WX6985), .IN2(n3032), .QN(n4465) );
  NAND2X0 U4946 ( .IN1(test_so65), .IN2(n3069), .QN(n4464) );
  NAND4X0 U4947 ( .IN1(n4470), .IN2(n4471), .IN3(n4472), .IN4(n4473), .QN(
        WX7145) );
  NAND2X0 U4948 ( .IN1(n4251), .IN2(n3100), .QN(n4473) );
  XOR3X1 U4949 ( .IN1(n2782), .IN2(n2603), .IN3(n4474), .Q(n4251) );
  XOR2X1 U4950 ( .IN1(WX8439), .IN2(test_so71), .Q(n4474) );
  NAND2X0 U4951 ( .IN1(n3003), .IN2(n4475), .QN(n4472) );
  NAND2X0 U4952 ( .IN1(WX6983), .IN2(n3032), .QN(n4471) );
  NAND2X0 U4953 ( .IN1(n3064), .IN2(CRC_OUT_4_13), .QN(n4470) );
  NAND4X0 U4954 ( .IN1(n4476), .IN2(n4477), .IN3(n4478), .IN4(n4479), .QN(
        WX7143) );
  NAND2X0 U4955 ( .IN1(n3092), .IN2(n4257), .QN(n4479) );
  XNOR3X1 U4956 ( .IN1(n2781), .IN2(n2604), .IN3(n4480), .Q(n4257) );
  XOR2X1 U4957 ( .IN1(WX8501), .IN2(n6032), .Q(n4480) );
  NAND2X0 U4958 ( .IN1(n3003), .IN2(n4481), .QN(n4478) );
  NAND2X0 U4959 ( .IN1(WX6981), .IN2(n3032), .QN(n4477) );
  NAND2X0 U4960 ( .IN1(n3064), .IN2(CRC_OUT_4_14), .QN(n4476) );
  NAND4X0 U4961 ( .IN1(n4482), .IN2(n4483), .IN3(n4484), .IN4(n4485), .QN(
        WX7141) );
  NAND2X0 U4962 ( .IN1(n4263), .IN2(n3100), .QN(n4485) );
  XOR3X1 U4963 ( .IN1(n3625), .IN2(n2780), .IN3(n4486), .Q(n4263) );
  XOR2X1 U4964 ( .IN1(WX8563), .IN2(test_so69), .Q(n4486) );
  NAND2X0 U4965 ( .IN1(n3003), .IN2(n4487), .QN(n4484) );
  NAND2X0 U4966 ( .IN1(WX6979), .IN2(n3032), .QN(n4483) );
  NAND2X0 U4967 ( .IN1(n3064), .IN2(CRC_OUT_4_15), .QN(n4482) );
  NAND4X0 U4968 ( .IN1(n4488), .IN2(n4489), .IN3(n4490), .IN4(n4491), .QN(
        WX7139) );
  NAND2X0 U4969 ( .IN1(n3092), .IN2(n4269), .QN(n4491) );
  XNOR3X1 U4970 ( .IN1(n2403), .IN2(n3568), .IN3(n4492), .Q(n4269) );
  XOR3X1 U4971 ( .IN1(n6033), .IN2(n2691), .IN3(WX8561), .Q(n4492) );
  NAND2X0 U4972 ( .IN1(n3003), .IN2(n4493), .QN(n4490) );
  NAND2X0 U4973 ( .IN1(WX6977), .IN2(n3032), .QN(n4489) );
  NAND2X0 U4974 ( .IN1(n3065), .IN2(CRC_OUT_4_16), .QN(n4488) );
  NAND4X0 U4975 ( .IN1(n4494), .IN2(n4495), .IN3(n4496), .IN4(n4497), .QN(
        WX7137) );
  NAND2X0 U4976 ( .IN1(n3093), .IN2(n4275), .QN(n4497) );
  XNOR3X1 U4977 ( .IN1(n2405), .IN2(n3568), .IN3(n4498), .Q(n4275) );
  XOR3X1 U4978 ( .IN1(n6034), .IN2(n2779), .IN3(WX8559), .Q(n4498) );
  NAND2X0 U4979 ( .IN1(n3003), .IN2(n4499), .QN(n4496) );
  NAND2X0 U4980 ( .IN1(WX6975), .IN2(n3032), .QN(n4495) );
  NAND2X0 U4981 ( .IN1(n3065), .IN2(CRC_OUT_4_17), .QN(n4494) );
  NAND4X0 U4982 ( .IN1(n4500), .IN2(n4501), .IN3(n4502), .IN4(n4503), .QN(
        WX7135) );
  NAND2X0 U4983 ( .IN1(n3092), .IN2(n4281), .QN(n4503) );
  XNOR3X1 U4984 ( .IN1(n2407), .IN2(n3568), .IN3(n4504), .Q(n4281) );
  XOR3X1 U4985 ( .IN1(n6035), .IN2(n2778), .IN3(WX8557), .Q(n4504) );
  NAND2X0 U4986 ( .IN1(n3003), .IN2(n4505), .QN(n4502) );
  NAND2X0 U4987 ( .IN1(WX6973), .IN2(n3032), .QN(n4501) );
  NAND2X0 U4988 ( .IN1(n3065), .IN2(CRC_OUT_4_18), .QN(n4500) );
  NAND4X0 U4989 ( .IN1(n4506), .IN2(n4507), .IN3(n4508), .IN4(n4509), .QN(
        WX7133) );
  NAND2X0 U4990 ( .IN1(n3093), .IN2(n4287), .QN(n4509) );
  XNOR3X1 U4991 ( .IN1(n2409), .IN2(n3568), .IN3(n4510), .Q(n4287) );
  XOR3X1 U4992 ( .IN1(n6036), .IN2(n2777), .IN3(WX8555), .Q(n4510) );
  NAND2X0 U4993 ( .IN1(n3002), .IN2(n4511), .QN(n4508) );
  NAND2X0 U4994 ( .IN1(WX6971), .IN2(n3032), .QN(n4507) );
  NAND2X0 U4995 ( .IN1(n3064), .IN2(CRC_OUT_4_19), .QN(n4506) );
  NAND4X0 U4996 ( .IN1(n4512), .IN2(n4513), .IN3(n4514), .IN4(n4515), .QN(
        WX7131) );
  NAND2X0 U4997 ( .IN1(n3093), .IN2(n4293), .QN(n4515) );
  XNOR3X1 U4998 ( .IN1(n2411), .IN2(n3568), .IN3(n4516), .Q(n4293) );
  XOR3X1 U4999 ( .IN1(n6037), .IN2(n2776), .IN3(WX8553), .Q(n4516) );
  NAND2X0 U5000 ( .IN1(n3002), .IN2(n4517), .QN(n4514) );
  NAND2X0 U5001 ( .IN1(WX6969), .IN2(n3032), .QN(n4513) );
  NAND2X0 U5002 ( .IN1(n3065), .IN2(CRC_OUT_4_20), .QN(n4512) );
  NAND4X0 U5003 ( .IN1(n4518), .IN2(n4519), .IN3(n4520), .IN4(n4521), .QN(
        WX7129) );
  NAND2X0 U5004 ( .IN1(n3092), .IN2(n4299), .QN(n4521) );
  XNOR3X1 U5005 ( .IN1(n2413), .IN2(n3568), .IN3(n4522), .Q(n4299) );
  XOR3X1 U5006 ( .IN1(n6038), .IN2(n2775), .IN3(WX8551), .Q(n4522) );
  NAND2X0 U5007 ( .IN1(n4523), .IN2(n3018), .QN(n4520) );
  NAND2X0 U5008 ( .IN1(WX6967), .IN2(n3032), .QN(n4519) );
  NAND2X0 U5009 ( .IN1(n3065), .IN2(CRC_OUT_4_21), .QN(n4518) );
  NAND4X0 U5010 ( .IN1(n4524), .IN2(n4525), .IN3(n4526), .IN4(n4527), .QN(
        WX7127) );
  NAND2X0 U5011 ( .IN1(n3093), .IN2(n4305), .QN(n4527) );
  XNOR3X1 U5012 ( .IN1(n2415), .IN2(n3568), .IN3(n4528), .Q(n4305) );
  XOR3X1 U5013 ( .IN1(n6039), .IN2(n2774), .IN3(WX8549), .Q(n4528) );
  NAND2X0 U5014 ( .IN1(n3002), .IN2(n4529), .QN(n4526) );
  NAND2X0 U5015 ( .IN1(WX6965), .IN2(n3033), .QN(n4525) );
  NAND2X0 U5016 ( .IN1(n3065), .IN2(CRC_OUT_4_22), .QN(n4524) );
  NAND4X0 U5017 ( .IN1(n4530), .IN2(n4531), .IN3(n4532), .IN4(n4533), .QN(
        WX7125) );
  NAND2X0 U5018 ( .IN1(n3092), .IN2(n4311), .QN(n4533) );
  XNOR3X1 U5019 ( .IN1(n2417), .IN2(n3568), .IN3(n4534), .Q(n4311) );
  XOR3X1 U5020 ( .IN1(n6040), .IN2(n2773), .IN3(WX8547), .Q(n4534) );
  NAND2X0 U5021 ( .IN1(n4535), .IN2(n3019), .QN(n4532) );
  NAND2X0 U5022 ( .IN1(WX6963), .IN2(n3033), .QN(n4531) );
  NAND2X0 U5023 ( .IN1(n3065), .IN2(CRC_OUT_4_23), .QN(n4530) );
  NAND4X0 U5024 ( .IN1(n4536), .IN2(n4537), .IN3(n4538), .IN4(n4539), .QN(
        WX7123) );
  NAND2X0 U5025 ( .IN1(n3093), .IN2(n4317), .QN(n4539) );
  XNOR3X1 U5026 ( .IN1(n2419), .IN2(n3568), .IN3(n4540), .Q(n4317) );
  XOR3X1 U5027 ( .IN1(n6041), .IN2(n2772), .IN3(WX8545), .Q(n4540) );
  NAND2X0 U5028 ( .IN1(n3002), .IN2(n4541), .QN(n4538) );
  NAND2X0 U5029 ( .IN1(WX6961), .IN2(n3033), .QN(n4537) );
  NAND2X0 U5030 ( .IN1(n3065), .IN2(CRC_OUT_4_24), .QN(n4536) );
  NAND4X0 U5031 ( .IN1(n4542), .IN2(n4543), .IN3(n4544), .IN4(n4545), .QN(
        WX7121) );
  NAND2X0 U5032 ( .IN1(n3093), .IN2(n4323), .QN(n4545) );
  XNOR3X1 U5033 ( .IN1(n2421), .IN2(n3568), .IN3(n4546), .Q(n4323) );
  XOR3X1 U5034 ( .IN1(n6042), .IN2(n2771), .IN3(WX8543), .Q(n4546) );
  NAND2X0 U5035 ( .IN1(n4547), .IN2(n3019), .QN(n4544) );
  NAND2X0 U5036 ( .IN1(WX6959), .IN2(n3033), .QN(n4543) );
  NAND2X0 U5037 ( .IN1(n3065), .IN2(CRC_OUT_4_25), .QN(n4542) );
  NAND4X0 U5038 ( .IN1(n4548), .IN2(n4549), .IN3(n4550), .IN4(n4551), .QN(
        WX7119) );
  NAND2X0 U5039 ( .IN1(n4329), .IN2(n3099), .QN(n4551) );
  XOR3X1 U5040 ( .IN1(n2423), .IN2(n3579), .IN3(n4552), .Q(n4329) );
  XOR3X1 U5041 ( .IN1(test_so74), .IN2(n6043), .IN3(WX8541), .Q(n4552) );
  NAND2X0 U5042 ( .IN1(n3002), .IN2(n4553), .QN(n4550) );
  NAND2X0 U5043 ( .IN1(WX6957), .IN2(n3033), .QN(n4549) );
  NAND2X0 U5044 ( .IN1(n3066), .IN2(CRC_OUT_4_26), .QN(n4548) );
  NAND4X0 U5045 ( .IN1(n4554), .IN2(n4555), .IN3(n4556), .IN4(n4557), .QN(
        WX7117) );
  NAND2X0 U5046 ( .IN1(n3094), .IN2(n4335), .QN(n4557) );
  XNOR3X1 U5047 ( .IN1(n2424), .IN2(n3568), .IN3(n4558), .Q(n4335) );
  XOR3X1 U5048 ( .IN1(n6044), .IN2(n2770), .IN3(WX8539), .Q(n4558) );
  NAND2X0 U5049 ( .IN1(n4559), .IN2(n3019), .QN(n4556) );
  NAND2X0 U5050 ( .IN1(WX6955), .IN2(n3033), .QN(n4555) );
  NAND2X0 U5051 ( .IN1(n3066), .IN2(CRC_OUT_4_27), .QN(n4554) );
  NAND4X0 U5052 ( .IN1(n4560), .IN2(n4561), .IN3(n4562), .IN4(n4563), .QN(
        WX7115) );
  NAND2X0 U5053 ( .IN1(n4341), .IN2(n3099), .QN(n4563) );
  XOR3X1 U5054 ( .IN1(n2426), .IN2(n3578), .IN3(n4564), .Q(n4341) );
  XNOR3X1 U5055 ( .IN1(test_so72), .IN2(n6045), .IN3(n2769), .Q(n4564) );
  NAND2X0 U5056 ( .IN1(n3002), .IN2(n4565), .QN(n4562) );
  NAND2X0 U5057 ( .IN1(WX6953), .IN2(n3033), .QN(n4561) );
  NAND2X0 U5058 ( .IN1(n3066), .IN2(CRC_OUT_4_28), .QN(n4560) );
  NAND4X0 U5059 ( .IN1(n4566), .IN2(n4567), .IN3(n4568), .IN4(n4569), .QN(
        WX7113) );
  NAND2X0 U5060 ( .IN1(n3093), .IN2(n4347), .QN(n4569) );
  XNOR3X1 U5061 ( .IN1(n2427), .IN2(n3568), .IN3(n4570), .Q(n4347) );
  XOR3X1 U5062 ( .IN1(n6046), .IN2(n2768), .IN3(WX8535), .Q(n4570) );
  NAND2X0 U5063 ( .IN1(n3002), .IN2(n4571), .QN(n4568) );
  NAND2X0 U5064 ( .IN1(WX6951), .IN2(n3033), .QN(n4567) );
  NAND2X0 U5065 ( .IN1(test_so66), .IN2(n3070), .QN(n4566) );
  NAND4X0 U5066 ( .IN1(n4572), .IN2(n4573), .IN3(n4574), .IN4(n4575), .QN(
        WX7111) );
  NAND2X0 U5067 ( .IN1(n4353), .IN2(n3098), .QN(n4575) );
  XOR3X1 U5068 ( .IN1(n2429), .IN2(n3578), .IN3(n4576), .Q(n4353) );
  XNOR3X1 U5069 ( .IN1(test_so70), .IN2(n6047), .IN3(n2767), .Q(n4576) );
  NAND2X0 U5070 ( .IN1(n3002), .IN2(n4577), .QN(n4574) );
  NAND2X0 U5071 ( .IN1(WX6949), .IN2(n3033), .QN(n4573) );
  NAND2X0 U5072 ( .IN1(n3066), .IN2(CRC_OUT_4_30), .QN(n4572) );
  NAND4X0 U5073 ( .IN1(n4578), .IN2(n4579), .IN3(n4580), .IN4(n4581), .QN(
        WX7109) );
  NAND2X0 U5074 ( .IN1(n3093), .IN2(n4359), .QN(n4581) );
  XNOR3X1 U5075 ( .IN1(n2338), .IN2(n3570), .IN3(n4582), .Q(n4359) );
  XOR3X1 U5076 ( .IN1(n6048), .IN2(n2766), .IN3(WX8531), .Q(n4582) );
  NAND2X0 U5077 ( .IN1(n3002), .IN2(n4583), .QN(n4580) );
  NAND2X0 U5078 ( .IN1(n3065), .IN2(CRC_OUT_4_31), .QN(n4579) );
  NAND2X0 U5079 ( .IN1(n2245), .IN2(WX6950), .QN(n4578) );
  NAND4X0 U5080 ( .IN1(n4584), .IN2(n4585), .IN3(n4586), .IN4(n4587), .QN(
        WX706) );
  NAND2X0 U5081 ( .IN1(n4588), .IN2(n3098), .QN(n4587) );
  NAND2X0 U5082 ( .IN1(n3002), .IN2(n4589), .QN(n4586) );
  NAND2X0 U5083 ( .IN1(WX544), .IN2(n3033), .QN(n4585) );
  NAND2X0 U5084 ( .IN1(n3066), .IN2(CRC_OUT_9_0), .QN(n4584) );
  NAND4X0 U5085 ( .IN1(n4590), .IN2(n4591), .IN3(n4592), .IN4(n4593), .QN(
        WX704) );
  NAND2X0 U5086 ( .IN1(n3094), .IN2(n4594), .QN(n4593) );
  NAND2X0 U5087 ( .IN1(n3002), .IN2(n4595), .QN(n4592) );
  NAND2X0 U5088 ( .IN1(WX542), .IN2(n3033), .QN(n4591) );
  NAND2X0 U5089 ( .IN1(test_so9), .IN2(n3070), .QN(n4590) );
  NAND4X0 U5090 ( .IN1(n4596), .IN2(n4597), .IN3(n4598), .IN4(n4599), .QN(
        WX702) );
  NAND2X0 U5091 ( .IN1(n3094), .IN2(n4600), .QN(n4599) );
  NAND2X0 U5092 ( .IN1(n4601), .IN2(n3020), .QN(n4598) );
  NAND2X0 U5093 ( .IN1(WX540), .IN2(n3033), .QN(n4597) );
  NAND2X0 U5094 ( .IN1(n3066), .IN2(CRC_OUT_9_2), .QN(n4596) );
  NOR2X0 U5095 ( .IN1(n3750), .IN2(WX6950), .QN(WX7011) );
  AND2X1 U5096 ( .IN1(n3623), .IN2(n8438), .Q(WX7009) );
  AND2X1 U5097 ( .IN1(n3623), .IN2(n8439), .Q(WX7007) );
  AND2X1 U5098 ( .IN1(n3623), .IN2(n8440), .Q(WX7005) );
  AND2X1 U5099 ( .IN1(n3622), .IN2(n8441), .Q(WX7003) );
  AND2X1 U5100 ( .IN1(n3622), .IN2(n8442), .Q(WX7001) );
  NAND4X0 U5101 ( .IN1(n4602), .IN2(n4603), .IN3(n4604), .IN4(n4605), .QN(
        WX700) );
  NAND2X0 U5102 ( .IN1(n3094), .IN2(n4606), .QN(n4605) );
  NAND2X0 U5103 ( .IN1(n3002), .IN2(n4607), .QN(n4604) );
  NAND2X0 U5104 ( .IN1(WX538), .IN2(n3033), .QN(n4603) );
  NAND2X0 U5105 ( .IN1(n3065), .IN2(CRC_OUT_9_3), .QN(n4602) );
  AND2X1 U5106 ( .IN1(n3622), .IN2(n8443), .Q(WX6999) );
  AND2X1 U5107 ( .IN1(n3622), .IN2(n8444), .Q(WX6997) );
  AND2X1 U5108 ( .IN1(n3622), .IN2(n8445), .Q(WX6995) );
  AND2X1 U5109 ( .IN1(n3622), .IN2(n8446), .Q(WX6993) );
  AND2X1 U5110 ( .IN1(n3622), .IN2(n8447), .Q(WX6991) );
  AND2X1 U5111 ( .IN1(n3622), .IN2(n8448), .Q(WX6989) );
  AND2X1 U5112 ( .IN1(n3622), .IN2(n8449), .Q(WX6987) );
  AND2X1 U5113 ( .IN1(test_so56), .IN2(n3598), .Q(WX6985) );
  AND2X1 U5114 ( .IN1(n3621), .IN2(n8452), .Q(WX6983) );
  AND2X1 U5115 ( .IN1(n3621), .IN2(n8453), .Q(WX6981) );
  NAND4X0 U5116 ( .IN1(n4608), .IN2(n4609), .IN3(n4610), .IN4(n4611), .QN(
        WX698) );
  NAND2X0 U5117 ( .IN1(n4612), .IN2(n3097), .QN(n4611) );
  NAND2X0 U5118 ( .IN1(n3001), .IN2(n4613), .QN(n4610) );
  NAND2X0 U5119 ( .IN1(WX536), .IN2(n3033), .QN(n4609) );
  NAND2X0 U5120 ( .IN1(n3066), .IN2(CRC_OUT_9_4), .QN(n4608) );
  AND2X1 U5121 ( .IN1(n3621), .IN2(n8454), .Q(WX6979) );
  AND2X1 U5122 ( .IN1(n3621), .IN2(n8455), .Q(WX6977) );
  AND2X1 U5123 ( .IN1(n3621), .IN2(n8456), .Q(WX6975) );
  AND2X1 U5124 ( .IN1(n3621), .IN2(n8457), .Q(WX6973) );
  AND2X1 U5125 ( .IN1(n3621), .IN2(n8458), .Q(WX6971) );
  AND2X1 U5126 ( .IN1(n3620), .IN2(n8459), .Q(WX6969) );
  AND2X1 U5127 ( .IN1(n3620), .IN2(n8460), .Q(WX6967) );
  AND2X1 U5128 ( .IN1(n3620), .IN2(n8461), .Q(WX6965) );
  AND2X1 U5129 ( .IN1(n3620), .IN2(n8462), .Q(WX6963) );
  AND2X1 U5130 ( .IN1(n3620), .IN2(n8463), .Q(WX6961) );
  NAND4X0 U5131 ( .IN1(n4614), .IN2(n4615), .IN3(n4616), .IN4(n4617), .QN(
        WX696) );
  NAND2X0 U5132 ( .IN1(n3094), .IN2(n4618), .QN(n4617) );
  NAND2X0 U5133 ( .IN1(n3001), .IN2(n4619), .QN(n4616) );
  NAND2X0 U5134 ( .IN1(WX534), .IN2(n3033), .QN(n4615) );
  NAND2X0 U5135 ( .IN1(n3067), .IN2(CRC_OUT_9_5), .QN(n4614) );
  AND2X1 U5136 ( .IN1(n3620), .IN2(n8464), .Q(WX6959) );
  AND2X1 U5137 ( .IN1(n3620), .IN2(n8465), .Q(WX6957) );
  AND2X1 U5138 ( .IN1(n3620), .IN2(n8466), .Q(WX6955) );
  AND2X1 U5139 ( .IN1(n3620), .IN2(n8467), .Q(WX6953) );
  AND2X1 U5140 ( .IN1(test_so55), .IN2(n3598), .Q(WX6951) );
  AND2X1 U5141 ( .IN1(n3619), .IN2(n8470), .Q(WX6949) );
  NAND4X0 U5142 ( .IN1(n4620), .IN2(n4621), .IN3(n4622), .IN4(n4623), .QN(
        WX694) );
  NAND2X0 U5143 ( .IN1(n3093), .IN2(n4624), .QN(n4623) );
  NAND2X0 U5144 ( .IN1(n4625), .IN2(n3020), .QN(n4622) );
  NAND2X0 U5145 ( .IN1(WX532), .IN2(n3033), .QN(n4621) );
  NAND2X0 U5146 ( .IN1(n3066), .IN2(CRC_OUT_9_6), .QN(n4620) );
  NAND4X0 U5147 ( .IN1(n4626), .IN2(n4627), .IN3(n4628), .IN4(n4629), .QN(
        WX692) );
  NAND2X0 U5148 ( .IN1(n3094), .IN2(n4630), .QN(n4629) );
  NAND2X0 U5149 ( .IN1(n3001), .IN2(n4631), .QN(n4628) );
  NAND2X0 U5150 ( .IN1(WX530), .IN2(n3033), .QN(n4627) );
  NAND2X0 U5151 ( .IN1(n3067), .IN2(CRC_OUT_9_7), .QN(n4626) );
  NAND4X0 U5152 ( .IN1(n4632), .IN2(n4633), .IN3(n4634), .IN4(n4635), .QN(
        WX690) );
  NAND2X0 U5153 ( .IN1(n3092), .IN2(n4636), .QN(n4635) );
  NAND2X0 U5154 ( .IN1(n3001), .IN2(n4637), .QN(n4634) );
  NAND2X0 U5155 ( .IN1(WX528), .IN2(n3034), .QN(n4633) );
  NAND2X0 U5156 ( .IN1(n3065), .IN2(CRC_OUT_9_8), .QN(n4632) );
  NAND4X0 U5157 ( .IN1(n4638), .IN2(n4639), .IN3(n4640), .IN4(n4641), .QN(
        WX688) );
  NAND2X0 U5158 ( .IN1(n3093), .IN2(n4642), .QN(n4641) );
  NAND2X0 U5159 ( .IN1(n3001), .IN2(n4643), .QN(n4640) );
  NAND2X0 U5160 ( .IN1(WX526), .IN2(n3034), .QN(n4639) );
  NAND2X0 U5161 ( .IN1(n3067), .IN2(CRC_OUT_9_9), .QN(n4638) );
  NAND4X0 U5162 ( .IN1(n4644), .IN2(n4645), .IN3(n4646), .IN4(n4647), .QN(
        WX686) );
  NAND2X0 U5163 ( .IN1(n4648), .IN2(n3097), .QN(n4647) );
  NAND2X0 U5164 ( .IN1(n4649), .IN2(n3020), .QN(n4646) );
  NAND2X0 U5165 ( .IN1(WX524), .IN2(n3034), .QN(n4645) );
  NAND2X0 U5166 ( .IN1(n3067), .IN2(CRC_OUT_9_10), .QN(n4644) );
  NAND4X0 U5167 ( .IN1(n4650), .IN2(n4651), .IN3(n4652), .IN4(n4653), .QN(
        WX684) );
  NAND2X0 U5168 ( .IN1(n3093), .IN2(n4654), .QN(n4653) );
  NAND2X0 U5169 ( .IN1(n3001), .IN2(n4655), .QN(n4652) );
  NAND2X0 U5170 ( .IN1(WX522), .IN2(n3034), .QN(n4651) );
  NAND2X0 U5171 ( .IN1(n3067), .IN2(CRC_OUT_9_11), .QN(n4650) );
  NAND4X0 U5172 ( .IN1(n4656), .IN2(n4657), .IN3(n4658), .IN4(n4659), .QN(
        WX682) );
  NAND2X0 U5173 ( .IN1(n3093), .IN2(n4660), .QN(n4659) );
  NAND2X0 U5174 ( .IN1(n3001), .IN2(n4661), .QN(n4658) );
  NAND2X0 U5175 ( .IN1(WX520), .IN2(n3034), .QN(n4657) );
  NAND2X0 U5176 ( .IN1(n3066), .IN2(CRC_OUT_9_12), .QN(n4656) );
  NAND4X0 U5177 ( .IN1(n4662), .IN2(n4663), .IN3(n4664), .IN4(n4665), .QN(
        WX680) );
  NAND2X0 U5178 ( .IN1(n3092), .IN2(n4666), .QN(n4665) );
  NAND2X0 U5179 ( .IN1(n3001), .IN2(n4667), .QN(n4664) );
  NAND2X0 U5180 ( .IN1(WX518), .IN2(n3034), .QN(n4663) );
  NAND2X0 U5181 ( .IN1(n3064), .IN2(CRC_OUT_9_13), .QN(n4662) );
  NAND4X0 U5182 ( .IN1(n4668), .IN2(n4669), .IN3(n4670), .IN4(n4671), .QN(
        WX678) );
  NAND2X0 U5183 ( .IN1(n4672), .IN2(n3096), .QN(n4671) );
  NAND2X0 U5184 ( .IN1(n3001), .IN2(n4673), .QN(n4670) );
  NAND2X0 U5185 ( .IN1(WX516), .IN2(n3034), .QN(n4669) );
  NAND2X0 U5186 ( .IN1(n3066), .IN2(CRC_OUT_9_14), .QN(n4668) );
  NAND4X0 U5187 ( .IN1(n4674), .IN2(n4675), .IN3(n4676), .IN4(n4677), .QN(
        WX676) );
  NAND2X0 U5188 ( .IN1(n3092), .IN2(n4678), .QN(n4677) );
  NAND2X0 U5189 ( .IN1(n3001), .IN2(n4679), .QN(n4676) );
  NAND2X0 U5190 ( .IN1(WX514), .IN2(n3034), .QN(n4675) );
  NAND2X0 U5191 ( .IN1(n3068), .IN2(CRC_OUT_9_15), .QN(n4674) );
  NAND4X0 U5192 ( .IN1(n4680), .IN2(n4681), .IN3(n4682), .IN4(n4683), .QN(
        WX674) );
  NAND2X0 U5193 ( .IN1(n3082), .IN2(n4684), .QN(n4683) );
  NAND2X0 U5194 ( .IN1(n4685), .IN2(n3018), .QN(n4682) );
  NAND2X0 U5195 ( .IN1(WX512), .IN2(n3034), .QN(n4681) );
  NAND2X0 U5196 ( .IN1(n3067), .IN2(CRC_OUT_9_16), .QN(n4680) );
  NAND4X0 U5197 ( .IN1(n4686), .IN2(n4687), .IN3(n4688), .IN4(n4689), .QN(
        WX672) );
  NAND2X0 U5198 ( .IN1(n3078), .IN2(n4690), .QN(n4689) );
  NAND2X0 U5199 ( .IN1(n3001), .IN2(n4691), .QN(n4688) );
  NAND2X0 U5200 ( .IN1(WX510), .IN2(n3034), .QN(n4687) );
  NAND2X0 U5201 ( .IN1(n3068), .IN2(CRC_OUT_9_17), .QN(n4686) );
  NAND4X0 U5202 ( .IN1(n4692), .IN2(n4693), .IN3(n4694), .IN4(n4695), .QN(
        WX670) );
  NAND2X0 U5203 ( .IN1(n4696), .IN2(n3096), .QN(n4695) );
  NAND2X0 U5204 ( .IN1(n3001), .IN2(n4697), .QN(n4694) );
  NAND2X0 U5205 ( .IN1(WX508), .IN2(n3034), .QN(n4693) );
  NAND2X0 U5206 ( .IN1(n3066), .IN2(CRC_OUT_9_18), .QN(n4692) );
  NAND4X0 U5207 ( .IN1(n4698), .IN2(n4699), .IN3(n4700), .IN4(n4701), .QN(
        WX668) );
  NAND2X0 U5208 ( .IN1(n3078), .IN2(n4702), .QN(n4701) );
  NAND2X0 U5209 ( .IN1(n3000), .IN2(n4703), .QN(n4700) );
  NAND2X0 U5210 ( .IN1(WX506), .IN2(n3034), .QN(n4699) );
  NAND2X0 U5211 ( .IN1(test_so10), .IN2(n3069), .QN(n4698) );
  NAND4X0 U5212 ( .IN1(n4704), .IN2(n4705), .IN3(n4706), .IN4(n4707), .QN(
        WX666) );
  NAND2X0 U5213 ( .IN1(n3078), .IN2(n4708), .QN(n4707) );
  NAND2X0 U5214 ( .IN1(n4709), .IN2(n3016), .QN(n4706) );
  NAND2X0 U5215 ( .IN1(WX504), .IN2(n3034), .QN(n4705) );
  NAND2X0 U5216 ( .IN1(n3068), .IN2(CRC_OUT_9_20), .QN(n4704) );
  NAND4X0 U5217 ( .IN1(n4710), .IN2(n4711), .IN3(n4712), .IN4(n4713), .QN(
        WX664) );
  NAND2X0 U5218 ( .IN1(n3078), .IN2(n4714), .QN(n4713) );
  NAND2X0 U5219 ( .IN1(n3000), .IN2(n4715), .QN(n4712) );
  NAND2X0 U5220 ( .IN1(WX502), .IN2(n3034), .QN(n4711) );
  NAND2X0 U5221 ( .IN1(n3067), .IN2(CRC_OUT_9_21), .QN(n4710) );
  NAND4X0 U5222 ( .IN1(n4716), .IN2(n4717), .IN3(n4718), .IN4(n4719), .QN(
        WX662) );
  NAND2X0 U5223 ( .IN1(n4720), .IN2(n3097), .QN(n4719) );
  NAND2X0 U5224 ( .IN1(n3000), .IN2(n4721), .QN(n4718) );
  NAND2X0 U5225 ( .IN1(WX500), .IN2(n3034), .QN(n4717) );
  NAND2X0 U5226 ( .IN1(n3068), .IN2(CRC_OUT_9_22), .QN(n4716) );
  NAND4X0 U5227 ( .IN1(n4722), .IN2(n4723), .IN3(n4724), .IN4(n4725), .QN(
        WX660) );
  NAND2X0 U5228 ( .IN1(n3078), .IN2(n4726), .QN(n4725) );
  NAND2X0 U5229 ( .IN1(n3000), .IN2(n4727), .QN(n4724) );
  NAND2X0 U5230 ( .IN1(WX498), .IN2(n3034), .QN(n4723) );
  NAND2X0 U5231 ( .IN1(n3066), .IN2(CRC_OUT_9_23), .QN(n4722) );
  NAND4X0 U5232 ( .IN1(n4728), .IN2(n4729), .IN3(n4730), .IN4(n4731), .QN(
        WX658) );
  NAND2X0 U5233 ( .IN1(n3078), .IN2(n4732), .QN(n4731) );
  NAND2X0 U5234 ( .IN1(n4733), .IN2(n3016), .QN(n4730) );
  NAND2X0 U5235 ( .IN1(WX496), .IN2(n3034), .QN(n4729) );
  NAND2X0 U5236 ( .IN1(n3068), .IN2(CRC_OUT_9_24), .QN(n4728) );
  NAND4X0 U5237 ( .IN1(n4734), .IN2(n4735), .IN3(n4736), .IN4(n4737), .QN(
        WX656) );
  NAND2X0 U5238 ( .IN1(n3078), .IN2(n4738), .QN(n4737) );
  NAND2X0 U5239 ( .IN1(n3000), .IN2(n4739), .QN(n4736) );
  NAND2X0 U5240 ( .IN1(WX494), .IN2(n3035), .QN(n4735) );
  NAND2X0 U5241 ( .IN1(n3067), .IN2(CRC_OUT_9_25), .QN(n4734) );
  NAND4X0 U5242 ( .IN1(n4740), .IN2(n4741), .IN3(n4742), .IN4(n4743), .QN(
        WX654) );
  NAND2X0 U5243 ( .IN1(n3078), .IN2(n4744), .QN(n4743) );
  NAND2X0 U5244 ( .IN1(n3000), .IN2(n4745), .QN(n4742) );
  NAND2X0 U5245 ( .IN1(WX492), .IN2(n3035), .QN(n4741) );
  NAND2X0 U5246 ( .IN1(n3068), .IN2(CRC_OUT_9_26), .QN(n4740) );
  NAND4X0 U5247 ( .IN1(n4746), .IN2(n4747), .IN3(n4748), .IN4(n4749), .QN(
        WX652) );
  NAND2X0 U5248 ( .IN1(n3078), .IN2(n4750), .QN(n4749) );
  NAND2X0 U5249 ( .IN1(n3000), .IN2(n4751), .QN(n4748) );
  NAND2X0 U5250 ( .IN1(WX490), .IN2(n3035), .QN(n4747) );
  NAND2X0 U5251 ( .IN1(n3067), .IN2(CRC_OUT_9_27), .QN(n4746) );
  NAND4X0 U5252 ( .IN1(n4752), .IN2(n4753), .IN3(n4754), .IN4(n4755), .QN(
        WX650) );
  NAND2X0 U5253 ( .IN1(n4756), .IN2(n3097), .QN(n4755) );
  NAND2X0 U5254 ( .IN1(n4757), .IN2(n3016), .QN(n4754) );
  NAND2X0 U5255 ( .IN1(WX488), .IN2(n3035), .QN(n4753) );
  NAND2X0 U5256 ( .IN1(n3067), .IN2(CRC_OUT_9_28), .QN(n4752) );
  NOR2X0 U5257 ( .IN1(n3750), .IN2(n4758), .QN(WX6498) );
  XOR2X1 U5258 ( .IN1(n2819), .IN2(DFF_958_n1), .Q(n4758) );
  NOR2X0 U5259 ( .IN1(n3750), .IN2(n4759), .QN(WX6496) );
  XOR2X1 U5260 ( .IN1(n2820), .IN2(DFF_957_n1), .Q(n4759) );
  NOR2X0 U5261 ( .IN1(n3750), .IN2(n4760), .QN(WX6494) );
  XOR2X1 U5262 ( .IN1(n2821), .IN2(DFF_956_n1), .Q(n4760) );
  NOR2X0 U5263 ( .IN1(n3750), .IN2(n4761), .QN(WX6492) );
  XOR2X1 U5264 ( .IN1(n2822), .IN2(DFF_955_n1), .Q(n4761) );
  NOR2X0 U5265 ( .IN1(n3750), .IN2(n4762), .QN(WX6490) );
  XOR2X1 U5266 ( .IN1(n2823), .IN2(DFF_954_n1), .Q(n4762) );
  NOR2X0 U5267 ( .IN1(n3750), .IN2(n4763), .QN(WX6488) );
  XOR2X1 U5268 ( .IN1(n2824), .IN2(DFF_953_n1), .Q(n4763) );
  NOR2X0 U5269 ( .IN1(n3750), .IN2(n4764), .QN(WX6486) );
  XOR2X1 U5270 ( .IN1(n2825), .IN2(DFF_952_n1), .Q(n4764) );
  NOR2X0 U5271 ( .IN1(n3750), .IN2(n4765), .QN(WX6484) );
  XOR2X1 U5272 ( .IN1(n2826), .IN2(DFF_951_n1), .Q(n4765) );
  NOR2X0 U5273 ( .IN1(n3750), .IN2(n4766), .QN(WX6482) );
  XOR2X1 U5274 ( .IN1(n2827), .IN2(DFF_950_n1), .Q(n4766) );
  NOR2X0 U5275 ( .IN1(n3750), .IN2(n4767), .QN(WX6480) );
  XOR2X1 U5276 ( .IN1(n2828), .IN2(DFF_949_n1), .Q(n4767) );
  NAND4X0 U5277 ( .IN1(n4768), .IN2(n4769), .IN3(n4770), .IN4(n4771), .QN(
        WX648) );
  NAND2X0 U5278 ( .IN1(n3078), .IN2(n4772), .QN(n4771) );
  NAND2X0 U5279 ( .IN1(n3000), .IN2(n4773), .QN(n4770) );
  NAND2X0 U5280 ( .IN1(WX486), .IN2(n3035), .QN(n4769) );
  NAND2X0 U5281 ( .IN1(n3068), .IN2(CRC_OUT_9_29), .QN(n4768) );
  NOR2X0 U5282 ( .IN1(n3750), .IN2(n4774), .QN(WX6478) );
  XOR2X1 U5283 ( .IN1(n2829), .IN2(DFF_948_n1), .Q(n4774) );
  NOR2X0 U5284 ( .IN1(n3751), .IN2(n4775), .QN(WX6476) );
  XOR2X1 U5285 ( .IN1(n2830), .IN2(DFF_947_n1), .Q(n4775) );
  NOR2X0 U5286 ( .IN1(n3751), .IN2(n4776), .QN(WX6474) );
  XOR2X1 U5287 ( .IN1(n2831), .IN2(DFF_946_n1), .Q(n4776) );
  NOR2X0 U5288 ( .IN1(n3751), .IN2(n4777), .QN(WX6472) );
  XNOR2X1 U5289 ( .IN1(n2832), .IN2(test_so54), .Q(n4777) );
  NOR2X0 U5290 ( .IN1(n3751), .IN2(n4778), .QN(WX6470) );
  XOR2X1 U5291 ( .IN1(n2833), .IN2(DFF_944_n1), .Q(n4778) );
  NOR2X0 U5292 ( .IN1(n3751), .IN2(n4779), .QN(WX6468) );
  XOR3X1 U5293 ( .IN1(test_so52), .IN2(DFF_959_n1), .IN3(DFF_943_n1), .Q(n4779) );
  NOR2X0 U5294 ( .IN1(n3751), .IN2(n4780), .QN(WX6466) );
  XOR2X1 U5295 ( .IN1(n2834), .IN2(DFF_942_n1), .Q(n4780) );
  NOR2X0 U5296 ( .IN1(n3751), .IN2(n4781), .QN(WX6464) );
  XOR2X1 U5297 ( .IN1(n2835), .IN2(DFF_941_n1), .Q(n4781) );
  NOR2X0 U5298 ( .IN1(n3751), .IN2(n4782), .QN(WX6462) );
  XOR2X1 U5299 ( .IN1(n2836), .IN2(DFF_940_n1), .Q(n4782) );
  NOR2X0 U5300 ( .IN1(n3751), .IN2(n4783), .QN(WX6460) );
  XOR2X1 U5301 ( .IN1(n2837), .IN2(DFF_939_n1), .Q(n4783) );
  NAND4X0 U5302 ( .IN1(n4784), .IN2(n4785), .IN3(n4786), .IN4(n4787), .QN(
        WX646) );
  NAND2X0 U5303 ( .IN1(n3078), .IN2(n4788), .QN(n4787) );
  NAND2X0 U5304 ( .IN1(n3000), .IN2(n4789), .QN(n4786) );
  NAND2X0 U5305 ( .IN1(WX484), .IN2(n3035), .QN(n4785) );
  NAND2X0 U5306 ( .IN1(n3069), .IN2(CRC_OUT_9_30), .QN(n4784) );
  NOR2X0 U5307 ( .IN1(n3751), .IN2(n4790), .QN(WX6458) );
  XOR3X1 U5308 ( .IN1(n2696), .IN2(DFF_959_n1), .IN3(CRC_OUT_5_10), .Q(n4790)
         );
  NOR2X0 U5309 ( .IN1(n3751), .IN2(n4791), .QN(WX6456) );
  XOR2X1 U5310 ( .IN1(n2838), .IN2(DFF_937_n1), .Q(n4791) );
  NOR2X0 U5311 ( .IN1(n3751), .IN2(n4792), .QN(WX6454) );
  XOR2X1 U5312 ( .IN1(n2839), .IN2(DFF_936_n1), .Q(n4792) );
  NOR2X0 U5313 ( .IN1(n3752), .IN2(n4793), .QN(WX6452) );
  XOR2X1 U5314 ( .IN1(n2840), .IN2(DFF_935_n1), .Q(n4793) );
  NOR2X0 U5315 ( .IN1(n3752), .IN2(n4794), .QN(WX6450) );
  XOR2X1 U5316 ( .IN1(n2841), .IN2(DFF_934_n1), .Q(n4794) );
  NOR2X0 U5317 ( .IN1(n3752), .IN2(n4795), .QN(WX6448) );
  XOR2X1 U5318 ( .IN1(n2842), .IN2(DFF_933_n1), .Q(n4795) );
  NOR2X0 U5319 ( .IN1(n3752), .IN2(n4796), .QN(WX6446) );
  XOR2X1 U5320 ( .IN1(n2843), .IN2(DFF_932_n1), .Q(n4796) );
  NOR2X0 U5321 ( .IN1(n3752), .IN2(n4797), .QN(WX6444) );
  XOR3X1 U5322 ( .IN1(n2697), .IN2(DFF_959_n1), .IN3(CRC_OUT_5_3), .Q(n4797)
         );
  NOR2X0 U5323 ( .IN1(n3752), .IN2(n4798), .QN(WX6442) );
  XOR2X1 U5324 ( .IN1(n2844), .IN2(DFF_930_n1), .Q(n4798) );
  NOR2X0 U5325 ( .IN1(n3752), .IN2(n4799), .QN(WX6440) );
  XOR2X1 U5326 ( .IN1(n2845), .IN2(DFF_929_n1), .Q(n4799) );
  NAND4X0 U5327 ( .IN1(n4800), .IN2(n4801), .IN3(n4802), .IN4(n4803), .QN(
        WX644) );
  NAND2X0 U5328 ( .IN1(n3079), .IN2(n4804), .QN(n4803) );
  NAND2X0 U5329 ( .IN1(n3000), .IN2(n4805), .QN(n4802) );
  NAND2X0 U5330 ( .IN1(n3068), .IN2(CRC_OUT_9_31), .QN(n4801) );
  NAND2X0 U5331 ( .IN1(n2245), .IN2(WX485), .QN(n4800) );
  NOR2X0 U5332 ( .IN1(n3752), .IN2(n4806), .QN(WX6438) );
  XNOR2X1 U5333 ( .IN1(n2846), .IN2(test_so53), .Q(n4806) );
  NOR2X0 U5334 ( .IN1(n3752), .IN2(n4807), .QN(WX6436) );
  XOR2X1 U5335 ( .IN1(n2710), .IN2(DFF_959_n1), .Q(n4807) );
  NOR2X0 U5336 ( .IN1(n6090), .IN2(n3655), .QN(WX5910) );
  NOR2X0 U5337 ( .IN1(n6091), .IN2(n3656), .QN(WX5908) );
  NOR2X0 U5338 ( .IN1(n6092), .IN2(n3656), .QN(WX5906) );
  NOR2X0 U5339 ( .IN1(n6093), .IN2(n3656), .QN(WX5904) );
  NOR2X0 U5340 ( .IN1(n6094), .IN2(n3656), .QN(WX5902) );
  NOR2X0 U5341 ( .IN1(n6095), .IN2(n3656), .QN(WX5900) );
  AND2X1 U5342 ( .IN1(n3619), .IN2(test_so46), .Q(WX5898) );
  NOR2X0 U5343 ( .IN1(n6097), .IN2(n3656), .QN(WX5896) );
  NOR2X0 U5344 ( .IN1(n6098), .IN2(n3656), .QN(WX5894) );
  NOR2X0 U5345 ( .IN1(n6099), .IN2(n3656), .QN(WX5892) );
  NOR2X0 U5346 ( .IN1(n6100), .IN2(n3656), .QN(WX5890) );
  NOR2X0 U5347 ( .IN1(n6101), .IN2(n3656), .QN(WX5888) );
  NOR2X0 U5348 ( .IN1(n6102), .IN2(n3656), .QN(WX5886) );
  NOR2X0 U5349 ( .IN1(n6103), .IN2(n3656), .QN(WX5884) );
  NOR2X0 U5350 ( .IN1(n6104), .IN2(n3657), .QN(WX5882) );
  NOR2X0 U5351 ( .IN1(n6105), .IN2(n3730), .QN(WX5880) );
  NAND4X0 U5352 ( .IN1(n4808), .IN2(n4809), .IN3(n4810), .IN4(n4811), .QN(
        WX5878) );
  NAND2X0 U5353 ( .IN1(n3079), .IN2(n4397), .QN(n4811) );
  XNOR3X1 U5354 ( .IN1(n2709), .IN2(n2605), .IN3(n4812), .Q(n4397) );
  XOR2X1 U5355 ( .IN1(WX7236), .IN2(n6049), .Q(n4812) );
  NAND2X0 U5356 ( .IN1(n3000), .IN2(n4813), .QN(n4810) );
  NAND2X0 U5357 ( .IN1(WX5716), .IN2(n3035), .QN(n4809) );
  NAND2X0 U5358 ( .IN1(test_so53), .IN2(n3070), .QN(n4808) );
  NAND4X0 U5359 ( .IN1(n4814), .IN2(n4815), .IN3(n4816), .IN4(n4817), .QN(
        WX5876) );
  NAND2X0 U5360 ( .IN1(n3079), .IN2(n4403), .QN(n4817) );
  XNOR3X1 U5361 ( .IN1(n2818), .IN2(n2606), .IN3(n4818), .Q(n4403) );
  XOR2X1 U5362 ( .IN1(WX7234), .IN2(n6050), .Q(n4818) );
  NAND2X0 U5363 ( .IN1(n4819), .IN2(n3017), .QN(n4816) );
  NAND2X0 U5364 ( .IN1(WX5714), .IN2(n3035), .QN(n4815) );
  NAND2X0 U5365 ( .IN1(n3067), .IN2(CRC_OUT_5_1), .QN(n4814) );
  NAND4X0 U5366 ( .IN1(n4820), .IN2(n4821), .IN3(n4822), .IN4(n4823), .QN(
        WX5874) );
  NAND2X0 U5367 ( .IN1(n3079), .IN2(n4409), .QN(n4823) );
  XNOR3X1 U5368 ( .IN1(n2817), .IN2(n2607), .IN3(n4824), .Q(n4409) );
  XOR2X1 U5369 ( .IN1(WX7232), .IN2(n6051), .Q(n4824) );
  NAND2X0 U5370 ( .IN1(n3000), .IN2(n4825), .QN(n4822) );
  NAND2X0 U5371 ( .IN1(WX5712), .IN2(n3035), .QN(n4821) );
  NAND2X0 U5372 ( .IN1(n3069), .IN2(CRC_OUT_5_2), .QN(n4820) );
  NAND4X0 U5373 ( .IN1(n4826), .IN2(n4827), .IN3(n4828), .IN4(n4829), .QN(
        WX5872) );
  NAND2X0 U5374 ( .IN1(n3079), .IN2(n4415), .QN(n4829) );
  XNOR3X1 U5375 ( .IN1(n2816), .IN2(n2608), .IN3(n4830), .Q(n4415) );
  XOR2X1 U5376 ( .IN1(WX7230), .IN2(n6052), .Q(n4830) );
  NAND2X0 U5377 ( .IN1(n4831), .IN2(n3018), .QN(n4828) );
  NAND2X0 U5378 ( .IN1(WX5710), .IN2(n3035), .QN(n4827) );
  NAND2X0 U5379 ( .IN1(n3068), .IN2(CRC_OUT_5_3), .QN(n4826) );
  NAND4X0 U5380 ( .IN1(n4832), .IN2(n4833), .IN3(n4834), .IN4(n4835), .QN(
        WX5870) );
  NAND2X0 U5381 ( .IN1(n4421), .IN2(n3098), .QN(n4835) );
  XOR3X1 U5382 ( .IN1(n3635), .IN2(n2609), .IN3(n4836), .Q(n4421) );
  XOR2X1 U5383 ( .IN1(WX7164), .IN2(test_so64), .Q(n4836) );
  NAND2X0 U5384 ( .IN1(n2999), .IN2(n4837), .QN(n4834) );
  NAND2X0 U5385 ( .IN1(WX5708), .IN2(n3035), .QN(n4833) );
  NAND2X0 U5386 ( .IN1(n3069), .IN2(CRC_OUT_5_4), .QN(n4832) );
  NAND4X0 U5387 ( .IN1(n4838), .IN2(n4839), .IN3(n4840), .IN4(n4841), .QN(
        WX5868) );
  NAND2X0 U5388 ( .IN1(n3079), .IN2(n4427), .QN(n4841) );
  XNOR3X1 U5389 ( .IN1(n2815), .IN2(n2610), .IN3(n4842), .Q(n4427) );
  XOR2X1 U5390 ( .IN1(WX7226), .IN2(n6053), .Q(n4842) );
  NAND2X0 U5391 ( .IN1(n4843), .IN2(n3018), .QN(n4840) );
  NAND2X0 U5392 ( .IN1(WX5706), .IN2(n3035), .QN(n4839) );
  NAND2X0 U5393 ( .IN1(n3068), .IN2(CRC_OUT_5_5), .QN(n4838) );
  NAND4X0 U5394 ( .IN1(n4844), .IN2(n4845), .IN3(n4846), .IN4(n4847), .QN(
        WX5866) );
  NAND2X0 U5395 ( .IN1(n4433), .IN2(n3098), .QN(n4847) );
  XOR3X1 U5396 ( .IN1(n3639), .IN2(n2814), .IN3(n4848), .Q(n4433) );
  XOR2X1 U5397 ( .IN1(WX7160), .IN2(test_so62), .Q(n4848) );
  NAND2X0 U5398 ( .IN1(n2999), .IN2(n4849), .QN(n4846) );
  NAND2X0 U5399 ( .IN1(WX5704), .IN2(n3035), .QN(n4845) );
  NAND2X0 U5400 ( .IN1(n3069), .IN2(CRC_OUT_5_6), .QN(n4844) );
  NAND4X0 U5401 ( .IN1(n4850), .IN2(n4851), .IN3(n4852), .IN4(n4853), .QN(
        WX5864) );
  NAND2X0 U5402 ( .IN1(n3079), .IN2(n4439), .QN(n4853) );
  XNOR3X1 U5403 ( .IN1(n2813), .IN2(n2611), .IN3(n4854), .Q(n4439) );
  XOR2X1 U5404 ( .IN1(WX7222), .IN2(n6054), .Q(n4854) );
  NAND2X0 U5405 ( .IN1(n2999), .IN2(n4855), .QN(n4852) );
  NAND2X0 U5406 ( .IN1(WX5702), .IN2(n3035), .QN(n4851) );
  NAND2X0 U5407 ( .IN1(n3069), .IN2(CRC_OUT_5_7), .QN(n4850) );
  NAND4X0 U5408 ( .IN1(n4856), .IN2(n4857), .IN3(n4858), .IN4(n4859), .QN(
        WX5862) );
  NAND2X0 U5409 ( .IN1(n4445), .IN2(n3098), .QN(n4859) );
  XOR3X1 U5410 ( .IN1(n2812), .IN2(n2612), .IN3(n4860), .Q(n4445) );
  XOR2X1 U5411 ( .IN1(WX7156), .IN2(test_so60), .Q(n4860) );
  NAND2X0 U5412 ( .IN1(n2999), .IN2(n4861), .QN(n4858) );
  NAND2X0 U5413 ( .IN1(WX5700), .IN2(n3035), .QN(n4857) );
  NAND2X0 U5414 ( .IN1(n3068), .IN2(CRC_OUT_5_8), .QN(n4856) );
  NAND4X0 U5415 ( .IN1(n4862), .IN2(n4863), .IN3(n4864), .IN4(n4865), .QN(
        WX5860) );
  NAND2X0 U5416 ( .IN1(n3079), .IN2(n4451), .QN(n4865) );
  XNOR3X1 U5417 ( .IN1(n2811), .IN2(n2613), .IN3(n4866), .Q(n4451) );
  XOR2X1 U5418 ( .IN1(WX7218), .IN2(n6055), .Q(n4866) );
  NAND2X0 U5419 ( .IN1(n2999), .IN2(n4867), .QN(n4864) );
  NAND2X0 U5420 ( .IN1(WX5698), .IN2(n3035), .QN(n4863) );
  NAND2X0 U5421 ( .IN1(n3069), .IN2(CRC_OUT_5_9), .QN(n4862) );
  NAND4X0 U5422 ( .IN1(n4868), .IN2(n4869), .IN3(n4870), .IN4(n4871), .QN(
        WX5858) );
  NAND2X0 U5423 ( .IN1(n4457), .IN2(n3099), .QN(n4871) );
  XOR3X1 U5424 ( .IN1(n3647), .IN2(n2810), .IN3(n4872), .Q(n4457) );
  XOR2X1 U5425 ( .IN1(WX7280), .IN2(test_so58), .Q(n4872) );
  NAND2X0 U5426 ( .IN1(n2999), .IN2(n4873), .QN(n4870) );
  NAND2X0 U5427 ( .IN1(WX5696), .IN2(n3035), .QN(n4869) );
  NAND2X0 U5428 ( .IN1(n3068), .IN2(CRC_OUT_5_10), .QN(n4868) );
  NAND4X0 U5429 ( .IN1(n4874), .IN2(n4875), .IN3(n4876), .IN4(n4877), .QN(
        WX5856) );
  NAND2X0 U5430 ( .IN1(n3079), .IN2(n4463), .QN(n4877) );
  XNOR3X1 U5431 ( .IN1(n2695), .IN2(n2614), .IN3(n4878), .Q(n4463) );
  XOR2X1 U5432 ( .IN1(WX7214), .IN2(n6056), .Q(n4878) );
  NAND2X0 U5433 ( .IN1(n2999), .IN2(n4879), .QN(n4876) );
  NAND2X0 U5434 ( .IN1(WX5694), .IN2(n3036), .QN(n4875) );
  NAND2X0 U5435 ( .IN1(n3067), .IN2(CRC_OUT_5_11), .QN(n4874) );
  NAND4X0 U5436 ( .IN1(n4880), .IN2(n4881), .IN3(n4882), .IN4(n4883), .QN(
        WX5854) );
  NAND2X0 U5437 ( .IN1(n3079), .IN2(n4469), .QN(n4883) );
  XNOR3X1 U5438 ( .IN1(n2809), .IN2(n2615), .IN3(n4884), .Q(n4469) );
  XOR2X1 U5439 ( .IN1(WX7212), .IN2(n6057), .Q(n4884) );
  NAND2X0 U5440 ( .IN1(n2999), .IN2(n4885), .QN(n4882) );
  NAND2X0 U5441 ( .IN1(WX5692), .IN2(n3036), .QN(n4881) );
  NAND2X0 U5442 ( .IN1(n3052), .IN2(CRC_OUT_5_12), .QN(n4880) );
  NAND4X0 U5443 ( .IN1(n4886), .IN2(n4887), .IN3(n4888), .IN4(n4889), .QN(
        WX5852) );
  NAND2X0 U5444 ( .IN1(n3079), .IN2(n4475), .QN(n4889) );
  XNOR3X1 U5445 ( .IN1(n2808), .IN2(n2616), .IN3(n4890), .Q(n4475) );
  XOR2X1 U5446 ( .IN1(WX7210), .IN2(n6058), .Q(n4890) );
  NAND2X0 U5447 ( .IN1(n2999), .IN2(n4891), .QN(n4888) );
  NAND2X0 U5448 ( .IN1(WX5690), .IN2(n3036), .QN(n4887) );
  NAND2X0 U5449 ( .IN1(n3047), .IN2(CRC_OUT_5_13), .QN(n4886) );
  NAND4X0 U5450 ( .IN1(n4892), .IN2(n4893), .IN3(n4894), .IN4(n4895), .QN(
        WX5850) );
  NAND2X0 U5451 ( .IN1(n3079), .IN2(n4481), .QN(n4895) );
  XNOR3X1 U5452 ( .IN1(n2807), .IN2(n2617), .IN3(n4896), .Q(n4481) );
  XOR2X1 U5453 ( .IN1(WX7208), .IN2(n6059), .Q(n4896) );
  NAND2X0 U5454 ( .IN1(n2999), .IN2(n4897), .QN(n4894) );
  NAND2X0 U5455 ( .IN1(WX5688), .IN2(n3036), .QN(n4893) );
  NAND2X0 U5456 ( .IN1(n3047), .IN2(CRC_OUT_5_14), .QN(n4892) );
  NAND4X0 U5457 ( .IN1(n4898), .IN2(n4899), .IN3(n4900), .IN4(n4901), .QN(
        WX5848) );
  NAND2X0 U5458 ( .IN1(n3080), .IN2(n4487), .QN(n4901) );
  XNOR3X1 U5459 ( .IN1(n2806), .IN2(n2618), .IN3(n4902), .Q(n4487) );
  XOR2X1 U5460 ( .IN1(WX7206), .IN2(n6060), .Q(n4902) );
  NAND2X0 U5461 ( .IN1(n2999), .IN2(n4903), .QN(n4900) );
  NAND2X0 U5462 ( .IN1(WX5686), .IN2(n3036), .QN(n4899) );
  NAND2X0 U5463 ( .IN1(n3047), .IN2(CRC_OUT_5_15), .QN(n4898) );
  NAND4X0 U5464 ( .IN1(n4904), .IN2(n4905), .IN3(n4906), .IN4(n4907), .QN(
        WX5846) );
  NAND2X0 U5465 ( .IN1(n3080), .IN2(n4493), .QN(n4907) );
  XNOR3X1 U5466 ( .IN1(n2430), .IN2(n3570), .IN3(n4908), .Q(n4493) );
  XOR3X1 U5467 ( .IN1(n6061), .IN2(n2694), .IN3(WX7268), .Q(n4908) );
  NAND2X0 U5468 ( .IN1(n4909), .IN2(n3019), .QN(n4906) );
  NAND2X0 U5469 ( .IN1(WX5684), .IN2(n3036), .QN(n4905) );
  NAND2X0 U5470 ( .IN1(n3047), .IN2(CRC_OUT_5_16), .QN(n4904) );
  NAND4X0 U5471 ( .IN1(n4910), .IN2(n4911), .IN3(n4912), .IN4(n4913), .QN(
        WX5844) );
  NAND2X0 U5472 ( .IN1(n3080), .IN2(n4499), .QN(n4913) );
  XNOR3X1 U5473 ( .IN1(n2432), .IN2(n3570), .IN3(n4914), .Q(n4499) );
  XOR3X1 U5474 ( .IN1(n6062), .IN2(n2805), .IN3(WX7266), .Q(n4914) );
  NAND2X0 U5475 ( .IN1(n2999), .IN2(n4915), .QN(n4912) );
  NAND2X0 U5476 ( .IN1(WX5682), .IN2(n3036), .QN(n4911) );
  NAND2X0 U5477 ( .IN1(test_so54), .IN2(n3070), .QN(n4910) );
  NAND4X0 U5478 ( .IN1(n4916), .IN2(n4917), .IN3(n4918), .IN4(n4919), .QN(
        WX5842) );
  NAND2X0 U5479 ( .IN1(n3080), .IN2(n4505), .QN(n4919) );
  XNOR3X1 U5480 ( .IN1(n2434), .IN2(n3570), .IN3(n4920), .Q(n4505) );
  XOR3X1 U5481 ( .IN1(n6063), .IN2(n2804), .IN3(WX7264), .Q(n4920) );
  NAND2X0 U5482 ( .IN1(n4921), .IN2(n3019), .QN(n4918) );
  NAND2X0 U5483 ( .IN1(WX5680), .IN2(n3036), .QN(n4917) );
  NAND2X0 U5484 ( .IN1(n3047), .IN2(CRC_OUT_5_18), .QN(n4916) );
  NAND4X0 U5485 ( .IN1(n4922), .IN2(n4923), .IN3(n4924), .IN4(n4925), .QN(
        WX5840) );
  NAND2X0 U5486 ( .IN1(n3080), .IN2(n4511), .QN(n4925) );
  XNOR3X1 U5487 ( .IN1(n2436), .IN2(n3570), .IN3(n4926), .Q(n4511) );
  XOR3X1 U5488 ( .IN1(n6064), .IN2(n2803), .IN3(WX7262), .Q(n4926) );
  NAND2X0 U5489 ( .IN1(n2998), .IN2(n4927), .QN(n4924) );
  NAND2X0 U5490 ( .IN1(WX5678), .IN2(n3036), .QN(n4923) );
  NAND2X0 U5491 ( .IN1(n3047), .IN2(CRC_OUT_5_19), .QN(n4922) );
  NAND4X0 U5492 ( .IN1(n4928), .IN2(n4929), .IN3(n4930), .IN4(n4931), .QN(
        WX5838) );
  NAND2X0 U5493 ( .IN1(n3080), .IN2(n4517), .QN(n4931) );
  XNOR3X1 U5494 ( .IN1(n2438), .IN2(n3570), .IN3(n4932), .Q(n4517) );
  XOR3X1 U5495 ( .IN1(n6065), .IN2(n2802), .IN3(WX7260), .Q(n4932) );
  NAND2X0 U5496 ( .IN1(n4933), .IN2(n3019), .QN(n4930) );
  NAND2X0 U5497 ( .IN1(WX5676), .IN2(n3036), .QN(n4929) );
  NAND2X0 U5498 ( .IN1(n3047), .IN2(CRC_OUT_5_20), .QN(n4928) );
  NAND4X0 U5499 ( .IN1(n4934), .IN2(n4935), .IN3(n4936), .IN4(n4937), .QN(
        WX5836) );
  NAND2X0 U5500 ( .IN1(n4523), .IN2(n3099), .QN(n4937) );
  XOR3X1 U5501 ( .IN1(n2440), .IN2(n3577), .IN3(n4938), .Q(n4523) );
  XOR3X1 U5502 ( .IN1(test_so63), .IN2(n6066), .IN3(WX7258), .Q(n4938) );
  NAND2X0 U5503 ( .IN1(n2998), .IN2(n4939), .QN(n4936) );
  NAND2X0 U5504 ( .IN1(WX5674), .IN2(n3036), .QN(n4935) );
  NAND2X0 U5505 ( .IN1(n3047), .IN2(CRC_OUT_5_21), .QN(n4934) );
  NAND4X0 U5506 ( .IN1(n4940), .IN2(n4941), .IN3(n4942), .IN4(n4943), .QN(
        WX5834) );
  NAND2X0 U5507 ( .IN1(n3080), .IN2(n4529), .QN(n4943) );
  XNOR3X1 U5508 ( .IN1(n2441), .IN2(n3570), .IN3(n4944), .Q(n4529) );
  XOR3X1 U5509 ( .IN1(n6067), .IN2(n2801), .IN3(WX7256), .Q(n4944) );
  NAND2X0 U5510 ( .IN1(n4945), .IN2(n3019), .QN(n4942) );
  NAND2X0 U5511 ( .IN1(WX5672), .IN2(n3036), .QN(n4941) );
  NAND2X0 U5512 ( .IN1(n3047), .IN2(CRC_OUT_5_22), .QN(n4940) );
  NAND4X0 U5513 ( .IN1(n4946), .IN2(n4947), .IN3(n4948), .IN4(n4949), .QN(
        WX5832) );
  NAND2X0 U5514 ( .IN1(n4535), .IN2(n3099), .QN(n4949) );
  XOR3X1 U5515 ( .IN1(n2443), .IN2(n3577), .IN3(n4950), .Q(n4535) );
  XNOR3X1 U5516 ( .IN1(test_so61), .IN2(n6068), .IN3(n2800), .Q(n4950) );
  NAND2X0 U5517 ( .IN1(n2998), .IN2(n4951), .QN(n4948) );
  NAND2X0 U5518 ( .IN1(WX5670), .IN2(n3036), .QN(n4947) );
  NAND2X0 U5519 ( .IN1(n3047), .IN2(CRC_OUT_5_23), .QN(n4946) );
  NAND4X0 U5520 ( .IN1(n4952), .IN2(n4953), .IN3(n4954), .IN4(n4955), .QN(
        WX5830) );
  NAND2X0 U5521 ( .IN1(n3080), .IN2(n4541), .QN(n4955) );
  XNOR3X1 U5522 ( .IN1(n2444), .IN2(n3570), .IN3(n4956), .Q(n4541) );
  XOR3X1 U5523 ( .IN1(n6069), .IN2(n2799), .IN3(WX7252), .Q(n4956) );
  NAND2X0 U5524 ( .IN1(n2998), .IN2(n4957), .QN(n4954) );
  NAND2X0 U5525 ( .IN1(WX5668), .IN2(n3036), .QN(n4953) );
  NAND2X0 U5526 ( .IN1(n3047), .IN2(CRC_OUT_5_24), .QN(n4952) );
  NAND4X0 U5527 ( .IN1(n4958), .IN2(n4959), .IN3(n4960), .IN4(n4961), .QN(
        WX5828) );
  NAND2X0 U5528 ( .IN1(n4547), .IN2(n3100), .QN(n4961) );
  XOR3X1 U5529 ( .IN1(n2446), .IN2(n3579), .IN3(n4962), .Q(n4547) );
  XNOR3X1 U5530 ( .IN1(test_so59), .IN2(n6070), .IN3(n2798), .Q(n4962) );
  NAND2X0 U5531 ( .IN1(n2998), .IN2(n4963), .QN(n4960) );
  NAND2X0 U5532 ( .IN1(WX5666), .IN2(n3036), .QN(n4959) );
  NAND2X0 U5533 ( .IN1(n3048), .IN2(CRC_OUT_5_25), .QN(n4958) );
  NAND4X0 U5534 ( .IN1(n4964), .IN2(n4965), .IN3(n4966), .IN4(n4967), .QN(
        WX5826) );
  NAND2X0 U5535 ( .IN1(n3080), .IN2(n4553), .QN(n4967) );
  XNOR3X1 U5536 ( .IN1(n2447), .IN2(n3570), .IN3(n4968), .Q(n4553) );
  XOR3X1 U5537 ( .IN1(n6071), .IN2(n2797), .IN3(WX7248), .Q(n4968) );
  NAND2X0 U5538 ( .IN1(n2998), .IN2(n4969), .QN(n4966) );
  NAND2X0 U5539 ( .IN1(WX5664), .IN2(n3036), .QN(n4965) );
  NAND2X0 U5540 ( .IN1(n3048), .IN2(CRC_OUT_5_26), .QN(n4964) );
  NAND4X0 U5541 ( .IN1(n4970), .IN2(n4971), .IN3(n4972), .IN4(n4973), .QN(
        WX5824) );
  NAND2X0 U5542 ( .IN1(n4559), .IN2(n3100), .QN(n4973) );
  XOR3X1 U5543 ( .IN1(n2449), .IN2(n3577), .IN3(n4974), .Q(n4559) );
  XNOR3X1 U5544 ( .IN1(test_so57), .IN2(n6072), .IN3(n2796), .Q(n4974) );
  NAND2X0 U5545 ( .IN1(n2998), .IN2(n4975), .QN(n4972) );
  NAND2X0 U5546 ( .IN1(WX5662), .IN2(n3036), .QN(n4971) );
  NAND2X0 U5547 ( .IN1(n3048), .IN2(CRC_OUT_5_27), .QN(n4970) );
  NAND4X0 U5548 ( .IN1(n4976), .IN2(n4977), .IN3(n4978), .IN4(n4979), .QN(
        WX5822) );
  NAND2X0 U5549 ( .IN1(n3080), .IN2(n4565), .QN(n4979) );
  XNOR3X1 U5550 ( .IN1(n2450), .IN2(n3570), .IN3(n4980), .Q(n4565) );
  XOR3X1 U5551 ( .IN1(n6073), .IN2(n2795), .IN3(WX7244), .Q(n4980) );
  NAND2X0 U5552 ( .IN1(n2998), .IN2(n4981), .QN(n4978) );
  NAND2X0 U5553 ( .IN1(WX5660), .IN2(n3037), .QN(n4977) );
  NAND2X0 U5554 ( .IN1(n3048), .IN2(CRC_OUT_5_28), .QN(n4976) );
  NAND4X0 U5555 ( .IN1(n4982), .IN2(n4983), .IN3(n4984), .IN4(n4985), .QN(
        WX5820) );
  NAND2X0 U5556 ( .IN1(n3080), .IN2(n4571), .QN(n4985) );
  XNOR3X1 U5557 ( .IN1(n2452), .IN2(n3570), .IN3(n4986), .Q(n4571) );
  XOR3X1 U5558 ( .IN1(n6074), .IN2(n2794), .IN3(WX7242), .Q(n4986) );
  NAND2X0 U5559 ( .IN1(n2998), .IN2(n4987), .QN(n4984) );
  NAND2X0 U5560 ( .IN1(WX5658), .IN2(n3037), .QN(n4983) );
  NAND2X0 U5561 ( .IN1(n3048), .IN2(CRC_OUT_5_29), .QN(n4982) );
  NAND4X0 U5562 ( .IN1(n4988), .IN2(n4989), .IN3(n4990), .IN4(n4991), .QN(
        WX5818) );
  NAND2X0 U5563 ( .IN1(n3080), .IN2(n4577), .QN(n4991) );
  XNOR3X1 U5564 ( .IN1(n2454), .IN2(n3570), .IN3(n4992), .Q(n4577) );
  XOR3X1 U5565 ( .IN1(n6075), .IN2(n2793), .IN3(WX7240), .Q(n4992) );
  NAND2X0 U5566 ( .IN1(n2998), .IN2(n4993), .QN(n4990) );
  NAND2X0 U5567 ( .IN1(WX5656), .IN2(n3037), .QN(n4989) );
  NAND2X0 U5568 ( .IN1(n3048), .IN2(CRC_OUT_5_30), .QN(n4988) );
  NAND4X0 U5569 ( .IN1(n4994), .IN2(n4995), .IN3(n4996), .IN4(n4997), .QN(
        WX5816) );
  NAND2X0 U5570 ( .IN1(n3081), .IN2(n4583), .QN(n4997) );
  XNOR3X1 U5571 ( .IN1(n2340), .IN2(n3571), .IN3(n4998), .Q(n4583) );
  XOR3X1 U5572 ( .IN1(n6076), .IN2(n2792), .IN3(WX7238), .Q(n4998) );
  NAND2X0 U5573 ( .IN1(n2998), .IN2(n4999), .QN(n4996) );
  NAND2X0 U5574 ( .IN1(n3048), .IN2(CRC_OUT_5_31), .QN(n4995) );
  NAND2X0 U5575 ( .IN1(n2245), .IN2(WX5657), .QN(n4994) );
  NOR2X0 U5576 ( .IN1(n3752), .IN2(WX5657), .QN(WX5718) );
  AND2X1 U5577 ( .IN1(n3619), .IN2(n8496), .Q(WX5716) );
  AND2X1 U5578 ( .IN1(n3619), .IN2(n8497), .Q(WX5714) );
  AND2X1 U5579 ( .IN1(n3619), .IN2(n8498), .Q(WX5712) );
  AND2X1 U5580 ( .IN1(n3619), .IN2(n8499), .Q(WX5710) );
  AND2X1 U5581 ( .IN1(n3619), .IN2(n8500), .Q(WX5708) );
  AND2X1 U5582 ( .IN1(n3619), .IN2(n8501), .Q(WX5706) );
  AND2X1 U5583 ( .IN1(n3619), .IN2(n8502), .Q(WX5704) );
  AND2X1 U5584 ( .IN1(test_so45), .IN2(n3598), .Q(WX5702) );
  AND2X1 U5585 ( .IN1(n3618), .IN2(n8505), .Q(WX5700) );
  AND2X1 U5586 ( .IN1(n3618), .IN2(n8506), .Q(WX5698) );
  AND2X1 U5587 ( .IN1(n3618), .IN2(n8507), .Q(WX5696) );
  AND2X1 U5588 ( .IN1(n3618), .IN2(n8508), .Q(WX5694) );
  AND2X1 U5589 ( .IN1(n3618), .IN2(n8509), .Q(WX5692) );
  AND2X1 U5590 ( .IN1(n3618), .IN2(n8510), .Q(WX5690) );
  AND2X1 U5591 ( .IN1(n3618), .IN2(n8511), .Q(WX5688) );
  AND2X1 U5592 ( .IN1(n3618), .IN2(n8512), .Q(WX5686) );
  AND2X1 U5593 ( .IN1(n3616), .IN2(n8513), .Q(WX5684) );
  AND2X1 U5594 ( .IN1(n3616), .IN2(n8514), .Q(WX5682) );
  AND2X1 U5595 ( .IN1(n3616), .IN2(n8515), .Q(WX5680) );
  AND2X1 U5596 ( .IN1(n3616), .IN2(n8516), .Q(WX5678) );
  AND2X1 U5597 ( .IN1(n3616), .IN2(n8517), .Q(WX5676) );
  AND2X1 U5598 ( .IN1(n3616), .IN2(n8518), .Q(WX5674) );
  AND2X1 U5599 ( .IN1(n3616), .IN2(n8519), .Q(WX5672) );
  AND2X1 U5600 ( .IN1(n3616), .IN2(n8520), .Q(WX5670) );
  AND2X1 U5601 ( .IN1(test_so44), .IN2(n3598), .Q(WX5668) );
  AND2X1 U5602 ( .IN1(n3615), .IN2(n8523), .Q(WX5666) );
  AND2X1 U5603 ( .IN1(n3615), .IN2(n8524), .Q(WX5664) );
  AND2X1 U5604 ( .IN1(n3615), .IN2(n8525), .Q(WX5662) );
  AND2X1 U5605 ( .IN1(n3615), .IN2(n8526), .Q(WX5660) );
  AND2X1 U5606 ( .IN1(n3615), .IN2(n8527), .Q(WX5658) );
  AND2X1 U5607 ( .IN1(n3615), .IN2(n8528), .Q(WX5656) );
  NOR2X0 U5608 ( .IN1(n3752), .IN2(WX485), .QN(WX546) );
  NOR2X0 U5609 ( .IN1(n3752), .IN2(n5000), .QN(WX5205) );
  XOR2X1 U5610 ( .IN1(n2847), .IN2(DFF_766_n1), .Q(n5000) );
  NOR2X0 U5611 ( .IN1(n3752), .IN2(n5001), .QN(WX5203) );
  XOR2X1 U5612 ( .IN1(n2848), .IN2(DFF_765_n1), .Q(n5001) );
  NOR2X0 U5613 ( .IN1(n3753), .IN2(n5002), .QN(WX5201) );
  XOR2X1 U5614 ( .IN1(n2849), .IN2(DFF_764_n1), .Q(n5002) );
  NOR2X0 U5615 ( .IN1(n3753), .IN2(n5003), .QN(WX5199) );
  XOR2X1 U5616 ( .IN1(CRC_OUT_6_27), .IN2(test_so40), .Q(n5003) );
  NOR2X0 U5617 ( .IN1(n3753), .IN2(n5004), .QN(WX5197) );
  XOR2X1 U5618 ( .IN1(n2850), .IN2(DFF_762_n1), .Q(n5004) );
  NOR2X0 U5619 ( .IN1(n3753), .IN2(n5005), .QN(WX5195) );
  XOR2X1 U5620 ( .IN1(n2851), .IN2(DFF_761_n1), .Q(n5005) );
  NOR2X0 U5621 ( .IN1(n3753), .IN2(n5006), .QN(WX5193) );
  XOR2X1 U5622 ( .IN1(n2852), .IN2(DFF_760_n1), .Q(n5006) );
  NOR2X0 U5623 ( .IN1(n3753), .IN2(n5007), .QN(WX5191) );
  XOR2X1 U5624 ( .IN1(n2853), .IN2(DFF_759_n1), .Q(n5007) );
  NOR2X0 U5625 ( .IN1(n3753), .IN2(n5008), .QN(WX5189) );
  XNOR2X1 U5626 ( .IN1(n2854), .IN2(test_so43), .Q(n5008) );
  NOR2X0 U5627 ( .IN1(n3753), .IN2(n5009), .QN(WX5187) );
  XOR2X1 U5628 ( .IN1(n2855), .IN2(DFF_757_n1), .Q(n5009) );
  NOR2X0 U5629 ( .IN1(n3753), .IN2(n5010), .QN(WX5185) );
  XOR2X1 U5630 ( .IN1(n2856), .IN2(DFF_756_n1), .Q(n5010) );
  NOR2X0 U5631 ( .IN1(n3753), .IN2(n5011), .QN(WX5183) );
  XOR2X1 U5632 ( .IN1(n2857), .IN2(DFF_755_n1), .Q(n5011) );
  NOR2X0 U5633 ( .IN1(n3753), .IN2(n5012), .QN(WX5181) );
  XOR2X1 U5634 ( .IN1(n2858), .IN2(DFF_754_n1), .Q(n5012) );
  NOR2X0 U5635 ( .IN1(n3753), .IN2(n5013), .QN(WX5179) );
  XOR2X1 U5636 ( .IN1(n2859), .IN2(DFF_753_n1), .Q(n5013) );
  NOR2X0 U5637 ( .IN1(n3753), .IN2(n5014), .QN(WX5177) );
  XOR2X1 U5638 ( .IN1(n2860), .IN2(DFF_752_n1), .Q(n5014) );
  NOR2X0 U5639 ( .IN1(n3754), .IN2(n5015), .QN(WX5175) );
  XOR3X1 U5640 ( .IN1(n2698), .IN2(DFF_767_n1), .IN3(CRC_OUT_6_15), .Q(n5015)
         );
  NOR2X0 U5641 ( .IN1(n3754), .IN2(n5016), .QN(WX5173) );
  XOR2X1 U5642 ( .IN1(n2861), .IN2(DFF_750_n1), .Q(n5016) );
  NOR2X0 U5643 ( .IN1(n3754), .IN2(n5017), .QN(WX5171) );
  XOR2X1 U5644 ( .IN1(n2862), .IN2(DFF_749_n1), .Q(n5017) );
  NOR2X0 U5645 ( .IN1(n3754), .IN2(n5018), .QN(WX5169) );
  XOR2X1 U5646 ( .IN1(n2863), .IN2(DFF_748_n1), .Q(n5018) );
  NOR2X0 U5647 ( .IN1(n3754), .IN2(n5019), .QN(WX5167) );
  XOR2X1 U5648 ( .IN1(n2864), .IN2(DFF_747_n1), .Q(n5019) );
  NOR2X0 U5649 ( .IN1(n3754), .IN2(n5020), .QN(WX5165) );
  XOR3X1 U5650 ( .IN1(test_so41), .IN2(DFF_767_n1), .IN3(DFF_746_n1), .Q(n5020) );
  NOR2X0 U5651 ( .IN1(n3754), .IN2(n5021), .QN(WX5163) );
  XOR2X1 U5652 ( .IN1(n2865), .IN2(DFF_745_n1), .Q(n5021) );
  NOR2X0 U5653 ( .IN1(n3754), .IN2(n5022), .QN(WX5161) );
  XOR2X1 U5654 ( .IN1(n2866), .IN2(DFF_744_n1), .Q(n5022) );
  NOR2X0 U5655 ( .IN1(n3754), .IN2(n5023), .QN(WX5159) );
  XOR2X1 U5656 ( .IN1(n2867), .IN2(DFF_743_n1), .Q(n5023) );
  NOR2X0 U5657 ( .IN1(n3754), .IN2(n5024), .QN(WX5157) );
  XOR2X1 U5658 ( .IN1(n2868), .IN2(DFF_742_n1), .Q(n5024) );
  NOR2X0 U5659 ( .IN1(n3754), .IN2(n5025), .QN(WX5155) );
  XNOR2X1 U5660 ( .IN1(n2869), .IN2(test_so42), .Q(n5025) );
  NOR2X0 U5661 ( .IN1(n3754), .IN2(n5026), .QN(WX5153) );
  XOR2X1 U5662 ( .IN1(n2870), .IN2(DFF_740_n1), .Q(n5026) );
  NOR2X0 U5663 ( .IN1(n3754), .IN2(n5027), .QN(WX5151) );
  XOR3X1 U5664 ( .IN1(n2699), .IN2(DFF_767_n1), .IN3(CRC_OUT_6_3), .Q(n5027)
         );
  NOR2X0 U5665 ( .IN1(n3755), .IN2(n5028), .QN(WX5149) );
  XOR2X1 U5666 ( .IN1(n2871), .IN2(DFF_738_n1), .Q(n5028) );
  NOR2X0 U5667 ( .IN1(n3755), .IN2(n5029), .QN(WX5147) );
  XOR2X1 U5668 ( .IN1(n2872), .IN2(DFF_737_n1), .Q(n5029) );
  NOR2X0 U5669 ( .IN1(n3755), .IN2(n5030), .QN(WX5145) );
  XOR2X1 U5670 ( .IN1(n2873), .IN2(DFF_736_n1), .Q(n5030) );
  NOR2X0 U5671 ( .IN1(n3755), .IN2(n5031), .QN(WX5143) );
  XOR2X1 U5672 ( .IN1(n2711), .IN2(DFF_767_n1), .Q(n5031) );
  NOR2X0 U5673 ( .IN1(n6118), .IN2(n3729), .QN(WX4617) );
  AND2X1 U5674 ( .IN1(n3615), .IN2(test_so35), .Q(WX4615) );
  NOR2X0 U5675 ( .IN1(n6120), .IN2(n3662), .QN(WX4613) );
  NOR2X0 U5676 ( .IN1(n6121), .IN2(n3662), .QN(WX4611) );
  NOR2X0 U5677 ( .IN1(n6122), .IN2(n3662), .QN(WX4609) );
  NOR2X0 U5678 ( .IN1(n6123), .IN2(n3662), .QN(WX4607) );
  NOR2X0 U5679 ( .IN1(n6124), .IN2(n3662), .QN(WX4605) );
  NOR2X0 U5680 ( .IN1(n6125), .IN2(n3662), .QN(WX4603) );
  NOR2X0 U5681 ( .IN1(n6126), .IN2(n3662), .QN(WX4601) );
  NOR2X0 U5682 ( .IN1(n6127), .IN2(n3662), .QN(WX4599) );
  NOR2X0 U5683 ( .IN1(n6128), .IN2(n3662), .QN(WX4597) );
  NOR2X0 U5684 ( .IN1(n6129), .IN2(n3662), .QN(WX4595) );
  NOR2X0 U5685 ( .IN1(n6130), .IN2(n3662), .QN(WX4593) );
  NOR2X0 U5686 ( .IN1(n6131), .IN2(n3662), .QN(WX4591) );
  NOR2X0 U5687 ( .IN1(n6132), .IN2(n3660), .QN(WX4589) );
  NOR2X0 U5688 ( .IN1(n6133), .IN2(n3660), .QN(WX4587) );
  NAND4X0 U5689 ( .IN1(n5032), .IN2(n5033), .IN3(n5034), .IN4(n5035), .QN(
        WX4585) );
  NAND2X0 U5690 ( .IN1(n3081), .IN2(n4813), .QN(n5035) );
  XNOR3X1 U5691 ( .IN1(n2710), .IN2(n2619), .IN3(n5036), .Q(n4813) );
  XOR2X1 U5692 ( .IN1(WX5943), .IN2(n6077), .Q(n5036) );
  NAND2X0 U5693 ( .IN1(n5037), .IN2(n3021), .QN(n5034) );
  NAND2X0 U5694 ( .IN1(WX4423), .IN2(n3037), .QN(n5033) );
  NAND2X0 U5695 ( .IN1(n3048), .IN2(CRC_OUT_6_0), .QN(n5032) );
  NAND4X0 U5696 ( .IN1(n5038), .IN2(n5039), .IN3(n5040), .IN4(n5041), .QN(
        WX4583) );
  NAND2X0 U5697 ( .IN1(n4819), .IN2(n3100), .QN(n5041) );
  XOR3X1 U5698 ( .IN1(n3661), .IN2(n2846), .IN3(n5042), .Q(n4819) );
  XOR2X1 U5699 ( .IN1(WX5877), .IN2(test_so51), .Q(n5042) );
  NAND2X0 U5700 ( .IN1(n3003), .IN2(n5043), .QN(n5040) );
  NAND2X0 U5701 ( .IN1(WX4421), .IN2(n3037), .QN(n5039) );
  NAND2X0 U5702 ( .IN1(n3048), .IN2(CRC_OUT_6_1), .QN(n5038) );
  NAND4X0 U5703 ( .IN1(n5044), .IN2(n5045), .IN3(n5046), .IN4(n5047), .QN(
        WX4581) );
  NAND2X0 U5704 ( .IN1(n3081), .IN2(n4825), .QN(n5047) );
  XNOR3X1 U5705 ( .IN1(n2845), .IN2(n2620), .IN3(n5048), .Q(n4825) );
  XOR2X1 U5706 ( .IN1(WX5939), .IN2(n6078), .Q(n5048) );
  NAND2X0 U5707 ( .IN1(n3013), .IN2(n5049), .QN(n5046) );
  NAND2X0 U5708 ( .IN1(WX4419), .IN2(n3037), .QN(n5045) );
  NAND2X0 U5709 ( .IN1(n3048), .IN2(CRC_OUT_6_2), .QN(n5044) );
  NAND4X0 U5710 ( .IN1(n5050), .IN2(n5051), .IN3(n5052), .IN4(n5053), .QN(
        WX4579) );
  NAND2X0 U5711 ( .IN1(n4831), .IN2(n3100), .QN(n5053) );
  XOR3X1 U5712 ( .IN1(n2844), .IN2(n2621), .IN3(n5054), .Q(n4831) );
  XOR2X1 U5713 ( .IN1(WX5873), .IN2(test_so49), .Q(n5054) );
  NAND2X0 U5714 ( .IN1(n3013), .IN2(n5055), .QN(n5052) );
  NAND2X0 U5715 ( .IN1(WX4417), .IN2(n3037), .QN(n5051) );
  NAND2X0 U6483 ( .IN1(n3048), .IN2(CRC_OUT_6_3), .QN(n5050) );
  NAND4X0 U6484 ( .IN1(n5056), .IN2(n5057), .IN3(n5058), .IN4(n5059), .QN(
        WX4577) );
  NAND2X0 U6485 ( .IN1(n3081), .IN2(n4837), .QN(n5059) );
  XNOR3X1 U6486 ( .IN1(n2697), .IN2(n2622), .IN3(n5060), .Q(n4837) );
  XOR2X1 U6487 ( .IN1(WX5935), .IN2(n6079), .Q(n5060) );
  NAND2X0 U6488 ( .IN1(n3013), .IN2(n5061), .QN(n5058) );
  NAND2X0 U6489 ( .IN1(WX4415), .IN2(n3037), .QN(n5057) );
  NAND2X0 U6490 ( .IN1(n3048), .IN2(CRC_OUT_6_4), .QN(n5056) );
  NAND4X0 U6491 ( .IN1(n5062), .IN2(n5063), .IN3(n5064), .IN4(n5065), .QN(
        WX4575) );
  NAND2X0 U6492 ( .IN1(n4843), .IN2(n3094), .QN(n5065) );
  XOR3X1 U6493 ( .IN1(n3669), .IN2(n2843), .IN3(n5066), .Q(n4843) );
  XOR2X1 U6494 ( .IN1(WX5997), .IN2(test_so47), .Q(n5066) );
  NAND2X0 U6495 ( .IN1(n3013), .IN2(n5067), .QN(n5064) );
  NAND2X0 U6496 ( .IN1(WX4413), .IN2(n3037), .QN(n5063) );
  NAND2X0 U6497 ( .IN1(test_so42), .IN2(n3070), .QN(n5062) );
  NAND4X0 U6498 ( .IN1(n5068), .IN2(n5069), .IN3(n5070), .IN4(n5071), .QN(
        WX4573) );
  NAND2X0 U6499 ( .IN1(n3081), .IN2(n4849), .QN(n5071) );
  XNOR3X1 U6500 ( .IN1(n2842), .IN2(n2623), .IN3(n5072), .Q(n4849) );
  XOR2X1 U6501 ( .IN1(WX5931), .IN2(n6080), .Q(n5072) );
  NAND2X0 U6502 ( .IN1(n3013), .IN2(n5073), .QN(n5070) );
  NAND2X0 U6503 ( .IN1(WX4411), .IN2(n3037), .QN(n5069) );
  NAND2X0 U6504 ( .IN1(n3049), .IN2(CRC_OUT_6_6), .QN(n5068) );
  NAND4X0 U6505 ( .IN1(n5074), .IN2(n5075), .IN3(n5076), .IN4(n5077), .QN(
        WX4571) );
  NAND2X0 U6506 ( .IN1(n3081), .IN2(n4855), .QN(n5077) );
  XNOR3X1 U6507 ( .IN1(n2841), .IN2(n2624), .IN3(n5078), .Q(n4855) );
  XOR2X1 U6508 ( .IN1(WX5929), .IN2(n6081), .Q(n5078) );
  NAND2X0 U6509 ( .IN1(n3013), .IN2(n5079), .QN(n5076) );
  NAND2X0 U6510 ( .IN1(WX4409), .IN2(n3037), .QN(n5075) );
  NAND2X0 U6511 ( .IN1(n3049), .IN2(CRC_OUT_6_7), .QN(n5074) );
  NAND4X0 U6512 ( .IN1(n5080), .IN2(n5081), .IN3(n5082), .IN4(n5083), .QN(
        WX4569) );
  NAND2X0 U6513 ( .IN1(n3081), .IN2(n4861), .QN(n5083) );
  XNOR3X1 U6514 ( .IN1(n2840), .IN2(n2625), .IN3(n5084), .Q(n4861) );
  XOR2X1 U6515 ( .IN1(WX5927), .IN2(n6082), .Q(n5084) );
  NAND2X0 U6516 ( .IN1(n3015), .IN2(n5085), .QN(n5082) );
  NAND2X0 U6517 ( .IN1(WX4407), .IN2(n3037), .QN(n5081) );
  NAND2X0 U6518 ( .IN1(n3049), .IN2(CRC_OUT_6_8), .QN(n5080) );
  NAND4X0 U6519 ( .IN1(n5086), .IN2(n5087), .IN3(n5088), .IN4(n5089), .QN(
        WX4567) );
  NAND2X0 U6520 ( .IN1(n3081), .IN2(n4867), .QN(n5089) );
  XNOR3X1 U6521 ( .IN1(n2839), .IN2(n2626), .IN3(n5090), .Q(n4867) );
  XOR2X1 U6522 ( .IN1(WX5925), .IN2(n6083), .Q(n5090) );
  NAND2X0 U6523 ( .IN1(n3014), .IN2(n5091), .QN(n5088) );
  NAND2X0 U6524 ( .IN1(WX4405), .IN2(n3037), .QN(n5087) );
  NAND2X0 U6525 ( .IN1(n3049), .IN2(CRC_OUT_6_9), .QN(n5086) );
  NAND4X0 U6526 ( .IN1(n5092), .IN2(n5093), .IN3(n5094), .IN4(n5095), .QN(
        WX4565) );
  NAND2X0 U6527 ( .IN1(n3081), .IN2(n4873), .QN(n5095) );
  XNOR3X1 U6528 ( .IN1(n2838), .IN2(n2627), .IN3(n5096), .Q(n4873) );
  XOR2X1 U6529 ( .IN1(WX5923), .IN2(n6084), .Q(n5096) );
  NAND2X0 U6530 ( .IN1(n3014), .IN2(n5097), .QN(n5094) );
  NAND2X0 U6531 ( .IN1(WX4403), .IN2(n3037), .QN(n5093) );
  NAND2X0 U6532 ( .IN1(n3049), .IN2(CRC_OUT_6_10), .QN(n5092) );
  NAND4X0 U6533 ( .IN1(n5098), .IN2(n5099), .IN3(n5100), .IN4(n5101), .QN(
        WX4563) );
  NAND2X0 U6534 ( .IN1(n3081), .IN2(n4879), .QN(n5101) );
  XNOR3X1 U6535 ( .IN1(n2696), .IN2(n2628), .IN3(n5102), .Q(n4879) );
  XOR2X1 U6536 ( .IN1(WX5921), .IN2(n6085), .Q(n5102) );
  NAND2X0 U6537 ( .IN1(n5103), .IN2(n3019), .QN(n5100) );
  NAND2X0 U6538 ( .IN1(WX4401), .IN2(n3037), .QN(n5099) );
  NAND2X0 U6539 ( .IN1(n3049), .IN2(CRC_OUT_6_11), .QN(n5098) );
  NAND4X0 U6540 ( .IN1(n5104), .IN2(n5105), .IN3(n5106), .IN4(n5107), .QN(
        WX4561) );
  NAND2X0 U6541 ( .IN1(n3081), .IN2(n4885), .QN(n5107) );
  XNOR3X1 U6542 ( .IN1(n2837), .IN2(n2629), .IN3(n5108), .Q(n4885) );
  XOR2X1 U6543 ( .IN1(WX5919), .IN2(n6086), .Q(n5108) );
  NAND2X0 U6544 ( .IN1(n3014), .IN2(n5109), .QN(n5106) );
  NAND2X0 U6545 ( .IN1(WX4399), .IN2(n3037), .QN(n5105) );
  NAND2X0 U6546 ( .IN1(n3049), .IN2(CRC_OUT_6_12), .QN(n5104) );
  NAND4X0 U6547 ( .IN1(n5110), .IN2(n5111), .IN3(n5112), .IN4(n5113), .QN(
        WX4559) );
  NAND2X0 U6548 ( .IN1(n3081), .IN2(n4891), .QN(n5113) );
  XNOR3X1 U6549 ( .IN1(n2836), .IN2(n2630), .IN3(n5114), .Q(n4891) );
  XOR2X1 U6550 ( .IN1(WX5917), .IN2(n6087), .Q(n5114) );
  NAND2X0 U6551 ( .IN1(n5115), .IN2(n3019), .QN(n5112) );
  NAND2X0 U6552 ( .IN1(WX4397), .IN2(n3037), .QN(n5111) );
  NAND2X0 U6553 ( .IN1(n3049), .IN2(CRC_OUT_6_13), .QN(n5110) );
  NAND4X0 U6554 ( .IN1(n5116), .IN2(n5117), .IN3(n5118), .IN4(n5119), .QN(
        WX4557) );
  NAND2X0 U6555 ( .IN1(n3082), .IN2(n4897), .QN(n5119) );
  XNOR3X1 U6556 ( .IN1(n2835), .IN2(n2631), .IN3(n5120), .Q(n4897) );
  XOR2X1 U6557 ( .IN1(WX5915), .IN2(n6088), .Q(n5120) );
  NAND2X0 U6558 ( .IN1(n3014), .IN2(n5121), .QN(n5118) );
  NAND2X0 U6559 ( .IN1(WX4395), .IN2(n3038), .QN(n5117) );
  NAND2X0 U6560 ( .IN1(n3049), .IN2(CRC_OUT_6_14), .QN(n5116) );
  NAND4X0 U6561 ( .IN1(n5122), .IN2(n5123), .IN3(n5124), .IN4(n5125), .QN(
        WX4555) );
  NAND2X0 U6562 ( .IN1(n3082), .IN2(n4903), .QN(n5125) );
  XNOR3X1 U6563 ( .IN1(n2834), .IN2(n2632), .IN3(n5126), .Q(n4903) );
  XOR2X1 U6564 ( .IN1(WX5913), .IN2(n6089), .Q(n5126) );
  NAND2X0 U6565 ( .IN1(n5127), .IN2(n3019), .QN(n5124) );
  NAND2X0 U6566 ( .IN1(WX4393), .IN2(n3038), .QN(n5123) );
  NAND2X0 U6567 ( .IN1(n3049), .IN2(CRC_OUT_6_15), .QN(n5122) );
  NAND4X0 U6568 ( .IN1(n5128), .IN2(n5129), .IN3(n5130), .IN4(n5131), .QN(
        WX4553) );
  NAND2X0 U6569 ( .IN1(n4909), .IN2(n3100), .QN(n5131) );
  XOR3X1 U6570 ( .IN1(n2456), .IN2(n3578), .IN3(n5132), .Q(n4909) );
  XOR3X1 U6571 ( .IN1(test_so52), .IN2(n6090), .IN3(WX5975), .Q(n5132) );
  NAND2X0 U6572 ( .IN1(n3014), .IN2(n5133), .QN(n5130) );
  NAND2X0 U6573 ( .IN1(WX4391), .IN2(n3038), .QN(n5129) );
  NAND2X0 U6574 ( .IN1(n3049), .IN2(CRC_OUT_6_16), .QN(n5128) );
  NAND4X0 U6575 ( .IN1(n5134), .IN2(n5135), .IN3(n5136), .IN4(n5137), .QN(
        WX4551) );
  NAND2X0 U6576 ( .IN1(n3082), .IN2(n4915), .QN(n5137) );
  XNOR3X1 U6577 ( .IN1(n2457), .IN2(n3571), .IN3(n5138), .Q(n4915) );
  XOR3X1 U6578 ( .IN1(n6091), .IN2(n2833), .IN3(WX5973), .Q(n5138) );
  NAND2X0 U6579 ( .IN1(n5139), .IN2(n3019), .QN(n5136) );
  NAND2X0 U6580 ( .IN1(WX4389), .IN2(n3038), .QN(n5135) );
  NAND2X0 U6581 ( .IN1(n3049), .IN2(CRC_OUT_6_17), .QN(n5134) );
  NAND4X0 U6582 ( .IN1(n5140), .IN2(n5141), .IN3(n5142), .IN4(n5143), .QN(
        WX4549) );
  NAND2X0 U6583 ( .IN1(n4921), .IN2(n3100), .QN(n5143) );
  XOR3X1 U6584 ( .IN1(n2459), .IN2(n3578), .IN3(n5144), .Q(n4921) );
  XNOR3X1 U6585 ( .IN1(test_so50), .IN2(n6092), .IN3(n2832), .Q(n5144) );
  NAND2X0 U6586 ( .IN1(n3014), .IN2(n5145), .QN(n5142) );
  NAND2X0 U6587 ( .IN1(WX4387), .IN2(n3038), .QN(n5141) );
  NAND2X0 U6588 ( .IN1(n3050), .IN2(CRC_OUT_6_18), .QN(n5140) );
  NAND4X0 U6589 ( .IN1(n5146), .IN2(n5147), .IN3(n5148), .IN4(n5149), .QN(
        WX4547) );
  NAND2X0 U6590 ( .IN1(n3082), .IN2(n4927), .QN(n5149) );
  XNOR3X1 U6591 ( .IN1(n2460), .IN2(n3571), .IN3(n5150), .Q(n4927) );
  XOR3X1 U6592 ( .IN1(n6093), .IN2(n2831), .IN3(WX5969), .Q(n5150) );
  NAND2X0 U6593 ( .IN1(n3014), .IN2(n5151), .QN(n5148) );
  NAND2X0 U6594 ( .IN1(WX4385), .IN2(n3038), .QN(n5147) );
  NAND2X0 U6595 ( .IN1(n3050), .IN2(CRC_OUT_6_19), .QN(n5146) );
  NAND4X0 U6596 ( .IN1(n5152), .IN2(n5153), .IN3(n5154), .IN4(n5155), .QN(
        WX4545) );
  NAND2X0 U6597 ( .IN1(n4933), .IN2(n3100), .QN(n5155) );
  XOR3X1 U6598 ( .IN1(n2462), .IN2(n3577), .IN3(n5156), .Q(n4933) );
  XNOR3X1 U6599 ( .IN1(test_so48), .IN2(n6094), .IN3(n2830), .Q(n5156) );
  NAND2X0 U6600 ( .IN1(n3014), .IN2(n5157), .QN(n5154) );
  NAND2X0 U6601 ( .IN1(WX4383), .IN2(n3038), .QN(n5153) );
  NAND2X0 U6602 ( .IN1(n3050), .IN2(CRC_OUT_6_20), .QN(n5152) );
  NAND4X0 U6603 ( .IN1(n5158), .IN2(n5159), .IN3(n5160), .IN4(n5161), .QN(
        WX4543) );
  NAND2X0 U6604 ( .IN1(n3082), .IN2(n4939), .QN(n5161) );
  XNOR3X1 U6605 ( .IN1(n2463), .IN2(n3571), .IN3(n5162), .Q(n4939) );
  XOR3X1 U6606 ( .IN1(n6095), .IN2(n2829), .IN3(WX5965), .Q(n5162) );
  NAND2X0 U6607 ( .IN1(n3014), .IN2(n5163), .QN(n5160) );
  NAND2X0 U6608 ( .IN1(WX4381), .IN2(n3038), .QN(n5159) );
  NAND2X0 U6609 ( .IN1(n3050), .IN2(CRC_OUT_6_21), .QN(n5158) );
  NAND4X0 U6610 ( .IN1(n5164), .IN2(n5165), .IN3(n5166), .IN4(n5167), .QN(
        WX4541) );
  NAND2X0 U6611 ( .IN1(n4945), .IN2(n3100), .QN(n5167) );
  XOR3X1 U6612 ( .IN1(n2465), .IN2(n3577), .IN3(n5168), .Q(n4945) );
  XNOR3X1 U6613 ( .IN1(test_so46), .IN2(n6096), .IN3(n2828), .Q(n5168) );
  NAND2X0 U6614 ( .IN1(n3014), .IN2(n5169), .QN(n5166) );
  NAND2X0 U6615 ( .IN1(WX4379), .IN2(n3038), .QN(n5165) );
  NAND2X0 U6616 ( .IN1(test_so43), .IN2(n3069), .QN(n5164) );
  NAND4X0 U6617 ( .IN1(n5170), .IN2(n5171), .IN3(n5172), .IN4(n5173), .QN(
        WX4539) );
  NAND2X0 U6618 ( .IN1(n3082), .IN2(n4951), .QN(n5173) );
  XNOR3X1 U6619 ( .IN1(n2466), .IN2(n3571), .IN3(n5174), .Q(n4951) );
  XOR3X1 U6620 ( .IN1(n6097), .IN2(n2827), .IN3(WX5961), .Q(n5174) );
  NAND2X0 U6621 ( .IN1(n3014), .IN2(n5175), .QN(n5172) );
  NAND2X0 U6622 ( .IN1(WX4377), .IN2(n3038), .QN(n5171) );
  NAND2X0 U6623 ( .IN1(n3050), .IN2(CRC_OUT_6_23), .QN(n5170) );
  NAND4X0 U6624 ( .IN1(n5176), .IN2(n5177), .IN3(n5178), .IN4(n5179), .QN(
        WX4537) );
  NAND2X0 U6625 ( .IN1(n3082), .IN2(n4957), .QN(n5179) );
  XNOR3X1 U6626 ( .IN1(n2468), .IN2(n3571), .IN3(n5180), .Q(n4957) );
  XOR3X1 U6627 ( .IN1(n6098), .IN2(n2826), .IN3(WX5959), .Q(n5180) );
  NAND2X0 U6628 ( .IN1(n3014), .IN2(n5181), .QN(n5178) );
  NAND2X0 U6629 ( .IN1(WX4375), .IN2(n3038), .QN(n5177) );
  NAND2X0 U6630 ( .IN1(n3050), .IN2(CRC_OUT_6_24), .QN(n5176) );
  NAND4X0 U6631 ( .IN1(n5182), .IN2(n5183), .IN3(n5184), .IN4(n5185), .QN(
        WX4535) );
  NAND2X0 U6632 ( .IN1(n3082), .IN2(n4963), .QN(n5185) );
  XNOR3X1 U6633 ( .IN1(n2470), .IN2(n3571), .IN3(n5186), .Q(n4963) );
  XOR3X1 U6634 ( .IN1(n6099), .IN2(n2825), .IN3(WX5957), .Q(n5186) );
  NAND2X0 U6635 ( .IN1(n3015), .IN2(n5187), .QN(n5184) );
  NAND2X0 U6636 ( .IN1(WX4373), .IN2(n3038), .QN(n5183) );
  NAND2X0 U6637 ( .IN1(n3050), .IN2(CRC_OUT_6_25), .QN(n5182) );
  NAND4X0 U6638 ( .IN1(n5188), .IN2(n5189), .IN3(n5190), .IN4(n5191), .QN(
        WX4533) );
  NAND2X0 U6639 ( .IN1(n3082), .IN2(n4969), .QN(n5191) );
  XNOR3X1 U6640 ( .IN1(n2472), .IN2(n3571), .IN3(n5192), .Q(n4969) );
  XOR3X1 U6641 ( .IN1(n6100), .IN2(n2824), .IN3(WX5955), .Q(n5192) );
  NAND2X0 U6642 ( .IN1(n3015), .IN2(n5193), .QN(n5190) );
  NAND2X0 U6643 ( .IN1(WX4371), .IN2(n3038), .QN(n5189) );
  NAND2X0 U6644 ( .IN1(n3050), .IN2(CRC_OUT_6_26), .QN(n5188) );
  NAND4X0 U6645 ( .IN1(n5194), .IN2(n5195), .IN3(n5196), .IN4(n5197), .QN(
        WX4531) );
  NAND2X0 U6646 ( .IN1(n3082), .IN2(n4975), .QN(n5197) );
  XNOR3X1 U6647 ( .IN1(n2474), .IN2(n3571), .IN3(n5198), .Q(n4975) );
  XOR3X1 U6648 ( .IN1(n6101), .IN2(n2823), .IN3(WX5953), .Q(n5198) );
  NAND2X0 U6649 ( .IN1(n3015), .IN2(n5199), .QN(n5196) );
  NAND2X0 U6650 ( .IN1(WX4369), .IN2(n3038), .QN(n5195) );
  NAND2X0 U6651 ( .IN1(n3050), .IN2(CRC_OUT_6_27), .QN(n5194) );
  NAND4X0 U6652 ( .IN1(n5200), .IN2(n5201), .IN3(n5202), .IN4(n5203), .QN(
        WX4529) );
  NAND2X0 U6653 ( .IN1(n3082), .IN2(n4981), .QN(n5203) );
  XNOR3X1 U6654 ( .IN1(n2476), .IN2(n3571), .IN3(n5204), .Q(n4981) );
  XOR3X1 U6655 ( .IN1(n6102), .IN2(n2822), .IN3(WX5951), .Q(n5204) );
  NAND2X0 U6656 ( .IN1(n5205), .IN2(n3018), .QN(n5202) );
  NAND2X0 U6657 ( .IN1(WX4367), .IN2(n3038), .QN(n5201) );
  NAND2X0 U6658 ( .IN1(n3050), .IN2(CRC_OUT_6_28), .QN(n5200) );
  NAND4X0 U6659 ( .IN1(n5206), .IN2(n5207), .IN3(n5208), .IN4(n5209), .QN(
        WX4527) );
  NAND2X0 U6660 ( .IN1(n3083), .IN2(n4987), .QN(n5209) );
  XNOR3X1 U6661 ( .IN1(n2478), .IN2(n3571), .IN3(n5210), .Q(n4987) );
  XOR3X1 U6662 ( .IN1(n6103), .IN2(n2821), .IN3(WX5949), .Q(n5210) );
  NAND2X0 U6663 ( .IN1(n3015), .IN2(n5211), .QN(n5208) );
  NAND2X0 U6664 ( .IN1(WX4365), .IN2(n3038), .QN(n5207) );
  NAND2X0 U6665 ( .IN1(n3050), .IN2(CRC_OUT_6_29), .QN(n5206) );
  NAND4X0 U6666 ( .IN1(n5212), .IN2(n5213), .IN3(n5214), .IN4(n5215), .QN(
        WX4525) );
  NAND2X0 U6667 ( .IN1(n3083), .IN2(n4993), .QN(n5215) );
  XNOR3X1 U6668 ( .IN1(n2480), .IN2(n3571), .IN3(n5216), .Q(n4993) );
  XOR3X1 U6669 ( .IN1(n6104), .IN2(n2820), .IN3(WX5947), .Q(n5216) );
  NAND2X0 U6670 ( .IN1(n5217), .IN2(n3017), .QN(n5214) );
  NAND2X0 U6671 ( .IN1(WX4363), .IN2(n3038), .QN(n5213) );
  NAND2X0 U6672 ( .IN1(n3050), .IN2(CRC_OUT_6_30), .QN(n5212) );
  NAND4X0 U6673 ( .IN1(n5218), .IN2(n5219), .IN3(n5220), .IN4(n5221), .QN(
        WX4523) );
  NAND2X0 U6674 ( .IN1(n3083), .IN2(n4999), .QN(n5221) );
  XNOR3X1 U6675 ( .IN1(n2342), .IN2(n3572), .IN3(n5222), .Q(n4999) );
  XOR3X1 U6676 ( .IN1(n6105), .IN2(n2819), .IN3(WX5945), .Q(n5222) );
  NAND2X0 U6677 ( .IN1(n3015), .IN2(n5223), .QN(n5220) );
  NAND2X0 U6678 ( .IN1(n3051), .IN2(CRC_OUT_6_31), .QN(n5219) );
  NAND2X0 U6679 ( .IN1(n2245), .IN2(WX4364), .QN(n5218) );
  NOR2X0 U6680 ( .IN1(n3755), .IN2(WX4364), .QN(WX4425) );
  AND2X1 U6681 ( .IN1(n3615), .IN2(n8554), .Q(WX4423) );
  AND2X1 U6682 ( .IN1(n3615), .IN2(n8555), .Q(WX4421) );
  AND2X1 U6683 ( .IN1(test_so34), .IN2(n3598), .Q(WX4419) );
  AND2X1 U6684 ( .IN1(n3614), .IN2(n8558), .Q(WX4417) );
  AND2X1 U6685 ( .IN1(n3614), .IN2(n8559), .Q(WX4415) );
  AND2X1 U6686 ( .IN1(n3614), .IN2(n8560), .Q(WX4413) );
  AND2X1 U6687 ( .IN1(n3614), .IN2(n8561), .Q(WX4411) );
  AND2X1 U6688 ( .IN1(n3614), .IN2(n8562), .Q(WX4409) );
  AND2X1 U6689 ( .IN1(n3614), .IN2(n8563), .Q(WX4407) );
  AND2X1 U6690 ( .IN1(n3614), .IN2(n8564), .Q(WX4405) );
  AND2X1 U6691 ( .IN1(n3614), .IN2(n8565), .Q(WX4403) );
  AND2X1 U6692 ( .IN1(n3612), .IN2(n8566), .Q(WX4401) );
  AND2X1 U6693 ( .IN1(n3612), .IN2(n8567), .Q(WX4399) );
  AND2X1 U6694 ( .IN1(n3612), .IN2(n8568), .Q(WX4397) );
  AND2X1 U6695 ( .IN1(n3621), .IN2(n8569), .Q(WX4395) );
  AND2X1 U6696 ( .IN1(n3599), .IN2(n8570), .Q(WX4393) );
  AND2X1 U6697 ( .IN1(n3614), .IN2(n8571), .Q(WX4391) );
  AND2X1 U6698 ( .IN1(n3616), .IN2(n8572), .Q(WX4389) );
  AND2X1 U6699 ( .IN1(n3618), .IN2(n8573), .Q(WX4387) );
  AND2X1 U6700 ( .IN1(test_so33), .IN2(n3599), .Q(WX4385) );
  AND2X1 U6701 ( .IN1(n3621), .IN2(n8576), .Q(WX4383) );
  AND2X1 U6702 ( .IN1(n3624), .IN2(n8577), .Q(WX4381) );
  AND2X1 U6703 ( .IN1(n3627), .IN2(n8578), .Q(WX4379) );
  AND2X1 U6704 ( .IN1(n3628), .IN2(n8579), .Q(WX4377) );
  AND2X1 U6705 ( .IN1(n3600), .IN2(n8580), .Q(WX4375) );
  AND2X1 U6706 ( .IN1(n3601), .IN2(n8581), .Q(WX4373) );
  AND2X1 U6707 ( .IN1(n3602), .IN2(n8582), .Q(WX4371) );
  AND2X1 U6708 ( .IN1(n3603), .IN2(n8583), .Q(WX4369) );
  AND2X1 U6709 ( .IN1(n3602), .IN2(n8584), .Q(WX4367) );
  AND2X1 U6710 ( .IN1(n3601), .IN2(n8585), .Q(WX4365) );
  AND2X1 U6711 ( .IN1(n3602), .IN2(n8586), .Q(WX4363) );
  NOR2X0 U6712 ( .IN1(n3755), .IN2(n5224), .QN(WX3912) );
  XOR2X1 U6713 ( .IN1(n2874), .IN2(DFF_574_n1), .Q(n5224) );
  NOR2X0 U6714 ( .IN1(n3755), .IN2(n5225), .QN(WX3910) );
  XOR2X1 U6715 ( .IN1(n2875), .IN2(DFF_573_n1), .Q(n5225) );
  NOR2X0 U6716 ( .IN1(n3755), .IN2(n5226), .QN(WX3908) );
  XOR2X1 U6717 ( .IN1(n2876), .IN2(DFF_572_n1), .Q(n5226) );
  NOR2X0 U6718 ( .IN1(n3755), .IN2(n5227), .QN(WX3906) );
  XNOR2X1 U6719 ( .IN1(n2877), .IN2(test_so32), .Q(n5227) );
  NOR2X0 U6720 ( .IN1(n3755), .IN2(n5228), .QN(WX3904) );
  XOR2X1 U6721 ( .IN1(n2878), .IN2(DFF_570_n1), .Q(n5228) );
  NOR2X0 U6722 ( .IN1(n3755), .IN2(n5229), .QN(WX3902) );
  XOR2X1 U6723 ( .IN1(n2879), .IN2(DFF_569_n1), .Q(n5229) );
  NOR2X0 U6724 ( .IN1(n3755), .IN2(n5230), .QN(WX3900) );
  XOR2X1 U6725 ( .IN1(n2880), .IN2(DFF_568_n1), .Q(n5230) );
  NOR2X0 U6726 ( .IN1(n3755), .IN2(n5231), .QN(WX3898) );
  XOR2X1 U6727 ( .IN1(n2881), .IN2(DFF_567_n1), .Q(n5231) );
  NOR2X0 U6728 ( .IN1(n3756), .IN2(n5232), .QN(WX3896) );
  XOR2X1 U6729 ( .IN1(CRC_OUT_7_22), .IN2(test_so29), .Q(n5232) );
  NOR2X0 U6730 ( .IN1(n3756), .IN2(n5233), .QN(WX3894) );
  XOR2X1 U6731 ( .IN1(n2882), .IN2(DFF_565_n1), .Q(n5233) );
  NOR2X0 U6732 ( .IN1(n3756), .IN2(n5234), .QN(WX3892) );
  XOR2X1 U6733 ( .IN1(n2883), .IN2(DFF_564_n1), .Q(n5234) );
  NOR2X0 U6734 ( .IN1(n3756), .IN2(n5235), .QN(WX3890) );
  XOR2X1 U6735 ( .IN1(n2884), .IN2(DFF_563_n1), .Q(n5235) );
  NOR2X0 U6736 ( .IN1(n3756), .IN2(n5236), .QN(WX3888) );
  XOR2X1 U6737 ( .IN1(n2885), .IN2(DFF_562_n1), .Q(n5236) );
  NOR2X0 U6738 ( .IN1(n3756), .IN2(n5237), .QN(WX3886) );
  XOR2X1 U6739 ( .IN1(n2886), .IN2(DFF_561_n1), .Q(n5237) );
  NOR2X0 U6740 ( .IN1(n3756), .IN2(n5238), .QN(WX3884) );
  XOR2X1 U6741 ( .IN1(n2887), .IN2(DFF_560_n1), .Q(n5238) );
  NOR2X0 U6742 ( .IN1(n3756), .IN2(n5239), .QN(WX3882) );
  XOR3X1 U6743 ( .IN1(n2700), .IN2(DFF_575_n1), .IN3(CRC_OUT_7_15), .Q(n5239)
         );
  NOR2X0 U6744 ( .IN1(n3756), .IN2(n5240), .QN(WX3880) );
  XOR2X1 U6745 ( .IN1(n2888), .IN2(DFF_558_n1), .Q(n5240) );
  NOR2X0 U6746 ( .IN1(n3756), .IN2(n5241), .QN(WX3878) );
  XOR2X1 U6747 ( .IN1(n2889), .IN2(DFF_557_n1), .Q(n5241) );
  NOR2X0 U6748 ( .IN1(n3756), .IN2(n5242), .QN(WX3876) );
  XOR2X1 U6749 ( .IN1(n2890), .IN2(DFF_556_n1), .Q(n5242) );
  NOR2X0 U6750 ( .IN1(n3756), .IN2(n5243), .QN(WX3874) );
  XOR2X1 U6751 ( .IN1(n2891), .IN2(DFF_555_n1), .Q(n5243) );
  NOR2X0 U6752 ( .IN1(n3756), .IN2(n5244), .QN(WX3872) );
  XOR3X1 U6753 ( .IN1(test_so31), .IN2(n2701), .IN3(DFF_575_n1), .Q(n5244) );
  NOR2X0 U6754 ( .IN1(n3693), .IN2(n5245), .QN(WX3870) );
  XOR2X1 U6755 ( .IN1(n2892), .IN2(DFF_553_n1), .Q(n5245) );
  NOR2X0 U6756 ( .IN1(n3694), .IN2(n5246), .QN(WX3868) );
  XOR2X1 U6757 ( .IN1(n2893), .IN2(DFF_552_n1), .Q(n5246) );
  NOR2X0 U6758 ( .IN1(n3695), .IN2(n5247), .QN(WX3866) );
  XOR2X1 U6759 ( .IN1(n2894), .IN2(DFF_551_n1), .Q(n5247) );
  NOR2X0 U6760 ( .IN1(n3696), .IN2(n5248), .QN(WX3864) );
  XOR2X1 U6761 ( .IN1(n2895), .IN2(DFF_550_n1), .Q(n5248) );
  NOR2X0 U6762 ( .IN1(n3697), .IN2(n5249), .QN(WX3862) );
  XOR2X1 U6763 ( .IN1(CRC_OUT_7_5), .IN2(test_so30), .Q(n5249) );
  NOR2X0 U6764 ( .IN1(n3681), .IN2(n5250), .QN(WX3860) );
  XOR2X1 U6765 ( .IN1(n2896), .IN2(DFF_548_n1), .Q(n5250) );
  NOR2X0 U6766 ( .IN1(n3682), .IN2(n5251), .QN(WX3858) );
  XOR3X1 U6767 ( .IN1(n2702), .IN2(DFF_575_n1), .IN3(CRC_OUT_7_3), .Q(n5251)
         );
  NOR2X0 U6768 ( .IN1(n3683), .IN2(n5252), .QN(WX3856) );
  XOR2X1 U6769 ( .IN1(n2897), .IN2(DFF_546_n1), .Q(n5252) );
  NOR2X0 U6770 ( .IN1(n3684), .IN2(n5253), .QN(WX3854) );
  XOR2X1 U6771 ( .IN1(n2898), .IN2(DFF_545_n1), .Q(n5253) );
  NOR2X0 U6772 ( .IN1(n3685), .IN2(n5254), .QN(WX3852) );
  XOR2X1 U6773 ( .IN1(n2899), .IN2(DFF_544_n1), .Q(n5254) );
  NOR2X0 U6774 ( .IN1(n3686), .IN2(n5255), .QN(WX3850) );
  XOR2X1 U6775 ( .IN1(n2712), .IN2(DFF_575_n1), .Q(n5255) );
  AND2X1 U6776 ( .IN1(n3602), .IN2(test_so24), .Q(WX3324) );
  NOR2X0 U6777 ( .IN1(n6161), .IN2(n3660), .QN(WX3322) );
  NOR2X0 U6778 ( .IN1(n6163), .IN2(n3660), .QN(WX3320) );
  NOR2X0 U6779 ( .IN1(n6165), .IN2(n3660), .QN(WX3318) );
  NOR2X0 U6780 ( .IN1(n6167), .IN2(n3660), .QN(WX3316) );
  NOR2X0 U6781 ( .IN1(n6169), .IN2(n3660), .QN(WX3314) );
  NOR2X0 U6782 ( .IN1(n6171), .IN2(n3660), .QN(WX3312) );
  NOR2X0 U6783 ( .IN1(n6173), .IN2(n3660), .QN(WX3310) );
  NOR2X0 U6784 ( .IN1(n6175), .IN2(n3660), .QN(WX3308) );
  NOR2X0 U6785 ( .IN1(n6177), .IN2(n3660), .QN(WX3306) );
  NOR2X0 U6786 ( .IN1(n6179), .IN2(n3660), .QN(WX3304) );
  NOR2X0 U6787 ( .IN1(n6181), .IN2(n3659), .QN(WX3302) );
  NOR2X0 U6788 ( .IN1(n6183), .IN2(n3659), .QN(WX3300) );
  NOR2X0 U6789 ( .IN1(n6185), .IN2(n3659), .QN(WX3298) );
  NOR2X0 U6790 ( .IN1(n6187), .IN2(n3659), .QN(WX3296) );
  NOR2X0 U6791 ( .IN1(n6190), .IN2(n3659), .QN(WX3294) );
  NAND4X0 U6792 ( .IN1(n5256), .IN2(n5257), .IN3(n5258), .IN4(n5259), .QN(
        WX3292) );
  NAND2X0 U6793 ( .IN1(n5037), .IN2(n3099), .QN(n5259) );
  XOR3X1 U6794 ( .IN1(n3691), .IN2(n2711), .IN3(n5260), .Q(n5037) );
  XOR2X1 U6795 ( .IN1(WX4714), .IN2(test_so36), .Q(n5260) );
  NAND2X0 U6796 ( .IN1(n3015), .IN2(n5261), .QN(n5258) );
  NAND2X0 U6797 ( .IN1(WX3130), .IN2(n3039), .QN(n5257) );
  NAND2X0 U6798 ( .IN1(n3051), .IN2(CRC_OUT_7_0), .QN(n5256) );
  NAND4X0 U6799 ( .IN1(n5262), .IN2(n5263), .IN3(n5264), .IN4(n5265), .QN(
        WX3290) );
  NAND2X0 U6800 ( .IN1(n3083), .IN2(n5043), .QN(n5265) );
  XNOR3X1 U6801 ( .IN1(n2873), .IN2(n2633), .IN3(n5266), .Q(n5043) );
  XOR2X1 U6802 ( .IN1(WX4648), .IN2(n6106), .Q(n5266) );
  NAND2X0 U6803 ( .IN1(n3015), .IN2(n5267), .QN(n5264) );
  NAND2X0 U6804 ( .IN1(WX3128), .IN2(n3039), .QN(n5263) );
  NAND2X0 U6805 ( .IN1(n3051), .IN2(CRC_OUT_7_1), .QN(n5262) );
  NAND4X0 U6806 ( .IN1(n5268), .IN2(n5269), .IN3(n5270), .IN4(n5271), .QN(
        WX3288) );
  NAND2X0 U6807 ( .IN1(n3083), .IN2(n5049), .QN(n5271) );
  XNOR3X1 U6808 ( .IN1(n2872), .IN2(n2634), .IN3(n5272), .Q(n5049) );
  XOR2X1 U6809 ( .IN1(WX4646), .IN2(n6107), .Q(n5272) );
  NAND2X0 U6810 ( .IN1(n3015), .IN2(n5273), .QN(n5270) );
  NAND2X0 U6811 ( .IN1(WX3126), .IN2(n3039), .QN(n5269) );
  NAND2X0 U6812 ( .IN1(n3051), .IN2(CRC_OUT_7_2), .QN(n5268) );
  NAND4X0 U6813 ( .IN1(n5274), .IN2(n5275), .IN3(n5276), .IN4(n5277), .QN(
        WX3286) );
  NAND2X0 U6814 ( .IN1(n3083), .IN2(n5055), .QN(n5277) );
  XNOR3X1 U6815 ( .IN1(n2871), .IN2(n2635), .IN3(n5278), .Q(n5055) );
  XOR2X1 U6816 ( .IN1(WX4644), .IN2(n6108), .Q(n5278) );
  NAND2X0 U6817 ( .IN1(n3015), .IN2(n5279), .QN(n5276) );
  NAND2X0 U6818 ( .IN1(WX3124), .IN2(n3039), .QN(n5275) );
  NAND2X0 U6819 ( .IN1(n3051), .IN2(CRC_OUT_7_3), .QN(n5274) );
  NAND4X0 U6820 ( .IN1(n5280), .IN2(n5281), .IN3(n5282), .IN4(n5283), .QN(
        WX3284) );
  NAND2X0 U6821 ( .IN1(n3083), .IN2(n5061), .QN(n5283) );
  XNOR3X1 U6822 ( .IN1(n2699), .IN2(n2636), .IN3(n5284), .Q(n5061) );
  XOR2X1 U6823 ( .IN1(WX4642), .IN2(n6109), .Q(n5284) );
  NAND2X0 U6824 ( .IN1(n3015), .IN2(n5285), .QN(n5282) );
  NAND2X0 U6825 ( .IN1(WX3122), .IN2(n3039), .QN(n5281) );
  NAND2X0 U6826 ( .IN1(n3051), .IN2(CRC_OUT_7_4), .QN(n5280) );
  NAND4X0 U6827 ( .IN1(n5286), .IN2(n5287), .IN3(n5288), .IN4(n5289), .QN(
        WX3282) );
  NAND2X0 U6828 ( .IN1(n3083), .IN2(n5067), .QN(n5289) );
  XNOR3X1 U6829 ( .IN1(n2870), .IN2(n2637), .IN3(n5290), .Q(n5067) );
  XOR2X1 U6830 ( .IN1(WX4640), .IN2(n6110), .Q(n5290) );
  NAND2X0 U6831 ( .IN1(n3015), .IN2(n5291), .QN(n5288) );
  NAND2X0 U6832 ( .IN1(WX3120), .IN2(n3039), .QN(n5287) );
  NAND2X0 U6833 ( .IN1(n3051), .IN2(CRC_OUT_7_5), .QN(n5286) );
  NAND4X0 U6834 ( .IN1(n5292), .IN2(n5293), .IN3(n5294), .IN4(n5295), .QN(
        WX3280) );
  NAND2X0 U6835 ( .IN1(n3083), .IN2(n5073), .QN(n5295) );
  XNOR3X1 U6836 ( .IN1(n2869), .IN2(n2638), .IN3(n5296), .Q(n5073) );
  XOR2X1 U6837 ( .IN1(WX4638), .IN2(n6111), .Q(n5296) );
  NAND2X0 U6838 ( .IN1(n5297), .IN2(n3017), .QN(n5294) );
  NAND2X0 U6839 ( .IN1(WX3118), .IN2(n3039), .QN(n5293) );
  NAND2X0 U6840 ( .IN1(n3051), .IN2(CRC_OUT_7_6), .QN(n5292) );
  NAND4X0 U6841 ( .IN1(n5298), .IN2(n5299), .IN3(n5300), .IN4(n5301), .QN(
        WX3278) );
  NAND2X0 U6842 ( .IN1(n3083), .IN2(n5079), .QN(n5301) );
  XNOR3X1 U6843 ( .IN1(n2868), .IN2(n2639), .IN3(n5302), .Q(n5079) );
  XOR2X1 U6844 ( .IN1(WX4636), .IN2(n6112), .Q(n5302) );
  NAND2X0 U6845 ( .IN1(n3016), .IN2(n5303), .QN(n5300) );
  NAND2X0 U6846 ( .IN1(WX3116), .IN2(n3039), .QN(n5299) );
  NAND2X0 U6847 ( .IN1(n3051), .IN2(CRC_OUT_7_7), .QN(n5298) );
  NAND4X0 U6848 ( .IN1(n5304), .IN2(n5305), .IN3(n5306), .IN4(n5307), .QN(
        WX3276) );
  NAND2X0 U6849 ( .IN1(n3083), .IN2(n5085), .QN(n5307) );
  XNOR3X1 U6850 ( .IN1(n2867), .IN2(n2640), .IN3(n5308), .Q(n5085) );
  XOR2X1 U6851 ( .IN1(WX4634), .IN2(n6113), .Q(n5308) );
  NAND2X0 U6852 ( .IN1(n5309), .IN2(n3018), .QN(n5306) );
  NAND2X0 U6853 ( .IN1(WX3114), .IN2(n3039), .QN(n5305) );
  NAND2X0 U6854 ( .IN1(n3051), .IN2(CRC_OUT_7_8), .QN(n5304) );
  NAND4X0 U6855 ( .IN1(n5310), .IN2(n5311), .IN3(n5312), .IN4(n5313), .QN(
        WX3274) );
  NAND2X0 U6856 ( .IN1(n3083), .IN2(n5091), .QN(n5313) );
  XNOR3X1 U6857 ( .IN1(n2866), .IN2(n2641), .IN3(n5314), .Q(n5091) );
  XOR2X1 U6858 ( .IN1(WX4632), .IN2(n6114), .Q(n5314) );
  NAND2X0 U6859 ( .IN1(n3016), .IN2(n5315), .QN(n5312) );
  NAND2X0 U6860 ( .IN1(WX3112), .IN2(n3039), .QN(n5311) );
  NAND2X0 U6861 ( .IN1(n3051), .IN2(CRC_OUT_7_9), .QN(n5310) );
  NAND4X0 U6862 ( .IN1(n5316), .IN2(n5317), .IN3(n5318), .IN4(n5319), .QN(
        WX3272) );
  NAND2X0 U6863 ( .IN1(n3084), .IN2(n5097), .QN(n5319) );
  XNOR3X1 U6864 ( .IN1(n2865), .IN2(n2642), .IN3(n5320), .Q(n5097) );
  XOR2X1 U6865 ( .IN1(WX4630), .IN2(n6115), .Q(n5320) );
  NAND2X0 U6866 ( .IN1(n3016), .IN2(n5321), .QN(n5318) );
  NAND2X0 U6867 ( .IN1(WX3110), .IN2(n3039), .QN(n5317) );
  NAND2X0 U6868 ( .IN1(test_so31), .IN2(n3070), .QN(n5316) );
  NAND4X0 U6869 ( .IN1(n5322), .IN2(n5323), .IN3(n5324), .IN4(n5325), .QN(
        WX3270) );
  NAND2X0 U6870 ( .IN1(n5103), .IN2(n3099), .QN(n5325) );
  XOR3X1 U6871 ( .IN1(n3713), .IN2(n2643), .IN3(n5326), .Q(n5103) );
  XOR2X1 U6872 ( .IN1(WX4564), .IN2(test_so41), .Q(n5326) );
  NAND2X0 U6873 ( .IN1(n3016), .IN2(n5327), .QN(n5324) );
  NAND2X0 U6874 ( .IN1(WX3108), .IN2(n3039), .QN(n5323) );
  NAND2X0 U6875 ( .IN1(n3051), .IN2(CRC_OUT_7_11), .QN(n5322) );
  NAND4X0 U6876 ( .IN1(n5328), .IN2(n5329), .IN3(n5330), .IN4(n5331), .QN(
        WX3268) );
  NAND2X0 U6877 ( .IN1(n3084), .IN2(n5109), .QN(n5331) );
  XNOR3X1 U6878 ( .IN1(n2864), .IN2(n2644), .IN3(n5332), .Q(n5109) );
  XOR2X1 U6879 ( .IN1(WX4626), .IN2(n6116), .Q(n5332) );
  NAND2X0 U6880 ( .IN1(n5333), .IN2(n3020), .QN(n5330) );
  NAND2X0 U6881 ( .IN1(WX3106), .IN2(n3039), .QN(n5329) );
  NAND2X0 U6882 ( .IN1(n3052), .IN2(CRC_OUT_7_12), .QN(n5328) );
  NAND4X0 U6883 ( .IN1(n5334), .IN2(n5335), .IN3(n5336), .IN4(n5337), .QN(
        WX3266) );
  NAND2X0 U6884 ( .IN1(n5115), .IN2(n3099), .QN(n5337) );
  XOR3X1 U6885 ( .IN1(n3717), .IN2(n2863), .IN3(n5338), .Q(n5115) );
  XOR2X1 U6886 ( .IN1(WX4560), .IN2(test_so39), .Q(n5338) );
  NAND2X0 U6887 ( .IN1(n3016), .IN2(n5339), .QN(n5336) );
  NAND2X0 U6888 ( .IN1(WX3104), .IN2(n3039), .QN(n5335) );
  NAND2X0 U6889 ( .IN1(n3052), .IN2(CRC_OUT_7_13), .QN(n5334) );
  NAND4X0 U6890 ( .IN1(n5340), .IN2(n5341), .IN3(n5342), .IN4(n5343), .QN(
        WX3264) );
  NAND2X0 U6891 ( .IN1(n3084), .IN2(n5121), .QN(n5343) );
  XNOR3X1 U6892 ( .IN1(n2862), .IN2(n2645), .IN3(n5344), .Q(n5121) );
  XOR2X1 U6893 ( .IN1(WX4622), .IN2(n6117), .Q(n5344) );
  NAND2X0 U6894 ( .IN1(n3016), .IN2(n5345), .QN(n5342) );
  NAND2X0 U6895 ( .IN1(WX3102), .IN2(n3039), .QN(n5341) );
  NAND2X0 U6896 ( .IN1(n3052), .IN2(CRC_OUT_7_14), .QN(n5340) );
  NAND4X0 U6897 ( .IN1(n5346), .IN2(n5347), .IN3(n5348), .IN4(n5349), .QN(
        WX3262) );
  NAND2X0 U6898 ( .IN1(n5127), .IN2(n3099), .QN(n5349) );
  XOR3X1 U6899 ( .IN1(n2861), .IN2(n2646), .IN3(n5350), .Q(n5127) );
  XOR2X1 U6900 ( .IN1(WX4556), .IN2(test_so37), .Q(n5350) );
  NAND2X0 U6901 ( .IN1(n3016), .IN2(n5351), .QN(n5348) );
  NAND2X0 U6902 ( .IN1(WX3100), .IN2(n3039), .QN(n5347) );
  NAND2X0 U6903 ( .IN1(n3052), .IN2(CRC_OUT_7_15), .QN(n5346) );
  NAND4X0 U6904 ( .IN1(n5352), .IN2(n5353), .IN3(n5354), .IN4(n5355), .QN(
        WX3260) );
  NAND2X0 U6905 ( .IN1(n3084), .IN2(n5133), .QN(n5355) );
  XNOR3X1 U6906 ( .IN1(n2482), .IN2(n3572), .IN3(n5356), .Q(n5133) );
  XOR3X1 U6907 ( .IN1(n6118), .IN2(n2698), .IN3(WX4682), .Q(n5356) );
  NAND2X0 U6908 ( .IN1(n5357), .IN2(n3021), .QN(n5354) );
  NAND2X0 U6909 ( .IN1(WX3098), .IN2(n3039), .QN(n5353) );
  NAND2X0 U6910 ( .IN1(n3052), .IN2(CRC_OUT_7_16), .QN(n5352) );
  NAND4X0 U6911 ( .IN1(n5358), .IN2(n5359), .IN3(n5360), .IN4(n5361), .QN(
        WX3258) );
  NAND2X0 U6912 ( .IN1(n5139), .IN2(n3099), .QN(n5361) );
  XOR3X1 U6913 ( .IN1(n2484), .IN2(n3578), .IN3(n5362), .Q(n5139) );
  XNOR3X1 U6914 ( .IN1(test_so35), .IN2(n6119), .IN3(n2860), .Q(n5362) );
  NAND2X0 U6915 ( .IN1(n3013), .IN2(n5363), .QN(n5360) );
  NAND2X0 U6916 ( .IN1(WX3096), .IN2(n3040), .QN(n5359) );
  NAND2X0 U6917 ( .IN1(n3052), .IN2(CRC_OUT_7_17), .QN(n5358) );
  NAND4X0 U6918 ( .IN1(n5364), .IN2(n5365), .IN3(n5366), .IN4(n5367), .QN(
        WX3256) );
  NAND2X0 U6919 ( .IN1(n3084), .IN2(n5145), .QN(n5367) );
  XNOR3X1 U6920 ( .IN1(n2485), .IN2(n3572), .IN3(n5368), .Q(n5145) );
  XOR3X1 U6921 ( .IN1(n6120), .IN2(n2859), .IN3(WX4678), .Q(n5368) );
  NAND2X0 U6922 ( .IN1(n3013), .IN2(n5369), .QN(n5366) );
  NAND2X0 U6923 ( .IN1(WX3094), .IN2(n3040), .QN(n5365) );
  NAND2X0 U6924 ( .IN1(n3052), .IN2(CRC_OUT_7_18), .QN(n5364) );
  NAND4X0 U6925 ( .IN1(n5370), .IN2(n5371), .IN3(n5372), .IN4(n5373), .QN(
        WX3254) );
  NAND2X0 U6926 ( .IN1(n3084), .IN2(n5151), .QN(n5373) );
  XNOR3X1 U6927 ( .IN1(n2487), .IN2(n3572), .IN3(n5374), .Q(n5151) );
  XOR3X1 U6928 ( .IN1(n6121), .IN2(n2858), .IN3(WX4676), .Q(n5374) );
  NAND2X0 U6929 ( .IN1(n3013), .IN2(n5375), .QN(n5372) );
  NAND2X0 U6930 ( .IN1(WX3092), .IN2(n3040), .QN(n5371) );
  NAND2X0 U6931 ( .IN1(n3052), .IN2(CRC_OUT_7_19), .QN(n5370) );
  NAND4X0 U6932 ( .IN1(n5376), .IN2(n5377), .IN3(n5378), .IN4(n5379), .QN(
        WX3252) );
  NAND2X0 U6933 ( .IN1(n3084), .IN2(n5157), .QN(n5379) );
  XNOR3X1 U6934 ( .IN1(n2489), .IN2(n3572), .IN3(n5380), .Q(n5157) );
  XOR3X1 U6935 ( .IN1(n6122), .IN2(n2857), .IN3(WX4674), .Q(n5380) );
  NAND2X0 U6936 ( .IN1(n3013), .IN2(n5381), .QN(n5378) );
  NAND2X0 U6937 ( .IN1(WX3090), .IN2(n3040), .QN(n5377) );
  NAND2X0 U6938 ( .IN1(n3052), .IN2(CRC_OUT_7_20), .QN(n5376) );
  NAND4X0 U6939 ( .IN1(n5382), .IN2(n5383), .IN3(n5384), .IN4(n5385), .QN(
        WX3250) );
  NAND2X0 U6940 ( .IN1(n3084), .IN2(n5163), .QN(n5385) );
  XNOR3X1 U6941 ( .IN1(n2491), .IN2(n3572), .IN3(n5386), .Q(n5163) );
  XOR3X1 U6942 ( .IN1(n6123), .IN2(n2856), .IN3(WX4672), .Q(n5386) );
  NAND2X0 U6943 ( .IN1(n3013), .IN2(n5387), .QN(n5384) );
  NAND2X0 U6944 ( .IN1(WX3088), .IN2(n3040), .QN(n5383) );
  NAND2X0 U6945 ( .IN1(n3052), .IN2(CRC_OUT_7_21), .QN(n5382) );
  NAND4X0 U6946 ( .IN1(n5388), .IN2(n5389), .IN3(n5390), .IN4(n5391), .QN(
        WX3248) );
  NAND2X0 U6947 ( .IN1(n3084), .IN2(n5169), .QN(n5391) );
  XNOR3X1 U6948 ( .IN1(n2493), .IN2(n3572), .IN3(n5392), .Q(n5169) );
  XOR3X1 U6949 ( .IN1(n6124), .IN2(n2855), .IN3(WX4670), .Q(n5392) );
  NAND2X0 U6950 ( .IN1(n3012), .IN2(n5393), .QN(n5390) );
  NAND2X0 U6951 ( .IN1(WX3086), .IN2(n3040), .QN(n5389) );
  NAND2X0 U6952 ( .IN1(n3052), .IN2(CRC_OUT_7_22), .QN(n5388) );
  NAND4X0 U6953 ( .IN1(n5394), .IN2(n5395), .IN3(n5396), .IN4(n5397), .QN(
        WX3246) );
  NAND2X0 U6954 ( .IN1(n3087), .IN2(n5175), .QN(n5397) );
  XNOR3X1 U6955 ( .IN1(n2495), .IN2(n3572), .IN3(n5398), .Q(n5175) );
  XOR3X1 U6956 ( .IN1(n6125), .IN2(n2854), .IN3(WX4668), .Q(n5398) );
  NAND2X0 U6957 ( .IN1(n5399), .IN2(n3020), .QN(n5396) );
  NAND2X0 U6958 ( .IN1(WX3084), .IN2(n3040), .QN(n5395) );
  NAND2X0 U6959 ( .IN1(n3058), .IN2(CRC_OUT_7_23), .QN(n5394) );
  NAND4X0 U6960 ( .IN1(n5400), .IN2(n5401), .IN3(n5402), .IN4(n5403), .QN(
        WX3244) );
  NAND2X0 U6961 ( .IN1(n3084), .IN2(n5181), .QN(n5403) );
  XNOR3X1 U6962 ( .IN1(n2497), .IN2(n3572), .IN3(n5404), .Q(n5181) );
  XOR3X1 U6963 ( .IN1(n6126), .IN2(n2853), .IN3(WX4666), .Q(n5404) );
  NAND2X0 U6964 ( .IN1(n3012), .IN2(n5405), .QN(n5402) );
  NAND2X0 U6965 ( .IN1(WX3082), .IN2(n3040), .QN(n5401) );
  NAND2X0 U6966 ( .IN1(n3053), .IN2(CRC_OUT_7_24), .QN(n5400) );
  NAND4X0 U6967 ( .IN1(n5406), .IN2(n5407), .IN3(n5408), .IN4(n5409), .QN(
        WX3242) );
  NAND2X0 U6968 ( .IN1(n3084), .IN2(n5187), .QN(n5409) );
  XNOR3X1 U6969 ( .IN1(n2499), .IN2(n3572), .IN3(n5410), .Q(n5187) );
  XOR3X1 U6970 ( .IN1(n6127), .IN2(n2852), .IN3(WX4664), .Q(n5410) );
  NAND2X0 U6971 ( .IN1(n3012), .IN2(n5411), .QN(n5408) );
  NAND2X0 U6972 ( .IN1(WX3080), .IN2(n3040), .QN(n5407) );
  NAND2X0 U6973 ( .IN1(n3053), .IN2(CRC_OUT_7_25), .QN(n5406) );
  NAND4X0 U6974 ( .IN1(n5412), .IN2(n5413), .IN3(n5414), .IN4(n5415), .QN(
        WX3240) );
  NAND2X0 U6975 ( .IN1(n3084), .IN2(n5193), .QN(n5415) );
  XNOR3X1 U6976 ( .IN1(n2501), .IN2(n3572), .IN3(n5416), .Q(n5193) );
  XOR3X1 U6977 ( .IN1(n6128), .IN2(n2851), .IN3(WX4662), .Q(n5416) );
  NAND2X0 U6978 ( .IN1(n5417), .IN2(n3018), .QN(n5414) );
  NAND2X0 U6979 ( .IN1(WX3078), .IN2(n3040), .QN(n5413) );
  NAND2X0 U6980 ( .IN1(n3053), .IN2(CRC_OUT_7_26), .QN(n5412) );
  NAND4X0 U6981 ( .IN1(n5418), .IN2(n5419), .IN3(n5420), .IN4(n5421), .QN(
        WX3238) );
  NAND2X0 U6982 ( .IN1(n3085), .IN2(n5199), .QN(n5421) );
  XNOR3X1 U6983 ( .IN1(n2503), .IN2(n3572), .IN3(n5422), .Q(n5199) );
  XOR3X1 U6984 ( .IN1(n6129), .IN2(n2850), .IN3(WX4660), .Q(n5422) );
  NAND2X0 U6985 ( .IN1(n3012), .IN2(n5423), .QN(n5420) );
  NAND2X0 U6986 ( .IN1(WX3076), .IN2(n3040), .QN(n5419) );
  NAND2X0 U6987 ( .IN1(test_so32), .IN2(n3069), .QN(n5418) );
  NAND4X0 U6988 ( .IN1(n5424), .IN2(n5425), .IN3(n5426), .IN4(n5427), .QN(
        WX3236) );
  NAND2X0 U6989 ( .IN1(n5205), .IN2(n3098), .QN(n5427) );
  XOR3X1 U6990 ( .IN1(n2505), .IN2(n3578), .IN3(n5428), .Q(n5205) );
  XOR3X1 U6991 ( .IN1(test_so40), .IN2(n6130), .IN3(WX4658), .Q(n5428) );
  NAND2X0 U6992 ( .IN1(n3012), .IN2(n5429), .QN(n5426) );
  NAND2X0 U6993 ( .IN1(WX3074), .IN2(n3040), .QN(n5425) );
  NAND2X0 U6994 ( .IN1(n3053), .IN2(CRC_OUT_7_28), .QN(n5424) );
  NAND4X0 U6995 ( .IN1(n5430), .IN2(n5431), .IN3(n5432), .IN4(n5433), .QN(
        WX3234) );
  NAND2X0 U6996 ( .IN1(n3085), .IN2(n5211), .QN(n5433) );
  XNOR3X1 U6997 ( .IN1(n2506), .IN2(n3573), .IN3(n5434), .Q(n5211) );
  XOR3X1 U6998 ( .IN1(n6131), .IN2(n2849), .IN3(WX4656), .Q(n5434) );
  NAND2X0 U6999 ( .IN1(n3012), .IN2(n5435), .QN(n5432) );
  NAND2X0 U7000 ( .IN1(WX3072), .IN2(n3040), .QN(n5431) );
  NAND2X0 U7001 ( .IN1(n3053), .IN2(CRC_OUT_7_29), .QN(n5430) );
  NAND4X0 U7002 ( .IN1(n5436), .IN2(n5437), .IN3(n5438), .IN4(n5439), .QN(
        WX3232) );
  NAND2X0 U7003 ( .IN1(n5217), .IN2(n3098), .QN(n5439) );
  XOR3X1 U7004 ( .IN1(n2508), .IN2(n3577), .IN3(n5440), .Q(n5217) );
  XNOR3X1 U7005 ( .IN1(test_so38), .IN2(n6132), .IN3(n2848), .Q(n5440) );
  NAND2X0 U7006 ( .IN1(n5441), .IN2(n3017), .QN(n5438) );
  NAND2X0 U7007 ( .IN1(WX3070), .IN2(n3040), .QN(n5437) );
  NAND2X0 U7008 ( .IN1(n3053), .IN2(CRC_OUT_7_30), .QN(n5436) );
  NAND4X0 U7009 ( .IN1(n5442), .IN2(n5443), .IN3(n5444), .IN4(n5445), .QN(
        WX3230) );
  NAND2X0 U7010 ( .IN1(n3085), .IN2(n5223), .QN(n5445) );
  XNOR3X1 U7011 ( .IN1(n2344), .IN2(n3573), .IN3(n5446), .Q(n5223) );
  XOR3X1 U7012 ( .IN1(n6133), .IN2(n2847), .IN3(WX4652), .Q(n5446) );
  NAND2X0 U7013 ( .IN1(n3012), .IN2(n5447), .QN(n5444) );
  NAND2X0 U7014 ( .IN1(n3053), .IN2(CRC_OUT_7_31), .QN(n5443) );
  NAND2X0 U7015 ( .IN1(n2245), .IN2(WX3071), .QN(n5442) );
  NOR2X0 U7016 ( .IN1(n3734), .IN2(WX3071), .QN(WX3132) );
  AND2X1 U7017 ( .IN1(n3602), .IN2(n8612), .Q(WX3130) );
  AND2X1 U7018 ( .IN1(n3602), .IN2(n8613), .Q(WX3128) );
  AND2X1 U7019 ( .IN1(test_so23), .IN2(n3599), .Q(WX3126) );
  AND2X1 U7020 ( .IN1(n3602), .IN2(n8616), .Q(WX3124) );
  AND2X1 U7021 ( .IN1(n3603), .IN2(n8617), .Q(WX3122) );
  AND2X1 U7022 ( .IN1(n3602), .IN2(n8618), .Q(WX3120) );
  AND2X1 U7023 ( .IN1(n3603), .IN2(n8619), .Q(WX3118) );
  AND2X1 U7024 ( .IN1(n3604), .IN2(n8620), .Q(WX3116) );
  AND2X1 U7025 ( .IN1(n3603), .IN2(n8621), .Q(WX3114) );
  AND2X1 U7026 ( .IN1(n3603), .IN2(n8622), .Q(WX3112) );
  AND2X1 U7027 ( .IN1(n3603), .IN2(n8623), .Q(WX3110) );
  AND2X1 U7028 ( .IN1(n3603), .IN2(n8624), .Q(WX3108) );
  AND2X1 U7029 ( .IN1(n3603), .IN2(n8625), .Q(WX3106) );
  AND2X1 U7030 ( .IN1(n3604), .IN2(n8626), .Q(WX3104) );
  AND2X1 U7031 ( .IN1(n3603), .IN2(n8627), .Q(WX3102) );
  AND2X1 U7032 ( .IN1(n3604), .IN2(n8628), .Q(WX3100) );
  AND2X1 U7033 ( .IN1(n3604), .IN2(n8629), .Q(WX3098) );
  AND2X1 U7034 ( .IN1(n3604), .IN2(n8630), .Q(WX3096) );
  AND2X1 U7035 ( .IN1(n3604), .IN2(n8631), .Q(WX3094) );
  AND2X1 U7036 ( .IN1(n3604), .IN2(n8632), .Q(WX3092) );
  AND2X1 U7037 ( .IN1(test_so22), .IN2(n3599), .Q(WX3090) );
  AND2X1 U7038 ( .IN1(n3604), .IN2(n8635), .Q(WX3088) );
  AND2X1 U7039 ( .IN1(n3605), .IN2(n8636), .Q(WX3086) );
  AND2X1 U7040 ( .IN1(n3604), .IN2(n8637), .Q(WX3084) );
  AND2X1 U7041 ( .IN1(n3605), .IN2(n8638), .Q(WX3082) );
  AND2X1 U7042 ( .IN1(n3605), .IN2(n8639), .Q(WX3080) );
  AND2X1 U7043 ( .IN1(n3605), .IN2(n8640), .Q(WX3078) );
  AND2X1 U7044 ( .IN1(n3605), .IN2(n8641), .Q(WX3076) );
  AND2X1 U7045 ( .IN1(n3605), .IN2(n8642), .Q(WX3074) );
  AND2X1 U7046 ( .IN1(n3605), .IN2(n8643), .Q(WX3072) );
  AND2X1 U7047 ( .IN1(n3605), .IN2(n8644), .Q(WX3070) );
  NOR2X0 U7048 ( .IN1(n3736), .IN2(n5448), .QN(WX2619) );
  XOR2X1 U7049 ( .IN1(n2900), .IN2(DFF_382_n1), .Q(n5448) );
  NOR2X0 U7050 ( .IN1(n3734), .IN2(n5449), .QN(WX2617) );
  XOR2X1 U7051 ( .IN1(n2901), .IN2(DFF_381_n1), .Q(n5449) );
  NOR2X0 U7052 ( .IN1(n3736), .IN2(n5450), .QN(WX2615) );
  XOR2X1 U7053 ( .IN1(n2902), .IN2(DFF_380_n1), .Q(n5450) );
  NOR2X0 U7054 ( .IN1(n3736), .IN2(n5451), .QN(WX2613) );
  XOR2X1 U7055 ( .IN1(CRC_OUT_8_27), .IN2(test_so18), .Q(n5451) );
  NOR2X0 U7056 ( .IN1(n3734), .IN2(n5452), .QN(WX2611) );
  XOR2X1 U7057 ( .IN1(n2903), .IN2(DFF_378_n1), .Q(n5452) );
  NOR2X0 U7058 ( .IN1(n3734), .IN2(n5453), .QN(WX2609) );
  XNOR2X1 U7059 ( .IN1(n2904), .IN2(test_so21), .Q(n5453) );
  NOR2X0 U7060 ( .IN1(n3736), .IN2(n5454), .QN(WX2607) );
  XOR2X1 U7061 ( .IN1(n2905), .IN2(DFF_376_n1), .Q(n5454) );
  NOR2X0 U7062 ( .IN1(n3734), .IN2(n5455), .QN(WX2605) );
  XOR2X1 U7063 ( .IN1(n2906), .IN2(DFF_375_n1), .Q(n5455) );
  NOR2X0 U7064 ( .IN1(n3734), .IN2(n5456), .QN(WX2603) );
  XOR2X1 U7065 ( .IN1(n2907), .IN2(DFF_374_n1), .Q(n5456) );
  NOR2X0 U7066 ( .IN1(n3736), .IN2(n5457), .QN(WX2601) );
  XOR2X1 U7067 ( .IN1(n2908), .IN2(DFF_373_n1), .Q(n5457) );
  NOR2X0 U7068 ( .IN1(n3734), .IN2(n5458), .QN(WX2599) );
  XOR2X1 U7069 ( .IN1(n2909), .IN2(DFF_372_n1), .Q(n5458) );
  NOR2X0 U7070 ( .IN1(n3734), .IN2(n5459), .QN(WX2597) );
  XOR2X1 U7071 ( .IN1(n2910), .IN2(DFF_371_n1), .Q(n5459) );
  NOR2X0 U7072 ( .IN1(n3733), .IN2(n5460), .QN(WX2595) );
  XOR2X1 U7073 ( .IN1(n2911), .IN2(DFF_370_n1), .Q(n5460) );
  NOR2X0 U7074 ( .IN1(n3733), .IN2(n5461), .QN(WX2593) );
  XOR2X1 U7075 ( .IN1(n2912), .IN2(DFF_369_n1), .Q(n5461) );
  NOR2X0 U7076 ( .IN1(n3734), .IN2(n5462), .QN(WX2591) );
  XOR2X1 U7077 ( .IN1(n2913), .IN2(DFF_368_n1), .Q(n5462) );
  NOR2X0 U7078 ( .IN1(n3733), .IN2(n5463), .QN(WX2589) );
  XOR3X1 U7079 ( .IN1(n2703), .IN2(DFF_383_n1), .IN3(CRC_OUT_8_15), .Q(n5463)
         );
  NOR2X0 U7080 ( .IN1(n3733), .IN2(n5464), .QN(WX2587) );
  XOR2X1 U7081 ( .IN1(n2914), .IN2(DFF_366_n1), .Q(n5464) );
  NOR2X0 U7082 ( .IN1(n3733), .IN2(n5465), .QN(WX2585) );
  XOR2X1 U7083 ( .IN1(n2915), .IN2(DFF_365_n1), .Q(n5465) );
  NOR2X0 U7084 ( .IN1(n3733), .IN2(n5466), .QN(WX2583) );
  XOR2X1 U7085 ( .IN1(n2916), .IN2(DFF_364_n1), .Q(n5466) );
  NOR2X0 U7086 ( .IN1(n3733), .IN2(n5467), .QN(WX2581) );
  XOR2X1 U7087 ( .IN1(n2917), .IN2(DFF_363_n1), .Q(n5467) );
  NOR2X0 U7088 ( .IN1(n3734), .IN2(n5468), .QN(WX2579) );
  XOR3X1 U7089 ( .IN1(n2704), .IN2(DFF_383_n1), .IN3(CRC_OUT_8_10), .Q(n5468)
         );
  NOR2X0 U7090 ( .IN1(n3734), .IN2(n5469), .QN(WX2577) );
  XOR2X1 U7091 ( .IN1(CRC_OUT_8_9), .IN2(test_so19), .Q(n5469) );
  NOR2X0 U7092 ( .IN1(n3733), .IN2(n5470), .QN(WX2575) );
  XOR2X1 U7093 ( .IN1(n2918), .IN2(DFF_360_n1), .Q(n5470) );
  NOR2X0 U7094 ( .IN1(n3734), .IN2(n5471), .QN(WX2573) );
  XNOR2X1 U7095 ( .IN1(n2919), .IN2(test_so20), .Q(n5471) );
  NOR2X0 U7096 ( .IN1(n3733), .IN2(n5472), .QN(WX2571) );
  XOR2X1 U7097 ( .IN1(n2920), .IN2(DFF_358_n1), .Q(n5472) );
  NOR2X0 U7098 ( .IN1(n3733), .IN2(n5473), .QN(WX2569) );
  XOR2X1 U7099 ( .IN1(n2921), .IN2(DFF_357_n1), .Q(n5473) );
  NOR2X0 U7100 ( .IN1(n3734), .IN2(n5474), .QN(WX2567) );
  XOR2X1 U7101 ( .IN1(n2922), .IN2(DFF_356_n1), .Q(n5474) );
  NOR2X0 U7102 ( .IN1(n3733), .IN2(n5475), .QN(WX2565) );
  XOR3X1 U7103 ( .IN1(n2705), .IN2(DFF_383_n1), .IN3(CRC_OUT_8_3), .Q(n5475)
         );
  NOR2X0 U7104 ( .IN1(n3733), .IN2(n5476), .QN(WX2563) );
  XOR2X1 U7105 ( .IN1(n2923), .IN2(DFF_354_n1), .Q(n5476) );
  NOR2X0 U7106 ( .IN1(n3737), .IN2(n5477), .QN(WX2561) );
  XOR2X1 U7107 ( .IN1(n2924), .IN2(DFF_353_n1), .Q(n5477) );
  NOR2X0 U7108 ( .IN1(n3733), .IN2(n5478), .QN(WX2559) );
  XOR2X1 U7109 ( .IN1(n2925), .IN2(DFF_352_n1), .Q(n5478) );
  NOR2X0 U7110 ( .IN1(n3737), .IN2(n5479), .QN(WX2557) );
  XOR2X1 U7111 ( .IN1(n2713), .IN2(DFF_383_n1), .Q(n5479) );
  NOR2X0 U7112 ( .IN1(n6160), .IN2(n3659), .QN(WX2031) );
  NOR2X0 U7113 ( .IN1(n6162), .IN2(n3659), .QN(WX2029) );
  NOR2X0 U7114 ( .IN1(n6164), .IN2(n3659), .QN(WX2027) );
  NOR2X0 U7115 ( .IN1(n6166), .IN2(n3659), .QN(WX2025) );
  NOR2X0 U7116 ( .IN1(n6168), .IN2(n3659), .QN(WX2023) );
  NOR2X0 U7117 ( .IN1(n6170), .IN2(n3659), .QN(WX2021) );
  AND2X1 U7118 ( .IN1(n3605), .IN2(test_so13), .Q(WX2019) );
  NOR2X0 U7119 ( .IN1(n6174), .IN2(n3658), .QN(WX2017) );
  NOR2X0 U7120 ( .IN1(n6176), .IN2(n3658), .QN(WX2015) );
  NOR2X0 U7121 ( .IN1(n6178), .IN2(n3658), .QN(WX2013) );
  NOR2X0 U7122 ( .IN1(n6180), .IN2(n3658), .QN(WX2011) );
  NOR2X0 U7123 ( .IN1(n6182), .IN2(n3658), .QN(WX2009) );
  NOR2X0 U7124 ( .IN1(n6184), .IN2(n3658), .QN(WX2007) );
  NOR2X0 U7125 ( .IN1(n6186), .IN2(n3658), .QN(WX2005) );
  NOR2X0 U7126 ( .IN1(n6188), .IN2(n3658), .QN(WX2003) );
  NOR2X0 U7127 ( .IN1(n6189), .IN2(n3658), .QN(WX2001) );
  NAND4X0 U7128 ( .IN1(n5480), .IN2(n5481), .IN3(n5482), .IN4(n5483), .QN(
        WX1999) );
  NAND2X0 U7129 ( .IN1(n3085), .IN2(n5261), .QN(n5483) );
  XNOR3X1 U7130 ( .IN1(n2712), .IN2(n2647), .IN3(n5484), .Q(n5261) );
  XOR2X1 U7131 ( .IN1(WX3357), .IN2(n6134), .Q(n5484) );
  NAND2X0 U7132 ( .IN1(n4588), .IN2(n3018), .QN(n5482) );
  XOR3X1 U7133 ( .IN1(n2713), .IN2(n2662), .IN3(n5485), .Q(n4588) );
  XOR2X1 U7134 ( .IN1(WX2000), .IN2(test_so16), .Q(n5485) );
  NAND2X0 U7135 ( .IN1(WX1837), .IN2(n3040), .QN(n5481) );
  NAND2X0 U7136 ( .IN1(n3053), .IN2(CRC_OUT_8_0), .QN(n5480) );
  NAND4X0 U7137 ( .IN1(n5486), .IN2(n5487), .IN3(n5488), .IN4(n5489), .QN(
        WX1997) );
  NAND2X0 U7138 ( .IN1(n3085), .IN2(n5267), .QN(n5489) );
  XNOR3X1 U7139 ( .IN1(n2899), .IN2(n2648), .IN3(n5490), .Q(n5267) );
  XOR2X1 U7140 ( .IN1(WX3355), .IN2(n6135), .Q(n5490) );
  NAND2X0 U7141 ( .IN1(n3012), .IN2(n4594), .QN(n5488) );
  XNOR3X1 U7142 ( .IN1(n2925), .IN2(n2663), .IN3(n5491), .Q(n4594) );
  XOR2X1 U7143 ( .IN1(WX2062), .IN2(n6136), .Q(n5491) );
  NAND2X0 U7144 ( .IN1(WX1835), .IN2(n3040), .QN(n5487) );
  NAND2X0 U7145 ( .IN1(n3053), .IN2(CRC_OUT_8_1), .QN(n5486) );
  NAND4X0 U7146 ( .IN1(n5492), .IN2(n5493), .IN3(n5494), .IN4(n5495), .QN(
        WX1995) );
  NAND2X0 U7147 ( .IN1(n3085), .IN2(n5273), .QN(n5495) );
  XNOR3X1 U7148 ( .IN1(n2898), .IN2(n2649), .IN3(n5496), .Q(n5273) );
  XOR2X1 U7149 ( .IN1(WX3353), .IN2(n6137), .Q(n5496) );
  NAND2X0 U7150 ( .IN1(n3012), .IN2(n4600), .QN(n5494) );
  XNOR3X1 U7151 ( .IN1(n2924), .IN2(n2664), .IN3(n5497), .Q(n4600) );
  XOR2X1 U7152 ( .IN1(WX2060), .IN2(n6138), .Q(n5497) );
  NAND2X0 U7153 ( .IN1(WX1833), .IN2(n3040), .QN(n5493) );
  NAND2X0 U7154 ( .IN1(n3053), .IN2(CRC_OUT_8_2), .QN(n5492) );
  NAND4X0 U7155 ( .IN1(n5498), .IN2(n5499), .IN3(n5500), .IN4(n5501), .QN(
        WX1993) );
  NAND2X0 U7156 ( .IN1(n3085), .IN2(n5279), .QN(n5501) );
  XNOR3X1 U7157 ( .IN1(n2897), .IN2(n2650), .IN3(n5502), .Q(n5279) );
  XOR2X1 U7158 ( .IN1(WX3351), .IN2(n6139), .Q(n5502) );
  NAND2X0 U7159 ( .IN1(n3012), .IN2(n4606), .QN(n5500) );
  XNOR3X1 U7160 ( .IN1(n2923), .IN2(n2665), .IN3(n5503), .Q(n4606) );
  XOR2X1 U7161 ( .IN1(WX2058), .IN2(n6140), .Q(n5503) );
  NAND2X0 U7162 ( .IN1(WX1831), .IN2(n3041), .QN(n5499) );
  NAND2X0 U7163 ( .IN1(n3053), .IN2(CRC_OUT_8_3), .QN(n5498) );
  NAND4X0 U7164 ( .IN1(n5504), .IN2(n5505), .IN3(n5506), .IN4(n5507), .QN(
        WX1991) );
  NAND2X0 U7165 ( .IN1(n3085), .IN2(n5285), .QN(n5507) );
  XNOR3X1 U7166 ( .IN1(n2702), .IN2(n2651), .IN3(n5508), .Q(n5285) );
  XOR2X1 U7167 ( .IN1(WX3349), .IN2(n6141), .Q(n5508) );
  NAND2X0 U7168 ( .IN1(n4612), .IN2(n3016), .QN(n5506) );
  XOR3X1 U7169 ( .IN1(n3763), .IN2(n2705), .IN3(n5509), .Q(n4612) );
  XOR2X1 U7170 ( .IN1(WX2120), .IN2(test_so14), .Q(n5509) );
  NAND2X0 U7171 ( .IN1(WX1829), .IN2(n3041), .QN(n5505) );
  NAND2X0 U7172 ( .IN1(n3053), .IN2(CRC_OUT_8_4), .QN(n5504) );
  NAND4X0 U7173 ( .IN1(n5510), .IN2(n5511), .IN3(n5512), .IN4(n5513), .QN(
        WX1989) );
  NAND2X0 U7174 ( .IN1(n3085), .IN2(n5291), .QN(n5513) );
  XNOR3X1 U7175 ( .IN1(n2896), .IN2(n2652), .IN3(n5514), .Q(n5291) );
  XOR2X1 U7176 ( .IN1(WX3347), .IN2(n6142), .Q(n5514) );
  NAND2X0 U7177 ( .IN1(n3012), .IN2(n4618), .QN(n5512) );
  XNOR3X1 U7178 ( .IN1(n2922), .IN2(n2666), .IN3(n5515), .Q(n4618) );
  XOR2X1 U7179 ( .IN1(WX2054), .IN2(n6143), .Q(n5515) );
  NAND2X0 U7180 ( .IN1(WX1827), .IN2(n3041), .QN(n5511) );
  NAND2X0 U7181 ( .IN1(n3054), .IN2(CRC_OUT_8_5), .QN(n5510) );
  NAND4X0 U7182 ( .IN1(n5516), .IN2(n5517), .IN3(n5518), .IN4(n5519), .QN(
        WX1987) );
  NAND2X0 U7183 ( .IN1(n5297), .IN2(n3098), .QN(n5519) );
  XOR3X1 U7184 ( .IN1(n3735), .IN2(n2653), .IN3(n5520), .Q(n5297) );
  XOR2X1 U7185 ( .IN1(WX3281), .IN2(test_so30), .Q(n5520) );
  NAND2X0 U7186 ( .IN1(n3012), .IN2(n4624), .QN(n5518) );
  XNOR3X1 U7187 ( .IN1(n2921), .IN2(n2667), .IN3(n5521), .Q(n4624) );
  XOR2X1 U7188 ( .IN1(WX2052), .IN2(n6144), .Q(n5521) );
  NAND2X0 U7189 ( .IN1(WX1825), .IN2(n3041), .QN(n5517) );
  NAND2X0 U7190 ( .IN1(n3054), .IN2(CRC_OUT_8_6), .QN(n5516) );
  NAND4X0 U7191 ( .IN1(n5522), .IN2(n5523), .IN3(n5524), .IN4(n5525), .QN(
        WX1985) );
  NAND2X0 U7192 ( .IN1(n3085), .IN2(n5303), .QN(n5525) );
  XNOR3X1 U7193 ( .IN1(n2895), .IN2(n2654), .IN3(n5526), .Q(n5303) );
  XOR2X1 U7194 ( .IN1(WX3343), .IN2(n6145), .Q(n5526) );
  NAND2X0 U7195 ( .IN1(n3011), .IN2(n4630), .QN(n5524) );
  XNOR3X1 U7196 ( .IN1(n2920), .IN2(n2668), .IN3(n5527), .Q(n4630) );
  XOR2X1 U7197 ( .IN1(WX2050), .IN2(n6146), .Q(n5527) );
  NAND2X0 U7198 ( .IN1(WX1823), .IN2(n3041), .QN(n5523) );
  NAND2X0 U7199 ( .IN1(test_so20), .IN2(n3070), .QN(n5522) );
  NAND4X0 U7200 ( .IN1(n5528), .IN2(n5529), .IN3(n5530), .IN4(n5531), .QN(
        WX1983) );
  NAND2X0 U7201 ( .IN1(n5309), .IN2(n3097), .QN(n5531) );
  XOR3X1 U7202 ( .IN1(n3739), .IN2(n2894), .IN3(n5532), .Q(n5309) );
  XOR2X1 U7203 ( .IN1(WX3277), .IN2(test_so28), .Q(n5532) );
  NAND2X0 U7204 ( .IN1(n3011), .IN2(n4636), .QN(n5530) );
  XNOR3X1 U7205 ( .IN1(n2919), .IN2(n2669), .IN3(n5533), .Q(n4636) );
  XOR2X1 U7206 ( .IN1(WX2048), .IN2(n6147), .Q(n5533) );
  NAND2X0 U7207 ( .IN1(WX1821), .IN2(n3041), .QN(n5529) );
  NAND2X0 U7208 ( .IN1(n3054), .IN2(CRC_OUT_8_8), .QN(n5528) );
  NAND4X0 U7209 ( .IN1(n5534), .IN2(n5535), .IN3(n5536), .IN4(n5537), .QN(
        WX1981) );
  NAND2X0 U7210 ( .IN1(n3085), .IN2(n5315), .QN(n5537) );
  XNOR3X1 U7211 ( .IN1(n2893), .IN2(n2655), .IN3(n5538), .Q(n5315) );
  XOR2X1 U7212 ( .IN1(WX3339), .IN2(n6148), .Q(n5538) );
  NAND2X0 U7213 ( .IN1(n3011), .IN2(n4642), .QN(n5536) );
  XNOR3X1 U7214 ( .IN1(n2918), .IN2(n2670), .IN3(n5539), .Q(n4642) );
  XOR2X1 U7215 ( .IN1(WX2046), .IN2(n6149), .Q(n5539) );
  NAND2X0 U7216 ( .IN1(WX1819), .IN2(n3041), .QN(n5535) );
  NAND2X0 U7217 ( .IN1(n3054), .IN2(CRC_OUT_8_9), .QN(n5534) );
  NAND4X0 U7218 ( .IN1(n5540), .IN2(n5541), .IN3(n5542), .IN4(n5543), .QN(
        WX1979) );
  NAND2X0 U7219 ( .IN1(n3085), .IN2(n5321), .QN(n5543) );
  XNOR3X1 U7220 ( .IN1(n2892), .IN2(n2656), .IN3(n5544), .Q(n5321) );
  XOR2X1 U7221 ( .IN1(WX3337), .IN2(n6150), .Q(n5544) );
  NAND2X0 U7222 ( .IN1(n4648), .IN2(n3017), .QN(n5542) );
  XOR3X1 U7223 ( .IN1(n3775), .IN2(n2671), .IN3(n5545), .Q(n4648) );
  XOR2X1 U7224 ( .IN1(WX1980), .IN2(test_so19), .Q(n5545) );
  NAND2X0 U7225 ( .IN1(WX1817), .IN2(n3041), .QN(n5541) );
  NAND2X0 U7226 ( .IN1(n3054), .IN2(CRC_OUT_8_10), .QN(n5540) );
  NAND4X0 U7227 ( .IN1(n5546), .IN2(n5547), .IN3(n5548), .IN4(n5549), .QN(
        WX1977) );
  NAND2X0 U7228 ( .IN1(n3086), .IN2(n5327), .QN(n5549) );
  XNOR3X1 U7229 ( .IN1(n2701), .IN2(n2657), .IN3(n5550), .Q(n5327) );
  XOR2X1 U7230 ( .IN1(WX3335), .IN2(n6151), .Q(n5550) );
  NAND2X0 U7231 ( .IN1(n3011), .IN2(n4654), .QN(n5548) );
  XNOR3X1 U7232 ( .IN1(n2704), .IN2(n2672), .IN3(n5551), .Q(n4654) );
  XOR2X1 U7233 ( .IN1(WX2042), .IN2(n6152), .Q(n5551) );
  NAND2X0 U7234 ( .IN1(WX1815), .IN2(n3041), .QN(n5547) );
  NAND2X0 U7235 ( .IN1(n3054), .IN2(CRC_OUT_8_11), .QN(n5546) );
  NAND4X0 U7236 ( .IN1(n5552), .IN2(n5553), .IN3(n5554), .IN4(n5555), .QN(
        WX1975) );
  NAND2X0 U7237 ( .IN1(n5333), .IN2(n3097), .QN(n5555) );
  XOR3X1 U7238 ( .IN1(n2891), .IN2(n2658), .IN3(n5556), .Q(n5333) );
  XOR2X1 U7239 ( .IN1(WX3269), .IN2(test_so26), .Q(n5556) );
  NAND2X0 U7240 ( .IN1(n3011), .IN2(n4660), .QN(n5554) );
  XNOR3X1 U7241 ( .IN1(n2917), .IN2(n2673), .IN3(n5557), .Q(n4660) );
  XOR2X1 U7242 ( .IN1(WX2040), .IN2(n6153), .Q(n5557) );
  NAND2X0 U7243 ( .IN1(WX1813), .IN2(n3041), .QN(n5553) );
  NAND2X0 U7244 ( .IN1(n3054), .IN2(CRC_OUT_8_12), .QN(n5552) );
  NAND4X0 U7245 ( .IN1(n5558), .IN2(n5559), .IN3(n5560), .IN4(n5561), .QN(
        WX1973) );
  NAND2X0 U7246 ( .IN1(n3086), .IN2(n5339), .QN(n5561) );
  XNOR3X1 U7247 ( .IN1(n2890), .IN2(n2659), .IN3(n5562), .Q(n5339) );
  XOR2X1 U7248 ( .IN1(WX3331), .IN2(n6154), .Q(n5562) );
  NAND2X0 U7249 ( .IN1(n3011), .IN2(n4666), .QN(n5560) );
  XNOR3X1 U7250 ( .IN1(n2916), .IN2(n2674), .IN3(n5563), .Q(n4666) );
  XOR2X1 U7251 ( .IN1(WX2038), .IN2(n6155), .Q(n5563) );
  NAND2X0 U7252 ( .IN1(WX1811), .IN2(n3041), .QN(n5559) );
  NAND2X0 U7253 ( .IN1(n3054), .IN2(CRC_OUT_8_13), .QN(n5558) );
  NAND4X0 U7254 ( .IN1(n5564), .IN2(n5565), .IN3(n5566), .IN4(n5567), .QN(
        WX1971) );
  NAND2X0 U7255 ( .IN1(n3086), .IN2(n5345), .QN(n5567) );
  XNOR3X1 U7256 ( .IN1(n2889), .IN2(n2660), .IN3(n5568), .Q(n5345) );
  XOR2X1 U7257 ( .IN1(WX3329), .IN2(n6156), .Q(n5568) );
  NAND2X0 U7258 ( .IN1(n4672), .IN2(n3016), .QN(n5566) );
  XOR3X1 U7259 ( .IN1(n3783), .IN2(n2915), .IN3(n5569), .Q(n4672) );
  XOR2X1 U7260 ( .IN1(WX1972), .IN2(test_so17), .Q(n5569) );
  NAND2X0 U7261 ( .IN1(WX1809), .IN2(n3041), .QN(n5565) );
  NAND2X0 U7262 ( .IN1(n3054), .IN2(CRC_OUT_8_14), .QN(n5564) );
  NAND4X0 U7263 ( .IN1(n5570), .IN2(n5571), .IN3(n5572), .IN4(n5573), .QN(
        WX1969) );
  NAND2X0 U7264 ( .IN1(n3086), .IN2(n5351), .QN(n5573) );
  XNOR3X1 U7265 ( .IN1(n2888), .IN2(n2661), .IN3(n5574), .Q(n5351) );
  XOR2X1 U7266 ( .IN1(WX3327), .IN2(n6157), .Q(n5574) );
  NAND2X0 U7267 ( .IN1(n3011), .IN2(n4678), .QN(n5572) );
  XNOR3X1 U7268 ( .IN1(n2914), .IN2(n2675), .IN3(n5575), .Q(n4678) );
  XOR2X1 U7269 ( .IN1(WX2034), .IN2(n6158), .Q(n5575) );
  NAND2X0 U7270 ( .IN1(WX1807), .IN2(n3041), .QN(n5571) );
  NAND2X0 U7271 ( .IN1(n3054), .IN2(CRC_OUT_8_15), .QN(n5570) );
  NAND4X0 U7272 ( .IN1(n5576), .IN2(n5577), .IN3(n5578), .IN4(n5579), .QN(
        WX1967) );
  NAND2X0 U7273 ( .IN1(n5357), .IN2(n3097), .QN(n5579) );
  XOR3X1 U7274 ( .IN1(n2509), .IN2(n3578), .IN3(n5580), .Q(n5357) );
  XNOR3X1 U7275 ( .IN1(test_so24), .IN2(n6159), .IN3(n2700), .Q(n5580) );
  NAND2X0 U7276 ( .IN1(n3011), .IN2(n4684), .QN(n5578) );
  XNOR3X1 U7277 ( .IN1(n2535), .IN2(n3573), .IN3(n5581), .Q(n4684) );
  XOR3X1 U7278 ( .IN1(n6160), .IN2(n2703), .IN3(WX2096), .Q(n5581) );
  NAND2X0 U7279 ( .IN1(WX1805), .IN2(n3041), .QN(n5577) );
  NAND2X0 U7280 ( .IN1(n3054), .IN2(CRC_OUT_8_16), .QN(n5576) );
  NAND4X0 U7281 ( .IN1(n5582), .IN2(n5583), .IN3(n5584), .IN4(n5585), .QN(
        WX1965) );
  NAND2X0 U7282 ( .IN1(n3086), .IN2(n5363), .QN(n5585) );
  XNOR3X1 U7283 ( .IN1(n2510), .IN2(n3573), .IN3(n5586), .Q(n5363) );
  XOR3X1 U7284 ( .IN1(n6161), .IN2(n2887), .IN3(WX3387), .Q(n5586) );
  NAND2X0 U7285 ( .IN1(n3011), .IN2(n4690), .QN(n5584) );
  XNOR3X1 U7286 ( .IN1(n2537), .IN2(n3573), .IN3(n5587), .Q(n4690) );
  XOR3X1 U7287 ( .IN1(n6162), .IN2(n2913), .IN3(WX2094), .Q(n5587) );
  NAND2X0 U7288 ( .IN1(WX1803), .IN2(n3041), .QN(n5583) );
  NAND2X0 U7289 ( .IN1(n3054), .IN2(CRC_OUT_8_17), .QN(n5582) );
  NAND4X0 U7290 ( .IN1(n5588), .IN2(n5589), .IN3(n5590), .IN4(n5591), .QN(
        WX1963) );
  NAND2X0 U7291 ( .IN1(n3086), .IN2(n5369), .QN(n5591) );
  XNOR3X1 U7292 ( .IN1(n2512), .IN2(n3573), .IN3(n5592), .Q(n5369) );
  XOR3X1 U7293 ( .IN1(n6163), .IN2(n2886), .IN3(WX3385), .Q(n5592) );
  NAND2X0 U7294 ( .IN1(n4696), .IN2(n3017), .QN(n5590) );
  XOR3X1 U7295 ( .IN1(n2539), .IN2(n3577), .IN3(n5593), .Q(n4696) );
  XNOR3X1 U7296 ( .IN1(test_so15), .IN2(n6164), .IN3(n2912), .Q(n5593) );
  NAND2X0 U7297 ( .IN1(WX1801), .IN2(n3041), .QN(n5589) );
  NAND2X0 U7298 ( .IN1(n3055), .IN2(CRC_OUT_8_18), .QN(n5588) );
  NAND4X0 U7299 ( .IN1(n5594), .IN2(n5595), .IN3(n5596), .IN4(n5597), .QN(
        WX1961) );
  NAND2X0 U7300 ( .IN1(n3086), .IN2(n5375), .QN(n5597) );
  XNOR3X1 U7301 ( .IN1(n2514), .IN2(n3573), .IN3(n5598), .Q(n5375) );
  XOR3X1 U7302 ( .IN1(n6165), .IN2(n2885), .IN3(WX3383), .Q(n5598) );
  NAND2X0 U7303 ( .IN1(n3011), .IN2(n4702), .QN(n5596) );
  XNOR3X1 U7304 ( .IN1(n2540), .IN2(n3573), .IN3(n5599), .Q(n4702) );
  XOR3X1 U7305 ( .IN1(n6166), .IN2(n2911), .IN3(WX2090), .Q(n5599) );
  NAND2X0 U7306 ( .IN1(WX1799), .IN2(n3041), .QN(n5595) );
  NAND2X0 U7307 ( .IN1(n3055), .IN2(CRC_OUT_8_19), .QN(n5594) );
  NAND4X0 U7308 ( .IN1(n5600), .IN2(n5601), .IN3(n5602), .IN4(n5603), .QN(
        WX1959) );
  NAND2X0 U7309 ( .IN1(n3086), .IN2(n5381), .QN(n5603) );
  XNOR3X1 U7310 ( .IN1(n2516), .IN2(n3573), .IN3(n5604), .Q(n5381) );
  XOR3X1 U7311 ( .IN1(n6167), .IN2(n2884), .IN3(WX3381), .Q(n5604) );
  NAND2X0 U7312 ( .IN1(n3011), .IN2(n4708), .QN(n5602) );
  XNOR3X1 U7313 ( .IN1(n2542), .IN2(n3573), .IN3(n5605), .Q(n4708) );
  XOR3X1 U7314 ( .IN1(n6168), .IN2(n2910), .IN3(WX2088), .Q(n5605) );
  NAND2X0 U7315 ( .IN1(WX1797), .IN2(n3042), .QN(n5601) );
  NAND2X0 U7316 ( .IN1(n3055), .IN2(CRC_OUT_8_20), .QN(n5600) );
  NAND4X0 U7317 ( .IN1(n5606), .IN2(n5607), .IN3(n5608), .IN4(n5609), .QN(
        WX1957) );
  NAND2X0 U7318 ( .IN1(n3086), .IN2(n5387), .QN(n5609) );
  XNOR3X1 U7319 ( .IN1(n2518), .IN2(n3573), .IN3(n5610), .Q(n5387) );
  XOR3X1 U7320 ( .IN1(n6169), .IN2(n2883), .IN3(WX3379), .Q(n5610) );
  NAND2X0 U7321 ( .IN1(n3011), .IN2(n4714), .QN(n5608) );
  XNOR3X1 U7322 ( .IN1(n2544), .IN2(n3573), .IN3(n5611), .Q(n4714) );
  XOR3X1 U7323 ( .IN1(n6170), .IN2(n2909), .IN3(WX2086), .Q(n5611) );
  NAND2X0 U7324 ( .IN1(WX1795), .IN2(n3042), .QN(n5607) );
  NAND2X0 U7325 ( .IN1(n3055), .IN2(CRC_OUT_8_21), .QN(n5606) );
  NAND4X0 U7326 ( .IN1(n5612), .IN2(n5613), .IN3(n5614), .IN4(n5615), .QN(
        WX1955) );
  NAND2X0 U7327 ( .IN1(n3086), .IN2(n5393), .QN(n5615) );
  XNOR3X1 U7328 ( .IN1(n2520), .IN2(n3574), .IN3(n5616), .Q(n5393) );
  XOR3X1 U7329 ( .IN1(n6171), .IN2(n2882), .IN3(WX3377), .Q(n5616) );
  NAND2X0 U7330 ( .IN1(n4720), .IN2(n3017), .QN(n5614) );
  XOR3X1 U7331 ( .IN1(n2546), .IN2(n3577), .IN3(n5617), .Q(n4720) );
  XNOR3X1 U7332 ( .IN1(test_so13), .IN2(n6172), .IN3(n2908), .Q(n5617) );
  NAND2X0 U7333 ( .IN1(WX1793), .IN2(n3042), .QN(n5613) );
  NAND2X0 U7334 ( .IN1(n3055), .IN2(CRC_OUT_8_22), .QN(n5612) );
  NAND4X0 U7335 ( .IN1(n5618), .IN2(n5619), .IN3(n5620), .IN4(n5621), .QN(
        WX1953) );
  NAND2X0 U7336 ( .IN1(n5399), .IN2(n3097), .QN(n5621) );
  XOR3X1 U7337 ( .IN1(n2522), .IN2(n3577), .IN3(n5622), .Q(n5399) );
  XOR3X1 U7338 ( .IN1(test_so29), .IN2(n6173), .IN3(WX3375), .Q(n5622) );
  NAND2X0 U7339 ( .IN1(n3010), .IN2(n4726), .QN(n5620) );
  XNOR3X1 U7340 ( .IN1(n2547), .IN2(n3574), .IN3(n5623), .Q(n4726) );
  XOR3X1 U7341 ( .IN1(n6174), .IN2(n2907), .IN3(WX2082), .Q(n5623) );
  NAND2X0 U7342 ( .IN1(WX1791), .IN2(n3042), .QN(n5619) );
  NAND2X0 U7343 ( .IN1(n3055), .IN2(CRC_OUT_8_23), .QN(n5618) );
  NAND4X0 U7344 ( .IN1(n5624), .IN2(n5625), .IN3(n5626), .IN4(n5627), .QN(
        WX1951) );
  NAND2X0 U7345 ( .IN1(n3086), .IN2(n5405), .QN(n5627) );
  XNOR3X1 U7346 ( .IN1(n2523), .IN2(n3574), .IN3(n5628), .Q(n5405) );
  XOR3X1 U7347 ( .IN1(n6175), .IN2(n2881), .IN3(WX3373), .Q(n5628) );
  NAND2X0 U7348 ( .IN1(n3010), .IN2(n4732), .QN(n5626) );
  XNOR3X1 U7349 ( .IN1(n2549), .IN2(n3574), .IN3(n5629), .Q(n4732) );
  XOR3X1 U7350 ( .IN1(n6176), .IN2(n2906), .IN3(WX2080), .Q(n5629) );
  NAND2X0 U7351 ( .IN1(WX1789), .IN2(n3042), .QN(n5625) );
  NAND2X0 U7352 ( .IN1(n3055), .IN2(CRC_OUT_8_24), .QN(n5624) );
  NAND4X0 U7353 ( .IN1(n5630), .IN2(n5631), .IN3(n5632), .IN4(n5633), .QN(
        WX1949) );
  NAND2X0 U7354 ( .IN1(n3086), .IN2(n5411), .QN(n5633) );
  XNOR3X1 U7355 ( .IN1(n2525), .IN2(n3574), .IN3(n5634), .Q(n5411) );
  XOR3X1 U7356 ( .IN1(n6177), .IN2(n2880), .IN3(WX3371), .Q(n5634) );
  NAND2X0 U7357 ( .IN1(n3010), .IN2(n4738), .QN(n5632) );
  XNOR3X1 U7358 ( .IN1(n2551), .IN2(n3574), .IN3(n5635), .Q(n4738) );
  XOR3X1 U7359 ( .IN1(n6178), .IN2(n2905), .IN3(WX2078), .Q(n5635) );
  NAND2X0 U7360 ( .IN1(WX1787), .IN2(n3042), .QN(n5631) );
  NAND2X0 U7361 ( .IN1(test_so21), .IN2(n3070), .QN(n5630) );
  NAND4X0 U7362 ( .IN1(n5636), .IN2(n5637), .IN3(n5638), .IN4(n5639), .QN(
        WX1947) );
  NAND2X0 U7363 ( .IN1(n5417), .IN2(n3096), .QN(n5639) );
  XOR3X1 U7364 ( .IN1(n2527), .IN2(n3578), .IN3(n5640), .Q(n5417) );
  XNOR3X1 U7365 ( .IN1(test_so27), .IN2(n6179), .IN3(n2879), .Q(n5640) );
  NAND2X0 U7366 ( .IN1(n3010), .IN2(n4744), .QN(n5638) );
  XNOR3X1 U7367 ( .IN1(n2553), .IN2(n3574), .IN3(n5641), .Q(n4744) );
  XOR3X1 U7368 ( .IN1(n6180), .IN2(n2904), .IN3(WX2076), .Q(n5641) );
  NAND2X0 U7369 ( .IN1(WX1785), .IN2(n3042), .QN(n5637) );
  NAND2X0 U7370 ( .IN1(n3055), .IN2(CRC_OUT_8_26), .QN(n5636) );
  NAND4X0 U7371 ( .IN1(n5642), .IN2(n5643), .IN3(n5644), .IN4(n5645), .QN(
        WX1945) );
  NAND2X0 U7372 ( .IN1(n3087), .IN2(n5423), .QN(n5645) );
  XNOR3X1 U7373 ( .IN1(n2528), .IN2(n3574), .IN3(n5646), .Q(n5423) );
  XOR3X1 U7374 ( .IN1(n6181), .IN2(n2878), .IN3(WX3367), .Q(n5646) );
  NAND2X0 U7375 ( .IN1(n3010), .IN2(n4750), .QN(n5644) );
  XNOR3X1 U7376 ( .IN1(n2555), .IN2(n3574), .IN3(n5647), .Q(n4750) );
  XOR3X1 U7377 ( .IN1(n6182), .IN2(n2903), .IN3(WX2074), .Q(n5647) );
  NAND2X0 U7378 ( .IN1(WX1783), .IN2(n3042), .QN(n5643) );
  NAND2X0 U7379 ( .IN1(n3055), .IN2(CRC_OUT_8_27), .QN(n5642) );
  NAND4X0 U7380 ( .IN1(n5648), .IN2(n5649), .IN3(n5650), .IN4(n5651), .QN(
        WX1943) );
  NAND2X0 U7381 ( .IN1(n3087), .IN2(n5429), .QN(n5651) );
  XNOR3X1 U7382 ( .IN1(n2530), .IN2(n3574), .IN3(n5652), .Q(n5429) );
  XOR3X1 U7383 ( .IN1(n6183), .IN2(n2877), .IN3(WX3365), .Q(n5652) );
  NAND2X0 U7384 ( .IN1(n4756), .IN2(n3018), .QN(n5650) );
  XOR3X1 U7385 ( .IN1(n2557), .IN2(n3578), .IN3(n5653), .Q(n4756) );
  XOR3X1 U7386 ( .IN1(test_so18), .IN2(n6184), .IN3(WX2072), .Q(n5653) );
  NAND2X0 U7387 ( .IN1(WX1781), .IN2(n3042), .QN(n5649) );
  NAND2X0 U7388 ( .IN1(n3055), .IN2(CRC_OUT_8_28), .QN(n5648) );
  NAND4X0 U7389 ( .IN1(n5654), .IN2(n5655), .IN3(n5656), .IN4(n5657), .QN(
        WX1941) );
  NAND2X0 U7390 ( .IN1(n3087), .IN2(n5435), .QN(n5657) );
  XNOR3X1 U7391 ( .IN1(n2532), .IN2(n3575), .IN3(n5658), .Q(n5435) );
  XOR3X1 U7392 ( .IN1(n6185), .IN2(n2876), .IN3(WX3363), .Q(n5658) );
  NAND2X0 U7393 ( .IN1(n3010), .IN2(n4772), .QN(n5656) );
  XNOR3X1 U7394 ( .IN1(n2558), .IN2(n3575), .IN3(n5659), .Q(n4772) );
  XOR3X1 U7395 ( .IN1(n6186), .IN2(n2902), .IN3(WX2070), .Q(n5659) );
  NAND2X0 U7396 ( .IN1(WX1779), .IN2(n3042), .QN(n5655) );
  NAND2X0 U7397 ( .IN1(n3055), .IN2(CRC_OUT_8_29), .QN(n5654) );
  NAND4X0 U7398 ( .IN1(n5660), .IN2(n5661), .IN3(n5662), .IN4(n5663), .QN(
        WX1939) );
  NAND2X0 U7399 ( .IN1(n5441), .IN2(n3096), .QN(n5663) );
  XOR3X1 U7400 ( .IN1(n2534), .IN2(n3578), .IN3(n5664), .Q(n5441) );
  XNOR3X1 U7401 ( .IN1(test_so25), .IN2(n6187), .IN3(n2875), .Q(n5664) );
  NAND2X0 U7402 ( .IN1(n3010), .IN2(n4788), .QN(n5662) );
  XNOR3X1 U7403 ( .IN1(n2560), .IN2(n3575), .IN3(n5665), .Q(n4788) );
  XOR3X1 U7404 ( .IN1(n6188), .IN2(n2901), .IN3(WX2068), .Q(n5665) );
  NAND2X0 U7405 ( .IN1(WX1777), .IN2(n3042), .QN(n5661) );
  NAND2X0 U7406 ( .IN1(n3055), .IN2(CRC_OUT_8_30), .QN(n5660) );
  NAND4X0 U7407 ( .IN1(n5666), .IN2(n5667), .IN3(n5668), .IN4(n5669), .QN(
        WX1937) );
  NAND2X0 U7408 ( .IN1(n3010), .IN2(n4804), .QN(n5669) );
  XNOR3X1 U7409 ( .IN1(n2348), .IN2(n3575), .IN3(n5670), .Q(n4804) );
  XOR3X1 U7410 ( .IN1(n6189), .IN2(n2900), .IN3(WX2066), .Q(n5670) );
  NAND2X0 U7411 ( .IN1(n3087), .IN2(n5447), .QN(n5668) );
  XNOR3X1 U7412 ( .IN1(n2346), .IN2(n3574), .IN3(n5671), .Q(n5447) );
  XOR3X1 U7413 ( .IN1(n6190), .IN2(n2874), .IN3(WX3359), .Q(n5671) );
  NAND2X0 U7414 ( .IN1(n3056), .IN2(CRC_OUT_8_31), .QN(n5667) );
  NAND2X0 U7415 ( .IN1(n2245), .IN2(WX1778), .QN(n5666) );
  NOR2X0 U7416 ( .IN1(n3736), .IN2(WX1778), .QN(WX1839) );
  AND2X1 U7417 ( .IN1(n3606), .IN2(n8670), .Q(WX1837) );
  AND2X1 U7418 ( .IN1(n3606), .IN2(n8671), .Q(WX1835) );
  AND2X1 U7419 ( .IN1(n3606), .IN2(n8672), .Q(WX1833) );
  AND2X1 U7420 ( .IN1(n3606), .IN2(n8673), .Q(WX1831) );
  AND2X1 U7421 ( .IN1(n3606), .IN2(n8674), .Q(WX1829) );
  AND2X1 U7422 ( .IN1(n3606), .IN2(n8675), .Q(WX1827) );
  AND2X1 U7423 ( .IN1(n3606), .IN2(n8676), .Q(WX1825) );
  AND2X1 U7424 ( .IN1(n3606), .IN2(n8677), .Q(WX1823) );
  AND2X1 U7425 ( .IN1(test_so12), .IN2(n3599), .Q(WX1821) );
  AND2X1 U7426 ( .IN1(n3607), .IN2(n8680), .Q(WX1819) );
  AND2X1 U7427 ( .IN1(n3607), .IN2(n8681), .Q(WX1817) );
  AND2X1 U7428 ( .IN1(n3607), .IN2(n8682), .Q(WX1815) );
  AND2X1 U7429 ( .IN1(n3607), .IN2(n8683), .Q(WX1813) );
  AND2X1 U7430 ( .IN1(n3607), .IN2(n8684), .Q(WX1811) );
  AND2X1 U7431 ( .IN1(n3607), .IN2(n8685), .Q(WX1809) );
  AND2X1 U7432 ( .IN1(n3607), .IN2(n8686), .Q(WX1807) );
  AND2X1 U7433 ( .IN1(n3607), .IN2(n8687), .Q(WX1805) );
  AND2X1 U7434 ( .IN1(n3607), .IN2(n8688), .Q(WX1803) );
  AND2X1 U7435 ( .IN1(n3608), .IN2(n8689), .Q(WX1801) );
  AND2X1 U7436 ( .IN1(n3608), .IN2(n8690), .Q(WX1799) );
  AND2X1 U7437 ( .IN1(n3608), .IN2(n8691), .Q(WX1797) );
  AND2X1 U7438 ( .IN1(n3608), .IN2(n8692), .Q(WX1795) );
  AND2X1 U7439 ( .IN1(n3608), .IN2(n8693), .Q(WX1793) );
  AND2X1 U7440 ( .IN1(n3608), .IN2(n8694), .Q(WX1791) );
  AND2X1 U7441 ( .IN1(n3608), .IN2(n8695), .Q(WX1789) );
  AND2X1 U7442 ( .IN1(n3608), .IN2(n8696), .Q(WX1787) );
  AND2X1 U7443 ( .IN1(test_so11), .IN2(n3599), .Q(WX1785) );
  AND2X1 U7444 ( .IN1(n3608), .IN2(n8699), .Q(WX1783) );
  AND2X1 U7445 ( .IN1(n3609), .IN2(n8700), .Q(WX1781) );
  AND2X1 U7446 ( .IN1(n3609), .IN2(n8701), .Q(WX1779) );
  AND2X1 U7447 ( .IN1(n3609), .IN2(n8702), .Q(WX1777) );
  NOR2X0 U7448 ( .IN1(n3736), .IN2(n5672), .QN(WX1326) );
  XOR2X1 U7449 ( .IN1(n2978), .IN2(DFF_190_n1), .Q(n5672) );
  NOR2X0 U7450 ( .IN1(n3736), .IN2(n5673), .QN(WX1324) );
  XOR2X1 U7451 ( .IN1(n2928), .IN2(DFF_189_n1), .Q(n5673) );
  NOR2X0 U7452 ( .IN1(n3736), .IN2(n5674), .QN(WX1322) );
  XOR2X1 U7453 ( .IN1(n2933), .IN2(DFF_188_n1), .Q(n5674) );
  NOR2X0 U7454 ( .IN1(n3736), .IN2(n5675), .QN(WX1320) );
  XOR2X1 U7455 ( .IN1(n2939), .IN2(DFF_187_n1), .Q(n5675) );
  NOR2X0 U7456 ( .IN1(n3736), .IN2(n5676), .QN(WX1318) );
  XOR2X1 U7457 ( .IN1(n2942), .IN2(DFF_186_n1), .Q(n5676) );
  NOR2X0 U7458 ( .IN1(n3737), .IN2(n5677), .QN(WX1316) );
  XOR2X1 U7459 ( .IN1(n2944), .IN2(DFF_185_n1), .Q(n5677) );
  NOR2X0 U7460 ( .IN1(n3737), .IN2(n5678), .QN(WX1314) );
  XOR2X1 U7461 ( .IN1(n2949), .IN2(DFF_184_n1), .Q(n5678) );
  NOR2X0 U7462 ( .IN1(n3737), .IN2(n5679), .QN(WX1312) );
  XOR2X1 U7463 ( .IN1(n2955), .IN2(DFF_183_n1), .Q(n5679) );
  NOR2X0 U7464 ( .IN1(n3736), .IN2(n5680), .QN(WX1310) );
  XOR2X1 U7465 ( .IN1(n2956), .IN2(DFF_182_n1), .Q(n5680) );
  NOR2X0 U7466 ( .IN1(n3737), .IN2(n5681), .QN(WX1308) );
  XOR2X1 U7467 ( .IN1(n2967), .IN2(DFF_181_n1), .Q(n5681) );
  NOR2X0 U7468 ( .IN1(n3737), .IN2(n5682), .QN(WX1306) );
  XOR2X1 U7469 ( .IN1(n2973), .IN2(DFF_180_n1), .Q(n5682) );
  NOR2X0 U7470 ( .IN1(n3737), .IN2(n5683), .QN(WX1304) );
  XNOR2X1 U7471 ( .IN1(n2976), .IN2(test_so10), .Q(n5683) );
  NOR2X0 U7472 ( .IN1(n3737), .IN2(n5684), .QN(WX1302) );
  XOR2X1 U7473 ( .IN1(n2931), .IN2(DFF_178_n1), .Q(n5684) );
  NOR2X0 U7474 ( .IN1(n3737), .IN2(n5685), .QN(WX1300) );
  XOR2X1 U7475 ( .IN1(n2940), .IN2(DFF_177_n1), .Q(n5685) );
  NOR2X0 U7476 ( .IN1(n3737), .IN2(n5686), .QN(WX1298) );
  XOR2X1 U7477 ( .IN1(n2947), .IN2(DFF_176_n1), .Q(n5686) );
  NOR2X0 U7478 ( .IN1(n3737), .IN2(n5687), .QN(WX1296) );
  XOR3X1 U7479 ( .IN1(test_so8), .IN2(DFF_191_n1), .IN3(DFF_175_n1), .Q(n5687)
         );
  NOR2X0 U7480 ( .IN1(n3737), .IN2(n5688), .QN(WX1294) );
  XOR2X1 U7481 ( .IN1(n2970), .IN2(DFF_174_n1), .Q(n5688) );
  NOR2X0 U7482 ( .IN1(n3738), .IN2(n5689), .QN(WX1292) );
  XOR2X1 U7483 ( .IN1(n2979), .IN2(DFF_173_n1), .Q(n5689) );
  NOR2X0 U7484 ( .IN1(n3738), .IN2(n5690), .QN(WX1290) );
  XOR2X1 U7485 ( .IN1(n2935), .IN2(DFF_172_n1), .Q(n5690) );
  NOR2X0 U7486 ( .IN1(n3738), .IN2(n5691), .QN(WX1288) );
  XOR2X1 U7487 ( .IN1(n2951), .IN2(DFF_171_n1), .Q(n5691) );
  NOR2X0 U7488 ( .IN1(n3738), .IN2(n5692), .QN(WX1286) );
  XOR3X1 U7489 ( .IN1(n2986), .IN2(DFF_191_n1), .IN3(CRC_OUT_9_10), .Q(n5692)
         );
  NOR2X0 U7490 ( .IN1(n3738), .IN2(n5693), .QN(WX1284) );
  XOR2X1 U7491 ( .IN1(n2946), .IN2(DFF_169_n1), .Q(n5693) );
  NOR2X0 U7492 ( .IN1(n3738), .IN2(n5694), .QN(WX1282) );
  XOR2X1 U7493 ( .IN1(n2954), .IN2(DFF_168_n1), .Q(n5694) );
  NOR2X0 U7494 ( .IN1(n3738), .IN2(n5695), .QN(WX1280) );
  XOR2X1 U7495 ( .IN1(n2959), .IN2(DFF_167_n1), .Q(n5695) );
  NOR2X0 U7496 ( .IN1(n3738), .IN2(n5696), .QN(WX1278) );
  XOR2X1 U7497 ( .IN1(n2985), .IN2(DFF_166_n1), .Q(n5696) );
  NOR2X0 U7498 ( .IN1(n3738), .IN2(n5697), .QN(WX1276) );
  XOR2X1 U7499 ( .IN1(n2975), .IN2(DFF_165_n1), .Q(n5697) );
  NOR2X0 U7500 ( .IN1(n3738), .IN2(n5698), .QN(WX1274) );
  XOR2X1 U7501 ( .IN1(n2961), .IN2(DFF_164_n1), .Q(n5698) );
  NOR2X0 U7502 ( .IN1(n3738), .IN2(n5699), .QN(WX1272) );
  XOR3X1 U7503 ( .IN1(n2963), .IN2(DFF_191_n1), .IN3(CRC_OUT_9_3), .Q(n5699)
         );
  NOR2X0 U7504 ( .IN1(n3738), .IN2(n5700), .QN(WX1270) );
  XOR2X1 U7505 ( .IN1(n2929), .IN2(DFF_162_n1), .Q(n5700) );
  NOR2X0 U7506 ( .IN1(n3738), .IN2(n5701), .QN(WX1268) );
  XNOR2X1 U7507 ( .IN1(n2982), .IN2(test_so9), .Q(n5701) );
  NOR2X0 U7508 ( .IN1(n3740), .IN2(n5702), .QN(WX1266) );
  XOR2X1 U7509 ( .IN1(n2937), .IN2(DFF_160_n1), .Q(n5702) );
  NOR2X0 U7510 ( .IN1(n3740), .IN2(n5703), .QN(WX1264) );
  XOR2X1 U7511 ( .IN1(n2990), .IN2(DFF_191_n1), .Q(n5703) );
  NOR2X0 U7512 ( .IN1(n3740), .IN2(n5704), .QN(WX11670) );
  XOR2X1 U7513 ( .IN1(n2714), .IN2(DFF_1726_n1), .Q(n5704) );
  NOR2X0 U7514 ( .IN1(n3740), .IN2(n5705), .QN(WX11668) );
  XOR2X1 U7515 ( .IN1(n2715), .IN2(DFF_1725_n1), .Q(n5705) );
  NOR2X0 U7516 ( .IN1(n3740), .IN2(n5706), .QN(WX11666) );
  XOR2X1 U7517 ( .IN1(n2716), .IN2(DFF_1724_n1), .Q(n5706) );
  NOR2X0 U7518 ( .IN1(n3740), .IN2(n5707), .QN(WX11664) );
  XOR2X1 U7519 ( .IN1(n2717), .IN2(DFF_1723_n1), .Q(n5707) );
  NOR2X0 U7520 ( .IN1(n3740), .IN2(n5708), .QN(WX11662) );
  XOR2X1 U7521 ( .IN1(n2718), .IN2(DFF_1722_n1), .Q(n5708) );
  NOR2X0 U7522 ( .IN1(n3740), .IN2(n5709), .QN(WX11660) );
  XOR2X1 U7523 ( .IN1(n2719), .IN2(DFF_1721_n1), .Q(n5709) );
  NOR2X0 U7524 ( .IN1(n3740), .IN2(n5710), .QN(WX11658) );
  XOR2X1 U7525 ( .IN1(n2720), .IN2(DFF_1720_n1), .Q(n5710) );
  NOR2X0 U7526 ( .IN1(n3740), .IN2(n5711), .QN(WX11656) );
  XOR2X1 U7527 ( .IN1(n2721), .IN2(DFF_1719_n1), .Q(n5711) );
  NOR2X0 U7528 ( .IN1(n3740), .IN2(n5712), .QN(WX11654) );
  XOR2X1 U7529 ( .IN1(n2722), .IN2(DFF_1718_n1), .Q(n5712) );
  NOR2X0 U7530 ( .IN1(n3740), .IN2(n5713), .QN(WX11652) );
  XOR2X1 U7531 ( .IN1(n2723), .IN2(DFF_1717_n1), .Q(n5713) );
  NOR2X0 U7532 ( .IN1(n3740), .IN2(n5714), .QN(WX11650) );
  XOR2X1 U7533 ( .IN1(n2724), .IN2(DFF_1716_n1), .Q(n5714) );
  NOR2X0 U7534 ( .IN1(n3741), .IN2(n5715), .QN(WX11648) );
  XOR2X1 U7535 ( .IN1(n2725), .IN2(DFF_1715_n1), .Q(n5715) );
  NOR2X0 U7536 ( .IN1(n3741), .IN2(n5716), .QN(WX11646) );
  XOR2X1 U7537 ( .IN1(CRC_OUT_1_18), .IN2(test_so97), .Q(n5716) );
  NOR2X0 U7538 ( .IN1(n3741), .IN2(n5717), .QN(WX11644) );
  XOR2X1 U7539 ( .IN1(n2726), .IN2(DFF_1713_n1), .Q(n5717) );
  NOR2X0 U7540 ( .IN1(n3741), .IN2(n5718), .QN(WX11642) );
  XOR2X1 U7541 ( .IN1(n2727), .IN2(DFF_1712_n1), .Q(n5718) );
  NOR2X0 U7542 ( .IN1(n3741), .IN2(n5719), .QN(WX11640) );
  XOR3X1 U7543 ( .IN1(test_so100), .IN2(n2685), .IN3(DFF_1711_n1), .Q(n5719)
         );
  NOR2X0 U7544 ( .IN1(n3741), .IN2(n5720), .QN(WX11638) );
  XNOR2X1 U7545 ( .IN1(n2728), .IN2(test_so99), .Q(n5720) );
  NOR2X0 U7546 ( .IN1(n3741), .IN2(n5721), .QN(WX11636) );
  XOR2X1 U7547 ( .IN1(n2729), .IN2(DFF_1709_n1), .Q(n5721) );
  NOR2X0 U7548 ( .IN1(n3741), .IN2(n5722), .QN(WX11634) );
  XOR2X1 U7549 ( .IN1(n2730), .IN2(DFF_1708_n1), .Q(n5722) );
  NOR2X0 U7550 ( .IN1(n3741), .IN2(n5723), .QN(WX11632) );
  XOR2X1 U7551 ( .IN1(n2731), .IN2(DFF_1707_n1), .Q(n5723) );
  NOR2X0 U7552 ( .IN1(n3741), .IN2(n5724), .QN(WX11630) );
  XOR3X1 U7553 ( .IN1(test_so100), .IN2(n2686), .IN3(DFF_1706_n1), .Q(n5724)
         );
  NOR2X0 U7554 ( .IN1(n3741), .IN2(n5725), .QN(WX11628) );
  XOR2X1 U7555 ( .IN1(n2732), .IN2(DFF_1705_n1), .Q(n5725) );
  NOR2X0 U7556 ( .IN1(n3741), .IN2(n5726), .QN(WX11626) );
  XOR2X1 U7557 ( .IN1(n2733), .IN2(DFF_1704_n1), .Q(n5726) );
  NOR2X0 U7558 ( .IN1(n3741), .IN2(n5727), .QN(WX11624) );
  XOR2X1 U7559 ( .IN1(n2734), .IN2(DFF_1703_n1), .Q(n5727) );
  NOR2X0 U7560 ( .IN1(n3742), .IN2(n5728), .QN(WX11622) );
  XOR2X1 U7561 ( .IN1(n2735), .IN2(DFF_1702_n1), .Q(n5728) );
  NOR2X0 U7562 ( .IN1(n3742), .IN2(n5729), .QN(WX11620) );
  XOR2X1 U7563 ( .IN1(n2736), .IN2(DFF_1701_n1), .Q(n5729) );
  NOR2X0 U7564 ( .IN1(n3742), .IN2(n5730), .QN(WX11618) );
  XOR2X1 U7565 ( .IN1(n2737), .IN2(DFF_1700_n1), .Q(n5730) );
  NOR2X0 U7566 ( .IN1(n3742), .IN2(n5731), .QN(WX11616) );
  XOR3X1 U7567 ( .IN1(test_so100), .IN2(n2687), .IN3(DFF_1699_n1), .Q(n5731)
         );
  NOR2X0 U7568 ( .IN1(n3742), .IN2(n5732), .QN(WX11614) );
  XOR2X1 U7569 ( .IN1(n2738), .IN2(DFF_1698_n1), .Q(n5732) );
  NOR2X0 U7570 ( .IN1(n3742), .IN2(n5733), .QN(WX11612) );
  XOR2X1 U7571 ( .IN1(CRC_OUT_1_1), .IN2(test_so98), .Q(n5733) );
  NOR2X0 U7572 ( .IN1(n3742), .IN2(n5734), .QN(WX11610) );
  XOR2X1 U7573 ( .IN1(n2739), .IN2(DFF_1696_n1), .Q(n5734) );
  NOR2X0 U7574 ( .IN1(n3742), .IN2(n5735), .QN(WX11608) );
  XNOR2X1 U7575 ( .IN1(n2706), .IN2(test_so100), .Q(n5735) );
  NOR2X0 U7576 ( .IN1(n6203), .IN2(n3658), .QN(WX11082) );
  NOR2X0 U7577 ( .IN1(n6204), .IN2(n3658), .QN(WX11080) );
  NOR2X0 U7578 ( .IN1(n6205), .IN2(n3658), .QN(WX11078) );
  NOR2X0 U7579 ( .IN1(n6206), .IN2(n3657), .QN(WX11076) );
  NOR2X0 U7580 ( .IN1(n6207), .IN2(n3657), .QN(WX11074) );
  NOR2X0 U7581 ( .IN1(n6208), .IN2(n3657), .QN(WX11072) );
  NOR2X0 U7582 ( .IN1(n6209), .IN2(n3657), .QN(WX11070) );
  NOR2X0 U7583 ( .IN1(n6210), .IN2(n3657), .QN(WX11068) );
  NOR2X0 U7584 ( .IN1(n6211), .IN2(n3657), .QN(WX11066) );
  AND2X1 U7585 ( .IN1(n3609), .IN2(test_so91), .Q(WX11064) );
  NOR2X0 U7586 ( .IN1(n6213), .IN2(n3657), .QN(WX11062) );
  NOR2X0 U7587 ( .IN1(n6214), .IN2(n3657), .QN(WX11060) );
  NOR2X0 U7588 ( .IN1(n6215), .IN2(n3657), .QN(WX11058) );
  NOR2X0 U7589 ( .IN1(n6216), .IN2(n3657), .QN(WX11056) );
  NOR2X0 U7590 ( .IN1(n6217), .IN2(n3657), .QN(WX11054) );
  NOR2X0 U7591 ( .IN1(n6218), .IN2(n3659), .QN(WX11052) );
  NAND4X0 U7592 ( .IN1(n5736), .IN2(n5737), .IN3(n5738), .IN4(n5739), .QN(
        WX11050) );
  NAND2X0 U7593 ( .IN1(n3010), .IN2(n3949), .QN(n5739) );
  XNOR3X1 U7594 ( .IN1(n2706), .IN2(n2562), .IN3(n5740), .Q(n3949) );
  XOR2X1 U7595 ( .IN1(WX11115), .IN2(n6191), .Q(n5740) );
  NAND2X0 U7596 ( .IN1(WX10888), .IN2(n3042), .QN(n5738) );
  NAND2X0 U7597 ( .IN1(DATA_0_0), .IN2(n3096), .QN(n5737) );
  NAND2X0 U7598 ( .IN1(n3056), .IN2(CRC_OUT_1_0), .QN(n5736) );
  NAND4X0 U7599 ( .IN1(n5741), .IN2(n5742), .IN3(n5743), .IN4(n5744), .QN(
        WX11048) );
  NAND2X0 U7600 ( .IN1(n3010), .IN2(n3955), .QN(n5744) );
  XNOR3X1 U7601 ( .IN1(n2739), .IN2(n2563), .IN3(n5745), .Q(n3955) );
  XOR2X1 U7602 ( .IN1(WX11113), .IN2(n6192), .Q(n5745) );
  NAND2X0 U7603 ( .IN1(WX10886), .IN2(n3042), .QN(n5743) );
  NAND2X0 U7604 ( .IN1(DATA_0_1), .IN2(n3097), .QN(n5742) );
  NAND2X0 U7605 ( .IN1(n3056), .IN2(CRC_OUT_1_1), .QN(n5741) );
  NAND4X0 U7606 ( .IN1(n5746), .IN2(n5747), .IN3(n5748), .IN4(n5749), .QN(
        WX11046) );
  NAND2X0 U7607 ( .IN1(n3961), .IN2(n3018), .QN(n5749) );
  XOR3X1 U7608 ( .IN1(n3535), .IN2(n2564), .IN3(n5750), .Q(n3961) );
  XOR2X1 U7609 ( .IN1(WX11047), .IN2(test_so98), .Q(n5750) );
  NAND2X0 U7610 ( .IN1(WX10884), .IN2(n3042), .QN(n5748) );
  NAND2X0 U7611 ( .IN1(DATA_0_2), .IN2(n3096), .QN(n5747) );
  NAND2X0 U7612 ( .IN1(n3056), .IN2(CRC_OUT_1_2), .QN(n5746) );
  NAND4X0 U7613 ( .IN1(n5751), .IN2(n5752), .IN3(n5753), .IN4(n5754), .QN(
        WX11044) );
  NAND2X0 U7614 ( .IN1(n3010), .IN2(n3967), .QN(n5754) );
  XNOR3X1 U7615 ( .IN1(n2738), .IN2(n2565), .IN3(n5755), .Q(n3967) );
  XOR2X1 U7616 ( .IN1(WX11109), .IN2(n6193), .Q(n5755) );
  NAND2X0 U7617 ( .IN1(WX10882), .IN2(n3042), .QN(n5753) );
  NAND2X0 U7618 ( .IN1(DATA_0_3), .IN2(n3095), .QN(n5752) );
  NAND2X0 U7619 ( .IN1(n3056), .IN2(CRC_OUT_1_3), .QN(n5751) );
  NAND4X0 U7620 ( .IN1(n5756), .IN2(n5757), .IN3(n5758), .IN4(n5759), .QN(
        WX11042) );
  NAND2X0 U7621 ( .IN1(n3973), .IN2(n3018), .QN(n5759) );
  XOR3X1 U7622 ( .IN1(n3539), .IN2(n2687), .IN3(n5760), .Q(n3973) );
  XOR2X1 U7623 ( .IN1(WX11043), .IN2(test_so96), .Q(n5760) );
  NAND2X0 U7624 ( .IN1(WX10880), .IN2(n3042), .QN(n5758) );
  NAND2X0 U7625 ( .IN1(DATA_0_4), .IN2(n3096), .QN(n5757) );
  NAND2X0 U7626 ( .IN1(n3056), .IN2(CRC_OUT_1_4), .QN(n5756) );
  NAND4X0 U7627 ( .IN1(n5761), .IN2(n5762), .IN3(n5763), .IN4(n5764), .QN(
        WX11040) );
  NAND2X0 U7628 ( .IN1(n3010), .IN2(n3979), .QN(n5764) );
  XNOR3X1 U7629 ( .IN1(n2737), .IN2(n2566), .IN3(n5765), .Q(n3979) );
  XOR2X1 U7630 ( .IN1(WX11105), .IN2(n6194), .Q(n5765) );
  NAND2X0 U7631 ( .IN1(WX10878), .IN2(n3042), .QN(n5763) );
  NAND2X0 U7632 ( .IN1(DATA_0_5), .IN2(n3095), .QN(n5762) );
  NAND2X0 U7633 ( .IN1(n3056), .IN2(CRC_OUT_1_5), .QN(n5761) );
  NAND4X0 U7634 ( .IN1(n5766), .IN2(n5767), .IN3(n5768), .IN4(n5769), .QN(
        WX11038) );
  NAND2X0 U7635 ( .IN1(n3985), .IN2(n3019), .QN(n5769) );
  XOR3X1 U7636 ( .IN1(n2736), .IN2(n2567), .IN3(n5770), .Q(n3985) );
  XOR2X1 U7637 ( .IN1(WX11039), .IN2(test_so94), .Q(n5770) );
  NAND2X0 U7638 ( .IN1(WX10876), .IN2(n3043), .QN(n5768) );
  NAND2X0 U7639 ( .IN1(DATA_0_6), .IN2(n3097), .QN(n5767) );
  NAND2X0 U7640 ( .IN1(n3056), .IN2(CRC_OUT_1_6), .QN(n5766) );
  NAND4X0 U7641 ( .IN1(n5771), .IN2(n5772), .IN3(n5773), .IN4(n5774), .QN(
        WX11036) );
  NAND2X0 U7642 ( .IN1(n3009), .IN2(n3991), .QN(n5774) );
  XNOR3X1 U7643 ( .IN1(n2735), .IN2(n2568), .IN3(n5775), .Q(n3991) );
  XOR2X1 U7644 ( .IN1(WX11101), .IN2(n6195), .Q(n5775) );
  NAND2X0 U7645 ( .IN1(WX10874), .IN2(n3043), .QN(n5773) );
  NAND2X0 U7646 ( .IN1(DATA_0_7), .IN2(n3097), .QN(n5772) );
  NAND2X0 U7647 ( .IN1(n3056), .IN2(CRC_OUT_1_7), .QN(n5771) );
  NAND4X0 U7648 ( .IN1(n5776), .IN2(n5777), .IN3(n5778), .IN4(n5779), .QN(
        WX11034) );
  NAND2X0 U7649 ( .IN1(n3997), .IN2(n3019), .QN(n5779) );
  XOR3X1 U7650 ( .IN1(n3547), .IN2(n2734), .IN3(n5780), .Q(n3997) );
  XOR2X1 U7651 ( .IN1(WX11163), .IN2(test_so92), .Q(n5780) );
  NAND2X0 U7652 ( .IN1(WX10872), .IN2(n3043), .QN(n5778) );
  NAND2X0 U7653 ( .IN1(DATA_0_8), .IN2(n3095), .QN(n5777) );
  NAND2X0 U7654 ( .IN1(n3056), .IN2(CRC_OUT_1_8), .QN(n5776) );
  NAND4X0 U7655 ( .IN1(n5781), .IN2(n5782), .IN3(n5783), .IN4(n5784), .QN(
        WX11032) );
  NAND2X0 U7656 ( .IN1(n3009), .IN2(n4003), .QN(n5784) );
  XNOR3X1 U7657 ( .IN1(n2733), .IN2(n2569), .IN3(n5785), .Q(n4003) );
  XOR2X1 U7658 ( .IN1(WX11097), .IN2(n6196), .Q(n5785) );
  NAND2X0 U7659 ( .IN1(WX10870), .IN2(n3043), .QN(n5783) );
  NAND2X0 U7660 ( .IN1(DATA_0_9), .IN2(n3096), .QN(n5782) );
  NAND2X0 U7661 ( .IN1(n3056), .IN2(CRC_OUT_1_9), .QN(n5781) );
  NAND4X0 U7662 ( .IN1(n5786), .IN2(n5787), .IN3(n5788), .IN4(n5789), .QN(
        WX11030) );
  NAND2X0 U7663 ( .IN1(n3009), .IN2(n4009), .QN(n5789) );
  XNOR3X1 U7664 ( .IN1(n2732), .IN2(n2570), .IN3(n5790), .Q(n4009) );
  XOR2X1 U7665 ( .IN1(WX11095), .IN2(n6197), .Q(n5790) );
  NAND2X0 U7666 ( .IN1(WX10868), .IN2(n3043), .QN(n5788) );
  NAND2X0 U7667 ( .IN1(DATA_0_10), .IN2(n3096), .QN(n5787) );
  NAND2X0 U7668 ( .IN1(n3056), .IN2(CRC_OUT_1_10), .QN(n5786) );
  NAND4X0 U7669 ( .IN1(n5791), .IN2(n5792), .IN3(n5793), .IN4(n5794), .QN(
        WX11028) );
  NAND2X0 U7670 ( .IN1(n3009), .IN2(n4015), .QN(n5794) );
  XNOR3X1 U7671 ( .IN1(n2686), .IN2(n2571), .IN3(n5795), .Q(n4015) );
  XOR2X1 U7672 ( .IN1(WX11093), .IN2(n6198), .Q(n5795) );
  NAND2X0 U7673 ( .IN1(WX10866), .IN2(n3043), .QN(n5793) );
  NAND2X0 U7674 ( .IN1(DATA_0_11), .IN2(n3096), .QN(n5792) );
  NAND2X0 U7675 ( .IN1(n3057), .IN2(CRC_OUT_1_11), .QN(n5791) );
  NAND4X0 U7676 ( .IN1(n5796), .IN2(n5797), .IN3(n5798), .IN4(n5799), .QN(
        WX11026) );
  NAND2X0 U7677 ( .IN1(n3009), .IN2(n4021), .QN(n5799) );
  XNOR3X1 U7678 ( .IN1(n2731), .IN2(n2572), .IN3(n5800), .Q(n4021) );
  XOR2X1 U7679 ( .IN1(WX11091), .IN2(n6199), .Q(n5800) );
  NAND2X0 U7680 ( .IN1(WX10864), .IN2(n3043), .QN(n5798) );
  NAND2X0 U7681 ( .IN1(DATA_0_12), .IN2(n3095), .QN(n5797) );
  NAND2X0 U7682 ( .IN1(n3057), .IN2(CRC_OUT_1_12), .QN(n5796) );
  NAND4X0 U7683 ( .IN1(n5801), .IN2(n5802), .IN3(n5803), .IN4(n5804), .QN(
        WX11024) );
  NAND2X0 U7684 ( .IN1(n3009), .IN2(n4027), .QN(n5804) );
  XNOR3X1 U7685 ( .IN1(n2730), .IN2(n2573), .IN3(n5805), .Q(n4027) );
  XOR2X1 U7686 ( .IN1(WX11089), .IN2(n6200), .Q(n5805) );
  NAND2X0 U7687 ( .IN1(WX10862), .IN2(n3043), .QN(n5803) );
  NAND2X0 U7688 ( .IN1(DATA_0_13), .IN2(n3095), .QN(n5802) );
  NAND2X0 U7689 ( .IN1(n3057), .IN2(CRC_OUT_1_13), .QN(n5801) );
  NAND4X0 U7690 ( .IN1(n5806), .IN2(n5807), .IN3(n5808), .IN4(n5809), .QN(
        WX11022) );
  NAND2X0 U7691 ( .IN1(n3009), .IN2(n4033), .QN(n5809) );
  XNOR3X1 U7692 ( .IN1(n2729), .IN2(n2574), .IN3(n5810), .Q(n4033) );
  XOR2X1 U7693 ( .IN1(WX11087), .IN2(n6201), .Q(n5810) );
  NAND2X0 U7694 ( .IN1(WX10860), .IN2(n3043), .QN(n5808) );
  NAND2X0 U7695 ( .IN1(DATA_0_14), .IN2(n3095), .QN(n5807) );
  NAND2X0 U7696 ( .IN1(test_so99), .IN2(n3069), .QN(n5806) );
  NAND4X0 U7697 ( .IN1(n5811), .IN2(n5812), .IN3(n5813), .IN4(n5814), .QN(
        WX11020) );
  NAND2X0 U7698 ( .IN1(n3009), .IN2(n4039), .QN(n5814) );
  XNOR3X1 U7699 ( .IN1(n2728), .IN2(n2575), .IN3(n5815), .Q(n4039) );
  XOR2X1 U7700 ( .IN1(WX11085), .IN2(n6202), .Q(n5815) );
  NAND2X0 U7701 ( .IN1(WX10858), .IN2(n3043), .QN(n5813) );
  NAND2X0 U7702 ( .IN1(DATA_0_15), .IN2(n3095), .QN(n5812) );
  NAND2X0 U7703 ( .IN1(n3057), .IN2(CRC_OUT_1_15), .QN(n5811) );
  NAND4X0 U7704 ( .IN1(n5816), .IN2(n5817), .IN3(n5818), .IN4(n5819), .QN(
        WX11018) );
  NAND2X0 U7705 ( .IN1(n3009), .IN2(n4045), .QN(n5819) );
  XNOR3X1 U7706 ( .IN1(n2350), .IN2(n3575), .IN3(n5820), .Q(n4045) );
  XOR3X1 U7707 ( .IN1(n6203), .IN2(n2685), .IN3(WX11147), .Q(n5820) );
  NAND2X0 U7708 ( .IN1(WX10856), .IN2(n3043), .QN(n5818) );
  NAND2X0 U7709 ( .IN1(DATA_0_16), .IN2(n3095), .QN(n5817) );
  NAND2X0 U7710 ( .IN1(n3057), .IN2(CRC_OUT_1_16), .QN(n5816) );
  NAND4X0 U7711 ( .IN1(n5821), .IN2(n5822), .IN3(n5823), .IN4(n5824), .QN(
        WX11016) );
  NAND2X0 U7712 ( .IN1(n3009), .IN2(n4051), .QN(n5824) );
  XNOR3X1 U7713 ( .IN1(n2352), .IN2(n3576), .IN3(n5825), .Q(n4051) );
  XOR3X1 U7714 ( .IN1(n6204), .IN2(n2727), .IN3(WX11145), .Q(n5825) );
  NAND2X0 U7715 ( .IN1(WX10854), .IN2(n3043), .QN(n5823) );
  NAND2X0 U7716 ( .IN1(DATA_0_17), .IN2(n3095), .QN(n5822) );
  NAND2X0 U7717 ( .IN1(n3057), .IN2(CRC_OUT_1_17), .QN(n5821) );
  NAND4X0 U7718 ( .IN1(n5826), .IN2(n5827), .IN3(n5828), .IN4(n5829), .QN(
        WX11014) );
  NAND2X0 U7719 ( .IN1(n3009), .IN2(n4057), .QN(n5829) );
  XNOR3X1 U7720 ( .IN1(n2354), .IN2(n3575), .IN3(n5830), .Q(n4057) );
  XOR3X1 U7721 ( .IN1(n6205), .IN2(n2726), .IN3(WX11143), .Q(n5830) );
  NAND2X0 U7722 ( .IN1(WX10852), .IN2(n3043), .QN(n5828) );
  NAND2X0 U7723 ( .IN1(DATA_0_18), .IN2(n3095), .QN(n5827) );
  NAND2X0 U7724 ( .IN1(n3057), .IN2(CRC_OUT_1_18), .QN(n5826) );
  NAND4X0 U7725 ( .IN1(n5831), .IN2(n5832), .IN3(n5833), .IN4(n5834), .QN(
        WX11012) );
  NAND2X0 U7726 ( .IN1(n4063), .IN2(n3020), .QN(n5834) );
  XOR3X1 U7727 ( .IN1(n2356), .IN2(n3577), .IN3(n5835), .Q(n4063) );
  XOR3X1 U7728 ( .IN1(test_so97), .IN2(n6206), .IN3(WX11141), .Q(n5835) );
  NAND2X0 U7729 ( .IN1(WX10850), .IN2(n3043), .QN(n5833) );
  NAND2X0 U7730 ( .IN1(DATA_0_19), .IN2(n3096), .QN(n5832) );
  NAND2X0 U7731 ( .IN1(n3057), .IN2(CRC_OUT_1_19), .QN(n5831) );
  NAND4X0 U7732 ( .IN1(n5836), .IN2(n5837), .IN3(n5838), .IN4(n5839), .QN(
        WX11010) );
  NAND2X0 U7733 ( .IN1(n3009), .IN2(n4069), .QN(n5839) );
  XNOR3X1 U7734 ( .IN1(n2357), .IN2(n3575), .IN3(n5840), .Q(n4069) );
  XOR3X1 U7735 ( .IN1(n6207), .IN2(n2725), .IN3(WX11139), .Q(n5840) );
  NAND2X0 U7736 ( .IN1(WX10848), .IN2(n3043), .QN(n5838) );
  NAND2X0 U7737 ( .IN1(DATA_0_20), .IN2(n3095), .QN(n5837) );
  NAND2X0 U7738 ( .IN1(n3057), .IN2(CRC_OUT_1_20), .QN(n5836) );
  NAND4X0 U7739 ( .IN1(n5841), .IN2(n5842), .IN3(n5843), .IN4(n5844), .QN(
        WX11008) );
  NAND2X0 U7740 ( .IN1(n4075), .IN2(n3020), .QN(n5844) );
  XOR3X1 U7741 ( .IN1(n2359), .IN2(n3579), .IN3(n5845), .Q(n4075) );
  XNOR3X1 U7742 ( .IN1(test_so95), .IN2(n6208), .IN3(n2724), .Q(n5845) );
  NAND2X0 U7743 ( .IN1(WX10846), .IN2(n3043), .QN(n5843) );
  NAND2X0 U7744 ( .IN1(DATA_0_21), .IN2(n3094), .QN(n5842) );
  NAND2X0 U7745 ( .IN1(n3057), .IN2(CRC_OUT_1_21), .QN(n5841) );
  NAND4X0 U7746 ( .IN1(n5846), .IN2(n5847), .IN3(n5848), .IN4(n5849), .QN(
        WX11006) );
  NAND2X0 U7747 ( .IN1(n3008), .IN2(n4081), .QN(n5849) );
  XNOR3X1 U7748 ( .IN1(n2360), .IN2(n3576), .IN3(n5850), .Q(n4081) );
  XOR3X1 U7749 ( .IN1(n6209), .IN2(n2723), .IN3(WX11135), .Q(n5850) );
  NAND2X0 U7750 ( .IN1(WX10844), .IN2(n3043), .QN(n5848) );
  NAND2X0 U7751 ( .IN1(DATA_0_22), .IN2(n3095), .QN(n5847) );
  NAND2X0 U7752 ( .IN1(n3057), .IN2(CRC_OUT_1_22), .QN(n5846) );
  NAND4X0 U7753 ( .IN1(n5851), .IN2(n5852), .IN3(n5853), .IN4(n5854), .QN(
        WX11004) );
  NAND2X0 U7754 ( .IN1(n4087), .IN2(n3020), .QN(n5854) );
  XOR3X1 U7755 ( .IN1(n2362), .IN2(n3578), .IN3(n5855), .Q(n4087) );
  XNOR3X1 U7756 ( .IN1(test_so93), .IN2(n6210), .IN3(n2722), .Q(n5855) );
  NAND2X0 U7757 ( .IN1(WX10842), .IN2(n3044), .QN(n5853) );
  NAND2X0 U7758 ( .IN1(DATA_0_23), .IN2(n3094), .QN(n5852) );
  NAND2X0 U7759 ( .IN1(n3057), .IN2(CRC_OUT_1_23), .QN(n5851) );
  NAND4X0 U7760 ( .IN1(n5856), .IN2(n5857), .IN3(n5858), .IN4(n5859), .QN(
        WX11002) );
  NAND2X0 U7761 ( .IN1(n3008), .IN2(n4093), .QN(n5859) );
  XNOR3X1 U7762 ( .IN1(n2363), .IN2(n3574), .IN3(n5860), .Q(n4093) );
  XOR3X1 U7763 ( .IN1(n6211), .IN2(n2721), .IN3(WX11131), .Q(n5860) );
  NAND2X0 U7764 ( .IN1(WX10840), .IN2(n3044), .QN(n5858) );
  NAND2X0 U7765 ( .IN1(DATA_0_24), .IN2(n3094), .QN(n5857) );
  NAND2X0 U7766 ( .IN1(n3058), .IN2(CRC_OUT_1_24), .QN(n5856) );
  NAND4X0 U7767 ( .IN1(n5861), .IN2(n5862), .IN3(n5863), .IN4(n5864), .QN(
        WX11000) );
  NAND2X0 U7768 ( .IN1(n4099), .IN2(n3020), .QN(n5864) );
  XOR3X1 U7769 ( .IN1(n2365), .IN2(n3578), .IN3(n5865), .Q(n4099) );
  XNOR3X1 U7770 ( .IN1(test_so91), .IN2(n6212), .IN3(n2720), .Q(n5865) );
  NAND2X0 U7771 ( .IN1(WX10838), .IN2(n3044), .QN(n5863) );
  NAND2X0 U7772 ( .IN1(DATA_0_25), .IN2(n3095), .QN(n5862) );
  NAND2X0 U7773 ( .IN1(n3058), .IN2(CRC_OUT_1_25), .QN(n5861) );
  NAND4X0 U7774 ( .IN1(n5866), .IN2(n5867), .IN3(n5868), .IN4(n5869), .QN(
        WX10998) );
  NAND2X0 U7775 ( .IN1(n3008), .IN2(n4105), .QN(n5869) );
  XNOR3X1 U7776 ( .IN1(n2366), .IN2(n3575), .IN3(n5870), .Q(n4105) );
  XOR3X1 U7777 ( .IN1(n6213), .IN2(n2719), .IN3(WX11127), .Q(n5870) );
  NAND2X0 U7778 ( .IN1(WX10836), .IN2(n3044), .QN(n5868) );
  NAND2X0 U7779 ( .IN1(DATA_0_26), .IN2(n3094), .QN(n5867) );
  NAND2X0 U7780 ( .IN1(n3058), .IN2(CRC_OUT_1_26), .QN(n5866) );
  NAND4X0 U7781 ( .IN1(n5871), .IN2(n5872), .IN3(n5873), .IN4(n5874), .QN(
        WX10996) );
  NAND2X0 U7782 ( .IN1(n3008), .IN2(n4111), .QN(n5874) );
  XNOR3X1 U7783 ( .IN1(n2368), .IN2(n3576), .IN3(n5875), .Q(n4111) );
  XOR3X1 U7784 ( .IN1(n6214), .IN2(n2718), .IN3(WX11125), .Q(n5875) );
  NAND2X0 U7785 ( .IN1(WX10834), .IN2(n3044), .QN(n5873) );
  NAND2X0 U7786 ( .IN1(DATA_0_27), .IN2(n3096), .QN(n5872) );
  NAND2X0 U7787 ( .IN1(n3058), .IN2(CRC_OUT_1_27), .QN(n5871) );
  NAND4X0 U7788 ( .IN1(n5876), .IN2(n5877), .IN3(n5878), .IN4(n5879), .QN(
        WX10994) );
  NAND2X0 U7789 ( .IN1(n3008), .IN2(n4117), .QN(n5879) );
  XNOR3X1 U7790 ( .IN1(n2370), .IN2(n3576), .IN3(n5880), .Q(n4117) );
  XOR3X1 U7791 ( .IN1(n6215), .IN2(n2717), .IN3(WX11123), .Q(n5880) );
  NAND2X0 U7792 ( .IN1(WX10832), .IN2(n3044), .QN(n5878) );
  NAND2X0 U7793 ( .IN1(DATA_0_28), .IN2(n3094), .QN(n5877) );
  NAND2X0 U7794 ( .IN1(n3058), .IN2(CRC_OUT_1_28), .QN(n5876) );
  NAND4X0 U7795 ( .IN1(n5881), .IN2(n5882), .IN3(n5883), .IN4(n5884), .QN(
        WX10992) );
  NAND2X0 U7796 ( .IN1(n3008), .IN2(n4123), .QN(n5884) );
  XNOR3X1 U7797 ( .IN1(n2372), .IN2(n3575), .IN3(n5885), .Q(n4123) );
  XOR3X1 U7798 ( .IN1(n6216), .IN2(n2716), .IN3(WX11121), .Q(n5885) );
  NAND2X0 U7799 ( .IN1(WX10830), .IN2(n3044), .QN(n5883) );
  NAND2X0 U7800 ( .IN1(DATA_0_29), .IN2(n3094), .QN(n5882) );
  NAND2X0 U7801 ( .IN1(n3058), .IN2(CRC_OUT_1_29), .QN(n5881) );
  NAND4X0 U7802 ( .IN1(n5886), .IN2(n5887), .IN3(n5888), .IN4(n5889), .QN(
        WX10990) );
  NAND2X0 U7803 ( .IN1(n3013), .IN2(n4129), .QN(n5889) );
  XNOR3X1 U7804 ( .IN1(n2374), .IN2(n3576), .IN3(n5890), .Q(n4129) );
  XOR3X1 U7805 ( .IN1(n6217), .IN2(n2715), .IN3(WX11119), .Q(n5890) );
  NAND2X0 U7806 ( .IN1(WX10828), .IN2(n3044), .QN(n5888) );
  AND2X1 U7807 ( .IN1(n3579), .IN2(TM0), .Q(n2148) );
  NAND2X0 U7808 ( .IN1(DATA_0_30), .IN2(n3095), .QN(n5887) );
  NAND2X0 U7809 ( .IN1(n3058), .IN2(CRC_OUT_1_30), .QN(n5886) );
  NAND4X0 U7810 ( .IN1(n5891), .IN2(n5892), .IN3(n5893), .IN4(n5894), .QN(
        WX10988) );
  NAND2X0 U7811 ( .IN1(n2998), .IN2(n4135), .QN(n5894) );
  XNOR3X1 U7812 ( .IN1(n2335), .IN2(n3575), .IN3(n5895), .Q(n4135) );
  XOR3X1 U7813 ( .IN1(n6218), .IN2(n2714), .IN3(WX11117), .Q(n5895) );
  AND3X1 U7814 ( .IN1(n3597), .IN2(n281), .IN3(n3579), .Q(n3947) );
  NAND2X0 U7815 ( .IN1(DATA_0_31), .IN2(n3098), .QN(n5893) );
  NAND2X0 U7816 ( .IN1(test_so100), .IN2(n3070), .QN(n5892) );
  NAND2X0 U7817 ( .IN1(n2245), .IN2(WX10829), .QN(n5891) );
  NOR2X0 U7818 ( .IN1(n3742), .IN2(WX10829), .QN(WX10890) );
  AND2X1 U7819 ( .IN1(n3609), .IN2(n8263), .Q(WX10888) );
  AND2X1 U7820 ( .IN1(n3609), .IN2(n8264), .Q(WX10886) );
  AND2X1 U7821 ( .IN1(n3609), .IN2(n8265), .Q(WX10884) );
  AND2X1 U7822 ( .IN1(n3609), .IN2(n8266), .Q(WX10882) );
  AND2X1 U7823 ( .IN1(n3609), .IN2(n8267), .Q(WX10880) );
  AND2X1 U7824 ( .IN1(n3610), .IN2(n8268), .Q(WX10878) );
  AND2X1 U7825 ( .IN1(n3610), .IN2(n8269), .Q(WX10876) );
  AND2X1 U7826 ( .IN1(n3610), .IN2(n8270), .Q(WX10874) );
  AND2X1 U7827 ( .IN1(n3610), .IN2(n8271), .Q(WX10872) );
  AND2X1 U7828 ( .IN1(n3610), .IN2(n8272), .Q(WX10870) );
  AND2X1 U7829 ( .IN1(test_so90), .IN2(n3599), .Q(WX10868) );
  AND2X1 U7830 ( .IN1(n3610), .IN2(n8275), .Q(WX10866) );
  AND2X1 U7831 ( .IN1(n3610), .IN2(n8276), .Q(WX10864) );
  AND2X1 U7832 ( .IN1(n3610), .IN2(n8277), .Q(WX10862) );
  AND2X1 U7833 ( .IN1(n3610), .IN2(n8278), .Q(WX10860) );
  AND2X1 U7834 ( .IN1(n3611), .IN2(n8279), .Q(WX10858) );
  AND2X1 U7835 ( .IN1(n3611), .IN2(n8280), .Q(WX10856) );
  AND2X1 U7836 ( .IN1(n3611), .IN2(n8281), .Q(WX10854) );
  AND2X1 U7837 ( .IN1(n3611), .IN2(n8282), .Q(WX10852) );
  AND2X1 U7838 ( .IN1(n3611), .IN2(n8283), .Q(WX10850) );
  AND2X1 U7839 ( .IN1(n3611), .IN2(n8284), .Q(WX10848) );
  AND2X1 U7840 ( .IN1(n3611), .IN2(n8285), .Q(WX10846) );
  AND2X1 U7841 ( .IN1(n3611), .IN2(n8286), .Q(WX10844) );
  AND2X1 U7842 ( .IN1(n3611), .IN2(n8287), .Q(WX10842) );
  AND2X1 U7843 ( .IN1(n3612), .IN2(n8288), .Q(WX10840) );
  AND2X1 U7844 ( .IN1(n3612), .IN2(n8289), .Q(WX10838) );
  AND2X1 U7845 ( .IN1(n3612), .IN2(n8290), .Q(WX10836) );
  AND2X1 U7846 ( .IN1(test_so89), .IN2(n3598), .Q(WX10834) );
  AND2X1 U7847 ( .IN1(n3612), .IN2(n8293), .Q(WX10832) );
  AND2X1 U7848 ( .IN1(n3612), .IN2(n8294), .Q(WX10830) );
  AND2X1 U7849 ( .IN1(n3612), .IN2(n8295), .Q(WX10828) );
  NOR2X0 U7850 ( .IN1(n3742), .IN2(n5896), .QN(WX10377) );
  XOR2X1 U7851 ( .IN1(CRC_OUT_2_30), .IN2(test_so85), .Q(n5896) );
  NOR2X0 U7852 ( .IN1(n3742), .IN2(n5897), .QN(WX10375) );
  XOR2X1 U7853 ( .IN1(n2740), .IN2(DFF_1533_n1), .Q(n5897) );
  NOR2X0 U7854 ( .IN1(n3742), .IN2(n5898), .QN(WX10373) );
  XOR2X1 U7855 ( .IN1(n2741), .IN2(DFF_1532_n1), .Q(n5898) );
  NOR2X0 U7856 ( .IN1(n3742), .IN2(n5899), .QN(WX10371) );
  XOR2X1 U7857 ( .IN1(n2742), .IN2(DFF_1531_n1), .Q(n5899) );
  NOR2X0 U7858 ( .IN1(n3743), .IN2(n5900), .QN(WX10369) );
  XOR2X1 U7859 ( .IN1(n2743), .IN2(DFF_1530_n1), .Q(n5900) );
  NOR2X0 U7860 ( .IN1(n3743), .IN2(n5901), .QN(WX10367) );
  XOR2X1 U7861 ( .IN1(n2744), .IN2(DFF_1529_n1), .Q(n5901) );
  NOR2X0 U7862 ( .IN1(n3743), .IN2(n5902), .QN(WX10365) );
  XOR2X1 U7863 ( .IN1(n2745), .IN2(DFF_1528_n1), .Q(n5902) );
  NOR2X0 U7864 ( .IN1(n3743), .IN2(n5903), .QN(WX10363) );
  XOR2X1 U7865 ( .IN1(n2746), .IN2(DFF_1527_n1), .Q(n5903) );
  NOR2X0 U7866 ( .IN1(n3743), .IN2(n5904), .QN(WX10361) );
  XOR2X1 U7867 ( .IN1(n2747), .IN2(DFF_1526_n1), .Q(n5904) );
  NOR2X0 U7868 ( .IN1(n3743), .IN2(n5905), .QN(WX10359) );
  XOR2X1 U7869 ( .IN1(n2748), .IN2(DFF_1525_n1), .Q(n5905) );
  NOR2X0 U7870 ( .IN1(n3743), .IN2(n5906), .QN(WX10357) );
  XOR2X1 U7871 ( .IN1(n2749), .IN2(DFF_1524_n1), .Q(n5906) );
  NOR2X0 U7872 ( .IN1(n3743), .IN2(n5907), .QN(WX10355) );
  XNOR2X1 U7873 ( .IN1(n2750), .IN2(test_so88), .Q(n5907) );
  NOR2X0 U7874 ( .IN1(n3743), .IN2(n5908), .QN(WX10353) );
  XOR2X1 U7875 ( .IN1(n2751), .IN2(DFF_1522_n1), .Q(n5908) );
  NOR2X0 U7876 ( .IN1(n3743), .IN2(n5909), .QN(WX10351) );
  XOR2X1 U7877 ( .IN1(n2752), .IN2(DFF_1521_n1), .Q(n5909) );
  NOR2X0 U7878 ( .IN1(n3743), .IN2(n5910), .QN(WX10349) );
  XOR2X1 U7879 ( .IN1(n2753), .IN2(DFF_1520_n1), .Q(n5910) );
  NOR2X0 U7880 ( .IN1(n3743), .IN2(n5911), .QN(WX10347) );
  XOR3X1 U7881 ( .IN1(n2688), .IN2(DFF_1535_n1), .IN3(CRC_OUT_2_15), .Q(n5911)
         );
  NOR2X0 U7882 ( .IN1(n3743), .IN2(n5912), .QN(WX10345) );
  XOR2X1 U7883 ( .IN1(n2754), .IN2(DFF_1518_n1), .Q(n5912) );
  NOR2X0 U7884 ( .IN1(n3744), .IN2(n5913), .QN(WX10343) );
  XOR2X1 U7885 ( .IN1(CRC_OUT_2_13), .IN2(test_so86), .Q(n5913) );
  NOR2X0 U7886 ( .IN1(n3744), .IN2(n5914), .QN(WX10341) );
  XOR2X1 U7887 ( .IN1(n2755), .IN2(DFF_1516_n1), .Q(n5914) );
  NOR2X0 U7888 ( .IN1(n3744), .IN2(n5915), .QN(WX10339) );
  XOR2X1 U7889 ( .IN1(n2756), .IN2(DFF_1515_n1), .Q(n5915) );
  NOR2X0 U7890 ( .IN1(n3744), .IN2(n5916), .QN(WX10337) );
  XOR3X1 U7891 ( .IN1(n2689), .IN2(DFF_1535_n1), .IN3(CRC_OUT_2_10), .Q(n5916)
         );
  NOR2X0 U7892 ( .IN1(n3744), .IN2(n5917), .QN(WX10335) );
  XOR2X1 U7893 ( .IN1(n2757), .IN2(DFF_1513_n1), .Q(n5917) );
  NOR2X0 U7894 ( .IN1(n3744), .IN2(n5918), .QN(WX10333) );
  XOR2X1 U7895 ( .IN1(n2758), .IN2(DFF_1512_n1), .Q(n5918) );
  NOR2X0 U7896 ( .IN1(n3744), .IN2(n5919), .QN(WX10331) );
  XOR2X1 U7897 ( .IN1(n2759), .IN2(DFF_1511_n1), .Q(n5919) );
  NOR2X0 U7898 ( .IN1(n3744), .IN2(n5920), .QN(WX10329) );
  XOR2X1 U7899 ( .IN1(n2760), .IN2(DFF_1510_n1), .Q(n5920) );
  NOR2X0 U7900 ( .IN1(n3744), .IN2(n5921), .QN(WX10327) );
  XOR2X1 U7901 ( .IN1(n2761), .IN2(DFF_1509_n1), .Q(n5921) );
  NOR2X0 U7902 ( .IN1(n3744), .IN2(n5922), .QN(WX10325) );
  XOR2X1 U7903 ( .IN1(n2762), .IN2(DFF_1508_n1), .Q(n5922) );
  NOR2X0 U7904 ( .IN1(n3744), .IN2(n5923), .QN(WX10323) );
  XOR3X1 U7905 ( .IN1(n2690), .IN2(DFF_1535_n1), .IN3(CRC_OUT_2_3), .Q(n5923)
         );
  NOR2X0 U7906 ( .IN1(n3744), .IN2(n5924), .QN(WX10321) );
  XNOR2X1 U7907 ( .IN1(n2763), .IN2(test_so87), .Q(n5924) );
  NOR2X0 U7908 ( .IN1(n3744), .IN2(n5925), .QN(WX10319) );
  XOR2X1 U7909 ( .IN1(n2764), .IN2(DFF_1505_n1), .Q(n5925) );
  NOR2X0 U7910 ( .IN1(n3745), .IN2(n5926), .QN(WX10317) );
  XOR2X1 U7911 ( .IN1(n2765), .IN2(DFF_1504_n1), .Q(n5926) );
  NOR2X0 U7912 ( .IN1(n3745), .IN2(n5927), .QN(WX10315) );
  XOR2X1 U7913 ( .IN1(n2707), .IN2(DFF_1535_n1), .Q(n5927) );
  XNOR2X1 U7914 ( .IN1(n5928), .IN2(n4643), .Q(DATA_9_9) );
  XNOR3X1 U7915 ( .IN1(n2953), .IN2(TM0), .IN3(n5929), .Q(n4643) );
  XNOR3X1 U7916 ( .IN1(n6219), .IN2(n3485), .IN3(n2954), .Q(n5929) );
  NAND2X0 U7917 ( .IN1(TM0), .IN2(WX529), .QN(n5928) );
  XNOR2X1 U7918 ( .IN1(n5930), .IN2(n4637), .Q(DATA_9_8) );
  XNOR3X1 U7919 ( .IN1(n2959), .IN2(TM0), .IN3(n5931), .Q(n4637) );
  XOR3X1 U7920 ( .IN1(n6220), .IN2(n3483), .IN3(WX755), .Q(n5931) );
  NAND2X0 U7921 ( .IN1(TM0), .IN2(WX531), .QN(n5930) );
  XNOR2X1 U7922 ( .IN1(n5932), .IN2(n4631), .Q(DATA_9_7) );
  XNOR3X1 U7923 ( .IN1(n2983), .IN2(TM0), .IN3(n5933), .Q(n4631) );
  XOR3X1 U7924 ( .IN1(n3481), .IN2(n2985), .IN3(WX821), .Q(n5933) );
  NAND2X0 U7925 ( .IN1(TM0), .IN2(WX533), .QN(n5932) );
  XNOR2X1 U7926 ( .IN1(n5934), .IN2(n4625), .Q(DATA_9_6) );
  XNOR3X1 U7927 ( .IN1(n2974), .IN2(n281), .IN3(n5935), .Q(n4625) );
  XNOR3X1 U7928 ( .IN1(test_so5), .IN2(n3479), .IN3(n2975), .Q(n5935) );
  NAND2X0 U7929 ( .IN1(TM0), .IN2(WX535), .QN(n5934) );
  XNOR2X1 U7930 ( .IN1(n5936), .IN2(n4619), .Q(DATA_9_5) );
  XNOR3X1 U7931 ( .IN1(n2961), .IN2(TM0), .IN3(n5937), .Q(n4619) );
  XOR3X1 U7932 ( .IN1(n6221), .IN2(n3477), .IN3(WX761), .Q(n5937) );
  NAND2X0 U7933 ( .IN1(TM0), .IN2(WX537), .QN(n5936) );
  XNOR2X1 U7934 ( .IN1(n5938), .IN2(n4613), .Q(DATA_9_4) );
  XNOR3X1 U7935 ( .IN1(n2963), .IN2(TM0), .IN3(n5939), .Q(n4613) );
  XOR3X1 U7936 ( .IN1(n6222), .IN2(n3475), .IN3(WX763), .Q(n5939) );
  NAND2X0 U7937 ( .IN1(TM0), .IN2(WX539), .QN(n5938) );
  XNOR2X1 U7938 ( .IN1(n5940), .IN2(n4805), .Q(DATA_9_31) );
  XNOR3X1 U7939 ( .IN1(n2977), .IN2(n3576), .IN3(n5941), .Q(n4805) );
  XNOR3X1 U7940 ( .IN1(n6223), .IN2(n3529), .IN3(n2978), .Q(n5941) );
  NAND2X0 U7941 ( .IN1(TM0), .IN2(WX485), .QN(n5940) );
  XNOR2X1 U7942 ( .IN1(n5942), .IN2(n4789), .Q(DATA_9_30) );
  XNOR3X1 U7943 ( .IN1(n2926), .IN2(n3575), .IN3(n5943), .Q(n4789) );
  XOR3X1 U7944 ( .IN1(n3527), .IN2(n2928), .IN3(WX775), .Q(n5943) );
  NAND2X0 U7945 ( .IN1(TM0), .IN2(WX487), .QN(n5942) );
  XNOR2X1 U7946 ( .IN1(n5944), .IN2(n4607), .Q(DATA_9_3) );
  XNOR3X1 U7947 ( .IN1(n2929), .IN2(TM0), .IN3(n5945), .Q(n4607) );
  XOR3X1 U7948 ( .IN1(n6224), .IN2(n3473), .IN3(WX765), .Q(n5945) );
  NAND2X0 U7949 ( .IN1(TM0), .IN2(WX541), .QN(n5944) );
  XNOR2X1 U7950 ( .IN1(n5946), .IN2(n4773), .Q(DATA_9_29) );
  XNOR3X1 U7951 ( .IN1(n2933), .IN2(n3576), .IN3(n5947), .Q(n4773) );
  XOR3X1 U7952 ( .IN1(n6225), .IN2(n3525), .IN3(WX713), .Q(n5947) );
  NAND2X0 U7953 ( .IN1(TM0), .IN2(WX489), .QN(n5946) );
  XNOR2X1 U7954 ( .IN1(n5948), .IN2(n4757), .Q(DATA_9_28) );
  XOR3X1 U7955 ( .IN1(n2939), .IN2(n3579), .IN3(n5949), .Q(n4757) );
  XOR3X1 U7956 ( .IN1(test_so2), .IN2(n6226), .IN3(WX779), .Q(n5949) );
  NAND2X0 U7957 ( .IN1(TM0), .IN2(WX491), .QN(n5948) );
  XNOR2X1 U7958 ( .IN1(n5950), .IN2(n4751), .Q(DATA_9_27) );
  XNOR3X1 U7959 ( .IN1(n2942), .IN2(n3575), .IN3(n5951), .Q(n4751) );
  XOR3X1 U7960 ( .IN1(n6227), .IN2(n3521), .IN3(WX717), .Q(n5951) );
  NAND2X0 U7961 ( .IN1(TM0), .IN2(WX493), .QN(n5950) );
  XNOR2X1 U7962 ( .IN1(n5952), .IN2(n4745), .Q(DATA_9_26) );
  XNOR3X1 U7963 ( .IN1(n2944), .IN2(n3576), .IN3(n5953), .Q(n4745) );
  XOR3X1 U7964 ( .IN1(n6228), .IN2(n3519), .IN3(WX719), .Q(n5953) );
  NAND2X0 U7965 ( .IN1(TM0), .IN2(WX495), .QN(n5952) );
  XNOR2X1 U7966 ( .IN1(n5954), .IN2(n4739), .Q(DATA_9_25) );
  XNOR3X1 U7967 ( .IN1(n2949), .IN2(n3576), .IN3(n5955), .Q(n4739) );
  XOR3X1 U7968 ( .IN1(n6229), .IN2(n3517), .IN3(WX721), .Q(n5955) );
  NAND2X0 U7969 ( .IN1(TM0), .IN2(WX497), .QN(n5954) );
  XNOR2X1 U7970 ( .IN1(n5956), .IN2(n4733), .Q(DATA_9_24) );
  XOR3X1 U7971 ( .IN1(n2955), .IN2(n3579), .IN3(n5957), .Q(n4733) );
  XOR3X1 U7972 ( .IN1(test_so4), .IN2(n6230), .IN3(WX659), .Q(n5957) );
  NAND2X0 U7973 ( .IN1(TM0), .IN2(WX499), .QN(n5956) );
  XNOR2X1 U7974 ( .IN1(n5958), .IN2(n4727), .Q(DATA_9_23) );
  XNOR3X1 U7975 ( .IN1(n2956), .IN2(n3576), .IN3(n5959), .Q(n4727) );
  XOR3X1 U7976 ( .IN1(n6231), .IN2(n3513), .IN3(WX725), .Q(n5959) );
  NAND2X0 U7977 ( .IN1(TM0), .IN2(WX501), .QN(n5958) );
  XNOR2X1 U7978 ( .IN1(n5960), .IN2(n4721), .Q(DATA_9_22) );
  XNOR3X1 U7979 ( .IN1(n2965), .IN2(n3576), .IN3(n5961), .Q(n4721) );
  XOR3X1 U7980 ( .IN1(n3511), .IN2(n2967), .IN3(WX791), .Q(n5961) );
  NAND2X0 U7981 ( .IN1(TM0), .IN2(WX503), .QN(n5960) );
  XNOR2X1 U7982 ( .IN1(n5962), .IN2(n4715), .Q(DATA_9_21) );
  XNOR3X1 U7983 ( .IN1(n2971), .IN2(n3577), .IN3(n5963), .Q(n4715) );
  XOR3X1 U7984 ( .IN1(n3509), .IN2(n2973), .IN3(WX793), .Q(n5963) );
  NAND2X0 U7985 ( .IN1(TM0), .IN2(WX505), .QN(n5962) );
  XNOR2X1 U7986 ( .IN1(n5964), .IN2(n4709), .Q(DATA_9_20) );
  XOR3X1 U7987 ( .IN1(n2976), .IN2(n3579), .IN3(n5965), .Q(n4709) );
  XOR3X1 U7988 ( .IN1(test_so6), .IN2(n6232), .IN3(WX667), .Q(n5965) );
  NAND2X0 U7989 ( .IN1(TM0), .IN2(WX507), .QN(n5964) );
  XNOR2X1 U7990 ( .IN1(n5966), .IN2(n4601), .Q(DATA_9_2) );
  XNOR3X1 U7991 ( .IN1(n2981), .IN2(n281), .IN3(n5967), .Q(n4601) );
  XNOR3X1 U7992 ( .IN1(test_so7), .IN2(n3471), .IN3(n2982), .Q(n5967) );
  NAND2X0 U7993 ( .IN1(TM0), .IN2(WX543), .QN(n5966) );
  XNOR2X1 U7994 ( .IN1(n5968), .IN2(n4703), .Q(DATA_9_19) );
  XNOR3X1 U7995 ( .IN1(n2931), .IN2(n3576), .IN3(n5969), .Q(n4703) );
  XOR3X1 U7996 ( .IN1(n6233), .IN2(n3505), .IN3(WX733), .Q(n5969) );
  NAND2X0 U7997 ( .IN1(TM0), .IN2(WX509), .QN(n5968) );
  XNOR2X1 U7998 ( .IN1(n5970), .IN2(n4697), .Q(DATA_9_18) );
  XNOR3X1 U7999 ( .IN1(n2940), .IN2(n3577), .IN3(n5971), .Q(n4697) );
  XOR3X1 U8000 ( .IN1(n6234), .IN2(n3503), .IN3(WX735), .Q(n5971) );
  NAND2X0 U8001 ( .IN1(TM0), .IN2(WX511), .QN(n5970) );
  XNOR2X1 U8002 ( .IN1(n5972), .IN2(n4691), .Q(DATA_9_17) );
  XNOR3X1 U8003 ( .IN1(n2947), .IN2(n3577), .IN3(n5973), .Q(n4691) );
  XOR3X1 U8004 ( .IN1(n6235), .IN2(n3501), .IN3(WX737), .Q(n5973) );
  NAND2X0 U8005 ( .IN1(TM0), .IN2(WX513), .QN(n5972) );
  XNOR2X1 U8006 ( .IN1(n5974), .IN2(n4685), .Q(DATA_9_16) );
  XOR3X1 U8007 ( .IN1(n2958), .IN2(n3579), .IN3(n5975), .Q(n4685) );
  XOR3X1 U8008 ( .IN1(test_so8), .IN2(n6236), .IN3(WX675), .Q(n5975) );
  NAND2X0 U8009 ( .IN1(TM0), .IN2(WX515), .QN(n5974) );
  XNOR2X1 U8010 ( .IN1(n5976), .IN2(n4679), .Q(DATA_9_15) );
  XNOR3X1 U8011 ( .IN1(n2968), .IN2(TM0), .IN3(n5977), .Q(n4679) );
  XOR3X1 U8012 ( .IN1(n3497), .IN2(n2970), .IN3(WX805), .Q(n5977) );
  NAND2X0 U8013 ( .IN1(TM0), .IN2(WX517), .QN(n5976) );
  XNOR2X1 U8014 ( .IN1(n5978), .IN2(n4673), .Q(DATA_9_14) );
  XNOR3X1 U8015 ( .IN1(n2979), .IN2(TM0), .IN3(n5979), .Q(n4673) );
  XOR3X1 U8016 ( .IN1(n6237), .IN2(n3495), .IN3(WX743), .Q(n5979) );
  NAND2X0 U8017 ( .IN1(test_so1), .IN2(TM0), .QN(n5978) );
  XNOR2X1 U8018 ( .IN1(n5980), .IN2(n4667), .Q(DATA_9_13) );
  XNOR3X1 U8019 ( .IN1(n2935), .IN2(TM0), .IN3(n5981), .Q(n4667) );
  XOR3X1 U8020 ( .IN1(n6238), .IN2(n3493), .IN3(WX745), .Q(n5981) );
  NAND2X0 U8021 ( .IN1(TM0), .IN2(WX521), .QN(n5980) );
  XNOR2X1 U8022 ( .IN1(n5982), .IN2(n4661), .Q(DATA_9_12) );
  XNOR3X1 U8023 ( .IN1(n2951), .IN2(TM0), .IN3(n5983), .Q(n4661) );
  XOR3X1 U8024 ( .IN1(n6239), .IN2(n3491), .IN3(WX747), .Q(n5983) );
  NAND2X0 U8025 ( .IN1(TM0), .IN2(WX523), .QN(n5982) );
  XNOR2X1 U8026 ( .IN1(n5984), .IN2(n4655), .Q(DATA_9_11) );
  XNOR3X1 U8027 ( .IN1(n2986), .IN2(TM0), .IN3(n5985), .Q(n4655) );
  XOR3X1 U8028 ( .IN1(n6240), .IN2(n3489), .IN3(WX749), .Q(n5985) );
  NAND2X0 U8029 ( .IN1(TM0), .IN2(WX525), .QN(n5984) );
  XNOR2X1 U8030 ( .IN1(n5986), .IN2(n4649), .Q(DATA_9_10) );
  XNOR3X1 U8031 ( .IN1(n2946), .IN2(n281), .IN3(n5987), .Q(n4649) );
  XOR3X1 U8032 ( .IN1(test_so3), .IN2(n6241), .IN3(WX815), .Q(n5987) );
  INVX0 U8033 ( .INP(TM0), .ZN(n281) );
  NAND2X0 U8034 ( .IN1(TM0), .IN2(WX527), .QN(n5986) );
  XNOR2X1 U8035 ( .IN1(n5988), .IN2(n4595), .Q(DATA_9_1) );
  XNOR3X1 U8036 ( .IN1(n2937), .IN2(TM0), .IN3(n5989), .Q(n4595) );
  XOR3X1 U8037 ( .IN1(n6242), .IN2(n3469), .IN3(WX769), .Q(n5989) );
  NAND2X0 U8038 ( .IN1(TM0), .IN2(WX545), .QN(n5988) );
  XNOR2X1 U8039 ( .IN1(n5990), .IN2(n4589), .Q(DATA_9_0) );
  XNOR3X1 U8040 ( .IN1(n2988), .IN2(TM0), .IN3(n5991), .Q(n4589) );
  XOR3X1 U8041 ( .IN1(n3467), .IN2(n2990), .IN3(WX835), .Q(n5991) );
  NAND2X0 U8042 ( .IN1(TM0), .IN2(WX547), .QN(n5990) );
  NOR2X0 U3558_U2 ( .IN1(n3704), .IN2(U3558_n1), .QN(n2245) );
  INVX0 U3558_U1 ( .INP(n3028), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(n3278), .ZN(U3871_n1) );
  NOR2X0 U3871_U1 ( .IN1(TM0), .IN2(U3871_n1), .QN(n2153) );
  INVX0 U3991_U2 ( .INP(n3278), .ZN(U3991_n1) );
  NOR2X0 U3991_U1 ( .IN1(n281), .IN2(U3991_n1), .QN(n2152) );
  INVX0 U5716_U2 ( .INP(WX547), .ZN(U5716_n1) );
  NOR2X0 U5716_U1 ( .IN1(n3689), .IN2(U5716_n1), .QN(WX544) );
  INVX0 U5717_U2 ( .INP(WX545), .ZN(U5717_n1) );
  NOR2X0 U5717_U1 ( .IN1(n3708), .IN2(U5717_n1), .QN(WX542) );
  INVX0 U5718_U2 ( .INP(WX543), .ZN(U5718_n1) );
  NOR2X0 U5718_U1 ( .IN1(n3708), .IN2(U5718_n1), .QN(WX540) );
  INVX0 U5719_U2 ( .INP(WX541), .ZN(U5719_n1) );
  NOR2X0 U5719_U1 ( .IN1(n3708), .IN2(U5719_n1), .QN(WX538) );
  INVX0 U5720_U2 ( .INP(WX539), .ZN(U5720_n1) );
  NOR2X0 U5720_U1 ( .IN1(n3708), .IN2(U5720_n1), .QN(WX536) );
  INVX0 U5721_U2 ( .INP(WX537), .ZN(U5721_n1) );
  NOR2X0 U5721_U1 ( .IN1(n3708), .IN2(U5721_n1), .QN(WX534) );
  INVX0 U5722_U2 ( .INP(WX535), .ZN(U5722_n1) );
  NOR2X0 U5722_U1 ( .IN1(n3708), .IN2(U5722_n1), .QN(WX532) );
  INVX0 U5723_U2 ( .INP(WX533), .ZN(U5723_n1) );
  NOR2X0 U5723_U1 ( .IN1(n3708), .IN2(U5723_n1), .QN(WX530) );
  INVX0 U5724_U2 ( .INP(WX531), .ZN(U5724_n1) );
  NOR2X0 U5724_U1 ( .IN1(n3708), .IN2(U5724_n1), .QN(WX528) );
  INVX0 U5725_U2 ( .INP(WX529), .ZN(U5725_n1) );
  NOR2X0 U5725_U1 ( .IN1(n3708), .IN2(U5725_n1), .QN(WX526) );
  INVX0 U5726_U2 ( .INP(WX527), .ZN(U5726_n1) );
  NOR2X0 U5726_U1 ( .IN1(n3707), .IN2(U5726_n1), .QN(WX524) );
  INVX0 U5727_U2 ( .INP(WX525), .ZN(U5727_n1) );
  NOR2X0 U5727_U1 ( .IN1(n3707), .IN2(U5727_n1), .QN(WX522) );
  INVX0 U5728_U2 ( .INP(WX523), .ZN(U5728_n1) );
  NOR2X0 U5728_U1 ( .IN1(n3707), .IN2(U5728_n1), .QN(WX520) );
  INVX0 U5729_U2 ( .INP(WX521), .ZN(U5729_n1) );
  NOR2X0 U5729_U1 ( .IN1(n3707), .IN2(U5729_n1), .QN(WX518) );
  INVX0 U5730_U2 ( .INP(test_so1), .ZN(U5730_n1) );
  NOR2X0 U5730_U1 ( .IN1(n3707), .IN2(U5730_n1), .QN(WX516) );
  INVX0 U5731_U2 ( .INP(WX517), .ZN(U5731_n1) );
  NOR2X0 U5731_U1 ( .IN1(n3707), .IN2(U5731_n1), .QN(WX514) );
  INVX0 U5732_U2 ( .INP(WX515), .ZN(U5732_n1) );
  NOR2X0 U5732_U1 ( .IN1(n3704), .IN2(U5732_n1), .QN(WX512) );
  INVX0 U5733_U2 ( .INP(WX513), .ZN(U5733_n1) );
  NOR2X0 U5733_U1 ( .IN1(n3704), .IN2(U5733_n1), .QN(WX510) );
  INVX0 U5734_U2 ( .INP(WX511), .ZN(U5734_n1) );
  NOR2X0 U5734_U1 ( .IN1(n3704), .IN2(U5734_n1), .QN(WX508) );
  INVX0 U5735_U2 ( .INP(WX509), .ZN(U5735_n1) );
  NOR2X0 U5735_U1 ( .IN1(n3704), .IN2(U5735_n1), .QN(WX506) );
  INVX0 U5736_U2 ( .INP(WX507), .ZN(U5736_n1) );
  NOR2X0 U5736_U1 ( .IN1(n3704), .IN2(U5736_n1), .QN(WX504) );
  INVX0 U5737_U2 ( .INP(WX505), .ZN(U5737_n1) );
  NOR2X0 U5737_U1 ( .IN1(n3704), .IN2(U5737_n1), .QN(WX502) );
  INVX0 U5738_U2 ( .INP(WX503), .ZN(U5738_n1) );
  NOR2X0 U5738_U1 ( .IN1(n3704), .IN2(U5738_n1), .QN(WX500) );
  INVX0 U5739_U2 ( .INP(WX501), .ZN(U5739_n1) );
  NOR2X0 U5739_U1 ( .IN1(n3703), .IN2(U5739_n1), .QN(WX498) );
  INVX0 U5740_U2 ( .INP(WX499), .ZN(U5740_n1) );
  NOR2X0 U5740_U1 ( .IN1(n3703), .IN2(U5740_n1), .QN(WX496) );
  INVX0 U5741_U2 ( .INP(WX497), .ZN(U5741_n1) );
  NOR2X0 U5741_U1 ( .IN1(n3703), .IN2(U5741_n1), .QN(WX494) );
  INVX0 U5742_U2 ( .INP(WX495), .ZN(U5742_n1) );
  NOR2X0 U5742_U1 ( .IN1(n3703), .IN2(U5742_n1), .QN(WX492) );
  INVX0 U5743_U2 ( .INP(WX493), .ZN(U5743_n1) );
  NOR2X0 U5743_U1 ( .IN1(n3703), .IN2(U5743_n1), .QN(WX490) );
  INVX0 U5744_U2 ( .INP(WX491), .ZN(U5744_n1) );
  NOR2X0 U5744_U1 ( .IN1(n3703), .IN2(U5744_n1), .QN(WX488) );
  INVX0 U5745_U2 ( .INP(WX489), .ZN(U5745_n1) );
  NOR2X0 U5745_U1 ( .IN1(n3703), .IN2(U5745_n1), .QN(WX486) );
  INVX0 U5746_U2 ( .INP(WX487), .ZN(U5746_n1) );
  NOR2X0 U5746_U1 ( .IN1(n3703), .IN2(U5746_n1), .QN(WX484) );
  INVX0 U5747_U2 ( .INP(WX5939), .ZN(U5747_n1) );
  NOR2X0 U5747_U1 ( .IN1(n3701), .IN2(U5747_n1), .QN(WX6002) );
  INVX0 U5748_U2 ( .INP(test_so49), .ZN(U5748_n1) );
  NOR2X0 U5748_U1 ( .IN1(n3701), .IN2(U5748_n1), .QN(WX6000) );
  INVX0 U5749_U2 ( .INP(WX5935), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n3701), .IN2(U5749_n1), .QN(WX5998) );
  INVX0 U5750_U2 ( .INP(WX5933), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n3701), .IN2(U5750_n1), .QN(WX5996) );
  INVX0 U5751_U2 ( .INP(WX5931), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n3701), .IN2(U5751_n1), .QN(WX5994) );
  INVX0 U5752_U2 ( .INP(WX3269), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n3710), .IN2(U5752_n1), .QN(WX3332) );
  INVX0 U5753_U2 ( .INP(WX3265), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n3705), .IN2(U5753_n1), .QN(WX3328) );
  INVX0 U5754_U2 ( .INP(WX3263), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n3700), .IN2(U5754_n1), .QN(WX3326) );
  INVX0 U5755_U2 ( .INP(WX11179), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n3700), .IN2(U5755_n1), .QN(WX11242) );
  INVX0 U5756_U2 ( .INP(WX11177), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n3700), .IN2(U5756_n1), .QN(WX11240) );
  INVX0 U5757_U2 ( .INP(WX11175), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n3701), .IN2(U5757_n1), .QN(WX11238) );
  INVX0 U5758_U2 ( .INP(WX11173), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n3701), .IN2(U5758_n1), .QN(WX11236) );
  INVX0 U5759_U2 ( .INP(test_so96), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n3701), .IN2(U5759_n1), .QN(WX11234) );
  INVX0 U5760_U2 ( .INP(WX11169), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n3701), .IN2(U5760_n1), .QN(WX11232) );
  INVX0 U5761_U2 ( .INP(WX11167), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n3701), .IN2(U5761_n1), .QN(WX11230) );
  INVX0 U5762_U2 ( .INP(WX11165), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n3701), .IN2(U5762_n1), .QN(WX11228) );
  INVX0 U5763_U2 ( .INP(WX11163), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n3702), .IN2(U5763_n1), .QN(WX11226) );
  INVX0 U5764_U2 ( .INP(WX11161), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n3702), .IN2(U5764_n1), .QN(WX11224) );
  INVX0 U5765_U2 ( .INP(WX11159), .ZN(U5765_n1) );
  NOR2X0 U5765_U1 ( .IN1(n3702), .IN2(U5765_n1), .QN(WX11222) );
  INVX0 U5766_U2 ( .INP(WX11157), .ZN(U5766_n1) );
  NOR2X0 U5766_U1 ( .IN1(n3702), .IN2(U5766_n1), .QN(WX11220) );
  INVX0 U5767_U2 ( .INP(WX11155), .ZN(U5767_n1) );
  NOR2X0 U5767_U1 ( .IN1(n3702), .IN2(U5767_n1), .QN(WX11218) );
  INVX0 U5768_U2 ( .INP(WX11153), .ZN(U5768_n1) );
  NOR2X0 U5768_U1 ( .IN1(n3702), .IN2(U5768_n1), .QN(WX11216) );
  INVX0 U5769_U2 ( .INP(WX11151), .ZN(U5769_n1) );
  NOR2X0 U5769_U1 ( .IN1(n3702), .IN2(U5769_n1), .QN(WX11214) );
  INVX0 U5770_U2 ( .INP(WX11149), .ZN(U5770_n1) );
  NOR2X0 U5770_U1 ( .IN1(n3702), .IN2(U5770_n1), .QN(WX11212) );
  INVX0 U5771_U2 ( .INP(WX11147), .ZN(U5771_n1) );
  NOR2X0 U5771_U1 ( .IN1(n3702), .IN2(U5771_n1), .QN(WX11210) );
  INVX0 U5772_U2 ( .INP(WX11145), .ZN(U5772_n1) );
  NOR2X0 U5772_U1 ( .IN1(n3702), .IN2(U5772_n1), .QN(WX11208) );
  INVX0 U5773_U2 ( .INP(WX11143), .ZN(U5773_n1) );
  NOR2X0 U5773_U1 ( .IN1(n3702), .IN2(U5773_n1), .QN(WX11206) );
  INVX0 U5774_U2 ( .INP(WX11141), .ZN(U5774_n1) );
  NOR2X0 U5774_U1 ( .IN1(n3703), .IN2(U5774_n1), .QN(WX11204) );
  INVX0 U5775_U2 ( .INP(WX11139), .ZN(U5775_n1) );
  NOR2X0 U5775_U1 ( .IN1(n3703), .IN2(U5775_n1), .QN(WX11202) );
  INVX0 U5776_U2 ( .INP(test_so95), .ZN(U5776_n1) );
  NOR2X0 U5776_U1 ( .IN1(n3703), .IN2(U5776_n1), .QN(WX11200) );
  INVX0 U5777_U2 ( .INP(WX11135), .ZN(U5777_n1) );
  NOR2X0 U5777_U1 ( .IN1(n3704), .IN2(U5777_n1), .QN(WX11198) );
  INVX0 U5778_U2 ( .INP(WX11133), .ZN(U5778_n1) );
  NOR2X0 U5778_U1 ( .IN1(n3704), .IN2(U5778_n1), .QN(WX11196) );
  INVX0 U5779_U2 ( .INP(WX11131), .ZN(U5779_n1) );
  NOR2X0 U5779_U1 ( .IN1(n3704), .IN2(U5779_n1), .QN(WX11194) );
  INVX0 U5780_U2 ( .INP(WX11129), .ZN(U5780_n1) );
  NOR2X0 U5780_U1 ( .IN1(n3704), .IN2(U5780_n1), .QN(WX11192) );
  INVX0 U5781_U2 ( .INP(WX11127), .ZN(U5781_n1) );
  NOR2X0 U5781_U1 ( .IN1(n3705), .IN2(U5781_n1), .QN(WX11190) );
  INVX0 U5782_U2 ( .INP(WX11125), .ZN(U5782_n1) );
  NOR2X0 U5782_U1 ( .IN1(n3705), .IN2(U5782_n1), .QN(WX11188) );
  INVX0 U5783_U2 ( .INP(WX11123), .ZN(U5783_n1) );
  NOR2X0 U5783_U1 ( .IN1(n3705), .IN2(U5783_n1), .QN(WX11186) );
  INVX0 U5784_U2 ( .INP(WX11121), .ZN(U5784_n1) );
  NOR2X0 U5784_U1 ( .IN1(n3705), .IN2(U5784_n1), .QN(WX11184) );
  INVX0 U5785_U2 ( .INP(WX11119), .ZN(U5785_n1) );
  NOR2X0 U5785_U1 ( .IN1(n3705), .IN2(U5785_n1), .QN(WX11182) );
  INVX0 U5786_U2 ( .INP(WX11117), .ZN(U5786_n1) );
  NOR2X0 U5786_U1 ( .IN1(n3705), .IN2(U5786_n1), .QN(WX11180) );
  INVX0 U5787_U2 ( .INP(WX11115), .ZN(U5787_n1) );
  NOR2X0 U5787_U1 ( .IN1(n3705), .IN2(U5787_n1), .QN(WX11178) );
  INVX0 U5788_U2 ( .INP(WX11113), .ZN(U5788_n1) );
  NOR2X0 U5788_U1 ( .IN1(n3705), .IN2(U5788_n1), .QN(WX11176) );
  INVX0 U5789_U2 ( .INP(WX11111), .ZN(U5789_n1) );
  NOR2X0 U5789_U1 ( .IN1(n3705), .IN2(U5789_n1), .QN(WX11174) );
  INVX0 U5790_U2 ( .INP(WX11109), .ZN(U5790_n1) );
  NOR2X0 U5790_U1 ( .IN1(n3705), .IN2(U5790_n1), .QN(WX11172) );
  INVX0 U5791_U2 ( .INP(WX11107), .ZN(U5791_n1) );
  NOR2X0 U5791_U1 ( .IN1(n3706), .IN2(U5791_n1), .QN(WX11170) );
  INVX0 U5792_U2 ( .INP(WX11105), .ZN(U5792_n1) );
  NOR2X0 U5792_U1 ( .IN1(n3706), .IN2(U5792_n1), .QN(WX11168) );
  INVX0 U5793_U2 ( .INP(test_so94), .ZN(U5793_n1) );
  NOR2X0 U5793_U1 ( .IN1(n3706), .IN2(U5793_n1), .QN(WX11166) );
  INVX0 U5794_U2 ( .INP(WX11101), .ZN(U5794_n1) );
  NOR2X0 U5794_U1 ( .IN1(n3706), .IN2(U5794_n1), .QN(WX11164) );
  INVX0 U5795_U2 ( .INP(WX11099), .ZN(U5795_n1) );
  NOR2X0 U5795_U1 ( .IN1(n3706), .IN2(U5795_n1), .QN(WX11162) );
  INVX0 U5796_U2 ( .INP(WX11097), .ZN(U5796_n1) );
  NOR2X0 U5796_U1 ( .IN1(n3706), .IN2(U5796_n1), .QN(WX11160) );
  INVX0 U5797_U2 ( .INP(WX11095), .ZN(U5797_n1) );
  NOR2X0 U5797_U1 ( .IN1(n3706), .IN2(U5797_n1), .QN(WX11158) );
  INVX0 U5798_U2 ( .INP(WX11093), .ZN(U5798_n1) );
  NOR2X0 U5798_U1 ( .IN1(n3706), .IN2(U5798_n1), .QN(WX11156) );
  INVX0 U5799_U2 ( .INP(WX11091), .ZN(U5799_n1) );
  NOR2X0 U5799_U1 ( .IN1(n3706), .IN2(U5799_n1), .QN(WX11154) );
  INVX0 U5800_U2 ( .INP(WX11089), .ZN(U5800_n1) );
  NOR2X0 U5800_U1 ( .IN1(n3706), .IN2(U5800_n1), .QN(WX11152) );
  INVX0 U5801_U2 ( .INP(WX11087), .ZN(U5801_n1) );
  NOR2X0 U5801_U1 ( .IN1(n3706), .IN2(U5801_n1), .QN(WX11150) );
  INVX0 U5802_U2 ( .INP(WX11085), .ZN(U5802_n1) );
  NOR2X0 U5802_U1 ( .IN1(n3707), .IN2(U5802_n1), .QN(WX11148) );
  INVX0 U5803_U2 ( .INP(WX11083), .ZN(U5803_n1) );
  NOR2X0 U5803_U1 ( .IN1(n3707), .IN2(U5803_n1), .QN(WX11146) );
  INVX0 U5804_U2 ( .INP(WX11081), .ZN(U5804_n1) );
  NOR2X0 U5804_U1 ( .IN1(n3707), .IN2(U5804_n1), .QN(WX11144) );
  INVX0 U5805_U2 ( .INP(WX11079), .ZN(U5805_n1) );
  NOR2X0 U5805_U1 ( .IN1(n3707), .IN2(U5805_n1), .QN(WX11142) );
  INVX0 U5806_U2 ( .INP(WX11077), .ZN(U5806_n1) );
  NOR2X0 U5806_U1 ( .IN1(n3707), .IN2(U5806_n1), .QN(WX11140) );
  INVX0 U5807_U2 ( .INP(WX11075), .ZN(U5807_n1) );
  NOR2X0 U5807_U1 ( .IN1(n3708), .IN2(U5807_n1), .QN(WX11138) );
  INVX0 U5808_U2 ( .INP(WX11073), .ZN(U5808_n1) );
  NOR2X0 U5808_U1 ( .IN1(n3708), .IN2(U5808_n1), .QN(WX11136) );
  INVX0 U5809_U2 ( .INP(WX11071), .ZN(U5809_n1) );
  NOR2X0 U5809_U1 ( .IN1(n3709), .IN2(U5809_n1), .QN(WX11134) );
  INVX0 U5810_U2 ( .INP(test_so93), .ZN(U5810_n1) );
  NOR2X0 U5810_U1 ( .IN1(n3709), .IN2(U5810_n1), .QN(WX11132) );
  INVX0 U5811_U2 ( .INP(WX11067), .ZN(U5811_n1) );
  NOR2X0 U5811_U1 ( .IN1(n3709), .IN2(U5811_n1), .QN(WX11130) );
  INVX0 U5812_U2 ( .INP(WX11065), .ZN(U5812_n1) );
  NOR2X0 U5812_U1 ( .IN1(n3709), .IN2(U5812_n1), .QN(WX11128) );
  INVX0 U5813_U2 ( .INP(WX11063), .ZN(U5813_n1) );
  NOR2X0 U5813_U1 ( .IN1(n3709), .IN2(U5813_n1), .QN(WX11126) );
  INVX0 U5814_U2 ( .INP(WX11061), .ZN(U5814_n1) );
  NOR2X0 U5814_U1 ( .IN1(n3709), .IN2(U5814_n1), .QN(WX11124) );
  INVX0 U5815_U2 ( .INP(WX11059), .ZN(U5815_n1) );
  NOR2X0 U5815_U1 ( .IN1(n3709), .IN2(U5815_n1), .QN(WX11122) );
  INVX0 U5816_U2 ( .INP(WX11057), .ZN(U5816_n1) );
  NOR2X0 U5816_U1 ( .IN1(n3709), .IN2(U5816_n1), .QN(WX11120) );
  INVX0 U5817_U2 ( .INP(WX11055), .ZN(U5817_n1) );
  NOR2X0 U5817_U1 ( .IN1(n3709), .IN2(U5817_n1), .QN(WX11118) );
  INVX0 U5818_U2 ( .INP(WX11053), .ZN(U5818_n1) );
  NOR2X0 U5818_U1 ( .IN1(n3709), .IN2(U5818_n1), .QN(WX11116) );
  INVX0 U5819_U2 ( .INP(WX11051), .ZN(U5819_n1) );
  NOR2X0 U5819_U1 ( .IN1(n3709), .IN2(U5819_n1), .QN(WX11114) );
  INVX0 U5820_U2 ( .INP(WX11049), .ZN(U5820_n1) );
  NOR2X0 U5820_U1 ( .IN1(n3710), .IN2(U5820_n1), .QN(WX11112) );
  INVX0 U5821_U2 ( .INP(WX11047), .ZN(U5821_n1) );
  NOR2X0 U5821_U1 ( .IN1(n3710), .IN2(U5821_n1), .QN(WX11110) );
  INVX0 U5822_U2 ( .INP(WX11045), .ZN(U5822_n1) );
  NOR2X0 U5822_U1 ( .IN1(n3710), .IN2(U5822_n1), .QN(WX11108) );
  INVX0 U5823_U2 ( .INP(WX11043), .ZN(U5823_n1) );
  NOR2X0 U5823_U1 ( .IN1(n3710), .IN2(U5823_n1), .QN(WX11106) );
  INVX0 U5824_U2 ( .INP(WX11041), .ZN(U5824_n1) );
  NOR2X0 U5824_U1 ( .IN1(n3710), .IN2(U5824_n1), .QN(WX11104) );
  INVX0 U5825_U2 ( .INP(WX11039), .ZN(U5825_n1) );
  NOR2X0 U5825_U1 ( .IN1(n3710), .IN2(U5825_n1), .QN(WX11102) );
  INVX0 U5826_U2 ( .INP(WX11037), .ZN(U5826_n1) );
  NOR2X0 U5826_U1 ( .IN1(n3710), .IN2(U5826_n1), .QN(WX11100) );
  INVX0 U5827_U2 ( .INP(test_so92), .ZN(U5827_n1) );
  NOR2X0 U5827_U1 ( .IN1(n3710), .IN2(U5827_n1), .QN(WX11098) );
  INVX0 U5828_U2 ( .INP(WX11033), .ZN(U5828_n1) );
  NOR2X0 U5828_U1 ( .IN1(n3695), .IN2(U5828_n1), .QN(WX11096) );
  INVX0 U5829_U2 ( .INP(WX11031), .ZN(U5829_n1) );
  NOR2X0 U5829_U1 ( .IN1(n3689), .IN2(U5829_n1), .QN(WX11094) );
  INVX0 U5830_U2 ( .INP(WX11029), .ZN(U5830_n1) );
  NOR2X0 U5830_U1 ( .IN1(n3689), .IN2(U5830_n1), .QN(WX11092) );
  INVX0 U5831_U2 ( .INP(WX11027), .ZN(U5831_n1) );
  NOR2X0 U5831_U1 ( .IN1(n3689), .IN2(U5831_n1), .QN(WX11090) );
  INVX0 U5832_U2 ( .INP(WX11025), .ZN(U5832_n1) );
  NOR2X0 U5832_U1 ( .IN1(n3689), .IN2(U5832_n1), .QN(WX11088) );
  INVX0 U5833_U2 ( .INP(WX11023), .ZN(U5833_n1) );
  NOR2X0 U5833_U1 ( .IN1(n3690), .IN2(U5833_n1), .QN(WX11086) );
  INVX0 U5834_U2 ( .INP(WX11021), .ZN(U5834_n1) );
  NOR2X0 U5834_U1 ( .IN1(n3690), .IN2(U5834_n1), .QN(WX11084) );
  INVX0 U5835_U2 ( .INP(WX9886), .ZN(U5835_n1) );
  NOR2X0 U5835_U1 ( .IN1(n3690), .IN2(U5835_n1), .QN(WX9949) );
  INVX0 U5836_U2 ( .INP(WX9884), .ZN(U5836_n1) );
  NOR2X0 U5836_U1 ( .IN1(n3690), .IN2(U5836_n1), .QN(WX9947) );
  INVX0 U5837_U2 ( .INP(WX9882), .ZN(U5837_n1) );
  NOR2X0 U5837_U1 ( .IN1(n3690), .IN2(U5837_n1), .QN(WX9945) );
  INVX0 U5838_U2 ( .INP(WX9880), .ZN(U5838_n1) );
  NOR2X0 U5838_U1 ( .IN1(n3690), .IN2(U5838_n1), .QN(WX9943) );
  INVX0 U5839_U2 ( .INP(WX9878), .ZN(U5839_n1) );
  NOR2X0 U5839_U1 ( .IN1(n3690), .IN2(U5839_n1), .QN(WX9941) );
  INVX0 U5840_U2 ( .INP(WX9876), .ZN(U5840_n1) );
  NOR2X0 U5840_U1 ( .IN1(n3690), .IN2(U5840_n1), .QN(WX9939) );
  INVX0 U5841_U2 ( .INP(WX9874), .ZN(U5841_n1) );
  NOR2X0 U5841_U1 ( .IN1(n3690), .IN2(U5841_n1), .QN(WX9937) );
  INVX0 U5842_U2 ( .INP(WX9872), .ZN(U5842_n1) );
  NOR2X0 U5842_U1 ( .IN1(n3690), .IN2(U5842_n1), .QN(WX9935) );
  INVX0 U5843_U2 ( .INP(WX9870), .ZN(U5843_n1) );
  NOR2X0 U5843_U1 ( .IN1(n3690), .IN2(U5843_n1), .QN(WX9933) );
  INVX0 U5844_U2 ( .INP(WX9868), .ZN(U5844_n1) );
  NOR2X0 U5844_U1 ( .IN1(n3692), .IN2(U5844_n1), .QN(WX9931) );
  INVX0 U5845_U2 ( .INP(WX9866), .ZN(U5845_n1) );
  NOR2X0 U5845_U1 ( .IN1(n3692), .IN2(U5845_n1), .QN(WX9929) );
  INVX0 U5846_U2 ( .INP(WX9864), .ZN(U5846_n1) );
  NOR2X0 U5846_U1 ( .IN1(n3692), .IN2(U5846_n1), .QN(WX9927) );
  INVX0 U5847_U2 ( .INP(WX9862), .ZN(U5847_n1) );
  NOR2X0 U5847_U1 ( .IN1(n3692), .IN2(U5847_n1), .QN(WX9925) );
  INVX0 U5848_U2 ( .INP(WX9860), .ZN(U5848_n1) );
  NOR2X0 U5848_U1 ( .IN1(n3692), .IN2(U5848_n1), .QN(WX9923) );
  INVX0 U5849_U2 ( .INP(WX9858), .ZN(U5849_n1) );
  NOR2X0 U5849_U1 ( .IN1(n3692), .IN2(U5849_n1), .QN(WX9921) );
  INVX0 U5850_U2 ( .INP(WX9856), .ZN(U5850_n1) );
  NOR2X0 U5850_U1 ( .IN1(n3692), .IN2(U5850_n1), .QN(WX9919) );
  INVX0 U5851_U2 ( .INP(test_so84), .ZN(U5851_n1) );
  NOR2X0 U5851_U1 ( .IN1(n3692), .IN2(U5851_n1), .QN(WX9917) );
  INVX0 U5852_U2 ( .INP(WX9852), .ZN(U5852_n1) );
  NOR2X0 U5852_U1 ( .IN1(n3692), .IN2(U5852_n1), .QN(WX9915) );
  INVX0 U5853_U2 ( .INP(WX9850), .ZN(U5853_n1) );
  NOR2X0 U5853_U1 ( .IN1(n3692), .IN2(U5853_n1), .QN(WX9913) );
  INVX0 U5854_U2 ( .INP(WX9848), .ZN(U5854_n1) );
  NOR2X0 U5854_U1 ( .IN1(n3692), .IN2(U5854_n1), .QN(WX9911) );
  INVX0 U5855_U2 ( .INP(WX9846), .ZN(U5855_n1) );
  NOR2X0 U5855_U1 ( .IN1(n3693), .IN2(U5855_n1), .QN(WX9909) );
  INVX0 U5856_U2 ( .INP(WX9844), .ZN(U5856_n1) );
  NOR2X0 U5856_U1 ( .IN1(n3693), .IN2(U5856_n1), .QN(WX9907) );
  INVX0 U5857_U2 ( .INP(WX9842), .ZN(U5857_n1) );
  NOR2X0 U5857_U1 ( .IN1(n3693), .IN2(U5857_n1), .QN(WX9905) );
  INVX0 U5858_U2 ( .INP(WX9840), .ZN(U5858_n1) );
  NOR2X0 U5858_U1 ( .IN1(n3693), .IN2(U5858_n1), .QN(WX9903) );
  INVX0 U5859_U2 ( .INP(WX9838), .ZN(U5859_n1) );
  NOR2X0 U5859_U1 ( .IN1(n3693), .IN2(U5859_n1), .QN(WX9901) );
  INVX0 U5860_U2 ( .INP(WX9836), .ZN(U5860_n1) );
  NOR2X0 U5860_U1 ( .IN1(n3693), .IN2(U5860_n1), .QN(WX9899) );
  INVX0 U5861_U2 ( .INP(WX9834), .ZN(U5861_n1) );
  NOR2X0 U5861_U1 ( .IN1(n3693), .IN2(U5861_n1), .QN(WX9897) );
  INVX0 U5862_U2 ( .INP(WX9832), .ZN(U5862_n1) );
  NOR2X0 U5862_U1 ( .IN1(n3693), .IN2(U5862_n1), .QN(WX9895) );
  INVX0 U5863_U2 ( .INP(WX9830), .ZN(U5863_n1) );
  NOR2X0 U5863_U1 ( .IN1(n3693), .IN2(U5863_n1), .QN(WX9893) );
  INVX0 U5864_U2 ( .INP(WX9828), .ZN(U5864_n1) );
  NOR2X0 U5864_U1 ( .IN1(n3693), .IN2(U5864_n1), .QN(WX9891) );
  INVX0 U5865_U2 ( .INP(WX9826), .ZN(U5865_n1) );
  NOR2X0 U5865_U1 ( .IN1(n3693), .IN2(U5865_n1), .QN(WX9889) );
  INVX0 U5866_U2 ( .INP(WX9824), .ZN(U5866_n1) );
  NOR2X0 U5866_U1 ( .IN1(n3694), .IN2(U5866_n1), .QN(WX9887) );
  INVX0 U5867_U2 ( .INP(WX9822), .ZN(U5867_n1) );
  NOR2X0 U5867_U1 ( .IN1(n3694), .IN2(U5867_n1), .QN(WX9885) );
  INVX0 U5868_U2 ( .INP(test_so83), .ZN(U5868_n1) );
  NOR2X0 U5868_U1 ( .IN1(n3694), .IN2(U5868_n1), .QN(WX9883) );
  INVX0 U5869_U2 ( .INP(WX9818), .ZN(U5869_n1) );
  NOR2X0 U5869_U1 ( .IN1(n3694), .IN2(U5869_n1), .QN(WX9881) );
  INVX0 U5870_U2 ( .INP(WX9816), .ZN(U5870_n1) );
  NOR2X0 U5870_U1 ( .IN1(n3694), .IN2(U5870_n1), .QN(WX9879) );
  INVX0 U5871_U2 ( .INP(WX9814), .ZN(U5871_n1) );
  NOR2X0 U5871_U1 ( .IN1(n3694), .IN2(U5871_n1), .QN(WX9877) );
  INVX0 U5872_U2 ( .INP(WX9812), .ZN(U5872_n1) );
  NOR2X0 U5872_U1 ( .IN1(n3694), .IN2(U5872_n1), .QN(WX9875) );
  INVX0 U5873_U2 ( .INP(WX9810), .ZN(U5873_n1) );
  NOR2X0 U5873_U1 ( .IN1(n3694), .IN2(U5873_n1), .QN(WX9873) );
  INVX0 U5874_U2 ( .INP(WX9808), .ZN(U5874_n1) );
  NOR2X0 U5874_U1 ( .IN1(n3694), .IN2(U5874_n1), .QN(WX9871) );
  INVX0 U5875_U2 ( .INP(WX9806), .ZN(U5875_n1) );
  NOR2X0 U5875_U1 ( .IN1(n3694), .IN2(U5875_n1), .QN(WX9869) );
  INVX0 U5876_U2 ( .INP(WX9804), .ZN(U5876_n1) );
  NOR2X0 U5876_U1 ( .IN1(n3694), .IN2(U5876_n1), .QN(WX9867) );
  INVX0 U5877_U2 ( .INP(WX9802), .ZN(U5877_n1) );
  NOR2X0 U5877_U1 ( .IN1(n3695), .IN2(U5877_n1), .QN(WX9865) );
  INVX0 U5878_U2 ( .INP(WX9800), .ZN(U5878_n1) );
  NOR2X0 U5878_U1 ( .IN1(n3695), .IN2(U5878_n1), .QN(WX9863) );
  INVX0 U5879_U2 ( .INP(WX9798), .ZN(U5879_n1) );
  NOR2X0 U5879_U1 ( .IN1(n3695), .IN2(U5879_n1), .QN(WX9861) );
  INVX0 U5880_U2 ( .INP(WX9796), .ZN(U5880_n1) );
  NOR2X0 U5880_U1 ( .IN1(n3695), .IN2(U5880_n1), .QN(WX9859) );
  INVX0 U5881_U2 ( .INP(WX9794), .ZN(U5881_n1) );
  NOR2X0 U5881_U1 ( .IN1(n3695), .IN2(U5881_n1), .QN(WX9857) );
  INVX0 U5882_U2 ( .INP(WX9792), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(n3695), .IN2(U5882_n1), .QN(WX9855) );
  INVX0 U5883_U2 ( .INP(WX9790), .ZN(U5883_n1) );
  NOR2X0 U5883_U1 ( .IN1(n3695), .IN2(U5883_n1), .QN(WX9853) );
  INVX0 U5884_U2 ( .INP(WX9788), .ZN(U5884_n1) );
  NOR2X0 U5884_U1 ( .IN1(n3695), .IN2(U5884_n1), .QN(WX9851) );
  INVX0 U5885_U2 ( .INP(test_so82), .ZN(U5885_n1) );
  NOR2X0 U5885_U1 ( .IN1(n3695), .IN2(U5885_n1), .QN(WX9849) );
  INVX0 U5886_U2 ( .INP(WX9784), .ZN(U5886_n1) );
  NOR2X0 U5886_U1 ( .IN1(n3695), .IN2(U5886_n1), .QN(WX9847) );
  INVX0 U5887_U2 ( .INP(WX9782), .ZN(U5887_n1) );
  NOR2X0 U5887_U1 ( .IN1(n3696), .IN2(U5887_n1), .QN(WX9845) );
  INVX0 U5888_U2 ( .INP(WX9780), .ZN(U5888_n1) );
  NOR2X0 U5888_U1 ( .IN1(n3696), .IN2(U5888_n1), .QN(WX9843) );
  INVX0 U5889_U2 ( .INP(WX9778), .ZN(U5889_n1) );
  NOR2X0 U5889_U1 ( .IN1(n3696), .IN2(U5889_n1), .QN(WX9841) );
  INVX0 U5890_U2 ( .INP(WX9776), .ZN(U5890_n1) );
  NOR2X0 U5890_U1 ( .IN1(n3696), .IN2(U5890_n1), .QN(WX9839) );
  INVX0 U5891_U2 ( .INP(WX9774), .ZN(U5891_n1) );
  NOR2X0 U5891_U1 ( .IN1(n3696), .IN2(U5891_n1), .QN(WX9837) );
  INVX0 U5892_U2 ( .INP(WX9772), .ZN(U5892_n1) );
  NOR2X0 U5892_U1 ( .IN1(n3696), .IN2(U5892_n1), .QN(WX9835) );
  INVX0 U5893_U2 ( .INP(WX9770), .ZN(U5893_n1) );
  NOR2X0 U5893_U1 ( .IN1(n3696), .IN2(U5893_n1), .QN(WX9833) );
  INVX0 U5894_U2 ( .INP(WX9768), .ZN(U5894_n1) );
  NOR2X0 U5894_U1 ( .IN1(n3696), .IN2(U5894_n1), .QN(WX9831) );
  INVX0 U5895_U2 ( .INP(WX9766), .ZN(U5895_n1) );
  NOR2X0 U5895_U1 ( .IN1(n3696), .IN2(U5895_n1), .QN(WX9829) );
  INVX0 U5896_U2 ( .INP(WX9764), .ZN(U5896_n1) );
  NOR2X0 U5896_U1 ( .IN1(n3696), .IN2(U5896_n1), .QN(WX9827) );
  INVX0 U5897_U2 ( .INP(WX9762), .ZN(U5897_n1) );
  NOR2X0 U5897_U1 ( .IN1(n3696), .IN2(U5897_n1), .QN(WX9825) );
  INVX0 U5898_U2 ( .INP(WX9760), .ZN(U5898_n1) );
  NOR2X0 U5898_U1 ( .IN1(n3697), .IN2(U5898_n1), .QN(WX9823) );
  INVX0 U5899_U2 ( .INP(WX9758), .ZN(U5899_n1) );
  NOR2X0 U5899_U1 ( .IN1(n3697), .IN2(U5899_n1), .QN(WX9821) );
  INVX0 U5900_U2 ( .INP(WX9756), .ZN(U5900_n1) );
  NOR2X0 U5900_U1 ( .IN1(n3697), .IN2(U5900_n1), .QN(WX9819) );
  INVX0 U5901_U2 ( .INP(WX9754), .ZN(U5901_n1) );
  NOR2X0 U5901_U1 ( .IN1(n3697), .IN2(U5901_n1), .QN(WX9817) );
  INVX0 U5902_U2 ( .INP(test_so81), .ZN(U5902_n1) );
  NOR2X0 U5902_U1 ( .IN1(n3697), .IN2(U5902_n1), .QN(WX9815) );
  INVX0 U5903_U2 ( .INP(WX9750), .ZN(U5903_n1) );
  NOR2X0 U5903_U1 ( .IN1(n3697), .IN2(U5903_n1), .QN(WX9813) );
  INVX0 U5904_U2 ( .INP(WX9748), .ZN(U5904_n1) );
  NOR2X0 U5904_U1 ( .IN1(n3697), .IN2(U5904_n1), .QN(WX9811) );
  INVX0 U5905_U2 ( .INP(WX9746), .ZN(U5905_n1) );
  NOR2X0 U5905_U1 ( .IN1(n3697), .IN2(U5905_n1), .QN(WX9809) );
  INVX0 U5906_U2 ( .INP(WX9744), .ZN(U5906_n1) );
  NOR2X0 U5906_U1 ( .IN1(n3697), .IN2(U5906_n1), .QN(WX9807) );
  INVX0 U5907_U2 ( .INP(WX9742), .ZN(U5907_n1) );
  NOR2X0 U5907_U1 ( .IN1(n3697), .IN2(U5907_n1), .QN(WX9805) );
  INVX0 U5908_U2 ( .INP(WX9740), .ZN(U5908_n1) );
  NOR2X0 U5908_U1 ( .IN1(n3697), .IN2(U5908_n1), .QN(WX9803) );
  INVX0 U5909_U2 ( .INP(WX9738), .ZN(U5909_n1) );
  NOR2X0 U5909_U1 ( .IN1(n3698), .IN2(U5909_n1), .QN(WX9801) );
  INVX0 U5910_U2 ( .INP(WX9736), .ZN(U5910_n1) );
  NOR2X0 U5910_U1 ( .IN1(n3698), .IN2(U5910_n1), .QN(WX9799) );
  INVX0 U5911_U2 ( .INP(WX9734), .ZN(U5911_n1) );
  NOR2X0 U5911_U1 ( .IN1(n3698), .IN2(U5911_n1), .QN(WX9797) );
  INVX0 U5912_U2 ( .INP(WX9732), .ZN(U5912_n1) );
  NOR2X0 U5912_U1 ( .IN1(n3698), .IN2(U5912_n1), .QN(WX9795) );
  INVX0 U5913_U2 ( .INP(WX9730), .ZN(U5913_n1) );
  NOR2X0 U5913_U1 ( .IN1(n3698), .IN2(U5913_n1), .QN(WX9793) );
  INVX0 U5914_U2 ( .INP(WX9728), .ZN(U5914_n1) );
  NOR2X0 U5914_U1 ( .IN1(n3698), .IN2(U5914_n1), .QN(WX9791) );
  INVX0 U5915_U2 ( .INP(WX8593), .ZN(U5915_n1) );
  NOR2X0 U5915_U1 ( .IN1(n3698), .IN2(U5915_n1), .QN(WX8656) );
  INVX0 U5916_U2 ( .INP(WX8591), .ZN(U5916_n1) );
  NOR2X0 U5916_U1 ( .IN1(n3698), .IN2(U5916_n1), .QN(WX8654) );
  INVX0 U5917_U2 ( .INP(WX8589), .ZN(U5917_n1) );
  NOR2X0 U5917_U1 ( .IN1(n3698), .IN2(U5917_n1), .QN(WX8652) );
  INVX0 U5918_U2 ( .INP(WX8587), .ZN(U5918_n1) );
  NOR2X0 U5918_U1 ( .IN1(n3698), .IN2(U5918_n1), .QN(WX8650) );
  INVX0 U5919_U2 ( .INP(WX8585), .ZN(U5919_n1) );
  NOR2X0 U5919_U1 ( .IN1(n3698), .IN2(U5919_n1), .QN(WX8648) );
  INVX0 U5920_U2 ( .INP(WX8583), .ZN(U5920_n1) );
  NOR2X0 U5920_U1 ( .IN1(n3699), .IN2(U5920_n1), .QN(WX8646) );
  INVX0 U5921_U2 ( .INP(WX8581), .ZN(U5921_n1) );
  NOR2X0 U5921_U1 ( .IN1(n3699), .IN2(U5921_n1), .QN(WX8644) );
  INVX0 U5922_U2 ( .INP(WX8579), .ZN(U5922_n1) );
  NOR2X0 U5922_U1 ( .IN1(n3699), .IN2(U5922_n1), .QN(WX8642) );
  INVX0 U5923_U2 ( .INP(WX8577), .ZN(U5923_n1) );
  NOR2X0 U5923_U1 ( .IN1(n3699), .IN2(U5923_n1), .QN(WX8640) );
  INVX0 U5924_U2 ( .INP(WX8575), .ZN(U5924_n1) );
  NOR2X0 U5924_U1 ( .IN1(n3699), .IN2(U5924_n1), .QN(WX8638) );
  INVX0 U5925_U2 ( .INP(WX8573), .ZN(U5925_n1) );
  NOR2X0 U5925_U1 ( .IN1(n3699), .IN2(U5925_n1), .QN(WX8636) );
  INVX0 U5926_U2 ( .INP(test_so73), .ZN(U5926_n1) );
  NOR2X0 U5926_U1 ( .IN1(n3699), .IN2(U5926_n1), .QN(WX8634) );
  INVX0 U5927_U2 ( .INP(WX8569), .ZN(U5927_n1) );
  NOR2X0 U5927_U1 ( .IN1(n3699), .IN2(U5927_n1), .QN(WX8632) );
  INVX0 U5928_U2 ( .INP(WX8567), .ZN(U5928_n1) );
  NOR2X0 U5928_U1 ( .IN1(n3699), .IN2(U5928_n1), .QN(WX8630) );
  INVX0 U5929_U2 ( .INP(WX8565), .ZN(U5929_n1) );
  NOR2X0 U5929_U1 ( .IN1(n3699), .IN2(U5929_n1), .QN(WX8628) );
  INVX0 U5930_U2 ( .INP(WX8563), .ZN(U5930_n1) );
  NOR2X0 U5930_U1 ( .IN1(n3699), .IN2(U5930_n1), .QN(WX8626) );
  INVX0 U5931_U2 ( .INP(WX8561), .ZN(U5931_n1) );
  NOR2X0 U5931_U1 ( .IN1(n3700), .IN2(U5931_n1), .QN(WX8624) );
  INVX0 U5932_U2 ( .INP(WX8559), .ZN(U5932_n1) );
  NOR2X0 U5932_U1 ( .IN1(n3700), .IN2(U5932_n1), .QN(WX8622) );
  INVX0 U5933_U2 ( .INP(WX8557), .ZN(U5933_n1) );
  NOR2X0 U5933_U1 ( .IN1(n3700), .IN2(U5933_n1), .QN(WX8620) );
  INVX0 U5934_U2 ( .INP(WX8555), .ZN(U5934_n1) );
  NOR2X0 U5934_U1 ( .IN1(n3700), .IN2(U5934_n1), .QN(WX8618) );
  INVX0 U5935_U2 ( .INP(WX8553), .ZN(U5935_n1) );
  NOR2X0 U5935_U1 ( .IN1(n3700), .IN2(U5935_n1), .QN(WX8616) );
  INVX0 U5936_U2 ( .INP(WX8551), .ZN(U5936_n1) );
  NOR2X0 U5936_U1 ( .IN1(n3700), .IN2(U5936_n1), .QN(WX8614) );
  INVX0 U5937_U2 ( .INP(WX8549), .ZN(U5937_n1) );
  NOR2X0 U5937_U1 ( .IN1(n3700), .IN2(U5937_n1), .QN(WX8612) );
  INVX0 U5938_U2 ( .INP(WX8547), .ZN(U5938_n1) );
  NOR2X0 U5938_U1 ( .IN1(n3700), .IN2(U5938_n1), .QN(WX8610) );
  INVX0 U5939_U2 ( .INP(WX8545), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n3725), .IN2(U5939_n1), .QN(WX8608) );
  INVX0 U5940_U2 ( .INP(WX8543), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n3731), .IN2(U5940_n1), .QN(WX8606) );
  INVX0 U5941_U2 ( .INP(WX8541), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n3732), .IN2(U5941_n1), .QN(WX8604) );
  INVX0 U5942_U2 ( .INP(WX8539), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n3732), .IN2(U5942_n1), .QN(WX8602) );
  INVX0 U5943_U2 ( .INP(test_so72), .ZN(U5943_n1) );
  NOR2X0 U5943_U1 ( .IN1(n3731), .IN2(U5943_n1), .QN(WX8600) );
  INVX0 U5944_U2 ( .INP(WX8535), .ZN(U5944_n1) );
  NOR2X0 U5944_U1 ( .IN1(n3732), .IN2(U5944_n1), .QN(WX8598) );
  INVX0 U5945_U2 ( .INP(WX8533), .ZN(U5945_n1) );
  NOR2X0 U5945_U1 ( .IN1(n3732), .IN2(U5945_n1), .QN(WX8596) );
  INVX0 U5946_U2 ( .INP(WX8531), .ZN(U5946_n1) );
  NOR2X0 U5946_U1 ( .IN1(n3731), .IN2(U5946_n1), .QN(WX8594) );
  INVX0 U5947_U2 ( .INP(WX8529), .ZN(U5947_n1) );
  NOR2X0 U5947_U1 ( .IN1(n3730), .IN2(U5947_n1), .QN(WX8592) );
  INVX0 U5948_U2 ( .INP(WX8527), .ZN(U5948_n1) );
  NOR2X0 U5948_U1 ( .IN1(n3732), .IN2(U5948_n1), .QN(WX8590) );
  INVX0 U5949_U2 ( .INP(WX8525), .ZN(U5949_n1) );
  NOR2X0 U5949_U1 ( .IN1(n3731), .IN2(U5949_n1), .QN(WX8588) );
  INVX0 U5950_U2 ( .INP(WX8523), .ZN(U5950_n1) );
  NOR2X0 U5950_U1 ( .IN1(n3732), .IN2(U5950_n1), .QN(WX8586) );
  INVX0 U5951_U2 ( .INP(WX8521), .ZN(U5951_n1) );
  NOR2X0 U5951_U1 ( .IN1(n3732), .IN2(U5951_n1), .QN(WX8584) );
  INVX0 U5952_U2 ( .INP(WX8519), .ZN(U5952_n1) );
  NOR2X0 U5952_U1 ( .IN1(n3728), .IN2(U5952_n1), .QN(WX8582) );
  INVX0 U5953_U2 ( .INP(WX8517), .ZN(U5953_n1) );
  NOR2X0 U5953_U1 ( .IN1(n3732), .IN2(U5953_n1), .QN(WX8580) );
  INVX0 U5954_U2 ( .INP(WX8515), .ZN(U5954_n1) );
  NOR2X0 U5954_U1 ( .IN1(n3728), .IN2(U5954_n1), .QN(WX8578) );
  INVX0 U5955_U2 ( .INP(WX8513), .ZN(U5955_n1) );
  NOR2X0 U5955_U1 ( .IN1(n3728), .IN2(U5955_n1), .QN(WX8576) );
  INVX0 U5956_U2 ( .INP(WX8511), .ZN(U5956_n1) );
  NOR2X0 U5956_U1 ( .IN1(n3728), .IN2(U5956_n1), .QN(WX8574) );
  INVX0 U5957_U2 ( .INP(WX8509), .ZN(U5957_n1) );
  NOR2X0 U5957_U1 ( .IN1(n3728), .IN2(U5957_n1), .QN(WX8572) );
  INVX0 U5958_U2 ( .INP(WX8507), .ZN(U5958_n1) );
  NOR2X0 U5958_U1 ( .IN1(n3728), .IN2(U5958_n1), .QN(WX8570) );
  INVX0 U5959_U2 ( .INP(WX8505), .ZN(U5959_n1) );
  NOR2X0 U5959_U1 ( .IN1(n3727), .IN2(U5959_n1), .QN(WX8568) );
  INVX0 U5960_U2 ( .INP(test_so71), .ZN(U5960_n1) );
  NOR2X0 U5960_U1 ( .IN1(n3727), .IN2(U5960_n1), .QN(WX8566) );
  INVX0 U5961_U2 ( .INP(WX8501), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n3727), .IN2(U5961_n1), .QN(WX8564) );
  INVX0 U5962_U2 ( .INP(WX8499), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n3726), .IN2(U5962_n1), .QN(WX8562) );
  INVX0 U5963_U2 ( .INP(WX8497), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n3726), .IN2(U5963_n1), .QN(WX8560) );
  INVX0 U5964_U2 ( .INP(WX8495), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n3726), .IN2(U5964_n1), .QN(WX8558) );
  INVX0 U5965_U2 ( .INP(WX8493), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n3726), .IN2(U5965_n1), .QN(WX8556) );
  INVX0 U5966_U2 ( .INP(WX8491), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n3725), .IN2(U5966_n1), .QN(WX8554) );
  INVX0 U5967_U2 ( .INP(WX8489), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n3725), .IN2(U5967_n1), .QN(WX8552) );
  INVX0 U5968_U2 ( .INP(WX8487), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n3725), .IN2(U5968_n1), .QN(WX8550) );
  INVX0 U5969_U2 ( .INP(WX8485), .ZN(U5969_n1) );
  NOR2X0 U5969_U1 ( .IN1(n3725), .IN2(U5969_n1), .QN(WX8548) );
  INVX0 U5970_U2 ( .INP(WX8483), .ZN(U5970_n1) );
  NOR2X0 U5970_U1 ( .IN1(n3725), .IN2(U5970_n1), .QN(WX8546) );
  INVX0 U5971_U2 ( .INP(WX8481), .ZN(U5971_n1) );
  NOR2X0 U5971_U1 ( .IN1(n3725), .IN2(U5971_n1), .QN(WX8544) );
  INVX0 U5972_U2 ( .INP(WX8479), .ZN(U5972_n1) );
  NOR2X0 U5972_U1 ( .IN1(n3725), .IN2(U5972_n1), .QN(WX8542) );
  INVX0 U5973_U2 ( .INP(WX8477), .ZN(U5973_n1) );
  NOR2X0 U5973_U1 ( .IN1(n3725), .IN2(U5973_n1), .QN(WX8540) );
  INVX0 U5974_U2 ( .INP(WX8475), .ZN(U5974_n1) );
  NOR2X0 U5974_U1 ( .IN1(n3725), .IN2(U5974_n1), .QN(WX8538) );
  INVX0 U5975_U2 ( .INP(WX8473), .ZN(U5975_n1) );
  NOR2X0 U5975_U1 ( .IN1(n3725), .IN2(U5975_n1), .QN(WX8536) );
  INVX0 U5976_U2 ( .INP(WX8471), .ZN(U5976_n1) );
  NOR2X0 U5976_U1 ( .IN1(n3724), .IN2(U5976_n1), .QN(WX8534) );
  INVX0 U5977_U2 ( .INP(test_so70), .ZN(U5977_n1) );
  NOR2X0 U5977_U1 ( .IN1(n3724), .IN2(U5977_n1), .QN(WX8532) );
  INVX0 U5978_U2 ( .INP(WX8467), .ZN(U5978_n1) );
  NOR2X0 U5978_U1 ( .IN1(n3724), .IN2(U5978_n1), .QN(WX8530) );
  INVX0 U5979_U2 ( .INP(WX8465), .ZN(U5979_n1) );
  NOR2X0 U5979_U1 ( .IN1(n3724), .IN2(U5979_n1), .QN(WX8528) );
  INVX0 U5980_U2 ( .INP(WX8463), .ZN(U5980_n1) );
  NOR2X0 U5980_U1 ( .IN1(n3724), .IN2(U5980_n1), .QN(WX8526) );
  INVX0 U5981_U2 ( .INP(WX8461), .ZN(U5981_n1) );
  NOR2X0 U5981_U1 ( .IN1(n3724), .IN2(U5981_n1), .QN(WX8524) );
  INVX0 U5982_U2 ( .INP(WX8459), .ZN(U5982_n1) );
  NOR2X0 U5982_U1 ( .IN1(n3724), .IN2(U5982_n1), .QN(WX8522) );
  INVX0 U5983_U2 ( .INP(WX8457), .ZN(U5983_n1) );
  NOR2X0 U5983_U1 ( .IN1(n3724), .IN2(U5983_n1), .QN(WX8520) );
  INVX0 U5984_U2 ( .INP(WX8455), .ZN(U5984_n1) );
  NOR2X0 U5984_U1 ( .IN1(n3722), .IN2(U5984_n1), .QN(WX8518) );
  INVX0 U5985_U2 ( .INP(WX8453), .ZN(U5985_n1) );
  NOR2X0 U5985_U1 ( .IN1(n3723), .IN2(U5985_n1), .QN(WX8516) );
  INVX0 U5986_U2 ( .INP(WX8451), .ZN(U5986_n1) );
  NOR2X0 U5986_U1 ( .IN1(n3723), .IN2(U5986_n1), .QN(WX8514) );
  INVX0 U5987_U2 ( .INP(WX8449), .ZN(U5987_n1) );
  NOR2X0 U5987_U1 ( .IN1(n3723), .IN2(U5987_n1), .QN(WX8512) );
  INVX0 U5988_U2 ( .INP(WX8447), .ZN(U5988_n1) );
  NOR2X0 U5988_U1 ( .IN1(n3723), .IN2(U5988_n1), .QN(WX8510) );
  INVX0 U5989_U2 ( .INP(WX8445), .ZN(U5989_n1) );
  NOR2X0 U5989_U1 ( .IN1(n3723), .IN2(U5989_n1), .QN(WX8508) );
  INVX0 U5990_U2 ( .INP(WX8443), .ZN(U5990_n1) );
  NOR2X0 U5990_U1 ( .IN1(n3723), .IN2(U5990_n1), .QN(WX8506) );
  INVX0 U5991_U2 ( .INP(WX8441), .ZN(U5991_n1) );
  NOR2X0 U5991_U1 ( .IN1(n3723), .IN2(U5991_n1), .QN(WX8504) );
  INVX0 U5992_U2 ( .INP(WX8439), .ZN(U5992_n1) );
  NOR2X0 U5992_U1 ( .IN1(n3723), .IN2(U5992_n1), .QN(WX8502) );
  INVX0 U5993_U2 ( .INP(WX8437), .ZN(U5993_n1) );
  NOR2X0 U5993_U1 ( .IN1(n3723), .IN2(U5993_n1), .QN(WX8500) );
  INVX0 U5994_U2 ( .INP(test_so69), .ZN(U5994_n1) );
  NOR2X0 U5994_U1 ( .IN1(n3723), .IN2(U5994_n1), .QN(WX8498) );
  INVX0 U5995_U2 ( .INP(WX7300), .ZN(U5995_n1) );
  NOR2X0 U5995_U1 ( .IN1(n3723), .IN2(U5995_n1), .QN(WX7363) );
  INVX0 U5996_U2 ( .INP(WX7298), .ZN(U5996_n1) );
  NOR2X0 U5996_U1 ( .IN1(n3724), .IN2(U5996_n1), .QN(WX7361) );
  INVX0 U5997_U2 ( .INP(WX7296), .ZN(U5997_n1) );
  NOR2X0 U5997_U1 ( .IN1(n3724), .IN2(U5997_n1), .QN(WX7359) );
  INVX0 U5998_U2 ( .INP(WX7294), .ZN(U5998_n1) );
  NOR2X0 U5998_U1 ( .IN1(n3724), .IN2(U5998_n1), .QN(WX7357) );
  INVX0 U5999_U2 ( .INP(WX7292), .ZN(U5999_n1) );
  NOR2X0 U5999_U1 ( .IN1(n3726), .IN2(U5999_n1), .QN(WX7355) );
  INVX0 U6000_U2 ( .INP(WX7290), .ZN(U6000_n1) );
  NOR2X0 U6000_U1 ( .IN1(n3726), .IN2(U6000_n1), .QN(WX7353) );
  INVX0 U6001_U2 ( .INP(test_so62), .ZN(U6001_n1) );
  NOR2X0 U6001_U1 ( .IN1(n3726), .IN2(U6001_n1), .QN(WX7351) );
  INVX0 U6002_U2 ( .INP(WX7286), .ZN(U6002_n1) );
  NOR2X0 U6002_U1 ( .IN1(n3726), .IN2(U6002_n1), .QN(WX7349) );
  INVX0 U6003_U2 ( .INP(WX7284), .ZN(U6003_n1) );
  NOR2X0 U6003_U1 ( .IN1(n3726), .IN2(U6003_n1), .QN(WX7347) );
  INVX0 U6004_U2 ( .INP(WX7282), .ZN(U6004_n1) );
  NOR2X0 U6004_U1 ( .IN1(n3726), .IN2(U6004_n1), .QN(WX7345) );
  INVX0 U6005_U2 ( .INP(WX7280), .ZN(U6005_n1) );
  NOR2X0 U6005_U1 ( .IN1(n3726), .IN2(U6005_n1), .QN(WX7343) );
  INVX0 U6006_U2 ( .INP(WX7278), .ZN(U6006_n1) );
  NOR2X0 U6006_U1 ( .IN1(n3727), .IN2(U6006_n1), .QN(WX7341) );
  INVX0 U6007_U2 ( .INP(WX7276), .ZN(U6007_n1) );
  NOR2X0 U6007_U1 ( .IN1(n3727), .IN2(U6007_n1), .QN(WX7339) );
  INVX0 U6008_U2 ( .INP(WX7274), .ZN(U6008_n1) );
  NOR2X0 U6008_U1 ( .IN1(n3727), .IN2(U6008_n1), .QN(WX7337) );
  INVX0 U6009_U2 ( .INP(WX7272), .ZN(U6009_n1) );
  NOR2X0 U6009_U1 ( .IN1(n3727), .IN2(U6009_n1), .QN(WX7335) );
  INVX0 U6010_U2 ( .INP(WX7270), .ZN(U6010_n1) );
  NOR2X0 U6010_U1 ( .IN1(n3727), .IN2(U6010_n1), .QN(WX7333) );
  INVX0 U6011_U2 ( .INP(WX7268), .ZN(U6011_n1) );
  NOR2X0 U6011_U1 ( .IN1(n3727), .IN2(U6011_n1), .QN(WX7331) );
  INVX0 U6012_U2 ( .INP(WX7266), .ZN(U6012_n1) );
  NOR2X0 U6012_U1 ( .IN1(n3727), .IN2(U6012_n1), .QN(WX7329) );
  INVX0 U6013_U2 ( .INP(WX7264), .ZN(U6013_n1) );
  NOR2X0 U6013_U1 ( .IN1(n3727), .IN2(U6013_n1), .QN(WX7327) );
  INVX0 U6014_U2 ( .INP(WX7262), .ZN(U6014_n1) );
  NOR2X0 U6014_U1 ( .IN1(n3728), .IN2(U6014_n1), .QN(WX7325) );
  INVX0 U6015_U2 ( .INP(WX7260), .ZN(U6015_n1) );
  NOR2X0 U6015_U1 ( .IN1(n3728), .IN2(U6015_n1), .QN(WX7323) );
  INVX0 U6016_U2 ( .INP(WX7258), .ZN(U6016_n1) );
  NOR2X0 U6016_U1 ( .IN1(n3728), .IN2(U6016_n1), .QN(WX7321) );
  INVX0 U6017_U2 ( .INP(WX7256), .ZN(U6017_n1) );
  NOR2X0 U6017_U1 ( .IN1(n3728), .IN2(U6017_n1), .QN(WX7319) );
  INVX0 U6018_U2 ( .INP(test_so61), .ZN(U6018_n1) );
  NOR2X0 U6018_U1 ( .IN1(n3728), .IN2(U6018_n1), .QN(WX7317) );
  INVX0 U6019_U2 ( .INP(WX7252), .ZN(U6019_n1) );
  NOR2X0 U6019_U1 ( .IN1(n3729), .IN2(U6019_n1), .QN(WX7315) );
  INVX0 U6020_U2 ( .INP(WX7250), .ZN(U6020_n1) );
  NOR2X0 U6020_U1 ( .IN1(n3729), .IN2(U6020_n1), .QN(WX7313) );
  INVX0 U6021_U2 ( .INP(WX7248), .ZN(U6021_n1) );
  NOR2X0 U6021_U1 ( .IN1(n3729), .IN2(U6021_n1), .QN(WX7311) );
  INVX0 U6022_U2 ( .INP(WX7246), .ZN(U6022_n1) );
  NOR2X0 U6022_U1 ( .IN1(n3729), .IN2(U6022_n1), .QN(WX7309) );
  INVX0 U6023_U2 ( .INP(WX7244), .ZN(U6023_n1) );
  NOR2X0 U6023_U1 ( .IN1(n3729), .IN2(U6023_n1), .QN(WX7307) );
  INVX0 U6024_U2 ( .INP(WX7242), .ZN(U6024_n1) );
  NOR2X0 U6024_U1 ( .IN1(n3729), .IN2(U6024_n1), .QN(WX7305) );
  INVX0 U6025_U2 ( .INP(WX7240), .ZN(U6025_n1) );
  NOR2X0 U6025_U1 ( .IN1(n3730), .IN2(U6025_n1), .QN(WX7303) );
  INVX0 U6026_U2 ( .INP(WX7238), .ZN(U6026_n1) );
  NOR2X0 U6026_U1 ( .IN1(n3729), .IN2(U6026_n1), .QN(WX7301) );
  INVX0 U6027_U2 ( .INP(WX7236), .ZN(U6027_n1) );
  NOR2X0 U6027_U1 ( .IN1(n3730), .IN2(U6027_n1), .QN(WX7299) );
  INVX0 U6028_U2 ( .INP(WX7234), .ZN(U6028_n1) );
  NOR2X0 U6028_U1 ( .IN1(n3730), .IN2(U6028_n1), .QN(WX7297) );
  INVX0 U6029_U2 ( .INP(WX7232), .ZN(U6029_n1) );
  NOR2X0 U6029_U1 ( .IN1(n3729), .IN2(U6029_n1), .QN(WX7295) );
  INVX0 U6030_U2 ( .INP(WX7230), .ZN(U6030_n1) );
  NOR2X0 U6030_U1 ( .IN1(n3730), .IN2(U6030_n1), .QN(WX7293) );
  INVX0 U6031_U2 ( .INP(WX7228), .ZN(U6031_n1) );
  NOR2X0 U6031_U1 ( .IN1(n3730), .IN2(U6031_n1), .QN(WX7291) );
  INVX0 U6032_U2 ( .INP(WX7226), .ZN(U6032_n1) );
  NOR2X0 U6032_U1 ( .IN1(n3729), .IN2(U6032_n1), .QN(WX7289) );
  INVX0 U6033_U2 ( .INP(WX7224), .ZN(U6033_n1) );
  NOR2X0 U6033_U1 ( .IN1(n3730), .IN2(U6033_n1), .QN(WX7287) );
  INVX0 U6034_U2 ( .INP(WX7222), .ZN(U6034_n1) );
  NOR2X0 U6034_U1 ( .IN1(n3730), .IN2(U6034_n1), .QN(WX7285) );
  INVX0 U6035_U2 ( .INP(test_so60), .ZN(U6035_n1) );
  NOR2X0 U6035_U1 ( .IN1(n3729), .IN2(U6035_n1), .QN(WX7283) );
  INVX0 U6036_U2 ( .INP(WX7218), .ZN(U6036_n1) );
  NOR2X0 U6036_U1 ( .IN1(n3731), .IN2(U6036_n1), .QN(WX7281) );
  INVX0 U6037_U2 ( .INP(WX7216), .ZN(U6037_n1) );
  NOR2X0 U6037_U1 ( .IN1(n3731), .IN2(U6037_n1), .QN(WX7279) );
  INVX0 U6038_U2 ( .INP(WX7214), .ZN(U6038_n1) );
  NOR2X0 U6038_U1 ( .IN1(n3730), .IN2(U6038_n1), .QN(WX7277) );
  INVX0 U6039_U2 ( .INP(WX7212), .ZN(U6039_n1) );
  NOR2X0 U6039_U1 ( .IN1(n3731), .IN2(U6039_n1), .QN(WX7275) );
  INVX0 U6040_U2 ( .INP(WX7210), .ZN(U6040_n1) );
  NOR2X0 U6040_U1 ( .IN1(n3731), .IN2(U6040_n1), .QN(WX7273) );
  INVX0 U6041_U2 ( .INP(WX7208), .ZN(U6041_n1) );
  NOR2X0 U6041_U1 ( .IN1(n3730), .IN2(U6041_n1), .QN(WX7271) );
  INVX0 U6042_U2 ( .INP(WX7206), .ZN(U6042_n1) );
  NOR2X0 U6042_U1 ( .IN1(n3731), .IN2(U6042_n1), .QN(WX7269) );
  INVX0 U6043_U2 ( .INP(WX7204), .ZN(U6043_n1) );
  NOR2X0 U6043_U1 ( .IN1(n3731), .IN2(U6043_n1), .QN(WX7267) );
  INVX0 U6044_U2 ( .INP(WX7202), .ZN(U6044_n1) );
  NOR2X0 U6044_U1 ( .IN1(n3730), .IN2(U6044_n1), .QN(WX7265) );
  INVX0 U6045_U2 ( .INP(WX7200), .ZN(U6045_n1) );
  NOR2X0 U6045_U1 ( .IN1(n3732), .IN2(U6045_n1), .QN(WX7263) );
  INVX0 U6046_U2 ( .INP(WX7198), .ZN(U6046_n1) );
  NOR2X0 U6046_U1 ( .IN1(n3731), .IN2(U6046_n1), .QN(WX7261) );
  INVX0 U6047_U2 ( .INP(WX7196), .ZN(U6047_n1) );
  NOR2X0 U6047_U1 ( .IN1(n3732), .IN2(U6047_n1), .QN(WX7259) );
  INVX0 U6048_U2 ( .INP(WX7194), .ZN(U6048_n1) );
  NOR2X0 U6048_U1 ( .IN1(n3732), .IN2(U6048_n1), .QN(WX7257) );
  INVX0 U6049_U2 ( .INP(WX7192), .ZN(U6049_n1) );
  NOR2X0 U6049_U1 ( .IN1(n3729), .IN2(U6049_n1), .QN(WX7255) );
  INVX0 U6050_U2 ( .INP(WX7190), .ZN(U6050_n1) );
  NOR2X0 U6050_U1 ( .IN1(n3716), .IN2(U6050_n1), .QN(WX7253) );
  INVX0 U6051_U2 ( .INP(WX7188), .ZN(U6051_n1) );
  NOR2X0 U6051_U1 ( .IN1(n3710), .IN2(U6051_n1), .QN(WX7251) );
  INVX0 U6052_U2 ( .INP(test_so59), .ZN(U6052_n1) );
  NOR2X0 U6052_U1 ( .IN1(n3710), .IN2(U6052_n1), .QN(WX7249) );
  INVX0 U6053_U2 ( .INP(WX7184), .ZN(U6053_n1) );
  NOR2X0 U6053_U1 ( .IN1(n3711), .IN2(U6053_n1), .QN(WX7247) );
  INVX0 U6054_U2 ( .INP(WX7182), .ZN(U6054_n1) );
  NOR2X0 U6054_U1 ( .IN1(n3711), .IN2(U6054_n1), .QN(WX7245) );
  INVX0 U6055_U2 ( .INP(WX7180), .ZN(U6055_n1) );
  NOR2X0 U6055_U1 ( .IN1(n3711), .IN2(U6055_n1), .QN(WX7243) );
  INVX0 U6056_U2 ( .INP(WX7178), .ZN(U6056_n1) );
  NOR2X0 U6056_U1 ( .IN1(n3711), .IN2(U6056_n1), .QN(WX7241) );
  INVX0 U6057_U2 ( .INP(WX7176), .ZN(U6057_n1) );
  NOR2X0 U6057_U1 ( .IN1(n3711), .IN2(U6057_n1), .QN(WX7239) );
  INVX0 U6058_U2 ( .INP(WX7174), .ZN(U6058_n1) );
  NOR2X0 U6058_U1 ( .IN1(n3711), .IN2(U6058_n1), .QN(WX7237) );
  INVX0 U6059_U2 ( .INP(WX7172), .ZN(U6059_n1) );
  NOR2X0 U6059_U1 ( .IN1(n3711), .IN2(U6059_n1), .QN(WX7235) );
  INVX0 U6060_U2 ( .INP(WX7170), .ZN(U6060_n1) );
  NOR2X0 U6060_U1 ( .IN1(n3711), .IN2(U6060_n1), .QN(WX7233) );
  INVX0 U6061_U2 ( .INP(WX7168), .ZN(U6061_n1) );
  NOR2X0 U6061_U1 ( .IN1(n3711), .IN2(U6061_n1), .QN(WX7231) );
  INVX0 U6062_U2 ( .INP(WX7166), .ZN(U6062_n1) );
  NOR2X0 U6062_U1 ( .IN1(n3711), .IN2(U6062_n1), .QN(WX7229) );
  INVX0 U6063_U2 ( .INP(WX7164), .ZN(U6063_n1) );
  NOR2X0 U6063_U1 ( .IN1(n3711), .IN2(U6063_n1), .QN(WX7227) );
  INVX0 U6064_U2 ( .INP(WX7162), .ZN(U6064_n1) );
  NOR2X0 U6064_U1 ( .IN1(n3712), .IN2(U6064_n1), .QN(WX7225) );
  INVX0 U6065_U2 ( .INP(WX7160), .ZN(U6065_n1) );
  NOR2X0 U6065_U1 ( .IN1(n3712), .IN2(U6065_n1), .QN(WX7223) );
  INVX0 U6066_U2 ( .INP(WX7158), .ZN(U6066_n1) );
  NOR2X0 U6066_U1 ( .IN1(n3712), .IN2(U6066_n1), .QN(WX7221) );
  INVX0 U6067_U2 ( .INP(WX7156), .ZN(U6067_n1) );
  NOR2X0 U6067_U1 ( .IN1(n3712), .IN2(U6067_n1), .QN(WX7219) );
  INVX0 U6068_U2 ( .INP(WX7154), .ZN(U6068_n1) );
  NOR2X0 U6068_U1 ( .IN1(n3712), .IN2(U6068_n1), .QN(WX7217) );
  INVX0 U6069_U2 ( .INP(test_so58), .ZN(U6069_n1) );
  NOR2X0 U6069_U1 ( .IN1(n3712), .IN2(U6069_n1), .QN(WX7215) );
  INVX0 U6070_U2 ( .INP(WX7150), .ZN(U6070_n1) );
  NOR2X0 U6070_U1 ( .IN1(n3712), .IN2(U6070_n1), .QN(WX7213) );
  INVX0 U6071_U2 ( .INP(WX7148), .ZN(U6071_n1) );
  NOR2X0 U6071_U1 ( .IN1(n3712), .IN2(U6071_n1), .QN(WX7211) );
  INVX0 U6072_U2 ( .INP(WX7146), .ZN(U6072_n1) );
  NOR2X0 U6072_U1 ( .IN1(n3712), .IN2(U6072_n1), .QN(WX7209) );
  INVX0 U6073_U2 ( .INP(WX7144), .ZN(U6073_n1) );
  NOR2X0 U6073_U1 ( .IN1(n3712), .IN2(U6073_n1), .QN(WX7207) );
  INVX0 U6074_U2 ( .INP(WX7142), .ZN(U6074_n1) );
  NOR2X0 U6074_U1 ( .IN1(n3712), .IN2(U6074_n1), .QN(WX7205) );
  INVX0 U6075_U2 ( .INP(WX6007), .ZN(U6075_n1) );
  NOR2X0 U6075_U1 ( .IN1(n3714), .IN2(U6075_n1), .QN(WX6070) );
  INVX0 U6076_U2 ( .INP(test_so51), .ZN(U6076_n1) );
  NOR2X0 U6076_U1 ( .IN1(n3714), .IN2(U6076_n1), .QN(WX6068) );
  INVX0 U6077_U2 ( .INP(WX6003), .ZN(U6077_n1) );
  NOR2X0 U6077_U1 ( .IN1(n3714), .IN2(U6077_n1), .QN(WX6066) );
  INVX0 U6078_U2 ( .INP(WX6001), .ZN(U6078_n1) );
  NOR2X0 U6078_U1 ( .IN1(n3714), .IN2(U6078_n1), .QN(WX6064) );
  INVX0 U6079_U2 ( .INP(WX5999), .ZN(U6079_n1) );
  NOR2X0 U6079_U1 ( .IN1(n3714), .IN2(U6079_n1), .QN(WX6062) );
  INVX0 U6080_U2 ( .INP(WX5997), .ZN(U6080_n1) );
  NOR2X0 U6080_U1 ( .IN1(n3714), .IN2(U6080_n1), .QN(WX6060) );
  INVX0 U6081_U2 ( .INP(WX5995), .ZN(U6081_n1) );
  NOR2X0 U6081_U1 ( .IN1(n3714), .IN2(U6081_n1), .QN(WX6058) );
  INVX0 U6082_U2 ( .INP(WX5993), .ZN(U6082_n1) );
  NOR2X0 U6082_U1 ( .IN1(n3714), .IN2(U6082_n1), .QN(WX6056) );
  INVX0 U6083_U2 ( .INP(WX5991), .ZN(U6083_n1) );
  NOR2X0 U6083_U1 ( .IN1(n3714), .IN2(U6083_n1), .QN(WX6054) );
  INVX0 U6084_U2 ( .INP(WX5989), .ZN(U6084_n1) );
  NOR2X0 U6084_U1 ( .IN1(n3714), .IN2(U6084_n1), .QN(WX6052) );
  INVX0 U6085_U2 ( .INP(WX5987), .ZN(U6085_n1) );
  NOR2X0 U6085_U1 ( .IN1(n3714), .IN2(U6085_n1), .QN(WX6050) );
  INVX0 U6086_U2 ( .INP(WX5985), .ZN(U6086_n1) );
  NOR2X0 U6086_U1 ( .IN1(n3715), .IN2(U6086_n1), .QN(WX6048) );
  INVX0 U6087_U2 ( .INP(WX5983), .ZN(U6087_n1) );
  NOR2X0 U6087_U1 ( .IN1(n3715), .IN2(U6087_n1), .QN(WX6046) );
  INVX0 U6088_U2 ( .INP(WX5981), .ZN(U6088_n1) );
  NOR2X0 U6088_U1 ( .IN1(n3715), .IN2(U6088_n1), .QN(WX6044) );
  INVX0 U6089_U2 ( .INP(WX5979), .ZN(U6089_n1) );
  NOR2X0 U6089_U1 ( .IN1(n3715), .IN2(U6089_n1), .QN(WX6042) );
  INVX0 U6090_U2 ( .INP(WX5977), .ZN(U6090_n1) );
  NOR2X0 U6090_U1 ( .IN1(n3715), .IN2(U6090_n1), .QN(WX6040) );
  INVX0 U6091_U2 ( .INP(WX5975), .ZN(U6091_n1) );
  NOR2X0 U6091_U1 ( .IN1(n3715), .IN2(U6091_n1), .QN(WX6038) );
  INVX0 U6092_U2 ( .INP(WX5973), .ZN(U6092_n1) );
  NOR2X0 U6092_U1 ( .IN1(n3715), .IN2(U6092_n1), .QN(WX6036) );
  INVX0 U6093_U2 ( .INP(test_so50), .ZN(U6093_n1) );
  NOR2X0 U6093_U1 ( .IN1(n3715), .IN2(U6093_n1), .QN(WX6034) );
  INVX0 U6094_U2 ( .INP(WX5969), .ZN(U6094_n1) );
  NOR2X0 U6094_U1 ( .IN1(n3715), .IN2(U6094_n1), .QN(WX6032) );
  INVX0 U6095_U2 ( .INP(WX5967), .ZN(U6095_n1) );
  NOR2X0 U6095_U1 ( .IN1(n3715), .IN2(U6095_n1), .QN(WX6030) );
  INVX0 U6096_U2 ( .INP(WX5965), .ZN(U6096_n1) );
  NOR2X0 U6096_U1 ( .IN1(n3715), .IN2(U6096_n1), .QN(WX6028) );
  INVX0 U6097_U2 ( .INP(WX5963), .ZN(U6097_n1) );
  NOR2X0 U6097_U1 ( .IN1(n3716), .IN2(U6097_n1), .QN(WX6026) );
  INVX0 U6098_U2 ( .INP(WX5961), .ZN(U6098_n1) );
  NOR2X0 U6098_U1 ( .IN1(n3716), .IN2(U6098_n1), .QN(WX6024) );
  INVX0 U6099_U2 ( .INP(WX5959), .ZN(U6099_n1) );
  NOR2X0 U6099_U1 ( .IN1(n3716), .IN2(U6099_n1), .QN(WX6022) );
  INVX0 U6100_U2 ( .INP(WX5957), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n3716), .IN2(U6100_n1), .QN(WX6020) );
  INVX0 U6101_U2 ( .INP(WX5955), .ZN(U6101_n1) );
  NOR2X0 U6101_U1 ( .IN1(n3716), .IN2(U6101_n1), .QN(WX6018) );
  INVX0 U6102_U2 ( .INP(WX5953), .ZN(U6102_n1) );
  NOR2X0 U6102_U1 ( .IN1(n3716), .IN2(U6102_n1), .QN(WX6016) );
  INVX0 U6103_U2 ( .INP(WX5951), .ZN(U6103_n1) );
  NOR2X0 U6103_U1 ( .IN1(n3716), .IN2(U6103_n1), .QN(WX6014) );
  INVX0 U6104_U2 ( .INP(WX5949), .ZN(U6104_n1) );
  NOR2X0 U6104_U1 ( .IN1(n3716), .IN2(U6104_n1), .QN(WX6012) );
  INVX0 U6105_U2 ( .INP(WX5947), .ZN(U6105_n1) );
  NOR2X0 U6105_U1 ( .IN1(n3716), .IN2(U6105_n1), .QN(WX6010) );
  INVX0 U6106_U2 ( .INP(WX5945), .ZN(U6106_n1) );
  NOR2X0 U6106_U1 ( .IN1(n3716), .IN2(U6106_n1), .QN(WX6008) );
  INVX0 U6107_U2 ( .INP(WX5943), .ZN(U6107_n1) );
  NOR2X0 U6107_U1 ( .IN1(n3718), .IN2(U6107_n1), .QN(WX6006) );
  INVX0 U6108_U2 ( .INP(WX5941), .ZN(U6108_n1) );
  NOR2X0 U6108_U1 ( .IN1(n3718), .IN2(U6108_n1), .QN(WX6004) );
  INVX0 U6109_U2 ( .INP(WX5929), .ZN(U6109_n1) );
  NOR2X0 U6109_U1 ( .IN1(n3718), .IN2(U6109_n1), .QN(WX5992) );
  INVX0 U6110_U2 ( .INP(WX5927), .ZN(U6110_n1) );
  NOR2X0 U6110_U1 ( .IN1(n3718), .IN2(U6110_n1), .QN(WX5990) );
  INVX0 U6111_U2 ( .INP(WX5925), .ZN(U6111_n1) );
  NOR2X0 U6111_U1 ( .IN1(n3718), .IN2(U6111_n1), .QN(WX5988) );
  INVX0 U6112_U2 ( .INP(WX5923), .ZN(U6112_n1) );
  NOR2X0 U6112_U1 ( .IN1(n3718), .IN2(U6112_n1), .QN(WX5986) );
  INVX0 U6113_U2 ( .INP(WX5921), .ZN(U6113_n1) );
  NOR2X0 U6113_U1 ( .IN1(n3718), .IN2(U6113_n1), .QN(WX5984) );
  INVX0 U6114_U2 ( .INP(WX5919), .ZN(U6114_n1) );
  NOR2X0 U6114_U1 ( .IN1(n3718), .IN2(U6114_n1), .QN(WX5982) );
  INVX0 U6115_U2 ( .INP(WX5917), .ZN(U6115_n1) );
  NOR2X0 U6115_U1 ( .IN1(n3718), .IN2(U6115_n1), .QN(WX5980) );
  INVX0 U6116_U2 ( .INP(WX5915), .ZN(U6116_n1) );
  NOR2X0 U6116_U1 ( .IN1(n3718), .IN2(U6116_n1), .QN(WX5978) );
  INVX0 U6117_U2 ( .INP(WX5913), .ZN(U6117_n1) );
  NOR2X0 U6117_U1 ( .IN1(n3718), .IN2(U6117_n1), .QN(WX5976) );
  INVX0 U6118_U2 ( .INP(WX5911), .ZN(U6118_n1) );
  NOR2X0 U6118_U1 ( .IN1(n3719), .IN2(U6118_n1), .QN(WX5974) );
  INVX0 U6119_U2 ( .INP(WX5909), .ZN(U6119_n1) );
  NOR2X0 U6119_U1 ( .IN1(n3719), .IN2(U6119_n1), .QN(WX5972) );
  INVX0 U6120_U2 ( .INP(WX5907), .ZN(U6120_n1) );
  NOR2X0 U6120_U1 ( .IN1(n3719), .IN2(U6120_n1), .QN(WX5970) );
  INVX0 U6121_U2 ( .INP(WX5905), .ZN(U6121_n1) );
  NOR2X0 U6121_U1 ( .IN1(n3719), .IN2(U6121_n1), .QN(WX5968) );
  INVX0 U6122_U2 ( .INP(test_so48), .ZN(U6122_n1) );
  NOR2X0 U6122_U1 ( .IN1(n3719), .IN2(U6122_n1), .QN(WX5966) );
  INVX0 U6123_U2 ( .INP(WX5901), .ZN(U6123_n1) );
  NOR2X0 U6123_U1 ( .IN1(n3719), .IN2(U6123_n1), .QN(WX5964) );
  INVX0 U6124_U2 ( .INP(WX5899), .ZN(U6124_n1) );
  NOR2X0 U6124_U1 ( .IN1(n3719), .IN2(U6124_n1), .QN(WX5962) );
  INVX0 U6125_U2 ( .INP(WX5897), .ZN(U6125_n1) );
  NOR2X0 U6125_U1 ( .IN1(n3719), .IN2(U6125_n1), .QN(WX5960) );
  INVX0 U6126_U2 ( .INP(WX5895), .ZN(U6126_n1) );
  NOR2X0 U6126_U1 ( .IN1(n3719), .IN2(U6126_n1), .QN(WX5958) );
  INVX0 U6127_U2 ( .INP(WX5893), .ZN(U6127_n1) );
  NOR2X0 U6127_U1 ( .IN1(n3719), .IN2(U6127_n1), .QN(WX5956) );
  INVX0 U6128_U2 ( .INP(WX5891), .ZN(U6128_n1) );
  NOR2X0 U6128_U1 ( .IN1(n3719), .IN2(U6128_n1), .QN(WX5954) );
  INVX0 U6129_U2 ( .INP(WX5889), .ZN(U6129_n1) );
  NOR2X0 U6129_U1 ( .IN1(n3720), .IN2(U6129_n1), .QN(WX5952) );
  INVX0 U6130_U2 ( .INP(WX5887), .ZN(U6130_n1) );
  NOR2X0 U6130_U1 ( .IN1(n3720), .IN2(U6130_n1), .QN(WX5950) );
  INVX0 U6131_U2 ( .INP(WX5885), .ZN(U6131_n1) );
  NOR2X0 U6131_U1 ( .IN1(n3720), .IN2(U6131_n1), .QN(WX5948) );
  INVX0 U6132_U2 ( .INP(WX5883), .ZN(U6132_n1) );
  NOR2X0 U6132_U1 ( .IN1(n3720), .IN2(U6132_n1), .QN(WX5946) );
  INVX0 U6133_U2 ( .INP(WX5881), .ZN(U6133_n1) );
  NOR2X0 U6133_U1 ( .IN1(n3720), .IN2(U6133_n1), .QN(WX5944) );
  INVX0 U6134_U2 ( .INP(WX5879), .ZN(U6134_n1) );
  NOR2X0 U6134_U1 ( .IN1(n3720), .IN2(U6134_n1), .QN(WX5942) );
  INVX0 U6135_U2 ( .INP(WX5877), .ZN(U6135_n1) );
  NOR2X0 U6135_U1 ( .IN1(n3720), .IN2(U6135_n1), .QN(WX5940) );
  INVX0 U6136_U2 ( .INP(WX5875), .ZN(U6136_n1) );
  NOR2X0 U6136_U1 ( .IN1(n3720), .IN2(U6136_n1), .QN(WX5938) );
  INVX0 U6137_U2 ( .INP(WX5873), .ZN(U6137_n1) );
  NOR2X0 U6137_U1 ( .IN1(n3720), .IN2(U6137_n1), .QN(WX5936) );
  INVX0 U6138_U2 ( .INP(WX5871), .ZN(U6138_n1) );
  NOR2X0 U6138_U1 ( .IN1(n3720), .IN2(U6138_n1), .QN(WX5934) );
  INVX0 U6139_U2 ( .INP(test_so47), .ZN(U6139_n1) );
  NOR2X0 U6139_U1 ( .IN1(n3720), .IN2(U6139_n1), .QN(WX5932) );
  INVX0 U6140_U2 ( .INP(WX5867), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n3721), .IN2(U6140_n1), .QN(WX5930) );
  INVX0 U6141_U2 ( .INP(WX5865), .ZN(U6141_n1) );
  NOR2X0 U6141_U1 ( .IN1(n3721), .IN2(U6141_n1), .QN(WX5928) );
  INVX0 U6142_U2 ( .INP(WX5863), .ZN(U6142_n1) );
  NOR2X0 U6142_U1 ( .IN1(n3721), .IN2(U6142_n1), .QN(WX5926) );
  INVX0 U6143_U2 ( .INP(WX5861), .ZN(U6143_n1) );
  NOR2X0 U6143_U1 ( .IN1(n3721), .IN2(U6143_n1), .QN(WX5924) );
  INVX0 U6144_U2 ( .INP(WX5859), .ZN(U6144_n1) );
  NOR2X0 U6144_U1 ( .IN1(n3722), .IN2(U6144_n1), .QN(WX5922) );
  INVX0 U6145_U2 ( .INP(WX5857), .ZN(U6145_n1) );
  NOR2X0 U6145_U1 ( .IN1(n3721), .IN2(U6145_n1), .QN(WX5920) );
  INVX0 U6146_U2 ( .INP(WX5855), .ZN(U6146_n1) );
  NOR2X0 U6146_U1 ( .IN1(n3721), .IN2(U6146_n1), .QN(WX5918) );
  INVX0 U6147_U2 ( .INP(WX5853), .ZN(U6147_n1) );
  NOR2X0 U6147_U1 ( .IN1(n3721), .IN2(U6147_n1), .QN(WX5916) );
  INVX0 U6148_U2 ( .INP(WX5851), .ZN(U6148_n1) );
  NOR2X0 U6148_U1 ( .IN1(n3721), .IN2(U6148_n1), .QN(WX5914) );
  INVX0 U6149_U2 ( .INP(WX5849), .ZN(U6149_n1) );
  NOR2X0 U6149_U1 ( .IN1(n3721), .IN2(U6149_n1), .QN(WX5912) );
  INVX0 U6150_U2 ( .INP(WX4714), .ZN(U6150_n1) );
  NOR2X0 U6150_U1 ( .IN1(n3721), .IN2(U6150_n1), .QN(WX4777) );
  INVX0 U6151_U2 ( .INP(WX4712), .ZN(U6151_n1) );
  NOR2X0 U6151_U1 ( .IN1(n3722), .IN2(U6151_n1), .QN(WX4775) );
  INVX0 U6152_U2 ( .INP(WX4710), .ZN(U6152_n1) );
  NOR2X0 U6152_U1 ( .IN1(n3722), .IN2(U6152_n1), .QN(WX4773) );
  INVX0 U6153_U2 ( .INP(WX4708), .ZN(U6153_n1) );
  NOR2X0 U6153_U1 ( .IN1(n3722), .IN2(U6153_n1), .QN(WX4771) );
  INVX0 U6154_U2 ( .INP(WX4706), .ZN(U6154_n1) );
  NOR2X0 U6154_U1 ( .IN1(n3722), .IN2(U6154_n1), .QN(WX4769) );
  INVX0 U6155_U2 ( .INP(WX4704), .ZN(U6155_n1) );
  NOR2X0 U6155_U1 ( .IN1(n3722), .IN2(U6155_n1), .QN(WX4767) );
  INVX0 U6156_U2 ( .INP(WX4702), .ZN(U6156_n1) );
  NOR2X0 U6156_U1 ( .IN1(n3722), .IN2(U6156_n1), .QN(WX4765) );
  INVX0 U6157_U2 ( .INP(WX4700), .ZN(U6157_n1) );
  NOR2X0 U6157_U1 ( .IN1(n3722), .IN2(U6157_n1), .QN(WX4763) );
  INVX0 U6158_U2 ( .INP(WX4698), .ZN(U6158_n1) );
  NOR2X0 U6158_U1 ( .IN1(n3722), .IN2(U6158_n1), .QN(WX4761) );
  INVX0 U6159_U2 ( .INP(WX4696), .ZN(U6159_n1) );
  NOR2X0 U6159_U1 ( .IN1(n3722), .IN2(U6159_n1), .QN(WX4759) );
  INVX0 U6160_U2 ( .INP(WX4694), .ZN(U6160_n1) );
  NOR2X0 U6160_U1 ( .IN1(n3721), .IN2(U6160_n1), .QN(WX4757) );
  INVX0 U6161_U2 ( .INP(WX4692), .ZN(U6161_n1) );
  NOR2X0 U6161_U1 ( .IN1(n3674), .IN2(U6161_n1), .QN(WX4755) );
  INVX0 U6162_U2 ( .INP(WX4690), .ZN(U6162_n1) );
  NOR2X0 U6162_U1 ( .IN1(n3674), .IN2(U6162_n1), .QN(WX4753) );
  INVX0 U6163_U2 ( .INP(test_so39), .ZN(U6163_n1) );
  NOR2X0 U6163_U1 ( .IN1(n3674), .IN2(U6163_n1), .QN(WX4751) );
  INVX0 U6164_U2 ( .INP(WX4686), .ZN(U6164_n1) );
  NOR2X0 U6164_U1 ( .IN1(n3674), .IN2(U6164_n1), .QN(WX4749) );
  INVX0 U6165_U2 ( .INP(WX4684), .ZN(U6165_n1) );
  NOR2X0 U6165_U1 ( .IN1(n3674), .IN2(U6165_n1), .QN(WX4747) );
  INVX0 U6166_U2 ( .INP(WX4682), .ZN(U6166_n1) );
  NOR2X0 U6166_U1 ( .IN1(n3674), .IN2(U6166_n1), .QN(WX4745) );
  INVX0 U6167_U2 ( .INP(WX4680), .ZN(U6167_n1) );
  NOR2X0 U6167_U1 ( .IN1(n3674), .IN2(U6167_n1), .QN(WX4743) );
  INVX0 U6168_U2 ( .INP(WX4678), .ZN(U6168_n1) );
  NOR2X0 U6168_U1 ( .IN1(n3674), .IN2(U6168_n1), .QN(WX4741) );
  INVX0 U6169_U2 ( .INP(WX4676), .ZN(U6169_n1) );
  NOR2X0 U6169_U1 ( .IN1(n3674), .IN2(U6169_n1), .QN(WX4739) );
  INVX0 U6170_U2 ( .INP(WX4674), .ZN(U6170_n1) );
  NOR2X0 U6170_U1 ( .IN1(n3674), .IN2(U6170_n1), .QN(WX4737) );
  INVX0 U6171_U2 ( .INP(WX4672), .ZN(U6171_n1) );
  NOR2X0 U6171_U1 ( .IN1(n3673), .IN2(U6171_n1), .QN(WX4735) );
  INVX0 U6172_U2 ( .INP(WX4670), .ZN(U6172_n1) );
  NOR2X0 U6172_U1 ( .IN1(n3673), .IN2(U6172_n1), .QN(WX4733) );
  INVX0 U6173_U2 ( .INP(WX4668), .ZN(U6173_n1) );
  NOR2X0 U6173_U1 ( .IN1(n3673), .IN2(U6173_n1), .QN(WX4731) );
  INVX0 U6174_U2 ( .INP(WX4666), .ZN(U6174_n1) );
  NOR2X0 U6174_U1 ( .IN1(n3673), .IN2(U6174_n1), .QN(WX4729) );
  INVX0 U6175_U2 ( .INP(WX4664), .ZN(U6175_n1) );
  NOR2X0 U6175_U1 ( .IN1(n3673), .IN2(U6175_n1), .QN(WX4727) );
  INVX0 U6176_U2 ( .INP(WX4662), .ZN(U6176_n1) );
  NOR2X0 U6176_U1 ( .IN1(n3673), .IN2(U6176_n1), .QN(WX4725) );
  INVX0 U6177_U2 ( .INP(WX4660), .ZN(U6177_n1) );
  NOR2X0 U6177_U1 ( .IN1(n3673), .IN2(U6177_n1), .QN(WX4723) );
  INVX0 U6178_U2 ( .INP(WX4658), .ZN(U6178_n1) );
  NOR2X0 U6178_U1 ( .IN1(n3673), .IN2(U6178_n1), .QN(WX4721) );
  INVX0 U6179_U2 ( .INP(WX4656), .ZN(U6179_n1) );
  NOR2X0 U6179_U1 ( .IN1(n3673), .IN2(U6179_n1), .QN(WX4719) );
  INVX0 U6180_U2 ( .INP(test_so38), .ZN(U6180_n1) );
  NOR2X0 U6180_U1 ( .IN1(n3673), .IN2(U6180_n1), .QN(WX4717) );
  INVX0 U6181_U2 ( .INP(WX4652), .ZN(U6181_n1) );
  NOR2X0 U6181_U1 ( .IN1(n3673), .IN2(U6181_n1), .QN(WX4715) );
  INVX0 U6182_U2 ( .INP(WX4650), .ZN(U6182_n1) );
  NOR2X0 U6182_U1 ( .IN1(n3672), .IN2(U6182_n1), .QN(WX4713) );
  INVX0 U6183_U2 ( .INP(WX4648), .ZN(U6183_n1) );
  NOR2X0 U6183_U1 ( .IN1(n3672), .IN2(U6183_n1), .QN(WX4711) );
  INVX0 U6184_U2 ( .INP(WX4646), .ZN(U6184_n1) );
  NOR2X0 U6184_U1 ( .IN1(n3672), .IN2(U6184_n1), .QN(WX4709) );
  INVX0 U6185_U2 ( .INP(WX4644), .ZN(U6185_n1) );
  NOR2X0 U6185_U1 ( .IN1(n3672), .IN2(U6185_n1), .QN(WX4707) );
  INVX0 U6186_U2 ( .INP(WX4642), .ZN(U6186_n1) );
  NOR2X0 U6186_U1 ( .IN1(n3672), .IN2(U6186_n1), .QN(WX4705) );
  INVX0 U6187_U2 ( .INP(WX4640), .ZN(U6187_n1) );
  NOR2X0 U6187_U1 ( .IN1(n3672), .IN2(U6187_n1), .QN(WX4703) );
  INVX0 U6188_U2 ( .INP(WX4638), .ZN(U6188_n1) );
  NOR2X0 U6188_U1 ( .IN1(n3672), .IN2(U6188_n1), .QN(WX4701) );
  INVX0 U6189_U2 ( .INP(WX4636), .ZN(U6189_n1) );
  NOR2X0 U6189_U1 ( .IN1(n3672), .IN2(U6189_n1), .QN(WX4699) );
  INVX0 U6190_U2 ( .INP(WX4634), .ZN(U6190_n1) );
  NOR2X0 U6190_U1 ( .IN1(n3672), .IN2(U6190_n1), .QN(WX4697) );
  INVX0 U6191_U2 ( .INP(WX4632), .ZN(U6191_n1) );
  NOR2X0 U6191_U1 ( .IN1(n3672), .IN2(U6191_n1), .QN(WX4695) );
  INVX0 U6192_U2 ( .INP(WX4630), .ZN(U6192_n1) );
  NOR2X0 U6192_U1 ( .IN1(n3672), .IN2(U6192_n1), .QN(WX4693) );
  INVX0 U6193_U2 ( .INP(WX4628), .ZN(U6193_n1) );
  NOR2X0 U6193_U1 ( .IN1(n3671), .IN2(U6193_n1), .QN(WX4691) );
  INVX0 U6194_U2 ( .INP(WX4626), .ZN(U6194_n1) );
  NOR2X0 U6194_U1 ( .IN1(n3671), .IN2(U6194_n1), .QN(WX4689) );
  INVX0 U6195_U2 ( .INP(WX4624), .ZN(U6195_n1) );
  NOR2X0 U6195_U1 ( .IN1(n3671), .IN2(U6195_n1), .QN(WX4687) );
  INVX0 U6196_U2 ( .INP(WX4622), .ZN(U6196_n1) );
  NOR2X0 U6196_U1 ( .IN1(n3671), .IN2(U6196_n1), .QN(WX4685) );
  INVX0 U6197_U2 ( .INP(test_so37), .ZN(U6197_n1) );
  NOR2X0 U6197_U1 ( .IN1(n3671), .IN2(U6197_n1), .QN(WX4683) );
  INVX0 U6198_U2 ( .INP(WX4618), .ZN(U6198_n1) );
  NOR2X0 U6198_U1 ( .IN1(n3671), .IN2(U6198_n1), .QN(WX4681) );
  INVX0 U6199_U2 ( .INP(WX4616), .ZN(U6199_n1) );
  NOR2X0 U6199_U1 ( .IN1(n3671), .IN2(U6199_n1), .QN(WX4679) );
  INVX0 U6200_U2 ( .INP(WX4614), .ZN(U6200_n1) );
  NOR2X0 U6200_U1 ( .IN1(n3671), .IN2(U6200_n1), .QN(WX4677) );
  INVX0 U6201_U2 ( .INP(WX4612), .ZN(U6201_n1) );
  NOR2X0 U6201_U1 ( .IN1(n3671), .IN2(U6201_n1), .QN(WX4675) );
  INVX0 U6202_U2 ( .INP(WX4610), .ZN(U6202_n1) );
  NOR2X0 U6202_U1 ( .IN1(n3671), .IN2(U6202_n1), .QN(WX4673) );
  INVX0 U6203_U2 ( .INP(WX4608), .ZN(U6203_n1) );
  NOR2X0 U6203_U1 ( .IN1(n3671), .IN2(U6203_n1), .QN(WX4671) );
  INVX0 U6204_U2 ( .INP(WX4606), .ZN(U6204_n1) );
  NOR2X0 U6204_U1 ( .IN1(n3670), .IN2(U6204_n1), .QN(WX4669) );
  INVX0 U6205_U2 ( .INP(WX4604), .ZN(U6205_n1) );
  NOR2X0 U6205_U1 ( .IN1(n3670), .IN2(U6205_n1), .QN(WX4667) );
  INVX0 U6206_U2 ( .INP(WX4602), .ZN(U6206_n1) );
  NOR2X0 U6206_U1 ( .IN1(n3670), .IN2(U6206_n1), .QN(WX4665) );
  INVX0 U6207_U2 ( .INP(WX4600), .ZN(U6207_n1) );
  NOR2X0 U6207_U1 ( .IN1(n3670), .IN2(U6207_n1), .QN(WX4663) );
  INVX0 U6208_U2 ( .INP(WX4598), .ZN(U6208_n1) );
  NOR2X0 U6208_U1 ( .IN1(n3670), .IN2(U6208_n1), .QN(WX4661) );
  INVX0 U6209_U2 ( .INP(WX4596), .ZN(U6209_n1) );
  NOR2X0 U6209_U1 ( .IN1(n3670), .IN2(U6209_n1), .QN(WX4659) );
  INVX0 U6210_U2 ( .INP(WX4594), .ZN(U6210_n1) );
  NOR2X0 U6210_U1 ( .IN1(n3670), .IN2(U6210_n1), .QN(WX4657) );
  INVX0 U6211_U2 ( .INP(WX4592), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n3670), .IN2(U6211_n1), .QN(WX4655) );
  INVX0 U6212_U2 ( .INP(WX4590), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n3670), .IN2(U6212_n1), .QN(WX4653) );
  INVX0 U6213_U2 ( .INP(WX4588), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n3670), .IN2(U6213_n1), .QN(WX4651) );
  INVX0 U6214_U2 ( .INP(test_so36), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n3670), .IN2(U6214_n1), .QN(WX4649) );
  INVX0 U6215_U2 ( .INP(WX4584), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n3668), .IN2(U6215_n1), .QN(WX4647) );
  INVX0 U6216_U2 ( .INP(WX4582), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n3668), .IN2(U6216_n1), .QN(WX4645) );
  INVX0 U6217_U2 ( .INP(WX4580), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n3668), .IN2(U6217_n1), .QN(WX4643) );
  INVX0 U6218_U2 ( .INP(WX4578), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n3668), .IN2(U6218_n1), .QN(WX4641) );
  INVX0 U6219_U2 ( .INP(WX4576), .ZN(U6219_n1) );
  NOR2X0 U6219_U1 ( .IN1(n3668), .IN2(U6219_n1), .QN(WX4639) );
  INVX0 U6220_U2 ( .INP(WX4574), .ZN(U6220_n1) );
  NOR2X0 U6220_U1 ( .IN1(n3668), .IN2(U6220_n1), .QN(WX4637) );
  INVX0 U6221_U2 ( .INP(WX4572), .ZN(U6221_n1) );
  NOR2X0 U6221_U1 ( .IN1(n3668), .IN2(U6221_n1), .QN(WX4635) );
  INVX0 U6222_U2 ( .INP(WX4570), .ZN(U6222_n1) );
  NOR2X0 U6222_U1 ( .IN1(n3668), .IN2(U6222_n1), .QN(WX4633) );
  INVX0 U6223_U2 ( .INP(WX4568), .ZN(U6223_n1) );
  NOR2X0 U6223_U1 ( .IN1(n3668), .IN2(U6223_n1), .QN(WX4631) );
  INVX0 U6224_U2 ( .INP(WX4566), .ZN(U6224_n1) );
  NOR2X0 U6224_U1 ( .IN1(n3668), .IN2(U6224_n1), .QN(WX4629) );
  INVX0 U6225_U2 ( .INP(WX4564), .ZN(U6225_n1) );
  NOR2X0 U6225_U1 ( .IN1(n3668), .IN2(U6225_n1), .QN(WX4627) );
  INVX0 U6226_U2 ( .INP(WX4562), .ZN(U6226_n1) );
  NOR2X0 U6226_U1 ( .IN1(n3667), .IN2(U6226_n1), .QN(WX4625) );
  INVX0 U6227_U2 ( .INP(WX4560), .ZN(U6227_n1) );
  NOR2X0 U6227_U1 ( .IN1(n3667), .IN2(U6227_n1), .QN(WX4623) );
  INVX0 U6228_U2 ( .INP(WX4558), .ZN(U6228_n1) );
  NOR2X0 U6228_U1 ( .IN1(n3667), .IN2(U6228_n1), .QN(WX4621) );
  INVX0 U6229_U2 ( .INP(WX4556), .ZN(U6229_n1) );
  NOR2X0 U6229_U1 ( .IN1(n3667), .IN2(U6229_n1), .QN(WX4619) );
  INVX0 U6230_U2 ( .INP(WX3421), .ZN(U6230_n1) );
  NOR2X0 U6230_U1 ( .IN1(n3667), .IN2(U6230_n1), .QN(WX3484) );
  INVX0 U6231_U2 ( .INP(WX3419), .ZN(U6231_n1) );
  NOR2X0 U6231_U1 ( .IN1(n3667), .IN2(U6231_n1), .QN(WX3482) );
  INVX0 U6232_U2 ( .INP(WX3417), .ZN(U6232_n1) );
  NOR2X0 U6232_U1 ( .IN1(n3667), .IN2(U6232_n1), .QN(WX3480) );
  INVX0 U6233_U2 ( .INP(WX3415), .ZN(U6233_n1) );
  NOR2X0 U6233_U1 ( .IN1(n3667), .IN2(U6233_n1), .QN(WX3478) );
  INVX0 U6234_U2 ( .INP(WX3413), .ZN(U6234_n1) );
  NOR2X0 U6234_U1 ( .IN1(n3667), .IN2(U6234_n1), .QN(WX3476) );
  INVX0 U6235_U2 ( .INP(WX3411), .ZN(U6235_n1) );
  NOR2X0 U6235_U1 ( .IN1(n3667), .IN2(U6235_n1), .QN(WX3474) );
  INVX0 U6236_U2 ( .INP(WX3409), .ZN(U6236_n1) );
  NOR2X0 U6236_U1 ( .IN1(n3667), .IN2(U6236_n1), .QN(WX3472) );
  INVX0 U6237_U2 ( .INP(WX3407), .ZN(U6237_n1) );
  NOR2X0 U6237_U1 ( .IN1(n3666), .IN2(U6237_n1), .QN(WX3470) );
  INVX0 U6238_U2 ( .INP(test_so28), .ZN(U6238_n1) );
  NOR2X0 U6238_U1 ( .IN1(n3666), .IN2(U6238_n1), .QN(WX3468) );
  INVX0 U6239_U2 ( .INP(WX3403), .ZN(U6239_n1) );
  NOR2X0 U6239_U1 ( .IN1(n3666), .IN2(U6239_n1), .QN(WX3466) );
  INVX0 U6240_U2 ( .INP(WX3401), .ZN(U6240_n1) );
  NOR2X0 U6240_U1 ( .IN1(n3666), .IN2(U6240_n1), .QN(WX3464) );
  INVX0 U6241_U2 ( .INP(WX3399), .ZN(U6241_n1) );
  NOR2X0 U6241_U1 ( .IN1(n3666), .IN2(U6241_n1), .QN(WX3462) );
  INVX0 U6242_U2 ( .INP(WX3397), .ZN(U6242_n1) );
  NOR2X0 U6242_U1 ( .IN1(n3702), .IN2(U6242_n1), .QN(WX3460) );
  INVX0 U6243_U2 ( .INP(WX3395), .ZN(U6243_n1) );
  NOR2X0 U6243_U1 ( .IN1(n3731), .IN2(U6243_n1), .QN(WX3458) );
  INVX0 U6244_U2 ( .INP(WX3393), .ZN(U6244_n1) );
  NOR2X0 U6244_U1 ( .IN1(n3732), .IN2(U6244_n1), .QN(WX3456) );
  INVX0 U6245_U2 ( .INP(WX3391), .ZN(U6245_n1) );
  NOR2X0 U6245_U1 ( .IN1(n3723), .IN2(U6245_n1), .QN(WX3454) );
  INVX0 U6246_U2 ( .INP(WX3389), .ZN(U6246_n1) );
  NOR2X0 U6246_U1 ( .IN1(n3724), .IN2(U6246_n1), .QN(WX3452) );
  INVX0 U6247_U2 ( .INP(WX3387), .ZN(U6247_n1) );
  NOR2X0 U6247_U1 ( .IN1(n3725), .IN2(U6247_n1), .QN(WX3450) );
  INVX0 U6248_U2 ( .INP(WX3385), .ZN(U6248_n1) );
  NOR2X0 U6248_U1 ( .IN1(n3726), .IN2(U6248_n1), .QN(WX3448) );
  INVX0 U6249_U2 ( .INP(WX3383), .ZN(U6249_n1) );
  NOR2X0 U6249_U1 ( .IN1(n3727), .IN2(U6249_n1), .QN(WX3446) );
  INVX0 U6250_U2 ( .INP(WX3381), .ZN(U6250_n1) );
  NOR2X0 U6250_U1 ( .IN1(n3728), .IN2(U6250_n1), .QN(WX3444) );
  INVX0 U6251_U2 ( .INP(WX3379), .ZN(U6251_n1) );
  NOR2X0 U6251_U1 ( .IN1(n3687), .IN2(U6251_n1), .QN(WX3442) );
  INVX0 U6252_U2 ( .INP(WX3377), .ZN(U6252_n1) );
  NOR2X0 U6252_U1 ( .IN1(n3688), .IN2(U6252_n1), .QN(WX3440) );
  INVX0 U6253_U2 ( .INP(WX3375), .ZN(U6253_n1) );
  NOR2X0 U6253_U1 ( .IN1(n3673), .IN2(U6253_n1), .QN(WX3438) );
  INVX0 U6254_U2 ( .INP(WX3373), .ZN(U6254_n1) );
  NOR2X0 U6254_U1 ( .IN1(n3674), .IN2(U6254_n1), .QN(WX3436) );
  INVX0 U6255_U2 ( .INP(WX3371), .ZN(U6255_n1) );
  NOR2X0 U6255_U1 ( .IN1(n3675), .IN2(U6255_n1), .QN(WX3434) );
  INVX0 U6256_U2 ( .INP(test_so27), .ZN(U6256_n1) );
  NOR2X0 U6256_U1 ( .IN1(n3676), .IN2(U6256_n1), .QN(WX3432) );
  INVX0 U6257_U2 ( .INP(WX3367), .ZN(U6257_n1) );
  NOR2X0 U6257_U1 ( .IN1(n3677), .IN2(U6257_n1), .QN(WX3430) );
  INVX0 U6258_U2 ( .INP(WX3365), .ZN(U6258_n1) );
  NOR2X0 U6258_U1 ( .IN1(n3678), .IN2(U6258_n1), .QN(WX3428) );
  INVX0 U6259_U2 ( .INP(WX3363), .ZN(U6259_n1) );
  NOR2X0 U6259_U1 ( .IN1(n3679), .IN2(U6259_n1), .QN(WX3426) );
  INVX0 U6260_U2 ( .INP(WX3361), .ZN(U6260_n1) );
  NOR2X0 U6260_U1 ( .IN1(n3680), .IN2(U6260_n1), .QN(WX3424) );
  INVX0 U6261_U2 ( .INP(WX3359), .ZN(U6261_n1) );
  NOR2X0 U6261_U1 ( .IN1(n3714), .IN2(U6261_n1), .QN(WX3422) );
  INVX0 U6262_U2 ( .INP(WX3357), .ZN(U6262_n1) );
  NOR2X0 U6262_U1 ( .IN1(n3715), .IN2(U6262_n1), .QN(WX3420) );
  INVX0 U6263_U2 ( .INP(WX3355), .ZN(U6263_n1) );
  NOR2X0 U6263_U1 ( .IN1(n3716), .IN2(U6263_n1), .QN(WX3418) );
  INVX0 U6264_U2 ( .INP(WX3353), .ZN(U6264_n1) );
  NOR2X0 U6264_U1 ( .IN1(n3718), .IN2(U6264_n1), .QN(WX3416) );
  INVX0 U6265_U2 ( .INP(WX3351), .ZN(U6265_n1) );
  NOR2X0 U6265_U1 ( .IN1(n3719), .IN2(U6265_n1), .QN(WX3414) );
  INVX0 U6266_U2 ( .INP(WX3349), .ZN(U6266_n1) );
  NOR2X0 U6266_U1 ( .IN1(n3720), .IN2(U6266_n1), .QN(WX3412) );
  INVX0 U6267_U2 ( .INP(WX3347), .ZN(U6267_n1) );
  NOR2X0 U6267_U1 ( .IN1(n3721), .IN2(U6267_n1), .QN(WX3410) );
  INVX0 U6268_U2 ( .INP(WX3345), .ZN(U6268_n1) );
  NOR2X0 U6268_U1 ( .IN1(n3722), .IN2(U6268_n1), .QN(WX3408) );
  INVX0 U6269_U2 ( .INP(WX3343), .ZN(U6269_n1) );
  NOR2X0 U6269_U1 ( .IN1(n3705), .IN2(U6269_n1), .QN(WX3406) );
  INVX0 U6270_U2 ( .INP(WX3341), .ZN(U6270_n1) );
  NOR2X0 U6270_U1 ( .IN1(n3706), .IN2(U6270_n1), .QN(WX3404) );
  INVX0 U6271_U2 ( .INP(WX3339), .ZN(U6271_n1) );
  NOR2X0 U6271_U1 ( .IN1(n3707), .IN2(U6271_n1), .QN(WX3402) );
  INVX0 U6272_U2 ( .INP(WX3337), .ZN(U6272_n1) );
  NOR2X0 U6272_U1 ( .IN1(n3708), .IN2(U6272_n1), .QN(WX3400) );
  INVX0 U6273_U2 ( .INP(WX3335), .ZN(U6273_n1) );
  NOR2X0 U6273_U1 ( .IN1(n3709), .IN2(U6273_n1), .QN(WX3398) );
  INVX0 U6274_U2 ( .INP(test_so26), .ZN(U6274_n1) );
  NOR2X0 U6274_U1 ( .IN1(n3710), .IN2(U6274_n1), .QN(WX3396) );
  INVX0 U6275_U2 ( .INP(WX3331), .ZN(U6275_n1) );
  NOR2X0 U6275_U1 ( .IN1(n3711), .IN2(U6275_n1), .QN(WX3394) );
  INVX0 U6276_U2 ( .INP(WX3329), .ZN(U6276_n1) );
  NOR2X0 U6276_U1 ( .IN1(n3712), .IN2(U6276_n1), .QN(WX3392) );
  INVX0 U6277_U2 ( .INP(WX3327), .ZN(U6277_n1) );
  NOR2X0 U6277_U1 ( .IN1(n3698), .IN2(U6277_n1), .QN(WX3390) );
  INVX0 U6278_U2 ( .INP(WX3325), .ZN(U6278_n1) );
  NOR2X0 U6278_U1 ( .IN1(n3699), .IN2(U6278_n1), .QN(WX3388) );
  INVX0 U6279_U2 ( .INP(WX3323), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n3700), .IN2(U6279_n1), .QN(WX3386) );
  INVX0 U6280_U2 ( .INP(WX3321), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n3666), .IN2(U6280_n1), .QN(WX3384) );
  INVX0 U6281_U2 ( .INP(WX3319), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n3701), .IN2(U6281_n1), .QN(WX3382) );
  INVX0 U6282_U2 ( .INP(WX3317), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n3703), .IN2(U6282_n1), .QN(WX3380) );
  INVX0 U6283_U2 ( .INP(WX3315), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n3663), .IN2(U6283_n1), .QN(WX3378) );
  INVX0 U6284_U2 ( .INP(WX3313), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n3663), .IN2(U6284_n1), .QN(WX3376) );
  INVX0 U6285_U2 ( .INP(WX3311), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n3663), .IN2(U6285_n1), .QN(WX3374) );
  INVX0 U6286_U2 ( .INP(WX3309), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n3663), .IN2(U6286_n1), .QN(WX3372) );
  INVX0 U6287_U2 ( .INP(WX3307), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n3663), .IN2(U6287_n1), .QN(WX3370) );
  INVX0 U6288_U2 ( .INP(WX3305), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n3663), .IN2(U6288_n1), .QN(WX3368) );
  INVX0 U6289_U2 ( .INP(WX3303), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n3663), .IN2(U6289_n1), .QN(WX3366) );
  INVX0 U6290_U2 ( .INP(WX3301), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n3663), .IN2(U6290_n1), .QN(WX3364) );
  INVX0 U6291_U2 ( .INP(WX3299), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n3663), .IN2(U6291_n1), .QN(WX3362) );
  INVX0 U6292_U2 ( .INP(test_so25), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n3663), .IN2(U6292_n1), .QN(WX3360) );
  INVX0 U6293_U2 ( .INP(WX3295), .ZN(U6293_n1) );
  NOR2X0 U6293_U1 ( .IN1(n3663), .IN2(U6293_n1), .QN(WX3358) );
  INVX0 U6294_U2 ( .INP(WX3293), .ZN(U6294_n1) );
  NOR2X0 U6294_U1 ( .IN1(n3664), .IN2(U6294_n1), .QN(WX3356) );
  INVX0 U6295_U2 ( .INP(WX3291), .ZN(U6295_n1) );
  NOR2X0 U6295_U1 ( .IN1(n3664), .IN2(U6295_n1), .QN(WX3354) );
  INVX0 U6296_U2 ( .INP(WX3289), .ZN(U6296_n1) );
  NOR2X0 U6296_U1 ( .IN1(n3664), .IN2(U6296_n1), .QN(WX3352) );
  INVX0 U6297_U2 ( .INP(WX3287), .ZN(U6297_n1) );
  NOR2X0 U6297_U1 ( .IN1(n3664), .IN2(U6297_n1), .QN(WX3350) );
  INVX0 U6298_U2 ( .INP(WX3285), .ZN(U6298_n1) );
  NOR2X0 U6298_U1 ( .IN1(n3664), .IN2(U6298_n1), .QN(WX3348) );
  INVX0 U6299_U2 ( .INP(WX3283), .ZN(U6299_n1) );
  NOR2X0 U6299_U1 ( .IN1(n3664), .IN2(U6299_n1), .QN(WX3346) );
  INVX0 U6300_U2 ( .INP(WX3281), .ZN(U6300_n1) );
  NOR2X0 U6300_U1 ( .IN1(n3664), .IN2(U6300_n1), .QN(WX3344) );
  INVX0 U6301_U2 ( .INP(WX3279), .ZN(U6301_n1) );
  NOR2X0 U6301_U1 ( .IN1(n3664), .IN2(U6301_n1), .QN(WX3342) );
  INVX0 U6302_U2 ( .INP(WX3277), .ZN(U6302_n1) );
  NOR2X0 U6302_U1 ( .IN1(n3664), .IN2(U6302_n1), .QN(WX3340) );
  INVX0 U6303_U2 ( .INP(WX3275), .ZN(U6303_n1) );
  NOR2X0 U6303_U1 ( .IN1(n3664), .IN2(U6303_n1), .QN(WX3338) );
  INVX0 U6304_U2 ( .INP(WX3273), .ZN(U6304_n1) );
  NOR2X0 U6304_U1 ( .IN1(n3664), .IN2(U6304_n1), .QN(WX3336) );
  INVX0 U6305_U2 ( .INP(WX3271), .ZN(U6305_n1) );
  NOR2X0 U6305_U1 ( .IN1(n3665), .IN2(U6305_n1), .QN(WX3334) );
  INVX0 U6306_U2 ( .INP(WX3267), .ZN(U6306_n1) );
  NOR2X0 U6306_U1 ( .IN1(n3665), .IN2(U6306_n1), .QN(WX3330) );
  INVX0 U6307_U2 ( .INP(WX2128), .ZN(U6307_n1) );
  NOR2X0 U6307_U1 ( .IN1(n3665), .IN2(U6307_n1), .QN(WX2191) );
  INVX0 U6308_U2 ( .INP(WX2126), .ZN(U6308_n1) );
  NOR2X0 U6308_U1 ( .IN1(n3665), .IN2(U6308_n1), .QN(WX2189) );
  INVX0 U6309_U2 ( .INP(WX2124), .ZN(U6309_n1) );
  NOR2X0 U6309_U1 ( .IN1(n3665), .IN2(U6309_n1), .QN(WX2187) );
  INVX0 U6310_U2 ( .INP(WX2122), .ZN(U6310_n1) );
  NOR2X0 U6310_U1 ( .IN1(n3665), .IN2(U6310_n1), .QN(WX2185) );
  INVX0 U6311_U2 ( .INP(WX2120), .ZN(U6311_n1) );
  NOR2X0 U6311_U1 ( .IN1(n3665), .IN2(U6311_n1), .QN(WX2183) );
  INVX0 U6312_U2 ( .INP(WX2118), .ZN(U6312_n1) );
  NOR2X0 U6312_U1 ( .IN1(n3665), .IN2(U6312_n1), .QN(WX2181) );
  INVX0 U6313_U2 ( .INP(WX2116), .ZN(U6313_n1) );
  NOR2X0 U6313_U1 ( .IN1(n3665), .IN2(U6313_n1), .QN(WX2179) );
  INVX0 U6314_U2 ( .INP(WX2114), .ZN(U6314_n1) );
  NOR2X0 U6314_U1 ( .IN1(n3665), .IN2(U6314_n1), .QN(WX2177) );
  INVX0 U6315_U2 ( .INP(WX2112), .ZN(U6315_n1) );
  NOR2X0 U6315_U1 ( .IN1(n3665), .IN2(U6315_n1), .QN(WX2175) );
  INVX0 U6316_U2 ( .INP(WX2110), .ZN(U6316_n1) );
  NOR2X0 U6316_U1 ( .IN1(n3666), .IN2(U6316_n1), .QN(WX2173) );
  INVX0 U6317_U2 ( .INP(WX2108), .ZN(U6317_n1) );
  NOR2X0 U6317_U1 ( .IN1(n3666), .IN2(U6317_n1), .QN(WX2171) );
  INVX0 U6318_U2 ( .INP(WX2106), .ZN(U6318_n1) );
  NOR2X0 U6318_U1 ( .IN1(n3666), .IN2(U6318_n1), .QN(WX2169) );
  INVX0 U6319_U2 ( .INP(WX2104), .ZN(U6319_n1) );
  NOR2X0 U6319_U1 ( .IN1(n3666), .IN2(U6319_n1), .QN(WX2167) );
  INVX0 U6320_U2 ( .INP(WX2102), .ZN(U6320_n1) );
  NOR2X0 U6320_U1 ( .IN1(n3666), .IN2(U6320_n1), .QN(WX2165) );
  INVX0 U6321_U2 ( .INP(test_so17), .ZN(U6321_n1) );
  NOR2X0 U6321_U1 ( .IN1(n3666), .IN2(U6321_n1), .QN(WX2163) );
  INVX0 U6322_U2 ( .INP(WX2098), .ZN(U6322_n1) );
  NOR2X0 U6322_U1 ( .IN1(n3689), .IN2(U6322_n1), .QN(WX2161) );
  INVX0 U6323_U2 ( .INP(WX2096), .ZN(U6323_n1) );
  NOR2X0 U6323_U1 ( .IN1(n3689), .IN2(U6323_n1), .QN(WX2159) );
  INVX0 U6324_U2 ( .INP(WX2094), .ZN(U6324_n1) );
  NOR2X0 U6324_U1 ( .IN1(n3689), .IN2(U6324_n1), .QN(WX2157) );
  INVX0 U6325_U2 ( .INP(WX2092), .ZN(U6325_n1) );
  NOR2X0 U6325_U1 ( .IN1(n3689), .IN2(U6325_n1), .QN(WX2155) );
  INVX0 U6326_U2 ( .INP(WX2090), .ZN(U6326_n1) );
  NOR2X0 U6326_U1 ( .IN1(n3689), .IN2(U6326_n1), .QN(WX2153) );
  INVX0 U6327_U2 ( .INP(WX2088), .ZN(U6327_n1) );
  NOR2X0 U6327_U1 ( .IN1(n3689), .IN2(U6327_n1), .QN(WX2151) );
  INVX0 U6328_U2 ( .INP(WX2086), .ZN(U6328_n1) );
  NOR2X0 U6328_U1 ( .IN1(n3688), .IN2(U6328_n1), .QN(WX2149) );
  INVX0 U6329_U2 ( .INP(WX2084), .ZN(U6329_n1) );
  NOR2X0 U6329_U1 ( .IN1(n3688), .IN2(U6329_n1), .QN(WX2147) );
  INVX0 U6330_U2 ( .INP(WX2082), .ZN(U6330_n1) );
  NOR2X0 U6330_U1 ( .IN1(n3688), .IN2(U6330_n1), .QN(WX2145) );
  INVX0 U6331_U2 ( .INP(WX2080), .ZN(U6331_n1) );
  NOR2X0 U6331_U1 ( .IN1(n3688), .IN2(U6331_n1), .QN(WX2143) );
  INVX0 U6332_U2 ( .INP(WX2078), .ZN(U6332_n1) );
  NOR2X0 U6332_U1 ( .IN1(n3688), .IN2(U6332_n1), .QN(WX2141) );
  INVX0 U6333_U2 ( .INP(WX2076), .ZN(U6333_n1) );
  NOR2X0 U6333_U1 ( .IN1(n3688), .IN2(U6333_n1), .QN(WX2139) );
  INVX0 U6334_U2 ( .INP(WX2074), .ZN(U6334_n1) );
  NOR2X0 U6334_U1 ( .IN1(n3688), .IN2(U6334_n1), .QN(WX2137) );
  INVX0 U6335_U2 ( .INP(WX2072), .ZN(U6335_n1) );
  NOR2X0 U6335_U1 ( .IN1(n3688), .IN2(U6335_n1), .QN(WX2135) );
  INVX0 U6336_U2 ( .INP(WX2070), .ZN(U6336_n1) );
  NOR2X0 U6336_U1 ( .IN1(n3688), .IN2(U6336_n1), .QN(WX2133) );
  INVX0 U6337_U2 ( .INP(WX2068), .ZN(U6337_n1) );
  NOR2X0 U6337_U1 ( .IN1(n3688), .IN2(U6337_n1), .QN(WX2131) );
  INVX0 U6338_U2 ( .INP(WX2066), .ZN(U6338_n1) );
  NOR2X0 U6338_U1 ( .IN1(n3688), .IN2(U6338_n1), .QN(WX2129) );
  INVX0 U6339_U2 ( .INP(test_so16), .ZN(U6339_n1) );
  NOR2X0 U6339_U1 ( .IN1(n3687), .IN2(U6339_n1), .QN(WX2127) );
  INVX0 U6340_U2 ( .INP(WX2062), .ZN(U6340_n1) );
  NOR2X0 U6340_U1 ( .IN1(n3687), .IN2(U6340_n1), .QN(WX2125) );
  INVX0 U6341_U2 ( .INP(WX2060), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n3687), .IN2(U6341_n1), .QN(WX2123) );
  INVX0 U6342_U2 ( .INP(WX2058), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n3687), .IN2(U6342_n1), .QN(WX2121) );
  INVX0 U6343_U2 ( .INP(WX2056), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n3687), .IN2(U6343_n1), .QN(WX2119) );
  INVX0 U6344_U2 ( .INP(WX2054), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n3687), .IN2(U6344_n1), .QN(WX2117) );
  INVX0 U6345_U2 ( .INP(WX2052), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n3687), .IN2(U6345_n1), .QN(WX2115) );
  INVX0 U6346_U2 ( .INP(WX2050), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n3687), .IN2(U6346_n1), .QN(WX2113) );
  INVX0 U6347_U2 ( .INP(WX2048), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n3687), .IN2(U6347_n1), .QN(WX2111) );
  INVX0 U6348_U2 ( .INP(WX2046), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n3687), .IN2(U6348_n1), .QN(WX2109) );
  INVX0 U6349_U2 ( .INP(WX2044), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n3687), .IN2(U6349_n1), .QN(WX2107) );
  INVX0 U6350_U2 ( .INP(WX2042), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n3686), .IN2(U6350_n1), .QN(WX2105) );
  INVX0 U6351_U2 ( .INP(WX2040), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n3686), .IN2(U6351_n1), .QN(WX2103) );
  INVX0 U6352_U2 ( .INP(WX2038), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n3686), .IN2(U6352_n1), .QN(WX2101) );
  INVX0 U6353_U2 ( .INP(WX2036), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n3686), .IN2(U6353_n1), .QN(WX2099) );
  INVX0 U6354_U2 ( .INP(WX2034), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n3686), .IN2(U6354_n1), .QN(WX2097) );
  INVX0 U6355_U2 ( .INP(WX2032), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n3686), .IN2(U6355_n1), .QN(WX2095) );
  INVX0 U6356_U2 ( .INP(WX2030), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n3686), .IN2(U6356_n1), .QN(WX2093) );
  INVX0 U6357_U2 ( .INP(test_so15), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n3686), .IN2(U6357_n1), .QN(WX2091) );
  INVX0 U6358_U2 ( .INP(WX2026), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n3686), .IN2(U6358_n1), .QN(WX2089) );
  INVX0 U6359_U2 ( .INP(WX2024), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n3686), .IN2(U6359_n1), .QN(WX2087) );
  INVX0 U6360_U2 ( .INP(WX2022), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n3686), .IN2(U6360_n1), .QN(WX2085) );
  INVX0 U6361_U2 ( .INP(WX2020), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n3685), .IN2(U6361_n1), .QN(WX2083) );
  INVX0 U6362_U2 ( .INP(WX2018), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n3685), .IN2(U6362_n1), .QN(WX2081) );
  INVX0 U6363_U2 ( .INP(WX2016), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n3685), .IN2(U6363_n1), .QN(WX2079) );
  INVX0 U6364_U2 ( .INP(WX2014), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n3685), .IN2(U6364_n1), .QN(WX2077) );
  INVX0 U6365_U2 ( .INP(WX2012), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n3685), .IN2(U6365_n1), .QN(WX2075) );
  INVX0 U6366_U2 ( .INP(WX2010), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n3685), .IN2(U6366_n1), .QN(WX2073) );
  INVX0 U6367_U2 ( .INP(WX2008), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n3685), .IN2(U6367_n1), .QN(WX2071) );
  INVX0 U6368_U2 ( .INP(WX2006), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n3685), .IN2(U6368_n1), .QN(WX2069) );
  INVX0 U6369_U2 ( .INP(WX2004), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n3685), .IN2(U6369_n1), .QN(WX2067) );
  INVX0 U6370_U2 ( .INP(WX2002), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n3685), .IN2(U6370_n1), .QN(WX2065) );
  INVX0 U6371_U2 ( .INP(WX2000), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n3685), .IN2(U6371_n1), .QN(WX2063) );
  INVX0 U6372_U2 ( .INP(WX1998), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n3684), .IN2(U6372_n1), .QN(WX2061) );
  INVX0 U6373_U2 ( .INP(WX1996), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n3684), .IN2(U6373_n1), .QN(WX2059) );
  INVX0 U6374_U2 ( .INP(WX1994), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n3684), .IN2(U6374_n1), .QN(WX2057) );
  INVX0 U6375_U2 ( .INP(test_so14), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n3684), .IN2(U6375_n1), .QN(WX2055) );
  INVX0 U6376_U2 ( .INP(WX1990), .ZN(U6376_n1) );
  NOR2X0 U6376_U1 ( .IN1(n3684), .IN2(U6376_n1), .QN(WX2053) );
  INVX0 U6377_U2 ( .INP(WX1988), .ZN(U6377_n1) );
  NOR2X0 U6377_U1 ( .IN1(n3684), .IN2(U6377_n1), .QN(WX2051) );
  INVX0 U6378_U2 ( .INP(WX1986), .ZN(U6378_n1) );
  NOR2X0 U6378_U1 ( .IN1(n3684), .IN2(U6378_n1), .QN(WX2049) );
  INVX0 U6379_U2 ( .INP(WX1984), .ZN(U6379_n1) );
  NOR2X0 U6379_U1 ( .IN1(n3684), .IN2(U6379_n1), .QN(WX2047) );
  INVX0 U6380_U2 ( .INP(WX1982), .ZN(U6380_n1) );
  NOR2X0 U6380_U1 ( .IN1(n3684), .IN2(U6380_n1), .QN(WX2045) );
  INVX0 U6381_U2 ( .INP(WX1980), .ZN(U6381_n1) );
  NOR2X0 U6381_U1 ( .IN1(n3684), .IN2(U6381_n1), .QN(WX2043) );
  INVX0 U6382_U2 ( .INP(WX1978), .ZN(U6382_n1) );
  NOR2X0 U6382_U1 ( .IN1(n3684), .IN2(U6382_n1), .QN(WX2041) );
  INVX0 U6383_U2 ( .INP(WX1976), .ZN(U6383_n1) );
  NOR2X0 U6383_U1 ( .IN1(n3683), .IN2(U6383_n1), .QN(WX2039) );
  INVX0 U6384_U2 ( .INP(WX1974), .ZN(U6384_n1) );
  NOR2X0 U6384_U1 ( .IN1(n3683), .IN2(U6384_n1), .QN(WX2037) );
  INVX0 U6385_U2 ( .INP(WX1972), .ZN(U6385_n1) );
  NOR2X0 U6385_U1 ( .IN1(n3683), .IN2(U6385_n1), .QN(WX2035) );
  INVX0 U6386_U2 ( .INP(WX1970), .ZN(U6386_n1) );
  NOR2X0 U6386_U1 ( .IN1(n3683), .IN2(U6386_n1), .QN(WX2033) );
  INVX0 U6387_U2 ( .INP(WX835), .ZN(U6387_n1) );
  NOR2X0 U6387_U1 ( .IN1(n3683), .IN2(U6387_n1), .QN(WX898) );
  INVX0 U6388_U2 ( .INP(WX833), .ZN(U6388_n1) );
  NOR2X0 U6388_U1 ( .IN1(n3683), .IN2(U6388_n1), .QN(WX896) );
  INVX0 U6389_U2 ( .INP(test_so7), .ZN(U6389_n1) );
  NOR2X0 U6389_U1 ( .IN1(n3683), .IN2(U6389_n1), .QN(WX894) );
  INVX0 U6390_U2 ( .INP(WX829), .ZN(U6390_n1) );
  NOR2X0 U6390_U1 ( .IN1(n3683), .IN2(U6390_n1), .QN(WX892) );
  INVX0 U6391_U2 ( .INP(WX827), .ZN(U6391_n1) );
  NOR2X0 U6391_U1 ( .IN1(n3683), .IN2(U6391_n1), .QN(WX890) );
  INVX0 U6392_U2 ( .INP(WX825), .ZN(U6392_n1) );
  NOR2X0 U6392_U1 ( .IN1(n3683), .IN2(U6392_n1), .QN(WX888) );
  INVX0 U6393_U2 ( .INP(WX823), .ZN(U6393_n1) );
  NOR2X0 U6393_U1 ( .IN1(n3683), .IN2(U6393_n1), .QN(WX886) );
  INVX0 U6394_U2 ( .INP(WX821), .ZN(U6394_n1) );
  NOR2X0 U6394_U1 ( .IN1(n3682), .IN2(U6394_n1), .QN(WX884) );
  INVX0 U6395_U2 ( .INP(WX819), .ZN(U6395_n1) );
  NOR2X0 U6395_U1 ( .IN1(n3682), .IN2(U6395_n1), .QN(WX882) );
  INVX0 U6396_U2 ( .INP(WX817), .ZN(U6396_n1) );
  NOR2X0 U6396_U1 ( .IN1(n3682), .IN2(U6396_n1), .QN(WX880) );
  INVX0 U6397_U2 ( .INP(WX815), .ZN(U6397_n1) );
  NOR2X0 U6397_U1 ( .IN1(n3682), .IN2(U6397_n1), .QN(WX878) );
  INVX0 U6398_U2 ( .INP(WX813), .ZN(U6398_n1) );
  NOR2X0 U6398_U1 ( .IN1(n3682), .IN2(U6398_n1), .QN(WX876) );
  INVX0 U6399_U2 ( .INP(WX811), .ZN(U6399_n1) );
  NOR2X0 U6399_U1 ( .IN1(n3682), .IN2(U6399_n1), .QN(WX874) );
  INVX0 U6400_U2 ( .INP(WX809), .ZN(U6400_n1) );
  NOR2X0 U6400_U1 ( .IN1(n3682), .IN2(U6400_n1), .QN(WX872) );
  INVX0 U6401_U2 ( .INP(WX807), .ZN(U6401_n1) );
  NOR2X0 U6401_U1 ( .IN1(n3682), .IN2(U6401_n1), .QN(WX870) );
  INVX0 U6402_U2 ( .INP(WX805), .ZN(U6402_n1) );
  NOR2X0 U6402_U1 ( .IN1(n3682), .IN2(U6402_n1), .QN(WX868) );
  INVX0 U6403_U2 ( .INP(WX803), .ZN(U6403_n1) );
  NOR2X0 U6403_U1 ( .IN1(n3682), .IN2(U6403_n1), .QN(WX866) );
  INVX0 U6404_U2 ( .INP(WX801), .ZN(U6404_n1) );
  NOR2X0 U6404_U1 ( .IN1(n3681), .IN2(U6404_n1), .QN(WX864) );
  INVX0 U6405_U2 ( .INP(WX799), .ZN(U6405_n1) );
  NOR2X0 U6405_U1 ( .IN1(n3681), .IN2(U6405_n1), .QN(WX862) );
  INVX0 U6406_U2 ( .INP(WX797), .ZN(U6406_n1) );
  NOR2X0 U6406_U1 ( .IN1(n3681), .IN2(U6406_n1), .QN(WX860) );
  INVX0 U6407_U2 ( .INP(test_so6), .ZN(U6407_n1) );
  NOR2X0 U6407_U1 ( .IN1(n3681), .IN2(U6407_n1), .QN(WX858) );
  INVX0 U6408_U2 ( .INP(WX793), .ZN(U6408_n1) );
  NOR2X0 U6408_U1 ( .IN1(n3681), .IN2(U6408_n1), .QN(WX856) );
  INVX0 U6409_U2 ( .INP(WX791), .ZN(U6409_n1) );
  NOR2X0 U6409_U1 ( .IN1(n3681), .IN2(U6409_n1), .QN(WX854) );
  INVX0 U6410_U2 ( .INP(WX789), .ZN(U6410_n1) );
  NOR2X0 U6410_U1 ( .IN1(n3681), .IN2(U6410_n1), .QN(WX852) );
  INVX0 U6411_U2 ( .INP(WX787), .ZN(U6411_n1) );
  NOR2X0 U6411_U1 ( .IN1(n3681), .IN2(U6411_n1), .QN(WX850) );
  INVX0 U6412_U2 ( .INP(WX785), .ZN(U6412_n1) );
  NOR2X0 U6412_U1 ( .IN1(n3681), .IN2(U6412_n1), .QN(WX848) );
  INVX0 U6413_U2 ( .INP(WX783), .ZN(U6413_n1) );
  NOR2X0 U6413_U1 ( .IN1(n3681), .IN2(U6413_n1), .QN(WX846) );
  INVX0 U6414_U2 ( .INP(WX781), .ZN(U6414_n1) );
  NOR2X0 U6414_U1 ( .IN1(n3681), .IN2(U6414_n1), .QN(WX844) );
  INVX0 U6415_U2 ( .INP(WX779), .ZN(U6415_n1) );
  NOR2X0 U6415_U1 ( .IN1(n3680), .IN2(U6415_n1), .QN(WX842) );
  INVX0 U6416_U2 ( .INP(WX777), .ZN(U6416_n1) );
  NOR2X0 U6416_U1 ( .IN1(n3680), .IN2(U6416_n1), .QN(WX840) );
  INVX0 U6417_U2 ( .INP(WX775), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n3680), .IN2(U6417_n1), .QN(WX838) );
  INVX0 U6418_U2 ( .INP(WX773), .ZN(U6418_n1) );
  NOR2X0 U6418_U1 ( .IN1(n3680), .IN2(U6418_n1), .QN(WX836) );
  INVX0 U6419_U2 ( .INP(WX771), .ZN(U6419_n1) );
  NOR2X0 U6419_U1 ( .IN1(n3680), .IN2(U6419_n1), .QN(WX834) );
  INVX0 U6420_U2 ( .INP(WX769), .ZN(U6420_n1) );
  NOR2X0 U6420_U1 ( .IN1(n3680), .IN2(U6420_n1), .QN(WX832) );
  INVX0 U6421_U2 ( .INP(WX767), .ZN(U6421_n1) );
  NOR2X0 U6421_U1 ( .IN1(n3680), .IN2(U6421_n1), .QN(WX830) );
  INVX0 U6422_U2 ( .INP(WX765), .ZN(U6422_n1) );
  NOR2X0 U6422_U1 ( .IN1(n3680), .IN2(U6422_n1), .QN(WX828) );
  INVX0 U6423_U2 ( .INP(WX763), .ZN(U6423_n1) );
  NOR2X0 U6423_U1 ( .IN1(n3680), .IN2(U6423_n1), .QN(WX826) );
  INVX0 U6424_U2 ( .INP(WX761), .ZN(U6424_n1) );
  NOR2X0 U6424_U1 ( .IN1(n3680), .IN2(U6424_n1), .QN(WX824) );
  INVX0 U6425_U2 ( .INP(test_so5), .ZN(U6425_n1) );
  NOR2X0 U6425_U1 ( .IN1(n3680), .IN2(U6425_n1), .QN(WX822) );
  INVX0 U6426_U2 ( .INP(WX757), .ZN(U6426_n1) );
  NOR2X0 U6426_U1 ( .IN1(n3679), .IN2(U6426_n1), .QN(WX820) );
  INVX0 U6427_U2 ( .INP(WX755), .ZN(U6427_n1) );
  NOR2X0 U6427_U1 ( .IN1(n3679), .IN2(U6427_n1), .QN(WX818) );
  INVX0 U6428_U2 ( .INP(WX753), .ZN(U6428_n1) );
  NOR2X0 U6428_U1 ( .IN1(n3679), .IN2(U6428_n1), .QN(WX816) );
  INVX0 U6429_U2 ( .INP(WX751), .ZN(U6429_n1) );
  NOR2X0 U6429_U1 ( .IN1(n3679), .IN2(U6429_n1), .QN(WX814) );
  INVX0 U6430_U2 ( .INP(WX749), .ZN(U6430_n1) );
  NOR2X0 U6430_U1 ( .IN1(n3679), .IN2(U6430_n1), .QN(WX812) );
  INVX0 U6431_U2 ( .INP(WX747), .ZN(U6431_n1) );
  NOR2X0 U6431_U1 ( .IN1(n3679), .IN2(U6431_n1), .QN(WX810) );
  INVX0 U6432_U2 ( .INP(WX745), .ZN(U6432_n1) );
  NOR2X0 U6432_U1 ( .IN1(n3679), .IN2(U6432_n1), .QN(WX808) );
  INVX0 U6433_U2 ( .INP(WX743), .ZN(U6433_n1) );
  NOR2X0 U6433_U1 ( .IN1(n3679), .IN2(U6433_n1), .QN(WX806) );
  INVX0 U6434_U2 ( .INP(WX741), .ZN(U6434_n1) );
  NOR2X0 U6434_U1 ( .IN1(n3679), .IN2(U6434_n1), .QN(WX804) );
  INVX0 U6435_U2 ( .INP(WX739), .ZN(U6435_n1) );
  NOR2X0 U6435_U1 ( .IN1(n3679), .IN2(U6435_n1), .QN(WX802) );
  INVX0 U6436_U2 ( .INP(WX737), .ZN(U6436_n1) );
  NOR2X0 U6436_U1 ( .IN1(n3679), .IN2(U6436_n1), .QN(WX800) );
  INVX0 U6437_U2 ( .INP(WX735), .ZN(U6437_n1) );
  NOR2X0 U6437_U1 ( .IN1(n3678), .IN2(U6437_n1), .QN(WX798) );
  INVX0 U6438_U2 ( .INP(WX733), .ZN(U6438_n1) );
  NOR2X0 U6438_U1 ( .IN1(n3678), .IN2(U6438_n1), .QN(WX796) );
  INVX0 U6439_U2 ( .INP(WX731), .ZN(U6439_n1) );
  NOR2X0 U6439_U1 ( .IN1(n3678), .IN2(U6439_n1), .QN(WX794) );
  INVX0 U6440_U2 ( .INP(WX729), .ZN(U6440_n1) );
  NOR2X0 U6440_U1 ( .IN1(n3678), .IN2(U6440_n1), .QN(WX792) );
  INVX0 U6441_U2 ( .INP(WX727), .ZN(U6441_n1) );
  NOR2X0 U6441_U1 ( .IN1(n3678), .IN2(U6441_n1), .QN(WX790) );
  INVX0 U6442_U2 ( .INP(WX725), .ZN(U6442_n1) );
  NOR2X0 U6442_U1 ( .IN1(n3678), .IN2(U6442_n1), .QN(WX788) );
  INVX0 U6443_U2 ( .INP(test_so4), .ZN(U6443_n1) );
  NOR2X0 U6443_U1 ( .IN1(n3678), .IN2(U6443_n1), .QN(WX786) );
  INVX0 U6444_U2 ( .INP(WX721), .ZN(U6444_n1) );
  NOR2X0 U6444_U1 ( .IN1(n3678), .IN2(U6444_n1), .QN(WX784) );
  INVX0 U6445_U2 ( .INP(WX719), .ZN(U6445_n1) );
  NOR2X0 U6445_U1 ( .IN1(n3678), .IN2(U6445_n1), .QN(WX782) );
  INVX0 U6446_U2 ( .INP(WX717), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n3678), .IN2(U6446_n1), .QN(WX780) );
  INVX0 U6447_U2 ( .INP(WX715), .ZN(U6447_n1) );
  NOR2X0 U6447_U1 ( .IN1(n3678), .IN2(U6447_n1), .QN(WX778) );
  INVX0 U6448_U2 ( .INP(WX713), .ZN(U6448_n1) );
  NOR2X0 U6448_U1 ( .IN1(n3677), .IN2(U6448_n1), .QN(WX776) );
  INVX0 U6449_U2 ( .INP(WX711), .ZN(U6449_n1) );
  NOR2X0 U6449_U1 ( .IN1(n3677), .IN2(U6449_n1), .QN(WX774) );
  INVX0 U6450_U2 ( .INP(WX709), .ZN(U6450_n1) );
  NOR2X0 U6450_U1 ( .IN1(n3677), .IN2(U6450_n1), .QN(WX772) );
  INVX0 U6451_U2 ( .INP(WX707), .ZN(U6451_n1) );
  NOR2X0 U6451_U1 ( .IN1(n3677), .IN2(U6451_n1), .QN(WX770) );
  INVX0 U6452_U2 ( .INP(WX705), .ZN(U6452_n1) );
  NOR2X0 U6452_U1 ( .IN1(n3677), .IN2(U6452_n1), .QN(WX768) );
  INVX0 U6453_U2 ( .INP(WX703), .ZN(U6453_n1) );
  NOR2X0 U6453_U1 ( .IN1(n3677), .IN2(U6453_n1), .QN(WX766) );
  INVX0 U6454_U2 ( .INP(WX701), .ZN(U6454_n1) );
  NOR2X0 U6454_U1 ( .IN1(n3677), .IN2(U6454_n1), .QN(WX764) );
  INVX0 U6455_U2 ( .INP(WX699), .ZN(U6455_n1) );
  NOR2X0 U6455_U1 ( .IN1(n3677), .IN2(U6455_n1), .QN(WX762) );
  INVX0 U6456_U2 ( .INP(WX697), .ZN(U6456_n1) );
  NOR2X0 U6456_U1 ( .IN1(n3677), .IN2(U6456_n1), .QN(WX760) );
  INVX0 U6457_U2 ( .INP(WX695), .ZN(U6457_n1) );
  NOR2X0 U6457_U1 ( .IN1(n3677), .IN2(U6457_n1), .QN(WX758) );
  INVX0 U6458_U2 ( .INP(WX693), .ZN(U6458_n1) );
  NOR2X0 U6458_U1 ( .IN1(n3677), .IN2(U6458_n1), .QN(WX756) );
  INVX0 U6459_U2 ( .INP(WX691), .ZN(U6459_n1) );
  NOR2X0 U6459_U1 ( .IN1(n3676), .IN2(U6459_n1), .QN(WX754) );
  INVX0 U6460_U2 ( .INP(WX689), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(n3676), .IN2(U6460_n1), .QN(WX752) );
  INVX0 U6461_U2 ( .INP(test_so3), .ZN(U6461_n1) );
  NOR2X0 U6461_U1 ( .IN1(n3676), .IN2(U6461_n1), .QN(WX750) );
  INVX0 U6462_U2 ( .INP(WX685), .ZN(U6462_n1) );
  NOR2X0 U6462_U1 ( .IN1(n3676), .IN2(U6462_n1), .QN(WX748) );
  INVX0 U6463_U2 ( .INP(WX683), .ZN(U6463_n1) );
  NOR2X0 U6463_U1 ( .IN1(n3676), .IN2(U6463_n1), .QN(WX746) );
  INVX0 U6464_U2 ( .INP(WX681), .ZN(U6464_n1) );
  NOR2X0 U6464_U1 ( .IN1(n3676), .IN2(U6464_n1), .QN(WX744) );
  INVX0 U6465_U2 ( .INP(WX679), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n3676), .IN2(U6465_n1), .QN(WX742) );
  INVX0 U6466_U2 ( .INP(WX677), .ZN(U6466_n1) );
  NOR2X0 U6466_U1 ( .IN1(n3676), .IN2(U6466_n1), .QN(WX740) );
  INVX0 U6467_U2 ( .INP(WX675), .ZN(U6467_n1) );
  NOR2X0 U6467_U1 ( .IN1(n3676), .IN2(U6467_n1), .QN(WX738) );
  INVX0 U6468_U2 ( .INP(WX673), .ZN(U6468_n1) );
  NOR2X0 U6468_U1 ( .IN1(n3676), .IN2(U6468_n1), .QN(WX736) );
  INVX0 U6469_U2 ( .INP(WX671), .ZN(U6469_n1) );
  NOR2X0 U6469_U1 ( .IN1(n3676), .IN2(U6469_n1), .QN(WX734) );
  INVX0 U6470_U2 ( .INP(WX669), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n3675), .IN2(U6470_n1), .QN(WX732) );
  INVX0 U6471_U2 ( .INP(WX667), .ZN(U6471_n1) );
  NOR2X0 U6471_U1 ( .IN1(n3675), .IN2(U6471_n1), .QN(WX730) );
  INVX0 U6472_U2 ( .INP(WX665), .ZN(U6472_n1) );
  NOR2X0 U6472_U1 ( .IN1(n3675), .IN2(U6472_n1), .QN(WX728) );
  INVX0 U6473_U2 ( .INP(WX663), .ZN(U6473_n1) );
  NOR2X0 U6473_U1 ( .IN1(n3675), .IN2(U6473_n1), .QN(WX726) );
  INVX0 U6474_U2 ( .INP(WX661), .ZN(U6474_n1) );
  NOR2X0 U6474_U1 ( .IN1(n3675), .IN2(U6474_n1), .QN(WX724) );
  INVX0 U6475_U2 ( .INP(WX659), .ZN(U6475_n1) );
  NOR2X0 U6475_U1 ( .IN1(n3675), .IN2(U6475_n1), .QN(WX722) );
  INVX0 U6476_U2 ( .INP(WX657), .ZN(U6476_n1) );
  NOR2X0 U6476_U1 ( .IN1(n3675), .IN2(U6476_n1), .QN(WX720) );
  INVX0 U6477_U2 ( .INP(WX655), .ZN(U6477_n1) );
  NOR2X0 U6477_U1 ( .IN1(n3675), .IN2(U6477_n1), .QN(WX718) );
  INVX0 U6478_U2 ( .INP(WX653), .ZN(U6478_n1) );
  NOR2X0 U6478_U1 ( .IN1(n3675), .IN2(U6478_n1), .QN(WX716) );
  INVX0 U6479_U2 ( .INP(test_so2), .ZN(U6479_n1) );
  NOR2X0 U6479_U1 ( .IN1(n3675), .IN2(U6479_n1), .QN(WX714) );
  INVX0 U6480_U2 ( .INP(WX649), .ZN(U6480_n1) );
  NOR2X0 U6480_U1 ( .IN1(n3675), .IN2(U6480_n1), .QN(WX712) );
  INVX0 U6481_U2 ( .INP(WX647), .ZN(U6481_n1) );
  NOR2X0 U6481_U1 ( .IN1(n3674), .IN2(U6481_n1), .QN(WX710) );
  INVX0 U6482_U2 ( .INP(WX645), .ZN(U6482_n1) );
  NOR2X0 U6482_U1 ( .IN1(n3682), .IN2(U6482_n1), .QN(WX708) );
endmodule

