module locked_c1908 (  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n272_, new_n273_, new_n274_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n301_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n310_, new_n311_, new_n313_, new_n314_, new_n315_, new_n316_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n349_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_;
  INV_X1 g000 ( .A(KEYINPUT19), .ZN(new_n123_) );
  XOR2_X1 g001 ( .A(G902), .B(KEYINPUT15), .Z(new_n124_) );
  INV_X1 g002 ( .A(new_n124_), .ZN(new_n125_) );
  XNOR2_X1 g003 ( .A(G113), .B(G116), .ZN(new_n126_) );
  XNOR2_X1 g004 ( .A(G119), .B(KEYINPUT3), .ZN(new_n127_) );
  XNOR2_X1 g005 ( .A(new_n126_), .B(new_n127_), .ZN(new_n128_) );
  XNOR2_X1 g006 ( .A(G122), .B(KEYINPUT16), .ZN(new_n129_) );
  XNOR2_X1 g007 ( .A(new_n128_), .B(new_n129_), .ZN(new_n130_) );
  XOR2_X1 g008 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(new_n131_) );
  INV_X1 g009 ( .A(G953), .ZN(new_n132_) );
  AND2_X1 g010 ( .A1(new_n132_), .A2(G224), .ZN(new_n133_) );
  XNOR2_X1 g011 ( .A(new_n131_), .B(new_n133_), .ZN(new_n134_) );
  XOR2_X1 g012 ( .A(G125), .B(G146), .Z(new_n135_) );
  XNOR2_X1 g013 ( .A(new_n134_), .B(new_n135_), .ZN(new_n136_) );
  XNOR2_X1 g014 ( .A(new_n136_), .B(new_n130_), .ZN(new_n137_) );
  INV_X1 g015 ( .A(KEYINPUT4), .ZN(new_n138_) );
  XOR2_X1 g016 ( .A(G128), .B(G143), .Z(new_n139_) );
  OR2_X1 g017 ( .A1(new_n139_), .A2(new_n138_), .ZN(new_n140_) );
  INV_X1 g018 ( .A(G128), .ZN(new_n141_) );
  INV_X1 g019 ( .A(G143), .ZN(new_n142_) );
  AND2_X1 g020 ( .A1(new_n141_), .A2(new_n142_), .ZN(new_n143_) );
  AND2_X1 g021 ( .A1(G128), .A2(G143), .ZN(new_n144_) );
  OR2_X1 g022 ( .A1(new_n144_), .A2(KEYINPUT4), .ZN(new_n145_) );
  OR2_X1 g023 ( .A1(new_n145_), .A2(new_n143_), .ZN(new_n146_) );
  AND2_X1 g024 ( .A1(new_n146_), .A2(new_n140_), .ZN(new_n147_) );
  XNOR2_X1 g025 ( .A(new_n147_), .B(G101), .ZN(new_n148_) );
  INV_X1 g026 ( .A(G107), .ZN(new_n149_) );
  XNOR2_X1 g027 ( .A(G104), .B(G110), .ZN(new_n150_) );
  XNOR2_X1 g028 ( .A(new_n150_), .B(new_n149_), .ZN(new_n151_) );
  XNOR2_X1 g029 ( .A(new_n148_), .B(new_n151_), .ZN(new_n152_) );
  XNOR2_X1 g030 ( .A(new_n152_), .B(new_n137_), .ZN(new_n153_) );
  AND2_X1 g031 ( .A1(new_n153_), .A2(new_n125_), .ZN(new_n154_) );
  INV_X1 g032 ( .A(G237), .ZN(new_n155_) );
  INV_X1 g033 ( .A(G902), .ZN(new_n156_) );
  AND2_X1 g034 ( .A1(new_n155_), .A2(new_n156_), .ZN(new_n157_) );
  INV_X1 g035 ( .A(new_n157_), .ZN(new_n158_) );
  AND2_X1 g036 ( .A1(new_n158_), .A2(G210), .ZN(new_n159_) );
  INV_X1 g037 ( .A(new_n159_), .ZN(new_n160_) );
  XNOR2_X1 g038 ( .A(new_n154_), .B(new_n160_), .ZN(new_n161_) );
  AND2_X1 g039 ( .A1(new_n158_), .A2(G214), .ZN(new_n162_) );
  INV_X1 g040 ( .A(new_n162_), .ZN(new_n163_) );
  AND2_X1 g041 ( .A1(new_n161_), .A2(new_n163_), .ZN(new_n164_) );
  XNOR2_X1 g042 ( .A(new_n164_), .B(new_n123_), .ZN(new_n165_) );
  AND2_X1 g043 ( .A1(G234), .A2(G237), .ZN(new_n166_) );
  XNOR2_X1 g044 ( .A(new_n166_), .B(KEYINPUT14), .ZN(new_n167_) );
  INV_X1 g045 ( .A(new_n167_), .ZN(new_n168_) );
  AND2_X1 g046 ( .A1(new_n168_), .A2(G952), .ZN(new_n169_) );
  AND2_X1 g047 ( .A1(new_n169_), .A2(new_n132_), .ZN(new_n170_) );
  AND2_X1 g048 ( .A1(new_n168_), .A2(G902), .ZN(new_n171_) );
  OR2_X1 g049 ( .A1(new_n132_), .A2(G898), .ZN(new_n172_) );
  INV_X1 g050 ( .A(new_n172_), .ZN(new_n173_) );
  AND2_X1 g051 ( .A1(new_n171_), .A2(new_n173_), .ZN(new_n174_) );
  OR2_X1 g052 ( .A1(new_n170_), .A2(new_n174_), .ZN(new_n175_) );
  AND2_X1 g053 ( .A1(new_n165_), .A2(new_n175_), .ZN(new_n176_) );
  XNOR2_X1 g054 ( .A(new_n176_), .B(KEYINPUT0), .ZN(new_n177_) );
  AND2_X1 g055 ( .A1(new_n125_), .A2(G234), .ZN(new_n178_) );
  XOR2_X1 g056 ( .A(new_n178_), .B(KEYINPUT20), .Z(new_n179_) );
  AND2_X1 g057 ( .A1(new_n179_), .A2(G221), .ZN(new_n180_) );
  XNOR2_X1 g058 ( .A(new_n180_), .B(KEYINPUT21), .ZN(new_n181_) );
  XOR2_X1 g059 ( .A(G125), .B(KEYINPUT10), .Z(new_n182_) );
  XNOR2_X1 g060 ( .A(G140), .B(KEYINPUT11), .ZN(new_n183_) );
  XNOR2_X1 g061 ( .A(G113), .B(G122), .ZN(new_n184_) );
  XOR2_X1 g062 ( .A(new_n183_), .B(new_n184_), .Z(new_n185_) );
  XNOR2_X1 g063 ( .A(new_n185_), .B(new_n182_), .ZN(new_n186_) );
  XOR2_X1 g064 ( .A(G104), .B(G143), .Z(new_n187_) );
  XNOR2_X1 g065 ( .A(new_n186_), .B(new_n187_), .ZN(new_n188_) );
  XNOR2_X1 g066 ( .A(G131), .B(G146), .ZN(new_n189_) );
  XNOR2_X1 g067 ( .A(new_n189_), .B(KEYINPUT12), .ZN(new_n190_) );
  OR2_X1 g068 ( .A1(G237), .A2(G953), .ZN(new_n191_) );
  INV_X1 g069 ( .A(new_n191_), .ZN(new_n192_) );
  AND2_X1 g070 ( .A1(new_n192_), .A2(G214), .ZN(new_n193_) );
  XNOR2_X1 g071 ( .A(new_n190_), .B(new_n193_), .ZN(new_n194_) );
  XOR2_X1 g072 ( .A(new_n188_), .B(new_n194_), .Z(new_n195_) );
  INV_X1 g073 ( .A(new_n195_), .ZN(new_n196_) );
  AND2_X1 g074 ( .A1(new_n196_), .A2(new_n156_), .ZN(new_n197_) );
  XOR2_X1 g075 ( .A(G475), .B(KEYINPUT13), .Z(new_n198_) );
  XNOR2_X1 g076 ( .A(new_n197_), .B(new_n198_), .ZN(new_n199_) );
  XNOR2_X1 g077 ( .A(new_n139_), .B(G107), .ZN(new_n200_) );
  AND2_X1 g078 ( .A1(new_n132_), .A2(G234), .ZN(new_n201_) );
  XNOR2_X1 g079 ( .A(new_n201_), .B(KEYINPUT8), .ZN(new_n202_) );
  AND2_X1 g080 ( .A1(new_n202_), .A2(G217), .ZN(new_n203_) );
  XNOR2_X1 g081 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(new_n204_) );
  XNOR2_X1 g082 ( .A(new_n203_), .B(new_n204_), .ZN(new_n205_) );
  XNOR2_X1 g083 ( .A(new_n205_), .B(G116), .ZN(new_n206_) );
  XNOR2_X1 g084 ( .A(new_n206_), .B(new_n200_), .ZN(new_n207_) );
  XOR2_X1 g085 ( .A(G122), .B(G134), .Z(new_n208_) );
  XNOR2_X1 g086 ( .A(new_n207_), .B(new_n208_), .ZN(new_n209_) );
  AND2_X1 g087 ( .A1(new_n209_), .A2(new_n156_), .ZN(new_n210_) );
  XNOR2_X1 g088 ( .A(new_n210_), .B(G478), .ZN(new_n211_) );
  AND2_X1 g089 ( .A1(new_n211_), .A2(new_n199_), .ZN(new_n212_) );
  AND2_X1 g090 ( .A1(new_n212_), .A2(new_n181_), .ZN(new_n213_) );
  AND2_X1 g091 ( .A1(new_n177_), .A2(new_n213_), .ZN(new_n214_) );
  XNOR2_X1 g092 ( .A(new_n214_), .B(KEYINPUT22), .ZN(new_n215_) );
  INV_X1 g093 ( .A(KEYINPUT1), .ZN(new_n216_) );
  XNOR2_X1 g094 ( .A(G137), .B(G140), .ZN(new_n217_) );
  INV_X1 g095 ( .A(G134), .ZN(new_n218_) );
  XNOR2_X1 g096 ( .A(new_n189_), .B(new_n218_), .ZN(new_n219_) );
  XNOR2_X1 g097 ( .A(new_n219_), .B(new_n217_), .ZN(new_n220_) );
  AND2_X1 g098 ( .A1(new_n132_), .A2(G227), .ZN(new_n221_) );
  XNOR2_X1 g099 ( .A(new_n220_), .B(new_n221_), .ZN(new_n222_) );
  XNOR2_X1 g100 ( .A(new_n152_), .B(new_n222_), .ZN(new_n223_) );
  AND2_X1 g101 ( .A1(new_n223_), .A2(new_n156_), .ZN(new_n224_) );
  XNOR2_X1 g102 ( .A(new_n224_), .B(G469), .ZN(new_n225_) );
  XNOR2_X1 g103 ( .A(new_n225_), .B(new_n216_), .ZN(new_n226_) );
  INV_X1 g104 ( .A(new_n226_), .ZN(new_n227_) );
  AND2_X1 g105 ( .A1(new_n215_), .A2(new_n227_), .ZN(new_n228_) );
  AND2_X1 g106 ( .A1(new_n202_), .A2(G221), .ZN(new_n229_) );
  XOR2_X1 g107 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(new_n230_) );
  XNOR2_X1 g108 ( .A(new_n229_), .B(new_n230_), .ZN(new_n231_) );
  XNOR2_X1 g109 ( .A(new_n182_), .B(new_n217_), .ZN(new_n232_) );
  XNOR2_X1 g110 ( .A(G119), .B(G146), .ZN(new_n233_) );
  XNOR2_X1 g111 ( .A(G110), .B(G128), .ZN(new_n234_) );
  XNOR2_X1 g112 ( .A(new_n233_), .B(new_n234_), .ZN(new_n235_) );
  XNOR2_X1 g113 ( .A(new_n232_), .B(new_n235_), .ZN(new_n236_) );
  XNOR2_X1 g114 ( .A(new_n231_), .B(new_n236_), .ZN(new_n237_) );
  AND2_X1 g115 ( .A1(new_n237_), .A2(new_n156_), .ZN(new_n238_) );
  AND2_X1 g116 ( .A1(new_n179_), .A2(G217), .ZN(new_n239_) );
  XNOR2_X1 g117 ( .A(new_n238_), .B(new_n239_), .ZN(new_n240_) );
  XOR2_X1 g118 ( .A(new_n240_), .B(KEYINPUT25), .Z(new_n241_) );
  INV_X1 g119 ( .A(G472), .ZN(new_n242_) );
  XNOR2_X1 g120 ( .A(G137), .B(KEYINPUT5), .ZN(new_n243_) );
  AND2_X1 g121 ( .A1(new_n192_), .A2(G210), .ZN(new_n244_) );
  XNOR2_X1 g122 ( .A(new_n244_), .B(new_n243_), .ZN(new_n245_) );
  XNOR2_X1 g123 ( .A(new_n245_), .B(new_n128_), .ZN(new_n246_) );
  XNOR2_X1 g124 ( .A(new_n246_), .B(new_n219_), .ZN(new_n247_) );
  XNOR2_X1 g125 ( .A(new_n247_), .B(new_n148_), .ZN(new_n248_) );
  AND2_X1 g126 ( .A1(new_n248_), .A2(new_n156_), .ZN(new_n249_) );
  XNOR2_X1 g127 ( .A(new_n249_), .B(new_n242_), .ZN(new_n250_) );
  XOR2_X1 g128 ( .A(new_n250_), .B(KEYINPUT6), .Z(new_n251_) );
  INV_X1 g129 ( .A(new_n251_), .ZN(new_n252_) );
  AND2_X1 g130 ( .A1(new_n252_), .A2(new_n241_), .ZN(new_n253_) );
  AND2_X1 g131 ( .A1(new_n228_), .A2(new_n253_), .ZN(new_n254_) );
  XOR2_X1 g132 ( .A(new_n254_), .B(G101), .Z(G3) );
  INV_X1 g133 ( .A(new_n250_), .ZN(new_n256_) );
  INV_X1 g134 ( .A(new_n225_), .ZN(new_n257_) );
  AND2_X1 g135 ( .A1(new_n241_), .A2(new_n181_), .ZN(new_n258_) );
  AND2_X1 g136 ( .A1(new_n258_), .A2(new_n257_), .ZN(new_n259_) );
  AND2_X1 g137 ( .A1(new_n259_), .A2(new_n256_), .ZN(new_n260_) );
  AND2_X1 g138 ( .A1(new_n177_), .A2(new_n260_), .ZN(new_n261_) );
  INV_X1 g139 ( .A(new_n199_), .ZN(new_n262_) );
  AND2_X1 g140 ( .A1(new_n211_), .A2(new_n262_), .ZN(new_n263_) );
  AND2_X1 g141 ( .A1(new_n261_), .A2(new_n263_), .ZN(new_n264_) );
  XOR2_X1 g142 ( .A(new_n264_), .B(G104), .Z(G6) );
  INV_X1 g143 ( .A(new_n211_), .ZN(new_n266_) );
  AND2_X1 g144 ( .A1(new_n266_), .A2(new_n199_), .ZN(new_n267_) );
  AND2_X1 g145 ( .A1(new_n261_), .A2(new_n267_), .ZN(new_n268_) );
  XOR2_X1 g146 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(new_n269_) );
  XNOR2_X1 g147 ( .A(new_n268_), .B(new_n269_), .ZN(new_n270_) );
  XNOR2_X1 g148 ( .A(new_n270_), .B(new_n149_), .ZN(G9) );
  INV_X1 g149 ( .A(new_n241_), .ZN(new_n272_) );
  AND2_X1 g150 ( .A1(new_n272_), .A2(new_n256_), .ZN(new_n273_) );
  AND2_X1 g151 ( .A1(new_n228_), .A2(new_n273_), .ZN(new_n274_) );
  XOR2_X1 g152 ( .A(new_n274_), .B(G110), .Z(G12) );
  INV_X1 g153 ( .A(G900), .ZN(new_n276_) );
  AND2_X1 g154 ( .A1(new_n276_), .A2(G953), .ZN(new_n277_) );
  AND2_X1 g155 ( .A1(new_n171_), .A2(new_n277_), .ZN(new_n278_) );
  OR2_X1 g156 ( .A1(new_n170_), .A2(new_n278_), .ZN(new_n279_) );
  AND2_X1 g157 ( .A1(new_n181_), .A2(new_n279_), .ZN(new_n280_) );
  AND2_X1 g158 ( .A1(new_n272_), .A2(new_n280_), .ZN(new_n281_) );
  AND2_X1 g159 ( .A1(new_n281_), .A2(new_n250_), .ZN(new_n282_) );
  INV_X1 g160 ( .A(new_n282_), .ZN(new_n283_) );
  OR2_X1 g161 ( .A1(new_n283_), .A2(KEYINPUT28), .ZN(new_n284_) );
  INV_X1 g162 ( .A(KEYINPUT28), .ZN(new_n285_) );
  OR2_X1 g163 ( .A1(new_n282_), .A2(new_n285_), .ZN(new_n286_) );
  AND2_X1 g164 ( .A1(new_n286_), .A2(new_n257_), .ZN(new_n287_) );
  AND2_X1 g165 ( .A1(new_n287_), .A2(new_n284_), .ZN(new_n288_) );
  AND2_X1 g166 ( .A1(new_n288_), .A2(new_n165_), .ZN(new_n289_) );
  AND2_X1 g167 ( .A1(new_n289_), .A2(new_n267_), .ZN(new_n290_) );
  XNOR2_X1 g168 ( .A(G128), .B(KEYINPUT29), .ZN(new_n291_) );
  XNOR2_X1 g169 ( .A(new_n290_), .B(new_n291_), .ZN(G30) );
  AND2_X1 g170 ( .A1(new_n250_), .A2(new_n163_), .ZN(new_n293_) );
  XNOR2_X1 g171 ( .A(new_n293_), .B(KEYINPUT30), .ZN(new_n294_) );
  AND2_X1 g172 ( .A1(new_n259_), .A2(new_n279_), .ZN(new_n295_) );
  AND2_X1 g173 ( .A1(new_n295_), .A2(new_n294_), .ZN(new_n296_) );
  AND2_X1 g174 ( .A1(new_n266_), .A2(new_n262_), .ZN(new_n297_) );
  AND2_X1 g175 ( .A1(new_n297_), .A2(new_n161_), .ZN(new_n298_) );
  AND2_X1 g176 ( .A1(new_n296_), .A2(new_n298_), .ZN(new_n299_) );
  XNOR2_X1 g177 ( .A(new_n299_), .B(new_n142_), .ZN(G45) );
  AND2_X1 g178 ( .A1(new_n289_), .A2(new_n263_), .ZN(new_n301_) );
  XOR2_X1 g179 ( .A(new_n301_), .B(G146), .Z(G48) );
  INV_X1 g180 ( .A(new_n263_), .ZN(new_n303_) );
  AND2_X1 g181 ( .A1(new_n226_), .A2(new_n258_), .ZN(new_n304_) );
  AND2_X1 g182 ( .A1(new_n304_), .A2(new_n250_), .ZN(new_n305_) );
  AND2_X1 g183 ( .A1(new_n177_), .A2(new_n305_), .ZN(new_n306_) );
  XNOR2_X1 g184 ( .A(new_n306_), .B(KEYINPUT31), .ZN(new_n307_) );
  OR2_X1 g185 ( .A1(new_n307_), .A2(new_n303_), .ZN(new_n308_) );
  XNOR2_X1 g186 ( .A(new_n308_), .B(G113), .ZN(G15) );
  INV_X1 g187 ( .A(new_n267_), .ZN(new_n310_) );
  OR2_X1 g188 ( .A1(new_n307_), .A2(new_n310_), .ZN(new_n311_) );
  XNOR2_X1 g189 ( .A(new_n311_), .B(G116), .ZN(G18) );
  AND2_X1 g190 ( .A1(new_n252_), .A2(new_n272_), .ZN(new_n313_) );
  AND2_X1 g191 ( .A1(new_n313_), .A2(new_n226_), .ZN(new_n314_) );
  AND2_X1 g192 ( .A1(new_n215_), .A2(new_n314_), .ZN(new_n315_) );
  XNOR2_X1 g193 ( .A(new_n315_), .B(KEYINPUT32), .ZN(new_n316_) );
  XOR2_X1 g194 ( .A(new_n316_), .B(G119), .Z(G21) );
  INV_X1 g195 ( .A(KEYINPUT33), .ZN(new_n318_) );
  AND2_X1 g196 ( .A1(new_n304_), .A2(new_n251_), .ZN(new_n319_) );
  XNOR2_X1 g197 ( .A(new_n319_), .B(new_n318_), .ZN(new_n320_) );
  AND2_X1 g198 ( .A1(new_n177_), .A2(new_n320_), .ZN(new_n321_) );
  INV_X1 g199 ( .A(new_n321_), .ZN(new_n322_) );
  AND2_X1 g200 ( .A1(new_n322_), .A2(KEYINPUT34), .ZN(new_n323_) );
  INV_X1 g201 ( .A(new_n297_), .ZN(new_n324_) );
  INV_X1 g202 ( .A(KEYINPUT34), .ZN(new_n325_) );
  AND2_X1 g203 ( .A1(new_n321_), .A2(new_n325_), .ZN(new_n326_) );
  OR2_X1 g204 ( .A1(new_n326_), .A2(new_n324_), .ZN(new_n327_) );
  OR2_X1 g205 ( .A1(new_n327_), .A2(new_n323_), .ZN(new_n328_) );
  XNOR2_X1 g206 ( .A(new_n328_), .B(KEYINPUT35), .ZN(new_n329_) );
  XOR2_X1 g207 ( .A(new_n329_), .B(G122), .Z(G24) );
  INV_X1 g208 ( .A(KEYINPUT36), .ZN(new_n331_) );
  AND2_X1 g209 ( .A1(new_n251_), .A2(new_n281_), .ZN(new_n332_) );
  AND2_X1 g210 ( .A1(new_n332_), .A2(new_n263_), .ZN(new_n333_) );
  AND2_X1 g211 ( .A1(new_n333_), .A2(new_n164_), .ZN(new_n334_) );
  AND2_X1 g212 ( .A1(new_n334_), .A2(new_n331_), .ZN(new_n335_) );
  INV_X1 g213 ( .A(new_n335_), .ZN(new_n336_) );
  OR2_X1 g214 ( .A1(new_n334_), .A2(new_n331_), .ZN(new_n337_) );
  AND2_X1 g215 ( .A1(new_n337_), .A2(new_n226_), .ZN(new_n338_) );
  AND2_X1 g216 ( .A1(new_n338_), .A2(new_n336_), .ZN(new_n339_) );
  XNOR2_X1 g217 ( .A(new_n339_), .B(G125), .ZN(new_n340_) );
  XNOR2_X1 g218 ( .A(new_n340_), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 g219 ( .A(KEYINPUT40), .ZN(new_n342_) );
  XOR2_X1 g220 ( .A(new_n161_), .B(KEYINPUT38), .Z(new_n343_) );
  AND2_X1 g221 ( .A1(new_n296_), .A2(new_n343_), .ZN(new_n344_) );
  XOR2_X1 g222 ( .A(new_n344_), .B(KEYINPUT39), .Z(new_n345_) );
  AND2_X1 g223 ( .A1(new_n345_), .A2(new_n263_), .ZN(new_n346_) );
  XNOR2_X1 g224 ( .A(new_n346_), .B(new_n342_), .ZN(new_n347_) );
  XNOR2_X1 g225 ( .A(new_n347_), .B(G131), .ZN(G33) );
  AND2_X1 g226 ( .A1(new_n345_), .A2(new_n267_), .ZN(new_n349_) );
  XNOR2_X1 g227 ( .A(new_n349_), .B(new_n218_), .ZN(G36) );
  INV_X1 g228 ( .A(KEYINPUT41), .ZN(new_n351_) );
  AND2_X1 g229 ( .A1(new_n212_), .A2(new_n343_), .ZN(new_n352_) );
  AND2_X1 g230 ( .A1(new_n352_), .A2(new_n163_), .ZN(new_n353_) );
  INV_X1 g231 ( .A(new_n353_), .ZN(new_n354_) );
  OR2_X1 g232 ( .A1(new_n354_), .A2(new_n351_), .ZN(new_n355_) );
  OR2_X1 g233 ( .A1(new_n353_), .A2(KEYINPUT41), .ZN(new_n356_) );
  AND2_X1 g234 ( .A1(new_n288_), .A2(new_n356_), .ZN(new_n357_) );
  AND2_X1 g235 ( .A1(new_n357_), .A2(new_n355_), .ZN(new_n358_) );
  XOR2_X1 g236 ( .A(new_n358_), .B(KEYINPUT42), .Z(new_n359_) );
  XNOR2_X1 g237 ( .A(new_n359_), .B(G137), .ZN(G39) );
  INV_X1 g238 ( .A(KEYINPUT43), .ZN(new_n361_) );
  AND2_X1 g239 ( .A1(new_n227_), .A2(new_n163_), .ZN(new_n362_) );
  AND2_X1 g240 ( .A1(new_n333_), .A2(new_n362_), .ZN(new_n363_) );
  INV_X1 g241 ( .A(new_n363_), .ZN(new_n364_) );
  AND2_X1 g242 ( .A1(new_n364_), .A2(new_n361_), .ZN(new_n365_) );
  AND2_X1 g243 ( .A1(new_n363_), .A2(KEYINPUT43), .ZN(new_n366_) );
  OR2_X1 g244 ( .A1(new_n366_), .A2(new_n161_), .ZN(new_n367_) );
  OR2_X1 g245 ( .A1(new_n367_), .A2(new_n365_), .ZN(new_n368_) );
  XNOR2_X1 g246 ( .A(new_n368_), .B(G140), .ZN(G42) );
  INV_X1 g247 ( .A(KEYINPUT2), .ZN(new_n370_) );
  INV_X1 g248 ( .A(KEYINPUT45), .ZN(new_n371_) );
  INV_X1 g249 ( .A(KEYINPUT44), .ZN(new_n372_) );
  INV_X1 g250 ( .A(new_n329_), .ZN(new_n373_) );
  OR2_X1 g251 ( .A1(new_n316_), .A2(new_n274_), .ZN(new_n374_) );
  INV_X1 g252 ( .A(new_n374_), .ZN(new_n375_) );
  AND2_X1 g253 ( .A1(new_n375_), .A2(new_n373_), .ZN(new_n376_) );
  OR2_X1 g254 ( .A1(new_n376_), .A2(new_n372_), .ZN(new_n377_) );
  OR2_X1 g255 ( .A1(new_n329_), .A2(KEYINPUT44), .ZN(new_n378_) );
  OR2_X1 g256 ( .A1(new_n378_), .A2(new_n374_), .ZN(new_n379_) );
  INV_X1 g257 ( .A(new_n254_), .ZN(new_n380_) );
  AND2_X1 g258 ( .A1(new_n310_), .A2(new_n303_), .ZN(new_n381_) );
  INV_X1 g259 ( .A(new_n261_), .ZN(new_n382_) );
  AND2_X1 g260 ( .A1(new_n307_), .A2(new_n382_), .ZN(new_n383_) );
  OR2_X1 g261 ( .A1(new_n383_), .A2(new_n381_), .ZN(new_n384_) );
  AND2_X1 g262 ( .A1(new_n380_), .A2(new_n384_), .ZN(new_n385_) );
  AND2_X1 g263 ( .A1(new_n379_), .A2(new_n385_), .ZN(new_n386_) );
  AND2_X1 g264 ( .A1(new_n386_), .A2(new_n377_), .ZN(new_n387_) );
  XNOR2_X1 g265 ( .A(new_n387_), .B(new_n371_), .ZN(new_n388_) );
  AND2_X1 g266 ( .A1(new_n347_), .A2(new_n359_), .ZN(new_n389_) );
  XNOR2_X1 g267 ( .A(new_n389_), .B(KEYINPUT46), .ZN(new_n390_) );
  OR2_X1 g268 ( .A1(new_n339_), .A2(new_n299_), .ZN(new_n391_) );
  INV_X1 g269 ( .A(new_n391_), .ZN(new_n392_) );
  INV_X1 g270 ( .A(new_n381_), .ZN(new_n393_) );
  AND2_X1 g271 ( .A1(new_n289_), .A2(new_n393_), .ZN(new_n394_) );
  XNOR2_X1 g272 ( .A(new_n394_), .B(KEYINPUT47), .ZN(new_n395_) );
  AND2_X1 g273 ( .A1(new_n392_), .A2(new_n395_), .ZN(new_n396_) );
  AND2_X1 g274 ( .A1(new_n390_), .A2(new_n396_), .ZN(new_n397_) );
  INV_X1 g275 ( .A(new_n397_), .ZN(new_n398_) );
  OR2_X1 g276 ( .A1(new_n398_), .A2(KEYINPUT48), .ZN(new_n399_) );
  INV_X1 g277 ( .A(KEYINPUT48), .ZN(new_n400_) );
  OR2_X1 g278 ( .A1(new_n397_), .A2(new_n400_), .ZN(new_n401_) );
  INV_X1 g279 ( .A(new_n349_), .ZN(new_n402_) );
  AND2_X1 g280 ( .A1(new_n402_), .A2(new_n368_), .ZN(new_n403_) );
  AND2_X1 g281 ( .A1(new_n401_), .A2(new_n403_), .ZN(new_n404_) );
  AND2_X1 g282 ( .A1(new_n404_), .A2(new_n399_), .ZN(new_n405_) );
  AND2_X1 g283 ( .A1(new_n388_), .A2(new_n405_), .ZN(new_n406_) );
  XNOR2_X1 g284 ( .A(new_n406_), .B(new_n370_), .ZN(new_n407_) );
  INV_X1 g285 ( .A(KEYINPUT52), .ZN(new_n408_) );
  INV_X1 g286 ( .A(KEYINPUT51), .ZN(new_n409_) );
  OR2_X1 g287 ( .A1(new_n226_), .A2(new_n258_), .ZN(new_n410_) );
  INV_X1 g288 ( .A(new_n410_), .ZN(new_n411_) );
  AND2_X1 g289 ( .A1(new_n411_), .A2(KEYINPUT50), .ZN(new_n412_) );
  INV_X1 g290 ( .A(new_n412_), .ZN(new_n413_) );
  OR2_X1 g291 ( .A1(new_n411_), .A2(KEYINPUT50), .ZN(new_n414_) );
  OR2_X1 g292 ( .A1(new_n241_), .A2(new_n181_), .ZN(new_n415_) );
  XNOR2_X1 g293 ( .A(new_n415_), .B(KEYINPUT49), .ZN(new_n416_) );
  OR2_X1 g294 ( .A1(new_n416_), .A2(new_n250_), .ZN(new_n417_) );
  INV_X1 g295 ( .A(new_n417_), .ZN(new_n418_) );
  AND2_X1 g296 ( .A1(new_n418_), .A2(new_n414_), .ZN(new_n419_) );
  AND2_X1 g297 ( .A1(new_n419_), .A2(new_n413_), .ZN(new_n420_) );
  OR2_X1 g298 ( .A1(new_n420_), .A2(new_n305_), .ZN(new_n421_) );
  INV_X1 g299 ( .A(new_n421_), .ZN(new_n422_) );
  AND2_X1 g300 ( .A1(new_n422_), .A2(new_n409_), .ZN(new_n423_) );
  AND2_X1 g301 ( .A1(new_n355_), .A2(new_n356_), .ZN(new_n424_) );
  INV_X1 g302 ( .A(new_n424_), .ZN(new_n425_) );
  AND2_X1 g303 ( .A1(new_n421_), .A2(KEYINPUT51), .ZN(new_n426_) );
  OR2_X1 g304 ( .A1(new_n426_), .A2(new_n425_), .ZN(new_n427_) );
  OR2_X1 g305 ( .A1(new_n427_), .A2(new_n423_), .ZN(new_n428_) );
  AND2_X1 g306 ( .A1(new_n393_), .A2(new_n343_), .ZN(new_n429_) );
  OR2_X1 g307 ( .A1(new_n429_), .A2(new_n212_), .ZN(new_n430_) );
  INV_X1 g308 ( .A(new_n320_), .ZN(new_n431_) );
  INV_X1 g309 ( .A(new_n352_), .ZN(new_n432_) );
  AND2_X1 g310 ( .A1(new_n432_), .A2(new_n162_), .ZN(new_n433_) );
  OR2_X1 g311 ( .A1(new_n431_), .A2(new_n433_), .ZN(new_n434_) );
  INV_X1 g312 ( .A(new_n434_), .ZN(new_n435_) );
  AND2_X1 g313 ( .A1(new_n435_), .A2(new_n430_), .ZN(new_n436_) );
  INV_X1 g314 ( .A(new_n436_), .ZN(new_n437_) );
  AND2_X1 g315 ( .A1(new_n428_), .A2(new_n437_), .ZN(new_n438_) );
  INV_X1 g316 ( .A(new_n438_), .ZN(new_n439_) );
  OR2_X1 g317 ( .A1(new_n439_), .A2(new_n408_), .ZN(new_n440_) );
  OR2_X1 g318 ( .A1(new_n438_), .A2(KEYINPUT52), .ZN(new_n441_) );
  AND2_X1 g319 ( .A1(new_n441_), .A2(new_n169_), .ZN(new_n442_) );
  AND2_X1 g320 ( .A1(new_n442_), .A2(new_n440_), .ZN(new_n443_) );
  AND2_X1 g321 ( .A1(new_n424_), .A2(new_n320_), .ZN(new_n444_) );
  OR2_X1 g322 ( .A1(new_n444_), .A2(G953), .ZN(new_n445_) );
  OR2_X1 g323 ( .A1(new_n443_), .A2(new_n445_), .ZN(new_n446_) );
  OR2_X1 g324 ( .A1(new_n407_), .A2(new_n446_), .ZN(new_n447_) );
  XOR2_X1 g325 ( .A(new_n447_), .B(KEYINPUT53), .Z(G75) );
  AND2_X1 g326 ( .A1(new_n124_), .A2(G210), .ZN(new_n449_) );
  AND2_X1 g327 ( .A1(new_n407_), .A2(new_n449_), .ZN(new_n450_) );
  INV_X1 g328 ( .A(new_n450_), .ZN(new_n451_) );
  XNOR2_X1 g329 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(new_n452_) );
  XNOR2_X1 g330 ( .A(new_n153_), .B(new_n452_), .ZN(new_n453_) );
  OR2_X1 g331 ( .A1(new_n451_), .A2(new_n453_), .ZN(new_n454_) );
  OR2_X1 g332 ( .A1(new_n132_), .A2(G952), .ZN(new_n455_) );
  INV_X1 g333 ( .A(new_n453_), .ZN(new_n456_) );
  OR2_X1 g334 ( .A1(new_n450_), .A2(new_n456_), .ZN(new_n457_) );
  AND2_X1 g335 ( .A1(new_n457_), .A2(new_n455_), .ZN(new_n458_) );
  AND2_X1 g336 ( .A1(new_n458_), .A2(new_n454_), .ZN(new_n459_) );
  XNOR2_X1 g337 ( .A(new_n459_), .B(KEYINPUT56), .ZN(G51) );
  AND2_X1 g338 ( .A1(new_n124_), .A2(G469), .ZN(new_n461_) );
  AND2_X1 g339 ( .A1(new_n407_), .A2(new_n461_), .ZN(new_n462_) );
  XOR2_X1 g340 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(new_n463_) );
  INV_X1 g341 ( .A(new_n463_), .ZN(new_n464_) );
  XNOR2_X1 g342 ( .A(new_n462_), .B(new_n464_), .ZN(new_n465_) );
  INV_X1 g343 ( .A(new_n465_), .ZN(new_n466_) );
  OR2_X1 g344 ( .A1(new_n466_), .A2(new_n223_), .ZN(new_n467_) );
  INV_X1 g345 ( .A(new_n223_), .ZN(new_n468_) );
  OR2_X1 g346 ( .A1(new_n465_), .A2(new_n468_), .ZN(new_n469_) );
  AND2_X1 g347 ( .A1(new_n469_), .A2(new_n455_), .ZN(new_n470_) );
  AND2_X1 g348 ( .A1(new_n470_), .A2(new_n467_), .ZN(G54) );
  XNOR2_X1 g349 ( .A(new_n406_), .B(KEYINPUT2), .ZN(new_n472_) );
  AND2_X1 g350 ( .A1(new_n124_), .A2(G475), .ZN(new_n473_) );
  INV_X1 g351 ( .A(new_n473_), .ZN(new_n474_) );
  OR2_X1 g352 ( .A1(new_n472_), .A2(new_n474_), .ZN(new_n475_) );
  INV_X1 g353 ( .A(new_n475_), .ZN(new_n476_) );
  XOR2_X1 g354 ( .A(new_n195_), .B(KEYINPUT59), .Z(new_n477_) );
  INV_X1 g355 ( .A(new_n477_), .ZN(new_n478_) );
  OR2_X1 g356 ( .A1(new_n476_), .A2(new_n478_), .ZN(new_n479_) );
  OR2_X1 g357 ( .A1(new_n475_), .A2(new_n477_), .ZN(new_n480_) );
  AND2_X1 g358 ( .A1(new_n480_), .A2(new_n455_), .ZN(new_n481_) );
  AND2_X1 g359 ( .A1(new_n481_), .A2(new_n479_), .ZN(new_n482_) );
  XNOR2_X1 g360 ( .A(new_n482_), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 g361 ( .A(new_n209_), .ZN(new_n484_) );
  AND2_X1 g362 ( .A1(new_n124_), .A2(G478), .ZN(new_n485_) );
  AND2_X1 g363 ( .A1(new_n407_), .A2(new_n485_), .ZN(new_n486_) );
  INV_X1 g364 ( .A(new_n486_), .ZN(new_n487_) );
  OR2_X1 g365 ( .A1(new_n487_), .A2(new_n484_), .ZN(new_n488_) );
  OR2_X1 g366 ( .A1(new_n486_), .A2(new_n209_), .ZN(new_n489_) );
  AND2_X1 g367 ( .A1(new_n489_), .A2(new_n455_), .ZN(new_n490_) );
  AND2_X1 g368 ( .A1(new_n490_), .A2(new_n488_), .ZN(G63) );
  AND2_X1 g369 ( .A1(new_n124_), .A2(G217), .ZN(new_n492_) );
  INV_X1 g370 ( .A(new_n492_), .ZN(new_n493_) );
  OR2_X1 g371 ( .A1(new_n472_), .A2(new_n493_), .ZN(new_n494_) );
  INV_X1 g372 ( .A(new_n494_), .ZN(new_n495_) );
  OR2_X1 g373 ( .A1(new_n495_), .A2(new_n237_), .ZN(new_n496_) );
  INV_X1 g374 ( .A(new_n237_), .ZN(new_n497_) );
  OR2_X1 g375 ( .A1(new_n494_), .A2(new_n497_), .ZN(new_n498_) );
  AND2_X1 g376 ( .A1(new_n498_), .A2(new_n455_), .ZN(new_n499_) );
  AND2_X1 g377 ( .A1(new_n499_), .A2(new_n496_), .ZN(G66) );
  AND2_X1 g378 ( .A1(new_n388_), .A2(new_n132_), .ZN(new_n501_) );
  AND2_X1 g379 ( .A1(G224), .A2(G953), .ZN(new_n502_) );
  OR2_X1 g380 ( .A1(new_n502_), .A2(KEYINPUT61), .ZN(new_n503_) );
  AND2_X1 g381 ( .A1(new_n502_), .A2(KEYINPUT61), .ZN(new_n504_) );
  INV_X1 g382 ( .A(new_n504_), .ZN(new_n505_) );
  AND2_X1 g383 ( .A1(new_n505_), .A2(G898), .ZN(new_n506_) );
  AND2_X1 g384 ( .A1(new_n506_), .A2(new_n503_), .ZN(new_n507_) );
  OR2_X1 g385 ( .A1(new_n501_), .A2(new_n507_), .ZN(new_n508_) );
  XNOR2_X1 g386 ( .A(new_n151_), .B(G101), .ZN(new_n509_) );
  INV_X1 g387 ( .A(new_n509_), .ZN(new_n510_) );
  OR2_X1 g388 ( .A1(new_n510_), .A2(new_n130_), .ZN(new_n511_) );
  INV_X1 g389 ( .A(new_n130_), .ZN(new_n512_) );
  OR2_X1 g390 ( .A1(new_n512_), .A2(new_n509_), .ZN(new_n513_) );
  AND2_X1 g391 ( .A1(new_n513_), .A2(new_n172_), .ZN(new_n514_) );
  AND2_X1 g392 ( .A1(new_n514_), .A2(new_n511_), .ZN(new_n515_) );
  XNOR2_X1 g393 ( .A(new_n508_), .B(new_n515_), .ZN(G69) );
  XNOR2_X1 g394 ( .A(new_n147_), .B(new_n182_), .ZN(new_n517_) );
  XOR2_X1 g395 ( .A(new_n517_), .B(new_n220_), .Z(new_n518_) );
  XNOR2_X1 g396 ( .A(new_n405_), .B(new_n518_), .ZN(new_n519_) );
  AND2_X1 g397 ( .A1(new_n519_), .A2(new_n132_), .ZN(new_n520_) );
  XNOR2_X1 g398 ( .A(new_n518_), .B(G227), .ZN(new_n521_) );
  OR2_X1 g399 ( .A1(new_n521_), .A2(new_n276_), .ZN(new_n522_) );
  AND2_X1 g400 ( .A1(new_n522_), .A2(G953), .ZN(new_n523_) );
  OR2_X1 g401 ( .A1(new_n520_), .A2(new_n523_), .ZN(G72) );
  INV_X1 g402 ( .A(KEYINPUT63), .ZN(new_n525_) );
  AND2_X1 g403 ( .A1(new_n124_), .A2(G472), .ZN(new_n526_) );
  INV_X1 g404 ( .A(new_n526_), .ZN(new_n527_) );
  OR2_X1 g405 ( .A1(new_n472_), .A2(new_n527_), .ZN(new_n528_) );
  INV_X1 g406 ( .A(new_n528_), .ZN(new_n529_) );
  XOR2_X1 g407 ( .A(new_n248_), .B(KEYINPUT62), .Z(new_n530_) );
  INV_X1 g408 ( .A(new_n530_), .ZN(new_n531_) );
  OR2_X1 g409 ( .A1(new_n529_), .A2(new_n531_), .ZN(new_n532_) );
  OR2_X1 g410 ( .A1(new_n528_), .A2(new_n530_), .ZN(new_n533_) );
  AND2_X1 g411 ( .A1(new_n533_), .A2(new_n455_), .ZN(new_n534_) );
  AND2_X1 g412 ( .A1(new_n534_), .A2(new_n532_), .ZN(new_n535_) );
  XNOR2_X1 g413 ( .A(new_n535_), .B(new_n525_), .ZN(G57) );
endmodule


