module locked_c2670 (  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n376_, new_n379_, new_n381_, new_n382_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n394_, new_n395_, new_n396_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n504_, new_n505_, new_n507_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n553_, new_n554_, new_n555_, new_n557_, new_n558_, new_n559_, new_n561_, new_n562_, new_n563_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_;
  XNOR2_X1 g000 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 g001 ( .A(G132), .ZN(G219) );
  INV_X1 g002 ( .A(G82), .ZN(G220) );
  INV_X1 g003 ( .A(G96), .ZN(G221) );
  INV_X1 g004 ( .A(G69), .ZN(G235) );
  INV_X1 g005 ( .A(G120), .ZN(G236) );
  INV_X1 g006 ( .A(G57), .ZN(G237) );
  INV_X1 g007 ( .A(G108), .ZN(G238) );
  NAND2_X1 g008 ( .A1(G2078), .A2(G2084), .ZN(new_n367_) );
  NOR2_X1 g009 ( .A1(new_n367_), .A2(KEYINPUT20), .ZN(new_n368_) );
  NAND2_X1 g010 ( .A1(new_n367_), .A2(KEYINPUT20), .ZN(new_n369_) );
  NAND2_X1 g011 ( .A1(new_n369_), .A2(G2090), .ZN(new_n370_) );
  NOR2_X1 g012 ( .A1(new_n370_), .A2(new_n368_), .ZN(new_n371_) );
  NAND2_X1 g013 ( .A1(new_n371_), .A2(KEYINPUT21), .ZN(new_n372_) );
  OR2_X1 g014 ( .A1(new_n371_), .A2(KEYINPUT21), .ZN(new_n373_) );
  AND2_X1 g015 ( .A1(new_n373_), .A2(G2072), .ZN(new_n374_) );
  NAND2_X1 g016 ( .A1(new_n374_), .A2(new_n372_), .ZN(G158) );
  AND2_X1 g017 ( .A1(G2), .A2(G15), .ZN(new_n376_) );
  NAND2_X1 g018 ( .A1(new_n376_), .A2(G661), .ZN(G259) );
  AND2_X1 g019 ( .A1(G94), .A2(G452), .ZN(G173) );
  NAND2_X1 g020 ( .A1(G7), .A2(G661), .ZN(new_n379_) );
  XNOR2_X1 g021 ( .A(new_n379_), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 g022 ( .A(G223), .ZN(new_n381_) );
  NAND2_X1 g023 ( .A1(new_n381_), .A2(G567), .ZN(new_n382_) );
  XOR2_X1 g024 ( .A(new_n382_), .B(KEYINPUT11), .Z(G234) );
  NAND2_X1 g025 ( .A1(new_n381_), .A2(G2106), .ZN(G217) );
  NAND2_X1 g026 ( .A1(G82), .A2(G132), .ZN(new_n385_) );
  XOR2_X1 g027 ( .A(new_n385_), .B(KEYINPUT22), .Z(new_n386_) );
  NOR2_X1 g028 ( .A1(G218), .A2(G221), .ZN(new_n387_) );
  NAND2_X1 g029 ( .A1(new_n386_), .A2(new_n387_), .ZN(new_n388_) );
  NOR2_X1 g030 ( .A1(G237), .A2(G235), .ZN(new_n389_) );
  NOR2_X1 g031 ( .A1(G238), .A2(G236), .ZN(new_n390_) );
  NAND2_X1 g032 ( .A1(new_n389_), .A2(new_n390_), .ZN(new_n391_) );
  NOR2_X1 g033 ( .A1(new_n388_), .A2(new_n391_), .ZN(G325) );
  INV_X1 g034 ( .A(G325), .ZN(G261) );
  NAND2_X1 g035 ( .A1(new_n388_), .A2(G2106), .ZN(new_n394_) );
  NAND2_X1 g036 ( .A1(new_n391_), .A2(G567), .ZN(new_n395_) );
  NAND2_X1 g037 ( .A1(new_n394_), .A2(new_n395_), .ZN(new_n396_) );
  INV_X1 g038 ( .A(new_n396_), .ZN(G319) );
  INV_X1 g039 ( .A(G137), .ZN(new_n398_) );
  NOR2_X1 g040 ( .A1(G2104), .A2(G2105), .ZN(new_n399_) );
  NAND2_X1 g041 ( .A1(new_n399_), .A2(KEYINPUT17), .ZN(new_n400_) );
  INV_X1 g042 ( .A(KEYINPUT17), .ZN(new_n401_) );
  INV_X1 g043 ( .A(G2104), .ZN(new_n402_) );
  INV_X1 g044 ( .A(G2105), .ZN(new_n403_) );
  NAND2_X1 g045 ( .A1(new_n402_), .A2(new_n403_), .ZN(new_n404_) );
  NAND2_X1 g046 ( .A1(new_n404_), .A2(new_n401_), .ZN(new_n405_) );
  NAND2_X1 g047 ( .A1(new_n405_), .A2(new_n400_), .ZN(new_n406_) );
  NOR2_X1 g048 ( .A1(new_n406_), .A2(new_n398_), .ZN(new_n407_) );
  INV_X1 g049 ( .A(KEYINPUT23), .ZN(new_n408_) );
  NAND2_X1 g050 ( .A1(G101), .A2(G2104), .ZN(new_n409_) );
  NOR2_X1 g051 ( .A1(new_n409_), .A2(G2105), .ZN(new_n410_) );
  XNOR2_X1 g052 ( .A(new_n410_), .B(new_n408_), .ZN(new_n411_) );
  NOR2_X1 g053 ( .A1(new_n407_), .A2(new_n411_), .ZN(new_n412_) );
  NAND2_X1 g054 ( .A1(new_n402_), .A2(G125), .ZN(new_n413_) );
  NAND2_X1 g055 ( .A1(G113), .A2(G2104), .ZN(new_n414_) );
  NAND2_X1 g056 ( .A1(new_n413_), .A2(new_n414_), .ZN(new_n415_) );
  NAND2_X1 g057 ( .A1(new_n415_), .A2(G2105), .ZN(new_n416_) );
  NAND2_X1 g058 ( .A1(new_n412_), .A2(new_n416_), .ZN(new_n417_) );
  INV_X1 g059 ( .A(new_n417_), .ZN(G160) );
  XNOR2_X1 g060 ( .A(new_n399_), .B(new_n401_), .ZN(new_n419_) );
  NAND2_X1 g061 ( .A1(new_n419_), .A2(G136), .ZN(new_n420_) );
  INV_X1 g062 ( .A(KEYINPUT44), .ZN(new_n421_) );
  NOR2_X1 g063 ( .A1(new_n403_), .A2(G2104), .ZN(new_n422_) );
  NAND2_X1 g064 ( .A1(new_n422_), .A2(G124), .ZN(new_n423_) );
  NOR2_X1 g065 ( .A1(new_n423_), .A2(new_n421_), .ZN(new_n424_) );
  NAND2_X1 g066 ( .A1(new_n423_), .A2(new_n421_), .ZN(new_n425_) );
  INV_X1 g067 ( .A(new_n425_), .ZN(new_n426_) );
  NOR2_X1 g068 ( .A1(new_n402_), .A2(G2105), .ZN(new_n427_) );
  NAND2_X1 g069 ( .A1(new_n427_), .A2(G100), .ZN(new_n428_) );
  AND2_X1 g070 ( .A1(G2104), .A2(G2105), .ZN(new_n429_) );
  NAND2_X1 g071 ( .A1(new_n429_), .A2(G112), .ZN(new_n430_) );
  NAND2_X1 g072 ( .A1(new_n428_), .A2(new_n430_), .ZN(new_n431_) );
  NOR2_X1 g073 ( .A1(new_n426_), .A2(new_n431_), .ZN(new_n432_) );
  INV_X1 g074 ( .A(new_n432_), .ZN(new_n433_) );
  NOR2_X1 g075 ( .A1(new_n433_), .A2(new_n424_), .ZN(new_n434_) );
  NAND2_X1 g076 ( .A1(new_n434_), .A2(new_n420_), .ZN(new_n435_) );
  INV_X1 g077 ( .A(new_n435_), .ZN(G162) );
  NAND2_X1 g078 ( .A1(new_n419_), .A2(G138), .ZN(new_n437_) );
  AND2_X1 g079 ( .A1(new_n427_), .A2(G102), .ZN(new_n438_) );
  NAND2_X1 g080 ( .A1(new_n429_), .A2(G114), .ZN(new_n439_) );
  NAND2_X1 g081 ( .A1(new_n422_), .A2(G126), .ZN(new_n440_) );
  NAND2_X1 g082 ( .A1(new_n440_), .A2(new_n439_), .ZN(new_n441_) );
  NOR2_X1 g083 ( .A1(new_n441_), .A2(new_n438_), .ZN(new_n442_) );
  NAND2_X1 g084 ( .A1(new_n442_), .A2(new_n437_), .ZN(new_n443_) );
  INV_X1 g085 ( .A(new_n443_), .ZN(G164) );
  INV_X1 g086 ( .A(G543), .ZN(new_n445_) );
  NAND2_X1 g087 ( .A1(new_n445_), .A2(G651), .ZN(new_n446_) );
  XNOR2_X1 g088 ( .A(new_n446_), .B(KEYINPUT1), .ZN(new_n447_) );
  NAND2_X1 g089 ( .A1(new_n447_), .A2(G62), .ZN(new_n448_) );
  NOR2_X1 g090 ( .A1(G543), .A2(G651), .ZN(new_n449_) );
  NAND2_X1 g091 ( .A1(new_n449_), .A2(G88), .ZN(new_n450_) );
  NAND2_X1 g092 ( .A1(new_n448_), .A2(new_n450_), .ZN(new_n451_) );
  INV_X1 g093 ( .A(KEYINPUT0), .ZN(new_n452_) );
  NAND2_X1 g094 ( .A1(new_n452_), .A2(G543), .ZN(new_n453_) );
  NAND2_X1 g095 ( .A1(new_n445_), .A2(KEYINPUT0), .ZN(new_n454_) );
  NAND2_X1 g096 ( .A1(new_n453_), .A2(new_n454_), .ZN(new_n455_) );
  NOR2_X1 g097 ( .A1(new_n455_), .A2(G651), .ZN(new_n456_) );
  NAND2_X1 g098 ( .A1(new_n456_), .A2(G50), .ZN(new_n457_) );
  INV_X1 g099 ( .A(G651), .ZN(new_n458_) );
  NOR2_X1 g100 ( .A1(new_n455_), .A2(new_n458_), .ZN(new_n459_) );
  NAND2_X1 g101 ( .A1(new_n459_), .A2(G75), .ZN(new_n460_) );
  NAND2_X1 g102 ( .A1(new_n457_), .A2(new_n460_), .ZN(new_n461_) );
  NOR2_X1 g103 ( .A1(new_n451_), .A2(new_n461_), .ZN(G166) );
  NAND2_X1 g104 ( .A1(new_n447_), .A2(G63), .ZN(new_n463_) );
  NAND2_X1 g105 ( .A1(new_n456_), .A2(G51), .ZN(new_n464_) );
  NAND2_X1 g106 ( .A1(new_n463_), .A2(new_n464_), .ZN(new_n465_) );
  XOR2_X1 g107 ( .A(new_n465_), .B(KEYINPUT6), .Z(new_n466_) );
  NAND2_X1 g108 ( .A1(new_n459_), .A2(G76), .ZN(new_n467_) );
  NAND2_X1 g109 ( .A1(new_n449_), .A2(G89), .ZN(new_n468_) );
  XNOR2_X1 g110 ( .A(new_n468_), .B(KEYINPUT4), .ZN(new_n469_) );
  NAND2_X1 g111 ( .A1(new_n467_), .A2(new_n469_), .ZN(new_n470_) );
  XNOR2_X1 g112 ( .A(new_n470_), .B(KEYINPUT5), .ZN(new_n471_) );
  NAND2_X1 g113 ( .A1(new_n466_), .A2(new_n471_), .ZN(new_n472_) );
  XNOR2_X1 g114 ( .A(new_n472_), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 g115 ( .A(KEYINPUT9), .ZN(new_n474_) );
  NAND2_X1 g116 ( .A1(new_n459_), .A2(G77), .ZN(new_n475_) );
  NAND2_X1 g117 ( .A1(new_n449_), .A2(G90), .ZN(new_n476_) );
  NAND2_X1 g118 ( .A1(new_n475_), .A2(new_n476_), .ZN(new_n477_) );
  NOR2_X1 g119 ( .A1(new_n477_), .A2(new_n474_), .ZN(new_n478_) );
  NAND2_X1 g120 ( .A1(new_n477_), .A2(new_n474_), .ZN(new_n479_) );
  NAND2_X1 g121 ( .A1(new_n447_), .A2(G64), .ZN(new_n480_) );
  NAND2_X1 g122 ( .A1(new_n456_), .A2(G52), .ZN(new_n481_) );
  AND2_X1 g123 ( .A1(new_n480_), .A2(new_n481_), .ZN(new_n482_) );
  NAND2_X1 g124 ( .A1(new_n479_), .A2(new_n482_), .ZN(new_n483_) );
  NOR2_X1 g125 ( .A1(new_n483_), .A2(new_n478_), .ZN(G171) );
  INV_X1 g126 ( .A(KEYINPUT14), .ZN(new_n485_) );
  NAND2_X1 g127 ( .A1(new_n447_), .A2(G56), .ZN(new_n486_) );
  NOR2_X1 g128 ( .A1(new_n486_), .A2(new_n485_), .ZN(new_n487_) );
  NAND2_X1 g129 ( .A1(new_n486_), .A2(new_n485_), .ZN(new_n488_) );
  NAND2_X1 g130 ( .A1(new_n456_), .A2(G43), .ZN(new_n489_) );
  NAND2_X1 g131 ( .A1(new_n488_), .A2(new_n489_), .ZN(new_n490_) );
  NOR2_X1 g132 ( .A1(new_n490_), .A2(new_n487_), .ZN(new_n491_) );
  NAND2_X1 g133 ( .A1(new_n459_), .A2(G68), .ZN(new_n492_) );
  NAND2_X1 g134 ( .A1(new_n449_), .A2(G81), .ZN(new_n493_) );
  NAND2_X1 g135 ( .A1(new_n493_), .A2(KEYINPUT12), .ZN(new_n494_) );
  INV_X1 g136 ( .A(KEYINPUT12), .ZN(new_n495_) );
  AND2_X1 g137 ( .A1(new_n449_), .A2(G81), .ZN(new_n496_) );
  NAND2_X1 g138 ( .A1(new_n496_), .A2(new_n495_), .ZN(new_n497_) );
  NAND2_X1 g139 ( .A1(new_n497_), .A2(new_n494_), .ZN(new_n498_) );
  NAND2_X1 g140 ( .A1(new_n492_), .A2(new_n498_), .ZN(new_n499_) );
  XNOR2_X1 g141 ( .A(new_n499_), .B(KEYINPUT13), .ZN(new_n500_) );
  NAND2_X1 g142 ( .A1(new_n500_), .A2(new_n491_), .ZN(new_n501_) );
  INV_X1 g143 ( .A(new_n501_), .ZN(new_n502_) );
  NAND2_X1 g144 ( .A1(new_n502_), .A2(G860), .ZN(G153) );
  NAND2_X1 g145 ( .A1(G483), .A2(G661), .ZN(new_n504_) );
  NOR2_X1 g146 ( .A1(new_n396_), .A2(new_n504_), .ZN(new_n505_) );
  NAND2_X1 g147 ( .A1(new_n505_), .A2(G36), .ZN(G176) );
  NAND2_X1 g148 ( .A1(G1), .A2(G3), .ZN(new_n507_) );
  NAND2_X1 g149 ( .A1(new_n505_), .A2(new_n507_), .ZN(G188) );
  NAND2_X1 g150 ( .A1(new_n447_), .A2(G65), .ZN(new_n509_) );
  NAND2_X1 g151 ( .A1(new_n449_), .A2(G91), .ZN(new_n510_) );
  NAND2_X1 g152 ( .A1(new_n509_), .A2(new_n510_), .ZN(new_n511_) );
  NAND2_X1 g153 ( .A1(new_n459_), .A2(G78), .ZN(new_n512_) );
  NAND2_X1 g154 ( .A1(new_n456_), .A2(G53), .ZN(new_n513_) );
  NAND2_X1 g155 ( .A1(new_n513_), .A2(new_n512_), .ZN(new_n514_) );
  NOR2_X1 g156 ( .A1(new_n511_), .A2(new_n514_), .ZN(new_n515_) );
  INV_X1 g157 ( .A(new_n515_), .ZN(G299) );
  INV_X1 g158 ( .A(G171), .ZN(G301) );
  XOR2_X1 g159 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 g160 ( .A(G166), .ZN(G303) );
  NAND2_X1 g161 ( .A1(new_n456_), .A2(G49), .ZN(new_n520_) );
  NAND2_X1 g162 ( .A1(new_n455_), .A2(G87), .ZN(new_n521_) );
  AND2_X1 g163 ( .A1(G74), .A2(G651), .ZN(new_n522_) );
  NOR2_X1 g164 ( .A1(new_n447_), .A2(new_n522_), .ZN(new_n523_) );
  AND2_X1 g165 ( .A1(new_n523_), .A2(new_n521_), .ZN(new_n524_) );
  NAND2_X1 g166 ( .A1(new_n524_), .A2(new_n520_), .ZN(G288) );
  NAND2_X1 g167 ( .A1(new_n459_), .A2(G73), .ZN(new_n526_) );
  XNOR2_X1 g168 ( .A(new_n526_), .B(KEYINPUT2), .ZN(new_n527_) );
  AND2_X1 g169 ( .A1(new_n456_), .A2(G48), .ZN(new_n528_) );
  NAND2_X1 g170 ( .A1(new_n447_), .A2(G61), .ZN(new_n529_) );
  NAND2_X1 g171 ( .A1(new_n449_), .A2(G86), .ZN(new_n530_) );
  NAND2_X1 g172 ( .A1(new_n529_), .A2(new_n530_), .ZN(new_n531_) );
  NOR2_X1 g173 ( .A1(new_n531_), .A2(new_n528_), .ZN(new_n532_) );
  NAND2_X1 g174 ( .A1(new_n527_), .A2(new_n532_), .ZN(G305) );
  NAND2_X1 g175 ( .A1(new_n447_), .A2(G60), .ZN(new_n534_) );
  NAND2_X1 g176 ( .A1(new_n449_), .A2(G85), .ZN(new_n535_) );
  NAND2_X1 g177 ( .A1(new_n534_), .A2(new_n535_), .ZN(new_n536_) );
  NAND2_X1 g178 ( .A1(new_n456_), .A2(G47), .ZN(new_n537_) );
  NAND2_X1 g179 ( .A1(new_n459_), .A2(G72), .ZN(new_n538_) );
  NAND2_X1 g180 ( .A1(new_n537_), .A2(new_n538_), .ZN(new_n539_) );
  NOR2_X1 g181 ( .A1(new_n536_), .A2(new_n539_), .ZN(new_n540_) );
  INV_X1 g182 ( .A(new_n540_), .ZN(G290) );
  NAND2_X1 g183 ( .A1(new_n447_), .A2(G66), .ZN(new_n542_) );
  NAND2_X1 g184 ( .A1(new_n449_), .A2(G92), .ZN(new_n543_) );
  NAND2_X1 g185 ( .A1(new_n542_), .A2(new_n543_), .ZN(new_n544_) );
  NAND2_X1 g186 ( .A1(new_n456_), .A2(G54), .ZN(new_n545_) );
  NAND2_X1 g187 ( .A1(new_n459_), .A2(G79), .ZN(new_n546_) );
  NAND2_X1 g188 ( .A1(new_n545_), .A2(new_n546_), .ZN(new_n547_) );
  OR2_X1 g189 ( .A1(new_n544_), .A2(new_n547_), .ZN(new_n548_) );
  XNOR2_X1 g190 ( .A(new_n548_), .B(KEYINPUT15), .ZN(new_n549_) );
  OR2_X1 g191 ( .A1(new_n549_), .A2(G868), .ZN(new_n550_) );
  NAND2_X1 g192 ( .A1(G301), .A2(G868), .ZN(new_n551_) );
  NAND2_X1 g193 ( .A1(new_n550_), .A2(new_n551_), .ZN(G284) );
  INV_X1 g194 ( .A(G868), .ZN(new_n553_) );
  NOR2_X1 g195 ( .A1(G286), .A2(new_n553_), .ZN(new_n554_) );
  NOR2_X1 g196 ( .A1(G299), .A2(G868), .ZN(new_n555_) );
  NOR2_X1 g197 ( .A1(new_n554_), .A2(new_n555_), .ZN(G297) );
  INV_X1 g198 ( .A(G860), .ZN(new_n557_) );
  NAND2_X1 g199 ( .A1(new_n557_), .A2(G559), .ZN(new_n558_) );
  NAND2_X1 g200 ( .A1(new_n549_), .A2(new_n558_), .ZN(new_n559_) );
  XNOR2_X1 g201 ( .A(new_n559_), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 g202 ( .A1(new_n553_), .A2(G559), .ZN(new_n561_) );
  NAND2_X1 g203 ( .A1(new_n549_), .A2(new_n561_), .ZN(new_n562_) );
  NAND2_X1 g204 ( .A1(new_n502_), .A2(new_n553_), .ZN(new_n563_) );
  AND2_X1 g205 ( .A1(new_n562_), .A2(new_n563_), .ZN(G282) );
  NAND2_X1 g206 ( .A1(new_n419_), .A2(G135), .ZN(new_n565_) );
  INV_X1 g207 ( .A(KEYINPUT18), .ZN(new_n566_) );
  NAND2_X1 g208 ( .A1(new_n422_), .A2(G123), .ZN(new_n567_) );
  NOR2_X1 g209 ( .A1(new_n567_), .A2(new_n566_), .ZN(new_n568_) );
  NAND2_X1 g210 ( .A1(new_n567_), .A2(new_n566_), .ZN(new_n569_) );
  INV_X1 g211 ( .A(new_n569_), .ZN(new_n570_) );
  NAND2_X1 g212 ( .A1(new_n427_), .A2(G99), .ZN(new_n571_) );
  NAND2_X1 g213 ( .A1(new_n429_), .A2(G111), .ZN(new_n572_) );
  NAND2_X1 g214 ( .A1(new_n571_), .A2(new_n572_), .ZN(new_n573_) );
  NOR2_X1 g215 ( .A1(new_n570_), .A2(new_n573_), .ZN(new_n574_) );
  INV_X1 g216 ( .A(new_n574_), .ZN(new_n575_) );
  NOR2_X1 g217 ( .A1(new_n575_), .A2(new_n568_), .ZN(new_n576_) );
  NAND2_X1 g218 ( .A1(new_n576_), .A2(new_n565_), .ZN(new_n577_) );
  NAND2_X1 g219 ( .A1(new_n577_), .A2(G2096), .ZN(new_n578_) );
  NOR2_X1 g220 ( .A1(new_n577_), .A2(G2096), .ZN(new_n579_) );
  NOR2_X1 g221 ( .A1(new_n579_), .A2(G2100), .ZN(new_n580_) );
  NAND2_X1 g222 ( .A1(new_n580_), .A2(new_n578_), .ZN(G156) );
  XNOR2_X1 g223 ( .A(G2430), .B(G2454), .ZN(new_n582_) );
  XNOR2_X1 g224 ( .A(G1341), .B(G1348), .ZN(new_n583_) );
  XNOR2_X1 g225 ( .A(new_n582_), .B(new_n583_), .ZN(new_n584_) );
  XNOR2_X1 g226 ( .A(G2435), .B(G2438), .ZN(new_n585_) );
  XNOR2_X1 g227 ( .A(new_n584_), .B(new_n585_), .ZN(new_n586_) );
  XOR2_X1 g228 ( .A(G2446), .B(G2451), .Z(new_n587_) );
  XNOR2_X1 g229 ( .A(G2427), .B(G2443), .ZN(new_n588_) );
  XNOR2_X1 g230 ( .A(new_n587_), .B(new_n588_), .ZN(new_n589_) );
  NOR2_X1 g231 ( .A1(new_n586_), .A2(new_n589_), .ZN(new_n590_) );
  NAND2_X1 g232 ( .A1(new_n586_), .A2(new_n589_), .ZN(new_n591_) );
  NAND2_X1 g233 ( .A1(new_n591_), .A2(G14), .ZN(new_n592_) );
  NOR2_X1 g234 ( .A1(new_n592_), .A2(new_n590_), .ZN(G401) );
  XNOR2_X1 g235 ( .A(G2096), .B(G2100), .ZN(new_n594_) );
  XNOR2_X1 g236 ( .A(G2678), .B(KEYINPUT43), .ZN(new_n595_) );
  XNOR2_X1 g237 ( .A(new_n594_), .B(new_n595_), .ZN(new_n596_) );
  XNOR2_X1 g238 ( .A(G2090), .B(KEYINPUT42), .ZN(new_n597_) );
  XNOR2_X1 g239 ( .A(G2067), .B(G2072), .ZN(new_n598_) );
  XNOR2_X1 g240 ( .A(new_n597_), .B(new_n598_), .ZN(new_n599_) );
  XNOR2_X1 g241 ( .A(new_n596_), .B(new_n599_), .ZN(new_n600_) );
  XOR2_X1 g242 ( .A(G2078), .B(G2084), .Z(new_n601_) );
  XNOR2_X1 g243 ( .A(new_n600_), .B(new_n601_), .ZN(G227) );
  XNOR2_X1 g244 ( .A(G1976), .B(G1981), .ZN(new_n603_) );
  XNOR2_X1 g245 ( .A(G1956), .B(G1966), .ZN(new_n604_) );
  XNOR2_X1 g246 ( .A(new_n603_), .B(new_n604_), .ZN(new_n605_) );
  XNOR2_X1 g247 ( .A(new_n605_), .B(G2474), .ZN(new_n606_) );
  XNOR2_X1 g248 ( .A(G1991), .B(G1996), .ZN(new_n607_) );
  XNOR2_X1 g249 ( .A(new_n606_), .B(new_n607_), .ZN(new_n608_) );
  XOR2_X1 g250 ( .A(G1971), .B(KEYINPUT41), .Z(new_n609_) );
  XNOR2_X1 g251 ( .A(G1961), .B(G1986), .ZN(new_n610_) );
  XNOR2_X1 g252 ( .A(new_n609_), .B(new_n610_), .ZN(new_n611_) );
  XNOR2_X1 g253 ( .A(new_n608_), .B(new_n611_), .ZN(G229) );
  INV_X1 g254 ( .A(G29), .ZN(new_n613_) );
  NAND2_X1 g255 ( .A1(new_n422_), .A2(G127), .ZN(new_n614_) );
  NAND2_X1 g256 ( .A1(new_n429_), .A2(G115), .ZN(new_n615_) );
  NAND2_X1 g257 ( .A1(new_n614_), .A2(new_n615_), .ZN(new_n616_) );
  INV_X1 g258 ( .A(new_n616_), .ZN(new_n617_) );
  OR2_X1 g259 ( .A1(new_n617_), .A2(KEYINPUT47), .ZN(new_n618_) );
  NAND2_X1 g260 ( .A1(new_n427_), .A2(G103), .ZN(new_n619_) );
  NAND2_X1 g261 ( .A1(new_n618_), .A2(new_n619_), .ZN(new_n620_) );
  NAND2_X1 g262 ( .A1(new_n419_), .A2(G139), .ZN(new_n621_) );
  NAND2_X1 g263 ( .A1(new_n617_), .A2(KEYINPUT47), .ZN(new_n622_) );
  NAND2_X1 g264 ( .A1(new_n622_), .A2(new_n621_), .ZN(new_n623_) );
  NOR2_X1 g265 ( .A1(new_n620_), .A2(new_n623_), .ZN(new_n624_) );
  XNOR2_X1 g266 ( .A(new_n624_), .B(G2072), .ZN(new_n625_) );
  XOR2_X1 g267 ( .A(new_n443_), .B(G2078), .Z(new_n626_) );
  NAND2_X1 g268 ( .A1(new_n625_), .A2(new_n626_), .ZN(new_n627_) );
  NOR2_X1 g269 ( .A1(new_n627_), .A2(KEYINPUT50), .ZN(new_n628_) );
  INV_X1 g270 ( .A(KEYINPUT51), .ZN(new_n629_) );
  INV_X1 g271 ( .A(G2090), .ZN(new_n630_) );
  XNOR2_X1 g272 ( .A(new_n435_), .B(new_n630_), .ZN(new_n631_) );
  NAND2_X1 g273 ( .A1(new_n419_), .A2(G141), .ZN(new_n632_) );
  INV_X1 g274 ( .A(KEYINPUT38), .ZN(new_n633_) );
  NAND2_X1 g275 ( .A1(new_n427_), .A2(G105), .ZN(new_n634_) );
  NOR2_X1 g276 ( .A1(new_n634_), .A2(new_n633_), .ZN(new_n635_) );
  NAND2_X1 g277 ( .A1(new_n634_), .A2(new_n633_), .ZN(new_n636_) );
  INV_X1 g278 ( .A(new_n636_), .ZN(new_n637_) );
  NAND2_X1 g279 ( .A1(new_n422_), .A2(G129), .ZN(new_n638_) );
  NAND2_X1 g280 ( .A1(new_n429_), .A2(G117), .ZN(new_n639_) );
  NAND2_X1 g281 ( .A1(new_n638_), .A2(new_n639_), .ZN(new_n640_) );
  NOR2_X1 g282 ( .A1(new_n637_), .A2(new_n640_), .ZN(new_n641_) );
  INV_X1 g283 ( .A(new_n641_), .ZN(new_n642_) );
  NOR2_X1 g284 ( .A1(new_n642_), .A2(new_n635_), .ZN(new_n643_) );
  NAND2_X1 g285 ( .A1(new_n643_), .A2(new_n632_), .ZN(new_n644_) );
  OR2_X1 g286 ( .A1(new_n644_), .A2(G1996), .ZN(new_n645_) );
  NAND2_X1 g287 ( .A1(new_n631_), .A2(new_n645_), .ZN(new_n646_) );
  NAND2_X1 g288 ( .A1(new_n646_), .A2(new_n629_), .ZN(new_n647_) );
  NAND2_X1 g289 ( .A1(new_n627_), .A2(KEYINPUT50), .ZN(new_n648_) );
  NAND2_X1 g290 ( .A1(new_n647_), .A2(new_n648_), .ZN(new_n649_) );
  NOR2_X1 g291 ( .A1(new_n649_), .A2(new_n628_), .ZN(new_n650_) );
  NAND2_X1 g292 ( .A1(new_n419_), .A2(G140), .ZN(new_n651_) );
  NAND2_X1 g293 ( .A1(new_n427_), .A2(G104), .ZN(new_n652_) );
  NAND2_X1 g294 ( .A1(new_n651_), .A2(new_n652_), .ZN(new_n653_) );
  NOR2_X1 g295 ( .A1(new_n653_), .A2(KEYINPUT34), .ZN(new_n654_) );
  NAND2_X1 g296 ( .A1(new_n653_), .A2(KEYINPUT34), .ZN(new_n655_) );
  NAND2_X1 g297 ( .A1(new_n422_), .A2(G128), .ZN(new_n656_) );
  NAND2_X1 g298 ( .A1(new_n429_), .A2(G116), .ZN(new_n657_) );
  NAND2_X1 g299 ( .A1(new_n656_), .A2(new_n657_), .ZN(new_n658_) );
  XNOR2_X1 g300 ( .A(new_n658_), .B(KEYINPUT35), .ZN(new_n659_) );
  NAND2_X1 g301 ( .A1(new_n655_), .A2(new_n659_), .ZN(new_n660_) );
  NOR2_X1 g302 ( .A1(new_n660_), .A2(new_n654_), .ZN(new_n661_) );
  XNOR2_X1 g303 ( .A(new_n661_), .B(KEYINPUT36), .ZN(new_n662_) );
  XNOR2_X1 g304 ( .A(G2067), .B(KEYINPUT37), .ZN(new_n663_) );
  NOR2_X1 g305 ( .A1(new_n662_), .A2(new_n663_), .ZN(new_n664_) );
  NAND2_X1 g306 ( .A1(new_n662_), .A2(new_n663_), .ZN(new_n665_) );
  NOR2_X1 g307 ( .A1(new_n646_), .A2(new_n629_), .ZN(new_n666_) );
  NAND2_X1 g308 ( .A1(new_n644_), .A2(G1996), .ZN(new_n667_) );
  NAND2_X1 g309 ( .A1(new_n419_), .A2(G131), .ZN(new_n668_) );
  NAND2_X1 g310 ( .A1(new_n422_), .A2(G119), .ZN(new_n669_) );
  INV_X1 g311 ( .A(new_n669_), .ZN(new_n670_) );
  NAND2_X1 g312 ( .A1(new_n427_), .A2(G95), .ZN(new_n671_) );
  NAND2_X1 g313 ( .A1(new_n429_), .A2(G107), .ZN(new_n672_) );
  NAND2_X1 g314 ( .A1(new_n671_), .A2(new_n672_), .ZN(new_n673_) );
  NOR2_X1 g315 ( .A1(new_n673_), .A2(new_n670_), .ZN(new_n674_) );
  NAND2_X1 g316 ( .A1(new_n674_), .A2(new_n668_), .ZN(new_n675_) );
  NAND2_X1 g317 ( .A1(new_n675_), .A2(G1991), .ZN(new_n676_) );
  NAND2_X1 g318 ( .A1(new_n667_), .A2(new_n676_), .ZN(new_n677_) );
  INV_X1 g319 ( .A(G2084), .ZN(new_n678_) );
  XNOR2_X1 g320 ( .A(new_n417_), .B(new_n678_), .ZN(new_n679_) );
  INV_X1 g321 ( .A(new_n577_), .ZN(new_n680_) );
  NOR2_X1 g322 ( .A1(new_n675_), .A2(G1991), .ZN(new_n681_) );
  NOR2_X1 g323 ( .A1(new_n680_), .A2(new_n681_), .ZN(new_n682_) );
  NAND2_X1 g324 ( .A1(new_n682_), .A2(new_n679_), .ZN(new_n683_) );
  OR2_X1 g325 ( .A1(new_n683_), .A2(new_n677_), .ZN(new_n684_) );
  NOR2_X1 g326 ( .A1(new_n666_), .A2(new_n684_), .ZN(new_n685_) );
  NAND2_X1 g327 ( .A1(new_n685_), .A2(new_n665_), .ZN(new_n686_) );
  NOR2_X1 g328 ( .A1(new_n686_), .A2(new_n664_), .ZN(new_n687_) );
  NAND2_X1 g329 ( .A1(new_n687_), .A2(new_n650_), .ZN(new_n688_) );
  NOR2_X1 g330 ( .A1(new_n688_), .A2(KEYINPUT52), .ZN(new_n689_) );
  AND2_X1 g331 ( .A1(new_n688_), .A2(KEYINPUT52), .ZN(new_n690_) );
  OR2_X1 g332 ( .A1(new_n690_), .A2(KEYINPUT55), .ZN(new_n691_) );
  NOR2_X1 g333 ( .A1(new_n691_), .A2(new_n689_), .ZN(new_n692_) );
  NOR2_X1 g334 ( .A1(new_n692_), .A2(new_n613_), .ZN(new_n693_) );
  INV_X1 g335 ( .A(G168), .ZN(new_n694_) );
  NAND2_X1 g336 ( .A1(new_n694_), .A2(G1966), .ZN(new_n695_) );
  NOR2_X1 g337 ( .A1(new_n694_), .A2(G1966), .ZN(new_n696_) );
  XNOR2_X1 g338 ( .A(G305), .B(G1981), .ZN(new_n697_) );
  NOR2_X1 g339 ( .A1(new_n696_), .A2(new_n697_), .ZN(new_n698_) );
  NAND2_X1 g340 ( .A1(new_n698_), .A2(new_n695_), .ZN(new_n699_) );
  XNOR2_X1 g341 ( .A(new_n699_), .B(KEYINPUT57), .ZN(new_n700_) );
  XNOR2_X1 g342 ( .A(new_n549_), .B(G1348), .ZN(new_n701_) );
  XNOR2_X1 g343 ( .A(new_n515_), .B(G1956), .ZN(new_n702_) );
  NAND2_X1 g344 ( .A1(G288), .A2(G1976), .ZN(new_n703_) );
  INV_X1 g345 ( .A(new_n703_), .ZN(new_n704_) );
  INV_X1 g346 ( .A(G1971), .ZN(new_n705_) );
  NOR2_X1 g347 ( .A1(G166), .A2(new_n705_), .ZN(new_n706_) );
  NOR2_X1 g348 ( .A1(new_n704_), .A2(new_n706_), .ZN(new_n707_) );
  NAND2_X1 g349 ( .A1(new_n707_), .A2(new_n702_), .ZN(new_n708_) );
  NOR2_X1 g350 ( .A1(G303), .A2(G1971), .ZN(new_n709_) );
  NOR2_X1 g351 ( .A1(G288), .A2(G1976), .ZN(new_n710_) );
  NOR2_X1 g352 ( .A1(new_n709_), .A2(new_n710_), .ZN(new_n711_) );
  XNOR2_X1 g353 ( .A(new_n540_), .B(G1986), .ZN(new_n712_) );
  NAND2_X1 g354 ( .A1(new_n711_), .A2(new_n712_), .ZN(new_n713_) );
  NOR2_X1 g355 ( .A1(new_n708_), .A2(new_n713_), .ZN(new_n714_) );
  NAND2_X1 g356 ( .A1(new_n714_), .A2(new_n701_), .ZN(new_n715_) );
  INV_X1 g357 ( .A(G1341), .ZN(new_n716_) );
  XNOR2_X1 g358 ( .A(new_n501_), .B(new_n716_), .ZN(new_n717_) );
  XNOR2_X1 g359 ( .A(G171), .B(G1961), .ZN(new_n718_) );
  NAND2_X1 g360 ( .A1(new_n717_), .A2(new_n718_), .ZN(new_n719_) );
  NOR2_X1 g361 ( .A1(new_n715_), .A2(new_n719_), .ZN(new_n720_) );
  NAND2_X1 g362 ( .A1(new_n700_), .A2(new_n720_), .ZN(new_n721_) );
  XNOR2_X1 g363 ( .A(G16), .B(KEYINPUT56), .ZN(new_n722_) );
  NAND2_X1 g364 ( .A1(new_n721_), .A2(new_n722_), .ZN(new_n723_) );
  INV_X1 g365 ( .A(KEYINPUT53), .ZN(new_n724_) );
  XNOR2_X1 g366 ( .A(G32), .B(G1996), .ZN(new_n725_) );
  OR2_X1 g367 ( .A1(G33), .A2(G2072), .ZN(new_n726_) );
  AND2_X1 g368 ( .A1(new_n726_), .A2(G28), .ZN(new_n727_) );
  XOR2_X1 g369 ( .A(G26), .B(G2067), .Z(new_n728_) );
  NAND2_X1 g370 ( .A1(new_n727_), .A2(new_n728_), .ZN(new_n729_) );
  NOR2_X1 g371 ( .A1(new_n729_), .A2(new_n725_), .ZN(new_n730_) );
  INV_X1 g372 ( .A(G27), .ZN(new_n731_) );
  XNOR2_X1 g373 ( .A(G2078), .B(KEYINPUT25), .ZN(new_n732_) );
  NOR2_X1 g374 ( .A1(new_n732_), .A2(new_n731_), .ZN(new_n733_) );
  NAND2_X1 g375 ( .A1(new_n732_), .A2(new_n731_), .ZN(new_n734_) );
  NOR2_X1 g376 ( .A1(G25), .A2(G1991), .ZN(new_n735_) );
  NAND2_X1 g377 ( .A1(G33), .A2(G2072), .ZN(new_n736_) );
  NAND2_X1 g378 ( .A1(G25), .A2(G1991), .ZN(new_n737_) );
  NAND2_X1 g379 ( .A1(new_n736_), .A2(new_n737_), .ZN(new_n738_) );
  NOR2_X1 g380 ( .A1(new_n738_), .A2(new_n735_), .ZN(new_n739_) );
  NAND2_X1 g381 ( .A1(new_n734_), .A2(new_n739_), .ZN(new_n740_) );
  NOR2_X1 g382 ( .A1(new_n740_), .A2(new_n733_), .ZN(new_n741_) );
  NAND2_X1 g383 ( .A1(new_n741_), .A2(new_n730_), .ZN(new_n742_) );
  NOR2_X1 g384 ( .A1(new_n742_), .A2(new_n724_), .ZN(new_n743_) );
  NAND2_X1 g385 ( .A1(new_n742_), .A2(new_n724_), .ZN(new_n744_) );
  XNOR2_X1 g386 ( .A(G2084), .B(KEYINPUT54), .ZN(new_n745_) );
  NOR2_X1 g387 ( .A1(new_n745_), .A2(G34), .ZN(new_n746_) );
  NAND2_X1 g388 ( .A1(new_n745_), .A2(G34), .ZN(new_n747_) );
  XOR2_X1 g389 ( .A(G35), .B(G2090), .Z(new_n748_) );
  NAND2_X1 g390 ( .A1(new_n747_), .A2(new_n748_), .ZN(new_n749_) );
  NOR2_X1 g391 ( .A1(new_n749_), .A2(new_n746_), .ZN(new_n750_) );
  NAND2_X1 g392 ( .A1(new_n744_), .A2(new_n750_), .ZN(new_n751_) );
  OR2_X1 g393 ( .A1(new_n751_), .A2(new_n743_), .ZN(new_n752_) );
  NOR2_X1 g394 ( .A1(new_n752_), .A2(KEYINPUT55), .ZN(new_n753_) );
  NAND2_X1 g395 ( .A1(new_n752_), .A2(KEYINPUT55), .ZN(new_n754_) );
  NAND2_X1 g396 ( .A1(new_n754_), .A2(new_n613_), .ZN(new_n755_) );
  NOR2_X1 g397 ( .A1(new_n755_), .A2(new_n753_), .ZN(new_n756_) );
  XNOR2_X1 g398 ( .A(G1348), .B(KEYINPUT59), .ZN(new_n757_) );
  XNOR2_X1 g399 ( .A(new_n757_), .B(G4), .ZN(new_n758_) );
  XNOR2_X1 g400 ( .A(G20), .B(G1956), .ZN(new_n759_) );
  XOR2_X1 g401 ( .A(G19), .B(G1341), .Z(new_n760_) );
  XOR2_X1 g402 ( .A(G6), .B(G1981), .Z(new_n761_) );
  NAND2_X1 g403 ( .A1(new_n760_), .A2(new_n761_), .ZN(new_n762_) );
  NOR2_X1 g404 ( .A1(new_n762_), .A2(new_n759_), .ZN(new_n763_) );
  NAND2_X1 g405 ( .A1(new_n763_), .A2(new_n758_), .ZN(new_n764_) );
  XNOR2_X1 g406 ( .A(new_n764_), .B(KEYINPUT60), .ZN(new_n765_) );
  XOR2_X1 g407 ( .A(G24), .B(G1986), .Z(new_n766_) );
  NOR2_X1 g408 ( .A1(G22), .A2(G1971), .ZN(new_n767_) );
  NOR2_X1 g409 ( .A1(G23), .A2(G1976), .ZN(new_n768_) );
  OR2_X1 g410 ( .A1(new_n767_), .A2(new_n768_), .ZN(new_n769_) );
  NAND2_X1 g411 ( .A1(G23), .A2(G1976), .ZN(new_n770_) );
  NAND2_X1 g412 ( .A1(G22), .A2(G1971), .ZN(new_n771_) );
  NAND2_X1 g413 ( .A1(new_n770_), .A2(new_n771_), .ZN(new_n772_) );
  NOR2_X1 g414 ( .A1(new_n769_), .A2(new_n772_), .ZN(new_n773_) );
  NAND2_X1 g415 ( .A1(new_n773_), .A2(new_n766_), .ZN(new_n774_) );
  NOR2_X1 g416 ( .A1(new_n774_), .A2(KEYINPUT58), .ZN(new_n775_) );
  NAND2_X1 g417 ( .A1(new_n774_), .A2(KEYINPUT58), .ZN(new_n776_) );
  NOR2_X1 g418 ( .A1(G21), .A2(G1966), .ZN(new_n777_) );
  NOR2_X1 g419 ( .A1(G5), .A2(G1961), .ZN(new_n778_) );
  OR2_X1 g420 ( .A1(new_n777_), .A2(new_n778_), .ZN(new_n779_) );
  NAND2_X1 g421 ( .A1(G5), .A2(G1961), .ZN(new_n780_) );
  NAND2_X1 g422 ( .A1(G21), .A2(G1966), .ZN(new_n781_) );
  NAND2_X1 g423 ( .A1(new_n780_), .A2(new_n781_), .ZN(new_n782_) );
  NOR2_X1 g424 ( .A1(new_n779_), .A2(new_n782_), .ZN(new_n783_) );
  NAND2_X1 g425 ( .A1(new_n776_), .A2(new_n783_), .ZN(new_n784_) );
  NOR2_X1 g426 ( .A1(new_n784_), .A2(new_n775_), .ZN(new_n785_) );
  INV_X1 g427 ( .A(new_n785_), .ZN(new_n786_) );
  NOR2_X1 g428 ( .A1(new_n786_), .A2(new_n765_), .ZN(new_n787_) );
  INV_X1 g429 ( .A(new_n787_), .ZN(new_n788_) );
  OR2_X1 g430 ( .A1(new_n788_), .A2(KEYINPUT61), .ZN(new_n789_) );
  AND2_X1 g431 ( .A1(new_n788_), .A2(KEYINPUT61), .ZN(new_n790_) );
  NOR2_X1 g432 ( .A1(new_n790_), .A2(G16), .ZN(new_n791_) );
  NAND2_X1 g433 ( .A1(new_n791_), .A2(new_n789_), .ZN(new_n792_) );
  NAND2_X1 g434 ( .A1(new_n792_), .A2(G11), .ZN(new_n793_) );
  NOR2_X1 g435 ( .A1(new_n793_), .A2(new_n756_), .ZN(new_n794_) );
  NAND2_X1 g436 ( .A1(new_n723_), .A2(new_n794_), .ZN(new_n795_) );
  NOR2_X1 g437 ( .A1(new_n693_), .A2(new_n795_), .ZN(new_n796_) );
  XNOR2_X1 g438 ( .A(new_n796_), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 g439 ( .A(G311), .ZN(G150) );
  NAND2_X1 g440 ( .A1(new_n549_), .A2(G559), .ZN(new_n799_) );
  NOR2_X1 g441 ( .A1(new_n799_), .A2(new_n501_), .ZN(new_n800_) );
  NAND2_X1 g442 ( .A1(new_n799_), .A2(new_n501_), .ZN(new_n801_) );
  NAND2_X1 g443 ( .A1(new_n801_), .A2(new_n557_), .ZN(new_n802_) );
  NOR2_X1 g444 ( .A1(new_n802_), .A2(new_n800_), .ZN(new_n803_) );
  NAND2_X1 g445 ( .A1(new_n447_), .A2(G67), .ZN(new_n804_) );
  NAND2_X1 g446 ( .A1(new_n449_), .A2(G93), .ZN(new_n805_) );
  NAND2_X1 g447 ( .A1(new_n804_), .A2(new_n805_), .ZN(new_n806_) );
  NAND2_X1 g448 ( .A1(new_n456_), .A2(G55), .ZN(new_n807_) );
  NAND2_X1 g449 ( .A1(new_n459_), .A2(G80), .ZN(new_n808_) );
  NAND2_X1 g450 ( .A1(new_n807_), .A2(new_n808_), .ZN(new_n809_) );
  NOR2_X1 g451 ( .A1(new_n806_), .A2(new_n809_), .ZN(new_n810_) );
  XNOR2_X1 g452 ( .A(new_n803_), .B(new_n810_), .ZN(G145) );
  XNOR2_X1 g453 ( .A(new_n624_), .B(new_n417_), .ZN(new_n812_) );
  XNOR2_X1 g454 ( .A(new_n662_), .B(new_n812_), .ZN(new_n813_) );
  INV_X1 g455 ( .A(KEYINPUT45), .ZN(new_n814_) );
  NAND2_X1 g456 ( .A1(new_n419_), .A2(G142), .ZN(new_n815_) );
  NAND2_X1 g457 ( .A1(new_n427_), .A2(G106), .ZN(new_n816_) );
  NAND2_X1 g458 ( .A1(new_n815_), .A2(new_n816_), .ZN(new_n817_) );
  NAND2_X1 g459 ( .A1(new_n817_), .A2(new_n814_), .ZN(new_n818_) );
  NOR2_X1 g460 ( .A1(new_n817_), .A2(new_n814_), .ZN(new_n819_) );
  NAND2_X1 g461 ( .A1(new_n422_), .A2(G130), .ZN(new_n820_) );
  NAND2_X1 g462 ( .A1(new_n429_), .A2(G118), .ZN(new_n821_) );
  NAND2_X1 g463 ( .A1(new_n820_), .A2(new_n821_), .ZN(new_n822_) );
  NOR2_X1 g464 ( .A1(new_n819_), .A2(new_n822_), .ZN(new_n823_) );
  NAND2_X1 g465 ( .A1(new_n823_), .A2(new_n818_), .ZN(new_n824_) );
  XNOR2_X1 g466 ( .A(new_n824_), .B(new_n644_), .ZN(new_n825_) );
  XNOR2_X1 g467 ( .A(new_n825_), .B(new_n435_), .ZN(new_n826_) );
  XNOR2_X1 g468 ( .A(new_n826_), .B(new_n813_), .ZN(new_n827_) );
  XNOR2_X1 g469 ( .A(new_n577_), .B(new_n675_), .ZN(new_n828_) );
  XNOR2_X1 g470 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(new_n829_) );
  XNOR2_X1 g471 ( .A(new_n828_), .B(new_n829_), .ZN(new_n830_) );
  XNOR2_X1 g472 ( .A(new_n830_), .B(G164), .ZN(new_n831_) );
  NOR2_X1 g473 ( .A1(new_n827_), .A2(new_n831_), .ZN(new_n832_) );
  INV_X1 g474 ( .A(G37), .ZN(new_n833_) );
  NAND2_X1 g475 ( .A1(new_n827_), .A2(new_n831_), .ZN(new_n834_) );
  NAND2_X1 g476 ( .A1(new_n834_), .A2(new_n833_), .ZN(new_n835_) );
  NOR2_X1 g477 ( .A1(new_n835_), .A2(new_n832_), .ZN(G395) );
  XNOR2_X1 g478 ( .A(new_n501_), .B(G290), .ZN(new_n837_) );
  XNOR2_X1 g479 ( .A(new_n837_), .B(G288), .ZN(new_n838_) );
  XOR2_X1 g480 ( .A(new_n515_), .B(KEYINPUT19), .Z(new_n839_) );
  XNOR2_X1 g481 ( .A(new_n839_), .B(G305), .ZN(new_n840_) );
  XNOR2_X1 g482 ( .A(new_n838_), .B(new_n840_), .ZN(new_n841_) );
  XNOR2_X1 g483 ( .A(G166), .B(new_n810_), .ZN(new_n842_) );
  XNOR2_X1 g484 ( .A(new_n841_), .B(new_n842_), .ZN(new_n843_) );
  XOR2_X1 g485 ( .A(new_n843_), .B(new_n799_), .Z(new_n844_) );
  NAND2_X1 g486 ( .A1(new_n844_), .A2(G868), .ZN(new_n845_) );
  OR2_X1 g487 ( .A1(new_n810_), .A2(G868), .ZN(new_n846_) );
  NAND2_X1 g488 ( .A1(new_n845_), .A2(new_n846_), .ZN(G295) );
  XNOR2_X1 g489 ( .A(G286), .B(new_n549_), .ZN(new_n848_) );
  XNOR2_X1 g490 ( .A(new_n843_), .B(new_n848_), .ZN(new_n849_) );
  NOR2_X1 g491 ( .A1(new_n849_), .A2(G171), .ZN(new_n850_) );
  NAND2_X1 g492 ( .A1(new_n849_), .A2(G171), .ZN(new_n851_) );
  NAND2_X1 g493 ( .A1(new_n851_), .A2(new_n833_), .ZN(new_n852_) );
  NOR2_X1 g494 ( .A1(new_n852_), .A2(new_n850_), .ZN(G397) );
  INV_X1 g495 ( .A(KEYINPUT40), .ZN(new_n854_) );
  INV_X1 g496 ( .A(KEYINPUT33), .ZN(new_n855_) );
  INV_X1 g497 ( .A(KEYINPUT32), .ZN(new_n856_) );
  INV_X1 g498 ( .A(KEYINPUT26), .ZN(new_n857_) );
  INV_X1 g499 ( .A(G1384), .ZN(new_n858_) );
  NAND2_X1 g500 ( .A1(new_n443_), .A2(new_n858_), .ZN(new_n859_) );
  AND2_X1 g501 ( .A1(new_n416_), .A2(G40), .ZN(new_n860_) );
  NAND2_X1 g502 ( .A1(new_n412_), .A2(new_n860_), .ZN(new_n861_) );
  NOR2_X1 g503 ( .A1(new_n861_), .A2(new_n859_), .ZN(new_n862_) );
  NAND2_X1 g504 ( .A1(new_n862_), .A2(G1996), .ZN(new_n863_) );
  NOR2_X1 g505 ( .A1(new_n863_), .A2(new_n857_), .ZN(new_n864_) );
  NAND2_X1 g506 ( .A1(new_n863_), .A2(new_n857_), .ZN(new_n865_) );
  NOR2_X1 g507 ( .A1(new_n862_), .A2(new_n716_), .ZN(new_n866_) );
  NOR2_X1 g508 ( .A1(new_n866_), .A2(new_n501_), .ZN(new_n867_) );
  NAND2_X1 g509 ( .A1(new_n867_), .A2(new_n865_), .ZN(new_n868_) );
  NOR2_X1 g510 ( .A1(new_n868_), .A2(new_n864_), .ZN(new_n869_) );
  NAND2_X1 g511 ( .A1(new_n869_), .A2(new_n549_), .ZN(new_n870_) );
  INV_X1 g512 ( .A(new_n862_), .ZN(new_n871_) );
  NAND2_X1 g513 ( .A1(new_n871_), .A2(G1348), .ZN(new_n872_) );
  NAND2_X1 g514 ( .A1(new_n862_), .A2(G2067), .ZN(new_n873_) );
  NAND2_X1 g515 ( .A1(new_n872_), .A2(new_n873_), .ZN(new_n874_) );
  NAND2_X1 g516 ( .A1(new_n870_), .A2(new_n874_), .ZN(new_n875_) );
  OR2_X1 g517 ( .A1(new_n869_), .A2(new_n549_), .ZN(new_n876_) );
  NAND2_X1 g518 ( .A1(new_n875_), .A2(new_n876_), .ZN(new_n877_) );
  NAND2_X1 g519 ( .A1(new_n862_), .A2(G2072), .ZN(new_n878_) );
  NOR2_X1 g520 ( .A1(new_n878_), .A2(KEYINPUT27), .ZN(new_n879_) );
  NAND2_X1 g521 ( .A1(new_n878_), .A2(KEYINPUT27), .ZN(new_n880_) );
  NAND2_X1 g522 ( .A1(new_n871_), .A2(G1956), .ZN(new_n881_) );
  NAND2_X1 g523 ( .A1(new_n880_), .A2(new_n881_), .ZN(new_n882_) );
  NOR2_X1 g524 ( .A1(new_n882_), .A2(new_n879_), .ZN(new_n883_) );
  NAND2_X1 g525 ( .A1(new_n883_), .A2(new_n515_), .ZN(new_n884_) );
  NAND2_X1 g526 ( .A1(new_n877_), .A2(new_n884_), .ZN(new_n885_) );
  OR2_X1 g527 ( .A1(new_n883_), .A2(new_n515_), .ZN(new_n886_) );
  XNOR2_X1 g528 ( .A(new_n886_), .B(KEYINPUT28), .ZN(new_n887_) );
  NAND2_X1 g529 ( .A1(new_n885_), .A2(new_n887_), .ZN(new_n888_) );
  OR2_X1 g530 ( .A1(new_n888_), .A2(KEYINPUT29), .ZN(new_n889_) );
  NAND2_X1 g531 ( .A1(new_n888_), .A2(KEYINPUT29), .ZN(new_n890_) );
  OR2_X1 g532 ( .A1(new_n862_), .A2(G1961), .ZN(new_n891_) );
  NAND2_X1 g533 ( .A1(new_n862_), .A2(new_n732_), .ZN(new_n892_) );
  NAND2_X1 g534 ( .A1(new_n891_), .A2(new_n892_), .ZN(new_n893_) );
  NAND2_X1 g535 ( .A1(new_n893_), .A2(G171), .ZN(new_n894_) );
  AND2_X1 g536 ( .A1(new_n890_), .A2(new_n894_), .ZN(new_n895_) );
  NAND2_X1 g537 ( .A1(new_n895_), .A2(new_n889_), .ZN(new_n896_) );
  INV_X1 g538 ( .A(KEYINPUT30), .ZN(new_n897_) );
  NAND2_X1 g539 ( .A1(new_n871_), .A2(G8), .ZN(new_n898_) );
  NOR2_X1 g540 ( .A1(new_n898_), .A2(G1966), .ZN(new_n899_) );
  NAND2_X1 g541 ( .A1(new_n862_), .A2(new_n678_), .ZN(new_n900_) );
  NAND2_X1 g542 ( .A1(new_n900_), .A2(G8), .ZN(new_n901_) );
  NOR2_X1 g543 ( .A1(new_n899_), .A2(new_n901_), .ZN(new_n902_) );
  NAND2_X1 g544 ( .A1(new_n902_), .A2(new_n897_), .ZN(new_n903_) );
  NOR2_X1 g545 ( .A1(new_n902_), .A2(new_n897_), .ZN(new_n904_) );
  NOR2_X1 g546 ( .A1(new_n904_), .A2(G168), .ZN(new_n905_) );
  AND2_X1 g547 ( .A1(new_n905_), .A2(new_n903_), .ZN(new_n906_) );
  NOR2_X1 g548 ( .A1(new_n893_), .A2(G171), .ZN(new_n907_) );
  NOR2_X1 g549 ( .A1(new_n906_), .A2(new_n907_), .ZN(new_n908_) );
  XOR2_X1 g550 ( .A(new_n908_), .B(KEYINPUT31), .Z(new_n909_) );
  NAND2_X1 g551 ( .A1(new_n896_), .A2(new_n909_), .ZN(new_n910_) );
  NAND2_X1 g552 ( .A1(new_n910_), .A2(G286), .ZN(new_n911_) );
  INV_X1 g553 ( .A(new_n898_), .ZN(new_n912_) );
  NAND2_X1 g554 ( .A1(new_n912_), .A2(new_n705_), .ZN(new_n913_) );
  NOR2_X1 g555 ( .A1(new_n871_), .A2(G2090), .ZN(new_n914_) );
  NOR2_X1 g556 ( .A1(new_n914_), .A2(G166), .ZN(new_n915_) );
  NAND2_X1 g557 ( .A1(new_n913_), .A2(new_n915_), .ZN(new_n916_) );
  NAND2_X1 g558 ( .A1(new_n911_), .A2(new_n916_), .ZN(new_n917_) );
  NAND2_X1 g559 ( .A1(new_n917_), .A2(G8), .ZN(new_n918_) );
  NOR2_X1 g560 ( .A1(new_n918_), .A2(new_n856_), .ZN(new_n919_) );
  INV_X1 g561 ( .A(new_n919_), .ZN(new_n920_) );
  NAND2_X1 g562 ( .A1(new_n918_), .A2(new_n856_), .ZN(new_n921_) );
  INV_X1 g563 ( .A(G8), .ZN(new_n922_) );
  NOR2_X1 g564 ( .A1(new_n900_), .A2(new_n922_), .ZN(new_n923_) );
  NOR2_X1 g565 ( .A1(new_n899_), .A2(new_n923_), .ZN(new_n924_) );
  NAND2_X1 g566 ( .A1(new_n910_), .A2(new_n924_), .ZN(new_n925_) );
  AND2_X1 g567 ( .A1(new_n921_), .A2(new_n925_), .ZN(new_n926_) );
  NAND2_X1 g568 ( .A1(new_n926_), .A2(new_n920_), .ZN(new_n927_) );
  NAND2_X1 g569 ( .A1(new_n927_), .A2(new_n711_), .ZN(new_n928_) );
  NOR2_X1 g570 ( .A1(new_n898_), .A2(new_n704_), .ZN(new_n929_) );
  NAND2_X1 g571 ( .A1(new_n928_), .A2(new_n929_), .ZN(new_n930_) );
  NAND2_X1 g572 ( .A1(new_n930_), .A2(new_n855_), .ZN(new_n931_) );
  NAND2_X1 g573 ( .A1(new_n710_), .A2(KEYINPUT33), .ZN(new_n932_) );
  NOR2_X1 g574 ( .A1(new_n898_), .A2(new_n932_), .ZN(new_n933_) );
  NOR2_X1 g575 ( .A1(new_n933_), .A2(new_n697_), .ZN(new_n934_) );
  NAND2_X1 g576 ( .A1(new_n931_), .A2(new_n934_), .ZN(new_n935_) );
  NAND2_X1 g577 ( .A1(new_n921_), .A2(new_n925_), .ZN(new_n936_) );
  NOR2_X1 g578 ( .A1(new_n936_), .A2(new_n919_), .ZN(new_n937_) );
  NAND2_X1 g579 ( .A1(new_n630_), .A2(G8), .ZN(new_n938_) );
  NOR2_X1 g580 ( .A1(G303), .A2(new_n938_), .ZN(new_n939_) );
  NOR2_X1 g581 ( .A1(new_n937_), .A2(new_n939_), .ZN(new_n940_) );
  NOR2_X1 g582 ( .A1(new_n940_), .A2(new_n912_), .ZN(new_n941_) );
  INV_X1 g583 ( .A(KEYINPUT24), .ZN(new_n942_) );
  NOR2_X1 g584 ( .A1(G305), .A2(G1981), .ZN(new_n943_) );
  NOR2_X1 g585 ( .A1(new_n943_), .A2(new_n942_), .ZN(new_n944_) );
  NAND2_X1 g586 ( .A1(new_n943_), .A2(new_n942_), .ZN(new_n945_) );
  NAND2_X1 g587 ( .A1(new_n912_), .A2(new_n945_), .ZN(new_n946_) );
  NOR2_X1 g588 ( .A1(new_n946_), .A2(new_n944_), .ZN(new_n947_) );
  NOR2_X1 g589 ( .A1(new_n941_), .A2(new_n947_), .ZN(new_n948_) );
  NAND2_X1 g590 ( .A1(new_n935_), .A2(new_n948_), .ZN(new_n949_) );
  INV_X1 g591 ( .A(new_n861_), .ZN(new_n950_) );
  NAND2_X1 g592 ( .A1(new_n950_), .A2(new_n859_), .ZN(new_n951_) );
  INV_X1 g593 ( .A(new_n951_), .ZN(new_n952_) );
  AND2_X1 g594 ( .A1(new_n664_), .A2(new_n952_), .ZN(new_n953_) );
  OR2_X1 g595 ( .A1(new_n712_), .A2(new_n951_), .ZN(new_n954_) );
  NAND2_X1 g596 ( .A1(new_n677_), .A2(new_n952_), .ZN(new_n955_) );
  NAND2_X1 g597 ( .A1(new_n954_), .A2(new_n955_), .ZN(new_n956_) );
  NOR2_X1 g598 ( .A1(new_n953_), .A2(new_n956_), .ZN(new_n957_) );
  NAND2_X1 g599 ( .A1(new_n949_), .A2(new_n957_), .ZN(new_n958_) );
  INV_X1 g600 ( .A(KEYINPUT39), .ZN(new_n959_) );
  NOR2_X1 g601 ( .A1(G290), .A2(G1986), .ZN(new_n960_) );
  OR2_X1 g602 ( .A1(new_n960_), .A2(new_n681_), .ZN(new_n961_) );
  NAND2_X1 g603 ( .A1(new_n955_), .A2(new_n961_), .ZN(new_n962_) );
  AND2_X1 g604 ( .A1(new_n962_), .A2(new_n645_), .ZN(new_n963_) );
  NAND2_X1 g605 ( .A1(new_n963_), .A2(new_n959_), .ZN(new_n964_) );
  NOR2_X1 g606 ( .A1(new_n963_), .A2(new_n959_), .ZN(new_n965_) );
  NOR2_X1 g607 ( .A1(new_n965_), .A2(new_n953_), .ZN(new_n966_) );
  NAND2_X1 g608 ( .A1(new_n966_), .A2(new_n964_), .ZN(new_n967_) );
  NAND2_X1 g609 ( .A1(new_n967_), .A2(new_n665_), .ZN(new_n968_) );
  NAND2_X1 g610 ( .A1(new_n968_), .A2(new_n952_), .ZN(new_n969_) );
  AND2_X1 g611 ( .A1(new_n958_), .A2(new_n969_), .ZN(new_n970_) );
  NAND2_X1 g612 ( .A1(new_n970_), .A2(new_n854_), .ZN(new_n971_) );
  NAND2_X1 g613 ( .A1(new_n958_), .A2(new_n969_), .ZN(new_n972_) );
  NAND2_X1 g614 ( .A1(new_n972_), .A2(KEYINPUT40), .ZN(new_n973_) );
  NAND2_X1 g615 ( .A1(new_n971_), .A2(new_n973_), .ZN(G329) );
  NOR2_X1 g616 ( .A1(G229), .A2(G227), .ZN(new_n976_) );
  NAND2_X1 g617 ( .A1(new_n976_), .A2(KEYINPUT49), .ZN(new_n977_) );
  NOR2_X1 g618 ( .A1(new_n976_), .A2(KEYINPUT49), .ZN(new_n978_) );
  OR2_X1 g619 ( .A1(G401), .A2(new_n396_), .ZN(new_n979_) );
  NOR2_X1 g620 ( .A1(new_n978_), .A2(new_n979_), .ZN(new_n980_) );
  NAND2_X1 g621 ( .A1(new_n980_), .A2(new_n977_), .ZN(new_n981_) );
  OR2_X1 g622 ( .A1(G395), .A2(new_n981_), .ZN(new_n982_) );
  NOR2_X1 g623 ( .A1(G397), .A2(new_n982_), .ZN(G308) );
  INV_X1 g624 ( .A(G308), .ZN(G225) );
  assign   G231 = 1'b0;
  BUF_X1 g625 ( .A(G452), .Z(G350) );
  BUF_X1 g626 ( .A(G452), .Z(G335) );
  BUF_X1 g627 ( .A(G452), .Z(G409) );
  BUF_X1 g628 ( .A(G1083), .Z(G369) );
  BUF_X1 g629 ( .A(G1083), .Z(G367) );
  BUF_X1 g630 ( .A(G2066), .Z(G411) );
  BUF_X1 g631 ( .A(G2066), .Z(G337) );
  BUF_X1 g632 ( .A(G2066), .Z(G384) );
  BUF_X1 g633 ( .A(G452), .Z(G391) );
  NAND2_X1 g634 ( .A1(new_n550_), .A2(new_n551_), .ZN(G321) );
  NOR2_X1 g635 ( .A1(new_n554_), .A2(new_n555_), .ZN(G280) );
  AND2_X1 g636 ( .A1(new_n562_), .A2(new_n563_), .ZN(G323) );
  NAND2_X1 g637 ( .A1(new_n845_), .A2(new_n846_), .ZN(G331) );
endmodule


