module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n1233_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n608_, new_n501_, new_n1157_, new_n421_, new_n777_, new_n1048_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n1327_, new_n566_, new_n641_, new_n339_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n728_, new_n1071_, new_n1294_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n1213_, new_n752_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n721_, new_n504_, new_n742_, new_n892_, new_n472_, new_n873_, new_n1167_, new_n774_, new_n792_, new_n953_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n655_, new_n1054_, new_n630_, new_n1288_, new_n385_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n297_, new_n565_, new_n1196_, new_n511_, new_n303_, new_n325_, new_n1285_, new_n1031_, new_n1216_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n324_, new_n960_, new_n491_, new_n549_, new_n676_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1062_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1275_, new_n1277_, new_n1198_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n1333_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n267_, new_n473_, new_n1147_, new_n1229_, new_n969_, new_n334_, new_n331_, new_n835_, new_n1234_, new_n378_, new_n621_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n1315_, new_n1003_, new_n696_, new_n1039_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n729_, new_n1111_, new_n1218_, new_n559_, new_n1282_, new_n762_, new_n1193_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n295_, new_n1256_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n1032_, new_n867_, new_n954_, new_n901_, new_n1171_, new_n276_, new_n688_, new_n1255_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n296_, new_n661_, new_n797_, new_n232_, new_n724_, new_n1070_, new_n1109_, new_n672_, new_n1269_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n604_, new_n1104_, new_n571_, new_n758_, new_n328_, new_n460_, new_n1267_, new_n268_, new_n1299_, new_n380_, new_n1079_, new_n861_, new_n1252_, new_n352_, new_n931_, new_n575_, new_n562_, new_n944_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n963_, new_n586_, new_n1325_, new_n993_, new_n1191_, new_n824_, new_n717_, new_n403_, new_n475_, new_n868_, new_n1242_, new_n858_, new_n1343_, new_n936_, new_n411_, new_n1016_, new_n673_, new_n1144_, new_n407_, new_n666_, new_n1290_, new_n736_, new_n879_, new_n513_, new_n558_, new_n219_, new_n313_, new_n382_, new_n239_, new_n718_, new_n1310_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n1040_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n255_, new_n533_, new_n1130_, new_n795_, new_n459_, new_n1122_, new_n1185_, new_n1240_, new_n1174_, new_n968_, new_n613_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n591_, new_n837_, new_n801_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1334_, new_n531_, new_n593_, new_n974_, new_n252_, new_n1248_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n470_, new_n769_, new_n433_, new_n871_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n1052_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1220_, new_n989_, new_n1117_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n1276_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n818_, new_n881_, new_n1268_, new_n640_, new_n684_, new_n1274_, new_n754_, new_n653_, new_n377_, new_n905_, new_n1258_, new_n375_, new_n962_, new_n760_, new_n627_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n1339_, new_n320_, new_n780_, new_n984_, new_n1183_, new_n643_, new_n1194_, new_n1316_, new_n1338_, new_n1230_, new_n1027_, new_n348_, new_n610_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1259_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n709_, new_n373_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n770_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n889_, new_n536_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n1249_, new_n955_, new_n847_, new_n250_, new_n888_, new_n288_, new_n1340_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n827_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1207_, new_n1176_, new_n601_, new_n842_, new_n1057_, new_n682_, new_n1075_, new_n812_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n1342_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n413_, new_n442_, new_n642_, new_n462_, new_n603_, new_n564_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n799_, new_n1304_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n1264_, new_n215_, new_n1319_, new_n626_, new_n959_, new_n990_, new_n716_, new_n701_, new_n1238_, new_n1058_, new_n1162_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n414_, new_n1101_, new_n1250_, new_n315_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n281_, new_n430_, new_n844_, new_n482_, new_n1302_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n1297_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n906_, new_n361_, new_n764_, new_n683_, new_n463_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n1292_, new_n517_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1051_, new_n899_, new_n1053_, new_n492_, new_n1200_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1219_, new_n920_, new_n1121_, new_n1341_, new_n820_, new_n771_, new_n979_, new_n508_, new_n714_, new_n1280_, new_n1007_, new_n1241_, new_n882_, new_n1145_, new_n929_, new_n986_, new_n314_, new_n1159_, new_n1337_, new_n216_, new_n917_, new_n1322_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n447_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n465_, new_n739_, new_n783_, new_n341_, new_n996_, new_n1318_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n848_, new_n277_, new_n1245_, new_n663_, new_n579_, new_n286_, new_n1254_, new_n438_, new_n939_, new_n632_, new_n1335_, new_n671_, new_n965_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n397_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n948_, new_n1231_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1301_, new_n1128_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1161_, new_n1329_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n784_, new_n1273_, new_n258_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n693_, new_n1272_, new_n1287_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1289_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n578_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1001_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n231_, new_n583_, new_n617_, new_n1080_, new_n1279_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n1155_, new_n1186_, new_n1261_, new_n225_, new_n1246_, new_n922_, new_n387_, new_n476_, new_n987_, new_n949_, new_n221_, new_n243_, new_n450_, new_n1179_, new_n298_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n623_, new_n446_, new_n316_, new_n590_, new_n826_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n307_, new_n1181_, new_n597_, new_n1093_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1296_, new_n435_, new_n1309_, new_n1010_, new_n776_, new_n687_, new_n370_, new_n1029_, new_n638_, new_n523_, new_n909_, new_n788_, new_n841_, new_n1204_, new_n1112_, new_n711_, new_n1156_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n645_, new_n1096_, new_n1087_, new_n723_, new_n756_, new_n823_, new_n574_, new_n928_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n1291_, new_n247_, new_n539_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n294_, new_n1295_, new_n1173_, new_n704_, new_n1189_, new_n1197_, new_n1312_, new_n474_, new_n1223_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1243_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n947_, new_n994_, new_n982_, new_n964_, new_n1078_, new_n551_, new_n279_, new_n455_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n573_, new_n765_, new_n1314_, new_n1103_;

not g0000 ( new_n215_, N75 );
nand g0001 ( new_n216_, N29, N42 );
nor g0002 ( N388, new_n216_, new_n215_ );
not g0003 ( new_n218_, N80 );
nand g0004 ( new_n219_, N29, N36 );
nor g0005 ( N389, new_n219_, new_n218_ );
not g0006 ( new_n221_, N42 );
nor g0007 ( N390, new_n219_, new_n221_ );
nand g0008 ( new_n223_, N85, N86 );
not g0009 ( N391, new_n223_ );
not g0010 ( new_n225_, N17 );
nand g0011 ( new_n226_, N1, N8 );
not g0012 ( new_n227_, new_n226_ );
nand g0013 ( new_n228_, new_n227_, N13 );
nor g0014 ( N418, new_n228_, new_n225_ );
not g0015 ( new_n230_, N390 );
nand g0016 ( new_n231_, N1, N26 );
nand g0017 ( new_n232_, N13, N17 );
nor g0018 ( new_n233_, new_n231_, new_n232_ );
nand g0019 ( N419, new_n230_, new_n233_ );
nand g0020 ( new_n235_, N59, N75 );
not g0021 ( new_n236_, new_n235_ );
nand g0022 ( N420, new_n236_, N80 );
nand g0023 ( new_n238_, N36, N59 );
not g0024 ( new_n239_, new_n238_ );
nand g0025 ( N421, new_n239_, N80 );
nand g0026 ( N422, new_n239_, N42 );
not g0027 ( new_n242_, N90 );
nor g0028 ( new_n243_, N87, N88 );
nor g0029 ( N423, new_n243_, new_n242_ );
nand g0030 ( N446, new_n233_, N390 );
not g0031 ( new_n246_, keyIn_0_0 );
not g0032 ( new_n247_, new_n231_ );
nand g0033 ( new_n248_, new_n247_, N51 );
nor g0034 ( new_n249_, new_n248_, new_n246_ );
not g0035 ( new_n250_, N51 );
nor g0036 ( new_n251_, new_n231_, new_n250_ );
nor g0037 ( new_n252_, new_n251_, keyIn_0_0 );
nor g0038 ( N447, new_n249_, new_n252_ );
not g0039 ( new_n254_, new_n228_ );
nand g0040 ( new_n255_, new_n254_, N55 );
nand g0041 ( new_n256_, N29, N68 );
nor g0042 ( N448, new_n255_, new_n256_ );
nand g0043 ( new_n258_, N59, N68 );
not g0044 ( new_n259_, new_n258_ );
nand g0045 ( new_n260_, new_n259_, N74 );
nor g0046 ( N449, new_n255_, new_n260_ );
not g0047 ( new_n262_, N89 );
nor g0048 ( N450, new_n243_, new_n262_ );
not g0049 ( new_n264_, N130 );
not g0050 ( new_n265_, keyIn_0_23 );
nand g0051 ( new_n266_, N91, N96 );
nor g0052 ( new_n267_, N91, N96 );
nor g0053 ( new_n268_, new_n267_, keyIn_0_12 );
nand g0054 ( new_n269_, new_n268_, new_n266_ );
not g0055 ( new_n270_, new_n269_ );
not g0056 ( new_n271_, keyIn_0_12 );
not g0057 ( new_n272_, new_n266_ );
nor g0058 ( new_n273_, new_n272_, new_n267_ );
nor g0059 ( new_n274_, new_n273_, new_n271_ );
nor g0060 ( new_n275_, new_n270_, new_n274_ );
not g0061 ( new_n276_, new_n275_ );
not g0062 ( new_n277_, N101 );
nor g0063 ( new_n278_, new_n277_, N106 );
nand g0064 ( new_n279_, new_n277_, N106 );
not g0065 ( new_n280_, new_n279_ );
nor g0066 ( new_n281_, new_n280_, new_n278_ );
not g0067 ( new_n282_, new_n281_ );
nand g0068 ( new_n283_, new_n282_, keyIn_0_13 );
not g0069 ( new_n284_, new_n283_ );
nor g0070 ( new_n285_, new_n282_, keyIn_0_13 );
nor g0071 ( new_n286_, new_n284_, new_n285_ );
nor g0072 ( new_n287_, new_n286_, new_n276_ );
not g0073 ( new_n288_, new_n287_ );
nand g0074 ( new_n289_, new_n288_, new_n265_ );
nand g0075 ( new_n290_, new_n287_, keyIn_0_23 );
nand g0076 ( new_n291_, new_n289_, new_n290_ );
not g0077 ( new_n292_, keyIn_0_28 );
nand g0078 ( new_n293_, new_n286_, new_n276_ );
nand g0079 ( new_n294_, new_n293_, new_n292_ );
not g0080 ( new_n295_, new_n293_ );
nand g0081 ( new_n296_, new_n295_, keyIn_0_28 );
nand g0082 ( new_n297_, new_n296_, new_n294_ );
nand g0083 ( new_n298_, new_n291_, new_n297_ );
nand g0084 ( new_n299_, new_n298_, keyIn_0_37 );
not g0085 ( new_n300_, new_n299_ );
nor g0086 ( new_n301_, new_n298_, keyIn_0_37 );
nor g0087 ( new_n302_, new_n300_, new_n301_ );
nor g0088 ( new_n303_, new_n302_, new_n264_ );
nand g0089 ( new_n304_, new_n302_, new_n264_ );
not g0090 ( new_n305_, new_n304_ );
nor g0091 ( new_n306_, new_n305_, new_n303_ );
not g0092 ( new_n307_, N135 );
not g0093 ( new_n308_, N111 );
nor g0094 ( new_n309_, new_n308_, N116 );
nand g0095 ( new_n310_, new_n308_, N116 );
not g0096 ( new_n311_, new_n310_ );
nor g0097 ( new_n312_, new_n311_, new_n309_ );
not g0098 ( new_n313_, new_n312_ );
nand g0099 ( new_n314_, new_n313_, keyIn_0_14 );
not g0100 ( new_n315_, new_n314_ );
nor g0101 ( new_n316_, new_n313_, keyIn_0_14 );
nor g0102 ( new_n317_, new_n315_, new_n316_ );
nand g0103 ( new_n318_, N121, N126 );
nor g0104 ( new_n319_, N121, N126 );
nor g0105 ( new_n320_, new_n319_, keyIn_0_15 );
nand g0106 ( new_n321_, new_n320_, new_n318_ );
not g0107 ( new_n322_, new_n321_ );
not g0108 ( new_n323_, keyIn_0_15 );
not g0109 ( new_n324_, new_n318_ );
nor g0110 ( new_n325_, new_n324_, new_n319_ );
nor g0111 ( new_n326_, new_n325_, new_n323_ );
nor g0112 ( new_n327_, new_n322_, new_n326_ );
not g0113 ( new_n328_, new_n327_ );
nor g0114 ( new_n329_, new_n317_, new_n328_ );
not g0115 ( new_n330_, new_n329_ );
nand g0116 ( new_n331_, new_n330_, keyIn_0_24 );
not g0117 ( new_n332_, keyIn_0_24 );
nand g0118 ( new_n333_, new_n329_, new_n332_ );
nand g0119 ( new_n334_, new_n331_, new_n333_ );
nand g0120 ( new_n335_, new_n317_, new_n328_ );
nand g0121 ( new_n336_, new_n335_, keyIn_0_29 );
not g0122 ( new_n337_, keyIn_0_29 );
not g0123 ( new_n338_, new_n335_ );
nand g0124 ( new_n339_, new_n338_, new_n337_ );
nand g0125 ( new_n340_, new_n339_, new_n336_ );
nand g0126 ( new_n341_, new_n334_, new_n340_ );
nand g0127 ( new_n342_, new_n341_, keyIn_0_38 );
not g0128 ( new_n343_, new_n342_ );
nor g0129 ( new_n344_, new_n341_, keyIn_0_38 );
nor g0130 ( new_n345_, new_n343_, new_n344_ );
nor g0131 ( new_n346_, new_n345_, new_n307_ );
nand g0132 ( new_n347_, new_n345_, new_n307_ );
not g0133 ( new_n348_, new_n347_ );
nor g0134 ( new_n349_, new_n348_, new_n346_ );
nand g0135 ( new_n350_, new_n306_, new_n349_ );
not g0136 ( new_n351_, new_n306_ );
not g0137 ( new_n352_, new_n349_ );
nand g0138 ( new_n353_, new_n351_, new_n352_ );
nand g0139 ( N767, new_n353_, new_n350_ );
not g0140 ( new_n355_, N207 );
not g0141 ( new_n356_, N195 );
nor g0142 ( new_n357_, new_n356_, N201 );
not g0143 ( new_n358_, N201 );
nor g0144 ( new_n359_, new_n358_, N195 );
nor g0145 ( new_n360_, new_n357_, new_n359_ );
not g0146 ( new_n361_, new_n360_ );
nand g0147 ( new_n362_, new_n361_, keyIn_0_21 );
not g0148 ( new_n363_, new_n362_ );
nor g0149 ( new_n364_, new_n361_, keyIn_0_21 );
nor g0150 ( new_n365_, new_n363_, new_n364_ );
nor g0151 ( new_n366_, N183, N189 );
nand g0152 ( new_n367_, N183, N189 );
not g0153 ( new_n368_, new_n367_ );
nor g0154 ( new_n369_, new_n368_, new_n366_ );
not g0155 ( new_n370_, new_n369_ );
nor g0156 ( new_n371_, new_n370_, keyIn_0_20 );
nand g0157 ( new_n372_, new_n370_, keyIn_0_20 );
not g0158 ( new_n373_, new_n372_ );
nor g0159 ( new_n374_, new_n373_, new_n371_ );
nor g0160 ( new_n375_, new_n365_, new_n374_ );
not g0161 ( new_n376_, new_n375_ );
nand g0162 ( new_n377_, new_n376_, keyIn_0_27 );
not g0163 ( new_n378_, new_n377_ );
nor g0164 ( new_n379_, new_n376_, keyIn_0_27 );
nor g0165 ( new_n380_, new_n378_, new_n379_ );
nand g0166 ( new_n381_, new_n365_, new_n374_ );
not g0167 ( new_n382_, new_n381_ );
nor g0168 ( new_n383_, new_n382_, keyIn_0_36 );
nand g0169 ( new_n384_, new_n382_, keyIn_0_36 );
not g0170 ( new_n385_, new_n384_ );
nor g0171 ( new_n386_, new_n385_, new_n383_ );
nor g0172 ( new_n387_, new_n380_, new_n386_ );
not g0173 ( new_n388_, new_n387_ );
nand g0174 ( new_n389_, new_n388_, keyIn_0_50 );
not g0175 ( new_n390_, new_n389_ );
nor g0176 ( new_n391_, new_n388_, keyIn_0_50 );
nor g0177 ( new_n392_, new_n390_, new_n391_ );
nor g0178 ( new_n393_, new_n392_, new_n355_ );
nand g0179 ( new_n394_, new_n392_, new_n355_ );
not g0180 ( new_n395_, new_n394_ );
nor g0181 ( new_n396_, new_n395_, new_n393_ );
not g0182 ( new_n397_, new_n396_ );
not g0183 ( new_n398_, keyIn_0_26 );
nor g0184 ( new_n399_, N171, N177 );
nand g0185 ( new_n400_, N171, N177 );
not g0186 ( new_n401_, new_n400_ );
nor g0187 ( new_n402_, new_n401_, new_n399_ );
not g0188 ( new_n403_, new_n402_ );
nor g0189 ( new_n404_, new_n403_, keyIn_0_19 );
nand g0190 ( new_n405_, new_n403_, keyIn_0_19 );
not g0191 ( new_n406_, new_n405_ );
nor g0192 ( new_n407_, new_n406_, new_n404_ );
not g0193 ( new_n408_, new_n407_ );
not g0194 ( new_n409_, N159 );
nor g0195 ( new_n410_, new_n409_, N165 );
not g0196 ( new_n411_, N165 );
nor g0197 ( new_n412_, new_n411_, N159 );
nor g0198 ( new_n413_, new_n410_, new_n412_ );
not g0199 ( new_n414_, new_n413_ );
nand g0200 ( new_n415_, new_n414_, keyIn_0_18 );
not g0201 ( new_n416_, new_n415_ );
nor g0202 ( new_n417_, new_n414_, keyIn_0_18 );
nor g0203 ( new_n418_, new_n416_, new_n417_ );
not g0204 ( new_n419_, new_n418_ );
nor g0205 ( new_n420_, new_n419_, new_n408_ );
nor g0206 ( new_n421_, new_n420_, new_n398_ );
nor g0207 ( new_n422_, new_n418_, new_n407_ );
not g0208 ( new_n423_, new_n422_ );
nand g0209 ( new_n424_, new_n423_, keyIn_0_35 );
not g0210 ( new_n425_, new_n424_ );
nor g0211 ( new_n426_, new_n425_, new_n421_ );
nand g0212 ( new_n427_, new_n420_, new_n398_ );
not g0213 ( new_n428_, new_n427_ );
nor g0214 ( new_n429_, new_n423_, keyIn_0_35 );
nor g0215 ( new_n430_, new_n428_, new_n429_ );
nand g0216 ( new_n431_, new_n426_, new_n430_ );
not g0217 ( new_n432_, new_n431_ );
nor g0218 ( new_n433_, new_n432_, keyIn_0_49 );
nand g0219 ( new_n434_, new_n432_, keyIn_0_49 );
not g0220 ( new_n435_, new_n434_ );
nor g0221 ( new_n436_, new_n435_, new_n433_ );
not g0222 ( new_n437_, new_n436_ );
nand g0223 ( new_n438_, new_n437_, N130 );
not g0224 ( new_n439_, new_n438_ );
nor g0225 ( new_n440_, new_n437_, N130 );
nor g0226 ( new_n441_, new_n439_, new_n440_ );
not g0227 ( new_n442_, new_n441_ );
nand g0228 ( new_n443_, new_n442_, new_n397_ );
nand g0229 ( new_n444_, new_n441_, new_n396_ );
nand g0230 ( N768, new_n443_, new_n444_ );
not g0231 ( new_n446_, keyIn_0_112 );
not g0232 ( new_n447_, N261 );
not g0233 ( new_n448_, keyIn_0_94 );
not g0234 ( new_n449_, keyIn_0_78 );
not g0235 ( new_n450_, keyIn_0_70 );
not g0236 ( new_n451_, keyIn_0_34 );
nand g0237 ( new_n452_, new_n251_, keyIn_0_0 );
nand g0238 ( new_n453_, new_n248_, new_n246_ );
nand g0239 ( new_n454_, new_n453_, new_n452_ );
nand g0240 ( new_n455_, new_n454_, keyIn_0_8 );
not g0241 ( new_n456_, keyIn_0_8 );
nand g0242 ( new_n457_, N447, new_n456_ );
nand g0243 ( new_n458_, new_n457_, new_n455_ );
nand g0244 ( new_n459_, new_n458_, keyIn_0_22 );
not g0245 ( new_n460_, keyIn_0_22 );
nor g0246 ( new_n461_, N447, new_n456_ );
nor g0247 ( new_n462_, new_n454_, keyIn_0_8 );
nor g0248 ( new_n463_, new_n461_, new_n462_ );
nand g0249 ( new_n464_, new_n463_, new_n460_ );
nand g0250 ( new_n465_, new_n464_, new_n459_ );
nand g0251 ( new_n466_, N59, N156 );
nand g0252 ( new_n467_, new_n466_, keyIn_0_5 );
not g0253 ( new_n468_, new_n467_ );
nor g0254 ( new_n469_, new_n466_, keyIn_0_5 );
nor g0255 ( new_n470_, new_n468_, new_n469_ );
nor g0256 ( new_n471_, new_n470_, new_n225_ );
not g0257 ( new_n472_, new_n471_ );
nor g0258 ( new_n473_, new_n465_, new_n472_ );
nand g0259 ( new_n474_, new_n473_, new_n451_ );
nor g0260 ( new_n475_, new_n463_, new_n460_ );
nor g0261 ( new_n476_, new_n458_, keyIn_0_22 );
nor g0262 ( new_n477_, new_n475_, new_n476_ );
nand g0263 ( new_n478_, new_n477_, new_n471_ );
nand g0264 ( new_n479_, new_n478_, keyIn_0_34 );
nand g0265 ( new_n480_, new_n479_, new_n474_ );
nand g0266 ( new_n481_, new_n480_, N1 );
not g0267 ( new_n482_, new_n481_ );
nand g0268 ( new_n483_, new_n482_, keyIn_0_44 );
not g0269 ( new_n484_, keyIn_0_44 );
nand g0270 ( new_n485_, new_n481_, new_n484_ );
nand g0271 ( new_n486_, new_n483_, new_n485_ );
nand g0272 ( new_n487_, new_n486_, N153 );
nand g0273 ( new_n488_, new_n487_, keyIn_0_61 );
not g0274 ( new_n489_, keyIn_0_39 );
not g0275 ( new_n490_, keyIn_0_33 );
not g0276 ( new_n491_, keyIn_0_17 );
nor g0277 ( new_n492_, N17, N42 );
nor g0278 ( new_n493_, new_n492_, keyIn_0_6 );
not g0279 ( new_n494_, new_n493_ );
nand g0280 ( new_n495_, new_n492_, keyIn_0_6 );
nand g0281 ( new_n496_, new_n494_, new_n495_ );
nand g0282 ( new_n497_, N17, N42 );
nor g0283 ( new_n498_, new_n497_, keyIn_0_7 );
not g0284 ( new_n499_, new_n498_ );
nand g0285 ( new_n500_, new_n497_, keyIn_0_7 );
nand g0286 ( new_n501_, new_n499_, new_n500_ );
nor g0287 ( new_n502_, new_n496_, new_n501_ );
not g0288 ( new_n503_, new_n502_ );
nor g0289 ( new_n504_, new_n503_, new_n491_ );
not g0290 ( new_n505_, new_n504_ );
nor g0291 ( new_n506_, new_n502_, keyIn_0_17 );
nor g0292 ( new_n507_, new_n506_, new_n466_ );
nand g0293 ( new_n508_, new_n505_, new_n507_ );
not g0294 ( new_n509_, new_n508_ );
nand g0295 ( new_n510_, new_n477_, new_n509_ );
nor g0296 ( new_n511_, new_n510_, new_n490_ );
nand g0297 ( new_n512_, new_n510_, new_n490_ );
not g0298 ( new_n513_, keyIn_0_1 );
nand g0299 ( new_n514_, N17, N51 );
nor g0300 ( new_n515_, new_n226_, new_n514_ );
nand g0301 ( new_n516_, new_n515_, new_n513_ );
nor g0302 ( new_n517_, new_n515_, new_n513_ );
not g0303 ( new_n518_, new_n517_ );
nand g0304 ( new_n519_, new_n518_, new_n516_ );
nand g0305 ( new_n520_, new_n519_, keyIn_0_9 );
not g0306 ( new_n521_, keyIn_0_9 );
not g0307 ( new_n522_, new_n516_ );
nor g0308 ( new_n523_, new_n522_, new_n517_ );
nand g0309 ( new_n524_, new_n523_, new_n521_ );
nand g0310 ( new_n525_, new_n524_, new_n520_ );
not g0311 ( new_n526_, keyIn_0_11 );
nand g0312 ( new_n527_, N42, N59 );
nor g0313 ( new_n528_, new_n527_, new_n215_ );
nand g0314 ( new_n529_, new_n528_, keyIn_0_3 );
nor g0315 ( new_n530_, new_n528_, keyIn_0_3 );
not g0316 ( new_n531_, new_n530_ );
nand g0317 ( new_n532_, new_n531_, new_n529_ );
nand g0318 ( new_n533_, new_n532_, new_n526_ );
not g0319 ( new_n534_, new_n532_ );
nand g0320 ( new_n535_, new_n534_, keyIn_0_11 );
nand g0321 ( new_n536_, new_n535_, new_n533_ );
nand g0322 ( new_n537_, new_n536_, new_n525_ );
nand g0323 ( new_n538_, new_n537_, keyIn_0_25 );
not g0324 ( new_n539_, new_n538_ );
nor g0325 ( new_n540_, new_n537_, keyIn_0_25 );
nor g0326 ( new_n541_, new_n539_, new_n540_ );
nand g0327 ( new_n542_, new_n512_, new_n541_ );
nor g0328 ( new_n543_, new_n542_, new_n511_ );
nand g0329 ( new_n544_, new_n543_, new_n489_ );
not g0330 ( new_n545_, new_n511_ );
nor g0331 ( new_n546_, new_n465_, new_n508_ );
nor g0332 ( new_n547_, new_n546_, keyIn_0_33 );
not g0333 ( new_n548_, keyIn_0_25 );
not g0334 ( new_n549_, new_n537_ );
nand g0335 ( new_n550_, new_n549_, new_n548_ );
nand g0336 ( new_n551_, new_n550_, new_n538_ );
nor g0337 ( new_n552_, new_n547_, new_n551_ );
nand g0338 ( new_n553_, new_n552_, new_n545_ );
nand g0339 ( new_n554_, new_n553_, keyIn_0_39 );
nand g0340 ( new_n555_, new_n544_, new_n554_ );
nand g0341 ( new_n556_, new_n555_, N126 );
nand g0342 ( new_n557_, new_n556_, keyIn_0_62 );
nand g0343 ( new_n558_, new_n488_, new_n557_ );
not g0344 ( new_n559_, keyIn_0_61 );
not g0345 ( new_n560_, N153 );
nor g0346 ( new_n561_, new_n481_, new_n484_ );
not g0347 ( new_n562_, new_n485_ );
nor g0348 ( new_n563_, new_n562_, new_n561_ );
nor g0349 ( new_n564_, new_n563_, new_n560_ );
nand g0350 ( new_n565_, new_n564_, new_n559_ );
not g0351 ( new_n566_, keyIn_0_62 );
not g0352 ( new_n567_, new_n556_ );
nand g0353 ( new_n568_, new_n567_, new_n566_ );
nand g0354 ( new_n569_, new_n565_, new_n568_ );
nor g0355 ( new_n570_, new_n569_, new_n558_ );
nand g0356 ( new_n571_, new_n570_, new_n450_ );
not g0357 ( new_n572_, new_n558_ );
nor g0358 ( new_n573_, new_n487_, keyIn_0_61 );
nor g0359 ( new_n574_, new_n556_, keyIn_0_62 );
nor g0360 ( new_n575_, new_n573_, new_n574_ );
nand g0361 ( new_n576_, new_n572_, new_n575_ );
nand g0362 ( new_n577_, new_n576_, keyIn_0_70 );
nand g0363 ( new_n578_, new_n577_, new_n571_ );
not g0364 ( new_n579_, keyIn_0_48 );
not g0365 ( new_n580_, N55 );
not g0366 ( new_n581_, keyIn_0_2 );
nand g0367 ( new_n582_, N29, N75 );
nor g0368 ( new_n583_, new_n582_, new_n218_ );
not g0369 ( new_n584_, new_n583_ );
nor g0370 ( new_n585_, new_n584_, new_n581_ );
nor g0371 ( new_n586_, new_n583_, keyIn_0_2 );
nor g0372 ( new_n587_, new_n585_, new_n586_ );
nor g0373 ( new_n588_, new_n465_, new_n587_ );
not g0374 ( new_n589_, new_n588_ );
nor g0375 ( new_n590_, new_n589_, new_n580_ );
not g0376 ( new_n591_, new_n590_ );
nand g0377 ( new_n592_, new_n591_, keyIn_0_32 );
not g0378 ( new_n593_, keyIn_0_32 );
nand g0379 ( new_n594_, new_n590_, new_n593_ );
nand g0380 ( new_n595_, new_n592_, new_n594_ );
not g0381 ( new_n596_, N268 );
nor g0382 ( new_n597_, new_n596_, keyIn_0_4 );
nand g0383 ( new_n598_, new_n596_, keyIn_0_4 );
not g0384 ( new_n599_, new_n598_ );
nor g0385 ( new_n600_, new_n599_, new_n597_ );
not g0386 ( new_n601_, new_n600_ );
nand g0387 ( new_n602_, new_n601_, keyIn_0_16 );
not g0388 ( new_n603_, new_n602_ );
nor g0389 ( new_n604_, new_n601_, keyIn_0_16 );
nor g0390 ( new_n605_, new_n603_, new_n604_ );
not g0391 ( new_n606_, new_n605_ );
nand g0392 ( new_n607_, new_n595_, new_n606_ );
not g0393 ( new_n608_, new_n607_ );
nand g0394 ( new_n609_, new_n608_, new_n579_ );
nand g0395 ( new_n610_, new_n607_, keyIn_0_48 );
nand g0396 ( new_n611_, new_n609_, new_n610_ );
nand g0397 ( new_n612_, new_n578_, new_n611_ );
nor g0398 ( new_n613_, new_n612_, new_n449_ );
nand g0399 ( new_n614_, new_n612_, new_n449_ );
not g0400 ( new_n615_, new_n614_ );
nor g0401 ( new_n616_, new_n615_, new_n613_ );
nand g0402 ( new_n617_, new_n616_, N201 );
nor g0403 ( new_n618_, new_n617_, keyIn_0_83 );
nand g0404 ( new_n619_, new_n617_, keyIn_0_83 );
not g0405 ( new_n620_, new_n619_ );
nor g0406 ( new_n621_, new_n620_, new_n618_ );
nor g0407 ( new_n622_, new_n616_, N201 );
nand g0408 ( new_n623_, new_n622_, keyIn_0_84 );
not g0409 ( new_n624_, keyIn_0_84 );
not g0410 ( new_n625_, new_n613_ );
nand g0411 ( new_n626_, new_n625_, new_n614_ );
nand g0412 ( new_n627_, new_n626_, new_n358_ );
nand g0413 ( new_n628_, new_n627_, new_n624_ );
nand g0414 ( new_n629_, new_n623_, new_n628_ );
nor g0415 ( new_n630_, new_n621_, new_n629_ );
nor g0416 ( new_n631_, new_n630_, new_n448_ );
nand g0417 ( new_n632_, new_n630_, new_n448_ );
not g0418 ( new_n633_, new_n632_ );
nor g0419 ( new_n634_, new_n633_, new_n631_ );
not g0420 ( new_n635_, new_n634_ );
nor g0421 ( new_n636_, new_n635_, new_n447_ );
nand g0422 ( new_n637_, new_n635_, new_n447_ );
nand g0423 ( new_n638_, new_n637_, N219 );
nor g0424 ( new_n639_, new_n638_, new_n636_ );
not g0425 ( new_n640_, N228 );
nor g0426 ( new_n641_, new_n635_, new_n640_ );
not g0427 ( new_n642_, keyIn_0_93 );
not g0428 ( new_n643_, keyIn_0_83 );
not g0429 ( new_n644_, new_n617_ );
nand g0430 ( new_n645_, new_n644_, new_n643_ );
nand g0431 ( new_n646_, new_n645_, new_n619_ );
nand g0432 ( new_n647_, new_n646_, new_n642_ );
nand g0433 ( new_n648_, new_n621_, keyIn_0_93 );
nand g0434 ( new_n649_, new_n648_, new_n647_ );
nand g0435 ( new_n650_, new_n649_, N237 );
not g0436 ( new_n651_, N246 );
nor g0437 ( new_n652_, new_n626_, new_n651_ );
not g0438 ( new_n653_, keyIn_0_10 );
not g0439 ( new_n654_, new_n527_ );
nand g0440 ( new_n655_, N68, N72 );
not g0441 ( new_n656_, new_n655_ );
nand g0442 ( new_n657_, new_n654_, new_n656_ );
nor g0443 ( new_n658_, new_n255_, new_n657_ );
nor g0444 ( new_n659_, new_n658_, new_n653_ );
nand g0445 ( new_n660_, new_n658_, new_n653_ );
nand g0446 ( new_n661_, new_n660_, N73 );
nor g0447 ( new_n662_, new_n661_, new_n659_ );
nand g0448 ( new_n663_, new_n662_, N201 );
nand g0449 ( new_n664_, N121, N210 );
nand g0450 ( new_n665_, N255, N267 );
nand g0451 ( new_n666_, new_n664_, new_n665_ );
not g0452 ( new_n667_, new_n666_ );
nand g0453 ( new_n668_, new_n663_, new_n667_ );
nor g0454 ( new_n669_, new_n652_, new_n668_ );
nand g0455 ( new_n670_, new_n650_, new_n669_ );
nor g0456 ( new_n671_, new_n641_, new_n670_ );
not g0457 ( new_n672_, new_n671_ );
nor g0458 ( new_n673_, new_n639_, new_n672_ );
not g0459 ( new_n674_, new_n673_ );
nand g0460 ( new_n675_, new_n674_, new_n446_ );
nand g0461 ( new_n676_, new_n673_, keyIn_0_112 );
nand g0462 ( N850, new_n675_, new_n676_ );
not g0463 ( new_n678_, keyIn_0_106 );
not g0464 ( new_n679_, keyIn_0_103 );
not g0465 ( new_n680_, keyIn_0_99 );
not g0466 ( new_n681_, keyIn_0_68 );
nand g0467 ( new_n682_, new_n486_, N146 );
nand g0468 ( new_n683_, new_n682_, keyIn_0_57 );
not g0469 ( new_n684_, keyIn_0_58 );
nand g0470 ( new_n685_, new_n555_, N116 );
nand g0471 ( new_n686_, new_n685_, new_n684_ );
nand g0472 ( new_n687_, new_n683_, new_n686_ );
not g0473 ( new_n688_, new_n687_ );
nor g0474 ( new_n689_, new_n682_, keyIn_0_57 );
nor g0475 ( new_n690_, new_n685_, new_n684_ );
nor g0476 ( new_n691_, new_n689_, new_n690_ );
nand g0477 ( new_n692_, new_n688_, new_n691_ );
nor g0478 ( new_n693_, new_n692_, new_n681_ );
not g0479 ( new_n694_, new_n693_ );
not g0480 ( new_n695_, keyIn_0_57 );
not g0481 ( new_n696_, N146 );
nor g0482 ( new_n697_, new_n563_, new_n696_ );
nand g0483 ( new_n698_, new_n697_, new_n695_ );
not g0484 ( new_n699_, new_n685_ );
nand g0485 ( new_n700_, new_n699_, keyIn_0_58 );
nand g0486 ( new_n701_, new_n698_, new_n700_ );
nor g0487 ( new_n702_, new_n701_, new_n687_ );
nor g0488 ( new_n703_, new_n702_, keyIn_0_68 );
not g0489 ( new_n704_, keyIn_0_46 );
nor g0490 ( new_n705_, new_n607_, new_n704_ );
not g0491 ( new_n706_, new_n705_ );
nand g0492 ( new_n707_, new_n607_, new_n704_ );
nand g0493 ( new_n708_, new_n706_, new_n707_ );
not g0494 ( new_n709_, new_n708_ );
nor g0495 ( new_n710_, new_n703_, new_n709_ );
nand g0496 ( new_n711_, new_n710_, new_n694_ );
nand g0497 ( new_n712_, new_n711_, keyIn_0_76 );
not g0498 ( new_n713_, keyIn_0_76 );
nand g0499 ( new_n714_, new_n692_, new_n681_ );
nand g0500 ( new_n715_, new_n714_, new_n708_ );
nor g0501 ( new_n716_, new_n715_, new_n693_ );
nand g0502 ( new_n717_, new_n716_, new_n713_ );
nand g0503 ( new_n718_, new_n712_, new_n717_ );
nor g0504 ( new_n719_, new_n718_, N189 );
nand g0505 ( new_n720_, new_n719_, keyIn_0_80 );
not g0506 ( new_n721_, keyIn_0_80 );
not g0507 ( new_n722_, N189 );
nor g0508 ( new_n723_, new_n716_, new_n713_ );
nor g0509 ( new_n724_, new_n711_, keyIn_0_76 );
nor g0510 ( new_n725_, new_n724_, new_n723_ );
nand g0511 ( new_n726_, new_n725_, new_n722_ );
nand g0512 ( new_n727_, new_n726_, new_n721_ );
nand g0513 ( new_n728_, new_n727_, new_n720_ );
not g0514 ( new_n729_, keyIn_0_82 );
not g0515 ( new_n730_, keyIn_0_60 );
nand g0516 ( new_n731_, new_n555_, N121 );
not g0517 ( new_n732_, new_n731_ );
nand g0518 ( new_n733_, new_n732_, new_n730_ );
nand g0519 ( new_n734_, new_n731_, keyIn_0_60 );
nand g0520 ( new_n735_, new_n733_, new_n734_ );
not g0521 ( new_n736_, keyIn_0_59 );
not g0522 ( new_n737_, N149 );
nor g0523 ( new_n738_, new_n563_, new_n737_ );
nand g0524 ( new_n739_, new_n738_, new_n736_ );
nand g0525 ( new_n740_, new_n486_, N149 );
nand g0526 ( new_n741_, new_n740_, keyIn_0_59 );
nand g0527 ( new_n742_, new_n739_, new_n741_ );
nand g0528 ( new_n743_, new_n742_, new_n735_ );
nor g0529 ( new_n744_, new_n743_, keyIn_0_69 );
not g0530 ( new_n745_, new_n744_ );
nand g0531 ( new_n746_, new_n743_, keyIn_0_69 );
nor g0532 ( new_n747_, new_n607_, keyIn_0_47 );
nand g0533 ( new_n748_, new_n607_, keyIn_0_47 );
not g0534 ( new_n749_, new_n748_ );
nor g0535 ( new_n750_, new_n749_, new_n747_ );
nand g0536 ( new_n751_, new_n746_, new_n750_ );
not g0537 ( new_n752_, new_n751_ );
nand g0538 ( new_n753_, new_n752_, new_n745_ );
nand g0539 ( new_n754_, new_n753_, keyIn_0_77 );
not g0540 ( new_n755_, keyIn_0_77 );
nor g0541 ( new_n756_, new_n751_, new_n744_ );
nand g0542 ( new_n757_, new_n756_, new_n755_ );
nand g0543 ( new_n758_, new_n754_, new_n757_ );
nor g0544 ( new_n759_, new_n758_, N195 );
nand g0545 ( new_n760_, new_n759_, new_n729_ );
nor g0546 ( new_n761_, new_n756_, new_n755_ );
not g0547 ( new_n762_, new_n757_ );
nor g0548 ( new_n763_, new_n762_, new_n761_ );
nand g0549 ( new_n764_, new_n763_, new_n356_ );
nand g0550 ( new_n765_, new_n764_, keyIn_0_82 );
nand g0551 ( new_n766_, new_n765_, new_n760_ );
nand g0552 ( new_n767_, new_n766_, new_n728_ );
not g0553 ( new_n768_, new_n767_ );
nand g0554 ( new_n769_, new_n649_, new_n768_ );
nor g0555 ( new_n770_, new_n769_, new_n680_ );
not g0556 ( new_n771_, new_n770_ );
nand g0557 ( new_n772_, new_n769_, new_n680_ );
nand g0558 ( new_n773_, new_n771_, new_n772_ );
not g0559 ( new_n774_, keyIn_0_96 );
nor g0560 ( new_n775_, new_n627_, new_n624_ );
nor g0561 ( new_n776_, new_n622_, keyIn_0_84 );
nor g0562 ( new_n777_, new_n776_, new_n775_ );
nand g0563 ( new_n778_, new_n777_, N261 );
nor g0564 ( new_n779_, new_n778_, new_n767_ );
nand g0565 ( new_n780_, new_n779_, new_n774_ );
nor g0566 ( new_n781_, new_n629_, new_n447_ );
nand g0567 ( new_n782_, new_n768_, new_n781_ );
nand g0568 ( new_n783_, new_n782_, keyIn_0_96 );
nand g0569 ( new_n784_, new_n780_, new_n783_ );
nor g0570 ( new_n785_, new_n725_, new_n722_ );
not g0571 ( new_n786_, new_n785_ );
nand g0572 ( new_n787_, new_n786_, keyIn_0_79 );
not g0573 ( new_n788_, new_n787_ );
nor g0574 ( new_n789_, new_n786_, keyIn_0_79 );
nor g0575 ( new_n790_, new_n788_, new_n789_ );
nand g0576 ( new_n791_, new_n784_, new_n790_ );
not g0577 ( new_n792_, keyIn_0_98 );
not g0578 ( new_n793_, keyIn_0_81 );
nand g0579 ( new_n794_, new_n758_, N195 );
nand g0580 ( new_n795_, new_n794_, new_n793_ );
not g0581 ( new_n796_, new_n795_ );
nor g0582 ( new_n797_, new_n794_, new_n793_ );
nor g0583 ( new_n798_, new_n796_, new_n797_ );
nor g0584 ( new_n799_, new_n798_, keyIn_0_91 );
not g0585 ( new_n800_, keyIn_0_91 );
not g0586 ( new_n801_, new_n794_ );
nand g0587 ( new_n802_, new_n801_, keyIn_0_81 );
nand g0588 ( new_n803_, new_n802_, new_n795_ );
nor g0589 ( new_n804_, new_n803_, new_n800_ );
nor g0590 ( new_n805_, new_n799_, new_n804_ );
nand g0591 ( new_n806_, new_n805_, new_n728_ );
nand g0592 ( new_n807_, new_n806_, new_n792_ );
not g0593 ( new_n808_, new_n728_ );
nand g0594 ( new_n809_, new_n803_, new_n800_ );
nand g0595 ( new_n810_, new_n798_, keyIn_0_91 );
nand g0596 ( new_n811_, new_n810_, new_n809_ );
nor g0597 ( new_n812_, new_n811_, new_n808_ );
nand g0598 ( new_n813_, new_n812_, keyIn_0_98 );
nand g0599 ( new_n814_, new_n807_, new_n813_ );
nor g0600 ( new_n815_, new_n791_, new_n814_ );
nand g0601 ( new_n816_, new_n815_, new_n773_ );
nand g0602 ( new_n817_, new_n816_, new_n679_ );
not g0603 ( new_n818_, new_n772_ );
nor g0604 ( new_n819_, new_n818_, new_n770_ );
not g0605 ( new_n820_, new_n791_ );
nor g0606 ( new_n821_, new_n812_, keyIn_0_98 );
nor g0607 ( new_n822_, new_n806_, new_n792_ );
nor g0608 ( new_n823_, new_n822_, new_n821_ );
nand g0609 ( new_n824_, new_n820_, new_n823_ );
nor g0610 ( new_n825_, new_n824_, new_n819_ );
nand g0611 ( new_n826_, new_n825_, keyIn_0_103 );
nand g0612 ( new_n827_, new_n826_, new_n817_ );
not g0613 ( new_n828_, keyIn_0_89 );
not g0614 ( new_n829_, keyIn_0_75 );
not g0615 ( new_n830_, N143 );
nor g0616 ( new_n831_, new_n563_, new_n830_ );
not g0617 ( new_n832_, new_n831_ );
nand g0618 ( new_n833_, new_n832_, keyIn_0_55 );
not g0619 ( new_n834_, keyIn_0_56 );
nand g0620 ( new_n835_, new_n555_, N111 );
nand g0621 ( new_n836_, new_n835_, new_n834_ );
nand g0622 ( new_n837_, new_n833_, new_n836_ );
nor g0623 ( new_n838_, new_n832_, keyIn_0_55 );
nor g0624 ( new_n839_, new_n835_, new_n834_ );
nor g0625 ( new_n840_, new_n838_, new_n839_ );
not g0626 ( new_n841_, new_n840_ );
nor g0627 ( new_n842_, new_n841_, new_n837_ );
nor g0628 ( new_n843_, new_n842_, keyIn_0_67 );
nand g0629 ( new_n844_, new_n842_, keyIn_0_67 );
not g0630 ( new_n845_, new_n844_ );
nor g0631 ( new_n846_, new_n607_, keyIn_0_45 );
nand g0632 ( new_n847_, new_n607_, keyIn_0_45 );
not g0633 ( new_n848_, new_n847_ );
nor g0634 ( new_n849_, new_n848_, new_n846_ );
nor g0635 ( new_n850_, new_n845_, new_n849_ );
not g0636 ( new_n851_, new_n850_ );
nor g0637 ( new_n852_, new_n851_, new_n843_ );
nor g0638 ( new_n853_, new_n852_, new_n829_ );
nand g0639 ( new_n854_, new_n852_, new_n829_ );
not g0640 ( new_n855_, new_n854_ );
nor g0641 ( new_n856_, new_n855_, new_n853_ );
nor g0642 ( new_n857_, new_n856_, N183 );
nand g0643 ( new_n858_, new_n856_, N183 );
not g0644 ( new_n859_, new_n858_ );
nor g0645 ( new_n860_, new_n859_, new_n857_ );
nor g0646 ( new_n861_, new_n860_, new_n828_ );
nand g0647 ( new_n862_, new_n860_, new_n828_ );
not g0648 ( new_n863_, new_n862_ );
nor g0649 ( new_n864_, new_n863_, new_n861_ );
not g0650 ( new_n865_, new_n864_ );
nor g0651 ( new_n866_, new_n827_, new_n865_ );
not g0652 ( new_n867_, new_n866_ );
nor g0653 ( new_n868_, new_n867_, new_n678_ );
nor g0654 ( new_n869_, new_n866_, keyIn_0_106 );
nand g0655 ( new_n870_, new_n827_, new_n865_ );
nand g0656 ( new_n871_, new_n870_, N219 );
nor g0657 ( new_n872_, new_n869_, new_n871_ );
not g0658 ( new_n873_, new_n872_ );
nor g0659 ( new_n874_, new_n873_, new_n868_ );
nor g0660 ( new_n875_, new_n865_, new_n640_ );
not g0661 ( new_n876_, N237 );
nor g0662 ( new_n877_, new_n858_, new_n876_ );
nand g0663 ( new_n878_, new_n856_, N246 );
not g0664 ( new_n879_, new_n878_ );
nand g0665 ( new_n880_, new_n662_, N183 );
nand g0666 ( new_n881_, N106, N210 );
nand g0667 ( new_n882_, new_n880_, new_n881_ );
nor g0668 ( new_n883_, new_n879_, new_n882_ );
not g0669 ( new_n884_, new_n883_ );
nor g0670 ( new_n885_, new_n884_, new_n877_ );
not g0671 ( new_n886_, new_n885_ );
nor g0672 ( new_n887_, new_n875_, new_n886_ );
not g0673 ( new_n888_, new_n887_ );
nor g0674 ( new_n889_, new_n874_, new_n888_ );
nand g0675 ( new_n890_, new_n889_, keyIn_0_121 );
not g0676 ( new_n891_, keyIn_0_121 );
not g0677 ( new_n892_, new_n889_ );
nand g0678 ( new_n893_, new_n892_, new_n891_ );
nand g0679 ( N863, new_n893_, new_n890_ );
not g0680 ( new_n895_, keyIn_0_122 );
not g0681 ( new_n896_, keyIn_0_104 );
not g0682 ( new_n897_, keyIn_0_97 );
not g0683 ( new_n898_, new_n649_ );
not g0684 ( new_n899_, new_n766_ );
nor g0685 ( new_n900_, new_n898_, new_n899_ );
not g0686 ( new_n901_, new_n900_ );
nand g0687 ( new_n902_, new_n901_, new_n897_ );
nand g0688 ( new_n903_, new_n902_, new_n811_ );
nor g0689 ( new_n904_, new_n901_, new_n897_ );
nor g0690 ( new_n905_, new_n778_, new_n899_ );
nor g0691 ( new_n906_, new_n905_, keyIn_0_95 );
nand g0692 ( new_n907_, new_n905_, keyIn_0_95 );
not g0693 ( new_n908_, new_n907_ );
nor g0694 ( new_n909_, new_n908_, new_n906_ );
nor g0695 ( new_n910_, new_n904_, new_n909_ );
not g0696 ( new_n911_, new_n910_ );
nor g0697 ( new_n912_, new_n911_, new_n903_ );
nor g0698 ( new_n913_, new_n912_, new_n896_ );
nand g0699 ( new_n914_, new_n912_, new_n896_ );
not g0700 ( new_n915_, new_n914_ );
nor g0701 ( new_n916_, new_n915_, new_n913_ );
not g0702 ( new_n917_, new_n916_ );
not g0703 ( new_n918_, keyIn_0_90 );
not g0704 ( new_n919_, new_n790_ );
nor g0705 ( new_n920_, new_n919_, new_n808_ );
nor g0706 ( new_n921_, new_n920_, new_n918_ );
nand g0707 ( new_n922_, new_n920_, new_n918_ );
not g0708 ( new_n923_, new_n922_ );
nor g0709 ( new_n924_, new_n923_, new_n921_ );
not g0710 ( new_n925_, new_n924_ );
nand g0711 ( new_n926_, new_n917_, new_n925_ );
nor g0712 ( new_n927_, new_n926_, keyIn_0_107 );
nand g0713 ( new_n928_, new_n926_, keyIn_0_107 );
not g0714 ( new_n929_, N219 );
nor g0715 ( new_n930_, new_n917_, new_n925_ );
nor g0716 ( new_n931_, new_n930_, new_n929_ );
nand g0717 ( new_n932_, new_n931_, new_n928_ );
nor g0718 ( new_n933_, new_n932_, new_n927_ );
nand g0719 ( new_n934_, new_n925_, N228 );
nor g0720 ( new_n935_, new_n790_, new_n876_ );
nand g0721 ( new_n936_, new_n718_, N246 );
nand g0722 ( new_n937_, new_n662_, N189 );
nand g0723 ( new_n938_, N111, N210 );
nand g0724 ( new_n939_, N255, N259 );
nand g0725 ( new_n940_, new_n938_, new_n939_ );
not g0726 ( new_n941_, new_n940_ );
nand g0727 ( new_n942_, new_n937_, new_n941_ );
not g0728 ( new_n943_, new_n942_ );
nand g0729 ( new_n944_, new_n936_, new_n943_ );
nor g0730 ( new_n945_, new_n935_, new_n944_ );
nand g0731 ( new_n946_, new_n934_, new_n945_ );
nor g0732 ( new_n947_, new_n933_, new_n946_ );
nand g0733 ( new_n948_, new_n947_, new_n895_ );
not g0734 ( new_n949_, new_n947_ );
nand g0735 ( new_n950_, new_n949_, keyIn_0_122 );
nand g0736 ( N864, new_n950_, new_n948_ );
not g0737 ( new_n952_, keyIn_0_123 );
not g0738 ( new_n953_, keyIn_0_105 );
nor g0739 ( new_n954_, new_n649_, new_n781_ );
nor g0740 ( new_n955_, new_n954_, new_n953_ );
nand g0741 ( new_n956_, new_n954_, new_n953_ );
not g0742 ( new_n957_, new_n956_ );
nor g0743 ( new_n958_, new_n957_, new_n955_ );
not g0744 ( new_n959_, new_n958_ );
not g0745 ( new_n960_, keyIn_0_92 );
nor g0746 ( new_n961_, new_n899_, new_n803_ );
nor g0747 ( new_n962_, new_n961_, new_n960_ );
nand g0748 ( new_n963_, new_n961_, new_n960_ );
not g0749 ( new_n964_, new_n963_ );
nor g0750 ( new_n965_, new_n964_, new_n962_ );
not g0751 ( new_n966_, new_n965_ );
nor g0752 ( new_n967_, new_n959_, new_n966_ );
nor g0753 ( new_n968_, new_n967_, keyIn_0_108 );
nand g0754 ( new_n969_, new_n967_, keyIn_0_108 );
not g0755 ( new_n970_, new_n969_ );
nand g0756 ( new_n971_, new_n959_, new_n966_ );
nand g0757 ( new_n972_, new_n971_, N219 );
nor g0758 ( new_n973_, new_n970_, new_n972_ );
not g0759 ( new_n974_, new_n973_ );
nor g0760 ( new_n975_, new_n974_, new_n968_ );
nor g0761 ( new_n976_, new_n966_, new_n640_ );
nor g0762 ( new_n977_, new_n811_, new_n876_ );
nand g0763 ( new_n978_, new_n758_, N246 );
nand g0764 ( new_n979_, new_n662_, N195 );
nand g0765 ( new_n980_, N116, N210 );
nand g0766 ( new_n981_, N255, N260 );
nand g0767 ( new_n982_, new_n980_, new_n981_ );
not g0768 ( new_n983_, new_n982_ );
nand g0769 ( new_n984_, new_n979_, new_n983_ );
not g0770 ( new_n985_, new_n984_ );
nand g0771 ( new_n986_, new_n978_, new_n985_ );
nor g0772 ( new_n987_, new_n977_, new_n986_ );
not g0773 ( new_n988_, new_n987_ );
nor g0774 ( new_n989_, new_n976_, new_n988_ );
not g0775 ( new_n990_, new_n989_ );
nor g0776 ( new_n991_, new_n975_, new_n990_ );
nand g0777 ( new_n992_, new_n991_, new_n952_ );
not g0778 ( new_n993_, new_n991_ );
nand g0779 ( new_n994_, new_n993_, keyIn_0_123 );
nand g0780 ( N865, new_n994_, new_n992_ );
not g0781 ( new_n996_, keyIn_0_116 );
not g0782 ( new_n997_, keyIn_0_110 );
nor g0783 ( new_n998_, new_n827_, new_n857_ );
nand g0784 ( new_n999_, new_n998_, keyIn_0_109 );
not g0785 ( new_n1000_, keyIn_0_109 );
not g0786 ( new_n1001_, new_n817_ );
nor g0787 ( new_n1002_, new_n816_, new_n679_ );
nor g0788 ( new_n1003_, new_n1001_, new_n1002_ );
not g0789 ( new_n1004_, new_n857_ );
nand g0790 ( new_n1005_, new_n1003_, new_n1004_ );
nand g0791 ( new_n1006_, new_n1005_, new_n1000_ );
nand g0792 ( new_n1007_, new_n1006_, new_n999_ );
nand g0793 ( new_n1008_, new_n1007_, new_n858_ );
nor g0794 ( new_n1009_, new_n1008_, new_n997_ );
nand g0795 ( new_n1010_, new_n1008_, new_n997_ );
not g0796 ( new_n1011_, new_n1010_ );
nor g0797 ( new_n1012_, new_n1011_, new_n1009_ );
nor g0798 ( new_n1013_, new_n589_, new_n225_ );
nor g0799 ( new_n1014_, new_n1013_, keyIn_0_31 );
nand g0800 ( new_n1015_, new_n1013_, keyIn_0_31 );
not g0801 ( new_n1016_, new_n1015_ );
nor g0802 ( new_n1017_, new_n1016_, new_n1014_ );
nor g0803 ( new_n1018_, new_n1017_, new_n600_ );
not g0804 ( new_n1019_, new_n1018_ );
nand g0805 ( new_n1020_, new_n1019_, keyIn_0_43 );
not g0806 ( new_n1021_, new_n1020_ );
nor g0807 ( new_n1022_, new_n1019_, keyIn_0_43 );
nor g0808 ( new_n1023_, new_n1021_, new_n1022_ );
nor g0809 ( new_n1024_, new_n470_, new_n580_ );
nand g0810 ( new_n1025_, new_n477_, new_n1024_ );
not g0811 ( new_n1026_, new_n1025_ );
nor g0812 ( new_n1027_, new_n1026_, keyIn_0_30 );
nand g0813 ( new_n1028_, new_n1026_, keyIn_0_30 );
not g0814 ( new_n1029_, new_n1028_ );
nor g0815 ( new_n1030_, new_n1029_, new_n1027_ );
nor g0816 ( new_n1031_, new_n1030_, new_n560_ );
nor g0817 ( new_n1032_, new_n1023_, new_n1031_ );
nor g0818 ( new_n1033_, new_n1032_, keyIn_0_54 );
nand g0819 ( new_n1034_, new_n1032_, keyIn_0_54 );
not g0820 ( new_n1035_, new_n1034_ );
nor g0821 ( new_n1036_, new_n1035_, new_n1033_ );
nand g0822 ( new_n1037_, new_n555_, N106 );
nand g0823 ( new_n1038_, N138, N152 );
nand g0824 ( new_n1039_, new_n1037_, new_n1038_ );
nand g0825 ( new_n1040_, new_n1039_, keyIn_0_66 );
not g0826 ( new_n1041_, new_n1040_ );
nor g0827 ( new_n1042_, new_n1039_, keyIn_0_66 );
nor g0828 ( new_n1043_, new_n1041_, new_n1042_ );
nor g0829 ( new_n1044_, new_n1036_, new_n1043_ );
not g0830 ( new_n1045_, new_n1044_ );
nand g0831 ( new_n1046_, new_n1045_, keyIn_0_74 );
not g0832 ( new_n1047_, new_n1046_ );
nor g0833 ( new_n1048_, new_n1045_, keyIn_0_74 );
nor g0834 ( new_n1049_, new_n1047_, new_n1048_ );
nor g0835 ( new_n1050_, new_n1049_, N177 );
not g0836 ( new_n1051_, new_n1050_ );
nand g0837 ( new_n1052_, new_n1012_, new_n1051_ );
not g0838 ( new_n1053_, keyIn_0_52 );
not g0839 ( new_n1054_, keyIn_0_41 );
nand g0840 ( new_n1055_, new_n1019_, new_n1054_ );
not g0841 ( new_n1056_, new_n1055_ );
nor g0842 ( new_n1057_, new_n1019_, new_n1054_ );
nor g0843 ( new_n1058_, new_n1056_, new_n1057_ );
nor g0844 ( new_n1059_, new_n1030_, new_n696_ );
nor g0845 ( new_n1060_, new_n1058_, new_n1059_ );
nor g0846 ( new_n1061_, new_n1060_, new_n1053_ );
nand g0847 ( new_n1062_, new_n1060_, new_n1053_ );
not g0848 ( new_n1063_, new_n1062_ );
nor g0849 ( new_n1064_, new_n1063_, new_n1061_ );
not g0850 ( new_n1065_, keyIn_0_64 );
nand g0851 ( new_n1066_, new_n555_, N96 );
nand g0852 ( new_n1067_, N51, N138 );
nand g0853 ( new_n1068_, new_n1066_, new_n1067_ );
nand g0854 ( new_n1069_, new_n1068_, new_n1065_ );
not g0855 ( new_n1070_, new_n1069_ );
nor g0856 ( new_n1071_, new_n1068_, new_n1065_ );
nor g0857 ( new_n1072_, new_n1070_, new_n1071_ );
nor g0858 ( new_n1073_, new_n1064_, new_n1072_ );
not g0859 ( new_n1074_, new_n1073_ );
nand g0860 ( new_n1075_, new_n1074_, keyIn_0_72 );
not g0861 ( new_n1076_, new_n1075_ );
nor g0862 ( new_n1077_, new_n1074_, keyIn_0_72 );
nor g0863 ( new_n1078_, new_n1076_, new_n1077_ );
nor g0864 ( new_n1079_, new_n1078_, N165 );
not g0865 ( new_n1080_, keyIn_0_73 );
nand g0866 ( new_n1081_, new_n1019_, keyIn_0_42 );
not g0867 ( new_n1082_, new_n1081_ );
nor g0868 ( new_n1083_, new_n1019_, keyIn_0_42 );
nor g0869 ( new_n1084_, new_n1082_, new_n1083_ );
nor g0870 ( new_n1085_, new_n1030_, new_n737_ );
nor g0871 ( new_n1086_, new_n1084_, new_n1085_ );
not g0872 ( new_n1087_, new_n1086_ );
nand g0873 ( new_n1088_, new_n1087_, keyIn_0_53 );
not g0874 ( new_n1089_, keyIn_0_65 );
nand g0875 ( new_n1090_, new_n555_, N101 );
nand g0876 ( new_n1091_, N17, N138 );
nand g0877 ( new_n1092_, new_n1090_, new_n1091_ );
nand g0878 ( new_n1093_, new_n1092_, new_n1089_ );
nand g0879 ( new_n1094_, new_n1088_, new_n1093_ );
nor g0880 ( new_n1095_, new_n1087_, keyIn_0_53 );
nor g0881 ( new_n1096_, new_n1092_, new_n1089_ );
nor g0882 ( new_n1097_, new_n1095_, new_n1096_ );
not g0883 ( new_n1098_, new_n1097_ );
nor g0884 ( new_n1099_, new_n1098_, new_n1094_ );
not g0885 ( new_n1100_, new_n1099_ );
nor g0886 ( new_n1101_, new_n1100_, new_n1080_ );
nor g0887 ( new_n1102_, new_n1099_, keyIn_0_73 );
nor g0888 ( new_n1103_, new_n1101_, new_n1102_ );
not g0889 ( new_n1104_, new_n1103_ );
nor g0890 ( new_n1105_, new_n1104_, N171 );
nor g0891 ( new_n1106_, new_n1105_, new_n1079_ );
not g0892 ( new_n1107_, new_n1106_ );
nor g0893 ( new_n1108_, new_n1052_, new_n1107_ );
nand g0894 ( new_n1109_, new_n1108_, keyIn_0_115 );
nor g0895 ( new_n1110_, new_n1108_, keyIn_0_115 );
not g0896 ( new_n1111_, new_n1110_ );
nand g0897 ( new_n1112_, new_n1111_, new_n1109_ );
nand g0898 ( new_n1113_, new_n1104_, N171 );
nor g0899 ( new_n1114_, new_n1113_, new_n1079_ );
not g0900 ( new_n1115_, new_n1114_ );
nor g0901 ( new_n1116_, new_n1115_, keyIn_0_101 );
nand g0902 ( new_n1117_, new_n1115_, keyIn_0_101 );
nand g0903 ( new_n1118_, new_n1078_, N165 );
nand g0904 ( new_n1119_, new_n1117_, new_n1118_ );
nor g0905 ( new_n1120_, new_n1119_, new_n1116_ );
nand g0906 ( new_n1121_, new_n1049_, N177 );
nor g0907 ( new_n1122_, new_n1107_, new_n1121_ );
nor g0908 ( new_n1123_, new_n1122_, keyIn_0_102 );
nand g0909 ( new_n1124_, new_n1122_, keyIn_0_102 );
not g0910 ( new_n1125_, new_n1124_ );
nor g0911 ( new_n1126_, new_n1125_, new_n1123_ );
nand g0912 ( new_n1127_, new_n1126_, new_n1120_ );
not g0913 ( new_n1128_, new_n1127_ );
nand g0914 ( new_n1129_, new_n1112_, new_n1128_ );
nand g0915 ( new_n1130_, new_n1129_, new_n996_ );
nor g0916 ( new_n1131_, new_n1129_, new_n996_ );
not g0917 ( new_n1132_, new_n1131_ );
nand g0918 ( new_n1133_, new_n1132_, new_n1130_ );
not g0919 ( new_n1134_, keyIn_0_71 );
not g0920 ( new_n1135_, keyIn_0_51 );
not g0921 ( new_n1136_, keyIn_0_40 );
nand g0922 ( new_n1137_, new_n1019_, new_n1136_ );
not g0923 ( new_n1138_, new_n1137_ );
nor g0924 ( new_n1139_, new_n1019_, new_n1136_ );
nor g0925 ( new_n1140_, new_n1138_, new_n1139_ );
nor g0926 ( new_n1141_, new_n1030_, new_n830_ );
nor g0927 ( new_n1142_, new_n1140_, new_n1141_ );
nor g0928 ( new_n1143_, new_n1142_, new_n1135_ );
nand g0929 ( new_n1144_, new_n1142_, new_n1135_ );
not g0930 ( new_n1145_, new_n1144_ );
nor g0931 ( new_n1146_, new_n1145_, new_n1143_ );
not g0932 ( new_n1147_, keyIn_0_63 );
nand g0933 ( new_n1148_, new_n555_, N91 );
nand g0934 ( new_n1149_, N8, N138 );
nand g0935 ( new_n1150_, new_n1148_, new_n1149_ );
nand g0936 ( new_n1151_, new_n1150_, new_n1147_ );
not g0937 ( new_n1152_, new_n1151_ );
nor g0938 ( new_n1153_, new_n1150_, new_n1147_ );
nor g0939 ( new_n1154_, new_n1152_, new_n1153_ );
nor g0940 ( new_n1155_, new_n1146_, new_n1154_ );
not g0941 ( new_n1156_, new_n1155_ );
nand g0942 ( new_n1157_, new_n1156_, new_n1134_ );
not g0943 ( new_n1158_, new_n1157_ );
nor g0944 ( new_n1159_, new_n1156_, new_n1134_ );
nor g0945 ( new_n1160_, new_n1158_, new_n1159_ );
nor g0946 ( new_n1161_, new_n1160_, N159 );
not g0947 ( new_n1162_, new_n1161_ );
nand g0948 ( new_n1163_, new_n1133_, new_n1162_ );
nand g0949 ( new_n1164_, new_n1160_, N159 );
nand g0950 ( N866, new_n1163_, new_n1164_ );
not g0951 ( new_n1166_, keyIn_0_111 );
not g0952 ( new_n1167_, new_n1009_ );
nand g0953 ( new_n1168_, new_n1167_, new_n1010_ );
not g0954 ( new_n1169_, keyIn_0_88 );
not g0955 ( new_n1170_, new_n1121_ );
nor g0956 ( new_n1171_, new_n1170_, new_n1050_ );
nor g0957 ( new_n1172_, new_n1171_, new_n1169_ );
nand g0958 ( new_n1173_, new_n1171_, new_n1169_ );
not g0959 ( new_n1174_, new_n1173_ );
nor g0960 ( new_n1175_, new_n1174_, new_n1172_ );
nor g0961 ( new_n1176_, new_n1168_, new_n1175_ );
not g0962 ( new_n1177_, new_n1176_ );
nand g0963 ( new_n1178_, new_n1177_, new_n1166_ );
nand g0964 ( new_n1179_, new_n1176_, keyIn_0_111 );
nand g0965 ( new_n1180_, new_n1178_, new_n1179_ );
not g0966 ( new_n1181_, new_n1175_ );
nor g0967 ( new_n1182_, new_n1012_, new_n1181_ );
nor g0968 ( new_n1183_, new_n1182_, new_n929_ );
nand g0969 ( new_n1184_, new_n1180_, new_n1183_ );
nand g0970 ( new_n1185_, new_n1181_, N228 );
nor g0971 ( new_n1186_, new_n1121_, new_n876_ );
nand g0972 ( new_n1187_, new_n1049_, N246 );
nand g0973 ( new_n1188_, new_n662_, N177 );
nand g0974 ( new_n1189_, N101, N210 );
nand g0975 ( new_n1190_, new_n1188_, new_n1189_ );
not g0976 ( new_n1191_, new_n1190_ );
nand g0977 ( new_n1192_, new_n1187_, new_n1191_ );
nor g0978 ( new_n1193_, new_n1186_, new_n1192_ );
nand g0979 ( new_n1194_, new_n1185_, new_n1193_ );
not g0980 ( new_n1195_, new_n1194_ );
nand g0981 ( new_n1196_, new_n1184_, new_n1195_ );
not g0982 ( new_n1197_, new_n1196_ );
nand g0983 ( new_n1198_, new_n1197_, keyIn_0_124 );
not g0984 ( new_n1199_, keyIn_0_124 );
nand g0985 ( new_n1200_, new_n1196_, new_n1199_ );
nand g0986 ( N874, new_n1198_, new_n1200_ );
not g0987 ( new_n1202_, keyIn_0_125 );
nand g0988 ( new_n1203_, new_n1162_, new_n1164_ );
not g0989 ( new_n1204_, new_n1203_ );
nor g0990 ( new_n1205_, new_n1204_, keyIn_0_85 );
nand g0991 ( new_n1206_, new_n1204_, keyIn_0_85 );
not g0992 ( new_n1207_, new_n1206_ );
nor g0993 ( new_n1208_, new_n1207_, new_n1205_ );
not g0994 ( new_n1209_, new_n1208_ );
nor g0995 ( new_n1210_, new_n1133_, new_n1209_ );
nand g0996 ( new_n1211_, new_n1133_, new_n1209_ );
nand g0997 ( new_n1212_, new_n1211_, N219 );
nor g0998 ( new_n1213_, new_n1212_, new_n1210_ );
nand g0999 ( new_n1214_, new_n1209_, N228 );
nor g1000 ( new_n1215_, new_n1164_, new_n876_ );
nand g1001 ( new_n1216_, new_n1160_, N246 );
nand g1002 ( new_n1217_, new_n662_, N159 );
nand g1003 ( new_n1218_, new_n605_, N210 );
nand g1004 ( new_n1219_, new_n1217_, new_n1218_ );
not g1005 ( new_n1220_, new_n1219_ );
nand g1006 ( new_n1221_, new_n1216_, new_n1220_ );
nor g1007 ( new_n1222_, new_n1215_, new_n1221_ );
nand g1008 ( new_n1223_, new_n1214_, new_n1222_ );
nor g1009 ( new_n1224_, new_n1213_, new_n1223_ );
nand g1010 ( new_n1225_, new_n1224_, new_n1202_ );
not g1011 ( new_n1226_, new_n1210_ );
not g1012 ( new_n1227_, new_n1130_ );
nor g1013 ( new_n1228_, new_n1227_, new_n1131_ );
nor g1014 ( new_n1229_, new_n1228_, new_n1208_ );
nor g1015 ( new_n1230_, new_n1229_, new_n929_ );
nand g1016 ( new_n1231_, new_n1230_, new_n1226_ );
not g1017 ( new_n1232_, new_n1223_ );
nand g1018 ( new_n1233_, new_n1231_, new_n1232_ );
nand g1019 ( new_n1234_, new_n1233_, keyIn_0_125 );
nand g1020 ( N878, new_n1234_, new_n1225_ );
not g1021 ( new_n1236_, keyIn_0_119 );
not g1022 ( new_n1237_, keyIn_0_114 );
nor g1023 ( new_n1238_, new_n1168_, new_n1050_ );
not g1024 ( new_n1239_, new_n1105_ );
nand g1025 ( new_n1240_, new_n1238_, new_n1239_ );
nor g1026 ( new_n1241_, new_n1240_, new_n1237_ );
nand g1027 ( new_n1242_, new_n1240_, new_n1237_ );
nor g1028 ( new_n1243_, new_n1105_, new_n1121_ );
not g1029 ( new_n1244_, new_n1243_ );
nor g1030 ( new_n1245_, new_n1244_, keyIn_0_100 );
nand g1031 ( new_n1246_, new_n1244_, keyIn_0_100 );
nand g1032 ( new_n1247_, new_n1246_, new_n1113_ );
nor g1033 ( new_n1248_, new_n1247_, new_n1245_ );
nand g1034 ( new_n1249_, new_n1242_, new_n1248_ );
nor g1035 ( new_n1250_, new_n1249_, new_n1241_ );
nor g1036 ( new_n1251_, new_n1250_, keyIn_0_117 );
not g1037 ( new_n1252_, keyIn_0_117 );
not g1038 ( new_n1253_, new_n1241_ );
nor g1039 ( new_n1254_, new_n1052_, new_n1105_ );
nor g1040 ( new_n1255_, new_n1254_, keyIn_0_114 );
not g1041 ( new_n1256_, new_n1248_ );
nor g1042 ( new_n1257_, new_n1255_, new_n1256_ );
nand g1043 ( new_n1258_, new_n1257_, new_n1253_ );
nor g1044 ( new_n1259_, new_n1258_, new_n1252_ );
nor g1045 ( new_n1260_, new_n1259_, new_n1251_ );
not g1046 ( new_n1261_, new_n1118_ );
nor g1047 ( new_n1262_, new_n1261_, new_n1079_ );
nor g1048 ( new_n1263_, new_n1262_, keyIn_0_86 );
nand g1049 ( new_n1264_, new_n1262_, keyIn_0_86 );
not g1050 ( new_n1265_, new_n1264_ );
nor g1051 ( new_n1266_, new_n1265_, new_n1263_ );
not g1052 ( new_n1267_, new_n1266_ );
nand g1053 ( new_n1268_, new_n1260_, new_n1267_ );
nor g1054 ( new_n1269_, new_n1268_, new_n1236_ );
nand g1055 ( new_n1270_, new_n1268_, new_n1236_ );
nand g1056 ( new_n1271_, new_n1258_, new_n1252_ );
nand g1057 ( new_n1272_, new_n1250_, keyIn_0_117 );
nand g1058 ( new_n1273_, new_n1271_, new_n1272_ );
nand g1059 ( new_n1274_, new_n1273_, new_n1266_ );
nand g1060 ( new_n1275_, new_n1274_, N219 );
not g1061 ( new_n1276_, new_n1275_ );
nand g1062 ( new_n1277_, new_n1276_, new_n1270_ );
nor g1063 ( new_n1278_, new_n1277_, new_n1269_ );
nand g1064 ( new_n1279_, new_n1267_, N228 );
nor g1065 ( new_n1280_, new_n1118_, new_n876_ );
nand g1066 ( new_n1281_, new_n1078_, N246 );
nand g1067 ( new_n1282_, new_n662_, N165 );
nand g1068 ( new_n1283_, N91, N210 );
nand g1069 ( new_n1284_, new_n1282_, new_n1283_ );
not g1070 ( new_n1285_, new_n1284_ );
nand g1071 ( new_n1286_, new_n1281_, new_n1285_ );
nor g1072 ( new_n1287_, new_n1280_, new_n1286_ );
nand g1073 ( new_n1288_, new_n1279_, new_n1287_ );
nor g1074 ( new_n1289_, new_n1278_, new_n1288_ );
nand g1075 ( new_n1290_, new_n1289_, keyIn_0_126 );
not g1076 ( new_n1291_, keyIn_0_126 );
not g1077 ( new_n1292_, new_n1269_ );
nor g1078 ( new_n1293_, new_n1273_, new_n1266_ );
nor g1079 ( new_n1294_, new_n1293_, keyIn_0_119 );
nor g1080 ( new_n1295_, new_n1294_, new_n1275_ );
nand g1081 ( new_n1296_, new_n1295_, new_n1292_ );
not g1082 ( new_n1297_, new_n1288_ );
nand g1083 ( new_n1298_, new_n1296_, new_n1297_ );
nand g1084 ( new_n1299_, new_n1298_, new_n1291_ );
nand g1085 ( N879, new_n1290_, new_n1299_ );
not g1086 ( new_n1301_, keyIn_0_118 );
nand g1087 ( new_n1302_, new_n1052_, keyIn_0_113 );
not g1088 ( new_n1303_, keyIn_0_113 );
nand g1089 ( new_n1304_, new_n1238_, new_n1303_ );
nand g1090 ( new_n1305_, new_n1304_, new_n1302_ );
nand g1091 ( new_n1306_, new_n1305_, new_n1121_ );
nand g1092 ( new_n1307_, new_n1306_, new_n1301_ );
not g1093 ( new_n1308_, new_n1307_ );
nor g1094 ( new_n1309_, new_n1306_, new_n1301_ );
nor g1095 ( new_n1310_, new_n1308_, new_n1309_ );
not g1096 ( new_n1311_, keyIn_0_87 );
not g1097 ( new_n1312_, new_n1113_ );
nor g1098 ( new_n1313_, new_n1312_, new_n1105_ );
nor g1099 ( new_n1314_, new_n1313_, new_n1311_ );
nand g1100 ( new_n1315_, new_n1313_, new_n1311_ );
not g1101 ( new_n1316_, new_n1315_ );
nor g1102 ( new_n1317_, new_n1316_, new_n1314_ );
nand g1103 ( new_n1318_, new_n1310_, new_n1317_ );
nor g1104 ( new_n1319_, new_n1318_, keyIn_0_120 );
nand g1105 ( new_n1320_, new_n1318_, keyIn_0_120 );
nor g1106 ( new_n1321_, new_n1310_, new_n1317_ );
nor g1107 ( new_n1322_, new_n1321_, new_n929_ );
nand g1108 ( new_n1323_, new_n1322_, new_n1320_ );
nor g1109 ( new_n1324_, new_n1323_, new_n1319_ );
not g1110 ( new_n1325_, new_n1317_ );
nor g1111 ( new_n1326_, new_n1325_, new_n640_ );
nor g1112 ( new_n1327_, new_n1113_, new_n876_ );
nand g1113 ( new_n1328_, new_n1104_, N246 );
nand g1114 ( new_n1329_, new_n662_, N171 );
nand g1115 ( new_n1330_, N96, N210 );
nand g1116 ( new_n1331_, new_n1329_, new_n1330_ );
not g1117 ( new_n1332_, new_n1331_ );
nand g1118 ( new_n1333_, new_n1328_, new_n1332_ );
nor g1119 ( new_n1334_, new_n1327_, new_n1333_ );
not g1120 ( new_n1335_, new_n1334_ );
nor g1121 ( new_n1336_, new_n1326_, new_n1335_ );
not g1122 ( new_n1337_, new_n1336_ );
nor g1123 ( new_n1338_, new_n1324_, new_n1337_ );
nand g1124 ( new_n1339_, new_n1338_, keyIn_0_127 );
not g1125 ( new_n1340_, keyIn_0_127 );
not g1126 ( new_n1341_, new_n1324_ );
nand g1127 ( new_n1342_, new_n1341_, new_n1336_ );
nand g1128 ( new_n1343_, new_n1342_, new_n1340_ );
nand g1129 ( N880, new_n1343_, new_n1339_ );
endmodule