module add_mul_sub_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        operation_0_, operation_1_, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, operation_0_,
         operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479;

  OR2_X1 U252 ( .A1(n244), .A2(n245), .ZN(Result_7_) );
  AND2_X1 U253 ( .A1(n246), .A2(n247), .ZN(n245) );
  OR2_X1 U254 ( .A1(n248), .A2(n249), .ZN(n246) );
  AND2_X1 U255 ( .A1(n250), .A2(n251), .ZN(n244) );
  OR3_X1 U256 ( .A1(n252), .A2(n253), .A3(n254), .ZN(Result_6_) );
  AND2_X1 U257 ( .A1(n251), .A2(n255), .ZN(n254) );
  OR4_X1 U258 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(n255) );
  AND2_X1 U259 ( .A1(n260), .A2(a_3_), .ZN(n259) );
  AND2_X1 U260 ( .A1(n261), .A2(b_3_), .ZN(n258) );
  AND2_X1 U261 ( .A1(n249), .A2(a_2_), .ZN(n257) );
  AND2_X1 U262 ( .A1(n248), .A2(b_2_), .ZN(n256) );
  AND2_X1 U263 ( .A1(n262), .A2(n263), .ZN(n253) );
  OR3_X1 U264 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n263) );
  AND2_X1 U265 ( .A1(n249), .A2(n267), .ZN(n266) );
  AND2_X1 U266 ( .A1(n248), .A2(n268), .ZN(n265) );
  AND2_X1 U267 ( .A1(n269), .A2(n250), .ZN(n264) );
  OR2_X1 U268 ( .A1(n270), .A2(n271), .ZN(n262) );
  AND2_X1 U269 ( .A1(n272), .A2(n273), .ZN(n252) );
  OR3_X1 U270 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n273) );
  AND2_X1 U271 ( .A1(n267), .A2(n277), .ZN(n276) );
  AND2_X1 U272 ( .A1(n268), .A2(n278), .ZN(n275) );
  AND2_X1 U273 ( .A1(n269), .A2(n279), .ZN(n274) );
  OR2_X1 U274 ( .A1(n261), .A2(n260), .ZN(n272) );
  INV_X1 U275 ( .A(n280), .ZN(n261) );
  OR3_X1 U276 ( .A1(n281), .A2(n282), .A3(n283), .ZN(Result_5_) );
  AND2_X1 U277 ( .A1(n251), .A2(n284), .ZN(n283) );
  OR2_X1 U278 ( .A1(n285), .A2(n286), .ZN(n284) );
  AND2_X1 U279 ( .A1(n287), .A2(n288), .ZN(n286) );
  INV_X1 U280 ( .A(n289), .ZN(n285) );
  OR2_X1 U281 ( .A1(n288), .A2(n287), .ZN(n289) );
  OR2_X1 U282 ( .A1(n290), .A2(n291), .ZN(n287) );
  AND2_X1 U283 ( .A1(n292), .A2(n293), .ZN(n291) );
  AND2_X1 U284 ( .A1(n294), .A2(n295), .ZN(n290) );
  INV_X1 U285 ( .A(n293), .ZN(n294) );
  AND2_X1 U286 ( .A1(n296), .A2(n297), .ZN(n282) );
  OR3_X1 U287 ( .A1(n298), .A2(n299), .A3(n300), .ZN(n297) );
  AND2_X1 U288 ( .A1(n267), .A2(n301), .ZN(n300) );
  AND2_X1 U289 ( .A1(n268), .A2(n302), .ZN(n299) );
  AND2_X1 U290 ( .A1(n303), .A2(n269), .ZN(n298) );
  INV_X1 U291 ( .A(n304), .ZN(n296) );
  AND2_X1 U292 ( .A1(n304), .A2(n305), .ZN(n281) );
  OR3_X1 U293 ( .A1(n306), .A2(n307), .A3(n308), .ZN(n305) );
  AND2_X1 U294 ( .A1(n309), .A2(n267), .ZN(n308) );
  INV_X1 U295 ( .A(n301), .ZN(n309) );
  AND2_X1 U296 ( .A1(n310), .A2(n268), .ZN(n307) );
  AND2_X1 U297 ( .A1(n269), .A2(n311), .ZN(n306) );
  OR2_X1 U298 ( .A1(n312), .A2(n313), .ZN(n304) );
  AND2_X1 U299 ( .A1(a_1_), .A2(n314), .ZN(n313) );
  AND2_X1 U300 ( .A1(b_1_), .A2(n315), .ZN(n312) );
  OR3_X1 U301 ( .A1(n316), .A2(n317), .A3(n318), .ZN(Result_4_) );
  AND2_X1 U302 ( .A1(n251), .A2(n319), .ZN(n318) );
  OR2_X1 U303 ( .A1(n320), .A2(n321), .ZN(n319) );
  AND2_X1 U304 ( .A1(n322), .A2(n323), .ZN(n321) );
  INV_X1 U305 ( .A(n324), .ZN(n320) );
  OR2_X1 U306 ( .A1(n323), .A2(n322), .ZN(n324) );
  OR2_X1 U307 ( .A1(n325), .A2(n326), .ZN(n322) );
  AND2_X1 U308 ( .A1(n327), .A2(n328), .ZN(n326) );
  INV_X1 U309 ( .A(n329), .ZN(n325) );
  OR2_X1 U310 ( .A1(n328), .A2(n327), .ZN(n329) );
  AND2_X1 U311 ( .A1(n330), .A2(n331), .ZN(n317) );
  OR3_X1 U312 ( .A1(n332), .A2(n333), .A3(n334), .ZN(n330) );
  AND2_X1 U313 ( .A1(n335), .A2(n267), .ZN(n334) );
  INV_X1 U314 ( .A(n336), .ZN(n335) );
  AND2_X1 U315 ( .A1(n337), .A2(n268), .ZN(n333) );
  INV_X1 U316 ( .A(n338), .ZN(n337) );
  AND2_X1 U317 ( .A1(n339), .A2(n269), .ZN(n332) );
  INV_X1 U318 ( .A(n340), .ZN(n339) );
  AND2_X1 U319 ( .A1(n341), .A2(n342), .ZN(n316) );
  OR3_X1 U320 ( .A1(n343), .A2(n344), .A3(n345), .ZN(n342) );
  AND2_X1 U321 ( .A1(n267), .A2(n336), .ZN(n345) );
  AND2_X1 U322 ( .A1(n268), .A2(n338), .ZN(n344) );
  AND2_X1 U323 ( .A1(n269), .A2(n340), .ZN(n343) );
  OR2_X1 U324 ( .A1(n346), .A2(n347), .ZN(n340) );
  AND2_X1 U325 ( .A1(n303), .A2(a_1_), .ZN(n347) );
  AND2_X1 U326 ( .A1(b_1_), .A2(n348), .ZN(n346) );
  OR2_X1 U327 ( .A1(n303), .A2(a_1_), .ZN(n348) );
  INV_X1 U328 ( .A(n311), .ZN(n303) );
  OR2_X1 U329 ( .A1(n349), .A2(n270), .ZN(n311) );
  AND2_X1 U330 ( .A1(n350), .A2(n351), .ZN(n270) );
  AND2_X1 U331 ( .A1(n352), .A2(n279), .ZN(n349) );
  AND2_X1 U332 ( .A1(n353), .A2(n354), .ZN(n269) );
  INV_X1 U333 ( .A(n331), .ZN(n341) );
  OR2_X1 U334 ( .A1(n355), .A2(n356), .ZN(n331) );
  OR2_X1 U335 ( .A1(n357), .A2(n358), .ZN(Result_3_) );
  AND3_X1 U336 ( .A1(n359), .A2(n360), .A3(n251), .ZN(n357) );
  OR2_X1 U337 ( .A1(n361), .A2(n362), .ZN(n360) );
  INV_X1 U338 ( .A(n363), .ZN(n362) );
  OR2_X1 U339 ( .A1(n364), .A2(n363), .ZN(n359) );
  OR2_X1 U340 ( .A1(n365), .A2(n358), .ZN(Result_2_) );
  AND3_X1 U341 ( .A1(n366), .A2(n367), .A3(n251), .ZN(n365) );
  INV_X1 U342 ( .A(n368), .ZN(n367) );
  OR2_X1 U343 ( .A1(n369), .A2(n370), .ZN(n366) );
  AND2_X1 U344 ( .A1(n364), .A2(n363), .ZN(n369) );
  OR2_X1 U345 ( .A1(n371), .A2(n358), .ZN(Result_1_) );
  AND3_X1 U346 ( .A1(n372), .A2(n373), .A3(n251), .ZN(n371) );
  INV_X1 U347 ( .A(n374), .ZN(n373) );
  OR2_X1 U348 ( .A1(n368), .A2(n375), .ZN(n372) );
  OR2_X1 U349 ( .A1(n376), .A2(n358), .ZN(Result_0_) );
  OR2_X1 U350 ( .A1(n377), .A2(n378), .ZN(n358) );
  AND2_X1 U351 ( .A1(n267), .A2(n379), .ZN(n378) );
  OR2_X1 U352 ( .A1(n380), .A2(n356), .ZN(n379) );
  INV_X1 U353 ( .A(n381), .ZN(n356) );
  AND2_X1 U354 ( .A1(n336), .A2(n382), .ZN(n380) );
  OR2_X1 U355 ( .A1(n383), .A2(n384), .ZN(n336) );
  AND2_X1 U356 ( .A1(n301), .A2(n315), .ZN(n384) );
  AND2_X1 U357 ( .A1(b_1_), .A2(n385), .ZN(n383) );
  OR2_X1 U358 ( .A1(n315), .A2(n301), .ZN(n385) );
  OR2_X1 U359 ( .A1(n386), .A2(n260), .ZN(n301) );
  AND2_X1 U360 ( .A1(n249), .A2(n280), .ZN(n386) );
  INV_X1 U361 ( .A(n277), .ZN(n249) );
  OR2_X1 U362 ( .A1(a_3_), .A2(n387), .ZN(n277) );
  AND2_X1 U363 ( .A1(n354), .A2(operation_1_), .ZN(n267) );
  AND3_X1 U364 ( .A1(n388), .A2(n381), .A3(n268), .ZN(n377) );
  AND2_X1 U365 ( .A1(n353), .A2(operation_0_), .ZN(n268) );
  OR2_X1 U366 ( .A1(a_0_), .A2(n389), .ZN(n381) );
  OR2_X1 U367 ( .A1(n355), .A2(n338), .ZN(n388) );
  OR2_X1 U368 ( .A1(n390), .A2(n391), .ZN(n338) );
  AND2_X1 U369 ( .A1(a_1_), .A2(n302), .ZN(n391) );
  AND2_X1 U370 ( .A1(n392), .A2(n314), .ZN(n390) );
  OR2_X1 U371 ( .A1(a_1_), .A2(n302), .ZN(n392) );
  INV_X1 U372 ( .A(n310), .ZN(n302) );
  AND2_X1 U373 ( .A1(n393), .A2(n280), .ZN(n310) );
  OR2_X1 U374 ( .A1(b_2_), .A2(n350), .ZN(n280) );
  OR2_X1 U375 ( .A1(n278), .A2(n260), .ZN(n393) );
  AND2_X1 U376 ( .A1(n350), .A2(b_2_), .ZN(n260) );
  INV_X1 U377 ( .A(n248), .ZN(n278) );
  AND2_X1 U378 ( .A1(n387), .A2(a_3_), .ZN(n248) );
  INV_X1 U379 ( .A(b_3_), .ZN(n387) );
  INV_X1 U380 ( .A(n382), .ZN(n355) );
  OR2_X1 U381 ( .A1(b_0_), .A2(n394), .ZN(n382) );
  AND2_X1 U382 ( .A1(n251), .A2(n395), .ZN(n376) );
  OR3_X1 U383 ( .A1(n396), .A2(n374), .A3(n397), .ZN(n395) );
  AND2_X1 U384 ( .A1(n375), .A2(n368), .ZN(n374) );
  AND3_X1 U385 ( .A1(n364), .A2(n363), .A3(n370), .ZN(n368) );
  AND2_X1 U386 ( .A1(n398), .A2(n399), .ZN(n370) );
  INV_X1 U387 ( .A(n400), .ZN(n399) );
  AND2_X1 U388 ( .A1(n401), .A2(n402), .ZN(n400) );
  AND2_X1 U389 ( .A1(n403), .A2(n404), .ZN(n363) );
  OR2_X1 U390 ( .A1(n405), .A2(n406), .ZN(n404) );
  INV_X1 U391 ( .A(n407), .ZN(n403) );
  AND2_X1 U392 ( .A1(n406), .A2(n405), .ZN(n407) );
  AND2_X1 U393 ( .A1(n408), .A2(n409), .ZN(n405) );
  OR2_X1 U394 ( .A1(n410), .A2(n411), .ZN(n409) );
  INV_X1 U395 ( .A(n412), .ZN(n411) );
  OR2_X1 U396 ( .A1(n412), .A2(n413), .ZN(n408) );
  INV_X1 U397 ( .A(n410), .ZN(n413) );
  INV_X1 U398 ( .A(n361), .ZN(n364) );
  OR2_X1 U399 ( .A1(n414), .A2(n415), .ZN(n361) );
  AND2_X1 U400 ( .A1(n416), .A2(n328), .ZN(n415) );
  AND2_X1 U401 ( .A1(n323), .A2(n417), .ZN(n414) );
  OR2_X1 U402 ( .A1(n328), .A2(n416), .ZN(n417) );
  INV_X1 U403 ( .A(n327), .ZN(n416) );
  AND2_X1 U404 ( .A1(b_3_), .A2(a_0_), .ZN(n327) );
  OR2_X1 U405 ( .A1(n418), .A2(n419), .ZN(n328) );
  AND2_X1 U406 ( .A1(n295), .A2(n293), .ZN(n419) );
  AND2_X1 U407 ( .A1(n288), .A2(n420), .ZN(n418) );
  OR2_X1 U408 ( .A1(n293), .A2(n295), .ZN(n420) );
  INV_X1 U409 ( .A(n292), .ZN(n295) );
  AND2_X1 U410 ( .A1(b_3_), .A2(a_1_), .ZN(n292) );
  OR2_X1 U411 ( .A1(n279), .A2(n352), .ZN(n293) );
  INV_X1 U412 ( .A(n250), .ZN(n279) );
  AND2_X1 U413 ( .A1(a_3_), .A2(b_3_), .ZN(n250) );
  AND2_X1 U414 ( .A1(n421), .A2(n422), .ZN(n288) );
  OR2_X1 U415 ( .A1(n352), .A2(n423), .ZN(n422) );
  OR2_X1 U416 ( .A1(n424), .A2(n271), .ZN(n421) );
  INV_X1 U417 ( .A(n352), .ZN(n271) );
  AND2_X1 U418 ( .A1(n425), .A2(n426), .ZN(n323) );
  INV_X1 U419 ( .A(n427), .ZN(n426) );
  AND2_X1 U420 ( .A1(n428), .A2(n429), .ZN(n427) );
  OR2_X1 U421 ( .A1(n429), .A2(n428), .ZN(n425) );
  OR2_X1 U422 ( .A1(n430), .A2(n431), .ZN(n428) );
  AND2_X1 U423 ( .A1(n432), .A2(n433), .ZN(n431) );
  INV_X1 U424 ( .A(n434), .ZN(n430) );
  OR2_X1 U425 ( .A1(n433), .A2(n432), .ZN(n434) );
  INV_X1 U426 ( .A(n435), .ZN(n375) );
  OR2_X1 U427 ( .A1(n436), .A2(n396), .ZN(n435) );
  AND2_X1 U428 ( .A1(n437), .A2(n398), .ZN(n436) );
  OR2_X1 U429 ( .A1(n401), .A2(n402), .ZN(n398) );
  INV_X1 U430 ( .A(n438), .ZN(n396) );
  OR3_X1 U431 ( .A1(n402), .A2(n401), .A3(n437), .ZN(n438) );
  OR2_X1 U432 ( .A1(n397), .A2(n439), .ZN(n437) );
  AND2_X1 U433 ( .A1(n440), .A2(n441), .ZN(n439) );
  OR2_X1 U434 ( .A1(n389), .A2(n394), .ZN(n440) );
  AND2_X1 U435 ( .A1(n442), .A2(a_0_), .ZN(n397) );
  INV_X1 U436 ( .A(n441), .ZN(n442) );
  OR2_X1 U437 ( .A1(n443), .A2(n444), .ZN(n441) );
  AND2_X1 U438 ( .A1(n445), .A2(n446), .ZN(n444) );
  AND2_X1 U439 ( .A1(n447), .A2(n448), .ZN(n443) );
  OR2_X1 U440 ( .A1(n446), .A2(n445), .ZN(n448) );
  OR2_X1 U441 ( .A1(n449), .A2(n450), .ZN(n401) );
  AND2_X1 U442 ( .A1(n451), .A2(n445), .ZN(n450) );
  INV_X1 U443 ( .A(n452), .ZN(n449) );
  OR2_X1 U444 ( .A1(n451), .A2(n445), .ZN(n452) );
  OR2_X1 U445 ( .A1(n314), .A2(n394), .ZN(n445) );
  OR2_X1 U446 ( .A1(n453), .A2(n454), .ZN(n451) );
  AND2_X1 U447 ( .A1(n447), .A2(n446), .ZN(n454) );
  INV_X1 U448 ( .A(n455), .ZN(n447) );
  AND2_X1 U449 ( .A1(n456), .A2(n455), .ZN(n453) );
  OR2_X1 U450 ( .A1(n457), .A2(n458), .ZN(n455) );
  AND2_X1 U451 ( .A1(n456), .A2(n459), .ZN(n457) );
  INV_X1 U452 ( .A(n446), .ZN(n456) );
  OR2_X1 U453 ( .A1(n315), .A2(n389), .ZN(n446) );
  OR2_X1 U454 ( .A1(n460), .A2(n461), .ZN(n402) );
  AND2_X1 U455 ( .A1(n410), .A2(n412), .ZN(n461) );
  AND2_X1 U456 ( .A1(n406), .A2(n462), .ZN(n460) );
  OR2_X1 U457 ( .A1(n412), .A2(n410), .ZN(n462) );
  OR2_X1 U458 ( .A1(n351), .A2(n394), .ZN(n410) );
  INV_X1 U459 ( .A(a_0_), .ZN(n394) );
  OR2_X1 U460 ( .A1(n463), .A2(n464), .ZN(n412) );
  AND2_X1 U461 ( .A1(n465), .A2(n433), .ZN(n464) );
  AND2_X1 U462 ( .A1(n429), .A2(n466), .ZN(n463) );
  OR2_X1 U463 ( .A1(n433), .A2(n465), .ZN(n466) );
  INV_X1 U464 ( .A(n432), .ZN(n465) );
  AND2_X1 U465 ( .A1(b_2_), .A2(a_1_), .ZN(n432) );
  OR2_X1 U466 ( .A1(n424), .A2(n352), .ZN(n433) );
  OR2_X1 U467 ( .A1(n350), .A2(n351), .ZN(n352) );
  INV_X1 U468 ( .A(b_2_), .ZN(n351) );
  INV_X1 U469 ( .A(n423), .ZN(n424) );
  AND2_X1 U470 ( .A1(a_3_), .A2(b_1_), .ZN(n423) );
  AND2_X1 U471 ( .A1(n467), .A2(n468), .ZN(n429) );
  OR2_X1 U472 ( .A1(n469), .A2(n470), .ZN(n468) );
  INV_X1 U473 ( .A(n471), .ZN(n467) );
  AND2_X1 U474 ( .A1(n470), .A2(n469), .ZN(n471) );
  OR2_X1 U475 ( .A1(n472), .A2(n473), .ZN(n406) );
  INV_X1 U476 ( .A(n474), .ZN(n473) );
  OR2_X1 U477 ( .A1(n475), .A2(n458), .ZN(n474) );
  AND2_X1 U478 ( .A1(n458), .A2(n475), .ZN(n472) );
  OR2_X1 U479 ( .A1(n476), .A2(n477), .ZN(n475) );
  AND3_X1 U480 ( .A1(a_2_), .A2(n478), .A3(b_0_), .ZN(n477) );
  OR2_X1 U481 ( .A1(n314), .A2(n315), .ZN(n478) );
  INV_X1 U482 ( .A(a_1_), .ZN(n315) );
  AND3_X1 U483 ( .A1(b_1_), .A2(n479), .A3(a_1_), .ZN(n476) );
  OR2_X1 U484 ( .A1(n350), .A2(n389), .ZN(n479) );
  INV_X1 U485 ( .A(b_0_), .ZN(n389) );
  AND2_X1 U486 ( .A1(n470), .A2(n459), .ZN(n458) );
  INV_X1 U487 ( .A(n469), .ZN(n459) );
  OR2_X1 U488 ( .A1(n350), .A2(n314), .ZN(n469) );
  INV_X1 U489 ( .A(b_1_), .ZN(n314) );
  INV_X1 U490 ( .A(a_2_), .ZN(n350) );
  AND2_X1 U491 ( .A1(a_3_), .A2(b_0_), .ZN(n470) );
  INV_X1 U492 ( .A(n247), .ZN(n251) );
  OR2_X1 U493 ( .A1(n354), .A2(n353), .ZN(n247) );
  INV_X1 U494 ( .A(operation_1_), .ZN(n353) );
  INV_X1 U495 ( .A(operation_0_), .ZN(n354) );
endmodule

