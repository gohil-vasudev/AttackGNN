module add_mul_mix_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        c_0_, c_1_, c_2_, c_3_, d_0_, d_1_, d_2_, d_3_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, c_0_, c_1_, c_2_, c_3_,
         d_0_, d_1_, d_2_, d_3_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227;

  XNOR2_X1 U115 ( .A(n108), .B(n109), .ZN(Result_6_) );
  NAND2_X1 U116 ( .A1(n110), .A2(n111), .ZN(n108) );
  XOR2_X1 U117 ( .A(n112), .B(n113), .Z(Result_5_) );
  XOR2_X1 U118 ( .A(n114), .B(n115), .Z(n113) );
  NOR2_X1 U119 ( .A1(n116), .A2(n117), .ZN(n115) );
  XNOR2_X1 U120 ( .A(n118), .B(n119), .ZN(Result_4_) );
  NAND2_X1 U121 ( .A1(n120), .A2(n121), .ZN(n118) );
  XOR2_X1 U122 ( .A(n122), .B(n123), .Z(Result_3_) );
  XNOR2_X1 U123 ( .A(n124), .B(n125), .ZN(Result_2_) );
  NAND2_X1 U124 ( .A1(n123), .A2(n122), .ZN(n125) );
  XOR2_X1 U125 ( .A(n126), .B(n127), .Z(Result_1_) );
  NAND2_X1 U126 ( .A1(n128), .A2(n129), .ZN(Result_0_) );
  NOR2_X1 U127 ( .A1(n130), .A2(n131), .ZN(n128) );
  NOR2_X1 U128 ( .A1(n126), .A2(n127), .ZN(n131) );
  NAND2_X1 U129 ( .A1(n132), .A2(n124), .ZN(n127) );
  AND2_X1 U130 ( .A1(n133), .A2(n134), .ZN(n124) );
  NAND2_X1 U131 ( .A1(n135), .A2(n136), .ZN(n134) );
  AND2_X1 U132 ( .A1(n122), .A2(n123), .ZN(n132) );
  XNOR2_X1 U133 ( .A(n137), .B(n138), .ZN(n123) );
  XNOR2_X1 U134 ( .A(n139), .B(n140), .ZN(n137) );
  NAND2_X1 U135 ( .A1(n120), .A2(n141), .ZN(n122) );
  NAND2_X1 U136 ( .A1(n119), .A2(n121), .ZN(n141) );
  NAND2_X1 U137 ( .A1(n142), .A2(n143), .ZN(n121) );
  NAND2_X1 U138 ( .A1(n144), .A2(n111), .ZN(n143) );
  INV_X1 U139 ( .A(n145), .ZN(n142) );
  XOR2_X1 U140 ( .A(n146), .B(n147), .Z(n119) );
  XNOR2_X1 U141 ( .A(n148), .B(n149), .ZN(n147) );
  NAND2_X1 U142 ( .A1(n150), .A2(n151), .ZN(n149) );
  NAND2_X1 U143 ( .A1(n144), .A2(n145), .ZN(n120) );
  NAND2_X1 U144 ( .A1(n152), .A2(n153), .ZN(n145) );
  NAND2_X1 U145 ( .A1(n154), .A2(n150), .ZN(n153) );
  NOR2_X1 U146 ( .A1(n155), .A2(n116), .ZN(n154) );
  NOR2_X1 U147 ( .A1(n114), .A2(n112), .ZN(n155) );
  NAND2_X1 U148 ( .A1(n114), .A2(n112), .ZN(n152) );
  XNOR2_X1 U149 ( .A(n156), .B(n157), .ZN(n112) );
  NAND2_X1 U150 ( .A1(n158), .A2(n159), .ZN(n156) );
  AND2_X1 U151 ( .A1(Result_7_), .A2(n157), .ZN(n114) );
  NOR2_X1 U152 ( .A1(n160), .A2(n161), .ZN(n157) );
  AND2_X1 U153 ( .A1(n111), .A2(n159), .ZN(Result_7_) );
  INV_X1 U154 ( .A(n116), .ZN(n111) );
  XOR2_X1 U155 ( .A(c_3_), .B(n162), .Z(n116) );
  OR2_X1 U156 ( .A1(n163), .A2(n130), .ZN(n126) );
  AND2_X1 U157 ( .A1(n164), .A2(n133), .ZN(n163) );
  NOR2_X1 U158 ( .A1(n133), .A2(n164), .ZN(n130) );
  NAND2_X1 U159 ( .A1(n129), .A2(n165), .ZN(n164) );
  NAND2_X1 U160 ( .A1(n166), .A2(n167), .ZN(n165) );
  NAND2_X1 U161 ( .A1(n168), .A2(n144), .ZN(n167) );
  INV_X1 U162 ( .A(n169), .ZN(n166) );
  NAND2_X1 U163 ( .A1(n144), .A2(n169), .ZN(n129) );
  NAND2_X1 U164 ( .A1(n170), .A2(n171), .ZN(n169) );
  NAND2_X1 U165 ( .A1(n168), .A2(n172), .ZN(n171) );
  NAND2_X1 U166 ( .A1(n173), .A2(n174), .ZN(n172) );
  NAND2_X1 U167 ( .A1(n175), .A2(n144), .ZN(n174) );
  NAND2_X1 U168 ( .A1(n150), .A2(n176), .ZN(n173) );
  OR2_X1 U169 ( .A1(n136), .A2(n135), .ZN(n133) );
  AND2_X1 U170 ( .A1(n177), .A2(n178), .ZN(n135) );
  NAND2_X1 U171 ( .A1(n140), .A2(n179), .ZN(n178) );
  NAND2_X1 U172 ( .A1(n138), .A2(n139), .ZN(n179) );
  NAND2_X1 U173 ( .A1(n180), .A2(n181), .ZN(n140) );
  NAND2_X1 U174 ( .A1(n182), .A2(n150), .ZN(n181) );
  NOR2_X1 U175 ( .A1(n183), .A2(n160), .ZN(n182) );
  INV_X1 U176 ( .A(n151), .ZN(n160) );
  NOR2_X1 U177 ( .A1(n148), .A2(n146), .ZN(n183) );
  NAND2_X1 U178 ( .A1(n148), .A2(n146), .ZN(n180) );
  XOR2_X1 U179 ( .A(n184), .B(n185), .Z(n146) );
  AND2_X1 U180 ( .A1(n185), .A2(n109), .ZN(n148) );
  AND2_X1 U181 ( .A1(n151), .A2(n159), .ZN(n109) );
  OR2_X1 U182 ( .A1(n139), .A2(n138), .ZN(n177) );
  XNOR2_X1 U183 ( .A(n186), .B(n187), .ZN(n138) );
  NAND2_X1 U184 ( .A1(n188), .A2(n189), .ZN(n186) );
  NAND2_X1 U185 ( .A1(n190), .A2(n191), .ZN(n189) );
  NAND2_X1 U186 ( .A1(n168), .A2(n110), .ZN(n190) );
  NAND2_X1 U187 ( .A1(n144), .A2(n151), .ZN(n139) );
  XNOR2_X1 U188 ( .A(n192), .B(n193), .ZN(n151) );
  XOR2_X1 U189 ( .A(d_2_), .B(c_2_), .Z(n193) );
  NAND2_X1 U190 ( .A1(c_3_), .A2(d_3_), .ZN(n192) );
  XOR2_X1 U191 ( .A(n194), .B(n195), .Z(n136) );
  NOR2_X1 U192 ( .A1(n196), .A2(n117), .ZN(n195) );
  NAND2_X1 U193 ( .A1(n170), .A2(n197), .ZN(n194) );
  NAND2_X1 U194 ( .A1(n198), .A2(n199), .ZN(n197) );
  NAND2_X1 U195 ( .A1(n158), .A2(n144), .ZN(n199) );
  INV_X1 U196 ( .A(n176), .ZN(n198) );
  NAND2_X1 U197 ( .A1(n144), .A2(n176), .ZN(n170) );
  NAND2_X1 U198 ( .A1(n187), .A2(n188), .ZN(n176) );
  NAND2_X1 U199 ( .A1(n200), .A2(n175), .ZN(n188) );
  INV_X1 U200 ( .A(n191), .ZN(n175) );
  NAND2_X1 U201 ( .A1(n150), .A2(n158), .ZN(n191) );
  INV_X1 U202 ( .A(n117), .ZN(n150) );
  XNOR2_X1 U203 ( .A(n201), .B(n202), .ZN(n117) );
  XNOR2_X1 U204 ( .A(n203), .B(a_1_), .ZN(n202) );
  NOR2_X1 U205 ( .A1(n161), .A2(n196), .ZN(n200) );
  INV_X1 U206 ( .A(n168), .ZN(n196) );
  INV_X1 U207 ( .A(n110), .ZN(n161) );
  NAND2_X1 U208 ( .A1(n184), .A2(n185), .ZN(n187) );
  AND2_X1 U209 ( .A1(n158), .A2(n110), .ZN(n185) );
  XNOR2_X1 U210 ( .A(n204), .B(n205), .ZN(n110) );
  XOR2_X1 U211 ( .A(b_2_), .B(a_2_), .Z(n205) );
  NAND2_X1 U212 ( .A1(a_3_), .A2(b_3_), .ZN(n204) );
  XOR2_X1 U213 ( .A(n206), .B(n207), .Z(n158) );
  XNOR2_X1 U214 ( .A(n208), .B(c_1_), .ZN(n207) );
  AND2_X1 U215 ( .A1(n168), .A2(n159), .ZN(n184) );
  XOR2_X1 U216 ( .A(a_3_), .B(b_3_), .Z(n159) );
  XNOR2_X1 U217 ( .A(n209), .B(n210), .ZN(n168) );
  XOR2_X1 U218 ( .A(d_0_), .B(c_0_), .Z(n210) );
  NAND2_X1 U219 ( .A1(n211), .A2(n212), .ZN(n209) );
  NAND2_X1 U220 ( .A1(n213), .A2(n208), .ZN(n212) );
  INV_X1 U221 ( .A(d_1_), .ZN(n208) );
  NAND2_X1 U222 ( .A1(c_1_), .A2(n206), .ZN(n213) );
  OR2_X1 U223 ( .A1(n206), .A2(c_1_), .ZN(n211) );
  NAND2_X1 U224 ( .A1(n214), .A2(n215), .ZN(n206) );
  NAND2_X1 U225 ( .A1(n216), .A2(c_3_), .ZN(n215) );
  NOR2_X1 U226 ( .A1(n217), .A2(n162), .ZN(n216) );
  INV_X1 U227 ( .A(d_3_), .ZN(n162) );
  NOR2_X1 U228 ( .A1(c_2_), .A2(d_2_), .ZN(n217) );
  NAND2_X1 U229 ( .A1(c_2_), .A2(d_2_), .ZN(n214) );
  XNOR2_X1 U230 ( .A(n218), .B(n219), .ZN(n144) );
  XOR2_X1 U231 ( .A(b_0_), .B(a_0_), .Z(n219) );
  NAND2_X1 U232 ( .A1(n220), .A2(n221), .ZN(n218) );
  NAND2_X1 U233 ( .A1(n222), .A2(n203), .ZN(n221) );
  INV_X1 U234 ( .A(b_1_), .ZN(n203) );
  NAND2_X1 U235 ( .A1(a_1_), .A2(n201), .ZN(n222) );
  OR2_X1 U236 ( .A1(n201), .A2(a_1_), .ZN(n220) );
  NAND2_X1 U237 ( .A1(n223), .A2(n224), .ZN(n201) );
  NAND2_X1 U238 ( .A1(n225), .A2(a_3_), .ZN(n224) );
  NOR2_X1 U239 ( .A1(n226), .A2(n227), .ZN(n225) );
  INV_X1 U240 ( .A(b_3_), .ZN(n227) );
  NOR2_X1 U241 ( .A1(a_2_), .A2(b_2_), .ZN(n226) );
  NAND2_X1 U242 ( .A1(a_2_), .A2(b_2_), .ZN(n223) );
endmodule

