module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n500_, new_n898_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n903_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n878_, new_n543_, new_n113_, new_n924_, new_n886_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n914_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n918_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n897_, new_n379_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n302_, new_n191_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, keyIn_0_24 );
not g001 ( new_n107_, keyIn_0_5 );
not g002 ( new_n108_, N81 );
or g003 ( new_n109_, new_n108_, N85 );
not g004 ( new_n110_, N85 );
or g005 ( new_n111_, new_n110_, N81 );
and g006 ( new_n112_, new_n109_, new_n111_ );
not g007 ( new_n113_, N93 );
and g008 ( new_n114_, new_n113_, N89 );
not g009 ( new_n115_, N89 );
and g010 ( new_n116_, new_n115_, N93 );
or g011 ( new_n117_, new_n114_, new_n116_ );
or g012 ( new_n118_, new_n117_, new_n112_ );
and g013 ( new_n119_, new_n110_, N81 );
and g014 ( new_n120_, new_n108_, N85 );
or g015 ( new_n121_, new_n119_, new_n120_ );
or g016 ( new_n122_, new_n115_, N93 );
or g017 ( new_n123_, new_n113_, N89 );
and g018 ( new_n124_, new_n122_, new_n123_ );
or g019 ( new_n125_, new_n121_, new_n124_ );
and g020 ( new_n126_, new_n118_, new_n125_ );
or g021 ( new_n127_, new_n126_, new_n107_ );
and g022 ( new_n128_, new_n121_, new_n124_ );
and g023 ( new_n129_, new_n117_, new_n112_ );
or g024 ( new_n130_, new_n128_, new_n129_ );
or g025 ( new_n131_, new_n130_, keyIn_0_5 );
and g026 ( new_n132_, new_n131_, new_n127_ );
not g027 ( new_n133_, keyIn_0_4 );
not g028 ( new_n134_, N77 );
and g029 ( new_n135_, new_n134_, N73 );
not g030 ( new_n136_, N73 );
and g031 ( new_n137_, new_n136_, N77 );
or g032 ( new_n138_, new_n135_, new_n137_ );
and g033 ( new_n139_, N65, N69 );
not g034 ( new_n140_, N65 );
not g035 ( new_n141_, N69 );
and g036 ( new_n142_, new_n140_, new_n141_ );
or g037 ( new_n143_, new_n142_, new_n139_ );
and g038 ( new_n144_, new_n138_, new_n143_ );
or g039 ( new_n145_, new_n136_, N77 );
or g040 ( new_n146_, new_n134_, N73 );
and g041 ( new_n147_, new_n145_, new_n146_ );
not g042 ( new_n148_, new_n139_ );
or g043 ( new_n149_, N65, N69 );
and g044 ( new_n150_, new_n148_, new_n149_ );
and g045 ( new_n151_, new_n147_, new_n150_ );
or g046 ( new_n152_, new_n144_, new_n151_ );
and g047 ( new_n153_, new_n152_, new_n133_ );
or g048 ( new_n154_, new_n147_, new_n150_ );
or g049 ( new_n155_, new_n138_, new_n143_ );
and g050 ( new_n156_, new_n155_, new_n154_ );
and g051 ( new_n157_, new_n156_, keyIn_0_4 );
or g052 ( new_n158_, new_n153_, new_n157_ );
or g053 ( new_n159_, new_n158_, new_n132_ );
and g054 ( new_n160_, new_n130_, keyIn_0_5 );
and g055 ( new_n161_, new_n126_, new_n107_ );
or g056 ( new_n162_, new_n160_, new_n161_ );
or g057 ( new_n163_, new_n156_, keyIn_0_4 );
or g058 ( new_n164_, new_n152_, new_n133_ );
and g059 ( new_n165_, new_n163_, new_n164_ );
or g060 ( new_n166_, new_n162_, new_n165_ );
and g061 ( new_n167_, new_n159_, new_n166_ );
or g062 ( new_n168_, new_n167_, keyIn_0_20 );
not g063 ( new_n169_, keyIn_0_20 );
and g064 ( new_n170_, new_n162_, new_n165_ );
and g065 ( new_n171_, new_n158_, new_n132_ );
or g066 ( new_n172_, new_n170_, new_n171_ );
or g067 ( new_n173_, new_n172_, new_n169_ );
and g068 ( new_n174_, new_n173_, new_n168_ );
and g069 ( new_n175_, N129, N137 );
not g070 ( new_n176_, new_n175_ );
or g071 ( new_n177_, new_n174_, new_n176_ );
and g072 ( new_n178_, new_n172_, new_n169_ );
and g073 ( new_n179_, new_n167_, keyIn_0_20 );
or g074 ( new_n180_, new_n178_, new_n179_ );
or g075 ( new_n181_, new_n180_, new_n175_ );
and g076 ( new_n182_, new_n181_, new_n177_ );
or g077 ( new_n183_, new_n182_, new_n106_ );
and g078 ( new_n184_, new_n180_, new_n175_ );
and g079 ( new_n185_, new_n174_, new_n176_ );
or g080 ( new_n186_, new_n184_, new_n185_ );
or g081 ( new_n187_, new_n186_, keyIn_0_24 );
and g082 ( new_n188_, new_n187_, new_n183_ );
not g083 ( new_n189_, keyIn_0_8 );
not g084 ( new_n190_, N17 );
and g085 ( new_n191_, new_n190_, N1 );
not g086 ( new_n192_, N1 );
and g087 ( new_n193_, new_n192_, N17 );
or g088 ( new_n194_, new_n191_, new_n193_ );
and g089 ( new_n195_, N33, N49 );
not g090 ( new_n196_, N33 );
not g091 ( new_n197_, N49 );
and g092 ( new_n198_, new_n196_, new_n197_ );
or g093 ( new_n199_, new_n198_, new_n195_ );
and g094 ( new_n200_, new_n194_, new_n199_ );
not g095 ( new_n201_, new_n200_ );
or g096 ( new_n202_, new_n194_, new_n199_ );
and g097 ( new_n203_, new_n201_, new_n202_ );
not g098 ( new_n204_, new_n203_ );
and g099 ( new_n205_, new_n204_, new_n189_ );
and g100 ( new_n206_, new_n203_, keyIn_0_8 );
or g101 ( new_n207_, new_n205_, new_n206_ );
not g102 ( new_n208_, new_n207_ );
or g103 ( new_n209_, new_n188_, new_n208_ );
and g104 ( new_n210_, new_n186_, keyIn_0_24 );
and g105 ( new_n211_, new_n182_, new_n106_ );
or g106 ( new_n212_, new_n210_, new_n211_ );
or g107 ( new_n213_, new_n212_, new_n207_ );
and g108 ( new_n214_, new_n213_, new_n209_ );
not g109 ( new_n215_, new_n214_ );
not g110 ( new_n216_, keyIn_0_25 );
not g111 ( new_n217_, keyIn_0_7 );
not g112 ( new_n218_, N117 );
and g113 ( new_n219_, new_n218_, N113 );
not g114 ( new_n220_, N113 );
and g115 ( new_n221_, new_n220_, N117 );
or g116 ( new_n222_, new_n219_, new_n221_ );
not g117 ( new_n223_, N125 );
and g118 ( new_n224_, new_n223_, N121 );
not g119 ( new_n225_, N121 );
and g120 ( new_n226_, new_n225_, N125 );
or g121 ( new_n227_, new_n224_, new_n226_ );
or g122 ( new_n228_, new_n222_, new_n227_ );
or g123 ( new_n229_, new_n220_, N117 );
or g124 ( new_n230_, new_n218_, N113 );
and g125 ( new_n231_, new_n229_, new_n230_ );
or g126 ( new_n232_, new_n225_, N125 );
or g127 ( new_n233_, new_n223_, N121 );
and g128 ( new_n234_, new_n232_, new_n233_ );
or g129 ( new_n235_, new_n231_, new_n234_ );
and g130 ( new_n236_, new_n228_, new_n235_ );
and g131 ( new_n237_, new_n236_, new_n217_ );
and g132 ( new_n238_, new_n231_, new_n234_ );
and g133 ( new_n239_, new_n222_, new_n227_ );
or g134 ( new_n240_, new_n239_, new_n238_ );
and g135 ( new_n241_, new_n240_, keyIn_0_7 );
or g136 ( new_n242_, new_n237_, new_n241_ );
not g137 ( new_n243_, keyIn_0_6 );
not g138 ( new_n244_, N101 );
and g139 ( new_n245_, new_n244_, N97 );
not g140 ( new_n246_, N97 );
and g141 ( new_n247_, new_n246_, N101 );
or g142 ( new_n248_, new_n245_, new_n247_ );
not g143 ( new_n249_, N109 );
and g144 ( new_n250_, new_n249_, N105 );
not g145 ( new_n251_, N105 );
and g146 ( new_n252_, new_n251_, N109 );
or g147 ( new_n253_, new_n250_, new_n252_ );
and g148 ( new_n254_, new_n248_, new_n253_ );
or g149 ( new_n255_, new_n246_, N101 );
or g150 ( new_n256_, new_n244_, N97 );
and g151 ( new_n257_, new_n255_, new_n256_ );
or g152 ( new_n258_, new_n251_, N109 );
or g153 ( new_n259_, new_n249_, N105 );
and g154 ( new_n260_, new_n258_, new_n259_ );
and g155 ( new_n261_, new_n257_, new_n260_ );
or g156 ( new_n262_, new_n254_, new_n261_ );
and g157 ( new_n263_, new_n262_, new_n243_ );
or g158 ( new_n264_, new_n257_, new_n260_ );
or g159 ( new_n265_, new_n248_, new_n253_ );
and g160 ( new_n266_, new_n265_, new_n264_ );
and g161 ( new_n267_, new_n266_, keyIn_0_6 );
or g162 ( new_n268_, new_n267_, new_n263_ );
and g163 ( new_n269_, new_n242_, new_n268_ );
or g164 ( new_n270_, new_n240_, keyIn_0_7 );
or g165 ( new_n271_, new_n236_, new_n217_ );
and g166 ( new_n272_, new_n271_, new_n270_ );
or g167 ( new_n273_, new_n266_, keyIn_0_6 );
or g168 ( new_n274_, new_n262_, new_n243_ );
and g169 ( new_n275_, new_n273_, new_n274_ );
and g170 ( new_n276_, new_n272_, new_n275_ );
or g171 ( new_n277_, new_n269_, new_n276_ );
and g172 ( new_n278_, new_n277_, keyIn_0_21 );
not g173 ( new_n279_, keyIn_0_21 );
or g174 ( new_n280_, new_n272_, new_n275_ );
or g175 ( new_n281_, new_n242_, new_n268_ );
and g176 ( new_n282_, new_n281_, new_n280_ );
and g177 ( new_n283_, new_n282_, new_n279_ );
or g178 ( new_n284_, new_n283_, new_n278_ );
and g179 ( new_n285_, N130, N137 );
not g180 ( new_n286_, new_n285_ );
and g181 ( new_n287_, new_n284_, new_n286_ );
or g182 ( new_n288_, new_n282_, new_n279_ );
or g183 ( new_n289_, new_n277_, keyIn_0_21 );
and g184 ( new_n290_, new_n288_, new_n289_ );
and g185 ( new_n291_, new_n290_, new_n285_ );
or g186 ( new_n292_, new_n287_, new_n291_ );
and g187 ( new_n293_, new_n292_, new_n216_ );
or g188 ( new_n294_, new_n290_, new_n285_ );
or g189 ( new_n295_, new_n284_, new_n286_ );
and g190 ( new_n296_, new_n295_, new_n294_ );
and g191 ( new_n297_, new_n296_, keyIn_0_25 );
or g192 ( new_n298_, new_n293_, new_n297_ );
not g193 ( new_n299_, N21 );
and g194 ( new_n300_, new_n299_, N5 );
not g195 ( new_n301_, N5 );
and g196 ( new_n302_, new_n301_, N21 );
or g197 ( new_n303_, new_n300_, new_n302_ );
and g198 ( new_n304_, N37, N53 );
not g199 ( new_n305_, N37 );
not g200 ( new_n306_, N53 );
and g201 ( new_n307_, new_n305_, new_n306_ );
or g202 ( new_n308_, new_n307_, new_n304_ );
and g203 ( new_n309_, new_n303_, new_n308_ );
not g204 ( new_n310_, new_n309_ );
or g205 ( new_n311_, new_n303_, new_n308_ );
and g206 ( new_n312_, new_n310_, new_n311_ );
not g207 ( new_n313_, new_n312_ );
and g208 ( new_n314_, new_n313_, keyIn_0_9 );
not g209 ( new_n315_, new_n314_ );
or g210 ( new_n316_, new_n313_, keyIn_0_9 );
and g211 ( new_n317_, new_n315_, new_n316_ );
and g212 ( new_n318_, new_n298_, new_n317_ );
or g213 ( new_n319_, new_n296_, keyIn_0_25 );
or g214 ( new_n320_, new_n292_, new_n216_ );
and g215 ( new_n321_, new_n320_, new_n319_ );
not g216 ( new_n322_, new_n317_ );
and g217 ( new_n323_, new_n321_, new_n322_ );
or g218 ( new_n324_, new_n318_, new_n323_ );
and g219 ( new_n325_, new_n215_, new_n324_ );
not g220 ( new_n326_, keyIn_0_23 );
or g221 ( new_n327_, new_n162_, new_n272_ );
or g222 ( new_n328_, new_n242_, new_n132_ );
and g223 ( new_n329_, new_n327_, new_n328_ );
or g224 ( new_n330_, new_n329_, new_n326_ );
and g225 ( new_n331_, new_n242_, new_n132_ );
and g226 ( new_n332_, new_n162_, new_n272_ );
or g227 ( new_n333_, new_n331_, new_n332_ );
or g228 ( new_n334_, new_n333_, keyIn_0_23 );
and g229 ( new_n335_, new_n334_, new_n330_ );
and g230 ( new_n336_, N132, N137 );
or g231 ( new_n337_, new_n335_, new_n336_ );
and g232 ( new_n338_, new_n333_, keyIn_0_23 );
and g233 ( new_n339_, new_n329_, new_n326_ );
or g234 ( new_n340_, new_n338_, new_n339_ );
not g235 ( new_n341_, new_n336_ );
or g236 ( new_n342_, new_n340_, new_n341_ );
and g237 ( new_n343_, new_n342_, new_n337_ );
or g238 ( new_n344_, new_n343_, keyIn_0_27 );
not g239 ( new_n345_, keyIn_0_27 );
and g240 ( new_n346_, new_n340_, new_n341_ );
and g241 ( new_n347_, new_n335_, new_n336_ );
or g242 ( new_n348_, new_n346_, new_n347_ );
or g243 ( new_n349_, new_n348_, new_n345_ );
and g244 ( new_n350_, new_n349_, new_n344_ );
not g245 ( new_n351_, N29 );
and g246 ( new_n352_, new_n351_, N13 );
not g247 ( new_n353_, N13 );
and g248 ( new_n354_, new_n353_, N29 );
or g249 ( new_n355_, new_n352_, new_n354_ );
and g250 ( new_n356_, N45, N61 );
not g251 ( new_n357_, N45 );
not g252 ( new_n358_, N61 );
and g253 ( new_n359_, new_n357_, new_n358_ );
or g254 ( new_n360_, new_n359_, new_n356_ );
and g255 ( new_n361_, new_n355_, new_n360_ );
not g256 ( new_n362_, new_n361_ );
or g257 ( new_n363_, new_n355_, new_n360_ );
and g258 ( new_n364_, new_n362_, new_n363_ );
not g259 ( new_n365_, new_n364_ );
and g260 ( new_n366_, new_n365_, keyIn_0_11 );
not g261 ( new_n367_, new_n366_ );
or g262 ( new_n368_, new_n365_, keyIn_0_11 );
and g263 ( new_n369_, new_n367_, new_n368_ );
not g264 ( new_n370_, new_n369_ );
or g265 ( new_n371_, new_n350_, new_n370_ );
and g266 ( new_n372_, new_n348_, new_n345_ );
and g267 ( new_n373_, new_n343_, keyIn_0_27 );
or g268 ( new_n374_, new_n372_, new_n373_ );
or g269 ( new_n375_, new_n374_, new_n369_ );
and g270 ( new_n376_, new_n375_, new_n371_ );
not g271 ( new_n377_, keyIn_0_26 );
or g272 ( new_n378_, new_n275_, new_n165_ );
or g273 ( new_n379_, new_n268_, new_n158_ );
and g274 ( new_n380_, new_n379_, new_n378_ );
or g275 ( new_n381_, new_n380_, keyIn_0_22 );
not g276 ( new_n382_, keyIn_0_22 );
and g277 ( new_n383_, new_n268_, new_n158_ );
and g278 ( new_n384_, new_n275_, new_n165_ );
or g279 ( new_n385_, new_n383_, new_n384_ );
or g280 ( new_n386_, new_n385_, new_n382_ );
and g281 ( new_n387_, new_n381_, new_n386_ );
and g282 ( new_n388_, N131, N137 );
not g283 ( new_n389_, new_n388_ );
or g284 ( new_n390_, new_n387_, new_n389_ );
and g285 ( new_n391_, new_n385_, new_n382_ );
and g286 ( new_n392_, new_n380_, keyIn_0_22 );
or g287 ( new_n393_, new_n392_, new_n391_ );
or g288 ( new_n394_, new_n393_, new_n388_ );
and g289 ( new_n395_, new_n394_, new_n390_ );
or g290 ( new_n396_, new_n395_, new_n377_ );
and g291 ( new_n397_, new_n393_, new_n388_ );
and g292 ( new_n398_, new_n387_, new_n389_ );
or g293 ( new_n399_, new_n397_, new_n398_ );
or g294 ( new_n400_, new_n399_, keyIn_0_26 );
and g295 ( new_n401_, new_n400_, new_n396_ );
not g296 ( new_n402_, keyIn_0_10 );
not g297 ( new_n403_, N25 );
and g298 ( new_n404_, new_n403_, N9 );
not g299 ( new_n405_, N9 );
and g300 ( new_n406_, new_n405_, N25 );
or g301 ( new_n407_, new_n404_, new_n406_ );
and g302 ( new_n408_, N41, N57 );
not g303 ( new_n409_, N41 );
not g304 ( new_n410_, N57 );
and g305 ( new_n411_, new_n409_, new_n410_ );
or g306 ( new_n412_, new_n411_, new_n408_ );
and g307 ( new_n413_, new_n407_, new_n412_ );
not g308 ( new_n414_, new_n413_ );
or g309 ( new_n415_, new_n407_, new_n412_ );
and g310 ( new_n416_, new_n414_, new_n415_ );
not g311 ( new_n417_, new_n416_ );
and g312 ( new_n418_, new_n417_, new_n402_ );
and g313 ( new_n419_, new_n416_, keyIn_0_10 );
or g314 ( new_n420_, new_n418_, new_n419_ );
or g315 ( new_n421_, new_n401_, new_n420_ );
and g316 ( new_n422_, new_n399_, keyIn_0_26 );
and g317 ( new_n423_, new_n395_, new_n377_ );
or g318 ( new_n424_, new_n422_, new_n423_ );
not g319 ( new_n425_, new_n420_ );
or g320 ( new_n426_, new_n424_, new_n425_ );
and g321 ( new_n427_, new_n426_, new_n421_ );
and g322 ( new_n428_, new_n376_, new_n427_ );
and g323 ( new_n429_, new_n325_, new_n428_ );
not g324 ( new_n430_, keyIn_0_16 );
and g325 ( new_n431_, new_n301_, N1 );
and g326 ( new_n432_, new_n192_, N5 );
or g327 ( new_n433_, new_n431_, new_n432_ );
and g328 ( new_n434_, new_n353_, N9 );
and g329 ( new_n435_, new_n405_, N13 );
or g330 ( new_n436_, new_n434_, new_n435_ );
and g331 ( new_n437_, new_n433_, new_n436_ );
or g332 ( new_n438_, new_n192_, N5 );
or g333 ( new_n439_, new_n301_, N1 );
and g334 ( new_n440_, new_n438_, new_n439_ );
or g335 ( new_n441_, new_n405_, N13 );
or g336 ( new_n442_, new_n353_, N9 );
and g337 ( new_n443_, new_n441_, new_n442_ );
and g338 ( new_n444_, new_n440_, new_n443_ );
or g339 ( new_n445_, new_n437_, new_n444_ );
and g340 ( new_n446_, new_n445_, keyIn_0_0 );
not g341 ( new_n447_, keyIn_0_0 );
or g342 ( new_n448_, new_n440_, new_n443_ );
or g343 ( new_n449_, new_n433_, new_n436_ );
and g344 ( new_n450_, new_n449_, new_n448_ );
and g345 ( new_n451_, new_n450_, new_n447_ );
or g346 ( new_n452_, new_n451_, new_n446_ );
not g347 ( new_n453_, keyIn_0_1 );
and g348 ( new_n454_, new_n299_, N17 );
and g349 ( new_n455_, new_n190_, N21 );
or g350 ( new_n456_, new_n454_, new_n455_ );
and g351 ( new_n457_, new_n351_, N25 );
and g352 ( new_n458_, new_n403_, N29 );
or g353 ( new_n459_, new_n457_, new_n458_ );
or g354 ( new_n460_, new_n456_, new_n459_ );
or g355 ( new_n461_, new_n190_, N21 );
or g356 ( new_n462_, new_n299_, N17 );
and g357 ( new_n463_, new_n461_, new_n462_ );
or g358 ( new_n464_, new_n403_, N29 );
or g359 ( new_n465_, new_n351_, N25 );
and g360 ( new_n466_, new_n464_, new_n465_ );
or g361 ( new_n467_, new_n463_, new_n466_ );
and g362 ( new_n468_, new_n460_, new_n467_ );
and g363 ( new_n469_, new_n468_, new_n453_ );
and g364 ( new_n470_, new_n463_, new_n466_ );
and g365 ( new_n471_, new_n456_, new_n459_ );
or g366 ( new_n472_, new_n471_, new_n470_ );
and g367 ( new_n473_, new_n472_, keyIn_0_1 );
or g368 ( new_n474_, new_n469_, new_n473_ );
and g369 ( new_n475_, new_n452_, new_n474_ );
or g370 ( new_n476_, new_n450_, new_n447_ );
or g371 ( new_n477_, new_n445_, keyIn_0_0 );
and g372 ( new_n478_, new_n476_, new_n477_ );
or g373 ( new_n479_, new_n472_, keyIn_0_1 );
or g374 ( new_n480_, new_n468_, new_n453_ );
and g375 ( new_n481_, new_n480_, new_n479_ );
and g376 ( new_n482_, new_n478_, new_n481_ );
or g377 ( new_n483_, new_n475_, new_n482_ );
and g378 ( new_n484_, new_n483_, new_n430_ );
or g379 ( new_n485_, new_n478_, new_n481_ );
or g380 ( new_n486_, new_n452_, new_n474_ );
and g381 ( new_n487_, new_n486_, new_n485_ );
and g382 ( new_n488_, new_n487_, keyIn_0_16 );
or g383 ( new_n489_, new_n488_, new_n484_ );
and g384 ( new_n490_, N133, N137 );
and g385 ( new_n491_, new_n489_, new_n490_ );
or g386 ( new_n492_, new_n487_, keyIn_0_16 );
or g387 ( new_n493_, new_n483_, new_n430_ );
and g388 ( new_n494_, new_n492_, new_n493_ );
not g389 ( new_n495_, new_n490_ );
and g390 ( new_n496_, new_n494_, new_n495_ );
or g391 ( new_n497_, new_n491_, new_n496_ );
and g392 ( new_n498_, new_n497_, keyIn_0_28 );
not g393 ( new_n499_, keyIn_0_28 );
or g394 ( new_n500_, new_n494_, new_n495_ );
or g395 ( new_n501_, new_n489_, new_n490_ );
and g396 ( new_n502_, new_n501_, new_n500_ );
and g397 ( new_n503_, new_n502_, new_n499_ );
or g398 ( new_n504_, new_n498_, new_n503_ );
and g399 ( new_n505_, new_n108_, N65 );
and g400 ( new_n506_, new_n140_, N81 );
or g401 ( new_n507_, new_n505_, new_n506_ );
and g402 ( new_n508_, N97, N113 );
and g403 ( new_n509_, new_n246_, new_n220_ );
or g404 ( new_n510_, new_n509_, new_n508_ );
and g405 ( new_n511_, new_n507_, new_n510_ );
not g406 ( new_n512_, new_n511_ );
or g407 ( new_n513_, new_n507_, new_n510_ );
and g408 ( new_n514_, new_n512_, new_n513_ );
not g409 ( new_n515_, new_n514_ );
and g410 ( new_n516_, new_n515_, keyIn_0_12 );
not g411 ( new_n517_, new_n516_ );
or g412 ( new_n518_, new_n515_, keyIn_0_12 );
and g413 ( new_n519_, new_n517_, new_n518_ );
and g414 ( new_n520_, new_n504_, new_n519_ );
or g415 ( new_n521_, new_n502_, new_n499_ );
or g416 ( new_n522_, new_n497_, keyIn_0_28 );
and g417 ( new_n523_, new_n522_, new_n521_ );
not g418 ( new_n524_, new_n519_ );
and g419 ( new_n525_, new_n523_, new_n524_ );
or g420 ( new_n526_, new_n520_, new_n525_ );
not g421 ( new_n527_, keyIn_0_2 );
and g422 ( new_n528_, new_n357_, N41 );
and g423 ( new_n529_, new_n409_, N45 );
or g424 ( new_n530_, new_n528_, new_n529_ );
and g425 ( new_n531_, N33, N37 );
and g426 ( new_n532_, new_n196_, new_n305_ );
or g427 ( new_n533_, new_n532_, new_n531_ );
and g428 ( new_n534_, new_n530_, new_n533_ );
or g429 ( new_n535_, new_n409_, N45 );
or g430 ( new_n536_, new_n357_, N41 );
and g431 ( new_n537_, new_n535_, new_n536_ );
not g432 ( new_n538_, new_n531_ );
or g433 ( new_n539_, N33, N37 );
and g434 ( new_n540_, new_n538_, new_n539_ );
and g435 ( new_n541_, new_n537_, new_n540_ );
or g436 ( new_n542_, new_n534_, new_n541_ );
and g437 ( new_n543_, new_n542_, new_n527_ );
or g438 ( new_n544_, new_n537_, new_n540_ );
or g439 ( new_n545_, new_n530_, new_n533_ );
and g440 ( new_n546_, new_n545_, new_n544_ );
and g441 ( new_n547_, new_n546_, keyIn_0_2 );
or g442 ( new_n548_, new_n543_, new_n547_ );
not g443 ( new_n549_, keyIn_0_3 );
and g444 ( new_n550_, new_n306_, N49 );
and g445 ( new_n551_, new_n197_, N53 );
or g446 ( new_n552_, new_n550_, new_n551_ );
and g447 ( new_n553_, new_n358_, N57 );
and g448 ( new_n554_, new_n410_, N61 );
or g449 ( new_n555_, new_n553_, new_n554_ );
and g450 ( new_n556_, new_n552_, new_n555_ );
or g451 ( new_n557_, new_n197_, N53 );
or g452 ( new_n558_, new_n306_, N49 );
and g453 ( new_n559_, new_n557_, new_n558_ );
or g454 ( new_n560_, new_n410_, N61 );
or g455 ( new_n561_, new_n358_, N57 );
and g456 ( new_n562_, new_n560_, new_n561_ );
and g457 ( new_n563_, new_n559_, new_n562_ );
or g458 ( new_n564_, new_n556_, new_n563_ );
and g459 ( new_n565_, new_n564_, new_n549_ );
or g460 ( new_n566_, new_n559_, new_n562_ );
or g461 ( new_n567_, new_n552_, new_n555_ );
and g462 ( new_n568_, new_n567_, new_n566_ );
and g463 ( new_n569_, new_n568_, keyIn_0_3 );
or g464 ( new_n570_, new_n569_, new_n565_ );
and g465 ( new_n571_, new_n570_, new_n548_ );
or g466 ( new_n572_, new_n546_, keyIn_0_2 );
or g467 ( new_n573_, new_n542_, new_n527_ );
and g468 ( new_n574_, new_n572_, new_n573_ );
or g469 ( new_n575_, new_n568_, keyIn_0_3 );
or g470 ( new_n576_, new_n564_, new_n549_ );
and g471 ( new_n577_, new_n575_, new_n576_ );
and g472 ( new_n578_, new_n577_, new_n574_ );
or g473 ( new_n579_, new_n571_, new_n578_ );
and g474 ( new_n580_, new_n579_, keyIn_0_17 );
not g475 ( new_n581_, keyIn_0_17 );
or g476 ( new_n582_, new_n577_, new_n574_ );
or g477 ( new_n583_, new_n570_, new_n548_ );
and g478 ( new_n584_, new_n583_, new_n582_ );
and g479 ( new_n585_, new_n584_, new_n581_ );
or g480 ( new_n586_, new_n585_, new_n580_ );
and g481 ( new_n587_, N134, N137 );
not g482 ( new_n588_, new_n587_ );
and g483 ( new_n589_, new_n586_, new_n588_ );
or g484 ( new_n590_, new_n584_, new_n581_ );
or g485 ( new_n591_, new_n579_, keyIn_0_17 );
and g486 ( new_n592_, new_n590_, new_n591_ );
and g487 ( new_n593_, new_n592_, new_n587_ );
or g488 ( new_n594_, new_n589_, new_n593_ );
and g489 ( new_n595_, new_n594_, keyIn_0_29 );
not g490 ( new_n596_, keyIn_0_29 );
or g491 ( new_n597_, new_n592_, new_n587_ );
or g492 ( new_n598_, new_n586_, new_n588_ );
and g493 ( new_n599_, new_n598_, new_n597_ );
and g494 ( new_n600_, new_n599_, new_n596_ );
or g495 ( new_n601_, new_n595_, new_n600_ );
and g496 ( new_n602_, new_n110_, N69 );
and g497 ( new_n603_, new_n141_, N85 );
or g498 ( new_n604_, new_n602_, new_n603_ );
and g499 ( new_n605_, N101, N117 );
and g500 ( new_n606_, new_n244_, new_n218_ );
or g501 ( new_n607_, new_n606_, new_n605_ );
and g502 ( new_n608_, new_n604_, new_n607_ );
not g503 ( new_n609_, new_n608_ );
or g504 ( new_n610_, new_n604_, new_n607_ );
and g505 ( new_n611_, new_n609_, new_n610_ );
not g506 ( new_n612_, new_n611_ );
and g507 ( new_n613_, new_n612_, keyIn_0_13 );
not g508 ( new_n614_, new_n613_ );
or g509 ( new_n615_, new_n612_, keyIn_0_13 );
and g510 ( new_n616_, new_n614_, new_n615_ );
and g511 ( new_n617_, new_n601_, new_n616_ );
or g512 ( new_n618_, new_n599_, new_n596_ );
or g513 ( new_n619_, new_n594_, keyIn_0_29 );
and g514 ( new_n620_, new_n619_, new_n618_ );
not g515 ( new_n621_, new_n616_ );
and g516 ( new_n622_, new_n620_, new_n621_ );
or g517 ( new_n623_, new_n617_, new_n622_ );
and g518 ( new_n624_, new_n526_, new_n623_ );
and g519 ( new_n625_, new_n452_, new_n574_ );
and g520 ( new_n626_, new_n548_, new_n478_ );
or g521 ( new_n627_, new_n625_, new_n626_ );
and g522 ( new_n628_, new_n627_, keyIn_0_18 );
not g523 ( new_n629_, keyIn_0_18 );
or g524 ( new_n630_, new_n548_, new_n478_ );
or g525 ( new_n631_, new_n452_, new_n574_ );
and g526 ( new_n632_, new_n630_, new_n631_ );
and g527 ( new_n633_, new_n632_, new_n629_ );
or g528 ( new_n634_, new_n628_, new_n633_ );
and g529 ( new_n635_, N135, N137 );
and g530 ( new_n636_, new_n634_, new_n635_ );
or g531 ( new_n637_, new_n632_, new_n629_ );
or g532 ( new_n638_, new_n627_, keyIn_0_18 );
and g533 ( new_n639_, new_n638_, new_n637_ );
not g534 ( new_n640_, new_n635_ );
and g535 ( new_n641_, new_n639_, new_n640_ );
or g536 ( new_n642_, new_n636_, new_n641_ );
and g537 ( new_n643_, new_n642_, keyIn_0_30 );
not g538 ( new_n644_, keyIn_0_30 );
or g539 ( new_n645_, new_n639_, new_n640_ );
or g540 ( new_n646_, new_n634_, new_n635_ );
and g541 ( new_n647_, new_n646_, new_n645_ );
and g542 ( new_n648_, new_n647_, new_n644_ );
or g543 ( new_n649_, new_n643_, new_n648_ );
not g544 ( new_n650_, keyIn_0_14 );
and g545 ( new_n651_, new_n115_, N73 );
and g546 ( new_n652_, new_n136_, N89 );
or g547 ( new_n653_, new_n651_, new_n652_ );
and g548 ( new_n654_, N105, N121 );
and g549 ( new_n655_, new_n251_, new_n225_ );
or g550 ( new_n656_, new_n655_, new_n654_ );
and g551 ( new_n657_, new_n653_, new_n656_ );
not g552 ( new_n658_, new_n657_ );
or g553 ( new_n659_, new_n653_, new_n656_ );
and g554 ( new_n660_, new_n658_, new_n659_ );
not g555 ( new_n661_, new_n660_ );
and g556 ( new_n662_, new_n661_, new_n650_ );
and g557 ( new_n663_, new_n660_, keyIn_0_14 );
or g558 ( new_n664_, new_n662_, new_n663_ );
and g559 ( new_n665_, new_n649_, new_n664_ );
or g560 ( new_n666_, new_n647_, new_n644_ );
or g561 ( new_n667_, new_n642_, keyIn_0_30 );
and g562 ( new_n668_, new_n667_, new_n666_ );
not g563 ( new_n669_, new_n664_ );
and g564 ( new_n670_, new_n668_, new_n669_ );
or g565 ( new_n671_, new_n665_, new_n670_ );
not g566 ( new_n672_, keyIn_0_31 );
not g567 ( new_n673_, keyIn_0_19 );
or g568 ( new_n674_, new_n570_, new_n481_ );
or g569 ( new_n675_, new_n474_, new_n577_ );
and g570 ( new_n676_, new_n674_, new_n675_ );
or g571 ( new_n677_, new_n676_, new_n673_ );
and g572 ( new_n678_, new_n474_, new_n577_ );
and g573 ( new_n679_, new_n570_, new_n481_ );
or g574 ( new_n680_, new_n678_, new_n679_ );
or g575 ( new_n681_, new_n680_, keyIn_0_19 );
and g576 ( new_n682_, new_n681_, new_n677_ );
and g577 ( new_n683_, N136, N137 );
or g578 ( new_n684_, new_n682_, new_n683_ );
and g579 ( new_n685_, new_n680_, keyIn_0_19 );
and g580 ( new_n686_, new_n676_, new_n673_ );
or g581 ( new_n687_, new_n685_, new_n686_ );
not g582 ( new_n688_, new_n683_ );
or g583 ( new_n689_, new_n687_, new_n688_ );
and g584 ( new_n690_, new_n689_, new_n684_ );
or g585 ( new_n691_, new_n690_, new_n672_ );
and g586 ( new_n692_, new_n687_, new_n688_ );
and g587 ( new_n693_, new_n682_, new_n683_ );
or g588 ( new_n694_, new_n692_, new_n693_ );
or g589 ( new_n695_, new_n694_, keyIn_0_31 );
and g590 ( new_n696_, new_n695_, new_n691_ );
not g591 ( new_n697_, keyIn_0_15 );
and g592 ( new_n698_, new_n113_, N77 );
and g593 ( new_n699_, new_n134_, N93 );
or g594 ( new_n700_, new_n698_, new_n699_ );
and g595 ( new_n701_, N109, N125 );
and g596 ( new_n702_, new_n249_, new_n223_ );
or g597 ( new_n703_, new_n702_, new_n701_ );
and g598 ( new_n704_, new_n700_, new_n703_ );
not g599 ( new_n705_, new_n704_ );
or g600 ( new_n706_, new_n700_, new_n703_ );
and g601 ( new_n707_, new_n705_, new_n706_ );
not g602 ( new_n708_, new_n707_ );
and g603 ( new_n709_, new_n708_, new_n697_ );
and g604 ( new_n710_, new_n707_, keyIn_0_15 );
or g605 ( new_n711_, new_n709_, new_n710_ );
or g606 ( new_n712_, new_n696_, new_n711_ );
and g607 ( new_n713_, new_n694_, keyIn_0_31 );
and g608 ( new_n714_, new_n690_, new_n672_ );
or g609 ( new_n715_, new_n713_, new_n714_ );
not g610 ( new_n716_, new_n711_ );
or g611 ( new_n717_, new_n715_, new_n716_ );
and g612 ( new_n718_, new_n717_, new_n712_ );
and g613 ( new_n719_, new_n671_, new_n718_ );
and g614 ( new_n720_, new_n624_, new_n719_ );
and g615 ( new_n721_, new_n429_, new_n720_ );
not g616 ( new_n722_, new_n721_ );
and g617 ( new_n723_, new_n722_, N1 );
and g618 ( new_n724_, new_n721_, new_n192_ );
or g619 ( N724, new_n723_, new_n724_ );
or g620 ( new_n726_, new_n321_, new_n322_ );
or g621 ( new_n727_, new_n298_, new_n317_ );
and g622 ( new_n728_, new_n727_, new_n726_ );
and g623 ( new_n729_, new_n728_, new_n214_ );
and g624 ( new_n730_, new_n428_, new_n729_ );
and g625 ( new_n731_, new_n720_, new_n730_ );
not g626 ( new_n732_, new_n731_ );
and g627 ( new_n733_, new_n732_, N5 );
and g628 ( new_n734_, new_n731_, new_n301_ );
or g629 ( N725, new_n733_, new_n734_ );
and g630 ( new_n736_, new_n424_, new_n425_ );
and g631 ( new_n737_, new_n401_, new_n420_ );
or g632 ( new_n738_, new_n736_, new_n737_ );
and g633 ( new_n739_, new_n376_, new_n738_ );
and g634 ( new_n740_, new_n739_, new_n324_ );
and g635 ( new_n741_, new_n740_, new_n214_ );
and g636 ( new_n742_, new_n741_, new_n720_ );
not g637 ( new_n743_, new_n742_ );
and g638 ( new_n744_, new_n743_, N9 );
and g639 ( new_n745_, new_n742_, new_n405_ );
or g640 ( N726, new_n744_, new_n745_ );
and g641 ( new_n747_, new_n374_, new_n369_ );
and g642 ( new_n748_, new_n350_, new_n370_ );
or g643 ( new_n749_, new_n747_, new_n748_ );
and g644 ( new_n750_, new_n749_, new_n427_ );
and g645 ( new_n751_, new_n324_, new_n214_ );
and g646 ( new_n752_, new_n750_, new_n751_ );
and g647 ( new_n753_, new_n720_, new_n752_ );
not g648 ( new_n754_, new_n753_ );
and g649 ( new_n755_, new_n754_, N13 );
and g650 ( new_n756_, new_n753_, new_n353_ );
or g651 ( N727, new_n755_, new_n756_ );
and g652 ( new_n758_, new_n715_, new_n716_ );
and g653 ( new_n759_, new_n696_, new_n711_ );
or g654 ( new_n760_, new_n758_, new_n759_ );
or g655 ( new_n761_, new_n668_, new_n669_ );
or g656 ( new_n762_, new_n649_, new_n664_ );
and g657 ( new_n763_, new_n762_, new_n761_ );
and g658 ( new_n764_, new_n624_, new_n763_ );
and g659 ( new_n765_, new_n764_, new_n760_ );
and g660 ( new_n766_, new_n765_, new_n429_ );
not g661 ( new_n767_, new_n766_ );
and g662 ( new_n768_, new_n767_, N17 );
and g663 ( new_n769_, new_n766_, new_n190_ );
or g664 ( N728, new_n768_, new_n769_ );
and g665 ( new_n771_, new_n765_, new_n730_ );
not g666 ( new_n772_, new_n771_ );
and g667 ( new_n773_, new_n772_, N21 );
and g668 ( new_n774_, new_n771_, new_n299_ );
or g669 ( N729, new_n773_, new_n774_ );
and g670 ( new_n776_, new_n741_, new_n765_ );
not g671 ( new_n777_, new_n776_ );
and g672 ( new_n778_, new_n777_, N25 );
and g673 ( new_n779_, new_n776_, new_n403_ );
or g674 ( N730, new_n778_, new_n779_ );
and g675 ( new_n781_, new_n765_, new_n752_ );
not g676 ( new_n782_, new_n781_ );
and g677 ( new_n783_, new_n782_, N29 );
and g678 ( new_n784_, new_n781_, new_n351_ );
or g679 ( N731, new_n783_, new_n784_ );
or g680 ( new_n786_, new_n620_, new_n621_ );
or g681 ( new_n787_, new_n601_, new_n616_ );
and g682 ( new_n788_, new_n787_, new_n786_ );
or g683 ( new_n789_, new_n523_, new_n524_ );
or g684 ( new_n790_, new_n504_, new_n519_ );
and g685 ( new_n791_, new_n790_, new_n789_ );
and g686 ( new_n792_, new_n719_, new_n791_ );
and g687 ( new_n793_, new_n792_, new_n788_ );
and g688 ( new_n794_, new_n793_, new_n429_ );
or g689 ( new_n795_, new_n794_, N33 );
and g690 ( new_n796_, new_n792_, N33 );
and g691 ( new_n797_, new_n429_, new_n788_ );
and g692 ( new_n798_, new_n797_, new_n796_ );
not g693 ( new_n799_, new_n798_ );
and g694 ( N732, new_n795_, new_n799_ );
and g695 ( new_n801_, new_n730_, new_n788_ );
and g696 ( new_n802_, new_n801_, new_n792_ );
not g697 ( new_n803_, new_n802_ );
and g698 ( new_n804_, new_n803_, N37 );
and g699 ( new_n805_, new_n802_, new_n305_ );
or g700 ( N733, new_n804_, new_n805_ );
and g701 ( new_n807_, new_n741_, new_n793_ );
or g702 ( new_n808_, new_n807_, N41 );
and g703 ( new_n809_, new_n792_, N41 );
and g704 ( new_n810_, new_n741_, new_n788_ );
and g705 ( new_n811_, new_n810_, new_n809_ );
not g706 ( new_n812_, new_n811_ );
and g707 ( N734, new_n812_, new_n808_ );
and g708 ( new_n814_, new_n752_, new_n788_ );
and g709 ( new_n815_, new_n814_, new_n792_ );
not g710 ( new_n816_, new_n815_ );
and g711 ( new_n817_, new_n816_, N45 );
and g712 ( new_n818_, new_n815_, new_n357_ );
or g713 ( N735, new_n817_, new_n818_ );
and g714 ( new_n820_, new_n791_, new_n763_ );
and g715 ( new_n821_, new_n820_, new_n760_ );
and g716 ( new_n822_, new_n821_, new_n788_ );
and g717 ( new_n823_, new_n822_, new_n429_ );
not g718 ( new_n824_, new_n823_ );
and g719 ( new_n825_, new_n824_, N49 );
and g720 ( new_n826_, new_n823_, new_n197_ );
or g721 ( N736, new_n825_, new_n826_ );
and g722 ( new_n828_, new_n822_, new_n730_ );
not g723 ( new_n829_, new_n828_ );
and g724 ( new_n830_, new_n829_, N53 );
and g725 ( new_n831_, new_n828_, new_n306_ );
or g726 ( N737, new_n830_, new_n831_ );
and g727 ( new_n833_, new_n741_, new_n822_ );
not g728 ( new_n834_, new_n833_ );
and g729 ( new_n835_, new_n834_, N57 );
and g730 ( new_n836_, new_n833_, new_n410_ );
or g731 ( N738, new_n835_, new_n836_ );
and g732 ( new_n838_, new_n822_, new_n752_ );
not g733 ( new_n839_, new_n838_ );
and g734 ( new_n840_, new_n839_, N61 );
and g735 ( new_n841_, new_n838_, new_n358_ );
or g736 ( N739, new_n840_, new_n841_ );
and g737 ( new_n843_, new_n740_, new_n215_ );
and g738 ( new_n844_, new_n764_, new_n718_ );
and g739 ( new_n845_, new_n843_, new_n844_ );
not g740 ( new_n846_, new_n845_ );
and g741 ( new_n847_, new_n846_, N65 );
and g742 ( new_n848_, new_n845_, new_n140_ );
or g743 ( N740, new_n847_, new_n848_ );
and g744 ( new_n850_, new_n718_, new_n788_ );
and g745 ( new_n851_, new_n820_, new_n850_ );
and g746 ( new_n852_, new_n843_, new_n851_ );
not g747 ( new_n853_, new_n852_ );
and g748 ( new_n854_, new_n853_, N69 );
and g749 ( new_n855_, new_n852_, new_n141_ );
or g750 ( N741, new_n854_, new_n855_ );
and g751 ( new_n857_, new_n792_, new_n623_ );
and g752 ( new_n858_, new_n843_, new_n857_ );
not g753 ( new_n859_, new_n858_ );
and g754 ( new_n860_, new_n859_, N73 );
and g755 ( new_n861_, new_n858_, new_n136_ );
or g756 ( N742, new_n860_, new_n861_ );
and g757 ( new_n863_, new_n821_, new_n623_ );
and g758 ( new_n864_, new_n843_, new_n863_ );
not g759 ( new_n865_, new_n864_ );
and g760 ( new_n866_, new_n865_, N77 );
and g761 ( new_n867_, new_n864_, new_n134_ );
or g762 ( N743, new_n866_, new_n867_ );
and g763 ( new_n869_, new_n325_, new_n750_ );
and g764 ( new_n870_, new_n844_, new_n869_ );
not g765 ( new_n871_, new_n870_ );
and g766 ( new_n872_, new_n871_, N81 );
and g767 ( new_n873_, new_n870_, new_n108_ );
or g768 ( N744, new_n872_, new_n873_ );
and g769 ( new_n875_, new_n869_, new_n851_ );
not g770 ( new_n876_, new_n875_ );
and g771 ( new_n877_, new_n876_, N85 );
and g772 ( new_n878_, new_n875_, new_n110_ );
or g773 ( N745, new_n877_, new_n878_ );
and g774 ( new_n880_, new_n857_, new_n869_ );
not g775 ( new_n881_, new_n880_ );
and g776 ( new_n882_, new_n881_, N89 );
and g777 ( new_n883_, new_n880_, new_n115_ );
or g778 ( N746, new_n882_, new_n883_ );
and g779 ( new_n885_, new_n863_, new_n869_ );
not g780 ( new_n886_, new_n885_ );
and g781 ( new_n887_, new_n886_, N93 );
and g782 ( new_n888_, new_n885_, new_n113_ );
or g783 ( N747, new_n887_, new_n888_ );
and g784 ( new_n890_, new_n739_, new_n729_ );
and g785 ( new_n891_, new_n844_, new_n890_ );
not g786 ( new_n892_, new_n891_ );
and g787 ( new_n893_, new_n892_, N97 );
and g788 ( new_n894_, new_n891_, new_n246_ );
or g789 ( N748, new_n893_, new_n894_ );
and g790 ( new_n896_, new_n851_, new_n890_ );
not g791 ( new_n897_, new_n896_ );
and g792 ( new_n898_, new_n897_, N101 );
and g793 ( new_n899_, new_n896_, new_n244_ );
or g794 ( N749, new_n898_, new_n899_ );
and g795 ( new_n901_, new_n857_, new_n890_ );
not g796 ( new_n902_, new_n901_ );
and g797 ( new_n903_, new_n902_, N105 );
and g798 ( new_n904_, new_n901_, new_n251_ );
or g799 ( N750, new_n903_, new_n904_ );
and g800 ( new_n906_, new_n863_, new_n890_ );
not g801 ( new_n907_, new_n906_ );
and g802 ( new_n908_, new_n907_, N109 );
and g803 ( new_n909_, new_n906_, new_n249_ );
or g804 ( N751, new_n908_, new_n909_ );
and g805 ( new_n911_, new_n750_, new_n729_ );
and g806 ( new_n912_, new_n844_, new_n911_ );
not g807 ( new_n913_, new_n912_ );
and g808 ( new_n914_, new_n913_, N113 );
and g809 ( new_n915_, new_n912_, new_n220_ );
or g810 ( N752, new_n914_, new_n915_ );
and g811 ( new_n917_, new_n851_, new_n911_ );
not g812 ( new_n918_, new_n917_ );
and g813 ( new_n919_, new_n918_, N117 );
and g814 ( new_n920_, new_n917_, new_n218_ );
or g815 ( N753, new_n919_, new_n920_ );
and g816 ( new_n922_, new_n857_, new_n911_ );
not g817 ( new_n923_, new_n922_ );
and g818 ( new_n924_, new_n923_, N121 );
and g819 ( new_n925_, new_n922_, new_n225_ );
or g820 ( N754, new_n924_, new_n925_ );
and g821 ( new_n927_, new_n863_, new_n911_ );
not g822 ( new_n928_, new_n927_ );
and g823 ( new_n929_, new_n928_, N125 );
and g824 ( new_n930_, new_n927_, new_n223_ );
or g825 ( N755, new_n929_, new_n930_ );
endmodule