module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n214_, new_n451_, new_n489_, new_n424_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n123_, new_n127_, new_n462_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n530_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n314_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n457_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n460_, new_n130_, new_n505_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n485_, new_n525_, new_n177_, new_n493_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n520_, new_n125_, new_n253_, new_n403_, new_n475_, new_n237_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n182_, new_n407_, new_n480_, new_n151_, new_n513_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n522_, new_n428_, new_n199_, new_n487_, new_n360_, new_n302_, new_n191_, new_n225_, new_n387_, new_n476_, new_n415_, new_n221_, new_n243_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n502_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n515_, new_n332_, new_n453_, new_n519_, new_n148_, new_n440_, new_n122_, new_n531_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n408_, new_n134_, new_n433_, new_n435_, new_n265_, new_n370_, new_n278_, new_n304_, new_n523_, new_n217_, new_n269_, new_n512_, new_n129_, new_n412_, new_n327_, new_n495_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n455_, new_n120_, new_n521_, new_n406_, new_n356_, new_n229_, new_n464_, new_n204_, new_n181_, new_n135_, new_n405_;

not g000 ( new_n119_, N75 );
nand g001 ( new_n120_, N29, N42 );
nor g002 ( N388, new_n120_, new_n119_ );
not g003 ( new_n122_, N80 );
nand g004 ( new_n123_, N29, N36 );
nor g005 ( N389, new_n123_, new_n122_ );
not g006 ( new_n125_, N42 );
nor g007 ( N390, new_n123_, new_n125_ );
nand g008 ( new_n127_, N85, N86 );
not g009 ( N391, new_n127_ );
not g010 ( new_n129_, N17 );
nand g011 ( new_n130_, N1, N8 );
not g012 ( new_n131_, new_n130_ );
nand g013 ( new_n132_, new_n131_, N13 );
nor g014 ( N418, new_n132_, new_n129_ );
xnor g015 ( new_n134_, N390, keyIn_0_0 );
not g016 ( new_n135_, new_n134_ );
nand g017 ( new_n136_, N1, N26 );
nand g018 ( new_n137_, N13, N17 );
nor g019 ( new_n138_, new_n136_, new_n137_ );
nand g020 ( N419, new_n135_, new_n138_ );
nand g021 ( new_n140_, N59, N75 );
not g022 ( new_n141_, new_n140_ );
nand g023 ( N420, new_n141_, N80 );
nand g024 ( new_n143_, N36, N59 );
not g025 ( new_n144_, new_n143_ );
nand g026 ( N421, new_n144_, N80 );
nand g027 ( N422, new_n144_, N42 );
not g028 ( new_n147_, N90 );
nor g029 ( new_n148_, N87, N88 );
nor g030 ( N423, new_n148_, new_n147_ );
nand g031 ( N446, new_n134_, new_n138_ );
not g032 ( new_n151_, N51 );
nor g033 ( N447, new_n136_, new_n151_ );
not g034 ( new_n153_, new_n132_ );
nand g035 ( new_n154_, new_n153_, N55 );
nand g036 ( new_n155_, N29, N68 );
xnor g037 ( new_n156_, new_n155_, keyIn_0_1 );
nor g038 ( N448, new_n154_, new_n156_ );
nand g039 ( new_n158_, N59, N68 );
not g040 ( new_n159_, new_n158_ );
nand g041 ( new_n160_, new_n159_, N74 );
nor g042 ( N449, new_n154_, new_n160_ );
not g043 ( new_n162_, N89 );
nor g044 ( N450, new_n148_, new_n162_ );
not g045 ( new_n164_, keyIn_0_7 );
nand g046 ( new_n165_, N101, N106 );
xnor g047 ( new_n166_, new_n165_, keyIn_0_2 );
nor g048 ( new_n167_, N101, N106 );
nor g049 ( new_n168_, new_n166_, new_n167_ );
xnor g050 ( new_n169_, N91, N96 );
not g051 ( new_n170_, new_n169_ );
nand g052 ( new_n171_, new_n168_, new_n170_ );
nor g053 ( new_n172_, new_n171_, new_n164_ );
nand g054 ( new_n173_, new_n171_, new_n164_ );
not g055 ( new_n174_, new_n168_ );
nand g056 ( new_n175_, new_n174_, new_n169_ );
nand g057 ( new_n176_, new_n173_, new_n175_ );
nor g058 ( new_n177_, new_n176_, new_n172_ );
nor g059 ( new_n178_, new_n177_, N130 );
xor g060 ( new_n179_, new_n178_, keyIn_0_10 );
nand g061 ( new_n180_, new_n177_, N130 );
xnor g062 ( new_n181_, new_n180_, keyIn_0_9 );
nand g063 ( new_n182_, new_n179_, new_n181_ );
xnor g064 ( new_n183_, N111, N116 );
xnor g065 ( new_n184_, N121, N126 );
xnor g066 ( new_n185_, new_n183_, new_n184_ );
xnor g067 ( new_n186_, new_n185_, N135 );
xnor g068 ( N767, new_n182_, new_n186_ );
not g069 ( new_n188_, keyIn_0_12 );
not g070 ( new_n189_, N130 );
xnor g071 ( new_n190_, N159, N165 );
xnor g072 ( new_n191_, N171, N177 );
xnor g073 ( new_n192_, new_n190_, new_n191_ );
nand g074 ( new_n193_, new_n192_, new_n189_ );
nor g075 ( new_n194_, new_n193_, new_n188_ );
nand g076 ( new_n195_, new_n193_, new_n188_ );
nor g077 ( new_n196_, new_n192_, new_n189_ );
nor g078 ( new_n197_, new_n196_, keyIn_0_15 );
nand g079 ( new_n198_, new_n197_, new_n195_ );
nor g080 ( new_n199_, new_n198_, new_n194_ );
not g081 ( new_n200_, keyIn_0_5 );
xor g082 ( new_n201_, N195, N201 );
not g083 ( new_n202_, new_n201_ );
nand g084 ( new_n203_, new_n202_, keyIn_0_6 );
nand g085 ( new_n204_, new_n203_, new_n200_ );
xor g086 ( new_n205_, N183, N189 );
nand g087 ( new_n206_, new_n204_, new_n205_ );
not g088 ( new_n207_, new_n205_ );
nand g089 ( new_n208_, new_n207_, new_n200_ );
nand g090 ( new_n209_, new_n208_, keyIn_0_6 );
nand g091 ( new_n210_, new_n209_, new_n201_ );
nand g092 ( new_n211_, new_n206_, new_n210_ );
xnor g093 ( new_n212_, new_n211_, N207 );
xnor g094 ( N768, new_n212_, new_n199_ );
not g095 ( new_n214_, keyIn_0_11 );
nand g096 ( new_n215_, N17, N51 );
nor g097 ( new_n216_, new_n130_, new_n215_ );
nor g098 ( new_n217_, new_n216_, keyIn_0_4 );
not g099 ( new_n218_, new_n217_ );
nand g100 ( new_n219_, new_n216_, keyIn_0_4 );
nand g101 ( new_n220_, new_n141_, N42 );
nand g102 ( new_n221_, new_n219_, new_n220_ );
not g103 ( new_n222_, new_n221_ );
nand g104 ( new_n223_, new_n222_, new_n218_ );
not g105 ( new_n224_, N447 );
nor g106 ( new_n225_, N17, N42 );
not g107 ( new_n226_, new_n225_ );
nand g108 ( new_n227_, N17, N42 );
not g109 ( new_n228_, new_n227_ );
nand g110 ( new_n229_, N59, N156 );
nor g111 ( new_n230_, new_n228_, new_n229_ );
nand g112 ( new_n231_, new_n230_, new_n226_ );
nor g113 ( new_n232_, new_n231_, new_n224_ );
not g114 ( new_n233_, new_n232_ );
nand g115 ( new_n234_, new_n223_, new_n233_ );
nand g116 ( new_n235_, new_n234_, N126 );
nand g117 ( new_n236_, new_n235_, new_n214_ );
not g118 ( new_n237_, N126 );
nor g119 ( new_n238_, new_n221_, new_n217_ );
nor g120 ( new_n239_, new_n238_, new_n232_ );
nor g121 ( new_n240_, new_n239_, new_n237_ );
nand g122 ( new_n241_, new_n240_, keyIn_0_11 );
nand g123 ( new_n242_, new_n236_, new_n241_ );
not g124 ( new_n243_, N153 );
not g125 ( new_n244_, N1 );
nand g126 ( new_n245_, N447, new_n229_ );
nor g127 ( new_n246_, new_n245_, new_n129_ );
nor g128 ( new_n247_, new_n246_, new_n244_ );
nor g129 ( new_n248_, new_n247_, new_n243_ );
nand g130 ( new_n249_, N29, N75 );
nor g131 ( new_n250_, new_n249_, new_n122_ );
nand g132 ( new_n251_, N447, new_n250_ );
not g133 ( new_n252_, N55 );
nor g134 ( new_n253_, new_n252_, N268 );
not g135 ( new_n254_, new_n253_ );
nor g136 ( new_n255_, new_n251_, new_n254_ );
nor g137 ( new_n256_, new_n248_, new_n255_ );
nand g138 ( new_n257_, new_n242_, new_n256_ );
nand g139 ( new_n258_, new_n257_, N201 );
not g140 ( new_n259_, new_n258_ );
nor g141 ( new_n260_, new_n257_, N201 );
nor g142 ( new_n261_, new_n259_, new_n260_ );
nand g143 ( new_n262_, new_n261_, N261 );
not g144 ( new_n263_, N219 );
nor g145 ( new_n264_, new_n261_, N261 );
nor g146 ( new_n265_, new_n264_, new_n263_ );
nand g147 ( new_n266_, new_n265_, new_n262_ );
nand g148 ( new_n267_, new_n261_, N228 );
not g149 ( new_n268_, N237 );
nor g150 ( new_n269_, new_n258_, new_n268_ );
not g151 ( new_n270_, N73 );
nand g152 ( new_n271_, N42, N72 );
nor g153 ( new_n272_, new_n271_, new_n270_ );
nand g154 ( new_n273_, new_n272_, new_n159_ );
nor g155 ( new_n274_, new_n154_, new_n273_ );
nand g156 ( new_n275_, new_n274_, N201 );
nand g157 ( new_n276_, N121, N210 );
nand g158 ( new_n277_, new_n275_, new_n276_ );
nor g159 ( new_n278_, new_n269_, new_n277_ );
nand g160 ( new_n279_, new_n267_, new_n278_ );
nand g161 ( new_n280_, new_n257_, N246 );
nand g162 ( new_n281_, N255, N267 );
nand g163 ( new_n282_, new_n280_, new_n281_ );
xnor g164 ( new_n283_, new_n282_, keyIn_0_19 );
nor g165 ( new_n284_, new_n279_, new_n283_ );
nand g166 ( N850, new_n266_, new_n284_ );
not g167 ( new_n286_, N261 );
nor g168 ( new_n287_, new_n260_, new_n286_ );
nor g169 ( new_n288_, new_n287_, new_n259_ );
nand g170 ( new_n289_, new_n234_, N121 );
not g171 ( new_n290_, N149 );
nor g172 ( new_n291_, new_n247_, new_n290_ );
nor g173 ( new_n292_, new_n291_, new_n255_ );
nand g174 ( new_n293_, new_n289_, new_n292_ );
xnor g175 ( new_n294_, new_n293_, keyIn_0_14 );
nor g176 ( new_n295_, new_n294_, N195 );
nor g177 ( new_n296_, new_n288_, new_n295_ );
not g178 ( new_n297_, keyIn_0_13 );
nand g179 ( new_n298_, new_n234_, N116 );
not g180 ( new_n299_, N146 );
nor g181 ( new_n300_, new_n247_, new_n299_ );
nor g182 ( new_n301_, new_n300_, new_n255_ );
nand g183 ( new_n302_, new_n298_, new_n301_ );
xnor g184 ( new_n303_, new_n302_, new_n297_ );
nor g185 ( new_n304_, new_n303_, N189 );
not g186 ( new_n305_, new_n304_ );
nand g187 ( new_n306_, new_n296_, new_n305_ );
nand g188 ( new_n307_, new_n303_, N189 );
xnor g189 ( new_n308_, new_n307_, keyIn_0_22 );
nand g190 ( new_n309_, new_n294_, N195 );
nor g191 ( new_n310_, new_n304_, new_n309_ );
nor g192 ( new_n311_, new_n308_, new_n310_ );
nand g193 ( new_n312_, new_n306_, new_n311_ );
xnor g194 ( new_n313_, new_n312_, keyIn_0_24 );
not g195 ( new_n314_, new_n313_ );
nand g196 ( new_n315_, new_n234_, N111 );
not g197 ( new_n316_, N143 );
nor g198 ( new_n317_, new_n247_, new_n316_ );
nor g199 ( new_n318_, new_n317_, new_n255_ );
nand g200 ( new_n319_, new_n315_, new_n318_ );
nor g201 ( new_n320_, new_n319_, N183 );
xor g202 ( new_n321_, new_n320_, keyIn_0_17 );
nand g203 ( new_n322_, new_n319_, N183 );
nand g204 ( new_n323_, new_n321_, new_n322_ );
nand g205 ( new_n324_, new_n314_, new_n323_ );
nor g206 ( new_n325_, new_n314_, new_n323_ );
nor g207 ( new_n326_, new_n325_, new_n263_ );
nand g208 ( new_n327_, new_n326_, new_n324_ );
not g209 ( new_n328_, N228 );
nor g210 ( new_n329_, new_n323_, new_n328_ );
xnor g211 ( new_n330_, new_n322_, keyIn_0_18 );
nand g212 ( new_n331_, new_n330_, N237 );
not g213 ( new_n332_, N246 );
not g214 ( new_n333_, new_n319_ );
nor g215 ( new_n334_, new_n333_, new_n332_ );
nand g216 ( new_n335_, new_n274_, N183 );
nand g217 ( new_n336_, N106, N210 );
xor g218 ( new_n337_, new_n336_, keyIn_0_3 );
nand g219 ( new_n338_, new_n335_, new_n337_ );
nor g220 ( new_n339_, new_n334_, new_n338_ );
nand g221 ( new_n340_, new_n331_, new_n339_ );
nor g222 ( new_n341_, new_n329_, new_n340_ );
nand g223 ( N863, new_n327_, new_n341_ );
not g224 ( new_n343_, new_n309_ );
nor g225 ( new_n344_, new_n296_, new_n343_ );
nand g226 ( new_n345_, new_n305_, new_n307_ );
nor g227 ( new_n346_, new_n344_, new_n345_ );
nand g228 ( new_n347_, new_n344_, new_n345_ );
nand g229 ( new_n348_, new_n347_, N219 );
nor g230 ( new_n349_, new_n348_, new_n346_ );
not g231 ( new_n350_, new_n345_ );
nand g232 ( new_n351_, new_n350_, N228 );
nor g233 ( new_n352_, new_n307_, new_n268_ );
nand g234 ( new_n353_, new_n303_, N246 );
nand g235 ( new_n354_, new_n274_, N189 );
nand g236 ( new_n355_, N111, N210 );
nand g237 ( new_n356_, N255, N259 );
nand g238 ( new_n357_, new_n355_, new_n356_ );
not g239 ( new_n358_, new_n357_ );
nand g240 ( new_n359_, new_n354_, new_n358_ );
not g241 ( new_n360_, new_n359_ );
nand g242 ( new_n361_, new_n353_, new_n360_ );
nor g243 ( new_n362_, new_n352_, new_n361_ );
nand g244 ( new_n363_, new_n351_, new_n362_ );
nor g245 ( new_n364_, new_n349_, new_n363_ );
xor g246 ( N864, new_n364_, keyIn_0_27 );
not g247 ( new_n366_, new_n288_ );
nor g248 ( new_n367_, new_n343_, new_n295_ );
nand g249 ( new_n368_, new_n366_, new_n367_ );
xnor g250 ( new_n369_, new_n368_, keyIn_0_25 );
nor g251 ( new_n370_, new_n366_, new_n367_ );
nor g252 ( new_n371_, new_n370_, new_n263_ );
nand g253 ( new_n372_, new_n369_, new_n371_ );
not g254 ( new_n373_, new_n367_ );
nor g255 ( new_n374_, new_n373_, new_n328_ );
nand g256 ( new_n375_, new_n343_, N237 );
not g257 ( new_n376_, new_n294_ );
nor g258 ( new_n377_, new_n376_, new_n332_ );
nand g259 ( new_n378_, new_n274_, N195 );
nand g260 ( new_n379_, N116, N210 );
nand g261 ( new_n380_, N255, N260 );
nand g262 ( new_n381_, new_n379_, new_n380_ );
not g263 ( new_n382_, new_n381_ );
nand g264 ( new_n383_, new_n378_, new_n382_ );
nor g265 ( new_n384_, new_n377_, new_n383_ );
nand g266 ( new_n385_, new_n384_, new_n375_ );
nor g267 ( new_n386_, new_n374_, new_n385_ );
nand g268 ( new_n387_, new_n372_, new_n386_ );
xnor g269 ( N865, new_n387_, keyIn_0_28 );
not g270 ( new_n389_, new_n330_ );
nand g271 ( new_n390_, new_n313_, new_n321_ );
nand g272 ( new_n391_, new_n390_, new_n389_ );
nand g273 ( new_n392_, new_n234_, N106 );
nor g274 ( new_n393_, new_n245_, new_n252_ );
not g275 ( new_n394_, new_n393_ );
nor g276 ( new_n395_, new_n394_, new_n243_ );
nor g277 ( new_n396_, new_n129_, N268 );
not g278 ( new_n397_, new_n396_ );
nor g279 ( new_n398_, new_n251_, new_n397_ );
not g280 ( new_n399_, new_n398_ );
nand g281 ( new_n400_, N138, N152 );
nand g282 ( new_n401_, new_n399_, new_n400_ );
nor g283 ( new_n402_, new_n395_, new_n401_ );
nand g284 ( new_n403_, new_n392_, new_n402_ );
nor g285 ( new_n404_, new_n403_, N177 );
not g286 ( new_n405_, new_n404_ );
nand g287 ( new_n406_, new_n391_, new_n405_ );
nand g288 ( new_n407_, new_n403_, N177 );
nand g289 ( new_n408_, new_n406_, new_n407_ );
not g290 ( new_n409_, N171 );
nand g291 ( new_n410_, new_n234_, N101 );
nor g292 ( new_n411_, new_n394_, new_n290_ );
nand g293 ( new_n412_, N17, N138 );
nand g294 ( new_n413_, new_n399_, new_n412_ );
nor g295 ( new_n414_, new_n411_, new_n413_ );
nand g296 ( new_n415_, new_n410_, new_n414_ );
not g297 ( new_n416_, new_n415_ );
nand g298 ( new_n417_, new_n416_, new_n409_ );
nand g299 ( new_n418_, new_n408_, new_n417_ );
nor g300 ( new_n419_, new_n416_, new_n409_ );
not g301 ( new_n420_, new_n419_ );
nand g302 ( new_n421_, new_n418_, new_n420_ );
nand g303 ( new_n422_, new_n234_, N96 );
nor g304 ( new_n423_, new_n394_, new_n299_ );
nand g305 ( new_n424_, N51, N138 );
nand g306 ( new_n425_, new_n399_, new_n424_ );
nor g307 ( new_n426_, new_n423_, new_n425_ );
nand g308 ( new_n427_, new_n422_, new_n426_ );
nor g309 ( new_n428_, new_n427_, N165 );
not g310 ( new_n429_, new_n428_ );
nand g311 ( new_n430_, new_n421_, new_n429_ );
nand g312 ( new_n431_, new_n427_, N165 );
xor g313 ( new_n432_, new_n431_, keyIn_0_16 );
nand g314 ( new_n433_, new_n430_, new_n432_ );
not g315 ( new_n434_, N159 );
nand g316 ( new_n435_, new_n234_, N91 );
nor g317 ( new_n436_, new_n398_, keyIn_0_8 );
nand g318 ( new_n437_, N8, N138 );
not g319 ( new_n438_, new_n437_ );
nor g320 ( new_n439_, new_n436_, new_n438_ );
not g321 ( new_n440_, new_n439_ );
nand g322 ( new_n441_, new_n393_, N143 );
nand g323 ( new_n442_, new_n398_, keyIn_0_8 );
nand g324 ( new_n443_, new_n442_, new_n441_ );
nor g325 ( new_n444_, new_n440_, new_n443_ );
nand g326 ( new_n445_, new_n444_, new_n435_ );
not g327 ( new_n446_, new_n445_ );
nand g328 ( new_n447_, new_n446_, new_n434_ );
nand g329 ( new_n448_, new_n433_, new_n447_ );
nand g330 ( new_n449_, new_n445_, N159 );
nand g331 ( N866, new_n448_, new_n449_ );
not g332 ( new_n451_, new_n407_ );
nor g333 ( new_n452_, new_n451_, new_n404_ );
nand g334 ( new_n453_, new_n391_, new_n452_ );
nor g335 ( new_n454_, new_n391_, new_n452_ );
nor g336 ( new_n455_, new_n454_, new_n263_ );
nand g337 ( new_n456_, new_n455_, new_n453_ );
nand g338 ( new_n457_, new_n452_, N228 );
nand g339 ( new_n458_, new_n451_, N237 );
nand g340 ( new_n459_, new_n457_, new_n458_ );
nor g341 ( new_n460_, new_n459_, keyIn_0_23 );
nand g342 ( new_n461_, new_n459_, keyIn_0_23 );
not g343 ( new_n462_, new_n403_ );
nor g344 ( new_n463_, new_n462_, new_n332_ );
nand g345 ( new_n464_, new_n274_, N177 );
nand g346 ( new_n465_, N101, N210 );
nand g347 ( new_n466_, new_n464_, new_n465_ );
nor g348 ( new_n467_, new_n463_, new_n466_ );
nand g349 ( new_n468_, new_n461_, new_n467_ );
nor g350 ( new_n469_, new_n468_, new_n460_ );
nand g351 ( N874, new_n456_, new_n469_ );
xnor g352 ( new_n471_, new_n445_, new_n434_ );
nand g353 ( new_n472_, new_n433_, new_n471_ );
nor g354 ( new_n473_, new_n433_, new_n471_ );
nor g355 ( new_n474_, new_n473_, new_n263_ );
nand g356 ( new_n475_, new_n474_, new_n472_ );
nand g357 ( new_n476_, new_n471_, N228 );
nor g358 ( new_n477_, new_n476_, keyIn_0_20 );
nand g359 ( new_n478_, new_n476_, keyIn_0_20 );
nor g360 ( new_n479_, new_n449_, new_n268_ );
nand g361 ( new_n480_, new_n445_, N246 );
nand g362 ( new_n481_, new_n274_, N159 );
nand g363 ( new_n482_, N210, N268 );
nand g364 ( new_n483_, new_n481_, new_n482_ );
not g365 ( new_n484_, new_n483_ );
nand g366 ( new_n485_, new_n480_, new_n484_ );
nor g367 ( new_n486_, new_n479_, new_n485_ );
nand g368 ( new_n487_, new_n478_, new_n486_ );
nor g369 ( new_n488_, new_n487_, new_n477_ );
nand g370 ( new_n489_, new_n475_, new_n488_ );
xnor g371 ( N878, new_n489_, keyIn_0_31 );
not g372 ( new_n491_, keyIn_0_29 );
nand g373 ( new_n492_, new_n432_, new_n429_ );
not g374 ( new_n493_, new_n492_ );
nand g375 ( new_n494_, new_n421_, new_n493_ );
nor g376 ( new_n495_, new_n421_, new_n493_ );
nor g377 ( new_n496_, new_n495_, new_n263_ );
nand g378 ( new_n497_, new_n496_, new_n494_ );
not g379 ( new_n498_, new_n497_ );
nand g380 ( new_n499_, new_n498_, new_n491_ );
nand g381 ( new_n500_, new_n497_, keyIn_0_29 );
nor g382 ( new_n501_, new_n492_, new_n328_ );
nor g383 ( new_n502_, new_n501_, keyIn_0_21 );
nand g384 ( new_n503_, new_n501_, keyIn_0_21 );
nor g385 ( new_n504_, new_n432_, new_n268_ );
nand g386 ( new_n505_, new_n427_, N246 );
nand g387 ( new_n506_, new_n274_, N165 );
nand g388 ( new_n507_, N91, N210 );
nand g389 ( new_n508_, new_n506_, new_n507_ );
not g390 ( new_n509_, new_n508_ );
nand g391 ( new_n510_, new_n505_, new_n509_ );
nor g392 ( new_n511_, new_n504_, new_n510_ );
nand g393 ( new_n512_, new_n503_, new_n511_ );
nor g394 ( new_n513_, new_n512_, new_n502_ );
nand g395 ( new_n514_, new_n500_, new_n513_ );
not g396 ( new_n515_, new_n514_ );
nand g397 ( N879, new_n515_, new_n499_ );
not g398 ( new_n517_, keyIn_0_26 );
nand g399 ( new_n518_, new_n420_, new_n417_ );
xor g400 ( new_n519_, new_n408_, new_n518_ );
nand g401 ( new_n520_, new_n519_, new_n517_ );
nor g402 ( new_n521_, new_n519_, new_n517_ );
nor g403 ( new_n522_, new_n521_, new_n263_ );
nand g404 ( new_n523_, new_n522_, new_n520_ );
nor g405 ( new_n524_, new_n518_, new_n328_ );
nand g406 ( new_n525_, new_n419_, N237 );
nor g407 ( new_n526_, new_n416_, new_n332_ );
nand g408 ( new_n527_, new_n274_, N171 );
nand g409 ( new_n528_, N96, N210 );
nand g410 ( new_n529_, new_n527_, new_n528_ );
nor g411 ( new_n530_, new_n526_, new_n529_ );
nand g412 ( new_n531_, new_n530_, new_n525_ );
nor g413 ( new_n532_, new_n524_, new_n531_ );
nand g414 ( new_n533_, new_n523_, new_n532_ );
xnor g415 ( N880, new_n533_, keyIn_0_30 );
endmodule