module add_mul_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, 
        b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, 
        b_15_, operation, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975;

  AND3_X1 U3525 ( .A1(n3493), .A2(n3494), .A3(operation), .ZN(Result_9_) );
  OR2_X1 U3526 ( .A1(n3495), .A2(n3496), .ZN(n3494) );
  INV_X1 U3527 ( .A(n3497), .ZN(n3493) );
  AND2_X1 U3528 ( .A1(n3496), .A2(n3495), .ZN(n3497) );
  OR2_X1 U3529 ( .A1(n3498), .A2(n3499), .ZN(n3495) );
  AND2_X1 U3530 ( .A1(n3500), .A2(n3501), .ZN(n3499) );
  INV_X1 U3531 ( .A(n3502), .ZN(n3498) );
  OR2_X1 U3532 ( .A1(n3501), .A2(n3500), .ZN(n3502) );
  AND3_X1 U3533 ( .A1(n3503), .A2(n3504), .A3(operation), .ZN(Result_8_) );
  OR3_X1 U3534 ( .A1(n3505), .A2(n3506), .A3(n3507), .ZN(n3504) );
  AND2_X1 U3535 ( .A1(n3508), .A2(n3509), .ZN(n3506) );
  AND2_X1 U3536 ( .A1(n3510), .A2(n3511), .ZN(n3505) );
  OR2_X1 U3537 ( .A1(n3511), .A2(n3512), .ZN(n3503) );
  AND2_X1 U3538 ( .A1(operation), .A2(n3513), .ZN(Result_7_) );
  OR2_X1 U3539 ( .A1(n3514), .A2(n3515), .ZN(n3513) );
  INV_X1 U3540 ( .A(n3516), .ZN(n3515) );
  OR2_X1 U3541 ( .A1(n3517), .A2(n3518), .ZN(n3516) );
  AND2_X1 U3542 ( .A1(n3518), .A2(n3517), .ZN(n3514) );
  OR2_X1 U3543 ( .A1(n3519), .A2(n3520), .ZN(n3517) );
  AND2_X1 U3544 ( .A1(n3521), .A2(n3522), .ZN(n3520) );
  OR2_X1 U3545 ( .A1(n3523), .A2(n3524), .ZN(n3522) );
  AND3_X1 U3546 ( .A1(n3525), .A2(n3526), .A3(operation), .ZN(Result_6_) );
  OR2_X1 U3547 ( .A1(n3527), .A2(n3528), .ZN(n3526) );
  INV_X1 U3548 ( .A(n3529), .ZN(n3527) );
  OR3_X1 U3549 ( .A1(n3530), .A2(n3531), .A3(n3529), .ZN(n3525) );
  AND2_X1 U3550 ( .A1(n3532), .A2(n3533), .ZN(n3531) );
  AND2_X1 U3551 ( .A1(n3534), .A2(n3528), .ZN(n3530) );
  AND2_X1 U3552 ( .A1(operation), .A2(n3535), .ZN(Result_5_) );
  OR2_X1 U3553 ( .A1(n3536), .A2(n3537), .ZN(n3535) );
  INV_X1 U3554 ( .A(n3538), .ZN(n3537) );
  OR2_X1 U3555 ( .A1(n3539), .A2(n3540), .ZN(n3538) );
  AND2_X1 U3556 ( .A1(n3540), .A2(n3539), .ZN(n3536) );
  OR2_X1 U3557 ( .A1(n3541), .A2(n3542), .ZN(n3539) );
  AND2_X1 U3558 ( .A1(n3543), .A2(n3544), .ZN(n3542) );
  OR2_X1 U3559 ( .A1(n3545), .A2(n3546), .ZN(n3544) );
  AND3_X1 U3560 ( .A1(n3547), .A2(n3548), .A3(operation), .ZN(Result_4_) );
  OR2_X1 U3561 ( .A1(n3549), .A2(n3550), .ZN(n3548) );
  INV_X1 U3562 ( .A(n3551), .ZN(n3549) );
  OR3_X1 U3563 ( .A1(n3552), .A2(n3553), .A3(n3551), .ZN(n3547) );
  AND2_X1 U3564 ( .A1(n3554), .A2(n3555), .ZN(n3553) );
  AND2_X1 U3565 ( .A1(n3556), .A2(n3550), .ZN(n3552) );
  AND2_X1 U3566 ( .A1(operation), .A2(n3557), .ZN(Result_3_) );
  OR2_X1 U3567 ( .A1(n3558), .A2(n3559), .ZN(n3557) );
  INV_X1 U3568 ( .A(n3560), .ZN(n3559) );
  OR2_X1 U3569 ( .A1(n3561), .A2(n3562), .ZN(n3560) );
  AND2_X1 U3570 ( .A1(n3562), .A2(n3561), .ZN(n3558) );
  OR2_X1 U3571 ( .A1(n3563), .A2(n3564), .ZN(n3561) );
  AND2_X1 U3572 ( .A1(n3565), .A2(n3566), .ZN(n3564) );
  OR2_X1 U3573 ( .A1(n3567), .A2(n3568), .ZN(n3566) );
  OR2_X1 U3574 ( .A1(n3569), .A2(n3570), .ZN(Result_31_) );
  AND2_X1 U3575 ( .A1(n3571), .A2(operation), .ZN(n3570) );
  AND2_X1 U3576 ( .A1(n3572), .A2(n3573), .ZN(n3569) );
  OR2_X1 U3577 ( .A1(n3574), .A2(n3575), .ZN(n3572) );
  AND2_X1 U3578 ( .A1(b_15_), .A2(n3576), .ZN(n3574) );
  OR2_X1 U3579 ( .A1(n3577), .A2(n3578), .ZN(Result_30_) );
  AND2_X1 U3580 ( .A1(n3579), .A2(n3573), .ZN(n3578) );
  OR2_X1 U3581 ( .A1(n3580), .A2(n3581), .ZN(n3579) );
  AND2_X1 U3582 ( .A1(n3582), .A2(n3583), .ZN(n3581) );
  INV_X1 U3583 ( .A(n3584), .ZN(n3580) );
  OR2_X1 U3584 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  OR2_X1 U3585 ( .A1(n3585), .A2(n3586), .ZN(n3582) );
  AND2_X1 U3586 ( .A1(b_14_), .A2(n3587), .ZN(n3585) );
  INV_X1 U3587 ( .A(n3571), .ZN(n3583) );
  AND2_X1 U3588 ( .A1(operation), .A2(n3588), .ZN(n3577) );
  OR2_X1 U3589 ( .A1(n3589), .A2(n3590), .ZN(n3588) );
  AND2_X1 U3590 ( .A1(b_15_), .A2(n3591), .ZN(n3590) );
  OR2_X1 U3591 ( .A1(n3586), .A2(n3592), .ZN(n3591) );
  AND2_X1 U3592 ( .A1(a_14_), .A2(n3593), .ZN(n3586) );
  AND2_X1 U3593 ( .A1(b_14_), .A2(n3594), .ZN(n3589) );
  OR2_X1 U3594 ( .A1(n3575), .A2(n3595), .ZN(n3594) );
  AND2_X1 U3595 ( .A1(a_15_), .A2(n3596), .ZN(n3575) );
  AND3_X1 U3596 ( .A1(n3597), .A2(n3598), .A3(operation), .ZN(Result_2_) );
  OR2_X1 U3597 ( .A1(n3599), .A2(n3600), .ZN(n3598) );
  OR3_X1 U3598 ( .A1(n3601), .A2(n3602), .A3(n3603), .ZN(n3597) );
  AND2_X1 U3599 ( .A1(n3604), .A2(n3605), .ZN(n3602) );
  INV_X1 U3600 ( .A(n3600), .ZN(n3604) );
  AND2_X1 U3601 ( .A1(n3606), .A2(n3600), .ZN(n3601) );
  OR2_X1 U3602 ( .A1(n3607), .A2(n3608), .ZN(Result_29_) );
  AND2_X1 U3603 ( .A1(n3609), .A2(operation), .ZN(n3608) );
  OR2_X1 U3604 ( .A1(n3610), .A2(n3611), .ZN(n3609) );
  AND2_X1 U3605 ( .A1(n3612), .A2(n3613), .ZN(n3611) );
  OR2_X1 U3606 ( .A1(n3614), .A2(n3615), .ZN(n3612) );
  AND2_X1 U3607 ( .A1(n3616), .A2(n3617), .ZN(n3615) );
  AND2_X1 U3608 ( .A1(n3618), .A2(n3619), .ZN(n3614) );
  AND3_X1 U3609 ( .A1(n3620), .A2(n3621), .A3(n3622), .ZN(n3610) );
  OR2_X1 U3610 ( .A1(n3616), .A2(n3617), .ZN(n3621) );
  OR2_X1 U3611 ( .A1(n3618), .A2(n3619), .ZN(n3620) );
  AND2_X1 U3612 ( .A1(n3623), .A2(n3573), .ZN(n3607) );
  OR2_X1 U3613 ( .A1(n3624), .A2(n3625), .ZN(n3623) );
  AND2_X1 U3614 ( .A1(n3626), .A2(n3627), .ZN(n3625) );
  OR2_X1 U3615 ( .A1(n3628), .A2(n3629), .ZN(n3626) );
  AND2_X1 U3616 ( .A1(a_13_), .A2(n3630), .ZN(n3629) );
  AND2_X1 U3617 ( .A1(b_13_), .A2(n3631), .ZN(n3628) );
  AND2_X1 U3618 ( .A1(n3632), .A2(n3633), .ZN(n3624) );
  OR2_X1 U3619 ( .A1(n3634), .A2(n3635), .ZN(n3632) );
  OR2_X1 U3620 ( .A1(n3636), .A2(n3637), .ZN(Result_28_) );
  AND3_X1 U3621 ( .A1(n3638), .A2(n3639), .A3(operation), .ZN(n3637) );
  INV_X1 U3622 ( .A(n3640), .ZN(n3639) );
  AND2_X1 U3623 ( .A1(n3641), .A2(n3642), .ZN(n3640) );
  OR2_X1 U3624 ( .A1(n3642), .A2(n3641), .ZN(n3638) );
  AND2_X1 U3625 ( .A1(n3643), .A2(n3644), .ZN(n3641) );
  INV_X1 U3626 ( .A(n3645), .ZN(n3644) );
  AND2_X1 U3627 ( .A1(n3646), .A2(n3647), .ZN(n3645) );
  OR2_X1 U3628 ( .A1(n3647), .A2(n3646), .ZN(n3643) );
  AND2_X1 U3629 ( .A1(n3648), .A2(n3573), .ZN(n3636) );
  OR2_X1 U3630 ( .A1(n3649), .A2(n3650), .ZN(n3648) );
  AND2_X1 U3631 ( .A1(n3651), .A2(n3652), .ZN(n3650) );
  AND2_X1 U3632 ( .A1(n3653), .A2(n3654), .ZN(n3649) );
  OR2_X1 U3633 ( .A1(n3655), .A2(n3656), .ZN(n3654) );
  INV_X1 U3634 ( .A(n3657), .ZN(n3653) );
  OR2_X1 U3635 ( .A1(n3658), .A2(n3659), .ZN(Result_27_) );
  AND3_X1 U3636 ( .A1(n3660), .A2(n3661), .A3(operation), .ZN(n3659) );
  INV_X1 U3637 ( .A(n3662), .ZN(n3661) );
  AND2_X1 U3638 ( .A1(n3663), .A2(n3664), .ZN(n3662) );
  OR2_X1 U3639 ( .A1(n3664), .A2(n3663), .ZN(n3660) );
  AND2_X1 U3640 ( .A1(n3665), .A2(n3666), .ZN(n3663) );
  OR2_X1 U3641 ( .A1(n3667), .A2(n3668), .ZN(n3666) );
  INV_X1 U3642 ( .A(n3669), .ZN(n3668) );
  OR2_X1 U3643 ( .A1(n3669), .A2(n3670), .ZN(n3665) );
  AND2_X1 U3644 ( .A1(n3671), .A2(n3573), .ZN(n3658) );
  OR3_X1 U3645 ( .A1(n3672), .A2(n3673), .A3(n3674), .ZN(n3671) );
  AND2_X1 U3646 ( .A1(n3675), .A2(n3676), .ZN(n3674) );
  AND2_X1 U3647 ( .A1(n3677), .A2(n3678), .ZN(n3673) );
  OR2_X1 U3648 ( .A1(n3679), .A2(n3680), .ZN(n3677) );
  AND2_X1 U3649 ( .A1(n3675), .A2(n3681), .ZN(n3680) );
  INV_X1 U3650 ( .A(n3682), .ZN(n3675) );
  AND2_X1 U3651 ( .A1(a_11_), .A2(n3682), .ZN(n3679) );
  AND3_X1 U3652 ( .A1(n3682), .A2(n3681), .A3(b_11_), .ZN(n3672) );
  OR2_X1 U3653 ( .A1(n3683), .A2(n3684), .ZN(Result_26_) );
  AND3_X1 U3654 ( .A1(n3685), .A2(n3686), .A3(operation), .ZN(n3684) );
  INV_X1 U3655 ( .A(n3687), .ZN(n3686) );
  AND2_X1 U3656 ( .A1(n3688), .A2(n3689), .ZN(n3687) );
  OR2_X1 U3657 ( .A1(n3689), .A2(n3688), .ZN(n3685) );
  AND2_X1 U3658 ( .A1(n3690), .A2(n3691), .ZN(n3688) );
  INV_X1 U3659 ( .A(n3692), .ZN(n3691) );
  AND2_X1 U3660 ( .A1(n3693), .A2(n3694), .ZN(n3692) );
  OR2_X1 U3661 ( .A1(n3694), .A2(n3693), .ZN(n3690) );
  INV_X1 U3662 ( .A(n3695), .ZN(n3693) );
  AND2_X1 U3663 ( .A1(n3696), .A2(n3573), .ZN(n3683) );
  OR2_X1 U3664 ( .A1(n3697), .A2(n3698), .ZN(n3696) );
  AND2_X1 U3665 ( .A1(n3699), .A2(n3700), .ZN(n3698) );
  INV_X1 U3666 ( .A(n3701), .ZN(n3697) );
  OR2_X1 U3667 ( .A1(n3700), .A2(n3699), .ZN(n3701) );
  INV_X1 U3668 ( .A(n3702), .ZN(n3699) );
  OR2_X1 U3669 ( .A1(n3703), .A2(n3704), .ZN(n3702) );
  OR2_X1 U3670 ( .A1(n3705), .A2(n3706), .ZN(Result_25_) );
  AND3_X1 U3671 ( .A1(n3707), .A2(n3708), .A3(operation), .ZN(n3706) );
  INV_X1 U3672 ( .A(n3709), .ZN(n3708) );
  AND2_X1 U3673 ( .A1(n3710), .A2(n3711), .ZN(n3709) );
  OR2_X1 U3674 ( .A1(n3711), .A2(n3710), .ZN(n3707) );
  AND2_X1 U3675 ( .A1(n3712), .A2(n3713), .ZN(n3710) );
  INV_X1 U3676 ( .A(n3714), .ZN(n3713) );
  AND2_X1 U3677 ( .A1(n3715), .A2(n3716), .ZN(n3714) );
  OR2_X1 U3678 ( .A1(n3716), .A2(n3715), .ZN(n3712) );
  AND2_X1 U3679 ( .A1(n3717), .A2(n3573), .ZN(n3705) );
  OR3_X1 U3680 ( .A1(n3718), .A2(n3719), .A3(n3720), .ZN(n3717) );
  AND2_X1 U3681 ( .A1(n3721), .A2(n3722), .ZN(n3720) );
  AND2_X1 U3682 ( .A1(n3723), .A2(n3724), .ZN(n3719) );
  OR2_X1 U3683 ( .A1(n3725), .A2(n3726), .ZN(n3723) );
  AND2_X1 U3684 ( .A1(n3721), .A2(n3727), .ZN(n3726) );
  INV_X1 U3685 ( .A(n3728), .ZN(n3721) );
  AND2_X1 U3686 ( .A1(a_9_), .A2(n3728), .ZN(n3725) );
  AND3_X1 U3687 ( .A1(n3728), .A2(n3727), .A3(b_9_), .ZN(n3718) );
  OR2_X1 U3688 ( .A1(n3729), .A2(n3730), .ZN(Result_24_) );
  AND3_X1 U3689 ( .A1(n3731), .A2(n3732), .A3(operation), .ZN(n3730) );
  INV_X1 U3690 ( .A(n3733), .ZN(n3732) );
  AND2_X1 U3691 ( .A1(n3734), .A2(n3735), .ZN(n3733) );
  OR2_X1 U3692 ( .A1(n3735), .A2(n3734), .ZN(n3731) );
  AND2_X1 U3693 ( .A1(n3736), .A2(n3737), .ZN(n3734) );
  INV_X1 U3694 ( .A(n3738), .ZN(n3737) );
  AND2_X1 U3695 ( .A1(n3739), .A2(n3740), .ZN(n3738) );
  OR2_X1 U3696 ( .A1(n3740), .A2(n3739), .ZN(n3736) );
  AND2_X1 U3697 ( .A1(n3741), .A2(n3573), .ZN(n3729) );
  OR2_X1 U3698 ( .A1(n3742), .A2(n3743), .ZN(n3741) );
  AND2_X1 U3699 ( .A1(n3744), .A2(n3745), .ZN(n3743) );
  INV_X1 U3700 ( .A(n3746), .ZN(n3742) );
  OR2_X1 U3701 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  AND2_X1 U3702 ( .A1(n3747), .A2(n3748), .ZN(n3744) );
  OR2_X1 U3703 ( .A1(n3749), .A2(n3750), .ZN(Result_23_) );
  AND3_X1 U3704 ( .A1(n3751), .A2(n3752), .A3(operation), .ZN(n3750) );
  INV_X1 U3705 ( .A(n3753), .ZN(n3752) );
  AND2_X1 U3706 ( .A1(n3754), .A2(n3755), .ZN(n3753) );
  OR2_X1 U3707 ( .A1(n3755), .A2(n3754), .ZN(n3751) );
  AND2_X1 U3708 ( .A1(n3756), .A2(n3757), .ZN(n3754) );
  INV_X1 U3709 ( .A(n3758), .ZN(n3757) );
  AND2_X1 U3710 ( .A1(n3759), .A2(n3760), .ZN(n3758) );
  OR2_X1 U3711 ( .A1(n3760), .A2(n3759), .ZN(n3756) );
  AND2_X1 U3712 ( .A1(n3761), .A2(n3573), .ZN(n3749) );
  OR3_X1 U3713 ( .A1(n3762), .A2(n3763), .A3(n3764), .ZN(n3761) );
  AND2_X1 U3714 ( .A1(n3765), .A2(n3766), .ZN(n3764) );
  AND2_X1 U3715 ( .A1(n3767), .A2(n3768), .ZN(n3763) );
  OR2_X1 U3716 ( .A1(n3769), .A2(n3770), .ZN(n3767) );
  AND2_X1 U3717 ( .A1(n3765), .A2(n3771), .ZN(n3770) );
  AND2_X1 U3718 ( .A1(a_7_), .A2(n3772), .ZN(n3769) );
  AND3_X1 U3719 ( .A1(n3772), .A2(n3771), .A3(b_7_), .ZN(n3762) );
  OR2_X1 U3720 ( .A1(n3773), .A2(n3774), .ZN(Result_22_) );
  AND3_X1 U3721 ( .A1(n3775), .A2(n3776), .A3(operation), .ZN(n3774) );
  INV_X1 U3722 ( .A(n3777), .ZN(n3776) );
  AND2_X1 U3723 ( .A1(n3778), .A2(n3779), .ZN(n3777) );
  OR2_X1 U3724 ( .A1(n3779), .A2(n3778), .ZN(n3775) );
  AND2_X1 U3725 ( .A1(n3780), .A2(n3781), .ZN(n3778) );
  INV_X1 U3726 ( .A(n3782), .ZN(n3781) );
  AND2_X1 U3727 ( .A1(n3783), .A2(n3784), .ZN(n3782) );
  OR2_X1 U3728 ( .A1(n3784), .A2(n3783), .ZN(n3780) );
  AND2_X1 U3729 ( .A1(n3785), .A2(n3573), .ZN(n3773) );
  OR2_X1 U3730 ( .A1(n3786), .A2(n3787), .ZN(n3785) );
  AND2_X1 U3731 ( .A1(n3788), .A2(n3789), .ZN(n3787) );
  INV_X1 U3732 ( .A(n3790), .ZN(n3786) );
  OR2_X1 U3733 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  AND2_X1 U3734 ( .A1(n3791), .A2(n3792), .ZN(n3788) );
  OR2_X1 U3735 ( .A1(n3793), .A2(n3794), .ZN(Result_21_) );
  AND3_X1 U3736 ( .A1(n3795), .A2(n3796), .A3(operation), .ZN(n3794) );
  INV_X1 U3737 ( .A(n3797), .ZN(n3796) );
  AND2_X1 U3738 ( .A1(n3798), .A2(n3799), .ZN(n3797) );
  OR2_X1 U3739 ( .A1(n3799), .A2(n3798), .ZN(n3795) );
  AND2_X1 U3740 ( .A1(n3800), .A2(n3801), .ZN(n3798) );
  INV_X1 U3741 ( .A(n3802), .ZN(n3801) );
  AND2_X1 U3742 ( .A1(n3803), .A2(n3804), .ZN(n3802) );
  OR2_X1 U3743 ( .A1(n3804), .A2(n3803), .ZN(n3800) );
  AND2_X1 U3744 ( .A1(n3805), .A2(n3573), .ZN(n3793) );
  OR3_X1 U3745 ( .A1(n3806), .A2(n3807), .A3(n3808), .ZN(n3805) );
  AND2_X1 U3746 ( .A1(n3809), .A2(n3810), .ZN(n3808) );
  AND2_X1 U3747 ( .A1(n3811), .A2(n3812), .ZN(n3807) );
  OR2_X1 U3748 ( .A1(n3813), .A2(n3814), .ZN(n3811) );
  AND2_X1 U3749 ( .A1(n3809), .A2(n3815), .ZN(n3814) );
  AND2_X1 U3750 ( .A1(a_5_), .A2(n3816), .ZN(n3813) );
  AND3_X1 U3751 ( .A1(n3816), .A2(n3815), .A3(b_5_), .ZN(n3806) );
  OR2_X1 U3752 ( .A1(n3817), .A2(n3818), .ZN(Result_20_) );
  AND3_X1 U3753 ( .A1(n3819), .A2(n3820), .A3(operation), .ZN(n3818) );
  INV_X1 U3754 ( .A(n3821), .ZN(n3820) );
  AND2_X1 U3755 ( .A1(n3822), .A2(n3823), .ZN(n3821) );
  OR2_X1 U3756 ( .A1(n3823), .A2(n3822), .ZN(n3819) );
  AND2_X1 U3757 ( .A1(n3824), .A2(n3825), .ZN(n3822) );
  INV_X1 U3758 ( .A(n3826), .ZN(n3825) );
  AND2_X1 U3759 ( .A1(n3827), .A2(n3828), .ZN(n3826) );
  OR2_X1 U3760 ( .A1(n3828), .A2(n3827), .ZN(n3824) );
  AND2_X1 U3761 ( .A1(n3829), .A2(n3573), .ZN(n3817) );
  OR2_X1 U3762 ( .A1(n3830), .A2(n3831), .ZN(n3829) );
  AND2_X1 U3763 ( .A1(n3832), .A2(n3833), .ZN(n3831) );
  INV_X1 U3764 ( .A(n3834), .ZN(n3830) );
  OR2_X1 U3765 ( .A1(n3833), .A2(n3832), .ZN(n3834) );
  AND2_X1 U3766 ( .A1(n3835), .A2(n3836), .ZN(n3832) );
  AND2_X1 U3767 ( .A1(operation), .A2(n3837), .ZN(Result_1_) );
  OR2_X1 U3768 ( .A1(n3838), .A2(n3839), .ZN(n3837) );
  INV_X1 U3769 ( .A(n3840), .ZN(n3839) );
  OR2_X1 U3770 ( .A1(n3841), .A2(n3842), .ZN(n3840) );
  AND2_X1 U3771 ( .A1(n3842), .A2(n3841), .ZN(n3838) );
  OR2_X1 U3772 ( .A1(n3843), .A2(n3844), .ZN(n3841) );
  INV_X1 U3773 ( .A(n3845), .ZN(n3844) );
  OR2_X1 U3774 ( .A1(n3846), .A2(n3847), .ZN(n3845) );
  OR2_X1 U3775 ( .A1(n3848), .A2(n3849), .ZN(Result_19_) );
  AND3_X1 U3776 ( .A1(n3850), .A2(n3851), .A3(operation), .ZN(n3849) );
  INV_X1 U3777 ( .A(n3852), .ZN(n3851) );
  AND2_X1 U3778 ( .A1(n3853), .A2(n3854), .ZN(n3852) );
  OR2_X1 U3779 ( .A1(n3854), .A2(n3853), .ZN(n3850) );
  AND2_X1 U3780 ( .A1(n3855), .A2(n3856), .ZN(n3853) );
  INV_X1 U3781 ( .A(n3857), .ZN(n3856) );
  AND2_X1 U3782 ( .A1(n3858), .A2(n3859), .ZN(n3857) );
  OR2_X1 U3783 ( .A1(n3859), .A2(n3858), .ZN(n3855) );
  AND2_X1 U3784 ( .A1(n3860), .A2(n3573), .ZN(n3848) );
  OR3_X1 U3785 ( .A1(n3861), .A2(n3862), .A3(n3863), .ZN(n3860) );
  AND2_X1 U3786 ( .A1(n3864), .A2(n3865), .ZN(n3863) );
  AND2_X1 U3787 ( .A1(n3866), .A2(n3867), .ZN(n3862) );
  OR2_X1 U3788 ( .A1(n3868), .A2(n3869), .ZN(n3866) );
  AND2_X1 U3789 ( .A1(n3864), .A2(n3870), .ZN(n3869) );
  AND2_X1 U3790 ( .A1(a_3_), .A2(n3871), .ZN(n3868) );
  AND3_X1 U3791 ( .A1(n3871), .A2(n3870), .A3(b_3_), .ZN(n3861) );
  OR2_X1 U3792 ( .A1(n3872), .A2(n3873), .ZN(Result_18_) );
  AND3_X1 U3793 ( .A1(n3874), .A2(n3875), .A3(operation), .ZN(n3873) );
  INV_X1 U3794 ( .A(n3876), .ZN(n3875) );
  AND2_X1 U3795 ( .A1(n3877), .A2(n3878), .ZN(n3876) );
  OR2_X1 U3796 ( .A1(n3878), .A2(n3877), .ZN(n3874) );
  AND2_X1 U3797 ( .A1(n3879), .A2(n3880), .ZN(n3877) );
  INV_X1 U3798 ( .A(n3881), .ZN(n3880) );
  AND2_X1 U3799 ( .A1(n3882), .A2(n3883), .ZN(n3881) );
  OR2_X1 U3800 ( .A1(n3883), .A2(n3882), .ZN(n3879) );
  AND2_X1 U3801 ( .A1(n3884), .A2(n3573), .ZN(n3872) );
  OR2_X1 U3802 ( .A1(n3885), .A2(n3886), .ZN(n3884) );
  AND2_X1 U3803 ( .A1(n3887), .A2(n3888), .ZN(n3886) );
  INV_X1 U3804 ( .A(n3889), .ZN(n3885) );
  OR2_X1 U3805 ( .A1(n3888), .A2(n3887), .ZN(n3889) );
  AND2_X1 U3806 ( .A1(n3890), .A2(n3891), .ZN(n3887) );
  OR2_X1 U3807 ( .A1(n3892), .A2(n3893), .ZN(Result_17_) );
  AND3_X1 U3808 ( .A1(n3894), .A2(n3895), .A3(operation), .ZN(n3893) );
  INV_X1 U3809 ( .A(n3896), .ZN(n3895) );
  AND2_X1 U3810 ( .A1(n3897), .A2(n3898), .ZN(n3896) );
  OR2_X1 U3811 ( .A1(n3898), .A2(n3897), .ZN(n3894) );
  AND2_X1 U3812 ( .A1(n3899), .A2(n3900), .ZN(n3897) );
  INV_X1 U3813 ( .A(n3901), .ZN(n3900) );
  AND2_X1 U3814 ( .A1(n3902), .A2(n3903), .ZN(n3901) );
  OR2_X1 U3815 ( .A1(n3903), .A2(n3902), .ZN(n3899) );
  AND2_X1 U3816 ( .A1(n3904), .A2(n3573), .ZN(n3892) );
  OR3_X1 U3817 ( .A1(n3905), .A2(n3906), .A3(n3907), .ZN(n3904) );
  AND2_X1 U3818 ( .A1(n3908), .A2(n3909), .ZN(n3907) );
  AND2_X1 U3819 ( .A1(n3910), .A2(n3911), .ZN(n3906) );
  OR2_X1 U3820 ( .A1(n3912), .A2(n3913), .ZN(n3910) );
  AND2_X1 U3821 ( .A1(n3908), .A2(n3914), .ZN(n3913) );
  AND2_X1 U3822 ( .A1(a_1_), .A2(n3915), .ZN(n3912) );
  AND3_X1 U3823 ( .A1(n3915), .A2(n3914), .A3(b_1_), .ZN(n3905) );
  OR2_X1 U3824 ( .A1(n3916), .A2(n3917), .ZN(Result_16_) );
  AND3_X1 U3825 ( .A1(n3918), .A2(n3919), .A3(operation), .ZN(n3917) );
  INV_X1 U3826 ( .A(n3920), .ZN(n3919) );
  AND2_X1 U3827 ( .A1(n3921), .A2(n3922), .ZN(n3920) );
  OR2_X1 U3828 ( .A1(n3922), .A2(n3921), .ZN(n3918) );
  AND2_X1 U3829 ( .A1(n3923), .A2(n3924), .ZN(n3921) );
  OR2_X1 U3830 ( .A1(n3925), .A2(n3926), .ZN(n3924) );
  INV_X1 U3831 ( .A(n3927), .ZN(n3923) );
  AND2_X1 U3832 ( .A1(n3926), .A2(n3925), .ZN(n3927) );
  INV_X1 U3833 ( .A(n3928), .ZN(n3926) );
  AND2_X1 U3834 ( .A1(n3929), .A2(n3573), .ZN(n3916) );
  INV_X1 U3835 ( .A(operation), .ZN(n3573) );
  OR2_X1 U3836 ( .A1(n3930), .A2(n3931), .ZN(n3929) );
  AND2_X1 U3837 ( .A1(n3932), .A2(n3933), .ZN(n3931) );
  INV_X1 U3838 ( .A(n3934), .ZN(n3932) );
  AND2_X1 U3839 ( .A1(n3935), .A2(n3934), .ZN(n3930) );
  AND2_X1 U3840 ( .A1(n3936), .A2(n3937), .ZN(n3934) );
  OR2_X1 U3841 ( .A1(n3938), .A2(b_0_), .ZN(n3937) );
  OR2_X1 U3842 ( .A1(n3939), .A2(a_0_), .ZN(n3936) );
  INV_X1 U3843 ( .A(n3933), .ZN(n3935) );
  OR2_X1 U3844 ( .A1(n3940), .A2(n3941), .ZN(n3933) );
  AND2_X1 U3845 ( .A1(n3914), .A2(n3911), .ZN(n3941) );
  AND2_X1 U3846 ( .A1(n3915), .A2(n3942), .ZN(n3940) );
  INV_X1 U3847 ( .A(n3908), .ZN(n3915) );
  AND2_X1 U3848 ( .A1(n3943), .A2(n3890), .ZN(n3908) );
  OR2_X1 U3849 ( .A1(a_2_), .A2(b_2_), .ZN(n3890) );
  INV_X1 U3850 ( .A(n3944), .ZN(n3943) );
  AND2_X1 U3851 ( .A1(n3888), .A2(n3891), .ZN(n3944) );
  OR2_X1 U3852 ( .A1(n3945), .A2(n3946), .ZN(n3888) );
  AND2_X1 U3853 ( .A1(n3870), .A2(n3867), .ZN(n3946) );
  AND2_X1 U3854 ( .A1(n3871), .A2(n3947), .ZN(n3945) );
  INV_X1 U3855 ( .A(n3864), .ZN(n3871) );
  AND2_X1 U3856 ( .A1(n3948), .A2(n3835), .ZN(n3864) );
  OR2_X1 U3857 ( .A1(a_4_), .A2(b_4_), .ZN(n3835) );
  INV_X1 U3858 ( .A(n3949), .ZN(n3948) );
  AND2_X1 U3859 ( .A1(n3833), .A2(n3836), .ZN(n3949) );
  OR2_X1 U3860 ( .A1(n3950), .A2(n3951), .ZN(n3833) );
  AND2_X1 U3861 ( .A1(n3815), .A2(n3812), .ZN(n3951) );
  AND2_X1 U3862 ( .A1(n3816), .A2(n3952), .ZN(n3950) );
  INV_X1 U3863 ( .A(n3809), .ZN(n3816) );
  AND2_X1 U3864 ( .A1(n3953), .A2(n3791), .ZN(n3809) );
  OR2_X1 U3865 ( .A1(a_6_), .A2(b_6_), .ZN(n3791) );
  INV_X1 U3866 ( .A(n3954), .ZN(n3953) );
  AND2_X1 U3867 ( .A1(n3789), .A2(n3792), .ZN(n3954) );
  OR2_X1 U3868 ( .A1(n3955), .A2(n3956), .ZN(n3789) );
  AND2_X1 U3869 ( .A1(n3771), .A2(n3768), .ZN(n3956) );
  AND2_X1 U3870 ( .A1(n3772), .A2(n3957), .ZN(n3955) );
  INV_X1 U3871 ( .A(n3765), .ZN(n3772) );
  AND2_X1 U3872 ( .A1(n3958), .A2(n3747), .ZN(n3765) );
  OR2_X1 U3873 ( .A1(a_8_), .A2(b_8_), .ZN(n3747) );
  INV_X1 U3874 ( .A(n3959), .ZN(n3958) );
  AND2_X1 U3875 ( .A1(n3745), .A2(n3748), .ZN(n3959) );
  OR2_X1 U3876 ( .A1(n3960), .A2(n3961), .ZN(n3745) );
  AND2_X1 U3877 ( .A1(n3727), .A2(n3724), .ZN(n3961) );
  AND2_X1 U3878 ( .A1(n3728), .A2(n3962), .ZN(n3960) );
  OR2_X1 U3879 ( .A1(n3963), .A2(n3703), .ZN(n3728) );
  AND2_X1 U3880 ( .A1(n3964), .A2(n3965), .ZN(n3703) );
  AND2_X1 U3881 ( .A1(n3700), .A2(n3966), .ZN(n3963) );
  OR2_X1 U3882 ( .A1(n3967), .A2(n3968), .ZN(n3700) );
  AND2_X1 U3883 ( .A1(n3681), .A2(n3678), .ZN(n3968) );
  AND2_X1 U3884 ( .A1(n3969), .A2(n3682), .ZN(n3967) );
  OR2_X1 U3885 ( .A1(n3655), .A2(n3651), .ZN(n3682) );
  AND2_X1 U3886 ( .A1(n3657), .A2(n3970), .ZN(n3651) );
  OR2_X1 U3887 ( .A1(n3635), .A2(n3971), .ZN(n3657) );
  AND2_X1 U3888 ( .A1(n3627), .A2(n3972), .ZN(n3971) );
  INV_X1 U3889 ( .A(n3633), .ZN(n3627) );
  OR2_X1 U3890 ( .A1(n3973), .A2(n3974), .ZN(n3633) );
  AND2_X1 U3891 ( .A1(b_15_), .A2(n3975), .ZN(n3974) );
  AND2_X1 U3892 ( .A1(b_14_), .A2(n3976), .ZN(n3973) );
  OR2_X1 U3893 ( .A1(n3571), .A2(a_14_), .ZN(n3976) );
  AND2_X1 U3894 ( .A1(a_15_), .A2(b_15_), .ZN(n3571) );
  AND2_X1 U3895 ( .A1(n3631), .A2(n3630), .ZN(n3635) );
  INV_X1 U3896 ( .A(n3652), .ZN(n3655) );
  OR2_X1 U3897 ( .A1(a_12_), .A2(b_12_), .ZN(n3652) );
  AND3_X1 U3898 ( .A1(n3977), .A2(n3978), .A3(operation), .ZN(Result_15_) );
  OR2_X1 U3899 ( .A1(n3979), .A2(n3980), .ZN(n3978) );
  OR2_X1 U3900 ( .A1(n3981), .A2(n3982), .ZN(n3977) );
  AND3_X1 U3901 ( .A1(n3983), .A2(n3984), .A3(operation), .ZN(Result_14_) );
  OR2_X1 U3902 ( .A1(n3985), .A2(n3986), .ZN(n3983) );
  AND2_X1 U3903 ( .A1(n3987), .A2(n3988), .ZN(n3986) );
  INV_X1 U3904 ( .A(n3989), .ZN(n3987) );
  AND2_X1 U3905 ( .A1(n3981), .A2(n3982), .ZN(n3985) );
  INV_X1 U3906 ( .A(n3979), .ZN(n3981) );
  AND2_X1 U3907 ( .A1(operation), .A2(n3990), .ZN(Result_13_) );
  OR2_X1 U3908 ( .A1(n3991), .A2(n3992), .ZN(n3990) );
  INV_X1 U3909 ( .A(n3993), .ZN(n3992) );
  OR2_X1 U3910 ( .A1(n3994), .A2(n3995), .ZN(n3993) );
  AND2_X1 U3911 ( .A1(n3995), .A2(n3994), .ZN(n3991) );
  OR2_X1 U3912 ( .A1(n3996), .A2(n3997), .ZN(n3994) );
  AND2_X1 U3913 ( .A1(n3988), .A2(n3998), .ZN(n3996) );
  AND3_X1 U3914 ( .A1(n3999), .A2(n4000), .A3(operation), .ZN(Result_12_) );
  INV_X1 U3915 ( .A(n4001), .ZN(n4000) );
  AND2_X1 U3916 ( .A1(n4002), .A2(n4003), .ZN(n4001) );
  OR2_X1 U3917 ( .A1(n4002), .A2(n4003), .ZN(n3999) );
  AND2_X1 U3918 ( .A1(n4004), .A2(n4005), .ZN(n4003) );
  OR2_X1 U3919 ( .A1(n4006), .A2(n4007), .ZN(n4005) );
  INV_X1 U3920 ( .A(n4008), .ZN(n4007) );
  OR2_X1 U3921 ( .A1(n4008), .A2(n4009), .ZN(n4004) );
  AND3_X1 U3922 ( .A1(n4010), .A2(n4011), .A3(operation), .ZN(Result_11_) );
  INV_X1 U3923 ( .A(n4012), .ZN(n4011) );
  AND2_X1 U3924 ( .A1(n4013), .A2(n4014), .ZN(n4012) );
  OR2_X1 U3925 ( .A1(n4013), .A2(n4014), .ZN(n4010) );
  AND2_X1 U3926 ( .A1(n4015), .A2(n4016), .ZN(n4014) );
  OR2_X1 U3927 ( .A1(n4017), .A2(n4018), .ZN(n4016) );
  INV_X1 U3928 ( .A(n4019), .ZN(n4018) );
  OR2_X1 U3929 ( .A1(n4019), .A2(n4020), .ZN(n4015) );
  AND3_X1 U3930 ( .A1(n4021), .A2(n4022), .A3(operation), .ZN(Result_10_) );
  OR2_X1 U3931 ( .A1(n4023), .A2(n4024), .ZN(n4022) );
  INV_X1 U3932 ( .A(n4025), .ZN(n4021) );
  AND2_X1 U3933 ( .A1(n4023), .A2(n4024), .ZN(n4025) );
  OR2_X1 U3934 ( .A1(n4026), .A2(n4027), .ZN(n4024) );
  INV_X1 U3935 ( .A(n4028), .ZN(n4026) );
  OR2_X1 U3936 ( .A1(n4029), .A2(n4030), .ZN(n4028) );
  AND2_X1 U3937 ( .A1(operation), .A2(n4031), .ZN(Result_0_) );
  OR3_X1 U3938 ( .A1(n3843), .A2(n4032), .A3(n4033), .ZN(n4031) );
  AND2_X1 U3939 ( .A1(n4034), .A2(a_0_), .ZN(n4033) );
  AND2_X1 U3940 ( .A1(n3842), .A2(n3846), .ZN(n4032) );
  INV_X1 U3941 ( .A(n4035), .ZN(n3842) );
  OR2_X1 U3942 ( .A1(n4036), .A2(n3600), .ZN(n4035) );
  OR2_X1 U3943 ( .A1(n4037), .A2(n3847), .ZN(n3600) );
  AND2_X1 U3944 ( .A1(n4038), .A2(n4039), .ZN(n4037) );
  AND2_X1 U3945 ( .A1(n3599), .A2(n3605), .ZN(n4036) );
  INV_X1 U3946 ( .A(n3603), .ZN(n3599) );
  OR2_X1 U3947 ( .A1(n4040), .A2(n3563), .ZN(n3603) );
  AND3_X1 U3948 ( .A1(n4041), .A2(n4042), .A3(n4043), .ZN(n3563) );
  AND2_X1 U3949 ( .A1(n3562), .A2(n4043), .ZN(n4040) );
  INV_X1 U3950 ( .A(n3565), .ZN(n4043) );
  OR2_X1 U3951 ( .A1(n3606), .A2(n4044), .ZN(n3565) );
  AND3_X1 U3952 ( .A1(n4045), .A2(n4046), .A3(n4047), .ZN(n4044) );
  INV_X1 U3953 ( .A(n3605), .ZN(n3606) );
  OR2_X1 U3954 ( .A1(n4048), .A2(n4047), .ZN(n3605) );
  OR2_X1 U3955 ( .A1(n4049), .A2(n4050), .ZN(n4047) );
  AND2_X1 U3956 ( .A1(n4051), .A2(n4052), .ZN(n4050) );
  AND2_X1 U3957 ( .A1(n4053), .A2(n4054), .ZN(n4049) );
  OR2_X1 U3958 ( .A1(n4052), .A2(n4051), .ZN(n4054) );
  AND2_X1 U3959 ( .A1(n4045), .A2(n4046), .ZN(n4048) );
  OR2_X1 U3960 ( .A1(n4055), .A2(n4056), .ZN(n4046) );
  OR2_X1 U3961 ( .A1(n4057), .A2(n4058), .ZN(n4045) );
  INV_X1 U3962 ( .A(n4055), .ZN(n4058) );
  OR2_X1 U3963 ( .A1(n4059), .A2(n4060), .ZN(n4055) );
  AND2_X1 U3964 ( .A1(n4061), .A2(n4062), .ZN(n4060) );
  INV_X1 U3965 ( .A(n4063), .ZN(n4059) );
  OR2_X1 U3966 ( .A1(n4062), .A2(n4061), .ZN(n4063) );
  INV_X1 U3967 ( .A(n4064), .ZN(n4061) );
  INV_X1 U3968 ( .A(n4056), .ZN(n4057) );
  AND2_X1 U3969 ( .A1(n4065), .A2(n3554), .ZN(n3562) );
  INV_X1 U3970 ( .A(n3550), .ZN(n3554) );
  AND2_X1 U3971 ( .A1(n4066), .A2(n4067), .ZN(n3550) );
  OR2_X1 U3972 ( .A1(n3567), .A2(n4042), .ZN(n4067) );
  INV_X1 U3973 ( .A(n3568), .ZN(n4042) );
  INV_X1 U3974 ( .A(n4041), .ZN(n3567) );
  OR2_X1 U3975 ( .A1(n4041), .A2(n3568), .ZN(n4066) );
  OR2_X1 U3976 ( .A1(n4068), .A2(n4069), .ZN(n3568) );
  AND2_X1 U3977 ( .A1(n4070), .A2(n4071), .ZN(n4069) );
  AND2_X1 U3978 ( .A1(n4072), .A2(n4073), .ZN(n4068) );
  OR2_X1 U3979 ( .A1(n4071), .A2(n4070), .ZN(n4073) );
  OR2_X1 U3980 ( .A1(n4074), .A2(n4075), .ZN(n4041) );
  AND2_X1 U3981 ( .A1(n4076), .A2(n4053), .ZN(n4075) );
  INV_X1 U3982 ( .A(n4077), .ZN(n4074) );
  OR2_X1 U3983 ( .A1(n4053), .A2(n4076), .ZN(n4077) );
  OR2_X1 U3984 ( .A1(n4078), .A2(n4079), .ZN(n4076) );
  INV_X1 U3985 ( .A(n4080), .ZN(n4079) );
  OR2_X1 U3986 ( .A1(n4051), .A2(n4081), .ZN(n4080) );
  AND2_X1 U3987 ( .A1(n4081), .A2(n4051), .ZN(n4078) );
  OR2_X1 U3988 ( .A1(n3867), .A2(n3938), .ZN(n4051) );
  INV_X1 U3989 ( .A(n4052), .ZN(n4081) );
  OR2_X1 U3990 ( .A1(n4082), .A2(n4083), .ZN(n4052) );
  AND2_X1 U3991 ( .A1(n4084), .A2(n4085), .ZN(n4083) );
  AND2_X1 U3992 ( .A1(n4086), .A2(n4087), .ZN(n4082) );
  OR2_X1 U3993 ( .A1(n4085), .A2(n4084), .ZN(n4087) );
  INV_X1 U3994 ( .A(n4088), .ZN(n4084) );
  AND2_X1 U3995 ( .A1(n4089), .A2(n4090), .ZN(n4053) );
  INV_X1 U3996 ( .A(n4091), .ZN(n4090) );
  AND2_X1 U3997 ( .A1(n4092), .A2(n4093), .ZN(n4091) );
  OR2_X1 U3998 ( .A1(n4093), .A2(n4092), .ZN(n4089) );
  OR2_X1 U3999 ( .A1(n4094), .A2(n4095), .ZN(n4092) );
  AND2_X1 U4000 ( .A1(n4096), .A2(n4097), .ZN(n4095) );
  INV_X1 U4001 ( .A(n4098), .ZN(n4094) );
  OR2_X1 U4002 ( .A1(n4097), .A2(n4096), .ZN(n4098) );
  OR2_X1 U4003 ( .A1(n3551), .A2(n3556), .ZN(n4065) );
  OR2_X1 U4004 ( .A1(n4099), .A2(n3541), .ZN(n3551) );
  AND3_X1 U4005 ( .A1(n4100), .A2(n4101), .A3(n4102), .ZN(n3541) );
  AND2_X1 U4006 ( .A1(n3540), .A2(n4102), .ZN(n4099) );
  INV_X1 U4007 ( .A(n3543), .ZN(n4102) );
  OR2_X1 U4008 ( .A1(n3556), .A2(n4103), .ZN(n3543) );
  AND3_X1 U4009 ( .A1(n4104), .A2(n4105), .A3(n4106), .ZN(n4103) );
  INV_X1 U4010 ( .A(n3555), .ZN(n3556) );
  OR2_X1 U4011 ( .A1(n4107), .A2(n4106), .ZN(n3555) );
  OR2_X1 U4012 ( .A1(n4108), .A2(n4109), .ZN(n4106) );
  AND2_X1 U4013 ( .A1(n4110), .A2(n4111), .ZN(n4109) );
  AND2_X1 U4014 ( .A1(n4112), .A2(n4113), .ZN(n4108) );
  OR2_X1 U4015 ( .A1(n4111), .A2(n4110), .ZN(n4113) );
  AND2_X1 U4016 ( .A1(n4104), .A2(n4105), .ZN(n4107) );
  OR2_X1 U4017 ( .A1(n4114), .A2(n4072), .ZN(n4105) );
  INV_X1 U4018 ( .A(n4115), .ZN(n4072) );
  OR2_X1 U4019 ( .A1(n4115), .A2(n4116), .ZN(n4104) );
  INV_X1 U4020 ( .A(n4114), .ZN(n4116) );
  OR2_X1 U4021 ( .A1(n4117), .A2(n4118), .ZN(n4114) );
  AND2_X1 U4022 ( .A1(n4119), .A2(n4071), .ZN(n4118) );
  INV_X1 U4023 ( .A(n4120), .ZN(n4117) );
  OR2_X1 U4024 ( .A1(n4071), .A2(n4119), .ZN(n4120) );
  INV_X1 U4025 ( .A(n4070), .ZN(n4119) );
  OR2_X1 U4026 ( .A1(n4121), .A2(n3938), .ZN(n4070) );
  OR2_X1 U4027 ( .A1(n4122), .A2(n4123), .ZN(n4071) );
  AND2_X1 U4028 ( .A1(n4124), .A2(n4125), .ZN(n4123) );
  AND2_X1 U4029 ( .A1(n4126), .A2(n4127), .ZN(n4122) );
  OR2_X1 U4030 ( .A1(n4125), .A2(n4124), .ZN(n4127) );
  INV_X1 U4031 ( .A(n4128), .ZN(n4124) );
  OR2_X1 U4032 ( .A1(n4129), .A2(n4130), .ZN(n4115) );
  AND2_X1 U4033 ( .A1(n4131), .A2(n4086), .ZN(n4130) );
  INV_X1 U4034 ( .A(n4132), .ZN(n4129) );
  OR2_X1 U4035 ( .A1(n4086), .A2(n4131), .ZN(n4132) );
  OR2_X1 U4036 ( .A1(n4133), .A2(n4134), .ZN(n4131) );
  AND2_X1 U4037 ( .A1(n4088), .A2(n4085), .ZN(n4134) );
  INV_X1 U4038 ( .A(n4135), .ZN(n4133) );
  OR2_X1 U4039 ( .A1(n4085), .A2(n4088), .ZN(n4135) );
  AND2_X1 U4040 ( .A1(b_3_), .A2(a_1_), .ZN(n4088) );
  OR2_X1 U4041 ( .A1(n4136), .A2(n4137), .ZN(n4085) );
  AND2_X1 U4042 ( .A1(n4138), .A2(n4139), .ZN(n4137) );
  AND2_X1 U4043 ( .A1(n4140), .A2(n4141), .ZN(n4136) );
  OR2_X1 U4044 ( .A1(n4139), .A2(n4138), .ZN(n4141) );
  INV_X1 U4045 ( .A(n4142), .ZN(n4138) );
  AND2_X1 U4046 ( .A1(n4143), .A2(n4144), .ZN(n4086) );
  INV_X1 U4047 ( .A(n4145), .ZN(n4144) );
  AND2_X1 U4048 ( .A1(n4146), .A2(n4147), .ZN(n4145) );
  OR2_X1 U4049 ( .A1(n4147), .A2(n4146), .ZN(n4143) );
  OR2_X1 U4050 ( .A1(n4148), .A2(n4149), .ZN(n4146) );
  INV_X1 U4051 ( .A(n4150), .ZN(n4149) );
  OR2_X1 U4052 ( .A1(n3891), .A2(n4151), .ZN(n4150) );
  AND2_X1 U4053 ( .A1(n4151), .A2(n3891), .ZN(n4148) );
  INV_X1 U4054 ( .A(n4152), .ZN(n4151) );
  AND2_X1 U4055 ( .A1(n4153), .A2(n3532), .ZN(n3540) );
  INV_X1 U4056 ( .A(n3528), .ZN(n3532) );
  AND2_X1 U4057 ( .A1(n4154), .A2(n4155), .ZN(n3528) );
  OR2_X1 U4058 ( .A1(n3545), .A2(n4101), .ZN(n4155) );
  INV_X1 U4059 ( .A(n3546), .ZN(n4101) );
  INV_X1 U4060 ( .A(n4100), .ZN(n3545) );
  OR2_X1 U4061 ( .A1(n4100), .A2(n3546), .ZN(n4154) );
  OR2_X1 U4062 ( .A1(n4156), .A2(n4157), .ZN(n3546) );
  AND2_X1 U4063 ( .A1(n4158), .A2(n4159), .ZN(n4157) );
  AND2_X1 U4064 ( .A1(n4160), .A2(n4161), .ZN(n4156) );
  OR2_X1 U4065 ( .A1(n4159), .A2(n4158), .ZN(n4161) );
  OR2_X1 U4066 ( .A1(n4162), .A2(n4163), .ZN(n4100) );
  AND2_X1 U4067 ( .A1(n4164), .A2(n4112), .ZN(n4163) );
  INV_X1 U4068 ( .A(n4165), .ZN(n4162) );
  OR2_X1 U4069 ( .A1(n4112), .A2(n4164), .ZN(n4165) );
  OR2_X1 U4070 ( .A1(n4166), .A2(n4167), .ZN(n4164) );
  INV_X1 U4071 ( .A(n4168), .ZN(n4167) );
  OR2_X1 U4072 ( .A1(n4110), .A2(n4169), .ZN(n4168) );
  AND2_X1 U4073 ( .A1(n4169), .A2(n4110), .ZN(n4166) );
  OR2_X1 U4074 ( .A1(n3812), .A2(n3938), .ZN(n4110) );
  INV_X1 U4075 ( .A(n4111), .ZN(n4169) );
  OR2_X1 U4076 ( .A1(n4170), .A2(n4171), .ZN(n4111) );
  AND2_X1 U4077 ( .A1(n4172), .A2(n4173), .ZN(n4171) );
  AND2_X1 U4078 ( .A1(n4174), .A2(n4175), .ZN(n4170) );
  OR2_X1 U4079 ( .A1(n4173), .A2(n4172), .ZN(n4175) );
  INV_X1 U4080 ( .A(n4176), .ZN(n4172) );
  AND2_X1 U4081 ( .A1(n4177), .A2(n4178), .ZN(n4112) );
  INV_X1 U4082 ( .A(n4179), .ZN(n4178) );
  AND2_X1 U4083 ( .A1(n4180), .A2(n4126), .ZN(n4179) );
  OR2_X1 U4084 ( .A1(n4126), .A2(n4180), .ZN(n4177) );
  OR2_X1 U4085 ( .A1(n4181), .A2(n4182), .ZN(n4180) );
  AND2_X1 U4086 ( .A1(n4128), .A2(n4125), .ZN(n4182) );
  INV_X1 U4087 ( .A(n4183), .ZN(n4181) );
  OR2_X1 U4088 ( .A1(n4125), .A2(n4128), .ZN(n4183) );
  AND2_X1 U4089 ( .A1(b_4_), .A2(a_1_), .ZN(n4128) );
  OR2_X1 U4090 ( .A1(n4184), .A2(n4185), .ZN(n4125) );
  AND2_X1 U4091 ( .A1(n4186), .A2(n4187), .ZN(n4185) );
  AND2_X1 U4092 ( .A1(n4188), .A2(n4189), .ZN(n4184) );
  OR2_X1 U4093 ( .A1(n4187), .A2(n4186), .ZN(n4189) );
  INV_X1 U4094 ( .A(n4190), .ZN(n4186) );
  AND2_X1 U4095 ( .A1(n4191), .A2(n4192), .ZN(n4126) );
  INV_X1 U4096 ( .A(n4193), .ZN(n4192) );
  AND2_X1 U4097 ( .A1(n4194), .A2(n4140), .ZN(n4193) );
  OR2_X1 U4098 ( .A1(n4140), .A2(n4194), .ZN(n4191) );
  OR2_X1 U4099 ( .A1(n4195), .A2(n4196), .ZN(n4194) );
  AND2_X1 U4100 ( .A1(n4142), .A2(n4139), .ZN(n4196) );
  INV_X1 U4101 ( .A(n4197), .ZN(n4195) );
  OR2_X1 U4102 ( .A1(n4139), .A2(n4142), .ZN(n4197) );
  AND2_X1 U4103 ( .A1(b_3_), .A2(a_2_), .ZN(n4142) );
  OR2_X1 U4104 ( .A1(n4198), .A2(n4199), .ZN(n4139) );
  AND2_X1 U4105 ( .A1(n3947), .A2(n4200), .ZN(n4199) );
  AND2_X1 U4106 ( .A1(n4201), .A2(n4202), .ZN(n4198) );
  OR2_X1 U4107 ( .A1(n4200), .A2(n3947), .ZN(n4202) );
  INV_X1 U4108 ( .A(n3865), .ZN(n3947) );
  AND2_X1 U4109 ( .A1(n4203), .A2(n4204), .ZN(n4140) );
  INV_X1 U4110 ( .A(n4205), .ZN(n4204) );
  AND2_X1 U4111 ( .A1(n4206), .A2(n4207), .ZN(n4205) );
  OR2_X1 U4112 ( .A1(n4207), .A2(n4206), .ZN(n4203) );
  OR2_X1 U4113 ( .A1(n4208), .A2(n4209), .ZN(n4206) );
  AND2_X1 U4114 ( .A1(n4210), .A2(n4211), .ZN(n4209) );
  INV_X1 U4115 ( .A(n4212), .ZN(n4208) );
  OR2_X1 U4116 ( .A1(n4211), .A2(n4210), .ZN(n4212) );
  OR2_X1 U4117 ( .A1(n3529), .A2(n3534), .ZN(n4153) );
  OR2_X1 U4118 ( .A1(n4213), .A2(n3519), .ZN(n3529) );
  AND3_X1 U4119 ( .A1(n4214), .A2(n4215), .A3(n4216), .ZN(n3519) );
  AND2_X1 U4120 ( .A1(n3518), .A2(n4216), .ZN(n4213) );
  INV_X1 U4121 ( .A(n3521), .ZN(n4216) );
  OR2_X1 U4122 ( .A1(n3534), .A2(n4217), .ZN(n3521) );
  AND3_X1 U4123 ( .A1(n4218), .A2(n4219), .A3(n4220), .ZN(n4217) );
  INV_X1 U4124 ( .A(n3533), .ZN(n3534) );
  OR2_X1 U4125 ( .A1(n4221), .A2(n4220), .ZN(n3533) );
  OR2_X1 U4126 ( .A1(n4222), .A2(n4223), .ZN(n4220) );
  AND2_X1 U4127 ( .A1(n4224), .A2(n4225), .ZN(n4223) );
  AND2_X1 U4128 ( .A1(n4226), .A2(n4227), .ZN(n4222) );
  OR2_X1 U4129 ( .A1(n4225), .A2(n4224), .ZN(n4227) );
  AND2_X1 U4130 ( .A1(n4218), .A2(n4219), .ZN(n4221) );
  OR2_X1 U4131 ( .A1(n4228), .A2(n4160), .ZN(n4219) );
  INV_X1 U4132 ( .A(n4229), .ZN(n4160) );
  OR2_X1 U4133 ( .A1(n4229), .A2(n4230), .ZN(n4218) );
  INV_X1 U4134 ( .A(n4228), .ZN(n4230) );
  OR2_X1 U4135 ( .A1(n4231), .A2(n4232), .ZN(n4228) );
  AND2_X1 U4136 ( .A1(n4233), .A2(n4159), .ZN(n4232) );
  INV_X1 U4137 ( .A(n4234), .ZN(n4231) );
  OR2_X1 U4138 ( .A1(n4159), .A2(n4233), .ZN(n4234) );
  INV_X1 U4139 ( .A(n4158), .ZN(n4233) );
  OR2_X1 U4140 ( .A1(n4235), .A2(n3938), .ZN(n4158) );
  OR2_X1 U4141 ( .A1(n4236), .A2(n4237), .ZN(n4159) );
  AND2_X1 U4142 ( .A1(n4238), .A2(n4239), .ZN(n4237) );
  AND2_X1 U4143 ( .A1(n4240), .A2(n4241), .ZN(n4236) );
  OR2_X1 U4144 ( .A1(n4239), .A2(n4238), .ZN(n4241) );
  INV_X1 U4145 ( .A(n4242), .ZN(n4238) );
  OR2_X1 U4146 ( .A1(n4243), .A2(n4244), .ZN(n4229) );
  AND2_X1 U4147 ( .A1(n4245), .A2(n4174), .ZN(n4244) );
  INV_X1 U4148 ( .A(n4246), .ZN(n4243) );
  OR2_X1 U4149 ( .A1(n4174), .A2(n4245), .ZN(n4246) );
  OR2_X1 U4150 ( .A1(n4247), .A2(n4248), .ZN(n4245) );
  AND2_X1 U4151 ( .A1(n4176), .A2(n4173), .ZN(n4248) );
  INV_X1 U4152 ( .A(n4249), .ZN(n4247) );
  OR2_X1 U4153 ( .A1(n4173), .A2(n4176), .ZN(n4249) );
  AND2_X1 U4154 ( .A1(b_5_), .A2(a_1_), .ZN(n4176) );
  OR2_X1 U4155 ( .A1(n4250), .A2(n4251), .ZN(n4173) );
  AND2_X1 U4156 ( .A1(n4252), .A2(n4253), .ZN(n4251) );
  AND2_X1 U4157 ( .A1(n4254), .A2(n4255), .ZN(n4250) );
  OR2_X1 U4158 ( .A1(n4253), .A2(n4252), .ZN(n4255) );
  INV_X1 U4159 ( .A(n4256), .ZN(n4252) );
  AND2_X1 U4160 ( .A1(n4257), .A2(n4258), .ZN(n4174) );
  INV_X1 U4161 ( .A(n4259), .ZN(n4258) );
  AND2_X1 U4162 ( .A1(n4260), .A2(n4188), .ZN(n4259) );
  OR2_X1 U4163 ( .A1(n4188), .A2(n4260), .ZN(n4257) );
  OR2_X1 U4164 ( .A1(n4261), .A2(n4262), .ZN(n4260) );
  AND2_X1 U4165 ( .A1(n4190), .A2(n4187), .ZN(n4262) );
  INV_X1 U4166 ( .A(n4263), .ZN(n4261) );
  OR2_X1 U4167 ( .A1(n4187), .A2(n4190), .ZN(n4263) );
  AND2_X1 U4168 ( .A1(b_4_), .A2(a_2_), .ZN(n4190) );
  OR2_X1 U4169 ( .A1(n4264), .A2(n4265), .ZN(n4187) );
  AND2_X1 U4170 ( .A1(n4266), .A2(n4267), .ZN(n4265) );
  AND2_X1 U4171 ( .A1(n4268), .A2(n4269), .ZN(n4264) );
  OR2_X1 U4172 ( .A1(n4267), .A2(n4266), .ZN(n4269) );
  INV_X1 U4173 ( .A(n4270), .ZN(n4266) );
  AND2_X1 U4174 ( .A1(n4271), .A2(n4272), .ZN(n4188) );
  INV_X1 U4175 ( .A(n4273), .ZN(n4272) );
  AND2_X1 U4176 ( .A1(n4274), .A2(n4201), .ZN(n4273) );
  OR2_X1 U4177 ( .A1(n4201), .A2(n4274), .ZN(n4271) );
  OR2_X1 U4178 ( .A1(n4275), .A2(n4276), .ZN(n4274) );
  AND2_X1 U4179 ( .A1(n3865), .A2(n4200), .ZN(n4276) );
  INV_X1 U4180 ( .A(n4277), .ZN(n4275) );
  OR2_X1 U4181 ( .A1(n4200), .A2(n3865), .ZN(n4277) );
  AND2_X1 U4182 ( .A1(b_3_), .A2(a_3_), .ZN(n3865) );
  OR2_X1 U4183 ( .A1(n4278), .A2(n4279), .ZN(n4200) );
  AND2_X1 U4184 ( .A1(n4280), .A2(n4281), .ZN(n4279) );
  AND2_X1 U4185 ( .A1(n4282), .A2(n4283), .ZN(n4278) );
  OR2_X1 U4186 ( .A1(n4281), .A2(n4280), .ZN(n4283) );
  INV_X1 U4187 ( .A(n4284), .ZN(n4280) );
  AND2_X1 U4188 ( .A1(n4285), .A2(n4286), .ZN(n4201) );
  INV_X1 U4189 ( .A(n4287), .ZN(n4286) );
  AND2_X1 U4190 ( .A1(n4288), .A2(n4289), .ZN(n4287) );
  OR2_X1 U4191 ( .A1(n4289), .A2(n4288), .ZN(n4285) );
  OR2_X1 U4192 ( .A1(n4290), .A2(n4291), .ZN(n4288) );
  AND2_X1 U4193 ( .A1(n4292), .A2(n4293), .ZN(n4291) );
  INV_X1 U4194 ( .A(n4294), .ZN(n4290) );
  OR2_X1 U4195 ( .A1(n4293), .A2(n4292), .ZN(n4294) );
  AND2_X1 U4196 ( .A1(n4295), .A2(n3508), .ZN(n3518) );
  INV_X1 U4197 ( .A(n3511), .ZN(n3508) );
  AND2_X1 U4198 ( .A1(n4296), .A2(n4297), .ZN(n3511) );
  OR2_X1 U4199 ( .A1(n3523), .A2(n4215), .ZN(n4297) );
  INV_X1 U4200 ( .A(n3524), .ZN(n4215) );
  INV_X1 U4201 ( .A(n4214), .ZN(n3523) );
  OR2_X1 U4202 ( .A1(n4214), .A2(n3524), .ZN(n4296) );
  OR2_X1 U4203 ( .A1(n4298), .A2(n4299), .ZN(n3524) );
  AND2_X1 U4204 ( .A1(n4300), .A2(n4301), .ZN(n4299) );
  AND2_X1 U4205 ( .A1(n4302), .A2(n4303), .ZN(n4298) );
  OR2_X1 U4206 ( .A1(n4301), .A2(n4300), .ZN(n4303) );
  OR2_X1 U4207 ( .A1(n4304), .A2(n4305), .ZN(n4214) );
  AND2_X1 U4208 ( .A1(n4306), .A2(n4226), .ZN(n4305) );
  INV_X1 U4209 ( .A(n4307), .ZN(n4304) );
  OR2_X1 U4210 ( .A1(n4226), .A2(n4306), .ZN(n4307) );
  OR2_X1 U4211 ( .A1(n4308), .A2(n4309), .ZN(n4306) );
  INV_X1 U4212 ( .A(n4310), .ZN(n4309) );
  OR2_X1 U4213 ( .A1(n4224), .A2(n4311), .ZN(n4310) );
  AND2_X1 U4214 ( .A1(n4311), .A2(n4224), .ZN(n4308) );
  OR2_X1 U4215 ( .A1(n3768), .A2(n3938), .ZN(n4224) );
  INV_X1 U4216 ( .A(n4225), .ZN(n4311) );
  OR2_X1 U4217 ( .A1(n4312), .A2(n4313), .ZN(n4225) );
  AND2_X1 U4218 ( .A1(n4314), .A2(n4315), .ZN(n4313) );
  AND2_X1 U4219 ( .A1(n4316), .A2(n4317), .ZN(n4312) );
  OR2_X1 U4220 ( .A1(n4315), .A2(n4314), .ZN(n4317) );
  INV_X1 U4221 ( .A(n4318), .ZN(n4314) );
  AND2_X1 U4222 ( .A1(n4319), .A2(n4320), .ZN(n4226) );
  INV_X1 U4223 ( .A(n4321), .ZN(n4320) );
  AND2_X1 U4224 ( .A1(n4322), .A2(n4240), .ZN(n4321) );
  OR2_X1 U4225 ( .A1(n4240), .A2(n4322), .ZN(n4319) );
  OR2_X1 U4226 ( .A1(n4323), .A2(n4324), .ZN(n4322) );
  AND2_X1 U4227 ( .A1(n4242), .A2(n4239), .ZN(n4324) );
  INV_X1 U4228 ( .A(n4325), .ZN(n4323) );
  OR2_X1 U4229 ( .A1(n4239), .A2(n4242), .ZN(n4325) );
  AND2_X1 U4230 ( .A1(b_6_), .A2(a_1_), .ZN(n4242) );
  OR2_X1 U4231 ( .A1(n4326), .A2(n4327), .ZN(n4239) );
  AND2_X1 U4232 ( .A1(n4328), .A2(n4329), .ZN(n4327) );
  AND2_X1 U4233 ( .A1(n4330), .A2(n4331), .ZN(n4326) );
  OR2_X1 U4234 ( .A1(n4329), .A2(n4328), .ZN(n4331) );
  INV_X1 U4235 ( .A(n4332), .ZN(n4328) );
  AND2_X1 U4236 ( .A1(n4333), .A2(n4334), .ZN(n4240) );
  INV_X1 U4237 ( .A(n4335), .ZN(n4334) );
  AND2_X1 U4238 ( .A1(n4336), .A2(n4254), .ZN(n4335) );
  OR2_X1 U4239 ( .A1(n4254), .A2(n4336), .ZN(n4333) );
  OR2_X1 U4240 ( .A1(n4337), .A2(n4338), .ZN(n4336) );
  AND2_X1 U4241 ( .A1(n4256), .A2(n4253), .ZN(n4338) );
  INV_X1 U4242 ( .A(n4339), .ZN(n4337) );
  OR2_X1 U4243 ( .A1(n4253), .A2(n4256), .ZN(n4339) );
  AND2_X1 U4244 ( .A1(b_5_), .A2(a_2_), .ZN(n4256) );
  OR2_X1 U4245 ( .A1(n4340), .A2(n4341), .ZN(n4253) );
  AND2_X1 U4246 ( .A1(n4342), .A2(n4343), .ZN(n4341) );
  AND2_X1 U4247 ( .A1(n4344), .A2(n4345), .ZN(n4340) );
  OR2_X1 U4248 ( .A1(n4343), .A2(n4342), .ZN(n4345) );
  INV_X1 U4249 ( .A(n4346), .ZN(n4342) );
  AND2_X1 U4250 ( .A1(n4347), .A2(n4348), .ZN(n4254) );
  INV_X1 U4251 ( .A(n4349), .ZN(n4348) );
  AND2_X1 U4252 ( .A1(n4350), .A2(n4268), .ZN(n4349) );
  OR2_X1 U4253 ( .A1(n4268), .A2(n4350), .ZN(n4347) );
  OR2_X1 U4254 ( .A1(n4351), .A2(n4352), .ZN(n4350) );
  AND2_X1 U4255 ( .A1(n4270), .A2(n4267), .ZN(n4352) );
  INV_X1 U4256 ( .A(n4353), .ZN(n4351) );
  OR2_X1 U4257 ( .A1(n4267), .A2(n4270), .ZN(n4353) );
  AND2_X1 U4258 ( .A1(b_4_), .A2(a_3_), .ZN(n4270) );
  OR2_X1 U4259 ( .A1(n4354), .A2(n4355), .ZN(n4267) );
  AND2_X1 U4260 ( .A1(n3836), .A2(n4356), .ZN(n4355) );
  AND2_X1 U4261 ( .A1(n4357), .A2(n4358), .ZN(n4354) );
  OR2_X1 U4262 ( .A1(n4356), .A2(n3836), .ZN(n4358) );
  AND2_X1 U4263 ( .A1(n4359), .A2(n4360), .ZN(n4268) );
  INV_X1 U4264 ( .A(n4361), .ZN(n4360) );
  AND2_X1 U4265 ( .A1(n4362), .A2(n4282), .ZN(n4361) );
  OR2_X1 U4266 ( .A1(n4282), .A2(n4362), .ZN(n4359) );
  OR2_X1 U4267 ( .A1(n4363), .A2(n4364), .ZN(n4362) );
  AND2_X1 U4268 ( .A1(n4284), .A2(n4281), .ZN(n4364) );
  INV_X1 U4269 ( .A(n4365), .ZN(n4363) );
  OR2_X1 U4270 ( .A1(n4281), .A2(n4284), .ZN(n4365) );
  AND2_X1 U4271 ( .A1(b_3_), .A2(a_4_), .ZN(n4284) );
  OR2_X1 U4272 ( .A1(n4366), .A2(n4367), .ZN(n4281) );
  AND2_X1 U4273 ( .A1(n4368), .A2(n4369), .ZN(n4367) );
  AND2_X1 U4274 ( .A1(n4370), .A2(n4371), .ZN(n4366) );
  OR2_X1 U4275 ( .A1(n4369), .A2(n4368), .ZN(n4371) );
  INV_X1 U4276 ( .A(n4372), .ZN(n4368) );
  AND2_X1 U4277 ( .A1(n4373), .A2(n4374), .ZN(n4282) );
  INV_X1 U4278 ( .A(n4375), .ZN(n4374) );
  AND2_X1 U4279 ( .A1(n4376), .A2(n4377), .ZN(n4375) );
  OR2_X1 U4280 ( .A1(n4377), .A2(n4376), .ZN(n4373) );
  OR2_X1 U4281 ( .A1(n4378), .A2(n4379), .ZN(n4376) );
  AND2_X1 U4282 ( .A1(n4380), .A2(n4381), .ZN(n4379) );
  INV_X1 U4283 ( .A(n4382), .ZN(n4378) );
  OR2_X1 U4284 ( .A1(n4381), .A2(n4380), .ZN(n4382) );
  OR2_X1 U4285 ( .A1(n3510), .A2(n3507), .ZN(n4295) );
  INV_X1 U4286 ( .A(n3512), .ZN(n3507) );
  OR2_X1 U4287 ( .A1(n4383), .A2(n3501), .ZN(n3512) );
  OR2_X1 U4288 ( .A1(n3510), .A2(n4384), .ZN(n3501) );
  AND3_X1 U4289 ( .A1(n4385), .A2(n4386), .A3(n4387), .ZN(n4384) );
  AND2_X1 U4290 ( .A1(n3500), .A2(n3496), .ZN(n4383) );
  INV_X1 U4291 ( .A(n4388), .ZN(n3500) );
  OR2_X1 U4292 ( .A1(n4027), .A2(n4389), .ZN(n4388) );
  AND2_X1 U4293 ( .A1(n4390), .A2(n4030), .ZN(n4389) );
  AND2_X1 U4294 ( .A1(n4030), .A2(n4029), .ZN(n4027) );
  OR2_X1 U4295 ( .A1(n4391), .A2(n4392), .ZN(n4029) );
  AND2_X1 U4296 ( .A1(n4013), .A2(n4020), .ZN(n4392) );
  AND2_X1 U4297 ( .A1(n4020), .A2(n4019), .ZN(n4391) );
  OR2_X1 U4298 ( .A1(n4393), .A2(n4394), .ZN(n4019) );
  AND2_X1 U4299 ( .A1(n4002), .A2(n4009), .ZN(n4394) );
  AND2_X1 U4300 ( .A1(n4009), .A2(n4008), .ZN(n4393) );
  OR2_X1 U4301 ( .A1(n3997), .A2(n4395), .ZN(n4008) );
  AND2_X1 U4302 ( .A1(n3995), .A2(n4396), .ZN(n4395) );
  INV_X1 U4303 ( .A(n3984), .ZN(n3995) );
  OR4_X1 U4304 ( .A1(n3979), .A2(n3980), .A3(n4397), .A4(n3989), .ZN(n3984) );
  AND2_X1 U4305 ( .A1(n4398), .A2(n4399), .ZN(n3989) );
  INV_X1 U4306 ( .A(n3982), .ZN(n3980) );
  AND2_X1 U4307 ( .A1(n4400), .A2(n4401), .ZN(n3982) );
  OR2_X1 U4308 ( .A1(n4402), .A2(n4403), .ZN(n4401) );
  INV_X1 U4309 ( .A(n4404), .ZN(n4400) );
  AND2_X1 U4310 ( .A1(n4403), .A2(n4402), .ZN(n4404) );
  AND2_X1 U4311 ( .A1(n4405), .A2(n4406), .ZN(n4402) );
  OR2_X1 U4312 ( .A1(n4407), .A2(n4408), .ZN(n4406) );
  INV_X1 U4313 ( .A(n4409), .ZN(n4405) );
  AND2_X1 U4314 ( .A1(n4408), .A2(n4407), .ZN(n4409) );
  INV_X1 U4315 ( .A(n4410), .ZN(n4408) );
  OR2_X1 U4316 ( .A1(n4411), .A2(n4412), .ZN(n3979) );
  AND2_X1 U4317 ( .A1(n3925), .A2(n3928), .ZN(n4412) );
  AND2_X1 U4318 ( .A1(n3922), .A2(n4413), .ZN(n4411) );
  OR2_X1 U4319 ( .A1(n3925), .A2(n3928), .ZN(n4413) );
  OR2_X1 U4320 ( .A1(n4414), .A2(n4415), .ZN(n3928) );
  AND2_X1 U4321 ( .A1(n4416), .A2(n3903), .ZN(n4415) );
  AND2_X1 U4322 ( .A1(n3898), .A2(n4417), .ZN(n4414) );
  OR2_X1 U4323 ( .A1(n4416), .A2(n3903), .ZN(n4417) );
  OR2_X1 U4324 ( .A1(n4418), .A2(n4419), .ZN(n3903) );
  AND2_X1 U4325 ( .A1(n4420), .A2(n3883), .ZN(n4419) );
  AND2_X1 U4326 ( .A1(n3878), .A2(n4421), .ZN(n4418) );
  OR2_X1 U4327 ( .A1(n4420), .A2(n3883), .ZN(n4421) );
  OR2_X1 U4328 ( .A1(n4422), .A2(n4423), .ZN(n3883) );
  AND2_X1 U4329 ( .A1(n4424), .A2(n3859), .ZN(n4423) );
  AND2_X1 U4330 ( .A1(n3854), .A2(n4425), .ZN(n4422) );
  OR2_X1 U4331 ( .A1(n4424), .A2(n3859), .ZN(n4425) );
  OR2_X1 U4332 ( .A1(n4426), .A2(n4427), .ZN(n3859) );
  AND2_X1 U4333 ( .A1(n4428), .A2(n3828), .ZN(n4427) );
  AND2_X1 U4334 ( .A1(n3823), .A2(n4429), .ZN(n4426) );
  OR2_X1 U4335 ( .A1(n4428), .A2(n3828), .ZN(n4429) );
  OR2_X1 U4336 ( .A1(n4430), .A2(n4431), .ZN(n3828) );
  AND2_X1 U4337 ( .A1(n4432), .A2(n3804), .ZN(n4431) );
  AND2_X1 U4338 ( .A1(n3799), .A2(n4433), .ZN(n4430) );
  OR2_X1 U4339 ( .A1(n4432), .A2(n3804), .ZN(n4433) );
  OR2_X1 U4340 ( .A1(n4434), .A2(n4435), .ZN(n3804) );
  AND2_X1 U4341 ( .A1(n4436), .A2(n3784), .ZN(n4435) );
  AND2_X1 U4342 ( .A1(n3779), .A2(n4437), .ZN(n4434) );
  OR2_X1 U4343 ( .A1(n4436), .A2(n3784), .ZN(n4437) );
  OR2_X1 U4344 ( .A1(n4438), .A2(n4439), .ZN(n3784) );
  AND2_X1 U4345 ( .A1(n4440), .A2(n3760), .ZN(n4439) );
  AND2_X1 U4346 ( .A1(n3755), .A2(n4441), .ZN(n4438) );
  OR2_X1 U4347 ( .A1(n4440), .A2(n3760), .ZN(n4441) );
  OR2_X1 U4348 ( .A1(n4442), .A2(n4443), .ZN(n3760) );
  AND2_X1 U4349 ( .A1(n4444), .A2(n3740), .ZN(n4443) );
  AND2_X1 U4350 ( .A1(n3735), .A2(n4445), .ZN(n4442) );
  OR2_X1 U4351 ( .A1(n4444), .A2(n3740), .ZN(n4445) );
  OR2_X1 U4352 ( .A1(n4446), .A2(n4447), .ZN(n3740) );
  AND2_X1 U4353 ( .A1(n4448), .A2(n3716), .ZN(n4447) );
  AND2_X1 U4354 ( .A1(n3711), .A2(n4449), .ZN(n4446) );
  OR2_X1 U4355 ( .A1(n4448), .A2(n3716), .ZN(n4449) );
  OR2_X1 U4356 ( .A1(n4450), .A2(n4451), .ZN(n3716) );
  AND2_X1 U4357 ( .A1(n3695), .A2(n3694), .ZN(n4451) );
  AND2_X1 U4358 ( .A1(n3689), .A2(n4452), .ZN(n4450) );
  OR2_X1 U4359 ( .A1(n3695), .A2(n3694), .ZN(n4452) );
  OR2_X1 U4360 ( .A1(n4453), .A2(n4454), .ZN(n3694) );
  AND2_X1 U4361 ( .A1(n3667), .A2(n3669), .ZN(n4454) );
  AND2_X1 U4362 ( .A1(n3664), .A2(n4455), .ZN(n4453) );
  OR2_X1 U4363 ( .A1(n3667), .A2(n3669), .ZN(n4455) );
  OR2_X1 U4364 ( .A1(n4456), .A2(n4457), .ZN(n3669) );
  AND2_X1 U4365 ( .A1(n4458), .A2(n3647), .ZN(n4457) );
  AND2_X1 U4366 ( .A1(n3642), .A2(n4459), .ZN(n4456) );
  OR2_X1 U4367 ( .A1(n4458), .A2(n3647), .ZN(n4459) );
  OR2_X1 U4368 ( .A1(n4460), .A2(n4461), .ZN(n3647) );
  AND2_X1 U4369 ( .A1(n3619), .A2(n3617), .ZN(n4461) );
  AND2_X1 U4370 ( .A1(n3613), .A2(n4462), .ZN(n4460) );
  OR2_X1 U4371 ( .A1(n3619), .A2(n3617), .ZN(n4462) );
  INV_X1 U4372 ( .A(n3618), .ZN(n3617) );
  AND3_X1 U4373 ( .A1(n3975), .A2(b_14_), .A3(b_15_), .ZN(n3618) );
  INV_X1 U4374 ( .A(n3616), .ZN(n3619) );
  AND2_X1 U4375 ( .A1(a_13_), .A2(b_15_), .ZN(n3616) );
  INV_X1 U4376 ( .A(n3622), .ZN(n3613) );
  OR2_X1 U4377 ( .A1(n4463), .A2(n4464), .ZN(n3622) );
  AND2_X1 U4378 ( .A1(b_14_), .A2(n4465), .ZN(n4464) );
  OR2_X1 U4379 ( .A1(n4466), .A2(n3592), .ZN(n4465) );
  AND2_X1 U4380 ( .A1(a_14_), .A2(n3630), .ZN(n4466) );
  AND2_X1 U4381 ( .A1(b_13_), .A2(n4467), .ZN(n4463) );
  OR2_X1 U4382 ( .A1(n4468), .A2(n3595), .ZN(n4467) );
  AND2_X1 U4383 ( .A1(a_15_), .A2(n3593), .ZN(n4468) );
  INV_X1 U4384 ( .A(n3646), .ZN(n4458) );
  AND2_X1 U4385 ( .A1(a_12_), .A2(b_15_), .ZN(n3646) );
  OR2_X1 U4386 ( .A1(n4469), .A2(n4470), .ZN(n3642) );
  AND2_X1 U4387 ( .A1(n4471), .A2(n4472), .ZN(n4470) );
  INV_X1 U4388 ( .A(n4473), .ZN(n4469) );
  OR2_X1 U4389 ( .A1(n4471), .A2(n4472), .ZN(n4473) );
  OR2_X1 U4390 ( .A1(n4474), .A2(n4475), .ZN(n4471) );
  AND2_X1 U4391 ( .A1(n4476), .A2(n4477), .ZN(n4475) );
  AND2_X1 U4392 ( .A1(n4478), .A2(n4479), .ZN(n4474) );
  INV_X1 U4393 ( .A(n3670), .ZN(n3667) );
  AND2_X1 U4394 ( .A1(a_11_), .A2(b_15_), .ZN(n3670) );
  OR2_X1 U4395 ( .A1(n4480), .A2(n4481), .ZN(n3664) );
  INV_X1 U4396 ( .A(n4482), .ZN(n4481) );
  OR2_X1 U4397 ( .A1(n4483), .A2(n4484), .ZN(n4482) );
  AND2_X1 U4398 ( .A1(n4484), .A2(n4483), .ZN(n4480) );
  AND2_X1 U4399 ( .A1(n4485), .A2(n4486), .ZN(n4483) );
  OR2_X1 U4400 ( .A1(n4487), .A2(n4488), .ZN(n4486) );
  INV_X1 U4401 ( .A(n4489), .ZN(n4488) );
  OR2_X1 U4402 ( .A1(n4489), .A2(n4490), .ZN(n4485) );
  OR2_X1 U4403 ( .A1(n3964), .A2(n3596), .ZN(n3695) );
  OR2_X1 U4404 ( .A1(n4491), .A2(n4492), .ZN(n3689) );
  INV_X1 U4405 ( .A(n4493), .ZN(n4492) );
  OR2_X1 U4406 ( .A1(n4494), .A2(n4495), .ZN(n4493) );
  AND2_X1 U4407 ( .A1(n4495), .A2(n4494), .ZN(n4491) );
  AND2_X1 U4408 ( .A1(n4496), .A2(n4497), .ZN(n4494) );
  INV_X1 U4409 ( .A(n4498), .ZN(n4497) );
  AND2_X1 U4410 ( .A1(n4499), .A2(n4500), .ZN(n4498) );
  OR2_X1 U4411 ( .A1(n4500), .A2(n4499), .ZN(n4496) );
  INV_X1 U4412 ( .A(n3715), .ZN(n4448) );
  AND2_X1 U4413 ( .A1(a_9_), .A2(b_15_), .ZN(n3715) );
  OR2_X1 U4414 ( .A1(n4501), .A2(n4502), .ZN(n3711) );
  INV_X1 U4415 ( .A(n4503), .ZN(n4502) );
  OR2_X1 U4416 ( .A1(n4504), .A2(n4505), .ZN(n4503) );
  AND2_X1 U4417 ( .A1(n4505), .A2(n4504), .ZN(n4501) );
  AND2_X1 U4418 ( .A1(n4506), .A2(n4507), .ZN(n4504) );
  INV_X1 U4419 ( .A(n4508), .ZN(n4507) );
  AND2_X1 U4420 ( .A1(n4509), .A2(n4510), .ZN(n4508) );
  OR2_X1 U4421 ( .A1(n4510), .A2(n4509), .ZN(n4506) );
  INV_X1 U4422 ( .A(n4511), .ZN(n4509) );
  INV_X1 U4423 ( .A(n3739), .ZN(n4444) );
  AND2_X1 U4424 ( .A1(a_8_), .A2(b_15_), .ZN(n3739) );
  OR2_X1 U4425 ( .A1(n4512), .A2(n4513), .ZN(n3735) );
  INV_X1 U4426 ( .A(n4514), .ZN(n4513) );
  OR2_X1 U4427 ( .A1(n4515), .A2(n4516), .ZN(n4514) );
  AND2_X1 U4428 ( .A1(n4516), .A2(n4515), .ZN(n4512) );
  AND2_X1 U4429 ( .A1(n4517), .A2(n4518), .ZN(n4515) );
  INV_X1 U4430 ( .A(n4519), .ZN(n4518) );
  AND2_X1 U4431 ( .A1(n4520), .A2(n4521), .ZN(n4519) );
  OR2_X1 U4432 ( .A1(n4521), .A2(n4520), .ZN(n4517) );
  INV_X1 U4433 ( .A(n3759), .ZN(n4440) );
  AND2_X1 U4434 ( .A1(a_7_), .A2(b_15_), .ZN(n3759) );
  OR2_X1 U4435 ( .A1(n4522), .A2(n4523), .ZN(n3755) );
  INV_X1 U4436 ( .A(n4524), .ZN(n4523) );
  OR2_X1 U4437 ( .A1(n4525), .A2(n4526), .ZN(n4524) );
  AND2_X1 U4438 ( .A1(n4526), .A2(n4525), .ZN(n4522) );
  AND2_X1 U4439 ( .A1(n4527), .A2(n4528), .ZN(n4525) );
  INV_X1 U4440 ( .A(n4529), .ZN(n4528) );
  AND2_X1 U4441 ( .A1(n4530), .A2(n4531), .ZN(n4529) );
  OR2_X1 U4442 ( .A1(n4531), .A2(n4530), .ZN(n4527) );
  INV_X1 U4443 ( .A(n3783), .ZN(n4436) );
  AND2_X1 U4444 ( .A1(a_6_), .A2(b_15_), .ZN(n3783) );
  OR2_X1 U4445 ( .A1(n4532), .A2(n4533), .ZN(n3779) );
  INV_X1 U4446 ( .A(n4534), .ZN(n4533) );
  OR2_X1 U4447 ( .A1(n4535), .A2(n4536), .ZN(n4534) );
  AND2_X1 U4448 ( .A1(n4536), .A2(n4535), .ZN(n4532) );
  AND2_X1 U4449 ( .A1(n4537), .A2(n4538), .ZN(n4535) );
  INV_X1 U4450 ( .A(n4539), .ZN(n4538) );
  AND2_X1 U4451 ( .A1(n4540), .A2(n4541), .ZN(n4539) );
  OR2_X1 U4452 ( .A1(n4541), .A2(n4540), .ZN(n4537) );
  INV_X1 U4453 ( .A(n3803), .ZN(n4432) );
  AND2_X1 U4454 ( .A1(a_5_), .A2(b_15_), .ZN(n3803) );
  OR2_X1 U4455 ( .A1(n4542), .A2(n4543), .ZN(n3799) );
  INV_X1 U4456 ( .A(n4544), .ZN(n4543) );
  OR2_X1 U4457 ( .A1(n4545), .A2(n4546), .ZN(n4544) );
  AND2_X1 U4458 ( .A1(n4546), .A2(n4545), .ZN(n4542) );
  AND2_X1 U4459 ( .A1(n4547), .A2(n4548), .ZN(n4545) );
  INV_X1 U4460 ( .A(n4549), .ZN(n4548) );
  AND2_X1 U4461 ( .A1(n4550), .A2(n4551), .ZN(n4549) );
  OR2_X1 U4462 ( .A1(n4551), .A2(n4550), .ZN(n4547) );
  INV_X1 U4463 ( .A(n3827), .ZN(n4428) );
  AND2_X1 U4464 ( .A1(a_4_), .A2(b_15_), .ZN(n3827) );
  OR2_X1 U4465 ( .A1(n4552), .A2(n4553), .ZN(n3823) );
  INV_X1 U4466 ( .A(n4554), .ZN(n4553) );
  OR2_X1 U4467 ( .A1(n4555), .A2(n4556), .ZN(n4554) );
  AND2_X1 U4468 ( .A1(n4556), .A2(n4555), .ZN(n4552) );
  AND2_X1 U4469 ( .A1(n4557), .A2(n4558), .ZN(n4555) );
  INV_X1 U4470 ( .A(n4559), .ZN(n4558) );
  AND2_X1 U4471 ( .A1(n4560), .A2(n4561), .ZN(n4559) );
  OR2_X1 U4472 ( .A1(n4561), .A2(n4560), .ZN(n4557) );
  INV_X1 U4473 ( .A(n3858), .ZN(n4424) );
  AND2_X1 U4474 ( .A1(a_3_), .A2(b_15_), .ZN(n3858) );
  OR2_X1 U4475 ( .A1(n4562), .A2(n4563), .ZN(n3854) );
  INV_X1 U4476 ( .A(n4564), .ZN(n4563) );
  OR2_X1 U4477 ( .A1(n4565), .A2(n4566), .ZN(n4564) );
  AND2_X1 U4478 ( .A1(n4566), .A2(n4565), .ZN(n4562) );
  AND2_X1 U4479 ( .A1(n4567), .A2(n4568), .ZN(n4565) );
  INV_X1 U4480 ( .A(n4569), .ZN(n4568) );
  AND2_X1 U4481 ( .A1(n4570), .A2(n4571), .ZN(n4569) );
  OR2_X1 U4482 ( .A1(n4571), .A2(n4570), .ZN(n4567) );
  INV_X1 U4483 ( .A(n3882), .ZN(n4420) );
  AND2_X1 U4484 ( .A1(a_2_), .A2(b_15_), .ZN(n3882) );
  OR2_X1 U4485 ( .A1(n4572), .A2(n4573), .ZN(n3878) );
  INV_X1 U4486 ( .A(n4574), .ZN(n4573) );
  OR2_X1 U4487 ( .A1(n4575), .A2(n4576), .ZN(n4574) );
  AND2_X1 U4488 ( .A1(n4576), .A2(n4575), .ZN(n4572) );
  AND2_X1 U4489 ( .A1(n4577), .A2(n4578), .ZN(n4575) );
  INV_X1 U4490 ( .A(n4579), .ZN(n4578) );
  AND2_X1 U4491 ( .A1(n4580), .A2(n4581), .ZN(n4579) );
  OR2_X1 U4492 ( .A1(n4581), .A2(n4580), .ZN(n4577) );
  INV_X1 U4493 ( .A(n3902), .ZN(n4416) );
  AND2_X1 U4494 ( .A1(a_1_), .A2(b_15_), .ZN(n3902) );
  OR2_X1 U4495 ( .A1(n4582), .A2(n4583), .ZN(n3898) );
  INV_X1 U4496 ( .A(n4584), .ZN(n4583) );
  OR2_X1 U4497 ( .A1(n4585), .A2(n4586), .ZN(n4584) );
  AND2_X1 U4498 ( .A1(n4586), .A2(n4585), .ZN(n4582) );
  AND2_X1 U4499 ( .A1(n4587), .A2(n4588), .ZN(n4585) );
  INV_X1 U4500 ( .A(n4589), .ZN(n4588) );
  AND2_X1 U4501 ( .A1(n4590), .A2(n4591), .ZN(n4589) );
  OR2_X1 U4502 ( .A1(n4591), .A2(n4590), .ZN(n4587) );
  OR2_X1 U4503 ( .A1(n3938), .A2(n3596), .ZN(n3925) );
  INV_X1 U4504 ( .A(b_15_), .ZN(n3596) );
  OR2_X1 U4505 ( .A1(n4592), .A2(n4593), .ZN(n3922) );
  INV_X1 U4506 ( .A(n4594), .ZN(n4593) );
  OR2_X1 U4507 ( .A1(n4595), .A2(n4596), .ZN(n4594) );
  AND2_X1 U4508 ( .A1(n4596), .A2(n4595), .ZN(n4592) );
  AND2_X1 U4509 ( .A1(n4597), .A2(n4598), .ZN(n4595) );
  INV_X1 U4510 ( .A(n4599), .ZN(n4598) );
  AND2_X1 U4511 ( .A1(n4600), .A2(n4601), .ZN(n4599) );
  OR2_X1 U4512 ( .A1(n4601), .A2(n4600), .ZN(n4597) );
  AND2_X1 U4513 ( .A1(n4397), .A2(n4396), .ZN(n3997) );
  INV_X1 U4514 ( .A(n3998), .ZN(n4396) );
  OR2_X1 U4515 ( .A1(n4602), .A2(n4002), .ZN(n3998) );
  INV_X1 U4516 ( .A(n4603), .ZN(n4002) );
  OR2_X1 U4517 ( .A1(n4604), .A2(n4605), .ZN(n4603) );
  AND2_X1 U4518 ( .A1(n4604), .A2(n4605), .ZN(n4602) );
  OR2_X1 U4519 ( .A1(n4606), .A2(n4607), .ZN(n4605) );
  AND2_X1 U4520 ( .A1(n4608), .A2(n4609), .ZN(n4607) );
  AND2_X1 U4521 ( .A1(n4610), .A2(n4611), .ZN(n4606) );
  OR2_X1 U4522 ( .A1(n4608), .A2(n4609), .ZN(n4611) );
  AND2_X1 U4523 ( .A1(n4612), .A2(n4613), .ZN(n4604) );
  INV_X1 U4524 ( .A(n4614), .ZN(n4613) );
  AND2_X1 U4525 ( .A1(n4615), .A2(n4616), .ZN(n4614) );
  OR2_X1 U4526 ( .A1(n4616), .A2(n4615), .ZN(n4612) );
  OR2_X1 U4527 ( .A1(n4617), .A2(n4618), .ZN(n4615) );
  INV_X1 U4528 ( .A(n4619), .ZN(n4618) );
  OR2_X1 U4529 ( .A1(n4620), .A2(n4621), .ZN(n4619) );
  AND2_X1 U4530 ( .A1(n4621), .A2(n4620), .ZN(n4617) );
  INV_X1 U4531 ( .A(n4622), .ZN(n4621) );
  INV_X1 U4532 ( .A(n3988), .ZN(n4397) );
  OR2_X1 U4533 ( .A1(n4398), .A2(n4399), .ZN(n3988) );
  OR2_X1 U4534 ( .A1(n4623), .A2(n4624), .ZN(n4399) );
  INV_X1 U4535 ( .A(n4625), .ZN(n4624) );
  OR2_X1 U4536 ( .A1(n4626), .A2(n4610), .ZN(n4625) );
  AND2_X1 U4537 ( .A1(n4610), .A2(n4626), .ZN(n4623) );
  AND2_X1 U4538 ( .A1(n4627), .A2(n4628), .ZN(n4626) );
  OR2_X1 U4539 ( .A1(n4608), .A2(n4629), .ZN(n4628) );
  INV_X1 U4540 ( .A(n4630), .ZN(n4627) );
  AND2_X1 U4541 ( .A1(n4629), .A2(n4608), .ZN(n4630) );
  OR2_X1 U4542 ( .A1(n3938), .A2(n3630), .ZN(n4608) );
  INV_X1 U4543 ( .A(n4609), .ZN(n4629) );
  OR2_X1 U4544 ( .A1(n4631), .A2(n4632), .ZN(n4609) );
  AND2_X1 U4545 ( .A1(n4633), .A2(n4634), .ZN(n4632) );
  AND2_X1 U4546 ( .A1(n4635), .A2(n4636), .ZN(n4631) );
  OR2_X1 U4547 ( .A1(n4633), .A2(n4634), .ZN(n4636) );
  INV_X1 U4548 ( .A(n4637), .ZN(n4633) );
  OR2_X1 U4549 ( .A1(n4638), .A2(n4639), .ZN(n4610) );
  INV_X1 U4550 ( .A(n4640), .ZN(n4639) );
  OR2_X1 U4551 ( .A1(n4641), .A2(n4642), .ZN(n4640) );
  AND2_X1 U4552 ( .A1(n4642), .A2(n4641), .ZN(n4638) );
  AND2_X1 U4553 ( .A1(n4643), .A2(n4644), .ZN(n4641) );
  INV_X1 U4554 ( .A(n4645), .ZN(n4644) );
  AND2_X1 U4555 ( .A1(n4646), .A2(n4647), .ZN(n4645) );
  OR2_X1 U4556 ( .A1(n4647), .A2(n4646), .ZN(n4643) );
  OR2_X1 U4557 ( .A1(n4648), .A2(n4649), .ZN(n4398) );
  AND2_X1 U4558 ( .A1(n4407), .A2(n4410), .ZN(n4649) );
  AND2_X1 U4559 ( .A1(n4403), .A2(n4650), .ZN(n4648) );
  OR2_X1 U4560 ( .A1(n4407), .A2(n4410), .ZN(n4650) );
  OR2_X1 U4561 ( .A1(n4651), .A2(n4652), .ZN(n4410) );
  AND2_X1 U4562 ( .A1(n4653), .A2(n4601), .ZN(n4652) );
  AND2_X1 U4563 ( .A1(n4596), .A2(n4654), .ZN(n4651) );
  OR2_X1 U4564 ( .A1(n4653), .A2(n4601), .ZN(n4654) );
  OR2_X1 U4565 ( .A1(n4655), .A2(n4656), .ZN(n4601) );
  AND2_X1 U4566 ( .A1(n4657), .A2(n4591), .ZN(n4656) );
  AND2_X1 U4567 ( .A1(n4586), .A2(n4658), .ZN(n4655) );
  OR2_X1 U4568 ( .A1(n4657), .A2(n4591), .ZN(n4658) );
  OR2_X1 U4569 ( .A1(n4659), .A2(n4660), .ZN(n4591) );
  AND2_X1 U4570 ( .A1(n4661), .A2(n4581), .ZN(n4660) );
  AND2_X1 U4571 ( .A1(n4576), .A2(n4662), .ZN(n4659) );
  OR2_X1 U4572 ( .A1(n4661), .A2(n4581), .ZN(n4662) );
  OR2_X1 U4573 ( .A1(n4663), .A2(n4664), .ZN(n4581) );
  AND2_X1 U4574 ( .A1(n4665), .A2(n4571), .ZN(n4664) );
  AND2_X1 U4575 ( .A1(n4566), .A2(n4666), .ZN(n4663) );
  OR2_X1 U4576 ( .A1(n4665), .A2(n4571), .ZN(n4666) );
  OR2_X1 U4577 ( .A1(n4667), .A2(n4668), .ZN(n4571) );
  AND2_X1 U4578 ( .A1(n4669), .A2(n4561), .ZN(n4668) );
  AND2_X1 U4579 ( .A1(n4556), .A2(n4670), .ZN(n4667) );
  OR2_X1 U4580 ( .A1(n4669), .A2(n4561), .ZN(n4670) );
  OR2_X1 U4581 ( .A1(n4671), .A2(n4672), .ZN(n4561) );
  AND2_X1 U4582 ( .A1(n4673), .A2(n4551), .ZN(n4672) );
  AND2_X1 U4583 ( .A1(n4546), .A2(n4674), .ZN(n4671) );
  OR2_X1 U4584 ( .A1(n4673), .A2(n4551), .ZN(n4674) );
  OR2_X1 U4585 ( .A1(n4675), .A2(n4676), .ZN(n4551) );
  AND2_X1 U4586 ( .A1(n4677), .A2(n4541), .ZN(n4676) );
  AND2_X1 U4587 ( .A1(n4536), .A2(n4678), .ZN(n4675) );
  OR2_X1 U4588 ( .A1(n4677), .A2(n4541), .ZN(n4678) );
  OR2_X1 U4589 ( .A1(n4679), .A2(n4680), .ZN(n4541) );
  AND2_X1 U4590 ( .A1(n4681), .A2(n4531), .ZN(n4680) );
  AND2_X1 U4591 ( .A1(n4526), .A2(n4682), .ZN(n4679) );
  OR2_X1 U4592 ( .A1(n4681), .A2(n4531), .ZN(n4682) );
  OR2_X1 U4593 ( .A1(n4683), .A2(n4684), .ZN(n4531) );
  AND2_X1 U4594 ( .A1(n4685), .A2(n4521), .ZN(n4684) );
  AND2_X1 U4595 ( .A1(n4516), .A2(n4686), .ZN(n4683) );
  OR2_X1 U4596 ( .A1(n4685), .A2(n4521), .ZN(n4686) );
  OR2_X1 U4597 ( .A1(n4687), .A2(n4688), .ZN(n4521) );
  AND2_X1 U4598 ( .A1(n4511), .A2(n4510), .ZN(n4688) );
  AND2_X1 U4599 ( .A1(n4505), .A2(n4689), .ZN(n4687) );
  OR2_X1 U4600 ( .A1(n4511), .A2(n4510), .ZN(n4689) );
  OR2_X1 U4601 ( .A1(n4690), .A2(n4691), .ZN(n4510) );
  AND2_X1 U4602 ( .A1(n4692), .A2(n4500), .ZN(n4691) );
  AND2_X1 U4603 ( .A1(n4495), .A2(n4693), .ZN(n4690) );
  OR2_X1 U4604 ( .A1(n4692), .A2(n4500), .ZN(n4693) );
  OR2_X1 U4605 ( .A1(n4694), .A2(n4695), .ZN(n4500) );
  AND2_X1 U4606 ( .A1(n4487), .A2(n4489), .ZN(n4695) );
  AND2_X1 U4607 ( .A1(n4484), .A2(n4696), .ZN(n4694) );
  OR2_X1 U4608 ( .A1(n4487), .A2(n4489), .ZN(n4696) );
  OR2_X1 U4609 ( .A1(n4697), .A2(n4698), .ZN(n4489) );
  AND2_X1 U4610 ( .A1(n4472), .A2(n4477), .ZN(n4698) );
  AND2_X1 U4611 ( .A1(n4476), .A2(n4699), .ZN(n4697) );
  OR2_X1 U4612 ( .A1(n4472), .A2(n4477), .ZN(n4699) );
  INV_X1 U4613 ( .A(n4478), .ZN(n4477) );
  AND3_X1 U4614 ( .A1(n3975), .A2(b_13_), .A3(b_14_), .ZN(n4478) );
  OR2_X1 U4615 ( .A1(n3631), .A2(n3593), .ZN(n4472) );
  INV_X1 U4616 ( .A(n4479), .ZN(n4476) );
  OR2_X1 U4617 ( .A1(n4700), .A2(n4701), .ZN(n4479) );
  AND2_X1 U4618 ( .A1(b_13_), .A2(n4702), .ZN(n4701) );
  OR2_X1 U4619 ( .A1(n4703), .A2(n3592), .ZN(n4702) );
  AND2_X1 U4620 ( .A1(a_14_), .A2(n4704), .ZN(n4703) );
  AND2_X1 U4621 ( .A1(b_12_), .A2(n4705), .ZN(n4700) );
  OR2_X1 U4622 ( .A1(n4706), .A2(n3595), .ZN(n4705) );
  AND2_X1 U4623 ( .A1(a_15_), .A2(n3630), .ZN(n4706) );
  INV_X1 U4624 ( .A(n4490), .ZN(n4487) );
  AND2_X1 U4625 ( .A1(a_12_), .A2(b_14_), .ZN(n4490) );
  OR2_X1 U4626 ( .A1(n4707), .A2(n4708), .ZN(n4484) );
  AND2_X1 U4627 ( .A1(n4709), .A2(n3972), .ZN(n4708) );
  INV_X1 U4628 ( .A(n4710), .ZN(n4707) );
  OR2_X1 U4629 ( .A1(n4709), .A2(n3972), .ZN(n4710) );
  OR2_X1 U4630 ( .A1(n4711), .A2(n4712), .ZN(n4709) );
  AND2_X1 U4631 ( .A1(n4713), .A2(n4714), .ZN(n4712) );
  AND2_X1 U4632 ( .A1(n4715), .A2(n4716), .ZN(n4711) );
  INV_X1 U4633 ( .A(n4499), .ZN(n4692) );
  AND2_X1 U4634 ( .A1(a_11_), .A2(b_14_), .ZN(n4499) );
  OR2_X1 U4635 ( .A1(n4717), .A2(n4718), .ZN(n4495) );
  INV_X1 U4636 ( .A(n4719), .ZN(n4718) );
  OR2_X1 U4637 ( .A1(n4720), .A2(n4721), .ZN(n4719) );
  AND2_X1 U4638 ( .A1(n4721), .A2(n4720), .ZN(n4717) );
  AND2_X1 U4639 ( .A1(n4722), .A2(n4723), .ZN(n4720) );
  INV_X1 U4640 ( .A(n4724), .ZN(n4723) );
  AND2_X1 U4641 ( .A1(n4725), .A2(n4726), .ZN(n4724) );
  OR2_X1 U4642 ( .A1(n4726), .A2(n4725), .ZN(n4722) );
  OR2_X1 U4643 ( .A1(n3964), .A2(n3593), .ZN(n4511) );
  OR2_X1 U4644 ( .A1(n4727), .A2(n4728), .ZN(n4505) );
  INV_X1 U4645 ( .A(n4729), .ZN(n4728) );
  OR2_X1 U4646 ( .A1(n4730), .A2(n4731), .ZN(n4729) );
  AND2_X1 U4647 ( .A1(n4731), .A2(n4730), .ZN(n4727) );
  AND2_X1 U4648 ( .A1(n4732), .A2(n4733), .ZN(n4730) );
  INV_X1 U4649 ( .A(n4734), .ZN(n4733) );
  AND2_X1 U4650 ( .A1(n4735), .A2(n4736), .ZN(n4734) );
  OR2_X1 U4651 ( .A1(n4736), .A2(n4735), .ZN(n4732) );
  INV_X1 U4652 ( .A(n4520), .ZN(n4685) );
  AND2_X1 U4653 ( .A1(a_9_), .A2(b_14_), .ZN(n4520) );
  OR2_X1 U4654 ( .A1(n4737), .A2(n4738), .ZN(n4516) );
  INV_X1 U4655 ( .A(n4739), .ZN(n4738) );
  OR2_X1 U4656 ( .A1(n4740), .A2(n4741), .ZN(n4739) );
  AND2_X1 U4657 ( .A1(n4741), .A2(n4740), .ZN(n4737) );
  AND2_X1 U4658 ( .A1(n4742), .A2(n4743), .ZN(n4740) );
  INV_X1 U4659 ( .A(n4744), .ZN(n4743) );
  AND2_X1 U4660 ( .A1(n4745), .A2(n4746), .ZN(n4744) );
  OR2_X1 U4661 ( .A1(n4746), .A2(n4745), .ZN(n4742) );
  INV_X1 U4662 ( .A(n4747), .ZN(n4745) );
  INV_X1 U4663 ( .A(n4530), .ZN(n4681) );
  AND2_X1 U4664 ( .A1(a_8_), .A2(b_14_), .ZN(n4530) );
  OR2_X1 U4665 ( .A1(n4748), .A2(n4749), .ZN(n4526) );
  INV_X1 U4666 ( .A(n4750), .ZN(n4749) );
  OR2_X1 U4667 ( .A1(n4751), .A2(n4752), .ZN(n4750) );
  AND2_X1 U4668 ( .A1(n4752), .A2(n4751), .ZN(n4748) );
  AND2_X1 U4669 ( .A1(n4753), .A2(n4754), .ZN(n4751) );
  INV_X1 U4670 ( .A(n4755), .ZN(n4754) );
  AND2_X1 U4671 ( .A1(n4756), .A2(n4757), .ZN(n4755) );
  OR2_X1 U4672 ( .A1(n4757), .A2(n4756), .ZN(n4753) );
  INV_X1 U4673 ( .A(n4540), .ZN(n4677) );
  AND2_X1 U4674 ( .A1(a_7_), .A2(b_14_), .ZN(n4540) );
  OR2_X1 U4675 ( .A1(n4758), .A2(n4759), .ZN(n4536) );
  INV_X1 U4676 ( .A(n4760), .ZN(n4759) );
  OR2_X1 U4677 ( .A1(n4761), .A2(n4762), .ZN(n4760) );
  AND2_X1 U4678 ( .A1(n4762), .A2(n4761), .ZN(n4758) );
  AND2_X1 U4679 ( .A1(n4763), .A2(n4764), .ZN(n4761) );
  INV_X1 U4680 ( .A(n4765), .ZN(n4764) );
  AND2_X1 U4681 ( .A1(n4766), .A2(n4767), .ZN(n4765) );
  OR2_X1 U4682 ( .A1(n4767), .A2(n4766), .ZN(n4763) );
  INV_X1 U4683 ( .A(n4550), .ZN(n4673) );
  AND2_X1 U4684 ( .A1(a_6_), .A2(b_14_), .ZN(n4550) );
  OR2_X1 U4685 ( .A1(n4768), .A2(n4769), .ZN(n4546) );
  INV_X1 U4686 ( .A(n4770), .ZN(n4769) );
  OR2_X1 U4687 ( .A1(n4771), .A2(n4772), .ZN(n4770) );
  AND2_X1 U4688 ( .A1(n4772), .A2(n4771), .ZN(n4768) );
  AND2_X1 U4689 ( .A1(n4773), .A2(n4774), .ZN(n4771) );
  INV_X1 U4690 ( .A(n4775), .ZN(n4774) );
  AND2_X1 U4691 ( .A1(n4776), .A2(n4777), .ZN(n4775) );
  OR2_X1 U4692 ( .A1(n4777), .A2(n4776), .ZN(n4773) );
  INV_X1 U4693 ( .A(n4560), .ZN(n4669) );
  AND2_X1 U4694 ( .A1(a_5_), .A2(b_14_), .ZN(n4560) );
  OR2_X1 U4695 ( .A1(n4778), .A2(n4779), .ZN(n4556) );
  INV_X1 U4696 ( .A(n4780), .ZN(n4779) );
  OR2_X1 U4697 ( .A1(n4781), .A2(n4782), .ZN(n4780) );
  AND2_X1 U4698 ( .A1(n4782), .A2(n4781), .ZN(n4778) );
  AND2_X1 U4699 ( .A1(n4783), .A2(n4784), .ZN(n4781) );
  INV_X1 U4700 ( .A(n4785), .ZN(n4784) );
  AND2_X1 U4701 ( .A1(n4786), .A2(n4787), .ZN(n4785) );
  OR2_X1 U4702 ( .A1(n4787), .A2(n4786), .ZN(n4783) );
  INV_X1 U4703 ( .A(n4570), .ZN(n4665) );
  AND2_X1 U4704 ( .A1(a_4_), .A2(b_14_), .ZN(n4570) );
  OR2_X1 U4705 ( .A1(n4788), .A2(n4789), .ZN(n4566) );
  INV_X1 U4706 ( .A(n4790), .ZN(n4789) );
  OR2_X1 U4707 ( .A1(n4791), .A2(n4792), .ZN(n4790) );
  AND2_X1 U4708 ( .A1(n4792), .A2(n4791), .ZN(n4788) );
  AND2_X1 U4709 ( .A1(n4793), .A2(n4794), .ZN(n4791) );
  INV_X1 U4710 ( .A(n4795), .ZN(n4794) );
  AND2_X1 U4711 ( .A1(n4796), .A2(n4797), .ZN(n4795) );
  OR2_X1 U4712 ( .A1(n4797), .A2(n4796), .ZN(n4793) );
  INV_X1 U4713 ( .A(n4580), .ZN(n4661) );
  AND2_X1 U4714 ( .A1(a_3_), .A2(b_14_), .ZN(n4580) );
  OR2_X1 U4715 ( .A1(n4798), .A2(n4799), .ZN(n4576) );
  INV_X1 U4716 ( .A(n4800), .ZN(n4799) );
  OR2_X1 U4717 ( .A1(n4801), .A2(n4802), .ZN(n4800) );
  AND2_X1 U4718 ( .A1(n4802), .A2(n4801), .ZN(n4798) );
  AND2_X1 U4719 ( .A1(n4803), .A2(n4804), .ZN(n4801) );
  INV_X1 U4720 ( .A(n4805), .ZN(n4804) );
  AND2_X1 U4721 ( .A1(n4806), .A2(n4807), .ZN(n4805) );
  OR2_X1 U4722 ( .A1(n4807), .A2(n4806), .ZN(n4803) );
  INV_X1 U4723 ( .A(n4590), .ZN(n4657) );
  AND2_X1 U4724 ( .A1(a_2_), .A2(b_14_), .ZN(n4590) );
  OR2_X1 U4725 ( .A1(n4808), .A2(n4809), .ZN(n4586) );
  INV_X1 U4726 ( .A(n4810), .ZN(n4809) );
  OR2_X1 U4727 ( .A1(n4811), .A2(n4812), .ZN(n4810) );
  AND2_X1 U4728 ( .A1(n4812), .A2(n4811), .ZN(n4808) );
  AND2_X1 U4729 ( .A1(n4813), .A2(n4814), .ZN(n4811) );
  INV_X1 U4730 ( .A(n4815), .ZN(n4814) );
  AND2_X1 U4731 ( .A1(n4816), .A2(n4817), .ZN(n4815) );
  OR2_X1 U4732 ( .A1(n4817), .A2(n4816), .ZN(n4813) );
  INV_X1 U4733 ( .A(n4600), .ZN(n4653) );
  AND2_X1 U4734 ( .A1(a_1_), .A2(b_14_), .ZN(n4600) );
  OR2_X1 U4735 ( .A1(n4818), .A2(n4819), .ZN(n4596) );
  INV_X1 U4736 ( .A(n4820), .ZN(n4819) );
  OR2_X1 U4737 ( .A1(n4821), .A2(n4822), .ZN(n4820) );
  AND2_X1 U4738 ( .A1(n4822), .A2(n4821), .ZN(n4818) );
  AND2_X1 U4739 ( .A1(n4823), .A2(n4824), .ZN(n4821) );
  INV_X1 U4740 ( .A(n4825), .ZN(n4824) );
  AND2_X1 U4741 ( .A1(n4826), .A2(n4827), .ZN(n4825) );
  OR2_X1 U4742 ( .A1(n4827), .A2(n4826), .ZN(n4823) );
  OR2_X1 U4743 ( .A1(n3938), .A2(n3593), .ZN(n4407) );
  INV_X1 U4744 ( .A(b_14_), .ZN(n3593) );
  OR2_X1 U4745 ( .A1(n4828), .A2(n4829), .ZN(n4403) );
  INV_X1 U4746 ( .A(n4830), .ZN(n4829) );
  OR2_X1 U4747 ( .A1(n4831), .A2(n4635), .ZN(n4830) );
  AND2_X1 U4748 ( .A1(n4635), .A2(n4831), .ZN(n4828) );
  AND2_X1 U4749 ( .A1(n4832), .A2(n4833), .ZN(n4831) );
  INV_X1 U4750 ( .A(n4834), .ZN(n4833) );
  AND2_X1 U4751 ( .A1(n4637), .A2(n4634), .ZN(n4834) );
  OR2_X1 U4752 ( .A1(n4634), .A2(n4637), .ZN(n4832) );
  AND2_X1 U4753 ( .A1(a_1_), .A2(b_13_), .ZN(n4637) );
  OR2_X1 U4754 ( .A1(n4835), .A2(n4836), .ZN(n4634) );
  AND2_X1 U4755 ( .A1(n4837), .A2(n4827), .ZN(n4836) );
  AND2_X1 U4756 ( .A1(n4822), .A2(n4838), .ZN(n4835) );
  OR2_X1 U4757 ( .A1(n4837), .A2(n4827), .ZN(n4838) );
  OR2_X1 U4758 ( .A1(n4839), .A2(n4840), .ZN(n4827) );
  AND2_X1 U4759 ( .A1(n4841), .A2(n4817), .ZN(n4840) );
  AND2_X1 U4760 ( .A1(n4812), .A2(n4842), .ZN(n4839) );
  OR2_X1 U4761 ( .A1(n4841), .A2(n4817), .ZN(n4842) );
  OR2_X1 U4762 ( .A1(n4843), .A2(n4844), .ZN(n4817) );
  AND2_X1 U4763 ( .A1(n4845), .A2(n4807), .ZN(n4844) );
  AND2_X1 U4764 ( .A1(n4802), .A2(n4846), .ZN(n4843) );
  OR2_X1 U4765 ( .A1(n4845), .A2(n4807), .ZN(n4846) );
  OR2_X1 U4766 ( .A1(n4847), .A2(n4848), .ZN(n4807) );
  AND2_X1 U4767 ( .A1(n4849), .A2(n4797), .ZN(n4848) );
  AND2_X1 U4768 ( .A1(n4792), .A2(n4850), .ZN(n4847) );
  OR2_X1 U4769 ( .A1(n4849), .A2(n4797), .ZN(n4850) );
  OR2_X1 U4770 ( .A1(n4851), .A2(n4852), .ZN(n4797) );
  AND2_X1 U4771 ( .A1(n4853), .A2(n4787), .ZN(n4852) );
  AND2_X1 U4772 ( .A1(n4782), .A2(n4854), .ZN(n4851) );
  OR2_X1 U4773 ( .A1(n4853), .A2(n4787), .ZN(n4854) );
  OR2_X1 U4774 ( .A1(n4855), .A2(n4856), .ZN(n4787) );
  AND2_X1 U4775 ( .A1(n4857), .A2(n4777), .ZN(n4856) );
  AND2_X1 U4776 ( .A1(n4772), .A2(n4858), .ZN(n4855) );
  OR2_X1 U4777 ( .A1(n4857), .A2(n4777), .ZN(n4858) );
  OR2_X1 U4778 ( .A1(n4859), .A2(n4860), .ZN(n4777) );
  AND2_X1 U4779 ( .A1(n4861), .A2(n4767), .ZN(n4860) );
  AND2_X1 U4780 ( .A1(n4762), .A2(n4862), .ZN(n4859) );
  OR2_X1 U4781 ( .A1(n4861), .A2(n4767), .ZN(n4862) );
  OR2_X1 U4782 ( .A1(n4863), .A2(n4864), .ZN(n4767) );
  AND2_X1 U4783 ( .A1(n4865), .A2(n4757), .ZN(n4864) );
  AND2_X1 U4784 ( .A1(n4752), .A2(n4866), .ZN(n4863) );
  OR2_X1 U4785 ( .A1(n4865), .A2(n4757), .ZN(n4866) );
  OR2_X1 U4786 ( .A1(n4867), .A2(n4868), .ZN(n4757) );
  AND2_X1 U4787 ( .A1(n4747), .A2(n4746), .ZN(n4868) );
  AND2_X1 U4788 ( .A1(n4741), .A2(n4869), .ZN(n4867) );
  OR2_X1 U4789 ( .A1(n4747), .A2(n4746), .ZN(n4869) );
  OR2_X1 U4790 ( .A1(n4870), .A2(n4871), .ZN(n4746) );
  AND2_X1 U4791 ( .A1(n4872), .A2(n4736), .ZN(n4871) );
  AND2_X1 U4792 ( .A1(n4731), .A2(n4873), .ZN(n4870) );
  OR2_X1 U4793 ( .A1(n4872), .A2(n4736), .ZN(n4873) );
  OR2_X1 U4794 ( .A1(n4874), .A2(n4875), .ZN(n4736) );
  AND2_X1 U4795 ( .A1(n4876), .A2(n4726), .ZN(n4875) );
  AND2_X1 U4796 ( .A1(n4721), .A2(n4877), .ZN(n4874) );
  OR2_X1 U4797 ( .A1(n4876), .A2(n4726), .ZN(n4877) );
  OR2_X1 U4798 ( .A1(n4878), .A2(n4879), .ZN(n4726) );
  AND2_X1 U4799 ( .A1(n3972), .A2(n4714), .ZN(n4879) );
  AND2_X1 U4800 ( .A1(n4713), .A2(n4880), .ZN(n4878) );
  OR2_X1 U4801 ( .A1(n3972), .A2(n4714), .ZN(n4880) );
  INV_X1 U4802 ( .A(n4715), .ZN(n4714) );
  AND3_X1 U4803 ( .A1(n3975), .A2(b_12_), .A3(b_13_), .ZN(n4715) );
  INV_X1 U4804 ( .A(n3634), .ZN(n3972) );
  AND2_X1 U4805 ( .A1(a_13_), .A2(b_13_), .ZN(n3634) );
  INV_X1 U4806 ( .A(n4716), .ZN(n4713) );
  OR2_X1 U4807 ( .A1(n4881), .A2(n4882), .ZN(n4716) );
  AND2_X1 U4808 ( .A1(b_12_), .A2(n4883), .ZN(n4882) );
  OR2_X1 U4809 ( .A1(n4884), .A2(n3592), .ZN(n4883) );
  AND2_X1 U4810 ( .A1(a_14_), .A2(n3678), .ZN(n4884) );
  AND2_X1 U4811 ( .A1(b_11_), .A2(n4885), .ZN(n4881) );
  OR2_X1 U4812 ( .A1(n4886), .A2(n3595), .ZN(n4885) );
  AND2_X1 U4813 ( .A1(a_15_), .A2(n4704), .ZN(n4886) );
  INV_X1 U4814 ( .A(n4725), .ZN(n4876) );
  AND2_X1 U4815 ( .A1(a_12_), .A2(b_13_), .ZN(n4725) );
  OR2_X1 U4816 ( .A1(n4887), .A2(n4888), .ZN(n4721) );
  AND2_X1 U4817 ( .A1(n4889), .A2(n4890), .ZN(n4888) );
  INV_X1 U4818 ( .A(n4891), .ZN(n4887) );
  OR2_X1 U4819 ( .A1(n4889), .A2(n4890), .ZN(n4891) );
  OR2_X1 U4820 ( .A1(n4892), .A2(n4893), .ZN(n4889) );
  AND2_X1 U4821 ( .A1(n4894), .A2(n4895), .ZN(n4893) );
  AND2_X1 U4822 ( .A1(n4896), .A2(n4897), .ZN(n4892) );
  INV_X1 U4823 ( .A(n4735), .ZN(n4872) );
  AND2_X1 U4824 ( .A1(a_11_), .A2(b_13_), .ZN(n4735) );
  OR2_X1 U4825 ( .A1(n4898), .A2(n4899), .ZN(n4731) );
  INV_X1 U4826 ( .A(n4900), .ZN(n4899) );
  OR2_X1 U4827 ( .A1(n4901), .A2(n4902), .ZN(n4900) );
  AND2_X1 U4828 ( .A1(n4902), .A2(n4901), .ZN(n4898) );
  AND2_X1 U4829 ( .A1(n4903), .A2(n4904), .ZN(n4901) );
  INV_X1 U4830 ( .A(n4905), .ZN(n4904) );
  AND2_X1 U4831 ( .A1(n3656), .A2(n4906), .ZN(n4905) );
  OR2_X1 U4832 ( .A1(n4906), .A2(n3656), .ZN(n4903) );
  OR2_X1 U4833 ( .A1(n3964), .A2(n3630), .ZN(n4747) );
  INV_X1 U4834 ( .A(b_13_), .ZN(n3630) );
  OR2_X1 U4835 ( .A1(n4907), .A2(n4908), .ZN(n4741) );
  INV_X1 U4836 ( .A(n4909), .ZN(n4908) );
  OR2_X1 U4837 ( .A1(n4910), .A2(n4911), .ZN(n4909) );
  AND2_X1 U4838 ( .A1(n4911), .A2(n4910), .ZN(n4907) );
  AND2_X1 U4839 ( .A1(n4912), .A2(n4913), .ZN(n4910) );
  INV_X1 U4840 ( .A(n4914), .ZN(n4913) );
  AND2_X1 U4841 ( .A1(n4915), .A2(n4916), .ZN(n4914) );
  OR2_X1 U4842 ( .A1(n4916), .A2(n4915), .ZN(n4912) );
  INV_X1 U4843 ( .A(n4756), .ZN(n4865) );
  AND2_X1 U4844 ( .A1(a_9_), .A2(b_13_), .ZN(n4756) );
  OR2_X1 U4845 ( .A1(n4917), .A2(n4918), .ZN(n4752) );
  INV_X1 U4846 ( .A(n4919), .ZN(n4918) );
  OR2_X1 U4847 ( .A1(n4920), .A2(n4921), .ZN(n4919) );
  AND2_X1 U4848 ( .A1(n4921), .A2(n4920), .ZN(n4917) );
  AND2_X1 U4849 ( .A1(n4922), .A2(n4923), .ZN(n4920) );
  INV_X1 U4850 ( .A(n4924), .ZN(n4923) );
  AND2_X1 U4851 ( .A1(n4925), .A2(n4926), .ZN(n4924) );
  OR2_X1 U4852 ( .A1(n4926), .A2(n4925), .ZN(n4922) );
  INV_X1 U4853 ( .A(n4927), .ZN(n4925) );
  INV_X1 U4854 ( .A(n4766), .ZN(n4861) );
  AND2_X1 U4855 ( .A1(a_8_), .A2(b_13_), .ZN(n4766) );
  OR2_X1 U4856 ( .A1(n4928), .A2(n4929), .ZN(n4762) );
  INV_X1 U4857 ( .A(n4930), .ZN(n4929) );
  OR2_X1 U4858 ( .A1(n4931), .A2(n4932), .ZN(n4930) );
  AND2_X1 U4859 ( .A1(n4932), .A2(n4931), .ZN(n4928) );
  AND2_X1 U4860 ( .A1(n4933), .A2(n4934), .ZN(n4931) );
  INV_X1 U4861 ( .A(n4935), .ZN(n4934) );
  AND2_X1 U4862 ( .A1(n4936), .A2(n4937), .ZN(n4935) );
  OR2_X1 U4863 ( .A1(n4937), .A2(n4936), .ZN(n4933) );
  INV_X1 U4864 ( .A(n4776), .ZN(n4857) );
  AND2_X1 U4865 ( .A1(a_7_), .A2(b_13_), .ZN(n4776) );
  OR2_X1 U4866 ( .A1(n4938), .A2(n4939), .ZN(n4772) );
  INV_X1 U4867 ( .A(n4940), .ZN(n4939) );
  OR2_X1 U4868 ( .A1(n4941), .A2(n4942), .ZN(n4940) );
  AND2_X1 U4869 ( .A1(n4942), .A2(n4941), .ZN(n4938) );
  AND2_X1 U4870 ( .A1(n4943), .A2(n4944), .ZN(n4941) );
  INV_X1 U4871 ( .A(n4945), .ZN(n4944) );
  AND2_X1 U4872 ( .A1(n4946), .A2(n4947), .ZN(n4945) );
  OR2_X1 U4873 ( .A1(n4947), .A2(n4946), .ZN(n4943) );
  INV_X1 U4874 ( .A(n4786), .ZN(n4853) );
  AND2_X1 U4875 ( .A1(a_6_), .A2(b_13_), .ZN(n4786) );
  OR2_X1 U4876 ( .A1(n4948), .A2(n4949), .ZN(n4782) );
  INV_X1 U4877 ( .A(n4950), .ZN(n4949) );
  OR2_X1 U4878 ( .A1(n4951), .A2(n4952), .ZN(n4950) );
  AND2_X1 U4879 ( .A1(n4952), .A2(n4951), .ZN(n4948) );
  AND2_X1 U4880 ( .A1(n4953), .A2(n4954), .ZN(n4951) );
  INV_X1 U4881 ( .A(n4955), .ZN(n4954) );
  AND2_X1 U4882 ( .A1(n4956), .A2(n4957), .ZN(n4955) );
  OR2_X1 U4883 ( .A1(n4957), .A2(n4956), .ZN(n4953) );
  INV_X1 U4884 ( .A(n4796), .ZN(n4849) );
  AND2_X1 U4885 ( .A1(a_5_), .A2(b_13_), .ZN(n4796) );
  OR2_X1 U4886 ( .A1(n4958), .A2(n4959), .ZN(n4792) );
  INV_X1 U4887 ( .A(n4960), .ZN(n4959) );
  OR2_X1 U4888 ( .A1(n4961), .A2(n4962), .ZN(n4960) );
  AND2_X1 U4889 ( .A1(n4962), .A2(n4961), .ZN(n4958) );
  AND2_X1 U4890 ( .A1(n4963), .A2(n4964), .ZN(n4961) );
  INV_X1 U4891 ( .A(n4965), .ZN(n4964) );
  AND2_X1 U4892 ( .A1(n4966), .A2(n4967), .ZN(n4965) );
  OR2_X1 U4893 ( .A1(n4967), .A2(n4966), .ZN(n4963) );
  INV_X1 U4894 ( .A(n4806), .ZN(n4845) );
  AND2_X1 U4895 ( .A1(a_4_), .A2(b_13_), .ZN(n4806) );
  OR2_X1 U4896 ( .A1(n4968), .A2(n4969), .ZN(n4802) );
  INV_X1 U4897 ( .A(n4970), .ZN(n4969) );
  OR2_X1 U4898 ( .A1(n4971), .A2(n4972), .ZN(n4970) );
  AND2_X1 U4899 ( .A1(n4972), .A2(n4971), .ZN(n4968) );
  AND2_X1 U4900 ( .A1(n4973), .A2(n4974), .ZN(n4971) );
  INV_X1 U4901 ( .A(n4975), .ZN(n4974) );
  AND2_X1 U4902 ( .A1(n4976), .A2(n4977), .ZN(n4975) );
  OR2_X1 U4903 ( .A1(n4977), .A2(n4976), .ZN(n4973) );
  INV_X1 U4904 ( .A(n4816), .ZN(n4841) );
  AND2_X1 U4905 ( .A1(a_3_), .A2(b_13_), .ZN(n4816) );
  OR2_X1 U4906 ( .A1(n4978), .A2(n4979), .ZN(n4812) );
  INV_X1 U4907 ( .A(n4980), .ZN(n4979) );
  OR2_X1 U4908 ( .A1(n4981), .A2(n4982), .ZN(n4980) );
  AND2_X1 U4909 ( .A1(n4982), .A2(n4981), .ZN(n4978) );
  AND2_X1 U4910 ( .A1(n4983), .A2(n4984), .ZN(n4981) );
  INV_X1 U4911 ( .A(n4985), .ZN(n4984) );
  AND2_X1 U4912 ( .A1(n4986), .A2(n4987), .ZN(n4985) );
  OR2_X1 U4913 ( .A1(n4987), .A2(n4986), .ZN(n4983) );
  INV_X1 U4914 ( .A(n4826), .ZN(n4837) );
  AND2_X1 U4915 ( .A1(a_2_), .A2(b_13_), .ZN(n4826) );
  OR2_X1 U4916 ( .A1(n4988), .A2(n4989), .ZN(n4822) );
  INV_X1 U4917 ( .A(n4990), .ZN(n4989) );
  OR2_X1 U4918 ( .A1(n4991), .A2(n4992), .ZN(n4990) );
  AND2_X1 U4919 ( .A1(n4992), .A2(n4991), .ZN(n4988) );
  AND2_X1 U4920 ( .A1(n4993), .A2(n4994), .ZN(n4991) );
  INV_X1 U4921 ( .A(n4995), .ZN(n4994) );
  AND2_X1 U4922 ( .A1(n4996), .A2(n4997), .ZN(n4995) );
  OR2_X1 U4923 ( .A1(n4997), .A2(n4996), .ZN(n4993) );
  OR2_X1 U4924 ( .A1(n4998), .A2(n4999), .ZN(n4635) );
  INV_X1 U4925 ( .A(n5000), .ZN(n4999) );
  OR2_X1 U4926 ( .A1(n5001), .A2(n5002), .ZN(n5000) );
  AND2_X1 U4927 ( .A1(n5002), .A2(n5001), .ZN(n4998) );
  AND2_X1 U4928 ( .A1(n5003), .A2(n5004), .ZN(n5001) );
  INV_X1 U4929 ( .A(n5005), .ZN(n5004) );
  AND2_X1 U4930 ( .A1(n5006), .A2(n5007), .ZN(n5005) );
  OR2_X1 U4931 ( .A1(n5007), .A2(n5006), .ZN(n5003) );
  INV_X1 U4932 ( .A(n4006), .ZN(n4009) );
  OR2_X1 U4933 ( .A1(n5008), .A2(n4013), .ZN(n4006) );
  INV_X1 U4934 ( .A(n5009), .ZN(n4013) );
  OR2_X1 U4935 ( .A1(n5010), .A2(n5011), .ZN(n5009) );
  AND2_X1 U4936 ( .A1(n5010), .A2(n5011), .ZN(n5008) );
  OR2_X1 U4937 ( .A1(n5012), .A2(n5013), .ZN(n5011) );
  AND2_X1 U4938 ( .A1(n4620), .A2(n4622), .ZN(n5013) );
  AND2_X1 U4939 ( .A1(n4616), .A2(n5014), .ZN(n5012) );
  OR2_X1 U4940 ( .A1(n4622), .A2(n4620), .ZN(n5014) );
  OR2_X1 U4941 ( .A1(n3938), .A2(n4704), .ZN(n4620) );
  OR2_X1 U4942 ( .A1(n5015), .A2(n5016), .ZN(n4622) );
  AND2_X1 U4943 ( .A1(n5017), .A2(n4647), .ZN(n5016) );
  AND2_X1 U4944 ( .A1(n4642), .A2(n5018), .ZN(n5015) );
  OR2_X1 U4945 ( .A1(n4647), .A2(n5017), .ZN(n5018) );
  INV_X1 U4946 ( .A(n4646), .ZN(n5017) );
  AND2_X1 U4947 ( .A1(a_1_), .A2(b_12_), .ZN(n4646) );
  OR2_X1 U4948 ( .A1(n5019), .A2(n5020), .ZN(n4647) );
  AND2_X1 U4949 ( .A1(n5021), .A2(n5007), .ZN(n5020) );
  AND2_X1 U4950 ( .A1(n5002), .A2(n5022), .ZN(n5019) );
  OR2_X1 U4951 ( .A1(n5007), .A2(n5021), .ZN(n5022) );
  INV_X1 U4952 ( .A(n5006), .ZN(n5021) );
  AND2_X1 U4953 ( .A1(a_2_), .A2(b_12_), .ZN(n5006) );
  OR2_X1 U4954 ( .A1(n5023), .A2(n5024), .ZN(n5007) );
  AND2_X1 U4955 ( .A1(n5025), .A2(n4997), .ZN(n5024) );
  AND2_X1 U4956 ( .A1(n4992), .A2(n5026), .ZN(n5023) );
  OR2_X1 U4957 ( .A1(n4997), .A2(n5025), .ZN(n5026) );
  INV_X1 U4958 ( .A(n4996), .ZN(n5025) );
  AND2_X1 U4959 ( .A1(a_3_), .A2(b_12_), .ZN(n4996) );
  OR2_X1 U4960 ( .A1(n5027), .A2(n5028), .ZN(n4997) );
  AND2_X1 U4961 ( .A1(n5029), .A2(n4987), .ZN(n5028) );
  AND2_X1 U4962 ( .A1(n4982), .A2(n5030), .ZN(n5027) );
  OR2_X1 U4963 ( .A1(n4987), .A2(n5029), .ZN(n5030) );
  INV_X1 U4964 ( .A(n4986), .ZN(n5029) );
  AND2_X1 U4965 ( .A1(a_4_), .A2(b_12_), .ZN(n4986) );
  OR2_X1 U4966 ( .A1(n5031), .A2(n5032), .ZN(n4987) );
  AND2_X1 U4967 ( .A1(n5033), .A2(n4977), .ZN(n5032) );
  AND2_X1 U4968 ( .A1(n4972), .A2(n5034), .ZN(n5031) );
  OR2_X1 U4969 ( .A1(n4977), .A2(n5033), .ZN(n5034) );
  INV_X1 U4970 ( .A(n4976), .ZN(n5033) );
  AND2_X1 U4971 ( .A1(a_5_), .A2(b_12_), .ZN(n4976) );
  OR2_X1 U4972 ( .A1(n5035), .A2(n5036), .ZN(n4977) );
  AND2_X1 U4973 ( .A1(n5037), .A2(n4967), .ZN(n5036) );
  AND2_X1 U4974 ( .A1(n4962), .A2(n5038), .ZN(n5035) );
  OR2_X1 U4975 ( .A1(n4967), .A2(n5037), .ZN(n5038) );
  INV_X1 U4976 ( .A(n4966), .ZN(n5037) );
  AND2_X1 U4977 ( .A1(a_6_), .A2(b_12_), .ZN(n4966) );
  OR2_X1 U4978 ( .A1(n5039), .A2(n5040), .ZN(n4967) );
  AND2_X1 U4979 ( .A1(n5041), .A2(n4957), .ZN(n5040) );
  AND2_X1 U4980 ( .A1(n4952), .A2(n5042), .ZN(n5039) );
  OR2_X1 U4981 ( .A1(n4957), .A2(n5041), .ZN(n5042) );
  INV_X1 U4982 ( .A(n4956), .ZN(n5041) );
  AND2_X1 U4983 ( .A1(a_7_), .A2(b_12_), .ZN(n4956) );
  OR2_X1 U4984 ( .A1(n5043), .A2(n5044), .ZN(n4957) );
  AND2_X1 U4985 ( .A1(n5045), .A2(n4947), .ZN(n5044) );
  AND2_X1 U4986 ( .A1(n4942), .A2(n5046), .ZN(n5043) );
  OR2_X1 U4987 ( .A1(n4947), .A2(n5045), .ZN(n5046) );
  INV_X1 U4988 ( .A(n4946), .ZN(n5045) );
  AND2_X1 U4989 ( .A1(a_8_), .A2(b_12_), .ZN(n4946) );
  OR2_X1 U4990 ( .A1(n5047), .A2(n5048), .ZN(n4947) );
  AND2_X1 U4991 ( .A1(n5049), .A2(n4937), .ZN(n5048) );
  AND2_X1 U4992 ( .A1(n4932), .A2(n5050), .ZN(n5047) );
  OR2_X1 U4993 ( .A1(n4937), .A2(n5049), .ZN(n5050) );
  INV_X1 U4994 ( .A(n4936), .ZN(n5049) );
  AND2_X1 U4995 ( .A1(a_9_), .A2(b_12_), .ZN(n4936) );
  OR2_X1 U4996 ( .A1(n5051), .A2(n5052), .ZN(n4937) );
  AND2_X1 U4997 ( .A1(n4927), .A2(n4926), .ZN(n5052) );
  AND2_X1 U4998 ( .A1(n4921), .A2(n5053), .ZN(n5051) );
  OR2_X1 U4999 ( .A1(n4926), .A2(n4927), .ZN(n5053) );
  OR2_X1 U5000 ( .A1(n3964), .A2(n4704), .ZN(n4927) );
  OR2_X1 U5001 ( .A1(n5054), .A2(n5055), .ZN(n4926) );
  AND2_X1 U5002 ( .A1(n5056), .A2(n4916), .ZN(n5055) );
  AND2_X1 U5003 ( .A1(n4911), .A2(n5057), .ZN(n5054) );
  OR2_X1 U5004 ( .A1(n4916), .A2(n5056), .ZN(n5057) );
  INV_X1 U5005 ( .A(n4915), .ZN(n5056) );
  AND2_X1 U5006 ( .A1(a_11_), .A2(b_12_), .ZN(n4915) );
  OR2_X1 U5007 ( .A1(n5058), .A2(n5059), .ZN(n4916) );
  AND2_X1 U5008 ( .A1(n3970), .A2(n4906), .ZN(n5059) );
  AND2_X1 U5009 ( .A1(n4902), .A2(n5060), .ZN(n5058) );
  OR2_X1 U5010 ( .A1(n4906), .A2(n3970), .ZN(n5060) );
  INV_X1 U5011 ( .A(n3656), .ZN(n3970) );
  AND2_X1 U5012 ( .A1(a_12_), .A2(b_12_), .ZN(n3656) );
  OR2_X1 U5013 ( .A1(n5061), .A2(n5062), .ZN(n4906) );
  AND2_X1 U5014 ( .A1(n4890), .A2(n4895), .ZN(n5062) );
  AND2_X1 U5015 ( .A1(n4894), .A2(n5063), .ZN(n5061) );
  OR2_X1 U5016 ( .A1(n4895), .A2(n4890), .ZN(n5063) );
  OR2_X1 U5017 ( .A1(n3631), .A2(n4704), .ZN(n4890) );
  INV_X1 U5018 ( .A(b_12_), .ZN(n4704) );
  INV_X1 U5019 ( .A(n4896), .ZN(n4895) );
  AND3_X1 U5020 ( .A1(n3975), .A2(b_11_), .A3(b_12_), .ZN(n4896) );
  INV_X1 U5021 ( .A(n4897), .ZN(n4894) );
  OR2_X1 U5022 ( .A1(n5064), .A2(n5065), .ZN(n4897) );
  AND2_X1 U5023 ( .A1(b_11_), .A2(n5066), .ZN(n5065) );
  OR2_X1 U5024 ( .A1(n5067), .A2(n3592), .ZN(n5066) );
  AND2_X1 U5025 ( .A1(a_14_), .A2(n3965), .ZN(n5067) );
  AND2_X1 U5026 ( .A1(b_10_), .A2(n5068), .ZN(n5064) );
  OR2_X1 U5027 ( .A1(n5069), .A2(n3595), .ZN(n5068) );
  AND2_X1 U5028 ( .A1(a_15_), .A2(n3678), .ZN(n5069) );
  OR2_X1 U5029 ( .A1(n5070), .A2(n5071), .ZN(n4902) );
  AND2_X1 U5030 ( .A1(n5072), .A2(n5073), .ZN(n5071) );
  INV_X1 U5031 ( .A(n5074), .ZN(n5070) );
  OR2_X1 U5032 ( .A1(n5072), .A2(n5073), .ZN(n5074) );
  OR2_X1 U5033 ( .A1(n5075), .A2(n5076), .ZN(n5072) );
  AND2_X1 U5034 ( .A1(n5077), .A2(n5078), .ZN(n5076) );
  AND2_X1 U5035 ( .A1(n5079), .A2(n5080), .ZN(n5075) );
  OR2_X1 U5036 ( .A1(n5081), .A2(n5082), .ZN(n4911) );
  INV_X1 U5037 ( .A(n5083), .ZN(n5082) );
  OR2_X1 U5038 ( .A1(n5084), .A2(n5085), .ZN(n5083) );
  AND2_X1 U5039 ( .A1(n5085), .A2(n5084), .ZN(n5081) );
  AND2_X1 U5040 ( .A1(n5086), .A2(n5087), .ZN(n5084) );
  INV_X1 U5041 ( .A(n5088), .ZN(n5087) );
  AND2_X1 U5042 ( .A1(n5089), .A2(n5090), .ZN(n5088) );
  OR2_X1 U5043 ( .A1(n5090), .A2(n5089), .ZN(n5086) );
  OR2_X1 U5044 ( .A1(n5091), .A2(n5092), .ZN(n4921) );
  INV_X1 U5045 ( .A(n5093), .ZN(n5092) );
  OR2_X1 U5046 ( .A1(n5094), .A2(n5095), .ZN(n5093) );
  AND2_X1 U5047 ( .A1(n5095), .A2(n5094), .ZN(n5091) );
  AND2_X1 U5048 ( .A1(n5096), .A2(n5097), .ZN(n5094) );
  INV_X1 U5049 ( .A(n5098), .ZN(n5097) );
  AND2_X1 U5050 ( .A1(n3676), .A2(n5099), .ZN(n5098) );
  OR2_X1 U5051 ( .A1(n5099), .A2(n3676), .ZN(n5096) );
  OR2_X1 U5052 ( .A1(n5100), .A2(n5101), .ZN(n4932) );
  INV_X1 U5053 ( .A(n5102), .ZN(n5101) );
  OR2_X1 U5054 ( .A1(n5103), .A2(n5104), .ZN(n5102) );
  AND2_X1 U5055 ( .A1(n5104), .A2(n5103), .ZN(n5100) );
  AND2_X1 U5056 ( .A1(n5105), .A2(n5106), .ZN(n5103) );
  INV_X1 U5057 ( .A(n5107), .ZN(n5106) );
  AND2_X1 U5058 ( .A1(n5108), .A2(n5109), .ZN(n5107) );
  OR2_X1 U5059 ( .A1(n5109), .A2(n5108), .ZN(n5105) );
  INV_X1 U5060 ( .A(n5110), .ZN(n5108) );
  OR2_X1 U5061 ( .A1(n5111), .A2(n5112), .ZN(n4942) );
  INV_X1 U5062 ( .A(n5113), .ZN(n5112) );
  OR2_X1 U5063 ( .A1(n5114), .A2(n5115), .ZN(n5113) );
  AND2_X1 U5064 ( .A1(n5115), .A2(n5114), .ZN(n5111) );
  AND2_X1 U5065 ( .A1(n5116), .A2(n5117), .ZN(n5114) );
  INV_X1 U5066 ( .A(n5118), .ZN(n5117) );
  AND2_X1 U5067 ( .A1(n5119), .A2(n5120), .ZN(n5118) );
  OR2_X1 U5068 ( .A1(n5120), .A2(n5119), .ZN(n5116) );
  OR2_X1 U5069 ( .A1(n5121), .A2(n5122), .ZN(n4952) );
  INV_X1 U5070 ( .A(n5123), .ZN(n5122) );
  OR2_X1 U5071 ( .A1(n5124), .A2(n5125), .ZN(n5123) );
  AND2_X1 U5072 ( .A1(n5125), .A2(n5124), .ZN(n5121) );
  AND2_X1 U5073 ( .A1(n5126), .A2(n5127), .ZN(n5124) );
  INV_X1 U5074 ( .A(n5128), .ZN(n5127) );
  AND2_X1 U5075 ( .A1(n5129), .A2(n5130), .ZN(n5128) );
  OR2_X1 U5076 ( .A1(n5130), .A2(n5129), .ZN(n5126) );
  OR2_X1 U5077 ( .A1(n5131), .A2(n5132), .ZN(n4962) );
  INV_X1 U5078 ( .A(n5133), .ZN(n5132) );
  OR2_X1 U5079 ( .A1(n5134), .A2(n5135), .ZN(n5133) );
  AND2_X1 U5080 ( .A1(n5135), .A2(n5134), .ZN(n5131) );
  AND2_X1 U5081 ( .A1(n5136), .A2(n5137), .ZN(n5134) );
  INV_X1 U5082 ( .A(n5138), .ZN(n5137) );
  AND2_X1 U5083 ( .A1(n5139), .A2(n5140), .ZN(n5138) );
  OR2_X1 U5084 ( .A1(n5140), .A2(n5139), .ZN(n5136) );
  OR2_X1 U5085 ( .A1(n5141), .A2(n5142), .ZN(n4972) );
  INV_X1 U5086 ( .A(n5143), .ZN(n5142) );
  OR2_X1 U5087 ( .A1(n5144), .A2(n5145), .ZN(n5143) );
  AND2_X1 U5088 ( .A1(n5145), .A2(n5144), .ZN(n5141) );
  AND2_X1 U5089 ( .A1(n5146), .A2(n5147), .ZN(n5144) );
  INV_X1 U5090 ( .A(n5148), .ZN(n5147) );
  AND2_X1 U5091 ( .A1(n5149), .A2(n5150), .ZN(n5148) );
  OR2_X1 U5092 ( .A1(n5150), .A2(n5149), .ZN(n5146) );
  OR2_X1 U5093 ( .A1(n5151), .A2(n5152), .ZN(n4982) );
  INV_X1 U5094 ( .A(n5153), .ZN(n5152) );
  OR2_X1 U5095 ( .A1(n5154), .A2(n5155), .ZN(n5153) );
  AND2_X1 U5096 ( .A1(n5155), .A2(n5154), .ZN(n5151) );
  AND2_X1 U5097 ( .A1(n5156), .A2(n5157), .ZN(n5154) );
  INV_X1 U5098 ( .A(n5158), .ZN(n5157) );
  AND2_X1 U5099 ( .A1(n5159), .A2(n5160), .ZN(n5158) );
  OR2_X1 U5100 ( .A1(n5160), .A2(n5159), .ZN(n5156) );
  OR2_X1 U5101 ( .A1(n5161), .A2(n5162), .ZN(n4992) );
  INV_X1 U5102 ( .A(n5163), .ZN(n5162) );
  OR2_X1 U5103 ( .A1(n5164), .A2(n5165), .ZN(n5163) );
  AND2_X1 U5104 ( .A1(n5165), .A2(n5164), .ZN(n5161) );
  AND2_X1 U5105 ( .A1(n5166), .A2(n5167), .ZN(n5164) );
  INV_X1 U5106 ( .A(n5168), .ZN(n5167) );
  AND2_X1 U5107 ( .A1(n5169), .A2(n5170), .ZN(n5168) );
  OR2_X1 U5108 ( .A1(n5170), .A2(n5169), .ZN(n5166) );
  OR2_X1 U5109 ( .A1(n5171), .A2(n5172), .ZN(n5002) );
  INV_X1 U5110 ( .A(n5173), .ZN(n5172) );
  OR2_X1 U5111 ( .A1(n5174), .A2(n5175), .ZN(n5173) );
  AND2_X1 U5112 ( .A1(n5175), .A2(n5174), .ZN(n5171) );
  AND2_X1 U5113 ( .A1(n5176), .A2(n5177), .ZN(n5174) );
  INV_X1 U5114 ( .A(n5178), .ZN(n5177) );
  AND2_X1 U5115 ( .A1(n5179), .A2(n5180), .ZN(n5178) );
  OR2_X1 U5116 ( .A1(n5180), .A2(n5179), .ZN(n5176) );
  OR2_X1 U5117 ( .A1(n5181), .A2(n5182), .ZN(n4642) );
  INV_X1 U5118 ( .A(n5183), .ZN(n5182) );
  OR2_X1 U5119 ( .A1(n5184), .A2(n5185), .ZN(n5183) );
  AND2_X1 U5120 ( .A1(n5185), .A2(n5184), .ZN(n5181) );
  AND2_X1 U5121 ( .A1(n5186), .A2(n5187), .ZN(n5184) );
  INV_X1 U5122 ( .A(n5188), .ZN(n5187) );
  AND2_X1 U5123 ( .A1(n5189), .A2(n5190), .ZN(n5188) );
  OR2_X1 U5124 ( .A1(n5190), .A2(n5189), .ZN(n5186) );
  AND2_X1 U5125 ( .A1(n5191), .A2(n5192), .ZN(n4616) );
  INV_X1 U5126 ( .A(n5193), .ZN(n5192) );
  AND2_X1 U5127 ( .A1(n5194), .A2(n5195), .ZN(n5193) );
  OR2_X1 U5128 ( .A1(n5195), .A2(n5194), .ZN(n5191) );
  OR2_X1 U5129 ( .A1(n5196), .A2(n5197), .ZN(n5194) );
  AND2_X1 U5130 ( .A1(n5198), .A2(n5199), .ZN(n5197) );
  INV_X1 U5131 ( .A(n5200), .ZN(n5196) );
  OR2_X1 U5132 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  AND2_X1 U5133 ( .A1(n5201), .A2(n5202), .ZN(n5010) );
  INV_X1 U5134 ( .A(n5203), .ZN(n5202) );
  AND2_X1 U5135 ( .A1(n5204), .A2(n5205), .ZN(n5203) );
  OR2_X1 U5136 ( .A1(n5205), .A2(n5204), .ZN(n5201) );
  OR2_X1 U5137 ( .A1(n5206), .A2(n5207), .ZN(n5204) );
  INV_X1 U5138 ( .A(n5208), .ZN(n5207) );
  OR2_X1 U5139 ( .A1(n5209), .A2(n5210), .ZN(n5208) );
  AND2_X1 U5140 ( .A1(n5210), .A2(n5209), .ZN(n5206) );
  INV_X1 U5141 ( .A(n5211), .ZN(n5210) );
  INV_X1 U5142 ( .A(n4017), .ZN(n4020) );
  OR2_X1 U5143 ( .A1(n5212), .A2(n4390), .ZN(n4017) );
  INV_X1 U5144 ( .A(n4023), .ZN(n4390) );
  OR2_X1 U5145 ( .A1(n5213), .A2(n5214), .ZN(n4023) );
  AND2_X1 U5146 ( .A1(n5213), .A2(n5214), .ZN(n5212) );
  OR2_X1 U5147 ( .A1(n5215), .A2(n5216), .ZN(n5214) );
  AND2_X1 U5148 ( .A1(n5209), .A2(n5211), .ZN(n5216) );
  AND2_X1 U5149 ( .A1(n5205), .A2(n5217), .ZN(n5215) );
  OR2_X1 U5150 ( .A1(n5211), .A2(n5209), .ZN(n5217) );
  OR2_X1 U5151 ( .A1(n3938), .A2(n3678), .ZN(n5209) );
  OR2_X1 U5152 ( .A1(n5218), .A2(n5219), .ZN(n5211) );
  AND2_X1 U5153 ( .A1(n5220), .A2(n5199), .ZN(n5219) );
  AND2_X1 U5154 ( .A1(n5195), .A2(n5221), .ZN(n5218) );
  OR2_X1 U5155 ( .A1(n5199), .A2(n5220), .ZN(n5221) );
  INV_X1 U5156 ( .A(n5198), .ZN(n5220) );
  AND2_X1 U5157 ( .A1(a_1_), .A2(b_11_), .ZN(n5198) );
  OR2_X1 U5158 ( .A1(n5222), .A2(n5223), .ZN(n5199) );
  AND2_X1 U5159 ( .A1(n5224), .A2(n5190), .ZN(n5223) );
  AND2_X1 U5160 ( .A1(n5185), .A2(n5225), .ZN(n5222) );
  OR2_X1 U5161 ( .A1(n5190), .A2(n5224), .ZN(n5225) );
  INV_X1 U5162 ( .A(n5189), .ZN(n5224) );
  AND2_X1 U5163 ( .A1(a_2_), .A2(b_11_), .ZN(n5189) );
  OR2_X1 U5164 ( .A1(n5226), .A2(n5227), .ZN(n5190) );
  AND2_X1 U5165 ( .A1(n5228), .A2(n5180), .ZN(n5227) );
  AND2_X1 U5166 ( .A1(n5175), .A2(n5229), .ZN(n5226) );
  OR2_X1 U5167 ( .A1(n5180), .A2(n5228), .ZN(n5229) );
  INV_X1 U5168 ( .A(n5179), .ZN(n5228) );
  AND2_X1 U5169 ( .A1(a_3_), .A2(b_11_), .ZN(n5179) );
  OR2_X1 U5170 ( .A1(n5230), .A2(n5231), .ZN(n5180) );
  AND2_X1 U5171 ( .A1(n5232), .A2(n5170), .ZN(n5231) );
  AND2_X1 U5172 ( .A1(n5165), .A2(n5233), .ZN(n5230) );
  OR2_X1 U5173 ( .A1(n5170), .A2(n5232), .ZN(n5233) );
  INV_X1 U5174 ( .A(n5169), .ZN(n5232) );
  AND2_X1 U5175 ( .A1(a_4_), .A2(b_11_), .ZN(n5169) );
  OR2_X1 U5176 ( .A1(n5234), .A2(n5235), .ZN(n5170) );
  AND2_X1 U5177 ( .A1(n5236), .A2(n5160), .ZN(n5235) );
  AND2_X1 U5178 ( .A1(n5155), .A2(n5237), .ZN(n5234) );
  OR2_X1 U5179 ( .A1(n5160), .A2(n5236), .ZN(n5237) );
  INV_X1 U5180 ( .A(n5159), .ZN(n5236) );
  AND2_X1 U5181 ( .A1(a_5_), .A2(b_11_), .ZN(n5159) );
  OR2_X1 U5182 ( .A1(n5238), .A2(n5239), .ZN(n5160) );
  AND2_X1 U5183 ( .A1(n5240), .A2(n5150), .ZN(n5239) );
  AND2_X1 U5184 ( .A1(n5145), .A2(n5241), .ZN(n5238) );
  OR2_X1 U5185 ( .A1(n5150), .A2(n5240), .ZN(n5241) );
  INV_X1 U5186 ( .A(n5149), .ZN(n5240) );
  AND2_X1 U5187 ( .A1(a_6_), .A2(b_11_), .ZN(n5149) );
  OR2_X1 U5188 ( .A1(n5242), .A2(n5243), .ZN(n5150) );
  AND2_X1 U5189 ( .A1(n5244), .A2(n5140), .ZN(n5243) );
  AND2_X1 U5190 ( .A1(n5135), .A2(n5245), .ZN(n5242) );
  OR2_X1 U5191 ( .A1(n5140), .A2(n5244), .ZN(n5245) );
  INV_X1 U5192 ( .A(n5139), .ZN(n5244) );
  AND2_X1 U5193 ( .A1(a_7_), .A2(b_11_), .ZN(n5139) );
  OR2_X1 U5194 ( .A1(n5246), .A2(n5247), .ZN(n5140) );
  AND2_X1 U5195 ( .A1(n5248), .A2(n5130), .ZN(n5247) );
  AND2_X1 U5196 ( .A1(n5125), .A2(n5249), .ZN(n5246) );
  OR2_X1 U5197 ( .A1(n5130), .A2(n5248), .ZN(n5249) );
  INV_X1 U5198 ( .A(n5129), .ZN(n5248) );
  AND2_X1 U5199 ( .A1(a_8_), .A2(b_11_), .ZN(n5129) );
  OR2_X1 U5200 ( .A1(n5250), .A2(n5251), .ZN(n5130) );
  AND2_X1 U5201 ( .A1(n5252), .A2(n5120), .ZN(n5251) );
  AND2_X1 U5202 ( .A1(n5115), .A2(n5253), .ZN(n5250) );
  OR2_X1 U5203 ( .A1(n5120), .A2(n5252), .ZN(n5253) );
  INV_X1 U5204 ( .A(n5119), .ZN(n5252) );
  AND2_X1 U5205 ( .A1(a_9_), .A2(b_11_), .ZN(n5119) );
  OR2_X1 U5206 ( .A1(n5254), .A2(n5255), .ZN(n5120) );
  AND2_X1 U5207 ( .A1(n5110), .A2(n5109), .ZN(n5255) );
  AND2_X1 U5208 ( .A1(n5104), .A2(n5256), .ZN(n5254) );
  OR2_X1 U5209 ( .A1(n5109), .A2(n5110), .ZN(n5256) );
  OR2_X1 U5210 ( .A1(n3964), .A2(n3678), .ZN(n5110) );
  OR2_X1 U5211 ( .A1(n5257), .A2(n5258), .ZN(n5109) );
  AND2_X1 U5212 ( .A1(n3969), .A2(n5099), .ZN(n5258) );
  AND2_X1 U5213 ( .A1(n5095), .A2(n5259), .ZN(n5257) );
  OR2_X1 U5214 ( .A1(n5099), .A2(n3969), .ZN(n5259) );
  INV_X1 U5215 ( .A(n3676), .ZN(n3969) );
  AND2_X1 U5216 ( .A1(a_11_), .A2(b_11_), .ZN(n3676) );
  OR2_X1 U5217 ( .A1(n5260), .A2(n5261), .ZN(n5099) );
  AND2_X1 U5218 ( .A1(n5262), .A2(n5090), .ZN(n5261) );
  AND2_X1 U5219 ( .A1(n5085), .A2(n5263), .ZN(n5260) );
  OR2_X1 U5220 ( .A1(n5090), .A2(n5262), .ZN(n5263) );
  INV_X1 U5221 ( .A(n5089), .ZN(n5262) );
  AND2_X1 U5222 ( .A1(a_12_), .A2(b_11_), .ZN(n5089) );
  OR2_X1 U5223 ( .A1(n5264), .A2(n5265), .ZN(n5090) );
  AND2_X1 U5224 ( .A1(n5073), .A2(n5078), .ZN(n5265) );
  AND2_X1 U5225 ( .A1(n5077), .A2(n5266), .ZN(n5264) );
  OR2_X1 U5226 ( .A1(n5078), .A2(n5073), .ZN(n5266) );
  OR2_X1 U5227 ( .A1(n3631), .A2(n3678), .ZN(n5073) );
  INV_X1 U5228 ( .A(b_11_), .ZN(n3678) );
  INV_X1 U5229 ( .A(n5079), .ZN(n5078) );
  AND3_X1 U5230 ( .A1(n3975), .A2(b_10_), .A3(b_11_), .ZN(n5079) );
  INV_X1 U5231 ( .A(n5080), .ZN(n5077) );
  OR2_X1 U5232 ( .A1(n5267), .A2(n5268), .ZN(n5080) );
  AND2_X1 U5233 ( .A1(b_9_), .A2(n5269), .ZN(n5268) );
  OR2_X1 U5234 ( .A1(n5270), .A2(n3595), .ZN(n5269) );
  AND2_X1 U5235 ( .A1(a_15_), .A2(n3965), .ZN(n5270) );
  AND2_X1 U5236 ( .A1(b_10_), .A2(n5271), .ZN(n5267) );
  OR2_X1 U5237 ( .A1(n5272), .A2(n3592), .ZN(n5271) );
  AND2_X1 U5238 ( .A1(a_14_), .A2(n3724), .ZN(n5272) );
  OR2_X1 U5239 ( .A1(n5273), .A2(n5274), .ZN(n5085) );
  AND2_X1 U5240 ( .A1(n5275), .A2(n5276), .ZN(n5274) );
  INV_X1 U5241 ( .A(n5277), .ZN(n5273) );
  OR2_X1 U5242 ( .A1(n5275), .A2(n5276), .ZN(n5277) );
  OR2_X1 U5243 ( .A1(n5278), .A2(n5279), .ZN(n5275) );
  AND2_X1 U5244 ( .A1(n5280), .A2(n5281), .ZN(n5279) );
  AND2_X1 U5245 ( .A1(n5282), .A2(n5283), .ZN(n5278) );
  OR2_X1 U5246 ( .A1(n5284), .A2(n5285), .ZN(n5095) );
  INV_X1 U5247 ( .A(n5286), .ZN(n5285) );
  OR2_X1 U5248 ( .A1(n5287), .A2(n5288), .ZN(n5286) );
  AND2_X1 U5249 ( .A1(n5288), .A2(n5287), .ZN(n5284) );
  AND2_X1 U5250 ( .A1(n5289), .A2(n5290), .ZN(n5287) );
  INV_X1 U5251 ( .A(n5291), .ZN(n5290) );
  AND2_X1 U5252 ( .A1(n5292), .A2(n5293), .ZN(n5291) );
  OR2_X1 U5253 ( .A1(n5293), .A2(n5292), .ZN(n5289) );
  OR2_X1 U5254 ( .A1(n5294), .A2(n5295), .ZN(n5104) );
  INV_X1 U5255 ( .A(n5296), .ZN(n5295) );
  OR2_X1 U5256 ( .A1(n5297), .A2(n5298), .ZN(n5296) );
  AND2_X1 U5257 ( .A1(n5298), .A2(n5297), .ZN(n5294) );
  AND2_X1 U5258 ( .A1(n5299), .A2(n5300), .ZN(n5297) );
  INV_X1 U5259 ( .A(n5301), .ZN(n5300) );
  AND2_X1 U5260 ( .A1(n5302), .A2(n5303), .ZN(n5301) );
  OR2_X1 U5261 ( .A1(n5303), .A2(n5302), .ZN(n5299) );
  OR2_X1 U5262 ( .A1(n5304), .A2(n5305), .ZN(n5115) );
  INV_X1 U5263 ( .A(n5306), .ZN(n5305) );
  OR2_X1 U5264 ( .A1(n5307), .A2(n5308), .ZN(n5306) );
  AND2_X1 U5265 ( .A1(n5308), .A2(n5307), .ZN(n5304) );
  AND2_X1 U5266 ( .A1(n5309), .A2(n5310), .ZN(n5307) );
  OR2_X1 U5267 ( .A1(n5311), .A2(n3704), .ZN(n5310) );
  INV_X1 U5268 ( .A(n5312), .ZN(n5309) );
  AND2_X1 U5269 ( .A1(n3704), .A2(n5311), .ZN(n5312) );
  INV_X1 U5270 ( .A(n3966), .ZN(n3704) );
  OR2_X1 U5271 ( .A1(n5313), .A2(n5314), .ZN(n5125) );
  INV_X1 U5272 ( .A(n5315), .ZN(n5314) );
  OR2_X1 U5273 ( .A1(n5316), .A2(n5317), .ZN(n5315) );
  AND2_X1 U5274 ( .A1(n5317), .A2(n5316), .ZN(n5313) );
  AND2_X1 U5275 ( .A1(n5318), .A2(n5319), .ZN(n5316) );
  INV_X1 U5276 ( .A(n5320), .ZN(n5319) );
  AND2_X1 U5277 ( .A1(n5321), .A2(n5322), .ZN(n5320) );
  OR2_X1 U5278 ( .A1(n5322), .A2(n5321), .ZN(n5318) );
  OR2_X1 U5279 ( .A1(n5323), .A2(n5324), .ZN(n5135) );
  INV_X1 U5280 ( .A(n5325), .ZN(n5324) );
  OR2_X1 U5281 ( .A1(n5326), .A2(n5327), .ZN(n5325) );
  AND2_X1 U5282 ( .A1(n5327), .A2(n5326), .ZN(n5323) );
  AND2_X1 U5283 ( .A1(n5328), .A2(n5329), .ZN(n5326) );
  INV_X1 U5284 ( .A(n5330), .ZN(n5329) );
  AND2_X1 U5285 ( .A1(n5331), .A2(n5332), .ZN(n5330) );
  OR2_X1 U5286 ( .A1(n5332), .A2(n5331), .ZN(n5328) );
  OR2_X1 U5287 ( .A1(n5333), .A2(n5334), .ZN(n5145) );
  INV_X1 U5288 ( .A(n5335), .ZN(n5334) );
  OR2_X1 U5289 ( .A1(n5336), .A2(n5337), .ZN(n5335) );
  AND2_X1 U5290 ( .A1(n5337), .A2(n5336), .ZN(n5333) );
  AND2_X1 U5291 ( .A1(n5338), .A2(n5339), .ZN(n5336) );
  INV_X1 U5292 ( .A(n5340), .ZN(n5339) );
  AND2_X1 U5293 ( .A1(n5341), .A2(n5342), .ZN(n5340) );
  OR2_X1 U5294 ( .A1(n5342), .A2(n5341), .ZN(n5338) );
  OR2_X1 U5295 ( .A1(n5343), .A2(n5344), .ZN(n5155) );
  INV_X1 U5296 ( .A(n5345), .ZN(n5344) );
  OR2_X1 U5297 ( .A1(n5346), .A2(n5347), .ZN(n5345) );
  AND2_X1 U5298 ( .A1(n5347), .A2(n5346), .ZN(n5343) );
  AND2_X1 U5299 ( .A1(n5348), .A2(n5349), .ZN(n5346) );
  INV_X1 U5300 ( .A(n5350), .ZN(n5349) );
  AND2_X1 U5301 ( .A1(n5351), .A2(n5352), .ZN(n5350) );
  OR2_X1 U5302 ( .A1(n5352), .A2(n5351), .ZN(n5348) );
  OR2_X1 U5303 ( .A1(n5353), .A2(n5354), .ZN(n5165) );
  INV_X1 U5304 ( .A(n5355), .ZN(n5354) );
  OR2_X1 U5305 ( .A1(n5356), .A2(n5357), .ZN(n5355) );
  AND2_X1 U5306 ( .A1(n5357), .A2(n5356), .ZN(n5353) );
  AND2_X1 U5307 ( .A1(n5358), .A2(n5359), .ZN(n5356) );
  INV_X1 U5308 ( .A(n5360), .ZN(n5359) );
  AND2_X1 U5309 ( .A1(n5361), .A2(n5362), .ZN(n5360) );
  OR2_X1 U5310 ( .A1(n5362), .A2(n5361), .ZN(n5358) );
  OR2_X1 U5311 ( .A1(n5363), .A2(n5364), .ZN(n5175) );
  INV_X1 U5312 ( .A(n5365), .ZN(n5364) );
  OR2_X1 U5313 ( .A1(n5366), .A2(n5367), .ZN(n5365) );
  AND2_X1 U5314 ( .A1(n5367), .A2(n5366), .ZN(n5363) );
  AND2_X1 U5315 ( .A1(n5368), .A2(n5369), .ZN(n5366) );
  INV_X1 U5316 ( .A(n5370), .ZN(n5369) );
  AND2_X1 U5317 ( .A1(n5371), .A2(n5372), .ZN(n5370) );
  OR2_X1 U5318 ( .A1(n5372), .A2(n5371), .ZN(n5368) );
  OR2_X1 U5319 ( .A1(n5373), .A2(n5374), .ZN(n5185) );
  INV_X1 U5320 ( .A(n5375), .ZN(n5374) );
  OR2_X1 U5321 ( .A1(n5376), .A2(n5377), .ZN(n5375) );
  AND2_X1 U5322 ( .A1(n5377), .A2(n5376), .ZN(n5373) );
  AND2_X1 U5323 ( .A1(n5378), .A2(n5379), .ZN(n5376) );
  INV_X1 U5324 ( .A(n5380), .ZN(n5379) );
  AND2_X1 U5325 ( .A1(n5381), .A2(n5382), .ZN(n5380) );
  OR2_X1 U5326 ( .A1(n5382), .A2(n5381), .ZN(n5378) );
  AND2_X1 U5327 ( .A1(n5383), .A2(n5384), .ZN(n5195) );
  INV_X1 U5328 ( .A(n5385), .ZN(n5384) );
  AND2_X1 U5329 ( .A1(n5386), .A2(n5387), .ZN(n5385) );
  OR2_X1 U5330 ( .A1(n5387), .A2(n5386), .ZN(n5383) );
  OR2_X1 U5331 ( .A1(n5388), .A2(n5389), .ZN(n5386) );
  AND2_X1 U5332 ( .A1(n5390), .A2(n5391), .ZN(n5389) );
  INV_X1 U5333 ( .A(n5392), .ZN(n5388) );
  OR2_X1 U5334 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  AND2_X1 U5335 ( .A1(n5393), .A2(n5394), .ZN(n5205) );
  INV_X1 U5336 ( .A(n5395), .ZN(n5394) );
  AND2_X1 U5337 ( .A1(n5396), .A2(n5397), .ZN(n5395) );
  OR2_X1 U5338 ( .A1(n5397), .A2(n5396), .ZN(n5393) );
  OR2_X1 U5339 ( .A1(n5398), .A2(n5399), .ZN(n5396) );
  AND2_X1 U5340 ( .A1(n5400), .A2(n5401), .ZN(n5399) );
  INV_X1 U5341 ( .A(n5402), .ZN(n5398) );
  OR2_X1 U5342 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  AND2_X1 U5343 ( .A1(n5403), .A2(n5404), .ZN(n5213) );
  INV_X1 U5344 ( .A(n5405), .ZN(n5404) );
  AND2_X1 U5345 ( .A1(n5406), .A2(n5407), .ZN(n5405) );
  OR2_X1 U5346 ( .A1(n5407), .A2(n5406), .ZN(n5403) );
  OR2_X1 U5347 ( .A1(n5408), .A2(n5409), .ZN(n5406) );
  INV_X1 U5348 ( .A(n5410), .ZN(n5409) );
  OR2_X1 U5349 ( .A1(n5411), .A2(n5412), .ZN(n5410) );
  AND2_X1 U5350 ( .A1(n5412), .A2(n5411), .ZN(n5408) );
  INV_X1 U5351 ( .A(n5413), .ZN(n5412) );
  AND2_X1 U5352 ( .A1(n5414), .A2(n3496), .ZN(n4030) );
  OR2_X1 U5353 ( .A1(n5415), .A2(n5416), .ZN(n3496) );
  INV_X1 U5354 ( .A(n5417), .ZN(n5414) );
  AND2_X1 U5355 ( .A1(n5415), .A2(n5416), .ZN(n5417) );
  OR2_X1 U5356 ( .A1(n5418), .A2(n5419), .ZN(n5416) );
  AND2_X1 U5357 ( .A1(n5411), .A2(n5413), .ZN(n5419) );
  AND2_X1 U5358 ( .A1(n5407), .A2(n5420), .ZN(n5418) );
  OR2_X1 U5359 ( .A1(n5411), .A2(n5413), .ZN(n5420) );
  OR2_X1 U5360 ( .A1(n5421), .A2(n5422), .ZN(n5413) );
  AND2_X1 U5361 ( .A1(n5423), .A2(n5401), .ZN(n5422) );
  AND2_X1 U5362 ( .A1(n5397), .A2(n5424), .ZN(n5421) );
  OR2_X1 U5363 ( .A1(n5423), .A2(n5401), .ZN(n5424) );
  OR2_X1 U5364 ( .A1(n5425), .A2(n5426), .ZN(n5401) );
  AND2_X1 U5365 ( .A1(n5427), .A2(n5391), .ZN(n5426) );
  AND2_X1 U5366 ( .A1(n5387), .A2(n5428), .ZN(n5425) );
  OR2_X1 U5367 ( .A1(n5427), .A2(n5391), .ZN(n5428) );
  OR2_X1 U5368 ( .A1(n5429), .A2(n5430), .ZN(n5391) );
  AND2_X1 U5369 ( .A1(n5377), .A2(n5431), .ZN(n5430) );
  AND2_X1 U5370 ( .A1(n5432), .A2(n5382), .ZN(n5429) );
  OR2_X1 U5371 ( .A1(n5433), .A2(n5434), .ZN(n5382) );
  AND2_X1 U5372 ( .A1(n5435), .A2(n5372), .ZN(n5434) );
  AND2_X1 U5373 ( .A1(n5367), .A2(n5436), .ZN(n5433) );
  OR2_X1 U5374 ( .A1(n5435), .A2(n5372), .ZN(n5436) );
  OR2_X1 U5375 ( .A1(n5437), .A2(n5438), .ZN(n5372) );
  AND2_X1 U5376 ( .A1(n5357), .A2(n5439), .ZN(n5438) );
  AND2_X1 U5377 ( .A1(n5440), .A2(n5362), .ZN(n5437) );
  OR2_X1 U5378 ( .A1(n5441), .A2(n5442), .ZN(n5362) );
  AND2_X1 U5379 ( .A1(n5347), .A2(n5443), .ZN(n5442) );
  AND2_X1 U5380 ( .A1(n5444), .A2(n5352), .ZN(n5441) );
  OR2_X1 U5381 ( .A1(n5445), .A2(n5446), .ZN(n5352) );
  AND2_X1 U5382 ( .A1(n5337), .A2(n5447), .ZN(n5446) );
  AND2_X1 U5383 ( .A1(n5448), .A2(n5342), .ZN(n5445) );
  OR2_X1 U5384 ( .A1(n5449), .A2(n5450), .ZN(n5342) );
  AND2_X1 U5385 ( .A1(n5327), .A2(n5451), .ZN(n5450) );
  AND2_X1 U5386 ( .A1(n5452), .A2(n5332), .ZN(n5449) );
  OR2_X1 U5387 ( .A1(n5453), .A2(n5454), .ZN(n5332) );
  AND2_X1 U5388 ( .A1(n5317), .A2(n5455), .ZN(n5454) );
  AND2_X1 U5389 ( .A1(n5456), .A2(n5322), .ZN(n5453) );
  OR2_X1 U5390 ( .A1(n5457), .A2(n5458), .ZN(n5322) );
  AND2_X1 U5391 ( .A1(n5308), .A2(n3966), .ZN(n5458) );
  AND2_X1 U5392 ( .A1(n5459), .A2(n5311), .ZN(n5457) );
  OR2_X1 U5393 ( .A1(n5460), .A2(n5461), .ZN(n5311) );
  AND2_X1 U5394 ( .A1(n5298), .A2(n5462), .ZN(n5461) );
  AND2_X1 U5395 ( .A1(n5463), .A2(n5303), .ZN(n5460) );
  OR2_X1 U5396 ( .A1(n5464), .A2(n5465), .ZN(n5303) );
  AND2_X1 U5397 ( .A1(n5288), .A2(n5466), .ZN(n5465) );
  AND2_X1 U5398 ( .A1(n5467), .A2(n5293), .ZN(n5464) );
  OR2_X1 U5399 ( .A1(n5468), .A2(n5469), .ZN(n5293) );
  AND2_X1 U5400 ( .A1(n5276), .A2(n5281), .ZN(n5469) );
  AND2_X1 U5401 ( .A1(n5280), .A2(n5470), .ZN(n5468) );
  OR2_X1 U5402 ( .A1(n5276), .A2(n5281), .ZN(n5470) );
  INV_X1 U5403 ( .A(n5282), .ZN(n5281) );
  AND3_X1 U5404 ( .A1(b_9_), .A2(n3975), .A3(b_10_), .ZN(n5282) );
  OR2_X1 U5405 ( .A1(n3965), .A2(n3631), .ZN(n5276) );
  INV_X1 U5406 ( .A(n5283), .ZN(n5280) );
  OR2_X1 U5407 ( .A1(n5471), .A2(n5472), .ZN(n5283) );
  AND2_X1 U5408 ( .A1(b_9_), .A2(n5473), .ZN(n5472) );
  OR2_X1 U5409 ( .A1(n5474), .A2(n3592), .ZN(n5473) );
  AND2_X1 U5410 ( .A1(a_14_), .A2(n5475), .ZN(n5474) );
  AND2_X1 U5411 ( .A1(b_8_), .A2(n5476), .ZN(n5471) );
  OR2_X1 U5412 ( .A1(n5477), .A2(n3595), .ZN(n5476) );
  AND2_X1 U5413 ( .A1(a_15_), .A2(n3724), .ZN(n5477) );
  OR2_X1 U5414 ( .A1(n5288), .A2(n5466), .ZN(n5467) );
  INV_X1 U5415 ( .A(n5292), .ZN(n5466) );
  AND2_X1 U5416 ( .A1(b_10_), .A2(a_12_), .ZN(n5292) );
  OR2_X1 U5417 ( .A1(n5478), .A2(n5479), .ZN(n5288) );
  AND2_X1 U5418 ( .A1(n5480), .A2(n5481), .ZN(n5479) );
  INV_X1 U5419 ( .A(n5482), .ZN(n5478) );
  OR2_X1 U5420 ( .A1(n5480), .A2(n5481), .ZN(n5482) );
  OR2_X1 U5421 ( .A1(n5483), .A2(n5484), .ZN(n5480) );
  AND2_X1 U5422 ( .A1(n5485), .A2(n5486), .ZN(n5484) );
  AND2_X1 U5423 ( .A1(n5487), .A2(n5488), .ZN(n5483) );
  OR2_X1 U5424 ( .A1(n5298), .A2(n5462), .ZN(n5463) );
  INV_X1 U5425 ( .A(n5302), .ZN(n5462) );
  AND2_X1 U5426 ( .A1(b_10_), .A2(a_11_), .ZN(n5302) );
  OR2_X1 U5427 ( .A1(n5489), .A2(n5490), .ZN(n5298) );
  INV_X1 U5428 ( .A(n5491), .ZN(n5490) );
  OR2_X1 U5429 ( .A1(n5492), .A2(n5493), .ZN(n5491) );
  AND2_X1 U5430 ( .A1(n5493), .A2(n5492), .ZN(n5489) );
  AND2_X1 U5431 ( .A1(n5494), .A2(n5495), .ZN(n5492) );
  INV_X1 U5432 ( .A(n5496), .ZN(n5495) );
  AND2_X1 U5433 ( .A1(n5497), .A2(n5498), .ZN(n5496) );
  OR2_X1 U5434 ( .A1(n5498), .A2(n5497), .ZN(n5494) );
  OR2_X1 U5435 ( .A1(n5308), .A2(n3966), .ZN(n5459) );
  OR2_X1 U5436 ( .A1(n3965), .A2(n3964), .ZN(n3966) );
  OR2_X1 U5437 ( .A1(n5499), .A2(n5500), .ZN(n5308) );
  INV_X1 U5438 ( .A(n5501), .ZN(n5500) );
  OR2_X1 U5439 ( .A1(n5502), .A2(n5503), .ZN(n5501) );
  AND2_X1 U5440 ( .A1(n5503), .A2(n5502), .ZN(n5499) );
  AND2_X1 U5441 ( .A1(n5504), .A2(n5505), .ZN(n5502) );
  INV_X1 U5442 ( .A(n5506), .ZN(n5505) );
  AND2_X1 U5443 ( .A1(n5507), .A2(n5508), .ZN(n5506) );
  OR2_X1 U5444 ( .A1(n5508), .A2(n5507), .ZN(n5504) );
  OR2_X1 U5445 ( .A1(n5317), .A2(n5455), .ZN(n5456) );
  INV_X1 U5446 ( .A(n5321), .ZN(n5455) );
  AND2_X1 U5447 ( .A1(b_10_), .A2(a_9_), .ZN(n5321) );
  OR2_X1 U5448 ( .A1(n5509), .A2(n5510), .ZN(n5317) );
  INV_X1 U5449 ( .A(n5511), .ZN(n5510) );
  OR2_X1 U5450 ( .A1(n5512), .A2(n5513), .ZN(n5511) );
  AND2_X1 U5451 ( .A1(n5513), .A2(n5512), .ZN(n5509) );
  AND2_X1 U5452 ( .A1(n5514), .A2(n5515), .ZN(n5512) );
  INV_X1 U5453 ( .A(n5516), .ZN(n5515) );
  AND2_X1 U5454 ( .A1(n5517), .A2(n5518), .ZN(n5516) );
  OR2_X1 U5455 ( .A1(n5518), .A2(n5517), .ZN(n5514) );
  INV_X1 U5456 ( .A(n5519), .ZN(n5517) );
  OR2_X1 U5457 ( .A1(n5327), .A2(n5451), .ZN(n5452) );
  INV_X1 U5458 ( .A(n5331), .ZN(n5451) );
  AND2_X1 U5459 ( .A1(b_10_), .A2(a_8_), .ZN(n5331) );
  OR2_X1 U5460 ( .A1(n5520), .A2(n5521), .ZN(n5327) );
  INV_X1 U5461 ( .A(n5522), .ZN(n5521) );
  OR2_X1 U5462 ( .A1(n5523), .A2(n5524), .ZN(n5522) );
  AND2_X1 U5463 ( .A1(n5524), .A2(n5523), .ZN(n5520) );
  AND2_X1 U5464 ( .A1(n5525), .A2(n5526), .ZN(n5523) );
  INV_X1 U5465 ( .A(n5527), .ZN(n5526) );
  AND2_X1 U5466 ( .A1(n3722), .A2(n5528), .ZN(n5527) );
  OR2_X1 U5467 ( .A1(n5528), .A2(n3722), .ZN(n5525) );
  OR2_X1 U5468 ( .A1(n5337), .A2(n5447), .ZN(n5448) );
  INV_X1 U5469 ( .A(n5341), .ZN(n5447) );
  AND2_X1 U5470 ( .A1(b_10_), .A2(a_7_), .ZN(n5341) );
  OR2_X1 U5471 ( .A1(n5529), .A2(n5530), .ZN(n5337) );
  INV_X1 U5472 ( .A(n5531), .ZN(n5530) );
  OR2_X1 U5473 ( .A1(n5532), .A2(n5533), .ZN(n5531) );
  AND2_X1 U5474 ( .A1(n5533), .A2(n5532), .ZN(n5529) );
  AND2_X1 U5475 ( .A1(n5534), .A2(n5535), .ZN(n5532) );
  INV_X1 U5476 ( .A(n5536), .ZN(n5535) );
  AND2_X1 U5477 ( .A1(n5537), .A2(n5538), .ZN(n5536) );
  OR2_X1 U5478 ( .A1(n5538), .A2(n5537), .ZN(n5534) );
  OR2_X1 U5479 ( .A1(n5347), .A2(n5443), .ZN(n5444) );
  INV_X1 U5480 ( .A(n5351), .ZN(n5443) );
  AND2_X1 U5481 ( .A1(b_10_), .A2(a_6_), .ZN(n5351) );
  OR2_X1 U5482 ( .A1(n5539), .A2(n5540), .ZN(n5347) );
  INV_X1 U5483 ( .A(n5541), .ZN(n5540) );
  OR2_X1 U5484 ( .A1(n5542), .A2(n5543), .ZN(n5541) );
  AND2_X1 U5485 ( .A1(n5543), .A2(n5542), .ZN(n5539) );
  AND2_X1 U5486 ( .A1(n5544), .A2(n5545), .ZN(n5542) );
  INV_X1 U5487 ( .A(n5546), .ZN(n5545) );
  AND2_X1 U5488 ( .A1(n5547), .A2(n5548), .ZN(n5546) );
  OR2_X1 U5489 ( .A1(n5548), .A2(n5547), .ZN(n5544) );
  OR2_X1 U5490 ( .A1(n5357), .A2(n5439), .ZN(n5440) );
  INV_X1 U5491 ( .A(n5361), .ZN(n5439) );
  AND2_X1 U5492 ( .A1(b_10_), .A2(a_5_), .ZN(n5361) );
  OR2_X1 U5493 ( .A1(n5549), .A2(n5550), .ZN(n5357) );
  INV_X1 U5494 ( .A(n5551), .ZN(n5550) );
  OR2_X1 U5495 ( .A1(n5552), .A2(n5553), .ZN(n5551) );
  AND2_X1 U5496 ( .A1(n5553), .A2(n5552), .ZN(n5549) );
  AND2_X1 U5497 ( .A1(n5554), .A2(n5555), .ZN(n5552) );
  INV_X1 U5498 ( .A(n5556), .ZN(n5555) );
  AND2_X1 U5499 ( .A1(n5557), .A2(n5558), .ZN(n5556) );
  OR2_X1 U5500 ( .A1(n5558), .A2(n5557), .ZN(n5554) );
  INV_X1 U5501 ( .A(n5371), .ZN(n5435) );
  AND2_X1 U5502 ( .A1(b_10_), .A2(a_4_), .ZN(n5371) );
  OR2_X1 U5503 ( .A1(n5559), .A2(n5560), .ZN(n5367) );
  INV_X1 U5504 ( .A(n5561), .ZN(n5560) );
  OR2_X1 U5505 ( .A1(n5562), .A2(n5563), .ZN(n5561) );
  AND2_X1 U5506 ( .A1(n5563), .A2(n5562), .ZN(n5559) );
  AND2_X1 U5507 ( .A1(n5564), .A2(n5565), .ZN(n5562) );
  INV_X1 U5508 ( .A(n5566), .ZN(n5565) );
  AND2_X1 U5509 ( .A1(n5567), .A2(n5568), .ZN(n5566) );
  OR2_X1 U5510 ( .A1(n5568), .A2(n5567), .ZN(n5564) );
  OR2_X1 U5511 ( .A1(n5377), .A2(n5431), .ZN(n5432) );
  INV_X1 U5512 ( .A(n5381), .ZN(n5431) );
  AND2_X1 U5513 ( .A1(b_10_), .A2(a_3_), .ZN(n5381) );
  OR2_X1 U5514 ( .A1(n5569), .A2(n5570), .ZN(n5377) );
  INV_X1 U5515 ( .A(n5571), .ZN(n5570) );
  OR2_X1 U5516 ( .A1(n5572), .A2(n5573), .ZN(n5571) );
  AND2_X1 U5517 ( .A1(n5573), .A2(n5572), .ZN(n5569) );
  AND2_X1 U5518 ( .A1(n5574), .A2(n5575), .ZN(n5572) );
  INV_X1 U5519 ( .A(n5576), .ZN(n5575) );
  AND2_X1 U5520 ( .A1(n5577), .A2(n5578), .ZN(n5576) );
  OR2_X1 U5521 ( .A1(n5578), .A2(n5577), .ZN(n5574) );
  INV_X1 U5522 ( .A(n5390), .ZN(n5427) );
  AND2_X1 U5523 ( .A1(b_10_), .A2(a_2_), .ZN(n5390) );
  AND2_X1 U5524 ( .A1(n5579), .A2(n5580), .ZN(n5387) );
  INV_X1 U5525 ( .A(n5581), .ZN(n5580) );
  AND2_X1 U5526 ( .A1(n5582), .A2(n5583), .ZN(n5581) );
  OR2_X1 U5527 ( .A1(n5583), .A2(n5582), .ZN(n5579) );
  OR2_X1 U5528 ( .A1(n5584), .A2(n5585), .ZN(n5582) );
  AND2_X1 U5529 ( .A1(n5586), .A2(n5587), .ZN(n5585) );
  INV_X1 U5530 ( .A(n5588), .ZN(n5584) );
  OR2_X1 U5531 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  INV_X1 U5532 ( .A(n5400), .ZN(n5423) );
  AND2_X1 U5533 ( .A1(b_10_), .A2(a_1_), .ZN(n5400) );
  AND2_X1 U5534 ( .A1(n5589), .A2(n5590), .ZN(n5397) );
  INV_X1 U5535 ( .A(n5591), .ZN(n5590) );
  AND2_X1 U5536 ( .A1(n5592), .A2(n5593), .ZN(n5591) );
  OR2_X1 U5537 ( .A1(n5593), .A2(n5592), .ZN(n5589) );
  OR2_X1 U5538 ( .A1(n5594), .A2(n5595), .ZN(n5592) );
  AND2_X1 U5539 ( .A1(n5596), .A2(n5597), .ZN(n5595) );
  INV_X1 U5540 ( .A(n5598), .ZN(n5594) );
  OR2_X1 U5541 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  OR2_X1 U5542 ( .A1(n3965), .A2(n3938), .ZN(n5411) );
  INV_X1 U5543 ( .A(b_10_), .ZN(n3965) );
  AND2_X1 U5544 ( .A1(n5599), .A2(n5600), .ZN(n5407) );
  INV_X1 U5545 ( .A(n5601), .ZN(n5600) );
  AND2_X1 U5546 ( .A1(n5602), .A2(n5603), .ZN(n5601) );
  OR2_X1 U5547 ( .A1(n5603), .A2(n5602), .ZN(n5599) );
  OR2_X1 U5548 ( .A1(n5604), .A2(n5605), .ZN(n5602) );
  AND2_X1 U5549 ( .A1(n5606), .A2(n5607), .ZN(n5605) );
  INV_X1 U5550 ( .A(n5608), .ZN(n5604) );
  OR2_X1 U5551 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  AND2_X1 U5552 ( .A1(n5609), .A2(n5610), .ZN(n5415) );
  INV_X1 U5553 ( .A(n5611), .ZN(n5610) );
  AND2_X1 U5554 ( .A1(n5612), .A2(n5613), .ZN(n5611) );
  OR2_X1 U5555 ( .A1(n5613), .A2(n5612), .ZN(n5609) );
  OR2_X1 U5556 ( .A1(n5614), .A2(n5615), .ZN(n5612) );
  INV_X1 U5557 ( .A(n5616), .ZN(n5615) );
  OR2_X1 U5558 ( .A1(n5617), .A2(n5618), .ZN(n5616) );
  AND2_X1 U5559 ( .A1(n5618), .A2(n5617), .ZN(n5614) );
  INV_X1 U5560 ( .A(n5619), .ZN(n5618) );
  INV_X1 U5561 ( .A(n3509), .ZN(n3510) );
  OR2_X1 U5562 ( .A1(n5620), .A2(n4387), .ZN(n3509) );
  OR2_X1 U5563 ( .A1(n5621), .A2(n5622), .ZN(n4387) );
  AND2_X1 U5564 ( .A1(n5617), .A2(n5619), .ZN(n5622) );
  AND2_X1 U5565 ( .A1(n5613), .A2(n5623), .ZN(n5621) );
  OR2_X1 U5566 ( .A1(n5619), .A2(n5617), .ZN(n5623) );
  OR2_X1 U5567 ( .A1(n3724), .A2(n3938), .ZN(n5617) );
  OR2_X1 U5568 ( .A1(n5624), .A2(n5625), .ZN(n5619) );
  AND2_X1 U5569 ( .A1(n5626), .A2(n5607), .ZN(n5625) );
  AND2_X1 U5570 ( .A1(n5603), .A2(n5627), .ZN(n5624) );
  OR2_X1 U5571 ( .A1(n5607), .A2(n5626), .ZN(n5627) );
  INV_X1 U5572 ( .A(n5606), .ZN(n5626) );
  AND2_X1 U5573 ( .A1(b_9_), .A2(a_1_), .ZN(n5606) );
  OR2_X1 U5574 ( .A1(n5628), .A2(n5629), .ZN(n5607) );
  AND2_X1 U5575 ( .A1(n5630), .A2(n5597), .ZN(n5629) );
  AND2_X1 U5576 ( .A1(n5593), .A2(n5631), .ZN(n5628) );
  OR2_X1 U5577 ( .A1(n5597), .A2(n5630), .ZN(n5631) );
  INV_X1 U5578 ( .A(n5596), .ZN(n5630) );
  AND2_X1 U5579 ( .A1(b_9_), .A2(a_2_), .ZN(n5596) );
  OR2_X1 U5580 ( .A1(n5632), .A2(n5633), .ZN(n5597) );
  AND2_X1 U5581 ( .A1(n5634), .A2(n5587), .ZN(n5633) );
  AND2_X1 U5582 ( .A1(n5583), .A2(n5635), .ZN(n5632) );
  OR2_X1 U5583 ( .A1(n5587), .A2(n5634), .ZN(n5635) );
  INV_X1 U5584 ( .A(n5586), .ZN(n5634) );
  AND2_X1 U5585 ( .A1(b_9_), .A2(a_3_), .ZN(n5586) );
  OR2_X1 U5586 ( .A1(n5636), .A2(n5637), .ZN(n5587) );
  AND2_X1 U5587 ( .A1(n5573), .A2(n5638), .ZN(n5637) );
  AND2_X1 U5588 ( .A1(n5639), .A2(n5578), .ZN(n5636) );
  OR2_X1 U5589 ( .A1(n5640), .A2(n5641), .ZN(n5578) );
  AND2_X1 U5590 ( .A1(n5642), .A2(n5568), .ZN(n5641) );
  AND2_X1 U5591 ( .A1(n5563), .A2(n5643), .ZN(n5640) );
  OR2_X1 U5592 ( .A1(n5568), .A2(n5642), .ZN(n5643) );
  INV_X1 U5593 ( .A(n5567), .ZN(n5642) );
  AND2_X1 U5594 ( .A1(b_9_), .A2(a_5_), .ZN(n5567) );
  OR2_X1 U5595 ( .A1(n5644), .A2(n5645), .ZN(n5568) );
  AND2_X1 U5596 ( .A1(n5553), .A2(n5646), .ZN(n5645) );
  AND2_X1 U5597 ( .A1(n5647), .A2(n5558), .ZN(n5644) );
  OR2_X1 U5598 ( .A1(n5648), .A2(n5649), .ZN(n5558) );
  AND2_X1 U5599 ( .A1(n5543), .A2(n5650), .ZN(n5649) );
  AND2_X1 U5600 ( .A1(n5651), .A2(n5548), .ZN(n5648) );
  OR2_X1 U5601 ( .A1(n5652), .A2(n5653), .ZN(n5548) );
  AND2_X1 U5602 ( .A1(n5533), .A2(n5654), .ZN(n5653) );
  AND2_X1 U5603 ( .A1(n5655), .A2(n5538), .ZN(n5652) );
  OR2_X1 U5604 ( .A1(n5656), .A2(n5657), .ZN(n5538) );
  AND2_X1 U5605 ( .A1(n5524), .A2(n3962), .ZN(n5657) );
  AND2_X1 U5606 ( .A1(n5658), .A2(n5528), .ZN(n5656) );
  OR2_X1 U5607 ( .A1(n5659), .A2(n5660), .ZN(n5528) );
  AND2_X1 U5608 ( .A1(n5513), .A2(n5519), .ZN(n5660) );
  AND2_X1 U5609 ( .A1(n5661), .A2(n5518), .ZN(n5659) );
  OR2_X1 U5610 ( .A1(n5662), .A2(n5663), .ZN(n5518) );
  AND2_X1 U5611 ( .A1(n5503), .A2(n5664), .ZN(n5663) );
  AND2_X1 U5612 ( .A1(n5665), .A2(n5508), .ZN(n5662) );
  OR2_X1 U5613 ( .A1(n5666), .A2(n5667), .ZN(n5508) );
  AND2_X1 U5614 ( .A1(n5493), .A2(n5668), .ZN(n5667) );
  AND2_X1 U5615 ( .A1(n5669), .A2(n5498), .ZN(n5666) );
  OR2_X1 U5616 ( .A1(n5670), .A2(n5671), .ZN(n5498) );
  AND2_X1 U5617 ( .A1(n5481), .A2(n5486), .ZN(n5671) );
  AND2_X1 U5618 ( .A1(n5485), .A2(n5672), .ZN(n5670) );
  OR2_X1 U5619 ( .A1(n5486), .A2(n5481), .ZN(n5672) );
  OR2_X1 U5620 ( .A1(n3724), .A2(n3631), .ZN(n5481) );
  INV_X1 U5621 ( .A(n5487), .ZN(n5486) );
  AND3_X1 U5622 ( .A1(b_8_), .A2(b_9_), .A3(n3975), .ZN(n5487) );
  INV_X1 U5623 ( .A(n5488), .ZN(n5485) );
  OR2_X1 U5624 ( .A1(n5673), .A2(n5674), .ZN(n5488) );
  AND2_X1 U5625 ( .A1(b_8_), .A2(n5675), .ZN(n5674) );
  OR2_X1 U5626 ( .A1(n5676), .A2(n3592), .ZN(n5675) );
  AND2_X1 U5627 ( .A1(a_14_), .A2(n3768), .ZN(n5676) );
  AND2_X1 U5628 ( .A1(b_7_), .A2(n5677), .ZN(n5673) );
  OR2_X1 U5629 ( .A1(n5678), .A2(n3595), .ZN(n5677) );
  AND2_X1 U5630 ( .A1(a_15_), .A2(n5475), .ZN(n5678) );
  OR2_X1 U5631 ( .A1(n5668), .A2(n5493), .ZN(n5669) );
  OR2_X1 U5632 ( .A1(n5679), .A2(n5680), .ZN(n5493) );
  AND2_X1 U5633 ( .A1(n5681), .A2(n5682), .ZN(n5680) );
  INV_X1 U5634 ( .A(n5683), .ZN(n5679) );
  OR2_X1 U5635 ( .A1(n5681), .A2(n5682), .ZN(n5683) );
  OR2_X1 U5636 ( .A1(n5684), .A2(n5685), .ZN(n5681) );
  AND2_X1 U5637 ( .A1(n5686), .A2(n5687), .ZN(n5685) );
  AND2_X1 U5638 ( .A1(n5688), .A2(n5689), .ZN(n5684) );
  INV_X1 U5639 ( .A(n5497), .ZN(n5668) );
  AND2_X1 U5640 ( .A1(b_9_), .A2(a_12_), .ZN(n5497) );
  OR2_X1 U5641 ( .A1(n5664), .A2(n5503), .ZN(n5665) );
  OR2_X1 U5642 ( .A1(n5690), .A2(n5691), .ZN(n5503) );
  INV_X1 U5643 ( .A(n5692), .ZN(n5691) );
  OR2_X1 U5644 ( .A1(n5693), .A2(n5694), .ZN(n5692) );
  AND2_X1 U5645 ( .A1(n5694), .A2(n5693), .ZN(n5690) );
  AND2_X1 U5646 ( .A1(n5695), .A2(n5696), .ZN(n5693) );
  INV_X1 U5647 ( .A(n5697), .ZN(n5696) );
  AND2_X1 U5648 ( .A1(n5698), .A2(n5699), .ZN(n5697) );
  OR2_X1 U5649 ( .A1(n5699), .A2(n5698), .ZN(n5695) );
  INV_X1 U5650 ( .A(n5507), .ZN(n5664) );
  AND2_X1 U5651 ( .A1(b_9_), .A2(a_11_), .ZN(n5507) );
  OR2_X1 U5652 ( .A1(n5519), .A2(n5513), .ZN(n5661) );
  OR2_X1 U5653 ( .A1(n5700), .A2(n5701), .ZN(n5513) );
  INV_X1 U5654 ( .A(n5702), .ZN(n5701) );
  OR2_X1 U5655 ( .A1(n5703), .A2(n5704), .ZN(n5702) );
  AND2_X1 U5656 ( .A1(n5704), .A2(n5703), .ZN(n5700) );
  AND2_X1 U5657 ( .A1(n5705), .A2(n5706), .ZN(n5703) );
  INV_X1 U5658 ( .A(n5707), .ZN(n5706) );
  AND2_X1 U5659 ( .A1(n5708), .A2(n5709), .ZN(n5707) );
  OR2_X1 U5660 ( .A1(n5709), .A2(n5708), .ZN(n5705) );
  OR2_X1 U5661 ( .A1(n3724), .A2(n3964), .ZN(n5519) );
  INV_X1 U5662 ( .A(b_9_), .ZN(n3724) );
  OR2_X1 U5663 ( .A1(n3962), .A2(n5524), .ZN(n5658) );
  OR2_X1 U5664 ( .A1(n5710), .A2(n5711), .ZN(n5524) );
  INV_X1 U5665 ( .A(n5712), .ZN(n5711) );
  OR2_X1 U5666 ( .A1(n5713), .A2(n5714), .ZN(n5712) );
  AND2_X1 U5667 ( .A1(n5714), .A2(n5713), .ZN(n5710) );
  AND2_X1 U5668 ( .A1(n5715), .A2(n5716), .ZN(n5713) );
  INV_X1 U5669 ( .A(n5717), .ZN(n5716) );
  AND2_X1 U5670 ( .A1(n5718), .A2(n5719), .ZN(n5717) );
  OR2_X1 U5671 ( .A1(n5719), .A2(n5718), .ZN(n5715) );
  INV_X1 U5672 ( .A(n5720), .ZN(n5718) );
  INV_X1 U5673 ( .A(n3722), .ZN(n3962) );
  AND2_X1 U5674 ( .A1(b_9_), .A2(a_9_), .ZN(n3722) );
  OR2_X1 U5675 ( .A1(n5654), .A2(n5533), .ZN(n5655) );
  OR2_X1 U5676 ( .A1(n5721), .A2(n5722), .ZN(n5533) );
  INV_X1 U5677 ( .A(n5723), .ZN(n5722) );
  OR2_X1 U5678 ( .A1(n5724), .A2(n5725), .ZN(n5723) );
  AND2_X1 U5679 ( .A1(n5725), .A2(n5724), .ZN(n5721) );
  AND2_X1 U5680 ( .A1(n5726), .A2(n5727), .ZN(n5724) );
  INV_X1 U5681 ( .A(n5728), .ZN(n5727) );
  AND2_X1 U5682 ( .A1(n5729), .A2(n5730), .ZN(n5728) );
  OR2_X1 U5683 ( .A1(n5730), .A2(n5729), .ZN(n5726) );
  INV_X1 U5684 ( .A(n5537), .ZN(n5654) );
  AND2_X1 U5685 ( .A1(b_9_), .A2(a_8_), .ZN(n5537) );
  OR2_X1 U5686 ( .A1(n5650), .A2(n5543), .ZN(n5651) );
  OR2_X1 U5687 ( .A1(n5731), .A2(n5732), .ZN(n5543) );
  INV_X1 U5688 ( .A(n5733), .ZN(n5732) );
  OR2_X1 U5689 ( .A1(n5734), .A2(n5735), .ZN(n5733) );
  AND2_X1 U5690 ( .A1(n5735), .A2(n5734), .ZN(n5731) );
  AND2_X1 U5691 ( .A1(n5736), .A2(n5737), .ZN(n5734) );
  INV_X1 U5692 ( .A(n5738), .ZN(n5737) );
  AND2_X1 U5693 ( .A1(n5739), .A2(n3748), .ZN(n5738) );
  OR2_X1 U5694 ( .A1(n3748), .A2(n5739), .ZN(n5736) );
  INV_X1 U5695 ( .A(n5740), .ZN(n5739) );
  INV_X1 U5696 ( .A(n5547), .ZN(n5650) );
  AND2_X1 U5697 ( .A1(b_9_), .A2(a_7_), .ZN(n5547) );
  OR2_X1 U5698 ( .A1(n5646), .A2(n5553), .ZN(n5647) );
  OR2_X1 U5699 ( .A1(n5741), .A2(n5742), .ZN(n5553) );
  INV_X1 U5700 ( .A(n5743), .ZN(n5742) );
  OR2_X1 U5701 ( .A1(n5744), .A2(n5745), .ZN(n5743) );
  AND2_X1 U5702 ( .A1(n5745), .A2(n5744), .ZN(n5741) );
  AND2_X1 U5703 ( .A1(n5746), .A2(n5747), .ZN(n5744) );
  INV_X1 U5704 ( .A(n5748), .ZN(n5747) );
  AND2_X1 U5705 ( .A1(n5749), .A2(n5750), .ZN(n5748) );
  OR2_X1 U5706 ( .A1(n5750), .A2(n5749), .ZN(n5746) );
  INV_X1 U5707 ( .A(n5557), .ZN(n5646) );
  AND2_X1 U5708 ( .A1(b_9_), .A2(a_6_), .ZN(n5557) );
  OR2_X1 U5709 ( .A1(n5751), .A2(n5752), .ZN(n5563) );
  INV_X1 U5710 ( .A(n5753), .ZN(n5752) );
  OR2_X1 U5711 ( .A1(n5754), .A2(n5755), .ZN(n5753) );
  AND2_X1 U5712 ( .A1(n5755), .A2(n5754), .ZN(n5751) );
  AND2_X1 U5713 ( .A1(n5756), .A2(n5757), .ZN(n5754) );
  INV_X1 U5714 ( .A(n5758), .ZN(n5757) );
  AND2_X1 U5715 ( .A1(n5759), .A2(n5760), .ZN(n5758) );
  OR2_X1 U5716 ( .A1(n5760), .A2(n5759), .ZN(n5756) );
  OR2_X1 U5717 ( .A1(n5638), .A2(n5573), .ZN(n5639) );
  OR2_X1 U5718 ( .A1(n5761), .A2(n5762), .ZN(n5573) );
  INV_X1 U5719 ( .A(n5763), .ZN(n5762) );
  OR2_X1 U5720 ( .A1(n5764), .A2(n5765), .ZN(n5763) );
  AND2_X1 U5721 ( .A1(n5765), .A2(n5764), .ZN(n5761) );
  AND2_X1 U5722 ( .A1(n5766), .A2(n5767), .ZN(n5764) );
  INV_X1 U5723 ( .A(n5768), .ZN(n5767) );
  AND2_X1 U5724 ( .A1(n5769), .A2(n5770), .ZN(n5768) );
  OR2_X1 U5725 ( .A1(n5770), .A2(n5769), .ZN(n5766) );
  INV_X1 U5726 ( .A(n5577), .ZN(n5638) );
  AND2_X1 U5727 ( .A1(b_9_), .A2(a_4_), .ZN(n5577) );
  AND2_X1 U5728 ( .A1(n5771), .A2(n5772), .ZN(n5583) );
  INV_X1 U5729 ( .A(n5773), .ZN(n5772) );
  AND2_X1 U5730 ( .A1(n5774), .A2(n5775), .ZN(n5773) );
  OR2_X1 U5731 ( .A1(n5775), .A2(n5774), .ZN(n5771) );
  OR2_X1 U5732 ( .A1(n5776), .A2(n5777), .ZN(n5774) );
  AND2_X1 U5733 ( .A1(n5778), .A2(n5779), .ZN(n5777) );
  INV_X1 U5734 ( .A(n5780), .ZN(n5776) );
  OR2_X1 U5735 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  AND2_X1 U5736 ( .A1(n5781), .A2(n5782), .ZN(n5593) );
  INV_X1 U5737 ( .A(n5783), .ZN(n5782) );
  AND2_X1 U5738 ( .A1(n5784), .A2(n5785), .ZN(n5783) );
  OR2_X1 U5739 ( .A1(n5785), .A2(n5784), .ZN(n5781) );
  OR2_X1 U5740 ( .A1(n5786), .A2(n5787), .ZN(n5784) );
  AND2_X1 U5741 ( .A1(n5788), .A2(n5789), .ZN(n5787) );
  INV_X1 U5742 ( .A(n5790), .ZN(n5786) );
  OR2_X1 U5743 ( .A1(n5789), .A2(n5788), .ZN(n5790) );
  AND2_X1 U5744 ( .A1(n5791), .A2(n5792), .ZN(n5603) );
  INV_X1 U5745 ( .A(n5793), .ZN(n5792) );
  AND2_X1 U5746 ( .A1(n5794), .A2(n5795), .ZN(n5793) );
  OR2_X1 U5747 ( .A1(n5795), .A2(n5794), .ZN(n5791) );
  OR2_X1 U5748 ( .A1(n5796), .A2(n5797), .ZN(n5794) );
  AND2_X1 U5749 ( .A1(n5798), .A2(n5799), .ZN(n5797) );
  INV_X1 U5750 ( .A(n5800), .ZN(n5796) );
  OR2_X1 U5751 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  AND2_X1 U5752 ( .A1(n5801), .A2(n5802), .ZN(n5613) );
  INV_X1 U5753 ( .A(n5803), .ZN(n5802) );
  AND2_X1 U5754 ( .A1(n5804), .A2(n5805), .ZN(n5803) );
  OR2_X1 U5755 ( .A1(n5805), .A2(n5804), .ZN(n5801) );
  OR2_X1 U5756 ( .A1(n5806), .A2(n5807), .ZN(n5804) );
  AND2_X1 U5757 ( .A1(n5808), .A2(n5809), .ZN(n5807) );
  INV_X1 U5758 ( .A(n5810), .ZN(n5806) );
  OR2_X1 U5759 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  AND2_X1 U5760 ( .A1(n4385), .A2(n4386), .ZN(n5620) );
  OR2_X1 U5761 ( .A1(n5811), .A2(n4302), .ZN(n4386) );
  INV_X1 U5762 ( .A(n5812), .ZN(n4302) );
  OR2_X1 U5763 ( .A1(n5812), .A2(n5813), .ZN(n4385) );
  INV_X1 U5764 ( .A(n5811), .ZN(n5813) );
  OR2_X1 U5765 ( .A1(n5814), .A2(n5815), .ZN(n5811) );
  AND2_X1 U5766 ( .A1(n5816), .A2(n4301), .ZN(n5815) );
  INV_X1 U5767 ( .A(n5817), .ZN(n5814) );
  OR2_X1 U5768 ( .A1(n4301), .A2(n5816), .ZN(n5817) );
  INV_X1 U5769 ( .A(n4300), .ZN(n5816) );
  OR2_X1 U5770 ( .A1(n5475), .A2(n3938), .ZN(n4300) );
  OR2_X1 U5771 ( .A1(n5818), .A2(n5819), .ZN(n4301) );
  AND2_X1 U5772 ( .A1(n5820), .A2(n5809), .ZN(n5819) );
  AND2_X1 U5773 ( .A1(n5805), .A2(n5821), .ZN(n5818) );
  OR2_X1 U5774 ( .A1(n5809), .A2(n5820), .ZN(n5821) );
  INV_X1 U5775 ( .A(n5808), .ZN(n5820) );
  AND2_X1 U5776 ( .A1(b_8_), .A2(a_1_), .ZN(n5808) );
  OR2_X1 U5777 ( .A1(n5822), .A2(n5823), .ZN(n5809) );
  AND2_X1 U5778 ( .A1(n5824), .A2(n5799), .ZN(n5823) );
  AND2_X1 U5779 ( .A1(n5795), .A2(n5825), .ZN(n5822) );
  OR2_X1 U5780 ( .A1(n5799), .A2(n5824), .ZN(n5825) );
  INV_X1 U5781 ( .A(n5798), .ZN(n5824) );
  AND2_X1 U5782 ( .A1(b_8_), .A2(a_2_), .ZN(n5798) );
  OR2_X1 U5783 ( .A1(n5826), .A2(n5827), .ZN(n5799) );
  AND2_X1 U5784 ( .A1(n5828), .A2(n5789), .ZN(n5827) );
  AND2_X1 U5785 ( .A1(n5785), .A2(n5829), .ZN(n5826) );
  OR2_X1 U5786 ( .A1(n5789), .A2(n5828), .ZN(n5829) );
  INV_X1 U5787 ( .A(n5788), .ZN(n5828) );
  AND2_X1 U5788 ( .A1(b_8_), .A2(a_3_), .ZN(n5788) );
  OR2_X1 U5789 ( .A1(n5830), .A2(n5831), .ZN(n5789) );
  AND2_X1 U5790 ( .A1(n5832), .A2(n5779), .ZN(n5831) );
  AND2_X1 U5791 ( .A1(n5775), .A2(n5833), .ZN(n5830) );
  OR2_X1 U5792 ( .A1(n5779), .A2(n5832), .ZN(n5833) );
  INV_X1 U5793 ( .A(n5778), .ZN(n5832) );
  AND2_X1 U5794 ( .A1(b_8_), .A2(a_4_), .ZN(n5778) );
  OR2_X1 U5795 ( .A1(n5834), .A2(n5835), .ZN(n5779) );
  AND2_X1 U5796 ( .A1(n5765), .A2(n5836), .ZN(n5835) );
  AND2_X1 U5797 ( .A1(n5837), .A2(n5770), .ZN(n5834) );
  OR2_X1 U5798 ( .A1(n5838), .A2(n5839), .ZN(n5770) );
  AND2_X1 U5799 ( .A1(n5840), .A2(n5760), .ZN(n5839) );
  AND2_X1 U5800 ( .A1(n5755), .A2(n5841), .ZN(n5838) );
  OR2_X1 U5801 ( .A1(n5760), .A2(n5840), .ZN(n5841) );
  INV_X1 U5802 ( .A(n5759), .ZN(n5840) );
  AND2_X1 U5803 ( .A1(b_8_), .A2(a_6_), .ZN(n5759) );
  OR2_X1 U5804 ( .A1(n5842), .A2(n5843), .ZN(n5760) );
  AND2_X1 U5805 ( .A1(n5745), .A2(n5844), .ZN(n5843) );
  AND2_X1 U5806 ( .A1(n5845), .A2(n5750), .ZN(n5842) );
  OR2_X1 U5807 ( .A1(n5846), .A2(n5847), .ZN(n5750) );
  AND2_X1 U5808 ( .A1(n5735), .A2(n3748), .ZN(n5847) );
  AND2_X1 U5809 ( .A1(n5848), .A2(n5740), .ZN(n5846) );
  OR2_X1 U5810 ( .A1(n5849), .A2(n5850), .ZN(n5740) );
  AND2_X1 U5811 ( .A1(n5725), .A2(n5851), .ZN(n5850) );
  AND2_X1 U5812 ( .A1(n5852), .A2(n5730), .ZN(n5849) );
  OR2_X1 U5813 ( .A1(n5853), .A2(n5854), .ZN(n5730) );
  AND2_X1 U5814 ( .A1(n5714), .A2(n5720), .ZN(n5854) );
  AND2_X1 U5815 ( .A1(n5855), .A2(n5719), .ZN(n5853) );
  OR2_X1 U5816 ( .A1(n5856), .A2(n5857), .ZN(n5719) );
  AND2_X1 U5817 ( .A1(n5704), .A2(n5858), .ZN(n5857) );
  AND2_X1 U5818 ( .A1(n5859), .A2(n5709), .ZN(n5856) );
  OR2_X1 U5819 ( .A1(n5860), .A2(n5861), .ZN(n5709) );
  AND2_X1 U5820 ( .A1(n5694), .A2(n5862), .ZN(n5861) );
  AND2_X1 U5821 ( .A1(n5863), .A2(n5699), .ZN(n5860) );
  OR2_X1 U5822 ( .A1(n5864), .A2(n5865), .ZN(n5699) );
  AND2_X1 U5823 ( .A1(n5682), .A2(n5687), .ZN(n5865) );
  AND2_X1 U5824 ( .A1(n5686), .A2(n5866), .ZN(n5864) );
  OR2_X1 U5825 ( .A1(n5687), .A2(n5682), .ZN(n5866) );
  OR2_X1 U5826 ( .A1(n5475), .A2(n3631), .ZN(n5682) );
  INV_X1 U5827 ( .A(n5688), .ZN(n5687) );
  AND3_X1 U5828 ( .A1(b_8_), .A2(n3975), .A3(b_7_), .ZN(n5688) );
  INV_X1 U5829 ( .A(n5689), .ZN(n5686) );
  OR2_X1 U5830 ( .A1(n5867), .A2(n5868), .ZN(n5689) );
  AND2_X1 U5831 ( .A1(b_7_), .A2(n5869), .ZN(n5868) );
  OR2_X1 U5832 ( .A1(n5870), .A2(n3592), .ZN(n5869) );
  AND2_X1 U5833 ( .A1(a_14_), .A2(n4235), .ZN(n5870) );
  AND2_X1 U5834 ( .A1(b_6_), .A2(n5871), .ZN(n5867) );
  OR2_X1 U5835 ( .A1(n5872), .A2(n3595), .ZN(n5871) );
  AND2_X1 U5836 ( .A1(a_15_), .A2(n3768), .ZN(n5872) );
  OR2_X1 U5837 ( .A1(n5862), .A2(n5694), .ZN(n5863) );
  OR2_X1 U5838 ( .A1(n5873), .A2(n5874), .ZN(n5694) );
  AND2_X1 U5839 ( .A1(n5875), .A2(n5876), .ZN(n5874) );
  INV_X1 U5840 ( .A(n5877), .ZN(n5873) );
  OR2_X1 U5841 ( .A1(n5875), .A2(n5876), .ZN(n5877) );
  OR2_X1 U5842 ( .A1(n5878), .A2(n5879), .ZN(n5875) );
  AND2_X1 U5843 ( .A1(n5880), .A2(n5881), .ZN(n5879) );
  AND2_X1 U5844 ( .A1(n5882), .A2(n5883), .ZN(n5878) );
  INV_X1 U5845 ( .A(n5698), .ZN(n5862) );
  AND2_X1 U5846 ( .A1(b_8_), .A2(a_12_), .ZN(n5698) );
  OR2_X1 U5847 ( .A1(n5858), .A2(n5704), .ZN(n5859) );
  OR2_X1 U5848 ( .A1(n5884), .A2(n5885), .ZN(n5704) );
  INV_X1 U5849 ( .A(n5886), .ZN(n5885) );
  OR2_X1 U5850 ( .A1(n5887), .A2(n5888), .ZN(n5886) );
  AND2_X1 U5851 ( .A1(n5888), .A2(n5887), .ZN(n5884) );
  AND2_X1 U5852 ( .A1(n5889), .A2(n5890), .ZN(n5887) );
  INV_X1 U5853 ( .A(n5891), .ZN(n5890) );
  AND2_X1 U5854 ( .A1(n5892), .A2(n5893), .ZN(n5891) );
  OR2_X1 U5855 ( .A1(n5893), .A2(n5892), .ZN(n5889) );
  INV_X1 U5856 ( .A(n5708), .ZN(n5858) );
  AND2_X1 U5857 ( .A1(b_8_), .A2(a_11_), .ZN(n5708) );
  OR2_X1 U5858 ( .A1(n5720), .A2(n5714), .ZN(n5855) );
  OR2_X1 U5859 ( .A1(n5894), .A2(n5895), .ZN(n5714) );
  INV_X1 U5860 ( .A(n5896), .ZN(n5895) );
  OR2_X1 U5861 ( .A1(n5897), .A2(n5898), .ZN(n5896) );
  AND2_X1 U5862 ( .A1(n5898), .A2(n5897), .ZN(n5894) );
  AND2_X1 U5863 ( .A1(n5899), .A2(n5900), .ZN(n5897) );
  INV_X1 U5864 ( .A(n5901), .ZN(n5900) );
  AND2_X1 U5865 ( .A1(n5902), .A2(n5903), .ZN(n5901) );
  OR2_X1 U5866 ( .A1(n5903), .A2(n5902), .ZN(n5899) );
  OR2_X1 U5867 ( .A1(n5475), .A2(n3964), .ZN(n5720) );
  OR2_X1 U5868 ( .A1(n5851), .A2(n5725), .ZN(n5852) );
  OR2_X1 U5869 ( .A1(n5904), .A2(n5905), .ZN(n5725) );
  INV_X1 U5870 ( .A(n5906), .ZN(n5905) );
  OR2_X1 U5871 ( .A1(n5907), .A2(n5908), .ZN(n5906) );
  AND2_X1 U5872 ( .A1(n5908), .A2(n5907), .ZN(n5904) );
  AND2_X1 U5873 ( .A1(n5909), .A2(n5910), .ZN(n5907) );
  INV_X1 U5874 ( .A(n5911), .ZN(n5910) );
  AND2_X1 U5875 ( .A1(n5912), .A2(n5913), .ZN(n5911) );
  OR2_X1 U5876 ( .A1(n5913), .A2(n5912), .ZN(n5909) );
  INV_X1 U5877 ( .A(n5914), .ZN(n5912) );
  INV_X1 U5878 ( .A(n5729), .ZN(n5851) );
  AND2_X1 U5879 ( .A1(b_8_), .A2(a_9_), .ZN(n5729) );
  OR2_X1 U5880 ( .A1(n3748), .A2(n5735), .ZN(n5848) );
  OR2_X1 U5881 ( .A1(n5915), .A2(n5916), .ZN(n5735) );
  INV_X1 U5882 ( .A(n5917), .ZN(n5916) );
  OR2_X1 U5883 ( .A1(n5918), .A2(n5919), .ZN(n5917) );
  AND2_X1 U5884 ( .A1(n5919), .A2(n5918), .ZN(n5915) );
  AND2_X1 U5885 ( .A1(n5920), .A2(n5921), .ZN(n5918) );
  INV_X1 U5886 ( .A(n5922), .ZN(n5921) );
  AND2_X1 U5887 ( .A1(n5923), .A2(n5924), .ZN(n5922) );
  OR2_X1 U5888 ( .A1(n5924), .A2(n5923), .ZN(n5920) );
  OR2_X1 U5889 ( .A1(n5475), .A2(n5925), .ZN(n3748) );
  INV_X1 U5890 ( .A(b_8_), .ZN(n5475) );
  OR2_X1 U5891 ( .A1(n5844), .A2(n5745), .ZN(n5845) );
  OR2_X1 U5892 ( .A1(n5926), .A2(n5927), .ZN(n5745) );
  INV_X1 U5893 ( .A(n5928), .ZN(n5927) );
  OR2_X1 U5894 ( .A1(n5929), .A2(n5930), .ZN(n5928) );
  AND2_X1 U5895 ( .A1(n5930), .A2(n5929), .ZN(n5926) );
  AND2_X1 U5896 ( .A1(n5931), .A2(n5932), .ZN(n5929) );
  INV_X1 U5897 ( .A(n5933), .ZN(n5932) );
  AND2_X1 U5898 ( .A1(n5934), .A2(n5935), .ZN(n5933) );
  OR2_X1 U5899 ( .A1(n5935), .A2(n5934), .ZN(n5931) );
  INV_X1 U5900 ( .A(n5749), .ZN(n5844) );
  AND2_X1 U5901 ( .A1(b_8_), .A2(a_7_), .ZN(n5749) );
  OR2_X1 U5902 ( .A1(n5936), .A2(n5937), .ZN(n5755) );
  INV_X1 U5903 ( .A(n5938), .ZN(n5937) );
  OR2_X1 U5904 ( .A1(n5939), .A2(n5940), .ZN(n5938) );
  AND2_X1 U5905 ( .A1(n5940), .A2(n5939), .ZN(n5936) );
  AND2_X1 U5906 ( .A1(n5941), .A2(n5942), .ZN(n5939) );
  INV_X1 U5907 ( .A(n5943), .ZN(n5942) );
  AND2_X1 U5908 ( .A1(n3766), .A2(n5944), .ZN(n5943) );
  OR2_X1 U5909 ( .A1(n5944), .A2(n3766), .ZN(n5941) );
  OR2_X1 U5910 ( .A1(n5836), .A2(n5765), .ZN(n5837) );
  OR2_X1 U5911 ( .A1(n5945), .A2(n5946), .ZN(n5765) );
  INV_X1 U5912 ( .A(n5947), .ZN(n5946) );
  OR2_X1 U5913 ( .A1(n5948), .A2(n5949), .ZN(n5947) );
  AND2_X1 U5914 ( .A1(n5949), .A2(n5948), .ZN(n5945) );
  AND2_X1 U5915 ( .A1(n5950), .A2(n5951), .ZN(n5948) );
  INV_X1 U5916 ( .A(n5952), .ZN(n5951) );
  AND2_X1 U5917 ( .A1(n5953), .A2(n5954), .ZN(n5952) );
  OR2_X1 U5918 ( .A1(n5954), .A2(n5953), .ZN(n5950) );
  INV_X1 U5919 ( .A(n5769), .ZN(n5836) );
  AND2_X1 U5920 ( .A1(b_8_), .A2(a_5_), .ZN(n5769) );
  AND2_X1 U5921 ( .A1(n5955), .A2(n5956), .ZN(n5775) );
  INV_X1 U5922 ( .A(n5957), .ZN(n5956) );
  AND2_X1 U5923 ( .A1(n5958), .A2(n5959), .ZN(n5957) );
  OR2_X1 U5924 ( .A1(n5959), .A2(n5958), .ZN(n5955) );
  OR2_X1 U5925 ( .A1(n5960), .A2(n5961), .ZN(n5958) );
  AND2_X1 U5926 ( .A1(n5962), .A2(n5963), .ZN(n5961) );
  INV_X1 U5927 ( .A(n5964), .ZN(n5960) );
  OR2_X1 U5928 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  AND2_X1 U5929 ( .A1(n5965), .A2(n5966), .ZN(n5785) );
  INV_X1 U5930 ( .A(n5967), .ZN(n5966) );
  AND2_X1 U5931 ( .A1(n5968), .A2(n5969), .ZN(n5967) );
  OR2_X1 U5932 ( .A1(n5969), .A2(n5968), .ZN(n5965) );
  OR2_X1 U5933 ( .A1(n5970), .A2(n5971), .ZN(n5968) );
  AND2_X1 U5934 ( .A1(n5972), .A2(n5973), .ZN(n5971) );
  INV_X1 U5935 ( .A(n5974), .ZN(n5970) );
  OR2_X1 U5936 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  AND2_X1 U5937 ( .A1(n5975), .A2(n5976), .ZN(n5795) );
  INV_X1 U5938 ( .A(n5977), .ZN(n5976) );
  AND2_X1 U5939 ( .A1(n5978), .A2(n5979), .ZN(n5977) );
  OR2_X1 U5940 ( .A1(n5979), .A2(n5978), .ZN(n5975) );
  OR2_X1 U5941 ( .A1(n5980), .A2(n5981), .ZN(n5978) );
  AND2_X1 U5942 ( .A1(n5982), .A2(n5983), .ZN(n5981) );
  INV_X1 U5943 ( .A(n5984), .ZN(n5980) );
  OR2_X1 U5944 ( .A1(n5983), .A2(n5982), .ZN(n5984) );
  AND2_X1 U5945 ( .A1(n5985), .A2(n5986), .ZN(n5805) );
  INV_X1 U5946 ( .A(n5987), .ZN(n5986) );
  AND2_X1 U5947 ( .A1(n5988), .A2(n5989), .ZN(n5987) );
  OR2_X1 U5948 ( .A1(n5989), .A2(n5988), .ZN(n5985) );
  OR2_X1 U5949 ( .A1(n5990), .A2(n5991), .ZN(n5988) );
  AND2_X1 U5950 ( .A1(n5992), .A2(n5993), .ZN(n5991) );
  INV_X1 U5951 ( .A(n5994), .ZN(n5990) );
  OR2_X1 U5952 ( .A1(n5993), .A2(n5992), .ZN(n5994) );
  OR2_X1 U5953 ( .A1(n5995), .A2(n5996), .ZN(n5812) );
  AND2_X1 U5954 ( .A1(n5997), .A2(n4316), .ZN(n5996) );
  INV_X1 U5955 ( .A(n5998), .ZN(n5995) );
  OR2_X1 U5956 ( .A1(n4316), .A2(n5997), .ZN(n5998) );
  OR2_X1 U5957 ( .A1(n5999), .A2(n6000), .ZN(n5997) );
  AND2_X1 U5958 ( .A1(n4318), .A2(n4315), .ZN(n6000) );
  INV_X1 U5959 ( .A(n6001), .ZN(n5999) );
  OR2_X1 U5960 ( .A1(n4315), .A2(n4318), .ZN(n6001) );
  AND2_X1 U5961 ( .A1(b_7_), .A2(a_1_), .ZN(n4318) );
  OR2_X1 U5962 ( .A1(n6002), .A2(n6003), .ZN(n4315) );
  AND2_X1 U5963 ( .A1(n6004), .A2(n5993), .ZN(n6003) );
  AND2_X1 U5964 ( .A1(n5989), .A2(n6005), .ZN(n6002) );
  OR2_X1 U5965 ( .A1(n5993), .A2(n6004), .ZN(n6005) );
  INV_X1 U5966 ( .A(n5992), .ZN(n6004) );
  AND2_X1 U5967 ( .A1(b_7_), .A2(a_2_), .ZN(n5992) );
  OR2_X1 U5968 ( .A1(n6006), .A2(n6007), .ZN(n5993) );
  AND2_X1 U5969 ( .A1(n6008), .A2(n5983), .ZN(n6007) );
  AND2_X1 U5970 ( .A1(n5979), .A2(n6009), .ZN(n6006) );
  OR2_X1 U5971 ( .A1(n5983), .A2(n6008), .ZN(n6009) );
  INV_X1 U5972 ( .A(n5982), .ZN(n6008) );
  AND2_X1 U5973 ( .A1(b_7_), .A2(a_3_), .ZN(n5982) );
  OR2_X1 U5974 ( .A1(n6010), .A2(n6011), .ZN(n5983) );
  AND2_X1 U5975 ( .A1(n6012), .A2(n5973), .ZN(n6011) );
  AND2_X1 U5976 ( .A1(n5969), .A2(n6013), .ZN(n6010) );
  OR2_X1 U5977 ( .A1(n5973), .A2(n6012), .ZN(n6013) );
  INV_X1 U5978 ( .A(n5972), .ZN(n6012) );
  AND2_X1 U5979 ( .A1(b_7_), .A2(a_4_), .ZN(n5972) );
  OR2_X1 U5980 ( .A1(n6014), .A2(n6015), .ZN(n5973) );
  AND2_X1 U5981 ( .A1(n6016), .A2(n5963), .ZN(n6015) );
  AND2_X1 U5982 ( .A1(n5959), .A2(n6017), .ZN(n6014) );
  OR2_X1 U5983 ( .A1(n5963), .A2(n6016), .ZN(n6017) );
  INV_X1 U5984 ( .A(n5962), .ZN(n6016) );
  AND2_X1 U5985 ( .A1(b_7_), .A2(a_5_), .ZN(n5962) );
  OR2_X1 U5986 ( .A1(n6018), .A2(n6019), .ZN(n5963) );
  AND2_X1 U5987 ( .A1(n5949), .A2(n6020), .ZN(n6019) );
  AND2_X1 U5988 ( .A1(n6021), .A2(n5954), .ZN(n6018) );
  OR2_X1 U5989 ( .A1(n6022), .A2(n6023), .ZN(n5954) );
  AND2_X1 U5990 ( .A1(n3957), .A2(n5944), .ZN(n6023) );
  AND2_X1 U5991 ( .A1(n5940), .A2(n6024), .ZN(n6022) );
  OR2_X1 U5992 ( .A1(n5944), .A2(n3957), .ZN(n6024) );
  INV_X1 U5993 ( .A(n3766), .ZN(n3957) );
  AND2_X1 U5994 ( .A1(b_7_), .A2(a_7_), .ZN(n3766) );
  OR2_X1 U5995 ( .A1(n6025), .A2(n6026), .ZN(n5944) );
  AND2_X1 U5996 ( .A1(n5930), .A2(n6027), .ZN(n6026) );
  AND2_X1 U5997 ( .A1(n6028), .A2(n5935), .ZN(n6025) );
  OR2_X1 U5998 ( .A1(n6029), .A2(n6030), .ZN(n5935) );
  AND2_X1 U5999 ( .A1(n5919), .A2(n6031), .ZN(n6030) );
  AND2_X1 U6000 ( .A1(n6032), .A2(n5924), .ZN(n6029) );
  OR2_X1 U6001 ( .A1(n6033), .A2(n6034), .ZN(n5924) );
  AND2_X1 U6002 ( .A1(n5908), .A2(n5914), .ZN(n6034) );
  AND2_X1 U6003 ( .A1(n6035), .A2(n5913), .ZN(n6033) );
  OR2_X1 U6004 ( .A1(n6036), .A2(n6037), .ZN(n5913) );
  AND2_X1 U6005 ( .A1(n5898), .A2(n6038), .ZN(n6037) );
  AND2_X1 U6006 ( .A1(n6039), .A2(n5903), .ZN(n6036) );
  OR2_X1 U6007 ( .A1(n6040), .A2(n6041), .ZN(n5903) );
  AND2_X1 U6008 ( .A1(n5888), .A2(n6042), .ZN(n6041) );
  AND2_X1 U6009 ( .A1(n6043), .A2(n5893), .ZN(n6040) );
  OR2_X1 U6010 ( .A1(n6044), .A2(n6045), .ZN(n5893) );
  AND2_X1 U6011 ( .A1(n5876), .A2(n5881), .ZN(n6045) );
  AND2_X1 U6012 ( .A1(n5880), .A2(n6046), .ZN(n6044) );
  OR2_X1 U6013 ( .A1(n5881), .A2(n5876), .ZN(n6046) );
  OR2_X1 U6014 ( .A1(n3631), .A2(n3768), .ZN(n5876) );
  INV_X1 U6015 ( .A(n5882), .ZN(n5881) );
  AND3_X1 U6016 ( .A1(n3975), .A2(b_7_), .A3(b_6_), .ZN(n5882) );
  INV_X1 U6017 ( .A(n5883), .ZN(n5880) );
  OR2_X1 U6018 ( .A1(n6047), .A2(n6048), .ZN(n5883) );
  AND2_X1 U6019 ( .A1(b_6_), .A2(n6049), .ZN(n6048) );
  OR2_X1 U6020 ( .A1(n6050), .A2(n3592), .ZN(n6049) );
  AND2_X1 U6021 ( .A1(a_14_), .A2(n3812), .ZN(n6050) );
  AND2_X1 U6022 ( .A1(b_5_), .A2(n6051), .ZN(n6047) );
  OR2_X1 U6023 ( .A1(n6052), .A2(n3595), .ZN(n6051) );
  AND2_X1 U6024 ( .A1(a_15_), .A2(n4235), .ZN(n6052) );
  OR2_X1 U6025 ( .A1(n6042), .A2(n5888), .ZN(n6043) );
  OR2_X1 U6026 ( .A1(n6053), .A2(n6054), .ZN(n5888) );
  AND2_X1 U6027 ( .A1(n6055), .A2(n6056), .ZN(n6054) );
  INV_X1 U6028 ( .A(n6057), .ZN(n6053) );
  OR2_X1 U6029 ( .A1(n6055), .A2(n6056), .ZN(n6057) );
  OR2_X1 U6030 ( .A1(n6058), .A2(n6059), .ZN(n6055) );
  AND2_X1 U6031 ( .A1(n6060), .A2(n6061), .ZN(n6059) );
  AND2_X1 U6032 ( .A1(n6062), .A2(n6063), .ZN(n6058) );
  INV_X1 U6033 ( .A(n5892), .ZN(n6042) );
  AND2_X1 U6034 ( .A1(a_12_), .A2(b_7_), .ZN(n5892) );
  OR2_X1 U6035 ( .A1(n6038), .A2(n5898), .ZN(n6039) );
  OR2_X1 U6036 ( .A1(n6064), .A2(n6065), .ZN(n5898) );
  INV_X1 U6037 ( .A(n6066), .ZN(n6065) );
  OR2_X1 U6038 ( .A1(n6067), .A2(n6068), .ZN(n6066) );
  AND2_X1 U6039 ( .A1(n6068), .A2(n6067), .ZN(n6064) );
  AND2_X1 U6040 ( .A1(n6069), .A2(n6070), .ZN(n6067) );
  INV_X1 U6041 ( .A(n6071), .ZN(n6070) );
  AND2_X1 U6042 ( .A1(n6072), .A2(n6073), .ZN(n6071) );
  OR2_X1 U6043 ( .A1(n6073), .A2(n6072), .ZN(n6069) );
  INV_X1 U6044 ( .A(n5902), .ZN(n6038) );
  AND2_X1 U6045 ( .A1(b_7_), .A2(a_11_), .ZN(n5902) );
  OR2_X1 U6046 ( .A1(n5914), .A2(n5908), .ZN(n6035) );
  OR2_X1 U6047 ( .A1(n6074), .A2(n6075), .ZN(n5908) );
  INV_X1 U6048 ( .A(n6076), .ZN(n6075) );
  OR2_X1 U6049 ( .A1(n6077), .A2(n6078), .ZN(n6076) );
  AND2_X1 U6050 ( .A1(n6078), .A2(n6077), .ZN(n6074) );
  AND2_X1 U6051 ( .A1(n6079), .A2(n6080), .ZN(n6077) );
  INV_X1 U6052 ( .A(n6081), .ZN(n6080) );
  AND2_X1 U6053 ( .A1(n6082), .A2(n6083), .ZN(n6081) );
  OR2_X1 U6054 ( .A1(n6083), .A2(n6082), .ZN(n6079) );
  OR2_X1 U6055 ( .A1(n3768), .A2(n3964), .ZN(n5914) );
  INV_X1 U6056 ( .A(b_7_), .ZN(n3768) );
  OR2_X1 U6057 ( .A1(n6031), .A2(n5919), .ZN(n6032) );
  OR2_X1 U6058 ( .A1(n6084), .A2(n6085), .ZN(n5919) );
  INV_X1 U6059 ( .A(n6086), .ZN(n6085) );
  OR2_X1 U6060 ( .A1(n6087), .A2(n6088), .ZN(n6086) );
  AND2_X1 U6061 ( .A1(n6088), .A2(n6087), .ZN(n6084) );
  AND2_X1 U6062 ( .A1(n6089), .A2(n6090), .ZN(n6087) );
  INV_X1 U6063 ( .A(n6091), .ZN(n6090) );
  AND2_X1 U6064 ( .A1(n6092), .A2(n6093), .ZN(n6091) );
  OR2_X1 U6065 ( .A1(n6093), .A2(n6092), .ZN(n6089) );
  INV_X1 U6066 ( .A(n6094), .ZN(n6092) );
  INV_X1 U6067 ( .A(n5923), .ZN(n6031) );
  AND2_X1 U6068 ( .A1(b_7_), .A2(a_9_), .ZN(n5923) );
  OR2_X1 U6069 ( .A1(n6027), .A2(n5930), .ZN(n6028) );
  OR2_X1 U6070 ( .A1(n6095), .A2(n6096), .ZN(n5930) );
  INV_X1 U6071 ( .A(n6097), .ZN(n6096) );
  OR2_X1 U6072 ( .A1(n6098), .A2(n6099), .ZN(n6097) );
  AND2_X1 U6073 ( .A1(n6099), .A2(n6098), .ZN(n6095) );
  AND2_X1 U6074 ( .A1(n6100), .A2(n6101), .ZN(n6098) );
  INV_X1 U6075 ( .A(n6102), .ZN(n6101) );
  AND2_X1 U6076 ( .A1(n6103), .A2(n6104), .ZN(n6102) );
  OR2_X1 U6077 ( .A1(n6104), .A2(n6103), .ZN(n6100) );
  INV_X1 U6078 ( .A(n5934), .ZN(n6027) );
  AND2_X1 U6079 ( .A1(b_7_), .A2(a_8_), .ZN(n5934) );
  OR2_X1 U6080 ( .A1(n6105), .A2(n6106), .ZN(n5940) );
  INV_X1 U6081 ( .A(n6107), .ZN(n6106) );
  OR2_X1 U6082 ( .A1(n6108), .A2(n6109), .ZN(n6107) );
  AND2_X1 U6083 ( .A1(n6109), .A2(n6108), .ZN(n6105) );
  AND2_X1 U6084 ( .A1(n6110), .A2(n6111), .ZN(n6108) );
  INV_X1 U6085 ( .A(n6112), .ZN(n6111) );
  AND2_X1 U6086 ( .A1(n6113), .A2(n6114), .ZN(n6112) );
  OR2_X1 U6087 ( .A1(n6114), .A2(n6113), .ZN(n6110) );
  OR2_X1 U6088 ( .A1(n6020), .A2(n5949), .ZN(n6021) );
  OR2_X1 U6089 ( .A1(n6115), .A2(n6116), .ZN(n5949) );
  INV_X1 U6090 ( .A(n6117), .ZN(n6116) );
  OR2_X1 U6091 ( .A1(n6118), .A2(n6119), .ZN(n6117) );
  AND2_X1 U6092 ( .A1(n6119), .A2(n6118), .ZN(n6115) );
  AND2_X1 U6093 ( .A1(n6120), .A2(n6121), .ZN(n6118) );
  INV_X1 U6094 ( .A(n6122), .ZN(n6121) );
  AND2_X1 U6095 ( .A1(n6123), .A2(n6124), .ZN(n6122) );
  OR2_X1 U6096 ( .A1(n6124), .A2(n6123), .ZN(n6120) );
  INV_X1 U6097 ( .A(n5953), .ZN(n6020) );
  AND2_X1 U6098 ( .A1(b_7_), .A2(a_6_), .ZN(n5953) );
  AND2_X1 U6099 ( .A1(n6125), .A2(n6126), .ZN(n5959) );
  INV_X1 U6100 ( .A(n6127), .ZN(n6126) );
  AND2_X1 U6101 ( .A1(n6128), .A2(n6129), .ZN(n6127) );
  OR2_X1 U6102 ( .A1(n6129), .A2(n6128), .ZN(n6125) );
  OR2_X1 U6103 ( .A1(n6130), .A2(n6131), .ZN(n6128) );
  INV_X1 U6104 ( .A(n6132), .ZN(n6131) );
  OR2_X1 U6105 ( .A1(n3792), .A2(n6133), .ZN(n6132) );
  AND2_X1 U6106 ( .A1(n6133), .A2(n3792), .ZN(n6130) );
  INV_X1 U6107 ( .A(n6134), .ZN(n6133) );
  AND2_X1 U6108 ( .A1(n6135), .A2(n6136), .ZN(n5969) );
  INV_X1 U6109 ( .A(n6137), .ZN(n6136) );
  AND2_X1 U6110 ( .A1(n6138), .A2(n6139), .ZN(n6137) );
  OR2_X1 U6111 ( .A1(n6139), .A2(n6138), .ZN(n6135) );
  OR2_X1 U6112 ( .A1(n6140), .A2(n6141), .ZN(n6138) );
  AND2_X1 U6113 ( .A1(n6142), .A2(n6143), .ZN(n6141) );
  INV_X1 U6114 ( .A(n6144), .ZN(n6140) );
  OR2_X1 U6115 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  AND2_X1 U6116 ( .A1(n6145), .A2(n6146), .ZN(n5979) );
  INV_X1 U6117 ( .A(n6147), .ZN(n6146) );
  AND2_X1 U6118 ( .A1(n6148), .A2(n6149), .ZN(n6147) );
  OR2_X1 U6119 ( .A1(n6149), .A2(n6148), .ZN(n6145) );
  OR2_X1 U6120 ( .A1(n6150), .A2(n6151), .ZN(n6148) );
  AND2_X1 U6121 ( .A1(n6152), .A2(n6153), .ZN(n6151) );
  INV_X1 U6122 ( .A(n6154), .ZN(n6150) );
  OR2_X1 U6123 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  AND2_X1 U6124 ( .A1(n6155), .A2(n6156), .ZN(n5989) );
  INV_X1 U6125 ( .A(n6157), .ZN(n6156) );
  AND2_X1 U6126 ( .A1(n6158), .A2(n6159), .ZN(n6157) );
  OR2_X1 U6127 ( .A1(n6159), .A2(n6158), .ZN(n6155) );
  OR2_X1 U6128 ( .A1(n6160), .A2(n6161), .ZN(n6158) );
  AND2_X1 U6129 ( .A1(n6162), .A2(n6163), .ZN(n6161) );
  INV_X1 U6130 ( .A(n6164), .ZN(n6160) );
  OR2_X1 U6131 ( .A1(n6163), .A2(n6162), .ZN(n6164) );
  AND2_X1 U6132 ( .A1(n6165), .A2(n6166), .ZN(n4316) );
  INV_X1 U6133 ( .A(n6167), .ZN(n6166) );
  AND2_X1 U6134 ( .A1(n6168), .A2(n4330), .ZN(n6167) );
  OR2_X1 U6135 ( .A1(n4330), .A2(n6168), .ZN(n6165) );
  OR2_X1 U6136 ( .A1(n6169), .A2(n6170), .ZN(n6168) );
  AND2_X1 U6137 ( .A1(n4332), .A2(n4329), .ZN(n6170) );
  INV_X1 U6138 ( .A(n6171), .ZN(n6169) );
  OR2_X1 U6139 ( .A1(n4329), .A2(n4332), .ZN(n6171) );
  AND2_X1 U6140 ( .A1(b_6_), .A2(a_2_), .ZN(n4332) );
  OR2_X1 U6141 ( .A1(n6172), .A2(n6173), .ZN(n4329) );
  AND2_X1 U6142 ( .A1(n6174), .A2(n6163), .ZN(n6173) );
  AND2_X1 U6143 ( .A1(n6159), .A2(n6175), .ZN(n6172) );
  OR2_X1 U6144 ( .A1(n6163), .A2(n6174), .ZN(n6175) );
  INV_X1 U6145 ( .A(n6162), .ZN(n6174) );
  AND2_X1 U6146 ( .A1(b_6_), .A2(a_3_), .ZN(n6162) );
  OR2_X1 U6147 ( .A1(n6176), .A2(n6177), .ZN(n6163) );
  AND2_X1 U6148 ( .A1(n6178), .A2(n6153), .ZN(n6177) );
  AND2_X1 U6149 ( .A1(n6149), .A2(n6179), .ZN(n6176) );
  OR2_X1 U6150 ( .A1(n6153), .A2(n6178), .ZN(n6179) );
  INV_X1 U6151 ( .A(n6152), .ZN(n6178) );
  AND2_X1 U6152 ( .A1(b_6_), .A2(a_4_), .ZN(n6152) );
  OR2_X1 U6153 ( .A1(n6180), .A2(n6181), .ZN(n6153) );
  AND2_X1 U6154 ( .A1(n6182), .A2(n6143), .ZN(n6181) );
  AND2_X1 U6155 ( .A1(n6139), .A2(n6183), .ZN(n6180) );
  OR2_X1 U6156 ( .A1(n6143), .A2(n6182), .ZN(n6183) );
  INV_X1 U6157 ( .A(n6142), .ZN(n6182) );
  AND2_X1 U6158 ( .A1(b_6_), .A2(a_5_), .ZN(n6142) );
  OR2_X1 U6159 ( .A1(n6184), .A2(n6185), .ZN(n6143) );
  AND2_X1 U6160 ( .A1(n3792), .A2(n6134), .ZN(n6185) );
  AND2_X1 U6161 ( .A1(n6129), .A2(n6186), .ZN(n6184) );
  OR2_X1 U6162 ( .A1(n6134), .A2(n3792), .ZN(n6186) );
  OR2_X1 U6163 ( .A1(n4235), .A2(n6187), .ZN(n3792) );
  OR2_X1 U6164 ( .A1(n6188), .A2(n6189), .ZN(n6134) );
  AND2_X1 U6165 ( .A1(n6119), .A2(n6190), .ZN(n6189) );
  AND2_X1 U6166 ( .A1(n6191), .A2(n6124), .ZN(n6188) );
  OR2_X1 U6167 ( .A1(n6192), .A2(n6193), .ZN(n6124) );
  AND2_X1 U6168 ( .A1(n6194), .A2(n6114), .ZN(n6193) );
  AND2_X1 U6169 ( .A1(n6109), .A2(n6195), .ZN(n6192) );
  OR2_X1 U6170 ( .A1(n6114), .A2(n6194), .ZN(n6195) );
  INV_X1 U6171 ( .A(n6113), .ZN(n6194) );
  AND2_X1 U6172 ( .A1(b_6_), .A2(a_8_), .ZN(n6113) );
  OR2_X1 U6173 ( .A1(n6196), .A2(n6197), .ZN(n6114) );
  AND2_X1 U6174 ( .A1(n6099), .A2(n6198), .ZN(n6197) );
  AND2_X1 U6175 ( .A1(n6199), .A2(n6104), .ZN(n6196) );
  OR2_X1 U6176 ( .A1(n6200), .A2(n6201), .ZN(n6104) );
  AND2_X1 U6177 ( .A1(n6088), .A2(n6094), .ZN(n6201) );
  AND2_X1 U6178 ( .A1(n6202), .A2(n6093), .ZN(n6200) );
  OR2_X1 U6179 ( .A1(n6203), .A2(n6204), .ZN(n6093) );
  AND2_X1 U6180 ( .A1(n6078), .A2(n6205), .ZN(n6204) );
  AND2_X1 U6181 ( .A1(n6206), .A2(n6083), .ZN(n6203) );
  OR2_X1 U6182 ( .A1(n6207), .A2(n6208), .ZN(n6083) );
  AND2_X1 U6183 ( .A1(n6068), .A2(n6209), .ZN(n6208) );
  AND2_X1 U6184 ( .A1(n6210), .A2(n6073), .ZN(n6207) );
  OR2_X1 U6185 ( .A1(n6211), .A2(n6212), .ZN(n6073) );
  AND2_X1 U6186 ( .A1(n6056), .A2(n6061), .ZN(n6212) );
  AND2_X1 U6187 ( .A1(n6060), .A2(n6213), .ZN(n6211) );
  OR2_X1 U6188 ( .A1(n6061), .A2(n6056), .ZN(n6213) );
  OR2_X1 U6189 ( .A1(n3631), .A2(n4235), .ZN(n6056) );
  INV_X1 U6190 ( .A(n6062), .ZN(n6061) );
  AND3_X1 U6191 ( .A1(n3975), .A2(b_6_), .A3(b_5_), .ZN(n6062) );
  INV_X1 U6192 ( .A(n6063), .ZN(n6060) );
  OR2_X1 U6193 ( .A1(n6214), .A2(n6215), .ZN(n6063) );
  AND2_X1 U6194 ( .A1(b_5_), .A2(n6216), .ZN(n6215) );
  OR2_X1 U6195 ( .A1(n6217), .A2(n3592), .ZN(n6216) );
  AND2_X1 U6196 ( .A1(a_14_), .A2(n4121), .ZN(n6217) );
  AND2_X1 U6197 ( .A1(b_4_), .A2(n6218), .ZN(n6214) );
  OR2_X1 U6198 ( .A1(n6219), .A2(n3595), .ZN(n6218) );
  AND2_X1 U6199 ( .A1(a_15_), .A2(n3812), .ZN(n6219) );
  OR2_X1 U6200 ( .A1(n6209), .A2(n6068), .ZN(n6210) );
  OR2_X1 U6201 ( .A1(n6220), .A2(n6221), .ZN(n6068) );
  AND2_X1 U6202 ( .A1(n6222), .A2(n6223), .ZN(n6221) );
  INV_X1 U6203 ( .A(n6224), .ZN(n6220) );
  OR2_X1 U6204 ( .A1(n6222), .A2(n6223), .ZN(n6224) );
  OR2_X1 U6205 ( .A1(n6225), .A2(n6226), .ZN(n6222) );
  AND2_X1 U6206 ( .A1(n6227), .A2(n6228), .ZN(n6226) );
  AND2_X1 U6207 ( .A1(n6229), .A2(n6230), .ZN(n6225) );
  INV_X1 U6208 ( .A(n6072), .ZN(n6209) );
  AND2_X1 U6209 ( .A1(a_12_), .A2(b_6_), .ZN(n6072) );
  OR2_X1 U6210 ( .A1(n6205), .A2(n6078), .ZN(n6206) );
  OR2_X1 U6211 ( .A1(n6231), .A2(n6232), .ZN(n6078) );
  INV_X1 U6212 ( .A(n6233), .ZN(n6232) );
  OR2_X1 U6213 ( .A1(n6234), .A2(n6235), .ZN(n6233) );
  AND2_X1 U6214 ( .A1(n6235), .A2(n6234), .ZN(n6231) );
  AND2_X1 U6215 ( .A1(n6236), .A2(n6237), .ZN(n6234) );
  INV_X1 U6216 ( .A(n6238), .ZN(n6237) );
  AND2_X1 U6217 ( .A1(n6239), .A2(n6240), .ZN(n6238) );
  OR2_X1 U6218 ( .A1(n6240), .A2(n6239), .ZN(n6236) );
  INV_X1 U6219 ( .A(n6082), .ZN(n6205) );
  AND2_X1 U6220 ( .A1(a_11_), .A2(b_6_), .ZN(n6082) );
  OR2_X1 U6221 ( .A1(n6094), .A2(n6088), .ZN(n6202) );
  OR2_X1 U6222 ( .A1(n6241), .A2(n6242), .ZN(n6088) );
  INV_X1 U6223 ( .A(n6243), .ZN(n6242) );
  OR2_X1 U6224 ( .A1(n6244), .A2(n6245), .ZN(n6243) );
  AND2_X1 U6225 ( .A1(n6245), .A2(n6244), .ZN(n6241) );
  AND2_X1 U6226 ( .A1(n6246), .A2(n6247), .ZN(n6244) );
  INV_X1 U6227 ( .A(n6248), .ZN(n6247) );
  AND2_X1 U6228 ( .A1(n6249), .A2(n6250), .ZN(n6248) );
  OR2_X1 U6229 ( .A1(n6250), .A2(n6249), .ZN(n6246) );
  OR2_X1 U6230 ( .A1(n4235), .A2(n3964), .ZN(n6094) );
  INV_X1 U6231 ( .A(b_6_), .ZN(n4235) );
  OR2_X1 U6232 ( .A1(n6198), .A2(n6099), .ZN(n6199) );
  OR2_X1 U6233 ( .A1(n6251), .A2(n6252), .ZN(n6099) );
  INV_X1 U6234 ( .A(n6253), .ZN(n6252) );
  OR2_X1 U6235 ( .A1(n6254), .A2(n6255), .ZN(n6253) );
  AND2_X1 U6236 ( .A1(n6255), .A2(n6254), .ZN(n6251) );
  AND2_X1 U6237 ( .A1(n6256), .A2(n6257), .ZN(n6254) );
  INV_X1 U6238 ( .A(n6258), .ZN(n6257) );
  AND2_X1 U6239 ( .A1(n6259), .A2(n6260), .ZN(n6258) );
  OR2_X1 U6240 ( .A1(n6260), .A2(n6259), .ZN(n6256) );
  INV_X1 U6241 ( .A(n6261), .ZN(n6259) );
  INV_X1 U6242 ( .A(n6103), .ZN(n6198) );
  AND2_X1 U6243 ( .A1(b_6_), .A2(a_9_), .ZN(n6103) );
  OR2_X1 U6244 ( .A1(n6262), .A2(n6263), .ZN(n6109) );
  INV_X1 U6245 ( .A(n6264), .ZN(n6263) );
  OR2_X1 U6246 ( .A1(n6265), .A2(n6266), .ZN(n6264) );
  AND2_X1 U6247 ( .A1(n6266), .A2(n6265), .ZN(n6262) );
  AND2_X1 U6248 ( .A1(n6267), .A2(n6268), .ZN(n6265) );
  INV_X1 U6249 ( .A(n6269), .ZN(n6268) );
  AND2_X1 U6250 ( .A1(n6270), .A2(n6271), .ZN(n6269) );
  OR2_X1 U6251 ( .A1(n6271), .A2(n6270), .ZN(n6267) );
  OR2_X1 U6252 ( .A1(n6190), .A2(n6119), .ZN(n6191) );
  OR2_X1 U6253 ( .A1(n6272), .A2(n6273), .ZN(n6119) );
  INV_X1 U6254 ( .A(n6274), .ZN(n6273) );
  OR2_X1 U6255 ( .A1(n6275), .A2(n6276), .ZN(n6274) );
  AND2_X1 U6256 ( .A1(n6276), .A2(n6275), .ZN(n6272) );
  AND2_X1 U6257 ( .A1(n6277), .A2(n6278), .ZN(n6275) );
  INV_X1 U6258 ( .A(n6279), .ZN(n6278) );
  AND2_X1 U6259 ( .A1(n6280), .A2(n6281), .ZN(n6279) );
  OR2_X1 U6260 ( .A1(n6281), .A2(n6280), .ZN(n6277) );
  INV_X1 U6261 ( .A(n6123), .ZN(n6190) );
  AND2_X1 U6262 ( .A1(b_6_), .A2(a_7_), .ZN(n6123) );
  AND2_X1 U6263 ( .A1(n6282), .A2(n6283), .ZN(n6129) );
  INV_X1 U6264 ( .A(n6284), .ZN(n6283) );
  AND2_X1 U6265 ( .A1(n6285), .A2(n6286), .ZN(n6284) );
  OR2_X1 U6266 ( .A1(n6286), .A2(n6285), .ZN(n6282) );
  OR2_X1 U6267 ( .A1(n6287), .A2(n6288), .ZN(n6285) );
  AND2_X1 U6268 ( .A1(n6289), .A2(n6290), .ZN(n6288) );
  INV_X1 U6269 ( .A(n6291), .ZN(n6287) );
  OR2_X1 U6270 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  AND2_X1 U6271 ( .A1(n6292), .A2(n6293), .ZN(n6139) );
  INV_X1 U6272 ( .A(n6294), .ZN(n6293) );
  AND2_X1 U6273 ( .A1(n6295), .A2(n6296), .ZN(n6294) );
  OR2_X1 U6274 ( .A1(n6296), .A2(n6295), .ZN(n6292) );
  OR2_X1 U6275 ( .A1(n6297), .A2(n6298), .ZN(n6295) );
  AND2_X1 U6276 ( .A1(n6299), .A2(n6300), .ZN(n6298) );
  INV_X1 U6277 ( .A(n6301), .ZN(n6297) );
  OR2_X1 U6278 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  AND2_X1 U6279 ( .A1(n6302), .A2(n6303), .ZN(n6149) );
  INV_X1 U6280 ( .A(n6304), .ZN(n6303) );
  AND2_X1 U6281 ( .A1(n6305), .A2(n6306), .ZN(n6304) );
  OR2_X1 U6282 ( .A1(n6306), .A2(n6305), .ZN(n6302) );
  OR2_X1 U6283 ( .A1(n6307), .A2(n6308), .ZN(n6305) );
  AND2_X1 U6284 ( .A1(n3810), .A2(n6309), .ZN(n6308) );
  INV_X1 U6285 ( .A(n6310), .ZN(n6307) );
  OR2_X1 U6286 ( .A1(n6309), .A2(n3810), .ZN(n6310) );
  AND2_X1 U6287 ( .A1(n6311), .A2(n6312), .ZN(n6159) );
  INV_X1 U6288 ( .A(n6313), .ZN(n6312) );
  AND2_X1 U6289 ( .A1(n6314), .A2(n6315), .ZN(n6313) );
  OR2_X1 U6290 ( .A1(n6315), .A2(n6314), .ZN(n6311) );
  OR2_X1 U6291 ( .A1(n6316), .A2(n6317), .ZN(n6314) );
  AND2_X1 U6292 ( .A1(n6318), .A2(n6319), .ZN(n6317) );
  INV_X1 U6293 ( .A(n6320), .ZN(n6316) );
  OR2_X1 U6294 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  AND2_X1 U6295 ( .A1(n6321), .A2(n6322), .ZN(n4330) );
  INV_X1 U6296 ( .A(n6323), .ZN(n6322) );
  AND2_X1 U6297 ( .A1(n6324), .A2(n4344), .ZN(n6323) );
  OR2_X1 U6298 ( .A1(n4344), .A2(n6324), .ZN(n6321) );
  OR2_X1 U6299 ( .A1(n6325), .A2(n6326), .ZN(n6324) );
  AND2_X1 U6300 ( .A1(n4346), .A2(n4343), .ZN(n6326) );
  INV_X1 U6301 ( .A(n6327), .ZN(n6325) );
  OR2_X1 U6302 ( .A1(n4343), .A2(n4346), .ZN(n6327) );
  AND2_X1 U6303 ( .A1(b_5_), .A2(a_3_), .ZN(n4346) );
  OR2_X1 U6304 ( .A1(n6328), .A2(n6329), .ZN(n4343) );
  AND2_X1 U6305 ( .A1(n6330), .A2(n6319), .ZN(n6329) );
  AND2_X1 U6306 ( .A1(n6315), .A2(n6331), .ZN(n6328) );
  OR2_X1 U6307 ( .A1(n6319), .A2(n6330), .ZN(n6331) );
  INV_X1 U6308 ( .A(n6318), .ZN(n6330) );
  AND2_X1 U6309 ( .A1(b_5_), .A2(a_4_), .ZN(n6318) );
  OR2_X1 U6310 ( .A1(n6332), .A2(n6333), .ZN(n6319) );
  AND2_X1 U6311 ( .A1(n3952), .A2(n6309), .ZN(n6333) );
  AND2_X1 U6312 ( .A1(n6306), .A2(n6334), .ZN(n6332) );
  OR2_X1 U6313 ( .A1(n6309), .A2(n3952), .ZN(n6334) );
  INV_X1 U6314 ( .A(n3810), .ZN(n3952) );
  AND2_X1 U6315 ( .A1(b_5_), .A2(a_5_), .ZN(n3810) );
  OR2_X1 U6316 ( .A1(n6335), .A2(n6336), .ZN(n6309) );
  AND2_X1 U6317 ( .A1(n6337), .A2(n6300), .ZN(n6336) );
  AND2_X1 U6318 ( .A1(n6296), .A2(n6338), .ZN(n6335) );
  OR2_X1 U6319 ( .A1(n6300), .A2(n6337), .ZN(n6338) );
  INV_X1 U6320 ( .A(n6299), .ZN(n6337) );
  AND2_X1 U6321 ( .A1(b_5_), .A2(a_6_), .ZN(n6299) );
  OR2_X1 U6322 ( .A1(n6339), .A2(n6340), .ZN(n6300) );
  AND2_X1 U6323 ( .A1(n6341), .A2(n6290), .ZN(n6340) );
  AND2_X1 U6324 ( .A1(n6286), .A2(n6342), .ZN(n6339) );
  OR2_X1 U6325 ( .A1(n6290), .A2(n6341), .ZN(n6342) );
  INV_X1 U6326 ( .A(n6289), .ZN(n6341) );
  AND2_X1 U6327 ( .A1(b_5_), .A2(a_7_), .ZN(n6289) );
  OR2_X1 U6328 ( .A1(n6343), .A2(n6344), .ZN(n6290) );
  AND2_X1 U6329 ( .A1(n6276), .A2(n6345), .ZN(n6344) );
  AND2_X1 U6330 ( .A1(n6346), .A2(n6281), .ZN(n6343) );
  OR2_X1 U6331 ( .A1(n6347), .A2(n6348), .ZN(n6281) );
  AND2_X1 U6332 ( .A1(n6349), .A2(n6271), .ZN(n6348) );
  AND2_X1 U6333 ( .A1(n6266), .A2(n6350), .ZN(n6347) );
  OR2_X1 U6334 ( .A1(n6271), .A2(n6349), .ZN(n6350) );
  INV_X1 U6335 ( .A(n6270), .ZN(n6349) );
  AND2_X1 U6336 ( .A1(b_5_), .A2(a_9_), .ZN(n6270) );
  OR2_X1 U6337 ( .A1(n6351), .A2(n6352), .ZN(n6271) );
  AND2_X1 U6338 ( .A1(n6255), .A2(n6261), .ZN(n6352) );
  AND2_X1 U6339 ( .A1(n6353), .A2(n6260), .ZN(n6351) );
  OR2_X1 U6340 ( .A1(n6354), .A2(n6355), .ZN(n6260) );
  AND2_X1 U6341 ( .A1(n6245), .A2(n6356), .ZN(n6355) );
  AND2_X1 U6342 ( .A1(n6357), .A2(n6250), .ZN(n6354) );
  OR2_X1 U6343 ( .A1(n6358), .A2(n6359), .ZN(n6250) );
  AND2_X1 U6344 ( .A1(n6235), .A2(n6360), .ZN(n6359) );
  AND2_X1 U6345 ( .A1(n6361), .A2(n6240), .ZN(n6358) );
  OR2_X1 U6346 ( .A1(n6362), .A2(n6363), .ZN(n6240) );
  AND2_X1 U6347 ( .A1(n6223), .A2(n6228), .ZN(n6363) );
  AND2_X1 U6348 ( .A1(n6227), .A2(n6364), .ZN(n6362) );
  OR2_X1 U6349 ( .A1(n6228), .A2(n6223), .ZN(n6364) );
  OR2_X1 U6350 ( .A1(n3631), .A2(n3812), .ZN(n6223) );
  INV_X1 U6351 ( .A(n6229), .ZN(n6228) );
  AND3_X1 U6352 ( .A1(n3975), .A2(b_5_), .A3(b_4_), .ZN(n6229) );
  INV_X1 U6353 ( .A(n6230), .ZN(n6227) );
  OR2_X1 U6354 ( .A1(n6365), .A2(n6366), .ZN(n6230) );
  AND2_X1 U6355 ( .A1(b_4_), .A2(n6367), .ZN(n6366) );
  OR2_X1 U6356 ( .A1(n6368), .A2(n3592), .ZN(n6367) );
  AND2_X1 U6357 ( .A1(a_14_), .A2(n3867), .ZN(n6368) );
  AND2_X1 U6358 ( .A1(b_3_), .A2(n6369), .ZN(n6365) );
  OR2_X1 U6359 ( .A1(n6370), .A2(n3595), .ZN(n6369) );
  AND2_X1 U6360 ( .A1(a_15_), .A2(n4121), .ZN(n6370) );
  OR2_X1 U6361 ( .A1(n6360), .A2(n6235), .ZN(n6361) );
  OR2_X1 U6362 ( .A1(n6371), .A2(n6372), .ZN(n6235) );
  AND2_X1 U6363 ( .A1(n6373), .A2(n6374), .ZN(n6372) );
  INV_X1 U6364 ( .A(n6375), .ZN(n6371) );
  OR2_X1 U6365 ( .A1(n6373), .A2(n6374), .ZN(n6375) );
  OR2_X1 U6366 ( .A1(n6376), .A2(n6377), .ZN(n6373) );
  AND2_X1 U6367 ( .A1(n6378), .A2(n6379), .ZN(n6377) );
  AND2_X1 U6368 ( .A1(n6380), .A2(n6381), .ZN(n6376) );
  INV_X1 U6369 ( .A(n6239), .ZN(n6360) );
  AND2_X1 U6370 ( .A1(a_12_), .A2(b_5_), .ZN(n6239) );
  OR2_X1 U6371 ( .A1(n6356), .A2(n6245), .ZN(n6357) );
  OR2_X1 U6372 ( .A1(n6382), .A2(n6383), .ZN(n6245) );
  INV_X1 U6373 ( .A(n6384), .ZN(n6383) );
  OR2_X1 U6374 ( .A1(n6385), .A2(n6386), .ZN(n6384) );
  AND2_X1 U6375 ( .A1(n6386), .A2(n6385), .ZN(n6382) );
  AND2_X1 U6376 ( .A1(n6387), .A2(n6388), .ZN(n6385) );
  INV_X1 U6377 ( .A(n6389), .ZN(n6388) );
  AND2_X1 U6378 ( .A1(n6390), .A2(n6391), .ZN(n6389) );
  OR2_X1 U6379 ( .A1(n6391), .A2(n6390), .ZN(n6387) );
  INV_X1 U6380 ( .A(n6249), .ZN(n6356) );
  AND2_X1 U6381 ( .A1(a_11_), .A2(b_5_), .ZN(n6249) );
  OR2_X1 U6382 ( .A1(n6261), .A2(n6255), .ZN(n6353) );
  OR2_X1 U6383 ( .A1(n6392), .A2(n6393), .ZN(n6255) );
  INV_X1 U6384 ( .A(n6394), .ZN(n6393) );
  OR2_X1 U6385 ( .A1(n6395), .A2(n6396), .ZN(n6394) );
  AND2_X1 U6386 ( .A1(n6396), .A2(n6395), .ZN(n6392) );
  AND2_X1 U6387 ( .A1(n6397), .A2(n6398), .ZN(n6395) );
  INV_X1 U6388 ( .A(n6399), .ZN(n6398) );
  AND2_X1 U6389 ( .A1(n6400), .A2(n6401), .ZN(n6399) );
  OR2_X1 U6390 ( .A1(n6401), .A2(n6400), .ZN(n6397) );
  OR2_X1 U6391 ( .A1(n3964), .A2(n3812), .ZN(n6261) );
  INV_X1 U6392 ( .A(b_5_), .ZN(n3812) );
  OR2_X1 U6393 ( .A1(n6402), .A2(n6403), .ZN(n6266) );
  INV_X1 U6394 ( .A(n6404), .ZN(n6403) );
  OR2_X1 U6395 ( .A1(n6405), .A2(n6406), .ZN(n6404) );
  AND2_X1 U6396 ( .A1(n6406), .A2(n6405), .ZN(n6402) );
  AND2_X1 U6397 ( .A1(n6407), .A2(n6408), .ZN(n6405) );
  INV_X1 U6398 ( .A(n6409), .ZN(n6408) );
  AND2_X1 U6399 ( .A1(n6410), .A2(n6411), .ZN(n6409) );
  OR2_X1 U6400 ( .A1(n6411), .A2(n6410), .ZN(n6407) );
  INV_X1 U6401 ( .A(n6412), .ZN(n6410) );
  OR2_X1 U6402 ( .A1(n6345), .A2(n6276), .ZN(n6346) );
  OR2_X1 U6403 ( .A1(n6413), .A2(n6414), .ZN(n6276) );
  INV_X1 U6404 ( .A(n6415), .ZN(n6414) );
  OR2_X1 U6405 ( .A1(n6416), .A2(n6417), .ZN(n6415) );
  AND2_X1 U6406 ( .A1(n6417), .A2(n6416), .ZN(n6413) );
  AND2_X1 U6407 ( .A1(n6418), .A2(n6419), .ZN(n6416) );
  INV_X1 U6408 ( .A(n6420), .ZN(n6419) );
  AND2_X1 U6409 ( .A1(n6421), .A2(n6422), .ZN(n6420) );
  OR2_X1 U6410 ( .A1(n6422), .A2(n6421), .ZN(n6418) );
  INV_X1 U6411 ( .A(n6280), .ZN(n6345) );
  AND2_X1 U6412 ( .A1(b_5_), .A2(a_8_), .ZN(n6280) );
  AND2_X1 U6413 ( .A1(n6423), .A2(n6424), .ZN(n6286) );
  INV_X1 U6414 ( .A(n6425), .ZN(n6424) );
  AND2_X1 U6415 ( .A1(n6426), .A2(n6427), .ZN(n6425) );
  OR2_X1 U6416 ( .A1(n6427), .A2(n6426), .ZN(n6423) );
  OR2_X1 U6417 ( .A1(n6428), .A2(n6429), .ZN(n6426) );
  AND2_X1 U6418 ( .A1(n6430), .A2(n6431), .ZN(n6429) );
  INV_X1 U6419 ( .A(n6432), .ZN(n6428) );
  OR2_X1 U6420 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  AND2_X1 U6421 ( .A1(n6433), .A2(n6434), .ZN(n6296) );
  INV_X1 U6422 ( .A(n6435), .ZN(n6434) );
  AND2_X1 U6423 ( .A1(n6436), .A2(n6437), .ZN(n6435) );
  OR2_X1 U6424 ( .A1(n6437), .A2(n6436), .ZN(n6433) );
  OR2_X1 U6425 ( .A1(n6438), .A2(n6439), .ZN(n6436) );
  AND2_X1 U6426 ( .A1(n6440), .A2(n6441), .ZN(n6439) );
  INV_X1 U6427 ( .A(n6442), .ZN(n6438) );
  OR2_X1 U6428 ( .A1(n6441), .A2(n6440), .ZN(n6442) );
  AND2_X1 U6429 ( .A1(n6443), .A2(n6444), .ZN(n6306) );
  INV_X1 U6430 ( .A(n6445), .ZN(n6444) );
  AND2_X1 U6431 ( .A1(n6446), .A2(n6447), .ZN(n6445) );
  OR2_X1 U6432 ( .A1(n6447), .A2(n6446), .ZN(n6443) );
  OR2_X1 U6433 ( .A1(n6448), .A2(n6449), .ZN(n6446) );
  AND2_X1 U6434 ( .A1(n6450), .A2(n6451), .ZN(n6449) );
  INV_X1 U6435 ( .A(n6452), .ZN(n6448) );
  OR2_X1 U6436 ( .A1(n6451), .A2(n6450), .ZN(n6452) );
  AND2_X1 U6437 ( .A1(n6453), .A2(n6454), .ZN(n6315) );
  INV_X1 U6438 ( .A(n6455), .ZN(n6454) );
  AND2_X1 U6439 ( .A1(n6456), .A2(n6457), .ZN(n6455) );
  OR2_X1 U6440 ( .A1(n6457), .A2(n6456), .ZN(n6453) );
  OR2_X1 U6441 ( .A1(n6458), .A2(n6459), .ZN(n6456) );
  AND2_X1 U6442 ( .A1(n6460), .A2(n6461), .ZN(n6459) );
  INV_X1 U6443 ( .A(n6462), .ZN(n6458) );
  OR2_X1 U6444 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  AND2_X1 U6445 ( .A1(n6463), .A2(n6464), .ZN(n4344) );
  INV_X1 U6446 ( .A(n6465), .ZN(n6464) );
  AND2_X1 U6447 ( .A1(n6466), .A2(n4357), .ZN(n6465) );
  OR2_X1 U6448 ( .A1(n4357), .A2(n6466), .ZN(n6463) );
  OR2_X1 U6449 ( .A1(n6467), .A2(n6468), .ZN(n6466) );
  INV_X1 U6450 ( .A(n6469), .ZN(n6468) );
  OR2_X1 U6451 ( .A1(n3836), .A2(n6470), .ZN(n6469) );
  AND2_X1 U6452 ( .A1(n6470), .A2(n3836), .ZN(n6467) );
  OR2_X1 U6453 ( .A1(n4121), .A2(n6471), .ZN(n3836) );
  INV_X1 U6454 ( .A(n4356), .ZN(n6470) );
  OR2_X1 U6455 ( .A1(n6472), .A2(n6473), .ZN(n4356) );
  AND2_X1 U6456 ( .A1(n6474), .A2(n6461), .ZN(n6473) );
  AND2_X1 U6457 ( .A1(n6457), .A2(n6475), .ZN(n6472) );
  OR2_X1 U6458 ( .A1(n6461), .A2(n6474), .ZN(n6475) );
  INV_X1 U6459 ( .A(n6460), .ZN(n6474) );
  AND2_X1 U6460 ( .A1(b_4_), .A2(a_5_), .ZN(n6460) );
  OR2_X1 U6461 ( .A1(n6476), .A2(n6477), .ZN(n6461) );
  AND2_X1 U6462 ( .A1(n6478), .A2(n6451), .ZN(n6477) );
  AND2_X1 U6463 ( .A1(n6447), .A2(n6479), .ZN(n6476) );
  OR2_X1 U6464 ( .A1(n6451), .A2(n6478), .ZN(n6479) );
  INV_X1 U6465 ( .A(n6450), .ZN(n6478) );
  AND2_X1 U6466 ( .A1(b_4_), .A2(a_6_), .ZN(n6450) );
  OR2_X1 U6467 ( .A1(n6480), .A2(n6481), .ZN(n6451) );
  AND2_X1 U6468 ( .A1(n6482), .A2(n6441), .ZN(n6481) );
  AND2_X1 U6469 ( .A1(n6437), .A2(n6483), .ZN(n6480) );
  OR2_X1 U6470 ( .A1(n6441), .A2(n6482), .ZN(n6483) );
  INV_X1 U6471 ( .A(n6440), .ZN(n6482) );
  AND2_X1 U6472 ( .A1(b_4_), .A2(a_7_), .ZN(n6440) );
  OR2_X1 U6473 ( .A1(n6484), .A2(n6485), .ZN(n6441) );
  AND2_X1 U6474 ( .A1(n6486), .A2(n6431), .ZN(n6485) );
  AND2_X1 U6475 ( .A1(n6427), .A2(n6487), .ZN(n6484) );
  OR2_X1 U6476 ( .A1(n6431), .A2(n6486), .ZN(n6487) );
  INV_X1 U6477 ( .A(n6430), .ZN(n6486) );
  AND2_X1 U6478 ( .A1(b_4_), .A2(a_8_), .ZN(n6430) );
  OR2_X1 U6479 ( .A1(n6488), .A2(n6489), .ZN(n6431) );
  AND2_X1 U6480 ( .A1(n6417), .A2(n6490), .ZN(n6489) );
  AND2_X1 U6481 ( .A1(n6491), .A2(n6422), .ZN(n6488) );
  OR2_X1 U6482 ( .A1(n6492), .A2(n6493), .ZN(n6422) );
  AND2_X1 U6483 ( .A1(n6412), .A2(n6411), .ZN(n6493) );
  AND2_X1 U6484 ( .A1(n6406), .A2(n6494), .ZN(n6492) );
  OR2_X1 U6485 ( .A1(n6411), .A2(n6412), .ZN(n6494) );
  OR2_X1 U6486 ( .A1(n3964), .A2(n4121), .ZN(n6412) );
  OR2_X1 U6487 ( .A1(n6495), .A2(n6496), .ZN(n6411) );
  AND2_X1 U6488 ( .A1(n6396), .A2(n6497), .ZN(n6496) );
  AND2_X1 U6489 ( .A1(n6498), .A2(n6401), .ZN(n6495) );
  OR2_X1 U6490 ( .A1(n6499), .A2(n6500), .ZN(n6401) );
  AND2_X1 U6491 ( .A1(n6386), .A2(n6501), .ZN(n6500) );
  AND2_X1 U6492 ( .A1(n6502), .A2(n6391), .ZN(n6499) );
  OR2_X1 U6493 ( .A1(n6503), .A2(n6504), .ZN(n6391) );
  AND2_X1 U6494 ( .A1(n6374), .A2(n6379), .ZN(n6504) );
  AND2_X1 U6495 ( .A1(n6378), .A2(n6505), .ZN(n6503) );
  OR2_X1 U6496 ( .A1(n6379), .A2(n6374), .ZN(n6505) );
  OR2_X1 U6497 ( .A1(n3631), .A2(n4121), .ZN(n6374) );
  INV_X1 U6498 ( .A(b_4_), .ZN(n4121) );
  INV_X1 U6499 ( .A(n6380), .ZN(n6379) );
  AND3_X1 U6500 ( .A1(n3975), .A2(b_4_), .A3(b_3_), .ZN(n6380) );
  INV_X1 U6501 ( .A(n6381), .ZN(n6378) );
  OR2_X1 U6502 ( .A1(n6506), .A2(n6507), .ZN(n6381) );
  AND2_X1 U6503 ( .A1(b_3_), .A2(n6508), .ZN(n6507) );
  OR2_X1 U6504 ( .A1(n6509), .A2(n3592), .ZN(n6508) );
  AND2_X1 U6505 ( .A1(a_14_), .A2(n6510), .ZN(n6509) );
  AND2_X1 U6506 ( .A1(b_2_), .A2(n6511), .ZN(n6506) );
  OR2_X1 U6507 ( .A1(n6512), .A2(n3595), .ZN(n6511) );
  AND2_X1 U6508 ( .A1(a_15_), .A2(n3867), .ZN(n6512) );
  OR2_X1 U6509 ( .A1(n6501), .A2(n6386), .ZN(n6502) );
  OR2_X1 U6510 ( .A1(n6513), .A2(n6514), .ZN(n6386) );
  AND2_X1 U6511 ( .A1(n6515), .A2(n6516), .ZN(n6514) );
  INV_X1 U6512 ( .A(n6517), .ZN(n6513) );
  OR2_X1 U6513 ( .A1(n6515), .A2(n6516), .ZN(n6517) );
  OR2_X1 U6514 ( .A1(n6518), .A2(n6519), .ZN(n6515) );
  AND2_X1 U6515 ( .A1(n6520), .A2(n6521), .ZN(n6519) );
  AND2_X1 U6516 ( .A1(n6522), .A2(n6523), .ZN(n6518) );
  INV_X1 U6517 ( .A(n6390), .ZN(n6501) );
  AND2_X1 U6518 ( .A1(a_12_), .A2(b_4_), .ZN(n6390) );
  OR2_X1 U6519 ( .A1(n6497), .A2(n6396), .ZN(n6498) );
  OR2_X1 U6520 ( .A1(n6524), .A2(n6525), .ZN(n6396) );
  INV_X1 U6521 ( .A(n6526), .ZN(n6525) );
  OR2_X1 U6522 ( .A1(n6527), .A2(n6528), .ZN(n6526) );
  AND2_X1 U6523 ( .A1(n6528), .A2(n6527), .ZN(n6524) );
  AND2_X1 U6524 ( .A1(n6529), .A2(n6530), .ZN(n6527) );
  INV_X1 U6525 ( .A(n6531), .ZN(n6530) );
  AND2_X1 U6526 ( .A1(n6532), .A2(n6533), .ZN(n6531) );
  OR2_X1 U6527 ( .A1(n6533), .A2(n6532), .ZN(n6529) );
  INV_X1 U6528 ( .A(n6400), .ZN(n6497) );
  AND2_X1 U6529 ( .A1(a_11_), .A2(b_4_), .ZN(n6400) );
  OR2_X1 U6530 ( .A1(n6534), .A2(n6535), .ZN(n6406) );
  INV_X1 U6531 ( .A(n6536), .ZN(n6535) );
  OR2_X1 U6532 ( .A1(n6537), .A2(n6538), .ZN(n6536) );
  AND2_X1 U6533 ( .A1(n6538), .A2(n6537), .ZN(n6534) );
  AND2_X1 U6534 ( .A1(n6539), .A2(n6540), .ZN(n6537) );
  INV_X1 U6535 ( .A(n6541), .ZN(n6540) );
  AND2_X1 U6536 ( .A1(n6542), .A2(n6543), .ZN(n6541) );
  OR2_X1 U6537 ( .A1(n6543), .A2(n6542), .ZN(n6539) );
  OR2_X1 U6538 ( .A1(n6490), .A2(n6417), .ZN(n6491) );
  OR2_X1 U6539 ( .A1(n6544), .A2(n6545), .ZN(n6417) );
  INV_X1 U6540 ( .A(n6546), .ZN(n6545) );
  OR2_X1 U6541 ( .A1(n6547), .A2(n6548), .ZN(n6546) );
  AND2_X1 U6542 ( .A1(n6548), .A2(n6547), .ZN(n6544) );
  AND2_X1 U6543 ( .A1(n6549), .A2(n6550), .ZN(n6547) );
  INV_X1 U6544 ( .A(n6551), .ZN(n6550) );
  AND2_X1 U6545 ( .A1(n6552), .A2(n6553), .ZN(n6551) );
  OR2_X1 U6546 ( .A1(n6553), .A2(n6552), .ZN(n6549) );
  INV_X1 U6547 ( .A(n6554), .ZN(n6552) );
  INV_X1 U6548 ( .A(n6421), .ZN(n6490) );
  AND2_X1 U6549 ( .A1(a_9_), .A2(b_4_), .ZN(n6421) );
  AND2_X1 U6550 ( .A1(n6555), .A2(n6556), .ZN(n6427) );
  INV_X1 U6551 ( .A(n6557), .ZN(n6556) );
  AND2_X1 U6552 ( .A1(n6558), .A2(n6559), .ZN(n6557) );
  OR2_X1 U6553 ( .A1(n6559), .A2(n6558), .ZN(n6555) );
  OR2_X1 U6554 ( .A1(n6560), .A2(n6561), .ZN(n6558) );
  AND2_X1 U6555 ( .A1(n6562), .A2(n6563), .ZN(n6561) );
  INV_X1 U6556 ( .A(n6564), .ZN(n6560) );
  OR2_X1 U6557 ( .A1(n6563), .A2(n6562), .ZN(n6564) );
  AND2_X1 U6558 ( .A1(n6565), .A2(n6566), .ZN(n6437) );
  INV_X1 U6559 ( .A(n6567), .ZN(n6566) );
  AND2_X1 U6560 ( .A1(n6568), .A2(n6569), .ZN(n6567) );
  OR2_X1 U6561 ( .A1(n6569), .A2(n6568), .ZN(n6565) );
  OR2_X1 U6562 ( .A1(n6570), .A2(n6571), .ZN(n6568) );
  AND2_X1 U6563 ( .A1(n6572), .A2(n6573), .ZN(n6571) );
  INV_X1 U6564 ( .A(n6574), .ZN(n6570) );
  OR2_X1 U6565 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  AND2_X1 U6566 ( .A1(n6575), .A2(n6576), .ZN(n6447) );
  INV_X1 U6567 ( .A(n6577), .ZN(n6576) );
  AND2_X1 U6568 ( .A1(n6578), .A2(n6579), .ZN(n6577) );
  OR2_X1 U6569 ( .A1(n6579), .A2(n6578), .ZN(n6575) );
  OR2_X1 U6570 ( .A1(n6580), .A2(n6581), .ZN(n6578) );
  AND2_X1 U6571 ( .A1(n6582), .A2(n6583), .ZN(n6581) );
  INV_X1 U6572 ( .A(n6584), .ZN(n6580) );
  OR2_X1 U6573 ( .A1(n6583), .A2(n6582), .ZN(n6584) );
  AND2_X1 U6574 ( .A1(n6585), .A2(n6586), .ZN(n6457) );
  INV_X1 U6575 ( .A(n6587), .ZN(n6586) );
  AND2_X1 U6576 ( .A1(n6588), .A2(n6589), .ZN(n6587) );
  OR2_X1 U6577 ( .A1(n6589), .A2(n6588), .ZN(n6585) );
  OR2_X1 U6578 ( .A1(n6590), .A2(n6591), .ZN(n6588) );
  AND2_X1 U6579 ( .A1(n6592), .A2(n6593), .ZN(n6591) );
  INV_X1 U6580 ( .A(n6594), .ZN(n6590) );
  OR2_X1 U6581 ( .A1(n6593), .A2(n6592), .ZN(n6594) );
  AND2_X1 U6582 ( .A1(n6595), .A2(n6596), .ZN(n4357) );
  INV_X1 U6583 ( .A(n6597), .ZN(n6596) );
  AND2_X1 U6584 ( .A1(n6598), .A2(n4370), .ZN(n6597) );
  OR2_X1 U6585 ( .A1(n4370), .A2(n6598), .ZN(n6595) );
  OR2_X1 U6586 ( .A1(n6599), .A2(n6600), .ZN(n6598) );
  AND2_X1 U6587 ( .A1(n4372), .A2(n4369), .ZN(n6600) );
  INV_X1 U6588 ( .A(n6601), .ZN(n6599) );
  OR2_X1 U6589 ( .A1(n4369), .A2(n4372), .ZN(n6601) );
  AND2_X1 U6590 ( .A1(b_3_), .A2(a_5_), .ZN(n4372) );
  OR2_X1 U6591 ( .A1(n6602), .A2(n6603), .ZN(n4369) );
  AND2_X1 U6592 ( .A1(n6604), .A2(n6593), .ZN(n6603) );
  AND2_X1 U6593 ( .A1(n6589), .A2(n6605), .ZN(n6602) );
  OR2_X1 U6594 ( .A1(n6593), .A2(n6604), .ZN(n6605) );
  INV_X1 U6595 ( .A(n6592), .ZN(n6604) );
  AND2_X1 U6596 ( .A1(b_3_), .A2(a_6_), .ZN(n6592) );
  OR2_X1 U6597 ( .A1(n6606), .A2(n6607), .ZN(n6593) );
  AND2_X1 U6598 ( .A1(n6608), .A2(n6583), .ZN(n6607) );
  AND2_X1 U6599 ( .A1(n6579), .A2(n6609), .ZN(n6606) );
  OR2_X1 U6600 ( .A1(n6583), .A2(n6608), .ZN(n6609) );
  INV_X1 U6601 ( .A(n6582), .ZN(n6608) );
  AND2_X1 U6602 ( .A1(b_3_), .A2(a_7_), .ZN(n6582) );
  OR2_X1 U6603 ( .A1(n6610), .A2(n6611), .ZN(n6583) );
  AND2_X1 U6604 ( .A1(n6612), .A2(n6573), .ZN(n6611) );
  AND2_X1 U6605 ( .A1(n6569), .A2(n6613), .ZN(n6610) );
  OR2_X1 U6606 ( .A1(n6573), .A2(n6612), .ZN(n6613) );
  INV_X1 U6607 ( .A(n6572), .ZN(n6612) );
  AND2_X1 U6608 ( .A1(a_8_), .A2(b_3_), .ZN(n6572) );
  OR2_X1 U6609 ( .A1(n6614), .A2(n6615), .ZN(n6573) );
  AND2_X1 U6610 ( .A1(n6616), .A2(n6563), .ZN(n6615) );
  AND2_X1 U6611 ( .A1(n6559), .A2(n6617), .ZN(n6614) );
  OR2_X1 U6612 ( .A1(n6563), .A2(n6616), .ZN(n6617) );
  INV_X1 U6613 ( .A(n6562), .ZN(n6616) );
  AND2_X1 U6614 ( .A1(a_9_), .A2(b_3_), .ZN(n6562) );
  OR2_X1 U6615 ( .A1(n6618), .A2(n6619), .ZN(n6563) );
  AND2_X1 U6616 ( .A1(n6548), .A2(n6554), .ZN(n6619) );
  AND2_X1 U6617 ( .A1(n6620), .A2(n6553), .ZN(n6618) );
  OR2_X1 U6618 ( .A1(n6621), .A2(n6622), .ZN(n6553) );
  AND2_X1 U6619 ( .A1(n6623), .A2(n6543), .ZN(n6622) );
  AND2_X1 U6620 ( .A1(n6538), .A2(n6624), .ZN(n6621) );
  OR2_X1 U6621 ( .A1(n6543), .A2(n6623), .ZN(n6624) );
  INV_X1 U6622 ( .A(n6542), .ZN(n6623) );
  AND2_X1 U6623 ( .A1(a_11_), .A2(b_3_), .ZN(n6542) );
  OR2_X1 U6624 ( .A1(n6625), .A2(n6626), .ZN(n6543) );
  AND2_X1 U6625 ( .A1(n6528), .A2(n6627), .ZN(n6626) );
  AND2_X1 U6626 ( .A1(n6628), .A2(n6533), .ZN(n6625) );
  OR2_X1 U6627 ( .A1(n6629), .A2(n6630), .ZN(n6533) );
  AND2_X1 U6628 ( .A1(n6516), .A2(n6521), .ZN(n6630) );
  AND2_X1 U6629 ( .A1(n6520), .A2(n6631), .ZN(n6629) );
  OR2_X1 U6630 ( .A1(n6521), .A2(n6516), .ZN(n6631) );
  OR2_X1 U6631 ( .A1(n3631), .A2(n3867), .ZN(n6516) );
  INV_X1 U6632 ( .A(n6522), .ZN(n6521) );
  AND3_X1 U6633 ( .A1(n3975), .A2(b_3_), .A3(b_2_), .ZN(n6522) );
  INV_X1 U6634 ( .A(n6523), .ZN(n6520) );
  OR2_X1 U6635 ( .A1(n6632), .A2(n6633), .ZN(n6523) );
  AND2_X1 U6636 ( .A1(b_2_), .A2(n6634), .ZN(n6633) );
  OR2_X1 U6637 ( .A1(n6635), .A2(n3592), .ZN(n6634) );
  AND2_X1 U6638 ( .A1(a_14_), .A2(n3911), .ZN(n6635) );
  AND2_X1 U6639 ( .A1(b_1_), .A2(n6636), .ZN(n6632) );
  OR2_X1 U6640 ( .A1(n6637), .A2(n3595), .ZN(n6636) );
  AND2_X1 U6641 ( .A1(a_15_), .A2(n6510), .ZN(n6637) );
  OR2_X1 U6642 ( .A1(n6627), .A2(n6528), .ZN(n6628) );
  OR2_X1 U6643 ( .A1(n6638), .A2(n6639), .ZN(n6528) );
  AND2_X1 U6644 ( .A1(n6640), .A2(n6641), .ZN(n6639) );
  INV_X1 U6645 ( .A(n6642), .ZN(n6638) );
  OR2_X1 U6646 ( .A1(n6640), .A2(n6641), .ZN(n6642) );
  OR2_X1 U6647 ( .A1(n6643), .A2(n6644), .ZN(n6640) );
  AND2_X1 U6648 ( .A1(n6645), .A2(n6646), .ZN(n6644) );
  AND2_X1 U6649 ( .A1(n6647), .A2(n6648), .ZN(n6643) );
  INV_X1 U6650 ( .A(n6532), .ZN(n6627) );
  AND2_X1 U6651 ( .A1(a_12_), .A2(b_3_), .ZN(n6532) );
  OR2_X1 U6652 ( .A1(n6649), .A2(n6650), .ZN(n6538) );
  INV_X1 U6653 ( .A(n6651), .ZN(n6650) );
  OR2_X1 U6654 ( .A1(n6652), .A2(n6653), .ZN(n6651) );
  AND2_X1 U6655 ( .A1(n6653), .A2(n6652), .ZN(n6649) );
  AND2_X1 U6656 ( .A1(n6654), .A2(n6655), .ZN(n6652) );
  INV_X1 U6657 ( .A(n6656), .ZN(n6655) );
  AND2_X1 U6658 ( .A1(n6657), .A2(n6658), .ZN(n6656) );
  OR2_X1 U6659 ( .A1(n6658), .A2(n6657), .ZN(n6654) );
  OR2_X1 U6660 ( .A1(n6554), .A2(n6548), .ZN(n6620) );
  OR2_X1 U6661 ( .A1(n6659), .A2(n6660), .ZN(n6548) );
  INV_X1 U6662 ( .A(n6661), .ZN(n6660) );
  OR2_X1 U6663 ( .A1(n6662), .A2(n6663), .ZN(n6661) );
  AND2_X1 U6664 ( .A1(n6663), .A2(n6662), .ZN(n6659) );
  AND2_X1 U6665 ( .A1(n6664), .A2(n6665), .ZN(n6662) );
  INV_X1 U6666 ( .A(n6666), .ZN(n6665) );
  AND2_X1 U6667 ( .A1(n6667), .A2(n6668), .ZN(n6666) );
  OR2_X1 U6668 ( .A1(n6668), .A2(n6667), .ZN(n6664) );
  OR2_X1 U6669 ( .A1(n3964), .A2(n3867), .ZN(n6554) );
  INV_X1 U6670 ( .A(b_3_), .ZN(n3867) );
  AND2_X1 U6671 ( .A1(n6669), .A2(n6670), .ZN(n6559) );
  INV_X1 U6672 ( .A(n6671), .ZN(n6670) );
  AND2_X1 U6673 ( .A1(n6672), .A2(n6673), .ZN(n6671) );
  OR2_X1 U6674 ( .A1(n6673), .A2(n6672), .ZN(n6669) );
  OR2_X1 U6675 ( .A1(n6674), .A2(n6675), .ZN(n6672) );
  AND2_X1 U6676 ( .A1(n6676), .A2(n6677), .ZN(n6675) );
  INV_X1 U6677 ( .A(n6678), .ZN(n6674) );
  OR2_X1 U6678 ( .A1(n6677), .A2(n6676), .ZN(n6678) );
  INV_X1 U6679 ( .A(n6679), .ZN(n6676) );
  AND2_X1 U6680 ( .A1(n6680), .A2(n6681), .ZN(n6569) );
  INV_X1 U6681 ( .A(n6682), .ZN(n6681) );
  AND2_X1 U6682 ( .A1(n6683), .A2(n6684), .ZN(n6682) );
  OR2_X1 U6683 ( .A1(n6684), .A2(n6683), .ZN(n6680) );
  OR2_X1 U6684 ( .A1(n6685), .A2(n6686), .ZN(n6683) );
  AND2_X1 U6685 ( .A1(n6687), .A2(n6688), .ZN(n6686) );
  INV_X1 U6686 ( .A(n6689), .ZN(n6685) );
  OR2_X1 U6687 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  AND2_X1 U6688 ( .A1(n6690), .A2(n6691), .ZN(n6579) );
  INV_X1 U6689 ( .A(n6692), .ZN(n6691) );
  AND2_X1 U6690 ( .A1(n6693), .A2(n6694), .ZN(n6692) );
  OR2_X1 U6691 ( .A1(n6694), .A2(n6693), .ZN(n6690) );
  OR2_X1 U6692 ( .A1(n6695), .A2(n6696), .ZN(n6693) );
  AND2_X1 U6693 ( .A1(n6697), .A2(n6698), .ZN(n6696) );
  INV_X1 U6694 ( .A(n6699), .ZN(n6695) );
  OR2_X1 U6695 ( .A1(n6698), .A2(n6697), .ZN(n6699) );
  AND2_X1 U6696 ( .A1(n6700), .A2(n6701), .ZN(n6589) );
  INV_X1 U6697 ( .A(n6702), .ZN(n6701) );
  AND2_X1 U6698 ( .A1(n6703), .A2(n6704), .ZN(n6702) );
  OR2_X1 U6699 ( .A1(n6704), .A2(n6703), .ZN(n6700) );
  OR2_X1 U6700 ( .A1(n6705), .A2(n6706), .ZN(n6703) );
  AND2_X1 U6701 ( .A1(n6707), .A2(n6708), .ZN(n6706) );
  INV_X1 U6702 ( .A(n6709), .ZN(n6705) );
  OR2_X1 U6703 ( .A1(n6708), .A2(n6707), .ZN(n6709) );
  AND2_X1 U6704 ( .A1(n6710), .A2(n6711), .ZN(n4370) );
  INV_X1 U6705 ( .A(n6712), .ZN(n6711) );
  AND2_X1 U6706 ( .A1(n6713), .A2(n6714), .ZN(n6712) );
  OR2_X1 U6707 ( .A1(n6714), .A2(n6713), .ZN(n6710) );
  OR2_X1 U6708 ( .A1(n6715), .A2(n6716), .ZN(n6713) );
  AND2_X1 U6709 ( .A1(n6717), .A2(n6718), .ZN(n6716) );
  INV_X1 U6710 ( .A(n6719), .ZN(n6715) );
  OR2_X1 U6711 ( .A1(n6718), .A2(n6717), .ZN(n6719) );
  AND2_X1 U6712 ( .A1(n3846), .A2(n3847), .ZN(n3843) );
  INV_X1 U6713 ( .A(n6720), .ZN(n3847) );
  OR2_X1 U6714 ( .A1(n4038), .A2(n4039), .ZN(n6720) );
  OR2_X1 U6715 ( .A1(n6721), .A2(n6722), .ZN(n4039) );
  AND2_X1 U6716 ( .A1(n4064), .A2(n4062), .ZN(n6722) );
  AND2_X1 U6717 ( .A1(n4056), .A2(n6723), .ZN(n6721) );
  OR2_X1 U6718 ( .A1(n4062), .A2(n4064), .ZN(n6723) );
  OR2_X1 U6719 ( .A1(n6510), .A2(n3938), .ZN(n4064) );
  OR2_X1 U6720 ( .A1(n6724), .A2(n6725), .ZN(n4062) );
  AND2_X1 U6721 ( .A1(n6726), .A2(n4097), .ZN(n6725) );
  AND2_X1 U6722 ( .A1(n4093), .A2(n6727), .ZN(n6724) );
  OR2_X1 U6723 ( .A1(n4097), .A2(n6726), .ZN(n6727) );
  INV_X1 U6724 ( .A(n4096), .ZN(n6726) );
  AND2_X1 U6725 ( .A1(b_2_), .A2(a_1_), .ZN(n4096) );
  OR2_X1 U6726 ( .A1(n6728), .A2(n6729), .ZN(n4097) );
  AND2_X1 U6727 ( .A1(n3891), .A2(n4152), .ZN(n6729) );
  AND2_X1 U6728 ( .A1(n4147), .A2(n6730), .ZN(n6728) );
  OR2_X1 U6729 ( .A1(n4152), .A2(n3891), .ZN(n6730) );
  OR2_X1 U6730 ( .A1(n6510), .A2(n6731), .ZN(n3891) );
  OR2_X1 U6731 ( .A1(n6732), .A2(n6733), .ZN(n4152) );
  AND2_X1 U6732 ( .A1(n6734), .A2(n4211), .ZN(n6733) );
  AND2_X1 U6733 ( .A1(n4207), .A2(n6735), .ZN(n6732) );
  OR2_X1 U6734 ( .A1(n4211), .A2(n6734), .ZN(n6735) );
  INV_X1 U6735 ( .A(n4210), .ZN(n6734) );
  AND2_X1 U6736 ( .A1(b_2_), .A2(a_3_), .ZN(n4210) );
  OR2_X1 U6737 ( .A1(n6736), .A2(n6737), .ZN(n4211) );
  AND2_X1 U6738 ( .A1(n6738), .A2(n4293), .ZN(n6737) );
  AND2_X1 U6739 ( .A1(n4289), .A2(n6739), .ZN(n6736) );
  OR2_X1 U6740 ( .A1(n4293), .A2(n6738), .ZN(n6739) );
  INV_X1 U6741 ( .A(n4292), .ZN(n6738) );
  AND2_X1 U6742 ( .A1(b_2_), .A2(a_4_), .ZN(n4292) );
  OR2_X1 U6743 ( .A1(n6740), .A2(n6741), .ZN(n4293) );
  AND2_X1 U6744 ( .A1(n6742), .A2(n4381), .ZN(n6741) );
  AND2_X1 U6745 ( .A1(n4377), .A2(n6743), .ZN(n6740) );
  OR2_X1 U6746 ( .A1(n4381), .A2(n6742), .ZN(n6743) );
  INV_X1 U6747 ( .A(n4380), .ZN(n6742) );
  AND2_X1 U6748 ( .A1(b_2_), .A2(a_5_), .ZN(n4380) );
  OR2_X1 U6749 ( .A1(n6744), .A2(n6745), .ZN(n4381) );
  AND2_X1 U6750 ( .A1(n6746), .A2(n6718), .ZN(n6745) );
  AND2_X1 U6751 ( .A1(n6714), .A2(n6747), .ZN(n6744) );
  OR2_X1 U6752 ( .A1(n6718), .A2(n6746), .ZN(n6747) );
  INV_X1 U6753 ( .A(n6717), .ZN(n6746) );
  AND2_X1 U6754 ( .A1(b_2_), .A2(a_6_), .ZN(n6717) );
  OR2_X1 U6755 ( .A1(n6748), .A2(n6749), .ZN(n6718) );
  AND2_X1 U6756 ( .A1(n6750), .A2(n6708), .ZN(n6749) );
  AND2_X1 U6757 ( .A1(n6704), .A2(n6751), .ZN(n6748) );
  OR2_X1 U6758 ( .A1(n6708), .A2(n6750), .ZN(n6751) );
  INV_X1 U6759 ( .A(n6707), .ZN(n6750) );
  AND2_X1 U6760 ( .A1(a_7_), .A2(b_2_), .ZN(n6707) );
  OR2_X1 U6761 ( .A1(n6752), .A2(n6753), .ZN(n6708) );
  AND2_X1 U6762 ( .A1(n6754), .A2(n6698), .ZN(n6753) );
  AND2_X1 U6763 ( .A1(n6694), .A2(n6755), .ZN(n6752) );
  OR2_X1 U6764 ( .A1(n6698), .A2(n6754), .ZN(n6755) );
  INV_X1 U6765 ( .A(n6697), .ZN(n6754) );
  AND2_X1 U6766 ( .A1(a_8_), .A2(b_2_), .ZN(n6697) );
  OR2_X1 U6767 ( .A1(n6756), .A2(n6757), .ZN(n6698) );
  AND2_X1 U6768 ( .A1(n6758), .A2(n6688), .ZN(n6757) );
  AND2_X1 U6769 ( .A1(n6684), .A2(n6759), .ZN(n6756) );
  OR2_X1 U6770 ( .A1(n6688), .A2(n6758), .ZN(n6759) );
  INV_X1 U6771 ( .A(n6687), .ZN(n6758) );
  AND2_X1 U6772 ( .A1(a_9_), .A2(b_2_), .ZN(n6687) );
  OR2_X1 U6773 ( .A1(n6760), .A2(n6761), .ZN(n6688) );
  AND2_X1 U6774 ( .A1(n6679), .A2(n6677), .ZN(n6761) );
  AND2_X1 U6775 ( .A1(n6673), .A2(n6762), .ZN(n6760) );
  OR2_X1 U6776 ( .A1(n6677), .A2(n6679), .ZN(n6762) );
  OR2_X1 U6777 ( .A1(n3964), .A2(n6510), .ZN(n6679) );
  OR2_X1 U6778 ( .A1(n6763), .A2(n6764), .ZN(n6677) );
  AND2_X1 U6779 ( .A1(n6663), .A2(n6765), .ZN(n6764) );
  AND2_X1 U6780 ( .A1(n6766), .A2(n6668), .ZN(n6763) );
  OR2_X1 U6781 ( .A1(n6767), .A2(n6768), .ZN(n6668) );
  AND2_X1 U6782 ( .A1(n6769), .A2(n6658), .ZN(n6768) );
  AND2_X1 U6783 ( .A1(n6653), .A2(n6770), .ZN(n6767) );
  OR2_X1 U6784 ( .A1(n6658), .A2(n6769), .ZN(n6770) );
  INV_X1 U6785 ( .A(n6657), .ZN(n6769) );
  AND2_X1 U6786 ( .A1(a_12_), .A2(b_2_), .ZN(n6657) );
  OR2_X1 U6787 ( .A1(n6771), .A2(n6772), .ZN(n6658) );
  AND2_X1 U6788 ( .A1(n6641), .A2(n6646), .ZN(n6772) );
  AND2_X1 U6789 ( .A1(n6645), .A2(n6773), .ZN(n6771) );
  OR2_X1 U6790 ( .A1(n6646), .A2(n6641), .ZN(n6773) );
  OR2_X1 U6791 ( .A1(n3631), .A2(n6510), .ZN(n6641) );
  INV_X1 U6792 ( .A(b_2_), .ZN(n6510) );
  INV_X1 U6793 ( .A(n6647), .ZN(n6646) );
  AND3_X1 U6794 ( .A1(n3975), .A2(b_2_), .A3(b_1_), .ZN(n6647) );
  INV_X1 U6795 ( .A(n6648), .ZN(n6645) );
  OR2_X1 U6796 ( .A1(n6774), .A2(n6775), .ZN(n6648) );
  AND2_X1 U6797 ( .A1(b_1_), .A2(n6776), .ZN(n6775) );
  OR2_X1 U6798 ( .A1(n6777), .A2(n3592), .ZN(n6776) );
  AND2_X1 U6799 ( .A1(n3576), .A2(a_14_), .ZN(n3592) );
  INV_X1 U6800 ( .A(a_15_), .ZN(n3576) );
  AND2_X1 U6801 ( .A1(a_14_), .A2(n3939), .ZN(n6777) );
  AND2_X1 U6802 ( .A1(b_0_), .A2(n6778), .ZN(n6774) );
  OR2_X1 U6803 ( .A1(n6779), .A2(n3595), .ZN(n6778) );
  AND2_X1 U6804 ( .A1(n3587), .A2(a_15_), .ZN(n3595) );
  AND2_X1 U6805 ( .A1(a_15_), .A2(n3911), .ZN(n6779) );
  OR2_X1 U6806 ( .A1(n6780), .A2(n6781), .ZN(n6653) );
  INV_X1 U6807 ( .A(n6782), .ZN(n6781) );
  OR2_X1 U6808 ( .A1(n6783), .A2(n6784), .ZN(n6782) );
  AND2_X1 U6809 ( .A1(n6784), .A2(n6783), .ZN(n6780) );
  OR2_X1 U6810 ( .A1(n6785), .A2(n6786), .ZN(n6783) );
  AND3_X1 U6811 ( .A1(a_13_), .A2(n6787), .A3(b_1_), .ZN(n6786) );
  OR2_X1 U6812 ( .A1(n3587), .A2(n3939), .ZN(n6787) );
  INV_X1 U6813 ( .A(a_14_), .ZN(n3587) );
  AND3_X1 U6814 ( .A1(a_14_), .A2(n6788), .A3(b_0_), .ZN(n6785) );
  OR2_X1 U6815 ( .A1(n3631), .A2(n3911), .ZN(n6788) );
  INV_X1 U6816 ( .A(a_13_), .ZN(n3631) );
  OR2_X1 U6817 ( .A1(n6765), .A2(n6663), .ZN(n6766) );
  OR2_X1 U6818 ( .A1(n6789), .A2(n6790), .ZN(n6663) );
  AND2_X1 U6819 ( .A1(n6791), .A2(n6792), .ZN(n6790) );
  INV_X1 U6820 ( .A(n6793), .ZN(n6789) );
  OR2_X1 U6821 ( .A1(n6791), .A2(n6792), .ZN(n6793) );
  OR2_X1 U6822 ( .A1(n6794), .A2(n6795), .ZN(n6791) );
  AND2_X1 U6823 ( .A1(n6796), .A2(n6797), .ZN(n6795) );
  AND2_X1 U6824 ( .A1(n6798), .A2(n6799), .ZN(n6794) );
  INV_X1 U6825 ( .A(n6667), .ZN(n6765) );
  AND2_X1 U6826 ( .A1(a_11_), .A2(b_2_), .ZN(n6667) );
  AND2_X1 U6827 ( .A1(n6800), .A2(n6801), .ZN(n6673) );
  INV_X1 U6828 ( .A(n6802), .ZN(n6801) );
  AND2_X1 U6829 ( .A1(n6803), .A2(n6804), .ZN(n6802) );
  OR2_X1 U6830 ( .A1(n6803), .A2(n6804), .ZN(n6800) );
  OR2_X1 U6831 ( .A1(n6805), .A2(n6806), .ZN(n6803) );
  AND2_X1 U6832 ( .A1(n6807), .A2(n6808), .ZN(n6806) );
  INV_X1 U6833 ( .A(n6809), .ZN(n6807) );
  AND2_X1 U6834 ( .A1(n6810), .A2(n6809), .ZN(n6805) );
  INV_X1 U6835 ( .A(n6808), .ZN(n6810) );
  AND2_X1 U6836 ( .A1(n6811), .A2(n6812), .ZN(n6684) );
  INV_X1 U6837 ( .A(n6813), .ZN(n6812) );
  AND2_X1 U6838 ( .A1(n6814), .A2(n6815), .ZN(n6813) );
  OR2_X1 U6839 ( .A1(n6814), .A2(n6815), .ZN(n6811) );
  OR2_X1 U6840 ( .A1(n6816), .A2(n6817), .ZN(n6814) );
  AND2_X1 U6841 ( .A1(n6818), .A2(n6819), .ZN(n6817) );
  INV_X1 U6842 ( .A(n6820), .ZN(n6818) );
  AND2_X1 U6843 ( .A1(n6821), .A2(n6820), .ZN(n6816) );
  INV_X1 U6844 ( .A(n6819), .ZN(n6821) );
  AND2_X1 U6845 ( .A1(n6822), .A2(n6823), .ZN(n6694) );
  INV_X1 U6846 ( .A(n6824), .ZN(n6823) );
  AND2_X1 U6847 ( .A1(n6825), .A2(n6826), .ZN(n6824) );
  OR2_X1 U6848 ( .A1(n6825), .A2(n6826), .ZN(n6822) );
  OR2_X1 U6849 ( .A1(n6827), .A2(n6828), .ZN(n6825) );
  AND2_X1 U6850 ( .A1(n6829), .A2(n6830), .ZN(n6828) );
  INV_X1 U6851 ( .A(n6831), .ZN(n6829) );
  AND2_X1 U6852 ( .A1(n6832), .A2(n6831), .ZN(n6827) );
  INV_X1 U6853 ( .A(n6830), .ZN(n6832) );
  AND2_X1 U6854 ( .A1(n6833), .A2(n6834), .ZN(n6704) );
  INV_X1 U6855 ( .A(n6835), .ZN(n6834) );
  AND2_X1 U6856 ( .A1(n6836), .A2(n6837), .ZN(n6835) );
  OR2_X1 U6857 ( .A1(n6836), .A2(n6837), .ZN(n6833) );
  OR2_X1 U6858 ( .A1(n6838), .A2(n6839), .ZN(n6836) );
  AND2_X1 U6859 ( .A1(n6840), .A2(n6841), .ZN(n6839) );
  INV_X1 U6860 ( .A(n6842), .ZN(n6840) );
  AND2_X1 U6861 ( .A1(n6843), .A2(n6842), .ZN(n6838) );
  INV_X1 U6862 ( .A(n6841), .ZN(n6843) );
  AND2_X1 U6863 ( .A1(n6844), .A2(n6845), .ZN(n6714) );
  INV_X1 U6864 ( .A(n6846), .ZN(n6845) );
  AND2_X1 U6865 ( .A1(n6847), .A2(n6848), .ZN(n6846) );
  OR2_X1 U6866 ( .A1(n6847), .A2(n6848), .ZN(n6844) );
  OR2_X1 U6867 ( .A1(n6849), .A2(n6850), .ZN(n6847) );
  AND2_X1 U6868 ( .A1(n6851), .A2(n6852), .ZN(n6850) );
  INV_X1 U6869 ( .A(n6853), .ZN(n6851) );
  AND2_X1 U6870 ( .A1(n6854), .A2(n6853), .ZN(n6849) );
  INV_X1 U6871 ( .A(n6852), .ZN(n6854) );
  AND2_X1 U6872 ( .A1(n6855), .A2(n6856), .ZN(n4377) );
  INV_X1 U6873 ( .A(n6857), .ZN(n6856) );
  AND2_X1 U6874 ( .A1(n6858), .A2(n6859), .ZN(n6857) );
  OR2_X1 U6875 ( .A1(n6858), .A2(n6859), .ZN(n6855) );
  OR2_X1 U6876 ( .A1(n6860), .A2(n6861), .ZN(n6858) );
  AND2_X1 U6877 ( .A1(n6862), .A2(n6863), .ZN(n6861) );
  INV_X1 U6878 ( .A(n6864), .ZN(n6862) );
  AND2_X1 U6879 ( .A1(n6865), .A2(n6864), .ZN(n6860) );
  INV_X1 U6880 ( .A(n6863), .ZN(n6865) );
  AND2_X1 U6881 ( .A1(n6866), .A2(n6867), .ZN(n4289) );
  INV_X1 U6882 ( .A(n6868), .ZN(n6867) );
  AND2_X1 U6883 ( .A1(n6869), .A2(n6870), .ZN(n6868) );
  OR2_X1 U6884 ( .A1(n6869), .A2(n6870), .ZN(n6866) );
  OR2_X1 U6885 ( .A1(n6871), .A2(n6872), .ZN(n6869) );
  AND2_X1 U6886 ( .A1(n6873), .A2(n6874), .ZN(n6872) );
  INV_X1 U6887 ( .A(n6875), .ZN(n6873) );
  AND2_X1 U6888 ( .A1(n6876), .A2(n6875), .ZN(n6871) );
  INV_X1 U6889 ( .A(n6874), .ZN(n6876) );
  AND2_X1 U6890 ( .A1(n6877), .A2(n6878), .ZN(n4207) );
  INV_X1 U6891 ( .A(n6879), .ZN(n6878) );
  AND2_X1 U6892 ( .A1(n6880), .A2(n6881), .ZN(n6879) );
  OR2_X1 U6893 ( .A1(n6880), .A2(n6881), .ZN(n6877) );
  OR2_X1 U6894 ( .A1(n6882), .A2(n6883), .ZN(n6880) );
  AND2_X1 U6895 ( .A1(n6884), .A2(n6885), .ZN(n6883) );
  INV_X1 U6896 ( .A(n6886), .ZN(n6884) );
  AND2_X1 U6897 ( .A1(n6887), .A2(n6886), .ZN(n6882) );
  INV_X1 U6898 ( .A(n6885), .ZN(n6887) );
  AND2_X1 U6899 ( .A1(n6888), .A2(n6889), .ZN(n4147) );
  INV_X1 U6900 ( .A(n6890), .ZN(n6889) );
  AND2_X1 U6901 ( .A1(n6891), .A2(n6892), .ZN(n6890) );
  OR2_X1 U6902 ( .A1(n6891), .A2(n6892), .ZN(n6888) );
  OR2_X1 U6903 ( .A1(n6893), .A2(n6894), .ZN(n6891) );
  AND2_X1 U6904 ( .A1(n6895), .A2(n6896), .ZN(n6894) );
  INV_X1 U6905 ( .A(n6897), .ZN(n6895) );
  AND2_X1 U6906 ( .A1(n6898), .A2(n6897), .ZN(n6893) );
  INV_X1 U6907 ( .A(n6896), .ZN(n6898) );
  AND2_X1 U6908 ( .A1(n6899), .A2(n6900), .ZN(n4093) );
  INV_X1 U6909 ( .A(n6901), .ZN(n6900) );
  AND2_X1 U6910 ( .A1(n6902), .A2(n6903), .ZN(n6901) );
  OR2_X1 U6911 ( .A1(n6902), .A2(n6903), .ZN(n6899) );
  OR2_X1 U6912 ( .A1(n6904), .A2(n6905), .ZN(n6902) );
  AND2_X1 U6913 ( .A1(n6906), .A2(n6907), .ZN(n6905) );
  INV_X1 U6914 ( .A(n6908), .ZN(n6906) );
  AND2_X1 U6915 ( .A1(n6909), .A2(n6908), .ZN(n6904) );
  INV_X1 U6916 ( .A(n6907), .ZN(n6909) );
  AND2_X1 U6917 ( .A1(n6910), .A2(n6911), .ZN(n4056) );
  INV_X1 U6918 ( .A(n6912), .ZN(n6911) );
  AND2_X1 U6919 ( .A1(n6913), .A2(n6914), .ZN(n6912) );
  OR2_X1 U6920 ( .A1(n6913), .A2(n6914), .ZN(n6910) );
  OR2_X1 U6921 ( .A1(n6915), .A2(n6916), .ZN(n6913) );
  INV_X1 U6922 ( .A(n6917), .ZN(n6916) );
  OR2_X1 U6923 ( .A1(n6918), .A2(n3909), .ZN(n6917) );
  AND2_X1 U6924 ( .A1(n3909), .A2(n6918), .ZN(n6915) );
  AND2_X1 U6925 ( .A1(n6919), .A2(n6920), .ZN(n4038) );
  INV_X1 U6926 ( .A(n6921), .ZN(n6920) );
  AND2_X1 U6927 ( .A1(n6922), .A2(n6923), .ZN(n6921) );
  OR2_X1 U6928 ( .A1(n6922), .A2(n6923), .ZN(n6919) );
  OR2_X1 U6929 ( .A1(n6924), .A2(n6925), .ZN(n6922) );
  INV_X1 U6930 ( .A(n6926), .ZN(n6925) );
  OR2_X1 U6931 ( .A1(n6927), .A2(n6928), .ZN(n6926) );
  AND2_X1 U6932 ( .A1(n6928), .A2(n6927), .ZN(n6924) );
  INV_X1 U6933 ( .A(n6929), .ZN(n6928) );
  OR2_X1 U6934 ( .A1(n6930), .A2(n6931), .ZN(n3846) );
  AND2_X1 U6935 ( .A1(n6932), .A2(n6933), .ZN(n6931) );
  INV_X1 U6936 ( .A(n6934), .ZN(n6932) );
  AND2_X1 U6937 ( .A1(n4034), .A2(n6934), .ZN(n6930) );
  OR2_X1 U6938 ( .A1(n3939), .A2(n3938), .ZN(n6934) );
  INV_X1 U6939 ( .A(n6933), .ZN(n4034) );
  OR2_X1 U6940 ( .A1(n6935), .A2(n6936), .ZN(n6933) );
  AND2_X1 U6941 ( .A1(n6923), .A2(n6927), .ZN(n6936) );
  AND2_X1 U6942 ( .A1(n6937), .A2(n6929), .ZN(n6935) );
  OR2_X1 U6943 ( .A1(n3911), .A2(n3938), .ZN(n6929) );
  INV_X1 U6944 ( .A(a_0_), .ZN(n3938) );
  OR2_X1 U6945 ( .A1(n6927), .A2(n6923), .ZN(n6937) );
  OR2_X1 U6946 ( .A1(n3939), .A2(n3914), .ZN(n6923) );
  INV_X1 U6947 ( .A(a_1_), .ZN(n3914) );
  OR2_X1 U6948 ( .A1(n6938), .A2(n6939), .ZN(n6927) );
  AND2_X1 U6949 ( .A1(n6914), .A2(n6918), .ZN(n6939) );
  AND2_X1 U6950 ( .A1(n6940), .A2(n3942), .ZN(n6938) );
  INV_X1 U6951 ( .A(n3909), .ZN(n3942) );
  AND2_X1 U6952 ( .A1(b_1_), .A2(a_1_), .ZN(n3909) );
  OR2_X1 U6953 ( .A1(n6918), .A2(n6914), .ZN(n6940) );
  OR2_X1 U6954 ( .A1(n3939), .A2(n6731), .ZN(n6914) );
  OR2_X1 U6955 ( .A1(n6941), .A2(n6942), .ZN(n6918) );
  AND2_X1 U6956 ( .A1(n6903), .A2(n6908), .ZN(n6942) );
  AND2_X1 U6957 ( .A1(n6943), .A2(n6907), .ZN(n6941) );
  OR2_X1 U6958 ( .A1(n3939), .A2(n3870), .ZN(n6907) );
  OR2_X1 U6959 ( .A1(n6908), .A2(n6903), .ZN(n6943) );
  OR2_X1 U6960 ( .A1(n3911), .A2(n6731), .ZN(n6903) );
  INV_X1 U6961 ( .A(a_2_), .ZN(n6731) );
  OR2_X1 U6962 ( .A1(n6944), .A2(n6945), .ZN(n6908) );
  AND2_X1 U6963 ( .A1(n6892), .A2(n6897), .ZN(n6945) );
  AND2_X1 U6964 ( .A1(n6946), .A2(n6896), .ZN(n6944) );
  OR2_X1 U6965 ( .A1(n3939), .A2(n6471), .ZN(n6896) );
  OR2_X1 U6966 ( .A1(n6897), .A2(n6892), .ZN(n6946) );
  OR2_X1 U6967 ( .A1(n3911), .A2(n3870), .ZN(n6892) );
  INV_X1 U6968 ( .A(a_3_), .ZN(n3870) );
  OR2_X1 U6969 ( .A1(n6947), .A2(n6948), .ZN(n6897) );
  AND2_X1 U6970 ( .A1(n6881), .A2(n6886), .ZN(n6948) );
  AND2_X1 U6971 ( .A1(n6949), .A2(n6885), .ZN(n6947) );
  OR2_X1 U6972 ( .A1(n3815), .A2(n3939), .ZN(n6885) );
  OR2_X1 U6973 ( .A1(n6886), .A2(n6881), .ZN(n6949) );
  OR2_X1 U6974 ( .A1(n3911), .A2(n6471), .ZN(n6881) );
  INV_X1 U6975 ( .A(a_4_), .ZN(n6471) );
  OR2_X1 U6976 ( .A1(n6950), .A2(n6951), .ZN(n6886) );
  AND2_X1 U6977 ( .A1(n6870), .A2(n6875), .ZN(n6951) );
  AND2_X1 U6978 ( .A1(n6952), .A2(n6874), .ZN(n6950) );
  OR2_X1 U6979 ( .A1(n6187), .A2(n3939), .ZN(n6874) );
  OR2_X1 U6980 ( .A1(n6875), .A2(n6870), .ZN(n6952) );
  OR2_X1 U6981 ( .A1(n3911), .A2(n3815), .ZN(n6870) );
  INV_X1 U6982 ( .A(a_5_), .ZN(n3815) );
  OR2_X1 U6983 ( .A1(n6953), .A2(n6954), .ZN(n6875) );
  AND2_X1 U6984 ( .A1(n6859), .A2(n6864), .ZN(n6954) );
  AND2_X1 U6985 ( .A1(n6955), .A2(n6863), .ZN(n6953) );
  OR2_X1 U6986 ( .A1(n3771), .A2(n3939), .ZN(n6863) );
  OR2_X1 U6987 ( .A1(n6864), .A2(n6859), .ZN(n6955) );
  OR2_X1 U6988 ( .A1(n6187), .A2(n3911), .ZN(n6859) );
  INV_X1 U6989 ( .A(a_6_), .ZN(n6187) );
  OR2_X1 U6990 ( .A1(n6956), .A2(n6957), .ZN(n6864) );
  AND2_X1 U6991 ( .A1(n6848), .A2(n6853), .ZN(n6957) );
  AND2_X1 U6992 ( .A1(n6958), .A2(n6852), .ZN(n6956) );
  OR2_X1 U6993 ( .A1(n5925), .A2(n3939), .ZN(n6852) );
  OR2_X1 U6994 ( .A1(n6853), .A2(n6848), .ZN(n6958) );
  OR2_X1 U6995 ( .A1(n3771), .A2(n3911), .ZN(n6848) );
  INV_X1 U6996 ( .A(a_7_), .ZN(n3771) );
  OR2_X1 U6997 ( .A1(n6959), .A2(n6960), .ZN(n6853) );
  AND2_X1 U6998 ( .A1(n6837), .A2(n6842), .ZN(n6960) );
  AND2_X1 U6999 ( .A1(n6961), .A2(n6841), .ZN(n6959) );
  OR2_X1 U7000 ( .A1(n3727), .A2(n3939), .ZN(n6841) );
  OR2_X1 U7001 ( .A1(n6842), .A2(n6837), .ZN(n6961) );
  OR2_X1 U7002 ( .A1(n5925), .A2(n3911), .ZN(n6837) );
  INV_X1 U7003 ( .A(a_8_), .ZN(n5925) );
  OR2_X1 U7004 ( .A1(n6962), .A2(n6963), .ZN(n6842) );
  AND2_X1 U7005 ( .A1(n6826), .A2(n6831), .ZN(n6963) );
  AND2_X1 U7006 ( .A1(n6964), .A2(n6830), .ZN(n6962) );
  OR2_X1 U7007 ( .A1(n3964), .A2(n3939), .ZN(n6830) );
  OR2_X1 U7008 ( .A1(n6831), .A2(n6826), .ZN(n6964) );
  OR2_X1 U7009 ( .A1(n3727), .A2(n3911), .ZN(n6826) );
  INV_X1 U7010 ( .A(a_9_), .ZN(n3727) );
  OR2_X1 U7011 ( .A1(n6965), .A2(n6966), .ZN(n6831) );
  AND2_X1 U7012 ( .A1(n6815), .A2(n6820), .ZN(n6966) );
  AND2_X1 U7013 ( .A1(n6967), .A2(n6819), .ZN(n6965) );
  OR2_X1 U7014 ( .A1(n3681), .A2(n3939), .ZN(n6819) );
  OR2_X1 U7015 ( .A1(n6820), .A2(n6815), .ZN(n6967) );
  OR2_X1 U7016 ( .A1(n3964), .A2(n3911), .ZN(n6815) );
  INV_X1 U7017 ( .A(a_10_), .ZN(n3964) );
  OR2_X1 U7018 ( .A1(n6968), .A2(n6969), .ZN(n6820) );
  AND2_X1 U7019 ( .A1(n6804), .A2(n6809), .ZN(n6969) );
  AND2_X1 U7020 ( .A1(n6970), .A2(n6808), .ZN(n6968) );
  OR2_X1 U7021 ( .A1(n6971), .A2(n3939), .ZN(n6808) );
  INV_X1 U7022 ( .A(b_0_), .ZN(n3939) );
  OR2_X1 U7023 ( .A1(n6809), .A2(n6804), .ZN(n6970) );
  OR2_X1 U7024 ( .A1(n3681), .A2(n3911), .ZN(n6804) );
  INV_X1 U7025 ( .A(a_11_), .ZN(n3681) );
  OR2_X1 U7026 ( .A1(n6972), .A2(n6973), .ZN(n6809) );
  AND2_X1 U7027 ( .A1(n6792), .A2(n6797), .ZN(n6973) );
  AND2_X1 U7028 ( .A1(n6796), .A2(n6974), .ZN(n6972) );
  OR2_X1 U7029 ( .A1(n6797), .A2(n6792), .ZN(n6974) );
  OR2_X1 U7030 ( .A1(n6971), .A2(n3911), .ZN(n6792) );
  INV_X1 U7031 ( .A(b_1_), .ZN(n3911) );
  INV_X1 U7032 ( .A(a_12_), .ZN(n6971) );
  INV_X1 U7033 ( .A(n6798), .ZN(n6797) );
  INV_X1 U7034 ( .A(n6799), .ZN(n6796) );
  OR2_X1 U7035 ( .A1(n6975), .A2(n6784), .ZN(n6799) );
  AND3_X1 U7036 ( .A1(n3975), .A2(b_1_), .A3(b_0_), .ZN(n6784) );
  AND2_X1 U7037 ( .A1(a_15_), .A2(a_14_), .ZN(n3975) );
  AND3_X1 U7038 ( .A1(b_1_), .A2(a_14_), .A3(n6798), .ZN(n6975) );
  AND2_X1 U7039 ( .A1(a_13_), .A2(b_0_), .ZN(n6798) );
endmodule

