module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n155_, new_n384_, new_n410_, new_n445_, new_n236_, new_n238_, new_n92_, new_n79_, new_n250_, new_n113_, new_n288_, new_n371_, new_n97_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n76_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n291_, new_n261_, new_n241_, new_n309_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n82_, new_n401_, new_n389_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n170_, new_n246_, new_n400_, new_n328_, new_n266_, new_n367_, new_n173_, new_n220_, new_n130_, new_n419_, new_n268_, new_n374_, new_n376_, new_n380_, new_n214_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n352_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n126_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n317_, new_n102_, new_n344_, new_n143_, new_n287_, new_n125_, new_n145_, new_n253_, new_n403_, new_n90_, new_n237_, new_n427_, new_n234_, new_n149_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n292_, new_n106_, new_n411_, new_n215_, new_n152_, new_n157_, new_n107_, new_n93_, new_n182_, new_n153_, new_n407_, new_n81_, new_n133_, new_n257_, new_n212_, new_n151_, new_n364_, new_n449_, new_n219_, new_n231_, new_n313_, new_n78_, new_n239_, new_n382_, new_n272_, new_n282_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n146_, new_n88_, new_n360_, new_n98_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n326_, new_n95_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n87_, new_n387_, new_n103_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n174_, new_n297_, new_n361_, new_n150_, new_n354_, new_n392_, new_n444_, new_n108_, new_n137_, new_n183_, new_n303_, new_n105_, new_n340_, new_n147_, new_n285_, new_n80_, new_n351_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n325_, new_n417_, new_n180_, new_n332_, new_n318_, new_n163_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n111_, new_n158_, new_n252_, new_n262_, new_n160_, new_n312_, new_n271_, new_n274_, new_n100_, new_n242_, new_n218_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n408_, new_n423_, new_n205_, new_n213_, new_n134_, new_n141_, new_n433_, new_n435_, new_n206_, new_n109_, new_n254_, new_n355_, new_n353_, new_n85_, new_n265_, new_n370_, new_n256_, new_n278_, new_n304_, new_n381_, new_n388_, new_n217_, new_n101_, new_n269_, new_n194_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n412_, new_n165_, new_n441_, new_n327_, new_n216_, new_n431_, new_n77_, new_n196_, new_n280_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n338_, new_n383_, new_n343_, new_n210_, new_n447_, new_n207_, new_n267_, new_n336_, new_n140_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n311_, new_n86_, new_n84_, new_n195_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n277_, new_n245_, new_n402_, new_n89_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n91_, new_n346_, new_n396_, new_n198_, new_n438_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n83_, new_n322_, new_n228_, new_n289_, new_n179_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n104_, new_n185_, new_n399_, new_n373_, new_n171_, new_n434_, new_n200_, new_n422_, new_n99_, new_n329_, new_n249_, new_n233_, new_n136_, new_n284_, new_n119_, new_n293_, new_n391_, new_n96_, new_n178_, new_n437_, new_n168_, new_n279_, new_n295_, new_n359_, new_n132_, new_n120_, new_n166_, new_n162_, new_n409_, new_n161_, new_n406_, new_n356_, new_n333_, new_n229_, new_n290_, new_n94_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n276_, new_n405_;

not g000 ( new_n76_, keyIn_0_10 );
not g001 ( new_n77_, N11 );
and g002 ( new_n78_, new_n77_, keyIn_0_1 );
not g003 ( new_n79_, keyIn_0_1 );
and g004 ( new_n80_, new_n79_, N11 );
or g005 ( new_n81_, new_n78_, new_n80_ );
and g006 ( new_n82_, new_n81_, N17 );
or g007 ( new_n83_, new_n82_, new_n76_ );
not g008 ( new_n84_, N17 );
not g009 ( new_n85_, new_n81_ );
or g010 ( new_n86_, new_n85_, keyIn_0_10, new_n84_ );
and g011 ( new_n87_, new_n83_, new_n86_ );
not g012 ( new_n88_, keyIn_0_13 );
and g013 ( new_n89_, keyIn_0_4, N50 );
not g014 ( new_n90_, keyIn_0_4 );
not g015 ( new_n91_, N50 );
and g016 ( new_n92_, new_n90_, new_n91_ );
or g017 ( new_n93_, new_n92_, new_n89_ );
and g018 ( new_n94_, new_n93_, N56 );
or g019 ( new_n95_, new_n94_, new_n88_ );
not g020 ( new_n96_, N56 );
not g021 ( new_n97_, new_n93_ );
or g022 ( new_n98_, new_n97_, keyIn_0_13, new_n96_ );
and g023 ( new_n99_, new_n95_, new_n98_ );
not g024 ( new_n100_, keyIn_0_14 );
not g025 ( new_n101_, N63 );
and g026 ( new_n102_, new_n101_, keyIn_0_5 );
not g027 ( new_n103_, new_n102_ );
or g028 ( new_n104_, new_n101_, keyIn_0_5 );
and g029 ( new_n105_, new_n103_, new_n104_, N69 );
or g030 ( new_n106_, new_n105_, new_n100_ );
not g031 ( new_n107_, N69 );
not g032 ( new_n108_, new_n104_ );
or g033 ( new_n109_, new_n108_, keyIn_0_14, new_n107_, new_n102_ );
and g034 ( new_n110_, new_n106_, new_n109_ );
and g035 ( new_n111_, new_n87_, new_n99_, new_n110_ );
not g036 ( new_n112_, keyIn_0_11 );
not g037 ( new_n113_, N24 );
and g038 ( new_n114_, new_n113_, keyIn_0_2 );
not g039 ( new_n115_, new_n114_ );
or g040 ( new_n116_, new_n113_, keyIn_0_2 );
and g041 ( new_n117_, new_n115_, new_n116_, N30 );
or g042 ( new_n118_, new_n117_, new_n112_ );
not g043 ( new_n119_, N30 );
not g044 ( new_n120_, new_n116_ );
or g045 ( new_n121_, new_n120_, keyIn_0_11, new_n119_, new_n114_ );
and g046 ( new_n122_, new_n118_, new_n121_ );
not g047 ( new_n123_, N95 );
and g048 ( new_n124_, keyIn_0_7, N89 );
not g049 ( new_n125_, new_n124_ );
or g050 ( new_n126_, keyIn_0_7, N89 );
and g051 ( new_n127_, new_n125_, new_n126_ );
or g052 ( new_n128_, new_n127_, new_n123_ );
and g053 ( new_n129_, new_n128_, keyIn_0_16 );
not g054 ( new_n130_, keyIn_0_16 );
not g055 ( new_n131_, new_n127_ );
and g056 ( new_n132_, new_n131_, new_n130_, N95 );
or g057 ( new_n133_, new_n129_, new_n132_ );
and g058 ( new_n134_, new_n133_, new_n122_ );
not g059 ( new_n135_, keyIn_0_17 );
not g060 ( new_n136_, N108 );
or g061 ( new_n137_, keyIn_0_8, N102 );
not g062 ( new_n138_, new_n137_ );
and g063 ( new_n139_, keyIn_0_8, N102 );
or g064 ( new_n140_, new_n138_, new_n136_, new_n139_ );
and g065 ( new_n141_, new_n140_, new_n135_ );
not g066 ( new_n142_, new_n139_ );
and g067 ( new_n143_, new_n142_, keyIn_0_17, N108, new_n137_ );
or g068 ( new_n144_, new_n141_, new_n143_ );
not g069 ( new_n145_, keyIn_0_0 );
and g070 ( new_n146_, new_n145_, N1 );
not g071 ( new_n147_, N1 );
and g072 ( new_n148_, new_n147_, keyIn_0_0 );
or g073 ( new_n149_, new_n146_, new_n148_ );
and g074 ( new_n150_, new_n149_, N4 );
or g075 ( new_n151_, new_n150_, keyIn_0_9 );
not g076 ( new_n152_, keyIn_0_9 );
not g077 ( new_n153_, N4 );
not g078 ( new_n154_, new_n149_ );
or g079 ( new_n155_, new_n154_, new_n152_, new_n153_ );
and g080 ( new_n156_, new_n151_, new_n155_ );
and g081 ( new_n157_, new_n156_, new_n144_ );
not g082 ( new_n158_, keyIn_0_12 );
and g083 ( new_n159_, keyIn_0_3, N37 );
not g084 ( new_n160_, keyIn_0_3 );
not g085 ( new_n161_, N37 );
and g086 ( new_n162_, new_n160_, new_n161_ );
or g087 ( new_n163_, new_n162_, new_n159_ );
and g088 ( new_n164_, new_n163_, N43 );
or g089 ( new_n165_, new_n164_, new_n158_ );
not g090 ( new_n166_, N43 );
not g091 ( new_n167_, new_n163_ );
or g092 ( new_n168_, new_n167_, keyIn_0_12, new_n166_ );
and g093 ( new_n169_, new_n165_, new_n168_ );
or g094 ( new_n170_, keyIn_0_6, N76 );
and g095 ( new_n171_, keyIn_0_6, N76 );
not g096 ( new_n172_, new_n171_ );
and g097 ( new_n173_, new_n172_, N82, new_n170_ );
or g098 ( new_n174_, new_n173_, keyIn_0_15 );
not g099 ( new_n175_, keyIn_0_15 );
not g100 ( new_n176_, N82 );
not g101 ( new_n177_, new_n170_ );
or g102 ( new_n178_, new_n177_, new_n171_, new_n175_, new_n176_ );
and g103 ( new_n179_, new_n174_, new_n178_ );
and g104 ( new_n180_, new_n169_, new_n179_ );
and g105 ( new_n181_, new_n111_, new_n134_, new_n157_, new_n180_ );
not g106 ( new_n182_, new_n181_ );
and g107 ( new_n183_, new_n182_, keyIn_0_18 );
not g108 ( new_n184_, keyIn_0_18 );
and g109 ( new_n185_, new_n156_, new_n169_, new_n144_, new_n179_ );
and g110 ( new_n186_, new_n185_, new_n184_, new_n111_, new_n134_ );
or g111 ( N223, new_n183_, new_n186_ );
not g112 ( new_n188_, keyIn_0_29 );
not g113 ( new_n189_, keyIn_0_26 );
not g114 ( new_n190_, new_n179_ );
not g115 ( new_n191_, keyIn_0_19 );
and g116 ( new_n192_, N223, new_n191_ );
or g117 ( new_n193_, new_n181_, new_n184_ );
not g118 ( new_n194_, new_n186_ );
and g119 ( new_n195_, new_n193_, keyIn_0_19, new_n194_ );
or g120 ( new_n196_, new_n192_, new_n195_ );
and g121 ( new_n197_, new_n196_, new_n190_ );
and g122 ( new_n198_, new_n193_, new_n194_ );
or g123 ( new_n199_, new_n198_, keyIn_0_19 );
not g124 ( new_n200_, new_n195_ );
and g125 ( new_n201_, new_n199_, new_n200_ );
and g126 ( new_n202_, new_n201_, new_n179_ );
or g127 ( new_n203_, new_n197_, new_n202_ );
and g128 ( new_n204_, new_n203_, new_n189_ );
or g129 ( new_n205_, new_n201_, new_n179_ );
not g130 ( new_n206_, new_n202_ );
and g131 ( new_n207_, new_n206_, keyIn_0_26, new_n205_ );
or g132 ( new_n208_, new_n204_, new_n176_, N86, new_n207_ );
not g133 ( new_n209_, keyIn_0_25 );
or g134 ( new_n210_, new_n201_, new_n110_ );
not g135 ( new_n211_, new_n210_ );
and g136 ( new_n212_, new_n199_, new_n110_, new_n200_ );
or g137 ( new_n213_, new_n211_, new_n212_ );
and g138 ( new_n214_, new_n213_, new_n209_ );
not g139 ( new_n215_, new_n212_ );
and g140 ( new_n216_, new_n210_, keyIn_0_25, new_n215_ );
or g141 ( new_n217_, new_n216_, N73 );
or g142 ( new_n218_, new_n214_, new_n217_, new_n107_ );
not g143 ( new_n219_, new_n99_ );
and g144 ( new_n220_, new_n196_, new_n219_ );
and g145 ( new_n221_, new_n199_, new_n99_, new_n200_ );
or g146 ( new_n222_, new_n220_, new_n221_ );
and g147 ( new_n223_, new_n222_, keyIn_0_24 );
not g148 ( new_n224_, keyIn_0_24 );
or g149 ( new_n225_, new_n201_, new_n99_ );
not g150 ( new_n226_, new_n221_ );
and g151 ( new_n227_, new_n225_, new_n224_, new_n226_ );
or g152 ( new_n228_, new_n227_, N60 );
or g153 ( new_n229_, new_n223_, new_n228_, new_n96_ );
not g154 ( new_n230_, new_n169_ );
and g155 ( new_n231_, new_n196_, new_n230_ );
and g156 ( new_n232_, new_n199_, new_n169_, new_n200_ );
or g157 ( new_n233_, new_n231_, new_n232_ );
and g158 ( new_n234_, new_n233_, keyIn_0_23 );
not g159 ( new_n235_, keyIn_0_23 );
or g160 ( new_n236_, new_n201_, new_n169_ );
not g161 ( new_n237_, new_n232_ );
and g162 ( new_n238_, new_n236_, new_n235_, new_n237_ );
or g163 ( new_n239_, new_n238_, N47 );
or g164 ( new_n240_, new_n234_, new_n239_, new_n166_ );
and g165 ( new_n241_, new_n208_, new_n218_, new_n229_, new_n240_ );
not g166 ( new_n242_, keyIn_0_27 );
or g167 ( new_n243_, new_n201_, new_n133_ );
and g168 ( new_n244_, new_n201_, new_n133_ );
not g169 ( new_n245_, new_n244_ );
and g170 ( new_n246_, new_n245_, new_n243_ );
or g171 ( new_n247_, new_n246_, new_n242_ );
and g172 ( new_n248_, new_n246_, new_n242_ );
not g173 ( new_n249_, new_n248_ );
and g174 ( new_n250_, new_n249_, new_n247_ );
or g175 ( new_n251_, new_n250_, new_n123_, N99 );
or g176 ( new_n252_, new_n201_, new_n87_ );
not g177 ( new_n253_, new_n252_ );
and g178 ( new_n254_, new_n199_, new_n87_, new_n200_ );
or g179 ( new_n255_, new_n253_, new_n254_ );
and g180 ( new_n256_, new_n255_, keyIn_0_21 );
not g181 ( new_n257_, keyIn_0_21 );
not g182 ( new_n258_, new_n254_ );
and g183 ( new_n259_, new_n252_, new_n257_, new_n258_ );
or g184 ( new_n260_, new_n259_, N21 );
or g185 ( new_n261_, new_n256_, new_n260_, new_n84_ );
not g186 ( new_n262_, keyIn_0_20 );
not g187 ( new_n263_, new_n156_ );
and g188 ( new_n264_, new_n196_, new_n263_ );
and g189 ( new_n265_, new_n199_, new_n156_, new_n200_ );
or g190 ( new_n266_, new_n264_, new_n265_ );
and g191 ( new_n267_, new_n266_, new_n262_ );
or g192 ( new_n268_, new_n201_, new_n156_ );
not g193 ( new_n269_, new_n265_ );
and g194 ( new_n270_, new_n268_, keyIn_0_20, new_n269_ );
or g195 ( new_n271_, new_n270_, N8 );
or g196 ( new_n272_, new_n267_, new_n271_, new_n153_ );
not g197 ( new_n273_, new_n122_ );
and g198 ( new_n274_, new_n196_, new_n273_ );
and g199 ( new_n275_, new_n199_, new_n122_, new_n200_ );
or g200 ( new_n276_, new_n274_, new_n275_ );
and g201 ( new_n277_, new_n276_, keyIn_0_22 );
not g202 ( new_n278_, keyIn_0_22 );
or g203 ( new_n279_, new_n201_, new_n122_ );
not g204 ( new_n280_, new_n275_ );
and g205 ( new_n281_, new_n279_, new_n278_, new_n280_ );
or g206 ( new_n282_, new_n281_, N34 );
or g207 ( new_n283_, new_n277_, new_n282_, new_n119_ );
not g208 ( new_n284_, new_n144_ );
and g209 ( new_n285_, new_n196_, new_n284_ );
and g210 ( new_n286_, new_n199_, new_n144_, new_n200_ );
or g211 ( new_n287_, new_n285_, new_n286_ );
and g212 ( new_n288_, new_n287_, keyIn_0_28 );
not g213 ( new_n289_, keyIn_0_28 );
or g214 ( new_n290_, new_n201_, new_n144_ );
not g215 ( new_n291_, new_n286_ );
and g216 ( new_n292_, new_n290_, new_n289_, new_n291_ );
or g217 ( new_n293_, new_n292_, N112 );
or g218 ( new_n294_, new_n288_, new_n293_, new_n136_ );
and g219 ( new_n295_, new_n261_, new_n272_, new_n283_, new_n294_ );
and g220 ( new_n296_, new_n241_, new_n295_, new_n251_ );
or g221 ( new_n297_, new_n296_, new_n188_ );
and g222 ( new_n298_, new_n241_, new_n295_, new_n188_, new_n251_ );
not g223 ( new_n299_, new_n298_ );
and g224 ( N329, new_n297_, new_n299_ );
not g225 ( new_n301_, new_n261_ );
or g226 ( new_n302_, N329, new_n301_ );
and g227 ( new_n303_, new_n297_, new_n301_, new_n299_ );
not g228 ( new_n304_, new_n303_ );
and g229 ( new_n305_, new_n302_, new_n304_ );
or g230 ( new_n306_, new_n256_, new_n84_, N27, new_n259_ );
or g231 ( new_n307_, new_n305_, new_n306_ );
not g232 ( new_n308_, new_n294_ );
or g233 ( new_n309_, N329, new_n308_ );
and g234 ( new_n310_, new_n297_, new_n308_, new_n299_ );
not g235 ( new_n311_, new_n310_ );
and g236 ( new_n312_, new_n309_, new_n311_ );
or g237 ( new_n313_, new_n288_, new_n136_, N115, new_n292_ );
or g238 ( new_n314_, new_n312_, new_n313_ );
not g239 ( new_n315_, new_n283_ );
or g240 ( new_n316_, N329, new_n315_ );
and g241 ( new_n317_, new_n297_, new_n315_, new_n299_ );
not g242 ( new_n318_, new_n317_ );
and g243 ( new_n319_, new_n316_, new_n318_ );
or g244 ( new_n320_, new_n277_, new_n119_, N40, new_n281_ );
or g245 ( new_n321_, new_n319_, new_n320_ );
and g246 ( new_n322_, new_n307_, new_n314_, new_n321_ );
not g247 ( new_n323_, new_n240_ );
or g248 ( new_n324_, N329, new_n323_ );
and g249 ( new_n325_, new_n297_, new_n323_, new_n299_ );
not g250 ( new_n326_, new_n325_ );
and g251 ( new_n327_, new_n324_, new_n326_ );
or g252 ( new_n328_, new_n234_, new_n166_, N53, new_n238_ );
or g253 ( new_n329_, new_n327_, new_n328_ );
not g254 ( new_n330_, new_n229_ );
or g255 ( new_n331_, N329, new_n330_ );
or g256 ( new_n332_, new_n229_, keyIn_0_29 );
and g257 ( new_n333_, new_n331_, new_n332_ );
or g258 ( new_n334_, new_n223_, new_n96_, N66, new_n227_ );
or g259 ( new_n335_, new_n333_, new_n334_ );
and g260 ( new_n336_, new_n329_, new_n335_ );
not g261 ( new_n337_, new_n218_ );
or g262 ( new_n338_, N329, new_n337_ );
and g263 ( new_n339_, new_n297_, new_n337_, new_n299_ );
not g264 ( new_n340_, new_n339_ );
and g265 ( new_n341_, new_n338_, new_n340_ );
or g266 ( new_n342_, new_n214_, new_n107_, N79, new_n216_ );
or g267 ( new_n343_, new_n341_, new_n342_ );
not g268 ( new_n344_, new_n251_ );
or g269 ( new_n345_, N329, new_n344_ );
and g270 ( new_n346_, new_n297_, new_n344_, new_n299_ );
not g271 ( new_n347_, new_n346_ );
and g272 ( new_n348_, new_n345_, new_n347_ );
or g273 ( new_n349_, new_n250_, new_n123_, N105 );
or g274 ( new_n350_, new_n348_, new_n349_ );
and g275 ( new_n351_, new_n343_, new_n350_ );
not g276 ( new_n352_, new_n208_ );
or g277 ( new_n353_, N329, new_n352_ );
and g278 ( new_n354_, new_n297_, new_n352_, new_n299_ );
not g279 ( new_n355_, new_n354_ );
and g280 ( new_n356_, new_n353_, new_n355_ );
or g281 ( new_n357_, new_n204_, new_n176_, N92, new_n207_ );
or g282 ( new_n358_, new_n356_, new_n357_ );
not g283 ( new_n359_, new_n272_ );
or g284 ( new_n360_, N329, new_n359_ );
and g285 ( new_n361_, new_n297_, new_n359_, new_n299_ );
not g286 ( new_n362_, new_n361_ );
and g287 ( new_n363_, new_n360_, new_n362_ );
or g288 ( new_n364_, new_n267_, new_n153_, N14, new_n270_ );
or g289 ( new_n365_, new_n363_, new_n364_ );
and g290 ( new_n366_, new_n358_, new_n365_ );
and g291 ( new_n367_, new_n322_, new_n336_, new_n351_, new_n366_ );
not g292 ( new_n368_, new_n367_ );
and g293 ( new_n369_, new_n368_, keyIn_0_30 );
not g294 ( new_n370_, keyIn_0_30 );
and g295 ( new_n371_, new_n367_, new_n370_ );
or g296 ( N370, new_n369_, new_n371_ );
and g297 ( new_n373_, N370, N27 );
and g298 ( new_n374_, N329, N21 );
and g299 ( new_n375_, N223, N11 );
or g300 ( new_n376_, new_n374_, new_n84_, new_n375_ );
or g301 ( new_n377_, new_n373_, new_n376_ );
and g302 ( new_n378_, N370, N40 );
and g303 ( new_n379_, N329, N34 );
and g304 ( new_n380_, N223, N24 );
or g305 ( new_n381_, new_n379_, new_n119_, new_n380_ );
or g306 ( new_n382_, new_n378_, new_n381_ );
and g307 ( new_n383_, new_n377_, new_n382_ );
and g308 ( new_n384_, N370, N66 );
and g309 ( new_n385_, N329, N60 );
and g310 ( new_n386_, N223, N50 );
or g311 ( new_n387_, new_n385_, new_n96_, new_n386_ );
or g312 ( new_n388_, new_n384_, new_n387_ );
and g313 ( new_n389_, N370, N53 );
and g314 ( new_n390_, N329, N47 );
and g315 ( new_n391_, N223, N37 );
or g316 ( new_n392_, new_n390_, new_n166_, new_n391_ );
or g317 ( new_n393_, new_n389_, new_n392_ );
and g318 ( new_n394_, new_n388_, new_n393_ );
and g319 ( new_n395_, N370, N79 );
and g320 ( new_n396_, N329, N73 );
and g321 ( new_n397_, N223, N63 );
or g322 ( new_n398_, new_n396_, new_n107_, new_n397_ );
or g323 ( new_n399_, new_n395_, new_n398_ );
and g324 ( new_n400_, N370, N92 );
and g325 ( new_n401_, N329, N86 );
and g326 ( new_n402_, N223, N76 );
or g327 ( new_n403_, new_n401_, new_n176_, new_n402_ );
or g328 ( new_n404_, new_n400_, new_n403_ );
and g329 ( new_n405_, N370, N105 );
and g330 ( new_n406_, N329, N99 );
and g331 ( new_n407_, N223, N89 );
or g332 ( new_n408_, new_n406_, new_n123_, new_n407_ );
or g333 ( new_n409_, new_n405_, new_n408_ );
and g334 ( new_n410_, N370, N115 );
and g335 ( new_n411_, N329, N112 );
and g336 ( new_n412_, N223, N102 );
or g337 ( new_n413_, new_n411_, new_n136_, new_n412_ );
or g338 ( new_n414_, new_n410_, new_n413_ );
and g339 ( new_n415_, new_n399_, new_n404_, new_n409_, new_n414_ );
and g340 ( new_n416_, new_n415_, keyIn_0_31, new_n383_, new_n394_ );
not g341 ( new_n417_, new_n416_ );
and g342 ( new_n418_, N370, N14 );
and g343 ( new_n419_, N329, N8 );
and g344 ( new_n420_, N223, N1 );
or g345 ( new_n421_, new_n418_, new_n153_, new_n419_, new_n420_ );
and g346 ( new_n422_, new_n399_, new_n404_ );
and g347 ( new_n423_, new_n409_, new_n414_ );
and g348 ( new_n424_, new_n383_, new_n394_, new_n422_, new_n423_ );
or g349 ( new_n425_, new_n424_, keyIn_0_31 );
and g350 ( N421, new_n425_, new_n417_, new_n421_ );
not g351 ( new_n427_, new_n383_ );
not g352 ( new_n428_, new_n394_ );
or g353 ( N430, new_n427_, new_n428_ );
not g354 ( new_n430_, new_n422_ );
and g355 ( new_n431_, new_n430_, new_n394_ );
or g356 ( N431, new_n431_, new_n427_ );
not g357 ( new_n433_, new_n377_ );
not g358 ( new_n434_, new_n393_ );
not g359 ( new_n435_, N79 );
or g360 ( new_n436_, new_n367_, new_n370_ );
not g361 ( new_n437_, new_n371_ );
and g362 ( new_n438_, new_n437_, new_n436_ );
or g363 ( new_n439_, new_n438_, new_n435_ );
not g364 ( new_n440_, new_n396_ );
not g365 ( new_n441_, new_n397_ );
and g366 ( new_n442_, new_n440_, N69, new_n441_ );
and g367 ( new_n443_, new_n388_, new_n439_, new_n442_ );
not g368 ( new_n444_, N105 );
or g369 ( new_n445_, new_n438_, new_n444_ );
not g370 ( new_n446_, new_n408_ );
and g371 ( new_n447_, new_n445_, new_n446_ );
and g372 ( new_n448_, new_n404_, new_n447_ );
or g373 ( new_n449_, new_n443_, new_n448_, new_n434_ );
and g374 ( new_n450_, new_n449_, new_n382_ );
or g375 ( N432, new_n450_, new_n433_ );
endmodule