module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n456_, new_n246_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n342_, new_n462_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n157_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n478_, new_n461_, new_n297_, new_n361_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n530_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n314_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n436_, new_n397_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n384_, new_n410_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n416_, new_n222_, new_n400_, new_n328_, new_n505_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n485_, new_n525_, new_n177_, new_n493_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n520_, new_n253_, new_n403_, new_n237_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n407_, new_n480_, new_n151_, new_n513_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n522_, new_n428_, new_n199_, new_n487_, new_n360_, new_n302_, new_n191_, new_n225_, new_n387_, new_n476_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n340_, new_n285_, new_n502_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n515_, new_n332_, new_n453_, new_n516_, new_n519_, new_n440_, new_n531_, new_n252_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n278_, new_n304_, new_n523_, new_n217_, new_n269_, new_n512_, new_n412_, new_n327_, new_n495_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n358_, new_n348_, new_n322_, new_n228_, new_n425_, new_n175_, new_n226_, new_n373_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n284_, new_n293_, new_n168_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n405_;

nand g000 ( new_n151_, N29, N42, N75 );
xor g001 ( N388, new_n151_, keyIn_0_3 );
and g002 ( N389, N29, N36, N80 );
nand g003 ( new_n154_, N29, N36, N42 );
xnor g004 ( N390, new_n154_, keyIn_0_4 );
and g005 ( N391, N85, N86 );
and g006 ( new_n157_, N1, N8 );
nand g007 ( new_n158_, new_n157_, N13, N17 );
xnor g008 ( N418, new_n158_, keyIn_0_0 );
xor g009 ( new_n160_, new_n154_, keyIn_0_1 );
not g010 ( new_n161_, new_n160_ );
and g011 ( new_n162_, N1, N13, N17, N26 );
nand g012 ( N419, new_n161_, new_n162_ );
nand g013 ( N420, N59, N75, N80 );
nand g014 ( N421, N36, N59, N80 );
nand g015 ( new_n166_, N36, N42, N59 );
xor g016 ( N422, new_n166_, keyIn_0_5 );
not g017 ( new_n168_, N90 );
nor g018 ( new_n169_, N87, N88 );
nor g019 ( N423, new_n169_, new_n168_ );
nand g020 ( N446, new_n160_, new_n162_ );
nand g021 ( new_n172_, keyIn_0_2, N1, N26, N51 );
not g022 ( new_n173_, keyIn_0_2 );
nand g023 ( new_n174_, N1, N26, N51 );
nand g024 ( new_n175_, new_n174_, new_n173_ );
and g025 ( N447, new_n175_, new_n172_ );
nand g026 ( new_n177_, new_n157_, N13, N55 );
not g027 ( new_n178_, new_n177_ );
and g028 ( N448, new_n178_, N29, N68 );
and g029 ( new_n180_, N59, N68 );
nand g030 ( new_n181_, new_n178_, N74, new_n180_ );
xor g031 ( N449, new_n181_, keyIn_0_12 );
not g032 ( new_n183_, N89 );
nor g033 ( new_n184_, new_n169_, new_n183_ );
xnor g034 ( N450, new_n184_, keyIn_0_9 );
not g035 ( new_n186_, N135 );
nor g036 ( new_n187_, N111, N116 );
xnor g037 ( new_n188_, new_n187_, keyIn_0_6 );
nand g038 ( new_n189_, N111, N116 );
nand g039 ( new_n190_, new_n188_, new_n189_ );
xnor g040 ( new_n191_, N121, N126 );
xnor g041 ( new_n192_, new_n190_, new_n191_ );
nand g042 ( new_n193_, new_n192_, new_n186_ );
or g043 ( new_n194_, new_n193_, keyIn_0_19 );
nand g044 ( new_n195_, new_n193_, keyIn_0_19 );
or g045 ( new_n196_, new_n192_, new_n186_ );
nand g046 ( new_n197_, new_n194_, new_n195_, new_n196_ );
xnor g047 ( new_n198_, N91, N96 );
xnor g048 ( new_n199_, N101, N106 );
xor g049 ( new_n200_, new_n198_, new_n199_ );
xnor g050 ( new_n201_, new_n200_, N130 );
or g051 ( new_n202_, new_n197_, new_n201_ );
nor g052 ( new_n203_, new_n202_, keyIn_0_32 );
and g053 ( new_n204_, new_n202_, keyIn_0_32 );
and g054 ( new_n205_, new_n197_, new_n201_ );
nor g055 ( N767, new_n204_, new_n203_, new_n205_ );
not g056 ( new_n207_, N207 );
xnor g057 ( new_n208_, N183, N189 );
xnor g058 ( new_n209_, N195, N201 );
xnor g059 ( new_n210_, new_n208_, new_n209_ );
nand g060 ( new_n211_, new_n210_, new_n207_ );
xor g061 ( new_n212_, new_n211_, keyIn_0_26 );
or g062 ( new_n213_, new_n210_, new_n207_ );
nand g063 ( new_n214_, new_n212_, new_n213_ );
nor g064 ( new_n215_, N159, N165 );
and g065 ( new_n216_, N159, N165 );
nor g066 ( new_n217_, new_n216_, new_n215_, keyIn_0_13 );
xor g067 ( new_n218_, N171, N177 );
xnor g068 ( new_n219_, new_n217_, new_n218_ );
not g069 ( new_n220_, new_n219_ );
nor g070 ( new_n221_, new_n220_, N130 );
not g071 ( new_n222_, new_n221_ );
or g072 ( new_n223_, new_n222_, keyIn_0_25 );
nand g073 ( new_n224_, new_n222_, keyIn_0_25 );
nand g074 ( new_n225_, new_n220_, N130 );
nand g075 ( new_n226_, new_n223_, keyIn_0_31, new_n224_, new_n225_ );
xor g076 ( N768, new_n226_, new_n214_ );
nand g077 ( new_n228_, N17, N42 );
nand g078 ( new_n229_, N59, N156 );
nor g079 ( new_n230_, N17, N42 );
nor g080 ( new_n231_, new_n230_, new_n229_ );
nand g081 ( new_n232_, new_n231_, new_n175_, new_n172_, new_n228_ );
nand g082 ( new_n233_, N42, N59, N75 );
nand g083 ( new_n234_, new_n157_, new_n233_, N17, N51 );
nand g084 ( new_n235_, new_n232_, new_n234_ );
nand g085 ( new_n236_, new_n235_, N126 );
nand g086 ( new_n237_, new_n236_, keyIn_0_24 );
not g087 ( new_n238_, keyIn_0_24 );
nand g088 ( new_n239_, new_n235_, new_n238_, N126 );
nand g089 ( new_n240_, new_n237_, new_n239_ );
not g090 ( new_n241_, keyIn_0_15 );
and g091 ( new_n242_, N29, N75, N80 );
nand g092 ( new_n243_, new_n175_, N55, new_n172_, new_n242_ );
xnor g093 ( new_n244_, new_n243_, new_n241_ );
xor g094 ( new_n245_, keyIn_0_10, N268 );
nand g095 ( new_n246_, new_n244_, new_n245_ );
nand g096 ( new_n247_, new_n175_, N17, new_n172_, new_n229_ );
nand g097 ( new_n248_, new_n247_, N1 );
nand g098 ( new_n249_, new_n248_, N153 );
nand g099 ( new_n250_, new_n240_, new_n246_, new_n249_ );
nand g100 ( new_n251_, new_n250_, keyIn_0_37, N201 );
not g101 ( new_n252_, keyIn_0_37 );
nand g102 ( new_n253_, new_n250_, N201 );
nand g103 ( new_n254_, new_n253_, new_n252_ );
nand g104 ( new_n255_, new_n254_, new_n251_ );
not g105 ( new_n256_, new_n255_ );
not g106 ( new_n257_, keyIn_0_38 );
not g107 ( new_n258_, N201 );
nand g108 ( new_n259_, new_n240_, new_n258_, new_n246_, new_n249_ );
xnor g109 ( new_n260_, new_n259_, new_n257_ );
nand g110 ( new_n261_, new_n256_, new_n260_ );
xor g111 ( new_n262_, new_n261_, N261 );
or g112 ( new_n263_, new_n262_, keyIn_0_52 );
nand g113 ( new_n264_, new_n262_, keyIn_0_52 );
nand g114 ( new_n265_, new_n263_, N219, new_n264_ );
nand g115 ( new_n266_, N121, N210 );
nand g116 ( new_n267_, new_n265_, new_n266_ );
xnor g117 ( new_n268_, new_n267_, keyIn_0_56 );
nand g118 ( new_n269_, new_n178_, N42, N72, new_n180_ );
not g119 ( new_n270_, new_n269_ );
or g120 ( new_n271_, new_n270_, keyIn_0_8 );
nand g121 ( new_n272_, new_n270_, keyIn_0_8 );
nand g122 ( new_n273_, new_n271_, N73, new_n272_ );
xnor g123 ( new_n274_, new_n273_, keyIn_0_11 );
xor g124 ( new_n275_, new_n274_, keyIn_0_14 );
xnor g125 ( new_n276_, new_n275_, keyIn_0_16 );
not g126 ( new_n277_, new_n276_ );
nand g127 ( new_n278_, new_n277_, N201 );
xnor g128 ( new_n279_, new_n278_, keyIn_0_28 );
nand g129 ( new_n280_, new_n250_, N246 );
nand g130 ( new_n281_, N255, N267 );
nand g131 ( new_n282_, new_n279_, new_n280_, new_n281_ );
nand g132 ( new_n283_, new_n255_, N237 );
and g133 ( new_n284_, new_n283_, keyIn_0_50 );
nor g134 ( new_n285_, new_n283_, keyIn_0_50 );
not g135 ( new_n286_, N228 );
nor g136 ( new_n287_, new_n261_, new_n286_ );
nor g137 ( new_n288_, new_n282_, new_n284_, new_n285_, new_n287_ );
nand g138 ( N850, new_n288_, new_n268_ );
not g139 ( new_n290_, keyIn_0_55 );
not g140 ( new_n291_, N189 );
not g141 ( new_n292_, keyIn_0_23 );
nand g142 ( new_n293_, new_n235_, N116 );
nand g143 ( new_n294_, new_n293_, new_n292_ );
nand g144 ( new_n295_, new_n248_, N146 );
nand g145 ( new_n296_, new_n235_, keyIn_0_23, N116 );
nand g146 ( new_n297_, new_n246_, new_n294_, new_n295_, new_n296_ );
nand g147 ( new_n298_, new_n297_, keyIn_0_30 );
not g148 ( new_n299_, keyIn_0_30 );
and g149 ( new_n300_, new_n296_, new_n295_ );
nand g150 ( new_n301_, new_n300_, new_n299_, new_n246_, new_n294_ );
nand g151 ( new_n302_, new_n298_, new_n301_ );
nand g152 ( new_n303_, new_n302_, new_n291_ );
nand g153 ( new_n304_, new_n248_, N149 );
nand g154 ( new_n305_, new_n235_, N121 );
nand g155 ( new_n306_, new_n246_, new_n304_, new_n305_ );
or g156 ( new_n307_, new_n306_, N195 );
nand g157 ( new_n308_, new_n255_, keyIn_0_51, new_n303_, new_n307_ );
not g158 ( new_n309_, keyIn_0_51 );
nand g159 ( new_n310_, new_n255_, new_n303_, new_n307_ );
nand g160 ( new_n311_, new_n310_, new_n309_ );
nand g161 ( new_n312_, new_n311_, new_n308_ );
nand g162 ( new_n313_, new_n260_, new_n303_, N261, new_n307_ );
or g163 ( new_n314_, new_n313_, keyIn_0_42 );
nand g164 ( new_n315_, new_n313_, keyIn_0_42 );
and g165 ( new_n316_, new_n306_, N195 );
nand g166 ( new_n317_, new_n303_, new_n316_ );
not g167 ( new_n318_, new_n302_ );
nand g168 ( new_n319_, new_n318_, N189 );
and g169 ( new_n320_, new_n317_, new_n319_ );
nand g170 ( new_n321_, new_n312_, new_n314_, new_n315_, new_n320_ );
nand g171 ( new_n322_, new_n235_, keyIn_0_22, N111 );
not g172 ( new_n323_, keyIn_0_22 );
nand g173 ( new_n324_, new_n235_, N111 );
nand g174 ( new_n325_, new_n324_, new_n323_ );
nand g175 ( new_n326_, new_n325_, new_n322_ );
nand g176 ( new_n327_, new_n248_, N143 );
nand g177 ( new_n328_, new_n326_, keyIn_0_29, new_n246_, new_n327_ );
not g178 ( new_n329_, keyIn_0_29 );
nand g179 ( new_n330_, new_n326_, new_n246_, new_n327_ );
nand g180 ( new_n331_, new_n330_, new_n329_ );
nand g181 ( new_n332_, new_n331_, new_n328_ );
nand g182 ( new_n333_, new_n332_, keyIn_0_36, N183 );
not g183 ( new_n334_, keyIn_0_36 );
nand g184 ( new_n335_, new_n332_, N183 );
nand g185 ( new_n336_, new_n335_, new_n334_ );
nand g186 ( new_n337_, new_n336_, new_n333_ );
or g187 ( new_n338_, new_n332_, N183 );
nand g188 ( new_n339_, new_n337_, new_n338_ );
not g189 ( new_n340_, new_n339_ );
and g190 ( new_n341_, new_n321_, new_n340_ );
or g191 ( new_n342_, new_n341_, keyIn_0_53 );
nand g192 ( new_n343_, new_n341_, keyIn_0_53 );
or g193 ( new_n344_, new_n321_, new_n340_ );
nand g194 ( new_n345_, new_n342_, new_n343_, new_n344_ );
nand g195 ( new_n346_, new_n345_, new_n290_ );
or g196 ( new_n347_, new_n345_, new_n290_ );
nand g197 ( new_n348_, new_n347_, N219, new_n346_ );
nor g198 ( new_n349_, new_n339_, new_n286_ );
nor g199 ( new_n350_, new_n349_, keyIn_0_47 );
nand g200 ( new_n351_, new_n277_, N183 );
xnor g201 ( new_n352_, new_n351_, keyIn_0_27 );
nand g202 ( new_n353_, new_n332_, N246 );
nand g203 ( new_n354_, N106, N210 );
nand g204 ( new_n355_, new_n352_, new_n353_, new_n354_ );
nor g205 ( new_n356_, new_n355_, new_n350_ );
not g206 ( new_n357_, keyIn_0_40 );
nand g207 ( new_n358_, new_n336_, new_n357_, new_n333_ );
nand g208 ( new_n359_, new_n337_, keyIn_0_40 );
and g209 ( new_n360_, new_n359_, new_n358_ );
nand g210 ( new_n361_, new_n360_, N237 );
nand g211 ( new_n362_, new_n349_, keyIn_0_47 );
nand g212 ( N863, new_n348_, new_n356_, new_n361_, new_n362_ );
nand g213 ( new_n364_, new_n260_, N261 );
nand g214 ( new_n365_, new_n364_, new_n256_ );
nand g215 ( new_n366_, new_n365_, new_n307_ );
xor g216 ( new_n367_, new_n316_, keyIn_0_49 );
nand g217 ( new_n368_, new_n366_, new_n367_ );
and g218 ( new_n369_, new_n319_, new_n303_ );
nand g219 ( new_n370_, new_n368_, new_n369_ );
or g220 ( new_n371_, new_n368_, new_n369_ );
nand g221 ( new_n372_, new_n371_, N219, new_n370_ );
nand g222 ( new_n373_, new_n318_, N246 );
nand g223 ( new_n374_, N255, N259 );
and g224 ( new_n375_, new_n373_, new_n374_ );
or g225 ( new_n376_, new_n375_, keyIn_0_41 );
and g226 ( new_n377_, new_n375_, keyIn_0_41 );
not g227 ( new_n378_, N237 );
nor g228 ( new_n379_, new_n319_, new_n378_ );
nor g229 ( new_n380_, new_n276_, new_n291_ );
and g230 ( new_n381_, N111, N210 );
nor g231 ( new_n382_, new_n380_, new_n377_, new_n379_, new_n381_ );
nand g232 ( new_n383_, new_n369_, N228 );
xnor g233 ( new_n384_, new_n383_, keyIn_0_48 );
nand g234 ( N864, new_n382_, new_n372_, new_n376_, new_n384_ );
not g235 ( new_n386_, new_n316_ );
nand g236 ( new_n387_, new_n365_, new_n307_, new_n386_ );
nand g237 ( new_n388_, new_n386_, new_n307_ );
nand g238 ( new_n389_, new_n364_, new_n256_, new_n388_ );
nand g239 ( new_n390_, new_n387_, N219, new_n389_ );
nand g240 ( new_n391_, new_n277_, N195 );
nor g241 ( new_n392_, new_n388_, new_n286_ );
nor g242 ( new_n393_, new_n386_, new_n378_ );
nand g243 ( new_n394_, new_n306_, N246 );
nand g244 ( new_n395_, N255, N260 );
nand g245 ( new_n396_, N116, N210 );
nand g246 ( new_n397_, new_n394_, new_n395_, new_n396_ );
nor g247 ( new_n398_, new_n392_, new_n393_, new_n397_ );
nand g248 ( N865, new_n391_, new_n390_, new_n398_ );
nand g249 ( new_n400_, new_n321_, new_n338_ );
nand g250 ( new_n401_, new_n360_, keyIn_0_46 );
not g251 ( new_n402_, keyIn_0_46 );
nand g252 ( new_n403_, new_n359_, new_n358_ );
nand g253 ( new_n404_, new_n403_, new_n402_ );
nand g254 ( new_n405_, new_n400_, new_n401_, new_n404_ );
nand g255 ( new_n406_, new_n405_, keyIn_0_54 );
not g256 ( new_n407_, keyIn_0_54 );
nand g257 ( new_n408_, new_n400_, new_n401_, new_n407_, new_n404_ );
nand g258 ( new_n409_, new_n406_, new_n408_ );
not g259 ( new_n410_, N268 );
nand g260 ( new_n411_, N447, N17, new_n410_, new_n242_ );
xor g261 ( new_n412_, new_n411_, keyIn_0_18 );
and g262 ( new_n413_, N447, N55, new_n229_ );
nand g263 ( new_n414_, new_n413_, N153 );
nand g264 ( new_n415_, new_n235_, N106 );
nand g265 ( new_n416_, N138, N152 );
nand g266 ( new_n417_, new_n412_, new_n414_, new_n415_, new_n416_ );
or g267 ( new_n418_, new_n417_, N177 );
nand g268 ( new_n419_, new_n409_, new_n418_ );
nand g269 ( new_n420_, new_n417_, N177 );
nand g270 ( new_n421_, new_n419_, new_n420_ );
nand g271 ( new_n422_, new_n413_, N149 );
xor g272 ( new_n423_, new_n422_, keyIn_0_17 );
nand g273 ( new_n424_, new_n235_, N101 );
nand g274 ( new_n425_, N17, N138 );
nand g275 ( new_n426_, new_n423_, new_n411_, new_n424_, new_n425_ );
nor g276 ( new_n427_, new_n426_, N171 );
not g277 ( new_n428_, new_n427_ );
nand g278 ( new_n429_, new_n421_, new_n428_ );
nand g279 ( new_n430_, new_n426_, N171 );
xnor g280 ( new_n431_, new_n430_, keyIn_0_35 );
nand g281 ( new_n432_, new_n429_, new_n431_ );
nand g282 ( new_n433_, new_n413_, N146 );
and g283 ( new_n434_, new_n433_, new_n411_ );
or g284 ( new_n435_, new_n434_, keyIn_0_21 );
nand g285 ( new_n436_, new_n434_, keyIn_0_21 );
nand g286 ( new_n437_, new_n235_, N96 );
nand g287 ( new_n438_, N51, N138 );
nand g288 ( new_n439_, new_n435_, new_n436_, new_n437_, new_n438_ );
or g289 ( new_n440_, new_n439_, N165 );
nand g290 ( new_n441_, new_n432_, new_n440_ );
nand g291 ( new_n442_, new_n439_, N165 );
nand g292 ( new_n443_, new_n441_, new_n442_ );
nand g293 ( new_n444_, new_n413_, N143 );
nand g294 ( new_n445_, new_n444_, new_n411_ );
or g295 ( new_n446_, new_n445_, keyIn_0_20 );
nand g296 ( new_n447_, new_n445_, keyIn_0_20 );
nand g297 ( new_n448_, new_n235_, N91 );
nand g298 ( new_n449_, N8, N138 );
nand g299 ( new_n450_, new_n446_, new_n447_, new_n448_, new_n449_ );
nor g300 ( new_n451_, new_n450_, N159 );
xor g301 ( new_n452_, new_n451_, keyIn_0_33 );
nand g302 ( new_n453_, new_n443_, new_n452_ );
nand g303 ( new_n454_, new_n450_, N159 );
xnor g304 ( new_n455_, new_n454_, keyIn_0_43 );
nand g305 ( new_n456_, new_n453_, new_n455_ );
nand g306 ( new_n457_, new_n456_, keyIn_0_59 );
not g307 ( new_n458_, keyIn_0_59 );
nand g308 ( new_n459_, new_n453_, new_n458_, new_n455_ );
nand g309 ( N866, new_n457_, new_n459_ );
nand g310 ( new_n461_, new_n418_, new_n420_ );
and g311 ( new_n462_, new_n406_, new_n408_, new_n461_ );
or g312 ( new_n463_, new_n462_, keyIn_0_57 );
nand g313 ( new_n464_, new_n462_, keyIn_0_57 );
nand g314 ( new_n465_, new_n409_, new_n418_, new_n420_ );
nand g315 ( new_n466_, new_n463_, new_n465_, N219, new_n464_ );
nand g316 ( new_n467_, new_n277_, N177 );
nor g317 ( new_n468_, new_n461_, new_n286_ );
nand g318 ( new_n469_, new_n417_, N177, N237 );
nand g319 ( new_n470_, new_n417_, N246 );
nand g320 ( new_n471_, N101, N210 );
nand g321 ( new_n472_, new_n469_, new_n470_, new_n471_ );
nor g322 ( new_n473_, new_n468_, new_n472_ );
nand g323 ( new_n474_, new_n466_, new_n467_, new_n473_ );
xor g324 ( N874, new_n474_, keyIn_0_62 );
and g325 ( new_n476_, new_n452_, new_n454_ );
nand g326 ( new_n477_, new_n443_, new_n476_ );
or g327 ( new_n478_, new_n443_, new_n476_ );
nand g328 ( new_n479_, new_n478_, N219, new_n477_ );
nand g329 ( new_n480_, new_n277_, N159 );
nand g330 ( new_n481_, new_n450_, N246 );
xor g331 ( new_n482_, new_n481_, keyIn_0_34 );
nand g332 ( new_n483_, new_n480_, new_n482_ );
xnor g333 ( new_n484_, new_n483_, keyIn_0_39 );
and g334 ( new_n485_, new_n476_, N228 );
nor g335 ( new_n486_, new_n454_, new_n378_ );
not g336 ( new_n487_, N210 );
nor g337 ( new_n488_, new_n245_, new_n487_ );
nor g338 ( new_n489_, new_n484_, new_n485_, new_n486_, new_n488_ );
nand g339 ( N878, new_n479_, new_n489_ );
nand g340 ( new_n491_, new_n409_, new_n418_, new_n428_ );
not g341 ( new_n492_, new_n431_ );
nor g342 ( new_n493_, new_n492_, keyIn_0_44 );
and g343 ( new_n494_, new_n492_, keyIn_0_44 );
nor g344 ( new_n495_, new_n427_, new_n420_ );
nor g345 ( new_n496_, new_n494_, new_n493_, new_n495_ );
nand g346 ( new_n497_, new_n440_, new_n442_ );
nand g347 ( new_n498_, new_n491_, new_n496_, new_n497_ );
nand g348 ( new_n499_, new_n498_, keyIn_0_58 );
not g349 ( new_n500_, keyIn_0_58 );
nand g350 ( new_n501_, new_n491_, new_n500_, new_n496_, new_n497_ );
nand g351 ( new_n502_, new_n499_, new_n501_ );
nand g352 ( new_n503_, new_n491_, new_n496_ );
nand g353 ( new_n504_, new_n503_, new_n440_, new_n442_ );
nand g354 ( new_n505_, new_n502_, N219, new_n504_ );
nand g355 ( new_n506_, N91, N210 );
xor g356 ( new_n507_, new_n506_, keyIn_0_7 );
nand g357 ( new_n508_, new_n505_, keyIn_0_60, new_n507_ );
not g358 ( new_n509_, keyIn_0_60 );
nand g359 ( new_n510_, new_n505_, new_n507_ );
nand g360 ( new_n511_, new_n510_, new_n509_ );
nand g361 ( new_n512_, new_n511_, new_n508_ );
nor g362 ( new_n513_, new_n497_, new_n286_ );
and g363 ( new_n514_, new_n277_, N165 );
nor g364 ( new_n515_, new_n442_, new_n378_ );
and g365 ( new_n516_, new_n439_, N246 );
nor g366 ( new_n517_, new_n514_, new_n513_, new_n515_, new_n516_ );
nand g367 ( N879, new_n512_, new_n517_ );
nor g368 ( new_n519_, new_n492_, new_n427_ );
nand g369 ( new_n520_, new_n421_, new_n519_ );
not g370 ( new_n521_, new_n519_ );
nand g371 ( new_n522_, new_n419_, new_n420_, new_n521_ );
nand g372 ( new_n523_, new_n520_, N219, new_n522_ );
nand g373 ( new_n524_, N96, N210 );
nand g374 ( new_n525_, new_n523_, keyIn_0_61, new_n524_ );
not g375 ( new_n526_, keyIn_0_61 );
nand g376 ( new_n527_, new_n523_, new_n524_ );
nand g377 ( new_n528_, new_n527_, new_n526_ );
nand g378 ( new_n529_, new_n528_, new_n525_ );
nand g379 ( new_n530_, new_n492_, N237 );
xnor g380 ( new_n531_, new_n530_, keyIn_0_45 );
nand g381 ( new_n532_, new_n519_, N228 );
nand g382 ( new_n533_, new_n277_, N171 );
nand g383 ( new_n534_, new_n426_, N246 );
and g384 ( new_n535_, new_n531_, new_n533_, new_n532_, new_n534_ );
nand g385 ( new_n536_, new_n529_, new_n535_ );
nand g386 ( new_n537_, new_n536_, keyIn_0_63 );
not g387 ( new_n538_, keyIn_0_63 );
nand g388 ( new_n539_, new_n529_, new_n538_, new_n535_ );
nand g389 ( N880, new_n537_, new_n539_ );
endmodule