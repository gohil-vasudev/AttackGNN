module add_mul_mix_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        c_0_, c_1_, c_2_, c_3_, d_0_, d_1_, d_2_, d_3_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, c_0_, c_1_, c_2_, c_3_,
         d_0_, d_1_, d_2_, d_3_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221;

  INV_X1 U116 ( .A(n109), .ZN(Result_7_) );
  XOR2_X1 U117 ( .A(n110), .B(n111), .Z(Result_6_) );
  OR2_X1 U118 ( .A1(n112), .A2(n113), .ZN(n111) );
  OR2_X1 U119 ( .A1(n114), .A2(n115), .ZN(n110) );
  XNOR2_X1 U120 ( .A(n116), .B(n117), .ZN(Result_5_) );
  XOR2_X1 U121 ( .A(n118), .B(n119), .Z(n117) );
  XOR2_X1 U122 ( .A(n120), .B(n121), .Z(Result_4_) );
  XNOR2_X1 U123 ( .A(n122), .B(n123), .ZN(n121) );
  XOR2_X1 U124 ( .A(n124), .B(n125), .Z(Result_3_) );
  XOR2_X1 U125 ( .A(n126), .B(n127), .Z(Result_2_) );
  OR2_X1 U126 ( .A1(n125), .A2(n124), .ZN(n126) );
  XNOR2_X1 U127 ( .A(n128), .B(n129), .ZN(Result_1_) );
  OR3_X1 U128 ( .A1(n130), .A2(n131), .A3(n132), .ZN(Result_0_) );
  INV_X1 U129 ( .A(n133), .ZN(n132) );
  OR2_X1 U130 ( .A1(n134), .A2(n135), .ZN(n133) );
  AND2_X1 U131 ( .A1(n136), .A2(n129), .ZN(n131) );
  XOR2_X1 U132 ( .A(n137), .B(n138), .Z(n129) );
  INV_X1 U133 ( .A(n128), .ZN(n136) );
  OR3_X1 U134 ( .A1(n125), .A2(n124), .A3(n127), .ZN(n128) );
  XNOR2_X1 U135 ( .A(n139), .B(n140), .ZN(n127) );
  OR2_X1 U136 ( .A1(n141), .A2(n142), .ZN(n124) );
  AND2_X1 U137 ( .A1(n123), .A2(n122), .ZN(n142) );
  AND2_X1 U138 ( .A1(n120), .A2(n143), .ZN(n141) );
  OR2_X1 U139 ( .A1(n122), .A2(n123), .ZN(n143) );
  OR2_X1 U140 ( .A1(n112), .A2(n135), .ZN(n123) );
  OR2_X1 U141 ( .A1(n144), .A2(n145), .ZN(n122) );
  AND2_X1 U142 ( .A1(n116), .A2(n119), .ZN(n145) );
  AND2_X1 U143 ( .A1(n146), .A2(n118), .ZN(n144) );
  OR2_X1 U144 ( .A1(n147), .A2(n148), .ZN(n118) );
  INV_X1 U145 ( .A(n149), .ZN(n148) );
  AND2_X1 U146 ( .A1(n150), .A2(n151), .ZN(n147) );
  OR2_X1 U147 ( .A1(n119), .A2(n116), .ZN(n146) );
  OR2_X1 U148 ( .A1(n151), .A2(n109), .ZN(n116) );
  OR2_X1 U149 ( .A1(n112), .A2(n114), .ZN(n109) );
  OR2_X1 U150 ( .A1(n152), .A2(n112), .ZN(n119) );
  INV_X1 U151 ( .A(n153), .ZN(n112) );
  AND2_X1 U152 ( .A1(n154), .A2(n155), .ZN(n153) );
  OR2_X1 U153 ( .A1(c_3_), .A2(d_3_), .ZN(n154) );
  XNOR2_X1 U154 ( .A(n156), .B(n157), .ZN(n120) );
  XNOR2_X1 U155 ( .A(n158), .B(n149), .ZN(n156) );
  XNOR2_X1 U156 ( .A(n159), .B(n160), .ZN(n125) );
  XNOR2_X1 U157 ( .A(n161), .B(n162), .ZN(n159) );
  AND2_X1 U158 ( .A1(n138), .A2(n137), .ZN(n130) );
  XOR2_X1 U159 ( .A(n163), .B(n134), .Z(n137) );
  OR2_X1 U160 ( .A1(n164), .A2(n165), .ZN(n134) );
  AND2_X1 U161 ( .A1(n166), .A2(n167), .ZN(n165) );
  AND2_X1 U162 ( .A1(n168), .A2(n169), .ZN(n164) );
  OR2_X1 U163 ( .A1(n167), .A2(n166), .ZN(n169) );
  OR2_X1 U164 ( .A1(n170), .A2(n135), .ZN(n163) );
  INV_X1 U165 ( .A(n171), .ZN(n138) );
  OR2_X1 U166 ( .A1(n139), .A2(n140), .ZN(n171) );
  OR2_X1 U167 ( .A1(n172), .A2(n173), .ZN(n140) );
  AND2_X1 U168 ( .A1(n161), .A2(n162), .ZN(n173) );
  AND2_X1 U169 ( .A1(n160), .A2(n174), .ZN(n172) );
  OR2_X1 U170 ( .A1(n162), .A2(n161), .ZN(n174) );
  OR2_X1 U171 ( .A1(n175), .A2(n176), .ZN(n161) );
  AND2_X1 U172 ( .A1(n157), .A2(n149), .ZN(n176) );
  AND2_X1 U173 ( .A1(n177), .A2(n158), .ZN(n175) );
  OR2_X1 U174 ( .A1(n178), .A2(n179), .ZN(n158) );
  AND2_X1 U175 ( .A1(n180), .A2(n181), .ZN(n178) );
  OR2_X1 U176 ( .A1(n149), .A2(n157), .ZN(n177) );
  OR2_X1 U177 ( .A1(n115), .A2(n152), .ZN(n157) );
  OR2_X1 U178 ( .A1(n151), .A2(n150), .ZN(n149) );
  OR2_X1 U179 ( .A1(n182), .A2(n114), .ZN(n150) );
  OR2_X1 U180 ( .A1(n115), .A2(n113), .ZN(n151) );
  OR2_X1 U181 ( .A1(n115), .A2(n135), .ZN(n162) );
  XNOR2_X1 U182 ( .A(n183), .B(n184), .ZN(n115) );
  XNOR2_X1 U183 ( .A(n185), .B(c_2_), .ZN(n184) );
  XNOR2_X1 U184 ( .A(n186), .B(n187), .ZN(n160) );
  OR2_X1 U185 ( .A1(n179), .A2(n188), .ZN(n186) );
  INV_X1 U186 ( .A(n189), .ZN(n179) );
  XOR2_X1 U187 ( .A(n190), .B(n166), .Z(n139) );
  OR2_X1 U188 ( .A1(n152), .A2(n170), .ZN(n166) );
  XOR2_X1 U189 ( .A(n168), .B(n167), .Z(n190) );
  OR2_X1 U190 ( .A1(n182), .A2(n135), .ZN(n167) );
  XNOR2_X1 U191 ( .A(n191), .B(n192), .ZN(n135) );
  XOR2_X1 U192 ( .A(b_0_), .B(a_0_), .Z(n192) );
  OR2_X1 U193 ( .A1(n193), .A2(n194), .ZN(n191) );
  AND2_X1 U194 ( .A1(n195), .A2(a_1_), .ZN(n194) );
  AND2_X1 U195 ( .A1(b_1_), .A2(n196), .ZN(n193) );
  OR2_X1 U196 ( .A1(n195), .A2(a_1_), .ZN(n196) );
  INV_X1 U197 ( .A(n197), .ZN(n195) );
  AND2_X1 U198 ( .A1(n189), .A2(n198), .ZN(n168) );
  OR2_X1 U199 ( .A1(n187), .A2(n188), .ZN(n198) );
  OR2_X1 U200 ( .A1(n113), .A2(n170), .ZN(n188) );
  OR2_X1 U201 ( .A1(n182), .A2(n152), .ZN(n187) );
  XNOR2_X1 U202 ( .A(n199), .B(n197), .ZN(n152) );
  OR2_X1 U203 ( .A1(n200), .A2(n201), .ZN(n197) );
  AND2_X1 U204 ( .A1(n202), .A2(n203), .ZN(n201) );
  AND2_X1 U205 ( .A1(n204), .A2(n205), .ZN(n200) );
  OR2_X1 U206 ( .A1(n203), .A2(n202), .ZN(n204) );
  INV_X1 U207 ( .A(n206), .ZN(n202) );
  INV_X1 U208 ( .A(a_2_), .ZN(n203) );
  XNOR2_X1 U209 ( .A(a_1_), .B(b_1_), .ZN(n199) );
  OR2_X1 U210 ( .A1(n180), .A2(n181), .ZN(n189) );
  OR2_X1 U211 ( .A1(n114), .A2(n170), .ZN(n181) );
  XNOR2_X1 U212 ( .A(n207), .B(n208), .ZN(n170) );
  XOR2_X1 U213 ( .A(d_0_), .B(c_0_), .Z(n208) );
  OR2_X1 U214 ( .A1(n209), .A2(n210), .ZN(n207) );
  AND2_X1 U215 ( .A1(n211), .A2(c_1_), .ZN(n210) );
  AND2_X1 U216 ( .A1(d_1_), .A2(n212), .ZN(n209) );
  OR2_X1 U217 ( .A1(n211), .A2(c_1_), .ZN(n212) );
  INV_X1 U218 ( .A(n213), .ZN(n211) );
  OR2_X1 U219 ( .A1(n214), .A2(n206), .ZN(n114) );
  INV_X1 U220 ( .A(n215), .ZN(n214) );
  OR2_X1 U221 ( .A1(a_3_), .A2(b_3_), .ZN(n215) );
  OR2_X1 U222 ( .A1(n113), .A2(n182), .ZN(n180) );
  XNOR2_X1 U223 ( .A(n216), .B(n213), .ZN(n182) );
  OR2_X1 U224 ( .A1(n217), .A2(n218), .ZN(n213) );
  AND2_X1 U225 ( .A1(n155), .A2(n219), .ZN(n218) );
  AND2_X1 U226 ( .A1(n220), .A2(n185), .ZN(n217) );
  INV_X1 U227 ( .A(d_2_), .ZN(n185) );
  OR2_X1 U228 ( .A1(n219), .A2(n155), .ZN(n220) );
  INV_X1 U229 ( .A(n183), .ZN(n155) );
  AND2_X1 U230 ( .A1(c_3_), .A2(d_3_), .ZN(n183) );
  INV_X1 U231 ( .A(c_2_), .ZN(n219) );
  XNOR2_X1 U232 ( .A(c_1_), .B(d_1_), .ZN(n216) );
  XNOR2_X1 U233 ( .A(n206), .B(n221), .ZN(n113) );
  XNOR2_X1 U234 ( .A(n205), .B(a_2_), .ZN(n221) );
  INV_X1 U235 ( .A(b_2_), .ZN(n205) );
  AND2_X1 U236 ( .A1(a_3_), .A2(b_3_), .ZN(n206) );
endmodule

