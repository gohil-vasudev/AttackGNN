module locked_c1908 (  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_;
  INV_X1 g000 ( .A(KEYINPUT22), .ZN(new_n123_) );
  INV_X1 g001 ( .A(G237), .ZN(new_n124_) );
  INV_X1 g002 ( .A(G902), .ZN(new_n125_) );
  AND2_X1 g003 ( .A1(new_n124_), .A2(new_n125_), .ZN(new_n126_) );
  INV_X1 g004 ( .A(new_n126_), .ZN(new_n127_) );
  AND2_X1 g005 ( .A1(new_n127_), .A2(G214), .ZN(new_n128_) );
  INV_X1 g006 ( .A(new_n128_), .ZN(new_n129_) );
  AND2_X1 g007 ( .A1(new_n127_), .A2(G210), .ZN(new_n130_) );
  INV_X1 g008 ( .A(new_n130_), .ZN(new_n131_) );
  AND2_X1 g009 ( .A1(G902), .A2(KEYINPUT15), .ZN(new_n132_) );
  INV_X1 g010 ( .A(new_n132_), .ZN(new_n133_) );
  OR2_X1 g011 ( .A1(G902), .A2(KEYINPUT15), .ZN(new_n134_) );
  AND2_X1 g012 ( .A1(new_n133_), .A2(new_n134_), .ZN(new_n135_) );
  INV_X1 g013 ( .A(G101), .ZN(new_n136_) );
  INV_X1 g014 ( .A(KEYINPUT4), .ZN(new_n137_) );
  AND2_X1 g015 ( .A1(G128), .A2(G143), .ZN(new_n138_) );
  INV_X1 g016 ( .A(new_n138_), .ZN(new_n139_) );
  OR2_X1 g017 ( .A1(G128), .A2(G143), .ZN(new_n140_) );
  AND2_X1 g018 ( .A1(new_n139_), .A2(new_n140_), .ZN(new_n141_) );
  OR2_X1 g019 ( .A1(new_n141_), .A2(new_n137_), .ZN(new_n142_) );
  INV_X1 g020 ( .A(G128), .ZN(new_n143_) );
  INV_X1 g021 ( .A(G143), .ZN(new_n144_) );
  AND2_X1 g022 ( .A1(new_n143_), .A2(new_n144_), .ZN(new_n145_) );
  OR2_X1 g023 ( .A1(new_n138_), .A2(KEYINPUT4), .ZN(new_n146_) );
  OR2_X1 g024 ( .A1(new_n146_), .A2(new_n145_), .ZN(new_n147_) );
  AND2_X1 g025 ( .A1(new_n142_), .A2(new_n147_), .ZN(new_n148_) );
  OR2_X1 g026 ( .A1(new_n148_), .A2(new_n136_), .ZN(new_n149_) );
  OR2_X1 g027 ( .A1(new_n145_), .A2(new_n138_), .ZN(new_n150_) );
  AND2_X1 g028 ( .A1(new_n150_), .A2(KEYINPUT4), .ZN(new_n151_) );
  INV_X1 g029 ( .A(new_n146_), .ZN(new_n152_) );
  AND2_X1 g030 ( .A1(new_n152_), .A2(new_n140_), .ZN(new_n153_) );
  OR2_X1 g031 ( .A1(new_n151_), .A2(new_n153_), .ZN(new_n154_) );
  OR2_X1 g032 ( .A1(new_n154_), .A2(G101), .ZN(new_n155_) );
  AND2_X1 g033 ( .A1(new_n155_), .A2(new_n149_), .ZN(new_n156_) );
  INV_X1 g034 ( .A(G107), .ZN(new_n157_) );
  AND2_X1 g035 ( .A1(G104), .A2(G110), .ZN(new_n158_) );
  INV_X1 g036 ( .A(G104), .ZN(new_n159_) );
  INV_X1 g037 ( .A(G110), .ZN(new_n160_) );
  AND2_X1 g038 ( .A1(new_n159_), .A2(new_n160_), .ZN(new_n161_) );
  OR2_X1 g039 ( .A1(new_n161_), .A2(new_n158_), .ZN(new_n162_) );
  AND2_X1 g040 ( .A1(new_n162_), .A2(new_n157_), .ZN(new_n163_) );
  INV_X1 g041 ( .A(new_n163_), .ZN(new_n164_) );
  OR2_X1 g042 ( .A1(new_n162_), .A2(new_n157_), .ZN(new_n165_) );
  AND2_X1 g043 ( .A1(new_n164_), .A2(new_n165_), .ZN(new_n166_) );
  INV_X1 g044 ( .A(new_n166_), .ZN(new_n167_) );
  OR2_X1 g045 ( .A1(new_n156_), .A2(new_n167_), .ZN(new_n168_) );
  AND2_X1 g046 ( .A1(new_n154_), .A2(G101), .ZN(new_n169_) );
  AND2_X1 g047 ( .A1(new_n148_), .A2(new_n136_), .ZN(new_n170_) );
  OR2_X1 g048 ( .A1(new_n169_), .A2(new_n170_), .ZN(new_n171_) );
  OR2_X1 g049 ( .A1(new_n171_), .A2(new_n166_), .ZN(new_n172_) );
  AND2_X1 g050 ( .A1(new_n168_), .A2(new_n172_), .ZN(new_n173_) );
  INV_X1 g051 ( .A(G116), .ZN(new_n174_) );
  AND2_X1 g052 ( .A1(new_n174_), .A2(G113), .ZN(new_n175_) );
  INV_X1 g053 ( .A(G113), .ZN(new_n176_) );
  AND2_X1 g054 ( .A1(new_n176_), .A2(G116), .ZN(new_n177_) );
  OR2_X1 g055 ( .A1(new_n175_), .A2(new_n177_), .ZN(new_n178_) );
  AND2_X1 g056 ( .A1(G119), .A2(KEYINPUT3), .ZN(new_n179_) );
  INV_X1 g057 ( .A(G119), .ZN(new_n180_) );
  INV_X1 g058 ( .A(KEYINPUT3), .ZN(new_n181_) );
  AND2_X1 g059 ( .A1(new_n180_), .A2(new_n181_), .ZN(new_n182_) );
  OR2_X1 g060 ( .A1(new_n182_), .A2(new_n179_), .ZN(new_n183_) );
  AND2_X1 g061 ( .A1(new_n178_), .A2(new_n183_), .ZN(new_n184_) );
  OR2_X1 g062 ( .A1(new_n176_), .A2(G116), .ZN(new_n185_) );
  OR2_X1 g063 ( .A1(new_n174_), .A2(G113), .ZN(new_n186_) );
  AND2_X1 g064 ( .A1(new_n185_), .A2(new_n186_), .ZN(new_n187_) );
  INV_X1 g065 ( .A(new_n179_), .ZN(new_n188_) );
  OR2_X1 g066 ( .A1(G119), .A2(KEYINPUT3), .ZN(new_n189_) );
  AND2_X1 g067 ( .A1(new_n188_), .A2(new_n189_), .ZN(new_n190_) );
  AND2_X1 g068 ( .A1(new_n187_), .A2(new_n190_), .ZN(new_n191_) );
  OR2_X1 g069 ( .A1(new_n184_), .A2(new_n191_), .ZN(new_n192_) );
  AND2_X1 g070 ( .A1(G122), .A2(KEYINPUT16), .ZN(new_n193_) );
  INV_X1 g071 ( .A(new_n193_), .ZN(new_n194_) );
  OR2_X1 g072 ( .A1(G122), .A2(KEYINPUT16), .ZN(new_n195_) );
  AND2_X1 g073 ( .A1(new_n194_), .A2(new_n195_), .ZN(new_n196_) );
  INV_X1 g074 ( .A(new_n196_), .ZN(new_n197_) );
  AND2_X1 g075 ( .A1(new_n192_), .A2(new_n197_), .ZN(new_n198_) );
  OR2_X1 g076 ( .A1(new_n187_), .A2(new_n190_), .ZN(new_n199_) );
  OR2_X1 g077 ( .A1(new_n178_), .A2(new_n183_), .ZN(new_n200_) );
  AND2_X1 g078 ( .A1(new_n200_), .A2(new_n199_), .ZN(new_n201_) );
  AND2_X1 g079 ( .A1(new_n201_), .A2(new_n196_), .ZN(new_n202_) );
  OR2_X1 g080 ( .A1(new_n198_), .A2(new_n202_), .ZN(new_n203_) );
  INV_X1 g081 ( .A(KEYINPUT17), .ZN(new_n204_) );
  OR2_X1 g082 ( .A1(new_n204_), .A2(KEYINPUT18), .ZN(new_n205_) );
  INV_X1 g083 ( .A(KEYINPUT18), .ZN(new_n206_) );
  OR2_X1 g084 ( .A1(new_n206_), .A2(KEYINPUT17), .ZN(new_n207_) );
  AND2_X1 g085 ( .A1(new_n205_), .A2(new_n207_), .ZN(new_n208_) );
  INV_X1 g086 ( .A(G953), .ZN(new_n209_) );
  AND2_X1 g087 ( .A1(new_n209_), .A2(G224), .ZN(new_n210_) );
  INV_X1 g088 ( .A(new_n210_), .ZN(new_n211_) );
  OR2_X1 g089 ( .A1(new_n208_), .A2(new_n211_), .ZN(new_n212_) );
  AND2_X1 g090 ( .A1(new_n206_), .A2(KEYINPUT17), .ZN(new_n213_) );
  AND2_X1 g091 ( .A1(new_n204_), .A2(KEYINPUT18), .ZN(new_n214_) );
  OR2_X1 g092 ( .A1(new_n213_), .A2(new_n214_), .ZN(new_n215_) );
  OR2_X1 g093 ( .A1(new_n215_), .A2(new_n210_), .ZN(new_n216_) );
  AND2_X1 g094 ( .A1(new_n216_), .A2(new_n212_), .ZN(new_n217_) );
  AND2_X1 g095 ( .A1(G125), .A2(G146), .ZN(new_n218_) );
  INV_X1 g096 ( .A(G125), .ZN(new_n219_) );
  INV_X1 g097 ( .A(G146), .ZN(new_n220_) );
  AND2_X1 g098 ( .A1(new_n219_), .A2(new_n220_), .ZN(new_n221_) );
  OR2_X1 g099 ( .A1(new_n221_), .A2(new_n218_), .ZN(new_n222_) );
  OR2_X1 g100 ( .A1(new_n217_), .A2(new_n222_), .ZN(new_n223_) );
  AND2_X1 g101 ( .A1(new_n215_), .A2(new_n210_), .ZN(new_n224_) );
  AND2_X1 g102 ( .A1(new_n208_), .A2(new_n211_), .ZN(new_n225_) );
  OR2_X1 g103 ( .A1(new_n224_), .A2(new_n225_), .ZN(new_n226_) );
  INV_X1 g104 ( .A(new_n222_), .ZN(new_n227_) );
  OR2_X1 g105 ( .A1(new_n226_), .A2(new_n227_), .ZN(new_n228_) );
  AND2_X1 g106 ( .A1(new_n228_), .A2(new_n223_), .ZN(new_n229_) );
  OR2_X1 g107 ( .A1(new_n203_), .A2(new_n229_), .ZN(new_n230_) );
  OR2_X1 g108 ( .A1(new_n201_), .A2(new_n196_), .ZN(new_n231_) );
  OR2_X1 g109 ( .A1(new_n192_), .A2(new_n197_), .ZN(new_n232_) );
  AND2_X1 g110 ( .A1(new_n231_), .A2(new_n232_), .ZN(new_n233_) );
  AND2_X1 g111 ( .A1(new_n226_), .A2(new_n227_), .ZN(new_n234_) );
  AND2_X1 g112 ( .A1(new_n217_), .A2(new_n222_), .ZN(new_n235_) );
  OR2_X1 g113 ( .A1(new_n234_), .A2(new_n235_), .ZN(new_n236_) );
  OR2_X1 g114 ( .A1(new_n236_), .A2(new_n233_), .ZN(new_n237_) );
  AND2_X1 g115 ( .A1(new_n237_), .A2(new_n230_), .ZN(new_n238_) );
  OR2_X1 g116 ( .A1(new_n238_), .A2(new_n173_), .ZN(new_n239_) );
  AND2_X1 g117 ( .A1(new_n171_), .A2(new_n166_), .ZN(new_n240_) );
  AND2_X1 g118 ( .A1(new_n156_), .A2(new_n167_), .ZN(new_n241_) );
  OR2_X1 g119 ( .A1(new_n240_), .A2(new_n241_), .ZN(new_n242_) );
  AND2_X1 g120 ( .A1(new_n236_), .A2(new_n233_), .ZN(new_n243_) );
  AND2_X1 g121 ( .A1(new_n203_), .A2(new_n229_), .ZN(new_n244_) );
  OR2_X1 g122 ( .A1(new_n244_), .A2(new_n243_), .ZN(new_n245_) );
  OR2_X1 g123 ( .A1(new_n245_), .A2(new_n242_), .ZN(new_n246_) );
  AND2_X1 g124 ( .A1(new_n246_), .A2(new_n239_), .ZN(new_n247_) );
  OR2_X1 g125 ( .A1(new_n247_), .A2(new_n135_), .ZN(new_n248_) );
  OR2_X1 g126 ( .A1(new_n248_), .A2(new_n131_), .ZN(new_n249_) );
  INV_X1 g127 ( .A(new_n135_), .ZN(new_n250_) );
  AND2_X1 g128 ( .A1(new_n245_), .A2(new_n242_), .ZN(new_n251_) );
  AND2_X1 g129 ( .A1(new_n238_), .A2(new_n173_), .ZN(new_n252_) );
  OR2_X1 g130 ( .A1(new_n251_), .A2(new_n252_), .ZN(new_n253_) );
  AND2_X1 g131 ( .A1(new_n253_), .A2(new_n250_), .ZN(new_n254_) );
  OR2_X1 g132 ( .A1(new_n254_), .A2(new_n130_), .ZN(new_n255_) );
  AND2_X1 g133 ( .A1(new_n249_), .A2(new_n255_), .ZN(new_n256_) );
  AND2_X1 g134 ( .A1(new_n256_), .A2(new_n129_), .ZN(new_n257_) );
  AND2_X1 g135 ( .A1(new_n257_), .A2(KEYINPUT19), .ZN(new_n258_) );
  INV_X1 g136 ( .A(KEYINPUT14), .ZN(new_n259_) );
  AND2_X1 g137 ( .A1(G234), .A2(G237), .ZN(new_n260_) );
  OR2_X1 g138 ( .A1(new_n260_), .A2(new_n259_), .ZN(new_n261_) );
  AND2_X1 g139 ( .A1(new_n260_), .A2(new_n259_), .ZN(new_n262_) );
  INV_X1 g140 ( .A(new_n262_), .ZN(new_n263_) );
  AND2_X1 g141 ( .A1(new_n263_), .A2(new_n261_), .ZN(new_n264_) );
  INV_X1 g142 ( .A(new_n264_), .ZN(new_n265_) );
  AND2_X1 g143 ( .A1(new_n265_), .A2(G952), .ZN(new_n266_) );
  AND2_X1 g144 ( .A1(new_n266_), .A2(new_n209_), .ZN(new_n267_) );
  AND2_X1 g145 ( .A1(new_n265_), .A2(G902), .ZN(new_n268_) );
  INV_X1 g146 ( .A(G898), .ZN(new_n269_) );
  AND2_X1 g147 ( .A1(new_n269_), .A2(G953), .ZN(new_n270_) );
  AND2_X1 g148 ( .A1(new_n268_), .A2(new_n270_), .ZN(new_n271_) );
  OR2_X1 g149 ( .A1(new_n267_), .A2(new_n271_), .ZN(new_n272_) );
  INV_X1 g150 ( .A(new_n272_), .ZN(new_n273_) );
  INV_X1 g151 ( .A(KEYINPUT19), .ZN(new_n274_) );
  AND2_X1 g152 ( .A1(new_n254_), .A2(new_n130_), .ZN(new_n275_) );
  AND2_X1 g153 ( .A1(new_n248_), .A2(new_n131_), .ZN(new_n276_) );
  OR2_X1 g154 ( .A1(new_n276_), .A2(new_n275_), .ZN(new_n277_) );
  OR2_X1 g155 ( .A1(new_n277_), .A2(new_n128_), .ZN(new_n278_) );
  AND2_X1 g156 ( .A1(new_n278_), .A2(new_n274_), .ZN(new_n279_) );
  OR2_X1 g157 ( .A1(new_n279_), .A2(new_n273_), .ZN(new_n280_) );
  OR2_X1 g158 ( .A1(new_n280_), .A2(new_n258_), .ZN(new_n281_) );
  AND2_X1 g159 ( .A1(new_n281_), .A2(KEYINPUT0), .ZN(new_n282_) );
  INV_X1 g160 ( .A(KEYINPUT0), .ZN(new_n283_) );
  INV_X1 g161 ( .A(new_n258_), .ZN(new_n284_) );
  OR2_X1 g162 ( .A1(new_n257_), .A2(KEYINPUT19), .ZN(new_n285_) );
  AND2_X1 g163 ( .A1(new_n285_), .A2(new_n272_), .ZN(new_n286_) );
  AND2_X1 g164 ( .A1(new_n286_), .A2(new_n284_), .ZN(new_n287_) );
  AND2_X1 g165 ( .A1(new_n287_), .A2(new_n283_), .ZN(new_n288_) );
  OR2_X1 g166 ( .A1(new_n282_), .A2(new_n288_), .ZN(new_n289_) );
  AND2_X1 g167 ( .A1(new_n250_), .A2(G234), .ZN(new_n290_) );
  INV_X1 g168 ( .A(new_n290_), .ZN(new_n291_) );
  AND2_X1 g169 ( .A1(new_n291_), .A2(KEYINPUT20), .ZN(new_n292_) );
  INV_X1 g170 ( .A(new_n292_), .ZN(new_n293_) );
  OR2_X1 g171 ( .A1(new_n291_), .A2(KEYINPUT20), .ZN(new_n294_) );
  AND2_X1 g172 ( .A1(new_n293_), .A2(new_n294_), .ZN(new_n295_) );
  INV_X1 g173 ( .A(new_n295_), .ZN(new_n296_) );
  AND2_X1 g174 ( .A1(new_n296_), .A2(G221), .ZN(new_n297_) );
  INV_X1 g175 ( .A(new_n297_), .ZN(new_n298_) );
  AND2_X1 g176 ( .A1(new_n298_), .A2(KEYINPUT21), .ZN(new_n299_) );
  INV_X1 g177 ( .A(new_n299_), .ZN(new_n300_) );
  OR2_X1 g178 ( .A1(new_n298_), .A2(KEYINPUT21), .ZN(new_n301_) );
  AND2_X1 g179 ( .A1(new_n300_), .A2(new_n301_), .ZN(new_n302_) );
  INV_X1 g180 ( .A(KEYINPUT10), .ZN(new_n303_) );
  AND2_X1 g181 ( .A1(new_n303_), .A2(G125), .ZN(new_n304_) );
  AND2_X1 g182 ( .A1(new_n219_), .A2(KEYINPUT10), .ZN(new_n305_) );
  OR2_X1 g183 ( .A1(new_n304_), .A2(new_n305_), .ZN(new_n306_) );
  INV_X1 g184 ( .A(new_n306_), .ZN(new_n307_) );
  AND2_X1 g185 ( .A1(G140), .A2(KEYINPUT11), .ZN(new_n308_) );
  INV_X1 g186 ( .A(new_n308_), .ZN(new_n309_) );
  OR2_X1 g187 ( .A1(G140), .A2(KEYINPUT11), .ZN(new_n310_) );
  AND2_X1 g188 ( .A1(new_n309_), .A2(new_n310_), .ZN(new_n311_) );
  AND2_X1 g189 ( .A1(G113), .A2(G122), .ZN(new_n312_) );
  INV_X1 g190 ( .A(G122), .ZN(new_n313_) );
  AND2_X1 g191 ( .A1(new_n176_), .A2(new_n313_), .ZN(new_n314_) );
  OR2_X1 g192 ( .A1(new_n314_), .A2(new_n312_), .ZN(new_n315_) );
  AND2_X1 g193 ( .A1(new_n315_), .A2(new_n311_), .ZN(new_n316_) );
  INV_X1 g194 ( .A(new_n316_), .ZN(new_n317_) );
  OR2_X1 g195 ( .A1(new_n315_), .A2(new_n311_), .ZN(new_n318_) );
  AND2_X1 g196 ( .A1(new_n317_), .A2(new_n318_), .ZN(new_n319_) );
  INV_X1 g197 ( .A(new_n319_), .ZN(new_n320_) );
  AND2_X1 g198 ( .A1(new_n320_), .A2(new_n307_), .ZN(new_n321_) );
  AND2_X1 g199 ( .A1(new_n319_), .A2(new_n306_), .ZN(new_n322_) );
  OR2_X1 g200 ( .A1(new_n321_), .A2(new_n322_), .ZN(new_n323_) );
  AND2_X1 g201 ( .A1(new_n144_), .A2(G104), .ZN(new_n324_) );
  AND2_X1 g202 ( .A1(new_n159_), .A2(G143), .ZN(new_n325_) );
  OR2_X1 g203 ( .A1(new_n324_), .A2(new_n325_), .ZN(new_n326_) );
  INV_X1 g204 ( .A(new_n326_), .ZN(new_n327_) );
  AND2_X1 g205 ( .A1(new_n323_), .A2(new_n327_), .ZN(new_n328_) );
  INV_X1 g206 ( .A(new_n328_), .ZN(new_n329_) );
  OR2_X1 g207 ( .A1(new_n323_), .A2(new_n327_), .ZN(new_n330_) );
  AND2_X1 g208 ( .A1(new_n329_), .A2(new_n330_), .ZN(new_n331_) );
  INV_X1 g209 ( .A(KEYINPUT12), .ZN(new_n332_) );
  INV_X1 g210 ( .A(G131), .ZN(new_n333_) );
  AND2_X1 g211 ( .A1(new_n333_), .A2(new_n220_), .ZN(new_n334_) );
  INV_X1 g212 ( .A(new_n334_), .ZN(new_n335_) );
  AND2_X1 g213 ( .A1(G131), .A2(G146), .ZN(new_n336_) );
  INV_X1 g214 ( .A(new_n336_), .ZN(new_n337_) );
  AND2_X1 g215 ( .A1(new_n335_), .A2(new_n337_), .ZN(new_n338_) );
  INV_X1 g216 ( .A(new_n338_), .ZN(new_n339_) );
  AND2_X1 g217 ( .A1(new_n339_), .A2(new_n332_), .ZN(new_n340_) );
  AND2_X1 g218 ( .A1(new_n338_), .A2(KEYINPUT12), .ZN(new_n341_) );
  OR2_X1 g219 ( .A1(new_n340_), .A2(new_n341_), .ZN(new_n342_) );
  AND2_X1 g220 ( .A1(new_n124_), .A2(G214), .ZN(new_n343_) );
  AND2_X1 g221 ( .A1(new_n343_), .A2(new_n209_), .ZN(new_n344_) );
  AND2_X1 g222 ( .A1(new_n342_), .A2(new_n344_), .ZN(new_n345_) );
  INV_X1 g223 ( .A(new_n345_), .ZN(new_n346_) );
  OR2_X1 g224 ( .A1(new_n342_), .A2(new_n344_), .ZN(new_n347_) );
  AND2_X1 g225 ( .A1(new_n346_), .A2(new_n347_), .ZN(new_n348_) );
  INV_X1 g226 ( .A(new_n348_), .ZN(new_n349_) );
  OR2_X1 g227 ( .A1(new_n331_), .A2(new_n349_), .ZN(new_n350_) );
  AND2_X1 g228 ( .A1(new_n331_), .A2(new_n349_), .ZN(new_n351_) );
  INV_X1 g229 ( .A(new_n351_), .ZN(new_n352_) );
  AND2_X1 g230 ( .A1(new_n352_), .A2(new_n350_), .ZN(new_n353_) );
  INV_X1 g231 ( .A(new_n353_), .ZN(new_n354_) );
  AND2_X1 g232 ( .A1(new_n354_), .A2(new_n125_), .ZN(new_n355_) );
  INV_X1 g233 ( .A(new_n355_), .ZN(new_n356_) );
  AND2_X1 g234 ( .A1(G475), .A2(KEYINPUT13), .ZN(new_n357_) );
  INV_X1 g235 ( .A(new_n357_), .ZN(new_n358_) );
  OR2_X1 g236 ( .A1(G475), .A2(KEYINPUT13), .ZN(new_n359_) );
  AND2_X1 g237 ( .A1(new_n358_), .A2(new_n359_), .ZN(new_n360_) );
  INV_X1 g238 ( .A(new_n360_), .ZN(new_n361_) );
  AND2_X1 g239 ( .A1(new_n356_), .A2(new_n361_), .ZN(new_n362_) );
  AND2_X1 g240 ( .A1(new_n355_), .A2(new_n360_), .ZN(new_n363_) );
  OR2_X1 g241 ( .A1(new_n362_), .A2(new_n363_), .ZN(new_n364_) );
  INV_X1 g242 ( .A(G478), .ZN(new_n365_) );
  INV_X1 g243 ( .A(KEYINPUT8), .ZN(new_n366_) );
  AND2_X1 g244 ( .A1(new_n209_), .A2(G234), .ZN(new_n367_) );
  INV_X1 g245 ( .A(new_n367_), .ZN(new_n368_) );
  AND2_X1 g246 ( .A1(new_n368_), .A2(new_n366_), .ZN(new_n369_) );
  AND2_X1 g247 ( .A1(new_n367_), .A2(KEYINPUT8), .ZN(new_n370_) );
  OR2_X1 g248 ( .A1(new_n369_), .A2(new_n370_), .ZN(new_n371_) );
  AND2_X1 g249 ( .A1(new_n371_), .A2(G217), .ZN(new_n372_) );
  INV_X1 g250 ( .A(KEYINPUT7), .ZN(new_n373_) );
  AND2_X1 g251 ( .A1(new_n373_), .A2(KEYINPUT9), .ZN(new_n374_) );
  INV_X1 g252 ( .A(new_n374_), .ZN(new_n375_) );
  OR2_X1 g253 ( .A1(new_n373_), .A2(KEYINPUT9), .ZN(new_n376_) );
  AND2_X1 g254 ( .A1(new_n375_), .A2(new_n376_), .ZN(new_n377_) );
  INV_X1 g255 ( .A(new_n377_), .ZN(new_n378_) );
  OR2_X1 g256 ( .A1(new_n372_), .A2(new_n378_), .ZN(new_n379_) );
  INV_X1 g257 ( .A(new_n379_), .ZN(new_n380_) );
  AND2_X1 g258 ( .A1(new_n372_), .A2(new_n378_), .ZN(new_n381_) );
  OR2_X1 g259 ( .A1(new_n380_), .A2(new_n381_), .ZN(new_n382_) );
  AND2_X1 g260 ( .A1(new_n382_), .A2(new_n174_), .ZN(new_n383_) );
  INV_X1 g261 ( .A(new_n381_), .ZN(new_n384_) );
  AND2_X1 g262 ( .A1(new_n384_), .A2(new_n379_), .ZN(new_n385_) );
  AND2_X1 g263 ( .A1(new_n385_), .A2(G116), .ZN(new_n386_) );
  OR2_X1 g264 ( .A1(new_n383_), .A2(new_n386_), .ZN(new_n387_) );
  AND2_X1 g265 ( .A1(new_n150_), .A2(G107), .ZN(new_n388_) );
  AND2_X1 g266 ( .A1(new_n141_), .A2(new_n157_), .ZN(new_n389_) );
  OR2_X1 g267 ( .A1(new_n388_), .A2(new_n389_), .ZN(new_n390_) );
  INV_X1 g268 ( .A(new_n390_), .ZN(new_n391_) );
  AND2_X1 g269 ( .A1(new_n387_), .A2(new_n391_), .ZN(new_n392_) );
  OR2_X1 g270 ( .A1(new_n385_), .A2(G116), .ZN(new_n393_) );
  INV_X1 g271 ( .A(new_n386_), .ZN(new_n394_) );
  AND2_X1 g272 ( .A1(new_n394_), .A2(new_n393_), .ZN(new_n395_) );
  AND2_X1 g273 ( .A1(new_n395_), .A2(new_n390_), .ZN(new_n396_) );
  OR2_X1 g274 ( .A1(new_n396_), .A2(new_n392_), .ZN(new_n397_) );
  AND2_X1 g275 ( .A1(G122), .A2(G134), .ZN(new_n398_) );
  INV_X1 g276 ( .A(G134), .ZN(new_n399_) );
  AND2_X1 g277 ( .A1(new_n313_), .A2(new_n399_), .ZN(new_n400_) );
  OR2_X1 g278 ( .A1(new_n400_), .A2(new_n398_), .ZN(new_n401_) );
  INV_X1 g279 ( .A(new_n401_), .ZN(new_n402_) );
  AND2_X1 g280 ( .A1(new_n397_), .A2(new_n402_), .ZN(new_n403_) );
  OR2_X1 g281 ( .A1(new_n395_), .A2(new_n390_), .ZN(new_n404_) );
  OR2_X1 g282 ( .A1(new_n387_), .A2(new_n391_), .ZN(new_n405_) );
  AND2_X1 g283 ( .A1(new_n404_), .A2(new_n405_), .ZN(new_n406_) );
  AND2_X1 g284 ( .A1(new_n406_), .A2(new_n401_), .ZN(new_n407_) );
  OR2_X1 g285 ( .A1(new_n403_), .A2(new_n407_), .ZN(new_n408_) );
  AND2_X1 g286 ( .A1(new_n408_), .A2(new_n125_), .ZN(new_n409_) );
  OR2_X1 g287 ( .A1(new_n409_), .A2(new_n365_), .ZN(new_n410_) );
  OR2_X1 g288 ( .A1(new_n406_), .A2(new_n401_), .ZN(new_n411_) );
  OR2_X1 g289 ( .A1(new_n397_), .A2(new_n402_), .ZN(new_n412_) );
  AND2_X1 g290 ( .A1(new_n412_), .A2(new_n411_), .ZN(new_n413_) );
  OR2_X1 g291 ( .A1(new_n413_), .A2(G902), .ZN(new_n414_) );
  OR2_X1 g292 ( .A1(new_n414_), .A2(G478), .ZN(new_n415_) );
  AND2_X1 g293 ( .A1(new_n415_), .A2(new_n410_), .ZN(new_n416_) );
  AND2_X1 g294 ( .A1(new_n416_), .A2(new_n364_), .ZN(new_n417_) );
  AND2_X1 g295 ( .A1(new_n417_), .A2(new_n302_), .ZN(new_n418_) );
  INV_X1 g296 ( .A(new_n418_), .ZN(new_n419_) );
  OR2_X1 g297 ( .A1(new_n289_), .A2(new_n419_), .ZN(new_n420_) );
  AND2_X1 g298 ( .A1(new_n420_), .A2(new_n123_), .ZN(new_n421_) );
  OR2_X1 g299 ( .A1(new_n287_), .A2(new_n283_), .ZN(new_n422_) );
  OR2_X1 g300 ( .A1(new_n281_), .A2(KEYINPUT0), .ZN(new_n423_) );
  AND2_X1 g301 ( .A1(new_n423_), .A2(new_n422_), .ZN(new_n424_) );
  AND2_X1 g302 ( .A1(new_n424_), .A2(new_n418_), .ZN(new_n425_) );
  AND2_X1 g303 ( .A1(new_n425_), .A2(KEYINPUT22), .ZN(new_n426_) );
  OR2_X1 g304 ( .A1(new_n421_), .A2(new_n426_), .ZN(new_n427_) );
  INV_X1 g305 ( .A(KEYINPUT1), .ZN(new_n428_) );
  OR2_X1 g306 ( .A1(new_n338_), .A2(new_n399_), .ZN(new_n429_) );
  AND2_X1 g307 ( .A1(new_n335_), .A2(new_n399_), .ZN(new_n430_) );
  AND2_X1 g308 ( .A1(new_n430_), .A2(new_n337_), .ZN(new_n431_) );
  INV_X1 g309 ( .A(new_n431_), .ZN(new_n432_) );
  AND2_X1 g310 ( .A1(new_n432_), .A2(new_n429_), .ZN(new_n433_) );
  AND2_X1 g311 ( .A1(G137), .A2(G140), .ZN(new_n434_) );
  INV_X1 g312 ( .A(G137), .ZN(new_n435_) );
  INV_X1 g313 ( .A(G140), .ZN(new_n436_) );
  AND2_X1 g314 ( .A1(new_n435_), .A2(new_n436_), .ZN(new_n437_) );
  OR2_X1 g315 ( .A1(new_n437_), .A2(new_n434_), .ZN(new_n438_) );
  OR2_X1 g316 ( .A1(new_n433_), .A2(new_n438_), .ZN(new_n439_) );
  INV_X1 g317 ( .A(new_n429_), .ZN(new_n440_) );
  OR2_X1 g318 ( .A1(new_n440_), .A2(new_n431_), .ZN(new_n441_) );
  INV_X1 g319 ( .A(new_n438_), .ZN(new_n442_) );
  OR2_X1 g320 ( .A1(new_n441_), .A2(new_n442_), .ZN(new_n443_) );
  AND2_X1 g321 ( .A1(new_n443_), .A2(new_n439_), .ZN(new_n444_) );
  AND2_X1 g322 ( .A1(new_n209_), .A2(G227), .ZN(new_n445_) );
  INV_X1 g323 ( .A(new_n445_), .ZN(new_n446_) );
  OR2_X1 g324 ( .A1(new_n444_), .A2(new_n446_), .ZN(new_n447_) );
  AND2_X1 g325 ( .A1(new_n441_), .A2(new_n442_), .ZN(new_n448_) );
  AND2_X1 g326 ( .A1(new_n433_), .A2(new_n438_), .ZN(new_n449_) );
  OR2_X1 g327 ( .A1(new_n448_), .A2(new_n449_), .ZN(new_n450_) );
  OR2_X1 g328 ( .A1(new_n450_), .A2(new_n445_), .ZN(new_n451_) );
  AND2_X1 g329 ( .A1(new_n451_), .A2(new_n447_), .ZN(new_n452_) );
  OR2_X1 g330 ( .A1(new_n452_), .A2(new_n173_), .ZN(new_n453_) );
  AND2_X1 g331 ( .A1(new_n450_), .A2(new_n445_), .ZN(new_n454_) );
  AND2_X1 g332 ( .A1(new_n444_), .A2(new_n446_), .ZN(new_n455_) );
  OR2_X1 g333 ( .A1(new_n454_), .A2(new_n455_), .ZN(new_n456_) );
  OR2_X1 g334 ( .A1(new_n456_), .A2(new_n242_), .ZN(new_n457_) );
  AND2_X1 g335 ( .A1(new_n457_), .A2(new_n453_), .ZN(new_n458_) );
  OR2_X1 g336 ( .A1(new_n458_), .A2(G902), .ZN(new_n459_) );
  AND2_X1 g337 ( .A1(new_n459_), .A2(G469), .ZN(new_n460_) );
  INV_X1 g338 ( .A(G469), .ZN(new_n461_) );
  AND2_X1 g339 ( .A1(new_n456_), .A2(new_n242_), .ZN(new_n462_) );
  AND2_X1 g340 ( .A1(new_n452_), .A2(new_n173_), .ZN(new_n463_) );
  OR2_X1 g341 ( .A1(new_n462_), .A2(new_n463_), .ZN(new_n464_) );
  AND2_X1 g342 ( .A1(new_n464_), .A2(new_n125_), .ZN(new_n465_) );
  AND2_X1 g343 ( .A1(new_n465_), .A2(new_n461_), .ZN(new_n466_) );
  OR2_X1 g344 ( .A1(new_n460_), .A2(new_n466_), .ZN(new_n467_) );
  AND2_X1 g345 ( .A1(new_n467_), .A2(new_n428_), .ZN(new_n468_) );
  OR2_X1 g346 ( .A1(new_n465_), .A2(new_n461_), .ZN(new_n469_) );
  OR2_X1 g347 ( .A1(new_n459_), .A2(G469), .ZN(new_n470_) );
  AND2_X1 g348 ( .A1(new_n470_), .A2(new_n469_), .ZN(new_n471_) );
  AND2_X1 g349 ( .A1(new_n471_), .A2(KEYINPUT1), .ZN(new_n472_) );
  OR2_X1 g350 ( .A1(new_n468_), .A2(new_n472_), .ZN(new_n473_) );
  AND2_X1 g351 ( .A1(new_n427_), .A2(new_n473_), .ZN(new_n474_) );
  INV_X1 g352 ( .A(KEYINPUT6), .ZN(new_n475_) );
  AND2_X1 g353 ( .A1(new_n171_), .A2(new_n441_), .ZN(new_n476_) );
  AND2_X1 g354 ( .A1(new_n156_), .A2(new_n433_), .ZN(new_n477_) );
  OR2_X1 g355 ( .A1(new_n476_), .A2(new_n477_), .ZN(new_n478_) );
  AND2_X1 g356 ( .A1(G137), .A2(KEYINPUT5), .ZN(new_n479_) );
  INV_X1 g357 ( .A(new_n479_), .ZN(new_n480_) );
  OR2_X1 g358 ( .A1(G137), .A2(KEYINPUT5), .ZN(new_n481_) );
  AND2_X1 g359 ( .A1(new_n480_), .A2(new_n481_), .ZN(new_n482_) );
  AND2_X1 g360 ( .A1(new_n124_), .A2(G210), .ZN(new_n483_) );
  AND2_X1 g361 ( .A1(new_n483_), .A2(new_n209_), .ZN(new_n484_) );
  OR2_X1 g362 ( .A1(new_n482_), .A2(new_n484_), .ZN(new_n485_) );
  AND2_X1 g363 ( .A1(new_n482_), .A2(new_n484_), .ZN(new_n486_) );
  INV_X1 g364 ( .A(new_n486_), .ZN(new_n487_) );
  AND2_X1 g365 ( .A1(new_n487_), .A2(new_n485_), .ZN(new_n488_) );
  OR2_X1 g366 ( .A1(new_n488_), .A2(new_n201_), .ZN(new_n489_) );
  AND2_X1 g367 ( .A1(new_n488_), .A2(new_n201_), .ZN(new_n490_) );
  INV_X1 g368 ( .A(new_n490_), .ZN(new_n491_) );
  AND2_X1 g369 ( .A1(new_n491_), .A2(new_n489_), .ZN(new_n492_) );
  INV_X1 g370 ( .A(new_n492_), .ZN(new_n493_) );
  AND2_X1 g371 ( .A1(new_n478_), .A2(new_n493_), .ZN(new_n494_) );
  OR2_X1 g372 ( .A1(new_n156_), .A2(new_n433_), .ZN(new_n495_) );
  OR2_X1 g373 ( .A1(new_n171_), .A2(new_n441_), .ZN(new_n496_) );
  AND2_X1 g374 ( .A1(new_n495_), .A2(new_n496_), .ZN(new_n497_) );
  AND2_X1 g375 ( .A1(new_n497_), .A2(new_n492_), .ZN(new_n498_) );
  OR2_X1 g376 ( .A1(new_n494_), .A2(new_n498_), .ZN(new_n499_) );
  AND2_X1 g377 ( .A1(new_n499_), .A2(new_n125_), .ZN(new_n500_) );
  OR2_X1 g378 ( .A1(new_n500_), .A2(G472), .ZN(new_n501_) );
  INV_X1 g379 ( .A(G472), .ZN(new_n502_) );
  OR2_X1 g380 ( .A1(new_n497_), .A2(new_n492_), .ZN(new_n503_) );
  OR2_X1 g381 ( .A1(new_n478_), .A2(new_n493_), .ZN(new_n504_) );
  AND2_X1 g382 ( .A1(new_n504_), .A2(new_n503_), .ZN(new_n505_) );
  OR2_X1 g383 ( .A1(new_n505_), .A2(G902), .ZN(new_n506_) );
  OR2_X1 g384 ( .A1(new_n506_), .A2(new_n502_), .ZN(new_n507_) );
  AND2_X1 g385 ( .A1(new_n507_), .A2(new_n501_), .ZN(new_n508_) );
  OR2_X1 g386 ( .A1(new_n508_), .A2(new_n475_), .ZN(new_n509_) );
  AND2_X1 g387 ( .A1(new_n506_), .A2(new_n502_), .ZN(new_n510_) );
  AND2_X1 g388 ( .A1(new_n500_), .A2(G472), .ZN(new_n511_) );
  OR2_X1 g389 ( .A1(new_n510_), .A2(new_n511_), .ZN(new_n512_) );
  OR2_X1 g390 ( .A1(new_n512_), .A2(KEYINPUT6), .ZN(new_n513_) );
  AND2_X1 g391 ( .A1(new_n513_), .A2(new_n509_), .ZN(new_n514_) );
  AND2_X1 g392 ( .A1(G110), .A2(G128), .ZN(new_n515_) );
  AND2_X1 g393 ( .A1(new_n160_), .A2(new_n143_), .ZN(new_n516_) );
  OR2_X1 g394 ( .A1(new_n516_), .A2(new_n515_), .ZN(new_n517_) );
  AND2_X1 g395 ( .A1(G119), .A2(G146), .ZN(new_n518_) );
  AND2_X1 g396 ( .A1(new_n180_), .A2(new_n220_), .ZN(new_n519_) );
  OR2_X1 g397 ( .A1(new_n519_), .A2(new_n518_), .ZN(new_n520_) );
  AND2_X1 g398 ( .A1(new_n517_), .A2(new_n520_), .ZN(new_n521_) );
  INV_X1 g399 ( .A(new_n521_), .ZN(new_n522_) );
  OR2_X1 g400 ( .A1(new_n517_), .A2(new_n520_), .ZN(new_n523_) );
  AND2_X1 g401 ( .A1(new_n522_), .A2(new_n523_), .ZN(new_n524_) );
  INV_X1 g402 ( .A(new_n524_), .ZN(new_n525_) );
  AND2_X1 g403 ( .A1(new_n307_), .A2(new_n442_), .ZN(new_n526_) );
  AND2_X1 g404 ( .A1(new_n306_), .A2(new_n438_), .ZN(new_n527_) );
  OR2_X1 g405 ( .A1(new_n526_), .A2(new_n527_), .ZN(new_n528_) );
  AND2_X1 g406 ( .A1(new_n525_), .A2(new_n528_), .ZN(new_n529_) );
  INV_X1 g407 ( .A(new_n526_), .ZN(new_n530_) );
  INV_X1 g408 ( .A(new_n527_), .ZN(new_n531_) );
  AND2_X1 g409 ( .A1(new_n530_), .A2(new_n531_), .ZN(new_n532_) );
  AND2_X1 g410 ( .A1(new_n532_), .A2(new_n524_), .ZN(new_n533_) );
  OR2_X1 g411 ( .A1(new_n533_), .A2(new_n529_), .ZN(new_n534_) );
  AND2_X1 g412 ( .A1(new_n371_), .A2(G221), .ZN(new_n535_) );
  INV_X1 g413 ( .A(KEYINPUT23), .ZN(new_n536_) );
  AND2_X1 g414 ( .A1(new_n536_), .A2(KEYINPUT24), .ZN(new_n537_) );
  INV_X1 g415 ( .A(new_n537_), .ZN(new_n538_) );
  OR2_X1 g416 ( .A1(new_n536_), .A2(KEYINPUT24), .ZN(new_n539_) );
  AND2_X1 g417 ( .A1(new_n538_), .A2(new_n539_), .ZN(new_n540_) );
  INV_X1 g418 ( .A(new_n540_), .ZN(new_n541_) );
  OR2_X1 g419 ( .A1(new_n535_), .A2(new_n541_), .ZN(new_n542_) );
  INV_X1 g420 ( .A(new_n542_), .ZN(new_n543_) );
  AND2_X1 g421 ( .A1(new_n535_), .A2(new_n541_), .ZN(new_n544_) );
  OR2_X1 g422 ( .A1(new_n543_), .A2(new_n544_), .ZN(new_n545_) );
  AND2_X1 g423 ( .A1(new_n534_), .A2(new_n545_), .ZN(new_n546_) );
  OR2_X1 g424 ( .A1(new_n532_), .A2(new_n524_), .ZN(new_n547_) );
  OR2_X1 g425 ( .A1(new_n525_), .A2(new_n528_), .ZN(new_n548_) );
  AND2_X1 g426 ( .A1(new_n547_), .A2(new_n548_), .ZN(new_n549_) );
  INV_X1 g427 ( .A(new_n544_), .ZN(new_n550_) );
  AND2_X1 g428 ( .A1(new_n550_), .A2(new_n542_), .ZN(new_n551_) );
  AND2_X1 g429 ( .A1(new_n549_), .A2(new_n551_), .ZN(new_n552_) );
  OR2_X1 g430 ( .A1(new_n546_), .A2(new_n552_), .ZN(new_n553_) );
  AND2_X1 g431 ( .A1(new_n553_), .A2(new_n125_), .ZN(new_n554_) );
  AND2_X1 g432 ( .A1(new_n296_), .A2(G217), .ZN(new_n555_) );
  INV_X1 g433 ( .A(new_n555_), .ZN(new_n556_) );
  OR2_X1 g434 ( .A1(new_n554_), .A2(new_n556_), .ZN(new_n557_) );
  OR2_X1 g435 ( .A1(new_n549_), .A2(new_n551_), .ZN(new_n558_) );
  OR2_X1 g436 ( .A1(new_n534_), .A2(new_n545_), .ZN(new_n559_) );
  AND2_X1 g437 ( .A1(new_n559_), .A2(new_n558_), .ZN(new_n560_) );
  OR2_X1 g438 ( .A1(new_n560_), .A2(G902), .ZN(new_n561_) );
  OR2_X1 g439 ( .A1(new_n561_), .A2(new_n555_), .ZN(new_n562_) );
  AND2_X1 g440 ( .A1(new_n562_), .A2(new_n557_), .ZN(new_n563_) );
  OR2_X1 g441 ( .A1(new_n563_), .A2(KEYINPUT25), .ZN(new_n564_) );
  AND2_X1 g442 ( .A1(new_n563_), .A2(KEYINPUT25), .ZN(new_n565_) );
  INV_X1 g443 ( .A(new_n565_), .ZN(new_n566_) );
  AND2_X1 g444 ( .A1(new_n566_), .A2(new_n564_), .ZN(new_n567_) );
  AND2_X1 g445 ( .A1(new_n514_), .A2(new_n567_), .ZN(new_n568_) );
  AND2_X1 g446 ( .A1(new_n474_), .A2(new_n568_), .ZN(new_n569_) );
  INV_X1 g447 ( .A(new_n569_), .ZN(new_n570_) );
  AND2_X1 g448 ( .A1(new_n570_), .A2(G101), .ZN(new_n571_) );
  AND2_X1 g449 ( .A1(new_n569_), .A2(new_n136_), .ZN(new_n572_) );
  OR2_X1 g450 ( .A1(new_n571_), .A2(new_n572_), .ZN(G3) );
  INV_X1 g451 ( .A(new_n364_), .ZN(new_n574_) );
  AND2_X1 g452 ( .A1(new_n416_), .A2(new_n574_), .ZN(new_n575_) );
  AND2_X1 g453 ( .A1(new_n567_), .A2(new_n302_), .ZN(new_n576_) );
  AND2_X1 g454 ( .A1(new_n576_), .A2(new_n467_), .ZN(new_n577_) );
  AND2_X1 g455 ( .A1(new_n577_), .A2(new_n512_), .ZN(new_n578_) );
  AND2_X1 g456 ( .A1(new_n424_), .A2(new_n578_), .ZN(new_n579_) );
  AND2_X1 g457 ( .A1(new_n579_), .A2(new_n575_), .ZN(new_n580_) );
  INV_X1 g458 ( .A(new_n580_), .ZN(new_n581_) );
  AND2_X1 g459 ( .A1(new_n581_), .A2(G104), .ZN(new_n582_) );
  AND2_X1 g460 ( .A1(new_n580_), .A2(new_n159_), .ZN(new_n583_) );
  OR2_X1 g461 ( .A1(new_n582_), .A2(new_n583_), .ZN(G6) );
  AND2_X1 g462 ( .A1(new_n414_), .A2(G478), .ZN(new_n585_) );
  AND2_X1 g463 ( .A1(new_n409_), .A2(new_n365_), .ZN(new_n586_) );
  OR2_X1 g464 ( .A1(new_n585_), .A2(new_n586_), .ZN(new_n587_) );
  AND2_X1 g465 ( .A1(new_n587_), .A2(new_n364_), .ZN(new_n588_) );
  AND2_X1 g466 ( .A1(new_n579_), .A2(new_n588_), .ZN(new_n589_) );
  INV_X1 g467 ( .A(KEYINPUT26), .ZN(new_n590_) );
  AND2_X1 g468 ( .A1(new_n590_), .A2(KEYINPUT27), .ZN(new_n591_) );
  INV_X1 g469 ( .A(new_n591_), .ZN(new_n592_) );
  OR2_X1 g470 ( .A1(new_n590_), .A2(KEYINPUT27), .ZN(new_n593_) );
  AND2_X1 g471 ( .A1(new_n592_), .A2(new_n593_), .ZN(new_n594_) );
  INV_X1 g472 ( .A(new_n594_), .ZN(new_n595_) );
  AND2_X1 g473 ( .A1(new_n589_), .A2(new_n595_), .ZN(new_n596_) );
  INV_X1 g474 ( .A(new_n596_), .ZN(new_n597_) );
  OR2_X1 g475 ( .A1(new_n589_), .A2(new_n595_), .ZN(new_n598_) );
  AND2_X1 g476 ( .A1(new_n597_), .A2(new_n598_), .ZN(new_n599_) );
  INV_X1 g477 ( .A(new_n599_), .ZN(new_n600_) );
  AND2_X1 g478 ( .A1(new_n600_), .A2(new_n157_), .ZN(new_n601_) );
  AND2_X1 g479 ( .A1(new_n599_), .A2(G107), .ZN(new_n602_) );
  OR2_X1 g480 ( .A1(new_n601_), .A2(new_n602_), .ZN(G9) );
  INV_X1 g481 ( .A(KEYINPUT25), .ZN(new_n604_) );
  AND2_X1 g482 ( .A1(new_n561_), .A2(new_n555_), .ZN(new_n605_) );
  AND2_X1 g483 ( .A1(new_n554_), .A2(new_n556_), .ZN(new_n606_) );
  OR2_X1 g484 ( .A1(new_n605_), .A2(new_n606_), .ZN(new_n607_) );
  AND2_X1 g485 ( .A1(new_n607_), .A2(new_n604_), .ZN(new_n608_) );
  OR2_X1 g486 ( .A1(new_n608_), .A2(new_n565_), .ZN(new_n609_) );
  AND2_X1 g487 ( .A1(new_n609_), .A2(new_n512_), .ZN(new_n610_) );
  AND2_X1 g488 ( .A1(new_n474_), .A2(new_n610_), .ZN(new_n611_) );
  INV_X1 g489 ( .A(new_n611_), .ZN(new_n612_) );
  AND2_X1 g490 ( .A1(new_n612_), .A2(G110), .ZN(new_n613_) );
  AND2_X1 g491 ( .A1(new_n611_), .A2(new_n160_), .ZN(new_n614_) );
  OR2_X1 g492 ( .A1(new_n613_), .A2(new_n614_), .ZN(G12) );
  INV_X1 g493 ( .A(KEYINPUT28), .ZN(new_n616_) );
  INV_X1 g494 ( .A(G900), .ZN(new_n617_) );
  AND2_X1 g495 ( .A1(new_n617_), .A2(G953), .ZN(new_n618_) );
  AND2_X1 g496 ( .A1(new_n268_), .A2(new_n618_), .ZN(new_n619_) );
  OR2_X1 g497 ( .A1(new_n267_), .A2(new_n619_), .ZN(new_n620_) );
  AND2_X1 g498 ( .A1(new_n302_), .A2(new_n620_), .ZN(new_n621_) );
  AND2_X1 g499 ( .A1(new_n508_), .A2(new_n621_), .ZN(new_n622_) );
  AND2_X1 g500 ( .A1(new_n622_), .A2(new_n609_), .ZN(new_n623_) );
  AND2_X1 g501 ( .A1(new_n623_), .A2(new_n616_), .ZN(new_n624_) );
  INV_X1 g502 ( .A(new_n624_), .ZN(new_n625_) );
  OR2_X1 g503 ( .A1(new_n623_), .A2(new_n616_), .ZN(new_n626_) );
  AND2_X1 g504 ( .A1(new_n626_), .A2(new_n467_), .ZN(new_n627_) );
  AND2_X1 g505 ( .A1(new_n627_), .A2(new_n625_), .ZN(new_n628_) );
  AND2_X1 g506 ( .A1(new_n284_), .A2(new_n285_), .ZN(new_n629_) );
  AND2_X1 g507 ( .A1(new_n628_), .A2(new_n629_), .ZN(new_n630_) );
  AND2_X1 g508 ( .A1(new_n630_), .A2(new_n588_), .ZN(new_n631_) );
  INV_X1 g509 ( .A(new_n631_), .ZN(new_n632_) );
  INV_X1 g510 ( .A(KEYINPUT29), .ZN(new_n633_) );
  AND2_X1 g511 ( .A1(new_n633_), .A2(G128), .ZN(new_n634_) );
  AND2_X1 g512 ( .A1(new_n143_), .A2(KEYINPUT29), .ZN(new_n635_) );
  OR2_X1 g513 ( .A1(new_n634_), .A2(new_n635_), .ZN(new_n636_) );
  AND2_X1 g514 ( .A1(new_n632_), .A2(new_n636_), .ZN(new_n637_) );
  INV_X1 g515 ( .A(new_n636_), .ZN(new_n638_) );
  AND2_X1 g516 ( .A1(new_n631_), .A2(new_n638_), .ZN(new_n639_) );
  OR2_X1 g517 ( .A1(new_n637_), .A2(new_n639_), .ZN(G30) );
  AND2_X1 g518 ( .A1(new_n577_), .A2(new_n620_), .ZN(new_n641_) );
  AND2_X1 g519 ( .A1(new_n641_), .A2(new_n256_), .ZN(new_n642_) );
  INV_X1 g520 ( .A(KEYINPUT30), .ZN(new_n643_) );
  AND2_X1 g521 ( .A1(new_n508_), .A2(new_n129_), .ZN(new_n644_) );
  INV_X1 g522 ( .A(new_n644_), .ZN(new_n645_) );
  AND2_X1 g523 ( .A1(new_n645_), .A2(new_n643_), .ZN(new_n646_) );
  AND2_X1 g524 ( .A1(new_n644_), .A2(KEYINPUT30), .ZN(new_n647_) );
  OR2_X1 g525 ( .A1(new_n646_), .A2(new_n647_), .ZN(new_n648_) );
  AND2_X1 g526 ( .A1(new_n587_), .A2(new_n574_), .ZN(new_n649_) );
  AND2_X1 g527 ( .A1(new_n649_), .A2(new_n648_), .ZN(new_n650_) );
  AND2_X1 g528 ( .A1(new_n642_), .A2(new_n650_), .ZN(new_n651_) );
  INV_X1 g529 ( .A(new_n651_), .ZN(new_n652_) );
  AND2_X1 g530 ( .A1(new_n652_), .A2(G143), .ZN(new_n653_) );
  AND2_X1 g531 ( .A1(new_n651_), .A2(new_n144_), .ZN(new_n654_) );
  OR2_X1 g532 ( .A1(new_n653_), .A2(new_n654_), .ZN(G45) );
  AND2_X1 g533 ( .A1(new_n630_), .A2(new_n575_), .ZN(new_n656_) );
  INV_X1 g534 ( .A(new_n656_), .ZN(new_n657_) );
  AND2_X1 g535 ( .A1(new_n657_), .A2(G146), .ZN(new_n658_) );
  AND2_X1 g536 ( .A1(new_n656_), .A2(new_n220_), .ZN(new_n659_) );
  OR2_X1 g537 ( .A1(new_n658_), .A2(new_n659_), .ZN(G48) );
  INV_X1 g538 ( .A(KEYINPUT31), .ZN(new_n661_) );
  INV_X1 g539 ( .A(new_n468_), .ZN(new_n662_) );
  INV_X1 g540 ( .A(new_n472_), .ZN(new_n663_) );
  AND2_X1 g541 ( .A1(new_n662_), .A2(new_n663_), .ZN(new_n664_) );
  AND2_X1 g542 ( .A1(new_n576_), .A2(new_n508_), .ZN(new_n665_) );
  AND2_X1 g543 ( .A1(new_n664_), .A2(new_n665_), .ZN(new_n666_) );
  AND2_X1 g544 ( .A1(new_n424_), .A2(new_n666_), .ZN(new_n667_) );
  AND2_X1 g545 ( .A1(new_n667_), .A2(new_n661_), .ZN(new_n668_) );
  INV_X1 g546 ( .A(new_n668_), .ZN(new_n669_) );
  OR2_X1 g547 ( .A1(new_n667_), .A2(new_n661_), .ZN(new_n670_) );
  AND2_X1 g548 ( .A1(new_n669_), .A2(new_n670_), .ZN(new_n671_) );
  INV_X1 g549 ( .A(new_n671_), .ZN(new_n672_) );
  AND2_X1 g550 ( .A1(new_n672_), .A2(new_n575_), .ZN(new_n673_) );
  INV_X1 g551 ( .A(new_n673_), .ZN(new_n674_) );
  AND2_X1 g552 ( .A1(new_n674_), .A2(G113), .ZN(new_n675_) );
  AND2_X1 g553 ( .A1(new_n673_), .A2(new_n176_), .ZN(new_n676_) );
  OR2_X1 g554 ( .A1(new_n675_), .A2(new_n676_), .ZN(G15) );
  AND2_X1 g555 ( .A1(new_n672_), .A2(new_n588_), .ZN(new_n678_) );
  INV_X1 g556 ( .A(new_n678_), .ZN(new_n679_) );
  AND2_X1 g557 ( .A1(new_n679_), .A2(G116), .ZN(new_n680_) );
  AND2_X1 g558 ( .A1(new_n678_), .A2(new_n174_), .ZN(new_n681_) );
  OR2_X1 g559 ( .A1(new_n680_), .A2(new_n681_), .ZN(G18) );
  OR2_X1 g560 ( .A1(new_n425_), .A2(KEYINPUT22), .ZN(new_n683_) );
  OR2_X1 g561 ( .A1(new_n420_), .A2(new_n123_), .ZN(new_n684_) );
  AND2_X1 g562 ( .A1(new_n684_), .A2(new_n683_), .ZN(new_n685_) );
  AND2_X1 g563 ( .A1(new_n514_), .A2(new_n609_), .ZN(new_n686_) );
  AND2_X1 g564 ( .A1(new_n664_), .A2(new_n686_), .ZN(new_n687_) );
  INV_X1 g565 ( .A(new_n687_), .ZN(new_n688_) );
  OR2_X1 g566 ( .A1(new_n685_), .A2(new_n688_), .ZN(new_n689_) );
  AND2_X1 g567 ( .A1(new_n689_), .A2(KEYINPUT32), .ZN(new_n690_) );
  INV_X1 g568 ( .A(KEYINPUT32), .ZN(new_n691_) );
  AND2_X1 g569 ( .A1(new_n427_), .A2(new_n687_), .ZN(new_n692_) );
  AND2_X1 g570 ( .A1(new_n692_), .A2(new_n691_), .ZN(new_n693_) );
  OR2_X1 g571 ( .A1(new_n690_), .A2(new_n693_), .ZN(new_n694_) );
  AND2_X1 g572 ( .A1(new_n694_), .A2(G119), .ZN(new_n695_) );
  OR2_X1 g573 ( .A1(new_n692_), .A2(new_n691_), .ZN(new_n696_) );
  OR2_X1 g574 ( .A1(new_n689_), .A2(KEYINPUT32), .ZN(new_n697_) );
  AND2_X1 g575 ( .A1(new_n697_), .A2(new_n696_), .ZN(new_n698_) );
  AND2_X1 g576 ( .A1(new_n698_), .A2(new_n180_), .ZN(new_n699_) );
  OR2_X1 g577 ( .A1(new_n695_), .A2(new_n699_), .ZN(G21) );
  INV_X1 g578 ( .A(new_n649_), .ZN(new_n701_) );
  INV_X1 g579 ( .A(new_n302_), .ZN(new_n702_) );
  OR2_X1 g580 ( .A1(new_n609_), .A2(new_n702_), .ZN(new_n703_) );
  OR2_X1 g581 ( .A1(new_n514_), .A2(new_n703_), .ZN(new_n704_) );
  OR2_X1 g582 ( .A1(new_n704_), .A2(new_n473_), .ZN(new_n705_) );
  AND2_X1 g583 ( .A1(new_n705_), .A2(KEYINPUT33), .ZN(new_n706_) );
  INV_X1 g584 ( .A(KEYINPUT33), .ZN(new_n707_) );
  AND2_X1 g585 ( .A1(new_n512_), .A2(KEYINPUT6), .ZN(new_n708_) );
  AND2_X1 g586 ( .A1(new_n508_), .A2(new_n475_), .ZN(new_n709_) );
  OR2_X1 g587 ( .A1(new_n708_), .A2(new_n709_), .ZN(new_n710_) );
  AND2_X1 g588 ( .A1(new_n710_), .A2(new_n576_), .ZN(new_n711_) );
  AND2_X1 g589 ( .A1(new_n664_), .A2(new_n711_), .ZN(new_n712_) );
  AND2_X1 g590 ( .A1(new_n712_), .A2(new_n707_), .ZN(new_n713_) );
  OR2_X1 g591 ( .A1(new_n706_), .A2(new_n713_), .ZN(new_n714_) );
  AND2_X1 g592 ( .A1(new_n424_), .A2(new_n714_), .ZN(new_n715_) );
  OR2_X1 g593 ( .A1(new_n715_), .A2(KEYINPUT34), .ZN(new_n716_) );
  INV_X1 g594 ( .A(KEYINPUT34), .ZN(new_n717_) );
  OR2_X1 g595 ( .A1(new_n712_), .A2(new_n707_), .ZN(new_n718_) );
  OR2_X1 g596 ( .A1(new_n705_), .A2(KEYINPUT33), .ZN(new_n719_) );
  AND2_X1 g597 ( .A1(new_n719_), .A2(new_n718_), .ZN(new_n720_) );
  OR2_X1 g598 ( .A1(new_n289_), .A2(new_n720_), .ZN(new_n721_) );
  OR2_X1 g599 ( .A1(new_n721_), .A2(new_n717_), .ZN(new_n722_) );
  AND2_X1 g600 ( .A1(new_n722_), .A2(new_n716_), .ZN(new_n723_) );
  OR2_X1 g601 ( .A1(new_n723_), .A2(new_n701_), .ZN(new_n724_) );
  AND2_X1 g602 ( .A1(new_n724_), .A2(KEYINPUT35), .ZN(new_n725_) );
  INV_X1 g603 ( .A(KEYINPUT35), .ZN(new_n726_) );
  AND2_X1 g604 ( .A1(new_n721_), .A2(new_n717_), .ZN(new_n727_) );
  AND2_X1 g605 ( .A1(new_n715_), .A2(KEYINPUT34), .ZN(new_n728_) );
  OR2_X1 g606 ( .A1(new_n727_), .A2(new_n728_), .ZN(new_n729_) );
  AND2_X1 g607 ( .A1(new_n729_), .A2(new_n649_), .ZN(new_n730_) );
  AND2_X1 g608 ( .A1(new_n730_), .A2(new_n726_), .ZN(new_n731_) );
  OR2_X1 g609 ( .A1(new_n725_), .A2(new_n731_), .ZN(new_n732_) );
  AND2_X1 g610 ( .A1(new_n732_), .A2(new_n313_), .ZN(new_n733_) );
  OR2_X1 g611 ( .A1(new_n730_), .A2(new_n726_), .ZN(new_n734_) );
  OR2_X1 g612 ( .A1(new_n724_), .A2(KEYINPUT35), .ZN(new_n735_) );
  AND2_X1 g613 ( .A1(new_n735_), .A2(new_n734_), .ZN(new_n736_) );
  AND2_X1 g614 ( .A1(new_n736_), .A2(G122), .ZN(new_n737_) );
  OR2_X1 g615 ( .A1(new_n733_), .A2(new_n737_), .ZN(G24) );
  INV_X1 g616 ( .A(KEYINPUT36), .ZN(new_n739_) );
  AND2_X1 g617 ( .A1(new_n621_), .A2(new_n129_), .ZN(new_n740_) );
  AND2_X1 g618 ( .A1(new_n609_), .A2(new_n740_), .ZN(new_n741_) );
  AND2_X1 g619 ( .A1(new_n710_), .A2(new_n741_), .ZN(new_n742_) );
  AND2_X1 g620 ( .A1(new_n575_), .A2(new_n742_), .ZN(new_n743_) );
  AND2_X1 g621 ( .A1(new_n743_), .A2(new_n256_), .ZN(new_n744_) );
  AND2_X1 g622 ( .A1(new_n744_), .A2(new_n739_), .ZN(new_n745_) );
  INV_X1 g623 ( .A(new_n745_), .ZN(new_n746_) );
  OR2_X1 g624 ( .A1(new_n744_), .A2(new_n739_), .ZN(new_n747_) );
  AND2_X1 g625 ( .A1(new_n747_), .A2(new_n664_), .ZN(new_n748_) );
  AND2_X1 g626 ( .A1(new_n748_), .A2(new_n746_), .ZN(new_n749_) );
  INV_X1 g627 ( .A(new_n749_), .ZN(new_n750_) );
  AND2_X1 g628 ( .A1(new_n750_), .A2(new_n219_), .ZN(new_n751_) );
  AND2_X1 g629 ( .A1(new_n749_), .A2(G125), .ZN(new_n752_) );
  OR2_X1 g630 ( .A1(new_n751_), .A2(new_n752_), .ZN(new_n753_) );
  AND2_X1 g631 ( .A1(new_n753_), .A2(KEYINPUT37), .ZN(new_n754_) );
  INV_X1 g632 ( .A(KEYINPUT37), .ZN(new_n755_) );
  INV_X1 g633 ( .A(new_n753_), .ZN(new_n756_) );
  AND2_X1 g634 ( .A1(new_n756_), .A2(new_n755_), .ZN(new_n757_) );
  OR2_X1 g635 ( .A1(new_n757_), .A2(new_n754_), .ZN(G27) );
  INV_X1 g636 ( .A(new_n575_), .ZN(new_n759_) );
  INV_X1 g637 ( .A(KEYINPUT39), .ZN(new_n760_) );
  AND2_X1 g638 ( .A1(new_n277_), .A2(KEYINPUT38), .ZN(new_n761_) );
  INV_X1 g639 ( .A(KEYINPUT38), .ZN(new_n762_) );
  AND2_X1 g640 ( .A1(new_n256_), .A2(new_n762_), .ZN(new_n763_) );
  OR2_X1 g641 ( .A1(new_n761_), .A2(new_n763_), .ZN(new_n764_) );
  AND2_X1 g642 ( .A1(new_n641_), .A2(new_n764_), .ZN(new_n765_) );
  AND2_X1 g643 ( .A1(new_n765_), .A2(new_n648_), .ZN(new_n766_) );
  OR2_X1 g644 ( .A1(new_n766_), .A2(new_n760_), .ZN(new_n767_) );
  AND2_X1 g645 ( .A1(new_n766_), .A2(new_n760_), .ZN(new_n768_) );
  INV_X1 g646 ( .A(new_n768_), .ZN(new_n769_) );
  AND2_X1 g647 ( .A1(new_n769_), .A2(new_n767_), .ZN(new_n770_) );
  OR2_X1 g648 ( .A1(new_n770_), .A2(new_n759_), .ZN(new_n771_) );
  AND2_X1 g649 ( .A1(new_n771_), .A2(KEYINPUT40), .ZN(new_n772_) );
  INV_X1 g650 ( .A(KEYINPUT40), .ZN(new_n773_) );
  INV_X1 g651 ( .A(new_n766_), .ZN(new_n774_) );
  AND2_X1 g652 ( .A1(new_n774_), .A2(KEYINPUT39), .ZN(new_n775_) );
  OR2_X1 g653 ( .A1(new_n775_), .A2(new_n768_), .ZN(new_n776_) );
  AND2_X1 g654 ( .A1(new_n776_), .A2(new_n575_), .ZN(new_n777_) );
  AND2_X1 g655 ( .A1(new_n777_), .A2(new_n773_), .ZN(new_n778_) );
  OR2_X1 g656 ( .A1(new_n772_), .A2(new_n778_), .ZN(new_n779_) );
  AND2_X1 g657 ( .A1(new_n779_), .A2(G131), .ZN(new_n780_) );
  OR2_X1 g658 ( .A1(new_n777_), .A2(new_n773_), .ZN(new_n781_) );
  OR2_X1 g659 ( .A1(new_n771_), .A2(KEYINPUT40), .ZN(new_n782_) );
  AND2_X1 g660 ( .A1(new_n781_), .A2(new_n782_), .ZN(new_n783_) );
  AND2_X1 g661 ( .A1(new_n783_), .A2(new_n333_), .ZN(new_n784_) );
  OR2_X1 g662 ( .A1(new_n780_), .A2(new_n784_), .ZN(G33) );
  AND2_X1 g663 ( .A1(new_n776_), .A2(new_n588_), .ZN(new_n786_) );
  INV_X1 g664 ( .A(new_n786_), .ZN(new_n787_) );
  AND2_X1 g665 ( .A1(new_n787_), .A2(G134), .ZN(new_n788_) );
  AND2_X1 g666 ( .A1(new_n786_), .A2(new_n399_), .ZN(new_n789_) );
  OR2_X1 g667 ( .A1(new_n788_), .A2(new_n789_), .ZN(G36) );
  INV_X1 g668 ( .A(new_n628_), .ZN(new_n791_) );
  INV_X1 g669 ( .A(KEYINPUT41), .ZN(new_n792_) );
  AND2_X1 g670 ( .A1(new_n417_), .A2(new_n764_), .ZN(new_n793_) );
  AND2_X1 g671 ( .A1(new_n793_), .A2(new_n129_), .ZN(new_n794_) );
  OR2_X1 g672 ( .A1(new_n794_), .A2(new_n792_), .ZN(new_n795_) );
  AND2_X1 g673 ( .A1(new_n794_), .A2(new_n792_), .ZN(new_n796_) );
  INV_X1 g674 ( .A(new_n796_), .ZN(new_n797_) );
  AND2_X1 g675 ( .A1(new_n797_), .A2(new_n795_), .ZN(new_n798_) );
  OR2_X1 g676 ( .A1(new_n798_), .A2(new_n791_), .ZN(new_n799_) );
  AND2_X1 g677 ( .A1(new_n799_), .A2(KEYINPUT42), .ZN(new_n800_) );
  INV_X1 g678 ( .A(KEYINPUT42), .ZN(new_n801_) );
  INV_X1 g679 ( .A(new_n794_), .ZN(new_n802_) );
  AND2_X1 g680 ( .A1(new_n802_), .A2(KEYINPUT41), .ZN(new_n803_) );
  OR2_X1 g681 ( .A1(new_n803_), .A2(new_n796_), .ZN(new_n804_) );
  AND2_X1 g682 ( .A1(new_n804_), .A2(new_n628_), .ZN(new_n805_) );
  AND2_X1 g683 ( .A1(new_n805_), .A2(new_n801_), .ZN(new_n806_) );
  OR2_X1 g684 ( .A1(new_n800_), .A2(new_n806_), .ZN(new_n807_) );
  AND2_X1 g685 ( .A1(new_n807_), .A2(G137), .ZN(new_n808_) );
  OR2_X1 g686 ( .A1(new_n805_), .A2(new_n801_), .ZN(new_n809_) );
  OR2_X1 g687 ( .A1(new_n799_), .A2(KEYINPUT42), .ZN(new_n810_) );
  AND2_X1 g688 ( .A1(new_n810_), .A2(new_n809_), .ZN(new_n811_) );
  AND2_X1 g689 ( .A1(new_n811_), .A2(new_n435_), .ZN(new_n812_) );
  OR2_X1 g690 ( .A1(new_n808_), .A2(new_n812_), .ZN(G39) );
  AND2_X1 g691 ( .A1(new_n743_), .A2(new_n473_), .ZN(new_n814_) );
  AND2_X1 g692 ( .A1(new_n814_), .A2(KEYINPUT43), .ZN(new_n815_) );
  INV_X1 g693 ( .A(new_n815_), .ZN(new_n816_) );
  OR2_X1 g694 ( .A1(new_n814_), .A2(KEYINPUT43), .ZN(new_n817_) );
  AND2_X1 g695 ( .A1(new_n817_), .A2(new_n277_), .ZN(new_n818_) );
  AND2_X1 g696 ( .A1(new_n818_), .A2(new_n816_), .ZN(new_n819_) );
  INV_X1 g697 ( .A(new_n819_), .ZN(new_n820_) );
  AND2_X1 g698 ( .A1(new_n820_), .A2(G140), .ZN(new_n821_) );
  AND2_X1 g699 ( .A1(new_n819_), .A2(new_n436_), .ZN(new_n822_) );
  OR2_X1 g700 ( .A1(new_n821_), .A2(new_n822_), .ZN(G42) );
  AND2_X1 g701 ( .A1(new_n694_), .A2(new_n612_), .ZN(new_n824_) );
  INV_X1 g702 ( .A(KEYINPUT44), .ZN(new_n825_) );
  AND2_X1 g703 ( .A1(new_n736_), .A2(new_n825_), .ZN(new_n826_) );
  AND2_X1 g704 ( .A1(new_n826_), .A2(new_n824_), .ZN(new_n827_) );
  OR2_X1 g705 ( .A1(new_n698_), .A2(new_n611_), .ZN(new_n828_) );
  AND2_X1 g706 ( .A1(new_n828_), .A2(KEYINPUT44), .ZN(new_n829_) );
  AND2_X1 g707 ( .A1(new_n732_), .A2(KEYINPUT44), .ZN(new_n830_) );
  OR2_X1 g708 ( .A1(new_n588_), .A2(new_n575_), .ZN(new_n831_) );
  INV_X1 g709 ( .A(new_n579_), .ZN(new_n832_) );
  AND2_X1 g710 ( .A1(new_n671_), .A2(new_n832_), .ZN(new_n833_) );
  INV_X1 g711 ( .A(new_n833_), .ZN(new_n834_) );
  AND2_X1 g712 ( .A1(new_n834_), .A2(new_n831_), .ZN(new_n835_) );
  OR2_X1 g713 ( .A1(new_n835_), .A2(new_n569_), .ZN(new_n836_) );
  OR2_X1 g714 ( .A1(new_n830_), .A2(new_n836_), .ZN(new_n837_) );
  OR2_X1 g715 ( .A1(new_n837_), .A2(new_n829_), .ZN(new_n838_) );
  OR2_X1 g716 ( .A1(new_n838_), .A2(new_n827_), .ZN(new_n839_) );
  AND2_X1 g717 ( .A1(new_n839_), .A2(KEYINPUT45), .ZN(new_n840_) );
  INV_X1 g718 ( .A(KEYINPUT45), .ZN(new_n841_) );
  INV_X1 g719 ( .A(new_n827_), .ZN(new_n842_) );
  OR2_X1 g720 ( .A1(new_n824_), .A2(new_n825_), .ZN(new_n843_) );
  OR2_X1 g721 ( .A1(new_n736_), .A2(new_n825_), .ZN(new_n844_) );
  INV_X1 g722 ( .A(new_n836_), .ZN(new_n845_) );
  AND2_X1 g723 ( .A1(new_n844_), .A2(new_n845_), .ZN(new_n846_) );
  AND2_X1 g724 ( .A1(new_n846_), .A2(new_n843_), .ZN(new_n847_) );
  AND2_X1 g725 ( .A1(new_n847_), .A2(new_n842_), .ZN(new_n848_) );
  AND2_X1 g726 ( .A1(new_n848_), .A2(new_n841_), .ZN(new_n849_) );
  OR2_X1 g727 ( .A1(new_n840_), .A2(new_n849_), .ZN(new_n850_) );
  INV_X1 g728 ( .A(KEYINPUT48), .ZN(new_n851_) );
  INV_X1 g729 ( .A(KEYINPUT46), .ZN(new_n852_) );
  OR2_X1 g730 ( .A1(new_n783_), .A2(new_n811_), .ZN(new_n853_) );
  AND2_X1 g731 ( .A1(new_n853_), .A2(new_n852_), .ZN(new_n854_) );
  AND2_X1 g732 ( .A1(new_n779_), .A2(new_n807_), .ZN(new_n855_) );
  AND2_X1 g733 ( .A1(new_n855_), .A2(KEYINPUT46), .ZN(new_n856_) );
  OR2_X1 g734 ( .A1(new_n854_), .A2(new_n856_), .ZN(new_n857_) );
  AND2_X1 g735 ( .A1(new_n750_), .A2(new_n652_), .ZN(new_n858_) );
  INV_X1 g736 ( .A(KEYINPUT47), .ZN(new_n859_) );
  AND2_X1 g737 ( .A1(new_n630_), .A2(new_n831_), .ZN(new_n860_) );
  OR2_X1 g738 ( .A1(new_n860_), .A2(new_n859_), .ZN(new_n861_) );
  AND2_X1 g739 ( .A1(new_n860_), .A2(new_n859_), .ZN(new_n862_) );
  INV_X1 g740 ( .A(new_n862_), .ZN(new_n863_) );
  AND2_X1 g741 ( .A1(new_n863_), .A2(new_n861_), .ZN(new_n864_) );
  AND2_X1 g742 ( .A1(new_n858_), .A2(new_n864_), .ZN(new_n865_) );
  AND2_X1 g743 ( .A1(new_n857_), .A2(new_n865_), .ZN(new_n866_) );
  AND2_X1 g744 ( .A1(new_n866_), .A2(new_n851_), .ZN(new_n867_) );
  INV_X1 g745 ( .A(new_n867_), .ZN(new_n868_) );
  OR2_X1 g746 ( .A1(new_n866_), .A2(new_n851_), .ZN(new_n869_) );
  AND2_X1 g747 ( .A1(new_n787_), .A2(new_n820_), .ZN(new_n870_) );
  AND2_X1 g748 ( .A1(new_n869_), .A2(new_n870_), .ZN(new_n871_) );
  AND2_X1 g749 ( .A1(new_n871_), .A2(new_n868_), .ZN(new_n872_) );
  AND2_X1 g750 ( .A1(new_n850_), .A2(new_n872_), .ZN(new_n873_) );
  OR2_X1 g751 ( .A1(new_n873_), .A2(KEYINPUT2), .ZN(new_n874_) );
  INV_X1 g752 ( .A(KEYINPUT2), .ZN(new_n875_) );
  OR2_X1 g753 ( .A1(new_n848_), .A2(new_n841_), .ZN(new_n876_) );
  OR2_X1 g754 ( .A1(new_n839_), .A2(KEYINPUT45), .ZN(new_n877_) );
  AND2_X1 g755 ( .A1(new_n877_), .A2(new_n876_), .ZN(new_n878_) );
  OR2_X1 g756 ( .A1(new_n855_), .A2(KEYINPUT46), .ZN(new_n879_) );
  OR2_X1 g757 ( .A1(new_n853_), .A2(new_n852_), .ZN(new_n880_) );
  AND2_X1 g758 ( .A1(new_n880_), .A2(new_n879_), .ZN(new_n881_) );
  INV_X1 g759 ( .A(new_n865_), .ZN(new_n882_) );
  OR2_X1 g760 ( .A1(new_n881_), .A2(new_n882_), .ZN(new_n883_) );
  AND2_X1 g761 ( .A1(new_n883_), .A2(KEYINPUT48), .ZN(new_n884_) );
  INV_X1 g762 ( .A(new_n870_), .ZN(new_n885_) );
  OR2_X1 g763 ( .A1(new_n884_), .A2(new_n885_), .ZN(new_n886_) );
  OR2_X1 g764 ( .A1(new_n886_), .A2(new_n867_), .ZN(new_n887_) );
  OR2_X1 g765 ( .A1(new_n878_), .A2(new_n887_), .ZN(new_n888_) );
  OR2_X1 g766 ( .A1(new_n888_), .A2(new_n875_), .ZN(new_n889_) );
  AND2_X1 g767 ( .A1(new_n889_), .A2(new_n874_), .ZN(new_n890_) );
  INV_X1 g768 ( .A(KEYINPUT52), .ZN(new_n891_) );
  INV_X1 g769 ( .A(KEYINPUT51), .ZN(new_n892_) );
  AND2_X1 g770 ( .A1(new_n473_), .A2(new_n703_), .ZN(new_n893_) );
  AND2_X1 g771 ( .A1(new_n893_), .A2(KEYINPUT50), .ZN(new_n894_) );
  INV_X1 g772 ( .A(new_n894_), .ZN(new_n895_) );
  OR2_X1 g773 ( .A1(new_n893_), .A2(KEYINPUT50), .ZN(new_n896_) );
  INV_X1 g774 ( .A(KEYINPUT49), .ZN(new_n897_) );
  AND2_X1 g775 ( .A1(new_n609_), .A2(new_n702_), .ZN(new_n898_) );
  AND2_X1 g776 ( .A1(new_n898_), .A2(new_n897_), .ZN(new_n899_) );
  INV_X1 g777 ( .A(new_n899_), .ZN(new_n900_) );
  OR2_X1 g778 ( .A1(new_n898_), .A2(new_n897_), .ZN(new_n901_) );
  AND2_X1 g779 ( .A1(new_n901_), .A2(new_n512_), .ZN(new_n902_) );
  AND2_X1 g780 ( .A1(new_n902_), .A2(new_n900_), .ZN(new_n903_) );
  AND2_X1 g781 ( .A1(new_n896_), .A2(new_n903_), .ZN(new_n904_) );
  AND2_X1 g782 ( .A1(new_n904_), .A2(new_n895_), .ZN(new_n905_) );
  OR2_X1 g783 ( .A1(new_n905_), .A2(new_n666_), .ZN(new_n906_) );
  INV_X1 g784 ( .A(new_n906_), .ZN(new_n907_) );
  AND2_X1 g785 ( .A1(new_n907_), .A2(new_n892_), .ZN(new_n908_) );
  AND2_X1 g786 ( .A1(new_n906_), .A2(KEYINPUT51), .ZN(new_n909_) );
  OR2_X1 g787 ( .A1(new_n909_), .A2(new_n798_), .ZN(new_n910_) );
  OR2_X1 g788 ( .A1(new_n910_), .A2(new_n908_), .ZN(new_n911_) );
  AND2_X1 g789 ( .A1(new_n831_), .A2(new_n764_), .ZN(new_n912_) );
  OR2_X1 g790 ( .A1(new_n912_), .A2(new_n417_), .ZN(new_n913_) );
  OR2_X1 g791 ( .A1(new_n587_), .A2(new_n574_), .ZN(new_n914_) );
  INV_X1 g792 ( .A(new_n764_), .ZN(new_n915_) );
  OR2_X1 g793 ( .A1(new_n914_), .A2(new_n915_), .ZN(new_n916_) );
  AND2_X1 g794 ( .A1(new_n916_), .A2(new_n128_), .ZN(new_n917_) );
  OR2_X1 g795 ( .A1(new_n720_), .A2(new_n917_), .ZN(new_n918_) );
  INV_X1 g796 ( .A(new_n918_), .ZN(new_n919_) );
  AND2_X1 g797 ( .A1(new_n919_), .A2(new_n913_), .ZN(new_n920_) );
  INV_X1 g798 ( .A(new_n920_), .ZN(new_n921_) );
  AND2_X1 g799 ( .A1(new_n911_), .A2(new_n921_), .ZN(new_n922_) );
  INV_X1 g800 ( .A(new_n922_), .ZN(new_n923_) );
  AND2_X1 g801 ( .A1(new_n923_), .A2(new_n891_), .ZN(new_n924_) );
  INV_X1 g802 ( .A(new_n924_), .ZN(new_n925_) );
  AND2_X1 g803 ( .A1(new_n922_), .A2(KEYINPUT52), .ZN(new_n926_) );
  INV_X1 g804 ( .A(new_n926_), .ZN(new_n927_) );
  AND2_X1 g805 ( .A1(new_n927_), .A2(new_n266_), .ZN(new_n928_) );
  AND2_X1 g806 ( .A1(new_n928_), .A2(new_n925_), .ZN(new_n929_) );
  AND2_X1 g807 ( .A1(new_n804_), .A2(new_n714_), .ZN(new_n930_) );
  OR2_X1 g808 ( .A1(new_n930_), .A2(G953), .ZN(new_n931_) );
  OR2_X1 g809 ( .A1(new_n929_), .A2(new_n931_), .ZN(new_n932_) );
  OR2_X1 g810 ( .A1(new_n890_), .A2(new_n932_), .ZN(new_n933_) );
  INV_X1 g811 ( .A(new_n933_), .ZN(new_n934_) );
  AND2_X1 g812 ( .A1(new_n934_), .A2(KEYINPUT53), .ZN(new_n935_) );
  INV_X1 g813 ( .A(KEYINPUT53), .ZN(new_n936_) );
  AND2_X1 g814 ( .A1(new_n933_), .A2(new_n936_), .ZN(new_n937_) );
  OR2_X1 g815 ( .A1(new_n935_), .A2(new_n937_), .ZN(G75) );
  INV_X1 g816 ( .A(KEYINPUT56), .ZN(new_n939_) );
  INV_X1 g817 ( .A(KEYINPUT54), .ZN(new_n940_) );
  AND2_X1 g818 ( .A1(new_n940_), .A2(KEYINPUT55), .ZN(new_n941_) );
  INV_X1 g819 ( .A(new_n941_), .ZN(new_n942_) );
  OR2_X1 g820 ( .A1(new_n940_), .A2(KEYINPUT55), .ZN(new_n943_) );
  AND2_X1 g821 ( .A1(new_n942_), .A2(new_n943_), .ZN(new_n944_) );
  INV_X1 g822 ( .A(new_n944_), .ZN(new_n945_) );
  AND2_X1 g823 ( .A1(new_n253_), .A2(new_n945_), .ZN(new_n946_) );
  AND2_X1 g824 ( .A1(new_n247_), .A2(new_n944_), .ZN(new_n947_) );
  OR2_X1 g825 ( .A1(new_n946_), .A2(new_n947_), .ZN(new_n948_) );
  INV_X1 g826 ( .A(new_n948_), .ZN(new_n949_) );
  INV_X1 g827 ( .A(G210), .ZN(new_n950_) );
  AND2_X1 g828 ( .A1(new_n888_), .A2(new_n875_), .ZN(new_n951_) );
  AND2_X1 g829 ( .A1(new_n873_), .A2(KEYINPUT2), .ZN(new_n952_) );
  OR2_X1 g830 ( .A1(new_n951_), .A2(new_n952_), .ZN(new_n953_) );
  OR2_X1 g831 ( .A1(new_n953_), .A2(new_n250_), .ZN(new_n954_) );
  OR2_X1 g832 ( .A1(new_n954_), .A2(new_n950_), .ZN(new_n955_) );
  AND2_X1 g833 ( .A1(new_n955_), .A2(new_n949_), .ZN(new_n956_) );
  OR2_X1 g834 ( .A1(new_n209_), .A2(G952), .ZN(new_n957_) );
  INV_X1 g835 ( .A(new_n957_), .ZN(new_n958_) );
  AND2_X1 g836 ( .A1(new_n890_), .A2(new_n135_), .ZN(new_n959_) );
  AND2_X1 g837 ( .A1(new_n959_), .A2(G210), .ZN(new_n960_) );
  AND2_X1 g838 ( .A1(new_n960_), .A2(new_n948_), .ZN(new_n961_) );
  OR2_X1 g839 ( .A1(new_n961_), .A2(new_n958_), .ZN(new_n962_) );
  OR2_X1 g840 ( .A1(new_n962_), .A2(new_n956_), .ZN(new_n963_) );
  AND2_X1 g841 ( .A1(new_n963_), .A2(new_n939_), .ZN(new_n964_) );
  INV_X1 g842 ( .A(new_n956_), .ZN(new_n965_) );
  OR2_X1 g843 ( .A1(new_n955_), .A2(new_n949_), .ZN(new_n966_) );
  AND2_X1 g844 ( .A1(new_n966_), .A2(new_n957_), .ZN(new_n967_) );
  AND2_X1 g845 ( .A1(new_n967_), .A2(new_n965_), .ZN(new_n968_) );
  AND2_X1 g846 ( .A1(new_n968_), .A2(KEYINPUT56), .ZN(new_n969_) );
  OR2_X1 g847 ( .A1(new_n969_), .A2(new_n964_), .ZN(G51) );
  AND2_X1 g848 ( .A1(KEYINPUT58), .A2(KEYINPUT57), .ZN(new_n971_) );
  INV_X1 g849 ( .A(new_n971_), .ZN(new_n972_) );
  OR2_X1 g850 ( .A1(KEYINPUT58), .A2(KEYINPUT57), .ZN(new_n973_) );
  AND2_X1 g851 ( .A1(new_n972_), .A2(new_n973_), .ZN(new_n974_) );
  INV_X1 g852 ( .A(new_n974_), .ZN(new_n975_) );
  OR2_X1 g853 ( .A1(new_n954_), .A2(new_n461_), .ZN(new_n976_) );
  OR2_X1 g854 ( .A1(new_n976_), .A2(new_n975_), .ZN(new_n977_) );
  AND2_X1 g855 ( .A1(new_n959_), .A2(G469), .ZN(new_n978_) );
  OR2_X1 g856 ( .A1(new_n978_), .A2(new_n974_), .ZN(new_n979_) );
  AND2_X1 g857 ( .A1(new_n977_), .A2(new_n979_), .ZN(new_n980_) );
  INV_X1 g858 ( .A(new_n980_), .ZN(new_n981_) );
  OR2_X1 g859 ( .A1(new_n981_), .A2(new_n464_), .ZN(new_n982_) );
  OR2_X1 g860 ( .A1(new_n980_), .A2(new_n458_), .ZN(new_n983_) );
  AND2_X1 g861 ( .A1(new_n983_), .A2(new_n957_), .ZN(new_n984_) );
  AND2_X1 g862 ( .A1(new_n984_), .A2(new_n982_), .ZN(G54) );
  INV_X1 g863 ( .A(KEYINPUT60), .ZN(new_n986_) );
  INV_X1 g864 ( .A(KEYINPUT59), .ZN(new_n987_) );
  AND2_X1 g865 ( .A1(new_n354_), .A2(new_n987_), .ZN(new_n988_) );
  AND2_X1 g866 ( .A1(new_n353_), .A2(KEYINPUT59), .ZN(new_n989_) );
  OR2_X1 g867 ( .A1(new_n988_), .A2(new_n989_), .ZN(new_n990_) );
  AND2_X1 g868 ( .A1(new_n959_), .A2(G475), .ZN(new_n991_) );
  AND2_X1 g869 ( .A1(new_n991_), .A2(new_n990_), .ZN(new_n992_) );
  INV_X1 g870 ( .A(new_n990_), .ZN(new_n993_) );
  INV_X1 g871 ( .A(G475), .ZN(new_n994_) );
  OR2_X1 g872 ( .A1(new_n954_), .A2(new_n994_), .ZN(new_n995_) );
  AND2_X1 g873 ( .A1(new_n995_), .A2(new_n993_), .ZN(new_n996_) );
  OR2_X1 g874 ( .A1(new_n996_), .A2(new_n958_), .ZN(new_n997_) );
  OR2_X1 g875 ( .A1(new_n997_), .A2(new_n992_), .ZN(new_n998_) );
  AND2_X1 g876 ( .A1(new_n998_), .A2(new_n986_), .ZN(new_n999_) );
  INV_X1 g877 ( .A(new_n992_), .ZN(new_n1000_) );
  OR2_X1 g878 ( .A1(new_n991_), .A2(new_n990_), .ZN(new_n1001_) );
  AND2_X1 g879 ( .A1(new_n1001_), .A2(new_n957_), .ZN(new_n1002_) );
  AND2_X1 g880 ( .A1(new_n1002_), .A2(new_n1000_), .ZN(new_n1003_) );
  AND2_X1 g881 ( .A1(new_n1003_), .A2(KEYINPUT60), .ZN(new_n1004_) );
  OR2_X1 g882 ( .A1(new_n999_), .A2(new_n1004_), .ZN(G60) );
  AND2_X1 g883 ( .A1(new_n959_), .A2(G478), .ZN(new_n1006_) );
  INV_X1 g884 ( .A(new_n1006_), .ZN(new_n1007_) );
  OR2_X1 g885 ( .A1(new_n1007_), .A2(new_n413_), .ZN(new_n1008_) );
  OR2_X1 g886 ( .A1(new_n1006_), .A2(new_n408_), .ZN(new_n1009_) );
  AND2_X1 g887 ( .A1(new_n1009_), .A2(new_n957_), .ZN(new_n1010_) );
  AND2_X1 g888 ( .A1(new_n1010_), .A2(new_n1008_), .ZN(G63) );
  AND2_X1 g889 ( .A1(new_n959_), .A2(G217), .ZN(new_n1012_) );
  INV_X1 g890 ( .A(new_n1012_), .ZN(new_n1013_) );
  OR2_X1 g891 ( .A1(new_n1013_), .A2(new_n560_), .ZN(new_n1014_) );
  OR2_X1 g892 ( .A1(new_n1012_), .A2(new_n553_), .ZN(new_n1015_) );
  AND2_X1 g893 ( .A1(new_n1015_), .A2(new_n957_), .ZN(new_n1016_) );
  AND2_X1 g894 ( .A1(new_n1016_), .A2(new_n1014_), .ZN(G66) );
  AND2_X1 g895 ( .A1(new_n850_), .A2(new_n209_), .ZN(new_n1018_) );
  AND2_X1 g896 ( .A1(G224), .A2(G953), .ZN(new_n1019_) );
  OR2_X1 g897 ( .A1(new_n1019_), .A2(KEYINPUT61), .ZN(new_n1020_) );
  AND2_X1 g898 ( .A1(new_n1019_), .A2(KEYINPUT61), .ZN(new_n1021_) );
  OR2_X1 g899 ( .A1(new_n1021_), .A2(new_n269_), .ZN(new_n1022_) );
  INV_X1 g900 ( .A(new_n1022_), .ZN(new_n1023_) );
  AND2_X1 g901 ( .A1(new_n1023_), .A2(new_n1020_), .ZN(new_n1024_) );
  OR2_X1 g902 ( .A1(new_n1018_), .A2(new_n1024_), .ZN(new_n1025_) );
  AND2_X1 g903 ( .A1(new_n167_), .A2(G101), .ZN(new_n1026_) );
  AND2_X1 g904 ( .A1(new_n166_), .A2(new_n136_), .ZN(new_n1027_) );
  OR2_X1 g905 ( .A1(new_n1026_), .A2(new_n1027_), .ZN(new_n1028_) );
  INV_X1 g906 ( .A(new_n1028_), .ZN(new_n1029_) );
  AND2_X1 g907 ( .A1(new_n1029_), .A2(new_n233_), .ZN(new_n1030_) );
  AND2_X1 g908 ( .A1(new_n1028_), .A2(new_n203_), .ZN(new_n1031_) );
  OR2_X1 g909 ( .A1(new_n1031_), .A2(new_n270_), .ZN(new_n1032_) );
  OR2_X1 g910 ( .A1(new_n1032_), .A2(new_n1030_), .ZN(new_n1033_) );
  INV_X1 g911 ( .A(new_n1033_), .ZN(new_n1034_) );
  AND2_X1 g912 ( .A1(new_n1025_), .A2(new_n1034_), .ZN(new_n1035_) );
  INV_X1 g913 ( .A(new_n1025_), .ZN(new_n1036_) );
  AND2_X1 g914 ( .A1(new_n1036_), .A2(new_n1033_), .ZN(new_n1037_) );
  OR2_X1 g915 ( .A1(new_n1037_), .A2(new_n1035_), .ZN(G69) );
  AND2_X1 g916 ( .A1(new_n154_), .A2(new_n306_), .ZN(new_n1039_) );
  AND2_X1 g917 ( .A1(new_n148_), .A2(new_n307_), .ZN(new_n1040_) );
  OR2_X1 g918 ( .A1(new_n1039_), .A2(new_n1040_), .ZN(new_n1041_) );
  AND2_X1 g919 ( .A1(new_n450_), .A2(new_n1041_), .ZN(new_n1042_) );
  INV_X1 g920 ( .A(new_n1042_), .ZN(new_n1043_) );
  OR2_X1 g921 ( .A1(new_n450_), .A2(new_n1041_), .ZN(new_n1044_) );
  AND2_X1 g922 ( .A1(new_n1043_), .A2(new_n1044_), .ZN(new_n1045_) );
  INV_X1 g923 ( .A(new_n1045_), .ZN(new_n1046_) );
  AND2_X1 g924 ( .A1(new_n872_), .A2(new_n1046_), .ZN(new_n1047_) );
  AND2_X1 g925 ( .A1(new_n887_), .A2(new_n1045_), .ZN(new_n1048_) );
  OR2_X1 g926 ( .A1(new_n1048_), .A2(new_n1047_), .ZN(new_n1049_) );
  AND2_X1 g927 ( .A1(new_n1049_), .A2(new_n209_), .ZN(new_n1050_) );
  OR2_X1 g928 ( .A1(new_n1045_), .A2(G227), .ZN(new_n1051_) );
  INV_X1 g929 ( .A(G227), .ZN(new_n1052_) );
  OR2_X1 g930 ( .A1(new_n1046_), .A2(new_n1052_), .ZN(new_n1053_) );
  AND2_X1 g931 ( .A1(new_n1053_), .A2(new_n1051_), .ZN(new_n1054_) );
  OR2_X1 g932 ( .A1(new_n1054_), .A2(new_n617_), .ZN(new_n1055_) );
  AND2_X1 g933 ( .A1(new_n1055_), .A2(G953), .ZN(new_n1056_) );
  OR2_X1 g934 ( .A1(new_n1050_), .A2(new_n1056_), .ZN(G72) );
  AND2_X1 g935 ( .A1(new_n499_), .A2(KEYINPUT62), .ZN(new_n1058_) );
  INV_X1 g936 ( .A(new_n1058_), .ZN(new_n1059_) );
  OR2_X1 g937 ( .A1(new_n499_), .A2(KEYINPUT62), .ZN(new_n1060_) );
  AND2_X1 g938 ( .A1(new_n1059_), .A2(new_n1060_), .ZN(new_n1061_) );
  INV_X1 g939 ( .A(new_n1061_), .ZN(new_n1062_) );
  AND2_X1 g940 ( .A1(new_n959_), .A2(G472), .ZN(new_n1063_) );
  AND2_X1 g941 ( .A1(new_n1063_), .A2(new_n1062_), .ZN(new_n1064_) );
  OR2_X1 g942 ( .A1(new_n954_), .A2(new_n502_), .ZN(new_n1065_) );
  AND2_X1 g943 ( .A1(new_n1065_), .A2(new_n1061_), .ZN(new_n1066_) );
  OR2_X1 g944 ( .A1(new_n1066_), .A2(new_n958_), .ZN(new_n1067_) );
  OR2_X1 g945 ( .A1(new_n1067_), .A2(new_n1064_), .ZN(new_n1068_) );
  AND2_X1 g946 ( .A1(new_n1068_), .A2(KEYINPUT63), .ZN(new_n1069_) );
  INV_X1 g947 ( .A(KEYINPUT63), .ZN(new_n1070_) );
  INV_X1 g948 ( .A(new_n1064_), .ZN(new_n1071_) );
  OR2_X1 g949 ( .A1(new_n1063_), .A2(new_n1062_), .ZN(new_n1072_) );
  AND2_X1 g950 ( .A1(new_n1072_), .A2(new_n957_), .ZN(new_n1073_) );
  AND2_X1 g951 ( .A1(new_n1073_), .A2(new_n1071_), .ZN(new_n1074_) );
  AND2_X1 g952 ( .A1(new_n1074_), .A2(new_n1070_), .ZN(new_n1075_) );
  OR2_X1 g953 ( .A1(new_n1069_), .A2(new_n1075_), .ZN(G57) );
endmodule


