module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n336_, new_n338_, new_n339_, new_n341_, new_n342_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n361_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n372_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n385_, new_n387_, new_n389_, new_n390_, new_n392_, new_n393_, new_n394_, new_n396_, new_n398_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n434_, new_n435_, new_n437_, new_n438_, new_n440_, new_n441_, new_n443_, new_n444_, new_n445_, new_n447_, new_n448_, new_n449_, new_n451_, new_n453_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n477_, new_n479_, new_n480_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n488_, new_n489_, new_n491_, new_n493_, new_n494_, new_n495_;
  XOR2_X1 g000 ( .A(G155GAT), .B(KEYINPUT3), .Z(new_n138_) );
  XNOR2_X1 g001 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n139_) );
  XNOR2_X1 g002 ( .A(new_n138_), .B(new_n139_), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(G57GAT), .B(KEYINPUT1), .ZN(new_n141_) );
  NAND2_X1 g004 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n142_) );
  XNOR2_X1 g005 ( .A(new_n141_), .B(new_n142_), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(new_n140_), .B(new_n143_), .ZN(new_n144_) );
  XNOR2_X1 g007 ( .A(G120GAT), .B(G127GAT), .ZN(new_n145_) );
  XNOR2_X1 g008 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n146_) );
  XNOR2_X1 g009 ( .A(new_n145_), .B(new_n146_), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n147_), .B(G1GAT), .ZN(new_n148_) );
  XNOR2_X1 g011 ( .A(new_n144_), .B(new_n148_), .ZN(new_n149_) );
  XNOR2_X1 g012 ( .A(G29GAT), .B(G134GAT), .ZN(new_n150_) );
  XNOR2_X1 g013 ( .A(new_n149_), .B(new_n150_), .ZN(new_n151_) );
  XNOR2_X1 g014 ( .A(G85GAT), .B(G162GAT), .ZN(new_n152_) );
  XNOR2_X1 g015 ( .A(new_n151_), .B(new_n152_), .ZN(new_n153_) );
  XOR2_X1 g016 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(new_n154_) );
  XNOR2_X1 g017 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n155_) );
  XNOR2_X1 g018 ( .A(new_n154_), .B(new_n155_), .ZN(new_n156_) );
  XOR2_X1 g019 ( .A(new_n153_), .B(new_n156_), .Z(new_n157_) );
  INV_X1 g020 ( .A(new_n157_), .ZN(new_n158_) );
  XOR2_X1 g021 ( .A(G211GAT), .B(G218GAT), .Z(new_n159_) );
  XNOR2_X1 g022 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n160_) );
  XNOR2_X1 g023 ( .A(new_n159_), .B(new_n160_), .ZN(new_n161_) );
  XNOR2_X1 g024 ( .A(new_n161_), .B(G197GAT), .ZN(new_n162_) );
  XNOR2_X1 g025 ( .A(new_n162_), .B(new_n140_), .ZN(new_n163_) );
  XNOR2_X1 g026 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(new_n164_) );
  XNOR2_X1 g027 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n165_) );
  XNOR2_X1 g028 ( .A(new_n164_), .B(new_n165_), .ZN(new_n166_) );
  INV_X1 g029 ( .A(G148GAT), .ZN(new_n167_) );
  NAND2_X1 g030 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n168_) );
  OR2_X1 g031 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n169_) );
  NAND2_X1 g032 ( .A1(new_n169_), .A2(new_n168_), .ZN(new_n170_) );
  NAND2_X1 g033 ( .A1(new_n170_), .A2(new_n167_), .ZN(new_n171_) );
  NAND3_X1 g034 ( .A1(new_n169_), .A2(G148GAT), .A3(new_n168_), .ZN(new_n172_) );
  NAND2_X1 g035 ( .A1(new_n171_), .A2(new_n172_), .ZN(new_n173_) );
  XNOR2_X1 g036 ( .A(new_n166_), .B(new_n173_), .ZN(new_n174_) );
  NAND2_X1 g037 ( .A1(new_n163_), .A2(new_n174_), .ZN(new_n175_) );
  OR2_X1 g038 ( .A1(new_n163_), .A2(new_n174_), .ZN(new_n176_) );
  NAND2_X1 g039 ( .A1(new_n176_), .A2(new_n175_), .ZN(new_n177_) );
  XNOR2_X1 g040 ( .A(G50GAT), .B(G162GAT), .ZN(new_n178_) );
  NAND2_X1 g041 ( .A1(new_n177_), .A2(new_n178_), .ZN(new_n179_) );
  INV_X1 g042 ( .A(new_n178_), .ZN(new_n180_) );
  NAND3_X1 g043 ( .A1(new_n176_), .A2(new_n175_), .A3(new_n180_), .ZN(new_n181_) );
  NAND2_X1 g044 ( .A1(new_n179_), .A2(new_n181_), .ZN(new_n182_) );
  NAND2_X1 g045 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n183_) );
  NAND2_X1 g046 ( .A1(new_n182_), .A2(new_n183_), .ZN(new_n184_) );
  NAND4_X1 g047 ( .A1(new_n179_), .A2(new_n181_), .A3(G228GAT), .A4(G233GAT), .ZN(new_n185_) );
  XNOR2_X1 g048 ( .A(new_n147_), .B(G15GAT), .ZN(new_n186_) );
  NAND2_X1 g049 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n187_) );
  XNOR2_X1 g050 ( .A(new_n186_), .B(new_n187_), .ZN(new_n188_) );
  XOR2_X1 g051 ( .A(G176GAT), .B(G183GAT), .Z(new_n189_) );
  XNOR2_X1 g052 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n190_) );
  XNOR2_X1 g053 ( .A(new_n189_), .B(new_n190_), .ZN(new_n191_) );
  XNOR2_X1 g054 ( .A(new_n188_), .B(new_n191_), .ZN(new_n192_) );
  XOR2_X1 g055 ( .A(G134GAT), .B(G190GAT), .Z(new_n193_) );
  XNOR2_X1 g056 ( .A(G43GAT), .B(G99GAT), .ZN(new_n194_) );
  XNOR2_X1 g057 ( .A(new_n193_), .B(new_n194_), .ZN(new_n195_) );
  XNOR2_X1 g058 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n196_) );
  XNOR2_X1 g059 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n197_) );
  XNOR2_X1 g060 ( .A(new_n196_), .B(new_n197_), .ZN(new_n198_) );
  XNOR2_X1 g061 ( .A(new_n195_), .B(new_n198_), .ZN(new_n199_) );
  XNOR2_X1 g062 ( .A(new_n192_), .B(new_n199_), .ZN(new_n200_) );
  NAND4_X1 g063 ( .A1(new_n184_), .A2(KEYINPUT26), .A3(new_n185_), .A4(new_n200_), .ZN(new_n201_) );
  INV_X1 g064 ( .A(KEYINPUT26), .ZN(new_n202_) );
  NAND3_X1 g065 ( .A1(new_n184_), .A2(new_n185_), .A3(new_n200_), .ZN(new_n203_) );
  NAND2_X1 g066 ( .A1(new_n203_), .A2(new_n202_), .ZN(new_n204_) );
  NAND2_X1 g067 ( .A1(new_n204_), .A2(new_n201_), .ZN(new_n205_) );
  XOR2_X1 g068 ( .A(G36GAT), .B(G190GAT), .Z(new_n206_) );
  XNOR2_X1 g069 ( .A(new_n162_), .B(new_n206_), .ZN(new_n207_) );
  XNOR2_X1 g070 ( .A(G64GAT), .B(G176GAT), .ZN(new_n208_) );
  XNOR2_X1 g071 ( .A(new_n208_), .B(G92GAT), .ZN(new_n209_) );
  NAND2_X1 g072 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n210_) );
  XNOR2_X1 g073 ( .A(new_n209_), .B(new_n210_), .ZN(new_n211_) );
  XNOR2_X1 g074 ( .A(G8GAT), .B(G183GAT), .ZN(new_n212_) );
  XNOR2_X1 g075 ( .A(new_n211_), .B(new_n212_), .ZN(new_n213_) );
  XNOR2_X1 g076 ( .A(new_n207_), .B(new_n213_), .ZN(new_n214_) );
  XNOR2_X1 g077 ( .A(new_n214_), .B(new_n198_), .ZN(new_n215_) );
  XNOR2_X1 g078 ( .A(new_n215_), .B(KEYINPUT27), .ZN(new_n216_) );
  NAND2_X1 g079 ( .A1(new_n205_), .A2(new_n216_), .ZN(new_n217_) );
  INV_X1 g080 ( .A(KEYINPUT25), .ZN(new_n218_) );
  NAND2_X1 g081 ( .A1(new_n184_), .A2(new_n185_), .ZN(new_n219_) );
  INV_X1 g082 ( .A(new_n200_), .ZN(new_n220_) );
  NAND2_X1 g083 ( .A1(new_n220_), .A2(new_n215_), .ZN(new_n221_) );
  NAND2_X1 g084 ( .A1(new_n219_), .A2(new_n221_), .ZN(new_n222_) );
  NAND2_X1 g085 ( .A1(new_n222_), .A2(new_n218_), .ZN(new_n223_) );
  NAND3_X1 g086 ( .A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT25), .ZN(new_n224_) );
  NAND2_X1 g087 ( .A1(new_n223_), .A2(new_n224_), .ZN(new_n225_) );
  NAND2_X1 g088 ( .A1(new_n217_), .A2(new_n225_), .ZN(new_n226_) );
  NAND2_X1 g089 ( .A1(new_n226_), .A2(new_n157_), .ZN(new_n227_) );
  XNOR2_X1 g090 ( .A(new_n219_), .B(KEYINPUT28), .ZN(new_n228_) );
  AND2_X1 g091 ( .A1(new_n158_), .A2(new_n216_), .ZN(new_n229_) );
  NAND3_X1 g092 ( .A1(new_n229_), .A2(new_n200_), .A3(new_n228_), .ZN(new_n230_) );
  NAND2_X1 g093 ( .A1(new_n227_), .A2(new_n230_), .ZN(new_n231_) );
  XNOR2_X1 g094 ( .A(G106GAT), .B(G218GAT), .ZN(new_n232_) );
  XOR2_X1 g095 ( .A(new_n150_), .B(new_n232_), .Z(new_n233_) );
  INV_X1 g096 ( .A(KEYINPUT7), .ZN(new_n234_) );
  XNOR2_X1 g097 ( .A(G43GAT), .B(KEYINPUT8), .ZN(new_n235_) );
  XNOR2_X1 g098 ( .A(new_n235_), .B(new_n234_), .ZN(new_n236_) );
  XNOR2_X1 g099 ( .A(G85GAT), .B(G99GAT), .ZN(new_n237_) );
  NAND2_X1 g100 ( .A1(new_n237_), .A2(G92GAT), .ZN(new_n238_) );
  INV_X1 g101 ( .A(G92GAT), .ZN(new_n239_) );
  NAND2_X1 g102 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n240_) );
  OR2_X1 g103 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n241_) );
  NAND3_X1 g104 ( .A1(new_n241_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n242_) );
  AND2_X1 g105 ( .A1(new_n238_), .A2(new_n242_), .ZN(new_n243_) );
  NAND2_X1 g106 ( .A1(new_n236_), .A2(new_n243_), .ZN(new_n244_) );
  OR2_X1 g107 ( .A1(new_n236_), .A2(new_n243_), .ZN(new_n245_) );
  NAND2_X1 g108 ( .A1(new_n245_), .A2(new_n244_), .ZN(new_n246_) );
  INV_X1 g109 ( .A(KEYINPUT9), .ZN(new_n247_) );
  XNOR2_X1 g110 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(new_n248_) );
  AND2_X1 g111 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n249_) );
  XNOR2_X1 g112 ( .A(new_n248_), .B(new_n249_), .ZN(new_n250_) );
  XNOR2_X1 g113 ( .A(new_n250_), .B(new_n247_), .ZN(new_n251_) );
  NAND2_X1 g114 ( .A1(new_n246_), .A2(new_n251_), .ZN(new_n252_) );
  XNOR2_X1 g115 ( .A(new_n250_), .B(KEYINPUT9), .ZN(new_n253_) );
  NAND3_X1 g116 ( .A1(new_n253_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n254_) );
  NAND3_X1 g117 ( .A1(new_n252_), .A2(new_n254_), .A3(new_n233_), .ZN(new_n255_) );
  INV_X1 g118 ( .A(new_n233_), .ZN(new_n256_) );
  NAND2_X1 g119 ( .A1(new_n252_), .A2(new_n254_), .ZN(new_n257_) );
  NAND2_X1 g120 ( .A1(new_n257_), .A2(new_n256_), .ZN(new_n258_) );
  NAND3_X1 g121 ( .A1(new_n258_), .A2(new_n180_), .A3(new_n255_), .ZN(new_n259_) );
  NAND2_X1 g122 ( .A1(new_n258_), .A2(new_n255_), .ZN(new_n260_) );
  NAND2_X1 g123 ( .A1(new_n260_), .A2(new_n178_), .ZN(new_n261_) );
  NAND3_X1 g124 ( .A1(new_n261_), .A2(new_n206_), .A3(new_n259_), .ZN(new_n262_) );
  INV_X1 g125 ( .A(new_n206_), .ZN(new_n263_) );
  NAND2_X1 g126 ( .A1(new_n261_), .A2(new_n259_), .ZN(new_n264_) );
  NAND2_X1 g127 ( .A1(new_n264_), .A2(new_n263_), .ZN(new_n265_) );
  NAND2_X1 g128 ( .A1(new_n265_), .A2(new_n262_), .ZN(new_n266_) );
  INV_X1 g129 ( .A(new_n266_), .ZN(new_n267_) );
  XNOR2_X1 g130 ( .A(G57GAT), .B(G71GAT), .ZN(new_n268_) );
  XNOR2_X1 g131 ( .A(new_n268_), .B(KEYINPUT13), .ZN(new_n269_) );
  INV_X1 g132 ( .A(new_n269_), .ZN(new_n270_) );
  XOR2_X1 g133 ( .A(G15GAT), .B(G22GAT), .Z(new_n271_) );
  XNOR2_X1 g134 ( .A(new_n271_), .B(G1GAT), .ZN(new_n272_) );
  XNOR2_X1 g135 ( .A(new_n270_), .B(new_n272_), .ZN(new_n273_) );
  XNOR2_X1 g136 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(new_n274_) );
  XNOR2_X1 g137 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n275_) );
  XNOR2_X1 g138 ( .A(new_n274_), .B(new_n275_), .ZN(new_n276_) );
  XNOR2_X1 g139 ( .A(G78GAT), .B(G155GAT), .ZN(new_n277_) );
  XNOR2_X1 g140 ( .A(G127GAT), .B(G211GAT), .ZN(new_n278_) );
  XNOR2_X1 g141 ( .A(new_n277_), .B(new_n278_), .ZN(new_n279_) );
  XNOR2_X1 g142 ( .A(new_n276_), .B(new_n279_), .ZN(new_n280_) );
  XNOR2_X1 g143 ( .A(new_n273_), .B(new_n280_), .ZN(new_n281_) );
  XNOR2_X1 g144 ( .A(new_n281_), .B(new_n212_), .ZN(new_n282_) );
  NAND2_X1 g145 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n283_) );
  XOR2_X1 g146 ( .A(new_n282_), .B(new_n283_), .Z(new_n284_) );
  NAND2_X1 g147 ( .A1(new_n267_), .A2(new_n284_), .ZN(new_n285_) );
  XOR2_X1 g148 ( .A(new_n285_), .B(KEYINPUT16), .Z(new_n286_) );
  AND2_X1 g149 ( .A1(new_n231_), .A2(new_n286_), .ZN(new_n287_) );
  XOR2_X1 g150 ( .A(G113GAT), .B(G197GAT), .Z(new_n288_) );
  XNOR2_X1 g151 ( .A(G29GAT), .B(G141GAT), .ZN(new_n289_) );
  XNOR2_X1 g152 ( .A(new_n288_), .B(new_n289_), .ZN(new_n290_) );
  XOR2_X1 g153 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(new_n291_) );
  XNOR2_X1 g154 ( .A(G8GAT), .B(G169GAT), .ZN(new_n292_) );
  XNOR2_X1 g155 ( .A(new_n291_), .B(new_n292_), .ZN(new_n293_) );
  XNOR2_X1 g156 ( .A(new_n290_), .B(new_n293_), .ZN(new_n294_) );
  XNOR2_X1 g157 ( .A(new_n272_), .B(new_n236_), .ZN(new_n295_) );
  XNOR2_X1 g158 ( .A(new_n294_), .B(new_n295_), .ZN(new_n296_) );
  XOR2_X1 g159 ( .A(G36GAT), .B(G50GAT), .Z(new_n297_) );
  NAND2_X1 g160 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n298_) );
  XNOR2_X1 g161 ( .A(new_n297_), .B(new_n298_), .ZN(new_n299_) );
  XNOR2_X1 g162 ( .A(new_n296_), .B(new_n299_), .ZN(new_n300_) );
  XNOR2_X1 g163 ( .A(G120GAT), .B(G204GAT), .ZN(new_n301_) );
  INV_X1 g164 ( .A(new_n301_), .ZN(new_n302_) );
  INV_X1 g165 ( .A(new_n208_), .ZN(new_n303_) );
  INV_X1 g166 ( .A(KEYINPUT32), .ZN(new_n304_) );
  NAND2_X1 g167 ( .A1(KEYINPUT33), .A2(KEYINPUT31), .ZN(new_n305_) );
  OR2_X1 g168 ( .A1(KEYINPUT33), .A2(KEYINPUT31), .ZN(new_n306_) );
  NAND2_X1 g169 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n307_) );
  NAND3_X1 g170 ( .A1(new_n306_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_) );
  XNOR2_X1 g171 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(new_n309_) );
  INV_X1 g172 ( .A(new_n307_), .ZN(new_n310_) );
  NAND2_X1 g173 ( .A1(new_n309_), .A2(new_n310_), .ZN(new_n311_) );
  NAND2_X1 g174 ( .A1(new_n311_), .A2(new_n308_), .ZN(new_n312_) );
  NAND2_X1 g175 ( .A1(new_n312_), .A2(new_n304_), .ZN(new_n313_) );
  NAND3_X1 g176 ( .A1(new_n311_), .A2(KEYINPUT32), .A3(new_n308_), .ZN(new_n314_) );
  NAND2_X1 g177 ( .A1(new_n238_), .A2(new_n242_), .ZN(new_n315_) );
  NAND2_X1 g178 ( .A1(new_n173_), .A2(new_n315_), .ZN(new_n316_) );
  NAND4_X1 g179 ( .A1(new_n171_), .A2(new_n238_), .A3(new_n172_), .A4(new_n242_), .ZN(new_n317_) );
  NAND4_X1 g180 ( .A1(new_n316_), .A2(new_n313_), .A3(new_n314_), .A4(new_n317_), .ZN(new_n318_) );
  NAND2_X1 g181 ( .A1(new_n313_), .A2(new_n314_), .ZN(new_n319_) );
  NAND2_X1 g182 ( .A1(new_n316_), .A2(new_n317_), .ZN(new_n320_) );
  NAND2_X1 g183 ( .A1(new_n320_), .A2(new_n319_), .ZN(new_n321_) );
  NAND3_X1 g184 ( .A1(new_n321_), .A2(new_n303_), .A3(new_n318_), .ZN(new_n322_) );
  NAND2_X1 g185 ( .A1(new_n321_), .A2(new_n318_), .ZN(new_n323_) );
  NAND2_X1 g186 ( .A1(new_n323_), .A2(new_n208_), .ZN(new_n324_) );
  NAND2_X1 g187 ( .A1(new_n324_), .A2(new_n322_), .ZN(new_n325_) );
  NAND2_X1 g188 ( .A1(new_n325_), .A2(new_n302_), .ZN(new_n326_) );
  NAND3_X1 g189 ( .A1(new_n324_), .A2(new_n301_), .A3(new_n322_), .ZN(new_n327_) );
  NAND2_X1 g190 ( .A1(new_n326_), .A2(new_n327_), .ZN(new_n328_) );
  NAND2_X1 g191 ( .A1(new_n328_), .A2(new_n269_), .ZN(new_n329_) );
  NAND3_X1 g192 ( .A1(new_n326_), .A2(new_n270_), .A3(new_n327_), .ZN(new_n330_) );
  AND3_X1 g193 ( .A1(new_n329_), .A2(new_n300_), .A3(new_n330_), .ZN(new_n331_) );
  AND2_X1 g194 ( .A1(new_n287_), .A2(new_n331_), .ZN(new_n332_) );
  NAND2_X1 g195 ( .A1(new_n332_), .A2(new_n158_), .ZN(new_n333_) );
  XNOR2_X1 g196 ( .A(new_n333_), .B(KEYINPUT34), .ZN(new_n334_) );
  XNOR2_X1 g197 ( .A(new_n334_), .B(G1GAT), .ZN(G1324GAT) );
  NAND2_X1 g198 ( .A1(new_n332_), .A2(new_n215_), .ZN(new_n336_) );
  XNOR2_X1 g199 ( .A(new_n336_), .B(G8GAT), .ZN(G1325GAT) );
  NAND2_X1 g200 ( .A1(new_n332_), .A2(new_n220_), .ZN(new_n338_) );
  XOR2_X1 g201 ( .A(G15GAT), .B(KEYINPUT35), .Z(new_n339_) );
  XNOR2_X1 g202 ( .A(new_n338_), .B(new_n339_), .ZN(G1326GAT) );
  INV_X1 g203 ( .A(new_n228_), .ZN(new_n341_) );
  NAND2_X1 g204 ( .A1(new_n332_), .A2(new_n341_), .ZN(new_n342_) );
  XNOR2_X1 g205 ( .A(new_n342_), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 g206 ( .A(KEYINPUT37), .ZN(new_n344_) );
  INV_X1 g207 ( .A(KEYINPUT36), .ZN(new_n345_) );
  NAND2_X1 g208 ( .A1(new_n266_), .A2(new_n345_), .ZN(new_n346_) );
  NAND3_X1 g209 ( .A1(new_n265_), .A2(KEYINPUT36), .A3(new_n262_), .ZN(new_n347_) );
  NAND2_X1 g210 ( .A1(new_n346_), .A2(new_n347_), .ZN(new_n348_) );
  NOR2_X1 g211 ( .A1(new_n348_), .A2(new_n284_), .ZN(new_n349_) );
  NAND2_X1 g212 ( .A1(new_n231_), .A2(new_n349_), .ZN(new_n350_) );
  NAND2_X1 g213 ( .A1(new_n350_), .A2(new_n344_), .ZN(new_n351_) );
  NAND3_X1 g214 ( .A1(new_n231_), .A2(KEYINPUT37), .A3(new_n349_), .ZN(new_n352_) );
  NAND4_X1 g215 ( .A1(new_n351_), .A2(KEYINPUT38), .A3(new_n331_), .A4(new_n352_), .ZN(new_n353_) );
  INV_X1 g216 ( .A(KEYINPUT38), .ZN(new_n354_) );
  NAND3_X1 g217 ( .A1(new_n351_), .A2(new_n331_), .A3(new_n352_), .ZN(new_n355_) );
  NAND2_X1 g218 ( .A1(new_n355_), .A2(new_n354_), .ZN(new_n356_) );
  NAND2_X1 g219 ( .A1(new_n356_), .A2(new_n353_), .ZN(new_n357_) );
  NAND2_X1 g220 ( .A1(new_n357_), .A2(new_n158_), .ZN(new_n358_) );
  XOR2_X1 g221 ( .A(G29GAT), .B(KEYINPUT39), .Z(new_n359_) );
  XNOR2_X1 g222 ( .A(new_n358_), .B(new_n359_), .ZN(G1328GAT) );
  NAND2_X1 g223 ( .A1(new_n357_), .A2(new_n215_), .ZN(new_n361_) );
  XNOR2_X1 g224 ( .A(new_n361_), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 g225 ( .A1(new_n357_), .A2(new_n220_), .ZN(new_n363_) );
  NAND2_X1 g226 ( .A1(new_n363_), .A2(KEYINPUT40), .ZN(new_n364_) );
  INV_X1 g227 ( .A(KEYINPUT40), .ZN(new_n365_) );
  NAND3_X1 g228 ( .A1(new_n357_), .A2(new_n365_), .A3(new_n220_), .ZN(new_n366_) );
  NAND2_X1 g229 ( .A1(new_n364_), .A2(new_n366_), .ZN(new_n367_) );
  NAND2_X1 g230 ( .A1(new_n367_), .A2(G43GAT), .ZN(new_n368_) );
  INV_X1 g231 ( .A(G43GAT), .ZN(new_n369_) );
  NAND3_X1 g232 ( .A1(new_n364_), .A2(new_n369_), .A3(new_n366_), .ZN(new_n370_) );
  NAND2_X1 g233 ( .A1(new_n368_), .A2(new_n370_), .ZN(G1330GAT) );
  NAND2_X1 g234 ( .A1(new_n357_), .A2(new_n341_), .ZN(new_n372_) );
  XNOR2_X1 g235 ( .A(new_n372_), .B(G50GAT), .ZN(G1331GAT) );
  NAND3_X1 g236 ( .A1(new_n329_), .A2(KEYINPUT41), .A3(new_n330_), .ZN(new_n374_) );
  INV_X1 g237 ( .A(KEYINPUT41), .ZN(new_n375_) );
  NAND2_X1 g238 ( .A1(new_n329_), .A2(new_n330_), .ZN(new_n376_) );
  NAND2_X1 g239 ( .A1(new_n376_), .A2(new_n375_), .ZN(new_n377_) );
  NAND2_X1 g240 ( .A1(new_n377_), .A2(new_n374_), .ZN(new_n378_) );
  INV_X1 g241 ( .A(new_n378_), .ZN(new_n379_) );
  NOR2_X1 g242 ( .A1(new_n379_), .A2(new_n300_), .ZN(new_n380_) );
  AND2_X1 g243 ( .A1(new_n287_), .A2(new_n380_), .ZN(new_n381_) );
  NAND2_X1 g244 ( .A1(new_n381_), .A2(new_n158_), .ZN(new_n382_) );
  XNOR2_X1 g245 ( .A(G57GAT), .B(KEYINPUT42), .ZN(new_n383_) );
  XNOR2_X1 g246 ( .A(new_n382_), .B(new_n383_), .ZN(G1332GAT) );
  NAND2_X1 g247 ( .A1(new_n381_), .A2(new_n215_), .ZN(new_n385_) );
  XNOR2_X1 g248 ( .A(new_n385_), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 g249 ( .A1(new_n381_), .A2(new_n220_), .ZN(new_n387_) );
  XNOR2_X1 g250 ( .A(new_n387_), .B(G71GAT), .ZN(G1334GAT) );
  NAND2_X1 g251 ( .A1(new_n381_), .A2(new_n341_), .ZN(new_n389_) );
  XOR2_X1 g252 ( .A(G78GAT), .B(KEYINPUT43), .Z(new_n390_) );
  XNOR2_X1 g253 ( .A(new_n389_), .B(new_n390_), .ZN(G1335GAT) );
  AND2_X1 g254 ( .A1(new_n351_), .A2(new_n352_), .ZN(new_n392_) );
  AND2_X1 g255 ( .A1(new_n392_), .A2(new_n380_), .ZN(new_n393_) );
  NAND2_X1 g256 ( .A1(new_n393_), .A2(new_n158_), .ZN(new_n394_) );
  XNOR2_X1 g257 ( .A(new_n394_), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 g258 ( .A1(new_n393_), .A2(new_n215_), .ZN(new_n396_) );
  XNOR2_X1 g259 ( .A(new_n396_), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 g260 ( .A1(new_n393_), .A2(new_n220_), .ZN(new_n398_) );
  XNOR2_X1 g261 ( .A(new_n398_), .B(G99GAT), .ZN(G1338GAT) );
  INV_X1 g262 ( .A(KEYINPUT44), .ZN(new_n400_) );
  AND3_X1 g263 ( .A1(new_n392_), .A2(new_n341_), .A3(new_n380_), .ZN(new_n401_) );
  OR2_X1 g264 ( .A1(new_n401_), .A2(new_n400_), .ZN(new_n402_) );
  NAND2_X1 g265 ( .A1(new_n401_), .A2(new_n400_), .ZN(new_n403_) );
  NAND2_X1 g266 ( .A1(new_n402_), .A2(new_n403_), .ZN(new_n404_) );
  NAND2_X1 g267 ( .A1(new_n404_), .A2(G106GAT), .ZN(new_n405_) );
  INV_X1 g268 ( .A(G106GAT), .ZN(new_n406_) );
  NAND3_X1 g269 ( .A1(new_n402_), .A2(new_n406_), .A3(new_n403_), .ZN(new_n407_) );
  NAND2_X1 g270 ( .A1(new_n405_), .A2(new_n407_), .ZN(G1339GAT) );
  INV_X1 g271 ( .A(KEYINPUT48), .ZN(new_n409_) );
  INV_X1 g272 ( .A(KEYINPUT47), .ZN(new_n410_) );
  NAND3_X1 g273 ( .A1(new_n378_), .A2(KEYINPUT46), .A3(new_n300_), .ZN(new_n411_) );
  INV_X1 g274 ( .A(KEYINPUT46), .ZN(new_n412_) );
  NAND2_X1 g275 ( .A1(new_n378_), .A2(new_n300_), .ZN(new_n413_) );
  NAND2_X1 g276 ( .A1(new_n413_), .A2(new_n412_), .ZN(new_n414_) );
  NOR2_X1 g277 ( .A1(new_n284_), .A2(new_n266_), .ZN(new_n415_) );
  NAND4_X1 g278 ( .A1(new_n414_), .A2(new_n410_), .A3(new_n411_), .A4(new_n415_), .ZN(new_n416_) );
  NAND3_X1 g279 ( .A1(new_n414_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n417_) );
  NAND2_X1 g280 ( .A1(new_n417_), .A2(KEYINPUT47), .ZN(new_n418_) );
  NAND3_X1 g281 ( .A1(new_n346_), .A2(new_n284_), .A3(new_n347_), .ZN(new_n419_) );
  NAND2_X1 g282 ( .A1(new_n419_), .A2(KEYINPUT45), .ZN(new_n420_) );
  INV_X1 g283 ( .A(KEYINPUT45), .ZN(new_n421_) );
  NAND4_X1 g284 ( .A1(new_n346_), .A2(new_n284_), .A3(new_n421_), .A4(new_n347_), .ZN(new_n422_) );
  NOR2_X1 g285 ( .A1(new_n376_), .A2(new_n300_), .ZN(new_n423_) );
  NAND3_X1 g286 ( .A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_) );
  NAND3_X1 g287 ( .A1(new_n418_), .A2(new_n416_), .A3(new_n424_), .ZN(new_n425_) );
  NAND2_X1 g288 ( .A1(new_n425_), .A2(new_n409_), .ZN(new_n426_) );
  NAND4_X1 g289 ( .A1(new_n418_), .A2(KEYINPUT48), .A3(new_n424_), .A4(new_n416_), .ZN(new_n427_) );
  AND3_X1 g290 ( .A1(new_n426_), .A2(new_n229_), .A3(new_n427_), .ZN(new_n428_) );
  NOR2_X1 g291 ( .A1(new_n341_), .A2(new_n200_), .ZN(new_n429_) );
  NAND2_X1 g292 ( .A1(new_n428_), .A2(new_n429_), .ZN(new_n430_) );
  INV_X1 g293 ( .A(new_n430_), .ZN(new_n431_) );
  NAND2_X1 g294 ( .A1(new_n431_), .A2(new_n300_), .ZN(new_n432_) );
  XNOR2_X1 g295 ( .A(new_n432_), .B(G113GAT), .ZN(G1340GAT) );
  NOR2_X1 g296 ( .A1(new_n430_), .A2(new_n379_), .ZN(new_n434_) );
  XNOR2_X1 g297 ( .A(G120GAT), .B(KEYINPUT49), .ZN(new_n435_) );
  XNOR2_X1 g298 ( .A(new_n434_), .B(new_n435_), .ZN(G1341GAT) );
  NAND2_X1 g299 ( .A1(new_n431_), .A2(new_n284_), .ZN(new_n437_) );
  XNOR2_X1 g300 ( .A(new_n437_), .B(KEYINPUT50), .ZN(new_n438_) );
  XNOR2_X1 g301 ( .A(new_n438_), .B(G127GAT), .ZN(G1342GAT) );
  NOR2_X1 g302 ( .A1(new_n430_), .A2(new_n267_), .ZN(new_n440_) );
  XNOR2_X1 g303 ( .A(G134GAT), .B(KEYINPUT51), .ZN(new_n441_) );
  XNOR2_X1 g304 ( .A(new_n440_), .B(new_n441_), .ZN(G1343GAT) );
  NAND2_X1 g305 ( .A1(new_n428_), .A2(new_n205_), .ZN(new_n443_) );
  INV_X1 g306 ( .A(new_n443_), .ZN(new_n444_) );
  NAND2_X1 g307 ( .A1(new_n444_), .A2(new_n300_), .ZN(new_n445_) );
  XNOR2_X1 g308 ( .A(new_n445_), .B(G141GAT), .ZN(G1344GAT) );
  NAND2_X1 g309 ( .A1(new_n444_), .A2(new_n378_), .ZN(new_n447_) );
  XNOR2_X1 g310 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(new_n448_) );
  XOR2_X1 g311 ( .A(new_n447_), .B(new_n448_), .Z(new_n449_) );
  XNOR2_X1 g312 ( .A(new_n449_), .B(G148GAT), .ZN(G1345GAT) );
  NAND2_X1 g313 ( .A1(new_n444_), .A2(new_n284_), .ZN(new_n451_) );
  XNOR2_X1 g314 ( .A(new_n451_), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 g315 ( .A1(new_n444_), .A2(new_n266_), .ZN(new_n453_) );
  XNOR2_X1 g316 ( .A(new_n453_), .B(G162GAT), .ZN(G1347GAT) );
  NAND3_X1 g317 ( .A1(new_n426_), .A2(new_n215_), .A3(new_n427_), .ZN(new_n455_) );
  NAND2_X1 g318 ( .A1(new_n455_), .A2(KEYINPUT54), .ZN(new_n456_) );
  INV_X1 g319 ( .A(KEYINPUT54), .ZN(new_n457_) );
  NAND4_X1 g320 ( .A1(new_n426_), .A2(new_n457_), .A3(new_n215_), .A4(new_n427_), .ZN(new_n458_) );
  NAND4_X1 g321 ( .A1(new_n456_), .A2(new_n157_), .A3(new_n219_), .A4(new_n458_), .ZN(new_n459_) );
  NAND2_X1 g322 ( .A1(new_n459_), .A2(KEYINPUT55), .ZN(new_n460_) );
  INV_X1 g323 ( .A(KEYINPUT55), .ZN(new_n461_) );
  AND2_X1 g324 ( .A1(new_n458_), .A2(new_n219_), .ZN(new_n462_) );
  NAND4_X1 g325 ( .A1(new_n462_), .A2(new_n461_), .A3(new_n157_), .A4(new_n456_), .ZN(new_n463_) );
  NAND2_X1 g326 ( .A1(new_n460_), .A2(new_n463_), .ZN(new_n464_) );
  NAND3_X1 g327 ( .A1(new_n464_), .A2(new_n220_), .A3(new_n300_), .ZN(new_n465_) );
  XNOR2_X1 g328 ( .A(new_n465_), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 g329 ( .A(G176GAT), .ZN(new_n467_) );
  NAND3_X1 g330 ( .A1(new_n464_), .A2(new_n220_), .A3(new_n378_), .ZN(new_n468_) );
  XOR2_X1 g331 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(new_n469_) );
  INV_X1 g332 ( .A(new_n469_), .ZN(new_n470_) );
  NAND2_X1 g333 ( .A1(new_n468_), .A2(new_n470_), .ZN(new_n471_) );
  NAND4_X1 g334 ( .A1(new_n464_), .A2(new_n220_), .A3(new_n378_), .A4(new_n469_), .ZN(new_n472_) );
  NAND2_X1 g335 ( .A1(new_n471_), .A2(new_n472_), .ZN(new_n473_) );
  NAND2_X1 g336 ( .A1(new_n473_), .A2(new_n467_), .ZN(new_n474_) );
  NAND3_X1 g337 ( .A1(new_n471_), .A2(G176GAT), .A3(new_n472_), .ZN(new_n475_) );
  NAND2_X1 g338 ( .A1(new_n474_), .A2(new_n475_), .ZN(G1349GAT) );
  NAND3_X1 g339 ( .A1(new_n464_), .A2(new_n220_), .A3(new_n284_), .ZN(new_n477_) );
  XNOR2_X1 g340 ( .A(new_n477_), .B(G183GAT), .ZN(G1350GAT) );
  NAND3_X1 g341 ( .A1(new_n464_), .A2(new_n220_), .A3(new_n266_), .ZN(new_n479_) );
  XNOR2_X1 g342 ( .A(G190GAT), .B(KEYINPUT58), .ZN(new_n480_) );
  XNOR2_X1 g343 ( .A(new_n479_), .B(new_n480_), .ZN(G1351GAT) );
  AND4_X1 g344 ( .A1(new_n157_), .A2(new_n456_), .A3(new_n205_), .A4(new_n458_), .ZN(new_n482_) );
  NAND2_X1 g345 ( .A1(new_n482_), .A2(new_n300_), .ZN(new_n483_) );
  XNOR2_X1 g346 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(new_n484_) );
  INV_X1 g347 ( .A(new_n484_), .ZN(new_n485_) );
  XNOR2_X1 g348 ( .A(new_n483_), .B(new_n485_), .ZN(new_n486_) );
  XNOR2_X1 g349 ( .A(new_n486_), .B(G197GAT), .ZN(G1352GAT) );
  NAND2_X1 g350 ( .A1(new_n482_), .A2(new_n376_), .ZN(new_n488_) );
  XOR2_X1 g351 ( .A(G204GAT), .B(KEYINPUT61), .Z(new_n489_) );
  XNOR2_X1 g352 ( .A(new_n488_), .B(new_n489_), .ZN(G1353GAT) );
  NAND2_X1 g353 ( .A1(new_n482_), .A2(new_n284_), .ZN(new_n491_) );
  XNOR2_X1 g354 ( .A(new_n491_), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 g355 ( .A(new_n348_), .ZN(new_n493_) );
  NAND2_X1 g356 ( .A1(new_n482_), .A2(new_n493_), .ZN(new_n494_) );
  XNOR2_X1 g357 ( .A(new_n494_), .B(KEYINPUT62), .ZN(new_n495_) );
  XNOR2_X1 g358 ( .A(new_n495_), .B(G218GAT), .ZN(G1355GAT) );
endmodule


