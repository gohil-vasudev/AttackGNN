module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n339_, new_n365_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n456_, new_n246_, new_n266_, new_n367_, new_n542_, new_n548_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n240_, new_n413_, new_n442_, new_n642_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n272_, new_n282_, new_n634_, new_n414_, new_n315_, new_n326_, new_n554_, new_n648_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n346_, new_n396_, new_n438_, new_n208_, new_n632_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n409_, new_n457_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n562_, new_n525_, new_n578_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n300_, new_n411_, new_n605_, new_n407_, new_n480_, new_n625_, new_n592_, new_n558_, new_n219_, new_n583_, new_n231_, new_n313_, new_n382_, new_n239_, new_n617_, new_n522_, new_n588_, new_n428_, new_n360_, new_n546_, new_n612_, new_n302_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n590_, new_n417_, new_n591_, new_n332_, new_n631_, new_n453_, new_n516_, new_n563_, new_n440_, new_n593_, new_n252_, new_n585_, new_n312_, new_n535_, new_n372_, new_n242_, new_n527_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n574_, new_n319_, new_n640_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n226_, new_n373_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n573_, new_n405_;

not g000 ( new_n202_, N1 );
not g001 ( new_n203_, keyIn_0_72 );
xnor g002 ( new_n204_, N1, N17 );
xnor g003 ( new_n205_, new_n204_, keyIn_0_24 );
xor g004 ( new_n206_, N33, N49 );
xnor g005 ( new_n207_, new_n206_, keyIn_0_25 );
xnor g006 ( new_n208_, new_n207_, new_n205_ );
xor g007 ( new_n209_, new_n208_, keyIn_0_48 );
and g008 ( new_n210_, N129, N137 );
xnor g009 ( new_n211_, new_n210_, keyIn_0_16 );
xnor g010 ( new_n212_, N73, N77 );
xnor g011 ( new_n213_, new_n212_, keyIn_0_8 );
xnor g012 ( new_n214_, N65, N69 );
xnor g013 ( new_n215_, new_n214_, keyIn_0_9 );
xor g014 ( new_n216_, new_n213_, new_n215_ );
xnor g015 ( new_n217_, new_n216_, keyIn_0_44 );
not g016 ( new_n218_, keyIn_0_10 );
xor g017 ( new_n219_, N81, N85 );
or g018 ( new_n220_, new_n219_, new_n218_ );
not g019 ( new_n221_, N81 );
not g020 ( new_n222_, N85 );
and g021 ( new_n223_, new_n221_, new_n222_ );
and g022 ( new_n224_, N81, N85 );
or g023 ( new_n225_, new_n224_, keyIn_0_10 );
or g024 ( new_n226_, new_n225_, new_n223_ );
and g025 ( new_n227_, new_n226_, new_n220_ );
not g026 ( new_n228_, keyIn_0_11 );
xor g027 ( new_n229_, N89, N93 );
or g028 ( new_n230_, new_n229_, new_n228_ );
not g029 ( new_n231_, N89 );
not g030 ( new_n232_, N93 );
and g031 ( new_n233_, new_n231_, new_n232_ );
and g032 ( new_n234_, N89, N93 );
or g033 ( new_n235_, new_n234_, keyIn_0_11 );
or g034 ( new_n236_, new_n235_, new_n233_ );
and g035 ( new_n237_, new_n236_, new_n230_ );
xnor g036 ( new_n238_, new_n227_, new_n237_ );
xnor g037 ( new_n239_, new_n238_, keyIn_0_45 );
xnor g038 ( new_n240_, new_n239_, new_n217_ );
xnor g039 ( new_n241_, new_n240_, keyIn_0_60 );
xnor g040 ( new_n242_, new_n241_, new_n211_ );
xnor g041 ( new_n243_, new_n242_, keyIn_0_64 );
xnor g042 ( new_n244_, new_n243_, new_n209_ );
xnor g043 ( new_n245_, new_n244_, new_n203_ );
not g044 ( new_n246_, keyIn_0_112 );
not g045 ( new_n247_, keyIn_0_105 );
xnor g046 ( new_n248_, N5, N21 );
xnor g047 ( new_n249_, new_n248_, keyIn_0_26 );
xor g048 ( new_n250_, N37, N53 );
xnor g049 ( new_n251_, new_n250_, keyIn_0_27 );
xnor g050 ( new_n252_, new_n251_, new_n249_ );
xnor g051 ( new_n253_, new_n252_, keyIn_0_49 );
xor g052 ( new_n254_, N113, N117 );
xnor g053 ( new_n255_, new_n254_, keyIn_0_14 );
xor g054 ( new_n256_, N121, N125 );
xnor g055 ( new_n257_, new_n256_, keyIn_0_15 );
xor g056 ( new_n258_, new_n255_, new_n257_ );
xnor g057 ( new_n259_, new_n258_, keyIn_0_47 );
not g058 ( new_n260_, keyIn_0_46 );
xnor g059 ( new_n261_, N97, N101 );
xnor g060 ( new_n262_, new_n261_, keyIn_0_12 );
xor g061 ( new_n263_, N105, N109 );
xnor g062 ( new_n264_, new_n263_, keyIn_0_13 );
xnor g063 ( new_n265_, new_n264_, new_n262_ );
xnor g064 ( new_n266_, new_n265_, new_n260_ );
xnor g065 ( new_n267_, new_n259_, new_n266_ );
xnor g066 ( new_n268_, new_n267_, keyIn_0_61 );
and g067 ( new_n269_, N130, N137 );
xnor g068 ( new_n270_, new_n269_, keyIn_0_17 );
xnor g069 ( new_n271_, new_n268_, new_n270_ );
xnor g070 ( new_n272_, new_n271_, keyIn_0_65 );
xnor g071 ( new_n273_, new_n272_, new_n253_ );
xnor g072 ( new_n274_, new_n273_, keyIn_0_73 );
and g073 ( new_n275_, new_n274_, keyIn_0_84 );
not g074 ( new_n276_, new_n275_ );
or g075 ( new_n277_, new_n274_, keyIn_0_84 );
not g076 ( new_n278_, keyIn_0_74 );
xor g077 ( new_n279_, N9, N25 );
xor g078 ( new_n280_, new_n279_, keyIn_0_28 );
xor g079 ( new_n281_, N41, N57 );
xnor g080 ( new_n282_, new_n281_, keyIn_0_29 );
xnor g081 ( new_n283_, new_n280_, new_n282_ );
xor g082 ( new_n284_, new_n283_, keyIn_0_50 );
and g083 ( new_n285_, N131, N137 );
xor g084 ( new_n286_, new_n285_, keyIn_0_18 );
xnor g085 ( new_n287_, new_n217_, new_n266_ );
xnor g086 ( new_n288_, new_n287_, keyIn_0_62 );
xnor g087 ( new_n289_, new_n288_, new_n286_ );
xnor g088 ( new_n290_, new_n289_, keyIn_0_66 );
xnor g089 ( new_n291_, new_n290_, new_n284_ );
xnor g090 ( new_n292_, new_n291_, new_n278_ );
and g091 ( new_n293_, new_n277_, new_n292_ );
and g092 ( new_n294_, new_n293_, new_n276_ );
xor g093 ( new_n295_, N13, N29 );
xnor g094 ( new_n296_, new_n295_, keyIn_0_30 );
xnor g095 ( new_n297_, N45, N61 );
xnor g096 ( new_n298_, new_n297_, keyIn_0_31 );
xnor g097 ( new_n299_, new_n296_, new_n298_ );
xnor g098 ( new_n300_, new_n299_, keyIn_0_51 );
xnor g099 ( new_n301_, new_n239_, new_n259_ );
xnor g100 ( new_n302_, new_n301_, keyIn_0_63 );
and g101 ( new_n303_, N132, N137 );
xnor g102 ( new_n304_, new_n303_, keyIn_0_19 );
xnor g103 ( new_n305_, new_n302_, new_n304_ );
xnor g104 ( new_n306_, new_n305_, keyIn_0_67 );
xnor g105 ( new_n307_, new_n306_, new_n300_ );
xnor g106 ( new_n308_, new_n307_, keyIn_0_75 );
xnor g107 ( new_n309_, new_n308_, keyIn_0_85 );
not g108 ( new_n310_, keyIn_0_83 );
xnor g109 ( new_n311_, new_n245_, new_n310_ );
not g110 ( new_n312_, new_n311_ );
and g111 ( new_n313_, new_n312_, new_n309_ );
and g112 ( new_n314_, new_n313_, new_n294_ );
or g113 ( new_n315_, new_n314_, new_n247_ );
not g114 ( new_n316_, new_n292_ );
and g115 ( new_n317_, new_n316_, keyIn_0_82 );
not g116 ( new_n318_, keyIn_0_82 );
and g117 ( new_n319_, new_n292_, new_n318_ );
or g118 ( new_n320_, new_n319_, new_n308_ );
or g119 ( new_n321_, new_n320_, new_n317_ );
not g120 ( new_n322_, keyIn_0_73 );
xnor g121 ( new_n323_, new_n273_, new_n322_ );
xnor g122 ( new_n324_, new_n323_, keyIn_0_81 );
xnor g123 ( new_n325_, new_n245_, keyIn_0_80 );
or g124 ( new_n326_, new_n325_, new_n324_ );
or g125 ( new_n327_, new_n326_, new_n321_ );
or g126 ( new_n328_, new_n327_, keyIn_0_104 );
and g127 ( new_n329_, new_n315_, new_n328_ );
not g128 ( new_n330_, keyIn_0_104 );
not g129 ( new_n331_, new_n321_ );
not g130 ( new_n332_, new_n326_ );
and g131 ( new_n333_, new_n332_, new_n331_ );
or g132 ( new_n334_, new_n333_, new_n330_ );
not g133 ( new_n335_, keyIn_0_84 );
and g134 ( new_n336_, new_n323_, new_n335_ );
or g135 ( new_n337_, new_n336_, new_n316_ );
or g136 ( new_n338_, new_n337_, new_n275_ );
xor g137 ( new_n339_, new_n307_, keyIn_0_75 );
xnor g138 ( new_n340_, new_n339_, keyIn_0_85 );
or g139 ( new_n341_, new_n340_, new_n311_ );
or g140 ( new_n342_, new_n341_, new_n338_ );
or g141 ( new_n343_, new_n342_, keyIn_0_105 );
and g142 ( new_n344_, new_n343_, new_n334_ );
and g143 ( new_n345_, new_n344_, new_n329_ );
and g144 ( new_n346_, new_n323_, keyIn_0_89 );
xor g145 ( new_n347_, new_n292_, keyIn_0_90 );
or g146 ( new_n348_, new_n347_, new_n346_ );
not g147 ( new_n349_, new_n245_ );
not g148 ( new_n350_, keyIn_0_89 );
and g149 ( new_n351_, new_n274_, new_n350_ );
or g150 ( new_n352_, new_n351_, new_n349_ );
xor g151 ( new_n353_, new_n308_, keyIn_0_91 );
or g152 ( new_n354_, new_n353_, new_n352_ );
or g153 ( new_n355_, new_n354_, new_n348_ );
xnor g154 ( new_n356_, new_n355_, keyIn_0_107 );
not g155 ( new_n357_, keyIn_0_88 );
or g156 ( new_n358_, new_n339_, new_n357_ );
xnor g157 ( new_n359_, new_n292_, keyIn_0_87 );
and g158 ( new_n360_, new_n358_, new_n359_ );
or g159 ( new_n361_, new_n308_, keyIn_0_88 );
and g160 ( new_n362_, new_n361_, new_n323_ );
xor g161 ( new_n363_, new_n245_, keyIn_0_86 );
and g162 ( new_n364_, new_n362_, new_n363_ );
and g163 ( new_n365_, new_n364_, new_n360_ );
xor g164 ( new_n366_, new_n365_, keyIn_0_106 );
and g165 ( new_n367_, new_n366_, new_n356_ );
and g166 ( new_n368_, new_n345_, new_n367_ );
xnor g167 ( new_n369_, new_n368_, new_n246_ );
not g168 ( new_n370_, keyIn_0_79 );
xnor g169 ( new_n371_, N77, N93 );
xnor g170 ( new_n372_, new_n371_, keyIn_0_38 );
xor g171 ( new_n373_, N109, N125 );
xnor g172 ( new_n374_, new_n373_, keyIn_0_39 );
xnor g173 ( new_n375_, new_n374_, new_n372_ );
xnor g174 ( new_n376_, new_n375_, keyIn_0_55 );
and g175 ( new_n377_, N136, N137 );
xor g176 ( new_n378_, new_n377_, keyIn_0_23 );
not g177 ( new_n379_, keyIn_0_7 );
xor g178 ( new_n380_, N57, N61 );
or g179 ( new_n381_, new_n380_, new_n379_ );
not g180 ( new_n382_, N57 );
not g181 ( new_n383_, N61 );
and g182 ( new_n384_, new_n382_, new_n383_ );
and g183 ( new_n385_, N57, N61 );
or g184 ( new_n386_, new_n385_, keyIn_0_7 );
or g185 ( new_n387_, new_n386_, new_n384_ );
and g186 ( new_n388_, new_n387_, new_n381_ );
xnor g187 ( new_n389_, N49, N53 );
xnor g188 ( new_n390_, new_n389_, keyIn_0_6 );
xnor g189 ( new_n391_, new_n388_, new_n390_ );
xnor g190 ( new_n392_, new_n391_, keyIn_0_43 );
xnor g191 ( new_n393_, N17, N21 );
xnor g192 ( new_n394_, new_n393_, keyIn_0_2 );
xor g193 ( new_n395_, N25, N29 );
xnor g194 ( new_n396_, new_n395_, keyIn_0_3 );
xnor g195 ( new_n397_, new_n396_, new_n394_ );
xor g196 ( new_n398_, new_n397_, keyIn_0_41 );
xnor g197 ( new_n399_, new_n392_, new_n398_ );
xnor g198 ( new_n400_, new_n399_, keyIn_0_59 );
xnor g199 ( new_n401_, new_n400_, new_n378_ );
xnor g200 ( new_n402_, new_n401_, keyIn_0_71 );
xnor g201 ( new_n403_, new_n402_, new_n376_ );
xnor g202 ( new_n404_, new_n403_, new_n370_ );
not g203 ( new_n405_, keyIn_0_78 );
xor g204 ( new_n406_, N73, N89 );
xnor g205 ( new_n407_, new_n406_, keyIn_0_36 );
xor g206 ( new_n408_, N105, N121 );
xnor g207 ( new_n409_, new_n408_, keyIn_0_37 );
xnor g208 ( new_n410_, new_n407_, new_n409_ );
xnor g209 ( new_n411_, new_n410_, keyIn_0_54 );
not g210 ( new_n412_, keyIn_0_58 );
not g211 ( new_n413_, N5 );
and g212 ( new_n414_, new_n202_, new_n413_ );
and g213 ( new_n415_, N1, N5 );
or g214 ( new_n416_, new_n415_, keyIn_0_0 );
or g215 ( new_n417_, new_n416_, new_n414_ );
not g216 ( new_n418_, keyIn_0_0 );
xor g217 ( new_n419_, N1, N5 );
or g218 ( new_n420_, new_n419_, new_n418_ );
and g219 ( new_n421_, new_n417_, new_n420_ );
xnor g220 ( new_n422_, N9, N13 );
xnor g221 ( new_n423_, new_n422_, keyIn_0_1 );
xnor g222 ( new_n424_, new_n421_, new_n423_ );
xnor g223 ( new_n425_, new_n424_, keyIn_0_40 );
not g224 ( new_n426_, keyIn_0_42 );
not g225 ( new_n427_, keyIn_0_5 );
xor g226 ( new_n428_, N41, N45 );
or g227 ( new_n429_, new_n428_, new_n427_ );
not g228 ( new_n430_, N41 );
not g229 ( new_n431_, N45 );
and g230 ( new_n432_, new_n430_, new_n431_ );
and g231 ( new_n433_, N41, N45 );
or g232 ( new_n434_, new_n433_, keyIn_0_5 );
or g233 ( new_n435_, new_n434_, new_n432_ );
and g234 ( new_n436_, new_n435_, new_n429_ );
xnor g235 ( new_n437_, N33, N37 );
xnor g236 ( new_n438_, new_n437_, keyIn_0_4 );
xnor g237 ( new_n439_, new_n436_, new_n438_ );
xnor g238 ( new_n440_, new_n439_, new_n426_ );
xnor g239 ( new_n441_, new_n425_, new_n440_ );
xnor g240 ( new_n442_, new_n441_, new_n412_ );
and g241 ( new_n443_, N135, N137 );
xor g242 ( new_n444_, new_n443_, keyIn_0_22 );
xnor g243 ( new_n445_, new_n442_, new_n444_ );
xnor g244 ( new_n446_, new_n445_, keyIn_0_70 );
xnor g245 ( new_n447_, new_n446_, new_n411_ );
xnor g246 ( new_n448_, new_n447_, new_n405_ );
and g247 ( new_n449_, new_n448_, new_n404_ );
and g248 ( new_n450_, new_n369_, new_n449_ );
not g249 ( new_n451_, keyIn_0_77 );
xor g250 ( new_n452_, N101, N117 );
xor g251 ( new_n453_, new_n452_, keyIn_0_35 );
xor g252 ( new_n454_, N69, N85 );
xnor g253 ( new_n455_, new_n454_, keyIn_0_34 );
xnor g254 ( new_n456_, new_n453_, new_n455_ );
xnor g255 ( new_n457_, new_n456_, keyIn_0_53 );
and g256 ( new_n458_, N134, N137 );
xnor g257 ( new_n459_, new_n458_, keyIn_0_21 );
xnor g258 ( new_n460_, new_n392_, new_n440_ );
xnor g259 ( new_n461_, new_n460_, keyIn_0_57 );
xnor g260 ( new_n462_, new_n461_, new_n459_ );
xnor g261 ( new_n463_, new_n462_, keyIn_0_69 );
xnor g262 ( new_n464_, new_n463_, new_n457_ );
xnor g263 ( new_n465_, new_n464_, new_n451_ );
not g264 ( new_n466_, new_n465_ );
and g265 ( new_n467_, N133, N137 );
xnor g266 ( new_n468_, new_n467_, keyIn_0_20 );
xnor g267 ( new_n469_, new_n425_, new_n398_ );
xnor g268 ( new_n470_, new_n469_, keyIn_0_56 );
xnor g269 ( new_n471_, new_n470_, new_n468_ );
xnor g270 ( new_n472_, new_n471_, keyIn_0_68 );
xor g271 ( new_n473_, N65, N81 );
xnor g272 ( new_n474_, new_n473_, keyIn_0_32 );
xor g273 ( new_n475_, N97, N113 );
xnor g274 ( new_n476_, new_n475_, keyIn_0_33 );
xnor g275 ( new_n477_, new_n474_, new_n476_ );
xnor g276 ( new_n478_, new_n477_, keyIn_0_52 );
xnor g277 ( new_n479_, new_n472_, new_n478_ );
xnor g278 ( new_n480_, new_n479_, keyIn_0_76 );
and g279 ( new_n481_, new_n466_, new_n480_ );
and g280 ( new_n482_, new_n450_, new_n481_ );
xor g281 ( new_n483_, new_n482_, keyIn_0_114 );
and g282 ( new_n484_, new_n483_, new_n245_ );
xnor g283 ( N724, new_n484_, new_n202_ );
and g284 ( new_n486_, new_n483_, new_n323_ );
xnor g285 ( N725, new_n486_, new_n413_ );
not g286 ( new_n488_, N9 );
and g287 ( new_n489_, new_n483_, new_n292_ );
xnor g288 ( N726, new_n489_, new_n488_ );
not g289 ( new_n491_, N13 );
and g290 ( new_n492_, new_n483_, new_n339_ );
xnor g291 ( N727, new_n492_, new_n491_ );
xnor g292 ( new_n494_, new_n403_, keyIn_0_79 );
xnor g293 ( new_n495_, new_n447_, keyIn_0_78 );
and g294 ( new_n496_, new_n495_, new_n494_ );
and g295 ( new_n497_, new_n481_, new_n496_ );
and g296 ( new_n498_, new_n369_, new_n497_ );
xnor g297 ( new_n499_, new_n498_, keyIn_0_115 );
and g298 ( new_n500_, new_n499_, new_n245_ );
xor g299 ( N728, new_n500_, N17 );
and g300 ( new_n502_, new_n499_, new_n323_ );
xor g301 ( N729, new_n502_, N21 );
and g302 ( new_n504_, new_n499_, new_n292_ );
xor g303 ( N730, new_n504_, N25 );
and g304 ( new_n506_, new_n499_, new_n339_ );
xor g305 ( N731, new_n506_, N29 );
not g306 ( new_n508_, new_n480_ );
and g307 ( new_n509_, new_n508_, new_n465_ );
and g308 ( new_n510_, new_n450_, new_n509_ );
xnor g309 ( new_n511_, new_n510_, keyIn_0_116 );
and g310 ( new_n512_, new_n511_, new_n245_ );
xor g311 ( N732, new_n512_, N33 );
and g312 ( new_n514_, new_n511_, new_n323_ );
xor g313 ( N733, new_n514_, N37 );
and g314 ( new_n516_, new_n511_, new_n292_ );
xnor g315 ( N734, new_n516_, new_n430_ );
and g316 ( new_n518_, new_n511_, new_n339_ );
xnor g317 ( N735, new_n518_, new_n431_ );
and g318 ( new_n520_, new_n509_, new_n496_ );
and g319 ( new_n521_, new_n369_, new_n520_ );
xnor g320 ( new_n522_, new_n521_, keyIn_0_117 );
and g321 ( new_n523_, new_n522_, new_n245_ );
xor g322 ( N736, new_n523_, N49 );
and g323 ( new_n525_, new_n522_, new_n323_ );
xor g324 ( N737, new_n525_, N53 );
and g325 ( new_n527_, new_n522_, new_n292_ );
xnor g326 ( N738, new_n527_, new_n382_ );
and g327 ( new_n529_, new_n522_, new_n339_ );
xnor g328 ( new_n530_, new_n529_, keyIn_0_122 );
xnor g329 ( N739, new_n530_, N61 );
not g330 ( new_n532_, N65 );
not g331 ( new_n533_, keyIn_0_118 );
and g332 ( new_n534_, new_n308_, new_n292_ );
and g333 ( new_n535_, new_n245_, new_n274_ );
and g334 ( new_n536_, new_n534_, new_n535_ );
not g335 ( new_n537_, keyIn_0_113 );
not g336 ( new_n538_, keyIn_0_97 );
and g337 ( new_n539_, new_n404_, new_n538_ );
not g338 ( new_n540_, new_n539_ );
or g339 ( new_n541_, new_n404_, new_n538_ );
and g340 ( new_n542_, new_n541_, new_n448_ );
and g341 ( new_n543_, new_n542_, new_n540_ );
xnor g342 ( new_n544_, new_n480_, keyIn_0_95 );
not g343 ( new_n545_, new_n544_ );
xnor g344 ( new_n546_, new_n465_, keyIn_0_96 );
not g345 ( new_n547_, new_n546_ );
and g346 ( new_n548_, new_n547_, new_n545_ );
and g347 ( new_n549_, new_n548_, new_n543_ );
or g348 ( new_n550_, new_n549_, keyIn_0_109 );
and g349 ( new_n551_, new_n495_, keyIn_0_99 );
not g350 ( new_n552_, new_n551_ );
or g351 ( new_n553_, new_n495_, keyIn_0_99 );
not g352 ( new_n554_, keyIn_0_100 );
or g353 ( new_n555_, new_n404_, new_n554_ );
and g354 ( new_n556_, new_n553_, new_n555_ );
and g355 ( new_n557_, new_n556_, new_n552_ );
or g356 ( new_n558_, new_n494_, keyIn_0_100 );
and g357 ( new_n559_, new_n558_, new_n465_ );
xnor g358 ( new_n560_, new_n480_, keyIn_0_98 );
not g359 ( new_n561_, new_n560_ );
and g360 ( new_n562_, new_n561_, new_n559_ );
and g361 ( new_n563_, new_n557_, new_n562_ );
or g362 ( new_n564_, new_n563_, keyIn_0_110 );
and g363 ( new_n565_, new_n550_, new_n564_ );
not g364 ( new_n566_, keyIn_0_109 );
and g365 ( new_n567_, new_n494_, keyIn_0_97 );
or g366 ( new_n568_, new_n567_, new_n495_ );
or g367 ( new_n569_, new_n568_, new_n539_ );
or g368 ( new_n570_, new_n546_, new_n544_ );
or g369 ( new_n571_, new_n569_, new_n570_ );
or g370 ( new_n572_, new_n571_, new_n566_ );
not g371 ( new_n573_, keyIn_0_110 );
not g372 ( new_n574_, keyIn_0_99 );
and g373 ( new_n575_, new_n448_, new_n574_ );
and g374 ( new_n576_, new_n494_, keyIn_0_100 );
or g375 ( new_n577_, new_n575_, new_n576_ );
or g376 ( new_n578_, new_n577_, new_n551_ );
and g377 ( new_n579_, new_n404_, new_n554_ );
or g378 ( new_n580_, new_n579_, new_n466_ );
or g379 ( new_n581_, new_n580_, new_n560_ );
or g380 ( new_n582_, new_n578_, new_n581_ );
or g381 ( new_n583_, new_n582_, new_n573_ );
and g382 ( new_n584_, new_n583_, new_n572_ );
and g383 ( new_n585_, new_n584_, new_n565_ );
or g384 ( new_n586_, new_n494_, keyIn_0_103 );
xor g385 ( new_n587_, new_n465_, keyIn_0_101 );
and g386 ( new_n588_, new_n587_, new_n586_ );
or g387 ( new_n589_, new_n495_, keyIn_0_102 );
and g388 ( new_n590_, new_n589_, new_n480_ );
not g389 ( new_n591_, keyIn_0_102 );
or g390 ( new_n592_, new_n448_, new_n591_ );
not g391 ( new_n593_, keyIn_0_103 );
or g392 ( new_n594_, new_n404_, new_n593_ );
and g393 ( new_n595_, new_n592_, new_n594_ );
and g394 ( new_n596_, new_n590_, new_n595_ );
and g395 ( new_n597_, new_n596_, new_n588_ );
xnor g396 ( new_n598_, new_n597_, keyIn_0_111 );
or g397 ( new_n599_, new_n508_, keyIn_0_92 );
not g398 ( new_n600_, keyIn_0_92 );
or g399 ( new_n601_, new_n480_, new_n600_ );
and g400 ( new_n602_, new_n601_, new_n494_ );
and g401 ( new_n603_, new_n602_, new_n599_ );
xnor g402 ( new_n604_, new_n495_, keyIn_0_94 );
xnor g403 ( new_n605_, new_n465_, keyIn_0_93 );
and g404 ( new_n606_, new_n604_, new_n605_ );
and g405 ( new_n607_, new_n603_, new_n606_ );
xor g406 ( new_n608_, new_n607_, keyIn_0_108 );
and g407 ( new_n609_, new_n608_, new_n598_ );
and g408 ( new_n610_, new_n585_, new_n609_ );
xnor g409 ( new_n611_, new_n610_, new_n537_ );
and g410 ( new_n612_, new_n611_, new_n536_ );
xnor g411 ( new_n613_, new_n612_, new_n533_ );
and g412 ( new_n614_, new_n613_, new_n480_ );
xnor g413 ( new_n615_, new_n614_, keyIn_0_123 );
xnor g414 ( N740, new_n615_, new_n532_ );
not g415 ( new_n617_, keyIn_0_124 );
and g416 ( new_n618_, new_n613_, new_n465_ );
xnor g417 ( new_n619_, new_n618_, new_n617_ );
xnor g418 ( N741, new_n619_, N69 );
and g419 ( new_n621_, new_n613_, new_n448_ );
xnor g420 ( new_n622_, new_n621_, keyIn_0_125 );
xnor g421 ( N742, new_n622_, N73 );
not g422 ( new_n624_, keyIn_0_126 );
and g423 ( new_n625_, new_n613_, new_n494_ );
xnor g424 ( new_n626_, new_n625_, new_n624_ );
xnor g425 ( N743, new_n626_, N77 );
not g426 ( new_n628_, keyIn_0_119 );
and g427 ( new_n629_, new_n339_, new_n316_ );
and g428 ( new_n630_, new_n629_, new_n535_ );
and g429 ( new_n631_, new_n611_, new_n630_ );
xnor g430 ( new_n632_, new_n631_, new_n628_ );
and g431 ( new_n633_, new_n632_, new_n480_ );
xnor g432 ( new_n634_, new_n633_, keyIn_0_127 );
xnor g433 ( N744, new_n634_, new_n221_ );
and g434 ( new_n636_, new_n632_, new_n465_ );
xnor g435 ( N745, new_n636_, new_n222_ );
and g436 ( new_n638_, new_n632_, new_n448_ );
xnor g437 ( N746, new_n638_, new_n231_ );
and g438 ( new_n640_, new_n632_, new_n494_ );
xnor g439 ( N747, new_n640_, new_n232_ );
and g440 ( new_n642_, new_n349_, new_n323_ );
and g441 ( new_n643_, new_n642_, new_n534_ );
and g442 ( new_n644_, new_n611_, new_n643_ );
xnor g443 ( new_n645_, new_n644_, keyIn_0_120 );
and g444 ( new_n646_, new_n645_, new_n480_ );
xor g445 ( N748, new_n646_, N97 );
and g446 ( new_n648_, new_n645_, new_n465_ );
xor g447 ( N749, new_n648_, N101 );
and g448 ( new_n650_, new_n645_, new_n448_ );
xor g449 ( N750, new_n650_, N105 );
and g450 ( new_n652_, new_n645_, new_n494_ );
xor g451 ( N751, new_n652_, N109 );
and g452 ( new_n654_, new_n642_, new_n629_ );
and g453 ( new_n655_, new_n611_, new_n654_ );
xor g454 ( new_n656_, new_n655_, keyIn_0_121 );
and g455 ( new_n657_, new_n656_, new_n480_ );
xor g456 ( N752, new_n657_, N113 );
and g457 ( new_n659_, new_n656_, new_n465_ );
xor g458 ( N753, new_n659_, N117 );
and g459 ( new_n661_, new_n656_, new_n448_ );
xor g460 ( N754, new_n661_, N121 );
and g461 ( new_n663_, new_n656_, new_n494_ );
xor g462 ( N755, new_n663_, N125 );
endmodule