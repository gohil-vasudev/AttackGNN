module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n1157_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n1058_, new_n953_, new_n257_, new_n1162_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n1145_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1159_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n1147_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n1158_, new_n572_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n923_, new_n233_, new_n469_, new_n391_, new_n1154_, new_n437_, new_n1085_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n543_, new_n924_, new_n886_, new_n371_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n1160_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n806_, new_n1016_, new_n605_, new_n1144_, new_n748_, new_n1137_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n1155_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1096_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n226_, new_n802_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n202_, keyIn_0_43 );
not g001 ( new_n203_, keyIn_0_10 );
not g002 ( new_n204_, N85 );
nand g003 ( new_n205_, new_n204_, N81 );
not g004 ( new_n206_, N81 );
nand g005 ( new_n207_, new_n206_, N85 );
nand g006 ( new_n208_, new_n205_, new_n207_ );
nand g007 ( new_n209_, new_n208_, new_n203_ );
nand g008 ( new_n210_, new_n205_, new_n207_, keyIn_0_10 );
nand g009 ( new_n211_, new_n209_, new_n210_ );
not g010 ( new_n212_, N93 );
nand g011 ( new_n213_, new_n212_, N89 );
not g012 ( new_n214_, N89 );
nand g013 ( new_n215_, new_n214_, N93 );
nand g014 ( new_n216_, new_n213_, new_n215_, keyIn_0_11 );
not g015 ( new_n217_, keyIn_0_11 );
nand g016 ( new_n218_, new_n213_, new_n215_ );
nand g017 ( new_n219_, new_n218_, new_n217_ );
nand g018 ( new_n220_, new_n211_, new_n216_, new_n219_ );
nand g019 ( new_n221_, new_n219_, new_n216_ );
nand g020 ( new_n222_, new_n221_, new_n209_, new_n210_ );
nand g021 ( new_n223_, new_n220_, new_n222_ );
nand g022 ( new_n224_, new_n223_, keyIn_0_33 );
not g023 ( new_n225_, keyIn_0_33 );
nand g024 ( new_n226_, new_n220_, new_n222_, new_n225_ );
nand g025 ( new_n227_, new_n224_, new_n226_ );
not g026 ( new_n228_, keyIn_0_32 );
not g027 ( new_n229_, N69 );
nand g028 ( new_n230_, new_n229_, N65 );
not g029 ( new_n231_, N65 );
nand g030 ( new_n232_, new_n231_, N69 );
nand g031 ( new_n233_, new_n230_, new_n232_ );
nand g032 ( new_n234_, new_n233_, keyIn_0_8 );
not g033 ( new_n235_, keyIn_0_8 );
nand g034 ( new_n236_, new_n230_, new_n232_, new_n235_ );
nand g035 ( new_n237_, new_n234_, new_n236_ );
not g036 ( new_n238_, keyIn_0_9 );
not g037 ( new_n239_, N77 );
nand g038 ( new_n240_, new_n239_, N73 );
not g039 ( new_n241_, N73 );
nand g040 ( new_n242_, new_n241_, N77 );
nand g041 ( new_n243_, new_n240_, new_n242_ );
nand g042 ( new_n244_, new_n243_, new_n238_ );
nand g043 ( new_n245_, new_n240_, new_n242_, keyIn_0_9 );
nand g044 ( new_n246_, new_n244_, new_n245_ );
nand g045 ( new_n247_, new_n237_, new_n246_ );
nand g046 ( new_n248_, new_n234_, new_n244_, new_n236_, new_n245_ );
nand g047 ( new_n249_, new_n247_, new_n248_ );
nand g048 ( new_n250_, new_n249_, new_n228_ );
nand g049 ( new_n251_, new_n247_, keyIn_0_32, new_n248_ );
nand g050 ( new_n252_, new_n250_, new_n251_ );
nand g051 ( new_n253_, new_n227_, new_n252_ );
not g052 ( new_n254_, new_n227_ );
not g053 ( new_n255_, new_n252_ );
nand g054 ( new_n256_, new_n254_, new_n255_ );
nand g055 ( new_n257_, new_n256_, new_n253_ );
nand g056 ( new_n258_, new_n257_, new_n202_ );
nand g057 ( new_n259_, new_n256_, keyIn_0_43, new_n253_ );
nand g058 ( new_n260_, N129, N137 );
nand g059 ( new_n261_, new_n258_, new_n259_, new_n260_ );
nand g060 ( new_n262_, new_n258_, new_n259_ );
nand g061 ( new_n263_, new_n262_, N129, N137 );
nand g062 ( new_n264_, new_n263_, new_n261_ );
nand g063 ( new_n265_, new_n264_, keyIn_0_47 );
not g064 ( new_n266_, keyIn_0_47 );
nand g065 ( new_n267_, new_n263_, new_n266_, new_n261_ );
nand g066 ( new_n268_, new_n265_, new_n267_ );
not g067 ( new_n269_, N49 );
nand g068 ( new_n270_, new_n269_, N33 );
not g069 ( new_n271_, N33 );
nand g070 ( new_n272_, new_n271_, N49 );
not g071 ( new_n273_, N17 );
nand g072 ( new_n274_, new_n273_, N1 );
not g073 ( new_n275_, N1 );
nand g074 ( new_n276_, new_n275_, N17 );
nand g075 ( new_n277_, new_n274_, new_n276_ );
nand g076 ( new_n278_, new_n277_, new_n270_, new_n272_ );
nand g077 ( new_n279_, new_n270_, new_n272_ );
nand g078 ( new_n280_, new_n279_, new_n274_, new_n276_ );
nand g079 ( new_n281_, new_n278_, new_n280_ );
nand g080 ( new_n282_, new_n268_, new_n281_ );
nand g081 ( new_n283_, new_n265_, new_n267_, new_n278_, new_n280_ );
nand g082 ( new_n284_, new_n282_, keyIn_0_55, new_n283_ );
not g083 ( new_n285_, keyIn_0_55 );
nand g084 ( new_n286_, new_n282_, new_n283_ );
nand g085 ( new_n287_, new_n286_, new_n285_ );
nand g086 ( new_n288_, new_n287_, new_n284_ );
not g087 ( new_n289_, keyIn_0_57 );
not g088 ( new_n290_, N101 );
nand g089 ( new_n291_, new_n290_, N97 );
not g090 ( new_n292_, N97 );
nand g091 ( new_n293_, new_n292_, N101 );
nand g092 ( new_n294_, new_n291_, new_n293_ );
nand g093 ( new_n295_, new_n294_, keyIn_0_12 );
not g094 ( new_n296_, keyIn_0_12 );
nand g095 ( new_n297_, new_n291_, new_n293_, new_n296_ );
nand g096 ( new_n298_, new_n295_, new_n297_ );
not g097 ( new_n299_, keyIn_0_13 );
not g098 ( new_n300_, N109 );
nand g099 ( new_n301_, new_n300_, N105 );
not g100 ( new_n302_, N105 );
nand g101 ( new_n303_, new_n302_, N109 );
nand g102 ( new_n304_, new_n301_, new_n303_ );
nand g103 ( new_n305_, new_n304_, new_n299_ );
nand g104 ( new_n306_, new_n301_, new_n303_, keyIn_0_13 );
nand g105 ( new_n307_, new_n305_, new_n306_ );
nand g106 ( new_n308_, new_n298_, new_n307_ );
nand g107 ( new_n309_, new_n295_, new_n305_, new_n297_, new_n306_ );
nand g108 ( new_n310_, new_n308_, new_n309_ );
nand g109 ( new_n311_, new_n310_, keyIn_0_34 );
not g110 ( new_n312_, keyIn_0_34 );
nand g111 ( new_n313_, new_n308_, new_n312_, new_n309_ );
nand g112 ( new_n314_, new_n311_, new_n313_ );
not g113 ( new_n315_, new_n314_ );
nand g114 ( new_n316_, new_n315_, new_n252_ );
nand g115 ( new_n317_, new_n255_, new_n314_ );
nand g116 ( new_n318_, new_n316_, new_n317_ );
nand g117 ( new_n319_, new_n318_, keyIn_0_45 );
not g118 ( new_n320_, keyIn_0_45 );
nand g119 ( new_n321_, new_n316_, new_n317_, new_n320_ );
nand g120 ( new_n322_, new_n319_, new_n321_ );
nand g121 ( new_n323_, new_n322_, keyIn_0_16 );
not g122 ( new_n324_, keyIn_0_16 );
nand g123 ( new_n325_, new_n319_, new_n324_, new_n321_ );
nand g124 ( new_n326_, new_n323_, N131, N137, new_n325_ );
nand g125 ( new_n327_, N131, N137 );
nand g126 ( new_n328_, new_n323_, new_n325_ );
nand g127 ( new_n329_, new_n328_, new_n327_ );
nand g128 ( new_n330_, new_n329_, new_n326_ );
nand g129 ( new_n331_, new_n330_, keyIn_0_49 );
not g130 ( new_n332_, keyIn_0_49 );
nand g131 ( new_n333_, new_n329_, new_n332_, new_n326_ );
nand g132 ( new_n334_, new_n331_, new_n333_ );
not g133 ( new_n335_, N25 );
nand g134 ( new_n336_, new_n335_, N9 );
not g135 ( new_n337_, N9 );
nand g136 ( new_n338_, new_n337_, N25 );
nand g137 ( new_n339_, new_n336_, new_n338_ );
nand g138 ( new_n340_, new_n339_, keyIn_0_21 );
not g139 ( new_n341_, keyIn_0_21 );
nand g140 ( new_n342_, new_n336_, new_n338_, new_n341_ );
nand g141 ( new_n343_, new_n340_, new_n342_ );
not g142 ( new_n344_, N57 );
nand g143 ( new_n345_, new_n344_, N41 );
not g144 ( new_n346_, N41 );
nand g145 ( new_n347_, new_n346_, N57 );
nand g146 ( new_n348_, new_n345_, new_n347_ );
nand g147 ( new_n349_, new_n348_, keyIn_0_22 );
not g148 ( new_n350_, keyIn_0_22 );
nand g149 ( new_n351_, new_n345_, new_n347_, new_n350_ );
nand g150 ( new_n352_, new_n343_, new_n349_, new_n351_ );
nand g151 ( new_n353_, new_n349_, new_n351_ );
nand g152 ( new_n354_, new_n353_, new_n340_, new_n342_ );
nand g153 ( new_n355_, new_n352_, new_n354_ );
nand g154 ( new_n356_, new_n355_, keyIn_0_36 );
not g155 ( new_n357_, keyIn_0_36 );
nand g156 ( new_n358_, new_n352_, new_n354_, new_n357_ );
nand g157 ( new_n359_, new_n356_, new_n358_ );
nand g158 ( new_n360_, new_n334_, new_n359_ );
nand g159 ( new_n361_, new_n331_, new_n333_, new_n356_, new_n358_ );
nand g160 ( new_n362_, new_n360_, new_n289_, new_n361_ );
nand g161 ( new_n363_, new_n360_, new_n361_ );
nand g162 ( new_n364_, new_n363_, keyIn_0_57 );
nand g163 ( new_n365_, new_n364_, new_n362_ );
nand g164 ( new_n366_, new_n365_, keyIn_0_63 );
not g165 ( new_n367_, keyIn_0_63 );
not g166 ( new_n368_, new_n365_ );
nand g167 ( new_n369_, new_n368_, new_n367_ );
not g168 ( new_n370_, keyIn_0_56 );
not g169 ( new_n371_, keyIn_0_35 );
not g170 ( new_n372_, keyIn_0_14 );
not g171 ( new_n373_, N117 );
nand g172 ( new_n374_, new_n373_, N113 );
not g173 ( new_n375_, N113 );
nand g174 ( new_n376_, new_n375_, N117 );
nand g175 ( new_n377_, new_n374_, new_n376_ );
nand g176 ( new_n378_, new_n377_, new_n372_ );
nand g177 ( new_n379_, new_n374_, new_n376_, keyIn_0_14 );
nand g178 ( new_n380_, new_n378_, new_n379_ );
not g179 ( new_n381_, keyIn_0_15 );
not g180 ( new_n382_, N125 );
nand g181 ( new_n383_, new_n382_, N121 );
not g182 ( new_n384_, N121 );
nand g183 ( new_n385_, new_n384_, N125 );
nand g184 ( new_n386_, new_n383_, new_n385_ );
nand g185 ( new_n387_, new_n386_, new_n381_ );
nand g186 ( new_n388_, new_n383_, new_n385_, keyIn_0_15 );
nand g187 ( new_n389_, new_n387_, new_n388_ );
nand g188 ( new_n390_, new_n380_, new_n389_ );
nand g189 ( new_n391_, new_n378_, new_n387_, new_n379_, new_n388_ );
nand g190 ( new_n392_, new_n390_, new_n391_ );
nand g191 ( new_n393_, new_n392_, new_n371_ );
nand g192 ( new_n394_, new_n390_, keyIn_0_35, new_n391_ );
nand g193 ( new_n395_, new_n393_, new_n394_ );
not g194 ( new_n396_, new_n395_ );
nand g195 ( new_n397_, new_n396_, new_n314_ );
nand g196 ( new_n398_, new_n315_, new_n395_ );
nand g197 ( new_n399_, new_n397_, new_n398_ );
nand g198 ( new_n400_, new_n399_, keyIn_0_44 );
not g199 ( new_n401_, keyIn_0_44 );
nand g200 ( new_n402_, new_n397_, new_n398_, new_n401_ );
nand g201 ( new_n403_, N130, N137 );
nand g202 ( new_n404_, new_n400_, new_n402_, new_n403_ );
nand g203 ( new_n405_, new_n400_, new_n402_ );
nand g204 ( new_n406_, new_n405_, N130, N137 );
nand g205 ( new_n407_, new_n406_, new_n404_ );
nand g206 ( new_n408_, new_n407_, keyIn_0_48 );
not g207 ( new_n409_, keyIn_0_48 );
nand g208 ( new_n410_, new_n406_, new_n409_, new_n404_ );
nand g209 ( new_n411_, new_n408_, new_n410_ );
not g210 ( new_n412_, N53 );
nand g211 ( new_n413_, new_n412_, N37 );
not g212 ( new_n414_, N37 );
nand g213 ( new_n415_, new_n414_, N53 );
not g214 ( new_n416_, N21 );
nand g215 ( new_n417_, new_n416_, N5 );
not g216 ( new_n418_, N5 );
nand g217 ( new_n419_, new_n418_, N21 );
nand g218 ( new_n420_, new_n417_, new_n419_ );
nand g219 ( new_n421_, new_n420_, new_n413_, new_n415_ );
nand g220 ( new_n422_, new_n413_, new_n415_ );
nand g221 ( new_n423_, new_n422_, new_n417_, new_n419_ );
nand g222 ( new_n424_, new_n421_, new_n423_ );
nand g223 ( new_n425_, new_n411_, new_n424_ );
nand g224 ( new_n426_, new_n408_, new_n410_, new_n421_, new_n423_ );
nand g225 ( new_n427_, new_n425_, new_n426_ );
nand g226 ( new_n428_, new_n427_, new_n370_ );
nand g227 ( new_n429_, new_n425_, keyIn_0_56, new_n426_ );
nand g228 ( new_n430_, new_n428_, new_n429_ );
nand g229 ( new_n431_, new_n288_, new_n430_ );
not g230 ( new_n432_, keyIn_0_50 );
not g231 ( new_n433_, keyIn_0_46 );
nand g232 ( new_n434_, new_n227_, new_n395_ );
nand g233 ( new_n435_, new_n254_, new_n396_ );
nand g234 ( new_n436_, new_n435_, new_n434_ );
nand g235 ( new_n437_, new_n436_, new_n433_ );
nand g236 ( new_n438_, new_n435_, keyIn_0_46, new_n434_ );
nand g237 ( new_n439_, new_n437_, N132, N137, new_n438_ );
nand g238 ( new_n440_, new_n437_, new_n438_ );
nand g239 ( new_n441_, N132, N137 );
nand g240 ( new_n442_, new_n440_, new_n441_ );
nand g241 ( new_n443_, new_n442_, new_n439_ );
nand g242 ( new_n444_, new_n443_, new_n432_ );
nand g243 ( new_n445_, new_n442_, keyIn_0_50, new_n439_ );
not g244 ( new_n446_, keyIn_0_23 );
not g245 ( new_n447_, N29 );
nand g246 ( new_n448_, new_n447_, N13 );
not g247 ( new_n449_, N13 );
nand g248 ( new_n450_, new_n449_, N29 );
nand g249 ( new_n451_, new_n448_, new_n450_ );
nand g250 ( new_n452_, new_n451_, new_n446_ );
nand g251 ( new_n453_, new_n448_, new_n450_, keyIn_0_23 );
nand g252 ( new_n454_, new_n452_, new_n453_ );
not g253 ( new_n455_, N45 );
nor g254 ( new_n456_, new_n455_, N61 );
not g255 ( new_n457_, N61 );
nor g256 ( new_n458_, new_n457_, N45 );
nor g257 ( new_n459_, new_n456_, new_n458_ );
nand g258 ( new_n460_, new_n454_, new_n459_ );
not g259 ( new_n461_, new_n459_ );
nand g260 ( new_n462_, new_n461_, new_n452_, new_n453_ );
nand g261 ( new_n463_, new_n460_, new_n462_ );
nand g262 ( new_n464_, new_n444_, new_n445_, new_n463_ );
nand g263 ( new_n465_, new_n444_, new_n445_ );
nand g264 ( new_n466_, new_n465_, new_n460_, new_n462_ );
nand g265 ( new_n467_, new_n466_, keyIn_0_58, new_n464_ );
not g266 ( new_n468_, keyIn_0_58 );
nand g267 ( new_n469_, new_n466_, new_n464_ );
nand g268 ( new_n470_, new_n469_, new_n468_ );
nand g269 ( new_n471_, new_n470_, new_n467_ );
nor g270 ( new_n472_, new_n431_, new_n471_ );
nand g271 ( new_n473_, new_n369_, new_n366_, new_n472_ );
not g272 ( new_n474_, new_n288_ );
not g273 ( new_n475_, new_n471_ );
nand g274 ( new_n476_, new_n368_, new_n430_, new_n475_ );
nand g275 ( new_n477_, new_n475_, new_n430_ );
nand g276 ( new_n478_, new_n477_, new_n365_ );
nor g277 ( new_n479_, new_n475_, new_n430_ );
not g278 ( new_n480_, new_n479_ );
nand g279 ( new_n481_, new_n476_, new_n474_, new_n478_, new_n480_ );
nand g280 ( new_n482_, new_n481_, new_n473_ );
not g281 ( new_n483_, keyIn_0_52 );
not g282 ( new_n484_, keyIn_0_40 );
not g283 ( new_n485_, keyIn_0_30 );
nand g284 ( new_n486_, new_n414_, N33 );
nand g285 ( new_n487_, new_n271_, N37 );
nand g286 ( new_n488_, new_n486_, new_n487_ );
nand g287 ( new_n489_, new_n488_, keyIn_0_4 );
not g288 ( new_n490_, keyIn_0_4 );
nand g289 ( new_n491_, new_n486_, new_n487_, new_n490_ );
nand g290 ( new_n492_, new_n489_, new_n491_ );
nand g291 ( new_n493_, new_n455_, N41 );
nand g292 ( new_n494_, new_n346_, N45 );
nand g293 ( new_n495_, new_n493_, new_n494_ );
nand g294 ( new_n496_, new_n495_, keyIn_0_5 );
not g295 ( new_n497_, keyIn_0_5 );
nand g296 ( new_n498_, new_n493_, new_n494_, new_n497_ );
nand g297 ( new_n499_, new_n496_, new_n498_ );
nand g298 ( new_n500_, new_n492_, new_n499_ );
nand g299 ( new_n501_, new_n489_, new_n496_, new_n491_, new_n498_ );
nand g300 ( new_n502_, new_n500_, new_n501_ );
nand g301 ( new_n503_, new_n502_, new_n485_ );
nand g302 ( new_n504_, new_n500_, keyIn_0_30, new_n501_ );
not g303 ( new_n505_, keyIn_0_31 );
not g304 ( new_n506_, keyIn_0_6 );
nand g305 ( new_n507_, new_n412_, N49 );
nand g306 ( new_n508_, new_n269_, N53 );
nand g307 ( new_n509_, new_n507_, new_n508_ );
nand g308 ( new_n510_, new_n509_, new_n506_ );
nand g309 ( new_n511_, new_n507_, new_n508_, keyIn_0_6 );
nand g310 ( new_n512_, new_n510_, new_n511_ );
nand g311 ( new_n513_, new_n457_, N57 );
nand g312 ( new_n514_, new_n344_, N61 );
nand g313 ( new_n515_, new_n513_, new_n514_ );
nand g314 ( new_n516_, new_n515_, keyIn_0_7 );
not g315 ( new_n517_, keyIn_0_7 );
nand g316 ( new_n518_, new_n513_, new_n514_, new_n517_ );
nand g317 ( new_n519_, new_n516_, new_n518_ );
nand g318 ( new_n520_, new_n512_, new_n519_ );
nand g319 ( new_n521_, new_n510_, new_n516_, new_n511_, new_n518_ );
nand g320 ( new_n522_, new_n520_, new_n521_ );
nand g321 ( new_n523_, new_n522_, new_n505_ );
nand g322 ( new_n524_, new_n520_, keyIn_0_31, new_n521_ );
nand g323 ( new_n525_, new_n503_, new_n523_, new_n504_, new_n524_ );
nand g324 ( new_n526_, new_n503_, new_n504_ );
nand g325 ( new_n527_, new_n523_, new_n524_ );
nand g326 ( new_n528_, new_n526_, new_n527_ );
nand g327 ( new_n529_, new_n528_, new_n484_, new_n525_ );
nand g328 ( new_n530_, new_n528_, new_n525_ );
nand g329 ( new_n531_, new_n530_, keyIn_0_40 );
nand g330 ( new_n532_, N134, N137 );
nand g331 ( new_n533_, new_n532_, keyIn_0_18 );
not g332 ( new_n534_, keyIn_0_18 );
nand g333 ( new_n535_, new_n534_, N134, N137 );
nand g334 ( new_n536_, new_n531_, new_n529_, new_n533_, new_n535_ );
nand g335 ( new_n537_, new_n531_, new_n529_ );
nand g336 ( new_n538_, new_n533_, new_n535_ );
nand g337 ( new_n539_, new_n537_, new_n538_ );
nand g338 ( new_n540_, new_n539_, new_n483_, new_n536_ );
nand g339 ( new_n541_, new_n539_, new_n536_ );
nand g340 ( new_n542_, new_n541_, keyIn_0_52 );
nand g341 ( new_n543_, new_n542_, new_n540_ );
not g342 ( new_n544_, keyIn_0_37 );
nand g343 ( new_n545_, new_n204_, N69 );
nand g344 ( new_n546_, new_n229_, N85 );
nand g345 ( new_n547_, new_n545_, new_n546_ );
nand g346 ( new_n548_, new_n547_, keyIn_0_24 );
not g347 ( new_n549_, keyIn_0_24 );
nand g348 ( new_n550_, new_n545_, new_n546_, new_n549_ );
nand g349 ( new_n551_, new_n548_, new_n550_ );
nand g350 ( new_n552_, new_n373_, N101 );
nand g351 ( new_n553_, new_n290_, N117 );
nand g352 ( new_n554_, new_n552_, new_n553_ );
nand g353 ( new_n555_, new_n554_, keyIn_0_25 );
not g354 ( new_n556_, keyIn_0_25 );
nand g355 ( new_n557_, new_n552_, new_n553_, new_n556_ );
nand g356 ( new_n558_, new_n555_, new_n557_ );
nand g357 ( new_n559_, new_n551_, new_n558_ );
nand g358 ( new_n560_, new_n548_, new_n555_, new_n550_, new_n557_ );
nand g359 ( new_n561_, new_n559_, new_n560_ );
nand g360 ( new_n562_, new_n561_, new_n544_ );
nand g361 ( new_n563_, new_n559_, keyIn_0_37, new_n560_ );
nand g362 ( new_n564_, new_n562_, new_n563_ );
not g363 ( new_n565_, new_n564_ );
nand g364 ( new_n566_, new_n543_, new_n565_ );
nand g365 ( new_n567_, new_n542_, new_n540_, new_n564_ );
nand g366 ( new_n568_, new_n566_, new_n567_ );
nand g367 ( new_n569_, new_n568_, keyIn_0_60 );
not g368 ( new_n570_, keyIn_0_60 );
nand g369 ( new_n571_, new_n566_, new_n570_, new_n567_ );
nand g370 ( new_n572_, new_n569_, new_n571_ );
not g371 ( new_n573_, new_n572_ );
not g372 ( new_n574_, keyIn_0_62 );
not g373 ( new_n575_, keyIn_0_2 );
nand g374 ( new_n576_, new_n416_, N17 );
nand g375 ( new_n577_, new_n273_, N21 );
nand g376 ( new_n578_, new_n576_, new_n577_ );
nand g377 ( new_n579_, new_n578_, new_n575_ );
nand g378 ( new_n580_, new_n576_, new_n577_, keyIn_0_2 );
nand g379 ( new_n581_, new_n579_, new_n580_ );
not g380 ( new_n582_, keyIn_0_3 );
nand g381 ( new_n583_, new_n447_, N25 );
nand g382 ( new_n584_, new_n335_, N29 );
nand g383 ( new_n585_, new_n583_, new_n584_, new_n582_ );
nand g384 ( new_n586_, new_n583_, new_n584_ );
nand g385 ( new_n587_, new_n586_, keyIn_0_3 );
nand g386 ( new_n588_, new_n581_, new_n585_, new_n587_ );
nand g387 ( new_n589_, new_n587_, new_n585_ );
nand g388 ( new_n590_, new_n589_, new_n579_, new_n580_ );
nand g389 ( new_n591_, new_n588_, new_n590_ );
nand g390 ( new_n592_, new_n591_, keyIn_0_29 );
not g391 ( new_n593_, keyIn_0_29 );
nand g392 ( new_n594_, new_n588_, new_n590_, new_n593_ );
nand g393 ( new_n595_, new_n592_, new_n594_ );
nand g394 ( new_n596_, new_n595_, new_n523_, new_n524_ );
nand g395 ( new_n597_, new_n527_, new_n592_, new_n594_ );
nand g396 ( new_n598_, new_n596_, new_n597_ );
nand g397 ( new_n599_, new_n598_, keyIn_0_42 );
not g398 ( new_n600_, keyIn_0_42 );
nand g399 ( new_n601_, new_n596_, new_n600_, new_n597_ );
nand g400 ( new_n602_, N136, N137 );
nand g401 ( new_n603_, new_n602_, keyIn_0_20 );
not g402 ( new_n604_, keyIn_0_20 );
nand g403 ( new_n605_, new_n604_, N136, N137 );
nand g404 ( new_n606_, new_n599_, new_n601_, new_n603_, new_n605_ );
nand g405 ( new_n607_, new_n599_, new_n601_ );
nand g406 ( new_n608_, new_n603_, new_n605_ );
nand g407 ( new_n609_, new_n607_, new_n608_ );
nand g408 ( new_n610_, new_n609_, keyIn_0_54, new_n606_ );
not g409 ( new_n611_, keyIn_0_54 );
nand g410 ( new_n612_, new_n609_, new_n606_ );
nand g411 ( new_n613_, new_n612_, new_n611_ );
nand g412 ( new_n614_, new_n613_, new_n610_ );
nand g413 ( new_n615_, new_n382_, N109 );
nand g414 ( new_n616_, new_n300_, N125 );
nand g415 ( new_n617_, new_n212_, N77 );
nand g416 ( new_n618_, new_n239_, N93 );
nand g417 ( new_n619_, new_n617_, new_n618_ );
nand g418 ( new_n620_, new_n619_, new_n615_, new_n616_ );
nand g419 ( new_n621_, new_n615_, new_n616_ );
nand g420 ( new_n622_, new_n621_, new_n617_, new_n618_ );
nand g421 ( new_n623_, new_n620_, new_n622_ );
nand g422 ( new_n624_, new_n614_, new_n623_ );
nand g423 ( new_n625_, new_n613_, new_n610_, new_n620_, new_n622_ );
nand g424 ( new_n626_, new_n624_, new_n574_, new_n625_ );
nand g425 ( new_n627_, new_n624_, new_n625_ );
nand g426 ( new_n628_, new_n627_, keyIn_0_62 );
nand g427 ( new_n629_, new_n628_, new_n626_ );
nor g428 ( new_n630_, new_n573_, new_n629_ );
not g429 ( new_n631_, keyIn_0_61 );
not g430 ( new_n632_, keyIn_0_53 );
nand g431 ( new_n633_, new_n418_, N1 );
nand g432 ( new_n634_, new_n275_, N5 );
nand g433 ( new_n635_, new_n633_, new_n634_ );
nand g434 ( new_n636_, new_n635_, keyIn_0_0 );
not g435 ( new_n637_, keyIn_0_0 );
nand g436 ( new_n638_, new_n633_, new_n634_, new_n637_ );
nand g437 ( new_n639_, new_n636_, new_n638_ );
not g438 ( new_n640_, keyIn_0_1 );
nand g439 ( new_n641_, new_n449_, N9 );
nand g440 ( new_n642_, new_n337_, N13 );
nand g441 ( new_n643_, new_n641_, new_n642_, new_n640_ );
nand g442 ( new_n644_, new_n641_, new_n642_ );
nand g443 ( new_n645_, new_n644_, keyIn_0_1 );
nand g444 ( new_n646_, new_n639_, new_n643_, new_n645_ );
nand g445 ( new_n647_, new_n645_, new_n643_ );
nand g446 ( new_n648_, new_n647_, new_n636_, new_n638_ );
nand g447 ( new_n649_, new_n646_, new_n648_ );
nand g448 ( new_n650_, new_n649_, keyIn_0_28 );
not g449 ( new_n651_, keyIn_0_28 );
nand g450 ( new_n652_, new_n646_, new_n648_, new_n651_ );
nand g451 ( new_n653_, new_n650_, new_n652_ );
nand g452 ( new_n654_, new_n653_, new_n503_, new_n504_ );
nand g453 ( new_n655_, new_n526_, new_n650_, new_n652_ );
nand g454 ( new_n656_, new_n654_, new_n655_ );
nand g455 ( new_n657_, new_n656_, keyIn_0_41 );
not g456 ( new_n658_, keyIn_0_41 );
nand g457 ( new_n659_, new_n654_, new_n658_, new_n655_ );
nand g458 ( new_n660_, N135, N137 );
nand g459 ( new_n661_, new_n660_, keyIn_0_19 );
not g460 ( new_n662_, keyIn_0_19 );
nand g461 ( new_n663_, new_n662_, N135, N137 );
nand g462 ( new_n664_, new_n657_, new_n659_, new_n661_, new_n663_ );
nand g463 ( new_n665_, new_n657_, new_n659_ );
nand g464 ( new_n666_, new_n661_, new_n663_ );
nand g465 ( new_n667_, new_n665_, new_n666_ );
nand g466 ( new_n668_, new_n667_, new_n632_, new_n664_ );
nand g467 ( new_n669_, new_n667_, new_n664_ );
nand g468 ( new_n670_, new_n669_, keyIn_0_53 );
nand g469 ( new_n671_, new_n670_, new_n668_ );
not g470 ( new_n672_, keyIn_0_26 );
nand g471 ( new_n673_, new_n214_, N73 );
nand g472 ( new_n674_, new_n241_, N89 );
nand g473 ( new_n675_, new_n673_, new_n674_ );
nand g474 ( new_n676_, new_n675_, new_n672_ );
nand g475 ( new_n677_, new_n673_, new_n674_, keyIn_0_26 );
nand g476 ( new_n678_, new_n676_, new_n677_ );
not g477 ( new_n679_, keyIn_0_27 );
nand g478 ( new_n680_, new_n384_, N105 );
nand g479 ( new_n681_, new_n302_, N121 );
nand g480 ( new_n682_, new_n680_, new_n681_ );
nand g481 ( new_n683_, new_n682_, new_n679_ );
nand g482 ( new_n684_, new_n680_, new_n681_, keyIn_0_27 );
nand g483 ( new_n685_, new_n683_, new_n684_ );
nand g484 ( new_n686_, new_n678_, new_n685_ );
nand g485 ( new_n687_, new_n676_, new_n683_, new_n677_, new_n684_ );
nand g486 ( new_n688_, new_n686_, new_n687_ );
nand g487 ( new_n689_, new_n688_, keyIn_0_38 );
not g488 ( new_n690_, keyIn_0_38 );
nand g489 ( new_n691_, new_n686_, new_n690_, new_n687_ );
nand g490 ( new_n692_, new_n689_, new_n691_ );
nand g491 ( new_n693_, new_n671_, new_n692_ );
nand g492 ( new_n694_, new_n670_, new_n668_, new_n689_, new_n691_ );
nand g493 ( new_n695_, new_n693_, new_n631_, new_n694_ );
nand g494 ( new_n696_, new_n693_, new_n694_ );
nand g495 ( new_n697_, new_n696_, keyIn_0_61 );
nand g496 ( new_n698_, new_n697_, new_n695_ );
not g497 ( new_n699_, new_n698_ );
not g498 ( new_n700_, keyIn_0_51 );
nand g499 ( new_n701_, new_n592_, new_n650_, new_n594_, new_n652_ );
nand g500 ( new_n702_, new_n595_, new_n653_ );
nand g501 ( new_n703_, new_n702_, keyIn_0_39, new_n701_ );
not g502 ( new_n704_, keyIn_0_39 );
nand g503 ( new_n705_, new_n702_, new_n701_ );
nand g504 ( new_n706_, new_n705_, new_n704_ );
nand g505 ( new_n707_, N133, N137 );
nand g506 ( new_n708_, new_n707_, keyIn_0_17 );
not g507 ( new_n709_, keyIn_0_17 );
nand g508 ( new_n710_, new_n709_, N133, N137 );
nand g509 ( new_n711_, new_n706_, new_n703_, new_n708_, new_n710_ );
nand g510 ( new_n712_, new_n706_, new_n703_ );
nand g511 ( new_n713_, new_n708_, new_n710_ );
nand g512 ( new_n714_, new_n712_, new_n713_ );
nand g513 ( new_n715_, new_n714_, new_n711_ );
nand g514 ( new_n716_, new_n715_, new_n700_ );
nand g515 ( new_n717_, new_n714_, keyIn_0_51, new_n711_ );
nand g516 ( new_n718_, new_n716_, new_n717_ );
nand g517 ( new_n719_, new_n375_, N97 );
nand g518 ( new_n720_, new_n292_, N113 );
nand g519 ( new_n721_, new_n206_, N65 );
nand g520 ( new_n722_, new_n231_, N81 );
nand g521 ( new_n723_, new_n721_, new_n722_ );
nand g522 ( new_n724_, new_n723_, new_n719_, new_n720_ );
nand g523 ( new_n725_, new_n719_, new_n720_ );
nand g524 ( new_n726_, new_n725_, new_n721_, new_n722_ );
nand g525 ( new_n727_, new_n724_, new_n726_ );
nand g526 ( new_n728_, new_n718_, new_n727_ );
nand g527 ( new_n729_, new_n716_, new_n717_, new_n724_, new_n726_ );
nand g528 ( new_n730_, new_n728_, keyIn_0_59, new_n729_ );
not g529 ( new_n731_, keyIn_0_59 );
nand g530 ( new_n732_, new_n728_, new_n729_ );
nand g531 ( new_n733_, new_n732_, new_n731_ );
nand g532 ( new_n734_, new_n733_, new_n730_ );
not g533 ( new_n735_, new_n734_ );
nand g534 ( new_n736_, new_n482_, new_n630_, new_n699_, new_n735_ );
not g535 ( new_n737_, new_n736_ );
nand g536 ( new_n738_, new_n737_, new_n288_ );
nand g537 ( new_n739_, new_n738_, N1 );
nand g538 ( new_n740_, new_n737_, new_n275_, new_n288_ );
nand g539 ( N724, new_n739_, new_n740_ );
not g540 ( new_n742_, new_n430_ );
nand g541 ( new_n743_, new_n737_, new_n742_ );
nand g542 ( new_n744_, new_n743_, N5 );
nand g543 ( new_n745_, new_n737_, new_n418_, new_n742_ );
nand g544 ( N725, new_n744_, new_n745_ );
nand g545 ( new_n747_, new_n737_, new_n365_ );
nand g546 ( new_n748_, new_n747_, N9 );
nand g547 ( new_n749_, new_n737_, new_n337_, new_n365_ );
nand g548 ( N726, new_n748_, new_n749_ );
nand g549 ( new_n751_, new_n737_, new_n471_ );
nand g550 ( new_n752_, new_n751_, N13 );
nand g551 ( new_n753_, new_n737_, new_n449_, new_n471_ );
nand g552 ( N727, new_n752_, new_n753_ );
not g553 ( new_n755_, keyIn_0_105 );
not g554 ( new_n756_, new_n629_ );
nor g555 ( new_n757_, new_n756_, new_n699_, new_n573_, new_n734_ );
nand g556 ( new_n758_, new_n482_, new_n757_ );
nand g557 ( new_n759_, new_n758_, keyIn_0_76 );
not g558 ( new_n760_, keyIn_0_76 );
nand g559 ( new_n761_, new_n482_, new_n760_, new_n757_ );
nand g560 ( new_n762_, new_n759_, new_n761_ );
not g561 ( new_n763_, new_n762_ );
nand g562 ( new_n764_, new_n763_, new_n288_ );
nand g563 ( new_n765_, new_n764_, keyIn_0_82 );
not g564 ( new_n766_, keyIn_0_82 );
nand g565 ( new_n767_, new_n763_, new_n766_, new_n288_ );
nand g566 ( new_n768_, new_n765_, new_n767_ );
nand g567 ( new_n769_, new_n768_, new_n273_ );
nand g568 ( new_n770_, new_n765_, N17, new_n767_ );
nand g569 ( new_n771_, new_n769_, new_n755_, new_n770_ );
nand g570 ( new_n772_, new_n769_, new_n770_ );
nand g571 ( new_n773_, new_n772_, keyIn_0_105 );
nand g572 ( new_n774_, new_n773_, new_n771_ );
not g573 ( N728, new_n774_ );
not g574 ( new_n776_, keyIn_0_83 );
nand g575 ( new_n777_, new_n763_, new_n742_ );
nand g576 ( new_n778_, new_n777_, new_n776_ );
nand g577 ( new_n779_, new_n763_, keyIn_0_83, new_n742_ );
nand g578 ( new_n780_, new_n778_, new_n779_ );
nand g579 ( new_n781_, new_n780_, N21 );
nand g580 ( new_n782_, new_n778_, new_n416_, new_n779_ );
nand g581 ( new_n783_, new_n781_, keyIn_0_106, new_n782_ );
not g582 ( new_n784_, keyIn_0_106 );
nand g583 ( new_n785_, new_n781_, new_n782_ );
nand g584 ( new_n786_, new_n785_, new_n784_ );
nand g585 ( new_n787_, new_n786_, new_n783_ );
not g586 ( N729, new_n787_ );
nand g587 ( new_n789_, new_n763_, new_n365_ );
nand g588 ( new_n790_, new_n789_, N25 );
nand g589 ( new_n791_, new_n763_, new_n335_, new_n365_ );
nand g590 ( N730, new_n790_, new_n791_ );
not g591 ( new_n793_, keyIn_0_84 );
nand g592 ( new_n794_, new_n763_, new_n471_ );
nand g593 ( new_n795_, new_n794_, new_n793_ );
nand g594 ( new_n796_, new_n763_, keyIn_0_84, new_n471_ );
nand g595 ( new_n797_, new_n795_, new_n796_ );
nand g596 ( new_n798_, new_n797_, new_n447_ );
nand g597 ( new_n799_, new_n795_, N29, new_n796_ );
nand g598 ( new_n800_, new_n798_, keyIn_0_107, new_n799_ );
not g599 ( new_n801_, keyIn_0_107 );
nand g600 ( new_n802_, new_n798_, new_n799_ );
nand g601 ( new_n803_, new_n802_, new_n801_ );
nand g602 ( new_n804_, new_n803_, new_n800_ );
not g603 ( N731, new_n804_ );
not g604 ( new_n806_, keyIn_0_108 );
not g605 ( new_n807_, keyIn_0_85 );
nor g606 ( new_n808_, new_n735_, new_n629_, new_n698_, new_n572_ );
nand g607 ( new_n809_, new_n482_, new_n808_ );
nand g608 ( new_n810_, new_n809_, keyIn_0_77 );
not g609 ( new_n811_, keyIn_0_77 );
nand g610 ( new_n812_, new_n482_, new_n811_, new_n808_ );
nand g611 ( new_n813_, new_n810_, new_n812_ );
not g612 ( new_n814_, new_n813_ );
nand g613 ( new_n815_, new_n814_, new_n288_ );
nand g614 ( new_n816_, new_n815_, new_n807_ );
nand g615 ( new_n817_, new_n814_, keyIn_0_85, new_n288_ );
nand g616 ( new_n818_, new_n816_, new_n817_ );
nand g617 ( new_n819_, new_n818_, N33 );
nand g618 ( new_n820_, new_n816_, new_n271_, new_n817_ );
nand g619 ( new_n821_, new_n819_, new_n806_, new_n820_ );
nand g620 ( new_n822_, new_n819_, new_n820_ );
nand g621 ( new_n823_, new_n822_, keyIn_0_108 );
nand g622 ( new_n824_, new_n823_, new_n821_ );
not g623 ( N732, new_n824_ );
nand g624 ( new_n826_, new_n814_, new_n742_ );
nand g625 ( new_n827_, new_n826_, keyIn_0_86 );
not g626 ( new_n828_, keyIn_0_86 );
nand g627 ( new_n829_, new_n814_, new_n828_, new_n742_ );
nand g628 ( new_n830_, new_n827_, new_n829_ );
nand g629 ( new_n831_, new_n830_, N37 );
nand g630 ( new_n832_, new_n827_, new_n414_, new_n829_ );
nand g631 ( new_n833_, new_n831_, keyIn_0_109, new_n832_ );
not g632 ( new_n834_, keyIn_0_109 );
nand g633 ( new_n835_, new_n831_, new_n832_ );
nand g634 ( new_n836_, new_n835_, new_n834_ );
nand g635 ( new_n837_, new_n836_, new_n833_ );
not g636 ( N733, new_n837_ );
not g637 ( new_n839_, keyIn_0_110 );
nand g638 ( new_n840_, new_n814_, new_n365_ );
nand g639 ( new_n841_, new_n840_, keyIn_0_87 );
not g640 ( new_n842_, keyIn_0_87 );
nand g641 ( new_n843_, new_n814_, new_n842_, new_n365_ );
nand g642 ( new_n844_, new_n841_, new_n843_ );
nand g643 ( new_n845_, new_n844_, new_n346_ );
nand g644 ( new_n846_, new_n841_, N41, new_n843_ );
nand g645 ( new_n847_, new_n845_, new_n846_ );
nand g646 ( new_n848_, new_n847_, new_n839_ );
nand g647 ( new_n849_, new_n845_, keyIn_0_110, new_n846_ );
nand g648 ( N734, new_n848_, new_n849_ );
not g649 ( new_n851_, keyIn_0_111 );
nand g650 ( new_n852_, new_n814_, new_n471_ );
nand g651 ( new_n853_, new_n852_, keyIn_0_88 );
not g652 ( new_n854_, keyIn_0_88 );
nand g653 ( new_n855_, new_n814_, new_n854_, new_n471_ );
nand g654 ( new_n856_, new_n853_, new_n855_ );
nand g655 ( new_n857_, new_n856_, new_n455_ );
nand g656 ( new_n858_, new_n853_, N45, new_n855_ );
nand g657 ( new_n859_, new_n857_, new_n851_, new_n858_ );
nand g658 ( new_n860_, new_n857_, new_n858_ );
nand g659 ( new_n861_, new_n860_, keyIn_0_111 );
nand g660 ( new_n862_, new_n861_, new_n859_ );
not g661 ( N735, new_n862_ );
nor g662 ( new_n864_, new_n735_, new_n572_ );
nand g663 ( new_n865_, new_n482_, new_n629_, new_n698_, new_n864_ );
not g664 ( new_n866_, new_n865_ );
nand g665 ( new_n867_, new_n866_, new_n288_ );
nand g666 ( new_n868_, new_n867_, N49 );
nand g667 ( new_n869_, new_n866_, new_n269_, new_n288_ );
nand g668 ( N736, new_n868_, new_n869_ );
nand g669 ( new_n871_, new_n866_, new_n742_ );
nand g670 ( new_n872_, new_n871_, N53 );
nand g671 ( new_n873_, new_n866_, new_n412_, new_n742_ );
nand g672 ( N737, new_n872_, new_n873_ );
nand g673 ( new_n875_, new_n866_, new_n365_ );
nand g674 ( new_n876_, new_n875_, N57 );
nand g675 ( new_n877_, new_n866_, new_n344_, new_n365_ );
nand g676 ( N738, new_n876_, new_n877_ );
nand g677 ( new_n879_, new_n866_, new_n471_ );
nand g678 ( new_n880_, new_n879_, N61 );
nand g679 ( new_n881_, new_n866_, new_n457_, new_n471_ );
nand g680 ( N739, new_n880_, new_n881_ );
not g681 ( new_n883_, keyIn_0_112 );
not g682 ( new_n884_, keyIn_0_78 );
nand g683 ( new_n885_, new_n629_, new_n734_, new_n572_ );
not g684 ( new_n886_, new_n885_ );
nand g685 ( new_n887_, new_n699_, keyIn_0_64 );
not g686 ( new_n888_, keyIn_0_64 );
nand g687 ( new_n889_, new_n698_, new_n888_ );
nand g688 ( new_n890_, new_n886_, new_n887_, new_n889_ );
nand g689 ( new_n891_, new_n890_, keyIn_0_71 );
not g690 ( new_n892_, keyIn_0_71 );
nand g691 ( new_n893_, new_n886_, new_n887_, new_n892_, new_n889_ );
nand g692 ( new_n894_, new_n891_, new_n893_ );
not g693 ( new_n895_, keyIn_0_65 );
nand g694 ( new_n896_, new_n697_, new_n895_, new_n695_ );
nand g695 ( new_n897_, new_n698_, keyIn_0_65 );
nand g696 ( new_n898_, new_n897_, new_n896_ );
nand g697 ( new_n899_, new_n898_, new_n864_, new_n756_ );
nand g698 ( new_n900_, new_n899_, keyIn_0_73 );
not g699 ( new_n901_, keyIn_0_73 );
nand g700 ( new_n902_, new_n898_, new_n864_, new_n901_, new_n756_ );
nand g701 ( new_n903_, new_n900_, new_n902_ );
not g702 ( new_n904_, new_n903_ );
not g703 ( new_n905_, keyIn_0_74 );
not g704 ( new_n906_, keyIn_0_66 );
nand g705 ( new_n907_, new_n697_, new_n906_, new_n695_ );
nand g706 ( new_n908_, new_n698_, keyIn_0_66 );
nand g707 ( new_n909_, new_n908_, new_n907_ );
nor g708 ( new_n910_, new_n573_, new_n629_, new_n734_ );
nand g709 ( new_n911_, new_n910_, new_n909_, new_n905_ );
nand g710 ( new_n912_, new_n910_, new_n909_ );
nand g711 ( new_n913_, new_n912_, keyIn_0_74 );
nand g712 ( new_n914_, new_n913_, new_n911_ );
nand g713 ( new_n915_, new_n756_, new_n699_, new_n572_, new_n734_ );
nand g714 ( new_n916_, new_n915_, keyIn_0_72 );
not g715 ( new_n917_, keyIn_0_72 );
nand g716 ( new_n918_, new_n630_, new_n917_, new_n699_, new_n734_ );
nand g717 ( new_n919_, new_n916_, new_n918_ );
nand g718 ( new_n920_, new_n914_, new_n919_ );
not g719 ( new_n921_, new_n920_ );
nand g720 ( new_n922_, new_n921_, keyIn_0_75, new_n894_, new_n904_ );
not g721 ( new_n923_, keyIn_0_75 );
nand g722 ( new_n924_, new_n904_, new_n894_, new_n914_, new_n919_ );
nand g723 ( new_n925_, new_n924_, new_n923_ );
nand g724 ( new_n926_, new_n925_, new_n922_ );
not g725 ( new_n927_, keyIn_0_67 );
nand g726 ( new_n928_, new_n430_, new_n927_ );
nand g727 ( new_n929_, new_n742_, keyIn_0_67 );
nand g728 ( new_n930_, new_n929_, new_n288_, new_n475_, new_n928_ );
nor g729 ( new_n931_, new_n930_, new_n368_ );
nand g730 ( new_n932_, new_n926_, new_n884_, new_n931_ );
nand g731 ( new_n933_, new_n926_, new_n931_ );
nand g732 ( new_n934_, new_n933_, keyIn_0_78 );
nand g733 ( new_n935_, new_n934_, new_n735_, new_n932_ );
nand g734 ( new_n936_, new_n935_, keyIn_0_89 );
not g735 ( new_n937_, keyIn_0_89 );
nand g736 ( new_n938_, new_n934_, new_n937_, new_n735_, new_n932_ );
nand g737 ( new_n939_, new_n936_, new_n938_ );
nand g738 ( new_n940_, new_n939_, new_n231_ );
nand g739 ( new_n941_, new_n936_, N65, new_n938_ );
nand g740 ( new_n942_, new_n940_, new_n941_ );
nand g741 ( new_n943_, new_n942_, new_n883_ );
nand g742 ( new_n944_, new_n940_, keyIn_0_112, new_n941_ );
nand g743 ( N740, new_n943_, new_n944_ );
not g744 ( new_n946_, keyIn_0_90 );
nand g745 ( new_n947_, new_n934_, new_n573_, new_n932_ );
nand g746 ( new_n948_, new_n947_, new_n946_ );
nand g747 ( new_n949_, new_n934_, keyIn_0_90, new_n573_, new_n932_ );
nand g748 ( new_n950_, new_n948_, new_n949_ );
nand g749 ( new_n951_, new_n950_, new_n229_ );
nand g750 ( new_n952_, new_n948_, N69, new_n949_ );
nand g751 ( new_n953_, new_n951_, keyIn_0_113, new_n952_ );
not g752 ( new_n954_, keyIn_0_113 );
nand g753 ( new_n955_, new_n951_, new_n952_ );
nand g754 ( new_n956_, new_n955_, new_n954_ );
nand g755 ( new_n957_, new_n956_, new_n953_ );
not g756 ( N741, new_n957_ );
not g757 ( new_n959_, keyIn_0_91 );
nand g758 ( new_n960_, new_n934_, new_n699_, new_n932_ );
nand g759 ( new_n961_, new_n960_, new_n959_ );
nand g760 ( new_n962_, new_n934_, keyIn_0_91, new_n699_, new_n932_ );
nand g761 ( new_n963_, new_n961_, new_n962_ );
nand g762 ( new_n964_, new_n963_, new_n241_ );
nand g763 ( new_n965_, new_n961_, N73, new_n962_ );
nand g764 ( new_n966_, new_n964_, new_n965_ );
nand g765 ( new_n967_, new_n966_, keyIn_0_114 );
not g766 ( new_n968_, keyIn_0_114 );
nand g767 ( new_n969_, new_n964_, new_n968_, new_n965_ );
nand g768 ( N742, new_n967_, new_n969_ );
nand g769 ( new_n971_, new_n934_, new_n629_, new_n932_ );
nand g770 ( new_n972_, new_n971_, keyIn_0_92 );
not g771 ( new_n973_, keyIn_0_92 );
nand g772 ( new_n974_, new_n934_, new_n973_, new_n629_, new_n932_ );
nand g773 ( new_n975_, new_n972_, new_n974_ );
nand g774 ( new_n976_, new_n975_, new_n239_ );
nand g775 ( new_n977_, new_n972_, N77, new_n974_ );
nand g776 ( new_n978_, new_n976_, new_n977_ );
nand g777 ( new_n979_, new_n978_, keyIn_0_115 );
not g778 ( new_n980_, keyIn_0_115 );
nand g779 ( new_n981_, new_n976_, new_n980_, new_n977_ );
nand g780 ( N743, new_n979_, new_n981_ );
not g781 ( new_n983_, keyIn_0_93 );
not g782 ( new_n984_, keyIn_0_68 );
nand g783 ( new_n985_, new_n365_, new_n984_ );
not g784 ( new_n986_, new_n985_ );
nand g785 ( new_n987_, new_n368_, keyIn_0_68 );
not g786 ( new_n988_, new_n987_ );
nor g787 ( new_n989_, new_n988_, new_n986_, new_n431_, new_n475_ );
nand g788 ( new_n990_, new_n926_, keyIn_0_79, new_n989_ );
not g789 ( new_n991_, keyIn_0_79 );
nand g790 ( new_n992_, new_n926_, new_n989_ );
nand g791 ( new_n993_, new_n992_, new_n991_ );
nand g792 ( new_n994_, new_n993_, new_n735_, new_n990_ );
nand g793 ( new_n995_, new_n994_, new_n983_ );
nand g794 ( new_n996_, new_n993_, keyIn_0_93, new_n735_, new_n990_ );
nand g795 ( new_n997_, new_n995_, new_n996_ );
nand g796 ( new_n998_, new_n997_, new_n206_ );
nand g797 ( new_n999_, new_n995_, N81, new_n996_ );
nand g798 ( new_n1000_, new_n998_, keyIn_0_116, new_n999_ );
not g799 ( new_n1001_, keyIn_0_116 );
nand g800 ( new_n1002_, new_n998_, new_n999_ );
nand g801 ( new_n1003_, new_n1002_, new_n1001_ );
nand g802 ( new_n1004_, new_n1003_, new_n1000_ );
not g803 ( N744, new_n1004_ );
nand g804 ( new_n1006_, new_n993_, new_n573_, new_n990_ );
nand g805 ( new_n1007_, new_n1006_, keyIn_0_94 );
not g806 ( new_n1008_, keyIn_0_94 );
nand g807 ( new_n1009_, new_n993_, new_n1008_, new_n573_, new_n990_ );
nand g808 ( new_n1010_, new_n1007_, new_n1009_ );
nand g809 ( new_n1011_, new_n1010_, new_n204_ );
nand g810 ( new_n1012_, new_n1007_, N85, new_n1009_ );
nand g811 ( new_n1013_, new_n1011_, keyIn_0_117, new_n1012_ );
not g812 ( new_n1014_, keyIn_0_117 );
nand g813 ( new_n1015_, new_n1011_, new_n1012_ );
nand g814 ( new_n1016_, new_n1015_, new_n1014_ );
nand g815 ( new_n1017_, new_n1016_, new_n1013_ );
not g816 ( N745, new_n1017_ );
nand g817 ( new_n1019_, new_n993_, new_n699_, new_n990_ );
nand g818 ( new_n1020_, new_n1019_, keyIn_0_95 );
not g819 ( new_n1021_, keyIn_0_95 );
nand g820 ( new_n1022_, new_n993_, new_n1021_, new_n699_, new_n990_ );
nand g821 ( new_n1023_, new_n1020_, new_n1022_ );
nand g822 ( new_n1024_, new_n1023_, N89 );
nand g823 ( new_n1025_, new_n1020_, new_n214_, new_n1022_ );
nand g824 ( new_n1026_, new_n1024_, keyIn_0_118, new_n1025_ );
not g825 ( new_n1027_, keyIn_0_118 );
nand g826 ( new_n1028_, new_n1024_, new_n1025_ );
nand g827 ( new_n1029_, new_n1028_, new_n1027_ );
nand g828 ( new_n1030_, new_n1029_, new_n1026_ );
not g829 ( N746, new_n1030_ );
nand g830 ( new_n1032_, new_n993_, new_n629_, new_n990_ );
nand g831 ( new_n1033_, new_n1032_, keyIn_0_96 );
not g832 ( new_n1034_, keyIn_0_96 );
nand g833 ( new_n1035_, new_n993_, new_n1034_, new_n629_, new_n990_ );
nand g834 ( new_n1036_, new_n1033_, new_n1035_ );
nand g835 ( new_n1037_, new_n1036_, N93 );
nand g836 ( new_n1038_, new_n1033_, new_n212_, new_n1035_ );
nand g837 ( new_n1039_, new_n1037_, new_n1038_ );
nand g838 ( new_n1040_, new_n1039_, keyIn_0_119 );
not g839 ( new_n1041_, keyIn_0_119 );
nand g840 ( new_n1042_, new_n1037_, new_n1041_, new_n1038_ );
nand g841 ( N747, new_n1040_, new_n1042_ );
not g842 ( new_n1044_, keyIn_0_97 );
not g843 ( new_n1045_, keyIn_0_80 );
nand g844 ( new_n1046_, new_n365_, new_n474_, new_n742_, new_n475_ );
not g845 ( new_n1047_, new_n1046_ );
nand g846 ( new_n1048_, new_n926_, new_n1045_, new_n1047_ );
nand g847 ( new_n1049_, new_n926_, new_n1047_ );
nand g848 ( new_n1050_, new_n1049_, keyIn_0_80 );
nand g849 ( new_n1051_, new_n1050_, new_n735_, new_n1048_ );
nand g850 ( new_n1052_, new_n1051_, new_n1044_ );
nand g851 ( new_n1053_, new_n1050_, keyIn_0_97, new_n735_, new_n1048_ );
nand g852 ( new_n1054_, new_n1052_, new_n1053_ );
nand g853 ( new_n1055_, new_n1054_, N97 );
nand g854 ( new_n1056_, new_n1052_, new_n292_, new_n1053_ );
nand g855 ( new_n1057_, new_n1055_, new_n1056_ );
nand g856 ( new_n1058_, new_n1057_, keyIn_0_120 );
not g857 ( new_n1059_, keyIn_0_120 );
nand g858 ( new_n1060_, new_n1055_, new_n1059_, new_n1056_ );
nand g859 ( N748, new_n1058_, new_n1060_ );
nand g860 ( new_n1062_, new_n1050_, new_n573_, new_n1048_ );
nand g861 ( new_n1063_, new_n1062_, keyIn_0_98 );
not g862 ( new_n1064_, keyIn_0_98 );
nand g863 ( new_n1065_, new_n1050_, new_n1064_, new_n573_, new_n1048_ );
nand g864 ( new_n1066_, new_n1063_, new_n1065_ );
nand g865 ( new_n1067_, new_n1066_, new_n290_ );
nand g866 ( new_n1068_, new_n1063_, N101, new_n1065_ );
nand g867 ( new_n1069_, new_n1067_, keyIn_0_121, new_n1068_ );
not g868 ( new_n1070_, keyIn_0_121 );
nand g869 ( new_n1071_, new_n1067_, new_n1068_ );
nand g870 ( new_n1072_, new_n1071_, new_n1070_ );
nand g871 ( new_n1073_, new_n1072_, new_n1069_ );
not g872 ( N749, new_n1073_ );
not g873 ( new_n1075_, keyIn_0_122 );
not g874 ( new_n1076_, keyIn_0_99 );
nand g875 ( new_n1077_, new_n1050_, new_n699_, new_n1048_ );
nand g876 ( new_n1078_, new_n1077_, new_n1076_ );
nand g877 ( new_n1079_, new_n1050_, keyIn_0_99, new_n699_, new_n1048_ );
nand g878 ( new_n1080_, new_n1078_, new_n1079_ );
nand g879 ( new_n1081_, new_n1080_, N105 );
nand g880 ( new_n1082_, new_n1078_, new_n302_, new_n1079_ );
nand g881 ( new_n1083_, new_n1081_, new_n1075_, new_n1082_ );
nand g882 ( new_n1084_, new_n1081_, new_n1082_ );
nand g883 ( new_n1085_, new_n1084_, keyIn_0_122 );
nand g884 ( new_n1086_, new_n1085_, new_n1083_ );
not g885 ( N750, new_n1086_ );
not g886 ( new_n1088_, keyIn_0_100 );
nand g887 ( new_n1089_, new_n1050_, new_n629_, new_n1048_ );
nand g888 ( new_n1090_, new_n1089_, new_n1088_ );
nand g889 ( new_n1091_, new_n1050_, keyIn_0_100, new_n629_, new_n1048_ );
nand g890 ( new_n1092_, new_n1090_, new_n1091_ );
nand g891 ( new_n1093_, new_n1092_, N109 );
nand g892 ( new_n1094_, new_n1090_, new_n300_, new_n1091_ );
nand g893 ( new_n1095_, new_n1093_, keyIn_0_123, new_n1094_ );
not g894 ( new_n1096_, keyIn_0_123 );
nand g895 ( new_n1097_, new_n1093_, new_n1094_ );
nand g896 ( new_n1098_, new_n1097_, new_n1096_ );
nand g897 ( new_n1099_, new_n1098_, new_n1095_ );
not g898 ( N751, new_n1099_ );
not g899 ( new_n1101_, keyIn_0_124 );
not g900 ( new_n1102_, keyIn_0_101 );
not g901 ( new_n1103_, keyIn_0_81 );
nand g902 ( new_n1104_, new_n365_, keyIn_0_70 );
not g903 ( new_n1105_, keyIn_0_70 );
nand g904 ( new_n1106_, new_n368_, new_n1105_ );
nand g905 ( new_n1107_, new_n1106_, new_n1104_ );
not g906 ( new_n1108_, keyIn_0_69 );
nand g907 ( new_n1109_, new_n474_, new_n1108_ );
nand g908 ( new_n1110_, new_n288_, keyIn_0_69 );
nand g909 ( new_n1111_, new_n1107_, new_n479_, new_n1109_, new_n1110_ );
not g910 ( new_n1112_, new_n1111_ );
nand g911 ( new_n1113_, new_n926_, new_n1103_, new_n1112_ );
nand g912 ( new_n1114_, new_n926_, new_n1112_ );
nand g913 ( new_n1115_, new_n1114_, keyIn_0_81 );
nand g914 ( new_n1116_, new_n1115_, new_n735_, new_n1113_ );
nand g915 ( new_n1117_, new_n1116_, new_n1102_ );
nand g916 ( new_n1118_, new_n1115_, keyIn_0_101, new_n735_, new_n1113_ );
nand g917 ( new_n1119_, new_n1117_, new_n1118_ );
nand g918 ( new_n1120_, new_n1119_, new_n375_ );
nand g919 ( new_n1121_, new_n1117_, N113, new_n1118_ );
nand g920 ( new_n1122_, new_n1120_, new_n1101_, new_n1121_ );
nand g921 ( new_n1123_, new_n1120_, new_n1121_ );
nand g922 ( new_n1124_, new_n1123_, keyIn_0_124 );
nand g923 ( new_n1125_, new_n1124_, new_n1122_ );
not g924 ( N752, new_n1125_ );
nand g925 ( new_n1127_, new_n1115_, new_n573_, new_n1113_ );
nand g926 ( new_n1128_, new_n1127_, keyIn_0_102 );
not g927 ( new_n1129_, keyIn_0_102 );
nand g928 ( new_n1130_, new_n1115_, new_n1129_, new_n573_, new_n1113_ );
nand g929 ( new_n1131_, new_n1128_, new_n1130_ );
nand g930 ( new_n1132_, new_n1131_, N117 );
nand g931 ( new_n1133_, new_n1128_, new_n373_, new_n1130_ );
nand g932 ( new_n1134_, new_n1132_, new_n1133_ );
nand g933 ( new_n1135_, new_n1134_, keyIn_0_125 );
not g934 ( new_n1136_, keyIn_0_125 );
nand g935 ( new_n1137_, new_n1132_, new_n1136_, new_n1133_ );
nand g936 ( N753, new_n1135_, new_n1137_ );
not g937 ( new_n1139_, keyIn_0_126 );
nand g938 ( new_n1140_, new_n1115_, new_n699_, new_n1113_ );
nand g939 ( new_n1141_, new_n1140_, keyIn_0_103 );
not g940 ( new_n1142_, keyIn_0_103 );
nand g941 ( new_n1143_, new_n1115_, new_n1142_, new_n699_, new_n1113_ );
nand g942 ( new_n1144_, new_n1141_, new_n1143_ );
nand g943 ( new_n1145_, new_n1144_, new_n384_ );
nand g944 ( new_n1146_, new_n1141_, N121, new_n1143_ );
nand g945 ( new_n1147_, new_n1145_, new_n1146_ );
nand g946 ( new_n1148_, new_n1147_, new_n1139_ );
nand g947 ( new_n1149_, new_n1145_, keyIn_0_126, new_n1146_ );
nand g948 ( N754, new_n1148_, new_n1149_ );
nand g949 ( new_n1151_, new_n1115_, new_n629_, new_n1113_ );
nand g950 ( new_n1152_, new_n1151_, keyIn_0_104 );
not g951 ( new_n1153_, keyIn_0_104 );
nand g952 ( new_n1154_, new_n1115_, new_n1153_, new_n629_, new_n1113_ );
nand g953 ( new_n1155_, new_n1152_, new_n1154_ );
nand g954 ( new_n1156_, new_n1155_, N125 );
nand g955 ( new_n1157_, new_n1152_, new_n382_, new_n1154_ );
nand g956 ( new_n1158_, new_n1156_, keyIn_0_127, new_n1157_ );
not g957 ( new_n1159_, keyIn_0_127 );
nand g958 ( new_n1160_, new_n1156_, new_n1157_ );
nand g959 ( new_n1161_, new_n1160_, new_n1159_ );
nand g960 ( new_n1162_, new_n1161_, new_n1158_ );
not g961 ( N755, new_n1162_ );
endmodule