module add_mul_comp_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, 
        b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, 
        b_13_, b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   Result_9_, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  AND2_X1 U316 ( .A1(n299), .A2(n300), .ZN(Result_9_) );
  OR2_X1 U317 ( .A1(n301), .A2(n302), .ZN(n299) );
  OR2_X1 U318 ( .A1(n303), .A2(n304), .ZN(Result_31_) );
  AND2_X1 U319 ( .A1(b_15_), .A2(n305), .ZN(n303) );
  OR2_X1 U320 ( .A1(n306), .A2(n307), .ZN(Result_30_) );
  OR2_X1 U321 ( .A1(n308), .A2(n309), .ZN(n307) );
  AND2_X1 U322 ( .A1(n310), .A2(b_14_), .ZN(n309) );
  OR2_X1 U323 ( .A1(n311), .A2(n312), .ZN(n310) );
  AND2_X1 U324 ( .A1(n313), .A2(n314), .ZN(n312) );
  AND2_X1 U325 ( .A1(a_14_), .A2(n315), .ZN(n311) );
  AND2_X1 U326 ( .A1(n316), .A2(n317), .ZN(n308) );
  AND2_X1 U327 ( .A1(a_14_), .A2(n313), .ZN(n316) );
  OR2_X1 U328 ( .A1(n318), .A2(n319), .ZN(n313) );
  AND2_X1 U329 ( .A1(n320), .A2(n321), .ZN(n319) );
  INV_X1 U330 ( .A(n304), .ZN(n321) );
  AND2_X1 U331 ( .A1(n322), .A2(n323), .ZN(n318) );
  OR2_X1 U332 ( .A1(n305), .A2(n324), .ZN(n323) );
  AND2_X1 U333 ( .A1(n325), .A2(n315), .ZN(n306) );
  OR2_X1 U334 ( .A1(n326), .A2(n327), .ZN(n315) );
  AND2_X1 U335 ( .A1(n320), .A2(n304), .ZN(n327) );
  AND2_X1 U336 ( .A1(n328), .A2(n322), .ZN(n326) );
  AND2_X1 U337 ( .A1(b_15_), .A2(a_15_), .ZN(n328) );
  OR2_X1 U338 ( .A1(n329), .A2(n330), .ZN(Result_29_) );
  AND2_X1 U339 ( .A1(n320), .A2(n331), .ZN(n330) );
  XOR2_X1 U340 ( .A(n332), .B(n333), .Z(n331) );
  AND2_X1 U341 ( .A1(n322), .A2(n334), .ZN(n329) );
  XNOR2_X1 U342 ( .A(n333), .B(n335), .ZN(n334) );
  OR2_X1 U343 ( .A1(n336), .A2(n337), .ZN(n333) );
  OR2_X1 U344 ( .A1(n338), .A2(n339), .ZN(Result_28_) );
  AND2_X1 U345 ( .A1(n320), .A2(n340), .ZN(n339) );
  XNOR2_X1 U346 ( .A(n341), .B(n342), .ZN(n340) );
  AND2_X1 U347 ( .A1(n343), .A2(n322), .ZN(n338) );
  XNOR2_X1 U348 ( .A(n342), .B(n344), .ZN(n343) );
  OR2_X1 U349 ( .A1(n345), .A2(n346), .ZN(n342) );
  OR2_X1 U350 ( .A1(n347), .A2(n348), .ZN(Result_27_) );
  AND2_X1 U351 ( .A1(n320), .A2(n349), .ZN(n348) );
  XOR2_X1 U352 ( .A(n350), .B(n351), .Z(n349) );
  AND2_X1 U353 ( .A1(n352), .A2(n322), .ZN(n347) );
  XNOR2_X1 U354 ( .A(n351), .B(n353), .ZN(n352) );
  OR2_X1 U355 ( .A1(n354), .A2(n355), .ZN(n351) );
  OR2_X1 U356 ( .A1(n356), .A2(n357), .ZN(Result_26_) );
  AND2_X1 U357 ( .A1(n320), .A2(n358), .ZN(n357) );
  XOR2_X1 U358 ( .A(n359), .B(n360), .Z(n358) );
  AND2_X1 U359 ( .A1(n361), .A2(n322), .ZN(n356) );
  XNOR2_X1 U360 ( .A(n360), .B(n362), .ZN(n361) );
  OR2_X1 U361 ( .A1(n363), .A2(n364), .ZN(n360) );
  OR2_X1 U362 ( .A1(n365), .A2(n366), .ZN(Result_25_) );
  AND2_X1 U363 ( .A1(n320), .A2(n367), .ZN(n366) );
  XOR2_X1 U364 ( .A(n368), .B(n369), .Z(n367) );
  AND2_X1 U365 ( .A1(n370), .A2(n322), .ZN(n365) );
  XNOR2_X1 U366 ( .A(n369), .B(n371), .ZN(n370) );
  OR2_X1 U367 ( .A1(n372), .A2(n373), .ZN(n369) );
  OR2_X1 U368 ( .A1(n374), .A2(n375), .ZN(Result_24_) );
  AND2_X1 U369 ( .A1(n320), .A2(n376), .ZN(n375) );
  XOR2_X1 U370 ( .A(n377), .B(n378), .Z(n376) );
  AND2_X1 U371 ( .A1(n379), .A2(n322), .ZN(n374) );
  XNOR2_X1 U372 ( .A(n378), .B(n380), .ZN(n379) );
  OR2_X1 U373 ( .A1(n381), .A2(n382), .ZN(n378) );
  OR2_X1 U374 ( .A1(n383), .A2(n384), .ZN(Result_23_) );
  AND2_X1 U375 ( .A1(n320), .A2(n385), .ZN(n384) );
  XOR2_X1 U376 ( .A(n386), .B(n387), .Z(n385) );
  AND2_X1 U377 ( .A1(n388), .A2(n322), .ZN(n383) );
  XNOR2_X1 U378 ( .A(n387), .B(n389), .ZN(n388) );
  OR2_X1 U379 ( .A1(n390), .A2(n391), .ZN(n387) );
  OR2_X1 U380 ( .A1(n392), .A2(n393), .ZN(Result_22_) );
  AND2_X1 U381 ( .A1(n320), .A2(n394), .ZN(n393) );
  XOR2_X1 U382 ( .A(n395), .B(n396), .Z(n394) );
  AND2_X1 U383 ( .A1(n397), .A2(n322), .ZN(n392) );
  XNOR2_X1 U384 ( .A(n396), .B(n398), .ZN(n397) );
  OR2_X1 U385 ( .A1(n399), .A2(n400), .ZN(n396) );
  OR2_X1 U386 ( .A1(n401), .A2(n402), .ZN(Result_21_) );
  AND2_X1 U387 ( .A1(n320), .A2(n403), .ZN(n402) );
  XOR2_X1 U388 ( .A(n404), .B(n405), .Z(n403) );
  AND2_X1 U389 ( .A1(n406), .A2(n322), .ZN(n401) );
  XNOR2_X1 U390 ( .A(n405), .B(n407), .ZN(n406) );
  OR2_X1 U391 ( .A1(n408), .A2(n409), .ZN(n405) );
  OR2_X1 U392 ( .A1(n410), .A2(n411), .ZN(Result_20_) );
  AND2_X1 U393 ( .A1(n320), .A2(n412), .ZN(n411) );
  XOR2_X1 U394 ( .A(n413), .B(n414), .Z(n412) );
  AND2_X1 U395 ( .A1(n415), .A2(n322), .ZN(n410) );
  XNOR2_X1 U396 ( .A(n414), .B(n416), .ZN(n415) );
  OR2_X1 U397 ( .A1(n417), .A2(n418), .ZN(n414) );
  OR2_X1 U398 ( .A1(n419), .A2(n420), .ZN(Result_19_) );
  AND2_X1 U399 ( .A1(n320), .A2(n421), .ZN(n420) );
  XOR2_X1 U400 ( .A(n422), .B(n423), .Z(n421) );
  AND2_X1 U401 ( .A1(n424), .A2(n322), .ZN(n419) );
  XNOR2_X1 U402 ( .A(n423), .B(n425), .ZN(n424) );
  OR2_X1 U403 ( .A1(n426), .A2(n427), .ZN(n423) );
  OR2_X1 U404 ( .A1(n428), .A2(n429), .ZN(Result_18_) );
  AND2_X1 U405 ( .A1(n320), .A2(n430), .ZN(n429) );
  XOR2_X1 U406 ( .A(n431), .B(n432), .Z(n430) );
  AND2_X1 U407 ( .A1(n433), .A2(n322), .ZN(n428) );
  XNOR2_X1 U408 ( .A(n432), .B(n434), .ZN(n433) );
  OR2_X1 U409 ( .A1(n435), .A2(n436), .ZN(n432) );
  AND2_X1 U410 ( .A1(b_2_), .A2(n437), .ZN(n435) );
  OR2_X1 U411 ( .A1(n438), .A2(n439), .ZN(Result_17_) );
  AND2_X1 U412 ( .A1(n320), .A2(n440), .ZN(n439) );
  XOR2_X1 U413 ( .A(n441), .B(n442), .Z(n440) );
  AND2_X1 U414 ( .A1(n443), .A2(n322), .ZN(n438) );
  XNOR2_X1 U415 ( .A(n441), .B(n444), .ZN(n443) );
  OR2_X1 U416 ( .A1(n445), .A2(n446), .ZN(n441) );
  INV_X1 U417 ( .A(n447), .ZN(n446) );
  OR2_X1 U418 ( .A1(n448), .A2(n449), .ZN(Result_16_) );
  AND2_X1 U419 ( .A1(n320), .A2(n450), .ZN(n449) );
  OR2_X1 U420 ( .A1(n451), .A2(n452), .ZN(n450) );
  INV_X1 U421 ( .A(n453), .ZN(n451) );
  OR2_X1 U422 ( .A1(n301), .A2(n445), .ZN(n453) );
  AND2_X1 U423 ( .A1(n447), .A2(n442), .ZN(n301) );
  OR2_X1 U424 ( .A1(n454), .A2(n436), .ZN(n442) );
  AND2_X1 U425 ( .A1(n455), .A2(n431), .ZN(n454) );
  OR2_X1 U426 ( .A1(n456), .A2(n426), .ZN(n431) );
  AND2_X1 U427 ( .A1(n422), .A2(n457), .ZN(n456) );
  OR2_X1 U428 ( .A1(n458), .A2(n417), .ZN(n422) );
  AND2_X1 U429 ( .A1(n413), .A2(n459), .ZN(n458) );
  OR2_X1 U430 ( .A1(n460), .A2(n408), .ZN(n413) );
  AND2_X1 U431 ( .A1(n404), .A2(n461), .ZN(n460) );
  OR2_X1 U432 ( .A1(n462), .A2(n399), .ZN(n404) );
  AND2_X1 U433 ( .A1(n395), .A2(n463), .ZN(n462) );
  OR2_X1 U434 ( .A1(n464), .A2(n390), .ZN(n395) );
  AND2_X1 U435 ( .A1(n386), .A2(n465), .ZN(n464) );
  OR2_X1 U436 ( .A1(n466), .A2(n381), .ZN(n386) );
  AND2_X1 U437 ( .A1(n377), .A2(n467), .ZN(n466) );
  OR2_X1 U438 ( .A1(n468), .A2(n372), .ZN(n377) );
  AND2_X1 U439 ( .A1(n368), .A2(n469), .ZN(n468) );
  OR2_X1 U440 ( .A1(n470), .A2(n363), .ZN(n368) );
  AND2_X1 U441 ( .A1(n359), .A2(n471), .ZN(n470) );
  OR2_X1 U442 ( .A1(n472), .A2(n354), .ZN(n359) );
  AND2_X1 U443 ( .A1(n350), .A2(n473), .ZN(n472) );
  OR2_X1 U444 ( .A1(n474), .A2(n345), .ZN(n350) );
  AND2_X1 U445 ( .A1(a_12_), .A2(n475), .ZN(n345) );
  AND2_X1 U446 ( .A1(n476), .A2(n477), .ZN(n474) );
  AND2_X1 U447 ( .A1(n478), .A2(n322), .ZN(n448) );
  INV_X1 U448 ( .A(n479), .ZN(n322) );
  OR2_X1 U449 ( .A1(n480), .A2(n320), .ZN(n479) );
  AND2_X1 U450 ( .A1(n300), .A2(n481), .ZN(n320) );
  OR2_X1 U451 ( .A1(n302), .A2(n482), .ZN(n481) );
  AND2_X1 U452 ( .A1(n483), .A2(n484), .ZN(n482) );
  OR2_X1 U453 ( .A1(n485), .A2(n486), .ZN(n483) );
  INV_X1 U454 ( .A(n487), .ZN(n486) );
  OR2_X1 U455 ( .A1(n488), .A2(n489), .ZN(n487) );
  OR2_X1 U456 ( .A1(n427), .A2(n418), .ZN(n489) );
  AND2_X1 U457 ( .A1(n490), .A2(n491), .ZN(n488) );
  OR2_X1 U458 ( .A1(n492), .A2(n493), .ZN(n491) );
  OR2_X1 U459 ( .A1(n409), .A2(n400), .ZN(n493) );
  AND2_X1 U460 ( .A1(n494), .A2(n495), .ZN(n492) );
  OR2_X1 U461 ( .A1(n496), .A2(n497), .ZN(n495) );
  OR2_X1 U462 ( .A1(n391), .A2(n382), .ZN(n497) );
  AND2_X1 U463 ( .A1(n498), .A2(n499), .ZN(n496) );
  OR2_X1 U464 ( .A1(n500), .A2(n501), .ZN(n499) );
  OR2_X1 U465 ( .A1(n373), .A2(n364), .ZN(n501) );
  AND2_X1 U466 ( .A1(n502), .A2(n503), .ZN(n500) );
  OR2_X1 U467 ( .A1(n504), .A2(n505), .ZN(n503) );
  OR2_X1 U468 ( .A1(n355), .A2(n346), .ZN(n505) );
  AND2_X1 U469 ( .A1(n341), .A2(n506), .ZN(n504) );
  OR2_X1 U470 ( .A1(b_12_), .A2(n507), .ZN(n506) );
  INV_X1 U471 ( .A(n476), .ZN(n341) );
  OR2_X1 U472 ( .A1(n508), .A2(n336), .ZN(n476) );
  AND2_X1 U473 ( .A1(a_13_), .A2(n509), .ZN(n336) );
  AND2_X1 U474 ( .A1(n510), .A2(n332), .ZN(n508) );
  OR2_X1 U475 ( .A1(n511), .A2(n512), .ZN(n332) );
  AND2_X1 U476 ( .A1(a_14_), .A2(n304), .ZN(n512) );
  AND2_X1 U477 ( .A1(n513), .A2(n317), .ZN(n511) );
  OR2_X1 U478 ( .A1(n304), .A2(a_14_), .ZN(n513) );
  AND2_X1 U479 ( .A1(n324), .A2(a_15_), .ZN(n304) );
  INV_X1 U480 ( .A(n514), .ZN(n502) );
  OR2_X1 U481 ( .A1(n363), .A2(n354), .ZN(n514) );
  AND2_X1 U482 ( .A1(n515), .A2(a_11_), .ZN(n354) );
  AND2_X1 U483 ( .A1(n516), .A2(a_10_), .ZN(n363) );
  INV_X1 U484 ( .A(n517), .ZN(n498) );
  OR2_X1 U485 ( .A1(n381), .A2(n372), .ZN(n517) );
  AND2_X1 U486 ( .A1(n518), .A2(a_9_), .ZN(n372) );
  AND2_X1 U487 ( .A1(n519), .A2(a_8_), .ZN(n381) );
  INV_X1 U488 ( .A(n520), .ZN(n494) );
  OR2_X1 U489 ( .A1(n399), .A2(n390), .ZN(n520) );
  AND2_X1 U490 ( .A1(n521), .A2(a_7_), .ZN(n390) );
  AND2_X1 U491 ( .A1(n522), .A2(a_6_), .ZN(n399) );
  INV_X1 U492 ( .A(n523), .ZN(n490) );
  OR2_X1 U493 ( .A1(n417), .A2(n408), .ZN(n523) );
  AND2_X1 U494 ( .A1(n524), .A2(a_5_), .ZN(n408) );
  AND2_X1 U495 ( .A1(n525), .A2(a_4_), .ZN(n417) );
  OR2_X1 U496 ( .A1(n436), .A2(n426), .ZN(n485) );
  AND2_X1 U497 ( .A1(n526), .A2(a_3_), .ZN(n426) );
  AND2_X1 U498 ( .A1(n527), .A2(a_2_), .ZN(n436) );
  OR2_X1 U499 ( .A1(n445), .A2(n528), .ZN(n302) );
  AND2_X1 U500 ( .A1(n529), .A2(a_1_), .ZN(n445) );
  AND2_X1 U501 ( .A1(n530), .A2(n531), .ZN(n480) );
  AND2_X1 U502 ( .A1(n532), .A2(n533), .ZN(n531) );
  AND2_X1 U503 ( .A1(n534), .A2(n535), .ZN(n533) );
  AND2_X1 U504 ( .A1(n457), .A2(n300), .ZN(n535) );
  INV_X1 U505 ( .A(n427), .ZN(n457) );
  AND2_X1 U506 ( .A1(n536), .A2(b_3_), .ZN(n427) );
  AND2_X1 U507 ( .A1(n461), .A2(n459), .ZN(n534) );
  INV_X1 U508 ( .A(n418), .ZN(n459) );
  AND2_X1 U509 ( .A1(n537), .A2(b_4_), .ZN(n418) );
  INV_X1 U510 ( .A(n409), .ZN(n461) );
  AND2_X1 U511 ( .A1(n538), .A2(b_5_), .ZN(n409) );
  AND2_X1 U512 ( .A1(n539), .A2(n540), .ZN(n532) );
  AND2_X1 U513 ( .A1(n465), .A2(n463), .ZN(n540) );
  INV_X1 U514 ( .A(n400), .ZN(n463) );
  AND2_X1 U515 ( .A1(n541), .A2(b_6_), .ZN(n400) );
  INV_X1 U516 ( .A(n391), .ZN(n465) );
  AND2_X1 U517 ( .A1(n542), .A2(b_7_), .ZN(n391) );
  AND2_X1 U518 ( .A1(n469), .A2(n467), .ZN(n539) );
  INV_X1 U519 ( .A(n382), .ZN(n467) );
  AND2_X1 U520 ( .A1(n543), .A2(b_8_), .ZN(n382) );
  INV_X1 U521 ( .A(n373), .ZN(n469) );
  AND2_X1 U522 ( .A1(n544), .A2(b_9_), .ZN(n373) );
  AND2_X1 U523 ( .A1(n545), .A2(n546), .ZN(n530) );
  AND2_X1 U524 ( .A1(n547), .A2(n548), .ZN(n546) );
  AND2_X1 U525 ( .A1(n473), .A2(n471), .ZN(n548) );
  INV_X1 U526 ( .A(n364), .ZN(n471) );
  AND2_X1 U527 ( .A1(n549), .A2(b_10_), .ZN(n364) );
  INV_X1 U528 ( .A(n355), .ZN(n473) );
  AND2_X1 U529 ( .A1(n550), .A2(b_11_), .ZN(n355) );
  AND2_X1 U530 ( .A1(n510), .A2(n477), .ZN(n547) );
  INV_X1 U531 ( .A(n346), .ZN(n477) );
  AND2_X1 U532 ( .A1(n507), .A2(b_12_), .ZN(n346) );
  INV_X1 U533 ( .A(n337), .ZN(n510) );
  AND2_X1 U534 ( .A1(n551), .A2(b_13_), .ZN(n337) );
  AND2_X1 U535 ( .A1(n552), .A2(n484), .ZN(n545) );
  AND2_X1 U536 ( .A1(n455), .A2(n447), .ZN(n484) );
  OR2_X1 U537 ( .A1(a_1_), .A2(n529), .ZN(n447) );
  INV_X1 U538 ( .A(b_1_), .ZN(n529) );
  OR2_X1 U539 ( .A1(n527), .A2(a_2_), .ZN(n455) );
  AND2_X1 U540 ( .A1(n553), .A2(n554), .ZN(n552) );
  OR2_X1 U541 ( .A1(a_14_), .A2(n317), .ZN(n554) );
  OR2_X1 U542 ( .A1(a_15_), .A2(n324), .ZN(n553) );
  XNOR2_X1 U543 ( .A(n452), .B(n555), .ZN(n478) );
  AND2_X1 U544 ( .A1(n556), .A2(n557), .ZN(n555) );
  OR2_X1 U545 ( .A1(b_1_), .A2(n558), .ZN(n557) );
  AND2_X1 U546 ( .A1(n559), .A2(a_1_), .ZN(n558) );
  OR2_X1 U547 ( .A1(a_1_), .A2(n559), .ZN(n556) );
  INV_X1 U548 ( .A(n444), .ZN(n559) );
  OR2_X1 U549 ( .A1(n560), .A2(n561), .ZN(n444) );
  AND2_X1 U550 ( .A1(n434), .A2(n437), .ZN(n561) );
  AND2_X1 U551 ( .A1(n562), .A2(n527), .ZN(n560) );
  INV_X1 U552 ( .A(b_2_), .ZN(n527) );
  OR2_X1 U553 ( .A1(n437), .A2(n434), .ZN(n562) );
  OR2_X1 U554 ( .A1(n563), .A2(n564), .ZN(n434) );
  AND2_X1 U555 ( .A1(n425), .A2(n536), .ZN(n564) );
  AND2_X1 U556 ( .A1(n565), .A2(n526), .ZN(n563) );
  INV_X1 U557 ( .A(b_3_), .ZN(n526) );
  OR2_X1 U558 ( .A1(n536), .A2(n425), .ZN(n565) );
  OR2_X1 U559 ( .A1(n566), .A2(n567), .ZN(n425) );
  AND2_X1 U560 ( .A1(n416), .A2(n537), .ZN(n567) );
  AND2_X1 U561 ( .A1(n568), .A2(n525), .ZN(n566) );
  INV_X1 U562 ( .A(b_4_), .ZN(n525) );
  OR2_X1 U563 ( .A1(n537), .A2(n416), .ZN(n568) );
  OR2_X1 U564 ( .A1(n569), .A2(n570), .ZN(n416) );
  AND2_X1 U565 ( .A1(n407), .A2(n538), .ZN(n570) );
  AND2_X1 U566 ( .A1(n571), .A2(n524), .ZN(n569) );
  INV_X1 U567 ( .A(b_5_), .ZN(n524) );
  OR2_X1 U568 ( .A1(n538), .A2(n407), .ZN(n571) );
  OR2_X1 U569 ( .A1(n572), .A2(n573), .ZN(n407) );
  AND2_X1 U570 ( .A1(n398), .A2(n541), .ZN(n573) );
  AND2_X1 U571 ( .A1(n574), .A2(n522), .ZN(n572) );
  INV_X1 U572 ( .A(b_6_), .ZN(n522) );
  OR2_X1 U573 ( .A1(n541), .A2(n398), .ZN(n574) );
  OR2_X1 U574 ( .A1(n575), .A2(n576), .ZN(n398) );
  AND2_X1 U575 ( .A1(n389), .A2(n542), .ZN(n576) );
  AND2_X1 U576 ( .A1(n577), .A2(n521), .ZN(n575) );
  INV_X1 U577 ( .A(b_7_), .ZN(n521) );
  OR2_X1 U578 ( .A1(n542), .A2(n389), .ZN(n577) );
  OR2_X1 U579 ( .A1(n578), .A2(n579), .ZN(n389) );
  AND2_X1 U580 ( .A1(n380), .A2(n543), .ZN(n579) );
  AND2_X1 U581 ( .A1(n580), .A2(n519), .ZN(n578) );
  INV_X1 U582 ( .A(b_8_), .ZN(n519) );
  OR2_X1 U583 ( .A1(n543), .A2(n380), .ZN(n580) );
  OR2_X1 U584 ( .A1(n581), .A2(n582), .ZN(n380) );
  AND2_X1 U585 ( .A1(n371), .A2(n544), .ZN(n582) );
  AND2_X1 U586 ( .A1(n583), .A2(n518), .ZN(n581) );
  INV_X1 U587 ( .A(b_9_), .ZN(n518) );
  OR2_X1 U588 ( .A1(n544), .A2(n371), .ZN(n583) );
  OR2_X1 U589 ( .A1(n584), .A2(n585), .ZN(n371) );
  AND2_X1 U590 ( .A1(n362), .A2(n549), .ZN(n585) );
  AND2_X1 U591 ( .A1(n586), .A2(n516), .ZN(n584) );
  INV_X1 U592 ( .A(b_10_), .ZN(n516) );
  OR2_X1 U593 ( .A1(n549), .A2(n362), .ZN(n586) );
  OR2_X1 U594 ( .A1(n587), .A2(n588), .ZN(n362) );
  AND2_X1 U595 ( .A1(n353), .A2(n550), .ZN(n588) );
  AND2_X1 U596 ( .A1(n589), .A2(n515), .ZN(n587) );
  INV_X1 U597 ( .A(b_11_), .ZN(n515) );
  OR2_X1 U598 ( .A1(n550), .A2(n353), .ZN(n589) );
  OR2_X1 U599 ( .A1(n590), .A2(n591), .ZN(n353) );
  AND2_X1 U600 ( .A1(n344), .A2(n507), .ZN(n591) );
  AND2_X1 U601 ( .A1(n592), .A2(n475), .ZN(n590) );
  INV_X1 U602 ( .A(b_12_), .ZN(n475) );
  OR2_X1 U603 ( .A1(n507), .A2(n344), .ZN(n592) );
  OR2_X1 U604 ( .A1(n593), .A2(n594), .ZN(n344) );
  AND2_X1 U605 ( .A1(n335), .A2(n551), .ZN(n594) );
  AND2_X1 U606 ( .A1(n595), .A2(n509), .ZN(n593) );
  INV_X1 U607 ( .A(b_13_), .ZN(n509) );
  OR2_X1 U608 ( .A1(n335), .A2(n551), .ZN(n595) );
  INV_X1 U609 ( .A(a_13_), .ZN(n551) );
  AND2_X1 U610 ( .A1(n596), .A2(n597), .ZN(n335) );
  OR2_X1 U611 ( .A1(n317), .A2(n314), .ZN(n597) );
  OR2_X1 U612 ( .A1(n598), .A2(n324), .ZN(n596) );
  INV_X1 U613 ( .A(b_15_), .ZN(n324) );
  OR2_X1 U614 ( .A1(n305), .A2(n325), .ZN(n598) );
  AND2_X1 U615 ( .A1(n314), .A2(n317), .ZN(n325) );
  INV_X1 U616 ( .A(b_14_), .ZN(n317) );
  INV_X1 U617 ( .A(a_14_), .ZN(n314) );
  INV_X1 U618 ( .A(a_15_), .ZN(n305) );
  INV_X1 U619 ( .A(a_12_), .ZN(n507) );
  INV_X1 U620 ( .A(a_11_), .ZN(n550) );
  INV_X1 U621 ( .A(a_10_), .ZN(n549) );
  INV_X1 U622 ( .A(a_9_), .ZN(n544) );
  INV_X1 U623 ( .A(a_8_), .ZN(n543) );
  INV_X1 U624 ( .A(a_7_), .ZN(n542) );
  INV_X1 U625 ( .A(a_6_), .ZN(n541) );
  INV_X1 U626 ( .A(a_5_), .ZN(n538) );
  INV_X1 U627 ( .A(a_4_), .ZN(n537) );
  INV_X1 U628 ( .A(a_3_), .ZN(n536) );
  INV_X1 U629 ( .A(a_2_), .ZN(n437) );
  AND2_X1 U630 ( .A1(n599), .A2(n300), .ZN(n452) );
  OR2_X1 U631 ( .A1(a_0_), .A2(n600), .ZN(n300) );
  INV_X1 U632 ( .A(n528), .ZN(n599) );
  AND2_X1 U633 ( .A1(n600), .A2(a_0_), .ZN(n528) );
  INV_X1 U634 ( .A(b_0_), .ZN(n600) );
endmodule

