module add_mul_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, operation_0_, operation_1_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_
 );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580;

  OR2_X1 U2190 ( .A1(n4493), .A2(operation_0_), .ZN(n2158) );
  INV_X2 U2191 ( .A(n2158), .ZN(n2159) );
  NAND2_X2 U2192 ( .A1(operation_0_), .A2(n4493), .ZN(n2237) );
  NOR2_X2 U2193 ( .A1(n4392), .A2(n2684), .ZN(n2685) );
  AND2_X2 U2194 ( .A1(operation_0_), .A2(operation_1_), .ZN(n2163) );
  NOR2_X2 U2195 ( .A1(operation_0_), .A2(operation_1_), .ZN(n2235) );
  NAND2_X1 U2196 ( .A1(n2160), .A2(n2161), .ZN(Result_9_) );
  NAND2_X1 U2197 ( .A1(n2162), .A2(n2163), .ZN(n2161) );
  XOR2_X1 U2198 ( .A(n2164), .B(n2165), .Z(n2162) );
  AND2_X1 U2199 ( .A1(n2166), .A2(n2167), .ZN(n2165) );
  NAND2_X1 U2200 ( .A1(n2160), .A2(n2168), .ZN(Result_8_) );
  NAND2_X1 U2201 ( .A1(n2169), .A2(n2163), .ZN(n2168) );
  XOR2_X1 U2202 ( .A(n2170), .B(n2171), .Z(n2169) );
  AND2_X1 U2203 ( .A1(n2172), .A2(n2173), .ZN(n2171) );
  NAND2_X1 U2204 ( .A1(n2160), .A2(n2174), .ZN(Result_7_) );
  NAND2_X1 U2205 ( .A1(n2175), .A2(n2163), .ZN(n2174) );
  XOR2_X1 U2206 ( .A(n2176), .B(n2177), .Z(n2175) );
  AND2_X1 U2207 ( .A1(n2178), .A2(n2179), .ZN(n2177) );
  NAND2_X1 U2208 ( .A1(n2160), .A2(n2180), .ZN(Result_6_) );
  NAND2_X1 U2209 ( .A1(n2181), .A2(n2163), .ZN(n2180) );
  XOR2_X1 U2210 ( .A(n2182), .B(n2183), .Z(n2181) );
  AND2_X1 U2211 ( .A1(n2184), .A2(n2185), .ZN(n2183) );
  NAND2_X1 U2212 ( .A1(n2160), .A2(n2186), .ZN(Result_5_) );
  NAND2_X1 U2213 ( .A1(n2187), .A2(n2163), .ZN(n2186) );
  XOR2_X1 U2214 ( .A(n2188), .B(n2189), .Z(n2187) );
  AND2_X1 U2215 ( .A1(n2190), .A2(n2191), .ZN(n2189) );
  NAND2_X1 U2216 ( .A1(n2160), .A2(n2192), .ZN(Result_4_) );
  NAND2_X1 U2217 ( .A1(n2193), .A2(n2163), .ZN(n2192) );
  XOR2_X1 U2218 ( .A(n2194), .B(n2195), .Z(n2193) );
  AND2_X1 U2219 ( .A1(n2196), .A2(n2197), .ZN(n2195) );
  NAND2_X1 U2220 ( .A1(n2160), .A2(n2198), .ZN(Result_3_) );
  NAND2_X1 U2221 ( .A1(n2199), .A2(n2163), .ZN(n2198) );
  XOR2_X1 U2222 ( .A(n2200), .B(n2201), .Z(n2199) );
  AND2_X1 U2223 ( .A1(n2202), .A2(n2203), .ZN(n2201) );
  NAND2_X1 U2224 ( .A1(n2204), .A2(n2205), .ZN(Result_31_) );
  NAND2_X1 U2225 ( .A1(n2206), .A2(n2163), .ZN(n2205) );
  NAND2_X1 U2226 ( .A1(n2207), .A2(n2208), .ZN(n2204) );
  NAND2_X1 U2227 ( .A1(n2209), .A2(n2210), .ZN(n2208) );
  NOR2_X1 U2228 ( .A1(n2211), .A2(n2159), .ZN(n2209) );
  NAND2_X1 U2229 ( .A1(n2212), .A2(n2213), .ZN(n2207) );
  NAND2_X1 U2230 ( .A1(n2214), .A2(n2215), .ZN(Result_30_) );
  NAND2_X1 U2231 ( .A1(n2163), .A2(n2216), .ZN(n2215) );
  NAND2_X1 U2232 ( .A1(n2217), .A2(n2218), .ZN(n2216) );
  NAND2_X1 U2233 ( .A1(n2219), .A2(a_14_), .ZN(n2218) );
  NOR2_X1 U2234 ( .A1(n2220), .A2(n2221), .ZN(n2217) );
  NOR2_X1 U2235 ( .A1(n2222), .A2(n2223), .ZN(n2221) );
  NOR2_X1 U2236 ( .A1(n2224), .A2(n2225), .ZN(n2220) );
  AND2_X1 U2237 ( .A1(n2226), .A2(n2212), .ZN(n2224) );
  NOR2_X1 U2238 ( .A1(n2227), .A2(n2228), .ZN(n2214) );
  NOR2_X1 U2239 ( .A1(n2229), .A2(n2230), .ZN(n2228) );
  NOR2_X1 U2240 ( .A1(n2231), .A2(n2232), .ZN(n2229) );
  NAND2_X1 U2241 ( .A1(n2233), .A2(n2234), .ZN(n2232) );
  NAND2_X1 U2242 ( .A1(n2235), .A2(n2206), .ZN(n2234) );
  INV_X1 U2243 ( .A(n2236), .ZN(n2206) );
  NAND2_X1 U2244 ( .A1(n2219), .A2(n2159), .ZN(n2233) );
  INV_X1 U2245 ( .A(n2213), .ZN(n2219) );
  NOR2_X1 U2246 ( .A1(n2237), .A2(n2212), .ZN(n2231) );
  NOR2_X1 U2247 ( .A1(n2238), .A2(n2239), .ZN(n2227) );
  NOR2_X1 U2248 ( .A1(n2240), .A2(n2241), .ZN(n2239) );
  NAND2_X1 U2249 ( .A1(n2242), .A2(n2243), .ZN(n2241) );
  NAND2_X1 U2250 ( .A1(n2235), .A2(n2236), .ZN(n2243) );
  NAND2_X1 U2251 ( .A1(n2159), .A2(n2213), .ZN(n2242) );
  AND2_X1 U2252 ( .A1(n2212), .A2(n2211), .ZN(n2240) );
  INV_X1 U2253 ( .A(n2230), .ZN(n2238) );
  NAND2_X1 U2254 ( .A1(n2223), .A2(n2244), .ZN(n2230) );
  NAND2_X1 U2255 ( .A1(n2160), .A2(n2245), .ZN(Result_2_) );
  NAND2_X1 U2256 ( .A1(n2246), .A2(n2163), .ZN(n2245) );
  XOR2_X1 U2257 ( .A(n2247), .B(n2248), .Z(n2246) );
  AND2_X1 U2258 ( .A1(n2249), .A2(n2250), .ZN(n2248) );
  NAND2_X1 U2259 ( .A1(n2251), .A2(n2252), .ZN(Result_29_) );
  NAND2_X1 U2260 ( .A1(n2253), .A2(n2163), .ZN(n2252) );
  XOR2_X1 U2261 ( .A(n2254), .B(n2255), .Z(n2253) );
  XOR2_X1 U2262 ( .A(n2256), .B(n2257), .Z(n2254) );
  NOR2_X1 U2263 ( .A1(n2258), .A2(n2259), .ZN(n2251) );
  NOR2_X1 U2264 ( .A1(n2260), .A2(n2261), .ZN(n2259) );
  NOR2_X1 U2265 ( .A1(n2262), .A2(n2263), .ZN(n2260) );
  NAND2_X1 U2266 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
  NAND2_X1 U2267 ( .A1(n2235), .A2(n2266), .ZN(n2265) );
  NAND2_X1 U2268 ( .A1(n2159), .A2(n2267), .ZN(n2264) );
  NOR2_X1 U2269 ( .A1(n2268), .A2(n2237), .ZN(n2262) );
  NOR2_X1 U2270 ( .A1(n2269), .A2(n2270), .ZN(n2258) );
  INV_X1 U2271 ( .A(n2261), .ZN(n2270) );
  XNOR2_X1 U2272 ( .A(n2271), .B(b_13_), .ZN(n2261) );
  NOR2_X1 U2273 ( .A1(n2272), .A2(n2273), .ZN(n2269) );
  NAND2_X1 U2274 ( .A1(n2274), .A2(n2275), .ZN(n2273) );
  OR2_X1 U2275 ( .A1(n2266), .A2(n2210), .ZN(n2275) );
  NAND2_X1 U2276 ( .A1(n2159), .A2(n2276), .ZN(n2274) );
  NOR2_X1 U2277 ( .A1(n2277), .A2(n2237), .ZN(n2272) );
  NAND2_X1 U2278 ( .A1(n2278), .A2(n2279), .ZN(Result_28_) );
  NAND2_X1 U2279 ( .A1(n2163), .A2(n2280), .ZN(n2279) );
  XNOR2_X1 U2280 ( .A(n2281), .B(n2282), .ZN(n2280) );
  XNOR2_X1 U2281 ( .A(n2283), .B(n2284), .ZN(n2282) );
  NOR2_X1 U2282 ( .A1(n2222), .A2(n2285), .ZN(n2284) );
  NOR2_X1 U2283 ( .A1(n2286), .A2(n2287), .ZN(n2278) );
  NOR2_X1 U2284 ( .A1(n2288), .A2(n2289), .ZN(n2287) );
  NOR2_X1 U2285 ( .A1(n2290), .A2(n2291), .ZN(n2288) );
  NAND2_X1 U2286 ( .A1(n2292), .A2(n2293), .ZN(n2291) );
  NAND2_X1 U2287 ( .A1(n2235), .A2(n2294), .ZN(n2293) );
  NAND2_X1 U2288 ( .A1(n2159), .A2(n2295), .ZN(n2292) );
  NOR2_X1 U2289 ( .A1(n2296), .A2(n2237), .ZN(n2290) );
  NOR2_X1 U2290 ( .A1(n2297), .A2(n2298), .ZN(n2286) );
  INV_X1 U2291 ( .A(n2289), .ZN(n2298) );
  XNOR2_X1 U2292 ( .A(n2299), .B(a_12_), .ZN(n2289) );
  NOR2_X1 U2293 ( .A1(n2300), .A2(n2301), .ZN(n2297) );
  NAND2_X1 U2294 ( .A1(n2302), .A2(n2303), .ZN(n2301) );
  NAND2_X1 U2295 ( .A1(n2304), .A2(n2235), .ZN(n2303) );
  NAND2_X1 U2296 ( .A1(n2159), .A2(n2305), .ZN(n2302) );
  NOR2_X1 U2297 ( .A1(n2306), .A2(n2237), .ZN(n2300) );
  NAND2_X1 U2298 ( .A1(n2307), .A2(n2308), .ZN(Result_27_) );
  NAND2_X1 U2299 ( .A1(n2309), .A2(n2163), .ZN(n2308) );
  XOR2_X1 U2300 ( .A(n2310), .B(n2311), .Z(n2309) );
  XOR2_X1 U2301 ( .A(n2312), .B(n2313), .Z(n2310) );
  NOR2_X1 U2302 ( .A1(n2222), .A2(n2314), .ZN(n2313) );
  NOR2_X1 U2303 ( .A1(n2315), .A2(n2316), .ZN(n2307) );
  NOR2_X1 U2304 ( .A1(n2317), .A2(n2318), .ZN(n2316) );
  NOR2_X1 U2305 ( .A1(n2319), .A2(n2320), .ZN(n2317) );
  NAND2_X1 U2306 ( .A1(n2321), .A2(n2322), .ZN(n2320) );
  NAND2_X1 U2307 ( .A1(n2235), .A2(n2323), .ZN(n2322) );
  NAND2_X1 U2308 ( .A1(n2159), .A2(n2324), .ZN(n2321) );
  NOR2_X1 U2309 ( .A1(n2325), .A2(n2237), .ZN(n2319) );
  NOR2_X1 U2310 ( .A1(n2326), .A2(n2327), .ZN(n2315) );
  INV_X1 U2311 ( .A(n2318), .ZN(n2327) );
  XNOR2_X1 U2312 ( .A(n2328), .B(a_11_), .ZN(n2318) );
  NOR2_X1 U2313 ( .A1(n2329), .A2(n2330), .ZN(n2326) );
  NAND2_X1 U2314 ( .A1(n2331), .A2(n2332), .ZN(n2330) );
  OR2_X1 U2315 ( .A1(n2323), .A2(n2210), .ZN(n2332) );
  NAND2_X1 U2316 ( .A1(n2159), .A2(n2333), .ZN(n2331) );
  NOR2_X1 U2317 ( .A1(n2334), .A2(n2237), .ZN(n2329) );
  NAND2_X1 U2318 ( .A1(n2335), .A2(n2336), .ZN(Result_26_) );
  NAND2_X1 U2319 ( .A1(n2163), .A2(n2337), .ZN(n2336) );
  XNOR2_X1 U2320 ( .A(n2338), .B(n2339), .ZN(n2337) );
  XOR2_X1 U2321 ( .A(n2340), .B(n2341), .Z(n2339) );
  NAND2_X1 U2322 ( .A1(a_10_), .A2(b_15_), .ZN(n2341) );
  NOR2_X1 U2323 ( .A1(n2342), .A2(n2343), .ZN(n2335) );
  NOR2_X1 U2324 ( .A1(n2344), .A2(n2345), .ZN(n2343) );
  NOR2_X1 U2325 ( .A1(n2346), .A2(n2347), .ZN(n2344) );
  NAND2_X1 U2326 ( .A1(n2348), .A2(n2349), .ZN(n2347) );
  NAND2_X1 U2327 ( .A1(n2235), .A2(n2350), .ZN(n2349) );
  NAND2_X1 U2328 ( .A1(n2159), .A2(n2351), .ZN(n2348) );
  NOR2_X1 U2329 ( .A1(n2352), .A2(n2237), .ZN(n2346) );
  NOR2_X1 U2330 ( .A1(n2353), .A2(n2354), .ZN(n2342) );
  INV_X1 U2331 ( .A(n2345), .ZN(n2354) );
  XNOR2_X1 U2332 ( .A(n2355), .B(a_10_), .ZN(n2345) );
  NOR2_X1 U2333 ( .A1(n2356), .A2(n2357), .ZN(n2353) );
  NAND2_X1 U2334 ( .A1(n2358), .A2(n2359), .ZN(n2357) );
  NAND2_X1 U2335 ( .A1(n2360), .A2(n2235), .ZN(n2359) );
  NAND2_X1 U2336 ( .A1(n2159), .A2(n2361), .ZN(n2358) );
  NOR2_X1 U2337 ( .A1(n2362), .A2(n2237), .ZN(n2356) );
  NAND2_X1 U2338 ( .A1(n2363), .A2(n2364), .ZN(Result_25_) );
  NAND2_X1 U2339 ( .A1(n2365), .A2(n2163), .ZN(n2364) );
  XNOR2_X1 U2340 ( .A(n2366), .B(n2367), .ZN(n2365) );
  NAND2_X1 U2341 ( .A1(n2368), .A2(n2369), .ZN(n2366) );
  NOR2_X1 U2342 ( .A1(n2370), .A2(n2371), .ZN(n2363) );
  NOR2_X1 U2343 ( .A1(n2372), .A2(n2373), .ZN(n2371) );
  NOR2_X1 U2344 ( .A1(n2374), .A2(n2375), .ZN(n2372) );
  NAND2_X1 U2345 ( .A1(n2376), .A2(n2377), .ZN(n2375) );
  NAND2_X1 U2346 ( .A1(n2235), .A2(n2378), .ZN(n2377) );
  NAND2_X1 U2347 ( .A1(n2159), .A2(n2379), .ZN(n2376) );
  NOR2_X1 U2348 ( .A1(n2380), .A2(n2237), .ZN(n2374) );
  NOR2_X1 U2349 ( .A1(n2381), .A2(n2382), .ZN(n2370) );
  INV_X1 U2350 ( .A(n2373), .ZN(n2382) );
  XNOR2_X1 U2351 ( .A(n2383), .B(b_9_), .ZN(n2373) );
  NOR2_X1 U2352 ( .A1(n2384), .A2(n2385), .ZN(n2381) );
  NAND2_X1 U2353 ( .A1(n2386), .A2(n2387), .ZN(n2385) );
  OR2_X1 U2354 ( .A1(n2378), .A2(n2210), .ZN(n2387) );
  NAND2_X1 U2355 ( .A1(n2159), .A2(n2388), .ZN(n2386) );
  NOR2_X1 U2356 ( .A1(n2389), .A2(n2237), .ZN(n2384) );
  NAND2_X1 U2357 ( .A1(n2390), .A2(n2391), .ZN(Result_24_) );
  NAND2_X1 U2358 ( .A1(n2163), .A2(n2392), .ZN(n2391) );
  XNOR2_X1 U2359 ( .A(n2393), .B(n2394), .ZN(n2392) );
  XOR2_X1 U2360 ( .A(n2395), .B(n2396), .Z(n2394) );
  NAND2_X1 U2361 ( .A1(a_8_), .A2(b_15_), .ZN(n2396) );
  NOR2_X1 U2362 ( .A1(n2397), .A2(n2398), .ZN(n2390) );
  NOR2_X1 U2363 ( .A1(n2399), .A2(n2400), .ZN(n2398) );
  NOR2_X1 U2364 ( .A1(n2401), .A2(n2402), .ZN(n2399) );
  NAND2_X1 U2365 ( .A1(n2403), .A2(n2404), .ZN(n2402) );
  NAND2_X1 U2366 ( .A1(n2235), .A2(n2405), .ZN(n2404) );
  NAND2_X1 U2367 ( .A1(n2159), .A2(n2406), .ZN(n2403) );
  NOR2_X1 U2368 ( .A1(n2407), .A2(n2237), .ZN(n2401) );
  NOR2_X1 U2369 ( .A1(n2408), .A2(n2409), .ZN(n2397) );
  INV_X1 U2370 ( .A(n2400), .ZN(n2409) );
  XNOR2_X1 U2371 ( .A(n2410), .B(a_8_), .ZN(n2400) );
  NOR2_X1 U2372 ( .A1(n2411), .A2(n2412), .ZN(n2408) );
  NAND2_X1 U2373 ( .A1(n2413), .A2(n2414), .ZN(n2412) );
  OR2_X1 U2374 ( .A1(n2405), .A2(n2210), .ZN(n2414) );
  NAND2_X1 U2375 ( .A1(n2159), .A2(n2415), .ZN(n2413) );
  NOR2_X1 U2376 ( .A1(n2416), .A2(n2237), .ZN(n2411) );
  NAND2_X1 U2377 ( .A1(n2417), .A2(n2418), .ZN(Result_23_) );
  NAND2_X1 U2378 ( .A1(n2419), .A2(n2163), .ZN(n2418) );
  XNOR2_X1 U2379 ( .A(n2420), .B(n2421), .ZN(n2419) );
  NAND2_X1 U2380 ( .A1(n2422), .A2(n2423), .ZN(n2420) );
  NOR2_X1 U2381 ( .A1(n2424), .A2(n2425), .ZN(n2417) );
  NOR2_X1 U2382 ( .A1(n2426), .A2(n2427), .ZN(n2425) );
  NOR2_X1 U2383 ( .A1(n2428), .A2(n2429), .ZN(n2426) );
  NAND2_X1 U2384 ( .A1(n2430), .A2(n2431), .ZN(n2429) );
  NAND2_X1 U2385 ( .A1(n2235), .A2(n2432), .ZN(n2431) );
  NAND2_X1 U2386 ( .A1(n2159), .A2(n2433), .ZN(n2430) );
  NOR2_X1 U2387 ( .A1(n2434), .A2(n2237), .ZN(n2428) );
  NOR2_X1 U2388 ( .A1(n2435), .A2(n2436), .ZN(n2424) );
  INV_X1 U2389 ( .A(n2427), .ZN(n2436) );
  XNOR2_X1 U2390 ( .A(n2437), .B(b_7_), .ZN(n2427) );
  NOR2_X1 U2391 ( .A1(n2438), .A2(n2439), .ZN(n2435) );
  NAND2_X1 U2392 ( .A1(n2440), .A2(n2441), .ZN(n2439) );
  OR2_X1 U2393 ( .A1(n2432), .A2(n2210), .ZN(n2441) );
  NAND2_X1 U2394 ( .A1(n2159), .A2(n2442), .ZN(n2440) );
  NOR2_X1 U2395 ( .A1(n2443), .A2(n2237), .ZN(n2438) );
  NAND2_X1 U2396 ( .A1(n2444), .A2(n2445), .ZN(Result_22_) );
  NAND2_X1 U2397 ( .A1(n2163), .A2(n2446), .ZN(n2445) );
  XNOR2_X1 U2398 ( .A(n2447), .B(n2448), .ZN(n2446) );
  XOR2_X1 U2399 ( .A(n2449), .B(n2450), .Z(n2448) );
  NAND2_X1 U2400 ( .A1(a_6_), .A2(b_15_), .ZN(n2450) );
  NOR2_X1 U2401 ( .A1(n2451), .A2(n2452), .ZN(n2444) );
  NOR2_X1 U2402 ( .A1(n2453), .A2(n2454), .ZN(n2452) );
  NOR2_X1 U2403 ( .A1(n2455), .A2(n2456), .ZN(n2453) );
  NAND2_X1 U2404 ( .A1(n2457), .A2(n2458), .ZN(n2456) );
  NAND2_X1 U2405 ( .A1(n2235), .A2(n2459), .ZN(n2458) );
  NAND2_X1 U2406 ( .A1(n2159), .A2(n2460), .ZN(n2457) );
  NOR2_X1 U2407 ( .A1(n2461), .A2(n2237), .ZN(n2455) );
  NOR2_X1 U2408 ( .A1(n2462), .A2(n2463), .ZN(n2451) );
  INV_X1 U2409 ( .A(n2454), .ZN(n2463) );
  XNOR2_X1 U2410 ( .A(n2464), .B(a_6_), .ZN(n2454) );
  NOR2_X1 U2411 ( .A1(n2465), .A2(n2466), .ZN(n2462) );
  NAND2_X1 U2412 ( .A1(n2467), .A2(n2468), .ZN(n2466) );
  NAND2_X1 U2413 ( .A1(n2469), .A2(n2235), .ZN(n2468) );
  NAND2_X1 U2414 ( .A1(n2159), .A2(n2470), .ZN(n2467) );
  NOR2_X1 U2415 ( .A1(n2471), .A2(n2237), .ZN(n2465) );
  NAND2_X1 U2416 ( .A1(n2472), .A2(n2473), .ZN(Result_21_) );
  NAND2_X1 U2417 ( .A1(n2474), .A2(n2163), .ZN(n2473) );
  XOR2_X1 U2418 ( .A(n2475), .B(n2476), .Z(n2474) );
  XOR2_X1 U2419 ( .A(n2477), .B(n2478), .Z(n2475) );
  NOR2_X1 U2420 ( .A1(n2222), .A2(n2479), .ZN(n2478) );
  NOR2_X1 U2421 ( .A1(n2480), .A2(n2481), .ZN(n2472) );
  NOR2_X1 U2422 ( .A1(n2482), .A2(n2483), .ZN(n2481) );
  NOR2_X1 U2423 ( .A1(n2484), .A2(n2485), .ZN(n2482) );
  NAND2_X1 U2424 ( .A1(n2486), .A2(n2487), .ZN(n2485) );
  NAND2_X1 U2425 ( .A1(n2235), .A2(n2488), .ZN(n2487) );
  NAND2_X1 U2426 ( .A1(n2159), .A2(n2489), .ZN(n2486) );
  NOR2_X1 U2427 ( .A1(n2490), .A2(n2237), .ZN(n2484) );
  NOR2_X1 U2428 ( .A1(n2491), .A2(n2492), .ZN(n2480) );
  INV_X1 U2429 ( .A(n2483), .ZN(n2492) );
  XNOR2_X1 U2430 ( .A(n2479), .B(b_5_), .ZN(n2483) );
  NOR2_X1 U2431 ( .A1(n2493), .A2(n2494), .ZN(n2491) );
  NAND2_X1 U2432 ( .A1(n2495), .A2(n2496), .ZN(n2494) );
  OR2_X1 U2433 ( .A1(n2488), .A2(n2210), .ZN(n2496) );
  NAND2_X1 U2434 ( .A1(n2159), .A2(n2497), .ZN(n2495) );
  NOR2_X1 U2435 ( .A1(n2498), .A2(n2237), .ZN(n2493) );
  NAND2_X1 U2436 ( .A1(n2499), .A2(n2500), .ZN(Result_20_) );
  NAND2_X1 U2437 ( .A1(n2501), .A2(n2163), .ZN(n2500) );
  XOR2_X1 U2438 ( .A(n2502), .B(n2503), .Z(n2501) );
  XOR2_X1 U2439 ( .A(n2504), .B(n2505), .Z(n2502) );
  NOR2_X1 U2440 ( .A1(n2222), .A2(n2506), .ZN(n2505) );
  NOR2_X1 U2441 ( .A1(n2507), .A2(n2508), .ZN(n2499) );
  NOR2_X1 U2442 ( .A1(n2509), .A2(n2510), .ZN(n2508) );
  NOR2_X1 U2443 ( .A1(n2511), .A2(n2512), .ZN(n2509) );
  NAND2_X1 U2444 ( .A1(n2513), .A2(n2514), .ZN(n2512) );
  NAND2_X1 U2445 ( .A1(n2235), .A2(n2515), .ZN(n2514) );
  NAND2_X1 U2446 ( .A1(n2159), .A2(n2516), .ZN(n2513) );
  NOR2_X1 U2447 ( .A1(n2517), .A2(n2237), .ZN(n2511) );
  NOR2_X1 U2448 ( .A1(n2518), .A2(n2519), .ZN(n2507) );
  INV_X1 U2449 ( .A(n2510), .ZN(n2519) );
  XNOR2_X1 U2450 ( .A(n2506), .B(b_4_), .ZN(n2510) );
  NOR2_X1 U2451 ( .A1(n2520), .A2(n2521), .ZN(n2518) );
  NAND2_X1 U2452 ( .A1(n2522), .A2(n2523), .ZN(n2521) );
  NAND2_X1 U2453 ( .A1(n2524), .A2(n2235), .ZN(n2523) );
  NAND2_X1 U2454 ( .A1(n2159), .A2(n2525), .ZN(n2522) );
  NOR2_X1 U2455 ( .A1(n2526), .A2(n2237), .ZN(n2520) );
  NAND2_X1 U2456 ( .A1(n2160), .A2(n2527), .ZN(Result_1_) );
  NAND2_X1 U2457 ( .A1(n2528), .A2(n2163), .ZN(n2527) );
  XNOR2_X1 U2458 ( .A(n2529), .B(n2530), .ZN(n2528) );
  NOR2_X1 U2459 ( .A1(n2531), .A2(n2532), .ZN(n2530) );
  NAND2_X1 U2460 ( .A1(n2533), .A2(n2534), .ZN(Result_19_) );
  NAND2_X1 U2461 ( .A1(n2535), .A2(n2163), .ZN(n2534) );
  XOR2_X1 U2462 ( .A(n2536), .B(n2537), .Z(n2535) );
  XOR2_X1 U2463 ( .A(n2538), .B(n2539), .Z(n2536) );
  NOR2_X1 U2464 ( .A1(n2540), .A2(n2541), .ZN(n2533) );
  NOR2_X1 U2465 ( .A1(n2542), .A2(n2543), .ZN(n2541) );
  NOR2_X1 U2466 ( .A1(n2544), .A2(n2545), .ZN(n2542) );
  NAND2_X1 U2467 ( .A1(n2546), .A2(n2547), .ZN(n2545) );
  NAND2_X1 U2468 ( .A1(n2235), .A2(n2548), .ZN(n2547) );
  NAND2_X1 U2469 ( .A1(n2159), .A2(n2549), .ZN(n2546) );
  NOR2_X1 U2470 ( .A1(n2550), .A2(n2237), .ZN(n2544) );
  NOR2_X1 U2471 ( .A1(n2551), .A2(n2552), .ZN(n2540) );
  INV_X1 U2472 ( .A(n2543), .ZN(n2552) );
  XNOR2_X1 U2473 ( .A(n2553), .B(b_3_), .ZN(n2543) );
  NOR2_X1 U2474 ( .A1(n2554), .A2(n2555), .ZN(n2551) );
  NAND2_X1 U2475 ( .A1(n2556), .A2(n2557), .ZN(n2555) );
  NAND2_X1 U2476 ( .A1(n2558), .A2(n2235), .ZN(n2557) );
  NAND2_X1 U2477 ( .A1(n2159), .A2(n2559), .ZN(n2556) );
  NOR2_X1 U2478 ( .A1(n2560), .A2(n2237), .ZN(n2554) );
  NAND2_X1 U2479 ( .A1(n2561), .A2(n2562), .ZN(Result_18_) );
  NAND2_X1 U2480 ( .A1(n2163), .A2(n2563), .ZN(n2562) );
  XNOR2_X1 U2481 ( .A(n2564), .B(n2565), .ZN(n2563) );
  XOR2_X1 U2482 ( .A(n2566), .B(n2567), .Z(n2565) );
  NAND2_X1 U2483 ( .A1(a_2_), .A2(b_15_), .ZN(n2567) );
  NOR2_X1 U2484 ( .A1(n2568), .A2(n2569), .ZN(n2561) );
  NOR2_X1 U2485 ( .A1(n2570), .A2(n2571), .ZN(n2569) );
  NOR2_X1 U2486 ( .A1(n2572), .A2(n2573), .ZN(n2570) );
  NAND2_X1 U2487 ( .A1(n2574), .A2(n2575), .ZN(n2573) );
  NAND2_X1 U2488 ( .A1(n2235), .A2(n2576), .ZN(n2575) );
  NAND2_X1 U2489 ( .A1(n2159), .A2(n2577), .ZN(n2574) );
  NOR2_X1 U2490 ( .A1(n2578), .A2(n2237), .ZN(n2572) );
  NOR2_X1 U2491 ( .A1(n2579), .A2(n2580), .ZN(n2568) );
  INV_X1 U2492 ( .A(n2571), .ZN(n2580) );
  XNOR2_X1 U2493 ( .A(n2581), .B(a_2_), .ZN(n2571) );
  NOR2_X1 U2494 ( .A1(n2582), .A2(n2583), .ZN(n2579) );
  NAND2_X1 U2495 ( .A1(n2584), .A2(n2585), .ZN(n2583) );
  NAND2_X1 U2496 ( .A1(n2586), .A2(n2235), .ZN(n2585) );
  NAND2_X1 U2497 ( .A1(n2159), .A2(n2587), .ZN(n2584) );
  NOR2_X1 U2498 ( .A1(n2588), .A2(n2237), .ZN(n2582) );
  NAND2_X1 U2499 ( .A1(n2589), .A2(n2590), .ZN(Result_17_) );
  NAND2_X1 U2500 ( .A1(n2163), .A2(n2591), .ZN(n2590) );
  XOR2_X1 U2501 ( .A(n2592), .B(n2593), .Z(n2591) );
  XOR2_X1 U2502 ( .A(n2594), .B(n2595), .Z(n2593) );
  NOR2_X1 U2503 ( .A1(n2596), .A2(n2597), .ZN(n2589) );
  NOR2_X1 U2504 ( .A1(n2598), .A2(n2599), .ZN(n2597) );
  NOR2_X1 U2505 ( .A1(n2600), .A2(n2601), .ZN(n2598) );
  NAND2_X1 U2506 ( .A1(n2602), .A2(n2603), .ZN(n2601) );
  NAND2_X1 U2507 ( .A1(n2235), .A2(n2604), .ZN(n2603) );
  NAND2_X1 U2508 ( .A1(n2159), .A2(n2605), .ZN(n2602) );
  NOR2_X1 U2509 ( .A1(n2606), .A2(n2237), .ZN(n2600) );
  NOR2_X1 U2510 ( .A1(n2607), .A2(n2608), .ZN(n2596) );
  INV_X1 U2511 ( .A(n2599), .ZN(n2608) );
  XNOR2_X1 U2512 ( .A(n2609), .B(b_1_), .ZN(n2599) );
  NOR2_X1 U2513 ( .A1(n2610), .A2(n2611), .ZN(n2607) );
  NAND2_X1 U2514 ( .A1(n2612), .A2(n2613), .ZN(n2611) );
  OR2_X1 U2515 ( .A1(n2604), .A2(n2210), .ZN(n2613) );
  NAND2_X1 U2516 ( .A1(n2159), .A2(n2614), .ZN(n2612) );
  NOR2_X1 U2517 ( .A1(n2615), .A2(n2237), .ZN(n2610) );
  NAND2_X1 U2518 ( .A1(n2616), .A2(n2617), .ZN(Result_16_) );
  NAND2_X1 U2519 ( .A1(n2618), .A2(n2163), .ZN(n2617) );
  XOR2_X1 U2520 ( .A(n2619), .B(n2620), .Z(n2618) );
  XOR2_X1 U2521 ( .A(n2621), .B(n2622), .Z(n2619) );
  NOR2_X1 U2522 ( .A1(n2222), .A2(n2623), .ZN(n2622) );
  NOR2_X1 U2523 ( .A1(n2624), .A2(n2625), .ZN(n2616) );
  NOR2_X1 U2524 ( .A1(n2626), .A2(n2627), .ZN(n2625) );
  NOR2_X1 U2525 ( .A1(n2628), .A2(n2629), .ZN(n2626) );
  NAND2_X1 U2526 ( .A1(n2630), .A2(n2631), .ZN(n2629) );
  OR2_X1 U2527 ( .A1(n2632), .A2(n2210), .ZN(n2631) );
  INV_X1 U2528 ( .A(n2235), .ZN(n2210) );
  NAND2_X1 U2529 ( .A1(n2159), .A2(n2633), .ZN(n2630) );
  NOR2_X1 U2530 ( .A1(n2634), .A2(n2237), .ZN(n2628) );
  NOR2_X1 U2531 ( .A1(n2635), .A2(n2636), .ZN(n2624) );
  INV_X1 U2532 ( .A(n2627), .ZN(n2636) );
  XNOR2_X1 U2533 ( .A(n2637), .B(a_0_), .ZN(n2627) );
  NOR2_X1 U2534 ( .A1(n2638), .A2(n2639), .ZN(n2635) );
  NAND2_X1 U2535 ( .A1(n2640), .A2(n2641), .ZN(n2639) );
  NAND2_X1 U2536 ( .A1(n2235), .A2(n2632), .ZN(n2641) );
  NAND2_X1 U2537 ( .A1(n2642), .A2(n2643), .ZN(n2632) );
  OR2_X1 U2538 ( .A1(n2604), .A2(n2644), .ZN(n2643) );
  NAND2_X1 U2539 ( .A1(n2645), .A2(n2646), .ZN(n2604) );
  NAND2_X1 U2540 ( .A1(n2647), .A2(n2576), .ZN(n2646) );
  INV_X1 U2541 ( .A(n2586), .ZN(n2576) );
  NOR2_X1 U2542 ( .A1(n2648), .A2(n2649), .ZN(n2586) );
  AND2_X1 U2543 ( .A1(n2650), .A2(n2548), .ZN(n2649) );
  INV_X1 U2544 ( .A(n2558), .ZN(n2548) );
  NOR2_X1 U2545 ( .A1(n2651), .A2(n2652), .ZN(n2558) );
  AND2_X1 U2546 ( .A1(n2653), .A2(n2515), .ZN(n2652) );
  INV_X1 U2547 ( .A(n2524), .ZN(n2515) );
  NOR2_X1 U2548 ( .A1(n2654), .A2(n2655), .ZN(n2524) );
  AND2_X1 U2549 ( .A1(n2656), .A2(n2488), .ZN(n2655) );
  NAND2_X1 U2550 ( .A1(n2657), .A2(n2658), .ZN(n2488) );
  NAND2_X1 U2551 ( .A1(n2659), .A2(n2459), .ZN(n2658) );
  INV_X1 U2552 ( .A(n2469), .ZN(n2459) );
  NOR2_X1 U2553 ( .A1(n2660), .A2(n2661), .ZN(n2469) );
  AND2_X1 U2554 ( .A1(n2662), .A2(n2432), .ZN(n2661) );
  NAND2_X1 U2555 ( .A1(n2663), .A2(n2664), .ZN(n2432) );
  NAND2_X1 U2556 ( .A1(n2665), .A2(n2405), .ZN(n2664) );
  NAND2_X1 U2557 ( .A1(n2666), .A2(n2667), .ZN(n2405) );
  NAND2_X1 U2558 ( .A1(n2668), .A2(n2378), .ZN(n2667) );
  NAND2_X1 U2559 ( .A1(n2669), .A2(n2670), .ZN(n2378) );
  NAND2_X1 U2560 ( .A1(n2671), .A2(n2350), .ZN(n2670) );
  INV_X1 U2561 ( .A(n2360), .ZN(n2350) );
  NOR2_X1 U2562 ( .A1(n2672), .A2(n2673), .ZN(n2360) );
  AND2_X1 U2563 ( .A1(n2674), .A2(n2323), .ZN(n2673) );
  NAND2_X1 U2564 ( .A1(n2675), .A2(n2676), .ZN(n2323) );
  NAND2_X1 U2565 ( .A1(n2677), .A2(n2294), .ZN(n2676) );
  INV_X1 U2566 ( .A(n2304), .ZN(n2294) );
  NOR2_X1 U2567 ( .A1(n2678), .A2(n2679), .ZN(n2304) );
  AND2_X1 U2568 ( .A1(n2680), .A2(n2266), .ZN(n2679) );
  NAND2_X1 U2569 ( .A1(n2681), .A2(n2682), .ZN(n2266) );
  NAND2_X1 U2570 ( .A1(b_14_), .A2(n2683), .ZN(n2682) );
  NAND2_X1 U2571 ( .A1(n2684), .A2(n2236), .ZN(n2683) );
  NAND2_X1 U2572 ( .A1(a_15_), .A2(b_15_), .ZN(n2236) );
  NAND2_X1 U2573 ( .A1(n2685), .A2(b_15_), .ZN(n2681) );
  NAND2_X1 U2574 ( .A1(n2686), .A2(n2271), .ZN(n2680) );
  NAND2_X1 U2575 ( .A1(n2299), .A2(n2285), .ZN(n2677) );
  NAND2_X1 U2576 ( .A1(n2328), .A2(n2314), .ZN(n2674) );
  NAND2_X1 U2577 ( .A1(n2355), .A2(n2687), .ZN(n2671) );
  NAND2_X1 U2578 ( .A1(n2688), .A2(n2383), .ZN(n2668) );
  NAND2_X1 U2579 ( .A1(n2410), .A2(n2689), .ZN(n2665) );
  NAND2_X1 U2580 ( .A1(n2690), .A2(n2437), .ZN(n2662) );
  NAND2_X1 U2581 ( .A1(n2464), .A2(n2691), .ZN(n2659) );
  NAND2_X1 U2582 ( .A1(n2692), .A2(n2479), .ZN(n2656) );
  NAND2_X1 U2583 ( .A1(n2693), .A2(n2506), .ZN(n2653) );
  NAND2_X1 U2584 ( .A1(n2694), .A2(n2553), .ZN(n2650) );
  NAND2_X1 U2585 ( .A1(n2581), .A2(n2695), .ZN(n2647) );
  NAND2_X1 U2586 ( .A1(n2696), .A2(n2609), .ZN(n2642) );
  NAND2_X1 U2587 ( .A1(n2159), .A2(n2697), .ZN(n2640) );
  NOR2_X1 U2588 ( .A1(n2698), .A2(n2237), .ZN(n2638) );
  NAND2_X1 U2589 ( .A1(n2160), .A2(n2699), .ZN(Result_15_) );
  NAND2_X1 U2590 ( .A1(n2163), .A2(n2700), .ZN(n2699) );
  XOR2_X1 U2591 ( .A(n2701), .B(n2702), .Z(n2700) );
  NAND2_X1 U2592 ( .A1(n2160), .A2(n2703), .ZN(Result_14_) );
  NAND2_X1 U2593 ( .A1(n2704), .A2(n2163), .ZN(n2703) );
  NOR2_X1 U2594 ( .A1(n2705), .A2(n2706), .ZN(n2704) );
  NOR2_X1 U2595 ( .A1(n2707), .A2(n2708), .ZN(n2706) );
  AND2_X1 U2596 ( .A1(n2701), .A2(n2702), .ZN(n2707) );
  NAND2_X1 U2597 ( .A1(n2160), .A2(n2709), .ZN(Result_13_) );
  NAND2_X1 U2598 ( .A1(n2163), .A2(n2710), .ZN(n2709) );
  XNOR2_X1 U2599 ( .A(n2705), .B(n2711), .ZN(n2710) );
  NAND2_X1 U2600 ( .A1(n2712), .A2(n2713), .ZN(n2711) );
  NAND2_X1 U2601 ( .A1(n2714), .A2(n2715), .ZN(n2713) );
  INV_X1 U2602 ( .A(n2716), .ZN(n2715) );
  NAND2_X1 U2603 ( .A1(n2717), .A2(n2718), .ZN(n2714) );
  NAND2_X1 U2604 ( .A1(n2160), .A2(n2719), .ZN(Result_12_) );
  NAND2_X1 U2605 ( .A1(n2720), .A2(n2163), .ZN(n2719) );
  XOR2_X1 U2606 ( .A(n2721), .B(n2722), .Z(n2720) );
  NAND2_X1 U2607 ( .A1(n2160), .A2(n2723), .ZN(Result_11_) );
  NAND2_X1 U2608 ( .A1(n2163), .A2(n2724), .ZN(n2723) );
  XNOR2_X1 U2609 ( .A(n2725), .B(n2726), .ZN(n2724) );
  NAND2_X1 U2610 ( .A1(n2727), .A2(n2728), .ZN(n2726) );
  NAND2_X1 U2611 ( .A1(n2160), .A2(n2729), .ZN(Result_10_) );
  NAND2_X1 U2612 ( .A1(n2730), .A2(n2163), .ZN(n2729) );
  XNOR2_X1 U2613 ( .A(n2731), .B(n2732), .ZN(n2730) );
  NAND2_X1 U2614 ( .A1(n2733), .A2(n2734), .ZN(n2731) );
  NAND2_X1 U2615 ( .A1(n2160), .A2(n2735), .ZN(Result_0_) );
  NAND2_X1 U2616 ( .A1(n2163), .A2(n2736), .ZN(n2735) );
  NAND2_X1 U2617 ( .A1(n2737), .A2(n2738), .ZN(n2736) );
  NAND2_X1 U2618 ( .A1(a_0_), .A2(n2739), .ZN(n2738) );
  NOR2_X1 U2619 ( .A1(n2532), .A2(n2740), .ZN(n2737) );
  NOR2_X1 U2620 ( .A1(n2529), .A2(n2531), .ZN(n2740) );
  AND2_X1 U2621 ( .A1(n2741), .A2(n2742), .ZN(n2531) );
  XOR2_X1 U2622 ( .A(n2739), .B(n2743), .Z(n2741) );
  NAND2_X1 U2623 ( .A1(b_0_), .A2(a_0_), .ZN(n2743) );
  AND2_X1 U2624 ( .A1(n2250), .A2(n2744), .ZN(n2529) );
  NAND2_X1 U2625 ( .A1(n2249), .A2(n2247), .ZN(n2744) );
  NAND2_X1 U2626 ( .A1(n2203), .A2(n2745), .ZN(n2247) );
  NAND2_X1 U2627 ( .A1(n2202), .A2(n2200), .ZN(n2745) );
  NAND2_X1 U2628 ( .A1(n2197), .A2(n2746), .ZN(n2200) );
  NAND2_X1 U2629 ( .A1(n2196), .A2(n2194), .ZN(n2746) );
  NAND2_X1 U2630 ( .A1(n2191), .A2(n2747), .ZN(n2194) );
  NAND2_X1 U2631 ( .A1(n2190), .A2(n2188), .ZN(n2747) );
  NAND2_X1 U2632 ( .A1(n2185), .A2(n2748), .ZN(n2188) );
  NAND2_X1 U2633 ( .A1(n2184), .A2(n2182), .ZN(n2748) );
  NAND2_X1 U2634 ( .A1(n2179), .A2(n2749), .ZN(n2182) );
  NAND2_X1 U2635 ( .A1(n2178), .A2(n2176), .ZN(n2749) );
  NAND2_X1 U2636 ( .A1(n2173), .A2(n2750), .ZN(n2176) );
  NAND2_X1 U2637 ( .A1(n2172), .A2(n2170), .ZN(n2750) );
  NAND2_X1 U2638 ( .A1(n2167), .A2(n2751), .ZN(n2170) );
  NAND2_X1 U2639 ( .A1(n2166), .A2(n2164), .ZN(n2751) );
  NAND2_X1 U2640 ( .A1(n2733), .A2(n2752), .ZN(n2164) );
  NAND2_X1 U2641 ( .A1(n2732), .A2(n2734), .ZN(n2752) );
  NAND2_X1 U2642 ( .A1(n2753), .A2(n2754), .ZN(n2734) );
  XOR2_X1 U2643 ( .A(n2755), .B(n2756), .Z(n2753) );
  NAND2_X1 U2644 ( .A1(n2727), .A2(n2757), .ZN(n2732) );
  NAND2_X1 U2645 ( .A1(n2725), .A2(n2728), .ZN(n2757) );
  NAND2_X1 U2646 ( .A1(n2758), .A2(n2759), .ZN(n2728) );
  NAND2_X1 U2647 ( .A1(n2760), .A2(n2754), .ZN(n2759) );
  NAND2_X1 U2648 ( .A1(n2761), .A2(n2762), .ZN(n2760) );
  NAND2_X1 U2649 ( .A1(n2763), .A2(n2764), .ZN(n2758) );
  NOR2_X1 U2650 ( .A1(n2721), .A2(n2722), .ZN(n2725) );
  AND2_X1 U2651 ( .A1(n2765), .A2(n2766), .ZN(n2722) );
  NAND2_X1 U2652 ( .A1(n2705), .A2(n2716), .ZN(n2766) );
  AND2_X1 U2653 ( .A1(n2767), .A2(n2702), .ZN(n2705) );
  XOR2_X1 U2654 ( .A(n2768), .B(n2769), .Z(n2702) );
  XOR2_X1 U2655 ( .A(n2770), .B(n2771), .Z(n2768) );
  NOR2_X1 U2656 ( .A1(n2225), .A2(n2623), .ZN(n2771) );
  AND2_X1 U2657 ( .A1(n2701), .A2(n2708), .ZN(n2767) );
  XOR2_X1 U2658 ( .A(n2718), .B(n2717), .Z(n2708) );
  NAND2_X1 U2659 ( .A1(n2772), .A2(n2773), .ZN(n2701) );
  NAND2_X1 U2660 ( .A1(n2774), .A2(a_0_), .ZN(n2773) );
  NOR2_X1 U2661 ( .A1(n2775), .A2(n2222), .ZN(n2774) );
  NOR2_X1 U2662 ( .A1(n2620), .A2(n2621), .ZN(n2775) );
  NAND2_X1 U2663 ( .A1(n2620), .A2(n2621), .ZN(n2772) );
  NAND2_X1 U2664 ( .A1(n2776), .A2(n2777), .ZN(n2621) );
  NAND2_X1 U2665 ( .A1(n2595), .A2(n2778), .ZN(n2777) );
  NAND2_X1 U2666 ( .A1(n2594), .A2(n2592), .ZN(n2778) );
  NOR2_X1 U2667 ( .A1(n2609), .A2(n2222), .ZN(n2595) );
  OR2_X1 U2668 ( .A1(n2592), .A2(n2594), .ZN(n2776) );
  AND2_X1 U2669 ( .A1(n2779), .A2(n2780), .ZN(n2594) );
  NAND2_X1 U2670 ( .A1(n2781), .A2(a_2_), .ZN(n2780) );
  NOR2_X1 U2671 ( .A1(n2782), .A2(n2222), .ZN(n2781) );
  NOR2_X1 U2672 ( .A1(n2564), .A2(n2566), .ZN(n2782) );
  NAND2_X1 U2673 ( .A1(n2564), .A2(n2566), .ZN(n2779) );
  NAND2_X1 U2674 ( .A1(n2783), .A2(n2784), .ZN(n2566) );
  NAND2_X1 U2675 ( .A1(n2537), .A2(n2785), .ZN(n2784) );
  OR2_X1 U2676 ( .A1(n2538), .A2(n2539), .ZN(n2785) );
  XNOR2_X1 U2677 ( .A(n2786), .B(n2787), .ZN(n2537) );
  XOR2_X1 U2678 ( .A(n2788), .B(n2789), .Z(n2787) );
  NAND2_X1 U2679 ( .A1(a_4_), .A2(b_14_), .ZN(n2789) );
  NAND2_X1 U2680 ( .A1(n2539), .A2(n2538), .ZN(n2783) );
  NAND2_X1 U2681 ( .A1(n2790), .A2(n2791), .ZN(n2538) );
  NAND2_X1 U2682 ( .A1(n2792), .A2(a_4_), .ZN(n2791) );
  NOR2_X1 U2683 ( .A1(n2793), .A2(n2222), .ZN(n2792) );
  NOR2_X1 U2684 ( .A1(n2503), .A2(n2504), .ZN(n2793) );
  NAND2_X1 U2685 ( .A1(n2503), .A2(n2504), .ZN(n2790) );
  NAND2_X1 U2686 ( .A1(n2794), .A2(n2795), .ZN(n2504) );
  NAND2_X1 U2687 ( .A1(n2796), .A2(a_5_), .ZN(n2795) );
  NOR2_X1 U2688 ( .A1(n2797), .A2(n2222), .ZN(n2796) );
  NOR2_X1 U2689 ( .A1(n2476), .A2(n2477), .ZN(n2797) );
  NAND2_X1 U2690 ( .A1(n2476), .A2(n2477), .ZN(n2794) );
  NAND2_X1 U2691 ( .A1(n2798), .A2(n2799), .ZN(n2477) );
  NAND2_X1 U2692 ( .A1(n2800), .A2(a_6_), .ZN(n2799) );
  NOR2_X1 U2693 ( .A1(n2801), .A2(n2222), .ZN(n2800) );
  NOR2_X1 U2694 ( .A1(n2447), .A2(n2449), .ZN(n2801) );
  NAND2_X1 U2695 ( .A1(n2447), .A2(n2449), .ZN(n2798) );
  NAND2_X1 U2696 ( .A1(n2422), .A2(n2802), .ZN(n2449) );
  NAND2_X1 U2697 ( .A1(n2421), .A2(n2423), .ZN(n2802) );
  NAND2_X1 U2698 ( .A1(n2803), .A2(n2804), .ZN(n2423) );
  NAND2_X1 U2699 ( .A1(a_7_), .A2(b_15_), .ZN(n2804) );
  INV_X1 U2700 ( .A(n2805), .ZN(n2803) );
  XOR2_X1 U2701 ( .A(n2806), .B(n2807), .Z(n2421) );
  XNOR2_X1 U2702 ( .A(n2808), .B(n2809), .ZN(n2806) );
  NAND2_X1 U2703 ( .A1(a_8_), .A2(b_14_), .ZN(n2808) );
  NAND2_X1 U2704 ( .A1(a_7_), .A2(n2805), .ZN(n2422) );
  NAND2_X1 U2705 ( .A1(n2810), .A2(n2811), .ZN(n2805) );
  NAND2_X1 U2706 ( .A1(n2812), .A2(a_8_), .ZN(n2811) );
  NOR2_X1 U2707 ( .A1(n2813), .A2(n2222), .ZN(n2812) );
  NOR2_X1 U2708 ( .A1(n2393), .A2(n2395), .ZN(n2813) );
  NAND2_X1 U2709 ( .A1(n2393), .A2(n2395), .ZN(n2810) );
  NAND2_X1 U2710 ( .A1(n2368), .A2(n2814), .ZN(n2395) );
  NAND2_X1 U2711 ( .A1(n2367), .A2(n2369), .ZN(n2814) );
  NAND2_X1 U2712 ( .A1(n2815), .A2(n2816), .ZN(n2369) );
  NAND2_X1 U2713 ( .A1(a_9_), .A2(b_15_), .ZN(n2816) );
  INV_X1 U2714 ( .A(n2817), .ZN(n2815) );
  XOR2_X1 U2715 ( .A(n2818), .B(n2819), .Z(n2367) );
  XOR2_X1 U2716 ( .A(n2820), .B(n2821), .Z(n2818) );
  NOR2_X1 U2717 ( .A1(n2225), .A2(n2687), .ZN(n2821) );
  NAND2_X1 U2718 ( .A1(a_9_), .A2(n2817), .ZN(n2368) );
  NAND2_X1 U2719 ( .A1(n2822), .A2(n2823), .ZN(n2817) );
  NAND2_X1 U2720 ( .A1(n2824), .A2(a_10_), .ZN(n2823) );
  NOR2_X1 U2721 ( .A1(n2825), .A2(n2222), .ZN(n2824) );
  NOR2_X1 U2722 ( .A1(n2338), .A2(n2340), .ZN(n2825) );
  NAND2_X1 U2723 ( .A1(n2338), .A2(n2340), .ZN(n2822) );
  NAND2_X1 U2724 ( .A1(n2826), .A2(n2827), .ZN(n2340) );
  NAND2_X1 U2725 ( .A1(n2828), .A2(a_11_), .ZN(n2827) );
  NOR2_X1 U2726 ( .A1(n2829), .A2(n2222), .ZN(n2828) );
  NOR2_X1 U2727 ( .A1(n2311), .A2(n2312), .ZN(n2829) );
  NAND2_X1 U2728 ( .A1(n2311), .A2(n2312), .ZN(n2826) );
  NAND2_X1 U2729 ( .A1(n2830), .A2(n2831), .ZN(n2312) );
  NAND2_X1 U2730 ( .A1(n2832), .A2(a_12_), .ZN(n2831) );
  NOR2_X1 U2731 ( .A1(n2833), .A2(n2222), .ZN(n2832) );
  NOR2_X1 U2732 ( .A1(n2281), .A2(n2283), .ZN(n2833) );
  NAND2_X1 U2733 ( .A1(n2281), .A2(n2283), .ZN(n2830) );
  NAND2_X1 U2734 ( .A1(n2834), .A2(n2835), .ZN(n2283) );
  NAND2_X1 U2735 ( .A1(n2257), .A2(n2836), .ZN(n2835) );
  OR2_X1 U2736 ( .A1(n2256), .A2(n2255), .ZN(n2836) );
  AND2_X1 U2737 ( .A1(n2837), .A2(n2685), .ZN(n2257) );
  NOR2_X1 U2738 ( .A1(n2222), .A2(n2225), .ZN(n2837) );
  NAND2_X1 U2739 ( .A1(n2255), .A2(n2256), .ZN(n2834) );
  NAND2_X1 U2740 ( .A1(n2838), .A2(n2839), .ZN(n2256) );
  NAND2_X1 U2741 ( .A1(b_13_), .A2(n2840), .ZN(n2839) );
  NAND2_X1 U2742 ( .A1(n2226), .A2(n2841), .ZN(n2840) );
  NAND2_X1 U2743 ( .A1(a_15_), .A2(n2225), .ZN(n2841) );
  NAND2_X1 U2744 ( .A1(b_14_), .A2(n2842), .ZN(n2838) );
  NAND2_X1 U2745 ( .A1(n2843), .A2(n2844), .ZN(n2842) );
  NAND2_X1 U2746 ( .A1(a_14_), .A2(n2686), .ZN(n2844) );
  NOR2_X1 U2747 ( .A1(n2271), .A2(n2222), .ZN(n2255) );
  XNOR2_X1 U2748 ( .A(n2845), .B(n2846), .ZN(n2281) );
  XNOR2_X1 U2749 ( .A(n2847), .B(n2848), .ZN(n2846) );
  XOR2_X1 U2750 ( .A(n2849), .B(n2850), .Z(n2311) );
  XNOR2_X1 U2751 ( .A(n2851), .B(n2852), .ZN(n2849) );
  NAND2_X1 U2752 ( .A1(a_12_), .A2(b_14_), .ZN(n2851) );
  XNOR2_X1 U2753 ( .A(n2853), .B(n2854), .ZN(n2338) );
  XNOR2_X1 U2754 ( .A(n2855), .B(n2856), .ZN(n2854) );
  XNOR2_X1 U2755 ( .A(n2857), .B(n2858), .ZN(n2393) );
  XNOR2_X1 U2756 ( .A(n2859), .B(n2860), .ZN(n2858) );
  XOR2_X1 U2757 ( .A(n2861), .B(n2862), .Z(n2447) );
  XOR2_X1 U2758 ( .A(n2863), .B(n2864), .Z(n2861) );
  XOR2_X1 U2759 ( .A(n2865), .B(n2866), .Z(n2476) );
  XOR2_X1 U2760 ( .A(n2867), .B(n2868), .Z(n2865) );
  NOR2_X1 U2761 ( .A1(n2225), .A2(n2691), .ZN(n2868) );
  XNOR2_X1 U2762 ( .A(n2869), .B(n2870), .ZN(n2503) );
  XNOR2_X1 U2763 ( .A(n2871), .B(n2872), .ZN(n2870) );
  NOR2_X1 U2764 ( .A1(n2553), .A2(n2222), .ZN(n2539) );
  XNOR2_X1 U2765 ( .A(n2873), .B(n2874), .ZN(n2564) );
  XNOR2_X1 U2766 ( .A(n2875), .B(n2876), .ZN(n2874) );
  XNOR2_X1 U2767 ( .A(n2877), .B(n2878), .ZN(n2592) );
  XOR2_X1 U2768 ( .A(n2879), .B(n2880), .Z(n2877) );
  NOR2_X1 U2769 ( .A1(n2225), .A2(n2695), .ZN(n2880) );
  XNOR2_X1 U2770 ( .A(n2881), .B(n2882), .ZN(n2620) );
  XOR2_X1 U2771 ( .A(n2883), .B(n2884), .Z(n2882) );
  NAND2_X1 U2772 ( .A1(a_1_), .A2(b_14_), .ZN(n2884) );
  NOR2_X1 U2773 ( .A1(n2885), .A2(n2886), .ZN(n2765) );
  INV_X1 U2774 ( .A(n2712), .ZN(n2885) );
  NAND2_X1 U2775 ( .A1(n2887), .A2(n2716), .ZN(n2712) );
  NOR2_X1 U2776 ( .A1(n2886), .A2(n2888), .ZN(n2716) );
  AND2_X1 U2777 ( .A1(n2889), .A2(n2890), .ZN(n2888) );
  NOR2_X1 U2778 ( .A1(n2890), .A2(n2889), .ZN(n2886) );
  XNOR2_X1 U2779 ( .A(n2891), .B(n2892), .ZN(n2889) );
  XOR2_X1 U2780 ( .A(n2893), .B(n2894), .Z(n2891) );
  NOR2_X1 U2781 ( .A1(n2623), .A2(n2299), .ZN(n2894) );
  NAND2_X1 U2782 ( .A1(n2895), .A2(n2896), .ZN(n2890) );
  NAND2_X1 U2783 ( .A1(n2897), .A2(n2898), .ZN(n2896) );
  NAND2_X1 U2784 ( .A1(n2899), .A2(n2900), .ZN(n2898) );
  OR2_X1 U2785 ( .A1(n2900), .A2(n2899), .ZN(n2895) );
  AND2_X1 U2786 ( .A1(n2718), .A2(n2717), .ZN(n2887) );
  XNOR2_X1 U2787 ( .A(n2900), .B(n2901), .ZN(n2717) );
  XOR2_X1 U2788 ( .A(n2897), .B(n2899), .Z(n2901) );
  NOR2_X1 U2789 ( .A1(n2686), .A2(n2623), .ZN(n2899) );
  AND2_X1 U2790 ( .A1(n2902), .A2(n2903), .ZN(n2897) );
  NAND2_X1 U2791 ( .A1(n2904), .A2(n2905), .ZN(n2903) );
  OR2_X1 U2792 ( .A1(n2906), .A2(n2907), .ZN(n2905) );
  NAND2_X1 U2793 ( .A1(n2907), .A2(n2906), .ZN(n2902) );
  XNOR2_X1 U2794 ( .A(n2908), .B(n2909), .ZN(n2900) );
  XNOR2_X1 U2795 ( .A(n2910), .B(n2911), .ZN(n2908) );
  NAND2_X1 U2796 ( .A1(n2912), .A2(n2913), .ZN(n2718) );
  NAND2_X1 U2797 ( .A1(n2914), .A2(a_0_), .ZN(n2913) );
  NOR2_X1 U2798 ( .A1(n2915), .A2(n2225), .ZN(n2914) );
  NOR2_X1 U2799 ( .A1(n2769), .A2(n2770), .ZN(n2915) );
  NAND2_X1 U2800 ( .A1(n2769), .A2(n2770), .ZN(n2912) );
  NAND2_X1 U2801 ( .A1(n2916), .A2(n2917), .ZN(n2770) );
  NAND2_X1 U2802 ( .A1(n2918), .A2(a_1_), .ZN(n2917) );
  NOR2_X1 U2803 ( .A1(n2919), .A2(n2225), .ZN(n2918) );
  NOR2_X1 U2804 ( .A1(n2881), .A2(n2883), .ZN(n2919) );
  NAND2_X1 U2805 ( .A1(n2881), .A2(n2883), .ZN(n2916) );
  NAND2_X1 U2806 ( .A1(n2920), .A2(n2921), .ZN(n2883) );
  NAND2_X1 U2807 ( .A1(n2922), .A2(a_2_), .ZN(n2921) );
  NOR2_X1 U2808 ( .A1(n2923), .A2(n2225), .ZN(n2922) );
  NOR2_X1 U2809 ( .A1(n2878), .A2(n2879), .ZN(n2923) );
  NAND2_X1 U2810 ( .A1(n2878), .A2(n2879), .ZN(n2920) );
  NAND2_X1 U2811 ( .A1(n2924), .A2(n2925), .ZN(n2879) );
  NAND2_X1 U2812 ( .A1(n2876), .A2(n2926), .ZN(n2925) );
  OR2_X1 U2813 ( .A1(n2875), .A2(n2873), .ZN(n2926) );
  NOR2_X1 U2814 ( .A1(n2553), .A2(n2225), .ZN(n2876) );
  NAND2_X1 U2815 ( .A1(n2873), .A2(n2875), .ZN(n2924) );
  NAND2_X1 U2816 ( .A1(n2927), .A2(n2928), .ZN(n2875) );
  NAND2_X1 U2817 ( .A1(n2929), .A2(a_4_), .ZN(n2928) );
  NOR2_X1 U2818 ( .A1(n2930), .A2(n2225), .ZN(n2929) );
  NOR2_X1 U2819 ( .A1(n2786), .A2(n2788), .ZN(n2930) );
  NAND2_X1 U2820 ( .A1(n2786), .A2(n2788), .ZN(n2927) );
  NAND2_X1 U2821 ( .A1(n2931), .A2(n2932), .ZN(n2788) );
  NAND2_X1 U2822 ( .A1(n2872), .A2(n2933), .ZN(n2932) );
  OR2_X1 U2823 ( .A1(n2871), .A2(n2869), .ZN(n2933) );
  NOR2_X1 U2824 ( .A1(n2479), .A2(n2225), .ZN(n2872) );
  NAND2_X1 U2825 ( .A1(n2869), .A2(n2871), .ZN(n2931) );
  NAND2_X1 U2826 ( .A1(n2934), .A2(n2935), .ZN(n2871) );
  NAND2_X1 U2827 ( .A1(n2936), .A2(a_6_), .ZN(n2935) );
  NOR2_X1 U2828 ( .A1(n2937), .A2(n2225), .ZN(n2936) );
  NOR2_X1 U2829 ( .A1(n2866), .A2(n2867), .ZN(n2937) );
  NAND2_X1 U2830 ( .A1(n2866), .A2(n2867), .ZN(n2934) );
  NAND2_X1 U2831 ( .A1(n2938), .A2(n2939), .ZN(n2867) );
  NAND2_X1 U2832 ( .A1(n2864), .A2(n2940), .ZN(n2939) );
  OR2_X1 U2833 ( .A1(n2863), .A2(n2862), .ZN(n2940) );
  NOR2_X1 U2834 ( .A1(n2437), .A2(n2225), .ZN(n2864) );
  NAND2_X1 U2835 ( .A1(n2862), .A2(n2863), .ZN(n2938) );
  NAND2_X1 U2836 ( .A1(n2941), .A2(n2942), .ZN(n2863) );
  NAND2_X1 U2837 ( .A1(n2943), .A2(a_8_), .ZN(n2942) );
  NOR2_X1 U2838 ( .A1(n2944), .A2(n2225), .ZN(n2943) );
  NOR2_X1 U2839 ( .A1(n2807), .A2(n2809), .ZN(n2944) );
  NAND2_X1 U2840 ( .A1(n2807), .A2(n2809), .ZN(n2941) );
  NAND2_X1 U2841 ( .A1(n2945), .A2(n2946), .ZN(n2809) );
  NAND2_X1 U2842 ( .A1(n2860), .A2(n2947), .ZN(n2946) );
  OR2_X1 U2843 ( .A1(n2859), .A2(n2857), .ZN(n2947) );
  NOR2_X1 U2844 ( .A1(n2383), .A2(n2225), .ZN(n2860) );
  NAND2_X1 U2845 ( .A1(n2857), .A2(n2859), .ZN(n2945) );
  NAND2_X1 U2846 ( .A1(n2948), .A2(n2949), .ZN(n2859) );
  NAND2_X1 U2847 ( .A1(n2950), .A2(a_10_), .ZN(n2949) );
  NOR2_X1 U2848 ( .A1(n2951), .A2(n2225), .ZN(n2950) );
  NOR2_X1 U2849 ( .A1(n2819), .A2(n2820), .ZN(n2951) );
  NAND2_X1 U2850 ( .A1(n2819), .A2(n2820), .ZN(n2948) );
  NAND2_X1 U2851 ( .A1(n2952), .A2(n2953), .ZN(n2820) );
  NAND2_X1 U2852 ( .A1(n2856), .A2(n2954), .ZN(n2953) );
  OR2_X1 U2853 ( .A1(n2855), .A2(n2853), .ZN(n2954) );
  NOR2_X1 U2854 ( .A1(n2314), .A2(n2225), .ZN(n2856) );
  NAND2_X1 U2855 ( .A1(n2853), .A2(n2855), .ZN(n2952) );
  NAND2_X1 U2856 ( .A1(n2955), .A2(n2956), .ZN(n2855) );
  NAND2_X1 U2857 ( .A1(n2957), .A2(a_12_), .ZN(n2956) );
  NOR2_X1 U2858 ( .A1(n2958), .A2(n2225), .ZN(n2957) );
  NOR2_X1 U2859 ( .A1(n2850), .A2(n2852), .ZN(n2958) );
  NAND2_X1 U2860 ( .A1(n2850), .A2(n2852), .ZN(n2955) );
  NAND2_X1 U2861 ( .A1(n2959), .A2(n2960), .ZN(n2852) );
  NAND2_X1 U2862 ( .A1(n2845), .A2(n2961), .ZN(n2960) );
  NAND2_X1 U2863 ( .A1(n2848), .A2(n2847), .ZN(n2961) );
  NOR2_X1 U2864 ( .A1(n2271), .A2(n2225), .ZN(n2845) );
  OR2_X1 U2865 ( .A1(n2847), .A2(n2848), .ZN(n2959) );
  AND2_X1 U2866 ( .A1(n2962), .A2(n2963), .ZN(n2848) );
  NAND2_X1 U2867 ( .A1(b_12_), .A2(n2964), .ZN(n2963) );
  NAND2_X1 U2868 ( .A1(n2226), .A2(n2965), .ZN(n2964) );
  NAND2_X1 U2869 ( .A1(a_15_), .A2(n2686), .ZN(n2965) );
  NAND2_X1 U2870 ( .A1(b_13_), .A2(n2966), .ZN(n2962) );
  NAND2_X1 U2871 ( .A1(n2843), .A2(n2967), .ZN(n2966) );
  NAND2_X1 U2872 ( .A1(a_14_), .A2(n2299), .ZN(n2967) );
  NAND2_X1 U2873 ( .A1(n2968), .A2(n2685), .ZN(n2847) );
  NOR2_X1 U2874 ( .A1(n2225), .A2(n2686), .ZN(n2968) );
  XNOR2_X1 U2875 ( .A(n2678), .B(n2969), .ZN(n2850) );
  XNOR2_X1 U2876 ( .A(n2970), .B(n2971), .ZN(n2969) );
  XOR2_X1 U2877 ( .A(n2972), .B(n2973), .Z(n2853) );
  XNOR2_X1 U2878 ( .A(n2974), .B(n2975), .ZN(n2972) );
  NAND2_X1 U2879 ( .A1(b_13_), .A2(a_12_), .ZN(n2974) );
  XNOR2_X1 U2880 ( .A(n2976), .B(n2977), .ZN(n2819) );
  NAND2_X1 U2881 ( .A1(n2978), .A2(n2979), .ZN(n2976) );
  XNOR2_X1 U2882 ( .A(n2980), .B(n2981), .ZN(n2857) );
  NAND2_X1 U2883 ( .A1(n2982), .A2(n2983), .ZN(n2980) );
  XNOR2_X1 U2884 ( .A(n2984), .B(n2985), .ZN(n2807) );
  XNOR2_X1 U2885 ( .A(n2986), .B(n2987), .ZN(n2984) );
  XNOR2_X1 U2886 ( .A(n2988), .B(n2989), .ZN(n2862) );
  XOR2_X1 U2887 ( .A(n2990), .B(n2991), .Z(n2989) );
  NAND2_X1 U2888 ( .A1(b_13_), .A2(a_8_), .ZN(n2991) );
  XNOR2_X1 U2889 ( .A(n2992), .B(n2993), .ZN(n2866) );
  XOR2_X1 U2890 ( .A(n2994), .B(n2995), .Z(n2993) );
  NAND2_X1 U2891 ( .A1(b_13_), .A2(a_7_), .ZN(n2995) );
  XNOR2_X1 U2892 ( .A(n2996), .B(n2997), .ZN(n2869) );
  NAND2_X1 U2893 ( .A1(n2998), .A2(n2999), .ZN(n2996) );
  XNOR2_X1 U2894 ( .A(n3000), .B(n3001), .ZN(n2786) );
  XNOR2_X1 U2895 ( .A(n3002), .B(n3003), .ZN(n3001) );
  XNOR2_X1 U2896 ( .A(n3004), .B(n3005), .ZN(n2873) );
  XOR2_X1 U2897 ( .A(n3006), .B(n3007), .Z(n3005) );
  NAND2_X1 U2898 ( .A1(b_13_), .A2(a_4_), .ZN(n3007) );
  XNOR2_X1 U2899 ( .A(n3008), .B(n3009), .ZN(n2878) );
  XOR2_X1 U2900 ( .A(n3010), .B(n3011), .Z(n3009) );
  NAND2_X1 U2901 ( .A1(b_13_), .A2(a_3_), .ZN(n3011) );
  XNOR2_X1 U2902 ( .A(n3012), .B(n3013), .ZN(n2881) );
  NAND2_X1 U2903 ( .A1(n3014), .A2(n3015), .ZN(n3012) );
  XNOR2_X1 U2904 ( .A(n2907), .B(n3016), .ZN(n2769) );
  XNOR2_X1 U2905 ( .A(n2906), .B(n2904), .ZN(n3016) );
  NOR2_X1 U2906 ( .A1(n2686), .A2(n2609), .ZN(n2904) );
  NAND2_X1 U2907 ( .A1(n3014), .A2(n3017), .ZN(n2906) );
  NAND2_X1 U2908 ( .A1(n3013), .A2(n3015), .ZN(n3017) );
  NAND2_X1 U2909 ( .A1(n3018), .A2(n3019), .ZN(n3015) );
  NAND2_X1 U2910 ( .A1(b_13_), .A2(a_2_), .ZN(n3019) );
  INV_X1 U2911 ( .A(n3020), .ZN(n3018) );
  XOR2_X1 U2912 ( .A(n3021), .B(n3022), .Z(n3013) );
  XOR2_X1 U2913 ( .A(n3023), .B(n3024), .Z(n3021) );
  NOR2_X1 U2914 ( .A1(n2553), .A2(n2299), .ZN(n3024) );
  NAND2_X1 U2915 ( .A1(a_2_), .A2(n3020), .ZN(n3014) );
  NAND2_X1 U2916 ( .A1(n3025), .A2(n3026), .ZN(n3020) );
  NAND2_X1 U2917 ( .A1(n3027), .A2(b_13_), .ZN(n3026) );
  NOR2_X1 U2918 ( .A1(n3028), .A2(n2553), .ZN(n3027) );
  NOR2_X1 U2919 ( .A1(n3008), .A2(n3010), .ZN(n3028) );
  NAND2_X1 U2920 ( .A1(n3008), .A2(n3010), .ZN(n3025) );
  NAND2_X1 U2921 ( .A1(n3029), .A2(n3030), .ZN(n3010) );
  NAND2_X1 U2922 ( .A1(n3031), .A2(b_13_), .ZN(n3030) );
  NOR2_X1 U2923 ( .A1(n3032), .A2(n2506), .ZN(n3031) );
  NOR2_X1 U2924 ( .A1(n3004), .A2(n3006), .ZN(n3032) );
  NAND2_X1 U2925 ( .A1(n3004), .A2(n3006), .ZN(n3029) );
  NAND2_X1 U2926 ( .A1(n3033), .A2(n3034), .ZN(n3006) );
  NAND2_X1 U2927 ( .A1(n3003), .A2(n3035), .ZN(n3034) );
  OR2_X1 U2928 ( .A1(n3002), .A2(n3000), .ZN(n3035) );
  NOR2_X1 U2929 ( .A1(n2686), .A2(n2479), .ZN(n3003) );
  NAND2_X1 U2930 ( .A1(n3000), .A2(n3002), .ZN(n3033) );
  NAND2_X1 U2931 ( .A1(n2998), .A2(n3036), .ZN(n3002) );
  NAND2_X1 U2932 ( .A1(n2997), .A2(n2999), .ZN(n3036) );
  NAND2_X1 U2933 ( .A1(n3037), .A2(n3038), .ZN(n2999) );
  NAND2_X1 U2934 ( .A1(b_13_), .A2(a_6_), .ZN(n3038) );
  INV_X1 U2935 ( .A(n3039), .ZN(n3037) );
  XNOR2_X1 U2936 ( .A(n3040), .B(n3041), .ZN(n2997) );
  XNOR2_X1 U2937 ( .A(n3042), .B(n3043), .ZN(n3041) );
  NAND2_X1 U2938 ( .A1(a_6_), .A2(n3039), .ZN(n2998) );
  NAND2_X1 U2939 ( .A1(n3044), .A2(n3045), .ZN(n3039) );
  NAND2_X1 U2940 ( .A1(n3046), .A2(b_13_), .ZN(n3045) );
  NOR2_X1 U2941 ( .A1(n3047), .A2(n2437), .ZN(n3046) );
  NOR2_X1 U2942 ( .A1(n2992), .A2(n2994), .ZN(n3047) );
  NAND2_X1 U2943 ( .A1(n2992), .A2(n2994), .ZN(n3044) );
  NAND2_X1 U2944 ( .A1(n3048), .A2(n3049), .ZN(n2994) );
  NAND2_X1 U2945 ( .A1(n3050), .A2(b_13_), .ZN(n3049) );
  NOR2_X1 U2946 ( .A1(n3051), .A2(n2689), .ZN(n3050) );
  NOR2_X1 U2947 ( .A1(n2988), .A2(n2990), .ZN(n3051) );
  NAND2_X1 U2948 ( .A1(n2988), .A2(n2990), .ZN(n3048) );
  NAND2_X1 U2949 ( .A1(n3052), .A2(n3053), .ZN(n2990) );
  NAND2_X1 U2950 ( .A1(n2987), .A2(n3054), .ZN(n3053) );
  NAND2_X1 U2951 ( .A1(n2986), .A2(n2985), .ZN(n3054) );
  NOR2_X1 U2952 ( .A1(n2686), .A2(n2383), .ZN(n2987) );
  OR2_X1 U2953 ( .A1(n2985), .A2(n2986), .ZN(n3052) );
  AND2_X1 U2954 ( .A1(n2982), .A2(n3055), .ZN(n2986) );
  NAND2_X1 U2955 ( .A1(n2981), .A2(n2983), .ZN(n3055) );
  NAND2_X1 U2956 ( .A1(n3056), .A2(n3057), .ZN(n2983) );
  NAND2_X1 U2957 ( .A1(b_13_), .A2(a_10_), .ZN(n3057) );
  INV_X1 U2958 ( .A(n3058), .ZN(n3056) );
  XNOR2_X1 U2959 ( .A(n3059), .B(n3060), .ZN(n2981) );
  NAND2_X1 U2960 ( .A1(n3061), .A2(n3062), .ZN(n3059) );
  NAND2_X1 U2961 ( .A1(a_10_), .A2(n3058), .ZN(n2982) );
  NAND2_X1 U2962 ( .A1(n2978), .A2(n3063), .ZN(n3058) );
  NAND2_X1 U2963 ( .A1(n2977), .A2(n2979), .ZN(n3063) );
  NAND2_X1 U2964 ( .A1(n3064), .A2(n3065), .ZN(n2979) );
  NAND2_X1 U2965 ( .A1(b_13_), .A2(a_11_), .ZN(n3065) );
  INV_X1 U2966 ( .A(n3066), .ZN(n3064) );
  XOR2_X1 U2967 ( .A(n3067), .B(n3068), .Z(n2977) );
  XOR2_X1 U2968 ( .A(n2675), .B(n3069), .Z(n3067) );
  NAND2_X1 U2969 ( .A1(a_11_), .A2(n3066), .ZN(n2978) );
  NAND2_X1 U2970 ( .A1(n3070), .A2(n3071), .ZN(n3066) );
  NAND2_X1 U2971 ( .A1(n3072), .A2(b_13_), .ZN(n3071) );
  NOR2_X1 U2972 ( .A1(n3073), .A2(n2285), .ZN(n3072) );
  NOR2_X1 U2973 ( .A1(n2973), .A2(n2975), .ZN(n3073) );
  NAND2_X1 U2974 ( .A1(n2973), .A2(n2975), .ZN(n3070) );
  NAND2_X1 U2975 ( .A1(n3074), .A2(n3075), .ZN(n2975) );
  NAND2_X1 U2976 ( .A1(n2678), .A2(n3076), .ZN(n3075) );
  NAND2_X1 U2977 ( .A1(n2971), .A2(n2970), .ZN(n3076) );
  NOR2_X1 U2978 ( .A1(n2686), .A2(n2271), .ZN(n2678) );
  OR2_X1 U2979 ( .A1(n2970), .A2(n2971), .ZN(n3074) );
  AND2_X1 U2980 ( .A1(n3077), .A2(n3078), .ZN(n2971) );
  NAND2_X1 U2981 ( .A1(b_11_), .A2(n3079), .ZN(n3078) );
  NAND2_X1 U2982 ( .A1(n2226), .A2(n3080), .ZN(n3079) );
  NAND2_X1 U2983 ( .A1(a_15_), .A2(n2299), .ZN(n3080) );
  NAND2_X1 U2984 ( .A1(b_12_), .A2(n3081), .ZN(n3077) );
  NAND2_X1 U2985 ( .A1(n2843), .A2(n3082), .ZN(n3081) );
  NAND2_X1 U2986 ( .A1(a_14_), .A2(n2328), .ZN(n3082) );
  NAND2_X1 U2987 ( .A1(n3083), .A2(n2685), .ZN(n2970) );
  NOR2_X1 U2988 ( .A1(n2686), .A2(n2299), .ZN(n3083) );
  XNOR2_X1 U2989 ( .A(n3084), .B(n3085), .ZN(n2973) );
  XNOR2_X1 U2990 ( .A(n3086), .B(n3087), .ZN(n3085) );
  XOR2_X1 U2991 ( .A(n3088), .B(n3089), .Z(n2985) );
  NAND2_X1 U2992 ( .A1(n3090), .A2(n3091), .ZN(n3088) );
  XNOR2_X1 U2993 ( .A(n3092), .B(n3093), .ZN(n2988) );
  XNOR2_X1 U2994 ( .A(n3094), .B(n3095), .ZN(n3093) );
  XNOR2_X1 U2995 ( .A(n3096), .B(n3097), .ZN(n2992) );
  XOR2_X1 U2996 ( .A(n3098), .B(n3099), .Z(n3097) );
  NAND2_X1 U2997 ( .A1(b_12_), .A2(a_8_), .ZN(n3099) );
  XOR2_X1 U2998 ( .A(n3100), .B(n3101), .Z(n3000) );
  XOR2_X1 U2999 ( .A(n3102), .B(n3103), .Z(n3100) );
  NOR2_X1 U3000 ( .A1(n2691), .A2(n2299), .ZN(n3103) );
  XOR2_X1 U3001 ( .A(n3104), .B(n3105), .Z(n3004) );
  XOR2_X1 U3002 ( .A(n3106), .B(n3107), .Z(n3104) );
  XNOR2_X1 U3003 ( .A(n3108), .B(n3109), .ZN(n3008) );
  XOR2_X1 U3004 ( .A(n3110), .B(n3111), .Z(n3109) );
  NAND2_X1 U3005 ( .A1(b_12_), .A2(a_4_), .ZN(n3111) );
  XOR2_X1 U3006 ( .A(n3112), .B(n3113), .Z(n2907) );
  XOR2_X1 U3007 ( .A(n3114), .B(n3115), .Z(n3112) );
  XOR2_X1 U3008 ( .A(n2764), .B(n3116), .Z(n2721) );
  NAND2_X1 U3009 ( .A1(n3117), .A2(n3118), .ZN(n2727) );
  AND2_X1 U3010 ( .A1(n2754), .A2(n2764), .ZN(n3118) );
  NAND2_X1 U3011 ( .A1(n3119), .A2(n3120), .ZN(n2764) );
  NAND2_X1 U3012 ( .A1(n3121), .A2(b_12_), .ZN(n3120) );
  NOR2_X1 U3013 ( .A1(n3122), .A2(n2623), .ZN(n3121) );
  NOR2_X1 U3014 ( .A1(n2892), .A2(n2893), .ZN(n3122) );
  NAND2_X1 U3015 ( .A1(n2892), .A2(n2893), .ZN(n3119) );
  NAND2_X1 U3016 ( .A1(n3123), .A2(n3124), .ZN(n2893) );
  NAND2_X1 U3017 ( .A1(n2911), .A2(n3125), .ZN(n3124) );
  NAND2_X1 U3018 ( .A1(n2910), .A2(n2909), .ZN(n3125) );
  NOR2_X1 U3019 ( .A1(n2299), .A2(n2609), .ZN(n2911) );
  OR2_X1 U3020 ( .A1(n2909), .A2(n2910), .ZN(n3123) );
  AND2_X1 U3021 ( .A1(n3126), .A2(n3127), .ZN(n2910) );
  NAND2_X1 U3022 ( .A1(n3115), .A2(n3128), .ZN(n3127) );
  OR2_X1 U3023 ( .A1(n3114), .A2(n3113), .ZN(n3128) );
  NOR2_X1 U3024 ( .A1(n2299), .A2(n2695), .ZN(n3115) );
  NAND2_X1 U3025 ( .A1(n3113), .A2(n3114), .ZN(n3126) );
  NAND2_X1 U3026 ( .A1(n3129), .A2(n3130), .ZN(n3114) );
  NAND2_X1 U3027 ( .A1(n3131), .A2(b_12_), .ZN(n3130) );
  NOR2_X1 U3028 ( .A1(n3132), .A2(n2553), .ZN(n3131) );
  NOR2_X1 U3029 ( .A1(n3022), .A2(n3023), .ZN(n3132) );
  NAND2_X1 U3030 ( .A1(n3022), .A2(n3023), .ZN(n3129) );
  NAND2_X1 U3031 ( .A1(n3133), .A2(n3134), .ZN(n3023) );
  NAND2_X1 U3032 ( .A1(n3135), .A2(b_12_), .ZN(n3134) );
  NOR2_X1 U3033 ( .A1(n3136), .A2(n2506), .ZN(n3135) );
  NOR2_X1 U3034 ( .A1(n3108), .A2(n3110), .ZN(n3136) );
  NAND2_X1 U3035 ( .A1(n3108), .A2(n3110), .ZN(n3133) );
  NAND2_X1 U3036 ( .A1(n3137), .A2(n3138), .ZN(n3110) );
  NAND2_X1 U3037 ( .A1(n3107), .A2(n3139), .ZN(n3138) );
  OR2_X1 U3038 ( .A1(n3106), .A2(n3105), .ZN(n3139) );
  NOR2_X1 U3039 ( .A1(n2299), .A2(n2479), .ZN(n3107) );
  NAND2_X1 U3040 ( .A1(n3105), .A2(n3106), .ZN(n3137) );
  NAND2_X1 U3041 ( .A1(n3140), .A2(n3141), .ZN(n3106) );
  NAND2_X1 U3042 ( .A1(n3142), .A2(b_12_), .ZN(n3141) );
  NOR2_X1 U3043 ( .A1(n3143), .A2(n2691), .ZN(n3142) );
  NOR2_X1 U3044 ( .A1(n3101), .A2(n3102), .ZN(n3143) );
  NAND2_X1 U3045 ( .A1(n3101), .A2(n3102), .ZN(n3140) );
  NAND2_X1 U3046 ( .A1(n3144), .A2(n3145), .ZN(n3102) );
  NAND2_X1 U3047 ( .A1(n3043), .A2(n3146), .ZN(n3145) );
  OR2_X1 U3048 ( .A1(n3042), .A2(n3040), .ZN(n3146) );
  NOR2_X1 U3049 ( .A1(n2299), .A2(n2437), .ZN(n3043) );
  NAND2_X1 U3050 ( .A1(n3040), .A2(n3042), .ZN(n3144) );
  NAND2_X1 U3051 ( .A1(n3147), .A2(n3148), .ZN(n3042) );
  NAND2_X1 U3052 ( .A1(n3149), .A2(b_12_), .ZN(n3148) );
  NOR2_X1 U3053 ( .A1(n3150), .A2(n2689), .ZN(n3149) );
  NOR2_X1 U3054 ( .A1(n3096), .A2(n3098), .ZN(n3150) );
  NAND2_X1 U3055 ( .A1(n3096), .A2(n3098), .ZN(n3147) );
  NAND2_X1 U3056 ( .A1(n3151), .A2(n3152), .ZN(n3098) );
  NAND2_X1 U3057 ( .A1(n3095), .A2(n3153), .ZN(n3152) );
  OR2_X1 U3058 ( .A1(n3094), .A2(n3092), .ZN(n3153) );
  NOR2_X1 U3059 ( .A1(n2299), .A2(n2383), .ZN(n3095) );
  NAND2_X1 U3060 ( .A1(n3092), .A2(n3094), .ZN(n3151) );
  NAND2_X1 U3061 ( .A1(n3090), .A2(n3154), .ZN(n3094) );
  NAND2_X1 U3062 ( .A1(n3089), .A2(n3091), .ZN(n3154) );
  NAND2_X1 U3063 ( .A1(n3155), .A2(n3156), .ZN(n3091) );
  NAND2_X1 U3064 ( .A1(b_12_), .A2(a_10_), .ZN(n3156) );
  INV_X1 U3065 ( .A(n3157), .ZN(n3155) );
  XNOR2_X1 U3066 ( .A(n3158), .B(n3159), .ZN(n3089) );
  XNOR2_X1 U3067 ( .A(n3160), .B(n2672), .ZN(n3159) );
  NAND2_X1 U3068 ( .A1(a_10_), .A2(n3157), .ZN(n3090) );
  NAND2_X1 U3069 ( .A1(n3061), .A2(n3161), .ZN(n3157) );
  NAND2_X1 U3070 ( .A1(n3060), .A2(n3062), .ZN(n3161) );
  NAND2_X1 U3071 ( .A1(n3162), .A2(n3163), .ZN(n3062) );
  NAND2_X1 U3072 ( .A1(b_12_), .A2(a_11_), .ZN(n3163) );
  INV_X1 U3073 ( .A(n3164), .ZN(n3162) );
  XOR2_X1 U3074 ( .A(n3165), .B(n3166), .Z(n3060) );
  XNOR2_X1 U3075 ( .A(n3167), .B(n3168), .ZN(n3165) );
  NAND2_X1 U3076 ( .A1(b_11_), .A2(a_12_), .ZN(n3167) );
  NAND2_X1 U3077 ( .A1(a_11_), .A2(n3164), .ZN(n3061) );
  NAND2_X1 U3078 ( .A1(n3169), .A2(n3170), .ZN(n3164) );
  NAND2_X1 U3079 ( .A1(n3068), .A2(n3171), .ZN(n3170) );
  NAND2_X1 U3080 ( .A1(n3069), .A2(n2675), .ZN(n3171) );
  INV_X1 U3081 ( .A(n3172), .ZN(n3069) );
  XNOR2_X1 U3082 ( .A(n3173), .B(n3174), .ZN(n3068) );
  XNOR2_X1 U3083 ( .A(n3175), .B(n3176), .ZN(n3174) );
  NAND2_X1 U3084 ( .A1(n3177), .A2(n3172), .ZN(n3169) );
  NAND2_X1 U3085 ( .A1(n3178), .A2(n3179), .ZN(n3172) );
  NAND2_X1 U3086 ( .A1(n3084), .A2(n3180), .ZN(n3179) );
  NAND2_X1 U3087 ( .A1(n3087), .A2(n3086), .ZN(n3180) );
  NOR2_X1 U3088 ( .A1(n2299), .A2(n2271), .ZN(n3084) );
  OR2_X1 U3089 ( .A1(n3086), .A2(n3087), .ZN(n3178) );
  AND2_X1 U3090 ( .A1(n3181), .A2(n3182), .ZN(n3087) );
  NAND2_X1 U3091 ( .A1(b_10_), .A2(n3183), .ZN(n3182) );
  NAND2_X1 U3092 ( .A1(n2226), .A2(n3184), .ZN(n3183) );
  NAND2_X1 U3093 ( .A1(a_15_), .A2(n2328), .ZN(n3184) );
  NAND2_X1 U3094 ( .A1(b_11_), .A2(n3185), .ZN(n3181) );
  NAND2_X1 U3095 ( .A1(n2843), .A2(n3186), .ZN(n3185) );
  NAND2_X1 U3096 ( .A1(a_14_), .A2(n2355), .ZN(n3186) );
  NAND2_X1 U3097 ( .A1(n3187), .A2(n2685), .ZN(n3086) );
  NOR2_X1 U3098 ( .A1(n2299), .A2(n2328), .ZN(n3187) );
  INV_X1 U3099 ( .A(n2675), .ZN(n3177) );
  NAND2_X1 U3100 ( .A1(b_12_), .A2(a_12_), .ZN(n2675) );
  XOR2_X1 U3101 ( .A(n3188), .B(n3189), .Z(n3092) );
  XOR2_X1 U3102 ( .A(n3190), .B(n3191), .Z(n3188) );
  NOR2_X1 U3103 ( .A1(n2687), .A2(n2328), .ZN(n3191) );
  XOR2_X1 U3104 ( .A(n3192), .B(n3193), .Z(n3096) );
  XOR2_X1 U3105 ( .A(n3194), .B(n3195), .Z(n3192) );
  XOR2_X1 U3106 ( .A(n3196), .B(n3197), .Z(n3040) );
  XOR2_X1 U3107 ( .A(n3198), .B(n3199), .Z(n3196) );
  NOR2_X1 U3108 ( .A1(n2689), .A2(n2328), .ZN(n3199) );
  XNOR2_X1 U3109 ( .A(n3200), .B(n3201), .ZN(n3101) );
  XNOR2_X1 U3110 ( .A(n3202), .B(n3203), .ZN(n3201) );
  XOR2_X1 U3111 ( .A(n3204), .B(n3205), .Z(n3105) );
  XOR2_X1 U3112 ( .A(n3206), .B(n3207), .Z(n3204) );
  NOR2_X1 U3113 ( .A1(n2691), .A2(n2328), .ZN(n3207) );
  XNOR2_X1 U3114 ( .A(n3208), .B(n3209), .ZN(n3108) );
  XNOR2_X1 U3115 ( .A(n3210), .B(n3211), .ZN(n3209) );
  XNOR2_X1 U3116 ( .A(n3212), .B(n3213), .ZN(n3022) );
  XNOR2_X1 U3117 ( .A(n3214), .B(n3215), .ZN(n3212) );
  XNOR2_X1 U3118 ( .A(n3216), .B(n3217), .ZN(n3113) );
  XOR2_X1 U3119 ( .A(n3218), .B(n3219), .Z(n3217) );
  NAND2_X1 U3120 ( .A1(b_11_), .A2(a_3_), .ZN(n3219) );
  XOR2_X1 U3121 ( .A(n3220), .B(n3221), .Z(n2909) );
  NAND2_X1 U3122 ( .A1(n3222), .A2(n3223), .ZN(n3220) );
  XOR2_X1 U3123 ( .A(n3224), .B(n3225), .Z(n2892) );
  XOR2_X1 U3124 ( .A(n3226), .B(n3227), .Z(n3224) );
  NOR2_X1 U3125 ( .A1(n2609), .A2(n2328), .ZN(n3227) );
  INV_X1 U3126 ( .A(n3228), .ZN(n2754) );
  NOR2_X1 U3127 ( .A1(n3229), .A2(n3116), .ZN(n3117) );
  INV_X1 U3128 ( .A(n2763), .ZN(n3116) );
  XOR2_X1 U3129 ( .A(n3230), .B(n3231), .Z(n2763) );
  XNOR2_X1 U3130 ( .A(n3232), .B(n3233), .ZN(n3231) );
  AND2_X1 U3131 ( .A1(n2762), .A2(n2761), .ZN(n3229) );
  NAND2_X1 U3132 ( .A1(n3228), .A2(n3234), .ZN(n2733) );
  XOR2_X1 U3133 ( .A(n3235), .B(n2756), .Z(n3234) );
  INV_X1 U3134 ( .A(n3236), .ZN(n2756) );
  NOR2_X1 U3135 ( .A1(n2762), .A2(n2761), .ZN(n3228) );
  XOR2_X1 U3136 ( .A(n3237), .B(n3238), .Z(n2761) );
  NAND2_X1 U3137 ( .A1(n3239), .A2(n3240), .ZN(n3237) );
  NAND2_X1 U3138 ( .A1(n3241), .A2(n3242), .ZN(n2762) );
  NAND2_X1 U3139 ( .A1(n3230), .A2(n3243), .ZN(n3242) );
  NAND2_X1 U3140 ( .A1(n3233), .A2(n3232), .ZN(n3243) );
  XNOR2_X1 U3141 ( .A(n3244), .B(n3245), .ZN(n3230) );
  XOR2_X1 U3142 ( .A(n3246), .B(n3247), .Z(n3245) );
  OR2_X1 U3143 ( .A1(n3232), .A2(n3233), .ZN(n3241) );
  NOR2_X1 U3144 ( .A1(n2328), .A2(n2623), .ZN(n3233) );
  NAND2_X1 U3145 ( .A1(n3248), .A2(n3249), .ZN(n3232) );
  NAND2_X1 U3146 ( .A1(n3250), .A2(b_11_), .ZN(n3249) );
  NOR2_X1 U3147 ( .A1(n3251), .A2(n2609), .ZN(n3250) );
  NOR2_X1 U3148 ( .A1(n3225), .A2(n3226), .ZN(n3251) );
  NAND2_X1 U3149 ( .A1(n3225), .A2(n3226), .ZN(n3248) );
  NAND2_X1 U3150 ( .A1(n3222), .A2(n3252), .ZN(n3226) );
  NAND2_X1 U3151 ( .A1(n3221), .A2(n3223), .ZN(n3252) );
  NAND2_X1 U3152 ( .A1(n3253), .A2(n3254), .ZN(n3223) );
  NAND2_X1 U3153 ( .A1(b_11_), .A2(a_2_), .ZN(n3254) );
  INV_X1 U3154 ( .A(n3255), .ZN(n3253) );
  XOR2_X1 U3155 ( .A(n3256), .B(n3257), .Z(n3221) );
  XOR2_X1 U3156 ( .A(n3258), .B(n3259), .Z(n3256) );
  NAND2_X1 U3157 ( .A1(a_2_), .A2(n3255), .ZN(n3222) );
  NAND2_X1 U3158 ( .A1(n3260), .A2(n3261), .ZN(n3255) );
  NAND2_X1 U3159 ( .A1(n3262), .A2(b_11_), .ZN(n3261) );
  NOR2_X1 U3160 ( .A1(n3263), .A2(n2553), .ZN(n3262) );
  NOR2_X1 U3161 ( .A1(n3216), .A2(n3218), .ZN(n3263) );
  NAND2_X1 U3162 ( .A1(n3216), .A2(n3218), .ZN(n3260) );
  NAND2_X1 U3163 ( .A1(n3264), .A2(n3265), .ZN(n3218) );
  NAND2_X1 U3164 ( .A1(n3215), .A2(n3266), .ZN(n3265) );
  NAND2_X1 U3165 ( .A1(n3214), .A2(n3213), .ZN(n3266) );
  NOR2_X1 U3166 ( .A1(n2328), .A2(n2506), .ZN(n3215) );
  OR2_X1 U3167 ( .A1(n3213), .A2(n3214), .ZN(n3264) );
  AND2_X1 U3168 ( .A1(n3267), .A2(n3268), .ZN(n3214) );
  NAND2_X1 U3169 ( .A1(n3211), .A2(n3269), .ZN(n3268) );
  OR2_X1 U3170 ( .A1(n3210), .A2(n3208), .ZN(n3269) );
  NOR2_X1 U3171 ( .A1(n2328), .A2(n2479), .ZN(n3211) );
  NAND2_X1 U3172 ( .A1(n3208), .A2(n3210), .ZN(n3267) );
  NAND2_X1 U3173 ( .A1(n3270), .A2(n3271), .ZN(n3210) );
  NAND2_X1 U3174 ( .A1(n3272), .A2(b_11_), .ZN(n3271) );
  NOR2_X1 U3175 ( .A1(n3273), .A2(n2691), .ZN(n3272) );
  NOR2_X1 U3176 ( .A1(n3205), .A2(n3206), .ZN(n3273) );
  NAND2_X1 U3177 ( .A1(n3205), .A2(n3206), .ZN(n3270) );
  NAND2_X1 U3178 ( .A1(n3274), .A2(n3275), .ZN(n3206) );
  NAND2_X1 U3179 ( .A1(n3203), .A2(n3276), .ZN(n3275) );
  OR2_X1 U3180 ( .A1(n3202), .A2(n3200), .ZN(n3276) );
  NOR2_X1 U3181 ( .A1(n2328), .A2(n2437), .ZN(n3203) );
  NAND2_X1 U3182 ( .A1(n3200), .A2(n3202), .ZN(n3274) );
  NAND2_X1 U3183 ( .A1(n3277), .A2(n3278), .ZN(n3202) );
  NAND2_X1 U3184 ( .A1(n3279), .A2(b_11_), .ZN(n3278) );
  NOR2_X1 U3185 ( .A1(n3280), .A2(n2689), .ZN(n3279) );
  NOR2_X1 U3186 ( .A1(n3197), .A2(n3198), .ZN(n3280) );
  NAND2_X1 U3187 ( .A1(n3197), .A2(n3198), .ZN(n3277) );
  NAND2_X1 U3188 ( .A1(n3281), .A2(n3282), .ZN(n3198) );
  NAND2_X1 U3189 ( .A1(n3195), .A2(n3283), .ZN(n3282) );
  OR2_X1 U3190 ( .A1(n3194), .A2(n3193), .ZN(n3283) );
  NOR2_X1 U3191 ( .A1(n2328), .A2(n2383), .ZN(n3195) );
  NAND2_X1 U3192 ( .A1(n3193), .A2(n3194), .ZN(n3281) );
  NAND2_X1 U3193 ( .A1(n3284), .A2(n3285), .ZN(n3194) );
  NAND2_X1 U3194 ( .A1(n3286), .A2(b_11_), .ZN(n3285) );
  NOR2_X1 U3195 ( .A1(n3287), .A2(n2687), .ZN(n3286) );
  NOR2_X1 U3196 ( .A1(n3189), .A2(n3190), .ZN(n3287) );
  NAND2_X1 U3197 ( .A1(n3189), .A2(n3190), .ZN(n3284) );
  NAND2_X1 U3198 ( .A1(n3288), .A2(n3289), .ZN(n3190) );
  NAND2_X1 U3199 ( .A1(n2672), .A2(n3290), .ZN(n3289) );
  OR2_X1 U3200 ( .A1(n3160), .A2(n3158), .ZN(n3290) );
  NOR2_X1 U3201 ( .A1(n2328), .A2(n2314), .ZN(n2672) );
  NAND2_X1 U3202 ( .A1(n3158), .A2(n3160), .ZN(n3288) );
  NAND2_X1 U3203 ( .A1(n3291), .A2(n3292), .ZN(n3160) );
  NAND2_X1 U3204 ( .A1(n3293), .A2(b_11_), .ZN(n3292) );
  NOR2_X1 U3205 ( .A1(n3294), .A2(n2285), .ZN(n3293) );
  NOR2_X1 U3206 ( .A1(n3166), .A2(n3168), .ZN(n3294) );
  NAND2_X1 U3207 ( .A1(n3166), .A2(n3168), .ZN(n3291) );
  NAND2_X1 U3208 ( .A1(n3295), .A2(n3296), .ZN(n3168) );
  NAND2_X1 U3209 ( .A1(n3173), .A2(n3297), .ZN(n3296) );
  NAND2_X1 U3210 ( .A1(n3176), .A2(n3175), .ZN(n3297) );
  NOR2_X1 U3211 ( .A1(n2328), .A2(n2271), .ZN(n3173) );
  OR2_X1 U3212 ( .A1(n3175), .A2(n3176), .ZN(n3295) );
  AND2_X1 U3213 ( .A1(n3298), .A2(n3299), .ZN(n3176) );
  NAND2_X1 U3214 ( .A1(b_10_), .A2(n3300), .ZN(n3299) );
  NAND2_X1 U3215 ( .A1(n2843), .A2(n3301), .ZN(n3300) );
  NAND2_X1 U3216 ( .A1(a_14_), .A2(n2688), .ZN(n3301) );
  NAND2_X1 U3217 ( .A1(b_9_), .A2(n3302), .ZN(n3298) );
  NAND2_X1 U3218 ( .A1(n2226), .A2(n3303), .ZN(n3302) );
  NAND2_X1 U3219 ( .A1(a_15_), .A2(n2355), .ZN(n3303) );
  NAND2_X1 U3220 ( .A1(n3304), .A2(n2685), .ZN(n3175) );
  NOR2_X1 U3221 ( .A1(n2328), .A2(n2355), .ZN(n3304) );
  XNOR2_X1 U3222 ( .A(n3305), .B(n3306), .ZN(n3166) );
  XNOR2_X1 U3223 ( .A(n3307), .B(n3308), .ZN(n3306) );
  XOR2_X1 U3224 ( .A(n3309), .B(n3310), .Z(n3158) );
  XNOR2_X1 U3225 ( .A(n3311), .B(n3312), .ZN(n3309) );
  NAND2_X1 U3226 ( .A1(b_10_), .A2(a_12_), .ZN(n3311) );
  XNOR2_X1 U3227 ( .A(n3313), .B(n3314), .ZN(n3189) );
  XNOR2_X1 U3228 ( .A(n3315), .B(n3316), .ZN(n3314) );
  XOR2_X1 U3229 ( .A(n3317), .B(n3318), .Z(n3193) );
  XOR2_X1 U3230 ( .A(n3319), .B(n3320), .Z(n3317) );
  XNOR2_X1 U3231 ( .A(n3321), .B(n3322), .ZN(n3197) );
  XNOR2_X1 U3232 ( .A(n3323), .B(n3324), .ZN(n3322) );
  XNOR2_X1 U3233 ( .A(n3325), .B(n3326), .ZN(n3200) );
  XOR2_X1 U3234 ( .A(n3327), .B(n3328), .Z(n3326) );
  NAND2_X1 U3235 ( .A1(b_10_), .A2(a_8_), .ZN(n3328) );
  XNOR2_X1 U3236 ( .A(n3329), .B(n3330), .ZN(n3205) );
  XNOR2_X1 U3237 ( .A(n3331), .B(n3332), .ZN(n3330) );
  XOR2_X1 U3238 ( .A(n3333), .B(n3334), .Z(n3208) );
  XOR2_X1 U3239 ( .A(n3335), .B(n3336), .Z(n3333) );
  NOR2_X1 U3240 ( .A1(n2691), .A2(n2355), .ZN(n3336) );
  XOR2_X1 U3241 ( .A(n3337), .B(n3338), .Z(n3213) );
  XOR2_X1 U3242 ( .A(n3339), .B(n3340), .Z(n3338) );
  NAND2_X1 U3243 ( .A1(b_10_), .A2(a_5_), .ZN(n3340) );
  XNOR2_X1 U3244 ( .A(n3341), .B(n3342), .ZN(n3216) );
  XNOR2_X1 U3245 ( .A(n3343), .B(n3344), .ZN(n3342) );
  XOR2_X1 U3246 ( .A(n3345), .B(n3346), .Z(n3225) );
  XOR2_X1 U3247 ( .A(n3347), .B(n3348), .Z(n3345) );
  NOR2_X1 U3248 ( .A1(n2695), .A2(n2355), .ZN(n3348) );
  NAND2_X1 U3249 ( .A1(n3349), .A2(n3350), .ZN(n2166) );
  NAND2_X1 U3250 ( .A1(n3236), .A2(n2755), .ZN(n3350) );
  NAND2_X1 U3251 ( .A1(n3351), .A2(n3236), .ZN(n2167) );
  XNOR2_X1 U3252 ( .A(n3352), .B(n3353), .ZN(n3236) );
  XOR2_X1 U3253 ( .A(n3354), .B(n3355), .Z(n3353) );
  NAND2_X1 U3254 ( .A1(b_9_), .A2(a_0_), .ZN(n3355) );
  NOR2_X1 U3255 ( .A1(n3235), .A2(n3349), .ZN(n3351) );
  XOR2_X1 U3256 ( .A(n3356), .B(n3357), .Z(n3349) );
  INV_X1 U3257 ( .A(n3358), .ZN(n3357) );
  INV_X1 U3258 ( .A(n2755), .ZN(n3235) );
  NAND2_X1 U3259 ( .A1(n3239), .A2(n3359), .ZN(n2755) );
  NAND2_X1 U3260 ( .A1(n3238), .A2(n3240), .ZN(n3359) );
  NAND2_X1 U3261 ( .A1(n3360), .A2(n3361), .ZN(n3240) );
  NAND2_X1 U3262 ( .A1(b_10_), .A2(a_0_), .ZN(n3361) );
  INV_X1 U3263 ( .A(n3362), .ZN(n3360) );
  XNOR2_X1 U3264 ( .A(n3363), .B(n3364), .ZN(n3238) );
  XOR2_X1 U3265 ( .A(n3365), .B(n3366), .Z(n3364) );
  NAND2_X1 U3266 ( .A1(b_9_), .A2(a_1_), .ZN(n3366) );
  NAND2_X1 U3267 ( .A1(a_0_), .A2(n3362), .ZN(n3239) );
  NAND2_X1 U3268 ( .A1(n3367), .A2(n3368), .ZN(n3362) );
  NAND2_X1 U3269 ( .A1(n3247), .A2(n3369), .ZN(n3368) );
  NAND2_X1 U3270 ( .A1(n3246), .A2(n3244), .ZN(n3369) );
  NOR2_X1 U3271 ( .A1(n2355), .A2(n2609), .ZN(n3247) );
  OR2_X1 U3272 ( .A1(n3244), .A2(n3246), .ZN(n3367) );
  AND2_X1 U3273 ( .A1(n3370), .A2(n3371), .ZN(n3246) );
  NAND2_X1 U3274 ( .A1(n3372), .A2(b_10_), .ZN(n3371) );
  NOR2_X1 U3275 ( .A1(n3373), .A2(n2695), .ZN(n3372) );
  NOR2_X1 U3276 ( .A1(n3346), .A2(n3347), .ZN(n3373) );
  NAND2_X1 U3277 ( .A1(n3346), .A2(n3347), .ZN(n3370) );
  NAND2_X1 U3278 ( .A1(n3374), .A2(n3375), .ZN(n3347) );
  NAND2_X1 U3279 ( .A1(n3259), .A2(n3376), .ZN(n3375) );
  OR2_X1 U3280 ( .A1(n3257), .A2(n3258), .ZN(n3376) );
  NOR2_X1 U3281 ( .A1(n2355), .A2(n2553), .ZN(n3259) );
  NAND2_X1 U3282 ( .A1(n3257), .A2(n3258), .ZN(n3374) );
  NAND2_X1 U3283 ( .A1(n3377), .A2(n3378), .ZN(n3258) );
  NAND2_X1 U3284 ( .A1(n3344), .A2(n3379), .ZN(n3378) );
  OR2_X1 U3285 ( .A1(n3341), .A2(n3343), .ZN(n3379) );
  NOR2_X1 U3286 ( .A1(n2355), .A2(n2506), .ZN(n3344) );
  NAND2_X1 U3287 ( .A1(n3341), .A2(n3343), .ZN(n3377) );
  NAND2_X1 U3288 ( .A1(n3380), .A2(n3381), .ZN(n3343) );
  NAND2_X1 U3289 ( .A1(n3382), .A2(b_10_), .ZN(n3381) );
  NOR2_X1 U3290 ( .A1(n3383), .A2(n2479), .ZN(n3382) );
  NOR2_X1 U3291 ( .A1(n3339), .A2(n3337), .ZN(n3383) );
  NAND2_X1 U3292 ( .A1(n3337), .A2(n3339), .ZN(n3380) );
  NAND2_X1 U3293 ( .A1(n3384), .A2(n3385), .ZN(n3339) );
  NAND2_X1 U3294 ( .A1(n3386), .A2(b_10_), .ZN(n3385) );
  NOR2_X1 U3295 ( .A1(n3387), .A2(n2691), .ZN(n3386) );
  NOR2_X1 U3296 ( .A1(n3335), .A2(n3334), .ZN(n3387) );
  NAND2_X1 U3297 ( .A1(n3334), .A2(n3335), .ZN(n3384) );
  NAND2_X1 U3298 ( .A1(n3388), .A2(n3389), .ZN(n3335) );
  NAND2_X1 U3299 ( .A1(n3332), .A2(n3390), .ZN(n3389) );
  OR2_X1 U3300 ( .A1(n3329), .A2(n3331), .ZN(n3390) );
  NOR2_X1 U3301 ( .A1(n2355), .A2(n2437), .ZN(n3332) );
  NAND2_X1 U3302 ( .A1(n3329), .A2(n3331), .ZN(n3388) );
  NAND2_X1 U3303 ( .A1(n3391), .A2(n3392), .ZN(n3331) );
  NAND2_X1 U3304 ( .A1(n3393), .A2(b_10_), .ZN(n3392) );
  NOR2_X1 U3305 ( .A1(n3394), .A2(n2689), .ZN(n3393) );
  NOR2_X1 U3306 ( .A1(n3325), .A2(n3327), .ZN(n3394) );
  NAND2_X1 U3307 ( .A1(n3325), .A2(n3327), .ZN(n3391) );
  NAND2_X1 U3308 ( .A1(n3395), .A2(n3396), .ZN(n3327) );
  NAND2_X1 U3309 ( .A1(n3324), .A2(n3397), .ZN(n3396) );
  OR2_X1 U3310 ( .A1(n3321), .A2(n3323), .ZN(n3397) );
  NOR2_X1 U3311 ( .A1(n2355), .A2(n2383), .ZN(n3324) );
  NAND2_X1 U3312 ( .A1(n3321), .A2(n3323), .ZN(n3395) );
  NAND2_X1 U3313 ( .A1(n3398), .A2(n3399), .ZN(n3323) );
  NAND2_X1 U3314 ( .A1(n3318), .A2(n3400), .ZN(n3399) );
  OR2_X1 U3315 ( .A1(n3319), .A2(n3320), .ZN(n3400) );
  XNOR2_X1 U3316 ( .A(n3401), .B(n3402), .ZN(n3318) );
  XNOR2_X1 U3317 ( .A(n3403), .B(n3404), .ZN(n3402) );
  NAND2_X1 U3318 ( .A1(n3320), .A2(n3319), .ZN(n3398) );
  NAND2_X1 U3319 ( .A1(n3405), .A2(n3406), .ZN(n3319) );
  NAND2_X1 U3320 ( .A1(n3316), .A2(n3407), .ZN(n3406) );
  OR2_X1 U3321 ( .A1(n3313), .A2(n3315), .ZN(n3407) );
  NOR2_X1 U3322 ( .A1(n2355), .A2(n2314), .ZN(n3316) );
  NAND2_X1 U3323 ( .A1(n3313), .A2(n3315), .ZN(n3405) );
  NAND2_X1 U3324 ( .A1(n3408), .A2(n3409), .ZN(n3315) );
  NAND2_X1 U3325 ( .A1(n3410), .A2(b_10_), .ZN(n3409) );
  NOR2_X1 U3326 ( .A1(n3411), .A2(n2285), .ZN(n3410) );
  NOR2_X1 U3327 ( .A1(n3310), .A2(n3312), .ZN(n3411) );
  NAND2_X1 U3328 ( .A1(n3310), .A2(n3312), .ZN(n3408) );
  NAND2_X1 U3329 ( .A1(n3412), .A2(n3413), .ZN(n3312) );
  NAND2_X1 U3330 ( .A1(n3305), .A2(n3414), .ZN(n3413) );
  NAND2_X1 U3331 ( .A1(n3308), .A2(n3307), .ZN(n3414) );
  NOR2_X1 U3332 ( .A1(n2355), .A2(n2271), .ZN(n3305) );
  OR2_X1 U3333 ( .A1(n3307), .A2(n3308), .ZN(n3412) );
  AND2_X1 U3334 ( .A1(n3415), .A2(n3416), .ZN(n3308) );
  NAND2_X1 U3335 ( .A1(b_8_), .A2(n3417), .ZN(n3416) );
  NAND2_X1 U3336 ( .A1(n2226), .A2(n3418), .ZN(n3417) );
  NAND2_X1 U3337 ( .A1(a_15_), .A2(n2688), .ZN(n3418) );
  NAND2_X1 U3338 ( .A1(b_9_), .A2(n3419), .ZN(n3415) );
  NAND2_X1 U3339 ( .A1(n2843), .A2(n3420), .ZN(n3419) );
  NAND2_X1 U3340 ( .A1(a_14_), .A2(n2410), .ZN(n3420) );
  NAND2_X1 U3341 ( .A1(n3421), .A2(n2685), .ZN(n3307) );
  NOR2_X1 U3342 ( .A1(n2355), .A2(n2688), .ZN(n3421) );
  XNOR2_X1 U3343 ( .A(n3422), .B(n3423), .ZN(n3310) );
  XNOR2_X1 U3344 ( .A(n3424), .B(n3425), .ZN(n3423) );
  XOR2_X1 U3345 ( .A(n3426), .B(n3427), .Z(n3313) );
  XNOR2_X1 U3346 ( .A(n3428), .B(n3429), .ZN(n3426) );
  NAND2_X1 U3347 ( .A1(b_9_), .A2(a_12_), .ZN(n3428) );
  INV_X1 U3348 ( .A(n2669), .ZN(n3320) );
  NAND2_X1 U3349 ( .A1(b_10_), .A2(a_10_), .ZN(n2669) );
  XOR2_X1 U3350 ( .A(n3430), .B(n3431), .Z(n3321) );
  XOR2_X1 U3351 ( .A(n3432), .B(n3433), .Z(n3430) );
  NOR2_X1 U3352 ( .A1(n2687), .A2(n2688), .ZN(n3433) );
  XOR2_X1 U3353 ( .A(n3434), .B(n3435), .Z(n3325) );
  XOR2_X1 U3354 ( .A(n3436), .B(n3437), .Z(n3434) );
  XOR2_X1 U3355 ( .A(n3438), .B(n3439), .Z(n3329) );
  XOR2_X1 U3356 ( .A(n3440), .B(n3441), .Z(n3438) );
  NOR2_X1 U3357 ( .A1(n2689), .A2(n2688), .ZN(n3441) );
  XNOR2_X1 U3358 ( .A(n3442), .B(n3443), .ZN(n3334) );
  XNOR2_X1 U3359 ( .A(n3444), .B(n3445), .ZN(n3443) );
  XNOR2_X1 U3360 ( .A(n3446), .B(n3447), .ZN(n3337) );
  XNOR2_X1 U3361 ( .A(n3448), .B(n3449), .ZN(n3446) );
  XOR2_X1 U3362 ( .A(n3450), .B(n3451), .Z(n3341) );
  XOR2_X1 U3363 ( .A(n3452), .B(n3453), .Z(n3450) );
  NOR2_X1 U3364 ( .A1(n2479), .A2(n2688), .ZN(n3453) );
  XNOR2_X1 U3365 ( .A(n3454), .B(n3455), .ZN(n3257) );
  XOR2_X1 U3366 ( .A(n3456), .B(n3457), .Z(n3455) );
  NAND2_X1 U3367 ( .A1(b_9_), .A2(a_4_), .ZN(n3457) );
  XNOR2_X1 U3368 ( .A(n3458), .B(n3459), .ZN(n3346) );
  XOR2_X1 U3369 ( .A(n3460), .B(n3461), .Z(n3459) );
  NAND2_X1 U3370 ( .A1(b_9_), .A2(a_3_), .ZN(n3461) );
  XOR2_X1 U3371 ( .A(n3462), .B(n3463), .Z(n3244) );
  XOR2_X1 U3372 ( .A(n3464), .B(n3465), .Z(n3463) );
  NAND2_X1 U3373 ( .A1(b_9_), .A2(a_2_), .ZN(n3465) );
  NAND2_X1 U3374 ( .A1(n3466), .A2(n3467), .ZN(n2172) );
  NAND2_X1 U3375 ( .A1(n3358), .A2(n3356), .ZN(n3467) );
  NAND2_X1 U3376 ( .A1(n3468), .A2(n3358), .ZN(n2173) );
  XOR2_X1 U3377 ( .A(n3469), .B(n3470), .Z(n3358) );
  XOR2_X1 U3378 ( .A(n3471), .B(n3472), .Z(n3469) );
  NOR2_X1 U3379 ( .A1(n3473), .A2(n3466), .ZN(n3468) );
  XOR2_X1 U3380 ( .A(n3474), .B(n3475), .Z(n3466) );
  INV_X1 U3381 ( .A(n3476), .ZN(n3475) );
  INV_X1 U3382 ( .A(n3356), .ZN(n3473) );
  NAND2_X1 U3383 ( .A1(n3477), .A2(n3478), .ZN(n3356) );
  NAND2_X1 U3384 ( .A1(n3479), .A2(b_9_), .ZN(n3478) );
  NOR2_X1 U3385 ( .A1(n3480), .A2(n2623), .ZN(n3479) );
  NOR2_X1 U3386 ( .A1(n3354), .A2(n3352), .ZN(n3480) );
  NAND2_X1 U3387 ( .A1(n3352), .A2(n3354), .ZN(n3477) );
  NAND2_X1 U3388 ( .A1(n3481), .A2(n3482), .ZN(n3354) );
  NAND2_X1 U3389 ( .A1(n3483), .A2(b_9_), .ZN(n3482) );
  NOR2_X1 U3390 ( .A1(n3484), .A2(n2609), .ZN(n3483) );
  NOR2_X1 U3391 ( .A1(n3363), .A2(n3365), .ZN(n3484) );
  NAND2_X1 U3392 ( .A1(n3363), .A2(n3365), .ZN(n3481) );
  NAND2_X1 U3393 ( .A1(n3485), .A2(n3486), .ZN(n3365) );
  NAND2_X1 U3394 ( .A1(n3487), .A2(b_9_), .ZN(n3486) );
  NOR2_X1 U3395 ( .A1(n3488), .A2(n2695), .ZN(n3487) );
  NOR2_X1 U3396 ( .A1(n3464), .A2(n3462), .ZN(n3488) );
  NAND2_X1 U3397 ( .A1(n3462), .A2(n3464), .ZN(n3485) );
  NAND2_X1 U3398 ( .A1(n3489), .A2(n3490), .ZN(n3464) );
  NAND2_X1 U3399 ( .A1(n3491), .A2(b_9_), .ZN(n3490) );
  NOR2_X1 U3400 ( .A1(n3492), .A2(n2553), .ZN(n3491) );
  NOR2_X1 U3401 ( .A1(n3460), .A2(n3458), .ZN(n3492) );
  NAND2_X1 U3402 ( .A1(n3458), .A2(n3460), .ZN(n3489) );
  NAND2_X1 U3403 ( .A1(n3493), .A2(n3494), .ZN(n3460) );
  NAND2_X1 U3404 ( .A1(n3495), .A2(b_9_), .ZN(n3494) );
  NOR2_X1 U3405 ( .A1(n3496), .A2(n2506), .ZN(n3495) );
  NOR2_X1 U3406 ( .A1(n3454), .A2(n3456), .ZN(n3496) );
  NAND2_X1 U3407 ( .A1(n3454), .A2(n3456), .ZN(n3493) );
  NAND2_X1 U3408 ( .A1(n3497), .A2(n3498), .ZN(n3456) );
  NAND2_X1 U3409 ( .A1(n3499), .A2(b_9_), .ZN(n3498) );
  NOR2_X1 U3410 ( .A1(n3500), .A2(n2479), .ZN(n3499) );
  NOR2_X1 U3411 ( .A1(n3451), .A2(n3452), .ZN(n3500) );
  NAND2_X1 U3412 ( .A1(n3451), .A2(n3452), .ZN(n3497) );
  NAND2_X1 U3413 ( .A1(n3501), .A2(n3502), .ZN(n3452) );
  NAND2_X1 U3414 ( .A1(n3449), .A2(n3503), .ZN(n3502) );
  NAND2_X1 U3415 ( .A1(n3448), .A2(n3447), .ZN(n3503) );
  NOR2_X1 U3416 ( .A1(n2688), .A2(n2691), .ZN(n3449) );
  OR2_X1 U3417 ( .A1(n3447), .A2(n3448), .ZN(n3501) );
  AND2_X1 U3418 ( .A1(n3504), .A2(n3505), .ZN(n3448) );
  NAND2_X1 U3419 ( .A1(n3445), .A2(n3506), .ZN(n3505) );
  OR2_X1 U3420 ( .A1(n3444), .A2(n3442), .ZN(n3506) );
  NOR2_X1 U3421 ( .A1(n2688), .A2(n2437), .ZN(n3445) );
  NAND2_X1 U3422 ( .A1(n3442), .A2(n3444), .ZN(n3504) );
  NAND2_X1 U3423 ( .A1(n3507), .A2(n3508), .ZN(n3444) );
  NAND2_X1 U3424 ( .A1(n3509), .A2(b_9_), .ZN(n3508) );
  NOR2_X1 U3425 ( .A1(n3510), .A2(n2689), .ZN(n3509) );
  NOR2_X1 U3426 ( .A1(n3439), .A2(n3440), .ZN(n3510) );
  NAND2_X1 U3427 ( .A1(n3439), .A2(n3440), .ZN(n3507) );
  NAND2_X1 U3428 ( .A1(n3511), .A2(n3512), .ZN(n3440) );
  NAND2_X1 U3429 ( .A1(n3437), .A2(n3513), .ZN(n3512) );
  OR2_X1 U3430 ( .A1(n3435), .A2(n3436), .ZN(n3513) );
  INV_X1 U3431 ( .A(n2666), .ZN(n3437) );
  NAND2_X1 U3432 ( .A1(b_9_), .A2(a_9_), .ZN(n2666) );
  NAND2_X1 U3433 ( .A1(n3435), .A2(n3436), .ZN(n3511) );
  NAND2_X1 U3434 ( .A1(n3514), .A2(n3515), .ZN(n3436) );
  NAND2_X1 U3435 ( .A1(n3516), .A2(b_9_), .ZN(n3515) );
  NOR2_X1 U3436 ( .A1(n3517), .A2(n2687), .ZN(n3516) );
  NOR2_X1 U3437 ( .A1(n3431), .A2(n3432), .ZN(n3517) );
  NAND2_X1 U3438 ( .A1(n3431), .A2(n3432), .ZN(n3514) );
  NAND2_X1 U3439 ( .A1(n3518), .A2(n3519), .ZN(n3432) );
  NAND2_X1 U3440 ( .A1(n3404), .A2(n3520), .ZN(n3519) );
  OR2_X1 U3441 ( .A1(n3401), .A2(n3403), .ZN(n3520) );
  NOR2_X1 U3442 ( .A1(n2688), .A2(n2314), .ZN(n3404) );
  NAND2_X1 U3443 ( .A1(n3401), .A2(n3403), .ZN(n3518) );
  NAND2_X1 U3444 ( .A1(n3521), .A2(n3522), .ZN(n3403) );
  NAND2_X1 U3445 ( .A1(n3523), .A2(b_9_), .ZN(n3522) );
  NOR2_X1 U3446 ( .A1(n3524), .A2(n2285), .ZN(n3523) );
  NOR2_X1 U3447 ( .A1(n3427), .A2(n3429), .ZN(n3524) );
  NAND2_X1 U3448 ( .A1(n3427), .A2(n3429), .ZN(n3521) );
  NAND2_X1 U3449 ( .A1(n3525), .A2(n3526), .ZN(n3429) );
  NAND2_X1 U3450 ( .A1(n3422), .A2(n3527), .ZN(n3526) );
  NAND2_X1 U3451 ( .A1(n3425), .A2(n3424), .ZN(n3527) );
  NOR2_X1 U3452 ( .A1(n2688), .A2(n2271), .ZN(n3422) );
  OR2_X1 U3453 ( .A1(n3424), .A2(n3425), .ZN(n3525) );
  AND2_X1 U3454 ( .A1(n3528), .A2(n3529), .ZN(n3425) );
  NAND2_X1 U3455 ( .A1(b_7_), .A2(n3530), .ZN(n3529) );
  NAND2_X1 U3456 ( .A1(n2226), .A2(n3531), .ZN(n3530) );
  NAND2_X1 U3457 ( .A1(a_15_), .A2(n2410), .ZN(n3531) );
  NAND2_X1 U3458 ( .A1(b_8_), .A2(n3532), .ZN(n3528) );
  NAND2_X1 U3459 ( .A1(n2843), .A2(n3533), .ZN(n3532) );
  NAND2_X1 U3460 ( .A1(a_14_), .A2(n2690), .ZN(n3533) );
  NAND2_X1 U3461 ( .A1(n3534), .A2(n2685), .ZN(n3424) );
  NOR2_X1 U3462 ( .A1(n2688), .A2(n2410), .ZN(n3534) );
  XNOR2_X1 U3463 ( .A(n3535), .B(n3536), .ZN(n3427) );
  XNOR2_X1 U3464 ( .A(n3537), .B(n3538), .ZN(n3536) );
  XOR2_X1 U3465 ( .A(n3539), .B(n3540), .Z(n3401) );
  XNOR2_X1 U3466 ( .A(n3541), .B(n3542), .ZN(n3539) );
  NAND2_X1 U3467 ( .A1(b_8_), .A2(a_12_), .ZN(n3541) );
  XNOR2_X1 U3468 ( .A(n3543), .B(n3544), .ZN(n3431) );
  XNOR2_X1 U3469 ( .A(n3545), .B(n3546), .ZN(n3544) );
  XOR2_X1 U3470 ( .A(n3547), .B(n3548), .Z(n3435) );
  XOR2_X1 U3471 ( .A(n3549), .B(n3550), .Z(n3547) );
  NOR2_X1 U3472 ( .A1(n2687), .A2(n2410), .ZN(n3550) );
  XOR2_X1 U3473 ( .A(n3551), .B(n3552), .Z(n3439) );
  XOR2_X1 U3474 ( .A(n3553), .B(n3554), .Z(n3551) );
  XOR2_X1 U3475 ( .A(n3555), .B(n3556), .Z(n3442) );
  XOR2_X1 U3476 ( .A(n3557), .B(n3558), .Z(n3555) );
  XOR2_X1 U3477 ( .A(n3559), .B(n3560), .Z(n3447) );
  XOR2_X1 U3478 ( .A(n3561), .B(n3562), .Z(n3560) );
  NAND2_X1 U3479 ( .A1(b_8_), .A2(a_7_), .ZN(n3562) );
  XOR2_X1 U3480 ( .A(n3563), .B(n3564), .Z(n3451) );
  XNOR2_X1 U3481 ( .A(n3565), .B(n3566), .ZN(n3563) );
  NAND2_X1 U3482 ( .A1(b_8_), .A2(a_6_), .ZN(n3565) );
  XNOR2_X1 U3483 ( .A(n3567), .B(n3568), .ZN(n3454) );
  XOR2_X1 U3484 ( .A(n3569), .B(n3570), .Z(n3568) );
  NAND2_X1 U3485 ( .A1(b_8_), .A2(a_5_), .ZN(n3570) );
  XNOR2_X1 U3486 ( .A(n3571), .B(n3572), .ZN(n3458) );
  XOR2_X1 U3487 ( .A(n3573), .B(n3574), .Z(n3572) );
  NAND2_X1 U3488 ( .A1(b_8_), .A2(a_4_), .ZN(n3574) );
  XOR2_X1 U3489 ( .A(n3575), .B(n3576), .Z(n3462) );
  XOR2_X1 U3490 ( .A(n3577), .B(n3578), .Z(n3576) );
  XOR2_X1 U3491 ( .A(n3579), .B(n3580), .Z(n3363) );
  XOR2_X1 U3492 ( .A(n3581), .B(n3582), .Z(n3579) );
  XNOR2_X1 U3493 ( .A(n3583), .B(n3584), .ZN(n3352) );
  NAND2_X1 U3494 ( .A1(n3585), .A2(n3586), .ZN(n3583) );
  NAND2_X1 U3495 ( .A1(n3587), .A2(n3588), .ZN(n2178) );
  NAND2_X1 U3496 ( .A1(n3476), .A2(n3474), .ZN(n3588) );
  NAND2_X1 U3497 ( .A1(n3589), .A2(n3476), .ZN(n2179) );
  XNOR2_X1 U3498 ( .A(n3590), .B(n3591), .ZN(n3476) );
  XOR2_X1 U3499 ( .A(n3592), .B(n3593), .Z(n3591) );
  NAND2_X1 U3500 ( .A1(b_7_), .A2(a_0_), .ZN(n3593) );
  NOR2_X1 U3501 ( .A1(n3594), .A2(n3587), .ZN(n3589) );
  XOR2_X1 U3502 ( .A(n3595), .B(n3596), .Z(n3587) );
  INV_X1 U3503 ( .A(n3597), .ZN(n3596) );
  INV_X1 U3504 ( .A(n3474), .ZN(n3594) );
  NAND2_X1 U3505 ( .A1(n3598), .A2(n3599), .ZN(n3474) );
  NAND2_X1 U3506 ( .A1(n3472), .A2(n3600), .ZN(n3599) );
  OR2_X1 U3507 ( .A1(n3470), .A2(n3471), .ZN(n3600) );
  NOR2_X1 U3508 ( .A1(n2410), .A2(n2623), .ZN(n3472) );
  NAND2_X1 U3509 ( .A1(n3470), .A2(n3471), .ZN(n3598) );
  NAND2_X1 U3510 ( .A1(n3585), .A2(n3601), .ZN(n3471) );
  NAND2_X1 U3511 ( .A1(n3584), .A2(n3586), .ZN(n3601) );
  NAND2_X1 U3512 ( .A1(n3602), .A2(n3603), .ZN(n3586) );
  NAND2_X1 U3513 ( .A1(b_8_), .A2(a_1_), .ZN(n3603) );
  INV_X1 U3514 ( .A(n3604), .ZN(n3602) );
  XNOR2_X1 U3515 ( .A(n3605), .B(n3606), .ZN(n3584) );
  XOR2_X1 U3516 ( .A(n3607), .B(n3608), .Z(n3606) );
  NAND2_X1 U3517 ( .A1(b_7_), .A2(a_2_), .ZN(n3608) );
  NAND2_X1 U3518 ( .A1(a_1_), .A2(n3604), .ZN(n3585) );
  NAND2_X1 U3519 ( .A1(n3609), .A2(n3610), .ZN(n3604) );
  NAND2_X1 U3520 ( .A1(n3582), .A2(n3611), .ZN(n3610) );
  OR2_X1 U3521 ( .A1(n3580), .A2(n3581), .ZN(n3611) );
  NOR2_X1 U3522 ( .A1(n2410), .A2(n2695), .ZN(n3582) );
  NAND2_X1 U3523 ( .A1(n3580), .A2(n3581), .ZN(n3609) );
  NAND2_X1 U3524 ( .A1(n3612), .A2(n3613), .ZN(n3581) );
  NAND2_X1 U3525 ( .A1(n3578), .A2(n3614), .ZN(n3613) );
  NAND2_X1 U3526 ( .A1(n3577), .A2(n3575), .ZN(n3614) );
  NOR2_X1 U3527 ( .A1(n2410), .A2(n2553), .ZN(n3578) );
  OR2_X1 U3528 ( .A1(n3575), .A2(n3577), .ZN(n3612) );
  AND2_X1 U3529 ( .A1(n3615), .A2(n3616), .ZN(n3577) );
  NAND2_X1 U3530 ( .A1(n3617), .A2(b_8_), .ZN(n3616) );
  NOR2_X1 U3531 ( .A1(n3618), .A2(n2506), .ZN(n3617) );
  NOR2_X1 U3532 ( .A1(n3571), .A2(n3573), .ZN(n3618) );
  NAND2_X1 U3533 ( .A1(n3571), .A2(n3573), .ZN(n3615) );
  NAND2_X1 U3534 ( .A1(n3619), .A2(n3620), .ZN(n3573) );
  NAND2_X1 U3535 ( .A1(n3621), .A2(b_8_), .ZN(n3620) );
  NOR2_X1 U3536 ( .A1(n3622), .A2(n2479), .ZN(n3621) );
  NOR2_X1 U3537 ( .A1(n3569), .A2(n3567), .ZN(n3622) );
  NAND2_X1 U3538 ( .A1(n3567), .A2(n3569), .ZN(n3619) );
  NAND2_X1 U3539 ( .A1(n3623), .A2(n3624), .ZN(n3569) );
  NAND2_X1 U3540 ( .A1(n3625), .A2(b_8_), .ZN(n3624) );
  NOR2_X1 U3541 ( .A1(n3626), .A2(n2691), .ZN(n3625) );
  NOR2_X1 U3542 ( .A1(n3566), .A2(n3564), .ZN(n3626) );
  NAND2_X1 U3543 ( .A1(n3564), .A2(n3566), .ZN(n3623) );
  NAND2_X1 U3544 ( .A1(n3627), .A2(n3628), .ZN(n3566) );
  NAND2_X1 U3545 ( .A1(n3629), .A2(b_8_), .ZN(n3628) );
  NOR2_X1 U3546 ( .A1(n3630), .A2(n2437), .ZN(n3629) );
  NOR2_X1 U3547 ( .A1(n3561), .A2(n3559), .ZN(n3630) );
  NAND2_X1 U3548 ( .A1(n3559), .A2(n3561), .ZN(n3627) );
  NAND2_X1 U3549 ( .A1(n3631), .A2(n3632), .ZN(n3561) );
  NAND2_X1 U3550 ( .A1(n3556), .A2(n3633), .ZN(n3632) );
  OR2_X1 U3551 ( .A1(n3557), .A2(n3558), .ZN(n3633) );
  XNOR2_X1 U3552 ( .A(n3634), .B(n3635), .ZN(n3556) );
  XNOR2_X1 U3553 ( .A(n3636), .B(n3637), .ZN(n3634) );
  NAND2_X1 U3554 ( .A1(n3558), .A2(n3557), .ZN(n3631) );
  NAND2_X1 U3555 ( .A1(n3638), .A2(n3639), .ZN(n3557) );
  NAND2_X1 U3556 ( .A1(n3554), .A2(n3640), .ZN(n3639) );
  OR2_X1 U3557 ( .A1(n3552), .A2(n3553), .ZN(n3640) );
  NOR2_X1 U3558 ( .A1(n2410), .A2(n2383), .ZN(n3554) );
  NAND2_X1 U3559 ( .A1(n3552), .A2(n3553), .ZN(n3638) );
  NAND2_X1 U3560 ( .A1(n3641), .A2(n3642), .ZN(n3553) );
  NAND2_X1 U3561 ( .A1(n3643), .A2(b_8_), .ZN(n3642) );
  NOR2_X1 U3562 ( .A1(n3644), .A2(n2687), .ZN(n3643) );
  NOR2_X1 U3563 ( .A1(n3548), .A2(n3549), .ZN(n3644) );
  NAND2_X1 U3564 ( .A1(n3548), .A2(n3549), .ZN(n3641) );
  NAND2_X1 U3565 ( .A1(n3645), .A2(n3646), .ZN(n3549) );
  NAND2_X1 U3566 ( .A1(n3546), .A2(n3647), .ZN(n3646) );
  OR2_X1 U3567 ( .A1(n3543), .A2(n3545), .ZN(n3647) );
  NOR2_X1 U3568 ( .A1(n2410), .A2(n2314), .ZN(n3546) );
  NAND2_X1 U3569 ( .A1(n3543), .A2(n3545), .ZN(n3645) );
  NAND2_X1 U3570 ( .A1(n3648), .A2(n3649), .ZN(n3545) );
  NAND2_X1 U3571 ( .A1(n3650), .A2(b_8_), .ZN(n3649) );
  NOR2_X1 U3572 ( .A1(n3651), .A2(n2285), .ZN(n3650) );
  NOR2_X1 U3573 ( .A1(n3540), .A2(n3542), .ZN(n3651) );
  NAND2_X1 U3574 ( .A1(n3540), .A2(n3542), .ZN(n3648) );
  NAND2_X1 U3575 ( .A1(n3652), .A2(n3653), .ZN(n3542) );
  NAND2_X1 U3576 ( .A1(n3535), .A2(n3654), .ZN(n3653) );
  NAND2_X1 U3577 ( .A1(n3538), .A2(n3537), .ZN(n3654) );
  NOR2_X1 U3578 ( .A1(n2410), .A2(n2271), .ZN(n3535) );
  OR2_X1 U3579 ( .A1(n3537), .A2(n3538), .ZN(n3652) );
  AND2_X1 U3580 ( .A1(n3655), .A2(n3656), .ZN(n3538) );
  NAND2_X1 U3581 ( .A1(b_6_), .A2(n3657), .ZN(n3656) );
  NAND2_X1 U3582 ( .A1(n2226), .A2(n3658), .ZN(n3657) );
  NAND2_X1 U3583 ( .A1(a_15_), .A2(n2690), .ZN(n3658) );
  NAND2_X1 U3584 ( .A1(b_7_), .A2(n3659), .ZN(n3655) );
  NAND2_X1 U3585 ( .A1(n2843), .A2(n3660), .ZN(n3659) );
  NAND2_X1 U3586 ( .A1(a_14_), .A2(n2464), .ZN(n3660) );
  NAND2_X1 U3587 ( .A1(n3661), .A2(n2685), .ZN(n3537) );
  NOR2_X1 U3588 ( .A1(n2410), .A2(n2690), .ZN(n3661) );
  XNOR2_X1 U3589 ( .A(n3662), .B(n3663), .ZN(n3540) );
  XNOR2_X1 U3590 ( .A(n3664), .B(n3665), .ZN(n3663) );
  XOR2_X1 U3591 ( .A(n3666), .B(n3667), .Z(n3543) );
  XNOR2_X1 U3592 ( .A(n3668), .B(n3669), .ZN(n3666) );
  NAND2_X1 U3593 ( .A1(b_7_), .A2(a_12_), .ZN(n3668) );
  XNOR2_X1 U3594 ( .A(n3670), .B(n3671), .ZN(n3548) );
  XNOR2_X1 U3595 ( .A(n3672), .B(n3673), .ZN(n3671) );
  XOR2_X1 U3596 ( .A(n3674), .B(n3675), .Z(n3552) );
  XOR2_X1 U3597 ( .A(n3676), .B(n3677), .Z(n3674) );
  NOR2_X1 U3598 ( .A1(n2687), .A2(n2690), .ZN(n3677) );
  INV_X1 U3599 ( .A(n2663), .ZN(n3558) );
  NAND2_X1 U3600 ( .A1(b_8_), .A2(a_8_), .ZN(n2663) );
  XOR2_X1 U3601 ( .A(n3678), .B(n3679), .Z(n3559) );
  XOR2_X1 U3602 ( .A(n3680), .B(n3681), .Z(n3678) );
  NOR2_X1 U3603 ( .A1(n2689), .A2(n2690), .ZN(n3681) );
  XNOR2_X1 U3604 ( .A(n3682), .B(n3683), .ZN(n3564) );
  XNOR2_X1 U3605 ( .A(n2660), .B(n3684), .ZN(n3683) );
  XNOR2_X1 U3606 ( .A(n3685), .B(n3686), .ZN(n3567) );
  NAND2_X1 U3607 ( .A1(n3687), .A2(n3688), .ZN(n3685) );
  XNOR2_X1 U3608 ( .A(n3689), .B(n3690), .ZN(n3571) );
  XOR2_X1 U3609 ( .A(n3691), .B(n3692), .Z(n3690) );
  NAND2_X1 U3610 ( .A1(b_7_), .A2(a_5_), .ZN(n3692) );
  XOR2_X1 U3611 ( .A(n3693), .B(n3694), .Z(n3575) );
  XOR2_X1 U3612 ( .A(n3695), .B(n3696), .Z(n3694) );
  NAND2_X1 U3613 ( .A1(b_7_), .A2(a_4_), .ZN(n3696) );
  XNOR2_X1 U3614 ( .A(n3697), .B(n3698), .ZN(n3580) );
  XOR2_X1 U3615 ( .A(n3699), .B(n3700), .Z(n3698) );
  NAND2_X1 U3616 ( .A1(b_7_), .A2(a_3_), .ZN(n3700) );
  XNOR2_X1 U3617 ( .A(n3701), .B(n3702), .ZN(n3470) );
  XOR2_X1 U3618 ( .A(n3703), .B(n3704), .Z(n3702) );
  NAND2_X1 U3619 ( .A1(b_7_), .A2(a_1_), .ZN(n3704) );
  NAND2_X1 U3620 ( .A1(n3705), .A2(n3706), .ZN(n2184) );
  NAND2_X1 U3621 ( .A1(n3597), .A2(n3595), .ZN(n3706) );
  NAND2_X1 U3622 ( .A1(n3707), .A2(n3597), .ZN(n2185) );
  XNOR2_X1 U3623 ( .A(n3708), .B(n3709), .ZN(n3597) );
  XOR2_X1 U3624 ( .A(n3710), .B(n3711), .Z(n3709) );
  NAND2_X1 U3625 ( .A1(b_6_), .A2(a_0_), .ZN(n3711) );
  NOR2_X1 U3626 ( .A1(n3712), .A2(n3705), .ZN(n3707) );
  XNOR2_X1 U3627 ( .A(n3713), .B(n3714), .ZN(n3705) );
  INV_X1 U3628 ( .A(n3595), .ZN(n3712) );
  NAND2_X1 U3629 ( .A1(n3715), .A2(n3716), .ZN(n3595) );
  NAND2_X1 U3630 ( .A1(n3717), .A2(b_7_), .ZN(n3716) );
  NOR2_X1 U3631 ( .A1(n3718), .A2(n2623), .ZN(n3717) );
  NOR2_X1 U3632 ( .A1(n3592), .A2(n3590), .ZN(n3718) );
  NAND2_X1 U3633 ( .A1(n3590), .A2(n3592), .ZN(n3715) );
  NAND2_X1 U3634 ( .A1(n3719), .A2(n3720), .ZN(n3592) );
  NAND2_X1 U3635 ( .A1(n3721), .A2(b_7_), .ZN(n3720) );
  NOR2_X1 U3636 ( .A1(n3722), .A2(n2609), .ZN(n3721) );
  NOR2_X1 U3637 ( .A1(n3701), .A2(n3703), .ZN(n3722) );
  NAND2_X1 U3638 ( .A1(n3701), .A2(n3703), .ZN(n3719) );
  NAND2_X1 U3639 ( .A1(n3723), .A2(n3724), .ZN(n3703) );
  NAND2_X1 U3640 ( .A1(n3725), .A2(b_7_), .ZN(n3724) );
  NOR2_X1 U3641 ( .A1(n3726), .A2(n2695), .ZN(n3725) );
  NOR2_X1 U3642 ( .A1(n3605), .A2(n3607), .ZN(n3726) );
  NAND2_X1 U3643 ( .A1(n3605), .A2(n3607), .ZN(n3723) );
  NAND2_X1 U3644 ( .A1(n3727), .A2(n3728), .ZN(n3607) );
  NAND2_X1 U3645 ( .A1(n3729), .A2(b_7_), .ZN(n3728) );
  NOR2_X1 U3646 ( .A1(n3730), .A2(n2553), .ZN(n3729) );
  NOR2_X1 U3647 ( .A1(n3697), .A2(n3699), .ZN(n3730) );
  NAND2_X1 U3648 ( .A1(n3697), .A2(n3699), .ZN(n3727) );
  NAND2_X1 U3649 ( .A1(n3731), .A2(n3732), .ZN(n3699) );
  NAND2_X1 U3650 ( .A1(n3733), .A2(b_7_), .ZN(n3732) );
  NOR2_X1 U3651 ( .A1(n3734), .A2(n2506), .ZN(n3733) );
  NOR2_X1 U3652 ( .A1(n3695), .A2(n3693), .ZN(n3734) );
  NAND2_X1 U3653 ( .A1(n3693), .A2(n3695), .ZN(n3731) );
  NAND2_X1 U3654 ( .A1(n3735), .A2(n3736), .ZN(n3695) );
  NAND2_X1 U3655 ( .A1(n3737), .A2(b_7_), .ZN(n3736) );
  NOR2_X1 U3656 ( .A1(n3738), .A2(n2479), .ZN(n3737) );
  NOR2_X1 U3657 ( .A1(n3691), .A2(n3689), .ZN(n3738) );
  NAND2_X1 U3658 ( .A1(n3689), .A2(n3691), .ZN(n3735) );
  NAND2_X1 U3659 ( .A1(n3687), .A2(n3739), .ZN(n3691) );
  NAND2_X1 U3660 ( .A1(n3686), .A2(n3688), .ZN(n3739) );
  NAND2_X1 U3661 ( .A1(n3740), .A2(n3741), .ZN(n3688) );
  NAND2_X1 U3662 ( .A1(b_7_), .A2(a_6_), .ZN(n3741) );
  INV_X1 U3663 ( .A(n3742), .ZN(n3740) );
  XNOR2_X1 U3664 ( .A(n3743), .B(n3744), .ZN(n3686) );
  XOR2_X1 U3665 ( .A(n3745), .B(n3746), .Z(n3744) );
  NAND2_X1 U3666 ( .A1(b_6_), .A2(a_7_), .ZN(n3746) );
  NAND2_X1 U3667 ( .A1(a_6_), .A2(n3742), .ZN(n3687) );
  NAND2_X1 U3668 ( .A1(n3747), .A2(n3748), .ZN(n3742) );
  NAND2_X1 U3669 ( .A1(n3682), .A2(n3749), .ZN(n3748) );
  OR2_X1 U3670 ( .A1(n3684), .A2(n2660), .ZN(n3749) );
  XOR2_X1 U3671 ( .A(n3750), .B(n3751), .Z(n3682) );
  XOR2_X1 U3672 ( .A(n3752), .B(n3753), .Z(n3750) );
  NOR2_X1 U3673 ( .A1(n2689), .A2(n2464), .ZN(n3753) );
  NAND2_X1 U3674 ( .A1(n2660), .A2(n3684), .ZN(n3747) );
  NAND2_X1 U3675 ( .A1(n3754), .A2(n3755), .ZN(n3684) );
  NAND2_X1 U3676 ( .A1(n3756), .A2(b_7_), .ZN(n3755) );
  NOR2_X1 U3677 ( .A1(n3757), .A2(n2689), .ZN(n3756) );
  NOR2_X1 U3678 ( .A1(n3679), .A2(n3680), .ZN(n3757) );
  NAND2_X1 U3679 ( .A1(n3679), .A2(n3680), .ZN(n3754) );
  NAND2_X1 U3680 ( .A1(n3758), .A2(n3759), .ZN(n3680) );
  NAND2_X1 U3681 ( .A1(n3637), .A2(n3760), .ZN(n3759) );
  NAND2_X1 U3682 ( .A1(n3636), .A2(n3635), .ZN(n3760) );
  NOR2_X1 U3683 ( .A1(n2690), .A2(n2383), .ZN(n3637) );
  OR2_X1 U3684 ( .A1(n3635), .A2(n3636), .ZN(n3758) );
  AND2_X1 U3685 ( .A1(n3761), .A2(n3762), .ZN(n3636) );
  NAND2_X1 U3686 ( .A1(n3763), .A2(b_7_), .ZN(n3762) );
  NOR2_X1 U3687 ( .A1(n3764), .A2(n2687), .ZN(n3763) );
  NOR2_X1 U3688 ( .A1(n3675), .A2(n3676), .ZN(n3764) );
  NAND2_X1 U3689 ( .A1(n3675), .A2(n3676), .ZN(n3761) );
  NAND2_X1 U3690 ( .A1(n3765), .A2(n3766), .ZN(n3676) );
  NAND2_X1 U3691 ( .A1(n3673), .A2(n3767), .ZN(n3766) );
  OR2_X1 U3692 ( .A1(n3670), .A2(n3672), .ZN(n3767) );
  NOR2_X1 U3693 ( .A1(n2690), .A2(n2314), .ZN(n3673) );
  NAND2_X1 U3694 ( .A1(n3670), .A2(n3672), .ZN(n3765) );
  NAND2_X1 U3695 ( .A1(n3768), .A2(n3769), .ZN(n3672) );
  NAND2_X1 U3696 ( .A1(n3770), .A2(b_7_), .ZN(n3769) );
  NOR2_X1 U3697 ( .A1(n3771), .A2(n2285), .ZN(n3770) );
  NOR2_X1 U3698 ( .A1(n3667), .A2(n3669), .ZN(n3771) );
  NAND2_X1 U3699 ( .A1(n3667), .A2(n3669), .ZN(n3768) );
  NAND2_X1 U3700 ( .A1(n3772), .A2(n3773), .ZN(n3669) );
  NAND2_X1 U3701 ( .A1(n3662), .A2(n3774), .ZN(n3773) );
  NAND2_X1 U3702 ( .A1(n3665), .A2(n3664), .ZN(n3774) );
  NOR2_X1 U3703 ( .A1(n2690), .A2(n2271), .ZN(n3662) );
  OR2_X1 U3704 ( .A1(n3664), .A2(n3665), .ZN(n3772) );
  AND2_X1 U3705 ( .A1(n3775), .A2(n3776), .ZN(n3665) );
  NAND2_X1 U3706 ( .A1(b_5_), .A2(n3777), .ZN(n3776) );
  NAND2_X1 U3707 ( .A1(n2226), .A2(n3778), .ZN(n3777) );
  NAND2_X1 U3708 ( .A1(a_15_), .A2(n2464), .ZN(n3778) );
  NAND2_X1 U3709 ( .A1(b_6_), .A2(n3779), .ZN(n3775) );
  NAND2_X1 U3710 ( .A1(n2843), .A2(n3780), .ZN(n3779) );
  NAND2_X1 U3711 ( .A1(a_14_), .A2(n2692), .ZN(n3780) );
  NAND2_X1 U3712 ( .A1(n3781), .A2(n2685), .ZN(n3664) );
  NOR2_X1 U3713 ( .A1(n2690), .A2(n2464), .ZN(n3781) );
  XNOR2_X1 U3714 ( .A(n3782), .B(n3783), .ZN(n3667) );
  XNOR2_X1 U3715 ( .A(n3784), .B(n3785), .ZN(n3783) );
  XOR2_X1 U3716 ( .A(n3786), .B(n3787), .Z(n3670) );
  XNOR2_X1 U3717 ( .A(n3788), .B(n3789), .ZN(n3786) );
  NAND2_X1 U3718 ( .A1(b_6_), .A2(a_12_), .ZN(n3788) );
  XNOR2_X1 U3719 ( .A(n3790), .B(n3791), .ZN(n3675) );
  XNOR2_X1 U3720 ( .A(n3792), .B(n3793), .ZN(n3791) );
  XNOR2_X1 U3721 ( .A(n3794), .B(n3795), .ZN(n3635) );
  XOR2_X1 U3722 ( .A(n3796), .B(n3797), .Z(n3794) );
  NOR2_X1 U3723 ( .A1(n2687), .A2(n2464), .ZN(n3797) );
  XNOR2_X1 U3724 ( .A(n3798), .B(n3799), .ZN(n3679) );
  NAND2_X1 U3725 ( .A1(n3800), .A2(n3801), .ZN(n3798) );
  NOR2_X1 U3726 ( .A1(n2690), .A2(n2437), .ZN(n2660) );
  XOR2_X1 U3727 ( .A(n3802), .B(n3803), .Z(n3689) );
  XOR2_X1 U3728 ( .A(n3804), .B(n3805), .Z(n3803) );
  XOR2_X1 U3729 ( .A(n3806), .B(n3807), .Z(n3693) );
  XOR2_X1 U3730 ( .A(n3808), .B(n3809), .Z(n3806) );
  XNOR2_X1 U3731 ( .A(n3810), .B(n3811), .ZN(n3697) );
  XNOR2_X1 U3732 ( .A(n3812), .B(n3813), .ZN(n3811) );
  XNOR2_X1 U3733 ( .A(n3814), .B(n3815), .ZN(n3605) );
  NAND2_X1 U3734 ( .A1(n3816), .A2(n3817), .ZN(n3814) );
  XOR2_X1 U3735 ( .A(n3818), .B(n3819), .Z(n3701) );
  XOR2_X1 U3736 ( .A(n3820), .B(n3821), .Z(n3818) );
  NOR2_X1 U3737 ( .A1(n2695), .A2(n2464), .ZN(n3821) );
  XNOR2_X1 U3738 ( .A(n3822), .B(n3823), .ZN(n3590) );
  XOR2_X1 U3739 ( .A(n3824), .B(n3825), .Z(n3823) );
  NAND2_X1 U3740 ( .A1(b_6_), .A2(a_1_), .ZN(n3825) );
  NAND2_X1 U3741 ( .A1(n3826), .A2(n3827), .ZN(n2190) );
  OR2_X1 U3742 ( .A1(n3714), .A2(n3713), .ZN(n3827) );
  XNOR2_X1 U3743 ( .A(n3828), .B(n3829), .ZN(n3826) );
  NAND2_X1 U3744 ( .A1(n3830), .A2(n3831), .ZN(n2191) );
  XOR2_X1 U3745 ( .A(n3828), .B(n3829), .Z(n3831) );
  NOR2_X1 U3746 ( .A1(n3713), .A2(n3714), .ZN(n3830) );
  XOR2_X1 U3747 ( .A(n3832), .B(n3833), .Z(n3714) );
  XOR2_X1 U3748 ( .A(n3834), .B(n3835), .Z(n3833) );
  NAND2_X1 U3749 ( .A1(b_5_), .A2(a_0_), .ZN(n3835) );
  AND2_X1 U3750 ( .A1(n3836), .A2(n3837), .ZN(n3713) );
  NAND2_X1 U3751 ( .A1(n3838), .A2(b_6_), .ZN(n3837) );
  NOR2_X1 U3752 ( .A1(n3839), .A2(n2623), .ZN(n3838) );
  NOR2_X1 U3753 ( .A1(n3710), .A2(n3708), .ZN(n3839) );
  NAND2_X1 U3754 ( .A1(n3708), .A2(n3710), .ZN(n3836) );
  NAND2_X1 U3755 ( .A1(n3840), .A2(n3841), .ZN(n3710) );
  NAND2_X1 U3756 ( .A1(n3842), .A2(b_6_), .ZN(n3841) );
  NOR2_X1 U3757 ( .A1(n3843), .A2(n2609), .ZN(n3842) );
  NOR2_X1 U3758 ( .A1(n3822), .A2(n3824), .ZN(n3843) );
  NAND2_X1 U3759 ( .A1(n3822), .A2(n3824), .ZN(n3840) );
  NAND2_X1 U3760 ( .A1(n3844), .A2(n3845), .ZN(n3824) );
  NAND2_X1 U3761 ( .A1(n3846), .A2(b_6_), .ZN(n3845) );
  NOR2_X1 U3762 ( .A1(n3847), .A2(n2695), .ZN(n3846) );
  NOR2_X1 U3763 ( .A1(n3820), .A2(n3819), .ZN(n3847) );
  NAND2_X1 U3764 ( .A1(n3819), .A2(n3820), .ZN(n3844) );
  NAND2_X1 U3765 ( .A1(n3816), .A2(n3848), .ZN(n3820) );
  NAND2_X1 U3766 ( .A1(n3815), .A2(n3817), .ZN(n3848) );
  NAND2_X1 U3767 ( .A1(n3849), .A2(n3850), .ZN(n3817) );
  NAND2_X1 U3768 ( .A1(b_6_), .A2(a_3_), .ZN(n3850) );
  INV_X1 U3769 ( .A(n3851), .ZN(n3849) );
  XOR2_X1 U3770 ( .A(n3852), .B(n3853), .Z(n3815) );
  XNOR2_X1 U3771 ( .A(n3854), .B(n3855), .ZN(n3852) );
  NAND2_X1 U3772 ( .A1(b_5_), .A2(a_4_), .ZN(n3854) );
  NAND2_X1 U3773 ( .A1(a_3_), .A2(n3851), .ZN(n3816) );
  NAND2_X1 U3774 ( .A1(n3856), .A2(n3857), .ZN(n3851) );
  NAND2_X1 U3775 ( .A1(n3813), .A2(n3858), .ZN(n3857) );
  OR2_X1 U3776 ( .A1(n3810), .A2(n3812), .ZN(n3858) );
  NOR2_X1 U3777 ( .A1(n2464), .A2(n2506), .ZN(n3813) );
  NAND2_X1 U3778 ( .A1(n3810), .A2(n3812), .ZN(n3856) );
  NAND2_X1 U3779 ( .A1(n3859), .A2(n3860), .ZN(n3812) );
  NAND2_X1 U3780 ( .A1(n3809), .A2(n3861), .ZN(n3860) );
  OR2_X1 U3781 ( .A1(n3808), .A2(n3807), .ZN(n3861) );
  NOR2_X1 U3782 ( .A1(n2464), .A2(n2479), .ZN(n3809) );
  NAND2_X1 U3783 ( .A1(n3807), .A2(n3808), .ZN(n3859) );
  NAND2_X1 U3784 ( .A1(n3862), .A2(n3863), .ZN(n3808) );
  NAND2_X1 U3785 ( .A1(n3805), .A2(n3864), .ZN(n3863) );
  NAND2_X1 U3786 ( .A1(n3804), .A2(n3802), .ZN(n3864) );
  INV_X1 U3787 ( .A(n2657), .ZN(n3805) );
  NAND2_X1 U3788 ( .A1(b_6_), .A2(a_6_), .ZN(n2657) );
  OR2_X1 U3789 ( .A1(n3802), .A2(n3804), .ZN(n3862) );
  AND2_X1 U3790 ( .A1(n3865), .A2(n3866), .ZN(n3804) );
  NAND2_X1 U3791 ( .A1(n3867), .A2(b_6_), .ZN(n3866) );
  NOR2_X1 U3792 ( .A1(n3868), .A2(n2437), .ZN(n3867) );
  NOR2_X1 U3793 ( .A1(n3743), .A2(n3745), .ZN(n3868) );
  NAND2_X1 U3794 ( .A1(n3743), .A2(n3745), .ZN(n3865) );
  NAND2_X1 U3795 ( .A1(n3869), .A2(n3870), .ZN(n3745) );
  NAND2_X1 U3796 ( .A1(n3871), .A2(b_6_), .ZN(n3870) );
  NOR2_X1 U3797 ( .A1(n3872), .A2(n2689), .ZN(n3871) );
  NOR2_X1 U3798 ( .A1(n3752), .A2(n3751), .ZN(n3872) );
  NAND2_X1 U3799 ( .A1(n3751), .A2(n3752), .ZN(n3869) );
  NAND2_X1 U3800 ( .A1(n3800), .A2(n3873), .ZN(n3752) );
  NAND2_X1 U3801 ( .A1(n3799), .A2(n3801), .ZN(n3873) );
  NAND2_X1 U3802 ( .A1(n3874), .A2(n3875), .ZN(n3801) );
  NAND2_X1 U3803 ( .A1(b_6_), .A2(a_9_), .ZN(n3875) );
  INV_X1 U3804 ( .A(n3876), .ZN(n3874) );
  XNOR2_X1 U3805 ( .A(n3877), .B(n3878), .ZN(n3799) );
  XNOR2_X1 U3806 ( .A(n3879), .B(n3880), .ZN(n3877) );
  NAND2_X1 U3807 ( .A1(a_9_), .A2(n3876), .ZN(n3800) );
  NAND2_X1 U3808 ( .A1(n3881), .A2(n3882), .ZN(n3876) );
  NAND2_X1 U3809 ( .A1(n3883), .A2(b_6_), .ZN(n3882) );
  NOR2_X1 U3810 ( .A1(n3884), .A2(n2687), .ZN(n3883) );
  NOR2_X1 U3811 ( .A1(n3796), .A2(n3795), .ZN(n3884) );
  NAND2_X1 U3812 ( .A1(n3795), .A2(n3796), .ZN(n3881) );
  NAND2_X1 U3813 ( .A1(n3885), .A2(n3886), .ZN(n3796) );
  NAND2_X1 U3814 ( .A1(n3793), .A2(n3887), .ZN(n3886) );
  OR2_X1 U3815 ( .A1(n3790), .A2(n3792), .ZN(n3887) );
  NOR2_X1 U3816 ( .A1(n2464), .A2(n2314), .ZN(n3793) );
  NAND2_X1 U3817 ( .A1(n3790), .A2(n3792), .ZN(n3885) );
  NAND2_X1 U3818 ( .A1(n3888), .A2(n3889), .ZN(n3792) );
  NAND2_X1 U3819 ( .A1(n3890), .A2(b_6_), .ZN(n3889) );
  NOR2_X1 U3820 ( .A1(n3891), .A2(n2285), .ZN(n3890) );
  NOR2_X1 U3821 ( .A1(n3787), .A2(n3789), .ZN(n3891) );
  NAND2_X1 U3822 ( .A1(n3787), .A2(n3789), .ZN(n3888) );
  NAND2_X1 U3823 ( .A1(n3892), .A2(n3893), .ZN(n3789) );
  NAND2_X1 U3824 ( .A1(n3782), .A2(n3894), .ZN(n3893) );
  NAND2_X1 U3825 ( .A1(n3785), .A2(n3784), .ZN(n3894) );
  NOR2_X1 U3826 ( .A1(n2464), .A2(n2271), .ZN(n3782) );
  OR2_X1 U3827 ( .A1(n3784), .A2(n3785), .ZN(n3892) );
  AND2_X1 U3828 ( .A1(n3895), .A2(n3896), .ZN(n3785) );
  NAND2_X1 U3829 ( .A1(b_4_), .A2(n3897), .ZN(n3896) );
  NAND2_X1 U3830 ( .A1(n2226), .A2(n3898), .ZN(n3897) );
  NAND2_X1 U3831 ( .A1(a_15_), .A2(n2692), .ZN(n3898) );
  NAND2_X1 U3832 ( .A1(b_5_), .A2(n3899), .ZN(n3895) );
  NAND2_X1 U3833 ( .A1(n2843), .A2(n3900), .ZN(n3899) );
  NAND2_X1 U3834 ( .A1(a_14_), .A2(n2693), .ZN(n3900) );
  NAND2_X1 U3835 ( .A1(n3901), .A2(n2685), .ZN(n3784) );
  NOR2_X1 U3836 ( .A1(n2464), .A2(n2692), .ZN(n3901) );
  XNOR2_X1 U3837 ( .A(n3902), .B(n3903), .ZN(n3787) );
  XNOR2_X1 U3838 ( .A(n3904), .B(n3905), .ZN(n3903) );
  XOR2_X1 U3839 ( .A(n3906), .B(n3907), .Z(n3790) );
  XNOR2_X1 U3840 ( .A(n3908), .B(n3909), .ZN(n3906) );
  NAND2_X1 U3841 ( .A1(b_5_), .A2(a_12_), .ZN(n3908) );
  XNOR2_X1 U3842 ( .A(n3910), .B(n3911), .ZN(n3795) );
  NAND2_X1 U3843 ( .A1(n3912), .A2(n3913), .ZN(n3910) );
  XNOR2_X1 U3844 ( .A(n3914), .B(n3915), .ZN(n3751) );
  NAND2_X1 U3845 ( .A1(n3916), .A2(n3917), .ZN(n3914) );
  XOR2_X1 U3846 ( .A(n3918), .B(n3919), .Z(n3743) );
  XOR2_X1 U3847 ( .A(n3920), .B(n3921), .Z(n3918) );
  NOR2_X1 U3848 ( .A1(n2689), .A2(n2692), .ZN(n3921) );
  XOR2_X1 U3849 ( .A(n3922), .B(n3923), .Z(n3802) );
  XOR2_X1 U3850 ( .A(n3924), .B(n3925), .Z(n3923) );
  NAND2_X1 U3851 ( .A1(b_5_), .A2(a_7_), .ZN(n3925) );
  XNOR2_X1 U3852 ( .A(n3926), .B(n3927), .ZN(n3807) );
  XOR2_X1 U3853 ( .A(n3928), .B(n3929), .Z(n3927) );
  NAND2_X1 U3854 ( .A1(b_5_), .A2(a_6_), .ZN(n3929) );
  XNOR2_X1 U3855 ( .A(n3930), .B(n3931), .ZN(n3810) );
  XNOR2_X1 U3856 ( .A(n2654), .B(n3932), .ZN(n3931) );
  XNOR2_X1 U3857 ( .A(n3933), .B(n3934), .ZN(n3819) );
  XOR2_X1 U3858 ( .A(n3935), .B(n3936), .Z(n3934) );
  NAND2_X1 U3859 ( .A1(b_5_), .A2(a_3_), .ZN(n3936) );
  XNOR2_X1 U3860 ( .A(n3937), .B(n3938), .ZN(n3822) );
  XOR2_X1 U3861 ( .A(n3939), .B(n3940), .Z(n3938) );
  NAND2_X1 U3862 ( .A1(b_5_), .A2(a_2_), .ZN(n3940) );
  XNOR2_X1 U3863 ( .A(n3941), .B(n3942), .ZN(n3708) );
  XOR2_X1 U3864 ( .A(n3943), .B(n3944), .Z(n3942) );
  NAND2_X1 U3865 ( .A1(b_5_), .A2(a_1_), .ZN(n3944) );
  NAND2_X1 U3866 ( .A1(n3945), .A2(n3946), .ZN(n2196) );
  NAND2_X1 U3867 ( .A1(n3829), .A2(n3828), .ZN(n3946) );
  XOR2_X1 U3868 ( .A(n3947), .B(n3948), .Z(n3945) );
  NAND2_X1 U3869 ( .A1(n3949), .A2(n3950), .ZN(n2197) );
  XOR2_X1 U3870 ( .A(n3951), .B(n3948), .Z(n3950) );
  AND2_X1 U3871 ( .A1(n3828), .A2(n3829), .ZN(n3949) );
  XNOR2_X1 U3872 ( .A(n3952), .B(n3953), .ZN(n3829) );
  XOR2_X1 U3873 ( .A(n3954), .B(n3955), .Z(n3953) );
  NAND2_X1 U3874 ( .A1(b_4_), .A2(a_0_), .ZN(n3955) );
  NAND2_X1 U3875 ( .A1(n3956), .A2(n3957), .ZN(n3828) );
  NAND2_X1 U3876 ( .A1(n3958), .A2(b_5_), .ZN(n3957) );
  NOR2_X1 U3877 ( .A1(n3959), .A2(n2623), .ZN(n3958) );
  NOR2_X1 U3878 ( .A1(n3834), .A2(n3832), .ZN(n3959) );
  NAND2_X1 U3879 ( .A1(n3832), .A2(n3834), .ZN(n3956) );
  NAND2_X1 U3880 ( .A1(n3960), .A2(n3961), .ZN(n3834) );
  NAND2_X1 U3881 ( .A1(n3962), .A2(b_5_), .ZN(n3961) );
  NOR2_X1 U3882 ( .A1(n3963), .A2(n2609), .ZN(n3962) );
  NOR2_X1 U3883 ( .A1(n3941), .A2(n3943), .ZN(n3963) );
  NAND2_X1 U3884 ( .A1(n3941), .A2(n3943), .ZN(n3960) );
  NAND2_X1 U3885 ( .A1(n3964), .A2(n3965), .ZN(n3943) );
  NAND2_X1 U3886 ( .A1(n3966), .A2(b_5_), .ZN(n3965) );
  NOR2_X1 U3887 ( .A1(n3967), .A2(n2695), .ZN(n3966) );
  NOR2_X1 U3888 ( .A1(n3939), .A2(n3937), .ZN(n3967) );
  NAND2_X1 U3889 ( .A1(n3937), .A2(n3939), .ZN(n3964) );
  NAND2_X1 U3890 ( .A1(n3968), .A2(n3969), .ZN(n3939) );
  NAND2_X1 U3891 ( .A1(n3970), .A2(b_5_), .ZN(n3969) );
  NOR2_X1 U3892 ( .A1(n3971), .A2(n2553), .ZN(n3970) );
  NOR2_X1 U3893 ( .A1(n3933), .A2(n3935), .ZN(n3971) );
  NAND2_X1 U3894 ( .A1(n3933), .A2(n3935), .ZN(n3968) );
  NAND2_X1 U3895 ( .A1(n3972), .A2(n3973), .ZN(n3935) );
  NAND2_X1 U3896 ( .A1(n3974), .A2(b_5_), .ZN(n3973) );
  NOR2_X1 U3897 ( .A1(n3975), .A2(n2506), .ZN(n3974) );
  NOR2_X1 U3898 ( .A1(n3855), .A2(n3853), .ZN(n3975) );
  NAND2_X1 U3899 ( .A1(n3853), .A2(n3855), .ZN(n3972) );
  NAND2_X1 U3900 ( .A1(n3976), .A2(n3977), .ZN(n3855) );
  NAND2_X1 U3901 ( .A1(n3930), .A2(n3978), .ZN(n3977) );
  OR2_X1 U3902 ( .A1(n3932), .A2(n2654), .ZN(n3978) );
  XNOR2_X1 U3903 ( .A(n3979), .B(n3980), .ZN(n3930) );
  XOR2_X1 U3904 ( .A(n3981), .B(n3982), .Z(n3980) );
  NAND2_X1 U3905 ( .A1(b_4_), .A2(a_6_), .ZN(n3982) );
  NAND2_X1 U3906 ( .A1(n2654), .A2(n3932), .ZN(n3976) );
  NAND2_X1 U3907 ( .A1(n3983), .A2(n3984), .ZN(n3932) );
  NAND2_X1 U3908 ( .A1(n3985), .A2(b_5_), .ZN(n3984) );
  NOR2_X1 U3909 ( .A1(n3986), .A2(n2691), .ZN(n3985) );
  NOR2_X1 U3910 ( .A1(n3928), .A2(n3926), .ZN(n3986) );
  NAND2_X1 U3911 ( .A1(n3926), .A2(n3928), .ZN(n3983) );
  NAND2_X1 U3912 ( .A1(n3987), .A2(n3988), .ZN(n3928) );
  NAND2_X1 U3913 ( .A1(n3989), .A2(b_5_), .ZN(n3988) );
  NOR2_X1 U3914 ( .A1(n3990), .A2(n2437), .ZN(n3989) );
  NOR2_X1 U3915 ( .A1(n3924), .A2(n3922), .ZN(n3990) );
  NAND2_X1 U3916 ( .A1(n3922), .A2(n3924), .ZN(n3987) );
  NAND2_X1 U3917 ( .A1(n3991), .A2(n3992), .ZN(n3924) );
  NAND2_X1 U3918 ( .A1(n3993), .A2(b_5_), .ZN(n3992) );
  NOR2_X1 U3919 ( .A1(n3994), .A2(n2689), .ZN(n3993) );
  NOR2_X1 U3920 ( .A1(n3920), .A2(n3919), .ZN(n3994) );
  NAND2_X1 U3921 ( .A1(n3919), .A2(n3920), .ZN(n3991) );
  NAND2_X1 U3922 ( .A1(n3916), .A2(n3995), .ZN(n3920) );
  NAND2_X1 U3923 ( .A1(n3915), .A2(n3917), .ZN(n3995) );
  NAND2_X1 U3924 ( .A1(n3996), .A2(n3997), .ZN(n3917) );
  NAND2_X1 U3925 ( .A1(b_5_), .A2(a_9_), .ZN(n3997) );
  INV_X1 U3926 ( .A(n3998), .ZN(n3996) );
  XNOR2_X1 U3927 ( .A(n3999), .B(n4000), .ZN(n3915) );
  XNOR2_X1 U3928 ( .A(n4001), .B(n4002), .ZN(n3999) );
  NAND2_X1 U3929 ( .A1(a_9_), .A2(n3998), .ZN(n3916) );
  NAND2_X1 U3930 ( .A1(n4003), .A2(n4004), .ZN(n3998) );
  NAND2_X1 U3931 ( .A1(n3880), .A2(n4005), .ZN(n4004) );
  NAND2_X1 U3932 ( .A1(n3878), .A2(n3879), .ZN(n4005) );
  NOR2_X1 U3933 ( .A1(n2692), .A2(n2687), .ZN(n3880) );
  OR2_X1 U3934 ( .A1(n3878), .A2(n3879), .ZN(n4003) );
  AND2_X1 U3935 ( .A1(n3912), .A2(n4006), .ZN(n3879) );
  NAND2_X1 U3936 ( .A1(n3911), .A2(n3913), .ZN(n4006) );
  NAND2_X1 U3937 ( .A1(n4007), .A2(n4008), .ZN(n3913) );
  NAND2_X1 U3938 ( .A1(b_5_), .A2(a_11_), .ZN(n4008) );
  INV_X1 U3939 ( .A(n4009), .ZN(n4007) );
  XNOR2_X1 U3940 ( .A(n4010), .B(n4011), .ZN(n3911) );
  XOR2_X1 U3941 ( .A(n4012), .B(n4013), .Z(n4011) );
  NAND2_X1 U3942 ( .A1(b_4_), .A2(a_12_), .ZN(n4013) );
  NAND2_X1 U3943 ( .A1(a_11_), .A2(n4009), .ZN(n3912) );
  NAND2_X1 U3944 ( .A1(n4014), .A2(n4015), .ZN(n4009) );
  NAND2_X1 U3945 ( .A1(n4016), .A2(b_5_), .ZN(n4015) );
  NOR2_X1 U3946 ( .A1(n4017), .A2(n2285), .ZN(n4016) );
  NOR2_X1 U3947 ( .A1(n3907), .A2(n3909), .ZN(n4017) );
  NAND2_X1 U3948 ( .A1(n3907), .A2(n3909), .ZN(n4014) );
  NAND2_X1 U3949 ( .A1(n4018), .A2(n4019), .ZN(n3909) );
  NAND2_X1 U3950 ( .A1(n3902), .A2(n4020), .ZN(n4019) );
  NAND2_X1 U3951 ( .A1(n3905), .A2(n3904), .ZN(n4020) );
  NOR2_X1 U3952 ( .A1(n2692), .A2(n2271), .ZN(n3902) );
  OR2_X1 U3953 ( .A1(n3904), .A2(n3905), .ZN(n4018) );
  AND2_X1 U3954 ( .A1(n4021), .A2(n4022), .ZN(n3905) );
  NAND2_X1 U3955 ( .A1(b_3_), .A2(n4023), .ZN(n4022) );
  NAND2_X1 U3956 ( .A1(n2226), .A2(n4024), .ZN(n4023) );
  NAND2_X1 U3957 ( .A1(a_15_), .A2(n2693), .ZN(n4024) );
  NAND2_X1 U3958 ( .A1(b_4_), .A2(n4025), .ZN(n4021) );
  NAND2_X1 U3959 ( .A1(n2843), .A2(n4026), .ZN(n4025) );
  NAND2_X1 U3960 ( .A1(a_14_), .A2(n2694), .ZN(n4026) );
  NAND2_X1 U3961 ( .A1(n4027), .A2(n2685), .ZN(n3904) );
  NOR2_X1 U3962 ( .A1(n2692), .A2(n2693), .ZN(n4027) );
  XOR2_X1 U3963 ( .A(n4028), .B(n4029), .Z(n3907) );
  XNOR2_X1 U3964 ( .A(n4030), .B(n4031), .ZN(n4029) );
  NAND2_X1 U3965 ( .A1(b_4_), .A2(a_13_), .ZN(n4028) );
  XOR2_X1 U3966 ( .A(n4032), .B(n4033), .Z(n3878) );
  NAND2_X1 U3967 ( .A1(n4034), .A2(n4035), .ZN(n4032) );
  XNOR2_X1 U3968 ( .A(n4036), .B(n4037), .ZN(n3919) );
  NAND2_X1 U3969 ( .A1(n4038), .A2(n4039), .ZN(n4036) );
  XOR2_X1 U3970 ( .A(n4040), .B(n4041), .Z(n3922) );
  XOR2_X1 U3971 ( .A(n4042), .B(n4043), .Z(n4040) );
  NOR2_X1 U3972 ( .A1(n2689), .A2(n2693), .ZN(n4043) );
  XNOR2_X1 U3973 ( .A(n4044), .B(n4045), .ZN(n3926) );
  XOR2_X1 U3974 ( .A(n4046), .B(n4047), .Z(n4045) );
  NAND2_X1 U3975 ( .A1(b_4_), .A2(a_7_), .ZN(n4047) );
  NOR2_X1 U3976 ( .A1(n2692), .A2(n2479), .ZN(n2654) );
  XNOR2_X1 U3977 ( .A(n4048), .B(n4049), .ZN(n3853) );
  XOR2_X1 U3978 ( .A(n4050), .B(n4051), .Z(n4049) );
  NAND2_X1 U3979 ( .A1(b_4_), .A2(a_5_), .ZN(n4051) );
  XNOR2_X1 U3980 ( .A(n4052), .B(n4053), .ZN(n3933) );
  XNOR2_X1 U3981 ( .A(n2651), .B(n4054), .ZN(n4053) );
  XOR2_X1 U3982 ( .A(n4055), .B(n4056), .Z(n3937) );
  XNOR2_X1 U3983 ( .A(n4057), .B(n4058), .ZN(n4055) );
  NAND2_X1 U3984 ( .A1(b_4_), .A2(a_3_), .ZN(n4057) );
  XOR2_X1 U3985 ( .A(n4059), .B(n4060), .Z(n3941) );
  XOR2_X1 U3986 ( .A(n4061), .B(n4062), .Z(n4059) );
  NOR2_X1 U3987 ( .A1(n2695), .A2(n2693), .ZN(n4062) );
  XNOR2_X1 U3988 ( .A(n4063), .B(n4064), .ZN(n3832) );
  XOR2_X1 U3989 ( .A(n4065), .B(n4066), .Z(n4064) );
  NAND2_X1 U3990 ( .A1(b_4_), .A2(a_1_), .ZN(n4066) );
  NAND2_X1 U3991 ( .A1(n4067), .A2(n4068), .ZN(n2202) );
  NAND2_X1 U3992 ( .A1(n3948), .A2(n3951), .ZN(n4068) );
  NAND2_X1 U3993 ( .A1(n4069), .A2(n3948), .ZN(n2203) );
  XOR2_X1 U3994 ( .A(n4070), .B(n4071), .Z(n3948) );
  XOR2_X1 U3995 ( .A(n4072), .B(n4073), .Z(n4070) );
  NOR2_X1 U3996 ( .A1(n2623), .A2(n2694), .ZN(n4073) );
  NOR2_X1 U3997 ( .A1(n3947), .A2(n4067), .ZN(n4069) );
  XOR2_X1 U3998 ( .A(n4074), .B(n4075), .Z(n4067) );
  INV_X1 U3999 ( .A(n3951), .ZN(n3947) );
  NAND2_X1 U4000 ( .A1(n4076), .A2(n4077), .ZN(n3951) );
  NAND2_X1 U4001 ( .A1(n4078), .A2(b_4_), .ZN(n4077) );
  NOR2_X1 U4002 ( .A1(n4079), .A2(n2623), .ZN(n4078) );
  NOR2_X1 U4003 ( .A1(n3952), .A2(n3954), .ZN(n4079) );
  NAND2_X1 U4004 ( .A1(n3952), .A2(n3954), .ZN(n4076) );
  NAND2_X1 U4005 ( .A1(n4080), .A2(n4081), .ZN(n3954) );
  NAND2_X1 U4006 ( .A1(n4082), .A2(b_4_), .ZN(n4081) );
  NOR2_X1 U4007 ( .A1(n4083), .A2(n2609), .ZN(n4082) );
  NOR2_X1 U4008 ( .A1(n4063), .A2(n4065), .ZN(n4083) );
  NAND2_X1 U4009 ( .A1(n4063), .A2(n4065), .ZN(n4080) );
  NAND2_X1 U4010 ( .A1(n4084), .A2(n4085), .ZN(n4065) );
  NAND2_X1 U4011 ( .A1(n4086), .A2(b_4_), .ZN(n4085) );
  NOR2_X1 U4012 ( .A1(n4087), .A2(n2695), .ZN(n4086) );
  NOR2_X1 U4013 ( .A1(n4061), .A2(n4060), .ZN(n4087) );
  NAND2_X1 U4014 ( .A1(n4060), .A2(n4061), .ZN(n4084) );
  NAND2_X1 U4015 ( .A1(n4088), .A2(n4089), .ZN(n4061) );
  NAND2_X1 U4016 ( .A1(n4090), .A2(b_4_), .ZN(n4089) );
  NOR2_X1 U4017 ( .A1(n4091), .A2(n2553), .ZN(n4090) );
  NOR2_X1 U4018 ( .A1(n4056), .A2(n4058), .ZN(n4091) );
  NAND2_X1 U4019 ( .A1(n4056), .A2(n4058), .ZN(n4088) );
  NAND2_X1 U4020 ( .A1(n4092), .A2(n4093), .ZN(n4058) );
  NAND2_X1 U4021 ( .A1(n4052), .A2(n4094), .ZN(n4093) );
  OR2_X1 U4022 ( .A1(n4054), .A2(n2651), .ZN(n4094) );
  XNOR2_X1 U4023 ( .A(n4095), .B(n4096), .ZN(n4052) );
  XOR2_X1 U4024 ( .A(n4097), .B(n4098), .Z(n4096) );
  NAND2_X1 U4025 ( .A1(b_3_), .A2(a_5_), .ZN(n4098) );
  NAND2_X1 U4026 ( .A1(n2651), .A2(n4054), .ZN(n4092) );
  NAND2_X1 U4027 ( .A1(n4099), .A2(n4100), .ZN(n4054) );
  NAND2_X1 U4028 ( .A1(n4101), .A2(b_4_), .ZN(n4100) );
  NOR2_X1 U4029 ( .A1(n4102), .A2(n2479), .ZN(n4101) );
  NOR2_X1 U4030 ( .A1(n4048), .A2(n4050), .ZN(n4102) );
  NAND2_X1 U4031 ( .A1(n4048), .A2(n4050), .ZN(n4099) );
  NAND2_X1 U4032 ( .A1(n4103), .A2(n4104), .ZN(n4050) );
  NAND2_X1 U4033 ( .A1(n4105), .A2(b_4_), .ZN(n4104) );
  NOR2_X1 U4034 ( .A1(n4106), .A2(n2691), .ZN(n4105) );
  NOR2_X1 U4035 ( .A1(n3981), .A2(n3979), .ZN(n4106) );
  NAND2_X1 U4036 ( .A1(n3979), .A2(n3981), .ZN(n4103) );
  NAND2_X1 U4037 ( .A1(n4107), .A2(n4108), .ZN(n3981) );
  NAND2_X1 U4038 ( .A1(n4109), .A2(b_4_), .ZN(n4108) );
  NOR2_X1 U4039 ( .A1(n4110), .A2(n2437), .ZN(n4109) );
  NOR2_X1 U4040 ( .A1(n4044), .A2(n4046), .ZN(n4110) );
  NAND2_X1 U4041 ( .A1(n4044), .A2(n4046), .ZN(n4107) );
  NAND2_X1 U4042 ( .A1(n4111), .A2(n4112), .ZN(n4046) );
  NAND2_X1 U4043 ( .A1(n4113), .A2(b_4_), .ZN(n4112) );
  NOR2_X1 U4044 ( .A1(n4114), .A2(n2689), .ZN(n4113) );
  NOR2_X1 U4045 ( .A1(n4041), .A2(n4042), .ZN(n4114) );
  NAND2_X1 U4046 ( .A1(n4041), .A2(n4042), .ZN(n4111) );
  NAND2_X1 U4047 ( .A1(n4038), .A2(n4115), .ZN(n4042) );
  NAND2_X1 U4048 ( .A1(n4037), .A2(n4039), .ZN(n4115) );
  NAND2_X1 U4049 ( .A1(n4116), .A2(n4117), .ZN(n4039) );
  NAND2_X1 U4050 ( .A1(b_4_), .A2(a_9_), .ZN(n4117) );
  INV_X1 U4051 ( .A(n4118), .ZN(n4116) );
  XNOR2_X1 U4052 ( .A(n4119), .B(n4120), .ZN(n4037) );
  NAND2_X1 U4053 ( .A1(n4121), .A2(n4122), .ZN(n4119) );
  NAND2_X1 U4054 ( .A1(a_9_), .A2(n4118), .ZN(n4038) );
  NAND2_X1 U4055 ( .A1(n4123), .A2(n4124), .ZN(n4118) );
  NAND2_X1 U4056 ( .A1(n4002), .A2(n4125), .ZN(n4124) );
  NAND2_X1 U4057 ( .A1(n4001), .A2(n4000), .ZN(n4125) );
  NOR2_X1 U4058 ( .A1(n2693), .A2(n2687), .ZN(n4002) );
  OR2_X1 U4059 ( .A1(n4000), .A2(n4001), .ZN(n4123) );
  AND2_X1 U4060 ( .A1(n4034), .A2(n4126), .ZN(n4001) );
  NAND2_X1 U4061 ( .A1(n4033), .A2(n4035), .ZN(n4126) );
  NAND2_X1 U4062 ( .A1(n4127), .A2(n4128), .ZN(n4035) );
  NAND2_X1 U4063 ( .A1(b_4_), .A2(a_11_), .ZN(n4128) );
  INV_X1 U4064 ( .A(n4129), .ZN(n4127) );
  XNOR2_X1 U4065 ( .A(n4130), .B(n4131), .ZN(n4033) );
  XNOR2_X1 U4066 ( .A(n4132), .B(n4133), .ZN(n4131) );
  NAND2_X1 U4067 ( .A1(a_11_), .A2(n4129), .ZN(n4034) );
  NAND2_X1 U4068 ( .A1(n4134), .A2(n4135), .ZN(n4129) );
  NAND2_X1 U4069 ( .A1(n4136), .A2(b_4_), .ZN(n4135) );
  NOR2_X1 U4070 ( .A1(n4137), .A2(n2285), .ZN(n4136) );
  NOR2_X1 U4071 ( .A1(n4010), .A2(n4012), .ZN(n4137) );
  NAND2_X1 U4072 ( .A1(n4010), .A2(n4012), .ZN(n4134) );
  NAND2_X1 U4073 ( .A1(n4138), .A2(n4139), .ZN(n4012) );
  NAND2_X1 U4074 ( .A1(n4140), .A2(b_4_), .ZN(n4139) );
  NOR2_X1 U4075 ( .A1(n4141), .A2(n2271), .ZN(n4140) );
  NOR2_X1 U4076 ( .A1(n4030), .A2(n4031), .ZN(n4141) );
  NAND2_X1 U4077 ( .A1(n4030), .A2(n4031), .ZN(n4138) );
  NAND2_X1 U4078 ( .A1(n4142), .A2(n4143), .ZN(n4031) );
  NAND2_X1 U4079 ( .A1(b_2_), .A2(n4144), .ZN(n4143) );
  NAND2_X1 U4080 ( .A1(n2226), .A2(n4145), .ZN(n4144) );
  NAND2_X1 U4081 ( .A1(a_15_), .A2(n2694), .ZN(n4145) );
  NAND2_X1 U4082 ( .A1(b_3_), .A2(n4146), .ZN(n4142) );
  NAND2_X1 U4083 ( .A1(n2843), .A2(n4147), .ZN(n4146) );
  NAND2_X1 U4084 ( .A1(a_14_), .A2(n2581), .ZN(n4147) );
  AND2_X1 U4085 ( .A1(n4148), .A2(n2685), .ZN(n4030) );
  NOR2_X1 U4086 ( .A1(n2693), .A2(n2694), .ZN(n4148) );
  XOR2_X1 U4087 ( .A(n4149), .B(n4150), .Z(n4010) );
  XNOR2_X1 U4088 ( .A(n4151), .B(n4152), .ZN(n4150) );
  NAND2_X1 U4089 ( .A1(b_3_), .A2(a_13_), .ZN(n4149) );
  XOR2_X1 U4090 ( .A(n4153), .B(n4154), .Z(n4000) );
  NAND2_X1 U4091 ( .A1(n4155), .A2(n4156), .ZN(n4153) );
  XNOR2_X1 U4092 ( .A(n4157), .B(n4158), .ZN(n4041) );
  NAND2_X1 U4093 ( .A1(n4159), .A2(n4160), .ZN(n4157) );
  XOR2_X1 U4094 ( .A(n4161), .B(n4162), .Z(n4044) );
  XOR2_X1 U4095 ( .A(n4163), .B(n4164), .Z(n4161) );
  NOR2_X1 U4096 ( .A1(n2689), .A2(n2694), .ZN(n4164) );
  XNOR2_X1 U4097 ( .A(n4165), .B(n4166), .ZN(n3979) );
  XOR2_X1 U4098 ( .A(n4167), .B(n4168), .Z(n4166) );
  NAND2_X1 U4099 ( .A1(b_3_), .A2(a_7_), .ZN(n4168) );
  XNOR2_X1 U4100 ( .A(n4169), .B(n4170), .ZN(n4048) );
  XOR2_X1 U4101 ( .A(n4171), .B(n4172), .Z(n4170) );
  NAND2_X1 U4102 ( .A1(b_3_), .A2(a_6_), .ZN(n4172) );
  NOR2_X1 U4103 ( .A1(n2693), .A2(n2506), .ZN(n2651) );
  XNOR2_X1 U4104 ( .A(n4173), .B(n4174), .ZN(n4056) );
  XOR2_X1 U4105 ( .A(n4175), .B(n4176), .Z(n4174) );
  NAND2_X1 U4106 ( .A1(b_3_), .A2(a_4_), .ZN(n4176) );
  XNOR2_X1 U4107 ( .A(n4177), .B(n4178), .ZN(n4060) );
  XNOR2_X1 U4108 ( .A(n2648), .B(n4179), .ZN(n4178) );
  XOR2_X1 U4109 ( .A(n4180), .B(n4181), .Z(n4063) );
  XNOR2_X1 U4110 ( .A(n4182), .B(n4183), .ZN(n4180) );
  NAND2_X1 U4111 ( .A1(b_3_), .A2(a_2_), .ZN(n4182) );
  XOR2_X1 U4112 ( .A(n4184), .B(n4185), .Z(n3952) );
  XOR2_X1 U4113 ( .A(n4186), .B(n4187), .Z(n4184) );
  NOR2_X1 U4114 ( .A1(n2609), .A2(n2694), .ZN(n4187) );
  NAND2_X1 U4115 ( .A1(n4188), .A2(n4189), .ZN(n2249) );
  NAND2_X1 U4116 ( .A1(n4190), .A2(n4074), .ZN(n4189) );
  INV_X1 U4117 ( .A(n4075), .ZN(n4190) );
  XNOR2_X1 U4118 ( .A(n4191), .B(n4192), .ZN(n4188) );
  NAND2_X1 U4119 ( .A1(n4193), .A2(n4194), .ZN(n2250) );
  AND2_X1 U4120 ( .A1(n2742), .A2(n4074), .ZN(n4194) );
  NAND2_X1 U4121 ( .A1(n4195), .A2(n4196), .ZN(n4074) );
  NAND2_X1 U4122 ( .A1(n4197), .A2(b_3_), .ZN(n4196) );
  NOR2_X1 U4123 ( .A1(n4198), .A2(n2623), .ZN(n4197) );
  NOR2_X1 U4124 ( .A1(n4072), .A2(n4071), .ZN(n4198) );
  NAND2_X1 U4125 ( .A1(n4071), .A2(n4072), .ZN(n4195) );
  NAND2_X1 U4126 ( .A1(n4199), .A2(n4200), .ZN(n4072) );
  NAND2_X1 U4127 ( .A1(n4201), .A2(b_3_), .ZN(n4200) );
  NOR2_X1 U4128 ( .A1(n4202), .A2(n2609), .ZN(n4201) );
  NOR2_X1 U4129 ( .A1(n4186), .A2(n4185), .ZN(n4202) );
  NAND2_X1 U4130 ( .A1(n4185), .A2(n4186), .ZN(n4199) );
  NAND2_X1 U4131 ( .A1(n4203), .A2(n4204), .ZN(n4186) );
  NAND2_X1 U4132 ( .A1(n4205), .A2(b_3_), .ZN(n4204) );
  NOR2_X1 U4133 ( .A1(n4206), .A2(n2695), .ZN(n4205) );
  NOR2_X1 U4134 ( .A1(n4183), .A2(n4181), .ZN(n4206) );
  NAND2_X1 U4135 ( .A1(n4181), .A2(n4183), .ZN(n4203) );
  NAND2_X1 U4136 ( .A1(n4207), .A2(n4208), .ZN(n4183) );
  NAND2_X1 U4137 ( .A1(n4177), .A2(n4209), .ZN(n4208) );
  OR2_X1 U4138 ( .A1(n4179), .A2(n2648), .ZN(n4209) );
  XNOR2_X1 U4139 ( .A(n4210), .B(n4211), .ZN(n4177) );
  NAND2_X1 U4140 ( .A1(n4212), .A2(n4213), .ZN(n4210) );
  NAND2_X1 U4141 ( .A1(n2648), .A2(n4179), .ZN(n4207) );
  NAND2_X1 U4142 ( .A1(n4214), .A2(n4215), .ZN(n4179) );
  NAND2_X1 U4143 ( .A1(n4216), .A2(b_3_), .ZN(n4215) );
  NOR2_X1 U4144 ( .A1(n4217), .A2(n2506), .ZN(n4216) );
  NOR2_X1 U4145 ( .A1(n4175), .A2(n4173), .ZN(n4217) );
  NAND2_X1 U4146 ( .A1(n4173), .A2(n4175), .ZN(n4214) );
  NAND2_X1 U4147 ( .A1(n4218), .A2(n4219), .ZN(n4175) );
  NAND2_X1 U4148 ( .A1(n4220), .A2(b_3_), .ZN(n4219) );
  NOR2_X1 U4149 ( .A1(n4221), .A2(n2479), .ZN(n4220) );
  NOR2_X1 U4150 ( .A1(n4095), .A2(n4097), .ZN(n4221) );
  NAND2_X1 U4151 ( .A1(n4095), .A2(n4097), .ZN(n4218) );
  NAND2_X1 U4152 ( .A1(n4222), .A2(n4223), .ZN(n4097) );
  NAND2_X1 U4153 ( .A1(n4224), .A2(b_3_), .ZN(n4223) );
  NOR2_X1 U4154 ( .A1(n4225), .A2(n2691), .ZN(n4224) );
  NOR2_X1 U4155 ( .A1(n4171), .A2(n4169), .ZN(n4225) );
  NAND2_X1 U4156 ( .A1(n4169), .A2(n4171), .ZN(n4222) );
  NAND2_X1 U4157 ( .A1(n4226), .A2(n4227), .ZN(n4171) );
  NAND2_X1 U4158 ( .A1(n4228), .A2(b_3_), .ZN(n4227) );
  NOR2_X1 U4159 ( .A1(n4229), .A2(n2437), .ZN(n4228) );
  NOR2_X1 U4160 ( .A1(n4165), .A2(n4167), .ZN(n4229) );
  NAND2_X1 U4161 ( .A1(n4165), .A2(n4167), .ZN(n4226) );
  NAND2_X1 U4162 ( .A1(n4230), .A2(n4231), .ZN(n4167) );
  NAND2_X1 U4163 ( .A1(n4232), .A2(b_3_), .ZN(n4231) );
  NOR2_X1 U4164 ( .A1(n4233), .A2(n2689), .ZN(n4232) );
  NOR2_X1 U4165 ( .A1(n4163), .A2(n4162), .ZN(n4233) );
  NAND2_X1 U4166 ( .A1(n4162), .A2(n4163), .ZN(n4230) );
  NAND2_X1 U4167 ( .A1(n4159), .A2(n4234), .ZN(n4163) );
  NAND2_X1 U4168 ( .A1(n4158), .A2(n4160), .ZN(n4234) );
  NAND2_X1 U4169 ( .A1(n4235), .A2(n4236), .ZN(n4160) );
  NAND2_X1 U4170 ( .A1(b_3_), .A2(a_9_), .ZN(n4236) );
  INV_X1 U4171 ( .A(n4237), .ZN(n4235) );
  XNOR2_X1 U4172 ( .A(n4238), .B(n4239), .ZN(n4158) );
  NAND2_X1 U4173 ( .A1(n4240), .A2(n4241), .ZN(n4238) );
  NAND2_X1 U4174 ( .A1(a_9_), .A2(n4237), .ZN(n4159) );
  NAND2_X1 U4175 ( .A1(n4121), .A2(n4242), .ZN(n4237) );
  NAND2_X1 U4176 ( .A1(n4120), .A2(n4122), .ZN(n4242) );
  NAND2_X1 U4177 ( .A1(n4243), .A2(n4244), .ZN(n4122) );
  NAND2_X1 U4178 ( .A1(b_3_), .A2(a_10_), .ZN(n4244) );
  INV_X1 U4179 ( .A(n4245), .ZN(n4243) );
  XNOR2_X1 U4180 ( .A(n4246), .B(n4247), .ZN(n4120) );
  XNOR2_X1 U4181 ( .A(n4248), .B(n4249), .ZN(n4246) );
  NAND2_X1 U4182 ( .A1(a_10_), .A2(n4245), .ZN(n4121) );
  NAND2_X1 U4183 ( .A1(n4155), .A2(n4250), .ZN(n4245) );
  NAND2_X1 U4184 ( .A1(n4154), .A2(n4156), .ZN(n4250) );
  NAND2_X1 U4185 ( .A1(n4251), .A2(n4252), .ZN(n4156) );
  NAND2_X1 U4186 ( .A1(b_3_), .A2(a_11_), .ZN(n4252) );
  INV_X1 U4187 ( .A(n4253), .ZN(n4251) );
  XNOR2_X1 U4188 ( .A(n4254), .B(n4255), .ZN(n4154) );
  XNOR2_X1 U4189 ( .A(n4256), .B(n4257), .ZN(n4255) );
  NAND2_X1 U4190 ( .A1(a_11_), .A2(n4253), .ZN(n4155) );
  NAND2_X1 U4191 ( .A1(n4258), .A2(n4259), .ZN(n4253) );
  NAND2_X1 U4192 ( .A1(n4133), .A2(n4260), .ZN(n4259) );
  OR2_X1 U4193 ( .A1(n4132), .A2(n4130), .ZN(n4260) );
  NOR2_X1 U4194 ( .A1(n2694), .A2(n2285), .ZN(n4133) );
  NAND2_X1 U4195 ( .A1(n4130), .A2(n4132), .ZN(n4258) );
  NAND2_X1 U4196 ( .A1(n4261), .A2(n4262), .ZN(n4132) );
  NAND2_X1 U4197 ( .A1(n4263), .A2(b_3_), .ZN(n4262) );
  NOR2_X1 U4198 ( .A1(n4264), .A2(n2271), .ZN(n4263) );
  NOR2_X1 U4199 ( .A1(n4152), .A2(n4151), .ZN(n4264) );
  NAND2_X1 U4200 ( .A1(n4152), .A2(n4151), .ZN(n4261) );
  NAND2_X1 U4201 ( .A1(n4265), .A2(n4266), .ZN(n4151) );
  NAND2_X1 U4202 ( .A1(b_1_), .A2(n4267), .ZN(n4266) );
  NAND2_X1 U4203 ( .A1(n4268), .A2(n2226), .ZN(n4267) );
  NAND2_X1 U4204 ( .A1(a_15_), .A2(n2581), .ZN(n4268) );
  NAND2_X1 U4205 ( .A1(b_2_), .A2(n4269), .ZN(n4265) );
  NAND2_X1 U4206 ( .A1(n4270), .A2(n2843), .ZN(n4269) );
  NAND2_X1 U4207 ( .A1(a_14_), .A2(n2696), .ZN(n4270) );
  AND2_X1 U4208 ( .A1(n4271), .A2(n2685), .ZN(n4152) );
  NOR2_X1 U4209 ( .A1(n2694), .A2(n2581), .ZN(n4271) );
  XOR2_X1 U4210 ( .A(n4272), .B(n4273), .Z(n4130) );
  XNOR2_X1 U4211 ( .A(n4274), .B(n4275), .ZN(n4273) );
  NAND2_X1 U4212 ( .A1(b_2_), .A2(a_13_), .ZN(n4272) );
  XNOR2_X1 U4213 ( .A(n4276), .B(n4277), .ZN(n4162) );
  XNOR2_X1 U4214 ( .A(n4278), .B(n4279), .ZN(n4276) );
  XNOR2_X1 U4215 ( .A(n4280), .B(n4281), .ZN(n4165) );
  NAND2_X1 U4216 ( .A1(n4282), .A2(n4283), .ZN(n4280) );
  XOR2_X1 U4217 ( .A(n4284), .B(n4285), .Z(n4169) );
  XOR2_X1 U4218 ( .A(n4286), .B(n4287), .Z(n4285) );
  XNOR2_X1 U4219 ( .A(n4288), .B(n4289), .ZN(n4095) );
  NAND2_X1 U4220 ( .A1(n4290), .A2(n4291), .ZN(n4288) );
  XOR2_X1 U4221 ( .A(n4292), .B(n4293), .Z(n4173) );
  XOR2_X1 U4222 ( .A(n4294), .B(n4295), .Z(n4292) );
  NOR2_X1 U4223 ( .A1(n2694), .A2(n2553), .ZN(n2648) );
  XNOR2_X1 U4224 ( .A(n4296), .B(n4297), .ZN(n4181) );
  XNOR2_X1 U4225 ( .A(n4298), .B(n4299), .ZN(n4296) );
  XOR2_X1 U4226 ( .A(n4300), .B(n4301), .Z(n4185) );
  XOR2_X1 U4227 ( .A(n4302), .B(n4303), .Z(n4300) );
  XNOR2_X1 U4228 ( .A(n4304), .B(n4305), .ZN(n4071) );
  XNOR2_X1 U4229 ( .A(n4306), .B(n4307), .ZN(n4304) );
  NOR2_X1 U4230 ( .A1(n4308), .A2(n4075), .ZN(n4193) );
  XOR2_X1 U4231 ( .A(n4309), .B(n4310), .Z(n4075) );
  NAND2_X1 U4232 ( .A1(n4311), .A2(n4312), .ZN(n4309) );
  NOR2_X1 U4233 ( .A1(n4192), .A2(n4191), .ZN(n4308) );
  AND2_X1 U4234 ( .A1(n4313), .A2(n4314), .ZN(n2532) );
  NOR2_X1 U4235 ( .A1(n2623), .A2(n2637), .ZN(n4314) );
  NOR2_X1 U4236 ( .A1(n2739), .A2(n2742), .ZN(n4313) );
  NAND2_X1 U4237 ( .A1(n4192), .A2(n4191), .ZN(n2742) );
  NAND2_X1 U4238 ( .A1(n4311), .A2(n4315), .ZN(n4191) );
  NAND2_X1 U4239 ( .A1(n4310), .A2(n4312), .ZN(n4315) );
  NAND2_X1 U4240 ( .A1(n4316), .A2(n4317), .ZN(n4312) );
  NAND2_X1 U4241 ( .A1(b_2_), .A2(a_0_), .ZN(n4317) );
  INV_X1 U4242 ( .A(n4318), .ZN(n4316) );
  XOR2_X1 U4243 ( .A(n4319), .B(n4320), .Z(n4310) );
  XNOR2_X1 U4244 ( .A(n2644), .B(n4321), .ZN(n4320) );
  NAND2_X1 U4245 ( .A1(b_0_), .A2(a_2_), .ZN(n4319) );
  NAND2_X1 U4246 ( .A1(a_0_), .A2(n4318), .ZN(n4311) );
  NAND2_X1 U4247 ( .A1(n4322), .A2(n4323), .ZN(n4318) );
  NAND2_X1 U4248 ( .A1(n4307), .A2(n4324), .ZN(n4323) );
  NAND2_X1 U4249 ( .A1(n4306), .A2(n4305), .ZN(n4324) );
  NOR2_X1 U4250 ( .A1(n2581), .A2(n2609), .ZN(n4307) );
  OR2_X1 U4251 ( .A1(n4305), .A2(n4306), .ZN(n4322) );
  AND2_X1 U4252 ( .A1(n4325), .A2(n4326), .ZN(n4306) );
  NAND2_X1 U4253 ( .A1(n4301), .A2(n4327), .ZN(n4326) );
  OR2_X1 U4254 ( .A1(n4302), .A2(n4303), .ZN(n4327) );
  XOR2_X1 U4255 ( .A(n4328), .B(n4329), .Z(n4301) );
  XNOR2_X1 U4256 ( .A(n4330), .B(n4331), .ZN(n4329) );
  NAND2_X1 U4257 ( .A1(b_1_), .A2(a_3_), .ZN(n4328) );
  NAND2_X1 U4258 ( .A1(n4303), .A2(n4302), .ZN(n4325) );
  NAND2_X1 U4259 ( .A1(n4332), .A2(n4333), .ZN(n4302) );
  NAND2_X1 U4260 ( .A1(n4299), .A2(n4334), .ZN(n4333) );
  NAND2_X1 U4261 ( .A1(n4298), .A2(n4297), .ZN(n4334) );
  NOR2_X1 U4262 ( .A1(n2581), .A2(n2553), .ZN(n4299) );
  OR2_X1 U4263 ( .A1(n4297), .A2(n4298), .ZN(n4332) );
  AND2_X1 U4264 ( .A1(n4212), .A2(n4335), .ZN(n4298) );
  NAND2_X1 U4265 ( .A1(n4211), .A2(n4213), .ZN(n4335) );
  NAND2_X1 U4266 ( .A1(n4336), .A2(n4337), .ZN(n4213) );
  NAND2_X1 U4267 ( .A1(b_2_), .A2(a_4_), .ZN(n4337) );
  INV_X1 U4268 ( .A(n4338), .ZN(n4336) );
  XOR2_X1 U4269 ( .A(n4339), .B(n4340), .Z(n4211) );
  XNOR2_X1 U4270 ( .A(n4341), .B(n4342), .ZN(n4340) );
  NAND2_X1 U4271 ( .A1(b_1_), .A2(a_5_), .ZN(n4339) );
  NAND2_X1 U4272 ( .A1(a_4_), .A2(n4338), .ZN(n4212) );
  NAND2_X1 U4273 ( .A1(n4343), .A2(n4344), .ZN(n4338) );
  NAND2_X1 U4274 ( .A1(n4295), .A2(n4345), .ZN(n4344) );
  OR2_X1 U4275 ( .A1(n4294), .A2(n4293), .ZN(n4345) );
  NOR2_X1 U4276 ( .A1(n2581), .A2(n2479), .ZN(n4295) );
  NAND2_X1 U4277 ( .A1(n4293), .A2(n4294), .ZN(n4343) );
  NAND2_X1 U4278 ( .A1(n4290), .A2(n4346), .ZN(n4294) );
  NAND2_X1 U4279 ( .A1(n4289), .A2(n4291), .ZN(n4346) );
  NAND2_X1 U4280 ( .A1(n4347), .A2(n4348), .ZN(n4291) );
  NAND2_X1 U4281 ( .A1(b_2_), .A2(a_6_), .ZN(n4348) );
  INV_X1 U4282 ( .A(n4349), .ZN(n4347) );
  XOR2_X1 U4283 ( .A(n4350), .B(n4351), .Z(n4289) );
  XNOR2_X1 U4284 ( .A(n4352), .B(n4353), .ZN(n4351) );
  NAND2_X1 U4285 ( .A1(b_1_), .A2(a_7_), .ZN(n4350) );
  NAND2_X1 U4286 ( .A1(a_6_), .A2(n4349), .ZN(n4290) );
  NAND2_X1 U4287 ( .A1(n4354), .A2(n4355), .ZN(n4349) );
  NAND2_X1 U4288 ( .A1(n4287), .A2(n4356), .ZN(n4355) );
  NAND2_X1 U4289 ( .A1(n4286), .A2(n4284), .ZN(n4356) );
  NOR2_X1 U4290 ( .A1(n2581), .A2(n2437), .ZN(n4287) );
  OR2_X1 U4291 ( .A1(n4284), .A2(n4286), .ZN(n4354) );
  AND2_X1 U4292 ( .A1(n4282), .A2(n4357), .ZN(n4286) );
  NAND2_X1 U4293 ( .A1(n4281), .A2(n4283), .ZN(n4357) );
  NAND2_X1 U4294 ( .A1(n4358), .A2(n4359), .ZN(n4283) );
  NAND2_X1 U4295 ( .A1(b_2_), .A2(a_8_), .ZN(n4359) );
  INV_X1 U4296 ( .A(n4360), .ZN(n4358) );
  XOR2_X1 U4297 ( .A(n4361), .B(n4362), .Z(n4281) );
  XNOR2_X1 U4298 ( .A(n4363), .B(n4364), .ZN(n4362) );
  NAND2_X1 U4299 ( .A1(b_1_), .A2(a_9_), .ZN(n4361) );
  NAND2_X1 U4300 ( .A1(a_8_), .A2(n4360), .ZN(n4282) );
  NAND2_X1 U4301 ( .A1(n4365), .A2(n4366), .ZN(n4360) );
  NAND2_X1 U4302 ( .A1(n4278), .A2(n4367), .ZN(n4366) );
  NAND2_X1 U4303 ( .A1(n4279), .A2(n4277), .ZN(n4367) );
  NOR2_X1 U4304 ( .A1(n2581), .A2(n2383), .ZN(n4278) );
  OR2_X1 U4305 ( .A1(n4277), .A2(n4279), .ZN(n4365) );
  AND2_X1 U4306 ( .A1(n4240), .A2(n4368), .ZN(n4279) );
  NAND2_X1 U4307 ( .A1(n4239), .A2(n4241), .ZN(n4368) );
  NAND2_X1 U4308 ( .A1(n4369), .A2(n4370), .ZN(n4241) );
  NAND2_X1 U4309 ( .A1(b_2_), .A2(a_10_), .ZN(n4370) );
  INV_X1 U4310 ( .A(n4371), .ZN(n4369) );
  XOR2_X1 U4311 ( .A(n4372), .B(n4373), .Z(n4239) );
  XNOR2_X1 U4312 ( .A(n4374), .B(n4375), .ZN(n4373) );
  NAND2_X1 U4313 ( .A1(b_1_), .A2(a_11_), .ZN(n4372) );
  NAND2_X1 U4314 ( .A1(a_10_), .A2(n4371), .ZN(n4240) );
  NAND2_X1 U4315 ( .A1(n4376), .A2(n4377), .ZN(n4371) );
  NAND2_X1 U4316 ( .A1(n4248), .A2(n4378), .ZN(n4377) );
  NAND2_X1 U4317 ( .A1(n4249), .A2(n4247), .ZN(n4378) );
  NOR2_X1 U4318 ( .A1(n2581), .A2(n2314), .ZN(n4248) );
  OR2_X1 U4319 ( .A1(n4247), .A2(n4249), .ZN(n4376) );
  AND2_X1 U4320 ( .A1(n4379), .A2(n4380), .ZN(n4249) );
  NAND2_X1 U4321 ( .A1(n4257), .A2(n4381), .ZN(n4380) );
  OR2_X1 U4322 ( .A1(n4254), .A2(n4256), .ZN(n4381) );
  NOR2_X1 U4323 ( .A1(n2581), .A2(n2285), .ZN(n4257) );
  NAND2_X1 U4324 ( .A1(n4254), .A2(n4256), .ZN(n4379) );
  NAND2_X1 U4325 ( .A1(n4382), .A2(n4383), .ZN(n4256) );
  NAND2_X1 U4326 ( .A1(n4384), .A2(b_2_), .ZN(n4383) );
  NOR2_X1 U4327 ( .A1(n4385), .A2(n2271), .ZN(n4384) );
  NOR2_X1 U4328 ( .A1(n4275), .A2(n4274), .ZN(n4385) );
  NAND2_X1 U4329 ( .A1(n4275), .A2(n4274), .ZN(n4382) );
  NAND2_X1 U4330 ( .A1(n4386), .A2(n4387), .ZN(n4274) );
  NAND2_X1 U4331 ( .A1(b_0_), .A2(n4388), .ZN(n4387) );
  NAND2_X1 U4332 ( .A1(n4389), .A2(n2226), .ZN(n4388) );
  NAND2_X1 U4333 ( .A1(a_15_), .A2(n2684), .ZN(n2226) );
  NAND2_X1 U4334 ( .A1(a_15_), .A2(n2696), .ZN(n4389) );
  NAND2_X1 U4335 ( .A1(b_1_), .A2(n4390), .ZN(n4386) );
  NAND2_X1 U4336 ( .A1(n4391), .A2(n2843), .ZN(n4390) );
  NAND2_X1 U4337 ( .A1(a_14_), .A2(n4392), .ZN(n2843) );
  NAND2_X1 U4338 ( .A1(a_14_), .A2(n2637), .ZN(n4391) );
  AND2_X1 U4339 ( .A1(n4393), .A2(n2685), .ZN(n4275) );
  NOR2_X1 U4340 ( .A1(n2581), .A2(n2696), .ZN(n4393) );
  XNOR2_X1 U4341 ( .A(n4394), .B(n4395), .ZN(n4254) );
  XOR2_X1 U4342 ( .A(n4396), .B(n4397), .Z(n4394) );
  XNOR2_X1 U4343 ( .A(n4398), .B(n4399), .ZN(n4247) );
  NOR2_X1 U4344 ( .A1(n2285), .A2(n2696), .ZN(n4399) );
  XOR2_X1 U4345 ( .A(n4400), .B(n4401), .Z(n4398) );
  XOR2_X1 U4346 ( .A(n4402), .B(n4403), .Z(n4277) );
  NAND2_X1 U4347 ( .A1(n4404), .A2(n4405), .ZN(n4402) );
  NAND2_X1 U4348 ( .A1(n4406), .A2(n4407), .ZN(n4405) );
  NAND2_X1 U4349 ( .A1(b_1_), .A2(a_10_), .ZN(n4406) );
  XOR2_X1 U4350 ( .A(n4408), .B(n4409), .Z(n4284) );
  NAND2_X1 U4351 ( .A1(n4410), .A2(n4411), .ZN(n4408) );
  NAND2_X1 U4352 ( .A1(n4412), .A2(n4413), .ZN(n4411) );
  NAND2_X1 U4353 ( .A1(b_1_), .A2(a_8_), .ZN(n4412) );
  XNOR2_X1 U4354 ( .A(n4414), .B(n4415), .ZN(n4293) );
  NAND2_X1 U4355 ( .A1(n4416), .A2(n4417), .ZN(n4414) );
  NAND2_X1 U4356 ( .A1(n4418), .A2(n4419), .ZN(n4417) );
  NAND2_X1 U4357 ( .A1(b_1_), .A2(a_6_), .ZN(n4418) );
  XOR2_X1 U4358 ( .A(n4420), .B(n4421), .Z(n4297) );
  NAND2_X1 U4359 ( .A1(n4422), .A2(n4423), .ZN(n4420) );
  NAND2_X1 U4360 ( .A1(n4424), .A2(n4425), .ZN(n4423) );
  NAND2_X1 U4361 ( .A1(b_1_), .A2(a_4_), .ZN(n4424) );
  INV_X1 U4362 ( .A(n2645), .ZN(n4303) );
  NAND2_X1 U4363 ( .A1(b_2_), .A2(a_2_), .ZN(n2645) );
  XNOR2_X1 U4364 ( .A(n4426), .B(n4427), .ZN(n4305) );
  NOR2_X1 U4365 ( .A1(n4428), .A2(n4429), .ZN(n4427) );
  INV_X1 U4366 ( .A(n4430), .ZN(n4429) );
  NOR2_X1 U4367 ( .A1(n4431), .A2(n4432), .ZN(n4428) );
  XOR2_X1 U4368 ( .A(n4433), .B(n4434), .Z(n4192) );
  NOR2_X1 U4369 ( .A1(n4435), .A2(n4436), .ZN(n4434) );
  INV_X1 U4370 ( .A(n4437), .ZN(n4436) );
  NOR2_X1 U4371 ( .A1(n4438), .A2(n4439), .ZN(n4435) );
  NAND2_X1 U4372 ( .A1(n4437), .A2(n4440), .ZN(n2739) );
  NAND2_X1 U4373 ( .A1(n4441), .A2(n4433), .ZN(n4440) );
  NAND2_X1 U4374 ( .A1(n4442), .A2(n4443), .ZN(n4433) );
  NAND2_X1 U4375 ( .A1(n4444), .A2(b_0_), .ZN(n4443) );
  NOR2_X1 U4376 ( .A1(n4445), .A2(n2695), .ZN(n4444) );
  NOR2_X1 U4377 ( .A1(n2644), .A2(n4321), .ZN(n4445) );
  NAND2_X1 U4378 ( .A1(n2644), .A2(n4321), .ZN(n4442) );
  NAND2_X1 U4379 ( .A1(n4430), .A2(n4446), .ZN(n4321) );
  NAND2_X1 U4380 ( .A1(n4447), .A2(n4426), .ZN(n4446) );
  NAND2_X1 U4381 ( .A1(n4448), .A2(n4449), .ZN(n4426) );
  NAND2_X1 U4382 ( .A1(n4450), .A2(b_1_), .ZN(n4449) );
  NOR2_X1 U4383 ( .A1(n4451), .A2(n2553), .ZN(n4450) );
  NOR2_X1 U4384 ( .A1(n4330), .A2(n4331), .ZN(n4451) );
  NAND2_X1 U4385 ( .A1(n4330), .A2(n4331), .ZN(n4448) );
  NAND2_X1 U4386 ( .A1(n4422), .A2(n4452), .ZN(n4331) );
  NAND2_X1 U4387 ( .A1(n4453), .A2(n4421), .ZN(n4452) );
  NAND2_X1 U4388 ( .A1(n4454), .A2(n4455), .ZN(n4421) );
  NAND2_X1 U4389 ( .A1(n4456), .A2(b_1_), .ZN(n4455) );
  NOR2_X1 U4390 ( .A1(n4457), .A2(n2479), .ZN(n4456) );
  NOR2_X1 U4391 ( .A1(n4341), .A2(n4342), .ZN(n4457) );
  NAND2_X1 U4392 ( .A1(n4341), .A2(n4342), .ZN(n4454) );
  NAND2_X1 U4393 ( .A1(n4416), .A2(n4458), .ZN(n4342) );
  NAND2_X1 U4394 ( .A1(n4459), .A2(n4415), .ZN(n4458) );
  NAND2_X1 U4395 ( .A1(n4460), .A2(n4461), .ZN(n4415) );
  NAND2_X1 U4396 ( .A1(n4462), .A2(b_1_), .ZN(n4461) );
  NOR2_X1 U4397 ( .A1(n4463), .A2(n2437), .ZN(n4462) );
  NOR2_X1 U4398 ( .A1(n4352), .A2(n4353), .ZN(n4463) );
  NAND2_X1 U4399 ( .A1(n4352), .A2(n4353), .ZN(n4460) );
  NAND2_X1 U4400 ( .A1(n4410), .A2(n4464), .ZN(n4353) );
  NAND2_X1 U4401 ( .A1(n4465), .A2(n4409), .ZN(n4464) );
  NAND2_X1 U4402 ( .A1(n4466), .A2(n4467), .ZN(n4409) );
  NAND2_X1 U4403 ( .A1(n4468), .A2(b_1_), .ZN(n4467) );
  NOR2_X1 U4404 ( .A1(n4469), .A2(n2383), .ZN(n4468) );
  NOR2_X1 U4405 ( .A1(n4363), .A2(n4364), .ZN(n4469) );
  NAND2_X1 U4406 ( .A1(n4363), .A2(n4364), .ZN(n4466) );
  NAND2_X1 U4407 ( .A1(n4404), .A2(n4470), .ZN(n4364) );
  NAND2_X1 U4408 ( .A1(n4471), .A2(n4403), .ZN(n4470) );
  NAND2_X1 U4409 ( .A1(n4472), .A2(n4473), .ZN(n4403) );
  NAND2_X1 U4410 ( .A1(n4474), .A2(b_1_), .ZN(n4473) );
  NOR2_X1 U4411 ( .A1(n4475), .A2(n2314), .ZN(n4474) );
  NOR2_X1 U4412 ( .A1(n4374), .A2(n4375), .ZN(n4475) );
  NAND2_X1 U4413 ( .A1(n4374), .A2(n4375), .ZN(n4472) );
  NAND2_X1 U4414 ( .A1(n4476), .A2(n4477), .ZN(n4375) );
  NAND2_X1 U4415 ( .A1(n4478), .A2(b_1_), .ZN(n4477) );
  NOR2_X1 U4416 ( .A1(n4479), .A2(n2285), .ZN(n4478) );
  NOR2_X1 U4417 ( .A1(n4400), .A2(n4401), .ZN(n4479) );
  NAND2_X1 U4418 ( .A1(n4400), .A2(n4401), .ZN(n4476) );
  NAND2_X1 U4419 ( .A1(n4397), .A2(n4480), .ZN(n4401) );
  NAND2_X1 U4420 ( .A1(n4395), .A2(n4396), .ZN(n4480) );
  NOR2_X1 U4421 ( .A1(n2696), .A2(n2271), .ZN(n4396) );
  NOR2_X1 U4422 ( .A1(n2684), .A2(n2637), .ZN(n4395) );
  NAND2_X1 U4423 ( .A1(n4481), .A2(n2685), .ZN(n4397) );
  NOR2_X1 U4424 ( .A1(n2696), .A2(n2637), .ZN(n4481) );
  NOR2_X1 U4425 ( .A1(n2637), .A2(n2271), .ZN(n4400) );
  NOR2_X1 U4426 ( .A1(n2637), .A2(n2285), .ZN(n4374) );
  NAND2_X1 U4427 ( .A1(n4407), .A2(n2687), .ZN(n4471) );
  NAND2_X1 U4428 ( .A1(n4482), .A2(n4483), .ZN(n4404) );
  INV_X1 U4429 ( .A(n4407), .ZN(n4483) );
  NAND2_X1 U4430 ( .A1(b_0_), .A2(a_11_), .ZN(n4407) );
  NOR2_X1 U4431 ( .A1(n2687), .A2(n2696), .ZN(n4482) );
  NOR2_X1 U4432 ( .A1(n2637), .A2(n2687), .ZN(n4363) );
  NAND2_X1 U4433 ( .A1(n4413), .A2(n2689), .ZN(n4465) );
  NAND2_X1 U4434 ( .A1(n4484), .A2(n4485), .ZN(n4410) );
  INV_X1 U4435 ( .A(n4413), .ZN(n4485) );
  NAND2_X1 U4436 ( .A1(b_0_), .A2(a_9_), .ZN(n4413) );
  NOR2_X1 U4437 ( .A1(n2689), .A2(n2696), .ZN(n4484) );
  NOR2_X1 U4438 ( .A1(n2637), .A2(n2689), .ZN(n4352) );
  NAND2_X1 U4439 ( .A1(n4419), .A2(n2691), .ZN(n4459) );
  NAND2_X1 U4440 ( .A1(n4486), .A2(n4487), .ZN(n4416) );
  INV_X1 U4441 ( .A(n4419), .ZN(n4487) );
  NAND2_X1 U4442 ( .A1(b_0_), .A2(a_7_), .ZN(n4419) );
  NOR2_X1 U4443 ( .A1(n2691), .A2(n2696), .ZN(n4486) );
  NOR2_X1 U4444 ( .A1(n2637), .A2(n2691), .ZN(n4341) );
  NAND2_X1 U4445 ( .A1(n4425), .A2(n2506), .ZN(n4453) );
  NAND2_X1 U4446 ( .A1(n4488), .A2(n4489), .ZN(n4422) );
  INV_X1 U4447 ( .A(n4425), .ZN(n4489) );
  NAND2_X1 U4448 ( .A1(b_0_), .A2(a_5_), .ZN(n4425) );
  NOR2_X1 U4449 ( .A1(n2506), .A2(n2696), .ZN(n4488) );
  NOR2_X1 U4450 ( .A1(n2637), .A2(n2506), .ZN(n4330) );
  OR2_X1 U4451 ( .A1(n4431), .A2(a_2_), .ZN(n4447) );
  NAND2_X1 U4452 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  NOR2_X1 U4453 ( .A1(n2637), .A2(n2553), .ZN(n4431) );
  NOR2_X1 U4454 ( .A1(n2695), .A2(n2696), .ZN(n4432) );
  NOR2_X1 U4455 ( .A1(n2696), .A2(n2609), .ZN(n2644) );
  OR2_X1 U4456 ( .A1(n4438), .A2(a_0_), .ZN(n4441) );
  NAND2_X1 U4457 ( .A1(n4439), .A2(n4438), .ZN(n4437) );
  NOR2_X1 U4458 ( .A1(n2637), .A2(n2609), .ZN(n4438) );
  NOR2_X1 U4459 ( .A1(n2623), .A2(n2696), .ZN(n4439) );
  AND2_X1 U4460 ( .A1(n4490), .A2(n4491), .ZN(n2160) );
  NAND2_X1 U4461 ( .A1(n4492), .A2(n2159), .ZN(n4491) );
  NOR2_X1 U4462 ( .A1(n4494), .A2(n4495), .ZN(n4492) );
  NOR2_X1 U4463 ( .A1(n2633), .A2(n2623), .ZN(n4495) );
  INV_X1 U4464 ( .A(n2697), .ZN(n2633) );
  NOR2_X1 U4465 ( .A1(b_0_), .A2(n4496), .ZN(n4494) );
  NOR2_X1 U4466 ( .A1(a_0_), .A2(n2697), .ZN(n4496) );
  NAND2_X1 U4467 ( .A1(n4497), .A2(n4498), .ZN(n2697) );
  NAND2_X1 U4468 ( .A1(n4499), .A2(n2696), .ZN(n4498) );
  INV_X1 U4469 ( .A(b_1_), .ZN(n2696) );
  NAND2_X1 U4470 ( .A1(n2605), .A2(n2609), .ZN(n4499) );
  INV_X1 U4471 ( .A(n2614), .ZN(n2605) );
  NAND2_X1 U4472 ( .A1(a_1_), .A2(n2614), .ZN(n4497) );
  NAND2_X1 U4473 ( .A1(n4500), .A2(n4501), .ZN(n2614) );
  NAND2_X1 U4474 ( .A1(n4502), .A2(n2581), .ZN(n4501) );
  INV_X1 U4475 ( .A(b_2_), .ZN(n2581) );
  NAND2_X1 U4476 ( .A1(n2577), .A2(n2695), .ZN(n4502) );
  INV_X1 U4477 ( .A(n2587), .ZN(n2577) );
  NAND2_X1 U4478 ( .A1(a_2_), .A2(n2587), .ZN(n4500) );
  NAND2_X1 U4479 ( .A1(n4503), .A2(n4504), .ZN(n2587) );
  NAND2_X1 U4480 ( .A1(n4505), .A2(n2694), .ZN(n4504) );
  INV_X1 U4481 ( .A(b_3_), .ZN(n2694) );
  NAND2_X1 U4482 ( .A1(n2549), .A2(n2553), .ZN(n4505) );
  INV_X1 U4483 ( .A(n2559), .ZN(n2549) );
  NAND2_X1 U4484 ( .A1(a_3_), .A2(n2559), .ZN(n4503) );
  NAND2_X1 U4485 ( .A1(n4506), .A2(n4507), .ZN(n2559) );
  NAND2_X1 U4486 ( .A1(n4508), .A2(n2693), .ZN(n4507) );
  INV_X1 U4487 ( .A(b_4_), .ZN(n2693) );
  NAND2_X1 U4488 ( .A1(n2516), .A2(n2506), .ZN(n4508) );
  INV_X1 U4489 ( .A(n2525), .ZN(n2516) );
  NAND2_X1 U4490 ( .A1(a_4_), .A2(n2525), .ZN(n4506) );
  NAND2_X1 U4491 ( .A1(n4509), .A2(n4510), .ZN(n2525) );
  NAND2_X1 U4492 ( .A1(n4511), .A2(n2692), .ZN(n4510) );
  INV_X1 U4493 ( .A(b_5_), .ZN(n2692) );
  NAND2_X1 U4494 ( .A1(n2489), .A2(n2479), .ZN(n4511) );
  INV_X1 U4495 ( .A(n2497), .ZN(n2489) );
  NAND2_X1 U4496 ( .A1(a_5_), .A2(n2497), .ZN(n4509) );
  NAND2_X1 U4497 ( .A1(n4512), .A2(n4513), .ZN(n2497) );
  NAND2_X1 U4498 ( .A1(n4514), .A2(n2464), .ZN(n4513) );
  INV_X1 U4499 ( .A(b_6_), .ZN(n2464) );
  NAND2_X1 U4500 ( .A1(n2460), .A2(n2691), .ZN(n4514) );
  INV_X1 U4501 ( .A(n2470), .ZN(n2460) );
  NAND2_X1 U4502 ( .A1(a_6_), .A2(n2470), .ZN(n4512) );
  NAND2_X1 U4503 ( .A1(n4515), .A2(n4516), .ZN(n2470) );
  NAND2_X1 U4504 ( .A1(n4517), .A2(n2690), .ZN(n4516) );
  INV_X1 U4505 ( .A(b_7_), .ZN(n2690) );
  NAND2_X1 U4506 ( .A1(n2433), .A2(n2437), .ZN(n4517) );
  INV_X1 U4507 ( .A(n2442), .ZN(n2433) );
  NAND2_X1 U4508 ( .A1(a_7_), .A2(n2442), .ZN(n4515) );
  NAND2_X1 U4509 ( .A1(n4518), .A2(n4519), .ZN(n2442) );
  NAND2_X1 U4510 ( .A1(n4520), .A2(n2410), .ZN(n4519) );
  INV_X1 U4511 ( .A(b_8_), .ZN(n2410) );
  NAND2_X1 U4512 ( .A1(n2406), .A2(n2689), .ZN(n4520) );
  INV_X1 U4513 ( .A(n2415), .ZN(n2406) );
  NAND2_X1 U4514 ( .A1(a_8_), .A2(n2415), .ZN(n4518) );
  NAND2_X1 U4515 ( .A1(n4521), .A2(n4522), .ZN(n2415) );
  NAND2_X1 U4516 ( .A1(n4523), .A2(n2688), .ZN(n4522) );
  INV_X1 U4517 ( .A(b_9_), .ZN(n2688) );
  NAND2_X1 U4518 ( .A1(n2379), .A2(n2383), .ZN(n4523) );
  INV_X1 U4519 ( .A(n2388), .ZN(n2379) );
  NAND2_X1 U4520 ( .A1(a_9_), .A2(n2388), .ZN(n4521) );
  NAND2_X1 U4521 ( .A1(n4524), .A2(n4525), .ZN(n2388) );
  NAND2_X1 U4522 ( .A1(n4526), .A2(n2355), .ZN(n4525) );
  INV_X1 U4523 ( .A(b_10_), .ZN(n2355) );
  NAND2_X1 U4524 ( .A1(n2351), .A2(n2687), .ZN(n4526) );
  INV_X1 U4525 ( .A(n2361), .ZN(n2351) );
  NAND2_X1 U4526 ( .A1(a_10_), .A2(n2361), .ZN(n4524) );
  NAND2_X1 U4527 ( .A1(n4527), .A2(n4528), .ZN(n2361) );
  NAND2_X1 U4528 ( .A1(n4529), .A2(n2328), .ZN(n4528) );
  INV_X1 U4529 ( .A(b_11_), .ZN(n2328) );
  NAND2_X1 U4530 ( .A1(n2324), .A2(n2314), .ZN(n4529) );
  INV_X1 U4531 ( .A(n2333), .ZN(n2324) );
  NAND2_X1 U4532 ( .A1(a_11_), .A2(n2333), .ZN(n4527) );
  NAND2_X1 U4533 ( .A1(n4530), .A2(n4531), .ZN(n2333) );
  NAND2_X1 U4534 ( .A1(n4532), .A2(n2299), .ZN(n4531) );
  INV_X1 U4535 ( .A(b_12_), .ZN(n2299) );
  NAND2_X1 U4536 ( .A1(n2295), .A2(n2285), .ZN(n4532) );
  INV_X1 U4537 ( .A(n2305), .ZN(n2295) );
  NAND2_X1 U4538 ( .A1(a_12_), .A2(n2305), .ZN(n4530) );
  NAND2_X1 U4539 ( .A1(n4533), .A2(n4534), .ZN(n2305) );
  NAND2_X1 U4540 ( .A1(n4535), .A2(n2686), .ZN(n4534) );
  INV_X1 U4541 ( .A(b_13_), .ZN(n2686) );
  NAND2_X1 U4542 ( .A1(n2267), .A2(n2271), .ZN(n4535) );
  INV_X1 U4543 ( .A(n2276), .ZN(n2267) );
  NAND2_X1 U4544 ( .A1(a_13_), .A2(n2276), .ZN(n4533) );
  NAND2_X1 U4545 ( .A1(n2223), .A2(n4536), .ZN(n2276) );
  NAND2_X1 U4546 ( .A1(n2244), .A2(n2213), .ZN(n4536) );
  NAND2_X1 U4547 ( .A1(b_15_), .A2(n4392), .ZN(n2213) );
  INV_X1 U4548 ( .A(a_15_), .ZN(n4392) );
  NAND2_X1 U4549 ( .A1(n4537), .A2(n2211), .ZN(n4490) );
  INV_X1 U4550 ( .A(n2237), .ZN(n2211) );
  INV_X1 U4551 ( .A(operation_1_), .ZN(n4493) );
  NOR2_X1 U4552 ( .A1(n4538), .A2(n4539), .ZN(n4537) );
  NOR2_X1 U4553 ( .A1(a_0_), .A2(n2698), .ZN(n4539) );
  INV_X1 U4554 ( .A(n2634), .ZN(n2698) );
  NOR2_X1 U4555 ( .A1(n4540), .A2(n2637), .ZN(n4538) );
  INV_X1 U4556 ( .A(b_0_), .ZN(n2637) );
  NOR2_X1 U4557 ( .A1(n2623), .A2(n2634), .ZN(n4540) );
  NAND2_X1 U4558 ( .A1(n4541), .A2(n4542), .ZN(n2634) );
  NAND2_X1 U4559 ( .A1(b_1_), .A2(n4543), .ZN(n4542) );
  NAND2_X1 U4560 ( .A1(n2615), .A2(a_1_), .ZN(n4543) );
  INV_X1 U4561 ( .A(n2606), .ZN(n2615) );
  NAND2_X1 U4562 ( .A1(n2606), .A2(n2609), .ZN(n4541) );
  INV_X1 U4563 ( .A(a_1_), .ZN(n2609) );
  NAND2_X1 U4564 ( .A1(n4544), .A2(n4545), .ZN(n2606) );
  NAND2_X1 U4565 ( .A1(b_2_), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U4566 ( .A1(n2588), .A2(a_2_), .ZN(n4546) );
  INV_X1 U4567 ( .A(n2578), .ZN(n2588) );
  NAND2_X1 U4568 ( .A1(n2578), .A2(n2695), .ZN(n4544) );
  INV_X1 U4569 ( .A(a_2_), .ZN(n2695) );
  NAND2_X1 U4570 ( .A1(n4547), .A2(n4548), .ZN(n2578) );
  NAND2_X1 U4571 ( .A1(b_3_), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U4572 ( .A1(n2560), .A2(a_3_), .ZN(n4549) );
  INV_X1 U4573 ( .A(n2550), .ZN(n2560) );
  NAND2_X1 U4574 ( .A1(n2550), .A2(n2553), .ZN(n4547) );
  INV_X1 U4575 ( .A(a_3_), .ZN(n2553) );
  NAND2_X1 U4576 ( .A1(n4550), .A2(n4551), .ZN(n2550) );
  NAND2_X1 U4577 ( .A1(b_4_), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U4578 ( .A1(n2526), .A2(a_4_), .ZN(n4552) );
  INV_X1 U4579 ( .A(n2517), .ZN(n2526) );
  NAND2_X1 U4580 ( .A1(n2517), .A2(n2506), .ZN(n4550) );
  INV_X1 U4581 ( .A(a_4_), .ZN(n2506) );
  NAND2_X1 U4582 ( .A1(n4553), .A2(n4554), .ZN(n2517) );
  NAND2_X1 U4583 ( .A1(b_5_), .A2(n4555), .ZN(n4554) );
  NAND2_X1 U4584 ( .A1(n2498), .A2(a_5_), .ZN(n4555) );
  INV_X1 U4585 ( .A(n2490), .ZN(n2498) );
  NAND2_X1 U4586 ( .A1(n2490), .A2(n2479), .ZN(n4553) );
  INV_X1 U4587 ( .A(a_5_), .ZN(n2479) );
  NAND2_X1 U4588 ( .A1(n4556), .A2(n4557), .ZN(n2490) );
  NAND2_X1 U4589 ( .A1(b_6_), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U4590 ( .A1(n2471), .A2(a_6_), .ZN(n4558) );
  INV_X1 U4591 ( .A(n2461), .ZN(n2471) );
  NAND2_X1 U4592 ( .A1(n2461), .A2(n2691), .ZN(n4556) );
  INV_X1 U4593 ( .A(a_6_), .ZN(n2691) );
  NAND2_X1 U4594 ( .A1(n4559), .A2(n4560), .ZN(n2461) );
  NAND2_X1 U4595 ( .A1(b_7_), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U4596 ( .A1(n2443), .A2(a_7_), .ZN(n4561) );
  INV_X1 U4597 ( .A(n2434), .ZN(n2443) );
  NAND2_X1 U4598 ( .A1(n2434), .A2(n2437), .ZN(n4559) );
  INV_X1 U4599 ( .A(a_7_), .ZN(n2437) );
  NAND2_X1 U4600 ( .A1(n4562), .A2(n4563), .ZN(n2434) );
  NAND2_X1 U4601 ( .A1(b_8_), .A2(n4564), .ZN(n4563) );
  NAND2_X1 U4602 ( .A1(n2416), .A2(a_8_), .ZN(n4564) );
  INV_X1 U4603 ( .A(n2407), .ZN(n2416) );
  NAND2_X1 U4604 ( .A1(n2407), .A2(n2689), .ZN(n4562) );
  INV_X1 U4605 ( .A(a_8_), .ZN(n2689) );
  NAND2_X1 U4606 ( .A1(n4565), .A2(n4566), .ZN(n2407) );
  NAND2_X1 U4607 ( .A1(b_9_), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U4608 ( .A1(n2389), .A2(a_9_), .ZN(n4567) );
  INV_X1 U4609 ( .A(n2380), .ZN(n2389) );
  NAND2_X1 U4610 ( .A1(n2380), .A2(n2383), .ZN(n4565) );
  INV_X1 U4611 ( .A(a_9_), .ZN(n2383) );
  NAND2_X1 U4612 ( .A1(n4568), .A2(n4569), .ZN(n2380) );
  NAND2_X1 U4613 ( .A1(b_10_), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U4614 ( .A1(n2362), .A2(a_10_), .ZN(n4570) );
  INV_X1 U4615 ( .A(n2352), .ZN(n2362) );
  NAND2_X1 U4616 ( .A1(n2352), .A2(n2687), .ZN(n4568) );
  INV_X1 U4617 ( .A(a_10_), .ZN(n2687) );
  NAND2_X1 U4618 ( .A1(n4571), .A2(n4572), .ZN(n2352) );
  NAND2_X1 U4619 ( .A1(b_11_), .A2(n4573), .ZN(n4572) );
  NAND2_X1 U4620 ( .A1(n2334), .A2(a_11_), .ZN(n4573) );
  INV_X1 U4621 ( .A(n2325), .ZN(n2334) );
  NAND2_X1 U4622 ( .A1(n2325), .A2(n2314), .ZN(n4571) );
  INV_X1 U4623 ( .A(a_11_), .ZN(n2314) );
  NAND2_X1 U4624 ( .A1(n4574), .A2(n4575), .ZN(n2325) );
  NAND2_X1 U4625 ( .A1(b_12_), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U4626 ( .A1(n2306), .A2(a_12_), .ZN(n4576) );
  INV_X1 U4627 ( .A(n2296), .ZN(n2306) );
  NAND2_X1 U4628 ( .A1(n2296), .A2(n2285), .ZN(n4574) );
  INV_X1 U4629 ( .A(a_12_), .ZN(n2285) );
  NAND2_X1 U4630 ( .A1(n4577), .A2(n4578), .ZN(n2296) );
  NAND2_X1 U4631 ( .A1(b_13_), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U4632 ( .A1(n2277), .A2(a_13_), .ZN(n4579) );
  INV_X1 U4633 ( .A(n2268), .ZN(n2277) );
  NAND2_X1 U4634 ( .A1(n2268), .A2(n2271), .ZN(n4577) );
  INV_X1 U4635 ( .A(a_13_), .ZN(n2271) );
  NAND2_X1 U4636 ( .A1(n2244), .A2(n4580), .ZN(n2268) );
  NAND2_X1 U4637 ( .A1(n2212), .A2(n2223), .ZN(n4580) );
  NAND2_X1 U4638 ( .A1(a_14_), .A2(n2225), .ZN(n2223) );
  INV_X1 U4639 ( .A(b_14_), .ZN(n2225) );
  NAND2_X1 U4640 ( .A1(a_15_), .A2(n2222), .ZN(n2212) );
  INV_X1 U4641 ( .A(b_15_), .ZN(n2222) );
  NAND2_X1 U4642 ( .A1(b_14_), .A2(n2684), .ZN(n2244) );
  INV_X1 U4643 ( .A(a_14_), .ZN(n2684) );
  INV_X1 U4644 ( .A(a_0_), .ZN(n2623) );
endmodule

