module add_mul_mix_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, 
        c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_,
         c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919;

  XOR2_X2 U457 ( .A(n900), .B(n901), .Z(n449) );
  XNOR2_X1 U458 ( .A(n441), .B(n442), .ZN(Result_9_) );
  XNOR2_X1 U459 ( .A(n443), .B(n444), .ZN(n442) );
  XNOR2_X1 U460 ( .A(n445), .B(n446), .ZN(Result_8_) );
  XOR2_X1 U461 ( .A(n447), .B(n448), .Z(n446) );
  NAND2_X1 U462 ( .A1(n449), .A2(n450), .ZN(n448) );
  XOR2_X1 U463 ( .A(n451), .B(n452), .Z(Result_7_) );
  NOR2_X1 U464 ( .A1(n453), .A2(n454), .ZN(Result_6_) );
  NOR2_X1 U465 ( .A1(n455), .A2(n456), .ZN(n454) );
  AND2_X1 U466 ( .A1(n452), .A2(n451), .ZN(n455) );
  XNOR2_X1 U467 ( .A(n453), .B(n457), .ZN(Result_5_) );
  NAND2_X1 U468 ( .A1(n458), .A2(n459), .ZN(n457) );
  NAND2_X1 U469 ( .A1(n460), .A2(n461), .ZN(n459) );
  NAND2_X1 U470 ( .A1(n462), .A2(n463), .ZN(n460) );
  XOR2_X1 U471 ( .A(n464), .B(n465), .Z(Result_4_) );
  XOR2_X1 U472 ( .A(n466), .B(n467), .Z(Result_3_) );
  AND2_X1 U473 ( .A1(n468), .A2(n469), .ZN(n467) );
  XOR2_X1 U474 ( .A(n470), .B(n471), .Z(Result_2_) );
  AND2_X1 U475 ( .A1(n472), .A2(n473), .ZN(n471) );
  XOR2_X1 U476 ( .A(n474), .B(n475), .Z(Result_1_) );
  NOR2_X1 U477 ( .A1(n476), .A2(n477), .ZN(n475) );
  INV_X1 U478 ( .A(n478), .ZN(n477) );
  NOR2_X1 U479 ( .A1(n479), .A2(n480), .ZN(n476) );
  XOR2_X1 U480 ( .A(n481), .B(n482), .Z(Result_14_) );
  NOR2_X1 U481 ( .A1(n483), .A2(n484), .ZN(n482) );
  XOR2_X1 U482 ( .A(n485), .B(n486), .Z(Result_13_) );
  XOR2_X1 U483 ( .A(n487), .B(n488), .Z(n486) );
  NOR2_X1 U484 ( .A1(n484), .A2(n489), .ZN(n488) );
  XNOR2_X1 U485 ( .A(n490), .B(n491), .ZN(Result_12_) );
  XNOR2_X1 U486 ( .A(n492), .B(n493), .ZN(n491) );
  XOR2_X1 U487 ( .A(n494), .B(n495), .Z(Result_11_) );
  NOR2_X1 U488 ( .A1(n496), .A2(n497), .ZN(n495) );
  NOR2_X1 U489 ( .A1(n498), .A2(n499), .ZN(n496) );
  NOR2_X1 U490 ( .A1(n484), .A2(n500), .ZN(n498) );
  XNOR2_X1 U491 ( .A(n501), .B(n502), .ZN(Result_10_) );
  XNOR2_X1 U492 ( .A(n503), .B(n504), .ZN(n502) );
  NAND3_X1 U493 ( .A1(n505), .A2(n480), .A3(n506), .ZN(Result_0_) );
  NAND2_X1 U494 ( .A1(n449), .A2(n479), .ZN(n506) );
  NAND3_X1 U495 ( .A1(n449), .A2(n507), .A3(n508), .ZN(n480) );
  NAND2_X1 U496 ( .A1(n478), .A2(n474), .ZN(n505) );
  NAND2_X1 U497 ( .A1(n473), .A2(n509), .ZN(n474) );
  NAND2_X1 U498 ( .A1(n472), .A2(n470), .ZN(n509) );
  NAND2_X1 U499 ( .A1(n469), .A2(n510), .ZN(n470) );
  NAND2_X1 U500 ( .A1(n466), .A2(n468), .ZN(n510) );
  NAND2_X1 U501 ( .A1(n511), .A2(n512), .ZN(n468) );
  NAND2_X1 U502 ( .A1(n513), .A2(n514), .ZN(n512) );
  XOR2_X1 U503 ( .A(n515), .B(n516), .Z(n511) );
  AND2_X1 U504 ( .A1(n464), .A2(n465), .ZN(n466) );
  NAND3_X1 U505 ( .A1(n517), .A2(n458), .A3(n518), .ZN(n465) );
  NAND2_X1 U506 ( .A1(n453), .A2(n519), .ZN(n518) );
  AND3_X1 U507 ( .A1(n451), .A2(n452), .A3(n456), .ZN(n453) );
  XOR2_X1 U508 ( .A(n463), .B(n462), .Z(n456) );
  NAND2_X1 U509 ( .A1(n520), .A2(n521), .ZN(n452) );
  NAND3_X1 U510 ( .A1(n450), .A2(n522), .A3(n449), .ZN(n521) );
  OR2_X1 U511 ( .A1(n447), .A2(n445), .ZN(n522) );
  NAND2_X1 U512 ( .A1(n445), .A2(n447), .ZN(n520) );
  NAND2_X1 U513 ( .A1(n523), .A2(n524), .ZN(n447) );
  NAND2_X1 U514 ( .A1(n444), .A2(n525), .ZN(n524) );
  NAND2_X1 U515 ( .A1(n443), .A2(n441), .ZN(n525) );
  NOR2_X1 U516 ( .A1(n526), .A2(n484), .ZN(n444) );
  OR2_X1 U517 ( .A1(n441), .A2(n443), .ZN(n523) );
  AND2_X1 U518 ( .A1(n527), .A2(n528), .ZN(n443) );
  NAND2_X1 U519 ( .A1(n504), .A2(n529), .ZN(n528) );
  NAND2_X1 U520 ( .A1(n503), .A2(n501), .ZN(n529) );
  NOR2_X1 U521 ( .A1(n530), .A2(n484), .ZN(n504) );
  OR2_X1 U522 ( .A1(n501), .A2(n503), .ZN(n527) );
  NOR2_X1 U523 ( .A1(n497), .A2(n531), .ZN(n503) );
  AND2_X1 U524 ( .A1(n494), .A2(n532), .ZN(n531) );
  NAND2_X1 U525 ( .A1(n533), .A2(n534), .ZN(n532) );
  NAND2_X1 U526 ( .A1(n535), .A2(n450), .ZN(n534) );
  XOR2_X1 U527 ( .A(n536), .B(n537), .Z(n494) );
  XOR2_X1 U528 ( .A(n538), .B(n539), .Z(n536) );
  NOR2_X1 U529 ( .A1(n500), .A2(n533), .ZN(n497) );
  INV_X1 U530 ( .A(n499), .ZN(n533) );
  NAND2_X1 U531 ( .A1(n540), .A2(n541), .ZN(n499) );
  NAND2_X1 U532 ( .A1(n493), .A2(n542), .ZN(n541) );
  OR2_X1 U533 ( .A1(n492), .A2(n490), .ZN(n542) );
  NOR2_X1 U534 ( .A1(n543), .A2(n484), .ZN(n493) );
  NAND2_X1 U535 ( .A1(n490), .A2(n492), .ZN(n540) );
  NAND2_X1 U536 ( .A1(n544), .A2(n545), .ZN(n492) );
  NAND3_X1 U537 ( .A1(n450), .A2(n546), .A3(n547), .ZN(n545) );
  NAND2_X1 U538 ( .A1(n485), .A2(n487), .ZN(n546) );
  INV_X1 U539 ( .A(n484), .ZN(n450) );
  OR2_X1 U540 ( .A1(n487), .A2(n485), .ZN(n544) );
  XNOR2_X1 U541 ( .A(n548), .B(n549), .ZN(n485) );
  NOR2_X1 U542 ( .A1(n550), .A2(n551), .ZN(n549) );
  NAND2_X1 U543 ( .A1(Result_15_), .A2(n548), .ZN(n487) );
  NOR2_X1 U544 ( .A1(n552), .A2(n483), .ZN(n548) );
  NOR2_X1 U545 ( .A1(n484), .A2(n550), .ZN(Result_15_) );
  XNOR2_X1 U546 ( .A(c_7_), .B(d_7_), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n553), .B(n554), .ZN(n490) );
  XOR2_X1 U548 ( .A(n555), .B(n556), .Z(n554) );
  NAND2_X1 U549 ( .A1(n547), .A2(n557), .ZN(n556) );
  XNOR2_X1 U550 ( .A(n558), .B(n559), .ZN(n501) );
  XOR2_X1 U551 ( .A(n560), .B(n561), .Z(n558) );
  NOR2_X1 U552 ( .A1(n552), .A2(n500), .ZN(n561) );
  XNOR2_X1 U553 ( .A(n562), .B(n563), .ZN(n441) );
  XOR2_X1 U554 ( .A(n564), .B(n565), .Z(n562) );
  NOR2_X1 U555 ( .A1(n552), .A2(n530), .ZN(n565) );
  XNOR2_X1 U556 ( .A(n566), .B(n567), .ZN(n445) );
  XOR2_X1 U557 ( .A(n568), .B(n569), .Z(n567) );
  NAND2_X1 U558 ( .A1(n570), .A2(n557), .ZN(n569) );
  XOR2_X1 U559 ( .A(n571), .B(n572), .Z(n451) );
  XOR2_X1 U560 ( .A(n573), .B(n574), .Z(n571) );
  NOR2_X1 U561 ( .A1(n552), .A2(n575), .ZN(n574) );
  NAND3_X1 U562 ( .A1(n462), .A2(n463), .A3(n519), .ZN(n458) );
  INV_X1 U563 ( .A(n461), .ZN(n519) );
  NAND2_X1 U564 ( .A1(n517), .A2(n576), .ZN(n461) );
  OR2_X1 U565 ( .A1(n577), .A2(n578), .ZN(n576) );
  NAND2_X1 U566 ( .A1(n579), .A2(n580), .ZN(n463) );
  NAND3_X1 U567 ( .A1(n557), .A2(n581), .A3(n449), .ZN(n580) );
  OR2_X1 U568 ( .A1(n573), .A2(n572), .ZN(n581) );
  NAND2_X1 U569 ( .A1(n572), .A2(n573), .ZN(n579) );
  NAND2_X1 U570 ( .A1(n582), .A2(n583), .ZN(n573) );
  NAND3_X1 U571 ( .A1(n557), .A2(n584), .A3(n570), .ZN(n583) );
  OR2_X1 U572 ( .A1(n566), .A2(n568), .ZN(n584) );
  NAND2_X1 U573 ( .A1(n566), .A2(n568), .ZN(n582) );
  NAND2_X1 U574 ( .A1(n585), .A2(n586), .ZN(n568) );
  NAND3_X1 U575 ( .A1(n557), .A2(n587), .A3(n588), .ZN(n586) );
  OR2_X1 U576 ( .A1(n563), .A2(n564), .ZN(n587) );
  NAND2_X1 U577 ( .A1(n563), .A2(n564), .ZN(n585) );
  NAND2_X1 U578 ( .A1(n589), .A2(n590), .ZN(n564) );
  NAND3_X1 U579 ( .A1(n557), .A2(n591), .A3(n535), .ZN(n590) );
  OR2_X1 U580 ( .A1(n560), .A2(n559), .ZN(n591) );
  NAND2_X1 U581 ( .A1(n559), .A2(n560), .ZN(n589) );
  NAND2_X1 U582 ( .A1(n592), .A2(n593), .ZN(n560) );
  NAND2_X1 U583 ( .A1(n539), .A2(n594), .ZN(n593) );
  OR2_X1 U584 ( .A1(n538), .A2(n537), .ZN(n594) );
  NOR2_X1 U585 ( .A1(n543), .A2(n552), .ZN(n539) );
  NAND2_X1 U586 ( .A1(n537), .A2(n538), .ZN(n592) );
  NAND2_X1 U587 ( .A1(n595), .A2(n596), .ZN(n538) );
  NAND3_X1 U588 ( .A1(n557), .A2(n597), .A3(n547), .ZN(n596) );
  NAND2_X1 U589 ( .A1(n553), .A2(n555), .ZN(n597) );
  INV_X1 U590 ( .A(n552), .ZN(n557) );
  OR2_X1 U591 ( .A1(n555), .A2(n553), .ZN(n595) );
  XNOR2_X1 U592 ( .A(n598), .B(n599), .ZN(n553) );
  NAND2_X1 U593 ( .A1(n481), .A2(n598), .ZN(n555) );
  NOR2_X1 U594 ( .A1(n552), .A2(n550), .ZN(n481) );
  XOR2_X1 U595 ( .A(n600), .B(n601), .Z(n552) );
  XOR2_X1 U596 ( .A(d_6_), .B(c_6_), .Z(n601) );
  NAND2_X1 U597 ( .A1(d_7_), .A2(c_7_), .ZN(n600) );
  XNOR2_X1 U598 ( .A(n602), .B(n603), .ZN(n537) );
  XOR2_X1 U599 ( .A(n604), .B(n605), .Z(n603) );
  NAND2_X1 U600 ( .A1(n606), .A2(n547), .ZN(n602) );
  XNOR2_X1 U601 ( .A(n607), .B(n608), .ZN(n559) );
  NAND2_X1 U602 ( .A1(n609), .A2(n610), .ZN(n607) );
  XOR2_X1 U603 ( .A(n611), .B(n612), .Z(n563) );
  XOR2_X1 U604 ( .A(n613), .B(n614), .Z(n611) );
  NOR2_X1 U605 ( .A1(n551), .A2(n500), .ZN(n614) );
  XOR2_X1 U606 ( .A(n615), .B(n616), .Z(n566) );
  XOR2_X1 U607 ( .A(n617), .B(n618), .Z(n615) );
  NOR2_X1 U608 ( .A1(n551), .A2(n530), .ZN(n618) );
  XNOR2_X1 U609 ( .A(n619), .B(n620), .ZN(n572) );
  XOR2_X1 U610 ( .A(n621), .B(n622), .Z(n620) );
  NAND2_X1 U611 ( .A1(n570), .A2(n606), .ZN(n622) );
  XNOR2_X1 U612 ( .A(n623), .B(n624), .ZN(n462) );
  XOR2_X1 U613 ( .A(n625), .B(n626), .Z(n624) );
  NAND2_X1 U614 ( .A1(n449), .A2(n606), .ZN(n626) );
  NAND2_X1 U615 ( .A1(n578), .A2(n577), .ZN(n517) );
  NAND2_X1 U616 ( .A1(n627), .A2(n628), .ZN(n577) );
  NAND3_X1 U617 ( .A1(n606), .A2(n629), .A3(n449), .ZN(n628) );
  OR2_X1 U618 ( .A1(n623), .A2(n625), .ZN(n629) );
  NAND2_X1 U619 ( .A1(n623), .A2(n625), .ZN(n627) );
  NAND2_X1 U620 ( .A1(n630), .A2(n631), .ZN(n625) );
  NAND3_X1 U621 ( .A1(n606), .A2(n632), .A3(n570), .ZN(n631) );
  OR2_X1 U622 ( .A1(n619), .A2(n621), .ZN(n632) );
  NAND2_X1 U623 ( .A1(n619), .A2(n621), .ZN(n630) );
  NAND2_X1 U624 ( .A1(n633), .A2(n634), .ZN(n621) );
  NAND3_X1 U625 ( .A1(n606), .A2(n635), .A3(n588), .ZN(n634) );
  OR2_X1 U626 ( .A1(n617), .A2(n616), .ZN(n635) );
  NAND2_X1 U627 ( .A1(n616), .A2(n617), .ZN(n633) );
  NAND2_X1 U628 ( .A1(n636), .A2(n637), .ZN(n617) );
  NAND3_X1 U629 ( .A1(n606), .A2(n638), .A3(n535), .ZN(n637) );
  OR2_X1 U630 ( .A1(n613), .A2(n612), .ZN(n638) );
  NAND2_X1 U631 ( .A1(n612), .A2(n613), .ZN(n636) );
  NAND2_X1 U632 ( .A1(n609), .A2(n639), .ZN(n613) );
  NAND2_X1 U633 ( .A1(n608), .A2(n610), .ZN(n639) );
  NAND2_X1 U634 ( .A1(n640), .A2(n641), .ZN(n610) );
  NAND2_X1 U635 ( .A1(n606), .A2(n642), .ZN(n641) );
  INV_X1 U636 ( .A(n643), .ZN(n640) );
  XNOR2_X1 U637 ( .A(n644), .B(n645), .ZN(n608) );
  XOR2_X1 U638 ( .A(n646), .B(n647), .Z(n644) );
  NOR2_X1 U639 ( .A1(n489), .A2(n648), .ZN(n647) );
  NAND2_X1 U640 ( .A1(n642), .A2(n643), .ZN(n609) );
  NAND2_X1 U641 ( .A1(n649), .A2(n650), .ZN(n643) );
  NAND3_X1 U642 ( .A1(n547), .A2(n651), .A3(n606), .ZN(n650) );
  NAND2_X1 U643 ( .A1(n604), .A2(n605), .ZN(n651) );
  OR2_X1 U644 ( .A1(n604), .A2(n605), .ZN(n649) );
  NAND2_X1 U645 ( .A1(n646), .A2(n652), .ZN(n605) );
  NAND2_X1 U646 ( .A1(n653), .A2(n654), .ZN(n652) );
  NAND2_X1 U647 ( .A1(n655), .A2(n656), .ZN(n654) );
  NAND2_X1 U648 ( .A1(n657), .A2(n658), .ZN(n653) );
  NAND2_X1 U649 ( .A1(n598), .A2(n599), .ZN(n604) );
  NOR2_X1 U650 ( .A1(n551), .A2(n483), .ZN(n598) );
  INV_X1 U651 ( .A(n606), .ZN(n551) );
  XOR2_X1 U652 ( .A(n659), .B(n660), .Z(n606) );
  XOR2_X1 U653 ( .A(d_5_), .B(c_5_), .Z(n660) );
  XNOR2_X1 U654 ( .A(n661), .B(n662), .ZN(n612) );
  XOR2_X1 U655 ( .A(n663), .B(n664), .Z(n661) );
  XOR2_X1 U656 ( .A(n665), .B(n666), .Z(n616) );
  XNOR2_X1 U657 ( .A(n667), .B(n668), .ZN(n665) );
  XOR2_X1 U658 ( .A(n669), .B(n670), .Z(n619) );
  NOR2_X1 U659 ( .A1(n671), .A2(n672), .ZN(n670) );
  NOR2_X1 U660 ( .A1(n673), .A2(n674), .ZN(n671) );
  NOR2_X1 U661 ( .A1(n648), .A2(n530), .ZN(n674) );
  INV_X1 U662 ( .A(n675), .ZN(n673) );
  XOR2_X1 U663 ( .A(n676), .B(n677), .Z(n623) );
  XNOR2_X1 U664 ( .A(n678), .B(n679), .ZN(n677) );
  NAND2_X1 U665 ( .A1(n570), .A2(n657), .ZN(n679) );
  XOR2_X1 U666 ( .A(n680), .B(n681), .Z(n578) );
  XOR2_X1 U667 ( .A(n682), .B(n683), .Z(n680) );
  NOR2_X1 U668 ( .A1(n648), .A2(n575), .ZN(n683) );
  XOR2_X1 U669 ( .A(n514), .B(n513), .Z(n464) );
  NAND3_X1 U670 ( .A1(n513), .A2(n514), .A3(n684), .ZN(n469) );
  XOR2_X1 U671 ( .A(n516), .B(n685), .Z(n684) );
  NAND2_X1 U672 ( .A1(n686), .A2(n687), .ZN(n514) );
  NAND3_X1 U673 ( .A1(n657), .A2(n688), .A3(n449), .ZN(n687) );
  OR2_X1 U674 ( .A1(n682), .A2(n681), .ZN(n688) );
  NAND2_X1 U675 ( .A1(n681), .A2(n682), .ZN(n686) );
  NAND2_X1 U676 ( .A1(n689), .A2(n690), .ZN(n682) );
  NAND3_X1 U677 ( .A1(n657), .A2(n691), .A3(n570), .ZN(n690) );
  NAND2_X1 U678 ( .A1(n678), .A2(n676), .ZN(n691) );
  OR2_X1 U679 ( .A1(n676), .A2(n678), .ZN(n689) );
  NOR2_X1 U680 ( .A1(n672), .A2(n692), .ZN(n678) );
  AND2_X1 U681 ( .A1(n669), .A2(n693), .ZN(n692) );
  NAND2_X1 U682 ( .A1(n675), .A2(n694), .ZN(n693) );
  NAND2_X1 U683 ( .A1(n588), .A2(n657), .ZN(n694) );
  XOR2_X1 U684 ( .A(n695), .B(n696), .Z(n669) );
  XNOR2_X1 U685 ( .A(n697), .B(n698), .ZN(n696) );
  NOR2_X1 U686 ( .A1(n675), .A2(n530), .ZN(n672) );
  NAND2_X1 U687 ( .A1(n699), .A2(n700), .ZN(n675) );
  NAND2_X1 U688 ( .A1(n666), .A2(n701), .ZN(n700) );
  NAND2_X1 U689 ( .A1(n668), .A2(n667), .ZN(n701) );
  XNOR2_X1 U690 ( .A(n702), .B(n703), .ZN(n666) );
  XOR2_X1 U691 ( .A(n704), .B(n705), .Z(n702) );
  NOR2_X1 U692 ( .A1(n706), .A2(n543), .ZN(n705) );
  OR2_X1 U693 ( .A1(n668), .A2(n667), .ZN(n699) );
  AND2_X1 U694 ( .A1(n707), .A2(n708), .ZN(n667) );
  NAND2_X1 U695 ( .A1(n662), .A2(n709), .ZN(n708) );
  NAND2_X1 U696 ( .A1(n664), .A2(n663), .ZN(n709) );
  XOR2_X1 U697 ( .A(n710), .B(n711), .Z(n662) );
  XOR2_X1 U698 ( .A(n712), .B(n713), .Z(n711) );
  NAND2_X1 U699 ( .A1(n655), .A2(n547), .ZN(n710) );
  OR2_X1 U700 ( .A1(n663), .A2(n664), .ZN(n707) );
  NOR2_X1 U701 ( .A1(n543), .A2(n648), .ZN(n664) );
  NAND2_X1 U702 ( .A1(n714), .A2(n715), .ZN(n663) );
  NAND3_X1 U703 ( .A1(n547), .A2(n716), .A3(n657), .ZN(n715) );
  OR2_X1 U704 ( .A1(n645), .A2(n717), .ZN(n716) );
  NAND2_X1 U705 ( .A1(n717), .A2(n645), .ZN(n714) );
  XOR2_X1 U706 ( .A(n718), .B(n719), .Z(n645) );
  NOR2_X1 U707 ( .A1(n550), .A2(n720), .ZN(n719) );
  INV_X1 U708 ( .A(n646), .ZN(n717) );
  NAND2_X1 U709 ( .A1(n599), .A2(n718), .ZN(n646) );
  NOR2_X1 U710 ( .A1(n648), .A2(n550), .ZN(n599) );
  NOR2_X1 U711 ( .A1(n500), .A2(n648), .ZN(n668) );
  INV_X1 U712 ( .A(n657), .ZN(n648) );
  XOR2_X1 U713 ( .A(n721), .B(n722), .Z(n657) );
  XOR2_X1 U714 ( .A(d_4_), .B(c_4_), .Z(n722) );
  XNOR2_X1 U715 ( .A(n723), .B(n724), .ZN(n676) );
  NOR2_X1 U716 ( .A1(n725), .A2(n726), .ZN(n724) );
  NOR2_X1 U717 ( .A1(n727), .A2(n728), .ZN(n725) );
  NOR2_X1 U718 ( .A1(n706), .A2(n530), .ZN(n728) );
  INV_X1 U719 ( .A(n729), .ZN(n727) );
  XNOR2_X1 U720 ( .A(n730), .B(n731), .ZN(n681) );
  XOR2_X1 U721 ( .A(n732), .B(n733), .Z(n731) );
  XOR2_X1 U722 ( .A(n734), .B(n735), .Z(n513) );
  NOR2_X1 U723 ( .A1(n736), .A2(n737), .ZN(n735) );
  NOR2_X1 U724 ( .A1(n738), .A2(n739), .ZN(n736) );
  NOR2_X1 U725 ( .A1(n706), .A2(n575), .ZN(n739) );
  INV_X1 U726 ( .A(n740), .ZN(n738) );
  NAND2_X1 U727 ( .A1(n741), .A2(n742), .ZN(n472) );
  NAND2_X1 U728 ( .A1(n743), .A2(n515), .ZN(n742) );
  XNOR2_X1 U729 ( .A(n744), .B(n745), .ZN(n741) );
  NAND4_X1 U730 ( .A1(n743), .A2(n746), .A3(n515), .A4(n747), .ZN(n473) );
  INV_X1 U731 ( .A(n685), .ZN(n515) );
  NOR2_X1 U732 ( .A1(n737), .A2(n748), .ZN(n685) );
  AND2_X1 U733 ( .A1(n734), .A2(n749), .ZN(n748) );
  NAND2_X1 U734 ( .A1(n740), .A2(n750), .ZN(n749) );
  NAND2_X1 U735 ( .A1(n449), .A2(n655), .ZN(n750) );
  XNOR2_X1 U736 ( .A(n751), .B(n752), .ZN(n734) );
  NAND2_X1 U737 ( .A1(n753), .A2(n754), .ZN(n751) );
  NOR2_X1 U738 ( .A1(n740), .A2(n575), .ZN(n737) );
  NAND2_X1 U739 ( .A1(n755), .A2(n756), .ZN(n740) );
  NAND2_X1 U740 ( .A1(n732), .A2(n757), .ZN(n756) );
  NAND2_X1 U741 ( .A1(n733), .A2(n730), .ZN(n757) );
  NOR2_X1 U742 ( .A1(n726), .A2(n758), .ZN(n732) );
  AND2_X1 U743 ( .A1(n723), .A2(n759), .ZN(n758) );
  NAND2_X1 U744 ( .A1(n729), .A2(n760), .ZN(n759) );
  NAND2_X1 U745 ( .A1(n588), .A2(n655), .ZN(n760) );
  XNOR2_X1 U746 ( .A(n761), .B(n762), .ZN(n723) );
  NAND2_X1 U747 ( .A1(n763), .A2(n764), .ZN(n761) );
  NOR2_X1 U748 ( .A1(n729), .A2(n530), .ZN(n726) );
  NAND2_X1 U749 ( .A1(n765), .A2(n766), .ZN(n729) );
  NAND2_X1 U750 ( .A1(n697), .A2(n767), .ZN(n766) );
  OR2_X1 U751 ( .A1(n695), .A2(n698), .ZN(n767) );
  AND2_X1 U752 ( .A1(n768), .A2(n769), .ZN(n697) );
  NAND3_X1 U753 ( .A1(n655), .A2(n770), .A3(n642), .ZN(n769) );
  OR2_X1 U754 ( .A1(n703), .A2(n704), .ZN(n770) );
  NAND2_X1 U755 ( .A1(n703), .A2(n704), .ZN(n768) );
  NAND2_X1 U756 ( .A1(n771), .A2(n772), .ZN(n704) );
  NAND3_X1 U757 ( .A1(n547), .A2(n773), .A3(n655), .ZN(n772) );
  NAND2_X1 U758 ( .A1(n713), .A2(n712), .ZN(n773) );
  OR2_X1 U759 ( .A1(n713), .A2(n712), .ZN(n771) );
  NAND3_X1 U760 ( .A1(n774), .A2(n656), .A3(n718), .ZN(n712) );
  NOR2_X1 U761 ( .A1(n706), .A2(n483), .ZN(n718) );
  NAND2_X1 U762 ( .A1(n775), .A2(n776), .ZN(n713) );
  NAND2_X1 U763 ( .A1(n777), .A2(n778), .ZN(n776) );
  XNOR2_X1 U764 ( .A(n779), .B(n780), .ZN(n703) );
  XOR2_X1 U765 ( .A(n775), .B(n781), .Z(n780) );
  NAND2_X1 U766 ( .A1(n774), .A2(n547), .ZN(n779) );
  NAND2_X1 U767 ( .A1(n695), .A2(n698), .ZN(n765) );
  NAND2_X1 U768 ( .A1(n535), .A2(n655), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n782), .B(n783), .ZN(n695) );
  XOR2_X1 U770 ( .A(n784), .B(n785), .Z(n782) );
  OR2_X1 U771 ( .A1(n730), .A2(n733), .ZN(n755) );
  NOR2_X1 U772 ( .A1(n526), .A2(n706), .ZN(n733) );
  INV_X1 U773 ( .A(n655), .ZN(n706) );
  XOR2_X1 U774 ( .A(n786), .B(n787), .Z(n655) );
  XOR2_X1 U775 ( .A(d_3_), .B(c_3_), .Z(n787) );
  XOR2_X1 U776 ( .A(n788), .B(n789), .Z(n730) );
  XOR2_X1 U777 ( .A(n790), .B(n791), .Z(n788) );
  NOR2_X1 U778 ( .A1(n720), .A2(n530), .ZN(n791) );
  NAND2_X1 U779 ( .A1(n745), .A2(n744), .ZN(n746) );
  INV_X1 U780 ( .A(n516), .ZN(n743) );
  XNOR2_X1 U781 ( .A(n792), .B(n793), .ZN(n516) );
  XOR2_X1 U782 ( .A(n794), .B(n795), .Z(n792) );
  NOR2_X1 U783 ( .A1(n720), .A2(n575), .ZN(n795) );
  INV_X1 U784 ( .A(n449), .ZN(n575) );
  NAND2_X1 U785 ( .A1(n796), .A2(n747), .ZN(n478) );
  INV_X1 U786 ( .A(n508), .ZN(n747) );
  NOR2_X1 U787 ( .A1(n744), .A2(n745), .ZN(n508) );
  AND2_X1 U788 ( .A1(n797), .A2(n798), .ZN(n745) );
  NAND3_X1 U789 ( .A1(n774), .A2(n799), .A3(n449), .ZN(n798) );
  OR2_X1 U790 ( .A1(n794), .A2(n793), .ZN(n799) );
  NAND2_X1 U791 ( .A1(n793), .A2(n794), .ZN(n797) );
  NAND2_X1 U792 ( .A1(n753), .A2(n800), .ZN(n794) );
  NAND2_X1 U793 ( .A1(n752), .A2(n754), .ZN(n800) );
  NAND2_X1 U794 ( .A1(n801), .A2(n802), .ZN(n754) );
  NAND2_X1 U795 ( .A1(n570), .A2(n774), .ZN(n802) );
  INV_X1 U796 ( .A(n803), .ZN(n801) );
  XOR2_X1 U797 ( .A(n804), .B(n805), .Z(n752) );
  XOR2_X1 U798 ( .A(n806), .B(n807), .Z(n804) );
  NAND2_X1 U799 ( .A1(n570), .A2(n803), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n808), .A2(n809), .ZN(n803) );
  NAND3_X1 U801 ( .A1(n774), .A2(n810), .A3(n588), .ZN(n809) );
  OR2_X1 U802 ( .A1(n790), .A2(n789), .ZN(n810) );
  NAND2_X1 U803 ( .A1(n789), .A2(n790), .ZN(n808) );
  NAND2_X1 U804 ( .A1(n763), .A2(n811), .ZN(n790) );
  NAND2_X1 U805 ( .A1(n762), .A2(n764), .ZN(n811) );
  NAND2_X1 U806 ( .A1(n812), .A2(n813), .ZN(n764) );
  NAND2_X1 U807 ( .A1(n535), .A2(n774), .ZN(n813) );
  INV_X1 U808 ( .A(n814), .ZN(n812) );
  XNOR2_X1 U809 ( .A(n815), .B(n816), .ZN(n762) );
  XNOR2_X1 U810 ( .A(n817), .B(n818), .ZN(n816) );
  NAND2_X1 U811 ( .A1(n535), .A2(n814), .ZN(n763) );
  NAND2_X1 U812 ( .A1(n819), .A2(n820), .ZN(n814) );
  NAND2_X1 U813 ( .A1(n785), .A2(n821), .ZN(n820) );
  OR2_X1 U814 ( .A1(n783), .A2(n784), .ZN(n821) );
  NOR2_X1 U815 ( .A1(n543), .A2(n720), .ZN(n785) );
  INV_X1 U816 ( .A(n774), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n783), .A2(n784), .ZN(n819) );
  NAND2_X1 U818 ( .A1(n822), .A2(n823), .ZN(n784) );
  NAND3_X1 U819 ( .A1(n547), .A2(n824), .A3(n774), .ZN(n823) );
  NAND2_X1 U820 ( .A1(n775), .A2(n781), .ZN(n824) );
  OR2_X1 U821 ( .A1(n781), .A2(n775), .ZN(n822) );
  OR2_X1 U822 ( .A1(n778), .A2(n777), .ZN(n775) );
  NAND2_X1 U823 ( .A1(n825), .A2(n656), .ZN(n777) );
  NAND2_X1 U824 ( .A1(n774), .A2(n658), .ZN(n778) );
  XOR2_X1 U825 ( .A(n826), .B(n827), .Z(n774) );
  XOR2_X1 U826 ( .A(d_2_), .B(c_2_), .Z(n827) );
  NAND2_X1 U827 ( .A1(n828), .A2(n829), .ZN(n781) );
  NAND2_X1 U828 ( .A1(n830), .A2(n831), .ZN(n829) );
  XOR2_X1 U829 ( .A(n832), .B(n828), .Z(n783) );
  NAND2_X1 U830 ( .A1(n833), .A2(n834), .ZN(n832) );
  NAND2_X1 U831 ( .A1(n835), .A2(n836), .ZN(n834) );
  NAND2_X1 U832 ( .A1(n507), .A2(n658), .ZN(n835) );
  XOR2_X1 U833 ( .A(n837), .B(n838), .Z(n789) );
  XOR2_X1 U834 ( .A(n839), .B(n840), .Z(n837) );
  XOR2_X1 U835 ( .A(n841), .B(n842), .Z(n793) );
  XOR2_X1 U836 ( .A(n843), .B(n844), .Z(n841) );
  XNOR2_X1 U837 ( .A(n845), .B(n846), .ZN(n744) );
  NOR2_X1 U838 ( .A1(n526), .A2(n847), .ZN(n846) );
  INV_X1 U839 ( .A(n570), .ZN(n526) );
  XOR2_X1 U840 ( .A(n848), .B(n849), .Z(n845) );
  XOR2_X1 U841 ( .A(n479), .B(n850), .Z(n796) );
  NAND2_X1 U842 ( .A1(n449), .A2(n507), .ZN(n850) );
  NAND2_X1 U843 ( .A1(n851), .A2(n852), .ZN(n479) );
  NAND3_X1 U844 ( .A1(n570), .A2(n853), .A3(n507), .ZN(n852) );
  OR2_X1 U845 ( .A1(n848), .A2(n849), .ZN(n853) );
  NAND2_X1 U846 ( .A1(n849), .A2(n848), .ZN(n851) );
  NAND2_X1 U847 ( .A1(n854), .A2(n855), .ZN(n848) );
  NAND2_X1 U848 ( .A1(n842), .A2(n856), .ZN(n855) );
  OR2_X1 U849 ( .A1(n843), .A2(n844), .ZN(n856) );
  NOR2_X1 U850 ( .A1(n847), .A2(n530), .ZN(n842) );
  INV_X1 U851 ( .A(n588), .ZN(n530) );
  NAND2_X1 U852 ( .A1(n844), .A2(n843), .ZN(n854) );
  NAND2_X1 U853 ( .A1(n857), .A2(n858), .ZN(n843) );
  NAND2_X1 U854 ( .A1(n805), .A2(n859), .ZN(n858) );
  OR2_X1 U855 ( .A1(n806), .A2(n807), .ZN(n859) );
  AND2_X1 U856 ( .A1(n588), .A2(n825), .ZN(n805) );
  XOR2_X1 U857 ( .A(n860), .B(n861), .Z(n588) );
  XOR2_X1 U858 ( .A(b_2_), .B(a_2_), .Z(n861) );
  NAND2_X1 U859 ( .A1(n807), .A2(n806), .ZN(n857) );
  NAND2_X1 U860 ( .A1(n862), .A2(n863), .ZN(n806) );
  NAND2_X1 U861 ( .A1(n838), .A2(n864), .ZN(n863) );
  NAND2_X1 U862 ( .A1(n840), .A2(n839), .ZN(n864) );
  NOR2_X1 U863 ( .A1(n847), .A2(n543), .ZN(n838) );
  INV_X1 U864 ( .A(n642), .ZN(n543) );
  OR2_X1 U865 ( .A1(n839), .A2(n840), .ZN(n862) );
  AND2_X1 U866 ( .A1(n865), .A2(n866), .ZN(n840) );
  NAND2_X1 U867 ( .A1(n815), .A2(n867), .ZN(n866) );
  OR2_X1 U868 ( .A1(n818), .A2(n817), .ZN(n867) );
  NOR2_X1 U869 ( .A1(n847), .A2(n489), .ZN(n815) );
  INV_X1 U870 ( .A(n547), .ZN(n489) );
  NAND2_X1 U871 ( .A1(n817), .A2(n818), .ZN(n865) );
  NAND2_X1 U872 ( .A1(n828), .A2(n833), .ZN(n818) );
  OR3_X1 U873 ( .A1(n847), .A2(n483), .A3(n836), .ZN(n833) );
  NAND2_X1 U874 ( .A1(n825), .A2(n547), .ZN(n836) );
  XOR2_X1 U875 ( .A(n868), .B(n869), .Z(n547) );
  XOR2_X1 U876 ( .A(b_5_), .B(a_5_), .Z(n869) );
  OR2_X1 U877 ( .A1(n831), .A2(n830), .ZN(n828) );
  NAND2_X1 U878 ( .A1(n825), .A2(n658), .ZN(n830) );
  INV_X1 U879 ( .A(n483), .ZN(n658) );
  XOR2_X1 U880 ( .A(n870), .B(n871), .Z(n483) );
  XOR2_X1 U881 ( .A(b_6_), .B(a_6_), .Z(n871) );
  NAND2_X1 U882 ( .A1(b_7_), .A2(a_7_), .ZN(n870) );
  NAND2_X1 U883 ( .A1(n507), .A2(n656), .ZN(n831) );
  INV_X1 U884 ( .A(n550), .ZN(n656) );
  XNOR2_X1 U885 ( .A(a_7_), .B(b_7_), .ZN(n550) );
  AND2_X1 U886 ( .A1(n642), .A2(n825), .ZN(n817) );
  XOR2_X1 U887 ( .A(n872), .B(n873), .Z(n642) );
  XOR2_X1 U888 ( .A(b_4_), .B(a_4_), .Z(n873) );
  NAND2_X1 U889 ( .A1(n535), .A2(n825), .ZN(n839) );
  NOR2_X1 U890 ( .A1(n847), .A2(n500), .ZN(n807) );
  INV_X1 U891 ( .A(n535), .ZN(n500) );
  XOR2_X1 U892 ( .A(n874), .B(n875), .Z(n535) );
  XOR2_X1 U893 ( .A(b_3_), .B(a_3_), .Z(n875) );
  INV_X1 U894 ( .A(n507), .ZN(n847) );
  XOR2_X1 U895 ( .A(n876), .B(n877), .Z(n507) );
  XOR2_X1 U896 ( .A(d_0_), .B(c_0_), .Z(n877) );
  NAND2_X1 U897 ( .A1(n878), .A2(n879), .ZN(n876) );
  NAND2_X1 U898 ( .A1(d_1_), .A2(n880), .ZN(n879) );
  OR2_X1 U899 ( .A1(n881), .A2(c_1_), .ZN(n880) );
  NAND2_X1 U900 ( .A1(c_1_), .A2(n881), .ZN(n878) );
  AND2_X1 U901 ( .A1(n570), .A2(n825), .ZN(n844) );
  XOR2_X1 U902 ( .A(n882), .B(n883), .Z(n570) );
  XOR2_X1 U903 ( .A(b_1_), .B(a_1_), .Z(n883) );
  AND2_X1 U904 ( .A1(n449), .A2(n825), .ZN(n849) );
  XOR2_X1 U905 ( .A(n881), .B(n884), .Z(n825) );
  XOR2_X1 U906 ( .A(d_1_), .B(c_1_), .Z(n884) );
  NAND2_X1 U907 ( .A1(n885), .A2(n886), .ZN(n881) );
  NAND2_X1 U908 ( .A1(d_2_), .A2(n887), .ZN(n886) );
  OR2_X1 U909 ( .A1(n826), .A2(c_2_), .ZN(n887) );
  NAND2_X1 U910 ( .A1(c_2_), .A2(n826), .ZN(n885) );
  NAND2_X1 U911 ( .A1(n888), .A2(n889), .ZN(n826) );
  NAND2_X1 U912 ( .A1(d_3_), .A2(n890), .ZN(n889) );
  OR2_X1 U913 ( .A1(n786), .A2(c_3_), .ZN(n890) );
  NAND2_X1 U914 ( .A1(c_3_), .A2(n786), .ZN(n888) );
  NAND2_X1 U915 ( .A1(n891), .A2(n892), .ZN(n786) );
  NAND2_X1 U916 ( .A1(d_4_), .A2(n893), .ZN(n892) );
  OR2_X1 U917 ( .A1(n721), .A2(c_4_), .ZN(n893) );
  NAND2_X1 U918 ( .A1(c_4_), .A2(n721), .ZN(n891) );
  NAND2_X1 U919 ( .A1(n894), .A2(n895), .ZN(n721) );
  NAND2_X1 U920 ( .A1(d_5_), .A2(n896), .ZN(n895) );
  OR2_X1 U921 ( .A1(n659), .A2(c_5_), .ZN(n896) );
  NAND2_X1 U922 ( .A1(c_5_), .A2(n659), .ZN(n894) );
  NAND2_X1 U923 ( .A1(n897), .A2(n898), .ZN(n659) );
  NAND3_X1 U924 ( .A1(c_7_), .A2(n899), .A3(d_7_), .ZN(n898) );
  OR2_X1 U925 ( .A1(d_6_), .A2(c_6_), .ZN(n899) );
  NAND2_X1 U926 ( .A1(d_6_), .A2(c_6_), .ZN(n897) );
  XOR2_X1 U927 ( .A(b_0_), .B(a_0_), .Z(n901) );
  NAND2_X1 U928 ( .A1(n902), .A2(n903), .ZN(n900) );
  NAND2_X1 U929 ( .A1(b_1_), .A2(n904), .ZN(n903) );
  OR2_X1 U930 ( .A1(n882), .A2(a_1_), .ZN(n904) );
  NAND2_X1 U931 ( .A1(a_1_), .A2(n882), .ZN(n902) );
  NAND2_X1 U932 ( .A1(n905), .A2(n906), .ZN(n882) );
  NAND2_X1 U933 ( .A1(b_2_), .A2(n907), .ZN(n906) );
  OR2_X1 U934 ( .A1(n860), .A2(a_2_), .ZN(n907) );
  NAND2_X1 U935 ( .A1(a_2_), .A2(n860), .ZN(n905) );
  NAND2_X1 U936 ( .A1(n908), .A2(n909), .ZN(n860) );
  NAND2_X1 U937 ( .A1(b_3_), .A2(n910), .ZN(n909) );
  OR2_X1 U938 ( .A1(n874), .A2(a_3_), .ZN(n910) );
  NAND2_X1 U939 ( .A1(a_3_), .A2(n874), .ZN(n908) );
  NAND2_X1 U940 ( .A1(n911), .A2(n912), .ZN(n874) );
  NAND2_X1 U941 ( .A1(b_4_), .A2(n913), .ZN(n912) );
  OR2_X1 U942 ( .A1(n872), .A2(a_4_), .ZN(n913) );
  NAND2_X1 U943 ( .A1(a_4_), .A2(n872), .ZN(n911) );
  NAND2_X1 U944 ( .A1(n914), .A2(n915), .ZN(n872) );
  NAND2_X1 U945 ( .A1(b_5_), .A2(n916), .ZN(n915) );
  OR2_X1 U946 ( .A1(n868), .A2(a_5_), .ZN(n916) );
  NAND2_X1 U947 ( .A1(a_5_), .A2(n868), .ZN(n914) );
  NAND2_X1 U948 ( .A1(n917), .A2(n918), .ZN(n868) );
  NAND3_X1 U949 ( .A1(a_7_), .A2(n919), .A3(b_7_), .ZN(n918) );
  OR2_X1 U950 ( .A1(b_6_), .A2(a_6_), .ZN(n919) );
  NAND2_X1 U951 ( .A1(b_6_), .A2(a_6_), .ZN(n917) );
endmodule

