module add_mul_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, 
        b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, operation, Result_0_, 
        Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, 
        Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, 
        Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;

  NAND2_X1 U516 ( .A1(n500), .A2(n501), .ZN(Result_9_) );
  NAND2_X1 U517 ( .A1(n502), .A2(operation), .ZN(n501) );
  XNOR2_X1 U518 ( .A(n503), .B(n504), .ZN(n502) );
  XNOR2_X1 U519 ( .A(n505), .B(n506), .ZN(n503) );
  NOR2_X1 U520 ( .A1(n507), .A2(n508), .ZN(n506) );
  NAND2_X1 U521 ( .A1(n509), .A2(n510), .ZN(n500) );
  NAND2_X1 U522 ( .A1(n511), .A2(n512), .ZN(n509) );
  INV_X1 U523 ( .A(n513), .ZN(n512) );
  NOR2_X1 U524 ( .A1(n514), .A2(n515), .ZN(n513) );
  NOR2_X1 U525 ( .A1(n516), .A2(n517), .ZN(n514) );
  NAND2_X1 U526 ( .A1(n518), .A2(n515), .ZN(n511) );
  INV_X1 U527 ( .A(n519), .ZN(n515) );
  XOR2_X1 U528 ( .A(b_1_), .B(a_1_), .Z(n518) );
  NAND2_X1 U529 ( .A1(n520), .A2(n521), .ZN(Result_8_) );
  NAND2_X1 U530 ( .A1(n522), .A2(n510), .ZN(n521) );
  XOR2_X1 U531 ( .A(n523), .B(n524), .Z(n522) );
  NOR2_X1 U532 ( .A1(n525), .A2(n526), .ZN(n524) );
  NOR2_X1 U533 ( .A1(b_0_), .A2(a_0_), .ZN(n525) );
  NOR2_X1 U534 ( .A1(n517), .A2(n527), .ZN(n523) );
  NOR2_X1 U535 ( .A1(n516), .A2(n519), .ZN(n527) );
  NAND2_X1 U536 ( .A1(n528), .A2(n529), .ZN(n519) );
  NAND2_X1 U537 ( .A1(n530), .A2(n531), .ZN(n529) );
  NOR2_X1 U538 ( .A1(b_1_), .A2(a_1_), .ZN(n517) );
  NAND2_X1 U539 ( .A1(n532), .A2(operation), .ZN(n520) );
  XOR2_X1 U540 ( .A(n533), .B(n534), .Z(n532) );
  XNOR2_X1 U541 ( .A(n535), .B(n536), .ZN(n534) );
  NOR2_X1 U542 ( .A1(n537), .A2(n510), .ZN(Result_7_) );
  XOR2_X1 U543 ( .A(n538), .B(n539), .Z(n537) );
  NOR2_X1 U544 ( .A1(n510), .A2(n540), .ZN(Result_6_) );
  NAND2_X1 U545 ( .A1(n541), .A2(n542), .ZN(n540) );
  NAND2_X1 U546 ( .A1(n543), .A2(n544), .ZN(n541) );
  NAND2_X1 U547 ( .A1(n538), .A2(n545), .ZN(n544) );
  INV_X1 U548 ( .A(n539), .ZN(n545) );
  NOR2_X1 U549 ( .A1(n546), .A2(n510), .ZN(Result_5_) );
  XOR2_X1 U550 ( .A(n542), .B(n547), .Z(n546) );
  NOR2_X1 U551 ( .A1(n548), .A2(n549), .ZN(n547) );
  NOR2_X1 U552 ( .A1(n550), .A2(n551), .ZN(n549) );
  NOR2_X1 U553 ( .A1(n552), .A2(n510), .ZN(Result_4_) );
  XOR2_X1 U554 ( .A(n553), .B(n554), .Z(n552) );
  NOR2_X1 U555 ( .A1(n555), .A2(n510), .ZN(Result_3_) );
  XNOR2_X1 U556 ( .A(n556), .B(n557), .ZN(n555) );
  NOR2_X1 U557 ( .A1(n558), .A2(n553), .ZN(n557) );
  INV_X1 U558 ( .A(n554), .ZN(n558) );
  NOR2_X1 U559 ( .A1(n559), .A2(n560), .ZN(n556) );
  NOR2_X1 U560 ( .A1(n561), .A2(n562), .ZN(n559) );
  NOR2_X1 U561 ( .A1(n510), .A2(n563), .ZN(Result_2_) );
  XNOR2_X1 U562 ( .A(n564), .B(n565), .ZN(n563) );
  NOR2_X1 U563 ( .A1(n566), .A2(n510), .ZN(Result_1_) );
  XNOR2_X1 U564 ( .A(n567), .B(n568), .ZN(n566) );
  NAND2_X1 U565 ( .A1(n564), .A2(n565), .ZN(n568) );
  NAND2_X1 U566 ( .A1(n569), .A2(n570), .ZN(n567) );
  NAND2_X1 U567 ( .A1(n571), .A2(n572), .ZN(Result_15_) );
  NAND2_X1 U568 ( .A1(n573), .A2(n510), .ZN(n572) );
  XOR2_X1 U569 ( .A(b_7_), .B(a_7_), .Z(n573) );
  NAND2_X1 U570 ( .A1(operation), .A2(n574), .ZN(n571) );
  NAND2_X1 U571 ( .A1(n575), .A2(n576), .ZN(Result_14_) );
  NAND2_X1 U572 ( .A1(n577), .A2(n510), .ZN(n576) );
  NAND2_X1 U573 ( .A1(n578), .A2(n579), .ZN(n577) );
  NOR2_X1 U574 ( .A1(n580), .A2(n581), .ZN(n578) );
  NOR2_X1 U575 ( .A1(n582), .A2(n583), .ZN(n581) );
  NAND2_X1 U576 ( .A1(n584), .A2(n585), .ZN(n583) );
  NOR2_X1 U577 ( .A1(b_6_), .A2(n586), .ZN(n580) );
  XOR2_X1 U578 ( .A(n584), .B(a_6_), .Z(n586) );
  NAND2_X1 U579 ( .A1(n587), .A2(operation), .ZN(n575) );
  XNOR2_X1 U580 ( .A(n588), .B(n589), .ZN(n587) );
  NAND2_X1 U581 ( .A1(a_6_), .A2(b_7_), .ZN(n589) );
  NAND2_X1 U582 ( .A1(n590), .A2(n591), .ZN(Result_13_) );
  NAND2_X1 U583 ( .A1(n592), .A2(n510), .ZN(n591) );
  NAND2_X1 U584 ( .A1(n593), .A2(n594), .ZN(n592) );
  NAND2_X1 U585 ( .A1(n595), .A2(n596), .ZN(n594) );
  NOR2_X1 U586 ( .A1(n597), .A2(n598), .ZN(n593) );
  NOR2_X1 U587 ( .A1(b_5_), .A2(n599), .ZN(n598) );
  XOR2_X1 U588 ( .A(a_5_), .B(n600), .Z(n599) );
  NOR2_X1 U589 ( .A1(n601), .A2(n602), .ZN(n597) );
  NAND2_X1 U590 ( .A1(n600), .A2(n603), .ZN(n602) );
  INV_X1 U591 ( .A(n596), .ZN(n600) );
  NAND2_X1 U592 ( .A1(n604), .A2(operation), .ZN(n590) );
  XOR2_X1 U593 ( .A(n605), .B(n606), .Z(n604) );
  XOR2_X1 U594 ( .A(n607), .B(n608), .Z(n606) );
  NAND2_X1 U595 ( .A1(n609), .A2(n610), .ZN(Result_12_) );
  NAND2_X1 U596 ( .A1(n611), .A2(n510), .ZN(n610) );
  XNOR2_X1 U597 ( .A(n612), .B(n613), .ZN(n611) );
  NAND2_X1 U598 ( .A1(n614), .A2(n615), .ZN(n612) );
  NAND2_X1 U599 ( .A1(n616), .A2(operation), .ZN(n609) );
  XNOR2_X1 U600 ( .A(n617), .B(n618), .ZN(n616) );
  NAND2_X1 U601 ( .A1(n619), .A2(n620), .ZN(n617) );
  NAND2_X1 U602 ( .A1(n621), .A2(n622), .ZN(Result_11_) );
  NAND2_X1 U603 ( .A1(n623), .A2(n510), .ZN(n622) );
  NAND2_X1 U604 ( .A1(n624), .A2(n625), .ZN(n623) );
  NAND2_X1 U605 ( .A1(n626), .A2(n627), .ZN(n625) );
  NOR2_X1 U606 ( .A1(n628), .A2(n629), .ZN(n624) );
  NOR2_X1 U607 ( .A1(b_3_), .A2(n630), .ZN(n629) );
  XOR2_X1 U608 ( .A(n631), .B(n627), .Z(n630) );
  NOR2_X1 U609 ( .A1(n632), .A2(n633), .ZN(n628) );
  INV_X1 U610 ( .A(n634), .ZN(n633) );
  NOR2_X1 U611 ( .A1(n627), .A2(a_3_), .ZN(n634) );
  NAND2_X1 U612 ( .A1(n635), .A2(operation), .ZN(n621) );
  XOR2_X1 U613 ( .A(n636), .B(n637), .Z(n635) );
  XOR2_X1 U614 ( .A(n638), .B(n639), .Z(n636) );
  NOR2_X1 U615 ( .A1(n507), .A2(n631), .ZN(n639) );
  NAND2_X1 U616 ( .A1(n640), .A2(n641), .ZN(Result_10_) );
  NAND2_X1 U617 ( .A1(n642), .A2(n510), .ZN(n641) );
  XNOR2_X1 U618 ( .A(n531), .B(n643), .ZN(n642) );
  NAND2_X1 U619 ( .A1(n530), .A2(n528), .ZN(n643) );
  NAND2_X1 U620 ( .A1(n644), .A2(n645), .ZN(n530) );
  NAND2_X1 U621 ( .A1(n646), .A2(n647), .ZN(n531) );
  NAND2_X1 U622 ( .A1(n648), .A2(n627), .ZN(n647) );
  NAND2_X1 U623 ( .A1(n614), .A2(n649), .ZN(n627) );
  NAND2_X1 U624 ( .A1(n615), .A2(n613), .ZN(n649) );
  NAND2_X1 U625 ( .A1(n650), .A2(n651), .ZN(n613) );
  NAND2_X1 U626 ( .A1(n652), .A2(n596), .ZN(n651) );
  NAND2_X1 U627 ( .A1(n653), .A2(n654), .ZN(n596) );
  NAND2_X1 U628 ( .A1(n574), .A2(n655), .ZN(n654) );
  NAND2_X1 U629 ( .A1(n582), .A2(n585), .ZN(n655) );
  INV_X1 U630 ( .A(n584), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n601), .A2(n603), .ZN(n652) );
  NAND2_X1 U632 ( .A1(n656), .A2(n657), .ZN(n615) );
  NAND2_X1 U633 ( .A1(n632), .A2(n631), .ZN(n648) );
  NAND2_X1 U634 ( .A1(n658), .A2(operation), .ZN(n640) );
  XOR2_X1 U635 ( .A(n659), .B(n660), .Z(n658) );
  XNOR2_X1 U636 ( .A(n661), .B(n662), .ZN(n660) );
  NOR2_X1 U637 ( .A1(n663), .A2(n510), .ZN(Result_0_) );
  INV_X1 U638 ( .A(operation), .ZN(n510) );
  NOR2_X1 U639 ( .A1(n664), .A2(n665), .ZN(n663) );
  NAND2_X1 U640 ( .A1(n666), .A2(n570), .ZN(n665) );
  INV_X1 U641 ( .A(n667), .ZN(n570) );
  NOR2_X1 U642 ( .A1(n668), .A2(n669), .ZN(n667) );
  NAND2_X1 U643 ( .A1(n670), .A2(n526), .ZN(n668) );
  NAND2_X1 U644 ( .A1(n671), .A2(n565), .ZN(n666) );
  XOR2_X1 U645 ( .A(n672), .B(n673), .Z(n565) );
  INV_X1 U646 ( .A(n674), .ZN(n671) );
  NAND2_X1 U647 ( .A1(n564), .A2(n569), .ZN(n674) );
  NAND2_X1 U648 ( .A1(n675), .A2(n669), .ZN(n569) );
  NAND2_X1 U649 ( .A1(n672), .A2(n673), .ZN(n669) );
  XOR2_X1 U650 ( .A(n676), .B(n677), .Z(n673) );
  NOR2_X1 U651 ( .A1(n508), .A2(n678), .ZN(n677) );
  XOR2_X1 U652 ( .A(n679), .B(n680), .Z(n676) );
  NAND2_X1 U653 ( .A1(n681), .A2(n682), .ZN(n672) );
  NAND2_X1 U654 ( .A1(n683), .A2(n684), .ZN(n682) );
  INV_X1 U655 ( .A(n685), .ZN(n684) );
  NOR2_X1 U656 ( .A1(n686), .A2(n687), .ZN(n685) );
  NAND2_X1 U657 ( .A1(n686), .A2(n687), .ZN(n681) );
  XOR2_X1 U658 ( .A(n526), .B(n670), .Z(n675) );
  NOR2_X1 U659 ( .A1(n688), .A2(n678), .ZN(n526) );
  NAND2_X1 U660 ( .A1(n689), .A2(n690), .ZN(n564) );
  NAND2_X1 U661 ( .A1(n691), .A2(n692), .ZN(n690) );
  NOR2_X1 U662 ( .A1(n560), .A2(n693), .ZN(n689) );
  NOR2_X1 U663 ( .A1(n553), .A2(n694), .ZN(n693) );
  NAND2_X1 U664 ( .A1(n561), .A2(n554), .ZN(n694) );
  NAND2_X1 U665 ( .A1(n695), .A2(n696), .ZN(n554) );
  NAND2_X1 U666 ( .A1(n697), .A2(n551), .ZN(n696) );
  INV_X1 U667 ( .A(n542), .ZN(n697) );
  NAND2_X1 U668 ( .A1(n698), .A2(n538), .ZN(n542) );
  NOR2_X1 U669 ( .A1(n699), .A2(n700), .ZN(n538) );
  INV_X1 U670 ( .A(n701), .ZN(n700) );
  NAND2_X1 U671 ( .A1(n533), .A2(n702), .ZN(n701) );
  NAND2_X1 U672 ( .A1(n536), .A2(n535), .ZN(n702) );
  XNOR2_X1 U673 ( .A(n703), .B(n704), .ZN(n533) );
  XOR2_X1 U674 ( .A(n705), .B(n706), .Z(n703) );
  NOR2_X1 U675 ( .A1(n582), .A2(n508), .ZN(n706) );
  NOR2_X1 U676 ( .A1(n535), .A2(n536), .ZN(n699) );
  NOR2_X1 U677 ( .A1(n688), .A2(n507), .ZN(n536) );
  NAND2_X1 U678 ( .A1(n707), .A2(n708), .ZN(n535) );
  NAND2_X1 U679 ( .A1(n709), .A2(a_1_), .ZN(n708) );
  NOR2_X1 U680 ( .A1(n710), .A2(n507), .ZN(n709) );
  NOR2_X1 U681 ( .A1(n505), .A2(n504), .ZN(n710) );
  NAND2_X1 U682 ( .A1(n504), .A2(n505), .ZN(n707) );
  NOR2_X1 U683 ( .A1(n711), .A2(n712), .ZN(n505) );
  INV_X1 U684 ( .A(n713), .ZN(n712) );
  NAND2_X1 U685 ( .A1(n659), .A2(n714), .ZN(n713) );
  NAND2_X1 U686 ( .A1(n662), .A2(n661), .ZN(n714) );
  XNOR2_X1 U687 ( .A(n715), .B(n716), .ZN(n659) );
  XOR2_X1 U688 ( .A(n717), .B(n718), .Z(n715) );
  NOR2_X1 U689 ( .A1(n661), .A2(n662), .ZN(n711) );
  NOR2_X1 U690 ( .A1(n645), .A2(n507), .ZN(n662) );
  NAND2_X1 U691 ( .A1(n719), .A2(n720), .ZN(n661) );
  NAND2_X1 U692 ( .A1(n721), .A2(a_3_), .ZN(n720) );
  NOR2_X1 U693 ( .A1(n722), .A2(n507), .ZN(n721) );
  NOR2_X1 U694 ( .A1(n637), .A2(n638), .ZN(n722) );
  NAND2_X1 U695 ( .A1(n637), .A2(n638), .ZN(n719) );
  NAND2_X1 U696 ( .A1(n619), .A2(n723), .ZN(n638) );
  NAND2_X1 U697 ( .A1(n618), .A2(n620), .ZN(n723) );
  NAND2_X1 U698 ( .A1(n724), .A2(n725), .ZN(n620) );
  NAND2_X1 U699 ( .A1(a_4_), .A2(b_7_), .ZN(n725) );
  XNOR2_X1 U700 ( .A(n726), .B(n727), .ZN(n618) );
  XOR2_X1 U701 ( .A(n728), .B(n729), .Z(n726) );
  INV_X1 U702 ( .A(n730), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n657), .A2(n724), .ZN(n730) );
  NOR2_X1 U704 ( .A1(n731), .A2(n732), .ZN(n724) );
  NOR2_X1 U705 ( .A1(n579), .A2(n733), .ZN(n732) );
  NOR2_X1 U706 ( .A1(n605), .A2(n608), .ZN(n733) );
  INV_X1 U707 ( .A(n607), .ZN(n579) );
  NOR2_X1 U708 ( .A1(n653), .A2(n584), .ZN(n607) );
  NAND2_X1 U709 ( .A1(b_7_), .A2(a_7_), .ZN(n584) );
  INV_X1 U710 ( .A(n734), .ZN(n731) );
  NAND2_X1 U711 ( .A1(n608), .A2(n605), .ZN(n734) );
  XNOR2_X1 U712 ( .A(n653), .B(n735), .ZN(n605) );
  NOR2_X1 U713 ( .A1(n736), .A2(n601), .ZN(n735) );
  NAND2_X1 U714 ( .A1(b_6_), .A2(a_6_), .ZN(n653) );
  NOR2_X1 U715 ( .A1(n603), .A2(n507), .ZN(n608) );
  INV_X1 U716 ( .A(b_7_), .ZN(n507) );
  XNOR2_X1 U717 ( .A(n737), .B(n738), .ZN(n637) );
  XNOR2_X1 U718 ( .A(n739), .B(n740), .ZN(n738) );
  XOR2_X1 U719 ( .A(n741), .B(n742), .Z(n504) );
  XOR2_X1 U720 ( .A(n743), .B(n744), .Z(n741) );
  NOR2_X1 U721 ( .A1(n539), .A2(n543), .ZN(n698) );
  XNOR2_X1 U722 ( .A(n745), .B(n746), .ZN(n543) );
  XNOR2_X1 U723 ( .A(n747), .B(n748), .ZN(n539) );
  XNOR2_X1 U724 ( .A(n749), .B(n750), .ZN(n748) );
  NOR2_X1 U725 ( .A1(n548), .A2(n751), .ZN(n695) );
  NOR2_X1 U726 ( .A1(n752), .A2(n753), .ZN(n751) );
  INV_X1 U727 ( .A(n754), .ZN(n548) );
  NAND2_X1 U728 ( .A1(n550), .A2(n551), .ZN(n754) );
  XOR2_X1 U729 ( .A(n753), .B(n752), .Z(n551) );
  XOR2_X1 U730 ( .A(n755), .B(n756), .Z(n752) );
  XOR2_X1 U731 ( .A(n757), .B(n758), .Z(n756) );
  NAND2_X1 U732 ( .A1(n759), .A2(n760), .ZN(n753) );
  NAND2_X1 U733 ( .A1(n761), .A2(n762), .ZN(n760) );
  NAND2_X1 U734 ( .A1(n763), .A2(n764), .ZN(n762) );
  INV_X1 U735 ( .A(n765), .ZN(n759) );
  NOR2_X1 U736 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U737 ( .A1(n746), .A2(n745), .ZN(n550) );
  NAND2_X1 U738 ( .A1(n766), .A2(n767), .ZN(n745) );
  NAND2_X1 U739 ( .A1(n747), .A2(n768), .ZN(n767) );
  NAND2_X1 U740 ( .A1(n750), .A2(n749), .ZN(n768) );
  XOR2_X1 U741 ( .A(n769), .B(n770), .Z(n747) );
  XOR2_X1 U742 ( .A(n771), .B(n772), .Z(n770) );
  NAND2_X1 U743 ( .A1(a_1_), .A2(b_5_), .ZN(n772) );
  INV_X1 U744 ( .A(n773), .ZN(n766) );
  NOR2_X1 U745 ( .A1(n749), .A2(n750), .ZN(n773) );
  NOR2_X1 U746 ( .A1(n688), .A2(n582), .ZN(n750) );
  NAND2_X1 U747 ( .A1(n774), .A2(n775), .ZN(n749) );
  NAND2_X1 U748 ( .A1(n776), .A2(a_1_), .ZN(n775) );
  NOR2_X1 U749 ( .A1(n777), .A2(n582), .ZN(n776) );
  NOR2_X1 U750 ( .A1(n705), .A2(n704), .ZN(n777) );
  NAND2_X1 U751 ( .A1(n704), .A2(n705), .ZN(n774) );
  NAND2_X1 U752 ( .A1(n778), .A2(n779), .ZN(n705) );
  NAND2_X1 U753 ( .A1(n744), .A2(n780), .ZN(n779) );
  INV_X1 U754 ( .A(n781), .ZN(n780) );
  NOR2_X1 U755 ( .A1(n742), .A2(n743), .ZN(n781) );
  NOR2_X1 U756 ( .A1(n645), .A2(n582), .ZN(n744) );
  NAND2_X1 U757 ( .A1(n742), .A2(n743), .ZN(n778) );
  NAND2_X1 U758 ( .A1(n782), .A2(n783), .ZN(n743) );
  NAND2_X1 U759 ( .A1(n718), .A2(n784), .ZN(n783) );
  INV_X1 U760 ( .A(n785), .ZN(n784) );
  NOR2_X1 U761 ( .A1(n717), .A2(n716), .ZN(n785) );
  NOR2_X1 U762 ( .A1(n631), .A2(n582), .ZN(n718) );
  NAND2_X1 U763 ( .A1(n716), .A2(n717), .ZN(n782) );
  NAND2_X1 U764 ( .A1(n786), .A2(n787), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n740), .A2(n788), .ZN(n787) );
  NAND2_X1 U766 ( .A1(n737), .A2(n739), .ZN(n788) );
  NOR2_X1 U767 ( .A1(n657), .A2(n582), .ZN(n740) );
  INV_X1 U768 ( .A(n789), .ZN(n786) );
  NOR2_X1 U769 ( .A1(n739), .A2(n737), .ZN(n789) );
  XNOR2_X1 U770 ( .A(n790), .B(n791), .ZN(n737) );
  XOR2_X1 U771 ( .A(n595), .B(n792), .Z(n790) );
  NAND2_X1 U772 ( .A1(n793), .A2(n794), .ZN(n739) );
  NAND2_X1 U773 ( .A1(n795), .A2(n729), .ZN(n794) );
  NAND2_X1 U774 ( .A1(n588), .A2(n796), .ZN(n729) );
  NOR2_X1 U775 ( .A1(n582), .A2(n736), .ZN(n588) );
  NAND2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n795) );
  INV_X1 U777 ( .A(n797), .ZN(n793) );
  NOR2_X1 U778 ( .A1(n727), .A2(n728), .ZN(n797) );
  NOR2_X1 U779 ( .A1(n603), .A2(n582), .ZN(n728) );
  INV_X1 U780 ( .A(b_6_), .ZN(n582) );
  XOR2_X1 U781 ( .A(n796), .B(n798), .Z(n727) );
  XNOR2_X1 U782 ( .A(n799), .B(n800), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n801), .A2(n802), .ZN(n799) );
  XNOR2_X1 U784 ( .A(n803), .B(n804), .ZN(n742) );
  XOR2_X1 U785 ( .A(n805), .B(n806), .Z(n804) );
  NAND2_X1 U786 ( .A1(a_3_), .A2(b_5_), .ZN(n806) );
  XNOR2_X1 U787 ( .A(n807), .B(n808), .ZN(n704) );
  XOR2_X1 U788 ( .A(n809), .B(n810), .Z(n808) );
  NAND2_X1 U789 ( .A1(a_2_), .A2(b_5_), .ZN(n810) );
  XNOR2_X1 U790 ( .A(n761), .B(n811), .ZN(n746) );
  XNOR2_X1 U791 ( .A(n764), .B(n763), .ZN(n811) );
  NOR2_X1 U792 ( .A1(n688), .A2(n601), .ZN(n763) );
  NAND2_X1 U793 ( .A1(n812), .A2(n813), .ZN(n764) );
  NAND2_X1 U794 ( .A1(n814), .A2(a_1_), .ZN(n813) );
  NOR2_X1 U795 ( .A1(n815), .A2(n601), .ZN(n814) );
  NOR2_X1 U796 ( .A1(n771), .A2(n769), .ZN(n815) );
  NAND2_X1 U797 ( .A1(n769), .A2(n771), .ZN(n812) );
  NAND2_X1 U798 ( .A1(n816), .A2(n817), .ZN(n771) );
  NAND2_X1 U799 ( .A1(n818), .A2(a_2_), .ZN(n817) );
  NOR2_X1 U800 ( .A1(n819), .A2(n601), .ZN(n818) );
  NOR2_X1 U801 ( .A1(n807), .A2(n809), .ZN(n819) );
  NAND2_X1 U802 ( .A1(n807), .A2(n809), .ZN(n816) );
  NAND2_X1 U803 ( .A1(n820), .A2(n821), .ZN(n809) );
  NAND2_X1 U804 ( .A1(n822), .A2(a_3_), .ZN(n821) );
  NOR2_X1 U805 ( .A1(n823), .A2(n601), .ZN(n822) );
  NOR2_X1 U806 ( .A1(n803), .A2(n805), .ZN(n823) );
  NAND2_X1 U807 ( .A1(n803), .A2(n805), .ZN(n820) );
  NAND2_X1 U808 ( .A1(n801), .A2(n824), .ZN(n805) );
  NAND2_X1 U809 ( .A1(n800), .A2(n802), .ZN(n824) );
  NAND2_X1 U810 ( .A1(n825), .A2(n826), .ZN(n802) );
  NAND2_X1 U811 ( .A1(a_4_), .A2(b_5_), .ZN(n826) );
  XNOR2_X1 U812 ( .A(n827), .B(n828), .ZN(n800) );
  NAND2_X1 U813 ( .A1(n829), .A2(n830), .ZN(n827) );
  NAND2_X1 U814 ( .A1(n831), .A2(a_4_), .ZN(n801) );
  INV_X1 U815 ( .A(n825), .ZN(n831) );
  NAND2_X1 U816 ( .A1(n832), .A2(n833), .ZN(n825) );
  NAND2_X1 U817 ( .A1(n834), .A2(n792), .ZN(n833) );
  NAND2_X1 U818 ( .A1(n796), .A2(n798), .ZN(n792) );
  NOR2_X1 U819 ( .A1(n656), .A2(n736), .ZN(n798) );
  NOR2_X1 U820 ( .A1(n601), .A2(n585), .ZN(n796) );
  INV_X1 U821 ( .A(a_6_), .ZN(n585) );
  INV_X1 U822 ( .A(b_5_), .ZN(n601) );
  NAND2_X1 U823 ( .A1(n595), .A2(n835), .ZN(n834) );
  INV_X1 U824 ( .A(n791), .ZN(n835) );
  INV_X1 U825 ( .A(n650), .ZN(n595) );
  NAND2_X1 U826 ( .A1(n791), .A2(n650), .ZN(n832) );
  NAND2_X1 U827 ( .A1(b_5_), .A2(a_5_), .ZN(n650) );
  NAND2_X1 U828 ( .A1(n836), .A2(n837), .ZN(n791) );
  NAND2_X1 U829 ( .A1(n838), .A2(n839), .ZN(n837) );
  XNOR2_X1 U830 ( .A(n840), .B(n841), .ZN(n803) );
  XOR2_X1 U831 ( .A(n614), .B(n842), .Z(n840) );
  XNOR2_X1 U832 ( .A(n843), .B(n844), .ZN(n807) );
  XNOR2_X1 U833 ( .A(n845), .B(n846), .ZN(n844) );
  XOR2_X1 U834 ( .A(n847), .B(n848), .Z(n769) );
  XOR2_X1 U835 ( .A(n849), .B(n850), .Z(n848) );
  XOR2_X1 U836 ( .A(n851), .B(n852), .Z(n761) );
  XNOR2_X1 U837 ( .A(n853), .B(n854), .ZN(n851) );
  XOR2_X1 U838 ( .A(n855), .B(n856), .Z(n553) );
  INV_X1 U839 ( .A(n857), .ZN(n560) );
  NAND2_X1 U840 ( .A1(n562), .A2(n561), .ZN(n857) );
  XOR2_X1 U841 ( .A(n692), .B(n691), .Z(n561) );
  XNOR2_X1 U842 ( .A(n686), .B(n858), .ZN(n691) );
  XNOR2_X1 U843 ( .A(n687), .B(n683), .ZN(n858) );
  NOR2_X1 U844 ( .A1(n688), .A2(n644), .ZN(n683) );
  NAND2_X1 U845 ( .A1(n859), .A2(n860), .ZN(n687) );
  NAND2_X1 U846 ( .A1(n861), .A2(n862), .ZN(n860) );
  INV_X1 U847 ( .A(n863), .ZN(n862) );
  NOR2_X1 U848 ( .A1(n864), .A2(n865), .ZN(n863) );
  NAND2_X1 U849 ( .A1(n864), .A2(n865), .ZN(n859) );
  XOR2_X1 U850 ( .A(n866), .B(n867), .Z(n686) );
  XOR2_X1 U851 ( .A(n516), .B(n868), .Z(n867) );
  NAND2_X1 U852 ( .A1(n869), .A2(n870), .ZN(n692) );
  NAND2_X1 U853 ( .A1(n871), .A2(n872), .ZN(n870) );
  INV_X1 U854 ( .A(n873), .ZN(n872) );
  NOR2_X1 U855 ( .A1(n874), .A2(n875), .ZN(n873) );
  NAND2_X1 U856 ( .A1(n875), .A2(n874), .ZN(n869) );
  NOR2_X1 U857 ( .A1(n876), .A2(n856), .ZN(n562) );
  XOR2_X1 U858 ( .A(n877), .B(n878), .Z(n856) );
  INV_X1 U859 ( .A(n871), .ZN(n878) );
  XNOR2_X1 U860 ( .A(n879), .B(n864), .ZN(n871) );
  XNOR2_X1 U861 ( .A(n880), .B(n881), .ZN(n864) );
  XOR2_X1 U862 ( .A(n882), .B(n883), .Z(n880) );
  XNOR2_X1 U863 ( .A(n865), .B(n861), .ZN(n879) );
  NOR2_X1 U864 ( .A1(n508), .A2(n644), .ZN(n861) );
  INV_X1 U865 ( .A(b_2_), .ZN(n644) );
  NOR2_X1 U866 ( .A1(n884), .A2(n885), .ZN(n865) );
  NOR2_X1 U867 ( .A1(n886), .A2(n887), .ZN(n885) );
  INV_X1 U868 ( .A(n528), .ZN(n887) );
  NOR2_X1 U869 ( .A1(n888), .A2(n889), .ZN(n886) );
  INV_X1 U870 ( .A(n890), .ZN(n884) );
  NAND2_X1 U871 ( .A1(n888), .A2(n889), .ZN(n890) );
  XOR2_X1 U872 ( .A(n875), .B(n874), .Z(n877) );
  NAND2_X1 U873 ( .A1(n891), .A2(n892), .ZN(n874) );
  NAND2_X1 U874 ( .A1(n893), .A2(n894), .ZN(n892) );
  INV_X1 U875 ( .A(n895), .ZN(n894) );
  NOR2_X1 U876 ( .A1(n896), .A2(n897), .ZN(n895) );
  NAND2_X1 U877 ( .A1(n897), .A2(n896), .ZN(n891) );
  NOR2_X1 U878 ( .A1(n688), .A2(n632), .ZN(n875) );
  INV_X1 U879 ( .A(n855), .ZN(n876) );
  NAND2_X1 U880 ( .A1(n898), .A2(n899), .ZN(n855) );
  NAND2_X1 U881 ( .A1(n758), .A2(n900), .ZN(n899) );
  NAND2_X1 U882 ( .A1(n901), .A2(n757), .ZN(n900) );
  INV_X1 U883 ( .A(n902), .ZN(n757) );
  NOR2_X1 U884 ( .A1(n688), .A2(n656), .ZN(n758) );
  NAND2_X1 U885 ( .A1(n755), .A2(n902), .ZN(n898) );
  NAND2_X1 U886 ( .A1(n903), .A2(n904), .ZN(n902) );
  NAND2_X1 U887 ( .A1(n854), .A2(n905), .ZN(n904) );
  NAND2_X1 U888 ( .A1(n852), .A2(n853), .ZN(n905) );
  NOR2_X1 U889 ( .A1(n508), .A2(n656), .ZN(n854) );
  INV_X1 U890 ( .A(n906), .ZN(n903) );
  NOR2_X1 U891 ( .A1(n852), .A2(n853), .ZN(n906) );
  NOR2_X1 U892 ( .A1(n907), .A2(n908), .ZN(n853) );
  INV_X1 U893 ( .A(n909), .ZN(n908) );
  NAND2_X1 U894 ( .A1(n850), .A2(n910), .ZN(n909) );
  NAND2_X1 U895 ( .A1(n849), .A2(n847), .ZN(n910) );
  NOR2_X1 U896 ( .A1(n645), .A2(n656), .ZN(n850) );
  NOR2_X1 U897 ( .A1(n847), .A2(n849), .ZN(n907) );
  NOR2_X1 U898 ( .A1(n911), .A2(n912), .ZN(n849) );
  INV_X1 U899 ( .A(n913), .ZN(n912) );
  NAND2_X1 U900 ( .A1(n846), .A2(n914), .ZN(n913) );
  NAND2_X1 U901 ( .A1(n843), .A2(n845), .ZN(n914) );
  NOR2_X1 U902 ( .A1(n631), .A2(n656), .ZN(n846) );
  INV_X1 U903 ( .A(b_4_), .ZN(n656) );
  INV_X1 U904 ( .A(a_3_), .ZN(n631) );
  NOR2_X1 U905 ( .A1(n843), .A2(n845), .ZN(n911) );
  NAND2_X1 U906 ( .A1(n915), .A2(n916), .ZN(n845) );
  NAND2_X1 U907 ( .A1(n841), .A2(n917), .ZN(n916) );
  INV_X1 U908 ( .A(n918), .ZN(n917) );
  NOR2_X1 U909 ( .A1(n614), .A2(n842), .ZN(n918) );
  XOR2_X1 U910 ( .A(n919), .B(n920), .Z(n841) );
  XNOR2_X1 U911 ( .A(n921), .B(n922), .ZN(n920) );
  NAND2_X1 U912 ( .A1(n842), .A2(n614), .ZN(n915) );
  NAND2_X1 U913 ( .A1(b_4_), .A2(a_4_), .ZN(n614) );
  INV_X1 U914 ( .A(n923), .ZN(n842) );
  NAND2_X1 U915 ( .A1(n829), .A2(n924), .ZN(n923) );
  NAND2_X1 U916 ( .A1(n828), .A2(n830), .ZN(n924) );
  NAND2_X1 U917 ( .A1(n836), .A2(n925), .ZN(n830) );
  NAND2_X1 U918 ( .A1(b_4_), .A2(a_5_), .ZN(n925) );
  INV_X1 U919 ( .A(n926), .ZN(n836) );
  NOR2_X1 U920 ( .A1(n922), .A2(n927), .ZN(n828) );
  INV_X1 U921 ( .A(n928), .ZN(n927) );
  NAND2_X1 U922 ( .A1(n929), .A2(n930), .ZN(n928) );
  NAND2_X1 U923 ( .A1(n926), .A2(a_5_), .ZN(n829) );
  NOR2_X1 U924 ( .A1(n839), .A2(n838), .ZN(n926) );
  NAND2_X1 U925 ( .A1(b_4_), .A2(a_6_), .ZN(n838) );
  NAND2_X1 U926 ( .A1(b_3_), .A2(a_7_), .ZN(n839) );
  XNOR2_X1 U927 ( .A(n931), .B(n932), .ZN(n843) );
  XOR2_X1 U928 ( .A(n933), .B(n934), .Z(n931) );
  XOR2_X1 U929 ( .A(n935), .B(n936), .Z(n847) );
  XOR2_X1 U930 ( .A(n937), .B(n646), .Z(n935) );
  XOR2_X1 U931 ( .A(n938), .B(n939), .Z(n852) );
  XNOR2_X1 U932 ( .A(n940), .B(n941), .ZN(n938) );
  INV_X1 U933 ( .A(n901), .ZN(n755) );
  XOR2_X1 U934 ( .A(n893), .B(n942), .Z(n901) );
  XNOR2_X1 U935 ( .A(n896), .B(n897), .ZN(n942) );
  NOR2_X1 U936 ( .A1(n508), .A2(n632), .ZN(n897) );
  NAND2_X1 U937 ( .A1(n943), .A2(n944), .ZN(n896) );
  NAND2_X1 U938 ( .A1(n939), .A2(n945), .ZN(n944) );
  INV_X1 U939 ( .A(n946), .ZN(n945) );
  NOR2_X1 U940 ( .A1(n941), .A2(n940), .ZN(n946) );
  XNOR2_X1 U941 ( .A(n947), .B(n948), .ZN(n939) );
  XOR2_X1 U942 ( .A(n949), .B(n950), .Z(n948) );
  NAND2_X1 U943 ( .A1(n941), .A2(n940), .ZN(n943) );
  NOR2_X1 U944 ( .A1(n951), .A2(n952), .ZN(n940) );
  NOR2_X1 U945 ( .A1(n953), .A2(n626), .ZN(n952) );
  INV_X1 U946 ( .A(n646), .ZN(n626) );
  NAND2_X1 U947 ( .A1(b_3_), .A2(a_3_), .ZN(n646) );
  NOR2_X1 U948 ( .A1(n936), .A2(n937), .ZN(n953) );
  INV_X1 U949 ( .A(n954), .ZN(n951) );
  NAND2_X1 U950 ( .A1(n936), .A2(n937), .ZN(n954) );
  NOR2_X1 U951 ( .A1(n955), .A2(n956), .ZN(n937) );
  INV_X1 U952 ( .A(n957), .ZN(n956) );
  NAND2_X1 U953 ( .A1(n932), .A2(n958), .ZN(n957) );
  NAND2_X1 U954 ( .A1(n933), .A2(n934), .ZN(n958) );
  XNOR2_X1 U955 ( .A(n959), .B(n960), .ZN(n932) );
  NAND2_X1 U956 ( .A1(n961), .A2(n962), .ZN(n959) );
  NOR2_X1 U957 ( .A1(n934), .A2(n933), .ZN(n955) );
  NOR2_X1 U958 ( .A1(n963), .A2(n964), .ZN(n933) );
  INV_X1 U959 ( .A(n965), .ZN(n964) );
  NAND2_X1 U960 ( .A1(n922), .A2(n966), .ZN(n965) );
  NAND2_X1 U961 ( .A1(n921), .A2(n919), .ZN(n966) );
  NOR2_X1 U962 ( .A1(n929), .A2(n930), .ZN(n922) );
  NAND2_X1 U963 ( .A1(b_3_), .A2(a_6_), .ZN(n929) );
  NOR2_X1 U964 ( .A1(n919), .A2(n921), .ZN(n963) );
  NAND2_X1 U965 ( .A1(n967), .A2(n968), .ZN(n921) );
  NAND2_X1 U966 ( .A1(n969), .A2(n970), .ZN(n968) );
  NAND2_X1 U967 ( .A1(b_2_), .A2(a_6_), .ZN(n969) );
  NAND2_X1 U968 ( .A1(b_3_), .A2(a_5_), .ZN(n919) );
  NAND2_X1 U969 ( .A1(b_3_), .A2(a_4_), .ZN(n934) );
  XOR2_X1 U970 ( .A(n971), .B(n972), .Z(n936) );
  NAND2_X1 U971 ( .A1(n973), .A2(n974), .ZN(n971) );
  NOR2_X1 U972 ( .A1(n645), .A2(n632), .ZN(n941) );
  INV_X1 U973 ( .A(b_3_), .ZN(n632) );
  XNOR2_X1 U974 ( .A(n888), .B(n975), .ZN(n893) );
  XOR2_X1 U975 ( .A(n528), .B(n889), .Z(n975) );
  NAND2_X1 U976 ( .A1(n976), .A2(n977), .ZN(n889) );
  NAND2_X1 U977 ( .A1(n978), .A2(n949), .ZN(n977) );
  NAND2_X1 U978 ( .A1(b_2_), .A2(a_3_), .ZN(n949) );
  NAND2_X1 U979 ( .A1(n947), .A2(n950), .ZN(n978) );
  INV_X1 U980 ( .A(n979), .ZN(n976) );
  NOR2_X1 U981 ( .A1(n950), .A2(n947), .ZN(n979) );
  XOR2_X1 U982 ( .A(n980), .B(n981), .Z(n947) );
  XOR2_X1 U983 ( .A(n982), .B(n983), .Z(n980) );
  NAND2_X1 U984 ( .A1(n973), .A2(n984), .ZN(n950) );
  NAND2_X1 U985 ( .A1(n972), .A2(n974), .ZN(n984) );
  NAND2_X1 U986 ( .A1(n985), .A2(n986), .ZN(n974) );
  NAND2_X1 U987 ( .A1(b_2_), .A2(a_4_), .ZN(n986) );
  INV_X1 U988 ( .A(n987), .ZN(n985) );
  XNOR2_X1 U989 ( .A(n988), .B(n989), .ZN(n972) );
  NOR2_X1 U990 ( .A1(n990), .A2(n991), .ZN(n989) );
  NAND2_X1 U991 ( .A1(a_4_), .A2(n987), .ZN(n973) );
  NAND2_X1 U992 ( .A1(n961), .A2(n992), .ZN(n987) );
  NAND2_X1 U993 ( .A1(n960), .A2(n962), .ZN(n992) );
  NAND2_X1 U994 ( .A1(n967), .A2(n993), .ZN(n962) );
  NAND2_X1 U995 ( .A1(b_2_), .A2(a_5_), .ZN(n993) );
  INV_X1 U996 ( .A(n994), .ZN(n967) );
  XNOR2_X1 U997 ( .A(n995), .B(n996), .ZN(n960) );
  NOR2_X1 U998 ( .A1(n736), .A2(n678), .ZN(n996) );
  INV_X1 U999 ( .A(a_7_), .ZN(n736) );
  NAND2_X1 U1000 ( .A1(n994), .A2(a_5_), .ZN(n961) );
  NOR2_X1 U1001 ( .A1(n930), .A2(n995), .ZN(n994) );
  NAND2_X1 U1002 ( .A1(b_1_), .A2(a_6_), .ZN(n995) );
  NAND2_X1 U1003 ( .A1(b_2_), .A2(a_7_), .ZN(n930) );
  NAND2_X1 U1004 ( .A1(b_2_), .A2(a_2_), .ZN(n528) );
  XOR2_X1 U1005 ( .A(n997), .B(n998), .Z(n888) );
  XNOR2_X1 U1006 ( .A(n999), .B(n1000), .ZN(n998) );
  NOR2_X1 U1007 ( .A1(n670), .A2(n688), .ZN(n664) );
  INV_X1 U1008 ( .A(n1001), .ZN(n670) );
  NAND2_X1 U1009 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
  NAND2_X1 U1010 ( .A1(n1004), .A2(b_0_), .ZN(n1003) );
  NOR2_X1 U1011 ( .A1(n1005), .A2(n508), .ZN(n1004) );
  INV_X1 U1012 ( .A(a_1_), .ZN(n508) );
  NOR2_X1 U1013 ( .A1(n680), .A2(n679), .ZN(n1005) );
  NAND2_X1 U1014 ( .A1(n680), .A2(n679), .ZN(n1002) );
  NAND2_X1 U1015 ( .A1(n1006), .A2(n1007), .ZN(n679) );
  NAND2_X1 U1016 ( .A1(n866), .A2(n1008), .ZN(n1007) );
  NAND2_X1 U1017 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
  NOR2_X1 U1018 ( .A1(n678), .A2(n645), .ZN(n866) );
  INV_X1 U1019 ( .A(a_2_), .ZN(n645) );
  NAND2_X1 U1020 ( .A1(n868), .A2(n516), .ZN(n1006) );
  INV_X1 U1021 ( .A(n1010), .ZN(n516) );
  NAND2_X1 U1022 ( .A1(a_1_), .A2(b_1_), .ZN(n1010) );
  INV_X1 U1023 ( .A(n1009), .ZN(n868) );
  NAND2_X1 U1024 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
  NAND2_X1 U1025 ( .A1(n1013), .A2(n882), .ZN(n1012) );
  NAND2_X1 U1026 ( .A1(b_0_), .A2(a_3_), .ZN(n882) );
  INV_X1 U1027 ( .A(n1014), .ZN(n1013) );
  NOR2_X1 U1028 ( .A1(n881), .A2(n883), .ZN(n1014) );
  NAND2_X1 U1029 ( .A1(n883), .A2(n881), .ZN(n1011) );
  NAND2_X1 U1030 ( .A1(b_1_), .A2(a_2_), .ZN(n881) );
  NOR2_X1 U1031 ( .A1(n1015), .A2(n1016), .ZN(n883) );
  INV_X1 U1032 ( .A(n1017), .ZN(n1016) );
  NAND2_X1 U1033 ( .A1(n997), .A2(n1018), .ZN(n1017) );
  NAND2_X1 U1034 ( .A1(n999), .A2(n1000), .ZN(n1018) );
  NOR2_X1 U1035 ( .A1(n678), .A2(n657), .ZN(n997) );
  INV_X1 U1036 ( .A(a_4_), .ZN(n657) );
  NOR2_X1 U1037 ( .A1(n1000), .A2(n999), .ZN(n1015) );
  NOR2_X1 U1038 ( .A1(n1019), .A2(n1020), .ZN(n999) );
  INV_X1 U1039 ( .A(n1021), .ZN(n1020) );
  NAND2_X1 U1040 ( .A1(n981), .A2(n1022), .ZN(n1021) );
  NAND2_X1 U1041 ( .A1(n983), .A2(n982), .ZN(n1022) );
  NOR2_X1 U1042 ( .A1(n678), .A2(n603), .ZN(n981) );
  INV_X1 U1043 ( .A(a_5_), .ZN(n603) );
  INV_X1 U1044 ( .A(b_0_), .ZN(n678) );
  NOR2_X1 U1045 ( .A1(n982), .A2(n983), .ZN(n1019) );
  NOR2_X1 U1046 ( .A1(n1023), .A2(n990), .ZN(n983) );
  NOR2_X1 U1047 ( .A1(n970), .A2(n991), .ZN(n990) );
  NAND2_X1 U1048 ( .A1(b_1_), .A2(a_7_), .ZN(n970) );
  NOR2_X1 U1049 ( .A1(n988), .A2(n991), .ZN(n1023) );
  NAND2_X1 U1050 ( .A1(b_0_), .A2(a_6_), .ZN(n991) );
  NAND2_X1 U1051 ( .A1(b_1_), .A2(a_5_), .ZN(n988) );
  NAND2_X1 U1052 ( .A1(b_1_), .A2(a_4_), .ZN(n982) );
  NAND2_X1 U1053 ( .A1(b_1_), .A2(a_3_), .ZN(n1000) );
  NOR2_X1 U1054 ( .A1(n688), .A2(n1024), .ZN(n680) );
  INV_X1 U1055 ( .A(b_1_), .ZN(n1024) );
  INV_X1 U1056 ( .A(a_0_), .ZN(n688) );
endmodule

