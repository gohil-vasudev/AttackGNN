module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g18881, g23612, g23652, g73, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29219, g29220, g29221, g30327, g30331,
         g30332, g31656, g31665, g34435, g34788, g34839, g36, g44, g53, g54,
         g56, g57, g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751,
         g6753, g84, g90, g91, g92, g99, test_so10, test_so26, test_so35,
         test_so39, test_so42, test_so44, test_so46, test_so80, test_so86,
         test_so92, test_so100, g34783, n4836, n4896, n4895, n4837, n4921,
         n4920, n2787, n4411, n5045, g559, n4959, g33046, g5057, n5615, g34441,
         g2771, n5544, g33982, g1882, g34007, g2299, g24276, g4040, n5530,
         g30381, g2547, n5782, g30405, g3243, g25604, g452, g30416, g3542,
         g30466, g5232, g25736, g5813, g34617, g33974, g1744, g30505, g5909,
         g33554, g1802, n5536, g30432, g3554, g33064, g6219, n5385, g34881,
         g807, n5479, g6031, g24216, g847, n5709, g24232, n9367, g34733, g4172,
         g34882, g4372, g33026, g3512, g31867, n5471, g25668, g3490, n5454,
         g24344, n5432, g4235, g33966, g1600, g33550, g1714, n5460, g30393,
         g3155, n5366, g29248, g2236, g4571, g4555, g24274, g3698, g33973,
         g1736, g30360, g1968, n5664, g34460, g30494, g5607, g30384, g2657,
         g24340, n5439, g29223, g490, n5708, g26881, g311, n5317, g34252, g772,
         n5334, g30489, g5587, g29301, g6177, n5874, g6377, g33022, g3167,
         n5652, g30496, g5615, g33043, g4567, g29263, g30533, g6287, g24256,
         n5302, g34015, g2563, g34031, g4776, n5707, g34452, g4593, n5303,
         g34646, g6199, g34001, g2295, g25633, g1384, g24259, g1339, n5381,
         g33049, g5180, n5384, g34609, g2844, g31869, g1024, g30490, g30427,
         g3598, g21894, g4264, n5823, g33965, g767, n5333, g34645, g5853,
         g33571, g2089, g34267, g4933, n5878, g26971, g4521, n5752, g34644,
         g5507, g30534, g6291, g33535, g294, n5680, g30498, g25728, g25743,
         g25684, g3813, g25613, g562, g34438, g608, n5475, g24244, g1205,
         n5547, g30439, g3909, g30541, g6259, g30519, g5905, g25621, g921,
         g34807, g2955, g25599, g203, g24235, g34036, g4878, n5283, g30476,
         g5204, g30429, g3606, g32997, g1926, n5510, g33063, g6215, n5651,
         g30424, g3586, g32977, g291, n5679, g34026, g4674, n5440, g30420,
         g3570, g33560, g29226, g676, n5751, g25619, g843, g34455, g4332,
         n5540, g30457, g4153, g33625, g6336, n5592, g34790, g622, n5672,
         g30414, g3506, n5576, g26966, g4558, g25656, g3111, g30390, g25688,
         g34727, g939, g25594, g278, g26963, g4492, g34034, g4864, n5318,
         g33541, g1036, g28093, g24236, g1178, g30404, g3239, g28051, g718,
         g29303, g6195, n5741, g26917, g1135, n5328, g33624, g6395, n5396,
         g24337, g34911, g554, g33963, g496, g34627, g3853, g29282, g5134,
         n5807, g25676, g33013, g2485, n5509, g32981, g925, n5725, g34976,
         n9357, g30483, g5555, g32994, g1798, g28070, g34806, g2941, g30453,
         g3905, g33539, g763, n5332, g30526, g6255, g26951, g4375, g34035,
         g4871, n5443, g34636, g4722, g32978, g590, n5472, g30348, g1632,
         n5836, g24336, n5438, g3100, g24250, g29236, g1437, n5696, g29298,
         g6154, n5747, g1579, g30499, g5567, g33976, g1752, g32996, g1917,
         g30335, g744, n5470, g34637, g4737, n5867, g25694, g30528, g6267,
         g24251, g1442, g30521, g26960, g4477, n5849, g24239, g34259, g4643,
         n5382, g30474, g5264, n5703, g33016, g2610, g34643, g5160, g30510,
         g5933, g29239, g1454, n5866, g26897, g753, g34729, g1296, g34625,
         g3151, g34800, g24353, g6727, n5531, g33029, g3530, n5569, g4104,
         g24253, g1532, g24281, g33997, n9352, g34971, n9351, g34263, g4754,
         n5877, g24237, g1189, g33584, g2287, n5353, g24280, g4273, n5764,
         g26920, g1389, g33548, g29296, g5835, n5663, g30338, g1171, n5363,
         g21895, g4269, n5763, g33588, g2399, n5762, g34041, g4983, n5367,
         g30495, g5611, g29279, g4572, g25655, g3143, n5882, g34795, g2898,
         g24269, g3343, g30403, g3235, g33042, g30419, g3566, g34023, n9348,
         g28090, g4961, g34642, g4927, n5879, g30370, g2259, n5419, g34448,
         g2819, n5609, g26946, g5802, g34610, g2852, g24209, g417, n5358,
         g28047, g681, g24206, g437, g26891, g30504, g5901, g34798, g2886,
         g25669, g3494, n5889, g30480, g5511, n5575, g33027, g3518, n5645,
         g33972, g1604, g25697, g5092, g28099, g4831, g26947, g4382, n5714,
         g24350, g6386, g24210, g479, g30455, g3965, g28084, g33993, g2008,
         g736, g30444, g3933, g33537, g222, g25650, g3050, g25625, g1052,
         g30366, g2122, n5784, g33593, g2465, n5523, g30502, g5889, g33036,
         g4495, g25595, g34462, g33024, g3179, n5390, g33552, g1728, n5352,
         g34014, g2433, g29273, g3835, n5662, g25748, g6187, n5453, g34638,
         g4917, g30341, g1070, g26899, g822, n5422, g30336, g914, n5560, g5339,
         g26940, g4164, g25622, g34447, g2807, n5379, g33613, g4054, n5395,
         g25749, g6191, n5888, g25704, g5077, n5455, g33053, g5523, n5647,
         g3680, g30555, g6637, g25601, g174, g33971, g1682, g26892, g355,
         g1087, g26915, g1105, n5478, g33008, g30538, g6307, g3802, g25750,
         g6159, g30369, g2255, g34446, g2815, n5404, g29230, g911, n5559, g43,
         g33975, g1748, g30497, g5551, g30418, g3558, g25721, g5499, n5885,
         g34622, g30438, g3901, g34266, g4888, n5863, g30540, g6251, g32986,
         g1373, g25648, g33960, g157, n5678, g34442, g2783, n5403, g4281,
         g30421, g3574, g33573, g2112, g34730, g1283, g24205, g10122_Tj, g4297,
         n5698, g32979, g758, n5331, g34025, g4639, n5727, g25763, g6537,
         n5884, g30481, g5543, g30517, g5961, g30539, g6243, g34880, n9340,
         g24242, n5654, g30436, g29265, g3476, n5786, g32990, g1664, g24245,
         g1246, n5756, g30553, g6629, g26907, g246, n6008, g24278, g4049,
         g26955, g24282, g2932, g29276, g4575, g31894, g4098, n5350, g33037,
         g4498, g26894, g528, n5327, g34977, n5477, g25654, g3139, n5447,
         g33962, g34451, g4584, n5539, g34250, g142, n5724, g29295, g5831,
         n5873, g26905, g239, g25629, g1216, n5442, g34792, g2848, g25703,
         g5022, g32983, g1030, g30402, g3231, g25757, g1430, n9336, g33999,
         g2241, g24262, g1564, g25729, g6148, g30558, g6649, g34781, g110,
         g26901, g225, n5597, g26961, g33039, g4504, g33059, g5873, n5388,
         g31899, g5037, n5611, g33007, g2319, n5375, g25720, g5495, n5446,
         g21891, g30462, g5208, g30487, g5579, g33058, g5869, n5649, g24261,
         g1589, n5755, g25730, g5752, g30531, g6279, g30506, g34804, g2975,
         n5750, g25747, g6167, n5430, n5701, g33601, g2599, n5524, g26922,
         g1448, n5343, g29250, g2370, g30459, g5164, n5570, g1333, n5616,
         g33534, g153, n5677, g30543, g6549, n5571, g29275, g4087, n5480,
         g34030, g34980, g2984, g30451, g3961, g25627, g962, n5630, g34657,
         g101, g30552, g6625, g34979, n9332, g30337, g1018, g24254, g24277,
         g4045, g29237, g1467, n5693, g30378, g2461, n5840, g33019, n5300,
         g33623, g5990, n5589, g29235, g1256, n5558, g31902, g5029, n5601,
         g29306, g6519, n5806, g25689, g4169, n5729, g33978, g1816, g26970,
         g4369, g29278, g4578, g34253, g4459, n5765, g29272, g3831, n5872,
         g33595, g2514, g33610, g3288, n5400, g33589, g34605, g2145, n5307,
         g30350, g1700, n5417, g25611, g513, n5548, g2841, n5963, g33619,
         g5297, n5588, g34022, g2763, g34033, g4793, n5368, g34726, g952,
         g31870, g1263, n5674, g33985, g1950, g29283, g5138, n5871, g34003,
         g2307, g25677, g34463, g4664, g33006, g2223, g29292, g5808, n5749,
         g30557, g6645, g33989, g2016, g33033, g3873, n5387, n5699, g34005,
         g2315, g26932, g2811, g30516, g5957, g33575, g2047, g33032, g30486,
         g5575, g34974, n9327, g25678, g3752, g30440, g3917, DFF_480_n1, g1585,
         n5757, g26949, g4388, g30530, g6275, g30542, g6311, g25624, g1041,
         g30383, g33597, g2537, g34598, g26957, g4430, g26967, n9325, g28102,
         g4826, g30524, g6239, g26903, g232, g30475, g5268, g34647, g6545,
         g30377, n9324, g33553, g1772, n5504, g31903, g5052, n5607, g25715,
         g33984, g1890, n5799, g33602, g2629, n5521, g28045, g572, n5337,
         g34603, g2130, g33035, g4108, n5715, g4308, g24208, g475, g990, n5622,
         g31, n5469, g34970, n9322, g24213, g33614, g3990, n5594, g33060,
         g30362, g1992, g33023, g3171, n5603, g26898, g812, n5733, g25618,
         g832, g30518, g5897, g4570, n5702, g26959, g4455, g34801, g2902,
         g26884, g333, g25600, g168, g26933, g28066, g3684, g33612, g3639,
         n5591, g24268, g3338, n5527, g25716, g5406, g26906, g269, g24203,
         g401, g24346, g6040, g24207, g441, g25701, n5690, g29269, g3808,
         n5745, g9, n5468, g34255, g30450, g3957, g30456, g4093, n5340, g32991,
         g1760, n5602, g24348, n5437, g34249, g160, n5843, g30371, g2279,
         n5778, g29268, g3498, n5740, g29224, g586, n5336, g33017, g2619,
         n5508, g30339, g1183, n5599, g33967, g1608, g33559, g1779, g29255,
         g2652, g30368, g2193, n5839, g30375, g2393, n5421, g28052, g661,
         g28089, g4950, g33055, g5535, n5566, g30392, g2834, g30343, g1361,
         g30523, g6235, g24233, g1146, n5851, g33018, g32976, g150, n5676,
         g30349, g1696, g33067, g6555, g26900, g33034, g3881, n5564, g30551,
         g6621, g25667, g3470, n5424, g30452, g3897, g34719, g518, g538,
         g33607, g2606, g26923, g1472, n5290, g24211, g33050, g5188, n5567,
         g24341, g5689, n5529, g24201, g405, g30463, g5216, g6494, g34464,
         g4669, g24243, g996, g24335, g4531, g34611, g2860, g34262, g4743,
         n5876, g30546, g6593, g25591, g4411, g30347, g1413, g30556, g6641, g6,
         g33562, g1936, n5534, g55, g25610, g504, n5519, g33015, g2587, n5372,
         g31896, g4480, g34004, n9314, g30428, g30485, g5571, g30422, g3578,
         g25714, g29294, g5827, n5809, g30423, g3582, g30529, g6271, g34028,
         g4688, n5656, g33587, g2380, g30460, g5196, g30401, g3227, g33990,
         n9312, g29309, g6541, n5739, g30411, g3203, g33546, g1668, n5598,
         g28085, g4760, g26904, g262, g33556, g1840, n5451, g25722, g5467,
         g25605, g460, g33062, g6209, g26893, n5704, g28050, g655, g34626,
         g33583, g2204, g30472, g5256, g34454, g4608, n5274, g34850, g794,
         n5291, g4423, g24272, g3689, n5532, g5685, g24214, g703, n5821,
         g26909, g862, n5682, g30406, g3247, g33569, g2040, n5505, g34628,
         g4146, n5981, g34458, g4633, n5844, g24240, n5304, g34634, g4732,
         g25700, n5689, g29293, g5817, g33009, g2351, n5511, g33603, g2648,
         g24355, g6736, g34268, g4944, n5875, g25691, g4072, g26890, g29264,
         g3466, g28072, g4116, g31900, g5041, n5605, g26956, g4434, g29271,
         g3827, n5808, g29304, g6500, n5748, g29261, g3133, n5661, g28063,
         g3333, g979, n5320, g34027, g4681, g33961, g298, n5675, g33604,
         g32995, g1894, n5374, g34624, g2988, g30415, g3538, g33536, g301,
         g26888, n9306, DFF_709_n1, g28055, g827, n5728, g24238, g33600, g2555,
         n5351, g28105, g5011, g34721, g199, g29307, g6523, n5870, g30345,
         g34453, g4601, n5365, g32980, g854, g29238, g1484, n5865, g34639,
         g4922, g25695, g5080, n5893, g33057, g5863, g26969, g4581, n5670,
         g29253, g2518, g34021, g2567, g26895, g568, n5335, g30413, g3263,
         g30549, g6613, g24347, g25758, g6444, g34808, g2965, g30501, g5857,
         n5573, g33969, n9303, g34440, g890, n5305, g30433, g3562, g21900,
         g26921, g1404, g29270, g3817, n9302, g33038, g4501, g31865, g26926,
         g2724, n5301, g28083, g4704, g34797, g22, g2878, g30478, g5220,
         g34724, g617, n5339, g24212, g26883, g316, g32985, g1277, g25761,
         g6513, n5426, g26886, g336, n5824, g34796, g2882, g32982, g33561,
         g1906, n5503, g26880, g305, n5282, g34975, g8, g26931, g2799, g34641,
         g4912, g34629, g4157, n5983, g33598, g2541, n5461, g33576, g2153,
         n5356, g34720, g550, g26902, g255, g29244, g30468, g5240, g26924,
         g1478, n5289, g33031, g3863, g29245, g1959, g29266, g3480, n5868,
         g30559, g6653, g34794, g2864, g28087, g4894, g30435, g3857, n5572,
         g25609, g28057, g1002, g34439, g776, n5330, g28, n5324, g1236, g34260,
         g4646, n5712, g33012, g2476, g32989, g1657, n5525, g34006, g2375, g63,
         g358, g26910, g896, n5431, g28043, g33021, g3161, g29251, g2384,
         n5700, g34456, g4616, n5608, g26968, g4561, g33991, g2024, g3451,
         g26930, g2795, g34599, g613, n5474, g28082, g4527, g33557, g1844,
         g30511, g5937, g33045, g30379, g2523, g24267, n5436, g34020, g2643,
         g24249, g1489, n5850, g25592, g30382, n9295, g29285, g5156, n5734,
         n5526, n9294, g25662, g21896, g33563, g1955, g33622, g33582, g2273,
         n5458, g28086, g4771, g25744, g6098, g29262, g3147, n5738, g24270,
         g3347, g33581, g2269, g191, g24266, g2712, g34849, g626, n5288,
         g33618, g2729, g5357, n5393, g34038, g34032, g4709, n5518, g34803,
         g2927, g34459, g4340, n5653, g30509, g5929, g34640, g4907, g28069,
         g4035, g21899, g2946, g31868, g918, n5673, g26938, g4082, g25756,
         g30363, g30334, g577, n5294, g33970, g1620, g30391, g2831, g25615,
         g667, g33540, g930, n5731, g30445, g3937, g25617, g817, n5822, g24247,
         g1249, g24215, g837, n5562, g33964, g599, n5550, g25719, g5475, n5425,
         g29228, g30514, g5949, g33627, g6682, n5590, g24231, g904, g34615,
         g2873, n5488, g30356, g1854, n5785, g25696, g5084, n5681, g30493,
         g5603, n5726, g33594, g2495, n5522, g34009, g2437, g30365, g2102,
         n5666, g33004, g2208, g34018, g25685, g4064, n5416, g34040, g4899,
         n5517, g25639, g2719, n5465, g34029, g4785, n5361, g30488, g5583,
         g34600, g781, n5551, g29300, g6173, n5810, g34802, g2917, g25614,
         g686, g28058, g1252, n5554, g29225, g671, g33580, g30532, g6283,
         DFF_909_n1, g33054, g5527, n5389, g26962, g4489, g33564, g1974, n5450,
         g32984, g1270, n5716, g34039, g4966, n5706, g33065, g6227, n5568,
         g30443, g3929, g29291, g5503, n5737, g24279, g30508, g5925, g29232,
         g1124, n5692, g34269, g4955, n5614, g30464, g5224, g33988, g2012,
         g30522, g6203, n5574, g25708, g5120, g30374, g2389, g26953, g4438,
         g34008, g2429, g34444, g2787, n5610, g34731, g33606, g2675, n5457,
         g24334, g34265, g4836, n5713, g30340, g1199, g24257, n5401, g30482,
         g5547, g34604, g2138, n5275, g33591, g2338, g30525, g6247, g26929,
         g2791, g30448, g34602, g1291, n2549, g30513, g5945, g30469, g5244,
         g33608, g2759, g33626, g6741, n5398, g34725, g785, n5293, g30342,
         g1259, n5553, g29267, g3484, n5668, g25593, g209, n5595, g30548,
         g6609, g33052, g5517, g34012, g2449, g34017, n9281, DFF_961_n1,
         g24263, g2715, n5299, g26912, g936, n5557, g30364, g2098, g34254,
         g4462, n5671, g34251, g604, n5473, g30560, g6589, g33983, n9280,
         g24204, g429, g33980, g1870, g34631, g29243, g1825, g25623, g1008,
         n5321, g26950, g4392, n5710, g30431, g3546, g30467, g5236, g30353,
         g1768, n5834, g34467, g4854, g30442, g3925, g29305, g6509, g25616,
         g732, n5732, g29252, g2504, g4519, g4520, g33003, g2185, n5376,
         g34613, g37, g4031, g33570, g2070, n5535, g34734, g4176, g24275,
         n5435, g4405, g872, g29302, g6181, n5667, g24349, g34264, g4765,
         n5613, g30484, g5563, g25634, g1395, g33567, g1913, g33585, g2331,
         n5513, g30527, g6263, g34978, n9276, g30447, g3945, g347, n5860,
         g34256, g4473, g25630, g1266, g29290, g5489, n5660, g29227, g31872,
         g2748, n5516, g29287, g5471, g31897, g4540, g6723, g30562, g6605,
         g34011, n9274, g33996, g2173, g21898, g33014, g2491, g34465, g4849,
         g33995, g2169, g30372, n9273, g30545, g30389, g33590, g2407, n5459,
         g34616, g2868, g26927, g2767, g32992, g1783, n5596, g25631, g1312,
         n5466, g30477, g5212, g34632, g4245, g28046, g645, g4291, g26896,
         n5657, g25602, g26916, g1129, n5329, g33578, g2227, n5538, g33579,
         g2246, g30354, g1830, g30425, g3590, g24200, g392, g33544, g1592,
         n5362, g25764, g6505, g24246, g1221, g30507, g5921, g26889, g30333,
         g218, g32998, g1932, g32987, g1624, n5370, g25702, g5062, g29286,
         g5462, n5744, g34606, g2689, g33070, g6573, n5563, g29240, g1677,
         g32999, g2028, n5371, g33605, g2671, g24255, g26945, g33558, g1848,
         n5464, g25699, n5669, g29289, g5485, n5869, g30388, g2741, n5349,
         n5482, g29254, g2638, g28074, g4122, g34450, g4322, n5506, g30512,
         g5941, g33572, g2108, n5452, g25, g33551, g33538, g595, n5476, g33005,
         g2217, n5512, g24248, n9267, g33002, g2066, g24234, g1152, n5618,
         g30471, g5252, g34000, g2165, g34016, g2571, g33048, g5176, n5650,
         g25628, g26934, g2827, g34468, g4859, g24202, g424, g33542, g1274,
         n5730, n9265, n6006, g34445, g2803, n5545, g33555, g1821, g34013,
         g2509, g28091, g5073, g26919, n5556, g30554, g6633, g29281, g5124,
         g30537, g6303, g28092, g5069, g34732, g2994, n5634, g28049, g650,
         g33545, g1636, n5549, g30441, g3921, g29247, g24354, g6732, g25636,
         g1306, n5796, g26914, g1061, g25670, g3462, g33998, g2181, g25626,
         g956, n5341, g33977, g1756, g29297, g5849, n5736, g28071, g4112,
         g30387, n9262, g33577, g2197, n5514, g33592, g26913, g1046, g28044,
         g482, n5820, g26948, g4401, g30344, g1514, n5364, g26885, g329, n5766,
         g33069, g6565, n5386, g34621, g2950, g28059, g1345, g25762, g6533,
         n5445, g34633, g4727, g24352, g26925, g1536, g30446, g3941, g25597,
         g370, g24342, g5694, g30357, g1858, g26908, g446, g30399, g3219,
         g29242, g1811, g30547, g6601, g34010, g2441, g33986, g1874, g34257,
         g30544, g6581, g30561, g6597, g5008, g30430, g3610, g34799, g2890,
         g33565, g1978, g33968, g1612, g34843, g112, g34793, g2856, g33566,
         g1982, n5462, g30465, g28073, g4119, g24351, g6390, g30346, g1542,
         g21893, g4258, g4818, g31904, g5033, g34635, g4717, g25637, g1554,
         n5768, g29274, g3849, n5735, g30396, g3199, g25735, g34037, g4975,
         n5360, g34791, g790, n5292, g30520, g5913, g30358, g1902, n5837,
         g29299, g6163, g25690, g4125, g28096, g4821, n5880, g28088, g4939,
         g24241, n5392, g30397, g3207, g4483, g30409, g29284, g5142, n5658,
         g30470, g5248, g30367, g2126, g24273, g3694, g29288, g5481, n5805,
         g30359, g1964, g25698, g5097, n5753, g30398, g3215, n9255, n6005,
         g26952, g4427, g26928, g2779, n5694, g26954, g30351, g1720, n5780,
         g31871, g1367, g5112, g19, g26939, g4145, g33994, g2161, g25596, g376,
         n5633, g33586, g2361, n5537, g21901, DFF_1234_n1, g31866, g582, n5552,
         g33000, g2051, g26918, g1193, g30373, g2327, n5841, g28056, g907,
         n5555, g34601, g947, n5286, g30355, g1834, n5665, g30426, g3594,
         g34805, g2999, g34002, g2303, g28053, g29229, g723, n5826, g33620,
         g5703, n5397, g34722, g546, g33599, g2472, g30515, g5953, g25649,
         g33979, g1740, g30417, g3550, g25683, g3845, n5886, g33574, g2116,
         n5463, g30410, g30454, g3913, g34024, g33547, g1687, g30386, g2681,
         n5777, g33596, g2533, n5761, g26887, g324, n5827, g34607, g2697,
         n5308, g31895, g4417, g33068, g6561, n5646, g29233, g1141, n5691,
         g24258, n5655, g30376, g33549, g1710, g29308, g6527, n5659, g30408,
         g3255, g29241, g1691, g34620, g2936, g33621, g5644, n5593, g25707,
         g5152, n5883, g24339, g5352, g34443, g2775, n5378, g34619, g2922,
         g29234, g30503, g5893, g30550, g6617, g33001, g2060, n5507, g33040,
         g4512, g30492, g5599, g25664, g3401, g26944, g4366, g34614, g29260,
         g3129, n5861, g33047, g5170, g24298, g25733, g5821, n5429, g30536,
         g6299, g29246, g2079, g34261, g4698, n5862, g33611, g3703, n5399,
         g25638, g1559, n5441, g34728, n9247, g29222, g411, g25742, g30449,
         g3953, g34608, g2704, n5377, g24345, g6035, n5528, n9245, g25635,
         g1300, n5483, g25686, g4057, n5711, g30461, g5200, g34466, g4843,
         g31901, g5046, n5578, g29249, g2250, g26882, n5456, g33041, g33011,
         g2453, n5373, g25734, g5841, n5449, n5705, g34618, g2912, g33010,
         g2357, g31864, g164, n5561, g34630, g4253, n5484, g31898, g5016,
         n5369, g25653, g3119, n5423, g25632, g1351, n5322, g32988, g33616,
         g29280, g5115, n5743, g33609, g3352, n5604, g30563, g6657, g33044,
         g4552, g30437, g3893, g30412, g3211, g30491, g5595, g30434, g3614,
         g34612, g29259, g3125, n5781, g25681, g3821, n5428, g25687, g4141,
         n5612, g33617, g30479, g5272, g29256, g2735, n5600, g28054, g728,
         g30535, g6295, g30385, g2661, n5418, g30361, g1988, n5783, g25705,
         g24260, g1548, n5546, g29257, g3106, n5742, g34461, g4659, g34258,
         g4358, n5348, g32993, g1792, n5359, g33992, g2084, g30394, g3187,
         g34449, g4311, n5323, g34019, g2583, g18597, n9240, g29231, g1094,
         n5697, g25682, g21897, g4284, g30395, g3191, g21892, g4239, g4180,
         n5380, g28048, g691, n5520, g34723, g534, g25598, g385, n5632, g33987,
         g2004, g30380, g2527, n5420, g5456, g26965, n6007, g25706, g30458,
         g4507, n5846, g24338, g5348, g30400, g3223, g34623, g2970, g24343,
         g5698, g30473, g5260, g24252, g1521, n5577, g33028, g3522, n5383,
         g29258, g3115, g30407, g3251, g26958, g34457, g33568, g1996, n5355,
         g25663, g26964, g4515, g34735, g4300, g30352, n9236, g33543, g1379,
         g24271, n5433, g33981, g1878, g30500, g5619, g34649, g71, g29277,
         g25612, n5287, g28060, n2505, n2499, n2461, n2396, n2668, g72, n5960,
         n4689, n5961, n4708, n3593, n3595, n3574, n3576, n3517, n3519, n3628,
         n3630, n3555, n3557, n3646, n3648, n3536, n3538, n3611, n3613, n3006,
         n3765, n3525, n3635, n4888, n3550, n2595, n2527, n3524, n3005, n3623,
         n3549, n3003, n3007, n3569, n3606, n3588, n3165, n3799, n3033, n3622,
         n3587, n3586, n3605, n3604, n3568, n3567, n3548, n3512, n3511, n3531,
         n3530, n3641, n3640, n3131, n3111, n3907, n3773, n3807, n3950, n3841,
         n3983, n3874, n4014, n4537, n4201, n3745, n3684, n3274, n2982, n2706,
         n2649, n2556, n2509, n2487, n2427, n2423, n4826, n2421, n4172, n4173,
         n4190, n4191, n4388, n4210, n3951, n3404, n3774, n3424, n3842, n3414,
         n3808, n3444, n3908, n3489, n3984, n3434, n3875, n3500, n4015, n3446,
         n3914, n3406, n3780, n3481, n3957, n3426, n3848, n3491, n3990, n3416,
         n3814, n3436, n3881, n3502, n4022, n3501, n4027, n3407, n3785, n3482,
         n3962, n3427, n3853, n3437, n3886, n3417, n3819, n3492, n3995, n3447,
         n3919, n3682, n3272, n2980, n2704, n2647, n2554, n2507, n2485, n2425,
         n2419, n2405, n2760, n2552, n4946, n4198, n2404, n4962, n4948, n2726,
         n2727, n3195, n3116, n4945, n4525, n4518, n3281, n3277, n3276, n2989,
         n2991, n3687, n2710, n2707, n3174, n3362, n3676, n2644, n3146, n3115,
         n3833, n3023, n3933, n3729, n4723, n3664, n3662, n3673, n3671, n2607,
         n3506, n2790, n4490, n4178, n4514, n4196, n3736, n3741, n2598, n4814,
         n4519, n2594, n3084, n2590, n4722, n3125, n3105, n3145, n3164, n3910,
         n3776, n3877, n3810, n4017, n3953, n3986, n3844, n3770, n3904, n3804,
         n3947, n3838, n3871, n3980, n4020, n3495, n3945, n3836, n3768, n3869,
         n3978, n3802, n3902, n2422, n5121, n4037, n4034, n4039, n3972, n3969,
         n3929, n3926, n3863, n3860, n4003, n4002, n4032, n4035, n3797, n3792,
         n3790, n3795, n3891, n3893, n3827, n3826, n3896, n4007, n3931, n3793,
         n3924, n3831, n3829, n3927, n3974, n3898, n3970, n4000, n3865, n3861,
         n3824, n3894, n3967, n3858, n4005, n3395, n4956, n5026, n3941, n3733,
         n4798, n4805, n4175, n4193, n3738, n4721, n4523, n4524, n4526, n2573,
         n2577, n2563, n2567, n4938, n4940, n4913, n4915, n4714, n4516, n4517,
         n5111, n3730, n3121, n3180, n4305, n4283, n2608, n4447, n4448, n4402,
         n4403, n4425, n4426, n4436, n4437, n4391, n4392, n4379, n4380, n4414,
         n4415, n4458, n4459, n5016, n5014, n3064, n3065, n4535, n5112, n3675,
         counter_31, counter_30, counter_29, counter_28, counter_27,
         counter_26, counter_25, counter_24, counter_23, counter_22,
         counter_21, counter_20, counter_19, counter_18, counter_17,
         counter_16, counter_15, counter_14, counter_13, counter_12,
         counter_11, counter_10, counter_9, counter_8, counter_7, counter_6,
         counter_5, counter_4, counter_3, counter_2, counter_1, counter_0,
         carry_31, carry_30, carry_29, carry_28, carry_27, carry_26, carry_25,
         carry_24, carry_23, carry_22, carry_21, carry_20, carry_19, carry_18,
         carry_17, carry_16, carry_15, carry_14, carry_13, carry_12, carry_11,
         carry_10, carry_9, carry_8, carry_7, carry_6, carry_5, carry_4,
         carry_3, carry_2, N31, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14,
         N15, N23, N24, N25, N26, N2, N3, N4, N16, N17, N18, N19, N20, N21,
         N22, N27, N28, N29, N30, N1, N32, n37, n87, n73, n86, n85, n84, n83,
         n82, n81, n80, n79, n78, n77, n76, n75, n74, n58, n59, n60, n61, n62,
         n63, n64, Trigger_out, n65, n66, n67, n68, n69, n70, n71, n72, n44,
         n53, n108, n120, g33959, n173, n174, g33533, n251, n286, n290, n333,
         n346, n515, n516, n646, n658, n662, n725, n727, n735, n736, n760,
         n879, n1075, g25167, n1156, n1282, n1284, n1285, n1287, n1289, n1340,
         n1643, n1645, n1698, n10006, n10007, n10008, n10010, n10011, n10012,
         n10018, n10019, n10021, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10035, n10036, n10037, n10041, n10042, n10045,
         n10046, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10057, n10058, n10059, n10060, n10061, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10074, n10076,
         n10077, n10078, n10080, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10104,
         n10109, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10121, n10122, n10123, n10124, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10152, n10153, n10155,
         n10156, n10159, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10233, n10235, n10237, n10239, n10241, n10243, n10245,
         n10246, n10248, n10250, n10252, n10254, n10255, n10257, n10259,
         n10261, n10263, n10264, n10265, n10266, n10267, n10268, n10270,
         n10271, n10274, n10275, n10276, n10302, n10305, n10306, n10308,
         n10310, n10312, n10313, n10315, n10317, n10319, n10320, n10323,
         n10324, n10327, n10328, n10331, n10332, n10335, n10338, n10339,
         n10342, n10343, n10346, n10347, n10350, n10351, n10352, n10353,
         n10356, n10357, n10360, n10361, n10364, n10365, n10368, n10369,
         n10372, n10373, n10376, n10377, n10380, n10381, n10385, n10386,
         n10387, n10388, n10389, n10391, n10392, n10397, n10398, n10399,
         n10400, n10401, n10402, n10413, n10416, n10417, n10418, n10419,
         n10421, n10422, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10452, n10455, n10456,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10481, n10482, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10519, n10520, n10521, n10522, n10523, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         g32975, n10537, n10538, n10539, n10540, n10541, n10542, g31860,
         n10544, g31862, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         U5353_n1, U5355_n1, U5961_n1, U5962_n1, U5963_n1, U5964_n1, U5965_n1,
         U5966_n1, U5967_n1, U5968_n1, U6100_n1, U6211_n1, U6212_n1, U6213_n1,
         U6214_n1, U6215_n1, U6216_n1, U6217_n1, U6218_n1, U6279_n1, U6280_n1,
         U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1, U6286_n1, U6287_n1,
         U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1, U6338_n1, U6341_n1,
         U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1,
         U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1,
         U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1,
         U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1,
         U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6417_n1,
         U6446_n1, U6465_n1, U6497_n1, U6523_n1, U6542_n1, U6552_n1, U6553_n1,
         U6554_n1, U6555_n1, U6556_n1, U6559_n1, U6560_n1, U6561_n1, U6570_n1,
         U6911_n1, U6912_n1, U6917_n1, U6926_n1, U6927_n1, U6929_n1, U6931_n1,
         U6932_n1, U6933_n1, U6934_n1, U6935_n1, U6936_n1, U6937_n1, U6938_n1,
         U6939_n1, U6940_n1, U6941_n1, U6944_n1, U6950_n1, U6954_n1, U6955_n1,
         U6956_n1, U6957_n1, U7174_n1, U7248_n1, U7249_n1, U7402_n1, U7405_n1,
         U7413_n1, U7416_n1, U7427_n1, U7438_n1, U7449_n1, U7455_n1, U7464_n1,
         U7467_n1, U7482_n1, U7492_n1, U7513_n1, U7516_n1, U7549_n1, U7561_n1,
         U7574_n1, U7577_n1, U7585_n1, U7595_n1, U7614_n1, U7621_n1, U7629_n1,
         U7636_n1, U7639_n1, U7649_n1, U7652_n1, U7668_n1, U7673_n1, U7690_n1,
         U7707_n1, U7712_n1, U7792_n1, U7794_n1, U7895_n1, U7897_n1, U7977_n1,
         U8034_n1, U8036_n1, U8050_n1, U8055_n1, U8060_n1, U8070_n1, U8074_n1,
         U8088_n1, U8112_n1, U8113_n1, U8147_n1, U8165_n1, U8185_n1, U8192_n1,
         U8210_n1, U8223_n1, U8224_n1, U8281_n1, U8307_n1, U8974_n1, U8975_n1,
         U9065_n1, U9070_n1, U9075_n1, U9076_n1, U9080_n1, U9084_n1, U9085_n1,
         U9086_n1, U9090_n1, U9098_n1, U9099_n1, U9101_n1, U9107_n1, U9111_n1,
         U9116_n1, U9120_n1, U9124_n1, U9128_n1, U9132_n1, U9136_n1, U9315_n1,
         U9453_n1, U9825_n1, U9886_n1, U9927_n1, U9953_n1, U9957_n1, U9958_n1,
         U9968_n1, U9972_n1, U9992_n1, U10314_n1, U10318_n1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g34597 = 1'b0;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g29218 = g18881;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g24167 = g73;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20557 = g29213;
  assign g20652 = g29214;
  assign g20901 = g29215;
  assign g21176 = g29216;
  assign g21270 = g29217;
  assign g20654 = g29219;
  assign g21245 = g29220;
  assign g21292 = g29221;
  assign g23002 = g30327;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g31521 = g34435;
  assign g33894 = g34788;
  assign g34956 = g34839;
  assign g21698 = g36;
  assign g24185 = g44;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18101 = g6746;
  assign g18097 = g6747;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18100 = g6751;
  assign g18092 = g6753;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g31861 = test_so10;
  assign g25219 = test_so10;
  assign g13881 = test_so26;
  assign g9615 = test_so35;
  assign g8785 = test_so39;
  assign g8291 = test_so42;
  assign g17316 = test_so44;
  assign g8178 = test_so46;
  assign g12470 = test_so80;
  assign g11447 = test_so86;
  assign g9682 = test_so92;
  assign g29210 = test_so100;
  assign g20049 = test_so100;
  assign g24166 = g72;
  assign g28753 = g33959;
  assign g27831 = g33533;
  assign g31863 = g25167;
  assign g26801 = g32975;
  assign g25114 = g31860;
  assign g25259 = g31862;

  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(n10597), .CLK(n10933), 
        .Q(g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(n10605), .CLK(n10941), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(n10697), .CLK(n11033), .Q(
        g1882) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(n10652), .CLK(n10988), .Q(
        g2299) );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(n10635), .CLK(n10971), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(n10663), .CLK(n10999), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(n10692), .CLK(n11028), .Q(
        g559) );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(n10622), .CLK(n10958), .Q(
        g3243) );
  SDFFX1 DFF_10_Q_reg ( .D(g25604), .SI(g3243), .SE(n10616), .CLK(n10952), .Q(
        g452), .QN(n10275) );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(n10691), .CLK(n11027), .Q(
        g3542) );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(n10626), .CLK(n10962), .Q(
        g5232) );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(n10665), .CLK(n11001), .Q(
        g5813), .QN(n10102) );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(n10686), .CLK(n11022), .Q(
        test_so1) );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(n10648), .CLK(n10984), 
        .Q(g1744) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(n10678), .CLK(n11014), .Q(
        g5909) );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(n10690), .CLK(n11026), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(n10653), .CLK(n10989), .Q(
        g3554), .QN(n10347) );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(n10653), .CLK(n10989), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(n10623), .CLK(n10959), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(n10675), .CLK(n11011), .Q(
        g6031) );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(n10616), .CLK(n10952), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(n10686), .CLK(n11022), .Q(
        n9367) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(n10626), .CLK(n10962), .Q(
        g4172) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(n10618), .CLK(n10954), .Q(
        g4372) );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(n10618), .CLK(n10954), .Q(
        g3512), .QN(n10427) );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(n10675), .CLK(n11011), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(g25668), .SI(test_si3), .SE(n10618), .CLK(n10954), 
        .Q(g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(n10656), .CLK(n10992), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(n10696), .CLK(n11032), .Q(
        g4235), .QN(n10455) );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(n10651), .CLK(n10987), .Q(
        g1600) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(n10611), .CLK(n10947), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(n10633), .CLK(n10969), .Q(
        g14451), .QN(n10373) );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(n10666), .CLK(n11002), 
        .Q(g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(n10642), .CLK(n10978), .Q(
        g2236), .QN(n10191) );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(n10677), .CLK(n11013), .Q(
        g4555) );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(n10633), .CLK(n10969), .Q(
        g3698), .QN(n10498) );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(n10648), .CLK(n10984), .Q(
        g1736) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(n10636), .CLK(n10972), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(n10674), .CLK(n11010), .Q(
        test_so3), .QN(n10575) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(n10603), .CLK(n10939), 
        .Q(g5607) );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(n10603), .CLK(n10939), .Q(
        g2657) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(n10657), .CLK(n10993), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(n10657), .CLK(n10993), 
        .Q(g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(n10661), .CLK(n10997), .Q(
        g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(n10691), .CLK(n11027), .Q(
        g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(n10602), .CLK(n10938), .Q(
        g5587) );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(n10608), .CLK(n10944), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(n10651), .CLK(n10987), .Q(
        g6377) );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(n10651), .CLK(n10987), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(n10599), .CLK(n10935), .Q(
        g5615) );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(n10698), .CLK(n11034), .Q(
        g4567) );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(n10619), .CLK(n10955), .Q(
        test_so4), .QN(n10573) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(n10664), .CLK(n11000), 
        .Q(g6287) );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(n10612), .CLK(n10948), .Q(
        g7946), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g7946), .SE(n10613), .CLK(n10949), .Q(
        g2563) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(n10684), .CLK(n11020), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(n10684), .CLK(n11020), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(n10684), .CLK(n11020), .Q(
        g6199) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(n10652), .CLK(n10988), .Q(
        g2295) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(n10611), .CLK(n10947), .Q(
        g1384), .QN(n10504) );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(n10637), .CLK(n10973), .Q(
        g1339), .QN(n5381) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(n10637), .CLK(n10973), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(n10649), .CLK(n10985), .Q(
        g2844) );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(n10610), .CLK(n10946), .Q(
        g1024), .QN(n10122) );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(n10603), .CLK(n10939), .Q(
        test_so5) );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(n10670), .CLK(n11006), 
        .Q(g3598) );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(n10670), .CLK(n11006), .Q(
        g4264), .QN(n5823) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(n10672), .CLK(n11008), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(n10672), .CLK(n11008), .Q(
        g5853) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(n10672), .CLK(n11008), .Q(
        g13865) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(n10655), .CLK(n10991), 
        .Q(g2089), .QN(n10065) );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(n10633), .CLK(n10969), .Q(
        g4933), .QN(n5878) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(n10633), .CLK(n10969), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(n10633), .CLK(n10969), .Q(
        g5507) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(n10633), .CLK(n10969), .Q(
        g16656), .QN(n10346) );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(n10653), .CLK(n10989), 
        .Q(g6291) );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(n10621), .CLK(n10957), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(n10703), .CLK(n11039), .Q(
        test_so6) );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(n10693), .CLK(n11029), 
        .Q(g9617) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(n10607), .CLK(n10943), .Q(
        g9741), .QN(n10045) );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(n10607), .CLK(n10943), .Q(
        g3813), .QN(n10087) );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(n10607), .CLK(n10943), .Q(
        g562) );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(n10643), .CLK(n10979), .Q(
        g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(n10655), .CLK(n10991), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(n10615), .CLK(n10951), .Q(
        g3909) );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(n10653), .CLK(n10989), .Q(
        g6259), .QN(n10376) );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(n10678), .CLK(n11014), .Q(
        g5905), .QN(n10332) );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(n10640), .CLK(n10976), .Q(
        g921), .QN(n10132) );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(n10598), .CLK(n10934), .Q(
        g2955), .QN(n10127) );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(n10672), .CLK(n11008), .Q(
        g203), .QN(n10136) );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(n10687), .CLK(n11023), .Q(
        test_so7), .QN(n10583) );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(n10661), .CLK(n10997), 
        .Q(g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(n10629), .CLK(n10965), 
        .Q(g5204), .QN(n10305) );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(n10681), .CLK(n11017), 
        .Q(g17604), .QN(n10335) );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(n10699), .CLK(n11035), 
        .Q(g3606) );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(n10649), .CLK(n10985), 
        .Q(g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(n10676), .CLK(n11012), 
        .Q(g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(n10692), .CLK(n11028), 
        .Q(g3586) );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(n10621), .CLK(n10957), 
        .Q(g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(n10674), .CLK(n11010), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(n10691), .CLK(n11027), 
        .Q(g3570) );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(n10692), .CLK(n11028), 
        .Q(g9048), .QN(n10006) );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(n10692), .CLK(n11028), 
        .Q(g17607), .QN(n10237) );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(n10661), .CLK(n10997), 
        .Q(test_so8), .QN(n10570) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(n10605), .CLK(n10941), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(n10671), .CLK(n11007), .Q(
        g843), .QN(n10109) );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(n10674), .CLK(n11010), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(n10626), .CLK(n10962), 
        .Q(g4153) );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(n10657), .CLK(n10993), 
        .Q(g17711), .QN(n10254) );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(n10607), .CLK(n10943), 
        .Q(g6336), .QN(n5592) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(n10644), .CLK(n10980), 
        .Q(g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(n10667), .CLK(n11003), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(n10677), .CLK(n11013), 
        .Q(g4558) );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(n10689), .CLK(n11025), 
        .Q(g17685), .QN(n10350) );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(n10689), .CLK(n11025), 
        .Q(g3111), .QN(n10084) );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(n10613), .CLK(n10949), 
        .Q(g29217) );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g29217), .SE(n10613), .CLK(n10949), 
        .Q(test_so9) );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(n10701), .CLK(n11037), 
        .Q(g939) );
  SDFFX1 DFF_128_Q_reg ( .D(g25594), .SI(g939), .SE(n10632), .CLK(n10968), .Q(
        g278) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(n10632), .CLK(n10968), .Q(
        g4492) );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(n10633), .CLK(n10969), 
        .Q(g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(n10622), .CLK(n10958), 
        .Q(g1036), .QN(n10090) );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(n10628), .CLK(n10964), 
        .Q(g29220) );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g29220), .SE(n10687), .CLK(n11023), 
        .Q(g1178), .QN(n10137) );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(n10636), .CLK(n10972), 
        .Q(g3239) );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(n10636), .CLK(n10972), 
        .Q(g718), .QN(n10188) );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(n10676), .CLK(n11012), .Q(
        g6195), .QN(n5741) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(n10611), .CLK(n10947), 
        .Q(g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(n10651), .CLK(n10987), 
        .Q(g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(n10634), .CLK(n10970), 
        .Q(test_so10), .QN(n10562) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(n10623), .CLK(n10959), 
        .Q(g554) );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(n10609), .CLK(n10945), .Q(
        g496) );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(n10609), .CLK(n10945), .Q(
        g3853) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(n10628), .CLK(n10964), 
        .Q(g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(n10628), .CLK(n10964), 
        .Q(g17404), .QN(n10129) );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(n10658), .CLK(n10994), 
        .Q(g8344) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(n10647), .CLK(n10983), 
        .Q(g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(n10701), .CLK(n11037), 
        .Q(g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(n10598), .CLK(n10934), .Q(
        n9357) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(n10598), .CLK(n10934), 
        .Q(g5555) );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(n10694), .CLK(n11030), 
        .Q(g14096) );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(n10630), .CLK(n10966), 
        .Q(g1798) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(n10641), .CLK(n10977), 
        .Q(test_so11), .QN(n10554) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(n10702), .CLK(n11038), 
        .Q(g2941), .QN(n10402) );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(n10615), .CLK(n10951), 
        .Q(g3905), .QN(n10339) );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(n10672), .CLK(n11008), 
        .Q(g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(n10653), .CLK(n10989), .Q(
        g6255) );
  SDFFX1 DFF_159_Q_reg ( .D(g26951), .SI(g6255), .SE(n10606), .CLK(n10942), 
        .Q(g4375), .QN(n10012) );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(n10661), .CLK(n10997), 
        .Q(g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(n10683), .CLK(n11019), 
        .Q(g4722) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(n10643), .CLK(n10979), 
        .Q(g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(n10682), .CLK(n11018), .Q(
        g13099), .QN(n10369) );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(n10650), .CLK(n10986), 
        .Q(g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(n10648), .CLK(n10984), 
        .Q(g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(n10648), .CLK(n10984), 
        .Q(g3100), .QN(n10060) );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(n10680), .CLK(n11016), 
        .Q(test_so12) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(n10692), .CLK(n11028), 
        .Q(g1437), .QN(n5696) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(n10608), .CLK(n10944), 
        .Q(g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(n10637), .CLK(n10973), 
        .Q(g1579), .QN(n10118) );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(n10598), .CLK(n10934), 
        .Q(g5567), .QN(n10360) );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(n10648), .CLK(n10984), 
        .Q(g1752) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(n10649), .CLK(n10985), 
        .Q(g1917), .QN(n10469) );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(n10610), .CLK(n10946), 
        .Q(g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(n10683), .CLK(n11019), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(n10683), .CLK(n11019), 
        .Q(g8132) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(n10679), .CLK(n11015), 
        .Q(g6267) );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(n10679), .CLK(n11015), 
        .Q(g16659), .QN(n10241) );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(n10680), .CLK(n11016), 
        .Q(g1442), .QN(n10433) );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(n10665), .CLK(n11001), 
        .Q(test_so13) );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(n10656), .CLK(n10992), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(n10644), .CLK(n10980), 
        .Q(g10500) );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(n10644), .CLK(n10980), 
        .Q(g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(n10626), .CLK(n10962), 
        .Q(g5264) );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(n10650), .CLK(n10986), 
        .Q(g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(n10630), .CLK(n10966), 
        .Q(g2610), .QN(n10468) );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(n10630), .CLK(n10966), 
        .Q(g5160) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(n10677), .CLK(n11013), 
        .Q(g5933) );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(n10693), .CLK(n11029), 
        .Q(g1454), .QN(n5866) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(n10631), .CLK(n10967), 
        .Q(g753), .QN(n10082) );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(n10632), .CLK(n10968), .Q(
        g1296), .QN(n10010) );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(n10632), .CLK(n10968), 
        .Q(g3151) );
  SDFFX1 DFF_197_Q_reg ( .D(g34800), .SI(g3151), .SE(n10686), .CLK(n11022), 
        .Q(test_so14) );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(n10645), .CLK(n10981), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(n10618), .CLK(n10954), 
        .Q(g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(n346), .SI(g3530), .SE(n10641), .CLK(n10977), .Q(
        g4104), .QN(n10274) );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(n10629), .CLK(n10965), 
        .Q(g1532) );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(n10654), .CLK(n10990), 
        .Q(g9251), .QN(n10389) );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(n10642), .CLK(n10978), 
        .Q(n9352) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(n10607), .CLK(n10943), 
        .Q(n9351) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(n10607), .CLK(n10943), 
        .Q(g4754), .QN(n5877) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(n10687), .CLK(n11023), 
        .Q(g1189) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(n10661), .CLK(n10997), 
        .Q(g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(n10670), .CLK(n11006), 
        .Q(g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(n10611), .CLK(n10947), 
        .Q(g1389), .QN(n10460) );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(n10651), .CLK(n10987), 
        .Q(test_so15), .QN(n10587) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(n10657), .CLK(n10993), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(n10687), .CLK(n11023), 
        .Q(g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(n10687), .CLK(n11023), 
        .Q(g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(g33588), .SI(g4269), .SE(n10687), .CLK(n11023), 
        .Q(g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(n10662), .CLK(n10998), 
        .Q(g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(n10598), .CLK(n10934), 
        .Q(g5611) );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(n10658), .CLK(n10994), 
        .Q(g16627), .QN(n10245) );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(n10601), .CLK(n10937), 
        .Q(g4572) );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(n10703), .CLK(n11039), 
        .Q(g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(n10599), .CLK(n10935), 
        .Q(g2898) );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(n10673), .CLK(n11009), 
        .Q(g3343), .QN(n10263) );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(n10673), .CLK(n11009), 
        .Q(g3235) );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(n10691), .CLK(n11027), 
        .Q(test_so16) );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(n10667), .CLK(n11003), 
        .Q(g3566) );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(n10640), .CLK(n10976), 
        .Q(n9348) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(n10601), .CLK(n10937), 
        .Q(g4961) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(n10601), .CLK(n10937), 
        .Q(g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(n10638), .CLK(n10974), 
        .Q(g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(n10604), .CLK(n10940), 
        .Q(g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(n10606), .CLK(n10942), 
        .Q(g7257) );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(n10606), .CLK(n10942), .Q(
        g5802), .QN(n10058) );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(n10649), .CLK(n10985), 
        .Q(g2852) );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(n10649), .CLK(n10985), 
        .Q(g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(n10650), .CLK(n10986), .Q(
        g681), .QN(n10128) );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(n10672), .CLK(n11008), .Q(
        g437) );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(n10654), .CLK(n10990), .Q(
        test_so17), .QN(n10578) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(n10678), .CLK(n11014), 
        .Q(g5901) );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(n10685), .CLK(n11021), 
        .Q(g2886) );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(n10602), .CLK(n10938), 
        .Q(g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(n10602), .CLK(n10938), 
        .Q(g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(n10618), .CLK(n10954), 
        .Q(g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(n10675), .CLK(n11011), 
        .Q(g1604) );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(n10608), .CLK(n10944), 
        .Q(g5092) );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(n10665), .CLK(n11001), 
        .Q(g4831), .QN(n10076) );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(n10665), .CLK(n11001), 
        .Q(g4382), .QN(n5714) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(n10700), .CLK(n11036), 
        .Q(g6386), .QN(n10264) );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(n10702), .CLK(n11038), 
        .Q(g479), .QN(n10116) );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(n10600), .CLK(n10936), .Q(
        g3965) );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(n10620), .CLK(n10956), 
        .Q(test_so18) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(n10675), .CLK(n11011), 
        .Q(g2008) );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(n10675), .CLK(n11011), 
        .Q(g736) );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(n10697), .CLK(n11033), .Q(
        g3933) );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(n10621), .CLK(n10957), 
        .Q(g222) );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(n10648), .CLK(n10984), .Q(
        g3050) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(n10681), .CLK(n11017), 
        .Q(g1052), .QN(n10320) );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(n10681), .CLK(n11017), 
        .Q(g17580), .QN(n10239) );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(n10681), .CLK(n11017), 
        .Q(g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(n10646), .CLK(n10982), 
        .Q(g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(n10667), .CLK(n11003), 
        .Q(g5889) );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(n10667), .CLK(n11003), 
        .Q(g4495) );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(n10671), .CLK(n11007), 
        .Q(g8719), .QN(n10155) );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(n10618), .CLK(n10954), 
        .Q(test_so19), .QN(n10567) );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(n10636), .CLK(n10972), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(n10690), .CLK(n11026), 
        .Q(g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(n10659), .CLK(n10995), 
        .Q(g2433) );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(n10600), .CLK(n10936), 
        .Q(g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(g25748), .SI(g3835), .SE(n10676), .CLK(n11012), 
        .Q(g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(n10676), .CLK(n11012), 
        .Q(g4917) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(n10675), .CLK(n11011), 
        .Q(g1070), .QN(n10529) );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(n10675), .CLK(n11011), 
        .Q(g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(n10675), .CLK(n11011), .Q(
        g17715) );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(n10641), .CLK(n10977), 
        .Q(g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(n10634), .CLK(n10970), .Q(
        g5339) );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(n10626), .CLK(n10962), 
        .Q(g4164), .QN(n10392) );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(n10610), .CLK(n10946), 
        .Q(test_so20) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(n10604), .CLK(n10940), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(n10674), .CLK(n11010), 
        .Q(g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(n10608), .CLK(n10944), 
        .Q(g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(n10608), .CLK(n10944), 
        .Q(g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(n10669), .CLK(n11005), 
        .Q(g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(n10685), .CLK(n11021), 
        .Q(g3680) );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(n10639), .CLK(n10975), 
        .Q(g6637) );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(n10616), .CLK(n10952), 
        .Q(g174) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(n10611), .CLK(n10947), .Q(
        g1682), .QN(n10099) );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(n10654), .CLK(n10990), 
        .Q(g355) );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(n10655), .CLK(n10991), .Q(
        g1087), .QN(n10388) );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(n10688), .CLK(n11024), 
        .Q(g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(n10597), .CLK(n10933), 
        .Q(test_so21), .QN(n10555) );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(n10653), .CLK(n10989), 
        .Q(g6307) );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(n10658), .CLK(n10994), .Q(
        g3802), .QN(n10054) );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(n10676), .CLK(n11012), 
        .Q(g6159), .QN(n10100) );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(n10638), .CLK(n10974), 
        .Q(g2255) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(n10604), .CLK(n10940), 
        .Q(g2815), .QN(n5404) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(n10641), .CLK(n10977), 
        .Q(g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n10533), .SI(g911), .SE(n10658), .CLK(n10994), .Q(
        g43) );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(n10658), .CLK(n10994), .Q(
        g16775), .QN(n10255) );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(n10700), .CLK(n11036), 
        .Q(g1748) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(n10602), .CLK(n10938), 
        .Q(g5551), .QN(n10310) );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(n10619), .CLK(n10955), 
        .Q(g3558) );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(n10702), .CLK(n11038), 
        .Q(g5499), .QN(n5885) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(n10620), .CLK(n10956), 
        .Q(test_so22) );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(n10615), .CLK(n10951), 
        .Q(g3901) );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(n10640), .CLK(n10976), 
        .Q(g4888), .QN(n5863) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(n10689), .CLK(n11025), 
        .Q(g6251), .QN(n10351) );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(n10689), .CLK(n11025), 
        .Q(g17649), .QN(n10246) );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(n10612), .CLK(n10948), 
        .Q(g1373), .QN(n10462) );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(n10636), .CLK(n10972), 
        .Q(g8215) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(n10617), .CLK(n10953), 
        .Q(g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(n10605), .CLK(n10941), .Q(
        g2783), .QN(n5403) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(n10625), .CLK(n10961), .Q(
        g4281), .QN(n10417) );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(n10698), .CLK(n11034), 
        .Q(g3574) );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(n10699), .CLK(n11035), 
        .Q(g2112) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(n10632), .CLK(n10968), 
        .Q(g1283) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(n10632), .CLK(n10968), 
        .Q(test_so23) );
  SDFFX1 DFF_325_Q_reg ( .D(g10122_Tj), .SI(test_si24), .SE(n10670), .CLK(
        n11006), .Q(g4297), .QN(n10492) );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(n10670), .CLK(n11006), 
        .Q(g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(n10672), .CLK(n11008), 
        .Q(g13272), .QN(n10474) );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(n10672), .CLK(n11008), 
        .Q(g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(g34025), .SI(g758), .SE(n10674), .CLK(n11010), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(n10612), .CLK(n10948), 
        .Q(g6537), .QN(n5884) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(n10612), .CLK(n10948), 
        .Q(g5543) );
  SDFFX1 DFF_334_Q_reg ( .D(g7946), .SI(g5543), .SE(n10612), .CLK(n10948), .Q(
        g8475), .QN(n10061) );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(n10665), .CLK(n11001), 
        .Q(g5961) );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(n10679), .CLK(n11015), 
        .Q(g6243), .QN(n10317) );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(n10644), .CLK(n10980), 
        .Q(n9340), .QN(n19032) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(n10644), .CLK(n10980), 
        .Q(g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(n10697), .CLK(n11033), 
        .Q(test_so24) );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(n10619), .CLK(n10955), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(n10619), .CLK(n10955), 
        .Q(g1664) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(n10647), .CLK(n10983), 
        .Q(g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(n10639), .CLK(n10975), 
        .Q(g6629) );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(n10631), .CLK(n10967), 
        .Q(g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(n10658), .CLK(n10994), .Q(
        g4049), .QN(n10490) );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(n10698), .CLK(n11034), 
        .Q(g7260) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(n10698), .CLK(n11034), 
        .Q(g2932) );
  SDFFX1 DFF_350_Q_reg ( .D(g29276), .SI(g2932), .SE(n10654), .CLK(n10990), 
        .Q(g4575) );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(n10654), .CLK(n10990), 
        .Q(g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(n10667), .CLK(n11003), 
        .Q(g4498) );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(n10679), .CLK(n11015), 
        .Q(g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(n10598), .CLK(n10934), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(g25654), .SI(test_si26), .SE(n10609), .CLK(n10945), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(n10609), .CLK(n10945), 
        .Q(g29215) );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g29215), .SE(n10684), .CLK(n11020), 
        .Q(g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(n10621), .CLK(n10957), 
        .Q(g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(n10634), .CLK(n10970), .Q(
        g17639) );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(n10657), .CLK(n10993), 
        .Q(g5831), .QN(n5873) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(n10632), .CLK(n10968), 
        .Q(g239), .QN(n10271) );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(n10668), .CLK(n11004), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(n10685), .CLK(n11021), 
        .Q(g2848) );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(n10634), .CLK(n10970), 
        .Q(g5022), .QN(n10507) );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(n10634), .CLK(n10970), 
        .Q(g16955) );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(n10622), .CLK(n10958), 
        .Q(g1030), .QN(n10461) );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(n10633), .CLK(n10969), 
        .Q(test_so26) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(n10608), .CLK(n10944), 
        .Q(g3231) );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(n10645), .CLK(n10981), 
        .Q(g9817), .QN(n10048) );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(n10645), .CLK(n10981), 
        .Q(g1430), .QN(n10386) );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(n10698), .CLK(n11034), .Q(
        n9336) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(n10638), .CLK(n10974), 
        .Q(g2241), .QN(n10098) );
  SDFFX1 DFF_375_Q_reg ( .D(g24262), .SI(g2241), .SE(n10646), .CLK(n10982), 
        .Q(g1564), .QN(n10385) );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(n10607), .CLK(n10943), 
        .Q(g9680), .QN(n10057) );
  SDFFX1 DFF_377_Q_reg ( .D(test_so92), .SI(g9680), .SE(n10607), .CLK(n10943), 
        .Q(g6148), .QN(n10046) );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(n10639), .CLK(n10975), 
        .Q(g6649) );
  SDFFX1 DFF_379_Q_reg ( .D(g34781), .SI(g6649), .SE(n10630), .CLK(n10966), 
        .Q(g110), .QN(n10531) );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(n10694), .CLK(n11030), .Q(
        g14147) );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(n10694), .CLK(n11030), 
        .Q(g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(n10694), .CLK(n11030), .Q(
        test_so27) );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(n10654), .CLK(n10990), 
        .Q(g4504) );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(n10665), .CLK(n11001), 
        .Q(g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(n10597), .CLK(n10933), 
        .Q(g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(n10597), .CLK(n10933), 
        .Q(g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(g25720), .SI(g2319), .SE(n10701), .CLK(n11037), 
        .Q(g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(n10626), .CLK(n10962), 
        .Q(g11770), .QN(n19035) );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(n10626), .CLK(n10962), 
        .Q(g5208) );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(n10598), .CLK(n10934), 
        .Q(g5579) );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(n10665), .CLK(n11001), 
        .Q(g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(n10689), .CLK(n11025), 
        .Q(g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(n10607), .CLK(n10943), 
        .Q(g5752) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(n10676), .CLK(n11012), 
        .Q(g6279) );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(n10677), .CLK(n11013), 
        .Q(test_so28) );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(n10610), .CLK(n10946), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(n10608), .CLK(n10944), 
        .Q(g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(n10658), .CLK(n10994), 
        .Q(g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(n10646), .CLK(n10982), 
        .Q(g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(n10693), .CLK(n11029), 
        .Q(g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(n10694), .CLK(n11030), 
        .Q(g14125) );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(n10597), .CLK(n10933), 
        .Q(g2370), .QN(n10195) );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(n10667), .CLK(n11003), 
        .Q(g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(n10667), .CLK(n11003), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(n10617), .CLK(n10953), 
        .Q(g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(n10666), .CLK(n11002), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(n10666), .CLK(n11002), 
        .Q(g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(n10684), .CLK(n11020), 
        .Q(test_so29), .QN(n10561) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(n10686), .CLK(n11022), 
        .Q(g2984) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(n10600), .CLK(n10936), 
        .Q(g3961) );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(n10687), .CLK(n11023), 
        .Q(g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(n10607), .CLK(n10943), .Q(
        g101) );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(n10624), .CLK(n10960), .Q(
        g8918), .QN(n19037) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(n10692), .CLK(n11028), 
        .Q(g6625) );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(n10610), .CLK(n10946), 
        .Q(n9332) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(n10610), .CLK(n10946), 
        .Q(g1018), .QN(n10458) );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(n10628), .CLK(n10964), 
        .Q(g17320), .QN(n10130) );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(n10658), .CLK(n10994), 
        .Q(g4045), .QN(n10268) );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(n10658), .CLK(n10994), 
        .Q(g1467), .QN(n5693) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(n10646), .CLK(n10982), 
        .Q(g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(n10663), .CLK(n10999), 
        .Q(test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(n10692), .CLK(n11028), 
        .Q(g5990), .QN(n5589) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(n10637), .CLK(n10973), 
        .Q(g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(n10702), .CLK(n11038), 
        .Q(g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(g29306), .SI(g5029), .SE(n10625), .CLK(n10961), 
        .Q(g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(n10625), .CLK(n10961), 
        .Q(g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(n10690), .CLK(n11026), 
        .Q(g1816), .QN(n10035) );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(n10690), .CLK(n11026), 
        .Q(g4369) );
  SDFFX1 DFF_439_Q_reg ( .D(g29278), .SI(g4369), .SE(n10690), .CLK(n11026), 
        .Q(g4578) );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(n10690), .CLK(n11026), 
        .Q(g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(n10600), .CLK(n10936), 
        .Q(g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(n10659), .CLK(n10995), 
        .Q(g2514), .QN(n10067) );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(n10633), .CLK(n10969), 
        .Q(g3288), .QN(n5400) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(n10598), .CLK(n10934), 
        .Q(test_so31) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(n10643), .CLK(n10979), 
        .Q(g2145), .QN(n5307) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(n10611), .CLK(n10947), 
        .Q(g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(n10679), .CLK(n11015), 
        .Q(g513), .QN(n5548) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(n10613), .CLK(n10949), 
        .Q(g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(n10628), .CLK(n10964), 
        .Q(g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(n10663), .CLK(n10999), 
        .Q(g2763), .QN(n10019) );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(n10684), .CLK(n11020), 
        .Q(g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(n10687), .CLK(n11023), 
        .Q(g952), .QN(n10011) );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(n10637), .CLK(n10973), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(n10691), .CLK(n11027), 
        .Q(g1950), .QN(n10097) );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(n10627), .CLK(n10963), 
        .Q(g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(n10699), .CLK(n11035), 
        .Q(g2307) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(n10699), .CLK(n11035), .Q(
        test_so32) );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(n10617), .CLK(n10953), 
        .Q(g8398), .QN(n10053) );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(n10618), .CLK(n10954), 
        .Q(g4664), .QN(n10055) );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(n10696), .CLK(n11032), 
        .Q(g2223) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(n10656), .CLK(n10992), 
        .Q(g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(n10639), .CLK(n10975), 
        .Q(g6645) );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(n10657), .CLK(n10993), 
        .Q(g2016) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(n10657), .CLK(n10993), 
        .Q(g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(n10657), .CLK(n10993), 
        .Q(g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(n10652), .CLK(n10988), 
        .Q(g2315) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(n10603), .CLK(n10939), 
        .Q(g2811), .QN(n10030) );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(n10678), .CLK(n11014), 
        .Q(g5957) );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(n10655), .CLK(n10991), 
        .Q(g2047) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(n10666), .CLK(n11002), 
        .Q(test_so33), .QN(n10553) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(n10650), .CLK(n10986), 
        .Q(g17760), .QN(n10261) );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(n10602), .CLK(n10938), 
        .Q(g5575) );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(n10617), .CLK(n10953), 
        .Q(n9327) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(n10617), .CLK(n10953), 
        .Q(g3752) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(n10697), .CLK(n11033), 
        .Q(g3917) );
  SDFFX1 DFF_480_Q_reg ( .D(test_so86), .SI(g3917), .SE(n10652), .CLK(n10988), 
        .Q(g8783), .QN(DFF_480_n1) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(n10652), .CLK(n10988), 
        .Q(g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(n10693), .CLK(n11029), 
        .Q(g4388), .QN(n10482) );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(n10653), .CLK(n10989), 
        .Q(g6275) );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(n10653), .CLK(n10989), 
        .Q(g6311) );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(n10653), .CLK(n10989), .Q(
        g8916), .QN(n19034) );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(n10622), .CLK(n10958), 
        .Q(g1041), .QN(n10505) );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(n10630), .CLK(n10966), 
        .Q(test_so34), .QN(n10589) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(n10647), .CLK(n10983), 
        .Q(g2537) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(n10606), .CLK(n10942), 
        .Q(g29221), .QN(g23612) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g29221), .SE(n10606), .CLK(n10942), 
        .Q(g4430), .QN(n10083) );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(n10684), .CLK(n11020), 
        .Q(n9325) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(n10653), .CLK(n10989), 
        .Q(g4826), .QN(n10074) );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(n10679), .CLK(n11015), 
        .Q(g6239) );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(n10695), .CLK(n11031), 
        .Q(g232), .QN(n10270) );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(n10627), .CLK(n10963), .Q(
        g5268) );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(n10627), .CLK(n10963), 
        .Q(g6545) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(n10614), .CLK(n10950), 
        .Q(n9324) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(n10614), .CLK(n10950), 
        .Q(g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(n10597), .CLK(n10933), 
        .Q(g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(n10673), .CLK(n11009), 
        .Q(test_so35), .QN(n10051) );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(n10660), .CLK(n10996), 
        .Q(g1890), .QN(n5799) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(n10646), .CLK(n10982), 
        .Q(g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(n10642), .CLK(n10978), 
        .Q(g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(n10643), .CLK(n10979), .Q(
        g2130) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(n10654), .CLK(n10990), 
        .Q(g4108), .QN(n5715) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(n10654), .CLK(n10990), .Q(
        g4308), .QN(n10418) );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(n10671), .CLK(n11007), 
        .Q(g475) );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(n10681), .CLK(n11017), .Q(
        g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(n10681), .CLK(n11017), .Q(
        g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(n10609), .CLK(n10945), .Q(
        n9322) );
  SDFFX1 DFF_515_Q_reg ( .D(g24213), .SI(n9322), .SE(n10610), .CLK(n10946), 
        .Q(g12184) );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(n10601), .CLK(n10937), 
        .Q(g3990), .QN(n5594) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(n10665), .CLK(n11001), 
        .Q(test_so36), .QN(n10576) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(n10636), .CLK(n10972), 
        .Q(g1992) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(n10636), .CLK(n10972), 
        .Q(g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(n10671), .CLK(n11007), 
        .Q(g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(n10672), .CLK(n11008), .Q(
        g832), .QN(n10419) );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(n10677), .CLK(n11013), .Q(
        g5897), .QN(n10308) );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(n10677), .CLK(n11013), 
        .Q(g25689) );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(n10677), .CLK(n11013), 
        .Q(g4571) );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(n10686), .CLK(n11022), 
        .Q(g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(n10686), .CLK(n11022), 
        .Q(g4455) );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(n10617), .CLK(n10953), 
        .Q(g2902) );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(n10642), .CLK(n10978), 
        .Q(g333) );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(n10616), .CLK(n10952), .Q(
        g168) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(n10603), .CLK(n10939), .Q(
        test_so37), .QN(n10584) );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(n10697), .CLK(n11033), 
        .Q(g3684) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(n10634), .CLK(n10970), 
        .Q(g3639), .QN(n5591) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(n10634), .CLK(n10970), 
        .Q(g14597) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(n10673), .CLK(n11009), 
        .Q(g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(n10673), .CLK(n11009), 
        .Q(g5406) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(n10694), .CLK(n11030), 
        .Q(g269) );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(n10632), .CLK(n10968), .Q(
        g401) );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(n10632), .CLK(n10968), .Q(
        g6040), .QN(n10265) );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(n10672), .CLK(n11008), 
        .Q(g441) );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(n10634), .CLK(n10970), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(n10600), .CLK(n10936), 
        .Q(g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(n10600), .CLK(n10936), 
        .Q(g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(n10655), .CLK(n10991), .Q(
        test_so38), .QN(n10566) );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(n10615), .CLK(n10951), 
        .Q(g3957) );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(n10666), .CLK(n11002), 
        .Q(g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(n10650), .CLK(n10986), 
        .Q(g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(n10650), .CLK(n10986), 
        .Q(g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(n10617), .CLK(n10953), 
        .Q(g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(n10696), .CLK(n11032), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(n10696), .CLK(n11032), 
        .Q(g3498), .QN(n5740) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(n10643), .CLK(n10979), 
        .Q(g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(n10693), .CLK(n11029), .Q(
        g14201) );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(n10663), .CLK(n10999), 
        .Q(g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(n10687), .CLK(n11023), 
        .Q(g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(n10651), .CLK(n10987), 
        .Q(g1608) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(n10652), .CLK(n10988), .Q(
        test_so39), .QN(n10141) );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(n10660), .CLK(n10996), 
        .Q(g17577), .QN(n10327) );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(n10697), .CLK(n11033), 
        .Q(g1779) );
  SDFFX1 DFF_568_Q_reg ( .D(g29255), .SI(g1779), .SE(n10702), .CLK(n11038), 
        .Q(g2652), .QN(n10202) );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(n10603), .CLK(n10939), 
        .Q(g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(n10598), .CLK(n10934), 
        .Q(g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(n10636), .CLK(n10972), 
        .Q(g661) );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(n10601), .CLK(n10937), .Q(
        g4950) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(n10670), .CLK(n11006), 
        .Q(g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(n10604), .CLK(n10940), 
        .Q(g2834), .QN(g23652) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(n10604), .CLK(n10940), 
        .Q(g1361), .QN(n10459) );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(n10676), .CLK(n11012), 
        .Q(g6235) );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(n10687), .CLK(n11023), 
        .Q(g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(n10663), .CLK(n10999), 
        .Q(test_so40) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(n10617), .CLK(n10953), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(n10611), .CLK(n10947), .Q(
        g1696) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(n10667), .CLK(n11003), 
        .Q(g6555), .QN(n10431) );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(n10693), .CLK(n11029), 
        .Q(g14189) );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(n10658), .CLK(n10994), 
        .Q(g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(n10639), .CLK(n10975), 
        .Q(g6621) );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(n10619), .CLK(n10955), 
        .Q(g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(n10614), .CLK(n10950), 
        .Q(g3897), .QN(n10312) );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(n10680), .CLK(n11016), .Q(
        g538) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(n10646), .CLK(n10982), .Q(
        g2606) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(n10659), .CLK(n10995), 
        .Q(g1472), .QN(n5290) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(n10606), .CLK(n10942), 
        .Q(test_so41) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(n10637), .CLK(n10973), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(n10635), .CLK(n10971), 
        .Q(g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(n10681), .CLK(n11017), 
        .Q(g13259), .QN(n10475) );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(n10681), .CLK(n11017), 
        .Q(g405), .QN(n10466) );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(n10627), .CLK(n10963), .Q(
        g5216) );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(n10669), .CLK(n11005), .Q(
        g6494), .QN(n10049) );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(n10618), .CLK(n10954), 
        .Q(g4669), .QN(n10021) );
  SDFFX1 DFF_606_Q_reg ( .D(g24243), .SI(g4669), .SE(n10644), .CLK(n10980), 
        .Q(g996), .QN(n10138) );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(n10645), .CLK(n10981), .Q(
        g4531), .QN(n10486) );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(n10645), .CLK(n10981), 
        .Q(g2860) );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(n10620), .CLK(n10956), 
        .Q(g4743), .QN(n5876) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(n10639), .CLK(n10975), 
        .Q(g6593) );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(n10680), .CLK(n11016), 
        .Q(test_so42), .QN(n10421) );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(n10606), .CLK(n10942), 
        .Q(g4411) );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(n10612), .CLK(n10948), 
        .Q(g1413), .QN(n10528) );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(n10656), .CLK(n10992), 
        .Q(g26960) );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(n10660), .CLK(n10996), 
        .Q(g13039), .QN(n10306) );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(n10660), .CLK(n10996), 
        .Q(g6641) );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(n10660), .CLK(n10996), 
        .Q(g6) );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(n10660), .CLK(n10996), .Q(
        g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n10532), .SI(g1936), .SE(n10660), .CLK(n10996), 
        .Q(g55), .QN(n10008) );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(n10679), .CLK(n11015), .Q(
        g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(n10630), .CLK(n10966), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(n10656), .CLK(n10992), 
        .Q(g4480) );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(n10652), .CLK(n10988), 
        .Q(n9314) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(n10652), .CLK(n10988), 
        .Q(test_so43) );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(n10602), .CLK(n10938), 
        .Q(g5571) );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(n10619), .CLK(n10955), 
        .Q(g3578) );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(n10670), .CLK(n11006), 
        .Q(g9555) );
  SDFFX1 DFF_632_Q_reg ( .D(g29294), .SI(g9555), .SE(n10670), .CLK(n11006), 
        .Q(g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(n10670), .CLK(n11006), 
        .Q(g3582) );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(n10664), .CLK(n11000), 
        .Q(g6271) );
  SDFFX1 DFF_635_Q_reg ( .D(g34028), .SI(g6271), .SE(n10674), .CLK(n11010), 
        .Q(g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(n10697), .CLK(n11033), 
        .Q(g2380), .QN(n10066) );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(n10637), .CLK(n10973), 
        .Q(g5196) );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(n10622), .CLK(n10958), 
        .Q(g3227) );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(n10690), .CLK(n11026), 
        .Q(n9312) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(n10690), .CLK(n11026), 
        .Q(g14518), .QN(n10365) );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(n10690), .CLK(n11026), 
        .Q(test_so44), .QN(n10574) );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(n10625), .CLK(n10961), 
        .Q(g6541), .QN(n5739) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(n10651), .CLK(n10987), 
        .Q(g3203), .QN(n10324) );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(n10651), .CLK(n10987), 
        .Q(g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(n10632), .CLK(n10968), 
        .Q(g4760) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(n10632), .CLK(n10968), 
        .Q(g262), .QN(n10153) );
  SDFFX1 DFF_649_Q_reg ( .D(g33556), .SI(g262), .SE(n10690), .CLK(n11026), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(n10615), .CLK(n10951), 
        .Q(g5467), .QN(n10086) );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(n10615), .CLK(n10951), 
        .Q(g460) );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(n10676), .CLK(n11012), .Q(
        g6209), .QN(n10428) );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(n10642), .CLK(n10978), 
        .Q(g29211), .QN(n10477) );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g29211), .SE(n10648), .CLK(n10984), 
        .Q(g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(n10700), .CLK(n11036), 
        .Q(g655), .QN(n10189) );
  SDFFX1 DFF_657_Q_reg ( .D(g34626), .SI(g655), .SE(n10700), .CLK(n11036), .Q(
        test_so45) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(n10629), .CLK(n10965), 
        .Q(g2204) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(n10629), .CLK(n10965), 
        .Q(g5256) );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(n10684), .CLK(n11020), 
        .Q(g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(n10623), .CLK(n10959), 
        .Q(g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(n10634), .CLK(n10970), .Q(
        g13906) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(n10601), .CLK(n10937), 
        .Q(g4423) );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(n10602), .CLK(n10938), 
        .Q(g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(n10635), .CLK(n10971), 
        .Q(g5685) );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(n10616), .CLK(n10952), 
        .Q(g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(n10671), .CLK(n11007), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(n10609), .CLK(n10945), .Q(
        g3247) );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(n10655), .CLK(n10991), 
        .Q(g2040), .QN(n5505) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(n10655), .CLK(n10991), 
        .Q(test_so46) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(n10626), .CLK(n10962), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(n10673), .CLK(n11009), 
        .Q(g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(n10681), .CLK(n11017), 
        .Q(g7916), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g7916), .SE(n10682), .CLK(n11018), 
        .Q(g4732) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(n10682), .CLK(n11018), 
        .Q(g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(n10656), .CLK(n10992), 
        .Q(g5817), .QN(n10523) );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(n10695), .CLK(n11031), 
        .Q(g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(n10613), .CLK(n10949), 
        .Q(g2648), .QN(n10070) );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(n10683), .CLK(n11019), 
        .Q(g6736), .QN(n10495) );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(n10601), .CLK(n10937), 
        .Q(g4944), .QN(n5875) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(n10654), .CLK(n10990), 
        .Q(g4072) );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(n10654), .CLK(n10990), 
        .Q(g7540) );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(n10697), .CLK(n11033), .Q(
        test_so47) );
  SDFFX1 DFF_688_Q_reg ( .D(g29264), .SI(test_si48), .SE(n10619), .CLK(n10955), 
        .Q(g3466), .QN(n10503) );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(n10701), .CLK(n11037), 
        .Q(g4116) );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(n10597), .CLK(n10933), 
        .Q(g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(n10606), .CLK(n10942), 
        .Q(g4434) );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(n10635), .CLK(n10971), 
        .Q(g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(n10635), .CLK(n10971), 
        .Q(g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(n10635), .CLK(n10971), 
        .Q(g17813) );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(n10609), .CLK(n10945), 
        .Q(g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(n10622), .CLK(n10958), 
        .Q(g3333), .QN(n10077) );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(n10622), .CLK(n10958), 
        .Q(g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(n10674), .CLK(n11010), .Q(
        g4681), .QN(n10435) );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(n10621), .CLK(n10957), 
        .Q(g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(n10700), .CLK(n11036), .Q(
        test_so48), .QN(n10585) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(n10688), .CLK(n11024), 
        .Q(g8789), .QN(n10144) );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(n10649), .CLK(n10985), 
        .Q(g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(n10649), .CLK(n10985), 
        .Q(g2988) );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(n10667), .CLK(n11003), 
        .Q(g3538) );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(n10617), .CLK(n10953), 
        .Q(g301) );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(n10695), .CLK(n11031), .Q(
        n9306), .QN(DFF_709_n1) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(n10695), .CLK(n11031), 
        .Q(g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(n10610), .CLK(n10946), .Q(
        g17291), .QN(n10111) );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(n10646), .CLK(n10982), 
        .Q(g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(n10701), .CLK(n11037), 
        .Q(g5011) );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(n10621), .CLK(n10957), 
        .Q(g199) );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(n10621), .CLK(n10957), .Q(
        g6523), .QN(n5870) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(n10629), .CLK(n10965), 
        .Q(test_so49), .QN(n10568) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(n10684), .CLK(n11020), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(n10616), .CLK(n10952), 
        .Q(g854) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(n10629), .CLK(n10965), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(n10676), .CLK(n11012), 
        .Q(g4922) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(n10665), .CLK(n11001), 
        .Q(g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(n10665), .CLK(n11001), 
        .Q(g5863), .QN(n10430) );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(n10645), .CLK(n10981), 
        .Q(g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(g29253), .SI(g4581), .SE(n10647), .CLK(n10983), 
        .Q(g2518), .QN(n10200) );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(n10613), .CLK(n10949), 
        .Q(g2567) );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(n10642), .CLK(n10978), 
        .Q(g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(n10622), .CLK(n10958), .Q(
        g3263) );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(n10638), .CLK(n10974), 
        .Q(g6613) );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(n10692), .CLK(n11028), 
        .Q(test_so50), .QN(n10579) );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(n10700), .CLK(n11036), 
        .Q(g6444) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(n10610), .CLK(n10946), 
        .Q(g2965) );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(n10667), .CLK(n11003), 
        .Q(g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(n10699), .CLK(n11035), 
        .Q(n9303) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(n10631), .CLK(n10967), 
        .Q(g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(n10692), .CLK(n11028), .Q(
        g17646), .QN(n10331) );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(n10618), .CLK(n10954), 
        .Q(g3562), .QN(n10372) );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(n10670), .CLK(n11006), 
        .Q(g10122_Tj), .QN(n10491) );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122_Tj), .SE(n10689), .CLK(n11025), 
        .Q(g1404), .QN(n10500) );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(n10600), .CLK(n10936), 
        .Q(g3817), .QN(n10502) );
  SDFFX1 DFF_743_Q_reg ( .D(n10537), .SI(g3817), .SE(n10620), .CLK(n10956), 
        .Q(n9302) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(n10620), .CLK(n10956), 
        .Q(g4501) );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(n10621), .CLK(n10957), 
        .Q(test_so51), .QN(n10571) );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(n10662), .CLK(n10998), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(n10628), .CLK(n10964), 
        .Q(g4704) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(n10599), .CLK(n10935), .Q(
        g2878) );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(n10627), .CLK(n10963), 
        .Q(g5220), .QN(n10276) );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(n10644), .CLK(n10980), 
        .Q(g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(n10644), .CLK(n10980), .Q(
        g12368) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(n10693), .CLK(n11029), 
        .Q(g316) );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(n10701), .CLK(n11037), .Q(
        g1277) );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(n10625), .CLK(n10961), 
        .Q(g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(n10693), .CLK(n11029), 
        .Q(g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(n10599), .CLK(n10935), .Q(
        g2882) );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(n10701), .CLK(n11037), 
        .Q(test_so52) );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(n10661), .CLK(n10997), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(n10661), .CLK(n10997), 
        .Q(g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(g34975), .SI(g305), .SE(n10702), .CLK(n11038), .Q(
        g8) );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(n10603), .CLK(n10939), .Q(
        g2799), .QN(n10027) );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(n10694), .CLK(n11030), 
        .Q(g14167) );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(n10694), .CLK(n11030), 
        .Q(g17787) );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(n10694), .CLK(n11030), 
        .Q(g4912) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(n10626), .CLK(n10962), 
        .Q(g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(n10647), .CLK(n10983), 
        .Q(g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(n10688), .CLK(n11024), 
        .Q(g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(n10606), .CLK(n10942), 
        .Q(g550), .QN(n10413) );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(n10695), .CLK(n11031), .Q(
        g255), .QN(n10152) );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(n10700), .CLK(n11036), .Q(
        test_so53), .QN(n10572) );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(n10638), .CLK(n10974), 
        .Q(g5240) );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(n10638), .CLK(n10974), 
        .Q(g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(n10666), .CLK(n11002), 
        .Q(g3863), .QN(n10432) );
  SDFFX1 DFF_777_Q_reg ( .D(g29245), .SI(g3863), .SE(n10700), .CLK(n11036), 
        .Q(g1959), .QN(n10199) );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(n10602), .CLK(n10938), 
        .Q(g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(n10639), .CLK(n10975), 
        .Q(g6653) );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(n10683), .CLK(n11019), 
        .Q(g17764) );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(n10640), .CLK(n10976), 
        .Q(g2864) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(n10640), .CLK(n10976), 
        .Q(g4894) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(n10635), .CLK(n10971), 
        .Q(g17678) );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(n10666), .CLK(n11002), 
        .Q(g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(n10679), .CLK(n11015), 
        .Q(g16693), .QN(n10338) );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(n10679), .CLK(n11015), 
        .Q(test_so54), .QN(n10581) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(n10622), .CLK(n10958), 
        .Q(g1002), .QN(n10510) );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(n10623), .CLK(n10959), 
        .Q(g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(n10623), .CLK(n10959), .Q(
        g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(n10644), .CLK(n10980), .Q(
        g1236), .QN(n10117) );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(n10674), .CLK(n11010), 
        .Q(g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(n10646), .CLK(n10982), 
        .Q(g2476), .QN(n10470) );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(n10619), .CLK(n10955), 
        .Q(g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(n10661), .CLK(n10997), 
        .Q(g2375), .QN(n10096) );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(n10661), .CLK(n10997), 
        .Q(g63), .QN(n10131) );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(n10671), .CLK(n11007), .Q(
        g17739), .QN(n10252) );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(n10671), .CLK(n11007), 
        .Q(g358), .QN(n10526) );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(n10671), .CLK(n11007), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(g28043), .SI(g896), .SE(n10702), .CLK(n11038), .Q(
        test_so55), .QN(n10558) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(n10666), .CLK(n11002), 
        .Q(g3161), .QN(n10425) );
  SDFFX1 DFF_804_Q_reg ( .D(g29251), .SI(g3161), .SE(n10597), .CLK(n10933), 
        .Q(g2384), .QN(n10194) );
  SDFFX1 DFF_806_Q_reg ( .D(test_so80), .SI(g2384), .SE(n10683), .CLK(n11019), 
        .Q(g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(n10684), .CLK(n11020), 
        .Q(g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(n10684), .CLK(n11020), 
        .Q(g4561) );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(n10690), .CLK(n11026), 
        .Q(g2024) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(n10623), .CLK(n10959), .Q(
        g3451), .QN(n10037) );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(n10605), .CLK(n10941), 
        .Q(g2795), .QN(n10028) );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(n10643), .CLK(n10979), 
        .Q(g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(n10702), .CLK(n11038), .Q(
        g4527) );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(n10631), .CLK(n10967), 
        .Q(g1844) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(n10678), .CLK(n11014), 
        .Q(g5937) );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(n10698), .CLK(n11034), 
        .Q(test_so56) );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(n10647), .CLK(n10983), 
        .Q(g2523) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(n10686), .CLK(n11022), 
        .Q(g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(n10613), .CLK(n10949), 
        .Q(g2643), .QN(n10095) );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(n10680), .CLK(n11016), 
        .Q(g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(n10680), .CLK(n11016), 
        .Q(g8358), .QN(n10139) );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(n10647), .CLK(n10983), 
        .Q(n9295) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(n10647), .CLK(n10983), 
        .Q(g5156), .QN(n5734) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(n10647), .CLK(n10983), 
        .Q(g30332), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(g34975), .SI(g30332), .SE(n10623), .CLK(n10959), 
        .Q(n9294) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(n10623), .CLK(n10959), 
        .Q(g8279) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(n10625), .CLK(n10961), 
        .Q(g8839) );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(n10691), .CLK(n11027), 
        .Q(g1955), .QN(n10063) );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(n10692), .CLK(n11028), 
        .Q(test_so57), .QN(n10559) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(n10638), .CLK(n10974), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(n10683), .CLK(n11019), 
        .Q(g14749) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(n10700), .CLK(n11036), 
        .Q(g4771) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(n10607), .CLK(n10943), 
        .Q(g6098) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(n10651), .CLK(n10987), 
        .Q(g3147), .QN(n5738) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(n10691), .CLK(n11027), 
        .Q(g3347), .QN(n10487) );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(n10638), .CLK(n10974), 
        .Q(g2269) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(n10680), .CLK(n11016), .Q(
        g191), .QN(n10140) );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(n10680), .CLK(n11016), .Q(
        g2712), .QN(n10493) );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(n10644), .CLK(n10980), 
        .Q(g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(n10628), .CLK(n10964), 
        .Q(g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(n10662), .CLK(n10998), 
        .Q(test_so58), .QN(n10560) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(n10656), .CLK(n10992), 
        .Q(g17819) );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(n10685), .CLK(n11021), 
        .Q(g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(n10698), .CLK(n11034), 
        .Q(g2927), .QN(n10123) );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(n10644), .CLK(n10980), 
        .Q(g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(n10678), .CLK(n11014), 
        .Q(g5929) );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(n10678), .CLK(n11014), 
        .Q(g4907) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(n10685), .CLK(n11021), 
        .Q(g16874) );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(n10685), .CLK(n11021), 
        .Q(g4035), .QN(n10078) );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(n10685), .CLK(n11021), 
        .Q(g2946) );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(n10641), .CLK(n10977), 
        .Q(g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(n10641), .CLK(n10977), .Q(
        g4082), .QN(n10467) );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(n10669), .CLK(n11005), 
        .Q(g9743) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(n10605), .CLK(n10941), 
        .Q(test_so59), .QN(n10590) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(n10643), .CLK(n10979), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(n10699), .CLK(n11035), .Q(
        g1620) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(n10605), .CLK(n10941), 
        .Q(g2831), .QN(g30331) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(n10605), .CLK(n10941), 
        .Q(g667) );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(n10701), .CLK(n11037), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(n10614), .CLK(n10950), .Q(
        g3937) );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(n10672), .CLK(n11008), 
        .Q(g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(n10689), .CLK(n11025), .Q(
        g1249), .QN(n10512) );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(n10616), .CLK(n10952), 
        .Q(g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(n10633), .CLK(n10969), .Q(
        g16924) );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(n10643), .CLK(n10979), 
        .Q(g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(n10599), .CLK(n10935), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(n10675), .CLK(n11011), 
        .Q(test_so60) );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(n10677), .CLK(n11013), 
        .Q(g5949) );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(n10640), .CLK(n10976), 
        .Q(g6682), .QN(n5590) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(n10640), .CLK(n10976), 
        .Q(g904), .QN(n10513) );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(n10649), .CLK(n10985), .Q(
        g2873), .QN(n5488) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(n10700), .CLK(n11036), 
        .Q(g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(n10608), .CLK(n10944), 
        .Q(g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(n10602), .CLK(n10938), 
        .Q(g5603) );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(n10624), .CLK(n10960), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(n10693), .CLK(n11029), 
        .Q(g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(n10659), .CLK(n10995), 
        .Q(g2437) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(n10656), .CLK(n10992), 
        .Q(g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(n10696), .CLK(n11032), 
        .Q(g2208), .QN(n10471) );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(n10613), .CLK(n10949), 
        .Q(test_so61) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(n10625), .CLK(n10961), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(n10662), .CLK(n10998), 
        .Q(g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(n10662), .CLK(n10998), 
        .Q(g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(n10685), .CLK(n11021), 
        .Q(g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(n10598), .CLK(n10934), 
        .Q(g5583) );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(n10623), .CLK(n10959), 
        .Q(g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(n10651), .CLK(n10987), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(n10651), .CLK(n10987), 
        .Q(g17743) );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(n10617), .CLK(n10953), 
        .Q(g2917), .QN(n10124) );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(n10636), .CLK(n10972), 
        .Q(g686) );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(n10636), .CLK(n10972), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(n10605), .CLK(n10941), 
        .Q(g671), .QN(n10042) );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(n10688), .CLK(n11024), .Q(
        test_so62), .QN(n10586) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(n10680), .CLK(n11016), 
        .Q(g6283) );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(n10660), .CLK(n10996), 
        .Q(g14705) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(n10660), .CLK(n10996), 
        .Q(g17519), .QN(n10235) );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(n10660), .CLK(n10996), 
        .Q(g8784), .QN(DFF_909_n1) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(n10669), .CLK(n11005), 
        .Q(g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(n10694), .CLK(n11030), 
        .Q(g4489) );
  SDFFX1 DFF_912_Q_reg ( .D(g33564), .SI(g4489), .SE(n10694), .CLK(n11030), 
        .Q(g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(n10637), .CLK(n10973), 
        .Q(g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(n10662), .CLK(n10998), 
        .Q(g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(n10653), .CLK(n10989), 
        .Q(g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(n10615), .CLK(n10951), 
        .Q(g3929) );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(n10615), .CLK(n10951), 
        .Q(g5503), .QN(n5737) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(n10624), .CLK(n10960), 
        .Q(test_so63) );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(n10678), .CLK(n11014), 
        .Q(g5925) );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(n10688), .CLK(n11024), 
        .Q(g1124), .QN(n5692) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(n10601), .CLK(n10937), 
        .Q(g4955), .QN(n5614) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(n10638), .CLK(n10974), 
        .Q(g5224) );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(n10676), .CLK(n11012), 
        .Q(g2012) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(n10676), .CLK(n11012), 
        .Q(g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(n10648), .CLK(n10984), 
        .Q(g5120), .QN(n10085) );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(n10648), .CLK(n10984), 
        .Q(g17674), .QN(n10250) );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(n10597), .CLK(n10933), 
        .Q(g2389) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(n10602), .CLK(n10938), 
        .Q(g4438) );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(n10659), .CLK(n10995), 
        .Q(g2429) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(n10605), .CLK(n10941), 
        .Q(g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(n10702), .CLK(n11038), 
        .Q(test_so64) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(n10603), .CLK(n10939), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(n10673), .CLK(n11009), 
        .Q(g18881) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g18881), .SE(n10674), .CLK(n11010), 
        .Q(g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(n10675), .CLK(n11011), 
        .Q(g1199) );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(n10604), .CLK(n10940), 
        .Q(g19357), .QN(n5401) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(n10602), .CLK(n10938), 
        .Q(g5547) );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(n10643), .CLK(n10979), 
        .Q(g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(n10657), .CLK(n10993), 
        .Q(g16744), .QN(n10259) );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(n10664), .CLK(n11000), 
        .Q(g2338) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(n10664), .CLK(n11000), .Q(
        g8919), .QN(n19038) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(n10664), .CLK(n11000), 
        .Q(g6247) );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(n10614), .CLK(n10950), 
        .Q(g2791), .QN(n10029) );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(n10614), .CLK(n10950), 
        .Q(test_so65) );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(n10597), .CLK(n10933), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(n10678), .CLK(n11014), 
        .Q(g5945) );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(n10629), .CLK(n10965), 
        .Q(g5244) );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(n10663), .CLK(n10999), 
        .Q(g2759), .QN(n10530) );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(n10640), .CLK(n10976), 
        .Q(g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(n10623), .CLK(n10959), 
        .Q(g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(n10637), .CLK(n10973), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(n10602), .CLK(n10938), 
        .Q(g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(n10680), .CLK(n11016), 
        .Q(g209), .QN(n5595) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(n10669), .CLK(n11005), .Q(
        g6609) );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(n10669), .CLK(n11005), 
        .Q(g5517), .QN(n10426) );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(n10659), .CLK(n10995), 
        .Q(g2449) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(n10630), .CLK(n10966), 
        .Q(test_so66) );
  SDFFX1 DFF_961_Q_reg ( .D(g18881), .SI(test_si67), .SE(n10674), .CLK(n11010), 
        .Q(n9281), .QN(DFF_961_n1) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(n10613), .CLK(n10949), 
        .Q(g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(n10641), .CLK(n10977), 
        .Q(g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(n10655), .CLK(n10991), .Q(
        g2098) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(n10655), .CLK(n10991), 
        .Q(g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(n10643), .CLK(n10979), 
        .Q(g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(n10697), .CLK(n11033), .Q(
        g6589), .QN(n10313) );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(n10660), .CLK(n10996), 
        .Q(n9280) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(n10660), .CLK(n10996), 
        .Q(g17845) );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(n10683), .CLK(n11019), 
        .Q(g17871) );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(n10632), .CLK(n10968), 
        .Q(g429) );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(n10659), .CLK(n10995), .Q(
        g1870) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(n10624), .CLK(n10960), 
        .Q(test_so67) );
  SDFFX1 DFF_977_Q_reg ( .D(g29243), .SI(test_si68), .SE(n10631), .CLK(n10967), 
        .Q(g1825), .QN(n10192) );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(n10622), .CLK(n10958), 
        .Q(g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(n10668), .CLK(n11004), 
        .Q(g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(test_so46), .SI(g4392), .SE(n10668), .CLK(n11004), 
        .Q(g8283), .QN(n10112) );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(n10691), .CLK(n11027), 
        .Q(g3546), .QN(n10315) );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(n10627), .CLK(n10963), 
        .Q(g5236) );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(n10614), .CLK(n10950), 
        .Q(g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(n10662), .CLK(n10998), 
        .Q(g4854), .QN(n10041) );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(n10615), .CLK(n10951), 
        .Q(g3925) );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(n10625), .CLK(n10961), 
        .Q(g6509), .QN(n10484) );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(n10631), .CLK(n10967), 
        .Q(g732), .QN(n5732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(n10647), .CLK(n10983), .Q(
        g2504), .QN(n10302) );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(n10672), .CLK(n11008), 
        .Q(test_so68), .QN(n10550) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(n10624), .CLK(n10960), 
        .Q(g4520) );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(n10624), .CLK(n10960), .Q(
        g8917), .QN(n19036) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(n10696), .CLK(n11032), 
        .Q(g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(n10645), .CLK(n10981), 
        .Q(g37), .QN(g30327) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(n10635), .CLK(n10971), .Q(
        g4031) );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(n10657), .CLK(n10993), 
        .Q(g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(n10683), .CLK(n11019), .Q(
        g8235), .QN(n10114) );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(n10626), .CLK(n10962), 
        .Q(g4176) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(n10658), .CLK(n10994), 
        .Q(g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(n10668), .CLK(n11004), 
        .Q(g4405) );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(n10694), .CLK(n11030), 
        .Q(g872) );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(n10608), .CLK(n10944), 
        .Q(g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(n10700), .CLK(n11036), 
        .Q(test_so69), .QN(n10563) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(n10607), .CLK(n10943), .Q(g4765), .QN(n5613) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(n10598), .CLK(n10934), 
        .Q(g5563) );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(n10689), .CLK(n11025), 
        .Q(g1395), .QN(n10319) );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(n10661), .CLK(n10997), 
        .Q(g1913) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(n10661), .CLK(n10997), 
        .Q(g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(n10676), .CLK(n11012), 
        .Q(g6263) );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(n10599), .CLK(n10935), 
        .Q(n9276) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(n10600), .CLK(n10936), 
        .Q(g3945) );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(n10654), .CLK(n10990), 
        .Q(g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(n10645), .CLK(n10981), 
        .Q(g4473), .QN(n10494) );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(n10689), .CLK(n11025), 
        .Q(g1266), .QN(n10133) );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(n10701), .CLK(n11037), 
        .Q(g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(n10605), .CLK(n10941), 
        .Q(test_so70), .QN(n10580) );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(n10663), .CLK(n10999), .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(n10599), .CLK(n10935), 
        .Q(g5471), .QN(n10521) );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(n10645), .CLK(n10981), 
        .Q(g4540) );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(n10645), .CLK(n10981), 
        .Q(g6723) );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(n10639), .CLK(n10975), 
        .Q(g6605), .QN(n10368) );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(n10659), .CLK(n10995), 
        .Q(n9274) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(n10642), .CLK(n10978), 
        .Q(g2173) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(n10642), .CLK(n10978), 
        .Q(g9019) );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(n10647), .CLK(n10983), 
        .Q(g2491) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(n10662), .CLK(n10998), 
        .Q(g4849), .QN(n10506) );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(n10641), .CLK(n10977), 
        .Q(g2169) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(n10638), .CLK(n10974), 
        .Q(n9273) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(n10638), .CLK(n10974), 
        .Q(test_so71) );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(n10614), .CLK(n10950), .Q(g29219) );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g29219), .SE(n10614), .CLK(n10950), 
        .Q(g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(n10649), .CLK(n10985), 
        .Q(g2868), .QN(n10476) );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(n10650), .CLK(n10986), 
        .Q(g2767), .QN(n10032) );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(n10650), .CLK(n10986), 
        .Q(g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(n10686), .CLK(n11022), 
        .Q(g16718), .QN(n10248) );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(n10604), .CLK(n10940), 
        .Q(g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(n10702), .CLK(n11038), 
        .Q(g5212), .QN(n10328) );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(n10625), .CLK(n10961), 
        .Q(g4245) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(n10631), .CLK(n10967), 
        .Q(g645) );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(n10642), .CLK(n10978), .Q(
        g4291), .QN(n10416) );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(n10616), .CLK(n10952), 
        .Q(g29212), .QN(n5657) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g29212), .SE(n10616), .CLK(n10952), 
        .Q(test_so72) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(n10688), .CLK(n11024), .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(n10688), .CLK(n11024), 
        .Q(g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(n10688), .CLK(n11024), 
        .Q(g8788), .QN(n10143) );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(n10638), .CLK(n10974), 
        .Q(g2246), .QN(n10069) );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(n10631), .CLK(n10967), 
        .Q(g1830) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(n10699), .CLK(n11035), 
        .Q(g3590) );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(n10616), .CLK(n10952), 
        .Q(g392), .QN(n10465) );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(n10651), .CLK(n10987), 
        .Q(g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(n10625), .CLK(n10961), 
        .Q(g6505), .QN(n10101) );
  SDFFX1 DFF_1057_Q_reg ( .D(g24246), .SI(g6505), .SE(n10655), .CLK(n10991), 
        .Q(g1221), .QN(n10387) );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(n10677), .CLK(n11013), 
        .Q(g5921) );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(n10693), .CLK(n11029), 
        .Q(g29216) );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g29216), .SE(n10695), .CLK(n11031), 
        .Q(test_so73) );
  SDFFX1 DFF_1061_Q_reg ( .D(test_so42), .SI(test_si74), .SE(n10680), .CLK(
        n11016), .Q(g218), .QN(n10422) );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(n10649), .CLK(n10985), 
        .Q(g1932) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(n10696), .CLK(n11032), 
        .Q(g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(n10702), .CLK(n11038), 
        .Q(g5062), .QN(n10508) );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(n10599), .CLK(n10935), 
        .Q(g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(n10599), .CLK(n10935), 
        .Q(g2689) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(n10669), .CLK(n11005), 
        .Q(g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(n10619), .CLK(n10955), 
        .Q(g1677), .QN(n10197) );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(n10663), .CLK(n10999), 
        .Q(g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(n10603), .CLK(n10939), 
        .Q(g2671) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(n10637), .CLK(n10973), 
        .Q(g10527) );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(n10668), .CLK(n11004), 
        .Q(g7243) );
  SDFFX1 DFF_1074_Q_reg ( .D(n10532), .SI(g7243), .SE(n10668), .CLK(n11004), 
        .Q(test_so74) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(n10631), .CLK(n10967), .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(n10703), .CLK(n11039), 
        .Q(g29213), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g29213), .SE(n10599), .CLK(n10935), 
        .Q(g5485), .QN(n5869) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(n10663), .CLK(n10999), 
        .Q(g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(n10610), .CLK(n10946), 
        .Q(g11678), .QN(n5482) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(n10613), .CLK(n10949), 
        .Q(g2638), .QN(n10201) );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(n10626), .CLK(n10962), 
        .Q(g4122) );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(n10674), .CLK(n11010), 
        .Q(g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(n10678), .CLK(n11014), 
        .Q(g5941) );
  SDFFX1 DFF_1086_Q_reg ( .D(g33572), .SI(g5941), .SE(n10656), .CLK(n10992), 
        .Q(g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(n10656), .CLK(n10992), 
        .Q(g13068), .QN(n10357) );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(n10656), .CLK(n10992), .Q(
        g25), .QN(n10473) );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(n10610), .CLK(n10946), .Q(
        test_so75) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(n10643), .CLK(n10979), .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(n10696), .CLK(n11032), 
        .Q(g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(n10604), .CLK(n10940), 
        .Q(n9267) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(n10604), .CLK(n10940), 
        .Q(g2066) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(n10687), .CLK(n11023), 
        .Q(g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(n10627), .CLK(n10963), 
        .Q(g5252) );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(n10688), .CLK(n11024), 
        .Q(g2165) );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(n10613), .CLK(n10949), 
        .Q(g2571) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(n10667), .CLK(n11003), 
        .Q(g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(n10668), .CLK(n11004), 
        .Q(g8403), .QN(n10113) );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(n10668), .CLK(n11004), 
        .Q(g14673) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(n10668), .CLK(n11004), 
        .Q(test_so76), .QN(n10565) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(n10604), .CLK(n10940), .Q(g2827), .QN(n10031) );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(n10693), .CLK(n11029), 
        .Q(g14217) );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(n10662), .CLK(n10998), 
        .Q(g4859), .QN(n10018) );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(n10671), .CLK(n11007), 
        .Q(g424) );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(n10637), .CLK(n10973), 
        .Q(g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(n10637), .CLK(n10973), 
        .Q(g17423), .QN(n10516) );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(n10696), .CLK(n11032), 
        .Q(n9265), .QN(n6006) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(n10604), .CLK(n10940), 
        .Q(g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(n10691), .CLK(n11027), 
        .Q(g1821), .QN(n10064) );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(n10659), .CLK(n10995), 
        .Q(g2509), .QN(n10094) );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(n10664), .CLK(n11000), 
        .Q(g5073), .QN(n10481) );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(n10689), .CLK(n11025), 
        .Q(test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(n10683), .CLK(n11019), 
        .Q(g8353), .QN(n10115) );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(n10689), .CLK(n11025), 
        .Q(g13085), .QN(n10377) );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(n10639), .CLK(n10975), 
        .Q(g6633) );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(n10627), .CLK(n10963), 
        .Q(g5124), .QN(n10525) );
  SDFFX1 DFF_1122_Q_reg ( .D(test_so44), .SI(g5124), .SE(n10691), .CLK(n11027), 
        .Q(g17400), .QN(n10515) );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(n10664), .CLK(n11000), 
        .Q(g6303) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(n10664), .CLK(n11000), 
        .Q(g5069), .QN(n10091) );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(n10698), .CLK(n11034), 
        .Q(g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(n10650), .CLK(n10986), 
        .Q(g650) );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(n10650), .CLK(n10986), 
        .Q(g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(n10614), .CLK(n10950), 
        .Q(g3921) );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(n10697), .CLK(n11033), 
        .Q(test_so78) );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(n10683), .CLK(n11019), .Q(g6732), .QN(n10380) );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(n10629), .CLK(n10965), 
        .Q(g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(n10686), .CLK(n11022), 
        .Q(g1061), .QN(n10499) );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(n10696), .CLK(n11032), 
        .Q(g3462), .QN(n10088) );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(n10642), .CLK(n10978), 
        .Q(g2181) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(n10689), .CLK(n11025), 
        .Q(g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(n10648), .CLK(n10984), 
        .Q(g1756) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(n10665), .CLK(n11001), 
        .Q(g5849), .QN(n5736) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(n10701), .CLK(n11037), 
        .Q(g4112) );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(n10603), .CLK(n10939), 
        .Q(n9262) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(n10603), .CLK(n10939), 
        .Q(g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(n10693), .CLK(n11029), 
        .Q(test_so79), .QN(n10569) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(n10622), .CLK(n10958), .Q(g1046), .QN(n10452) );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(n10679), .CLK(n11015), 
        .Q(g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(n10669), .CLK(n11005), 
        .Q(g4401), .QN(n10080) );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(n10669), .CLK(n11005), 
        .Q(g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(n10669), .CLK(n11005), 
        .Q(g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(n10669), .CLK(n11005), 
        .Q(g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(n10620), .CLK(n10956), 
        .Q(g2950), .QN(n10400) );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(n10612), .CLK(n10948), 
        .Q(g1345), .QN(n10511) );
  SDFFX1 DFF_1154_Q_reg ( .D(g25762), .SI(g1345), .SE(n10612), .CLK(n10948), 
        .Q(g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(n10682), .CLK(n11018), 
        .Q(g14421), .QN(n10353) );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(n10682), .CLK(n11018), 
        .Q(g4727) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(n10683), .CLK(n11019), 
        .Q(test_so80), .QN(n10557) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(n10612), .CLK(n10948), .Q(g1536) );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(n10615), .CLK(n10951), 
        .Q(g3941) );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(n10671), .CLK(n11007), 
        .Q(g370), .QN(n10156) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(n10620), .CLK(n10956), 
        .Q(g5694), .QN(n10267) );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(n10631), .CLK(n10967), 
        .Q(g1858) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(n10631), .CLK(n10967), 
        .Q(g446) );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(n10666), .CLK(n11002), 
        .Q(g3219) );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(n10630), .CLK(n10966), 
        .Q(g1811), .QN(n10193) );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(n10639), .CLK(n10975), 
        .Q(g6601) );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(n10659), .CLK(n10995), 
        .Q(g2441) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(n10659), .CLK(n10995), 
        .Q(g1874) );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(n10644), .CLK(n10980), 
        .Q(test_so81), .QN(n10552) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(n10669), .CLK(n11005), .Q(g6581) );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(n10639), .CLK(n10975), 
        .Q(g6597), .QN(n10343) );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(n10668), .CLK(n11004), 
        .Q(g5008) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(n10619), .CLK(n10955), 
        .Q(g3610) );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(n10649), .CLK(n10985), 
        .Q(g2890) );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(n10636), .CLK(n10972), 
        .Q(g1978) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(n10699), .CLK(n11035), 
        .Q(g1612) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(n10646), .CLK(n10982), 
        .Q(g112), .QN(n10463) );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(n10685), .CLK(n11021), 
        .Q(g2856) );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(n10636), .CLK(n10972), 
        .Q(g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(n10682), .CLK(n11018), 
        .Q(g17722), .QN(n10342) );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(n10629), .CLK(n10965), 
        .Q(test_so82) );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(n10625), .CLK(n10961), .Q(g4119) );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(n10650), .CLK(n10986), 
        .Q(g6390), .QN(n10488) );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(n10612), .CLK(n10948), 
        .Q(g1542) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(n10612), .CLK(n10948), 
        .Q(g4258), .QN(n10501) );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(n10684), .CLK(n11020), 
        .Q(g4818) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(n10597), .CLK(n10933), 
        .Q(g5033), .QN(n10464) );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(n10682), .CLK(n11018), 
        .Q(g4717) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(n10682), .CLK(n11018), 
        .Q(g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(n10682), .CLK(n11018), 
        .Q(g3849), .QN(n5735) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(n10682), .CLK(n11018), 
        .Q(g17778), .QN(n10257) );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(n10699), .CLK(n11035), 
        .Q(g3199) );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(n10699), .CLK(n11035), 
        .Q(test_so83), .QN(n10593) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(n10662), .CLK(n10998), .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(n10623), .CLK(n10959), 
        .Q(g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(n10678), .CLK(n11014), 
        .Q(g5913), .QN(n10356) );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(n10649), .CLK(n10985), 
        .Q(g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(n10608), .CLK(n10944), 
        .Q(g6163), .QN(n10522) );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(n10677), .CLK(n11013), 
        .Q(g4125), .QN(n10497) );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(n10677), .CLK(n11013), 
        .Q(g4821), .QN(n5880) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(n10633), .CLK(n10969), 
        .Q(g4939) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(n10681), .CLK(n11017), 
        .Q(g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(n10621), .CLK(n10957), 
        .Q(g3207) );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(n10624), .CLK(n10960), 
        .Q(g4483) );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(n10622), .CLK(n10958), 
        .Q(test_so84) );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(n10627), .CLK(n10963), .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(n10626), .CLK(n10962), 
        .Q(g5248) );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(n10600), .CLK(n10936), 
        .Q(g2126) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(n10601), .CLK(n10937), 
        .Q(g3694), .QN(n10266) );
  SDFFX1 DFF_1215_Q_reg ( .D(g29288), .SI(g3694), .SE(n10635), .CLK(n10971), 
        .Q(g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(n10635), .CLK(n10971), 
        .Q(g1964) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(n10608), .CLK(n10944), 
        .Q(g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(n10608), .CLK(n10944), 
        .Q(g3215) );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(n10635), .CLK(n10971), 
        .Q(g16748) );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(n10696), .CLK(n11032), 
        .Q(n9255), .QN(n6005) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(n10606), .CLK(n10942), 
        .Q(g4427), .QN(n10456) );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(n10617), .CLK(n10953), 
        .Q(test_so85) );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(n10614), .CLK(n10950), .Q(g2779), .QN(n10026) );
  SDFFX1 DFF_1224_Q_reg ( .D(test_so39), .SI(g2779), .SE(n10652), .CLK(n10988), 
        .Q(g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(n10697), .CLK(n11033), 
        .Q(g7245) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(n10698), .CLK(n11034), 
        .Q(g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(n10604), .CLK(n10940), 
        .Q(g1367), .QN(n10121) );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(n10634), .CLK(n10970), 
        .Q(g5112), .QN(n10489) );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(n10634), .CLK(n10970), 
        .Q(g19), .QN(n10519) );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(n10641), .CLK(n10977), .Q(
        g4145), .QN(n10391) );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(n10641), .CLK(n10977), 
        .Q(g2161) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(n10671), .CLK(n11007), 
        .Q(g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(n10664), .CLK(n11000), 
        .Q(g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(n10652), .CLK(n10988), 
        .Q(test_so86), .QN(DFF_1234_n1) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(n10643), .CLK(n10979), .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(n10663), .CLK(n10999), 
        .Q(g2051), .QN(n10472) );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(n10675), .CLK(n11011), 
        .Q(g1193) );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(n10699), .CLK(n11035), 
        .Q(g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(n10641), .CLK(n10977), 
        .Q(g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(n10641), .CLK(n10977), 
        .Q(g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(n10631), .CLK(n10967), 
        .Q(g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(n10619), .CLK(n10955), 
        .Q(g3594) );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(n10698), .CLK(n11034), 
        .Q(g2999) );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(n10652), .CLK(n10988), 
        .Q(g2303) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(n10682), .CLK(n11018), 
        .Q(g17688), .QN(n10243) );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(n10650), .CLK(n10986), 
        .Q(test_so87), .QN(n10582) );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(n10695), .CLK(n11031), .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(n10695), .CLK(n11031), 
        .Q(g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(n10695), .CLK(n11031), 
        .Q(g546) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(n10646), .CLK(n10982), 
        .Q(g2472) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(n10678), .CLK(n11014), 
        .Q(g5953) );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(n10648), .CLK(n10984), 
        .Q(g8277), .QN(n10059) );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(n10648), .CLK(n10984), 
        .Q(g1740) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(n10698), .CLK(n11034), 
        .Q(g3550) );
  SDFFX1 DFF_1260_Q_reg ( .D(g25683), .SI(g3550), .SE(n10600), .CLK(n10936), 
        .Q(g3845), .QN(n5886) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(n10600), .CLK(n10936), 
        .Q(g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(n10635), .CLK(n10971), 
        .Q(g14635) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(n10609), .CLK(n10945), 
        .Q(test_so88) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(n10615), .CLK(n10951), .Q(g3913), .QN(n10364) );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(n10601), .CLK(n10937), 
        .Q(g10306) );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(n10611), .CLK(n10947), 
        .Q(g1687), .QN(n10068) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(n10663), .CLK(n10999), 
        .Q(g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(g33596), .SI(g2681), .SE(n10663), .CLK(n10999), 
        .Q(g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(n10664), .CLK(n11000), 
        .Q(g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(n10664), .CLK(n11000), 
        .Q(g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(g31895), .SI(g2697), .SE(n10665), .CLK(n11001), 
        .Q(g4417), .QN(n10007) );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(n10666), .CLK(n11002), 
        .Q(g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(n10688), .CLK(n11024), 
        .Q(g1141), .QN(n5691) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(n10688), .CLK(n11024), 
        .Q(g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(n10695), .CLK(n11031), 
        .Q(test_so89), .QN(n10588) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(n10611), .CLK(n10947), .Q(g1710) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(n10621), .CLK(n10957), 
        .Q(g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(n10621), .CLK(n10957), 
        .Q(g3255) );
  SDFFX1 DFF_1281_Q_reg ( .D(g29241), .SI(g3255), .SE(n10620), .CLK(n10956), 
        .Q(g1691), .QN(n10196) );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(n10620), .CLK(n10956), 
        .Q(g2936), .QN(n10401) );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(n10620), .CLK(n10956), 
        .Q(g5644), .QN(n5593) );
  SDFFX1 DFF_1284_Q_reg ( .D(g25707), .SI(g5644), .SE(n10628), .CLK(n10964), 
        .Q(g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(n10628), .CLK(n10964), 
        .Q(g5352), .QN(n10514) );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(n10628), .CLK(n10964), 
        .Q(g8915), .QN(n19033) );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(n10605), .CLK(n10941), 
        .Q(g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(n10686), .CLK(n11022), 
        .Q(g2922), .QN(n10399) );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(n10687), .CLK(n11023), 
        .Q(test_so90) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(n10677), .CLK(n11013), .Q(g5893) );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(n10686), .CLK(n11022), 
        .Q(g16603), .QN(n10233) );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(n10639), .CLK(n10975), 
        .Q(g6617) );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(n10605), .CLK(n10941), 
        .Q(g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(n10601), .CLK(n10937), 
        .Q(g4512) );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(n10599), .CLK(n10935), 
        .Q(g5599) );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(n10623), .CLK(n10959), 
        .Q(g3401) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(n10685), .CLK(n11021), 
        .Q(g4366) );
  SDFFX1 DFF_1300_Q_reg ( .D(test_so26), .SI(g4366), .SE(n10685), .CLK(n11021), 
        .Q(g16722) );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(n10685), .CLK(n11021), 
        .Q(g29214) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g29214), .SE(n10609), .CLK(n10945), 
        .Q(g3129), .QN(n5861) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(n10673), .CLK(n11009), 
        .Q(test_so91) );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(n10667), .CLK(n11003), .Q(g5170), .QN(n10429) );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(n10668), .CLK(n11004), 
        .Q(g26959) );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(n10656), .CLK(n10992), 
        .Q(g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(n10680), .CLK(n11016), 
        .Q(g6299) );
  SDFFX1 DFF_1308_Q_reg ( .D(g7916), .SI(g6299), .SE(n10681), .CLK(n11017), 
        .Q(g8416), .QN(n10050) );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(n10697), .CLK(n11033), 
        .Q(g2079), .QN(n10198) );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(n10628), .CLK(n10964), 
        .Q(g4698), .QN(n5862) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(n10634), .CLK(n10970), 
        .Q(g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(n10646), .CLK(n10982), 
        .Q(g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(n10701), .CLK(n11037), 
        .Q(n9247) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(n10616), .CLK(n10952), 
        .Q(g411) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(n10653), .CLK(n10989), 
        .Q(test_so92) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(n10615), .CLK(n10951), .Q(g3953) );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(n10664), .CLK(n11000), 
        .Q(g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(n10692), .CLK(n11028), 
        .Q(g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(n10692), .CLK(n11028), 
        .Q(n9245) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(n10630), .CLK(n10966), 
        .Q(g1300), .QN(n5483) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(n10630), .CLK(n10966), 
        .Q(g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(n10629), .CLK(n10965), 
        .Q(g5200) );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(n10661), .CLK(n10997), 
        .Q(g4843), .QN(n10478) );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(n10597), .CLK(n10933), 
        .Q(g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(g29249), .SI(g5046), .SE(n10642), .CLK(n10978), 
        .Q(g2250), .QN(n10190) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(n10642), .CLK(n10978), 
        .Q(g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(n10698), .CLK(n11034), 
        .Q(test_so93) );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(n10646), .CLK(n10982), .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(g25734), .SI(g2453), .SE(n10657), .CLK(n10993), 
        .Q(g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(n10657), .CLK(n10993), 
        .Q(g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(n10686), .CLK(n11022), 
        .Q(g2912), .QN(n10398) );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(n10695), .CLK(n11031), 
        .Q(g2357) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(n10695), .CLK(n11031), 
        .Q(g8920), .QN(n19039) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(n10617), .CLK(n10953), 
        .Q(g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(n10624), .CLK(n10960), 
        .Q(g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(n10702), .CLK(n11038), 
        .Q(g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(n10609), .CLK(n10945), 
        .Q(g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(n10612), .CLK(n10948), 
        .Q(g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(n10696), .CLK(n11032), 
        .Q(test_so94), .QN(n10556) );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(n10624), .CLK(n10960), .Q(g4519) );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(n10627), .CLK(n10963), 
        .Q(g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(n10691), .CLK(n11027), 
        .Q(g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(n10640), .CLK(n10976), 
        .Q(g6657) );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(n10640), .CLK(n10976), 
        .Q(g4552) );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(n10614), .CLK(n10950), 
        .Q(g3893) );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(n10621), .CLK(n10957), 
        .Q(g3211), .QN(n10352) );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(n10681), .CLK(n11017), 
        .Q(g13049), .QN(n10361) );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(n10682), .CLK(n11018), 
        .Q(g16624), .QN(n10323) );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(n10598), .CLK(n10934), 
        .Q(g5595) );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(n10619), .CLK(n10955), 
        .Q(g3614) );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(n10645), .CLK(n10981), 
        .Q(test_so95) );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(n10691), .CLK(n11027), .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(n10673), .CLK(n11009), 
        .Q(g16686) );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(n10600), .CLK(n10936), 
        .Q(g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(n10630), .CLK(n10966), 
        .Q(g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(n10640), .CLK(n10976), 
        .Q(g4570) );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(n10627), .CLK(n10963), 
        .Q(g5272) );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(n10662), .CLK(n10998), 
        .Q(g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(n10616), .CLK(n10952), 
        .Q(g728), .QN(n10159) );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(n10679), .CLK(n11015), 
        .Q(g6295) );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(n10603), .CLK(n10939), 
        .Q(g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(n10700), .CLK(n11036), 
        .Q(g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(n10627), .CLK(n10963), 
        .Q(test_so96), .QN(n10577) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(n10645), .CLK(n10981), .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(n10609), .CLK(n10945), 
        .Q(g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(n10618), .CLK(n10954), 
        .Q(g4659), .QN(n10509) );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(n10618), .CLK(n10954), 
        .Q(g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(n10630), .CLK(n10966), 
        .Q(g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(n10655), .CLK(n10991), 
        .Q(g2084), .QN(n10093) );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(n10666), .CLK(n11002), 
        .Q(g3187) );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(n10674), .CLK(n11010), 
        .Q(g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(n10613), .CLK(n10949), 
        .Q(g2583) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(n10610), .CLK(n10946), 
        .Q(n9240) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(n10611), .CLK(n10947), 
        .Q(g1094), .QN(n5697) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(n10658), .CLK(n10994), 
        .Q(test_so97), .QN(n10592) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(n10625), .CLK(n10961), .Q(g4284) );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(n10666), .CLK(n11002), 
        .Q(g3191) );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(n10670), .CLK(n11006), 
        .Q(g4239), .QN(n10104) );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(n10688), .CLK(n11024), 
        .Q(g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(n10606), .CLK(n10942), 
        .Q(g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(n10606), .CLK(n10942), 
        .Q(g534) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(n10671), .CLK(n11007), 
        .Q(g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(n10675), .CLK(n11011), 
        .Q(g2004) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(n10647), .CLK(n10983), 
        .Q(g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(n10670), .CLK(n11006), 
        .Q(g5456), .QN(n10052) );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(n10640), .CLK(n10976), 
        .Q(n6007), .QN(n10564) );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(n10701), .CLK(n11037), 
        .Q(test_so98), .QN(n10591) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(n10690), .CLK(n11026), .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(n10628), .CLK(n10964), 
        .Q(g5348), .QN(n10381) );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(n10699), .CLK(n11035), 
        .Q(g3223) );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(n10620), .CLK(n10956), 
        .Q(g2970), .QN(n10397) );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(n10620), .CLK(n10956), 
        .Q(g5698), .QN(n10496) );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(n10629), .CLK(n10965), 
        .Q(g5260) );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(n10629), .CLK(n10965), 
        .Q(g1521), .QN(n5577) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(n10618), .CLK(n10954), 
        .Q(g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(n10609), .CLK(n10945), 
        .Q(g3115), .QN(n10485) );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(n10673), .CLK(n11009), 
        .Q(g3251) );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(n10673), .CLK(n11009), 
        .Q(g12832) );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(n10673), .CLK(n11009), 
        .Q(test_so99), .QN(n10551) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(n10655), .CLK(
        n10991), .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(n10624), .CLK(n10960), 
        .Q(g8342), .QN(n10036) );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(n10624), .CLK(n10960), 
        .Q(g4515), .QN(n10434) );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(n10652), .CLK(n10988), 
        .Q(g8787), .QN(n10142) );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(n10624), .CLK(n10960), 
        .Q(g4300) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(n10611), .CLK(n10947), 
        .Q(n9236) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(n10611), .CLK(n10947), 
        .Q(g1379), .QN(n10089) );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(n10633), .CLK(n10969), 
        .Q(g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(n10659), .CLK(n10995), 
        .Q(g1878) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(n10599), .CLK(n10935), 
        .Q(g5619) );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(n10601), .CLK(n10937), 
        .Q(g71) );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(n10654), .CLK(n10990), .Q(
        test_so100) );
  SDFFX1 DFF_748_Q_reg ( .D(n1340), .SI(g4704), .SE(n10668), .CLK(n11004), .Q(
        g22), .QN(n10527) );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(n10679), .CLK(n11015), 
        .Q(g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(n10662), .CLK(n10998), .Q(
        g2729), .QN(n10520) );
  HADDX1 Trojan_U1_1_30 ( .A0(counter_30), .B0(carry_30), .C1(carry_31), .SO(
        N31) );
  HADDX1 Trojan_U1_1_4 ( .A0(counter_4), .B0(carry_4), .C1(carry_5), .SO(N5)
         );
  HADDX1 Trojan_U1_1_5 ( .A0(counter_5), .B0(carry_5), .C1(carry_6), .SO(N6)
         );
  HADDX1 Trojan_U1_1_6 ( .A0(counter_6), .B0(carry_6), .C1(carry_7), .SO(N7)
         );
  HADDX1 Trojan_U1_1_7 ( .A0(counter_7), .B0(carry_7), .C1(carry_8), .SO(N8)
         );
  HADDX1 Trojan_U1_1_8 ( .A0(counter_8), .B0(carry_8), .C1(carry_9), .SO(N9)
         );
  HADDX1 Trojan_U1_1_9 ( .A0(counter_9), .B0(carry_9), .C1(carry_10), .SO(N10)
         );
  HADDX1 Trojan_U1_1_10 ( .A0(counter_10), .B0(carry_10), .C1(carry_11), .SO(
        N11) );
  HADDX1 Trojan_U1_1_11 ( .A0(counter_11), .B0(carry_11), .C1(carry_12), .SO(
        N12) );
  HADDX1 Trojan_U1_1_12 ( .A0(counter_12), .B0(carry_12), .C1(carry_13), .SO(
        N13) );
  HADDX1 Trojan_U1_1_13 ( .A0(counter_13), .B0(carry_13), .C1(carry_14), .SO(
        N14) );
  HADDX1 Trojan_U1_1_14 ( .A0(counter_14), .B0(carry_14), .C1(carry_15), .SO(
        N15) );
  HADDX1 Trojan_U1_1_22 ( .A0(counter_22), .B0(carry_22), .C1(carry_23), .SO(
        N23) );
  HADDX1 Trojan_U1_1_23 ( .A0(counter_23), .B0(carry_23), .C1(carry_24), .SO(
        N24) );
  HADDX1 Trojan_U1_1_24 ( .A0(counter_24), .B0(carry_24), .C1(carry_25), .SO(
        N25) );
  HADDX1 Trojan_U1_1_25 ( .A0(counter_25), .B0(carry_25), .C1(carry_26), .SO(
        N26) );
  HADDX1 Trojan_U1_1_1 ( .A0(counter_1), .B0(counter_0), .C1(carry_2), .SO(N2)
         );
  HADDX1 Trojan_U1_1_2 ( .A0(counter_2), .B0(carry_2), .C1(carry_3), .SO(N3)
         );
  HADDX1 Trojan_U1_1_3 ( .A0(counter_3), .B0(carry_3), .C1(carry_4), .SO(N4)
         );
  HADDX1 Trojan_U1_1_15 ( .A0(counter_15), .B0(carry_15), .C1(carry_16), .SO(
        N16) );
  HADDX1 Trojan_U1_1_16 ( .A0(counter_16), .B0(carry_16), .C1(carry_17), .SO(
        N17) );
  HADDX1 Trojan_U1_1_17 ( .A0(counter_17), .B0(carry_17), .C1(carry_18), .SO(
        N18) );
  HADDX1 Trojan_U1_1_18 ( .A0(counter_18), .B0(carry_18), .C1(carry_19), .SO(
        N19) );
  HADDX1 Trojan_U1_1_19 ( .A0(counter_19), .B0(carry_19), .C1(carry_20), .SO(
        N20) );
  HADDX1 Trojan_U1_1_20 ( .A0(counter_20), .B0(carry_20), .C1(carry_21), .SO(
        N21) );
  HADDX1 Trojan_U1_1_21 ( .A0(counter_21), .B0(carry_21), .C1(carry_22), .SO(
        N22) );
  HADDX1 Trojan_U1_1_26 ( .A0(counter_26), .B0(carry_26), .C1(carry_27), .SO(
        N27) );
  HADDX1 Trojan_U1_1_27 ( .A0(counter_27), .B0(carry_27), .C1(carry_28), .SO(
        N28) );
  HADDX1 Trojan_U1_1_28 ( .A0(counter_28), .B0(carry_28), .C1(carry_29), .SO(
        N29) );
  HADDX1 Trojan_U1_1_29 ( .A0(counter_29), .B0(carry_29), .C1(carry_30), .SO(
        N30) );
  INVX0 Trojan_U1 ( .INP(counter_0), .ZN(N1) );
  XOR2X1 Trojan_U2 ( .IN1(carry_31), .IN2(counter_31), .Q(N32) );
  DFFARX1 Trojan_counter_reg_31_ ( .D(N32), .CLK(n37), .RSTB(n10596), .Q(
        counter_31), .QN(n73) );
  DFFARX1 Trojan_counter_reg_1_ ( .D(N2), .CLK(n37), .RSTB(n10595), .Q(
        counter_1) );
  DFFARX1 Trojan_counter_reg_2_ ( .D(N3), .CLK(n37), .RSTB(n87), .Q(counter_2)
         );
  DFFARX1 Trojan_counter_reg_3_ ( .D(N4), .CLK(n37), .RSTB(n10596), .Q(
        counter_3), .QN(n86) );
  DFFARX1 Trojan_counter_reg_15_ ( .D(N16), .CLK(n37), .RSTB(n10595), .Q(
        counter_15), .QN(n85) );
  DFFARX1 Trojan_counter_reg_16_ ( .D(N17), .CLK(n37), .RSTB(n87), .Q(
        counter_16), .QN(n84) );
  DFFARX1 Trojan_counter_reg_17_ ( .D(N18), .CLK(n37), .RSTB(n10596), .Q(
        counter_17), .QN(n83) );
  DFFARX1 Trojan_counter_reg_18_ ( .D(N19), .CLK(n37), .RSTB(n10595), .Q(
        counter_18), .QN(n82) );
  DFFARX1 Trojan_counter_reg_19_ ( .D(N20), .CLK(n37), .RSTB(n87), .Q(
        counter_19), .QN(n81) );
  DFFARX1 Trojan_counter_reg_20_ ( .D(N21), .CLK(n37), .RSTB(n10596), .Q(
        counter_20), .QN(n80) );
  DFFARX1 Trojan_counter_reg_21_ ( .D(N22), .CLK(n37), .RSTB(n10595), .Q(
        counter_21), .QN(n79) );
  DFFARX1 Trojan_counter_reg_26_ ( .D(N27), .CLK(n37), .RSTB(n87), .Q(
        counter_26), .QN(n78) );
  DFFARX1 Trojan_counter_reg_27_ ( .D(N28), .CLK(n37), .RSTB(n10596), .Q(
        counter_27), .QN(n77) );
  DFFARX1 Trojan_counter_reg_28_ ( .D(N29), .CLK(n37), .RSTB(n10595), .Q(
        counter_28), .QN(n76) );
  DFFARX1 Trojan_counter_reg_29_ ( .D(N30), .CLK(n37), .RSTB(n87), .Q(
        counter_29), .QN(n75) );
  DFFARX1 Trojan_counter_reg_30_ ( .D(N31), .CLK(n37), .RSTB(n10596), .Q(
        counter_30), .QN(n74) );
  DFFARX1 Trojan_counter_reg_7_ ( .D(N8), .CLK(n37), .RSTB(n10595), .Q(
        counter_7) );
  DFFARX1 Trojan_counter_reg_11_ ( .D(N12), .CLK(n37), .RSTB(n87), .Q(
        counter_11) );
  DFFARX1 Trojan_counter_reg_25_ ( .D(N26), .CLK(n37), .RSTB(n10596), .Q(
        counter_25) );
  DFFARX1 Trojan_counter_reg_6_ ( .D(N7), .CLK(n37), .RSTB(n10595), .Q(
        counter_6) );
  DFFARX1 Trojan_counter_reg_10_ ( .D(N11), .CLK(n37), .RSTB(n87), .Q(
        counter_10) );
  DFFARX1 Trojan_counter_reg_12_ ( .D(N13), .CLK(n37), .RSTB(n10596), .Q(
        counter_12) );
  DFFARX1 Trojan_counter_reg_24_ ( .D(N25), .CLK(n37), .RSTB(n10595), .Q(
        counter_24) );
  DFFARX1 Trojan_counter_reg_4_ ( .D(N5), .CLK(n37), .RSTB(n87), .Q(counter_4)
         );
  DFFARX1 Trojan_counter_reg_5_ ( .D(N6), .CLK(n37), .RSTB(n10596), .Q(
        counter_5) );
  DFFARX1 Trojan_counter_reg_9_ ( .D(N10), .CLK(n37), .RSTB(n10595), .Q(
        counter_9) );
  DFFARX1 Trojan_counter_reg_14_ ( .D(N15), .CLK(n37), .RSTB(n87), .Q(
        counter_14) );
  DFFARX1 Trojan_counter_reg_23_ ( .D(N24), .CLK(n37), .RSTB(n10596), .Q(
        counter_23) );
  DFFARX1 Trojan_counter_reg_8_ ( .D(N9), .CLK(n37), .RSTB(n10595), .Q(
        counter_8) );
  DFFARX1 Trojan_counter_reg_13_ ( .D(N14), .CLK(n37), .RSTB(n87), .Q(
        counter_13) );
  DFFARX1 Trojan_counter_reg_22_ ( .D(N23), .CLK(n37), .RSTB(n10596), .Q(
        counter_22) );
  DFFARX1 Trojan_counter_reg_0_ ( .D(N1), .CLK(n37), .RSTB(n10595), .Q(
        counter_0) );
  NAND4X0 Trojan_U14 ( .IN1(n3180), .IN2(n3121), .IN3(n2461), .IN4(n58), .QN(
        n87) );
  INVX0 Trojan_U15 ( .INP(n59), .ZN(n58) );
  NOR4X0 Trojan_U16 ( .IN1(n3180), .IN2(n3121), .IN3(n2461), .IN4(n59), .QN(
        n37) );
  NAND3X0 Trojan_U17 ( .IN1(n108), .IN2(n5111), .IN3(n60), .QN(n59) );
  AND3X1 Trojan_U18 ( .IN1(n2396), .IN2(n44), .IN3(n10534), .Q(n60) );
  NOR4X0 Trojan_U19 ( .IN1(n61), .IN2(n62), .IN3(n63), .IN4(n64), .QN(
        Trigger_out) );
  NAND4X0 Trojan_U20 ( .IN1(n78), .IN2(n77), .IN3(n76), .IN4(n75), .QN(n64) );
  NAND4X0 Trojan_U21 ( .IN1(n74), .IN2(n73), .IN3(counter_6), .IN4(counter_5), 
        .QN(n63) );
  NAND4X0 Trojan_U22 ( .IN1(n80), .IN2(n79), .IN3(n81), .IN4(n65), .QN(n62) );
  NOR4X0 Trojan_U23 ( .IN1(counter_25), .IN2(counter_24), .IN3(counter_23), 
        .IN4(counter_22), .QN(n65) );
  NAND4X0 Trojan_U24 ( .IN1(n66), .IN2(n67), .IN3(n68), .IN4(n69), .QN(n61) );
  NOR4X0 Trojan_U25 ( .IN1(n70), .IN2(counter_12), .IN3(counter_14), .IN4(
        counter_13), .QN(n69) );
  NAND4X0 Trojan_U26 ( .IN1(n85), .IN2(n84), .IN3(n83), .IN4(n82), .QN(n70) );
  NOR4X0 Trojan_U27 ( .IN1(counter_11), .IN2(counter_10), .IN3(counter_9), 
        .IN4(counter_8), .QN(n68) );
  MUX21X1 Trojan_U28 ( .IN1(n71), .IN2(n72), .S(n86), .Q(n67) );
  OA21X1 Trojan_U29 ( .IN1(counter_1), .IN2(counter_0), .IN3(counter_2), .Q(
        n72) );
  NAND2X0 Trojan_U30 ( .IN1(counter_2), .IN2(counter_1), .QN(n71) );
  NOR2X0 Trojan_U31 ( .IN1(counter_7), .IN2(counter_4), .QN(n66) );
  MUX21X1 Trojan_Paylod ( .IN1(g10122_Tj), .IN2(g25715), .S(Trigger_out), .Q(
        g10122) );
  INVX0 U10532 ( .INP(n87), .ZN(n10594) );
  INVX0 U10533 ( .INP(n10594), .ZN(n10595) );
  INVX0 U10534 ( .INP(n10594), .ZN(n10596) );
  NBUFFX2 U10535 ( .INP(n10725), .Z(n10598) );
  NBUFFX2 U10536 ( .INP(n10725), .Z(n10597) );
  NBUFFX2 U10537 ( .INP(n10712), .Z(n10660) );
  NBUFFX2 U10538 ( .INP(n10721), .Z(n10614) );
  NBUFFX2 U10539 ( .INP(n10705), .Z(n10695) );
  NBUFFX2 U10540 ( .INP(n10719), .Z(n10627) );
  NBUFFX2 U10541 ( .INP(n10719), .Z(n10624) );
  NBUFFX2 U10542 ( .INP(n10711), .Z(n10668) );
  NBUFFX2 U10543 ( .INP(n10719), .Z(n10625) );
  NBUFFX2 U10544 ( .INP(n10721), .Z(n10617) );
  NBUFFX2 U10545 ( .INP(n10707), .Z(n10688) );
  NBUFFX2 U10546 ( .INP(n10716), .Z(n10639) );
  NBUFFX2 U10547 ( .INP(n10710), .Z(n10669) );
  NBUFFX2 U10548 ( .INP(n10712), .Z(n10659) );
  NBUFFX2 U10549 ( .INP(n10715), .Z(n10646) );
  NBUFFX2 U10550 ( .INP(n10720), .Z(n10620) );
  NBUFFX2 U10551 ( .INP(n10724), .Z(n10600) );
  NBUFFX2 U10552 ( .INP(n10707), .Z(n10685) );
  NBUFFX2 U10553 ( .INP(n10723), .Z(n10604) );
  NBUFFX2 U10554 ( .INP(n10717), .Z(n10638) );
  NBUFFX2 U10555 ( .INP(n10710), .Z(n10673) );
  NBUFFX2 U10556 ( .INP(n10724), .Z(n10601) );
  NBUFFX2 U10557 ( .INP(n10712), .Z(n10662) );
  NBUFFX2 U10558 ( .INP(n10713), .Z(n10654) );
  NBUFFX2 U10559 ( .INP(n10715), .Z(n10645) );
  NBUFFX2 U10560 ( .INP(n10718), .Z(n10631) );
  NBUFFX2 U10561 ( .INP(n10708), .Z(n10679) );
  NBUFFX2 U10562 ( .INP(n10708), .Z(n10680) );
  NBUFFX2 U10563 ( .INP(n10714), .Z(n10650) );
  NBUFFX2 U10564 ( .INP(n10708), .Z(n10682) );
  NBUFFX2 U10565 ( .INP(n10708), .Z(n10683) );
  NBUFFX2 U10566 ( .INP(n10723), .Z(n10606) );
  NBUFFX2 U10567 ( .INP(n10716), .Z(n10641) );
  NBUFFX2 U10568 ( .INP(n10718), .Z(n10630) );
  NBUFFX2 U10569 ( .INP(n10705), .Z(n10694) );
  NBUFFX2 U10570 ( .INP(n10715), .Z(n10647) );
  NBUFFX2 U10571 ( .INP(n10713), .Z(n10658) );
  NBUFFX2 U10572 ( .INP(n10722), .Z(n10609) );
  NBUFFX2 U10573 ( .INP(n10717), .Z(n10634) );
  NBUFFX2 U10574 ( .INP(n10719), .Z(n10628) );
  NBUFFX2 U10575 ( .INP(n10718), .Z(n10632) );
  NBUFFX2 U10576 ( .INP(n10706), .Z(n10689) );
  NBUFFX2 U10577 ( .INP(n10711), .Z(n10667) );
  NBUFFX2 U10578 ( .INP(n10715), .Z(n10644) );
  NBUFFX2 U10579 ( .INP(n10710), .Z(n10671) );
  NBUFFX2 U10580 ( .INP(n10709), .Z(n10676) );
  NBUFFX2 U10581 ( .INP(n10708), .Z(n10681) );
  NBUFFX2 U10582 ( .INP(n10718), .Z(n10629) );
  NBUFFX2 U10583 ( .INP(n10707), .Z(n10687) );
  NBUFFX2 U10584 ( .INP(n10716), .Z(n10640) );
  NBUFFX2 U10585 ( .INP(n10721), .Z(n10615) );
  NBUFFX2 U10586 ( .INP(n10716), .Z(n10643) );
  NBUFFX2 U10587 ( .INP(n10723), .Z(n10607) );
  NBUFFX2 U10588 ( .INP(n10706), .Z(n10693) );
  NBUFFX2 U10589 ( .INP(n10720), .Z(n10621) );
  NBUFFX2 U10590 ( .INP(n10713), .Z(n10655) );
  NBUFFX2 U10591 ( .INP(n10710), .Z(n10672) );
  NBUFFX2 U10592 ( .INP(n10710), .Z(n10670) );
  NBUFFX2 U10593 ( .INP(n10722), .Z(n10610) );
  NBUFFX2 U10594 ( .INP(n10714), .Z(n10649) );
  NBUFFX2 U10595 ( .INP(n10717), .Z(n10637) );
  NBUFFX2 U10596 ( .INP(n10707), .Z(n10684) );
  NBUFFX2 U10597 ( .INP(n10722), .Z(n10613) );
  NBUFFX2 U10598 ( .INP(n10722), .Z(n10612) );
  NBUFFX2 U10599 ( .INP(n10711), .Z(n10664) );
  NBUFFX2 U10600 ( .INP(n10720), .Z(n10619) );
  NBUFFX2 U10601 ( .INP(n10705), .Z(n10698) );
  NBUFFX2 U10602 ( .INP(n10724), .Z(n10599) );
  NBUFFX2 U10603 ( .INP(n10723), .Z(n10608) );
  NBUFFX2 U10604 ( .INP(n10724), .Z(n10602) );
  NBUFFX2 U10605 ( .INP(n10712), .Z(n10661) );
  NBUFFX2 U10606 ( .INP(n10713), .Z(n10657) );
  NBUFFX2 U10607 ( .INP(n10724), .Z(n10603) );
  NBUFFX2 U10608 ( .INP(n10709), .Z(n10674) );
  NBUFFX2 U10609 ( .INP(n10717), .Z(n10636) );
  NBUFFX2 U10610 ( .INP(n10709), .Z(n10677) );
  NBUFFX2 U10611 ( .INP(n10716), .Z(n10642) );
  NBUFFX2 U10612 ( .INP(n10711), .Z(n10666) );
  NBUFFX2 U10613 ( .INP(n10718), .Z(n10633) );
  NBUFFX2 U10614 ( .INP(n10722), .Z(n10611) );
  NBUFFX2 U10615 ( .INP(n10714), .Z(n10651) );
  NBUFFX2 U10616 ( .INP(n10705), .Z(n10696) );
  NBUFFX2 U10617 ( .INP(n10713), .Z(n10656) );
  NBUFFX2 U10618 ( .INP(n10721), .Z(n10618) );
  NBUFFX2 U10619 ( .INP(n10709), .Z(n10675) );
  NBUFFX2 U10620 ( .INP(n10720), .Z(n10623) );
  NBUFFX2 U10621 ( .INP(n10714), .Z(n10653) );
  NBUFFX2 U10622 ( .INP(n10706), .Z(n10690) );
  NBUFFX2 U10623 ( .INP(n10709), .Z(n10678) );
  NBUFFX2 U10624 ( .INP(n10715), .Z(n10648) );
  NBUFFX2 U10625 ( .INP(n10707), .Z(n10686) );
  NBUFFX2 U10626 ( .INP(n10711), .Z(n10665) );
  NBUFFX2 U10627 ( .INP(n10719), .Z(n10626) );
  NBUFFX2 U10628 ( .INP(n10706), .Z(n10691) );
  NBUFFX2 U10629 ( .INP(n10721), .Z(n10616) );
  NBUFFX2 U10630 ( .INP(n10720), .Z(n10622) );
  NBUFFX2 U10631 ( .INP(n10706), .Z(n10692) );
  NBUFFX2 U10632 ( .INP(n10712), .Z(n10663) );
  NBUFFX2 U10633 ( .INP(n10717), .Z(n10635) );
  NBUFFX2 U10634 ( .INP(n10714), .Z(n10652) );
  NBUFFX2 U10635 ( .INP(n10705), .Z(n10697) );
  NBUFFX2 U10636 ( .INP(n10723), .Z(n10605) );
  NBUFFX2 U10637 ( .INP(n11061), .Z(n10934) );
  NBUFFX2 U10638 ( .INP(n11061), .Z(n10933) );
  NBUFFX2 U10639 ( .INP(n11048), .Z(n10996) );
  NBUFFX2 U10640 ( .INP(n11057), .Z(n10950) );
  NBUFFX2 U10641 ( .INP(n11041), .Z(n11031) );
  NBUFFX2 U10642 ( .INP(n11055), .Z(n10963) );
  NBUFFX2 U10643 ( .INP(n11055), .Z(n10960) );
  NBUFFX2 U10644 ( .INP(n11047), .Z(n11004) );
  NBUFFX2 U10645 ( .INP(n11055), .Z(n10961) );
  NBUFFX2 U10646 ( .INP(n11057), .Z(n10953) );
  NBUFFX2 U10647 ( .INP(n11043), .Z(n11024) );
  NBUFFX2 U10648 ( .INP(n11052), .Z(n10975) );
  NBUFFX2 U10649 ( .INP(n11046), .Z(n11005) );
  NBUFFX2 U10650 ( .INP(n11048), .Z(n10995) );
  NBUFFX2 U10651 ( .INP(n11051), .Z(n10982) );
  NBUFFX2 U10652 ( .INP(n11056), .Z(n10956) );
  NBUFFX2 U10653 ( .INP(n11060), .Z(n10936) );
  NBUFFX2 U10654 ( .INP(n11043), .Z(n11021) );
  NBUFFX2 U10655 ( .INP(n11059), .Z(n10940) );
  NBUFFX2 U10656 ( .INP(n11053), .Z(n10974) );
  NBUFFX2 U10657 ( .INP(n11046), .Z(n11009) );
  NBUFFX2 U10658 ( .INP(n11060), .Z(n10937) );
  NBUFFX2 U10659 ( .INP(n11048), .Z(n10998) );
  NBUFFX2 U10660 ( .INP(n11049), .Z(n10990) );
  NBUFFX2 U10661 ( .INP(n11051), .Z(n10981) );
  NBUFFX2 U10662 ( .INP(n11054), .Z(n10967) );
  NBUFFX2 U10663 ( .INP(n11044), .Z(n11015) );
  NBUFFX2 U10664 ( .INP(n11044), .Z(n11016) );
  NBUFFX2 U10665 ( .INP(n11050), .Z(n10986) );
  NBUFFX2 U10666 ( .INP(n11044), .Z(n11018) );
  NBUFFX2 U10667 ( .INP(n11044), .Z(n11019) );
  NBUFFX2 U10668 ( .INP(n11059), .Z(n10942) );
  NBUFFX2 U10669 ( .INP(n11052), .Z(n10977) );
  NBUFFX2 U10670 ( .INP(n11054), .Z(n10966) );
  NBUFFX2 U10671 ( .INP(n11041), .Z(n11030) );
  NBUFFX2 U10672 ( .INP(n11051), .Z(n10983) );
  NBUFFX2 U10673 ( .INP(n11049), .Z(n10994) );
  NBUFFX2 U10674 ( .INP(n11058), .Z(n10945) );
  NBUFFX2 U10675 ( .INP(n11053), .Z(n10970) );
  NBUFFX2 U10676 ( .INP(n11055), .Z(n10964) );
  NBUFFX2 U10677 ( .INP(n11054), .Z(n10968) );
  NBUFFX2 U10678 ( .INP(n11042), .Z(n11025) );
  NBUFFX2 U10679 ( .INP(n11047), .Z(n11003) );
  NBUFFX2 U10680 ( .INP(n11051), .Z(n10980) );
  NBUFFX2 U10681 ( .INP(n11046), .Z(n11007) );
  NBUFFX2 U10682 ( .INP(n11045), .Z(n11012) );
  NBUFFX2 U10683 ( .INP(n11044), .Z(n11017) );
  NBUFFX2 U10684 ( .INP(n11054), .Z(n10965) );
  NBUFFX2 U10685 ( .INP(n11043), .Z(n11023) );
  NBUFFX2 U10686 ( .INP(n11052), .Z(n10976) );
  NBUFFX2 U10687 ( .INP(n11057), .Z(n10951) );
  NBUFFX2 U10688 ( .INP(n11052), .Z(n10979) );
  NBUFFX2 U10689 ( .INP(n11059), .Z(n10943) );
  NBUFFX2 U10690 ( .INP(n11042), .Z(n11029) );
  NBUFFX2 U10691 ( .INP(n11056), .Z(n10957) );
  NBUFFX2 U10692 ( .INP(n11049), .Z(n10991) );
  NBUFFX2 U10693 ( .INP(n11046), .Z(n11008) );
  NBUFFX2 U10694 ( .INP(n11046), .Z(n11006) );
  NBUFFX2 U10695 ( .INP(n11058), .Z(n10946) );
  NBUFFX2 U10696 ( .INP(n11050), .Z(n10985) );
  NBUFFX2 U10697 ( .INP(n11053), .Z(n10973) );
  NBUFFX2 U10698 ( .INP(n11043), .Z(n11020) );
  NBUFFX2 U10699 ( .INP(n11058), .Z(n10949) );
  NBUFFX2 U10700 ( .INP(n11058), .Z(n10948) );
  NBUFFX2 U10701 ( .INP(n11047), .Z(n11000) );
  NBUFFX2 U10702 ( .INP(n11056), .Z(n10955) );
  NBUFFX2 U10703 ( .INP(n11041), .Z(n11034) );
  NBUFFX2 U10704 ( .INP(n11060), .Z(n10935) );
  NBUFFX2 U10705 ( .INP(n11059), .Z(n10944) );
  NBUFFX2 U10706 ( .INP(n11060), .Z(n10938) );
  NBUFFX2 U10707 ( .INP(n11048), .Z(n10997) );
  NBUFFX2 U10708 ( .INP(n11049), .Z(n10993) );
  NBUFFX2 U10709 ( .INP(n11060), .Z(n10939) );
  NBUFFX2 U10710 ( .INP(n11045), .Z(n11010) );
  NBUFFX2 U10711 ( .INP(n11053), .Z(n10972) );
  NBUFFX2 U10712 ( .INP(n11045), .Z(n11013) );
  NBUFFX2 U10713 ( .INP(n11052), .Z(n10978) );
  NBUFFX2 U10714 ( .INP(n11047), .Z(n11002) );
  NBUFFX2 U10715 ( .INP(n11054), .Z(n10969) );
  NBUFFX2 U10716 ( .INP(n11058), .Z(n10947) );
  NBUFFX2 U10717 ( .INP(n11050), .Z(n10987) );
  NBUFFX2 U10718 ( .INP(n11041), .Z(n11032) );
  NBUFFX2 U10719 ( .INP(n11049), .Z(n10992) );
  NBUFFX2 U10720 ( .INP(n11057), .Z(n10954) );
  NBUFFX2 U10721 ( .INP(n11045), .Z(n11011) );
  NBUFFX2 U10722 ( .INP(n11056), .Z(n10959) );
  NBUFFX2 U10723 ( .INP(n11050), .Z(n10989) );
  NBUFFX2 U10724 ( .INP(n11042), .Z(n11026) );
  NBUFFX2 U10725 ( .INP(n11045), .Z(n11014) );
  NBUFFX2 U10726 ( .INP(n11051), .Z(n10984) );
  NBUFFX2 U10727 ( .INP(n11043), .Z(n11022) );
  NBUFFX2 U10728 ( .INP(n11047), .Z(n11001) );
  NBUFFX2 U10729 ( .INP(n11055), .Z(n10962) );
  NBUFFX2 U10730 ( .INP(n11042), .Z(n11027) );
  NBUFFX2 U10731 ( .INP(n11057), .Z(n10952) );
  NBUFFX2 U10732 ( .INP(n11056), .Z(n10958) );
  NBUFFX2 U10733 ( .INP(n11042), .Z(n11028) );
  NBUFFX2 U10734 ( .INP(n11048), .Z(n10999) );
  NBUFFX2 U10735 ( .INP(n11053), .Z(n10971) );
  NBUFFX2 U10736 ( .INP(n11050), .Z(n10988) );
  NBUFFX2 U10737 ( .INP(n11041), .Z(n11033) );
  NBUFFX2 U10738 ( .INP(n11059), .Z(n10941) );
  NBUFFX2 U10739 ( .INP(n10704), .Z(n10700) );
  NBUFFX2 U10740 ( .INP(n10704), .Z(n10702) );
  NBUFFX2 U10741 ( .INP(n10704), .Z(n10701) );
  NBUFFX2 U10742 ( .INP(n10704), .Z(n10699) );
  NBUFFX2 U10743 ( .INP(n11040), .Z(n11036) );
  NBUFFX2 U10744 ( .INP(n11040), .Z(n11038) );
  NBUFFX2 U10745 ( .INP(n11040), .Z(n11037) );
  NBUFFX2 U10746 ( .INP(n11040), .Z(n11035) );
  NBUFFX2 U10747 ( .INP(n10704), .Z(n10703) );
  NBUFFX2 U10748 ( .INP(n11040), .Z(n11039) );
  NBUFFX2 U10749 ( .INP(n10733), .Z(n10704) );
  NBUFFX2 U10750 ( .INP(n10732), .Z(n10705) );
  NBUFFX2 U10751 ( .INP(n10732), .Z(n10706) );
  NBUFFX2 U10752 ( .INP(n10732), .Z(n10707) );
  NBUFFX2 U10753 ( .INP(n10731), .Z(n10708) );
  NBUFFX2 U10754 ( .INP(n10731), .Z(n10709) );
  NBUFFX2 U10755 ( .INP(n10731), .Z(n10710) );
  NBUFFX2 U10756 ( .INP(n10730), .Z(n10711) );
  NBUFFX2 U10757 ( .INP(n10730), .Z(n10712) );
  NBUFFX2 U10758 ( .INP(n10730), .Z(n10713) );
  NBUFFX2 U10759 ( .INP(n10729), .Z(n10714) );
  NBUFFX2 U10760 ( .INP(n10729), .Z(n10715) );
  NBUFFX2 U10761 ( .INP(n10729), .Z(n10716) );
  NBUFFX2 U10762 ( .INP(n10728), .Z(n10717) );
  NBUFFX2 U10763 ( .INP(n10728), .Z(n10718) );
  NBUFFX2 U10764 ( .INP(n10728), .Z(n10719) );
  NBUFFX2 U10765 ( .INP(n10727), .Z(n10720) );
  NBUFFX2 U10766 ( .INP(n10727), .Z(n10721) );
  NBUFFX2 U10767 ( .INP(n10727), .Z(n10722) );
  NBUFFX2 U10768 ( .INP(n10726), .Z(n10723) );
  NBUFFX2 U10769 ( .INP(n10726), .Z(n10724) );
  NBUFFX2 U10770 ( .INP(n10726), .Z(n10725) );
  NBUFFX2 U10771 ( .INP(n10736), .Z(n10726) );
  NBUFFX2 U10772 ( .INP(n10736), .Z(n10727) );
  NBUFFX2 U10773 ( .INP(n10735), .Z(n10728) );
  NBUFFX2 U10774 ( .INP(n10735), .Z(n10729) );
  NBUFFX2 U10775 ( .INP(n10735), .Z(n10730) );
  NBUFFX2 U10776 ( .INP(n10734), .Z(n10731) );
  NBUFFX2 U10777 ( .INP(n10734), .Z(n10732) );
  NBUFFX2 U10778 ( .INP(n10734), .Z(n10733) );
  NBUFFX2 U10779 ( .INP(test_se), .Z(n10734) );
  NBUFFX2 U10780 ( .INP(test_se), .Z(n10735) );
  NBUFFX2 U10781 ( .INP(test_se), .Z(n10736) );
  NBUFFX2 U10782 ( .INP(n10858), .Z(n10737) );
  NBUFFX2 U10783 ( .INP(n10858), .Z(n10738) );
  NBUFFX2 U10784 ( .INP(n10857), .Z(n10739) );
  NBUFFX2 U10785 ( .INP(n10857), .Z(n10740) );
  NBUFFX2 U10786 ( .INP(n10857), .Z(n10741) );
  NBUFFX2 U10787 ( .INP(n10856), .Z(n10742) );
  NBUFFX2 U10788 ( .INP(n10856), .Z(n10743) );
  NBUFFX2 U10789 ( .INP(n10856), .Z(n10744) );
  NBUFFX2 U10790 ( .INP(n10855), .Z(n10745) );
  NBUFFX2 U10791 ( .INP(n10855), .Z(n10746) );
  NBUFFX2 U10792 ( .INP(n10855), .Z(n10747) );
  NBUFFX2 U10793 ( .INP(n10854), .Z(n10748) );
  NBUFFX2 U10794 ( .INP(n10854), .Z(n10749) );
  NBUFFX2 U10795 ( .INP(n10854), .Z(n10750) );
  NBUFFX2 U10796 ( .INP(n10853), .Z(n10751) );
  NBUFFX2 U10797 ( .INP(n10853), .Z(n10752) );
  NBUFFX2 U10798 ( .INP(n10853), .Z(n10753) );
  NBUFFX2 U10799 ( .INP(n10852), .Z(n10754) );
  NBUFFX2 U10800 ( .INP(n10852), .Z(n10755) );
  NBUFFX2 U10801 ( .INP(n10852), .Z(n10756) );
  NBUFFX2 U10802 ( .INP(n10851), .Z(n10757) );
  NBUFFX2 U10803 ( .INP(n10851), .Z(n10758) );
  NBUFFX2 U10804 ( .INP(n10851), .Z(n10759) );
  NBUFFX2 U10805 ( .INP(n10850), .Z(n10760) );
  NBUFFX2 U10806 ( .INP(n10850), .Z(n10761) );
  NBUFFX2 U10807 ( .INP(n10850), .Z(n10762) );
  NBUFFX2 U10808 ( .INP(n10849), .Z(n10763) );
  NBUFFX2 U10809 ( .INP(n10849), .Z(n10764) );
  NBUFFX2 U10810 ( .INP(n10849), .Z(n10765) );
  NBUFFX2 U10811 ( .INP(n10848), .Z(n10766) );
  NBUFFX2 U10812 ( .INP(n10848), .Z(n10767) );
  NBUFFX2 U10813 ( .INP(n10848), .Z(n10768) );
  NBUFFX2 U10814 ( .INP(n10847), .Z(n10769) );
  NBUFFX2 U10815 ( .INP(n10847), .Z(n10770) );
  NBUFFX2 U10816 ( .INP(n10847), .Z(n10771) );
  NBUFFX2 U10817 ( .INP(n10846), .Z(n10772) );
  NBUFFX2 U10818 ( .INP(n10846), .Z(n10773) );
  NBUFFX2 U10819 ( .INP(n10846), .Z(n10774) );
  NBUFFX2 U10820 ( .INP(n10845), .Z(n10775) );
  NBUFFX2 U10821 ( .INP(n10845), .Z(n10776) );
  NBUFFX2 U10822 ( .INP(n10845), .Z(n10777) );
  NBUFFX2 U10823 ( .INP(n10844), .Z(n10778) );
  NBUFFX2 U10824 ( .INP(n10844), .Z(n10779) );
  NBUFFX2 U10825 ( .INP(n10844), .Z(n10780) );
  NBUFFX2 U10826 ( .INP(n10843), .Z(n10781) );
  NBUFFX2 U10827 ( .INP(n10843), .Z(n10782) );
  NBUFFX2 U10828 ( .INP(n10843), .Z(n10783) );
  NBUFFX2 U10829 ( .INP(n10842), .Z(n10784) );
  NBUFFX2 U10830 ( .INP(n10842), .Z(n10785) );
  NBUFFX2 U10831 ( .INP(n10842), .Z(n10786) );
  NBUFFX2 U10832 ( .INP(n10841), .Z(n10787) );
  NBUFFX2 U10833 ( .INP(n10841), .Z(n10788) );
  NBUFFX2 U10834 ( .INP(n10841), .Z(n10789) );
  NBUFFX2 U10835 ( .INP(n10840), .Z(n10790) );
  NBUFFX2 U10836 ( .INP(n10840), .Z(n10791) );
  NBUFFX2 U10837 ( .INP(n10840), .Z(n10792) );
  NBUFFX2 U10838 ( .INP(n10839), .Z(n10793) );
  NBUFFX2 U10839 ( .INP(n10839), .Z(n10794) );
  NBUFFX2 U10840 ( .INP(n10839), .Z(n10795) );
  NBUFFX2 U10841 ( .INP(n10838), .Z(n10796) );
  NBUFFX2 U10842 ( .INP(n10838), .Z(n10797) );
  NBUFFX2 U10843 ( .INP(n10838), .Z(n10798) );
  NBUFFX2 U10844 ( .INP(n10837), .Z(n10799) );
  NBUFFX2 U10845 ( .INP(n10837), .Z(n10800) );
  NBUFFX2 U10846 ( .INP(n10837), .Z(n10801) );
  NBUFFX2 U10847 ( .INP(n10836), .Z(n10802) );
  NBUFFX2 U10848 ( .INP(n10836), .Z(n10803) );
  NBUFFX2 U10849 ( .INP(n10836), .Z(n10804) );
  NBUFFX2 U10850 ( .INP(n10835), .Z(n10805) );
  NBUFFX2 U10851 ( .INP(n10835), .Z(n10806) );
  NBUFFX2 U10852 ( .INP(n10835), .Z(n10807) );
  NBUFFX2 U10853 ( .INP(n10834), .Z(n10808) );
  NBUFFX2 U10854 ( .INP(n10834), .Z(n10809) );
  NBUFFX2 U10855 ( .INP(n10834), .Z(n10810) );
  NBUFFX2 U10856 ( .INP(n10833), .Z(n10811) );
  NBUFFX2 U10857 ( .INP(n10833), .Z(n10812) );
  NBUFFX2 U10858 ( .INP(n10833), .Z(n10813) );
  NBUFFX2 U10859 ( .INP(n10832), .Z(n10814) );
  NBUFFX2 U10860 ( .INP(n10832), .Z(n10815) );
  NBUFFX2 U10861 ( .INP(n10832), .Z(n10816) );
  NBUFFX2 U10862 ( .INP(n10831), .Z(n10817) );
  NBUFFX2 U10863 ( .INP(n10831), .Z(n10818) );
  NBUFFX2 U10864 ( .INP(n10831), .Z(n10819) );
  NBUFFX2 U10865 ( .INP(n10830), .Z(n10820) );
  NBUFFX2 U10866 ( .INP(n10830), .Z(n10821) );
  NBUFFX2 U10867 ( .INP(n10830), .Z(n10822) );
  NBUFFX2 U10868 ( .INP(n10829), .Z(n10823) );
  NBUFFX2 U10869 ( .INP(n10829), .Z(n10824) );
  NBUFFX2 U10870 ( .INP(n10829), .Z(n10825) );
  NBUFFX2 U10871 ( .INP(n10828), .Z(n10826) );
  NBUFFX2 U10872 ( .INP(n10828), .Z(n10827) );
  NBUFFX2 U10873 ( .INP(n10869), .Z(n10828) );
  NBUFFX2 U10874 ( .INP(n10868), .Z(n10829) );
  NBUFFX2 U10875 ( .INP(n10868), .Z(n10830) );
  NBUFFX2 U10876 ( .INP(n10868), .Z(n10831) );
  NBUFFX2 U10877 ( .INP(n10867), .Z(n10832) );
  NBUFFX2 U10878 ( .INP(n10867), .Z(n10833) );
  NBUFFX2 U10879 ( .INP(n10867), .Z(n10834) );
  NBUFFX2 U10880 ( .INP(n10866), .Z(n10835) );
  NBUFFX2 U10881 ( .INP(n10866), .Z(n10836) );
  NBUFFX2 U10882 ( .INP(n10866), .Z(n10837) );
  NBUFFX2 U10883 ( .INP(n10865), .Z(n10838) );
  NBUFFX2 U10884 ( .INP(n10865), .Z(n10839) );
  NBUFFX2 U10885 ( .INP(n10865), .Z(n10840) );
  NBUFFX2 U10886 ( .INP(n10864), .Z(n10841) );
  NBUFFX2 U10887 ( .INP(n10864), .Z(n10842) );
  NBUFFX2 U10888 ( .INP(n10864), .Z(n10843) );
  NBUFFX2 U10889 ( .INP(n10863), .Z(n10844) );
  NBUFFX2 U10890 ( .INP(n10863), .Z(n10845) );
  NBUFFX2 U10891 ( .INP(n10863), .Z(n10846) );
  NBUFFX2 U10892 ( .INP(n10862), .Z(n10847) );
  NBUFFX2 U10893 ( .INP(n10862), .Z(n10848) );
  NBUFFX2 U10894 ( .INP(n10862), .Z(n10849) );
  NBUFFX2 U10895 ( .INP(n10861), .Z(n10850) );
  NBUFFX2 U10896 ( .INP(n10861), .Z(n10851) );
  NBUFFX2 U10897 ( .INP(n10861), .Z(n10852) );
  NBUFFX2 U10898 ( .INP(n10860), .Z(n10853) );
  NBUFFX2 U10899 ( .INP(n10860), .Z(n10854) );
  NBUFFX2 U10900 ( .INP(n10860), .Z(n10855) );
  NBUFFX2 U10901 ( .INP(n10859), .Z(n10856) );
  NBUFFX2 U10902 ( .INP(n10859), .Z(n10857) );
  NBUFFX2 U10903 ( .INP(n10859), .Z(n10858) );
  NBUFFX2 U10904 ( .INP(n10873), .Z(n10859) );
  NBUFFX2 U10905 ( .INP(n10873), .Z(n10860) );
  NBUFFX2 U10906 ( .INP(n10872), .Z(n10861) );
  NBUFFX2 U10907 ( .INP(n10872), .Z(n10862) );
  NBUFFX2 U10908 ( .INP(n10872), .Z(n10863) );
  NBUFFX2 U10909 ( .INP(n10871), .Z(n10864) );
  NBUFFX2 U10910 ( .INP(n10871), .Z(n10865) );
  NBUFFX2 U10911 ( .INP(n10871), .Z(n10866) );
  NBUFFX2 U10912 ( .INP(n10870), .Z(n10867) );
  NBUFFX2 U10913 ( .INP(n10870), .Z(n10868) );
  NBUFFX2 U10914 ( .INP(n10870), .Z(n10869) );
  NBUFFX2 U10915 ( .INP(g35), .Z(n10870) );
  NBUFFX2 U10916 ( .INP(g35), .Z(n10871) );
  NBUFFX2 U10917 ( .INP(g35), .Z(n10872) );
  NBUFFX2 U10918 ( .INP(g35), .Z(n10873) );
  INVX0 U10919 ( .INP(n10740), .ZN(n10874) );
  INVX0 U10920 ( .INP(n10740), .ZN(n10875) );
  INVX0 U10921 ( .INP(n10740), .ZN(n10876) );
  INVX0 U10922 ( .INP(n10741), .ZN(n10877) );
  INVX0 U10923 ( .INP(n10741), .ZN(n10878) );
  INVX0 U10924 ( .INP(n10741), .ZN(n10879) );
  INVX0 U10925 ( .INP(n10741), .ZN(n10880) );
  INVX0 U10926 ( .INP(n10741), .ZN(n10881) );
  INVX0 U10927 ( .INP(n10741), .ZN(n10882) );
  INVX0 U10928 ( .INP(n10741), .ZN(n10883) );
  INVX0 U10929 ( .INP(n10741), .ZN(n10884) );
  INVX0 U10930 ( .INP(n10741), .ZN(n10885) );
  INVX0 U10931 ( .INP(n10742), .ZN(n10886) );
  INVX0 U10932 ( .INP(n10742), .ZN(n10887) );
  INVX0 U10933 ( .INP(n10742), .ZN(n10888) );
  INVX0 U10934 ( .INP(n10742), .ZN(n10889) );
  INVX0 U10935 ( .INP(n10742), .ZN(n10890) );
  INVX0 U10936 ( .INP(n10742), .ZN(n10891) );
  INVX0 U10937 ( .INP(n10742), .ZN(n10892) );
  INVX0 U10938 ( .INP(n10742), .ZN(n10893) );
  INVX0 U10939 ( .INP(n10743), .ZN(n10894) );
  INVX0 U10940 ( .INP(n10743), .ZN(n10895) );
  INVX0 U10941 ( .INP(n10743), .ZN(n10896) );
  INVX0 U10942 ( .INP(n10742), .ZN(n10897) );
  INVX0 U10943 ( .INP(n10743), .ZN(n10898) );
  INVX0 U10944 ( .INP(n10743), .ZN(n10899) );
  INVX0 U10945 ( .INP(n10743), .ZN(n10900) );
  INVX0 U10946 ( .INP(n10743), .ZN(n10901) );
  INVX0 U10947 ( .INP(n10743), .ZN(n10902) );
  INVX0 U10948 ( .INP(n10743), .ZN(n10903) );
  INVX0 U10949 ( .INP(n10744), .ZN(n10904) );
  INVX0 U10950 ( .INP(n10744), .ZN(n10905) );
  INVX0 U10951 ( .INP(n10744), .ZN(n10906) );
  INVX0 U10952 ( .INP(n10744), .ZN(n10907) );
  INVX0 U10953 ( .INP(n10744), .ZN(n10908) );
  INVX0 U10954 ( .INP(n10744), .ZN(n10909) );
  INVX0 U10955 ( .INP(n10744), .ZN(n10910) );
  INVX0 U10956 ( .INP(n10744), .ZN(n10911) );
  INVX0 U10957 ( .INP(n10744), .ZN(n10912) );
  INVX0 U10958 ( .INP(n10745), .ZN(n10913) );
  INVX0 U10959 ( .INP(n10746), .ZN(n10914) );
  INVX0 U10960 ( .INP(n10745), .ZN(n10915) );
  INVX0 U10961 ( .INP(n10745), .ZN(n10916) );
  INVX0 U10962 ( .INP(n10745), .ZN(n10917) );
  INVX0 U10963 ( .INP(n10746), .ZN(n10918) );
  INVX0 U10964 ( .INP(n10746), .ZN(n10919) );
  INVX0 U10965 ( .INP(n10747), .ZN(n10920) );
  INVX0 U10966 ( .INP(n10746), .ZN(n10921) );
  INVX0 U10967 ( .INP(n10746), .ZN(n10922) );
  INVX0 U10968 ( .INP(n10745), .ZN(n10923) );
  INVX0 U10969 ( .INP(n10745), .ZN(n10924) );
  INVX0 U10970 ( .INP(n10746), .ZN(n10925) );
  INVX0 U10971 ( .INP(n10746), .ZN(n10926) );
  INVX0 U10972 ( .INP(n10746), .ZN(n10927) );
  INVX0 U10973 ( .INP(n10745), .ZN(n10928) );
  INVX0 U10974 ( .INP(n10746), .ZN(n10929) );
  INVX0 U10975 ( .INP(n10745), .ZN(n10930) );
  INVX0 U10976 ( .INP(n10745), .ZN(n10931) );
  INVX0 U10977 ( .INP(n10740), .ZN(n10932) );
  NBUFFX2 U10978 ( .INP(n11069), .Z(n11040) );
  NBUFFX2 U10979 ( .INP(n11068), .Z(n11041) );
  NBUFFX2 U10980 ( .INP(n11068), .Z(n11042) );
  NBUFFX2 U10981 ( .INP(n11068), .Z(n11043) );
  NBUFFX2 U10982 ( .INP(n11067), .Z(n11044) );
  NBUFFX2 U10983 ( .INP(n11067), .Z(n11045) );
  NBUFFX2 U10984 ( .INP(n11067), .Z(n11046) );
  NBUFFX2 U10985 ( .INP(n11066), .Z(n11047) );
  NBUFFX2 U10986 ( .INP(n11066), .Z(n11048) );
  NBUFFX2 U10987 ( .INP(n11066), .Z(n11049) );
  NBUFFX2 U10988 ( .INP(n11065), .Z(n11050) );
  NBUFFX2 U10989 ( .INP(n11065), .Z(n11051) );
  NBUFFX2 U10990 ( .INP(n11065), .Z(n11052) );
  NBUFFX2 U10991 ( .INP(n11064), .Z(n11053) );
  NBUFFX2 U10992 ( .INP(n11064), .Z(n11054) );
  NBUFFX2 U10993 ( .INP(n11064), .Z(n11055) );
  NBUFFX2 U10994 ( .INP(n11063), .Z(n11056) );
  NBUFFX2 U10995 ( .INP(n11063), .Z(n11057) );
  NBUFFX2 U10996 ( .INP(n11063), .Z(n11058) );
  NBUFFX2 U10997 ( .INP(n11062), .Z(n11059) );
  NBUFFX2 U10998 ( .INP(n11062), .Z(n11060) );
  NBUFFX2 U10999 ( .INP(n11062), .Z(n11061) );
  NBUFFX2 U11000 ( .INP(n11072), .Z(n11062) );
  NBUFFX2 U11001 ( .INP(n11072), .Z(n11063) );
  NBUFFX2 U11002 ( .INP(n11071), .Z(n11064) );
  NBUFFX2 U11003 ( .INP(n11071), .Z(n11065) );
  NBUFFX2 U11004 ( .INP(n11071), .Z(n11066) );
  NBUFFX2 U11005 ( .INP(n11070), .Z(n11067) );
  NBUFFX2 U11006 ( .INP(n11070), .Z(n11068) );
  NBUFFX2 U11007 ( .INP(n11070), .Z(n11069) );
  NBUFFX2 U11008 ( .INP(CK), .Z(n11070) );
  NBUFFX2 U11009 ( .INP(CK), .Z(n11071) );
  NBUFFX2 U11010 ( .INP(CK), .Z(n11072) );
  INVX0 U11011 ( .INP(n11073), .ZN(n879) );
  INVX0 U11012 ( .INP(n11074), .ZN(n760) );
  INVX0 U11013 ( .INP(n11075), .ZN(n736) );
  INVX0 U11014 ( .INP(n11076), .ZN(n727) );
  INVX0 U11015 ( .INP(n11077), .ZN(n725) );
  OR2X1 U11016 ( .IN1(n11078), .IN2(n11079), .Q(n5961) );
  OR2X1 U11017 ( .IN1(n11080), .IN2(n11081), .Q(n11079) );
  AND2X1 U11018 ( .IN1(n10381), .IN2(n11082), .Q(n11081) );
  AND2X1 U11019 ( .IN1(n11083), .IN2(g5348), .Q(n11080) );
  OR2X1 U11020 ( .IN1(n11084), .IN2(n11085), .Q(n11078) );
  AND2X1 U11021 ( .IN1(n10514), .IN2(n11086), .Q(n11085) );
  AND2X1 U11022 ( .IN1(g31860), .IN2(g5352), .Q(n11084) );
  OR2X1 U11023 ( .IN1(n11087), .IN2(n11088), .Q(n5960) );
  OR2X1 U11024 ( .IN1(n11089), .IN2(n11090), .Q(n11088) );
  AND2X1 U11025 ( .IN1(n10380), .IN2(n11091), .Q(n11090) );
  AND2X1 U11026 ( .IN1(n11092), .IN2(g6732), .Q(n11089) );
  OR2X1 U11027 ( .IN1(n11093), .IN2(n11094), .Q(n11087) );
  AND2X1 U11028 ( .IN1(n10495), .IN2(n11095), .Q(n11094) );
  AND2X1 U11029 ( .IN1(n11096), .IN2(g6736), .Q(n11093) );
  INVX0 U11030 ( .INP(n11097), .ZN(n516) );
  INVX0 U11031 ( .INP(n11098), .ZN(n515) );
  INVX0 U11032 ( .INP(n11099), .ZN(n4722) );
  OR2X1 U11033 ( .IN1(n10197), .IN2(n11100), .Q(n4459) );
  OR2X1 U11034 ( .IN1(n10193), .IN2(n11101), .Q(n4448) );
  OR2X1 U11035 ( .IN1(n11102), .IN2(n10572), .Q(n4437) );
  OR2X1 U11036 ( .IN1(n10198), .IN2(n11103), .Q(n4426) );
  OR2X1 U11037 ( .IN1(n10191), .IN2(n11104), .Q(n4415) );
  OR2X1 U11038 ( .IN1(n10195), .IN2(n11105), .Q(n4403) );
  OR2X1 U11039 ( .IN1(n10302), .IN2(n11106), .Q(n4392) );
  OR2X1 U11040 ( .IN1(n10201), .IN2(n11107), .Q(n4380) );
  OR2X1 U11041 ( .IN1(n11108), .IN2(n11109), .Q(n4305) );
  OR2X1 U11042 ( .IN1(n11110), .IN2(n11111), .Q(n11109) );
  OR2X1 U11043 ( .IN1(n11112), .IN2(n11113), .Q(n11111) );
  AND2X1 U11044 ( .IN1(n11114), .IN2(n5656), .Q(n11113) );
  AND2X1 U11045 ( .IN1(n11115), .IN2(n11116), .Q(n11114) );
  OR2X1 U11046 ( .IN1(n11117), .IN2(n11118), .Q(n11116) );
  AND2X1 U11047 ( .IN1(n11119), .IN2(n11120), .Q(n11117) );
  OR2X1 U11048 ( .IN1(n11121), .IN2(n5707), .Q(n11120) );
  AND2X1 U11049 ( .IN1(n5368), .IN2(n11122), .Q(n11121) );
  XOR2X1 U11050 ( .IN1(g34657), .IN2(n11123), .Q(n11122) );
  OR2X1 U11051 ( .IN1(n11124), .IN2(n11125), .Q(n11123) );
  OR2X1 U11052 ( .IN1(n11126), .IN2(n11127), .Q(n11125) );
  AND2X1 U11053 ( .IN1(n11128), .IN2(g4727), .Q(n11127) );
  AND2X1 U11054 ( .IN1(n11129), .IN2(g4722), .Q(n11126) );
  OR2X1 U11055 ( .IN1(n11130), .IN2(n11131), .Q(n11124) );
  AND2X1 U11056 ( .IN1(n11132), .IN2(g4717), .Q(n11131) );
  AND2X1 U11057 ( .IN1(n11133), .IN2(g4732), .Q(n11130) );
  AND2X1 U11058 ( .IN1(n11134), .IN2(n11135), .Q(n11119) );
  OR2X1 U11059 ( .IN1(n11136), .IN2(g4793), .Q(n11135) );
  AND2X1 U11060 ( .IN1(n11137), .IN2(n10561), .Q(n11136) );
  OR2X1 U11061 ( .IN1(n11138), .IN2(n11139), .Q(n11137) );
  OR2X1 U11062 ( .IN1(n11140), .IN2(g4776), .Q(n11139) );
  AND2X1 U11063 ( .IN1(n5867), .IN2(n11128), .Q(n11140) );
  OR2X1 U11064 ( .IN1(n11132), .IN2(n11133), .Q(n11138) );
  OR2X1 U11065 ( .IN1(n5368), .IN2(g34657), .Q(n11134) );
  AND2X1 U11066 ( .IN1(n10074), .IN2(g4688), .Q(n11112) );
  AND2X1 U11067 ( .IN1(n5880), .IN2(g4674), .Q(n11110) );
  OR2X1 U11068 ( .IN1(n11141), .IN2(n11142), .Q(n11108) );
  INVX0 U11069 ( .INP(n11143), .ZN(n11142) );
  OR2X1 U11070 ( .IN1(n10076), .IN2(n10435), .Q(n11143) );
  AND2X1 U11071 ( .IN1(g29220), .IN2(g4646), .Q(n11141) );
  OR2X1 U11072 ( .IN1(n11144), .IN2(n11145), .Q(n4283) );
  OR2X1 U11073 ( .IN1(n11146), .IN2(n11147), .Q(n11145) );
  OR2X1 U11074 ( .IN1(n11148), .IN2(n11149), .Q(n11147) );
  AND2X1 U11075 ( .IN1(n11150), .IN2(n5283), .Q(n11149) );
  AND2X1 U11076 ( .IN1(n11151), .IN2(n11152), .Q(n11150) );
  OR2X1 U11077 ( .IN1(n11153), .IN2(n11154), .Q(n11152) );
  AND2X1 U11078 ( .IN1(n11155), .IN2(n11156), .Q(n11153) );
  OR2X1 U11079 ( .IN1(n11157), .IN2(n5706), .Q(n11156) );
  AND2X1 U11080 ( .IN1(n5367), .IN2(n11158), .Q(n11157) );
  XOR2X1 U11081 ( .IN1(g34649), .IN2(n11159), .Q(n11158) );
  OR2X1 U11082 ( .IN1(n11160), .IN2(n11161), .Q(n11159) );
  OR2X1 U11083 ( .IN1(n11162), .IN2(n11163), .Q(n11161) );
  AND2X1 U11084 ( .IN1(n11164), .IN2(g4907), .Q(n11163) );
  AND2X1 U11085 ( .IN1(n11165), .IN2(g4922), .Q(n11162) );
  OR2X1 U11086 ( .IN1(n11166), .IN2(n11167), .Q(n11160) );
  AND2X1 U11087 ( .IN1(n11168), .IN2(g4917), .Q(n11167) );
  AND2X1 U11088 ( .IN1(n11169), .IN2(g4912), .Q(n11166) );
  AND2X1 U11089 ( .IN1(n11170), .IN2(n11171), .Q(n11155) );
  OR2X1 U11090 ( .IN1(n11172), .IN2(g4983), .Q(n11171) );
  AND2X1 U11091 ( .IN1(n11173), .IN2(n10560), .Q(n11172) );
  OR2X1 U11092 ( .IN1(n11174), .IN2(n11175), .Q(n11173) );
  OR2X1 U11093 ( .IN1(n11176), .IN2(g4966), .Q(n11175) );
  AND2X1 U11094 ( .IN1(n5879), .IN2(n11168), .Q(n11176) );
  OR2X1 U11095 ( .IN1(n11164), .IN2(n11165), .Q(n11174) );
  OR2X1 U11096 ( .IN1(n5367), .IN2(g34649), .Q(n11170) );
  AND2X1 U11097 ( .IN1(n10078), .IN2(g4878), .Q(n11148) );
  AND2X1 U11098 ( .IN1(g4871), .IN2(g3684), .Q(n11146) );
  OR2X1 U11099 ( .IN1(n11177), .IN2(n11178), .Q(n11144) );
  AND2X1 U11100 ( .IN1(g5011), .IN2(g4836), .Q(n11178) );
  AND2X1 U11101 ( .IN1(n10077), .IN2(g4864), .Q(n11177) );
  AND2X1 U11102 ( .IN1(n11179), .IN2(n5652), .Q(n4034) );
  AND2X1 U11103 ( .IN1(n5366), .IN2(n10425), .Q(n11179) );
  AND2X1 U11104 ( .IN1(n11180), .IN2(n5645), .Q(n4002) );
  AND2X1 U11105 ( .IN1(n5576), .IN2(n10427), .Q(n11180) );
  AND2X1 U11106 ( .IN1(n11181), .IN2(n5572), .Q(n3969) );
  AND2X1 U11107 ( .IN1(n10432), .IN2(n10553), .Q(n11181) );
  AND2X1 U11108 ( .IN1(n11182), .IN2(n11183), .Q(n3933) );
  AND2X1 U11109 ( .IN1(n2760), .IN2(g43), .Q(n11183) );
  AND2X1 U11110 ( .IN1(n11184), .IN2(n5650), .Q(n3926) );
  AND2X1 U11111 ( .IN1(n5570), .IN2(n10429), .Q(n11184) );
  AND2X1 U11112 ( .IN1(n11185), .IN2(n5647), .Q(n3893) );
  AND2X1 U11113 ( .IN1(n5575), .IN2(n10426), .Q(n11185) );
  AND2X1 U11114 ( .IN1(n11186), .IN2(n5649), .Q(n3860) );
  AND2X1 U11115 ( .IN1(n5573), .IN2(n10430), .Q(n11186) );
  AND2X1 U11116 ( .IN1(n11187), .IN2(n5651), .Q(n3826) );
  AND2X1 U11117 ( .IN1(n5574), .IN2(n10428), .Q(n11187) );
  AND2X1 U11118 ( .IN1(n11188), .IN2(n5646), .Q(n3792) );
  AND2X1 U11119 ( .IN1(n5571), .IN2(n10431), .Q(n11188) );
  OR2X1 U11120 ( .IN1(n11189), .IN2(n11190), .Q(n3675) );
  OR2X1 U11121 ( .IN1(g691), .IN2(g417), .Q(n11190) );
  OR2X1 U11122 ( .IN1(n11191), .IN2(n11192), .Q(n11189) );
  AND2X1 U11123 ( .IN1(n11193), .IN2(g392), .Q(n11192) );
  OR2X1 U11124 ( .IN1(g441), .IN2(n11194), .Q(n11193) );
  XOR2X1 U11125 ( .IN1(test_so72), .IN2(n10275), .Q(n11194) );
  AND2X1 U11126 ( .IN1(n10465), .IN2(n11195), .Q(n11191) );
  OR2X1 U11127 ( .IN1(g411), .IN2(n11196), .Q(n11195) );
  XNOR2X1 U11128 ( .IN1(test_so72), .IN2(g174), .Q(n11196) );
  OR2X1 U11129 ( .IN1(n5349), .IN2(n11197), .Q(n3635) );
  INVX0 U11130 ( .INP(n11198), .ZN(n346) );
  AND2X1 U11131 ( .IN1(n3064), .IN2(n11199), .Q(n11198) );
  OR2X1 U11132 ( .IN1(n5715), .IN2(n11200), .Q(n11199) );
  AND2X1 U11133 ( .IN1(n11201), .IN2(n10771), .Q(n11200) );
  OR2X1 U11134 ( .IN1(g4104), .IN2(n11202), .Q(n11201) );
  AND2X1 U11135 ( .IN1(n11203), .IN2(n11204), .Q(n3174) );
  XNOR2X1 U11136 ( .IN1(g490), .IN2(g73), .Q(n11204) );
  XNOR2X1 U11137 ( .IN1(n11205), .IN2(n5820), .Q(n11203) );
  AND2X1 U11138 ( .IN1(n2760), .IN2(n9302), .Q(n3084) );
  OR2X1 U11139 ( .IN1(n11206), .IN2(n11207), .Q(n3065) );
  OR2X1 U11140 ( .IN1(n10274), .IN2(n10875), .Q(n11207) );
  AND2X1 U11141 ( .IN1(n11208), .IN2(g4108), .Q(n11206) );
  INVX0 U11142 ( .INP(n11209), .ZN(n290) );
  INVX0 U11143 ( .INP(n11210), .ZN(n286) );
  XNOR2X1 U11144 ( .IN1(g4311), .IN2(n2607), .Q(n2608) );
  INVX0 U11145 ( .INP(n11211), .ZN(n2461) );
  AND2X1 U11146 ( .IN1(g34979), .IN2(n11212), .Q(n11211) );
  AND2X1 U11147 ( .IN1(n11212), .IN2(g34971), .Q(n2396) );
  INVX0 U11148 ( .INP(n11213), .ZN(n174) );
  INVX0 U11149 ( .INP(n11214), .ZN(n173) );
  INVX0 U11150 ( .INP(n11215), .ZN(n1643) );
  INVX0 U11151 ( .INP(n11216), .ZN(n1289) );
  INVX0 U11152 ( .INP(n11217), .ZN(n1287) );
  INVX0 U11153 ( .INP(n11218), .ZN(n1285) );
  INVX0 U11154 ( .INP(n11219), .ZN(n1282) );
  INVX0 U11155 ( .INP(n11220), .ZN(n1156) );
  AND2X1 U11156 ( .IN1(n11182), .IN2(n11221), .Q(n10533) );
  OR2X1 U11157 ( .IN1(n11222), .IN2(n11223), .Q(g34980) );
  AND2X1 U11158 ( .IN1(n11224), .IN2(n10763), .Q(n11223) );
  OR2X1 U11159 ( .IN1(n11225), .IN2(g2984), .Q(n11224) );
  AND2X1 U11160 ( .IN1(n11226), .IN2(n11227), .Q(n11225) );
  INVX0 U11161 ( .INP(n11228), .ZN(n11227) );
  OR2X1 U11162 ( .IN1(g54), .IN2(g56), .Q(n11228) );
  AND2X1 U11163 ( .IN1(n10532), .IN2(n11229), .Q(n11226) );
  AND2X1 U11164 ( .IN1(test_so14), .IN2(n10895), .Q(n11222) );
  OR2X1 U11165 ( .IN1(n10527), .IN2(n10532), .Q(g34972) );
  XOR2X1 U11166 ( .IN1(n11230), .IN2(n11231), .Q(n10532) );
  XOR2X1 U11167 ( .IN1(n11232), .IN2(n11233), .Q(n11231) );
  XOR2X1 U11168 ( .IN1(n11234), .IN2(n11235), .Q(n11233) );
  XOR2X1 U11169 ( .IN1(g34978), .IN2(g34977), .Q(n11235) );
  XOR2X1 U11170 ( .IN1(g34976), .IN2(g34975), .Q(n11234) );
  XOR2X1 U11171 ( .IN1(n11236), .IN2(n11237), .Q(n11232) );
  XOR2X1 U11172 ( .IN1(g34974), .IN2(g34970), .Q(n11237) );
  XOR2X1 U11173 ( .IN1(g34979), .IN2(g34971), .Q(n11236) );
  OR2X1 U11174 ( .IN1(n11238), .IN2(n10008), .Q(n11230) );
  OR2X1 U11175 ( .IN1(n10527), .IN2(g34979), .Q(g34927) );
  OR2X1 U11176 ( .IN1(n11239), .IN2(n11240), .Q(g34979) );
  OR2X1 U11177 ( .IN1(n11241), .IN2(n11242), .Q(n11240) );
  OR2X1 U11178 ( .IN1(n11243), .IN2(n11244), .Q(n11242) );
  AND2X1 U11179 ( .IN1(n11245), .IN2(g1283), .Q(n11244) );
  AND2X1 U11180 ( .IN1(n11246), .IN2(g939), .Q(n11243) );
  OR2X1 U11181 ( .IN1(n11247), .IN2(n11248), .Q(n11241) );
  AND2X1 U11182 ( .IN1(n11249), .IN2(g2697), .Q(n11248) );
  AND2X1 U11183 ( .IN1(n11250), .IN2(n9332), .Q(n11247) );
  OR2X1 U11184 ( .IN1(n11251), .IN2(n11252), .Q(n11239) );
  OR2X1 U11185 ( .IN1(n11253), .IN2(n11254), .Q(n11252) );
  AND2X1 U11186 ( .IN1(n11255), .IN2(g2138), .Q(n11254) );
  AND2X1 U11187 ( .IN1(n1340), .IN2(n11256), .Q(n11253) );
  OR2X1 U11188 ( .IN1(n11257), .IN2(n11258), .Q(n11256) );
  OR2X1 U11189 ( .IN1(n11259), .IN2(n11260), .Q(n11258) );
  OR2X1 U11190 ( .IN1(n11261), .IN2(n11262), .Q(n11260) );
  OR2X1 U11191 ( .IN1(n11263), .IN2(n11264), .Q(n11262) );
  AND2X1 U11192 ( .IN1(n11265), .IN2(g604), .Q(n11264) );
  AND2X1 U11193 ( .IN1(n11266), .IN2(g744), .Q(n11263) );
  AND2X1 U11194 ( .IN1(n11267), .IN2(g568), .Q(n11261) );
  OR2X1 U11195 ( .IN1(n11268), .IN2(n11269), .Q(n11259) );
  OR2X1 U11196 ( .IN1(n11270), .IN2(n11271), .Q(n11269) );
  AND2X1 U11197 ( .IN1(n11272), .IN2(g2975), .Q(n11271) );
  AND2X1 U11198 ( .IN1(n11273), .IN2(g4146), .Q(n11270) );
  AND2X1 U11199 ( .IN1(g29221), .IN2(n11274), .Q(n11268) );
  OR2X1 U11200 ( .IN1(n11275), .IN2(n11276), .Q(n11257) );
  OR2X1 U11201 ( .IN1(n11277), .IN2(n11278), .Q(n11276) );
  OR2X1 U11202 ( .IN1(n11279), .IN2(n11280), .Q(n11278) );
  AND2X1 U11203 ( .IN1(n11281), .IN2(g2886), .Q(n11280) );
  AND2X1 U11204 ( .IN1(n11282), .IN2(g785), .Q(n11279) );
  AND2X1 U11205 ( .IN1(n11283), .IN2(g2970), .Q(n11277) );
  OR2X1 U11206 ( .IN1(n11284), .IN2(n11285), .Q(n11275) );
  OR2X1 U11207 ( .IN1(n11286), .IN2(n11287), .Q(n11285) );
  AND2X1 U11208 ( .IN1(g92), .IN2(n11288), .Q(n11287) );
  AND2X1 U11209 ( .IN1(g127), .IN2(n11289), .Q(n11286) );
  AND2X1 U11210 ( .IN1(test_so14), .IN2(n11212), .Q(n11284) );
  OR2X1 U11211 ( .IN1(n11290), .IN2(n11291), .Q(n11251) );
  AND2X1 U11212 ( .IN1(test_so67), .IN2(n11292), .Q(n11291) );
  OR2X1 U11213 ( .IN1(n10527), .IN2(g34978), .Q(g34925) );
  OR2X1 U11214 ( .IN1(n11293), .IN2(n11294), .Q(g34978) );
  OR2X1 U11215 ( .IN1(n11295), .IN2(n11296), .Q(n11294) );
  OR2X1 U11216 ( .IN1(n11297), .IN2(n11298), .Q(n11296) );
  AND2X1 U11217 ( .IN1(n10010), .IN2(n11245), .Q(n11298) );
  AND2X1 U11218 ( .IN1(n10011), .IN2(n11246), .Q(n11297) );
  OR2X1 U11219 ( .IN1(n11299), .IN2(n11300), .Q(n11295) );
  AND2X1 U11220 ( .IN1(n11249), .IN2(g2689), .Q(n11300) );
  AND2X1 U11221 ( .IN1(n11250), .IN2(n9276), .Q(n11299) );
  OR2X1 U11222 ( .IN1(n11301), .IN2(n11302), .Q(n11293) );
  OR2X1 U11223 ( .IN1(n11303), .IN2(n11304), .Q(n11302) );
  AND2X1 U11224 ( .IN1(n11255), .IN2(g2130), .Q(n11304) );
  AND2X1 U11225 ( .IN1(n1340), .IN2(n11305), .Q(n11303) );
  OR2X1 U11226 ( .IN1(n11306), .IN2(n11307), .Q(n11305) );
  OR2X1 U11227 ( .IN1(n11308), .IN2(n11309), .Q(n11307) );
  OR2X1 U11228 ( .IN1(n11310), .IN2(n11311), .Q(n11309) );
  AND2X1 U11229 ( .IN1(n11267), .IN2(g572), .Q(n11311) );
  AND2X1 U11230 ( .IN1(n11265), .IN2(g608), .Q(n11310) );
  OR2X1 U11231 ( .IN1(n11312), .IN2(n11313), .Q(n11308) );
  OR2X1 U11232 ( .IN1(n11314), .IN2(n11315), .Q(n11313) );
  AND2X1 U11233 ( .IN1(n10413), .IN2(n11274), .Q(n11315) );
  AND2X1 U11234 ( .IN1(n11272), .IN2(g2965), .Q(n11314) );
  AND2X1 U11235 ( .IN1(test_so2), .IN2(n11266), .Q(n11312) );
  OR2X1 U11236 ( .IN1(n11316), .IN2(n11317), .Q(n11306) );
  OR2X1 U11237 ( .IN1(n11318), .IN2(n11319), .Q(n11317) );
  OR2X1 U11238 ( .IN1(n11320), .IN2(n11321), .Q(n11319) );
  AND2X1 U11239 ( .IN1(test_so22), .IN2(n11283), .Q(n11321) );
  AND2X1 U11240 ( .IN1(n11281), .IN2(g2878), .Q(n11320) );
  AND2X1 U11241 ( .IN1(n11273), .IN2(g4176), .Q(n11318) );
  OR2X1 U11242 ( .IN1(n11322), .IN2(n11323), .Q(n11316) );
  OR2X1 U11243 ( .IN1(n11324), .IN2(n11325), .Q(n11323) );
  AND2X1 U11244 ( .IN1(n11288), .IN2(g29214), .Q(n11325) );
  AND2X1 U11245 ( .IN1(n11289), .IN2(g2873), .Q(n11324) );
  AND2X1 U11246 ( .IN1(n11282), .IN2(g790), .Q(n11322) );
  OR2X1 U11247 ( .IN1(n11290), .IN2(n11326), .Q(n11301) );
  AND2X1 U11248 ( .IN1(n11292), .IN2(g4253), .Q(n11326) );
  OR2X1 U11249 ( .IN1(n10527), .IN2(g34977), .Q(g34923) );
  OR2X1 U11250 ( .IN1(n11327), .IN2(n11328), .Q(g34977) );
  OR2X1 U11251 ( .IN1(n11329), .IN2(n11330), .Q(n11328) );
  OR2X1 U11252 ( .IN1(n11331), .IN2(n11332), .Q(n11330) );
  AND2X1 U11253 ( .IN1(n11245), .IN2(g1291), .Q(n11332) );
  AND2X1 U11254 ( .IN1(n11246), .IN2(g947), .Q(n11331) );
  OR2X1 U11255 ( .IN1(n11333), .IN2(n11334), .Q(n11329) );
  AND2X1 U11256 ( .IN1(n11335), .IN2(n5879), .Q(n11334) );
  AND2X1 U11257 ( .IN1(n11336), .IN2(n5867), .Q(n11333) );
  OR2X1 U11258 ( .IN1(n11337), .IN2(n11338), .Q(n11327) );
  OR2X1 U11259 ( .IN1(n11339), .IN2(n11340), .Q(n11338) );
  AND2X1 U11260 ( .IN1(n11250), .IN2(n9245), .Q(n11340) );
  AND2X1 U11261 ( .IN1(n1340), .IN2(n11341), .Q(n11339) );
  OR2X1 U11262 ( .IN1(n11342), .IN2(n11343), .Q(n11341) );
  OR2X1 U11263 ( .IN1(n11344), .IN2(n11345), .Q(n11343) );
  OR2X1 U11264 ( .IN1(n11346), .IN2(n11347), .Q(n11345) );
  OR2X1 U11265 ( .IN1(n11348), .IN2(n11349), .Q(n11347) );
  AND2X1 U11266 ( .IN1(n11265), .IN2(g613), .Q(n11349) );
  AND2X1 U11267 ( .IN1(n11266), .IN2(g758), .Q(n11348) );
  AND2X1 U11268 ( .IN1(n11267), .IN2(g586), .Q(n11346) );
  OR2X1 U11269 ( .IN1(n11350), .IN2(n11351), .Q(n11344) );
  OR2X1 U11270 ( .IN1(n11352), .IN2(n11353), .Q(n11351) );
  AND2X1 U11271 ( .IN1(n11272), .IN2(g2955), .Q(n11353) );
  AND2X1 U11272 ( .IN1(n11273), .IN2(g4172), .Q(n11352) );
  AND2X1 U11273 ( .IN1(n11274), .IN2(g534), .Q(n11350) );
  OR2X1 U11274 ( .IN1(n11354), .IN2(n11355), .Q(n11342) );
  OR2X1 U11275 ( .IN1(n11356), .IN2(n11357), .Q(n11355) );
  OR2X1 U11276 ( .IN1(n11358), .IN2(n11359), .Q(n11357) );
  AND2X1 U11277 ( .IN1(n11281), .IN2(g2882), .Q(n11359) );
  AND2X1 U11278 ( .IN1(n11282), .IN2(g794), .Q(n11358) );
  AND2X1 U11279 ( .IN1(n11283), .IN2(g2950), .Q(n11356) );
  OR2X1 U11280 ( .IN1(n11360), .IN2(n11361), .Q(n11354) );
  OR2X1 U11281 ( .IN1(n11362), .IN2(n11363), .Q(n11361) );
  AND2X1 U11282 ( .IN1(n11289), .IN2(g2868), .Q(n11363) );
  AND2X1 U11283 ( .IN1(n11288), .IN2(g37), .Q(n11360) );
  OR2X1 U11284 ( .IN1(n11290), .IN2(n11364), .Q(n11337) );
  AND2X1 U11285 ( .IN1(n11292), .IN2(g4300), .Q(n11364) );
  OR2X1 U11286 ( .IN1(n10527), .IN2(g34976), .Q(g34921) );
  OR2X1 U11287 ( .IN1(n11365), .IN2(n11366), .Q(g34976) );
  OR2X1 U11288 ( .IN1(n11367), .IN2(n11368), .Q(n11366) );
  OR2X1 U11289 ( .IN1(n11369), .IN2(n11370), .Q(n11368) );
  AND2X1 U11290 ( .IN1(n11335), .IN2(g4912), .Q(n11370) );
  AND2X1 U11291 ( .IN1(n11336), .IN2(g4722), .Q(n11369) );
  OR2X1 U11292 ( .IN1(n11371), .IN2(n11372), .Q(n11367) );
  AND2X1 U11293 ( .IN1(n11249), .IN2(g6545), .Q(n11372) );
  AND2X1 U11294 ( .IN1(n11250), .IN2(n9357), .Q(n11371) );
  OR2X1 U11295 ( .IN1(n11373), .IN2(n11374), .Q(n11365) );
  OR2X1 U11296 ( .IN1(n11375), .IN2(n11376), .Q(n11374) );
  AND2X1 U11297 ( .IN1(n11255), .IN2(g5160), .Q(n11376) );
  AND2X1 U11298 ( .IN1(n1340), .IN2(n11377), .Q(n11375) );
  OR2X1 U11299 ( .IN1(n11378), .IN2(n11379), .Q(n11377) );
  OR2X1 U11300 ( .IN1(n11380), .IN2(n11381), .Q(n11379) );
  OR2X1 U11301 ( .IN1(n11382), .IN2(n11383), .Q(n11381) );
  AND2X1 U11302 ( .IN1(n11267), .IN2(g577), .Q(n11383) );
  AND2X1 U11303 ( .IN1(n11265), .IN2(g617), .Q(n11382) );
  OR2X1 U11304 ( .IN1(n11384), .IN2(n11385), .Q(n11380) );
  OR2X1 U11305 ( .IN1(n11386), .IN2(n11387), .Q(n11385) );
  AND2X1 U11306 ( .IN1(test_so41), .IN2(n11274), .Q(n11387) );
  AND2X1 U11307 ( .IN1(n11272), .IN2(g2941), .Q(n11386) );
  AND2X1 U11308 ( .IN1(n11266), .IN2(g763), .Q(n11384) );
  OR2X1 U11309 ( .IN1(n11388), .IN2(n11389), .Q(n11378) );
  OR2X1 U11310 ( .IN1(n11390), .IN2(n11391), .Q(n11389) );
  OR2X1 U11311 ( .IN1(n11392), .IN2(n11393), .Q(n11391) );
  AND2X1 U11312 ( .IN1(n11283), .IN2(g2936), .Q(n11393) );
  AND2X1 U11313 ( .IN1(n11281), .IN2(g2898), .Q(n11392) );
  AND2X1 U11314 ( .IN1(test_so95), .IN2(n11273), .Q(n11390) );
  OR2X1 U11315 ( .IN1(n11394), .IN2(n11395), .Q(n11388) );
  OR2X1 U11316 ( .IN1(n11362), .IN2(n11396), .Q(n11395) );
  AND2X1 U11317 ( .IN1(n11289), .IN2(g2988), .Q(n11396) );
  AND2X1 U11318 ( .IN1(n11282), .IN2(g807), .Q(n11394) );
  OR2X1 U11319 ( .IN1(n11397), .IN2(n11398), .Q(n11373) );
  OR2X1 U11320 ( .IN1(n11290), .IN2(n11399), .Q(n11398) );
  AND2X1 U11321 ( .IN1(n11400), .IN2(g1478), .Q(n11399) );
  AND2X1 U11322 ( .IN1(n11401), .IN2(g1135), .Q(n11397) );
  OR2X1 U11323 ( .IN1(n10527), .IN2(g34975), .Q(g34919) );
  OR2X1 U11324 ( .IN1(n11402), .IN2(n11403), .Q(g34975) );
  OR2X1 U11325 ( .IN1(n11404), .IN2(n11405), .Q(n11403) );
  OR2X1 U11326 ( .IN1(n11406), .IN2(n11407), .Q(n11405) );
  AND2X1 U11327 ( .IN1(n11335), .IN2(g4907), .Q(n11407) );
  AND2X1 U11328 ( .IN1(n11336), .IN2(g4717), .Q(n11406) );
  OR2X1 U11329 ( .IN1(n11408), .IN2(n11409), .Q(n11404) );
  AND2X1 U11330 ( .IN1(n11249), .IN2(g3151), .Q(n11409) );
  AND2X1 U11331 ( .IN1(n11250), .IN2(n9294), .Q(n11408) );
  OR2X1 U11332 ( .IN1(n11410), .IN2(n11411), .Q(n11402) );
  OR2X1 U11333 ( .IN1(n11412), .IN2(n11413), .Q(n11411) );
  AND2X1 U11334 ( .IN1(n11255), .IN2(g5507), .Q(n11413) );
  AND2X1 U11335 ( .IN1(n1340), .IN2(n11414), .Q(n11412) );
  OR2X1 U11336 ( .IN1(n11415), .IN2(n11416), .Q(n11414) );
  OR2X1 U11337 ( .IN1(n11417), .IN2(n11418), .Q(n11416) );
  OR2X1 U11338 ( .IN1(n11419), .IN2(n11420), .Q(n11418) );
  AND2X1 U11339 ( .IN1(n11267), .IN2(g582), .Q(n11420) );
  AND2X1 U11340 ( .IN1(n11265), .IN2(g622), .Q(n11419) );
  OR2X1 U11341 ( .IN1(n11421), .IN2(n11422), .Q(n11417) );
  OR2X1 U11342 ( .IN1(n11423), .IN2(n11424), .Q(n11422) );
  AND2X1 U11343 ( .IN1(n11274), .IN2(g546), .Q(n11424) );
  AND2X1 U11344 ( .IN1(n11272), .IN2(g2927), .Q(n11423) );
  AND2X1 U11345 ( .IN1(n11266), .IN2(g767), .Q(n11421) );
  OR2X1 U11346 ( .IN1(n11425), .IN2(n11426), .Q(n11415) );
  OR2X1 U11347 ( .IN1(n11427), .IN2(n11428), .Q(n11426) );
  AND2X1 U11348 ( .IN1(n11273), .IN2(g2860), .Q(n11428) );
  AND2X1 U11349 ( .IN1(n11283), .IN2(g2922), .Q(n11427) );
  OR2X1 U11350 ( .IN1(n11429), .IN2(n11430), .Q(n11425) );
  OR2X1 U11351 ( .IN1(n11431), .IN2(n11432), .Q(n11430) );
  AND2X1 U11352 ( .IN1(n11282), .IN2(g554), .Q(n11432) );
  AND2X1 U11353 ( .IN1(n5634), .IN2(n11289), .Q(n11431) );
  AND2X1 U11354 ( .IN1(n11281), .IN2(g2864), .Q(n11429) );
  OR2X1 U11355 ( .IN1(n11433), .IN2(n11434), .Q(n11410) );
  OR2X1 U11356 ( .IN1(n11290), .IN2(n11435), .Q(n11434) );
  AND2X1 U11357 ( .IN1(n11400), .IN2(g1448), .Q(n11435) );
  AND2X1 U11358 ( .IN1(n11401), .IN2(g1105), .Q(n11433) );
  OR2X1 U11359 ( .IN1(n10527), .IN2(g34974), .Q(g34917) );
  OR2X1 U11360 ( .IN1(n11436), .IN2(n11437), .Q(g34974) );
  OR2X1 U11361 ( .IN1(n11438), .IN2(n11439), .Q(n11437) );
  OR2X1 U11362 ( .IN1(n11440), .IN2(n11441), .Q(n11439) );
  AND2X1 U11363 ( .IN1(n11335), .IN2(g4922), .Q(n11441) );
  AND2X1 U11364 ( .IN1(n11336), .IN2(g4732), .Q(n11440) );
  OR2X1 U11365 ( .IN1(n11442), .IN2(n11443), .Q(n11438) );
  AND2X1 U11366 ( .IN1(test_so45), .IN2(n11249), .Q(n11443) );
  AND2X1 U11367 ( .IN1(n11250), .IN2(n9327), .Q(n11442) );
  OR2X1 U11368 ( .IN1(n11444), .IN2(n11445), .Q(n11436) );
  OR2X1 U11369 ( .IN1(n11446), .IN2(n11447), .Q(n11445) );
  AND2X1 U11370 ( .IN1(n11255), .IN2(g5853), .Q(n11447) );
  AND2X1 U11371 ( .IN1(n1340), .IN2(n11448), .Q(n11446) );
  OR2X1 U11372 ( .IN1(n11449), .IN2(n11450), .Q(n11448) );
  OR2X1 U11373 ( .IN1(n11451), .IN2(n11452), .Q(n11450) );
  OR2X1 U11374 ( .IN1(n11453), .IN2(n11454), .Q(n11452) );
  AND2X1 U11375 ( .IN1(n11267), .IN2(g590), .Q(n11454) );
  AND2X1 U11376 ( .IN1(n11265), .IN2(g626), .Q(n11453) );
  OR2X1 U11377 ( .IN1(n11455), .IN2(n11456), .Q(n11451) );
  AND2X1 U11378 ( .IN1(n11266), .IN2(g772), .Q(n11456) );
  AND2X1 U11379 ( .IN1(n11272), .IN2(g2917), .Q(n11455) );
  OR2X1 U11380 ( .IN1(n11457), .IN2(n11458), .Q(n11449) );
  OR2X1 U11381 ( .IN1(n11459), .IN2(n11460), .Q(n11458) );
  AND2X1 U11382 ( .IN1(n11273), .IN2(g2852), .Q(n11460) );
  AND2X1 U11383 ( .IN1(n11283), .IN2(g2912), .Q(n11459) );
  OR2X1 U11384 ( .IN1(n11461), .IN2(n11462), .Q(n11457) );
  OR2X1 U11385 ( .IN1(n11463), .IN2(n11464), .Q(n11462) );
  AND2X1 U11386 ( .IN1(n11289), .IN2(g2999), .Q(n11464) );
  AND2X1 U11387 ( .IN1(n11281), .IN2(g2856), .Q(n11461) );
  OR2X1 U11388 ( .IN1(n11465), .IN2(n11466), .Q(n11444) );
  AND2X1 U11389 ( .IN1(n11401), .IN2(g1129), .Q(n11466) );
  AND2X1 U11390 ( .IN1(n11400), .IN2(g1472), .Q(n11465) );
  OR2X1 U11391 ( .IN1(n10527), .IN2(g34971), .Q(g34915) );
  OR2X1 U11392 ( .IN1(n11467), .IN2(n11468), .Q(g34971) );
  OR2X1 U11393 ( .IN1(n11469), .IN2(n11470), .Q(n11468) );
  OR2X1 U11394 ( .IN1(n11471), .IN2(n11472), .Q(n11470) );
  AND2X1 U11395 ( .IN1(test_so64), .IN2(n11245), .Q(n11472) );
  AND2X1 U11396 ( .IN1(n11246), .IN2(n9247), .Q(n11471) );
  OR2X1 U11397 ( .IN1(n11473), .IN2(n11474), .Q(n11469) );
  AND2X1 U11398 ( .IN1(n11249), .IN2(g2704), .Q(n11474) );
  AND2X1 U11399 ( .IN1(n11250), .IN2(n9351), .Q(n11473) );
  OR2X1 U11400 ( .IN1(n11475), .IN2(n11476), .Q(n11467) );
  OR2X1 U11401 ( .IN1(n11477), .IN2(n11478), .Q(n11476) );
  AND2X1 U11402 ( .IN1(n11255), .IN2(g2145), .Q(n11478) );
  AND2X1 U11403 ( .IN1(n1340), .IN2(n11479), .Q(n11477) );
  OR2X1 U11404 ( .IN1(n11480), .IN2(n11481), .Q(n11479) );
  OR2X1 U11405 ( .IN1(n11482), .IN2(n11483), .Q(n11481) );
  OR2X1 U11406 ( .IN1(n11484), .IN2(n11485), .Q(n11483) );
  AND2X1 U11407 ( .IN1(n11267), .IN2(g562), .Q(n11485) );
  AND2X1 U11408 ( .IN1(n11265), .IN2(g599), .Q(n11484) );
  OR2X1 U11409 ( .IN1(n11486), .IN2(n11487), .Q(n11482) );
  OR2X1 U11410 ( .IN1(n11488), .IN2(n11489), .Q(n11487) );
  AND2X1 U11411 ( .IN1(n11274), .IN2(g199), .Q(n11489) );
  AND2X1 U11412 ( .IN1(n11273), .IN2(g4157), .Q(n11488) );
  AND2X1 U11413 ( .IN1(n11266), .IN2(test_so60), .Q(n11486) );
  OR2X1 U11414 ( .IN1(n11490), .IN2(n11491), .Q(n11480) );
  OR2X1 U11415 ( .IN1(n11492), .IN2(n11493), .Q(n11491) );
  AND2X1 U11416 ( .IN1(n11282), .IN2(g781), .Q(n11493) );
  AND2X1 U11417 ( .IN1(n11212), .IN2(g2984), .Q(n11492) );
  AND2X1 U11418 ( .IN1(n11494), .IN2(n11495), .Q(n11212) );
  AND2X1 U11419 ( .IN1(n5324), .IN2(test_so25), .Q(n11495) );
  AND2X1 U11420 ( .IN1(n11496), .IN2(n10519), .Q(n11494) );
  OR2X1 U11421 ( .IN1(n11497), .IN2(n11498), .Q(n11490) );
  OR2X1 U11422 ( .IN1(n11362), .IN2(n11499), .Q(n11498) );
  AND2X1 U11423 ( .IN1(n11289), .IN2(g2890), .Q(n11499) );
  AND2X1 U11424 ( .IN1(n11500), .IN2(n11501), .Q(n11289) );
  INVX0 U11425 ( .INP(n11502), .ZN(n11362) );
  OR2X1 U11426 ( .IN1(n11503), .IN2(n11504), .Q(n11502) );
  OR2X1 U11427 ( .IN1(n10519), .IN2(n11505), .Q(n11504) );
  INVX0 U11428 ( .INP(n11496), .ZN(n11505) );
  OR2X1 U11429 ( .IN1(test_so25), .IN2(n5324), .Q(n11503) );
  AND2X1 U11430 ( .IN1(g100), .IN2(n11288), .Q(n11497) );
  AND2X1 U11431 ( .IN1(n11501), .IN2(n11506), .Q(n11288) );
  AND2X1 U11432 ( .IN1(g28), .IN2(n11507), .Q(n11506) );
  OR2X1 U11433 ( .IN1(n11290), .IN2(n11508), .Q(n11475) );
  AND2X1 U11434 ( .IN1(n11292), .IN2(g4245), .Q(n11508) );
  AND2X1 U11435 ( .IN1(n11500), .IN2(n11509), .Q(n11292) );
  AND2X1 U11436 ( .IN1(n1340), .IN2(n11510), .Q(n11290) );
  AND2X1 U11437 ( .IN1(n10902), .IN2(n11511), .Q(n11510) );
  OR2X1 U11438 ( .IN1(n11512), .IN2(n11282), .Q(n11511) );
  AND2X1 U11439 ( .IN1(n11513), .IN2(n11500), .Q(n11282) );
  OR2X1 U11440 ( .IN1(n10527), .IN2(g34970), .Q(g34913) );
  OR2X1 U11441 ( .IN1(n11514), .IN2(n11515), .Q(g34970) );
  OR2X1 U11442 ( .IN1(n11516), .IN2(n11517), .Q(n11515) );
  OR2X1 U11443 ( .IN1(n11518), .IN2(n11519), .Q(n11517) );
  AND2X1 U11444 ( .IN1(n1340), .IN2(n11520), .Q(n11519) );
  OR2X1 U11445 ( .IN1(n11521), .IN2(n11522), .Q(n11520) );
  OR2X1 U11446 ( .IN1(n11523), .IN2(n11524), .Q(n11522) );
  OR2X1 U11447 ( .IN1(n11525), .IN2(n11526), .Q(n11524) );
  AND2X1 U11448 ( .IN1(n11267), .IN2(g595), .Q(n11526) );
  AND2X1 U11449 ( .IN1(n11265), .IN2(n9340), .Q(n11525) );
  OR2X1 U11450 ( .IN1(n11527), .IN2(n11528), .Q(n11523) );
  AND2X1 U11451 ( .IN1(n11266), .IN2(g776), .Q(n11528) );
  AND2X1 U11452 ( .IN1(n11274), .IN2(g538), .Q(n11527) );
  AND2X1 U11453 ( .IN1(n11513), .IN2(n11529), .Q(n11274) );
  OR2X1 U11454 ( .IN1(n11530), .IN2(n11531), .Q(n11521) );
  OR2X1 U11455 ( .IN1(n11532), .IN2(n11533), .Q(n11531) );
  AND2X1 U11456 ( .IN1(n11272), .IN2(g2902), .Q(n11533) );
  AND2X1 U11457 ( .IN1(n11534), .IN2(n11535), .Q(n11272) );
  AND2X1 U11458 ( .IN1(n11496), .IN2(n5324), .Q(n11535) );
  AND2X1 U11459 ( .IN1(n11273), .IN2(g2844), .Q(n11532) );
  AND2X1 U11460 ( .IN1(n11529), .IN2(n11536), .Q(n11273) );
  OR2X1 U11461 ( .IN1(n11537), .IN2(n11538), .Q(n11530) );
  OR2X1 U11462 ( .IN1(n11463), .IN2(n11539), .Q(n11538) );
  AND2X1 U11463 ( .IN1(n11281), .IN2(g2848), .Q(n11539) );
  AND2X1 U11464 ( .IN1(n11500), .IN2(n11536), .Q(n11281) );
  AND2X1 U11465 ( .IN1(g9), .IN2(n11534), .Q(n11536) );
  AND2X1 U11466 ( .IN1(n11512), .IN2(n10895), .Q(n11463) );
  OR2X1 U11467 ( .IN1(n11266), .IN2(n11540), .Q(n11512) );
  OR2X1 U11468 ( .IN1(n11267), .IN2(n11265), .Q(n11540) );
  AND2X1 U11469 ( .IN1(n2552), .IN2(n11529), .Q(n11265) );
  AND2X1 U11470 ( .IN1(n2552), .IN2(n11541), .Q(n11267) );
  AND2X1 U11471 ( .IN1(n11507), .IN2(n11542), .Q(n11266) );
  AND2X1 U11472 ( .IN1(g28), .IN2(n11513), .Q(n11542) );
  AND2X1 U11473 ( .IN1(n11534), .IN2(n5468), .Q(n11513) );
  AND2X1 U11474 ( .IN1(test_so1), .IN2(n11283), .Q(n11537) );
  AND2X1 U11475 ( .IN1(n11534), .IN2(n11543), .Q(n11283) );
  AND2X1 U11476 ( .IN1(g28), .IN2(n11496), .Q(n11543) );
  AND2X1 U11477 ( .IN1(n11544), .IN2(n11545), .Q(n11496) );
  AND2X1 U11478 ( .IN1(test_so85), .IN2(n3395), .Q(n11545) );
  AND2X1 U11479 ( .IN1(g9), .IN2(g8), .Q(n11544) );
  AND2X1 U11480 ( .IN1(n5477), .IN2(n10519), .Q(n11534) );
  AND2X1 U11481 ( .IN1(n11335), .IN2(g4917), .Q(n11518) );
  AND2X1 U11482 ( .IN1(n2527), .IN2(n11546), .Q(n11335) );
  AND2X1 U11483 ( .IN1(n11500), .IN2(n1340), .Q(n11546) );
  OR2X1 U11484 ( .IN1(n11547), .IN2(n11548), .Q(n11516) );
  AND2X1 U11485 ( .IN1(n11336), .IN2(g4727), .Q(n11548) );
  AND2X1 U11486 ( .IN1(n2527), .IN2(n11549), .Q(n11336) );
  AND2X1 U11487 ( .IN1(n11249), .IN2(g3853), .Q(n11547) );
  AND2X1 U11488 ( .IN1(n11509), .IN2(n11541), .Q(n11249) );
  AND2X1 U11489 ( .IN1(n5324), .IN2(n11507), .Q(n11541) );
  INVX0 U11490 ( .INP(n11550), .ZN(n11507) );
  OR2X1 U11491 ( .IN1(n5469), .IN2(n11551), .Q(n11550) );
  OR2X1 U11492 ( .IN1(n11552), .IN2(n11553), .Q(n11514) );
  OR2X1 U11493 ( .IN1(n11554), .IN2(n11555), .Q(n11553) );
  AND2X1 U11494 ( .IN1(n11250), .IN2(n9322), .Q(n11555) );
  AND2X1 U11495 ( .IN1(n11229), .IN2(n11556), .Q(n11250) );
  AND2X1 U11496 ( .IN1(n11255), .IN2(g6199), .Q(n11554) );
  AND2X1 U11497 ( .IN1(n11529), .IN2(n11509), .Q(n11255) );
  INVX0 U11498 ( .INP(n11557), .ZN(n11509) );
  OR2X1 U11499 ( .IN1(n11558), .IN2(n11559), .Q(n11557) );
  OR2X1 U11500 ( .IN1(n10519), .IN2(n11556), .Q(n11559) );
  INVX0 U11501 ( .INP(n1340), .ZN(n11556) );
  OR2X1 U11502 ( .IN1(test_so25), .IN2(n5468), .Q(n11558) );
  OR2X1 U11503 ( .IN1(n11560), .IN2(n11561), .Q(n11552) );
  AND2X1 U11504 ( .IN1(n11401), .IN2(g956), .Q(n11561) );
  AND2X1 U11505 ( .IN1(n11246), .IN2(n5286), .Q(n11401) );
  AND2X1 U11506 ( .IN1(n1340), .IN2(n11562), .Q(n11246) );
  AND2X1 U11507 ( .IN1(n11500), .IN2(n2552), .Q(n11562) );
  AND2X1 U11508 ( .IN1(n5469), .IN2(n11563), .Q(n11500) );
  AND2X1 U11509 ( .IN1(g28), .IN2(n11564), .Q(n11563) );
  AND2X1 U11510 ( .IN1(n11400), .IN2(g1300), .Q(n11560) );
  AND2X1 U11511 ( .IN1(n11245), .IN2(n2549), .Q(n11400) );
  AND2X1 U11512 ( .IN1(n11501), .IN2(n11549), .Q(n11245) );
  AND2X1 U11513 ( .IN1(n11529), .IN2(n1340), .Q(n11549) );
  AND2X1 U11514 ( .IN1(n11565), .IN2(n11566), .Q(n1340) );
  AND2X1 U11515 ( .IN1(n11229), .IN2(n11238), .Q(n11566) );
  AND2X1 U11516 ( .IN1(n11567), .IN2(g54), .Q(n11238) );
  INVX0 U11517 ( .INP(g56), .ZN(n11567) );
  INVX0 U11518 ( .INP(g53), .ZN(n11229) );
  INVX0 U11519 ( .INP(n11568), .ZN(n11565) );
  OR2X1 U11520 ( .IN1(test_so74), .IN2(g57), .Q(n11568) );
  AND2X1 U11521 ( .IN1(n5469), .IN2(n11569), .Q(n11529) );
  AND2X1 U11522 ( .IN1(n5324), .IN2(n11564), .Q(n11569) );
  INVX0 U11523 ( .INP(n11551), .ZN(n11564) );
  OR2X1 U11524 ( .IN1(g6), .IN2(n11570), .Q(n11551) );
  OR2X1 U11525 ( .IN1(test_so85), .IN2(g8), .Q(n11570) );
  AND2X1 U11526 ( .IN1(n5468), .IN2(n11571), .Q(n11501) );
  AND2X1 U11527 ( .IN1(n10519), .IN2(test_so25), .Q(n11571) );
  OR2X1 U11528 ( .IN1(n11572), .IN2(n11573), .Q(g34911) );
  AND2X1 U11529 ( .IN1(n2404), .IN2(g554), .Q(n11573) );
  AND2X1 U11530 ( .IN1(n11574), .IN2(g807), .Q(n11572) );
  OR2X1 U11531 ( .IN1(n2405), .IN2(n10875), .Q(n11574) );
  OR2X1 U11532 ( .IN1(n11575), .IN2(n11576), .Q(g34882) );
  AND2X1 U11533 ( .IN1(n11577), .IN2(n10763), .Q(n11576) );
  OR2X1 U11534 ( .IN1(n11578), .IN2(n11579), .Q(n11577) );
  OR2X1 U11535 ( .IN1(n11580), .IN2(n11581), .Q(n11579) );
  AND2X1 U11536 ( .IN1(n11582), .IN2(n5348), .Q(n11581) );
  AND2X1 U11537 ( .IN1(n11583), .IN2(n10552), .Q(n11582) );
  AND2X1 U11538 ( .IN1(n11584), .IN2(g4358), .Q(n11580) );
  AND2X1 U11539 ( .IN1(test_so81), .IN2(g4340), .Q(n11584) );
  AND2X1 U11540 ( .IN1(n11585), .IN2(n11586), .Q(n11578) );
  AND2X1 U11541 ( .IN1(n5653), .IN2(n11587), .Q(n11585) );
  OR2X1 U11542 ( .IN1(g4358), .IN2(n11583), .Q(n11587) );
  OR2X1 U11543 ( .IN1(n11588), .IN2(n11589), .Q(n11583) );
  OR2X1 U11544 ( .IN1(test_so81), .IN2(g4340), .Q(n11589) );
  OR2X1 U11545 ( .IN1(n11590), .IN2(n11591), .Q(n11588) );
  AND2X1 U11546 ( .IN1(n11592), .IN2(g4332), .Q(n11591) );
  AND2X1 U11547 ( .IN1(n5506), .IN2(g4311), .Q(n11592) );
  AND2X1 U11548 ( .IN1(n5540), .IN2(n11593), .Q(n11590) );
  OR2X1 U11549 ( .IN1(n11594), .IN2(n11595), .Q(n11593) );
  OR2X1 U11550 ( .IN1(n11596), .IN2(n11597), .Q(n11595) );
  AND2X1 U11551 ( .IN1(n11598), .IN2(n5506), .Q(n11597) );
  AND2X1 U11552 ( .IN1(g90), .IN2(n5634), .Q(n11598) );
  AND2X1 U11553 ( .IN1(n10434), .IN2(g4322), .Q(n11596) );
  AND2X1 U11554 ( .IN1(n10921), .IN2(g4366), .Q(n11575) );
  OR2X1 U11555 ( .IN1(n11599), .IN2(n11600), .Q(g34881) );
  OR2X1 U11556 ( .IN1(n11601), .IN2(n11602), .Q(n11600) );
  AND2X1 U11557 ( .IN1(n2405), .IN2(n5479), .Q(n11602) );
  AND2X1 U11558 ( .IN1(n11603), .IN2(g807), .Q(n11601) );
  AND2X1 U11559 ( .IN1(n2404), .IN2(n11604), .Q(n11603) );
  INVX0 U11560 ( .INP(n2405), .ZN(n11604) );
  AND2X1 U11561 ( .IN1(n10918), .IN2(g794), .Q(n11599) );
  OR2X1 U11562 ( .IN1(n11605), .IN2(n11606), .Q(g34880) );
  OR2X1 U11563 ( .IN1(n11607), .IN2(n11608), .Q(n11606) );
  AND2X1 U11564 ( .IN1(n2422), .IN2(n19032), .Q(n11608) );
  AND2X1 U11565 ( .IN1(n11609), .IN2(n9340), .Q(n11607) );
  AND2X1 U11566 ( .IN1(n2421), .IN2(n11610), .Q(n11609) );
  INVX0 U11567 ( .INP(n2422), .ZN(n11610) );
  AND2X1 U11568 ( .IN1(n10916), .IN2(g626), .Q(n11605) );
  OR2X1 U11569 ( .IN1(n11611), .IN2(n11612), .Q(g34850) );
  OR2X1 U11570 ( .IN1(n11613), .IN2(n11614), .Q(n11612) );
  AND2X1 U11571 ( .IN1(n2419), .IN2(n5291), .Q(n11614) );
  AND2X1 U11572 ( .IN1(n11615), .IN2(g794), .Q(n11613) );
  AND2X1 U11573 ( .IN1(n2404), .IN2(n11616), .Q(n11615) );
  INVX0 U11574 ( .INP(n2419), .ZN(n11616) );
  AND2X1 U11575 ( .IN1(n10916), .IN2(g790), .Q(n11611) );
  OR2X1 U11576 ( .IN1(n11617), .IN2(n11618), .Q(g34849) );
  OR2X1 U11577 ( .IN1(n11619), .IN2(n11620), .Q(n11618) );
  AND2X1 U11578 ( .IN1(n2423), .IN2(n5288), .Q(n11620) );
  AND2X1 U11579 ( .IN1(n11621), .IN2(g626), .Q(n11619) );
  AND2X1 U11580 ( .IN1(n2421), .IN2(n11622), .Q(n11621) );
  INVX0 U11581 ( .INP(n2423), .ZN(n11622) );
  AND2X1 U11582 ( .IN1(n10916), .IN2(g622), .Q(n11617) );
  AND2X1 U11583 ( .IN1(n11623), .IN2(g4369), .Q(g34839) );
  OR2X1 U11584 ( .IN1(g4366), .IN2(n11624), .Q(n11623) );
  OR2X1 U11585 ( .IN1(n11625), .IN2(n11626), .Q(n11624) );
  AND2X1 U11586 ( .IN1(n11627), .IN2(g4332), .Q(n11626) );
  OR2X1 U11587 ( .IN1(n11628), .IN2(n11629), .Q(n11627) );
  OR2X1 U11588 ( .IN1(n11630), .IN2(g4311), .Q(n11629) );
  AND2X1 U11589 ( .IN1(n5540), .IN2(n11631), .Q(n11625) );
  OR2X1 U11590 ( .IN1(g4311), .IN2(n11632), .Q(n11631) );
  OR2X1 U11591 ( .IN1(g73), .IN2(n11630), .Q(n11632) );
  OR2X1 U11592 ( .IN1(n11633), .IN2(n11634), .Q(g34808) );
  AND2X1 U11593 ( .IN1(n11635), .IN2(n10763), .Q(n11634) );
  OR2X1 U11594 ( .IN1(g2965), .IN2(n11636), .Q(n11635) );
  OR2X1 U11595 ( .IN1(n11637), .IN2(n11638), .Q(n11636) );
  AND2X1 U11596 ( .IN1(n10916), .IN2(g2955), .Q(n11633) );
  OR2X1 U11597 ( .IN1(n11639), .IN2(n11640), .Q(g34807) );
  AND2X1 U11598 ( .IN1(n11641), .IN2(n10763), .Q(n11640) );
  OR2X1 U11599 ( .IN1(n11642), .IN2(n11643), .Q(n11641) );
  OR2X1 U11600 ( .IN1(g2946), .IN2(n11644), .Q(n11643) );
  OR2X1 U11601 ( .IN1(n11645), .IN2(g2955), .Q(n11644) );
  OR2X1 U11602 ( .IN1(n11646), .IN2(n11647), .Q(n11642) );
  OR2X1 U11603 ( .IN1(n11648), .IN2(n11649), .Q(n11647) );
  AND2X1 U11604 ( .IN1(n10916), .IN2(g2941), .Q(n11639) );
  OR2X1 U11605 ( .IN1(n11650), .IN2(n11651), .Q(g34806) );
  AND2X1 U11606 ( .IN1(n11652), .IN2(n10763), .Q(n11651) );
  OR2X1 U11607 ( .IN1(g4153), .IN2(n11653), .Q(n11652) );
  OR2X1 U11608 ( .IN1(g2941), .IN2(g4072), .Q(n11653) );
  AND2X1 U11609 ( .IN1(n10916), .IN2(g2927), .Q(n11650) );
  AND2X1 U11610 ( .IN1(n11654), .IN2(n10763), .Q(g34805) );
  OR2X1 U11611 ( .IN1(g2932), .IN2(g2999), .Q(n11654) );
  OR2X1 U11612 ( .IN1(n11655), .IN2(n11656), .Q(g34804) );
  AND2X1 U11613 ( .IN1(n11657), .IN2(n10763), .Q(n11656) );
  OR2X1 U11614 ( .IN1(g2975), .IN2(n11658), .Q(n11657) );
  OR2X1 U11615 ( .IN1(n5796), .IN2(n5630), .Q(n11658) );
  AND2X1 U11616 ( .IN1(n10916), .IN2(g2965), .Q(n11655) );
  OR2X1 U11617 ( .IN1(n11659), .IN2(n11660), .Q(g34803) );
  AND2X1 U11618 ( .IN1(n11661), .IN2(n10763), .Q(n11660) );
  OR2X1 U11619 ( .IN1(g2927), .IN2(n11662), .Q(n11661) );
  OR2X1 U11620 ( .IN1(g2932), .IN2(n11663), .Q(n11662) );
  AND2X1 U11621 ( .IN1(n10916), .IN2(g2917), .Q(n11659) );
  OR2X1 U11622 ( .IN1(n11664), .IN2(n11665), .Q(g34802) );
  AND2X1 U11623 ( .IN1(n11666), .IN2(n10763), .Q(n11665) );
  OR2X1 U11624 ( .IN1(g2917), .IN2(n11667), .Q(n11666) );
  OR2X1 U11625 ( .IN1(n11668), .IN2(n11669), .Q(n11667) );
  AND2X1 U11626 ( .IN1(n10916), .IN2(g2902), .Q(n11664) );
  OR2X1 U11627 ( .IN1(n11670), .IN2(n11671), .Q(g34801) );
  AND2X1 U11628 ( .IN1(n11672), .IN2(n10764), .Q(n11671) );
  OR2X1 U11629 ( .IN1(n11673), .IN2(n11674), .Q(n11672) );
  OR2X1 U11630 ( .IN1(g301), .IN2(g209), .Q(n11674) );
  OR2X1 U11631 ( .IN1(n5520), .IN2(g2902), .Q(n11673) );
  AND2X1 U11632 ( .IN1(n10916), .IN2(g2970), .Q(n11670) );
  OR2X1 U11633 ( .IN1(n11675), .IN2(n11676), .Q(g34800) );
  AND2X1 U11634 ( .IN1(n11677), .IN2(n10764), .Q(n11676) );
  OR2X1 U11635 ( .IN1(test_so14), .IN2(test_so74), .Q(n11677) );
  AND2X1 U11636 ( .IN1(n10916), .IN2(g2886), .Q(n11675) );
  OR2X1 U11637 ( .IN1(n11678), .IN2(n11679), .Q(g34799) );
  AND2X1 U11638 ( .IN1(n11680), .IN2(n10764), .Q(n11679) );
  OR2X1 U11639 ( .IN1(n11663), .IN2(g2890), .Q(n11680) );
  INVX0 U11640 ( .INP(g44), .ZN(n11663) );
  AND2X1 U11641 ( .IN1(n10916), .IN2(g2873), .Q(n11678) );
  OR2X1 U11642 ( .IN1(n11681), .IN2(n11682), .Q(g34798) );
  AND2X1 U11643 ( .IN1(n11683), .IN2(n10764), .Q(n11682) );
  OR2X1 U11644 ( .IN1(g2946), .IN2(g2886), .Q(n11683) );
  AND2X1 U11645 ( .IN1(n10916), .IN2(g2878), .Q(n11681) );
  OR2X1 U11646 ( .IN1(n11684), .IN2(n11685), .Q(g34797) );
  AND2X1 U11647 ( .IN1(n11686), .IN2(n10764), .Q(n11685) );
  OR2X1 U11648 ( .IN1(n11638), .IN2(g2878), .Q(n11686) );
  INVX0 U11649 ( .INP(g91), .ZN(n11638) );
  AND2X1 U11650 ( .IN1(n10916), .IN2(g2882), .Q(n11684) );
  OR2X1 U11651 ( .IN1(n11687), .IN2(n11688), .Q(g34796) );
  AND2X1 U11652 ( .IN1(n11689), .IN2(n10764), .Q(n11688) );
  OR2X1 U11653 ( .IN1(n11637), .IN2(g2882), .Q(n11689) );
  OR2X1 U11654 ( .IN1(n11690), .IN2(n11691), .Q(n11637) );
  AND2X1 U11655 ( .IN1(n10916), .IN2(g2898), .Q(n11687) );
  OR2X1 U11656 ( .IN1(n11692), .IN2(n11693), .Q(g34795) );
  AND2X1 U11657 ( .IN1(n11694), .IN2(n10764), .Q(n11693) );
  OR2X1 U11658 ( .IN1(n11646), .IN2(g2898), .Q(n11694) );
  INVX0 U11659 ( .INP(n11695), .ZN(n11646) );
  AND2X1 U11660 ( .IN1(n11696), .IN2(n11697), .Q(n11695) );
  AND2X1 U11661 ( .IN1(n11698), .IN2(n11699), .Q(n11697) );
  AND2X1 U11662 ( .IN1(n10916), .IN2(g2864), .Q(n11692) );
  OR2X1 U11663 ( .IN1(n11700), .IN2(n11701), .Q(g34794) );
  AND2X1 U11664 ( .IN1(n11702), .IN2(n10764), .Q(n11701) );
  OR2X1 U11665 ( .IN1(n11645), .IN2(g2864), .Q(n11702) );
  INVX0 U11666 ( .INP(n11703), .ZN(n11645) );
  AND2X1 U11667 ( .IN1(n11704), .IN2(n11705), .Q(n11703) );
  AND2X1 U11668 ( .IN1(n10484), .IN2(n11706), .Q(n11705) );
  AND2X1 U11669 ( .IN1(n11707), .IN2(n11708), .Q(n11704) );
  AND2X1 U11670 ( .IN1(n10564), .IN2(n11709), .Q(n11708) );
  AND2X1 U11671 ( .IN1(n10917), .IN2(g2856), .Q(n11700) );
  OR2X1 U11672 ( .IN1(n11710), .IN2(n11711), .Q(g34793) );
  AND2X1 U11673 ( .IN1(n11712), .IN2(n10764), .Q(n11711) );
  OR2X1 U11674 ( .IN1(n11649), .IN2(g2856), .Q(n11712) );
  OR2X1 U11675 ( .IN1(n11713), .IN2(n11714), .Q(n11649) );
  AND2X1 U11676 ( .IN1(n10917), .IN2(g2848), .Q(n11710) );
  OR2X1 U11677 ( .IN1(n11715), .IN2(n11716), .Q(g34792) );
  AND2X1 U11678 ( .IN1(n11717), .IN2(n10765), .Q(n11716) );
  OR2X1 U11679 ( .IN1(n11648), .IN2(g2848), .Q(n11717) );
  OR2X1 U11680 ( .IN1(n11718), .IN2(n11719), .Q(n11648) );
  AND2X1 U11681 ( .IN1(n10917), .IN2(g29214), .Q(n11715) );
  OR2X1 U11682 ( .IN1(n11720), .IN2(n11721), .Q(g34791) );
  OR2X1 U11683 ( .IN1(n11722), .IN2(n11723), .Q(n11721) );
  AND2X1 U11684 ( .IN1(n2425), .IN2(n5292), .Q(n11723) );
  AND2X1 U11685 ( .IN1(n11724), .IN2(g790), .Q(n11722) );
  AND2X1 U11686 ( .IN1(n2404), .IN2(n11725), .Q(n11724) );
  INVX0 U11687 ( .INP(n2425), .ZN(n11725) );
  AND2X1 U11688 ( .IN1(n10917), .IN2(g785), .Q(n11720) );
  OR2X1 U11689 ( .IN1(n11726), .IN2(n11727), .Q(g34790) );
  OR2X1 U11690 ( .IN1(n11728), .IN2(n11729), .Q(n11727) );
  AND2X1 U11691 ( .IN1(n2427), .IN2(n5672), .Q(n11729) );
  AND2X1 U11692 ( .IN1(n11730), .IN2(g622), .Q(n11728) );
  AND2X1 U11693 ( .IN1(n2421), .IN2(n11731), .Q(n11730) );
  INVX0 U11694 ( .INP(n2427), .ZN(n11731) );
  AND2X1 U11695 ( .IN1(n10917), .IN2(g617), .Q(n11726) );
  AND2X1 U11696 ( .IN1(n11732), .IN2(g890), .Q(g34788) );
  OR2X1 U11697 ( .IN1(n10116), .IN2(n11733), .Q(n11732) );
  OR2X1 U11698 ( .IN1(n11734), .IN2(n11735), .Q(g34783) );
  AND2X1 U11699 ( .IN1(n11736), .IN2(n11737), .Q(n11735) );
  AND2X1 U11700 ( .IN1(n11738), .IN2(n11739), .Q(n11736) );
  AND2X1 U11701 ( .IN1(n11740), .IN2(n11741), .Q(n11734) );
  AND2X1 U11702 ( .IN1(n11742), .IN2(n11743), .Q(n11740) );
  OR2X1 U11703 ( .IN1(n11744), .IN2(n11745), .Q(g34735) );
  AND2X1 U11704 ( .IN1(n11746), .IN2(n10765), .Q(n11745) );
  OR2X1 U11705 ( .IN1(test_so63), .IN2(g4300), .Q(n11746) );
  INVX0 U11706 ( .INP(n11747), .ZN(n11744) );
  OR2X1 U11707 ( .IN1(n10739), .IN2(n10492), .Q(n11747) );
  OR2X1 U11708 ( .IN1(n11748), .IN2(n11749), .Q(g34734) );
  AND2X1 U11709 ( .IN1(n11750), .IN2(n10765), .Q(n11749) );
  OR2X1 U11710 ( .IN1(g4072), .IN2(g4176), .Q(n11750) );
  AND2X1 U11711 ( .IN1(n10917), .IN2(g4172), .Q(n11748) );
  AND2X1 U11712 ( .IN1(n11751), .IN2(n10765), .Q(g34733) );
  OR2X1 U11713 ( .IN1(g4153), .IN2(g4172), .Q(n11751) );
  OR2X1 U11714 ( .IN1(n11752), .IN2(n11753), .Q(g34732) );
  AND2X1 U11715 ( .IN1(n10917), .IN2(g2999), .Q(n11753) );
  AND2X1 U11716 ( .IN1(n10811), .IN2(g2994), .Q(n11752) );
  OR2X1 U11717 ( .IN1(n11754), .IN2(n11755), .Q(g34731) );
  AND2X1 U11718 ( .IN1(n11756), .IN2(n10765), .Q(n11755) );
  OR2X1 U11719 ( .IN1(test_so64), .IN2(n11668), .Q(n11756) );
  AND2X1 U11720 ( .IN1(n10917), .IN2(g1283), .Q(n11754) );
  OR2X1 U11721 ( .IN1(n11757), .IN2(n11758), .Q(g34730) );
  AND2X1 U11722 ( .IN1(n11759), .IN2(n10765), .Q(n11758) );
  OR2X1 U11723 ( .IN1(g1283), .IN2(g1277), .Q(n11759) );
  INVX0 U11724 ( .INP(n11760), .ZN(n11757) );
  OR2X1 U11725 ( .IN1(n10739), .IN2(n10010), .Q(n11760) );
  OR2X1 U11726 ( .IN1(n2499), .IN2(n11761), .Q(g34729) );
  OR2X1 U11727 ( .IN1(n11762), .IN2(n11763), .Q(n11761) );
  AND2X1 U11728 ( .IN1(n10917), .IN2(g1291), .Q(n11763) );
  AND2X1 U11729 ( .IN1(n5796), .IN2(n10765), .Q(n11762) );
  OR2X1 U11730 ( .IN1(n11764), .IN2(n11765), .Q(g34728) );
  AND2X1 U11731 ( .IN1(n11766), .IN2(n10765), .Q(n11765) );
  OR2X1 U11732 ( .IN1(n11669), .IN2(n9247), .Q(n11766) );
  AND2X1 U11733 ( .IN1(n10917), .IN2(g939), .Q(n11764) );
  OR2X1 U11734 ( .IN1(n11767), .IN2(n11768), .Q(g34727) );
  AND2X1 U11735 ( .IN1(n11769), .IN2(n10765), .Q(n11768) );
  OR2X1 U11736 ( .IN1(test_so52), .IN2(g939), .Q(n11769) );
  INVX0 U11737 ( .INP(n11770), .ZN(n11767) );
  OR2X1 U11738 ( .IN1(n10739), .IN2(n10011), .Q(n11770) );
  OR2X1 U11739 ( .IN1(n2505), .IN2(n11771), .Q(g34726) );
  OR2X1 U11740 ( .IN1(n11772), .IN2(n11773), .Q(n11771) );
  AND2X1 U11741 ( .IN1(n10917), .IN2(g947), .Q(n11773) );
  AND2X1 U11742 ( .IN1(n5630), .IN2(n10766), .Q(n11772) );
  OR2X1 U11743 ( .IN1(n11774), .IN2(n11775), .Q(g34725) );
  OR2X1 U11744 ( .IN1(n11776), .IN2(n11777), .Q(n11775) );
  AND2X1 U11745 ( .IN1(n2485), .IN2(n5293), .Q(n11777) );
  AND2X1 U11746 ( .IN1(n11778), .IN2(g785), .Q(n11776) );
  AND2X1 U11747 ( .IN1(n2404), .IN2(n11779), .Q(n11778) );
  INVX0 U11748 ( .INP(n2485), .ZN(n11779) );
  AND2X1 U11749 ( .IN1(n10917), .IN2(g781), .Q(n11774) );
  OR2X1 U11750 ( .IN1(n11780), .IN2(n11781), .Q(g34724) );
  OR2X1 U11751 ( .IN1(n11782), .IN2(n11783), .Q(n11781) );
  AND2X1 U11752 ( .IN1(n2487), .IN2(n5339), .Q(n11783) );
  AND2X1 U11753 ( .IN1(n11784), .IN2(g617), .Q(n11782) );
  AND2X1 U11754 ( .IN1(n2421), .IN2(n11785), .Q(n11784) );
  INVX0 U11755 ( .INP(n2487), .ZN(n11785) );
  AND2X1 U11756 ( .IN1(n10917), .IN2(g613), .Q(n11780) );
  OR2X1 U11757 ( .IN1(n11786), .IN2(n11787), .Q(g34723) );
  AND2X1 U11758 ( .IN1(n11788), .IN2(n10766), .Q(n11787) );
  OR2X1 U11759 ( .IN1(g301), .IN2(g534), .Q(n11788) );
  AND2X1 U11760 ( .IN1(test_so41), .IN2(n10894), .Q(n11786) );
  OR2X1 U11761 ( .IN1(n11789), .IN2(n11790), .Q(g34722) );
  AND2X1 U11762 ( .IN1(n11791), .IN2(n10766), .Q(n11790) );
  OR2X1 U11763 ( .IN1(n5520), .IN2(g546), .Q(n11791) );
  AND2X1 U11764 ( .IN1(n10917), .IN2(g538), .Q(n11789) );
  OR2X1 U11765 ( .IN1(n11792), .IN2(n11793), .Q(g34721) );
  AND2X1 U11766 ( .IN1(n11794), .IN2(n10766), .Q(n11793) );
  OR2X1 U11767 ( .IN1(g199), .IN2(g222), .Q(n11794) );
  AND2X1 U11768 ( .IN1(g29221), .IN2(n10896), .Q(n11792) );
  OR2X1 U11769 ( .IN1(n11795), .IN2(n11796), .Q(g34720) );
  AND2X1 U11770 ( .IN1(n11797), .IN2(n10766), .Q(n11796) );
  OR2X1 U11771 ( .IN1(n5657), .IN2(g550), .Q(n11797) );
  AND2X1 U11772 ( .IN1(n10917), .IN2(g534), .Q(n11795) );
  AND2X1 U11773 ( .IN1(n11798), .IN2(n10766), .Q(g34719) );
  OR2X1 U11774 ( .IN1(g209), .IN2(g538), .Q(n11798) );
  AND2X1 U11775 ( .IN1(n10807), .IN2(g6545), .Q(g34647) );
  AND2X1 U11776 ( .IN1(n10807), .IN2(g6199), .Q(g34646) );
  AND2X1 U11777 ( .IN1(n10808), .IN2(g5853), .Q(g34645) );
  AND2X1 U11778 ( .IN1(n10807), .IN2(g5507), .Q(g34644) );
  AND2X1 U11779 ( .IN1(n10808), .IN2(g5160), .Q(g34643) );
  OR2X1 U11780 ( .IN1(n11799), .IN2(n11800), .Q(g34642) );
  AND2X1 U11781 ( .IN1(n10917), .IN2(g4912), .Q(n11800) );
  INVX0 U11782 ( .INP(n11801), .ZN(n11799) );
  OR2X1 U11783 ( .IN1(n10887), .IN2(n5879), .Q(n11801) );
  OR2X1 U11784 ( .IN1(n11802), .IN2(n11803), .Q(g34641) );
  AND2X1 U11785 ( .IN1(n10917), .IN2(g4907), .Q(n11803) );
  AND2X1 U11786 ( .IN1(n10807), .IN2(g4912), .Q(n11802) );
  OR2X1 U11787 ( .IN1(n11804), .IN2(n11805), .Q(g34640) );
  AND2X1 U11788 ( .IN1(n10917), .IN2(g4922), .Q(n11805) );
  AND2X1 U11789 ( .IN1(n10807), .IN2(g4907), .Q(n11804) );
  OR2X1 U11790 ( .IN1(n11806), .IN2(n11807), .Q(g34639) );
  AND2X1 U11791 ( .IN1(n10917), .IN2(g4917), .Q(n11807) );
  AND2X1 U11792 ( .IN1(n10808), .IN2(g4922), .Q(n11806) );
  AND2X1 U11793 ( .IN1(n10807), .IN2(g4917), .Q(g34638) );
  OR2X1 U11794 ( .IN1(n11808), .IN2(n11809), .Q(g34637) );
  AND2X1 U11795 ( .IN1(n10918), .IN2(g4722), .Q(n11809) );
  INVX0 U11796 ( .INP(n11810), .ZN(n11808) );
  OR2X1 U11797 ( .IN1(n10887), .IN2(n5867), .Q(n11810) );
  OR2X1 U11798 ( .IN1(n11811), .IN2(n11812), .Q(g34636) );
  AND2X1 U11799 ( .IN1(n10918), .IN2(g4717), .Q(n11812) );
  AND2X1 U11800 ( .IN1(n10809), .IN2(g4722), .Q(n11811) );
  OR2X1 U11801 ( .IN1(n11813), .IN2(n11814), .Q(g34635) );
  AND2X1 U11802 ( .IN1(n10918), .IN2(g4732), .Q(n11814) );
  AND2X1 U11803 ( .IN1(n10808), .IN2(g4717), .Q(n11813) );
  OR2X1 U11804 ( .IN1(n11815), .IN2(n11816), .Q(g34634) );
  AND2X1 U11805 ( .IN1(n10918), .IN2(g4727), .Q(n11816) );
  AND2X1 U11806 ( .IN1(n10808), .IN2(g4732), .Q(n11815) );
  AND2X1 U11807 ( .IN1(n10807), .IN2(g4727), .Q(g34633) );
  OR2X1 U11808 ( .IN1(n11817), .IN2(n11818), .Q(g34632) );
  AND2X1 U11809 ( .IN1(test_so67), .IN2(n10894), .Q(n11818) );
  AND2X1 U11810 ( .IN1(n10809), .IN2(g4245), .Q(n11817) );
  OR2X1 U11811 ( .IN1(n11819), .IN2(n11820), .Q(g34631) );
  AND2X1 U11812 ( .IN1(n10918), .IN2(g4253), .Q(n11820) );
  AND2X1 U11813 ( .IN1(test_so67), .IN2(n10766), .Q(n11819) );
  OR2X1 U11814 ( .IN1(n11821), .IN2(n11822), .Q(g34630) );
  AND2X1 U11815 ( .IN1(n10918), .IN2(g4300), .Q(n11822) );
  AND2X1 U11816 ( .IN1(n10809), .IN2(g4253), .Q(n11821) );
  OR2X1 U11817 ( .IN1(n11823), .IN2(n11824), .Q(g34629) );
  AND2X1 U11818 ( .IN1(n10918), .IN2(g4146), .Q(n11824) );
  AND2X1 U11819 ( .IN1(n10808), .IN2(g4157), .Q(n11823) );
  OR2X1 U11820 ( .IN1(n11825), .IN2(n11826), .Q(g34628) );
  AND2X1 U11821 ( .IN1(n10918), .IN2(g4176), .Q(n11826) );
  AND2X1 U11822 ( .IN1(n10809), .IN2(g4146), .Q(n11825) );
  AND2X1 U11823 ( .IN1(n10808), .IN2(g3853), .Q(g34627) );
  AND2X1 U11824 ( .IN1(test_so45), .IN2(n10766), .Q(g34626) );
  AND2X1 U11825 ( .IN1(n10809), .IN2(g3151), .Q(g34625) );
  OR2X1 U11826 ( .IN1(n11827), .IN2(n11828), .Q(g34624) );
  AND2X1 U11827 ( .IN1(n10918), .IN2(g2994), .Q(n11828) );
  AND2X1 U11828 ( .IN1(n10809), .IN2(g2988), .Q(n11827) );
  OR2X1 U11829 ( .IN1(n11829), .IN2(n11830), .Q(g34623) );
  AND2X1 U11830 ( .IN1(test_so22), .IN2(n10894), .Q(n11830) );
  AND2X1 U11831 ( .IN1(n10809), .IN2(g2970), .Q(n11829) );
  OR2X1 U11832 ( .IN1(n11831), .IN2(n11832), .Q(g34622) );
  AND2X1 U11833 ( .IN1(n10918), .IN2(g2950), .Q(n11832) );
  AND2X1 U11834 ( .IN1(test_so22), .IN2(n10766), .Q(n11831) );
  OR2X1 U11835 ( .IN1(n11833), .IN2(n11834), .Q(g34621) );
  AND2X1 U11836 ( .IN1(n10918), .IN2(g2936), .Q(n11834) );
  AND2X1 U11837 ( .IN1(n10810), .IN2(g2950), .Q(n11833) );
  OR2X1 U11838 ( .IN1(n11835), .IN2(n11836), .Q(g34620) );
  AND2X1 U11839 ( .IN1(n10918), .IN2(g2922), .Q(n11836) );
  AND2X1 U11840 ( .IN1(n10810), .IN2(g2936), .Q(n11835) );
  OR2X1 U11841 ( .IN1(n11837), .IN2(n11838), .Q(g34619) );
  AND2X1 U11842 ( .IN1(n10918), .IN2(g2912), .Q(n11838) );
  AND2X1 U11843 ( .IN1(n10810), .IN2(g2922), .Q(n11837) );
  OR2X1 U11844 ( .IN1(n11839), .IN2(n11840), .Q(g34618) );
  AND2X1 U11845 ( .IN1(test_so1), .IN2(n10893), .Q(n11840) );
  AND2X1 U11846 ( .IN1(n10810), .IN2(g2912), .Q(n11839) );
  OR2X1 U11847 ( .IN1(n11841), .IN2(n11842), .Q(g34617) );
  AND2X1 U11848 ( .IN1(n10918), .IN2(g2984), .Q(n11842) );
  AND2X1 U11849 ( .IN1(test_so1), .IN2(n10767), .Q(n11841) );
  OR2X1 U11850 ( .IN1(n11843), .IN2(n11844), .Q(g34616) );
  AND2X1 U11851 ( .IN1(n10918), .IN2(g2988), .Q(n11844) );
  AND2X1 U11852 ( .IN1(n10869), .IN2(g2868), .Q(n11843) );
  OR2X1 U11853 ( .IN1(n11845), .IN2(n11846), .Q(g34615) );
  AND2X1 U11854 ( .IN1(n10918), .IN2(g2868), .Q(n11846) );
  AND2X1 U11855 ( .IN1(n10827), .IN2(g2873), .Q(n11845) );
  OR2X1 U11856 ( .IN1(n11847), .IN2(n11848), .Q(g34614) );
  AND2X1 U11857 ( .IN1(g37), .IN2(n10893), .Q(n11848) );
  AND2X1 U11858 ( .IN1(n10827), .IN2(g29214), .Q(n11847) );
  OR2X1 U11859 ( .IN1(n11849), .IN2(n11850), .Q(g34613) );
  AND2X1 U11860 ( .IN1(g37), .IN2(n10767), .Q(n11850) );
  AND2X1 U11861 ( .IN1(test_so95), .IN2(n10894), .Q(n11849) );
  OR2X1 U11862 ( .IN1(n11851), .IN2(n11852), .Q(g34612) );
  AND2X1 U11863 ( .IN1(n10918), .IN2(g2860), .Q(n11852) );
  AND2X1 U11864 ( .IN1(test_so95), .IN2(n10767), .Q(n11851) );
  OR2X1 U11865 ( .IN1(n11853), .IN2(n11854), .Q(g34611) );
  AND2X1 U11866 ( .IN1(n10918), .IN2(g2852), .Q(n11854) );
  AND2X1 U11867 ( .IN1(n10827), .IN2(g2860), .Q(n11853) );
  OR2X1 U11868 ( .IN1(n11855), .IN2(n11856), .Q(g34610) );
  AND2X1 U11869 ( .IN1(n10919), .IN2(g2844), .Q(n11856) );
  AND2X1 U11870 ( .IN1(n10827), .IN2(g2852), .Q(n11855) );
  OR2X1 U11871 ( .IN1(n11857), .IN2(n11858), .Q(g34609) );
  AND2X1 U11872 ( .IN1(n10919), .IN2(g2890), .Q(n11858) );
  AND2X1 U11873 ( .IN1(n10827), .IN2(g2844), .Q(n11857) );
  OR2X1 U11874 ( .IN1(n11859), .IN2(n11860), .Q(g34608) );
  AND2X1 U11875 ( .IN1(n10919), .IN2(g2697), .Q(n11860) );
  AND2X1 U11876 ( .IN1(n10827), .IN2(g2704), .Q(n11859) );
  OR2X1 U11877 ( .IN1(n11861), .IN2(n11862), .Q(g34607) );
  AND2X1 U11878 ( .IN1(n10919), .IN2(g2689), .Q(n11862) );
  AND2X1 U11879 ( .IN1(n10827), .IN2(g2697), .Q(n11861) );
  AND2X1 U11880 ( .IN1(n10827), .IN2(g2689), .Q(g34606) );
  OR2X1 U11881 ( .IN1(n11863), .IN2(n11864), .Q(g34605) );
  AND2X1 U11882 ( .IN1(n10919), .IN2(g2138), .Q(n11864) );
  AND2X1 U11883 ( .IN1(n10826), .IN2(g2145), .Q(n11863) );
  OR2X1 U11884 ( .IN1(n11865), .IN2(n11866), .Q(g34604) );
  AND2X1 U11885 ( .IN1(n10919), .IN2(g2130), .Q(n11866) );
  AND2X1 U11886 ( .IN1(n10826), .IN2(g2138), .Q(n11865) );
  AND2X1 U11887 ( .IN1(n10826), .IN2(g2130), .Q(g34603) );
  AND2X1 U11888 ( .IN1(n10826), .IN2(g1291), .Q(g34602) );
  AND2X1 U11889 ( .IN1(n10826), .IN2(g947), .Q(g34601) );
  OR2X1 U11890 ( .IN1(n11867), .IN2(n11868), .Q(g34600) );
  OR2X1 U11891 ( .IN1(n11869), .IN2(n11870), .Q(n11868) );
  AND2X1 U11892 ( .IN1(n2507), .IN2(n5551), .Q(n11870) );
  AND2X1 U11893 ( .IN1(n11871), .IN2(g781), .Q(n11869) );
  AND2X1 U11894 ( .IN1(n2404), .IN2(n11872), .Q(n11871) );
  INVX0 U11895 ( .INP(n2507), .ZN(n11872) );
  AND2X1 U11896 ( .IN1(n10919), .IN2(g776), .Q(n11867) );
  OR2X1 U11897 ( .IN1(n11873), .IN2(n11874), .Q(g34599) );
  OR2X1 U11898 ( .IN1(n11875), .IN2(n11876), .Q(n11874) );
  AND2X1 U11899 ( .IN1(n2509), .IN2(n5474), .Q(n11876) );
  AND2X1 U11900 ( .IN1(n11877), .IN2(g613), .Q(n11875) );
  AND2X1 U11901 ( .IN1(n2421), .IN2(n11878), .Q(n11877) );
  INVX0 U11902 ( .INP(n2509), .ZN(n11878) );
  AND2X1 U11903 ( .IN1(n10919), .IN2(g608), .Q(n11873) );
  OR2X1 U11904 ( .IN1(n11879), .IN2(n11880), .Q(g34598) );
  AND2X1 U11905 ( .IN1(g29221), .IN2(n10767), .Q(n11880) );
  AND2X1 U11906 ( .IN1(n10919), .IN2(g550), .Q(n11879) );
  OR2X1 U11907 ( .IN1(n11881), .IN2(n11882), .Q(g34468) );
  AND2X1 U11908 ( .IN1(n11883), .IN2(g4859), .Q(n11882) );
  AND2X1 U11909 ( .IN1(n11884), .IN2(g4854), .Q(n11881) );
  OR2X1 U11910 ( .IN1(n10889), .IN2(n11885), .Q(n11884) );
  AND2X1 U11911 ( .IN1(n11886), .IN2(n11887), .Q(n11885) );
  OR2X1 U11912 ( .IN1(n11888), .IN2(n11889), .Q(g34467) );
  AND2X1 U11913 ( .IN1(n10919), .IN2(g4849), .Q(n11889) );
  AND2X1 U11914 ( .IN1(n11890), .IN2(n11883), .Q(n11888) );
  XNOR2X1 U11915 ( .IN1(n11887), .IN2(n10041), .Q(n11890) );
  AND2X1 U11916 ( .IN1(g4849), .IN2(n2563), .Q(n11887) );
  OR2X1 U11917 ( .IN1(n11891), .IN2(n11892), .Q(g34466) );
  AND2X1 U11918 ( .IN1(n11893), .IN2(n5283), .Q(n11892) );
  AND2X1 U11919 ( .IN1(n11883), .IN2(g4843), .Q(n11893) );
  AND2X1 U11920 ( .IN1(n11894), .IN2(g4878), .Q(n11891) );
  OR2X1 U11921 ( .IN1(n10889), .IN2(n11895), .Q(n11894) );
  AND2X1 U11922 ( .IN1(n10478), .IN2(n11886), .Q(n11895) );
  OR2X1 U11923 ( .IN1(n11896), .IN2(n11897), .Q(g34465) );
  OR2X1 U11924 ( .IN1(n11898), .IN2(n11899), .Q(n11897) );
  AND2X1 U11925 ( .IN1(n2567), .IN2(n11883), .Q(n11899) );
  AND2X1 U11926 ( .IN1(n11900), .IN2(n10506), .Q(n11898) );
  AND2X1 U11927 ( .IN1(n11886), .IN2(n2563), .Q(n11900) );
  AND2X1 U11928 ( .IN1(n10919), .IN2(g4843), .Q(n11896) );
  OR2X1 U11929 ( .IN1(n11901), .IN2(n11902), .Q(g34464) );
  AND2X1 U11930 ( .IN1(n11903), .IN2(g4669), .Q(n11902) );
  AND2X1 U11931 ( .IN1(n11904), .IN2(g4664), .Q(n11901) );
  OR2X1 U11932 ( .IN1(n10889), .IN2(n11905), .Q(n11904) );
  AND2X1 U11933 ( .IN1(n11906), .IN2(n11907), .Q(n11905) );
  OR2X1 U11934 ( .IN1(n11908), .IN2(n11909), .Q(g34463) );
  AND2X1 U11935 ( .IN1(n10919), .IN2(g4659), .Q(n11909) );
  AND2X1 U11936 ( .IN1(n11910), .IN2(n11903), .Q(n11908) );
  XNOR2X1 U11937 ( .IN1(n11907), .IN2(n10055), .Q(n11910) );
  AND2X1 U11938 ( .IN1(g4659), .IN2(n2573), .Q(n11907) );
  OR2X1 U11939 ( .IN1(n11911), .IN2(n11912), .Q(g34462) );
  AND2X1 U11940 ( .IN1(n11913), .IN2(n5656), .Q(n11912) );
  AND2X1 U11941 ( .IN1(n11903), .IN2(test_so19), .Q(n11913) );
  AND2X1 U11942 ( .IN1(n11914), .IN2(g4688), .Q(n11911) );
  OR2X1 U11943 ( .IN1(n10890), .IN2(n11915), .Q(n11914) );
  AND2X1 U11944 ( .IN1(n11906), .IN2(n10567), .Q(n11915) );
  OR2X1 U11945 ( .IN1(n11916), .IN2(n11917), .Q(g34461) );
  OR2X1 U11946 ( .IN1(n11918), .IN2(n11919), .Q(n11917) );
  AND2X1 U11947 ( .IN1(n2577), .IN2(n11903), .Q(n11919) );
  AND2X1 U11948 ( .IN1(n11920), .IN2(n10509), .Q(n11918) );
  AND2X1 U11949 ( .IN1(n11906), .IN2(n2573), .Q(n11920) );
  AND2X1 U11950 ( .IN1(test_so19), .IN2(n10894), .Q(n11916) );
  OR2X1 U11951 ( .IN1(n11921), .IN2(n11922), .Q(g34460) );
  AND2X1 U11952 ( .IN1(g34025), .IN2(test_so3), .Q(n11922) );
  AND2X1 U11953 ( .IN1(n11923), .IN2(g4639), .Q(n11921) );
  OR2X1 U11954 ( .IN1(n10890), .IN2(n11924), .Q(n11923) );
  AND2X1 U11955 ( .IN1(n11925), .IN2(n10575), .Q(n11924) );
  OR2X1 U11956 ( .IN1(n11926), .IN2(n11927), .Q(g34459) );
  AND2X1 U11957 ( .IN1(n11928), .IN2(n10767), .Q(n11927) );
  OR2X1 U11958 ( .IN1(n11929), .IN2(n11930), .Q(n11928) );
  AND2X1 U11959 ( .IN1(n11931), .IN2(n11932), .Q(n11929) );
  OR2X1 U11960 ( .IN1(n11933), .IN2(g4340), .Q(n11931) );
  AND2X1 U11961 ( .IN1(test_so99), .IN2(n11934), .Q(n11933) );
  AND2X1 U11962 ( .IN1(n10919), .IN2(g4643), .Q(n11926) );
  OR2X1 U11963 ( .IN1(n11935), .IN2(n11936), .Q(g34458) );
  AND2X1 U11964 ( .IN1(test_so99), .IN2(n11937), .Q(n11936) );
  OR2X1 U11965 ( .IN1(n10890), .IN2(n11938), .Q(n11937) );
  AND2X1 U11966 ( .IN1(n11939), .IN2(n11940), .Q(n11938) );
  AND2X1 U11967 ( .IN1(test_so3), .IN2(g4639), .Q(n11940) );
  AND2X1 U11968 ( .IN1(n5844), .IN2(n11925), .Q(n11939) );
  AND2X1 U11969 ( .IN1(n11941), .IN2(g4633), .Q(n11935) );
  OR2X1 U11970 ( .IN1(n11942), .IN2(n11943), .Q(n11941) );
  AND2X1 U11971 ( .IN1(n11944), .IN2(n11925), .Q(n11942) );
  AND2X1 U11972 ( .IN1(n10826), .IN2(n10551), .Q(n11944) );
  OR2X1 U11973 ( .IN1(n11945), .IN2(n11946), .Q(g34457) );
  AND2X1 U11974 ( .IN1(test_so99), .IN2(n11943), .Q(n11946) );
  OR2X1 U11975 ( .IN1(n11947), .IN2(g34025), .Q(n11943) );
  AND2X1 U11976 ( .IN1(n11948), .IN2(n11925), .Q(n11947) );
  AND2X1 U11977 ( .IN1(n10826), .IN2(n10575), .Q(n11948) );
  AND2X1 U11978 ( .IN1(test_so3), .IN2(n11949), .Q(n11945) );
  OR2X1 U11979 ( .IN1(n10890), .IN2(n11950), .Q(n11949) );
  AND2X1 U11980 ( .IN1(n11951), .IN2(n11925), .Q(n11950) );
  AND2X1 U11981 ( .IN1(g4639), .IN2(n10551), .Q(n11951) );
  OR2X1 U11982 ( .IN1(n11952), .IN2(n11953), .Q(g34456) );
  AND2X1 U11983 ( .IN1(n11954), .IN2(g4616), .Q(n11953) );
  AND2X1 U11984 ( .IN1(n11955), .IN2(g4608), .Q(n11952) );
  OR2X1 U11985 ( .IN1(n10890), .IN2(n11956), .Q(n11955) );
  AND2X1 U11986 ( .IN1(n2590), .IN2(n11957), .Q(n11956) );
  OR2X1 U11987 ( .IN1(n11958), .IN2(n11959), .Q(g34455) );
  AND2X1 U11988 ( .IN1(n2595), .IN2(g4332), .Q(n11959) );
  AND2X1 U11989 ( .IN1(n11960), .IN2(g4322), .Q(n11958) );
  OR2X1 U11990 ( .IN1(n10890), .IN2(n11961), .Q(n11960) );
  AND2X1 U11991 ( .IN1(n11962), .IN2(n2594), .Q(n11961) );
  AND2X1 U11992 ( .IN1(n11963), .IN2(n11964), .Q(n11962) );
  OR2X1 U11993 ( .IN1(n11965), .IN2(n11966), .Q(g34454) );
  AND2X1 U11994 ( .IN1(n10919), .IN2(g4601), .Q(n11966) );
  AND2X1 U11995 ( .IN1(n11967), .IN2(n11954), .Q(n11965) );
  XNOR2X1 U11996 ( .IN1(n2590), .IN2(n5274), .Q(n11967) );
  OR2X1 U11997 ( .IN1(n11968), .IN2(n11969), .Q(g34453) );
  OR2X1 U11998 ( .IN1(n11970), .IN2(n11971), .Q(n11969) );
  AND2X1 U11999 ( .IN1(n11972), .IN2(n5365), .Q(n11971) );
  AND2X1 U12000 ( .IN1(n2598), .IN2(n11957), .Q(n11972) );
  AND2X1 U12001 ( .IN1(n11973), .IN2(g4601), .Q(n11970) );
  AND2X1 U12002 ( .IN1(n11954), .IN2(n11974), .Q(n11973) );
  INVX0 U12003 ( .INP(n2598), .ZN(n11974) );
  AND2X1 U12004 ( .IN1(n10919), .IN2(g4593), .Q(n11968) );
  OR2X1 U12005 ( .IN1(n11975), .IN2(n11976), .Q(g34452) );
  AND2X1 U12006 ( .IN1(n10919), .IN2(g4584), .Q(n11976) );
  AND2X1 U12007 ( .IN1(n11977), .IN2(n11954), .Q(n11975) );
  XNOR2X1 U12008 ( .IN1(n5303), .IN2(n108), .Q(n11977) );
  OR2X1 U12009 ( .IN1(n11978), .IN2(n11979), .Q(g34451) );
  AND2X1 U12010 ( .IN1(n10919), .IN2(g4332), .Q(n11979) );
  AND2X1 U12011 ( .IN1(n11980), .IN2(n11954), .Q(n11978) );
  AND2X1 U12012 ( .IN1(n10826), .IN2(n11957), .Q(n11954) );
  INVX0 U12013 ( .INP(n11981), .ZN(n11957) );
  OR2X1 U12014 ( .IN1(n11930), .IN2(n11982), .Q(n11981) );
  AND2X1 U12015 ( .IN1(n108), .IN2(g4616), .Q(n11982) );
  AND2X1 U12016 ( .IN1(g4584), .IN2(n11983), .Q(n108) );
  INVX0 U12017 ( .INP(n11963), .ZN(n11930) );
  XNOR2X1 U12018 ( .IN1(n5539), .IN2(n11983), .Q(n11980) );
  OR2X1 U12019 ( .IN1(n11984), .IN2(n11985), .Q(g34450) );
  OR2X1 U12020 ( .IN1(n11986), .IN2(n11987), .Q(n11985) );
  AND2X1 U12021 ( .IN1(n11988), .IN2(n5506), .Q(n11987) );
  AND2X1 U12022 ( .IN1(n2594), .IN2(n11963), .Q(n11988) );
  AND2X1 U12023 ( .IN1(n11989), .IN2(g4322), .Q(n11986) );
  AND2X1 U12024 ( .IN1(n2595), .IN2(n11990), .Q(n11989) );
  INVX0 U12025 ( .INP(n2594), .ZN(n11990) );
  AND2X1 U12026 ( .IN1(n11964), .IN2(n11991), .Q(n2595) );
  INVX0 U12027 ( .INP(n11983), .ZN(n11964) );
  AND2X1 U12028 ( .IN1(n2607), .IN2(n11992), .Q(n11983) );
  AND2X1 U12029 ( .IN1(g4332), .IN2(g4322), .Q(n11992) );
  AND2X1 U12030 ( .IN1(g4358), .IN2(n11993), .Q(n2607) );
  AND2X1 U12031 ( .IN1(n10919), .IN2(g4311), .Q(n11984) );
  OR2X1 U12032 ( .IN1(n11994), .IN2(n11995), .Q(g34448) );
  OR2X1 U12033 ( .IN1(n11996), .IN2(n11997), .Q(n11995) );
  AND2X1 U12034 ( .IN1(n10919), .IN2(g2827), .Q(n11997) );
  AND2X1 U12035 ( .IN1(n11998), .IN2(n10767), .Q(n11996) );
  AND2X1 U12036 ( .IN1(n11999), .IN2(g2819), .Q(n11998) );
  AND2X1 U12037 ( .IN1(n12000), .IN2(n12001), .Q(n11994) );
  AND2X1 U12038 ( .IN1(n12002), .IN2(n12003), .Q(n12000) );
  OR2X1 U12039 ( .IN1(n12004), .IN2(n12005), .Q(n12002) );
  AND2X1 U12040 ( .IN1(n10031), .IN2(n10767), .Q(n12004) );
  OR2X1 U12041 ( .IN1(n12006), .IN2(n12007), .Q(g34447) );
  OR2X1 U12042 ( .IN1(n12008), .IN2(n12009), .Q(n12007) );
  AND2X1 U12043 ( .IN1(n10920), .IN2(g2815), .Q(n12009) );
  AND2X1 U12044 ( .IN1(n12010), .IN2(n10767), .Q(n12008) );
  AND2X1 U12045 ( .IN1(n12011), .IN2(g2807), .Q(n12010) );
  AND2X1 U12046 ( .IN1(n12012), .IN2(n12013), .Q(n12006) );
  AND2X1 U12047 ( .IN1(n12014), .IN2(n12003), .Q(n12012) );
  OR2X1 U12048 ( .IN1(n12015), .IN2(n12005), .Q(n12014) );
  AND2X1 U12049 ( .IN1(n10030), .IN2(n10767), .Q(n12015) );
  OR2X1 U12050 ( .IN1(n12016), .IN2(n12017), .Q(g34446) );
  OR2X1 U12051 ( .IN1(n12018), .IN2(n12019), .Q(n12017) );
  AND2X1 U12052 ( .IN1(n10920), .IN2(g2819), .Q(n12019) );
  AND2X1 U12053 ( .IN1(n12020), .IN2(n10768), .Q(n12018) );
  AND2X1 U12054 ( .IN1(n12021), .IN2(g2815), .Q(n12020) );
  AND2X1 U12055 ( .IN1(n12022), .IN2(n12023), .Q(n12016) );
  AND2X1 U12056 ( .IN1(n12024), .IN2(n12003), .Q(n12022) );
  OR2X1 U12057 ( .IN1(n12025), .IN2(n12005), .Q(n12024) );
  AND2X1 U12058 ( .IN1(n10825), .IN2(n10584), .Q(n12025) );
  OR2X1 U12059 ( .IN1(n12026), .IN2(n12027), .Q(g34445) );
  OR2X1 U12060 ( .IN1(n12028), .IN2(n12029), .Q(n12027) );
  AND2X1 U12061 ( .IN1(n10920), .IN2(g2807), .Q(n12029) );
  AND2X1 U12062 ( .IN1(n12030), .IN2(n10768), .Q(n12028) );
  AND2X1 U12063 ( .IN1(n12031), .IN2(g2803), .Q(n12030) );
  AND2X1 U12064 ( .IN1(n12032), .IN2(n12033), .Q(n12026) );
  AND2X1 U12065 ( .IN1(n12034), .IN2(n12003), .Q(n12032) );
  OR2X1 U12066 ( .IN1(n1698), .IN2(n6005), .Q(n12003) );
  OR2X1 U12067 ( .IN1(n12035), .IN2(n12005), .Q(n12034) );
  AND2X1 U12068 ( .IN1(n10027), .IN2(n10768), .Q(n12035) );
  OR2X1 U12069 ( .IN1(n12036), .IN2(n12037), .Q(g34444) );
  OR2X1 U12070 ( .IN1(n12038), .IN2(n12039), .Q(n12037) );
  AND2X1 U12071 ( .IN1(n10920), .IN2(g2795), .Q(n12039) );
  AND2X1 U12072 ( .IN1(n12040), .IN2(n10768), .Q(n12038) );
  AND2X1 U12073 ( .IN1(n11999), .IN2(g2787), .Q(n12040) );
  AND2X1 U12074 ( .IN1(n12041), .IN2(n12001), .Q(n12036) );
  INVX0 U12075 ( .INP(n11999), .ZN(n12001) );
  OR2X1 U12076 ( .IN1(n12042), .IN2(n12043), .Q(n11999) );
  AND2X1 U12077 ( .IN1(n12044), .IN2(n12045), .Q(n12041) );
  OR2X1 U12078 ( .IN1(n12046), .IN2(n12005), .Q(n12044) );
  AND2X1 U12079 ( .IN1(n10028), .IN2(n10768), .Q(n12046) );
  OR2X1 U12080 ( .IN1(n12047), .IN2(n12048), .Q(g34443) );
  OR2X1 U12081 ( .IN1(n12049), .IN2(n12050), .Q(n12048) );
  AND2X1 U12082 ( .IN1(n10920), .IN2(g2783), .Q(n12050) );
  AND2X1 U12083 ( .IN1(n12051), .IN2(n10768), .Q(n12049) );
  AND2X1 U12084 ( .IN1(n12011), .IN2(g2775), .Q(n12051) );
  AND2X1 U12085 ( .IN1(n12052), .IN2(n12013), .Q(n12047) );
  INVX0 U12086 ( .INP(n12011), .ZN(n12013) );
  OR2X1 U12087 ( .IN1(n12043), .IN2(n12053), .Q(n12011) );
  OR2X1 U12088 ( .IN1(n5301), .IN2(g2729), .Q(n12053) );
  AND2X1 U12089 ( .IN1(n12054), .IN2(n12045), .Q(n12052) );
  OR2X1 U12090 ( .IN1(n12055), .IN2(n12005), .Q(n12054) );
  AND2X1 U12091 ( .IN1(n10026), .IN2(n10768), .Q(n12055) );
  OR2X1 U12092 ( .IN1(n12056), .IN2(n12057), .Q(g34442) );
  OR2X1 U12093 ( .IN1(n12058), .IN2(n12059), .Q(n12057) );
  AND2X1 U12094 ( .IN1(n10920), .IN2(g2787), .Q(n12059) );
  AND2X1 U12095 ( .IN1(n12060), .IN2(n10768), .Q(n12058) );
  AND2X1 U12096 ( .IN1(n12021), .IN2(g2783), .Q(n12060) );
  AND2X1 U12097 ( .IN1(n12061), .IN2(n12023), .Q(n12056) );
  INVX0 U12098 ( .INP(n12021), .ZN(n12023) );
  OR2X1 U12099 ( .IN1(n12043), .IN2(n12062), .Q(n12021) );
  AND2X1 U12100 ( .IN1(n12063), .IN2(n12045), .Q(n12061) );
  OR2X1 U12101 ( .IN1(n12064), .IN2(n12005), .Q(n12063) );
  AND2X1 U12102 ( .IN1(n10029), .IN2(n10768), .Q(n12064) );
  OR2X1 U12103 ( .IN1(n12065), .IN2(n12066), .Q(g34441) );
  OR2X1 U12104 ( .IN1(n12067), .IN2(n12068), .Q(n12066) );
  AND2X1 U12105 ( .IN1(n10920), .IN2(g2775), .Q(n12068) );
  AND2X1 U12106 ( .IN1(n12069), .IN2(n10769), .Q(n12067) );
  AND2X1 U12107 ( .IN1(n12031), .IN2(g2771), .Q(n12069) );
  INVX0 U12108 ( .INP(n12033), .ZN(n12031) );
  AND2X1 U12109 ( .IN1(n12070), .IN2(n12033), .Q(n12065) );
  AND2X1 U12110 ( .IN1(n12071), .IN2(n12072), .Q(n12033) );
  AND2X1 U12111 ( .IN1(n12073), .IN2(n12045), .Q(n12070) );
  OR2X1 U12112 ( .IN1(n1698), .IN2(n6006), .Q(n12045) );
  OR2X1 U12113 ( .IN1(n12074), .IN2(n12005), .Q(n12073) );
  AND2X1 U12114 ( .IN1(n10032), .IN2(n10769), .Q(n12074) );
  OR2X1 U12115 ( .IN1(n12075), .IN2(n12076), .Q(g34440) );
  AND2X1 U12116 ( .IN1(n12077), .IN2(n10769), .Q(n12076) );
  OR2X1 U12117 ( .IN1(n12078), .IN2(n12079), .Q(n12077) );
  AND2X1 U12118 ( .IN1(g890), .IN2(g896), .Q(n12079) );
  AND2X1 U12119 ( .IN1(n12080), .IN2(g862), .Q(n12078) );
  OR2X1 U12120 ( .IN1(n12081), .IN2(n5431), .Q(n12080) );
  AND2X1 U12121 ( .IN1(n12082), .IN2(n12083), .Q(n12081) );
  OR2X1 U12122 ( .IN1(g703), .IN2(n12084), .Q(n12082) );
  OR2X1 U12123 ( .IN1(n2644), .IN2(n12085), .Q(n12084) );
  AND2X1 U12124 ( .IN1(n10920), .IN2(g446), .Q(n12075) );
  OR2X1 U12125 ( .IN1(n12086), .IN2(n12087), .Q(g34439) );
  OR2X1 U12126 ( .IN1(n12088), .IN2(n12089), .Q(n12087) );
  AND2X1 U12127 ( .IN1(n2554), .IN2(n5330), .Q(n12089) );
  AND2X1 U12128 ( .IN1(n12090), .IN2(g776), .Q(n12088) );
  AND2X1 U12129 ( .IN1(n2404), .IN2(n12091), .Q(n12090) );
  INVX0 U12130 ( .INP(n2554), .ZN(n12091) );
  AND2X1 U12131 ( .IN1(n10920), .IN2(g772), .Q(n12086) );
  OR2X1 U12132 ( .IN1(n12092), .IN2(n12093), .Q(g34438) );
  OR2X1 U12133 ( .IN1(n12094), .IN2(n12095), .Q(n12093) );
  AND2X1 U12134 ( .IN1(n2556), .IN2(n5475), .Q(n12095) );
  AND2X1 U12135 ( .IN1(n12096), .IN2(g608), .Q(n12094) );
  AND2X1 U12136 ( .IN1(n2421), .IN2(n12097), .Q(n12096) );
  INVX0 U12137 ( .INP(n2556), .ZN(n12097) );
  AND2X1 U12138 ( .IN1(n10920), .IN2(g604), .Q(n12092) );
  AND2X1 U12139 ( .IN1(n12098), .IN2(n12099), .Q(g34435) );
  AND2X1 U12140 ( .IN1(n10497), .IN2(n12100), .Q(n12099) );
  OR2X1 U12141 ( .IN1(g4141), .IN2(n12101), .Q(n12100) );
  OR2X1 U12142 ( .IN1(n12102), .IN2(g4082), .Q(n12101) );
  AND2X1 U12143 ( .IN1(n12103), .IN2(n12104), .Q(n12102) );
  AND2X1 U12144 ( .IN1(n12105), .IN2(g4112), .Q(n12104) );
  AND2X1 U12145 ( .IN1(test_so11), .IN2(n5350), .Q(n12103) );
  AND2X1 U12146 ( .IN1(n5711), .IN2(n5416), .Q(n12098) );
  OR2X1 U12147 ( .IN1(n10537), .IN2(n11210), .Q(g34425) );
  OR2X1 U12148 ( .IN1(n12106), .IN2(n12107), .Q(n11210) );
  AND2X1 U12149 ( .IN1(n12108), .IN2(n12109), .Q(n12106) );
  OR2X1 U12150 ( .IN1(n12110), .IN2(n12111), .Q(n10537) );
  AND2X1 U12151 ( .IN1(n12112), .IN2(test_so81), .Q(n12111) );
  OR2X1 U12152 ( .IN1(n12113), .IN2(n12114), .Q(n12112) );
  AND2X1 U12153 ( .IN1(n12115), .IN2(g4358), .Q(n12114) );
  OR2X1 U12154 ( .IN1(n12116), .IN2(n12117), .Q(n12115) );
  AND2X1 U12155 ( .IN1(n12118), .IN2(n11739), .Q(n12117) );
  AND2X1 U12156 ( .IN1(n12119), .IN2(n11743), .Q(n12116) );
  AND2X1 U12157 ( .IN1(n5348), .IN2(n12120), .Q(n12113) );
  OR2X1 U12158 ( .IN1(n12121), .IN2(n12122), .Q(n12120) );
  AND2X1 U12159 ( .IN1(n12123), .IN2(n11739), .Q(n12122) );
  AND2X1 U12160 ( .IN1(n12124), .IN2(n11743), .Q(n12121) );
  AND2X1 U12161 ( .IN1(n12125), .IN2(n10552), .Q(n12110) );
  OR2X1 U12162 ( .IN1(n12126), .IN2(n12127), .Q(n12125) );
  AND2X1 U12163 ( .IN1(n12128), .IN2(g4358), .Q(n12127) );
  OR2X1 U12164 ( .IN1(n12129), .IN2(n12130), .Q(n12128) );
  AND2X1 U12165 ( .IN1(n12131), .IN2(n11739), .Q(n12130) );
  AND2X1 U12166 ( .IN1(n12132), .IN2(n11743), .Q(n12129) );
  AND2X1 U12167 ( .IN1(n5348), .IN2(n12133), .Q(n12126) );
  OR2X1 U12168 ( .IN1(n12134), .IN2(n12135), .Q(n12133) );
  AND2X1 U12169 ( .IN1(n11739), .IN2(n11096), .Q(n12135) );
  INVX0 U12170 ( .INP(n12108), .ZN(n11739) );
  AND2X1 U12171 ( .IN1(n11743), .IN2(g31860), .Q(n12134) );
  INVX0 U12172 ( .INP(n12109), .ZN(n11743) );
  OR2X1 U12173 ( .IN1(n12107), .IN2(n12136), .Q(g34383) );
  OR2X1 U12174 ( .IN1(g34843), .IN2(n12137), .Q(n12136) );
  AND2X1 U12175 ( .IN1(n12138), .IN2(n12139), .Q(n12137) );
  AND2X1 U12176 ( .IN1(n12140), .IN2(n12141), .Q(n12139) );
  AND2X1 U12177 ( .IN1(n3165), .IN2(n12142), .Q(n12141) );
  AND2X1 U12178 ( .IN1(n12143), .IN2(n3146), .Q(n12140) );
  AND2X1 U12179 ( .IN1(n12144), .IN2(n12145), .Q(n12138) );
  AND2X1 U12180 ( .IN1(n12146), .IN2(n12147), .Q(n12144) );
  OR2X1 U12181 ( .IN1(n12148), .IN2(n12149), .Q(g34843) );
  OR2X1 U12182 ( .IN1(n12150), .IN2(n12151), .Q(n12149) );
  OR2X1 U12183 ( .IN1(n12152), .IN2(n12153), .Q(n12151) );
  AND2X1 U12184 ( .IN1(g31862), .IN2(n12154), .Q(n12153) );
  INVX0 U12185 ( .INP(n12155), .ZN(n12152) );
  OR2X1 U12186 ( .IN1(n12156), .IN2(n12142), .Q(n12155) );
  OR2X1 U12187 ( .IN1(n12157), .IN2(n12158), .Q(n12150) );
  INVX0 U12188 ( .INP(n12159), .ZN(n12158) );
  OR2X1 U12189 ( .IN1(n12160), .IN2(n2727), .Q(n12159) );
  AND2X1 U12190 ( .IN1(n12161), .IN2(n12162), .Q(n12157) );
  OR2X1 U12191 ( .IN1(n12163), .IN2(n12164), .Q(n12148) );
  OR2X1 U12192 ( .IN1(n12165), .IN2(n12166), .Q(n12164) );
  AND2X1 U12193 ( .IN1(n12167), .IN2(n5524), .Q(n12166) );
  OR2X1 U12194 ( .IN1(n12168), .IN2(n12169), .Q(n12163) );
  OR2X1 U12195 ( .IN1(n12170), .IN2(n12171), .Q(g34269) );
  AND2X1 U12196 ( .IN1(n12172), .IN2(n10769), .Q(n12171) );
  OR2X1 U12197 ( .IN1(n12173), .IN2(n12174), .Q(n12172) );
  AND2X1 U12198 ( .IN1(n12175), .IN2(n12176), .Q(n12174) );
  OR2X1 U12199 ( .IN1(n12177), .IN2(n12178), .Q(n12176) );
  AND2X1 U12200 ( .IN1(n12179), .IN2(g4961), .Q(n12178) );
  INVX0 U12201 ( .INP(n12180), .ZN(n12173) );
  OR2X1 U12202 ( .IN1(n12175), .IN2(n5614), .Q(n12180) );
  OR2X1 U12203 ( .IN1(n12181), .IN2(n12182), .Q(n12175) );
  AND2X1 U12204 ( .IN1(n10920), .IN2(g4961), .Q(n12170) );
  OR2X1 U12205 ( .IN1(n12183), .IN2(n12184), .Q(g34268) );
  AND2X1 U12206 ( .IN1(n12185), .IN2(n10769), .Q(n12184) );
  OR2X1 U12207 ( .IN1(n12186), .IN2(n12187), .Q(n12185) );
  AND2X1 U12208 ( .IN1(n12188), .IN2(n12189), .Q(n12187) );
  OR2X1 U12209 ( .IN1(n12177), .IN2(n12190), .Q(n12189) );
  AND2X1 U12210 ( .IN1(n12179), .IN2(g4950), .Q(n12190) );
  INVX0 U12211 ( .INP(n12191), .ZN(n12186) );
  OR2X1 U12212 ( .IN1(n12188), .IN2(n5875), .Q(n12191) );
  OR2X1 U12213 ( .IN1(n12192), .IN2(n12182), .Q(n12188) );
  AND2X1 U12214 ( .IN1(n10920), .IN2(g4950), .Q(n12183) );
  OR2X1 U12215 ( .IN1(n12193), .IN2(n12194), .Q(g34267) );
  AND2X1 U12216 ( .IN1(n12195), .IN2(n10769), .Q(n12194) );
  OR2X1 U12217 ( .IN1(n12196), .IN2(n12197), .Q(n12195) );
  AND2X1 U12218 ( .IN1(n12198), .IN2(n12199), .Q(n12197) );
  AND2X1 U12219 ( .IN1(n12200), .IN2(n12179), .Q(n12198) );
  OR2X1 U12220 ( .IN1(n12177), .IN2(g4939), .Q(n12200) );
  INVX0 U12221 ( .INP(n12201), .ZN(n12196) );
  OR2X1 U12222 ( .IN1(n12199), .IN2(n5878), .Q(n12201) );
  OR2X1 U12223 ( .IN1(n12202), .IN2(n12182), .Q(n12199) );
  AND2X1 U12224 ( .IN1(n10920), .IN2(g4939), .Q(n12193) );
  OR2X1 U12225 ( .IN1(n12203), .IN2(n12204), .Q(g34266) );
  AND2X1 U12226 ( .IN1(n12205), .IN2(n10769), .Q(n12204) );
  OR2X1 U12227 ( .IN1(n12206), .IN2(n12207), .Q(n12205) );
  AND2X1 U12228 ( .IN1(n12208), .IN2(n12209), .Q(n12207) );
  OR2X1 U12229 ( .IN1(n12177), .IN2(n12210), .Q(n12209) );
  AND2X1 U12230 ( .IN1(n12179), .IN2(g4894), .Q(n12210) );
  OR2X1 U12231 ( .IN1(n12177), .IN2(n12211), .Q(n12179) );
  AND2X1 U12232 ( .IN1(g71), .IN2(n12182), .Q(n12177) );
  INVX0 U12233 ( .INP(n12212), .ZN(n12206) );
  OR2X1 U12234 ( .IN1(n12208), .IN2(n5863), .Q(n12212) );
  OR2X1 U12235 ( .IN1(n11738), .IN2(n12182), .Q(n12208) );
  INVX0 U12236 ( .INP(n12211), .ZN(n12182) );
  OR2X1 U12237 ( .IN1(g5008), .IN2(n12213), .Q(n12211) );
  OR2X1 U12238 ( .IN1(test_so46), .IN2(n12214), .Q(n12213) );
  AND2X1 U12239 ( .IN1(n10920), .IN2(g4894), .Q(n12203) );
  AND2X1 U12240 ( .IN1(n11883), .IN2(n11151), .Q(g34265) );
  AND2X1 U12241 ( .IN1(n5713), .IN2(n12215), .Q(n11151) );
  AND2X1 U12242 ( .IN1(n5318), .IN2(n5443), .Q(n12215) );
  AND2X1 U12243 ( .IN1(n10824), .IN2(n11886), .Q(n11883) );
  AND2X1 U12244 ( .IN1(n12216), .IN2(n12217), .Q(n11886) );
  OR2X1 U12245 ( .IN1(n12218), .IN2(n12219), .Q(g34264) );
  AND2X1 U12246 ( .IN1(n12220), .IN2(n10769), .Q(n12219) );
  OR2X1 U12247 ( .IN1(n12221), .IN2(n12222), .Q(n12220) );
  AND2X1 U12248 ( .IN1(n12223), .IN2(n12224), .Q(n12222) );
  OR2X1 U12249 ( .IN1(n12225), .IN2(n12226), .Q(n12224) );
  AND2X1 U12250 ( .IN1(n12227), .IN2(g4771), .Q(n12226) );
  INVX0 U12251 ( .INP(n12228), .ZN(n12221) );
  OR2X1 U12252 ( .IN1(n12223), .IN2(n5613), .Q(n12228) );
  OR2X1 U12253 ( .IN1(n12229), .IN2(n12230), .Q(n12223) );
  AND2X1 U12254 ( .IN1(n10920), .IN2(g4771), .Q(n12218) );
  OR2X1 U12255 ( .IN1(n12231), .IN2(n12232), .Q(g34263) );
  AND2X1 U12256 ( .IN1(n12233), .IN2(n10769), .Q(n12232) );
  OR2X1 U12257 ( .IN1(n12234), .IN2(n12235), .Q(n12233) );
  AND2X1 U12258 ( .IN1(n12236), .IN2(n12237), .Q(n12235) );
  OR2X1 U12259 ( .IN1(n12225), .IN2(n12238), .Q(n12237) );
  AND2X1 U12260 ( .IN1(n12227), .IN2(g4760), .Q(n12238) );
  INVX0 U12261 ( .INP(n12239), .ZN(n12234) );
  OR2X1 U12262 ( .IN1(n12236), .IN2(n5877), .Q(n12239) );
  OR2X1 U12263 ( .IN1(n12240), .IN2(n12230), .Q(n12236) );
  AND2X1 U12264 ( .IN1(n10920), .IN2(g4760), .Q(n12231) );
  OR2X1 U12265 ( .IN1(n12241), .IN2(n12242), .Q(g34262) );
  AND2X1 U12266 ( .IN1(n12243), .IN2(n10770), .Q(n12242) );
  OR2X1 U12267 ( .IN1(n12244), .IN2(n12245), .Q(n12243) );
  AND2X1 U12268 ( .IN1(n12246), .IN2(n12247), .Q(n12245) );
  AND2X1 U12269 ( .IN1(n12248), .IN2(n12227), .Q(n12246) );
  OR2X1 U12270 ( .IN1(n12225), .IN2(test_so18), .Q(n12248) );
  INVX0 U12271 ( .INP(n12249), .ZN(n12244) );
  OR2X1 U12272 ( .IN1(n12247), .IN2(n5876), .Q(n12249) );
  OR2X1 U12273 ( .IN1(n12250), .IN2(n12230), .Q(n12247) );
  AND2X1 U12274 ( .IN1(test_so18), .IN2(n10894), .Q(n12241) );
  OR2X1 U12275 ( .IN1(n12251), .IN2(n12252), .Q(g34261) );
  AND2X1 U12276 ( .IN1(n12253), .IN2(n10770), .Q(n12252) );
  OR2X1 U12277 ( .IN1(n12254), .IN2(n12255), .Q(n12253) );
  AND2X1 U12278 ( .IN1(n12256), .IN2(n12257), .Q(n12255) );
  OR2X1 U12279 ( .IN1(n12225), .IN2(n12258), .Q(n12257) );
  AND2X1 U12280 ( .IN1(n12227), .IN2(g4704), .Q(n12258) );
  OR2X1 U12281 ( .IN1(n12225), .IN2(n12259), .Q(n12227) );
  AND2X1 U12282 ( .IN1(g101), .IN2(n12230), .Q(n12225) );
  INVX0 U12283 ( .INP(n12260), .ZN(n12254) );
  OR2X1 U12284 ( .IN1(n12256), .IN2(n5862), .Q(n12260) );
  OR2X1 U12285 ( .IN1(n11742), .IN2(n12230), .Q(n12256) );
  INVX0 U12286 ( .INP(n12259), .ZN(n12230) );
  OR2X1 U12287 ( .IN1(g8132), .IN2(n12261), .Q(n12259) );
  OR2X1 U12288 ( .IN1(n12214), .IN2(g4818), .Q(n12261) );
  AND2X1 U12289 ( .IN1(n10920), .IN2(g4704), .Q(n12251) );
  AND2X1 U12290 ( .IN1(n11903), .IN2(n11115), .Q(g34260) );
  AND2X1 U12291 ( .IN1(n5712), .IN2(n12262), .Q(n11115) );
  AND2X1 U12292 ( .IN1(n10435), .IN2(n5440), .Q(n12262) );
  AND2X1 U12293 ( .IN1(n10824), .IN2(n11906), .Q(n11903) );
  AND2X1 U12294 ( .IN1(n12263), .IN2(n12264), .Q(n11906) );
  AND2X1 U12295 ( .IN1(n12265), .IN2(g4633), .Q(g34259) );
  OR2X1 U12296 ( .IN1(n10880), .IN2(n12266), .Q(n12265) );
  AND2X1 U12297 ( .IN1(n11925), .IN2(n11934), .Q(n12266) );
  OR2X1 U12298 ( .IN1(n12267), .IN2(n12268), .Q(g34258) );
  OR2X1 U12299 ( .IN1(n12269), .IN2(n12270), .Q(n12268) );
  AND2X1 U12300 ( .IN1(n12271), .IN2(n5348), .Q(n12270) );
  AND2X1 U12301 ( .IN1(n11993), .IN2(n11963), .Q(n12271) );
  AND2X1 U12302 ( .IN1(n12272), .IN2(g4358), .Q(n12269) );
  AND2X1 U12303 ( .IN1(n11991), .IN2(n12273), .Q(n12272) );
  INVX0 U12304 ( .INP(n11993), .ZN(n12273) );
  AND2X1 U12305 ( .IN1(n12274), .IN2(test_so81), .Q(n11993) );
  AND2X1 U12306 ( .IN1(test_so81), .IN2(n10894), .Q(n12267) );
  OR2X1 U12307 ( .IN1(n12275), .IN2(n12276), .Q(g34257) );
  OR2X1 U12308 ( .IN1(n12277), .IN2(n12278), .Q(n12276) );
  AND2X1 U12309 ( .IN1(n12279), .IN2(n12274), .Q(n12278) );
  INVX0 U12310 ( .INP(n11932), .ZN(n12274) );
  AND2X1 U12311 ( .IN1(n11963), .IN2(n10552), .Q(n12279) );
  AND2X1 U12312 ( .IN1(n12280), .IN2(n11932), .Q(n12277) );
  OR2X1 U12313 ( .IN1(n10551), .IN2(n12281), .Q(n11932) );
  OR2X1 U12314 ( .IN1(n5653), .IN2(n12282), .Q(n12281) );
  AND2X1 U12315 ( .IN1(n11991), .IN2(test_so81), .Q(n12280) );
  AND2X1 U12316 ( .IN1(n10824), .IN2(n11963), .Q(n11991) );
  AND2X1 U12317 ( .IN1(n10920), .IN2(g4340), .Q(n12275) );
  OR2X1 U12318 ( .IN1(n12283), .IN2(n12284), .Q(g34256) );
  AND2X1 U12319 ( .IN1(n12285), .IN2(n10770), .Q(n12284) );
  OR2X1 U12320 ( .IN1(g4459), .IN2(n12286), .Q(n12285) );
  OR2X1 U12321 ( .IN1(n12287), .IN2(n12288), .Q(n12286) );
  AND2X1 U12322 ( .IN1(n5671), .IN2(g4473), .Q(n12288) );
  AND2X1 U12323 ( .IN1(n10920), .IN2(g4369), .Q(n12283) );
  OR2X1 U12324 ( .IN1(n12289), .IN2(n12290), .Q(g34255) );
  OR2X1 U12325 ( .IN1(n12291), .IN2(g4462), .Q(n12290) );
  AND2X1 U12326 ( .IN1(test_so38), .IN2(g4473), .Q(n12291) );
  OR2X1 U12327 ( .IN1(n10878), .IN2(n12287), .Q(n12289) );
  OR2X1 U12328 ( .IN1(n12292), .IN2(n12293), .Q(g34254) );
  AND2X1 U12329 ( .IN1(n12287), .IN2(n10770), .Q(n12293) );
  AND2X1 U12330 ( .IN1(n12294), .IN2(g4473), .Q(n12292) );
  OR2X1 U12331 ( .IN1(n12295), .IN2(n12296), .Q(n12294) );
  OR2X1 U12332 ( .IN1(n5382), .IN2(n10874), .Q(n12296) );
  OR2X1 U12333 ( .IN1(test_so38), .IN2(n5671), .Q(n12295) );
  AND2X1 U12334 ( .IN1(n12297), .IN2(n10770), .Q(g34253) );
  OR2X1 U12335 ( .IN1(n10566), .IN2(n12298), .Q(n12297) );
  OR2X1 U12336 ( .IN1(n5671), .IN2(n12287), .Q(n12298) );
  AND2X1 U12337 ( .IN1(n5849), .IN2(n12299), .Q(n12287) );
  AND2X1 U12338 ( .IN1(g26960), .IN2(n12300), .Q(n12299) );
  OR2X1 U12339 ( .IN1(n11594), .IN2(n12301), .Q(n12300) );
  AND2X1 U12340 ( .IN1(n2668), .IN2(n5846), .Q(n12301) );
  OR2X1 U12341 ( .IN1(n12302), .IN2(n12303), .Q(g34252) );
  OR2X1 U12342 ( .IN1(n12304), .IN2(n12305), .Q(n12303) );
  AND2X1 U12343 ( .IN1(n2647), .IN2(n5334), .Q(n12305) );
  AND2X1 U12344 ( .IN1(n12306), .IN2(g772), .Q(n12304) );
  AND2X1 U12345 ( .IN1(n2404), .IN2(n12307), .Q(n12306) );
  INVX0 U12346 ( .INP(n2647), .ZN(n12307) );
  AND2X1 U12347 ( .IN1(n10921), .IN2(g767), .Q(n12302) );
  OR2X1 U12348 ( .IN1(n12308), .IN2(n12309), .Q(g34251) );
  OR2X1 U12349 ( .IN1(n12310), .IN2(n12311), .Q(n12309) );
  AND2X1 U12350 ( .IN1(n2649), .IN2(n5473), .Q(n12311) );
  AND2X1 U12351 ( .IN1(n12312), .IN2(g604), .Q(n12310) );
  AND2X1 U12352 ( .IN1(n2421), .IN2(n12313), .Q(n12312) );
  INVX0 U12353 ( .INP(n2649), .ZN(n12313) );
  AND2X1 U12354 ( .IN1(n10921), .IN2(g599), .Q(n12308) );
  OR2X1 U12355 ( .IN1(n12314), .IN2(n12315), .Q(g34250) );
  OR2X1 U12356 ( .IN1(n12316), .IN2(n12317), .Q(n12315) );
  AND2X1 U12357 ( .IN1(n5724), .IN2(n2707), .Q(n12317) );
  AND2X1 U12358 ( .IN1(n12318), .IN2(g142), .Q(n12316) );
  AND2X1 U12359 ( .IN1(n10534), .IN2(n12319), .Q(n12318) );
  INVX0 U12360 ( .INP(n2707), .ZN(n12319) );
  AND2X1 U12361 ( .IN1(n10921), .IN2(g298), .Q(n12314) );
  OR2X1 U12362 ( .IN1(n12320), .IN2(n12321), .Q(g34249) );
  OR2X1 U12363 ( .IN1(n12322), .IN2(n12323), .Q(n12321) );
  AND2X1 U12364 ( .IN1(n2710), .IN2(n5843), .Q(n12323) );
  AND2X1 U12365 ( .IN1(n12324), .IN2(g160), .Q(n12322) );
  INVX0 U12366 ( .INP(n12325), .ZN(n12324) );
  OR2X1 U12367 ( .IN1(n12326), .IN2(n2710), .Q(n12325) );
  AND2X1 U12368 ( .IN1(n10921), .IN2(g157), .Q(n12320) );
  OR2X1 U12369 ( .IN1(n12107), .IN2(n12327), .Q(g34201) );
  OR2X1 U12370 ( .IN1(g34781), .IN2(n12328), .Q(n12327) );
  AND2X1 U12371 ( .IN1(n12329), .IN2(n12330), .Q(n12328) );
  AND2X1 U12372 ( .IN1(n12331), .IN2(n12332), .Q(n12330) );
  AND2X1 U12373 ( .IN1(n3003), .IN2(n1645), .Q(n12332) );
  AND2X1 U12374 ( .IN1(n3588), .IN2(n3606), .Q(n12331) );
  AND2X1 U12375 ( .IN1(n12333), .IN2(n12334), .Q(n12329) );
  AND2X1 U12376 ( .IN1(n3550), .IN2(n3569), .Q(n12334) );
  AND2X1 U12377 ( .IN1(n3006), .IN2(n3007), .Q(n12333) );
  OR2X1 U12378 ( .IN1(n12335), .IN2(n12336), .Q(g34781) );
  OR2X1 U12379 ( .IN1(n12337), .IN2(n12338), .Q(n12336) );
  OR2X1 U12380 ( .IN1(n12339), .IN2(n12340), .Q(n12338) );
  AND2X1 U12381 ( .IN1(g25167), .IN2(n12341), .Q(n12340) );
  AND2X1 U12382 ( .IN1(n12342), .IN2(n5359), .Q(n12339) );
  AND2X1 U12383 ( .IN1(n3005), .IN2(g1783), .Q(n12342) );
  OR2X1 U12384 ( .IN1(n12343), .IN2(n12344), .Q(n12337) );
  AND2X1 U12385 ( .IN1(n12345), .IN2(n5510), .Q(n12344) );
  AND2X1 U12386 ( .IN1(n12346), .IN2(g1917), .Q(n12345) );
  AND2X1 U12387 ( .IN1(n12347), .IN2(n5507), .Q(n12343) );
  AND2X1 U12388 ( .IN1(n12348), .IN2(g2051), .Q(n12347) );
  OR2X1 U12389 ( .IN1(n12349), .IN2(n12350), .Q(n12335) );
  OR2X1 U12390 ( .IN1(n12351), .IN2(n12352), .Q(n12350) );
  AND2X1 U12391 ( .IN1(n12353), .IN2(n5512), .Q(n12352) );
  AND2X1 U12392 ( .IN1(n12354), .IN2(g2208), .Q(n12353) );
  AND2X1 U12393 ( .IN1(n12355), .IN2(n5511), .Q(n12351) );
  AND2X1 U12394 ( .IN1(test_so21), .IN2(n12356), .Q(n12355) );
  OR2X1 U12395 ( .IN1(n12357), .IN2(n12358), .Q(n12349) );
  AND2X1 U12396 ( .IN1(n12359), .IN2(n5509), .Q(n12358) );
  AND2X1 U12397 ( .IN1(n12360), .IN2(g2476), .Q(n12359) );
  AND2X1 U12398 ( .IN1(n12361), .IN2(n5508), .Q(n12357) );
  AND2X1 U12399 ( .IN1(n12362), .IN2(g2610), .Q(n12361) );
  OR2X1 U12400 ( .IN1(n12363), .IN2(n12364), .Q(g34041) );
  AND2X1 U12401 ( .IN1(n10921), .IN2(g5008), .Q(n12364) );
  AND2X1 U12402 ( .IN1(n12365), .IN2(n12366), .Q(n12363) );
  XNOR2X1 U12403 ( .IN1(n11737), .IN2(n5367), .Q(n12365) );
  OR2X1 U12404 ( .IN1(n12367), .IN2(n12368), .Q(g34040) );
  OR2X1 U12405 ( .IN1(n12369), .IN2(n12370), .Q(n12368) );
  AND2X1 U12406 ( .IN1(n12366), .IN2(g4899), .Q(n12370) );
  AND2X1 U12407 ( .IN1(n12371), .IN2(n12217), .Q(n12369) );
  OR2X1 U12408 ( .IN1(n12372), .IN2(n12373), .Q(n12371) );
  AND2X1 U12409 ( .IN1(n11165), .IN2(n10770), .Q(n12373) );
  AND2X1 U12410 ( .IN1(n12374), .IN2(n11164), .Q(n12372) );
  AND2X1 U12411 ( .IN1(n10921), .IN2(g4975), .Q(n12367) );
  OR2X1 U12412 ( .IN1(n12375), .IN2(n12376), .Q(g34039) );
  AND2X1 U12413 ( .IN1(n12366), .IN2(g4966), .Q(n12376) );
  AND2X1 U12414 ( .IN1(test_so58), .IN2(n12377), .Q(n12375) );
  OR2X1 U12415 ( .IN1(n10877), .IN2(n12378), .Q(n12377) );
  OR2X1 U12416 ( .IN1(n12379), .IN2(n12380), .Q(g34038) );
  OR2X1 U12417 ( .IN1(n12381), .IN2(n12382), .Q(n12380) );
  AND2X1 U12418 ( .IN1(n12383), .IN2(test_so58), .Q(n12382) );
  AND2X1 U12419 ( .IN1(n12366), .IN2(n12384), .Q(n12383) );
  INVX0 U12420 ( .INP(n12385), .ZN(n12384) );
  AND2X1 U12421 ( .IN1(n12378), .IN2(n10560), .Q(n12381) );
  AND2X1 U12422 ( .IN1(n12386), .IN2(n12385), .Q(n12378) );
  AND2X1 U12423 ( .IN1(n10921), .IN2(g4983), .Q(n12379) );
  OR2X1 U12424 ( .IN1(n12387), .IN2(n12388), .Q(g34037) );
  OR2X1 U12425 ( .IN1(n12389), .IN2(n12390), .Q(n12388) );
  AND2X1 U12426 ( .IN1(n12391), .IN2(n5360), .Q(n12390) );
  AND2X1 U12427 ( .IN1(n12374), .IN2(n12217), .Q(n12391) );
  AND2X1 U12428 ( .IN1(n12366), .IN2(g4975), .Q(n12389) );
  AND2X1 U12429 ( .IN1(n10823), .IN2(n12386), .Q(n12366) );
  AND2X1 U12430 ( .IN1(n12217), .IN2(n12392), .Q(n12386) );
  INVX0 U12431 ( .INP(n12374), .ZN(n12392) );
  AND2X1 U12432 ( .IN1(g4966), .IN2(n12385), .Q(n12374) );
  AND2X1 U12433 ( .IN1(g4983), .IN2(n11737), .Q(n12385) );
  INVX0 U12434 ( .INP(n12216), .ZN(n11737) );
  OR2X1 U12435 ( .IN1(n5283), .IN2(n12393), .Q(n12216) );
  AND2X1 U12436 ( .IN1(n10921), .IN2(g4966), .Q(n12387) );
  AND2X1 U12437 ( .IN1(n12394), .IN2(g4871), .Q(g34036) );
  AND2X1 U12438 ( .IN1(n12394), .IN2(g4864), .Q(g34035) );
  AND2X1 U12439 ( .IN1(n12394), .IN2(g4836), .Q(g34034) );
  OR2X1 U12440 ( .IN1(n10879), .IN2(n12217), .Q(n12394) );
  OR2X1 U12441 ( .IN1(n12108), .IN2(n12395), .Q(n12217) );
  OR2X1 U12442 ( .IN1(n12396), .IN2(n12397), .Q(g34033) );
  AND2X1 U12443 ( .IN1(n10921), .IN2(g4818), .Q(n12397) );
  AND2X1 U12444 ( .IN1(n12398), .IN2(n12399), .Q(n12396) );
  XNOR2X1 U12445 ( .IN1(n11741), .IN2(n5368), .Q(n12398) );
  OR2X1 U12446 ( .IN1(n12400), .IN2(n12401), .Q(g34032) );
  OR2X1 U12447 ( .IN1(n12402), .IN2(n12403), .Q(n12401) );
  AND2X1 U12448 ( .IN1(n12399), .IN2(g4709), .Q(n12403) );
  AND2X1 U12449 ( .IN1(n12404), .IN2(n12263), .Q(n12402) );
  OR2X1 U12450 ( .IN1(n12405), .IN2(n12406), .Q(n12404) );
  AND2X1 U12451 ( .IN1(n11133), .IN2(n10770), .Q(n12406) );
  AND2X1 U12452 ( .IN1(n12407), .IN2(n11132), .Q(n12405) );
  AND2X1 U12453 ( .IN1(n10921), .IN2(g4785), .Q(n12400) );
  OR2X1 U12454 ( .IN1(n12408), .IN2(n12409), .Q(g34031) );
  AND2X1 U12455 ( .IN1(n12399), .IN2(g4776), .Q(n12409) );
  AND2X1 U12456 ( .IN1(test_so29), .IN2(n12410), .Q(n12408) );
  OR2X1 U12457 ( .IN1(n10878), .IN2(n12411), .Q(n12410) );
  OR2X1 U12458 ( .IN1(n12412), .IN2(n12413), .Q(g34030) );
  OR2X1 U12459 ( .IN1(n12414), .IN2(n12415), .Q(n12413) );
  AND2X1 U12460 ( .IN1(n12416), .IN2(test_so29), .Q(n12415) );
  AND2X1 U12461 ( .IN1(n12399), .IN2(n12417), .Q(n12416) );
  AND2X1 U12462 ( .IN1(n12411), .IN2(n10561), .Q(n12414) );
  AND2X1 U12463 ( .IN1(n12418), .IN2(n12419), .Q(n12411) );
  AND2X1 U12464 ( .IN1(n10921), .IN2(g4793), .Q(n12412) );
  OR2X1 U12465 ( .IN1(n12420), .IN2(n12421), .Q(g34029) );
  OR2X1 U12466 ( .IN1(n12422), .IN2(n12423), .Q(n12421) );
  AND2X1 U12467 ( .IN1(n12424), .IN2(n5361), .Q(n12423) );
  AND2X1 U12468 ( .IN1(n12407), .IN2(n12263), .Q(n12424) );
  INVX0 U12469 ( .INP(n12425), .ZN(n12407) );
  AND2X1 U12470 ( .IN1(n12399), .IN2(g4785), .Q(n12422) );
  AND2X1 U12471 ( .IN1(n10823), .IN2(n12418), .Q(n12399) );
  AND2X1 U12472 ( .IN1(n12425), .IN2(n12263), .Q(n12418) );
  OR2X1 U12473 ( .IN1(n5707), .IN2(n12417), .Q(n12425) );
  INVX0 U12474 ( .INP(n12419), .ZN(n12417) );
  AND2X1 U12475 ( .IN1(g4793), .IN2(n11741), .Q(n12419) );
  INVX0 U12476 ( .INP(n12264), .ZN(n11741) );
  OR2X1 U12477 ( .IN1(n5656), .IN2(n12426), .Q(n12264) );
  AND2X1 U12478 ( .IN1(n10913), .IN2(g4776), .Q(n12420) );
  AND2X1 U12479 ( .IN1(n11209), .IN2(g4674), .Q(g34027) );
  AND2X1 U12480 ( .IN1(n11209), .IN2(g4646), .Q(g34026) );
  OR2X1 U12481 ( .IN1(n10879), .IN2(n12263), .Q(n11209) );
  OR2X1 U12482 ( .IN1(n12109), .IN2(n12395), .Q(n12263) );
  OR2X1 U12483 ( .IN1(n10131), .IN2(n1698), .Q(n12395) );
  AND2X1 U12484 ( .IN1(n11925), .IN2(n12427), .Q(g34025) );
  AND2X1 U12485 ( .IN1(n10823), .IN2(n5727), .Q(n12427) );
  AND2X1 U12486 ( .IN1(n11963), .IN2(n5382), .Q(n11925) );
  OR2X1 U12487 ( .IN1(n12428), .IN2(DFF_961_n1), .Q(n11963) );
  AND2X1 U12488 ( .IN1(n12429), .IN2(n1698), .Q(n12428) );
  OR2X1 U12489 ( .IN1(n12430), .IN2(n12431), .Q(g34024) );
  AND2X1 U12490 ( .IN1(n12432), .IN2(n10770), .Q(n12431) );
  AND2X1 U12491 ( .IN1(n12433), .IN2(n12434), .Q(n12432) );
  OR2X1 U12492 ( .IN1(n12435), .IN2(n12436), .Q(n12434) );
  OR2X1 U12493 ( .IN1(n12429), .IN2(n12437), .Q(n12433) );
  AND2X1 U12494 ( .IN1(n10910), .IN2(g4492), .Q(n12430) );
  OR2X1 U12495 ( .IN1(n12438), .IN2(n12439), .Q(g34023) );
  AND2X1 U12496 ( .IN1(n12440), .IN2(n9325), .Q(n12439) );
  OR2X1 U12497 ( .IN1(n10880), .IN2(n12441), .Q(n12440) );
  AND2X1 U12498 ( .IN1(n12442), .IN2(n12443), .Q(n12441) );
  AND2X1 U12499 ( .IN1(g4558), .IN2(g4561), .Q(n12443) );
  AND2X1 U12500 ( .IN1(n12444), .IN2(g4555), .Q(n12442) );
  AND2X1 U12501 ( .IN1(n12445), .IN2(n12444), .Q(n12438) );
  OR2X1 U12502 ( .IN1(n12429), .IN2(n12446), .Q(n12444) );
  AND2X1 U12503 ( .IN1(n12436), .IN2(n10770), .Q(n12445) );
  OR2X1 U12504 ( .IN1(n11594), .IN2(g2988), .Q(n12436) );
  OR2X1 U12505 ( .IN1(n12447), .IN2(n12448), .Q(g34022) );
  OR2X1 U12506 ( .IN1(n2787), .IN2(n12449), .Q(n12448) );
  INVX0 U12507 ( .INP(n12450), .ZN(n12449) );
  OR2X1 U12508 ( .IN1(n12451), .IN2(g2763), .Q(n12450) );
  OR2X1 U12509 ( .IN1(n12452), .IN2(n12453), .Q(n12447) );
  AND2X1 U12510 ( .IN1(n10910), .IN2(g2759), .Q(n12453) );
  AND2X1 U12511 ( .IN1(n12454), .IN2(n10771), .Q(n12452) );
  AND2X1 U12512 ( .IN1(n12451), .IN2(g2763), .Q(n12454) );
  OR2X1 U12513 ( .IN1(n10530), .IN2(n12455), .Q(n12451) );
  OR2X1 U12514 ( .IN1(n12456), .IN2(n12457), .Q(g34021) );
  OR2X1 U12515 ( .IN1(n12458), .IN2(n12459), .Q(n12457) );
  AND2X1 U12516 ( .IN1(n12460), .IN2(g2567), .Q(n12459) );
  AND2X1 U12517 ( .IN1(n12461), .IN2(n12462), .Q(n12458) );
  AND2X1 U12518 ( .IN1(n10910), .IN2(g2648), .Q(n12456) );
  OR2X1 U12519 ( .IN1(n12463), .IN2(n12464), .Q(g34020) );
  AND2X1 U12520 ( .IN1(n12465), .IN2(n10771), .Q(n12464) );
  OR2X1 U12521 ( .IN1(n12466), .IN2(n12467), .Q(n12465) );
  AND2X1 U12522 ( .IN1(n12468), .IN2(g2643), .Q(n12467) );
  OR2X1 U12523 ( .IN1(n12469), .IN2(n12470), .Q(n12468) );
  AND2X1 U12524 ( .IN1(n12471), .IN2(g2555), .Q(n12469) );
  AND2X1 U12525 ( .IN1(n12472), .IN2(n12473), .Q(n12466) );
  INVX0 U12526 ( .INP(n12471), .ZN(n12473) );
  OR2X1 U12527 ( .IN1(n12474), .IN2(n12461), .Q(n12472) );
  AND2X1 U12528 ( .IN1(n10095), .IN2(n12475), .Q(n12474) );
  AND2X1 U12529 ( .IN1(n12476), .IN2(g2629), .Q(n12463) );
  OR2X1 U12530 ( .IN1(n10879), .IN2(n12477), .Q(n12476) );
  AND2X1 U12531 ( .IN1(n12471), .IN2(g2643), .Q(n12477) );
  AND2X1 U12532 ( .IN1(n12478), .IN2(n12479), .Q(n12471) );
  OR2X1 U12533 ( .IN1(g1589), .IN2(n12480), .Q(n12479) );
  OR2X1 U12534 ( .IN1(n12481), .IN2(n12482), .Q(g34019) );
  OR2X1 U12535 ( .IN1(n12483), .IN2(n12484), .Q(n12482) );
  AND2X1 U12536 ( .IN1(n10910), .IN2(g2571), .Q(n12484) );
  AND2X1 U12537 ( .IN1(n12485), .IN2(n10771), .Q(n12483) );
  AND2X1 U12538 ( .IN1(n12486), .IN2(g2583), .Q(n12485) );
  INVX0 U12539 ( .INP(n12487), .ZN(n12486) );
  AND2X1 U12540 ( .IN1(n12487), .IN2(n12462), .Q(n12481) );
  AND2X1 U12541 ( .IN1(g2629), .IN2(n12488), .Q(n12487) );
  OR2X1 U12542 ( .IN1(n12489), .IN2(n12490), .Q(g34018) );
  OR2X1 U12543 ( .IN1(n12491), .IN2(n12492), .Q(n12490) );
  AND2X1 U12544 ( .IN1(n10910), .IN2(g2583), .Q(n12492) );
  AND2X1 U12545 ( .IN1(n12493), .IN2(n10771), .Q(n12491) );
  AND2X1 U12546 ( .IN1(test_so61), .IN2(n12494), .Q(n12493) );
  INVX0 U12547 ( .INP(n12495), .ZN(n12494) );
  AND2X1 U12548 ( .IN1(n12495), .IN2(n12462), .Q(n12489) );
  AND2X1 U12549 ( .IN1(n5351), .IN2(n12496), .Q(n12495) );
  OR2X1 U12550 ( .IN1(n12497), .IN2(n12498), .Q(g34017) );
  OR2X1 U12551 ( .IN1(n12499), .IN2(n12500), .Q(n12498) );
  AND2X1 U12552 ( .IN1(test_so61), .IN2(n10895), .Q(n12500) );
  AND2X1 U12553 ( .IN1(n12501), .IN2(n10771), .Q(n12499) );
  AND2X1 U12554 ( .IN1(test_so66), .IN2(n12502), .Q(n12501) );
  AND2X1 U12555 ( .IN1(n12503), .IN2(n12462), .Q(n12497) );
  INVX0 U12556 ( .INP(n12502), .ZN(n12503) );
  OR2X1 U12557 ( .IN1(n12470), .IN2(n12504), .Q(n12502) );
  OR2X1 U12558 ( .IN1(n5521), .IN2(n5351), .Q(n12504) );
  OR2X1 U12559 ( .IN1(n12505), .IN2(n12506), .Q(g34016) );
  OR2X1 U12560 ( .IN1(n12507), .IN2(n12508), .Q(n12506) );
  AND2X1 U12561 ( .IN1(n10911), .IN2(g2563), .Q(n12508) );
  AND2X1 U12562 ( .IN1(n12509), .IN2(n10771), .Q(n12507) );
  AND2X1 U12563 ( .IN1(n12510), .IN2(g2571), .Q(n12509) );
  INVX0 U12564 ( .INP(n12511), .ZN(n12510) );
  AND2X1 U12565 ( .IN1(n12511), .IN2(n12462), .Q(n12505) );
  AND2X1 U12566 ( .IN1(n5521), .IN2(n12496), .Q(n12511) );
  OR2X1 U12567 ( .IN1(n12512), .IN2(n12513), .Q(g34015) );
  OR2X1 U12568 ( .IN1(n12514), .IN2(n12515), .Q(n12513) );
  AND2X1 U12569 ( .IN1(n10911), .IN2(g2567), .Q(n12515) );
  AND2X1 U12570 ( .IN1(n12516), .IN2(n10771), .Q(n12514) );
  AND2X1 U12571 ( .IN1(n12517), .IN2(g2563), .Q(n12516) );
  INVX0 U12572 ( .INP(n12518), .ZN(n12517) );
  AND2X1 U12573 ( .IN1(n12518), .IN2(n12462), .Q(n12512) );
  INVX0 U12574 ( .INP(n12519), .ZN(n12462) );
  OR2X1 U12575 ( .IN1(n10879), .IN2(n12520), .Q(n12519) );
  AND2X1 U12576 ( .IN1(n12521), .IN2(n12478), .Q(n12520) );
  OR2X1 U12577 ( .IN1(n12522), .IN2(n12523), .Q(n12478) );
  OR2X1 U12578 ( .IN1(n12524), .IN2(n12525), .Q(n12523) );
  INVX0 U12579 ( .INP(n12480), .ZN(n12525) );
  AND2X1 U12580 ( .IN1(n5483), .IN2(n12526), .Q(n12522) );
  OR2X1 U12581 ( .IN1(n12480), .IN2(g1585), .Q(n12521) );
  AND2X1 U12582 ( .IN1(g2555), .IN2(n12488), .Q(n12518) );
  OR2X1 U12583 ( .IN1(n12527), .IN2(n12528), .Q(g34014) );
  OR2X1 U12584 ( .IN1(n12529), .IN2(n12530), .Q(n12528) );
  AND2X1 U12585 ( .IN1(n12531), .IN2(g2433), .Q(n12530) );
  AND2X1 U12586 ( .IN1(n12532), .IN2(n12533), .Q(n12529) );
  AND2X1 U12587 ( .IN1(n10911), .IN2(g2514), .Q(n12527) );
  OR2X1 U12588 ( .IN1(n12534), .IN2(n12535), .Q(g34013) );
  AND2X1 U12589 ( .IN1(n12536), .IN2(n10771), .Q(n12535) );
  OR2X1 U12590 ( .IN1(n12537), .IN2(n12538), .Q(n12536) );
  AND2X1 U12591 ( .IN1(n12539), .IN2(g2509), .Q(n12538) );
  OR2X1 U12592 ( .IN1(n12540), .IN2(n12541), .Q(n12539) );
  AND2X1 U12593 ( .IN1(test_so79), .IN2(n12542), .Q(n12540) );
  AND2X1 U12594 ( .IN1(n12543), .IN2(n12544), .Q(n12537) );
  INVX0 U12595 ( .INP(n12542), .ZN(n12544) );
  OR2X1 U12596 ( .IN1(n12545), .IN2(n12532), .Q(n12543) );
  AND2X1 U12597 ( .IN1(n10094), .IN2(n12546), .Q(n12545) );
  AND2X1 U12598 ( .IN1(n12547), .IN2(g2495), .Q(n12534) );
  OR2X1 U12599 ( .IN1(n10880), .IN2(n12548), .Q(n12547) );
  AND2X1 U12600 ( .IN1(n12542), .IN2(g2509), .Q(n12548) );
  AND2X1 U12601 ( .IN1(n12549), .IN2(n12550), .Q(n12542) );
  OR2X1 U12602 ( .IN1(n12551), .IN2(n5755), .Q(n12550) );
  OR2X1 U12603 ( .IN1(n12552), .IN2(n12553), .Q(g34012) );
  OR2X1 U12604 ( .IN1(n12554), .IN2(n12555), .Q(n12553) );
  AND2X1 U12605 ( .IN1(n10911), .IN2(g2437), .Q(n12555) );
  AND2X1 U12606 ( .IN1(n12556), .IN2(n10772), .Q(n12554) );
  AND2X1 U12607 ( .IN1(n12557), .IN2(g2449), .Q(n12556) );
  AND2X1 U12608 ( .IN1(n12558), .IN2(n12533), .Q(n12552) );
  INVX0 U12609 ( .INP(n12557), .ZN(n12558) );
  OR2X1 U12610 ( .IN1(n12541), .IN2(n12160), .Q(n12557) );
  OR2X1 U12611 ( .IN1(n12559), .IN2(n12560), .Q(g34011) );
  OR2X1 U12612 ( .IN1(n12561), .IN2(n12562), .Q(n12560) );
  AND2X1 U12613 ( .IN1(n10911), .IN2(g2449), .Q(n12562) );
  AND2X1 U12614 ( .IN1(n12563), .IN2(n10772), .Q(n12561) );
  AND2X1 U12615 ( .IN1(n12564), .IN2(n9274), .Q(n12563) );
  INVX0 U12616 ( .INP(n12565), .ZN(n12564) );
  AND2X1 U12617 ( .IN1(n12565), .IN2(n12533), .Q(n12559) );
  AND2X1 U12618 ( .IN1(n10569), .IN2(n12566), .Q(n12565) );
  OR2X1 U12619 ( .IN1(n12567), .IN2(n12568), .Q(g34010) );
  OR2X1 U12620 ( .IN1(n12569), .IN2(n12570), .Q(n12568) );
  AND2X1 U12621 ( .IN1(n10911), .IN2(n9274), .Q(n12570) );
  AND2X1 U12622 ( .IN1(n12571), .IN2(n10772), .Q(n12569) );
  AND2X1 U12623 ( .IN1(n12572), .IN2(g2441), .Q(n12571) );
  INVX0 U12624 ( .INP(n12573), .ZN(n12572) );
  AND2X1 U12625 ( .IN1(n12573), .IN2(n12533), .Q(n12567) );
  AND2X1 U12626 ( .IN1(g2495), .IN2(n12574), .Q(n12573) );
  OR2X1 U12627 ( .IN1(n12575), .IN2(n12576), .Q(g34009) );
  OR2X1 U12628 ( .IN1(n12577), .IN2(n12578), .Q(n12576) );
  AND2X1 U12629 ( .IN1(n10911), .IN2(g2429), .Q(n12578) );
  AND2X1 U12630 ( .IN1(n12579), .IN2(n10772), .Q(n12577) );
  AND2X1 U12631 ( .IN1(n12580), .IN2(g2437), .Q(n12579) );
  INVX0 U12632 ( .INP(n12581), .ZN(n12580) );
  AND2X1 U12633 ( .IN1(n12581), .IN2(n12533), .Q(n12575) );
  AND2X1 U12634 ( .IN1(n5522), .IN2(n12566), .Q(n12581) );
  OR2X1 U12635 ( .IN1(n12582), .IN2(n12583), .Q(g34008) );
  OR2X1 U12636 ( .IN1(n12584), .IN2(n12585), .Q(n12583) );
  AND2X1 U12637 ( .IN1(n10911), .IN2(g2433), .Q(n12585) );
  AND2X1 U12638 ( .IN1(n12586), .IN2(n10772), .Q(n12584) );
  AND2X1 U12639 ( .IN1(n12587), .IN2(g2429), .Q(n12586) );
  INVX0 U12640 ( .INP(n12588), .ZN(n12587) );
  AND2X1 U12641 ( .IN1(n12588), .IN2(n12533), .Q(n12582) );
  AND2X1 U12642 ( .IN1(n10822), .IN2(n12589), .Q(n12533) );
  INVX0 U12643 ( .INP(n12590), .ZN(n12589) );
  AND2X1 U12644 ( .IN1(n12591), .IN2(n12549), .Q(n12590) );
  OR2X1 U12645 ( .IN1(n12592), .IN2(n12593), .Q(n12549) );
  OR2X1 U12646 ( .IN1(n12524), .IN2(n12594), .Q(n12593) );
  AND2X1 U12647 ( .IN1(n5290), .IN2(n12526), .Q(n12592) );
  OR2X1 U12648 ( .IN1(n5757), .IN2(n12551), .Q(n12591) );
  AND2X1 U12649 ( .IN1(n5523), .IN2(n12574), .Q(n12588) );
  OR2X1 U12650 ( .IN1(n12595), .IN2(n12596), .Q(g34007) );
  OR2X1 U12651 ( .IN1(n12597), .IN2(n12598), .Q(n12596) );
  AND2X1 U12652 ( .IN1(n12599), .IN2(g2299), .Q(n12598) );
  AND2X1 U12653 ( .IN1(n12600), .IN2(n12601), .Q(n12597) );
  AND2X1 U12654 ( .IN1(n10911), .IN2(g2380), .Q(n12595) );
  OR2X1 U12655 ( .IN1(n12602), .IN2(n12603), .Q(g34006) );
  AND2X1 U12656 ( .IN1(n12604), .IN2(n10772), .Q(n12603) );
  OR2X1 U12657 ( .IN1(n12605), .IN2(n12606), .Q(n12604) );
  AND2X1 U12658 ( .IN1(n12607), .IN2(g2375), .Q(n12606) );
  OR2X1 U12659 ( .IN1(n12608), .IN2(n12609), .Q(n12607) );
  AND2X1 U12660 ( .IN1(n12610), .IN2(g2287), .Q(n12608) );
  AND2X1 U12661 ( .IN1(n12611), .IN2(n12612), .Q(n12605) );
  INVX0 U12662 ( .INP(n12610), .ZN(n12612) );
  OR2X1 U12663 ( .IN1(n12613), .IN2(n12600), .Q(n12611) );
  AND2X1 U12664 ( .IN1(n10096), .IN2(n12614), .Q(n12613) );
  AND2X1 U12665 ( .IN1(n12615), .IN2(g2361), .Q(n12602) );
  OR2X1 U12666 ( .IN1(n10880), .IN2(n12616), .Q(n12615) );
  AND2X1 U12667 ( .IN1(n12610), .IN2(g2375), .Q(n12616) );
  AND2X1 U12668 ( .IN1(n12617), .IN2(n12618), .Q(n12610) );
  OR2X1 U12669 ( .IN1(n12619), .IN2(g1589), .Q(n12618) );
  OR2X1 U12670 ( .IN1(n12620), .IN2(n12621), .Q(g34005) );
  OR2X1 U12671 ( .IN1(n12622), .IN2(n12623), .Q(n12621) );
  AND2X1 U12672 ( .IN1(n10911), .IN2(g2303), .Q(n12623) );
  AND2X1 U12673 ( .IN1(n12624), .IN2(n10772), .Q(n12622) );
  AND2X1 U12674 ( .IN1(n12625), .IN2(g2315), .Q(n12624) );
  AND2X1 U12675 ( .IN1(n12626), .IN2(n12601), .Q(n12620) );
  INVX0 U12676 ( .INP(n12625), .ZN(n12626) );
  OR2X1 U12677 ( .IN1(g2331), .IN2(n12627), .Q(n12625) );
  OR2X1 U12678 ( .IN1(n12628), .IN2(n12629), .Q(g34004) );
  OR2X1 U12679 ( .IN1(n12630), .IN2(n12631), .Q(n12629) );
  AND2X1 U12680 ( .IN1(n10911), .IN2(g2315), .Q(n12631) );
  AND2X1 U12681 ( .IN1(n12632), .IN2(n10772), .Q(n12630) );
  AND2X1 U12682 ( .IN1(n12633), .IN2(n9314), .Q(n12632) );
  INVX0 U12683 ( .INP(n12634), .ZN(n12633) );
  AND2X1 U12684 ( .IN1(n12634), .IN2(n12601), .Q(n12628) );
  AND2X1 U12685 ( .IN1(n5353), .IN2(n12635), .Q(n12634) );
  OR2X1 U12686 ( .IN1(n12636), .IN2(n12637), .Q(g34003) );
  OR2X1 U12687 ( .IN1(n12638), .IN2(n12639), .Q(n12637) );
  AND2X1 U12688 ( .IN1(n10911), .IN2(n9314), .Q(n12639) );
  AND2X1 U12689 ( .IN1(n12640), .IN2(n10772), .Q(n12638) );
  AND2X1 U12690 ( .IN1(n12641), .IN2(g2307), .Q(n12640) );
  AND2X1 U12691 ( .IN1(n12642), .IN2(n12601), .Q(n12636) );
  INVX0 U12692 ( .INP(n12641), .ZN(n12642) );
  OR2X1 U12693 ( .IN1(n5353), .IN2(n12627), .Q(n12641) );
  OR2X1 U12694 ( .IN1(n12609), .IN2(n5537), .Q(n12627) );
  OR2X1 U12695 ( .IN1(n12643), .IN2(n12644), .Q(g34002) );
  OR2X1 U12696 ( .IN1(n12645), .IN2(n12646), .Q(n12644) );
  AND2X1 U12697 ( .IN1(n10911), .IN2(g2295), .Q(n12646) );
  AND2X1 U12698 ( .IN1(n12647), .IN2(n10773), .Q(n12645) );
  AND2X1 U12699 ( .IN1(n12648), .IN2(g2303), .Q(n12647) );
  INVX0 U12700 ( .INP(n12649), .ZN(n12648) );
  AND2X1 U12701 ( .IN1(n12649), .IN2(n12601), .Q(n12643) );
  AND2X1 U12702 ( .IN1(n5537), .IN2(n12635), .Q(n12649) );
  OR2X1 U12703 ( .IN1(n12650), .IN2(n12651), .Q(g34001) );
  OR2X1 U12704 ( .IN1(n12652), .IN2(n12653), .Q(n12651) );
  AND2X1 U12705 ( .IN1(n10911), .IN2(g2299), .Q(n12653) );
  AND2X1 U12706 ( .IN1(n12654), .IN2(n10773), .Q(n12652) );
  AND2X1 U12707 ( .IN1(n12655), .IN2(g2295), .Q(n12654) );
  AND2X1 U12708 ( .IN1(n12656), .IN2(n12601), .Q(n12650) );
  INVX0 U12709 ( .INP(n12657), .ZN(n12601) );
  OR2X1 U12710 ( .IN1(n10881), .IN2(n12658), .Q(n12657) );
  AND2X1 U12711 ( .IN1(n12659), .IN2(n12617), .Q(n12658) );
  OR2X1 U12712 ( .IN1(n12660), .IN2(n12661), .Q(n12617) );
  OR2X1 U12713 ( .IN1(n12524), .IN2(n12662), .Q(n12661) );
  AND2X1 U12714 ( .IN1(n5343), .IN2(n12526), .Q(n12660) );
  OR2X1 U12715 ( .IN1(g1585), .IN2(n12619), .Q(n12659) );
  INVX0 U12716 ( .INP(n12655), .ZN(n12656) );
  OR2X1 U12717 ( .IN1(g2331), .IN2(n12663), .Q(n12655) );
  OR2X1 U12718 ( .IN1(n5353), .IN2(n12609), .Q(n12663) );
  OR2X1 U12719 ( .IN1(n12664), .IN2(n12665), .Q(g34000) );
  OR2X1 U12720 ( .IN1(n12666), .IN2(n12667), .Q(n12665) );
  AND2X1 U12721 ( .IN1(n12668), .IN2(g2165), .Q(n12667) );
  AND2X1 U12722 ( .IN1(n12669), .IN2(n12670), .Q(n12666) );
  AND2X1 U12723 ( .IN1(n10911), .IN2(g2246), .Q(n12664) );
  OR2X1 U12724 ( .IN1(n12671), .IN2(n12672), .Q(g33999) );
  AND2X1 U12725 ( .IN1(n12673), .IN2(n10773), .Q(n12672) );
  OR2X1 U12726 ( .IN1(n12674), .IN2(n12675), .Q(n12673) );
  AND2X1 U12727 ( .IN1(n12676), .IN2(g2241), .Q(n12675) );
  OR2X1 U12728 ( .IN1(n12677), .IN2(n12678), .Q(n12676) );
  AND2X1 U12729 ( .IN1(n12679), .IN2(g2153), .Q(n12677) );
  AND2X1 U12730 ( .IN1(n12680), .IN2(n12681), .Q(n12674) );
  INVX0 U12731 ( .INP(n12679), .ZN(n12681) );
  OR2X1 U12732 ( .IN1(n12682), .IN2(n12669), .Q(n12680) );
  AND2X1 U12733 ( .IN1(n10098), .IN2(n12683), .Q(n12682) );
  AND2X1 U12734 ( .IN1(n12684), .IN2(g2227), .Q(n12671) );
  OR2X1 U12735 ( .IN1(n10881), .IN2(n12685), .Q(n12684) );
  AND2X1 U12736 ( .IN1(n12679), .IN2(g2241), .Q(n12685) );
  AND2X1 U12737 ( .IN1(n12686), .IN2(n12687), .Q(n12679) );
  OR2X1 U12738 ( .IN1(n12688), .IN2(n5755), .Q(n12687) );
  OR2X1 U12739 ( .IN1(n12689), .IN2(n12690), .Q(g33998) );
  OR2X1 U12740 ( .IN1(n12691), .IN2(n12692), .Q(n12690) );
  AND2X1 U12741 ( .IN1(n10911), .IN2(g2169), .Q(n12692) );
  AND2X1 U12742 ( .IN1(n12693), .IN2(n10779), .Q(n12691) );
  AND2X1 U12743 ( .IN1(n12694), .IN2(g2181), .Q(n12693) );
  AND2X1 U12744 ( .IN1(n12695), .IN2(n12670), .Q(n12689) );
  INVX0 U12745 ( .INP(n12694), .ZN(n12695) );
  OR2X1 U12746 ( .IN1(g2197), .IN2(n12696), .Q(n12694) );
  OR2X1 U12747 ( .IN1(n12697), .IN2(n12698), .Q(g33997) );
  OR2X1 U12748 ( .IN1(n12699), .IN2(n12700), .Q(n12698) );
  AND2X1 U12749 ( .IN1(n10911), .IN2(g2181), .Q(n12700) );
  AND2X1 U12750 ( .IN1(n12701), .IN2(n10773), .Q(n12699) );
  AND2X1 U12751 ( .IN1(n12702), .IN2(n9352), .Q(n12701) );
  INVX0 U12752 ( .INP(n12703), .ZN(n12702) );
  AND2X1 U12753 ( .IN1(n12703), .IN2(n12670), .Q(n12697) );
  AND2X1 U12754 ( .IN1(n5356), .IN2(n12704), .Q(n12703) );
  OR2X1 U12755 ( .IN1(n12705), .IN2(n12706), .Q(g33996) );
  OR2X1 U12756 ( .IN1(n12707), .IN2(n12708), .Q(n12706) );
  AND2X1 U12757 ( .IN1(n10911), .IN2(n9352), .Q(n12708) );
  AND2X1 U12758 ( .IN1(n12709), .IN2(n10773), .Q(n12707) );
  AND2X1 U12759 ( .IN1(n12710), .IN2(g2173), .Q(n12709) );
  AND2X1 U12760 ( .IN1(n12711), .IN2(n12670), .Q(n12705) );
  INVX0 U12761 ( .INP(n12710), .ZN(n12711) );
  OR2X1 U12762 ( .IN1(n5356), .IN2(n12696), .Q(n12710) );
  OR2X1 U12763 ( .IN1(n12678), .IN2(n5538), .Q(n12696) );
  OR2X1 U12764 ( .IN1(n12712), .IN2(n12713), .Q(g33995) );
  OR2X1 U12765 ( .IN1(n12714), .IN2(n12715), .Q(n12713) );
  AND2X1 U12766 ( .IN1(n10911), .IN2(g2161), .Q(n12715) );
  AND2X1 U12767 ( .IN1(n12716), .IN2(n10773), .Q(n12714) );
  AND2X1 U12768 ( .IN1(n12717), .IN2(g2169), .Q(n12716) );
  INVX0 U12769 ( .INP(n12718), .ZN(n12717) );
  AND2X1 U12770 ( .IN1(n12718), .IN2(n12670), .Q(n12712) );
  AND2X1 U12771 ( .IN1(n5538), .IN2(n12704), .Q(n12718) );
  OR2X1 U12772 ( .IN1(n12719), .IN2(n12720), .Q(g33994) );
  OR2X1 U12773 ( .IN1(n12721), .IN2(n12722), .Q(n12720) );
  AND2X1 U12774 ( .IN1(n10912), .IN2(g2165), .Q(n12722) );
  AND2X1 U12775 ( .IN1(n12723), .IN2(n10773), .Q(n12721) );
  AND2X1 U12776 ( .IN1(n12724), .IN2(g2161), .Q(n12723) );
  AND2X1 U12777 ( .IN1(n12725), .IN2(n12670), .Q(n12719) );
  INVX0 U12778 ( .INP(n12726), .ZN(n12670) );
  OR2X1 U12779 ( .IN1(n10881), .IN2(n12727), .Q(n12726) );
  AND2X1 U12780 ( .IN1(n12728), .IN2(n12686), .Q(n12727) );
  OR2X1 U12781 ( .IN1(n12729), .IN2(n12730), .Q(n12686) );
  OR2X1 U12782 ( .IN1(n12524), .IN2(n12731), .Q(n12730) );
  AND2X1 U12783 ( .IN1(g1291), .IN2(n12526), .Q(n12524) );
  AND2X1 U12784 ( .IN1(n5289), .IN2(n12526), .Q(n12729) );
  AND2X1 U12785 ( .IN1(g4180), .IN2(n12732), .Q(n12526) );
  OR2X1 U12786 ( .IN1(n5757), .IN2(n12688), .Q(n12728) );
  INVX0 U12787 ( .INP(n12724), .ZN(n12725) );
  OR2X1 U12788 ( .IN1(g2197), .IN2(n12733), .Q(n12724) );
  OR2X1 U12789 ( .IN1(n5356), .IN2(n12678), .Q(n12733) );
  OR2X1 U12790 ( .IN1(n12734), .IN2(n12735), .Q(g33993) );
  OR2X1 U12791 ( .IN1(n12736), .IN2(n12737), .Q(n12735) );
  AND2X1 U12792 ( .IN1(n12738), .IN2(g2008), .Q(n12737) );
  AND2X1 U12793 ( .IN1(n12739), .IN2(n12740), .Q(n12736) );
  AND2X1 U12794 ( .IN1(n10912), .IN2(g2089), .Q(n12734) );
  OR2X1 U12795 ( .IN1(n12741), .IN2(n12742), .Q(g33992) );
  AND2X1 U12796 ( .IN1(n12743), .IN2(n10773), .Q(n12742) );
  OR2X1 U12797 ( .IN1(n12744), .IN2(n12745), .Q(n12743) );
  AND2X1 U12798 ( .IN1(n12746), .IN2(g2084), .Q(n12745) );
  OR2X1 U12799 ( .IN1(n12747), .IN2(n12748), .Q(n12746) );
  AND2X1 U12800 ( .IN1(n12749), .IN2(g1996), .Q(n12747) );
  AND2X1 U12801 ( .IN1(n12750), .IN2(n12751), .Q(n12744) );
  INVX0 U12802 ( .INP(n12749), .ZN(n12751) );
  OR2X1 U12803 ( .IN1(n12752), .IN2(n12739), .Q(n12750) );
  AND2X1 U12804 ( .IN1(n10093), .IN2(n12753), .Q(n12752) );
  AND2X1 U12805 ( .IN1(n12754), .IN2(g2070), .Q(n12741) );
  OR2X1 U12806 ( .IN1(n10881), .IN2(n12755), .Q(n12754) );
  AND2X1 U12807 ( .IN1(n12749), .IN2(g2084), .Q(n12755) );
  AND2X1 U12808 ( .IN1(n12756), .IN2(n12757), .Q(n12749) );
  OR2X1 U12809 ( .IN1(g1246), .IN2(n12758), .Q(n12757) );
  OR2X1 U12810 ( .IN1(n12759), .IN2(n12760), .Q(g33991) );
  OR2X1 U12811 ( .IN1(n12761), .IN2(n12762), .Q(n12760) );
  AND2X1 U12812 ( .IN1(n10912), .IN2(g2012), .Q(n12762) );
  AND2X1 U12813 ( .IN1(n12763), .IN2(n10773), .Q(n12761) );
  AND2X1 U12814 ( .IN1(n12764), .IN2(g2024), .Q(n12763) );
  AND2X1 U12815 ( .IN1(n12765), .IN2(n12740), .Q(n12759) );
  INVX0 U12816 ( .INP(n12764), .ZN(n12765) );
  OR2X1 U12817 ( .IN1(n12748), .IN2(n12156), .Q(n12764) );
  OR2X1 U12818 ( .IN1(n12766), .IN2(n12767), .Q(g33990) );
  OR2X1 U12819 ( .IN1(n12768), .IN2(n12769), .Q(n12767) );
  AND2X1 U12820 ( .IN1(n10912), .IN2(g2024), .Q(n12769) );
  AND2X1 U12821 ( .IN1(n12770), .IN2(n10774), .Q(n12768) );
  AND2X1 U12822 ( .IN1(n12771), .IN2(n9312), .Q(n12770) );
  INVX0 U12823 ( .INP(n12772), .ZN(n12771) );
  AND2X1 U12824 ( .IN1(n12772), .IN2(n12740), .Q(n12766) );
  AND2X1 U12825 ( .IN1(n5355), .IN2(n12773), .Q(n12772) );
  OR2X1 U12826 ( .IN1(n12774), .IN2(n12775), .Q(g33989) );
  OR2X1 U12827 ( .IN1(n12776), .IN2(n12777), .Q(n12775) );
  AND2X1 U12828 ( .IN1(n10912), .IN2(n9312), .Q(n12777) );
  AND2X1 U12829 ( .IN1(n12778), .IN2(n10774), .Q(n12776) );
  AND2X1 U12830 ( .IN1(n12779), .IN2(g2016), .Q(n12778) );
  INVX0 U12831 ( .INP(n12780), .ZN(n12779) );
  AND2X1 U12832 ( .IN1(n12780), .IN2(n12740), .Q(n12774) );
  AND2X1 U12833 ( .IN1(g2070), .IN2(n12781), .Q(n12780) );
  OR2X1 U12834 ( .IN1(n12782), .IN2(n12783), .Q(g33988) );
  OR2X1 U12835 ( .IN1(n12784), .IN2(n12785), .Q(n12783) );
  AND2X1 U12836 ( .IN1(n10912), .IN2(g2004), .Q(n12785) );
  AND2X1 U12837 ( .IN1(n12786), .IN2(n10774), .Q(n12784) );
  AND2X1 U12838 ( .IN1(n12787), .IN2(g2012), .Q(n12786) );
  INVX0 U12839 ( .INP(n12788), .ZN(n12787) );
  AND2X1 U12840 ( .IN1(n12788), .IN2(n12740), .Q(n12782) );
  AND2X1 U12841 ( .IN1(n5535), .IN2(n12773), .Q(n12788) );
  OR2X1 U12842 ( .IN1(n12789), .IN2(n12790), .Q(g33987) );
  OR2X1 U12843 ( .IN1(n12791), .IN2(n12792), .Q(n12790) );
  AND2X1 U12844 ( .IN1(n10912), .IN2(g2008), .Q(n12792) );
  AND2X1 U12845 ( .IN1(n12793), .IN2(n10774), .Q(n12791) );
  AND2X1 U12846 ( .IN1(n12794), .IN2(g2004), .Q(n12793) );
  INVX0 U12847 ( .INP(n12795), .ZN(n12794) );
  AND2X1 U12848 ( .IN1(n12795), .IN2(n12740), .Q(n12789) );
  AND2X1 U12849 ( .IN1(n10820), .IN2(n12796), .Q(n12740) );
  INVX0 U12850 ( .INP(n12797), .ZN(n12796) );
  AND2X1 U12851 ( .IN1(n12798), .IN2(n12756), .Q(n12797) );
  OR2X1 U12852 ( .IN1(n12799), .IN2(n12800), .Q(n12756) );
  OR2X1 U12853 ( .IN1(n12801), .IN2(n12802), .Q(n12800) );
  AND2X1 U12854 ( .IN1(n5341), .IN2(n12803), .Q(n12799) );
  OR2X1 U12855 ( .IN1(n12758), .IN2(g30332), .Q(n12798) );
  AND2X1 U12856 ( .IN1(n5505), .IN2(n12781), .Q(n12795) );
  OR2X1 U12857 ( .IN1(n12804), .IN2(n12805), .Q(g33986) );
  OR2X1 U12858 ( .IN1(n12806), .IN2(n12807), .Q(n12805) );
  AND2X1 U12859 ( .IN1(n12808), .IN2(g1874), .Q(n12807) );
  AND2X1 U12860 ( .IN1(n12809), .IN2(n12810), .Q(n12806) );
  AND2X1 U12861 ( .IN1(n10912), .IN2(g1955), .Q(n12804) );
  OR2X1 U12862 ( .IN1(n12811), .IN2(n12812), .Q(g33985) );
  AND2X1 U12863 ( .IN1(n12813), .IN2(n10774), .Q(n12812) );
  OR2X1 U12864 ( .IN1(n12814), .IN2(n12815), .Q(n12813) );
  AND2X1 U12865 ( .IN1(n12816), .IN2(g1950), .Q(n12815) );
  OR2X1 U12866 ( .IN1(n12817), .IN2(n12818), .Q(n12816) );
  AND2X1 U12867 ( .IN1(test_so8), .IN2(n12819), .Q(n12817) );
  AND2X1 U12868 ( .IN1(n12820), .IN2(n12821), .Q(n12814) );
  INVX0 U12869 ( .INP(n12819), .ZN(n12821) );
  OR2X1 U12870 ( .IN1(n12822), .IN2(n12809), .Q(n12820) );
  AND2X1 U12871 ( .IN1(n10097), .IN2(n12823), .Q(n12822) );
  AND2X1 U12872 ( .IN1(n12824), .IN2(g1936), .Q(n12811) );
  OR2X1 U12873 ( .IN1(n10882), .IN2(n12825), .Q(n12824) );
  AND2X1 U12874 ( .IN1(n12819), .IN2(g1950), .Q(n12825) );
  AND2X1 U12875 ( .IN1(n12826), .IN2(n12827), .Q(n12819) );
  OR2X1 U12876 ( .IN1(n12828), .IN2(n5756), .Q(n12827) );
  OR2X1 U12877 ( .IN1(n12829), .IN2(n12830), .Q(g33984) );
  OR2X1 U12878 ( .IN1(n12831), .IN2(n12832), .Q(n12830) );
  AND2X1 U12879 ( .IN1(n10912), .IN2(g1878), .Q(n12832) );
  INVX0 U12880 ( .INP(n12833), .ZN(n12831) );
  OR2X1 U12881 ( .IN1(n12834), .IN2(n10875), .Q(n12833) );
  OR2X1 U12882 ( .IN1(n12835), .IN2(n5799), .Q(n12834) );
  AND2X1 U12883 ( .IN1(n12835), .IN2(n12810), .Q(n12829) );
  AND2X1 U12884 ( .IN1(n12823), .IN2(n12162), .Q(n12835) );
  OR2X1 U12885 ( .IN1(n12836), .IN2(n12837), .Q(g33983) );
  OR2X1 U12886 ( .IN1(n12838), .IN2(n12839), .Q(n12837) );
  AND2X1 U12887 ( .IN1(n10912), .IN2(g1890), .Q(n12839) );
  AND2X1 U12888 ( .IN1(n12840), .IN2(n10774), .Q(n12838) );
  AND2X1 U12889 ( .IN1(n12841), .IN2(n9280), .Q(n12840) );
  INVX0 U12890 ( .INP(n12842), .ZN(n12841) );
  AND2X1 U12891 ( .IN1(n12842), .IN2(n12810), .Q(n12836) );
  AND2X1 U12892 ( .IN1(n10570), .IN2(n12843), .Q(n12842) );
  OR2X1 U12893 ( .IN1(n12844), .IN2(n12845), .Q(g33982) );
  OR2X1 U12894 ( .IN1(n12846), .IN2(n12847), .Q(n12845) );
  AND2X1 U12895 ( .IN1(n10912), .IN2(n9280), .Q(n12847) );
  AND2X1 U12896 ( .IN1(n12848), .IN2(n10774), .Q(n12846) );
  AND2X1 U12897 ( .IN1(n12849), .IN2(g1882), .Q(n12848) );
  INVX0 U12898 ( .INP(n12850), .ZN(n12849) );
  AND2X1 U12899 ( .IN1(n12850), .IN2(n12810), .Q(n12844) );
  AND2X1 U12900 ( .IN1(g1936), .IN2(n12851), .Q(n12850) );
  OR2X1 U12901 ( .IN1(n12852), .IN2(n12853), .Q(g33981) );
  OR2X1 U12902 ( .IN1(n12854), .IN2(n12855), .Q(n12853) );
  AND2X1 U12903 ( .IN1(n10912), .IN2(g1870), .Q(n12855) );
  AND2X1 U12904 ( .IN1(n12856), .IN2(n10774), .Q(n12854) );
  AND2X1 U12905 ( .IN1(n12857), .IN2(g1878), .Q(n12856) );
  INVX0 U12906 ( .INP(n12858), .ZN(n12857) );
  AND2X1 U12907 ( .IN1(n12858), .IN2(n12810), .Q(n12852) );
  AND2X1 U12908 ( .IN1(n5534), .IN2(n12843), .Q(n12858) );
  OR2X1 U12909 ( .IN1(n12859), .IN2(n12860), .Q(g33980) );
  OR2X1 U12910 ( .IN1(n12861), .IN2(n12862), .Q(n12860) );
  AND2X1 U12911 ( .IN1(n10912), .IN2(g1874), .Q(n12862) );
  AND2X1 U12912 ( .IN1(n12863), .IN2(n10774), .Q(n12861) );
  AND2X1 U12913 ( .IN1(n12864), .IN2(g1870), .Q(n12863) );
  INVX0 U12914 ( .INP(n12865), .ZN(n12864) );
  AND2X1 U12915 ( .IN1(n12865), .IN2(n12810), .Q(n12859) );
  INVX0 U12916 ( .INP(n12866), .ZN(n12810) );
  OR2X1 U12917 ( .IN1(n10882), .IN2(n12867), .Q(n12866) );
  AND2X1 U12918 ( .IN1(n12868), .IN2(n12826), .Q(n12867) );
  OR2X1 U12919 ( .IN1(n12869), .IN2(n12870), .Q(n12826) );
  OR2X1 U12920 ( .IN1(n12801), .IN2(n12871), .Q(n12870) );
  AND2X1 U12921 ( .IN1(n5329), .IN2(n12803), .Q(n12869) );
  OR2X1 U12922 ( .IN1(n5526), .IN2(n12828), .Q(n12868) );
  AND2X1 U12923 ( .IN1(n5503), .IN2(n12851), .Q(n12865) );
  OR2X1 U12924 ( .IN1(n12872), .IN2(n12873), .Q(g33979) );
  OR2X1 U12925 ( .IN1(n12874), .IN2(n12875), .Q(n12873) );
  AND2X1 U12926 ( .IN1(n12876), .IN2(g1740), .Q(n12875) );
  AND2X1 U12927 ( .IN1(n12877), .IN2(n12878), .Q(n12874) );
  AND2X1 U12928 ( .IN1(n10912), .IN2(g1821), .Q(n12872) );
  OR2X1 U12929 ( .IN1(n12879), .IN2(n12880), .Q(g33978) );
  AND2X1 U12930 ( .IN1(n12881), .IN2(n10775), .Q(n12880) );
  OR2X1 U12931 ( .IN1(n12882), .IN2(n12883), .Q(n12881) );
  AND2X1 U12932 ( .IN1(n12884), .IN2(g1816), .Q(n12883) );
  OR2X1 U12933 ( .IN1(n12885), .IN2(n12886), .Q(n12884) );
  AND2X1 U12934 ( .IN1(n12887), .IN2(g1728), .Q(n12885) );
  AND2X1 U12935 ( .IN1(n12888), .IN2(n12889), .Q(n12882) );
  INVX0 U12936 ( .INP(n12887), .ZN(n12889) );
  OR2X1 U12937 ( .IN1(n12890), .IN2(n12877), .Q(n12888) );
  AND2X1 U12938 ( .IN1(n10035), .IN2(n12891), .Q(n12890) );
  AND2X1 U12939 ( .IN1(n12892), .IN2(g1802), .Q(n12879) );
  OR2X1 U12940 ( .IN1(n10883), .IN2(n12893), .Q(n12892) );
  AND2X1 U12941 ( .IN1(n12887), .IN2(g1816), .Q(n12893) );
  AND2X1 U12942 ( .IN1(n12894), .IN2(n12895), .Q(n12887) );
  OR2X1 U12943 ( .IN1(n12896), .IN2(g1246), .Q(n12895) );
  OR2X1 U12944 ( .IN1(n12897), .IN2(n12898), .Q(g33977) );
  OR2X1 U12945 ( .IN1(n12899), .IN2(n12900), .Q(n12898) );
  AND2X1 U12946 ( .IN1(n10912), .IN2(g1744), .Q(n12900) );
  AND2X1 U12947 ( .IN1(n12901), .IN2(n10775), .Q(n12899) );
  AND2X1 U12948 ( .IN1(n12902), .IN2(g1756), .Q(n12901) );
  AND2X1 U12949 ( .IN1(n12903), .IN2(n12878), .Q(n12897) );
  INVX0 U12950 ( .INP(n12902), .ZN(n12903) );
  OR2X1 U12951 ( .IN1(g1772), .IN2(n12904), .Q(n12902) );
  OR2X1 U12952 ( .IN1(n12905), .IN2(n12906), .Q(g33976) );
  OR2X1 U12953 ( .IN1(n12907), .IN2(n12908), .Q(n12906) );
  AND2X1 U12954 ( .IN1(n10912), .IN2(g1756), .Q(n12908) );
  AND2X1 U12955 ( .IN1(n12909), .IN2(n10775), .Q(n12907) );
  AND2X1 U12956 ( .IN1(n12910), .IN2(g1752), .Q(n12909) );
  INVX0 U12957 ( .INP(n12911), .ZN(n12910) );
  AND2X1 U12958 ( .IN1(n12911), .IN2(n12878), .Q(n12905) );
  AND2X1 U12959 ( .IN1(n5352), .IN2(n12912), .Q(n12911) );
  OR2X1 U12960 ( .IN1(n12913), .IN2(n12914), .Q(g33975) );
  OR2X1 U12961 ( .IN1(n12915), .IN2(n12916), .Q(n12914) );
  AND2X1 U12962 ( .IN1(n10912), .IN2(g1752), .Q(n12916) );
  AND2X1 U12963 ( .IN1(n12917), .IN2(n10775), .Q(n12915) );
  AND2X1 U12964 ( .IN1(n12918), .IN2(g1748), .Q(n12917) );
  AND2X1 U12965 ( .IN1(n12919), .IN2(n12878), .Q(n12913) );
  INVX0 U12966 ( .INP(n12918), .ZN(n12919) );
  OR2X1 U12967 ( .IN1(n5352), .IN2(n12904), .Q(n12918) );
  OR2X1 U12968 ( .IN1(n12886), .IN2(n5536), .Q(n12904) );
  OR2X1 U12969 ( .IN1(n12920), .IN2(n12921), .Q(g33974) );
  OR2X1 U12970 ( .IN1(n12922), .IN2(n12923), .Q(n12921) );
  AND2X1 U12971 ( .IN1(n10912), .IN2(g1736), .Q(n12923) );
  AND2X1 U12972 ( .IN1(n12924), .IN2(n10775), .Q(n12922) );
  AND2X1 U12973 ( .IN1(n12925), .IN2(g1744), .Q(n12924) );
  INVX0 U12974 ( .INP(n12926), .ZN(n12925) );
  AND2X1 U12975 ( .IN1(n12926), .IN2(n12878), .Q(n12920) );
  AND2X1 U12976 ( .IN1(n5536), .IN2(n12912), .Q(n12926) );
  OR2X1 U12977 ( .IN1(n12927), .IN2(n12928), .Q(g33973) );
  OR2X1 U12978 ( .IN1(n12929), .IN2(n12930), .Q(n12928) );
  AND2X1 U12979 ( .IN1(n10912), .IN2(g1740), .Q(n12930) );
  AND2X1 U12980 ( .IN1(n12931), .IN2(n10775), .Q(n12929) );
  AND2X1 U12981 ( .IN1(n12932), .IN2(g1736), .Q(n12931) );
  AND2X1 U12982 ( .IN1(n12933), .IN2(n12878), .Q(n12927) );
  INVX0 U12983 ( .INP(n12934), .ZN(n12878) );
  OR2X1 U12984 ( .IN1(n10883), .IN2(n12935), .Q(n12934) );
  AND2X1 U12985 ( .IN1(n12936), .IN2(n12894), .Q(n12935) );
  OR2X1 U12986 ( .IN1(n12937), .IN2(n12938), .Q(n12894) );
  OR2X1 U12987 ( .IN1(n12801), .IN2(n12939), .Q(n12938) );
  AND2X1 U12988 ( .IN1(n5478), .IN2(n12803), .Q(n12937) );
  OR2X1 U12989 ( .IN1(g30332), .IN2(n12896), .Q(n12936) );
  INVX0 U12990 ( .INP(n12932), .ZN(n12933) );
  OR2X1 U12991 ( .IN1(g1772), .IN2(n12940), .Q(n12932) );
  OR2X1 U12992 ( .IN1(n5352), .IN2(n12886), .Q(n12940) );
  OR2X1 U12993 ( .IN1(n12941), .IN2(n12942), .Q(g33972) );
  OR2X1 U12994 ( .IN1(n12943), .IN2(n12944), .Q(n12942) );
  AND2X1 U12995 ( .IN1(n12945), .IN2(g1604), .Q(n12944) );
  AND2X1 U12996 ( .IN1(n12946), .IN2(n12947), .Q(n12943) );
  AND2X1 U12997 ( .IN1(n10913), .IN2(g1687), .Q(n12941) );
  OR2X1 U12998 ( .IN1(n12948), .IN2(n12949), .Q(g33971) );
  AND2X1 U12999 ( .IN1(n12950), .IN2(n10775), .Q(n12949) );
  OR2X1 U13000 ( .IN1(n12951), .IN2(n12952), .Q(n12950) );
  AND2X1 U13001 ( .IN1(n12953), .IN2(g1682), .Q(n12952) );
  OR2X1 U13002 ( .IN1(n12954), .IN2(n12955), .Q(n12953) );
  AND2X1 U13003 ( .IN1(n12956), .IN2(g1592), .Q(n12954) );
  AND2X1 U13004 ( .IN1(n12957), .IN2(n12958), .Q(n12951) );
  INVX0 U13005 ( .INP(n12956), .ZN(n12958) );
  OR2X1 U13006 ( .IN1(n12959), .IN2(n12946), .Q(n12957) );
  AND2X1 U13007 ( .IN1(n10099), .IN2(n12960), .Q(n12959) );
  AND2X1 U13008 ( .IN1(n12961), .IN2(g1668), .Q(n12948) );
  OR2X1 U13009 ( .IN1(n10883), .IN2(n12962), .Q(n12961) );
  AND2X1 U13010 ( .IN1(n12956), .IN2(g1682), .Q(n12962) );
  AND2X1 U13011 ( .IN1(n12963), .IN2(n12964), .Q(n12956) );
  OR2X1 U13012 ( .IN1(n12965), .IN2(n5756), .Q(n12964) );
  OR2X1 U13013 ( .IN1(n12966), .IN2(n12967), .Q(g33970) );
  OR2X1 U13014 ( .IN1(n12968), .IN2(n12969), .Q(n12967) );
  AND2X1 U13015 ( .IN1(n10913), .IN2(g1608), .Q(n12969) );
  AND2X1 U13016 ( .IN1(n12970), .IN2(n10775), .Q(n12968) );
  AND2X1 U13017 ( .IN1(n12971), .IN2(g1620), .Q(n12970) );
  INVX0 U13018 ( .INP(n12972), .ZN(n12971) );
  AND2X1 U13019 ( .IN1(n12972), .IN2(n12947), .Q(n12966) );
  AND2X1 U13020 ( .IN1(n12960), .IN2(g31862), .Q(n12972) );
  OR2X1 U13021 ( .IN1(n12973), .IN2(n12974), .Q(g33969) );
  OR2X1 U13022 ( .IN1(n12975), .IN2(n12976), .Q(n12974) );
  AND2X1 U13023 ( .IN1(n10913), .IN2(g1620), .Q(n12976) );
  AND2X1 U13024 ( .IN1(n12977), .IN2(n10775), .Q(n12975) );
  AND2X1 U13025 ( .IN1(n12978), .IN2(n9303), .Q(n12977) );
  INVX0 U13026 ( .INP(n12979), .ZN(n12978) );
  AND2X1 U13027 ( .IN1(n12979), .IN2(n12947), .Q(n12973) );
  AND2X1 U13028 ( .IN1(n5362), .IN2(n12980), .Q(n12979) );
  OR2X1 U13029 ( .IN1(n12981), .IN2(n12982), .Q(g33968) );
  OR2X1 U13030 ( .IN1(n12983), .IN2(n12984), .Q(n12982) );
  AND2X1 U13031 ( .IN1(n10913), .IN2(n9303), .Q(n12984) );
  AND2X1 U13032 ( .IN1(n12985), .IN2(n10776), .Q(n12983) );
  AND2X1 U13033 ( .IN1(n12986), .IN2(g1612), .Q(n12985) );
  INVX0 U13034 ( .INP(n12987), .ZN(n12986) );
  AND2X1 U13035 ( .IN1(n12987), .IN2(n12947), .Q(n12981) );
  AND2X1 U13036 ( .IN1(g1668), .IN2(n12988), .Q(n12987) );
  OR2X1 U13037 ( .IN1(n12989), .IN2(n12990), .Q(g33967) );
  OR2X1 U13038 ( .IN1(n12991), .IN2(n12992), .Q(n12990) );
  AND2X1 U13039 ( .IN1(n10913), .IN2(g1600), .Q(n12992) );
  AND2X1 U13040 ( .IN1(n12993), .IN2(n10776), .Q(n12991) );
  AND2X1 U13041 ( .IN1(n12994), .IN2(g1608), .Q(n12993) );
  INVX0 U13042 ( .INP(n12995), .ZN(n12994) );
  AND2X1 U13043 ( .IN1(n12995), .IN2(n12947), .Q(n12989) );
  AND2X1 U13044 ( .IN1(n5598), .IN2(n12980), .Q(n12995) );
  OR2X1 U13045 ( .IN1(n12996), .IN2(n12997), .Q(g33966) );
  OR2X1 U13046 ( .IN1(n12998), .IN2(n12999), .Q(n12997) );
  AND2X1 U13047 ( .IN1(n10913), .IN2(g1604), .Q(n12999) );
  AND2X1 U13048 ( .IN1(n13000), .IN2(n10776), .Q(n12998) );
  AND2X1 U13049 ( .IN1(n13001), .IN2(g1600), .Q(n13000) );
  INVX0 U13050 ( .INP(n13002), .ZN(n13001) );
  AND2X1 U13051 ( .IN1(n13002), .IN2(n12947), .Q(n12996) );
  AND2X1 U13052 ( .IN1(n10819), .IN2(n13003), .Q(n12947) );
  INVX0 U13053 ( .INP(n13004), .ZN(n13003) );
  AND2X1 U13054 ( .IN1(n13005), .IN2(n12963), .Q(n13004) );
  OR2X1 U13055 ( .IN1(n13006), .IN2(n13007), .Q(n12963) );
  OR2X1 U13056 ( .IN1(n12801), .IN2(n13008), .Q(n13007) );
  AND2X1 U13057 ( .IN1(g947), .IN2(n12803), .Q(n12801) );
  AND2X1 U13058 ( .IN1(n5328), .IN2(n12803), .Q(n13006) );
  AND2X1 U13059 ( .IN1(g4180), .IN2(n13009), .Q(n12803) );
  OR2X1 U13060 ( .IN1(n5526), .IN2(n12965), .Q(n13005) );
  AND2X1 U13061 ( .IN1(n5549), .IN2(n12988), .Q(n13002) );
  OR2X1 U13062 ( .IN1(n13010), .IN2(n13011), .Q(g33965) );
  OR2X1 U13063 ( .IN1(n13012), .IN2(n13013), .Q(n13011) );
  AND2X1 U13064 ( .IN1(n2704), .IN2(n5333), .Q(n13013) );
  AND2X1 U13065 ( .IN1(n13014), .IN2(g767), .Q(n13012) );
  AND2X1 U13066 ( .IN1(n2404), .IN2(n13015), .Q(n13014) );
  INVX0 U13067 ( .INP(n2704), .ZN(n13015) );
  AND2X1 U13068 ( .IN1(n10913), .IN2(g763), .Q(n13010) );
  OR2X1 U13069 ( .IN1(n13016), .IN2(n13017), .Q(g33964) );
  OR2X1 U13070 ( .IN1(n13018), .IN2(n13019), .Q(n13017) );
  AND2X1 U13071 ( .IN1(n2706), .IN2(n5550), .Q(n13019) );
  AND2X1 U13072 ( .IN1(n13020), .IN2(g599), .Q(n13018) );
  AND2X1 U13073 ( .IN1(n2421), .IN2(n13021), .Q(n13020) );
  INVX0 U13074 ( .INP(n2706), .ZN(n13021) );
  AND2X1 U13075 ( .IN1(n10913), .IN2(g595), .Q(n13016) );
  OR2X1 U13076 ( .IN1(n13022), .IN2(n13023), .Q(g33963) );
  AND2X1 U13077 ( .IN1(n13024), .IN2(n10776), .Q(n13023) );
  AND2X1 U13078 ( .IN1(n13025), .IN2(n13026), .Q(n13024) );
  OR2X1 U13079 ( .IN1(n13027), .IN2(n13028), .Q(n13026) );
  OR2X1 U13080 ( .IN1(g73), .IN2(n13029), .Q(n13028) );
  AND2X1 U13081 ( .IN1(n13030), .IN2(g269), .Q(n13029) );
  AND2X1 U13082 ( .IN1(g72), .IN2(g262), .Q(n13027) );
  OR2X1 U13083 ( .IN1(n13031), .IN2(n11628), .Q(n13025) );
  AND2X1 U13084 ( .IN1(n13030), .IN2(g255), .Q(n13031) );
  AND2X1 U13085 ( .IN1(n10913), .IN2(g29215), .Q(n13022) );
  OR2X1 U13086 ( .IN1(n13032), .IN2(n13033), .Q(g33962) );
  AND2X1 U13087 ( .IN1(n13034), .IN2(n10776), .Q(n13033) );
  AND2X1 U13088 ( .IN1(n13035), .IN2(n13036), .Q(n13034) );
  OR2X1 U13089 ( .IN1(n13037), .IN2(n11628), .Q(n13036) );
  AND2X1 U13090 ( .IN1(n13038), .IN2(n13039), .Q(n13037) );
  OR2X1 U13091 ( .IN1(g225), .IN2(n13030), .Q(n13039) );
  OR2X1 U13092 ( .IN1(g72), .IN2(g232), .Q(n13038) );
  OR2X1 U13093 ( .IN1(n13040), .IN2(n13041), .Q(n13035) );
  OR2X1 U13094 ( .IN1(g73), .IN2(n13042), .Q(n13041) );
  AND2X1 U13095 ( .IN1(n13030), .IN2(g246), .Q(n13042) );
  AND2X1 U13096 ( .IN1(g72), .IN2(g239), .Q(n13040) );
  INVX0 U13097 ( .INP(n13043), .ZN(n13032) );
  OR2X1 U13098 ( .IN1(n10739), .IN2(n10116), .Q(n13043) );
  OR2X1 U13099 ( .IN1(n13044), .IN2(n13045), .Q(g33961) );
  OR2X1 U13100 ( .IN1(n13046), .IN2(n13047), .Q(n13045) );
  AND2X1 U13101 ( .IN1(n2989), .IN2(n5675), .Q(n13047) );
  AND2X1 U13102 ( .IN1(n13048), .IN2(g298), .Q(n13046) );
  AND2X1 U13103 ( .IN1(n10534), .IN2(n13049), .Q(n13048) );
  INVX0 U13104 ( .INP(n2989), .ZN(n13049) );
  AND2X1 U13105 ( .IN1(n10913), .IN2(g294), .Q(n13044) );
  OR2X1 U13106 ( .IN1(n13050), .IN2(n13051), .Q(g33960) );
  OR2X1 U13107 ( .IN1(n13052), .IN2(n13053), .Q(n13051) );
  AND2X1 U13108 ( .IN1(n2991), .IN2(n5678), .Q(n13053) );
  AND2X1 U13109 ( .IN1(n13054), .IN2(g157), .Q(n13052) );
  AND2X1 U13110 ( .IN1(n13055), .IN2(n13056), .Q(n13054) );
  INVX0 U13111 ( .INP(n2991), .ZN(n13056) );
  AND2X1 U13112 ( .IN1(n10913), .IN2(g153), .Q(n13050) );
  OR2X1 U13113 ( .IN1(n13057), .IN2(n13058), .Q(g33935) );
  OR2X1 U13114 ( .IN1(g34649), .IN2(n12214), .Q(n13058) );
  OR2X1 U13115 ( .IN1(n13059), .IN2(n13060), .Q(g34649) );
  OR2X1 U13116 ( .IN1(n13061), .IN2(n13062), .Q(n13060) );
  OR2X1 U13117 ( .IN1(n13063), .IN2(n13064), .Q(n13059) );
  OR2X1 U13118 ( .IN1(n10113), .IN2(n10112), .Q(n13057) );
  OR2X1 U13119 ( .IN1(g18881), .IN2(n13065), .Q(g33874) );
  OR2X1 U13120 ( .IN1(n5846), .IN2(n12214), .Q(n13065) );
  OR2X1 U13121 ( .IN1(n13066), .IN2(n13067), .Q(g33659) );
  OR2X1 U13122 ( .IN1(n12107), .IN2(n11221), .Q(n13067) );
  OR2X1 U13123 ( .IN1(n13068), .IN2(n13069), .Q(n11221) );
  AND2X1 U13124 ( .IN1(n13070), .IN2(g4098), .Q(n13069) );
  OR2X1 U13125 ( .IN1(n13071), .IN2(n13072), .Q(n13070) );
  OR2X1 U13126 ( .IN1(n13073), .IN2(n13074), .Q(n13072) );
  AND2X1 U13127 ( .IN1(n13075), .IN2(n12105), .Q(n13074) );
  AND2X1 U13128 ( .IN1(n13076), .IN2(g4093), .Q(n13073) );
  AND2X1 U13129 ( .IN1(n13077), .IN2(n13078), .Q(n13076) );
  OR2X1 U13130 ( .IN1(n13079), .IN2(g4087), .Q(n13078) );
  OR2X1 U13131 ( .IN1(n5480), .IN2(n13080), .Q(n13077) );
  AND2X1 U13132 ( .IN1(n13081), .IN2(n13082), .Q(n13071) );
  AND2X1 U13133 ( .IN1(n5350), .IN2(n13083), .Q(n13068) );
  OR2X1 U13134 ( .IN1(n13084), .IN2(n13085), .Q(n13083) );
  OR2X1 U13135 ( .IN1(n13086), .IN2(n13087), .Q(n13085) );
  AND2X1 U13136 ( .IN1(g32975), .IN2(n12105), .Q(n13087) );
  AND2X1 U13137 ( .IN1(n13088), .IN2(g4093), .Q(n13086) );
  AND2X1 U13138 ( .IN1(n13089), .IN2(n13090), .Q(n13088) );
  OR2X1 U13139 ( .IN1(n13091), .IN2(g4087), .Q(n13090) );
  OR2X1 U13140 ( .IN1(n5480), .IN2(n13092), .Q(n13089) );
  AND2X1 U13141 ( .IN1(n13093), .IN2(n13081), .Q(n13084) );
  OR2X1 U13142 ( .IN1(n12214), .IN2(n13094), .Q(n12107) );
  INVX0 U13143 ( .INP(n11182), .ZN(n13066) );
  AND2X1 U13144 ( .IN1(n13095), .IN2(n13096), .Q(n11182) );
  XNOR2X1 U13145 ( .IN1(n5715), .IN2(n11205), .Q(n13096) );
  XNOR2X1 U13146 ( .IN1(n10274), .IN2(n13097), .Q(n13095) );
  OR2X1 U13147 ( .IN1(n13098), .IN2(n13099), .Q(g33636) );
  OR2X1 U13148 ( .IN1(g34657), .IN2(n12214), .Q(n13099) );
  INVX0 U13149 ( .INP(n2668), .ZN(n12214) );
  OR2X1 U13150 ( .IN1(n13100), .IN2(g134), .Q(n2668) );
  AND2X1 U13151 ( .IN1(g99), .IN2(g37), .Q(n13100) );
  OR2X1 U13152 ( .IN1(n13101), .IN2(n13102), .Q(g34657) );
  OR2X1 U13153 ( .IN1(n13103), .IN2(n13104), .Q(n13102) );
  OR2X1 U13154 ( .IN1(n13105), .IN2(n13106), .Q(n13101) );
  OR2X1 U13155 ( .IN1(n10115), .IN2(n10114), .Q(n13098) );
  OR2X1 U13156 ( .IN1(n13107), .IN2(n13108), .Q(g33627) );
  AND2X1 U13157 ( .IN1(n10913), .IN2(g6741), .Q(n13108) );
  AND2X1 U13158 ( .IN1(n13109), .IN2(n13110), .Q(n13107) );
  OR2X1 U13159 ( .IN1(n13111), .IN2(n13112), .Q(n13109) );
  AND2X1 U13160 ( .IN1(n11095), .IN2(n13113), .Q(n13112) );
  AND2X1 U13161 ( .IN1(n13114), .IN2(n10776), .Q(n13111) );
  OR2X1 U13162 ( .IN1(n13115), .IN2(n11092), .Q(n13114) );
  AND2X1 U13163 ( .IN1(n10540), .IN2(g6682), .Q(n13115) );
  OR2X1 U13164 ( .IN1(n13116), .IN2(n13117), .Q(g33626) );
  OR2X1 U13165 ( .IN1(n13118), .IN2(n13119), .Q(n13117) );
  AND2X1 U13166 ( .IN1(n10913), .IN2(g6736), .Q(n13119) );
  AND2X1 U13167 ( .IN1(n13120), .IN2(n10776), .Q(n13118) );
  AND2X1 U13168 ( .IN1(n13121), .IN2(n5398), .Q(n13120) );
  AND2X1 U13169 ( .IN1(n13110), .IN2(n13113), .Q(n13121) );
  OR2X1 U13170 ( .IN1(n13122), .IN2(n13123), .Q(n13110) );
  OR2X1 U13171 ( .IN1(n12108), .IN2(n13124), .Q(n13123) );
  OR2X1 U13172 ( .IN1(test_so81), .IN2(n10540), .Q(n13122) );
  AND2X1 U13173 ( .IN1(n13125), .IN2(g6741), .Q(n13116) );
  OR2X1 U13174 ( .IN1(n13126), .IN2(n13127), .Q(g33625) );
  AND2X1 U13175 ( .IN1(n10913), .IN2(g6395), .Q(n13127) );
  AND2X1 U13176 ( .IN1(n13128), .IN2(n13129), .Q(n13126) );
  OR2X1 U13177 ( .IN1(n13130), .IN2(n13131), .Q(n13128) );
  AND2X1 U13178 ( .IN1(n13132), .IN2(n13133), .Q(n13131) );
  AND2X1 U13179 ( .IN1(n13134), .IN2(n10776), .Q(n13130) );
  OR2X1 U13180 ( .IN1(n13135), .IN2(n13136), .Q(n13134) );
  AND2X1 U13181 ( .IN1(n13137), .IN2(g6336), .Q(n13135) );
  OR2X1 U13182 ( .IN1(n13138), .IN2(n13139), .Q(g33624) );
  OR2X1 U13183 ( .IN1(n13140), .IN2(n13141), .Q(n13139) );
  AND2X1 U13184 ( .IN1(n13142), .IN2(n5396), .Q(n13141) );
  AND2X1 U13185 ( .IN1(n13143), .IN2(n13129), .Q(n13142) );
  OR2X1 U13186 ( .IN1(n13144), .IN2(n13145), .Q(n13129) );
  OR2X1 U13187 ( .IN1(n13137), .IN2(n13146), .Q(n13145) );
  AND2X1 U13188 ( .IN1(n13147), .IN2(g6395), .Q(n13140) );
  AND2X1 U13189 ( .IN1(n10913), .IN2(g6390), .Q(n13138) );
  OR2X1 U13190 ( .IN1(n13148), .IN2(n13149), .Q(g33623) );
  AND2X1 U13191 ( .IN1(test_so57), .IN2(n10897), .Q(n13149) );
  AND2X1 U13192 ( .IN1(n13150), .IN2(n13151), .Q(n13148) );
  OR2X1 U13193 ( .IN1(n13152), .IN2(n13153), .Q(n13150) );
  AND2X1 U13194 ( .IN1(n13154), .IN2(n13155), .Q(n13153) );
  AND2X1 U13195 ( .IN1(n13156), .IN2(n10776), .Q(n13152) );
  OR2X1 U13196 ( .IN1(n13157), .IN2(n13158), .Q(n13156) );
  AND2X1 U13197 ( .IN1(n13159), .IN2(g5990), .Q(n13157) );
  OR2X1 U13198 ( .IN1(n13160), .IN2(n13161), .Q(g33622) );
  OR2X1 U13199 ( .IN1(n13162), .IN2(n13163), .Q(n13161) );
  AND2X1 U13200 ( .IN1(n13164), .IN2(test_so57), .Q(n13163) );
  AND2X1 U13201 ( .IN1(n13165), .IN2(n10559), .Q(n13162) );
  AND2X1 U13202 ( .IN1(n13166), .IN2(n13151), .Q(n13165) );
  OR2X1 U13203 ( .IN1(n13167), .IN2(n13168), .Q(n13151) );
  OR2X1 U13204 ( .IN1(n13146), .IN2(n13159), .Q(n13168) );
  OR2X1 U13205 ( .IN1(test_so81), .IN2(n12109), .Q(n13167) );
  AND2X1 U13206 ( .IN1(test_so50), .IN2(n10896), .Q(n13160) );
  OR2X1 U13207 ( .IN1(n13169), .IN2(n13170), .Q(g33621) );
  AND2X1 U13208 ( .IN1(n10913), .IN2(g5703), .Q(n13170) );
  AND2X1 U13209 ( .IN1(n13171), .IN2(n13172), .Q(n13169) );
  OR2X1 U13210 ( .IN1(n13173), .IN2(n13174), .Q(n13171) );
  AND2X1 U13211 ( .IN1(n13175), .IN2(n13176), .Q(n13174) );
  AND2X1 U13212 ( .IN1(n13177), .IN2(n10777), .Q(n13173) );
  OR2X1 U13213 ( .IN1(n13178), .IN2(n13179), .Q(n13177) );
  AND2X1 U13214 ( .IN1(n13180), .IN2(g5644), .Q(n13178) );
  OR2X1 U13215 ( .IN1(n13181), .IN2(n13182), .Q(g33620) );
  OR2X1 U13216 ( .IN1(n13183), .IN2(n13184), .Q(n13182) );
  AND2X1 U13217 ( .IN1(n10913), .IN2(g5698), .Q(n13184) );
  AND2X1 U13218 ( .IN1(n13185), .IN2(n10777), .Q(n13183) );
  AND2X1 U13219 ( .IN1(n13186), .IN2(n5397), .Q(n13185) );
  AND2X1 U13220 ( .IN1(n13176), .IN2(n13172), .Q(n13186) );
  OR2X1 U13221 ( .IN1(n13144), .IN2(n13187), .Q(n13172) );
  OR2X1 U13222 ( .IN1(n13124), .IN2(n13180), .Q(n13187) );
  OR2X1 U13223 ( .IN1(n12109), .IN2(n10552), .Q(n13144) );
  AND2X1 U13224 ( .IN1(n13188), .IN2(g5703), .Q(n13181) );
  OR2X1 U13225 ( .IN1(n13189), .IN2(n13190), .Q(g33619) );
  AND2X1 U13226 ( .IN1(n10913), .IN2(g5357), .Q(n13190) );
  AND2X1 U13227 ( .IN1(n13191), .IN2(n13192), .Q(n13189) );
  OR2X1 U13228 ( .IN1(n13193), .IN2(n13194), .Q(n13191) );
  AND2X1 U13229 ( .IN1(n11086), .IN2(g33959), .Q(n13194) );
  AND2X1 U13230 ( .IN1(n13195), .IN2(n10777), .Q(n13193) );
  OR2X1 U13231 ( .IN1(n13196), .IN2(n11083), .Q(n13195) );
  AND2X1 U13232 ( .IN1(n10535), .IN2(g5297), .Q(n13196) );
  OR2X1 U13233 ( .IN1(n13197), .IN2(n13198), .Q(g33618) );
  OR2X1 U13234 ( .IN1(n13199), .IN2(n13200), .Q(n13198) );
  AND2X1 U13235 ( .IN1(n10914), .IN2(g5352), .Q(n13200) );
  AND2X1 U13236 ( .IN1(n13201), .IN2(n10777), .Q(n13199) );
  AND2X1 U13237 ( .IN1(n13202), .IN2(n5393), .Q(n13201) );
  AND2X1 U13238 ( .IN1(n13192), .IN2(g33959), .Q(n13202) );
  OR2X1 U13239 ( .IN1(n13203), .IN2(n13204), .Q(n13192) );
  OR2X1 U13240 ( .IN1(n12109), .IN2(n13124), .Q(n13204) );
  OR2X1 U13241 ( .IN1(n13205), .IN2(g4311), .Q(n12109) );
  OR2X1 U13242 ( .IN1(test_so81), .IN2(n10535), .Q(n13203) );
  AND2X1 U13243 ( .IN1(n13206), .IN2(g5357), .Q(n13197) );
  OR2X1 U13244 ( .IN1(n13207), .IN2(n13208), .Q(g33617) );
  AND2X1 U13245 ( .IN1(n12446), .IN2(n10777), .Q(n13208) );
  OR2X1 U13246 ( .IN1(n13209), .IN2(n13210), .Q(n12446) );
  AND2X1 U13247 ( .IN1(n13211), .IN2(g4581), .Q(n13210) );
  OR2X1 U13248 ( .IN1(n11594), .IN2(g4575), .Q(n13211) );
  AND2X1 U13249 ( .IN1(n5670), .IN2(g4552), .Q(n13209) );
  AND2X1 U13250 ( .IN1(n10914), .IN2(g4552), .Q(n13207) );
  OR2X1 U13251 ( .IN1(n13212), .IN2(n13213), .Q(g33616) );
  AND2X1 U13252 ( .IN1(n12437), .IN2(n10777), .Q(n13213) );
  OR2X1 U13253 ( .IN1(n13214), .IN2(n13215), .Q(n12437) );
  AND2X1 U13254 ( .IN1(n13216), .IN2(g4581), .Q(n13215) );
  OR2X1 U13255 ( .IN1(test_so100), .IN2(n11594), .Q(n13216) );
  AND2X1 U13256 ( .IN1(n5670), .IN2(g4512), .Q(n13214) );
  AND2X1 U13257 ( .IN1(n10914), .IN2(g4515), .Q(n13212) );
  OR2X1 U13258 ( .IN1(n13217), .IN2(n13218), .Q(g33614) );
  AND2X1 U13259 ( .IN1(n10914), .IN2(g4054), .Q(n13218) );
  AND2X1 U13260 ( .IN1(n13219), .IN2(n13220), .Q(n13217) );
  OR2X1 U13261 ( .IN1(n13221), .IN2(n13222), .Q(n13219) );
  AND2X1 U13262 ( .IN1(n13223), .IN2(n13224), .Q(n13222) );
  AND2X1 U13263 ( .IN1(n13225), .IN2(n10777), .Q(n13221) );
  OR2X1 U13264 ( .IN1(n13226), .IN2(n13227), .Q(n13225) );
  AND2X1 U13265 ( .IN1(n13228), .IN2(g3990), .Q(n13226) );
  OR2X1 U13266 ( .IN1(n13229), .IN2(n13230), .Q(g33613) );
  OR2X1 U13267 ( .IN1(n13231), .IN2(n13232), .Q(n13230) );
  AND2X1 U13268 ( .IN1(n13233), .IN2(n5395), .Q(n13232) );
  AND2X1 U13269 ( .IN1(n13234), .IN2(n13220), .Q(n13233) );
  OR2X1 U13270 ( .IN1(n13235), .IN2(n13236), .Q(n13220) );
  OR2X1 U13271 ( .IN1(n13146), .IN2(n13228), .Q(n13236) );
  AND2X1 U13272 ( .IN1(n13237), .IN2(g4054), .Q(n13231) );
  AND2X1 U13273 ( .IN1(n10914), .IN2(g4049), .Q(n13229) );
  OR2X1 U13274 ( .IN1(n13238), .IN2(n13239), .Q(g33612) );
  AND2X1 U13275 ( .IN1(n10914), .IN2(g3703), .Q(n13239) );
  AND2X1 U13276 ( .IN1(n13240), .IN2(n13241), .Q(n13238) );
  OR2X1 U13277 ( .IN1(n13242), .IN2(n13243), .Q(n13240) );
  AND2X1 U13278 ( .IN1(n13244), .IN2(n13245), .Q(n13243) );
  AND2X1 U13279 ( .IN1(n13246), .IN2(n10777), .Q(n13242) );
  OR2X1 U13280 ( .IN1(n13247), .IN2(n13248), .Q(n13246) );
  AND2X1 U13281 ( .IN1(n13249), .IN2(g3639), .Q(n13247) );
  OR2X1 U13282 ( .IN1(n13250), .IN2(n13251), .Q(g33611) );
  OR2X1 U13283 ( .IN1(n13252), .IN2(n13253), .Q(n13251) );
  AND2X1 U13284 ( .IN1(n13254), .IN2(n5399), .Q(n13253) );
  AND2X1 U13285 ( .IN1(n13255), .IN2(n13241), .Q(n13254) );
  OR2X1 U13286 ( .IN1(n13256), .IN2(n13257), .Q(n13241) );
  OR2X1 U13287 ( .IN1(n13146), .IN2(n13249), .Q(n13257) );
  INVX0 U13288 ( .INP(n3033), .ZN(n13146) );
  OR2X1 U13289 ( .IN1(test_so81), .IN2(n12108), .Q(n13256) );
  AND2X1 U13290 ( .IN1(n13258), .IN2(g3703), .Q(n13252) );
  AND2X1 U13291 ( .IN1(n10914), .IN2(g3698), .Q(n13250) );
  OR2X1 U13292 ( .IN1(n13259), .IN2(n13260), .Q(g33610) );
  AND2X1 U13293 ( .IN1(n13261), .IN2(n10777), .Q(n13260) );
  AND2X1 U13294 ( .IN1(n13262), .IN2(n13263), .Q(n13261) );
  OR2X1 U13295 ( .IN1(n13264), .IN2(n13265), .Q(n13262) );
  OR2X1 U13296 ( .IN1(n13266), .IN2(n13267), .Q(n13265) );
  AND2X1 U13297 ( .IN1(n13268), .IN2(g3288), .Q(n13267) );
  AND2X1 U13298 ( .IN1(n13269), .IN2(n13270), .Q(n13266) );
  AND2X1 U13299 ( .IN1(n10914), .IN2(g3352), .Q(n13259) );
  OR2X1 U13300 ( .IN1(n13271), .IN2(n13272), .Q(g33609) );
  OR2X1 U13301 ( .IN1(n13273), .IN2(n13274), .Q(n13272) );
  AND2X1 U13302 ( .IN1(n10914), .IN2(g3347), .Q(n13274) );
  AND2X1 U13303 ( .IN1(n13275), .IN2(n10778), .Q(n13273) );
  AND2X1 U13304 ( .IN1(n13276), .IN2(n5604), .Q(n13275) );
  AND2X1 U13305 ( .IN1(n13270), .IN2(n13263), .Q(n13276) );
  OR2X1 U13306 ( .IN1(n13235), .IN2(n13277), .Q(n13263) );
  OR2X1 U13307 ( .IN1(n13124), .IN2(n13268), .Q(n13277) );
  INVX0 U13308 ( .INP(n3023), .ZN(n13124) );
  OR2X1 U13309 ( .IN1(n10552), .IN2(n12108), .Q(n13235) );
  OR2X1 U13310 ( .IN1(n5323), .IN2(n13205), .Q(n12108) );
  OR2X1 U13311 ( .IN1(n11630), .IN2(n13278), .Q(n13205) );
  XNOR2X1 U13312 ( .IN1(g73), .IN2(n5540), .Q(n13278) );
  XNOR2X1 U13313 ( .IN1(g72), .IN2(n5506), .Q(n11630) );
  AND2X1 U13314 ( .IN1(n13279), .IN2(g3352), .Q(n13271) );
  OR2X1 U13315 ( .IN1(n13280), .IN2(n13281), .Q(g33608) );
  OR2X1 U13316 ( .IN1(n2787), .IN2(n13282), .Q(n13281) );
  AND2X1 U13317 ( .IN1(n13283), .IN2(n10530), .Q(n13282) );
  OR2X1 U13318 ( .IN1(n13284), .IN2(n13285), .Q(n13280) );
  AND2X1 U13319 ( .IN1(test_so30), .IN2(n10896), .Q(n13285) );
  AND2X1 U13320 ( .IN1(n13286), .IN2(n10778), .Q(n13284) );
  AND2X1 U13321 ( .IN1(n12455), .IN2(g2759), .Q(n13286) );
  INVX0 U13322 ( .INP(n13283), .ZN(n12455) );
  AND2X1 U13323 ( .IN1(test_so30), .IN2(n2790), .Q(n13283) );
  OR2X1 U13324 ( .IN1(n13287), .IN2(n13288), .Q(g33607) );
  OR2X1 U13325 ( .IN1(n13289), .IN2(n13290), .Q(n13288) );
  AND2X1 U13326 ( .IN1(n13291), .IN2(g2606), .Q(n13290) );
  OR2X1 U13327 ( .IN1(n13292), .IN2(n13293), .Q(n13291) );
  INVX0 U13328 ( .INP(n13294), .ZN(n13292) );
  OR2X1 U13329 ( .IN1(n10884), .IN2(n3105), .Q(n13294) );
  AND2X1 U13330 ( .IN1(n13295), .IN2(n646), .Q(n13289) );
  AND2X1 U13331 ( .IN1(n13296), .IN2(n13297), .Q(n13295) );
  OR2X1 U13332 ( .IN1(g2599), .IN2(n13298), .Q(n13297) );
  OR2X1 U13333 ( .IN1(n5521), .IN2(n10463), .Q(n13298) );
  OR2X1 U13334 ( .IN1(n13299), .IN2(n13300), .Q(n13296) );
  AND2X1 U13335 ( .IN1(n3111), .IN2(n10778), .Q(n13300) );
  AND2X1 U13336 ( .IN1(n13301), .IN2(n12167), .Q(n13299) );
  AND2X1 U13337 ( .IN1(n13302), .IN2(g2629), .Q(n12167) );
  INVX0 U13338 ( .INP(n2726), .ZN(n13302) );
  OR2X1 U13339 ( .IN1(g504), .IN2(n12143), .Q(n2726) );
  AND2X1 U13340 ( .IN1(n5524), .IN2(n12005), .Q(n13301) );
  AND2X1 U13341 ( .IN1(n10914), .IN2(g2555), .Q(n13287) );
  OR2X1 U13342 ( .IN1(n13303), .IN2(n13304), .Q(g33606) );
  OR2X1 U13343 ( .IN1(n13305), .IN2(n13306), .Q(n13304) );
  AND2X1 U13344 ( .IN1(n10914), .IN2(g2671), .Q(n13306) );
  AND2X1 U13345 ( .IN1(n13307), .IN2(n10778), .Q(n13305) );
  AND2X1 U13346 ( .IN1(n5457), .IN2(n12461), .Q(n13307) );
  AND2X1 U13347 ( .IN1(n12460), .IN2(g2675), .Q(n13303) );
  OR2X1 U13348 ( .IN1(n13308), .IN2(n13309), .Q(g33605) );
  OR2X1 U13349 ( .IN1(n13310), .IN2(n13311), .Q(n13309) );
  AND2X1 U13350 ( .IN1(n13312), .IN2(n10585), .Q(n13311) );
  AND2X1 U13351 ( .IN1(n13313), .IN2(n5418), .Q(n13312) );
  AND2X1 U13352 ( .IN1(n12461), .IN2(n10778), .Q(n13313) );
  AND2X1 U13353 ( .IN1(test_so48), .IN2(n13314), .Q(n13310) );
  OR2X1 U13354 ( .IN1(n10877), .IN2(n13315), .Q(n13314) );
  AND2X1 U13355 ( .IN1(n12461), .IN2(g2661), .Q(n13315) );
  AND2X1 U13356 ( .IN1(n12460), .IN2(g2671), .Q(n13308) );
  OR2X1 U13357 ( .IN1(n13316), .IN2(n13317), .Q(g33604) );
  AND2X1 U13358 ( .IN1(n13318), .IN2(g2661), .Q(n13317) );
  AND2X1 U13359 ( .IN1(test_so48), .IN2(n12460), .Q(n13316) );
  OR2X1 U13360 ( .IN1(n13319), .IN2(n13320), .Q(g33603) );
  AND2X1 U13361 ( .IN1(n13318), .IN2(g2643), .Q(n13320) );
  AND2X1 U13362 ( .IN1(n12460), .IN2(g2648), .Q(n13319) );
  INVX0 U13363 ( .INP(n13318), .ZN(n12460) );
  OR2X1 U13364 ( .IN1(n10884), .IN2(n12461), .Q(n13318) );
  AND2X1 U13365 ( .IN1(n5521), .IN2(n13321), .Q(n12461) );
  AND2X1 U13366 ( .IN1(n12475), .IN2(n5351), .Q(n13321) );
  OR2X1 U13367 ( .IN1(n13322), .IN2(n13323), .Q(g33602) );
  OR2X1 U13368 ( .IN1(n13324), .IN2(n13325), .Q(n13323) );
  AND2X1 U13369 ( .IN1(n12496), .IN2(n13326), .Q(n13325) );
  AND2X1 U13370 ( .IN1(n12475), .IN2(g2599), .Q(n12496) );
  AND2X1 U13371 ( .IN1(n13327), .IN2(g2629), .Q(n13324) );
  AND2X1 U13372 ( .IN1(n10914), .IN2(g2599), .Q(n13322) );
  OR2X1 U13373 ( .IN1(n13328), .IN2(n13329), .Q(g33601) );
  OR2X1 U13374 ( .IN1(n13330), .IN2(n13331), .Q(n13329) );
  AND2X1 U13375 ( .IN1(n13332), .IN2(n10778), .Q(n13331) );
  AND2X1 U13376 ( .IN1(n13333), .IN2(n12475), .Q(n13332) );
  AND2X1 U13377 ( .IN1(n13326), .IN2(g2555), .Q(n13333) );
  AND2X1 U13378 ( .IN1(n10914), .IN2(g2606), .Q(n13330) );
  AND2X1 U13379 ( .IN1(n13327), .IN2(g2599), .Q(n13328) );
  OR2X1 U13380 ( .IN1(n13334), .IN2(n13335), .Q(g33600) );
  AND2X1 U13381 ( .IN1(n13327), .IN2(g2555), .Q(n13335) );
  AND2X1 U13382 ( .IN1(n10818), .IN2(n12470), .Q(n13327) );
  INVX0 U13383 ( .INP(n12475), .ZN(n12470) );
  AND2X1 U13384 ( .IN1(n13336), .IN2(n13337), .Q(n13334) );
  AND2X1 U13385 ( .IN1(n10818), .IN2(n13326), .Q(n13337) );
  INVX0 U13386 ( .INP(n3111), .ZN(n13326) );
  AND2X1 U13387 ( .IN1(n5521), .IN2(n13338), .Q(n13336) );
  OR2X1 U13388 ( .IN1(n12488), .IN2(g2555), .Q(n13338) );
  AND2X1 U13389 ( .IN1(n12475), .IN2(n5524), .Q(n12488) );
  OR2X1 U13390 ( .IN1(n646), .IN2(n12480), .Q(n12475) );
  OR2X1 U13391 ( .IN1(n13339), .IN2(n13340), .Q(n12480) );
  OR2X1 U13392 ( .IN1(n13341), .IN2(n13342), .Q(n13340) );
  AND2X1 U13393 ( .IN1(n13343), .IN2(g2697), .Q(n13342) );
  AND2X1 U13394 ( .IN1(n2549), .IN2(g1300), .Q(n13339) );
  AND2X1 U13395 ( .IN1(n13344), .IN2(g1430), .Q(n646) );
  OR2X1 U13396 ( .IN1(n13345), .IN2(g1514), .Q(n13344) );
  OR2X1 U13397 ( .IN1(n13346), .IN2(test_so49), .Q(n13345) );
  OR2X1 U13398 ( .IN1(n13347), .IN2(n13348), .Q(g33599) );
  OR2X1 U13399 ( .IN1(n13349), .IN2(n13350), .Q(n13348) );
  AND2X1 U13400 ( .IN1(n13351), .IN2(g2472), .Q(n13350) );
  OR2X1 U13401 ( .IN1(n13352), .IN2(n13293), .Q(n13351) );
  INVX0 U13402 ( .INP(n13353), .ZN(n13352) );
  OR2X1 U13403 ( .IN1(n10884), .IN2(n3125), .Q(n13353) );
  INVX0 U13404 ( .INP(n3121), .ZN(n13349) );
  OR2X1 U13405 ( .IN1(n13354), .IN2(n13355), .Q(n3121) );
  OR2X1 U13406 ( .IN1(n12160), .IN2(n13356), .Q(n13355) );
  OR2X1 U13407 ( .IN1(g112), .IN2(n13357), .Q(n13354) );
  OR2X1 U13408 ( .IN1(n2727), .IN2(n13358), .Q(n13357) );
  OR2X1 U13409 ( .IN1(n5519), .IN2(n12143), .Q(n2727) );
  OR2X1 U13410 ( .IN1(n5287), .IN2(n13359), .Q(n12143) );
  OR2X1 U13411 ( .IN1(n13360), .IN2(n13361), .Q(n13347) );
  AND2X1 U13412 ( .IN1(n13362), .IN2(n10778), .Q(n13361) );
  AND2X1 U13413 ( .IN1(n13363), .IN2(n3131), .Q(n13362) );
  AND2X1 U13414 ( .IN1(n662), .IN2(n13364), .Q(n13363) );
  OR2X1 U13415 ( .IN1(n10463), .IN2(n12160), .Q(n13364) );
  OR2X1 U13416 ( .IN1(n5522), .IN2(g2465), .Q(n12160) );
  INVX0 U13417 ( .INP(n13356), .ZN(n662) );
  AND2X1 U13418 ( .IN1(test_so79), .IN2(n10896), .Q(n13360) );
  OR2X1 U13419 ( .IN1(n13365), .IN2(n13366), .Q(g33598) );
  OR2X1 U13420 ( .IN1(n13367), .IN2(n13368), .Q(n13366) );
  AND2X1 U13421 ( .IN1(n10914), .IN2(g2537), .Q(n13368) );
  AND2X1 U13422 ( .IN1(n13369), .IN2(n10778), .Q(n13367) );
  AND2X1 U13423 ( .IN1(n5461), .IN2(n12532), .Q(n13369) );
  AND2X1 U13424 ( .IN1(n12531), .IN2(g2541), .Q(n13365) );
  OR2X1 U13425 ( .IN1(n13370), .IN2(n13371), .Q(g33597) );
  OR2X1 U13426 ( .IN1(n13372), .IN2(n13373), .Q(n13371) );
  AND2X1 U13427 ( .IN1(n13374), .IN2(n5761), .Q(n13373) );
  AND2X1 U13428 ( .IN1(n13375), .IN2(n5420), .Q(n13374) );
  AND2X1 U13429 ( .IN1(n12532), .IN2(n10778), .Q(n13375) );
  AND2X1 U13430 ( .IN1(n13376), .IN2(g2533), .Q(n13372) );
  OR2X1 U13431 ( .IN1(n10884), .IN2(n13377), .Q(n13376) );
  AND2X1 U13432 ( .IN1(n12532), .IN2(g2527), .Q(n13377) );
  AND2X1 U13433 ( .IN1(n12531), .IN2(g2537), .Q(n13370) );
  OR2X1 U13434 ( .IN1(n13378), .IN2(n13379), .Q(g33596) );
  AND2X1 U13435 ( .IN1(n13380), .IN2(g2527), .Q(n13379) );
  AND2X1 U13436 ( .IN1(n12531), .IN2(g2533), .Q(n13378) );
  OR2X1 U13437 ( .IN1(n13381), .IN2(n13382), .Q(g33595) );
  AND2X1 U13438 ( .IN1(n13380), .IN2(g2509), .Q(n13382) );
  AND2X1 U13439 ( .IN1(n12531), .IN2(g2514), .Q(n13381) );
  INVX0 U13440 ( .INP(n13380), .ZN(n12531) );
  OR2X1 U13441 ( .IN1(n10884), .IN2(n12532), .Q(n13380) );
  AND2X1 U13442 ( .IN1(n5522), .IN2(n13383), .Q(n12532) );
  AND2X1 U13443 ( .IN1(n10569), .IN2(n12546), .Q(n13383) );
  OR2X1 U13444 ( .IN1(n13384), .IN2(n13385), .Q(g33594) );
  OR2X1 U13445 ( .IN1(n13386), .IN2(n13387), .Q(n13385) );
  AND2X1 U13446 ( .IN1(n12566), .IN2(n13388), .Q(n13387) );
  AND2X1 U13447 ( .IN1(n12546), .IN2(g2465), .Q(n12566) );
  AND2X1 U13448 ( .IN1(n13389), .IN2(g2495), .Q(n13386) );
  AND2X1 U13449 ( .IN1(n10914), .IN2(g2465), .Q(n13384) );
  OR2X1 U13450 ( .IN1(n13390), .IN2(n13391), .Q(g33593) );
  OR2X1 U13451 ( .IN1(n13392), .IN2(n13393), .Q(n13391) );
  AND2X1 U13452 ( .IN1(n13394), .IN2(n10779), .Q(n13393) );
  AND2X1 U13453 ( .IN1(n12574), .IN2(n13388), .Q(n13394) );
  AND2X1 U13454 ( .IN1(n12546), .IN2(test_so79), .Q(n12574) );
  AND2X1 U13455 ( .IN1(n10914), .IN2(g2472), .Q(n13392) );
  AND2X1 U13456 ( .IN1(n13389), .IN2(g2465), .Q(n13390) );
  OR2X1 U13457 ( .IN1(n13395), .IN2(n13396), .Q(g33592) );
  AND2X1 U13458 ( .IN1(n13389), .IN2(test_so79), .Q(n13396) );
  AND2X1 U13459 ( .IN1(n10817), .IN2(n12541), .Q(n13389) );
  AND2X1 U13460 ( .IN1(n13397), .IN2(n13398), .Q(n13395) );
  AND2X1 U13461 ( .IN1(n10817), .IN2(n13388), .Q(n13398) );
  INVX0 U13462 ( .INP(n3131), .ZN(n13388) );
  AND2X1 U13463 ( .IN1(n5522), .IN2(n13399), .Q(n13397) );
  OR2X1 U13464 ( .IN1(n13400), .IN2(test_so79), .Q(n13399) );
  AND2X1 U13465 ( .IN1(n5523), .IN2(n12546), .Q(n13400) );
  INVX0 U13466 ( .INP(n12541), .ZN(n12546) );
  AND2X1 U13467 ( .IN1(n13356), .IN2(n12594), .Q(n12541) );
  INVX0 U13468 ( .INP(n12551), .ZN(n12594) );
  OR2X1 U13469 ( .IN1(n13401), .IN2(n13402), .Q(n12551) );
  OR2X1 U13470 ( .IN1(n13341), .IN2(n13403), .Q(n13402) );
  AND2X1 U13471 ( .IN1(n13404), .IN2(n5377), .Q(n13403) );
  AND2X1 U13472 ( .IN1(g2697), .IN2(g2689), .Q(n13404) );
  AND2X1 U13473 ( .IN1(n2549), .IN2(g1472), .Q(n13401) );
  OR2X1 U13474 ( .IN1(n13405), .IN2(n10516), .Q(n13356) );
  AND2X1 U13475 ( .IN1(n13406), .IN2(n13407), .Q(n13405) );
  OR2X1 U13476 ( .IN1(n13408), .IN2(n13409), .Q(g33591) );
  OR2X1 U13477 ( .IN1(n13410), .IN2(n13411), .Q(n13409) );
  AND2X1 U13478 ( .IN1(n13412), .IN2(g2338), .Q(n13411) );
  OR2X1 U13479 ( .IN1(n13413), .IN2(n13293), .Q(n13412) );
  INVX0 U13480 ( .INP(n13414), .ZN(n13413) );
  OR2X1 U13481 ( .IN1(n10884), .IN2(n3145), .Q(n13414) );
  AND2X1 U13482 ( .IN1(n13415), .IN2(n333), .Q(n13410) );
  INVX0 U13483 ( .INP(n13416), .ZN(n333) );
  AND2X1 U13484 ( .IN1(n13417), .IN2(n13418), .Q(n13415) );
  OR2X1 U13485 ( .IN1(g2331), .IN2(n13419), .Q(n13418) );
  OR2X1 U13486 ( .IN1(n5537), .IN2(n10463), .Q(n13419) );
  OR2X1 U13487 ( .IN1(n13420), .IN2(n13421), .Q(n13417) );
  AND2X1 U13488 ( .IN1(n13422), .IN2(n10779), .Q(n13421) );
  INVX0 U13489 ( .INP(n13423), .ZN(n13422) );
  AND2X1 U13490 ( .IN1(n12169), .IN2(n12005), .Q(n13420) );
  AND2X1 U13491 ( .IN1(n5513), .IN2(n13424), .Q(n12169) );
  AND2X1 U13492 ( .IN1(g2361), .IN2(n13425), .Q(n13424) );
  INVX0 U13493 ( .INP(n3146), .ZN(n13425) );
  AND2X1 U13494 ( .IN1(n10914), .IN2(g2287), .Q(n13408) );
  OR2X1 U13495 ( .IN1(n13426), .IN2(n13427), .Q(g33590) );
  OR2X1 U13496 ( .IN1(n13428), .IN2(n13429), .Q(n13427) );
  AND2X1 U13497 ( .IN1(test_so31), .IN2(n10896), .Q(n13429) );
  AND2X1 U13498 ( .IN1(n13430), .IN2(n10779), .Q(n13428) );
  AND2X1 U13499 ( .IN1(n5459), .IN2(n12600), .Q(n13430) );
  AND2X1 U13500 ( .IN1(n12599), .IN2(g2407), .Q(n13426) );
  OR2X1 U13501 ( .IN1(n13431), .IN2(n13432), .Q(g33589) );
  OR2X1 U13502 ( .IN1(n13433), .IN2(n13434), .Q(n13432) );
  AND2X1 U13503 ( .IN1(n13435), .IN2(n5762), .Q(n13434) );
  AND2X1 U13504 ( .IN1(n13436), .IN2(n5421), .Q(n13435) );
  AND2X1 U13505 ( .IN1(n12600), .IN2(n10754), .Q(n13436) );
  AND2X1 U13506 ( .IN1(n13437), .IN2(g2399), .Q(n13433) );
  OR2X1 U13507 ( .IN1(n10884), .IN2(n13438), .Q(n13437) );
  AND2X1 U13508 ( .IN1(n12600), .IN2(g2393), .Q(n13438) );
  AND2X1 U13509 ( .IN1(test_so31), .IN2(n12599), .Q(n13431) );
  OR2X1 U13510 ( .IN1(n13439), .IN2(n13440), .Q(g33588) );
  AND2X1 U13511 ( .IN1(n13441), .IN2(g2393), .Q(n13440) );
  AND2X1 U13512 ( .IN1(n12599), .IN2(g2399), .Q(n13439) );
  OR2X1 U13513 ( .IN1(n13442), .IN2(n13443), .Q(g33587) );
  AND2X1 U13514 ( .IN1(n13441), .IN2(g2375), .Q(n13443) );
  AND2X1 U13515 ( .IN1(n12599), .IN2(g2380), .Q(n13442) );
  INVX0 U13516 ( .INP(n13441), .ZN(n12599) );
  OR2X1 U13517 ( .IN1(n10884), .IN2(n12600), .Q(n13441) );
  AND2X1 U13518 ( .IN1(n5537), .IN2(n13444), .Q(n12600) );
  AND2X1 U13519 ( .IN1(n12614), .IN2(n5353), .Q(n13444) );
  OR2X1 U13520 ( .IN1(n13445), .IN2(n13446), .Q(g33586) );
  OR2X1 U13521 ( .IN1(n13447), .IN2(n13448), .Q(n13446) );
  AND2X1 U13522 ( .IN1(n12635), .IN2(n13423), .Q(n13448) );
  AND2X1 U13523 ( .IN1(n12614), .IN2(g2331), .Q(n12635) );
  AND2X1 U13524 ( .IN1(n13449), .IN2(g2361), .Q(n13447) );
  AND2X1 U13525 ( .IN1(n10914), .IN2(g2331), .Q(n13445) );
  OR2X1 U13526 ( .IN1(n13450), .IN2(n13451), .Q(g33585) );
  OR2X1 U13527 ( .IN1(n13452), .IN2(n13453), .Q(n13451) );
  AND2X1 U13528 ( .IN1(n13454), .IN2(n10747), .Q(n13453) );
  AND2X1 U13529 ( .IN1(n13455), .IN2(n12614), .Q(n13454) );
  AND2X1 U13530 ( .IN1(n13423), .IN2(g2287), .Q(n13455) );
  AND2X1 U13531 ( .IN1(n10914), .IN2(g2338), .Q(n13452) );
  AND2X1 U13532 ( .IN1(n13449), .IN2(g2331), .Q(n13450) );
  OR2X1 U13533 ( .IN1(n13456), .IN2(n13457), .Q(g33584) );
  AND2X1 U13534 ( .IN1(n13449), .IN2(g2287), .Q(n13457) );
  AND2X1 U13535 ( .IN1(n10817), .IN2(n12609), .Q(n13449) );
  AND2X1 U13536 ( .IN1(n13458), .IN2(n13459), .Q(n13456) );
  AND2X1 U13537 ( .IN1(n13423), .IN2(n10754), .Q(n13459) );
  OR2X1 U13538 ( .IN1(n3146), .IN2(n13460), .Q(n13423) );
  OR2X1 U13539 ( .IN1(n13359), .IN2(n13461), .Q(n3146) );
  AND2X1 U13540 ( .IN1(n5537), .IN2(n13462), .Q(n13458) );
  OR2X1 U13541 ( .IN1(n13463), .IN2(g2287), .Q(n13462) );
  AND2X1 U13542 ( .IN1(n5513), .IN2(n12614), .Q(n13463) );
  INVX0 U13543 ( .INP(n12609), .ZN(n12614) );
  AND2X1 U13544 ( .IN1(n13416), .IN2(n12662), .Q(n12609) );
  INVX0 U13545 ( .INP(n12619), .ZN(n12662) );
  OR2X1 U13546 ( .IN1(n13464), .IN2(n13465), .Q(n12619) );
  OR2X1 U13547 ( .IN1(n13341), .IN2(n13466), .Q(n13465) );
  AND2X1 U13548 ( .IN1(n13343), .IN2(n5308), .Q(n13466) );
  AND2X1 U13549 ( .IN1(g2689), .IN2(g2704), .Q(n13343) );
  AND2X1 U13550 ( .IN1(n2549), .IN2(g1448), .Q(n13464) );
  OR2X1 U13551 ( .IN1(n13467), .IN2(n10129), .Q(n13416) );
  AND2X1 U13552 ( .IN1(n13468), .IN2(n13406), .Q(n13467) );
  OR2X1 U13553 ( .IN1(n13469), .IN2(n13470), .Q(g33583) );
  OR2X1 U13554 ( .IN1(n13471), .IN2(n13472), .Q(n13470) );
  AND2X1 U13555 ( .IN1(n13473), .IN2(g2204), .Q(n13472) );
  OR2X1 U13556 ( .IN1(n13474), .IN2(n13293), .Q(n13473) );
  INVX0 U13557 ( .INP(n13475), .ZN(n13474) );
  OR2X1 U13558 ( .IN1(n10884), .IN2(n3164), .Q(n13475) );
  AND2X1 U13559 ( .IN1(n13476), .IN2(n658), .Q(n13471) );
  INVX0 U13560 ( .INP(n13477), .ZN(n658) );
  AND2X1 U13561 ( .IN1(n13478), .IN2(n13479), .Q(n13476) );
  OR2X1 U13562 ( .IN1(g2197), .IN2(n13480), .Q(n13479) );
  OR2X1 U13563 ( .IN1(n5538), .IN2(n10463), .Q(n13480) );
  OR2X1 U13564 ( .IN1(n13481), .IN2(n13482), .Q(n13478) );
  AND2X1 U13565 ( .IN1(n13483), .IN2(n10754), .Q(n13482) );
  INVX0 U13566 ( .INP(n13484), .ZN(n13483) );
  AND2X1 U13567 ( .IN1(n12168), .IN2(n12005), .Q(n13481) );
  AND2X1 U13568 ( .IN1(n5514), .IN2(n13485), .Q(n12168) );
  AND2X1 U13569 ( .IN1(g2227), .IN2(n13486), .Q(n13485) );
  INVX0 U13570 ( .INP(n3165), .ZN(n13486) );
  AND2X1 U13571 ( .IN1(n10915), .IN2(g2153), .Q(n13469) );
  OR2X1 U13572 ( .IN1(n13487), .IN2(n13488), .Q(g33582) );
  OR2X1 U13573 ( .IN1(n13489), .IN2(n13490), .Q(n13488) );
  AND2X1 U13574 ( .IN1(n10915), .IN2(g2269), .Q(n13490) );
  AND2X1 U13575 ( .IN1(n13491), .IN2(n10754), .Q(n13489) );
  AND2X1 U13576 ( .IN1(n5458), .IN2(n12669), .Q(n13491) );
  AND2X1 U13577 ( .IN1(n12668), .IN2(g2273), .Q(n13487) );
  OR2X1 U13578 ( .IN1(n13492), .IN2(n13493), .Q(g33581) );
  OR2X1 U13579 ( .IN1(n13494), .IN2(n13495), .Q(n13493) );
  AND2X1 U13580 ( .IN1(n13496), .IN2(n10586), .Q(n13495) );
  AND2X1 U13581 ( .IN1(n13497), .IN2(n5419), .Q(n13496) );
  AND2X1 U13582 ( .IN1(n12669), .IN2(n10754), .Q(n13497) );
  AND2X1 U13583 ( .IN1(test_so62), .IN2(n13498), .Q(n13494) );
  OR2X1 U13584 ( .IN1(n10884), .IN2(n13499), .Q(n13498) );
  AND2X1 U13585 ( .IN1(n12669), .IN2(g2259), .Q(n13499) );
  AND2X1 U13586 ( .IN1(n12668), .IN2(g2269), .Q(n13492) );
  OR2X1 U13587 ( .IN1(n13500), .IN2(n13501), .Q(g33580) );
  AND2X1 U13588 ( .IN1(n13502), .IN2(g2259), .Q(n13501) );
  AND2X1 U13589 ( .IN1(test_so62), .IN2(n12668), .Q(n13500) );
  OR2X1 U13590 ( .IN1(n13503), .IN2(n13504), .Q(g33579) );
  AND2X1 U13591 ( .IN1(n13502), .IN2(g2241), .Q(n13504) );
  AND2X1 U13592 ( .IN1(n12668), .IN2(g2246), .Q(n13503) );
  INVX0 U13593 ( .INP(n13502), .ZN(n12668) );
  OR2X1 U13594 ( .IN1(n10884), .IN2(n12669), .Q(n13502) );
  AND2X1 U13595 ( .IN1(n5538), .IN2(n13505), .Q(n12669) );
  AND2X1 U13596 ( .IN1(n12683), .IN2(n5356), .Q(n13505) );
  OR2X1 U13597 ( .IN1(n13506), .IN2(n13507), .Q(g33578) );
  OR2X1 U13598 ( .IN1(n13508), .IN2(n13509), .Q(n13507) );
  AND2X1 U13599 ( .IN1(n12704), .IN2(n13484), .Q(n13509) );
  AND2X1 U13600 ( .IN1(n12683), .IN2(g2197), .Q(n12704) );
  AND2X1 U13601 ( .IN1(n13510), .IN2(g2227), .Q(n13508) );
  AND2X1 U13602 ( .IN1(n10915), .IN2(g2197), .Q(n13506) );
  OR2X1 U13603 ( .IN1(n13511), .IN2(n13512), .Q(g33577) );
  OR2X1 U13604 ( .IN1(n13513), .IN2(n13514), .Q(n13512) );
  AND2X1 U13605 ( .IN1(n13515), .IN2(n10753), .Q(n13514) );
  AND2X1 U13606 ( .IN1(n13516), .IN2(n12683), .Q(n13515) );
  AND2X1 U13607 ( .IN1(n13484), .IN2(g2153), .Q(n13516) );
  AND2X1 U13608 ( .IN1(n10915), .IN2(g2204), .Q(n13513) );
  AND2X1 U13609 ( .IN1(n13510), .IN2(g2197), .Q(n13511) );
  OR2X1 U13610 ( .IN1(n13517), .IN2(n13518), .Q(g33576) );
  AND2X1 U13611 ( .IN1(n13510), .IN2(g2153), .Q(n13518) );
  AND2X1 U13612 ( .IN1(n10816), .IN2(n12678), .Q(n13510) );
  AND2X1 U13613 ( .IN1(n13519), .IN2(n13520), .Q(n13517) );
  AND2X1 U13614 ( .IN1(n13484), .IN2(n10753), .Q(n13520) );
  OR2X1 U13615 ( .IN1(n3165), .IN2(n13460), .Q(n13484) );
  OR2X1 U13616 ( .IN1(n13359), .IN2(n13521), .Q(n3165) );
  INVX0 U13617 ( .INP(n3116), .ZN(n13359) );
  AND2X1 U13618 ( .IN1(n5538), .IN2(n13522), .Q(n13519) );
  OR2X1 U13619 ( .IN1(n13523), .IN2(g2153), .Q(n13522) );
  AND2X1 U13620 ( .IN1(n5514), .IN2(n12683), .Q(n13523) );
  INVX0 U13621 ( .INP(n12678), .ZN(n12683) );
  AND2X1 U13622 ( .IN1(n13477), .IN2(n12731), .Q(n12678) );
  INVX0 U13623 ( .INP(n12688), .ZN(n12731) );
  OR2X1 U13624 ( .IN1(n13524), .IN2(n13525), .Q(n12688) );
  OR2X1 U13625 ( .IN1(n13341), .IN2(n13526), .Q(n13525) );
  AND2X1 U13626 ( .IN1(n13527), .IN2(n5308), .Q(n13526) );
  AND2X1 U13627 ( .IN1(n5377), .IN2(g2689), .Q(n13527) );
  INVX0 U13628 ( .INP(n12732), .ZN(n13341) );
  OR2X1 U13629 ( .IN1(n13528), .IN2(g134), .Q(n12732) );
  AND2X1 U13630 ( .IN1(n13529), .IN2(n5595), .Q(n13528) );
  AND2X1 U13631 ( .IN1(n13530), .IN2(g691), .Q(n13529) );
  AND2X1 U13632 ( .IN1(n2549), .IN2(g1478), .Q(n13524) );
  OR2X1 U13633 ( .IN1(n13531), .IN2(n10130), .Q(n13477) );
  AND2X1 U13634 ( .IN1(n13532), .IN2(n13406), .Q(n13531) );
  INVX0 U13635 ( .INP(n13346), .ZN(n13406) );
  OR2X1 U13636 ( .IN1(n13533), .IN2(n13534), .Q(n13346) );
  OR2X1 U13637 ( .IN1(n10550), .IN2(n13535), .Q(n13534) );
  OR2X1 U13638 ( .IN1(g1548), .IN2(g1554), .Q(n13535) );
  OR2X1 U13639 ( .IN1(g1559), .IN2(n13536), .Q(n13533) );
  OR2X1 U13640 ( .IN1(n10500), .IN2(g1564), .Q(n13536) );
  AND2X1 U13641 ( .IN1(g1514), .IN2(n10568), .Q(n13532) );
  OR2X1 U13642 ( .IN1(n13537), .IN2(n13538), .Q(g33575) );
  OR2X1 U13643 ( .IN1(n13539), .IN2(n13540), .Q(n13538) );
  AND2X1 U13644 ( .IN1(n13541), .IN2(g2047), .Q(n13540) );
  OR2X1 U13645 ( .IN1(n13542), .IN2(n13293), .Q(n13541) );
  AND2X1 U13646 ( .IN1(n13543), .IN2(n10753), .Q(n13542) );
  INVX0 U13647 ( .INP(n3180), .ZN(n13539) );
  OR2X1 U13648 ( .IN1(n13544), .IN2(n13545), .Q(n3180) );
  OR2X1 U13649 ( .IN1(n13358), .IN2(g112), .Q(n13545) );
  INVX0 U13650 ( .INP(n12005), .ZN(n13358) );
  OR2X1 U13651 ( .IN1(n13543), .IN2(n12156), .Q(n13544) );
  OR2X1 U13652 ( .IN1(n12142), .IN2(n13546), .Q(n13543) );
  OR2X1 U13653 ( .IN1(n13547), .IN2(n13548), .Q(n13537) );
  AND2X1 U13654 ( .IN1(n13549), .IN2(n10753), .Q(n13548) );
  AND2X1 U13655 ( .IN1(n13550), .IN2(n13551), .Q(n13549) );
  INVX0 U13656 ( .INP(n13552), .ZN(n13551) );
  AND2X1 U13657 ( .IN1(n13553), .IN2(n13554), .Q(n13550) );
  OR2X1 U13658 ( .IN1(n10463), .IN2(n12156), .Q(n13554) );
  OR2X1 U13659 ( .IN1(n5535), .IN2(g2040), .Q(n12156) );
  INVX0 U13660 ( .INP(n13546), .ZN(n13553) );
  AND2X1 U13661 ( .IN1(n10915), .IN2(g1996), .Q(n13547) );
  OR2X1 U13662 ( .IN1(n13555), .IN2(n13556), .Q(g33574) );
  OR2X1 U13663 ( .IN1(n13557), .IN2(n13558), .Q(n13556) );
  AND2X1 U13664 ( .IN1(n10915), .IN2(g2112), .Q(n13558) );
  AND2X1 U13665 ( .IN1(n13559), .IN2(n10753), .Q(n13557) );
  AND2X1 U13666 ( .IN1(n5463), .IN2(n12739), .Q(n13559) );
  AND2X1 U13667 ( .IN1(n12738), .IN2(g2116), .Q(n13555) );
  OR2X1 U13668 ( .IN1(n13560), .IN2(n13561), .Q(g33573) );
  OR2X1 U13669 ( .IN1(n13562), .IN2(n13563), .Q(n13561) );
  AND2X1 U13670 ( .IN1(n13564), .IN2(n5452), .Q(n13563) );
  AND2X1 U13671 ( .IN1(n13565), .IN2(n5666), .Q(n13564) );
  AND2X1 U13672 ( .IN1(n12739), .IN2(n10753), .Q(n13565) );
  AND2X1 U13673 ( .IN1(n13566), .IN2(g2108), .Q(n13562) );
  OR2X1 U13674 ( .IN1(n10883), .IN2(n13567), .Q(n13566) );
  AND2X1 U13675 ( .IN1(n12739), .IN2(g2102), .Q(n13567) );
  AND2X1 U13676 ( .IN1(n12738), .IN2(g2112), .Q(n13560) );
  OR2X1 U13677 ( .IN1(n13568), .IN2(n13569), .Q(g33572) );
  AND2X1 U13678 ( .IN1(n13570), .IN2(g2102), .Q(n13569) );
  AND2X1 U13679 ( .IN1(n12738), .IN2(g2108), .Q(n13568) );
  OR2X1 U13680 ( .IN1(n13571), .IN2(n13572), .Q(g33571) );
  AND2X1 U13681 ( .IN1(n13570), .IN2(g2084), .Q(n13572) );
  AND2X1 U13682 ( .IN1(n12738), .IN2(g2089), .Q(n13571) );
  INVX0 U13683 ( .INP(n13570), .ZN(n12738) );
  OR2X1 U13684 ( .IN1(n10883), .IN2(n12739), .Q(n13570) );
  AND2X1 U13685 ( .IN1(n5535), .IN2(n13573), .Q(n12739) );
  AND2X1 U13686 ( .IN1(n12753), .IN2(n5355), .Q(n13573) );
  OR2X1 U13687 ( .IN1(n13574), .IN2(n13575), .Q(g33570) );
  OR2X1 U13688 ( .IN1(n13576), .IN2(n13577), .Q(n13575) );
  AND2X1 U13689 ( .IN1(n12773), .IN2(n13552), .Q(n13577) );
  AND2X1 U13690 ( .IN1(n12753), .IN2(g2040), .Q(n12773) );
  AND2X1 U13691 ( .IN1(n13578), .IN2(g2070), .Q(n13576) );
  AND2X1 U13692 ( .IN1(n10915), .IN2(g2040), .Q(n13574) );
  OR2X1 U13693 ( .IN1(n13579), .IN2(n13580), .Q(g33569) );
  OR2X1 U13694 ( .IN1(n13581), .IN2(n13582), .Q(n13580) );
  AND2X1 U13695 ( .IN1(n13583), .IN2(n10753), .Q(n13582) );
  AND2X1 U13696 ( .IN1(n12781), .IN2(n13552), .Q(n13583) );
  AND2X1 U13697 ( .IN1(n12753), .IN2(g1996), .Q(n12781) );
  AND2X1 U13698 ( .IN1(n10915), .IN2(g2047), .Q(n13581) );
  AND2X1 U13699 ( .IN1(n13578), .IN2(g2040), .Q(n13579) );
  OR2X1 U13700 ( .IN1(n13584), .IN2(n13585), .Q(g33568) );
  AND2X1 U13701 ( .IN1(n13578), .IN2(g1996), .Q(n13585) );
  AND2X1 U13702 ( .IN1(n10816), .IN2(n12748), .Q(n13578) );
  AND2X1 U13703 ( .IN1(n13586), .IN2(n13587), .Q(n13584) );
  AND2X1 U13704 ( .IN1(n13552), .IN2(n10753), .Q(n13587) );
  OR2X1 U13705 ( .IN1(n12142), .IN2(n13460), .Q(n13552) );
  OR2X1 U13706 ( .IN1(n11733), .IN2(n13588), .Q(n12142) );
  OR2X1 U13707 ( .IN1(n5287), .IN2(g504), .Q(n13588) );
  AND2X1 U13708 ( .IN1(n5535), .IN2(n13589), .Q(n13586) );
  OR2X1 U13709 ( .IN1(n13590), .IN2(g1996), .Q(n13589) );
  AND2X1 U13710 ( .IN1(n5505), .IN2(n12753), .Q(n13590) );
  INVX0 U13711 ( .INP(n12748), .ZN(n12753) );
  AND2X1 U13712 ( .IN1(n13546), .IN2(n12802), .Q(n12748) );
  INVX0 U13713 ( .INP(n12758), .ZN(n12802) );
  OR2X1 U13714 ( .IN1(n13591), .IN2(n13592), .Q(n12758) );
  OR2X1 U13715 ( .IN1(n13593), .IN2(n13594), .Q(n13592) );
  AND2X1 U13716 ( .IN1(n13595), .IN2(g2138), .Q(n13594) );
  AND2X1 U13717 ( .IN1(n5286), .IN2(g956), .Q(n13591) );
  OR2X1 U13718 ( .IN1(n13596), .IN2(n10388), .Q(n13546) );
  AND2X1 U13719 ( .IN1(n13597), .IN2(n5599), .Q(n13596) );
  AND2X1 U13720 ( .IN1(n5363), .IN2(n13598), .Q(n13597) );
  OR2X1 U13721 ( .IN1(n13599), .IN2(n13600), .Q(g33567) );
  OR2X1 U13722 ( .IN1(n13601), .IN2(n13602), .Q(n13600) );
  AND2X1 U13723 ( .IN1(n13603), .IN2(g1913), .Q(n13602) );
  OR2X1 U13724 ( .IN1(n13604), .IN2(n13293), .Q(n13603) );
  AND2X1 U13725 ( .IN1(n13605), .IN2(n10753), .Q(n13604) );
  OR2X1 U13726 ( .IN1(n12146), .IN2(n13606), .Q(n13605) );
  AND2X1 U13727 ( .IN1(n13607), .IN2(n13608), .Q(n13601) );
  OR2X1 U13728 ( .IN1(n13609), .IN2(n13610), .Q(n13608) );
  AND2X1 U13729 ( .IN1(n10463), .IN2(n13611), .Q(n13610) );
  OR2X1 U13730 ( .IN1(n13612), .IN2(n13613), .Q(n13611) );
  AND2X1 U13731 ( .IN1(n13614), .IN2(n10752), .Q(n13613) );
  AND2X1 U13732 ( .IN1(n13615), .IN2(n12161), .Q(n13612) );
  AND2X1 U13733 ( .IN1(n12162), .IN2(n12005), .Q(n13615) );
  AND2X1 U13734 ( .IN1(n13616), .IN2(n13614), .Q(n13609) );
  AND2X1 U13735 ( .IN1(n13617), .IN2(n10752), .Q(n13616) );
  INVX0 U13736 ( .INP(n12162), .ZN(n13617) );
  AND2X1 U13737 ( .IN1(g1936), .IN2(n5503), .Q(n12162) );
  INVX0 U13738 ( .INP(n13606), .ZN(n13607) );
  AND2X1 U13739 ( .IN1(test_so8), .IN2(n10896), .Q(n13599) );
  OR2X1 U13740 ( .IN1(n13618), .IN2(n13619), .Q(g33566) );
  OR2X1 U13741 ( .IN1(n13620), .IN2(n13621), .Q(n13619) );
  AND2X1 U13742 ( .IN1(n10915), .IN2(g1978), .Q(n13621) );
  AND2X1 U13743 ( .IN1(n13622), .IN2(n10752), .Q(n13620) );
  AND2X1 U13744 ( .IN1(n5462), .IN2(n12809), .Q(n13622) );
  AND2X1 U13745 ( .IN1(n12808), .IN2(g1982), .Q(n13618) );
  OR2X1 U13746 ( .IN1(n13623), .IN2(n13624), .Q(g33565) );
  OR2X1 U13747 ( .IN1(n13625), .IN2(n13626), .Q(n13624) );
  AND2X1 U13748 ( .IN1(n13627), .IN2(n5450), .Q(n13626) );
  AND2X1 U13749 ( .IN1(n13628), .IN2(n5664), .Q(n13627) );
  AND2X1 U13750 ( .IN1(n12809), .IN2(n10752), .Q(n13628) );
  AND2X1 U13751 ( .IN1(n13629), .IN2(g1974), .Q(n13625) );
  OR2X1 U13752 ( .IN1(n10883), .IN2(n13630), .Q(n13629) );
  AND2X1 U13753 ( .IN1(n12809), .IN2(g1968), .Q(n13630) );
  AND2X1 U13754 ( .IN1(n12808), .IN2(g1978), .Q(n13623) );
  OR2X1 U13755 ( .IN1(n13631), .IN2(n13632), .Q(g33564) );
  AND2X1 U13756 ( .IN1(n13633), .IN2(g1968), .Q(n13632) );
  AND2X1 U13757 ( .IN1(n12808), .IN2(g1974), .Q(n13631) );
  OR2X1 U13758 ( .IN1(n13634), .IN2(n13635), .Q(g33563) );
  AND2X1 U13759 ( .IN1(n13633), .IN2(g1950), .Q(n13635) );
  AND2X1 U13760 ( .IN1(n12808), .IN2(g1955), .Q(n13634) );
  INVX0 U13761 ( .INP(n13633), .ZN(n12808) );
  OR2X1 U13762 ( .IN1(n10883), .IN2(n12809), .Q(n13633) );
  AND2X1 U13763 ( .IN1(n5534), .IN2(n13636), .Q(n12809) );
  AND2X1 U13764 ( .IN1(n10570), .IN2(n12823), .Q(n13636) );
  OR2X1 U13765 ( .IN1(n13637), .IN2(n13638), .Q(g33562) );
  OR2X1 U13766 ( .IN1(n13639), .IN2(n13640), .Q(n13638) );
  AND2X1 U13767 ( .IN1(n12843), .IN2(n13641), .Q(n13640) );
  AND2X1 U13768 ( .IN1(n12823), .IN2(g1906), .Q(n12843) );
  AND2X1 U13769 ( .IN1(n13642), .IN2(g1936), .Q(n13639) );
  AND2X1 U13770 ( .IN1(n10915), .IN2(g1906), .Q(n13637) );
  OR2X1 U13771 ( .IN1(n13643), .IN2(n13644), .Q(g33561) );
  OR2X1 U13772 ( .IN1(n13645), .IN2(n13646), .Q(n13644) );
  AND2X1 U13773 ( .IN1(n13647), .IN2(n10752), .Q(n13646) );
  AND2X1 U13774 ( .IN1(n12851), .IN2(n13641), .Q(n13647) );
  AND2X1 U13775 ( .IN1(n12823), .IN2(test_so8), .Q(n12851) );
  AND2X1 U13776 ( .IN1(n10915), .IN2(g1913), .Q(n13645) );
  AND2X1 U13777 ( .IN1(n13642), .IN2(g1906), .Q(n13643) );
  OR2X1 U13778 ( .IN1(n13648), .IN2(n13649), .Q(g33560) );
  AND2X1 U13779 ( .IN1(n13642), .IN2(test_so8), .Q(n13649) );
  AND2X1 U13780 ( .IN1(n10815), .IN2(n12818), .Q(n13642) );
  AND2X1 U13781 ( .IN1(n13650), .IN2(n13651), .Q(n13648) );
  AND2X1 U13782 ( .IN1(n13641), .IN2(n10752), .Q(n13651) );
  INVX0 U13783 ( .INP(n13614), .ZN(n13641) );
  AND2X1 U13784 ( .IN1(n12161), .IN2(n3115), .Q(n13614) );
  INVX0 U13785 ( .INP(n12146), .ZN(n12161) );
  OR2X1 U13786 ( .IN1(n11733), .IN2(n13652), .Q(n12146) );
  OR2X1 U13787 ( .IN1(n5519), .IN2(n5287), .Q(n13652) );
  AND2X1 U13788 ( .IN1(n5534), .IN2(n13653), .Q(n13650) );
  OR2X1 U13789 ( .IN1(n13654), .IN2(test_so8), .Q(n13653) );
  AND2X1 U13790 ( .IN1(n5503), .IN2(n12823), .Q(n13654) );
  INVX0 U13791 ( .INP(n12818), .ZN(n12823) );
  AND2X1 U13792 ( .IN1(n13606), .IN2(n12871), .Q(n12818) );
  INVX0 U13793 ( .INP(n12828), .ZN(n12871) );
  OR2X1 U13794 ( .IN1(n13655), .IN2(n13656), .Q(n12828) );
  OR2X1 U13795 ( .IN1(n13593), .IN2(n13657), .Q(n13656) );
  AND2X1 U13796 ( .IN1(n13658), .IN2(n5307), .Q(n13657) );
  AND2X1 U13797 ( .IN1(g2138), .IN2(g2130), .Q(n13658) );
  AND2X1 U13798 ( .IN1(n5286), .IN2(g1129), .Q(n13655) );
  OR2X1 U13799 ( .IN1(n13659), .IN2(n10515), .Q(n13606) );
  AND2X1 U13800 ( .IN1(n13660), .IN2(n13598), .Q(n13659) );
  AND2X1 U13801 ( .IN1(g1171), .IN2(g1183), .Q(n13660) );
  OR2X1 U13802 ( .IN1(n13661), .IN2(n13662), .Q(g33559) );
  OR2X1 U13803 ( .IN1(n13663), .IN2(n13664), .Q(n13662) );
  AND2X1 U13804 ( .IN1(n13665), .IN2(g1779), .Q(n13664) );
  OR2X1 U13805 ( .IN1(n13666), .IN2(n13293), .Q(n13665) );
  AND2X1 U13806 ( .IN1(n13667), .IN2(n10752), .Q(n13666) );
  OR2X1 U13807 ( .IN1(n12145), .IN2(n13668), .Q(n13667) );
  AND2X1 U13808 ( .IN1(n13669), .IN2(n13670), .Q(n13663) );
  INVX0 U13809 ( .INP(n13668), .ZN(n13670) );
  AND2X1 U13810 ( .IN1(n13671), .IN2(n13672), .Q(n13669) );
  OR2X1 U13811 ( .IN1(g1772), .IN2(n13673), .Q(n13672) );
  OR2X1 U13812 ( .IN1(n5536), .IN2(n10463), .Q(n13673) );
  OR2X1 U13813 ( .IN1(n13674), .IN2(n13675), .Q(n13671) );
  AND2X1 U13814 ( .IN1(n13676), .IN2(n10752), .Q(n13675) );
  INVX0 U13815 ( .INP(n13677), .ZN(n13676) );
  AND2X1 U13816 ( .IN1(n12165), .IN2(n12005), .Q(n13674) );
  AND2X1 U13817 ( .IN1(n5504), .IN2(n13678), .Q(n12165) );
  AND2X1 U13818 ( .IN1(g1802), .IN2(n13679), .Q(n13678) );
  INVX0 U13819 ( .INP(n12145), .ZN(n13679) );
  AND2X1 U13820 ( .IN1(n10915), .IN2(g1728), .Q(n13661) );
  OR2X1 U13821 ( .IN1(n13680), .IN2(n13681), .Q(g33558) );
  OR2X1 U13822 ( .IN1(n13682), .IN2(n13683), .Q(n13681) );
  AND2X1 U13823 ( .IN1(n10915), .IN2(g1844), .Q(n13683) );
  AND2X1 U13824 ( .IN1(n13684), .IN2(n10752), .Q(n13682) );
  AND2X1 U13825 ( .IN1(n5464), .IN2(n12877), .Q(n13684) );
  AND2X1 U13826 ( .IN1(n12876), .IN2(g1848), .Q(n13680) );
  OR2X1 U13827 ( .IN1(n13685), .IN2(n13686), .Q(g33557) );
  OR2X1 U13828 ( .IN1(n13687), .IN2(n13688), .Q(n13686) );
  AND2X1 U13829 ( .IN1(n13689), .IN2(n5451), .Q(n13688) );
  AND2X1 U13830 ( .IN1(n13690), .IN2(n5665), .Q(n13689) );
  AND2X1 U13831 ( .IN1(n12877), .IN2(n10751), .Q(n13690) );
  AND2X1 U13832 ( .IN1(n13691), .IN2(g1840), .Q(n13687) );
  OR2X1 U13833 ( .IN1(n10883), .IN2(n13692), .Q(n13691) );
  AND2X1 U13834 ( .IN1(n12877), .IN2(g1834), .Q(n13692) );
  AND2X1 U13835 ( .IN1(n12876), .IN2(g1844), .Q(n13685) );
  OR2X1 U13836 ( .IN1(n13693), .IN2(n13694), .Q(g33556) );
  AND2X1 U13837 ( .IN1(n13695), .IN2(g1834), .Q(n13694) );
  AND2X1 U13838 ( .IN1(n12876), .IN2(g1840), .Q(n13693) );
  OR2X1 U13839 ( .IN1(n13696), .IN2(n13697), .Q(g33555) );
  AND2X1 U13840 ( .IN1(n13695), .IN2(g1816), .Q(n13697) );
  AND2X1 U13841 ( .IN1(n12876), .IN2(g1821), .Q(n13696) );
  INVX0 U13842 ( .INP(n13695), .ZN(n12876) );
  OR2X1 U13843 ( .IN1(n10883), .IN2(n12877), .Q(n13695) );
  AND2X1 U13844 ( .IN1(n5536), .IN2(n13698), .Q(n12877) );
  AND2X1 U13845 ( .IN1(n12891), .IN2(n5352), .Q(n13698) );
  OR2X1 U13846 ( .IN1(n13699), .IN2(n13700), .Q(g33554) );
  OR2X1 U13847 ( .IN1(n13701), .IN2(n13702), .Q(n13700) );
  AND2X1 U13848 ( .IN1(n12912), .IN2(n13677), .Q(n13702) );
  AND2X1 U13849 ( .IN1(n12891), .IN2(g1772), .Q(n12912) );
  AND2X1 U13850 ( .IN1(n13703), .IN2(g1802), .Q(n13701) );
  AND2X1 U13851 ( .IN1(n10915), .IN2(g1772), .Q(n13699) );
  OR2X1 U13852 ( .IN1(n13704), .IN2(n13705), .Q(g33553) );
  OR2X1 U13853 ( .IN1(n13706), .IN2(n13707), .Q(n13705) );
  AND2X1 U13854 ( .IN1(n13708), .IN2(n10751), .Q(n13707) );
  AND2X1 U13855 ( .IN1(n13709), .IN2(n12891), .Q(n13708) );
  AND2X1 U13856 ( .IN1(n13677), .IN2(g1728), .Q(n13709) );
  AND2X1 U13857 ( .IN1(n10915), .IN2(g1779), .Q(n13706) );
  AND2X1 U13858 ( .IN1(n13703), .IN2(g1772), .Q(n13704) );
  OR2X1 U13859 ( .IN1(n13710), .IN2(n13711), .Q(g33552) );
  AND2X1 U13860 ( .IN1(n13703), .IN2(g1728), .Q(n13711) );
  AND2X1 U13861 ( .IN1(n10817), .IN2(n12886), .Q(n13703) );
  AND2X1 U13862 ( .IN1(n13712), .IN2(n13713), .Q(n13710) );
  AND2X1 U13863 ( .IN1(n13677), .IN2(n10751), .Q(n13713) );
  OR2X1 U13864 ( .IN1(n12145), .IN2(n13460), .Q(n13677) );
  OR2X1 U13865 ( .IN1(n11733), .IN2(n13461), .Q(n12145) );
  OR2X1 U13866 ( .IN1(n5519), .IN2(g518), .Q(n13461) );
  AND2X1 U13867 ( .IN1(n5536), .IN2(n13714), .Q(n13712) );
  OR2X1 U13868 ( .IN1(n13715), .IN2(g1728), .Q(n13714) );
  AND2X1 U13869 ( .IN1(n5504), .IN2(n12891), .Q(n13715) );
  INVX0 U13870 ( .INP(n12886), .ZN(n12891) );
  AND2X1 U13871 ( .IN1(n13668), .IN2(n12939), .Q(n12886) );
  INVX0 U13872 ( .INP(n12896), .ZN(n12939) );
  OR2X1 U13873 ( .IN1(n13716), .IN2(n13717), .Q(n12896) );
  OR2X1 U13874 ( .IN1(n13593), .IN2(n13718), .Q(n13717) );
  AND2X1 U13875 ( .IN1(n13595), .IN2(n5275), .Q(n13718) );
  AND2X1 U13876 ( .IN1(g2145), .IN2(g2130), .Q(n13595) );
  AND2X1 U13877 ( .IN1(n5286), .IN2(g1105), .Q(n13716) );
  OR2X1 U13878 ( .IN1(n13719), .IN2(n10574), .Q(n13668) );
  AND2X1 U13879 ( .IN1(n13720), .IN2(n13598), .Q(n13719) );
  OR2X1 U13880 ( .IN1(n13721), .IN2(n13722), .Q(g33551) );
  OR2X1 U13881 ( .IN1(n13723), .IN2(n13724), .Q(n13722) );
  AND2X1 U13882 ( .IN1(test_so75), .IN2(n13293), .Q(n13724) );
  AND2X1 U13883 ( .IN1(n13725), .IN2(n13726), .Q(n13723) );
  AND2X1 U13884 ( .IN1(n13727), .IN2(n12154), .Q(n13726) );
  INVX0 U13885 ( .INP(n12147), .ZN(n12154) );
  AND2X1 U13886 ( .IN1(n10463), .IN2(n12005), .Q(n13727) );
  AND2X1 U13887 ( .IN1(g33533), .IN2(g31862), .Q(n13725) );
  OR2X1 U13888 ( .IN1(n13728), .IN2(n13729), .Q(n13721) );
  AND2X1 U13889 ( .IN1(n13730), .IN2(n10751), .Q(n13729) );
  OR2X1 U13890 ( .IN1(n13731), .IN2(n13732), .Q(n13730) );
  AND2X1 U13891 ( .IN1(test_so75), .IN2(n13733), .Q(n13732) );
  OR2X1 U13892 ( .IN1(n12147), .IN2(n13734), .Q(n13733) );
  INVX0 U13893 ( .INP(n13735), .ZN(n13731) );
  OR2X1 U13894 ( .IN1(n13736), .IN2(n13737), .Q(n13735) );
  OR2X1 U13895 ( .IN1(n13734), .IN2(n13738), .Q(n13736) );
  AND2X1 U13896 ( .IN1(g112), .IN2(g31862), .Q(n13738) );
  AND2X1 U13897 ( .IN1(n10915), .IN2(g1592), .Q(n13728) );
  OR2X1 U13898 ( .IN1(n13739), .IN2(n13740), .Q(g33550) );
  OR2X1 U13899 ( .IN1(n13741), .IN2(n13742), .Q(n13740) );
  AND2X1 U13900 ( .IN1(n10915), .IN2(g1710), .Q(n13742) );
  AND2X1 U13901 ( .IN1(n13743), .IN2(n10751), .Q(n13741) );
  AND2X1 U13902 ( .IN1(n5460), .IN2(n12946), .Q(n13743) );
  AND2X1 U13903 ( .IN1(n12945), .IN2(g1714), .Q(n13739) );
  OR2X1 U13904 ( .IN1(n13744), .IN2(n13745), .Q(g33549) );
  OR2X1 U13905 ( .IN1(n13746), .IN2(n13747), .Q(n13745) );
  AND2X1 U13906 ( .IN1(n13748), .IN2(n10587), .Q(n13747) );
  AND2X1 U13907 ( .IN1(n13749), .IN2(n5417), .Q(n13748) );
  AND2X1 U13908 ( .IN1(n12946), .IN2(n10751), .Q(n13749) );
  AND2X1 U13909 ( .IN1(test_so15), .IN2(n13750), .Q(n13746) );
  OR2X1 U13910 ( .IN1(n10883), .IN2(n13751), .Q(n13750) );
  AND2X1 U13911 ( .IN1(n12946), .IN2(g1700), .Q(n13751) );
  AND2X1 U13912 ( .IN1(n12945), .IN2(g1710), .Q(n13744) );
  OR2X1 U13913 ( .IN1(n13752), .IN2(n13753), .Q(g33548) );
  AND2X1 U13914 ( .IN1(n13754), .IN2(g1700), .Q(n13753) );
  AND2X1 U13915 ( .IN1(test_so15), .IN2(n12945), .Q(n13752) );
  OR2X1 U13916 ( .IN1(n13755), .IN2(n13756), .Q(g33547) );
  AND2X1 U13917 ( .IN1(n13754), .IN2(g1682), .Q(n13756) );
  AND2X1 U13918 ( .IN1(n12945), .IN2(g1687), .Q(n13755) );
  INVX0 U13919 ( .INP(n13754), .ZN(n12945) );
  OR2X1 U13920 ( .IN1(n10882), .IN2(n12946), .Q(n13754) );
  AND2X1 U13921 ( .IN1(n5598), .IN2(n13757), .Q(n12946) );
  AND2X1 U13922 ( .IN1(n12960), .IN2(n5362), .Q(n13757) );
  OR2X1 U13923 ( .IN1(n13758), .IN2(n13759), .Q(g33546) );
  OR2X1 U13924 ( .IN1(n13760), .IN2(n13761), .Q(n13759) );
  AND2X1 U13925 ( .IN1(n12980), .IN2(n13737), .Q(n13761) );
  AND2X1 U13926 ( .IN1(n12960), .IN2(g1636), .Q(n12980) );
  AND2X1 U13927 ( .IN1(n13762), .IN2(g1668), .Q(n13760) );
  AND2X1 U13928 ( .IN1(n10915), .IN2(g1636), .Q(n13758) );
  OR2X1 U13929 ( .IN1(n13763), .IN2(n13764), .Q(g33545) );
  OR2X1 U13930 ( .IN1(n13765), .IN2(n13766), .Q(n13764) );
  AND2X1 U13931 ( .IN1(n13767), .IN2(n10751), .Q(n13766) );
  AND2X1 U13932 ( .IN1(n12988), .IN2(n13737), .Q(n13767) );
  AND2X1 U13933 ( .IN1(n12960), .IN2(g1592), .Q(n12988) );
  AND2X1 U13934 ( .IN1(test_so75), .IN2(n10895), .Q(n13765) );
  AND2X1 U13935 ( .IN1(n13762), .IN2(g1636), .Q(n13763) );
  OR2X1 U13936 ( .IN1(n13768), .IN2(n13769), .Q(g33544) );
  AND2X1 U13937 ( .IN1(n13762), .IN2(g1592), .Q(n13769) );
  AND2X1 U13938 ( .IN1(n10818), .IN2(n12955), .Q(n13762) );
  AND2X1 U13939 ( .IN1(n13770), .IN2(n13771), .Q(n13768) );
  AND2X1 U13940 ( .IN1(n13737), .IN2(n10751), .Q(n13771) );
  OR2X1 U13941 ( .IN1(n12147), .IN2(n13460), .Q(n13737) );
  INVX0 U13942 ( .INP(n3115), .ZN(n13460) );
  OR2X1 U13943 ( .IN1(n11733), .IN2(n13521), .Q(n12147) );
  OR2X1 U13944 ( .IN1(g518), .IN2(g504), .Q(n13521) );
  INVX0 U13945 ( .INP(n3195), .ZN(n11733) );
  AND2X1 U13946 ( .IN1(n5598), .IN2(n13772), .Q(n13770) );
  OR2X1 U13947 ( .IN1(n13773), .IN2(g1592), .Q(n13772) );
  AND2X1 U13948 ( .IN1(n5549), .IN2(n12960), .Q(n13773) );
  INVX0 U13949 ( .INP(n12955), .ZN(n12960) );
  AND2X1 U13950 ( .IN1(n13734), .IN2(n13008), .Q(n12955) );
  INVX0 U13951 ( .INP(n12965), .ZN(n13008) );
  OR2X1 U13952 ( .IN1(n13774), .IN2(n13775), .Q(n12965) );
  OR2X1 U13953 ( .IN1(n13593), .IN2(n13776), .Q(n13775) );
  AND2X1 U13954 ( .IN1(n13777), .IN2(n5275), .Q(n13776) );
  AND2X1 U13955 ( .IN1(n5307), .IN2(g2130), .Q(n13777) );
  INVX0 U13956 ( .INP(n13009), .ZN(n13593) );
  OR2X1 U13957 ( .IN1(n13778), .IN2(g134), .Q(n13009) );
  AND2X1 U13958 ( .IN1(n13779), .IN2(n5595), .Q(n13778) );
  AND2X1 U13959 ( .IN1(n13780), .IN2(g691), .Q(n13779) );
  AND2X1 U13960 ( .IN1(n5286), .IN2(g1135), .Q(n13774) );
  OR2X1 U13961 ( .IN1(n13781), .IN2(n13782), .Q(g33543) );
  AND2X1 U13962 ( .IN1(n13783), .IN2(g1373), .Q(n13782) );
  OR2X1 U13963 ( .IN1(n10882), .IN2(n13784), .Q(n13783) );
  AND2X1 U13964 ( .IN1(n13785), .IN2(n10089), .Q(n13784) );
  AND2X1 U13965 ( .IN1(n13786), .IN2(n13787), .Q(n13785) );
  AND2X1 U13966 ( .IN1(n13788), .IN2(n13789), .Q(n13781) );
  OR2X1 U13967 ( .IN1(n13790), .IN2(n13791), .Q(n13789) );
  AND2X1 U13968 ( .IN1(n10462), .IN2(n13787), .Q(n13790) );
  AND2X1 U13969 ( .IN1(n10818), .IN2(g1379), .Q(n13788) );
  OR2X1 U13970 ( .IN1(n13792), .IN2(n13793), .Q(g33542) );
  OR2X1 U13971 ( .IN1(n13794), .IN2(n13795), .Q(n13793) );
  AND2X1 U13972 ( .IN1(n5730), .IN2(n13796), .Q(n13795) );
  INVX0 U13973 ( .INP(n13797), .ZN(n13794) );
  OR2X1 U13974 ( .IN1(n13798), .IN2(n5730), .Q(n13797) );
  OR2X1 U13975 ( .IN1(n13799), .IN2(n13796), .Q(n13798) );
  AND2X1 U13976 ( .IN1(n10915), .IN2(g1270), .Q(n13792) );
  OR2X1 U13977 ( .IN1(n13800), .IN2(n13801), .Q(g33541) );
  AND2X1 U13978 ( .IN1(n13802), .IN2(g1030), .Q(n13801) );
  OR2X1 U13979 ( .IN1(n10882), .IN2(n13803), .Q(n13802) );
  AND2X1 U13980 ( .IN1(n13804), .IN2(n10090), .Q(n13803) );
  AND2X1 U13981 ( .IN1(n13805), .IN2(n13806), .Q(n13804) );
  AND2X1 U13982 ( .IN1(n13807), .IN2(n13808), .Q(n13800) );
  OR2X1 U13983 ( .IN1(n13809), .IN2(n13810), .Q(n13808) );
  AND2X1 U13984 ( .IN1(n10461), .IN2(n13806), .Q(n13809) );
  AND2X1 U13985 ( .IN1(n10818), .IN2(g1036), .Q(n13807) );
  OR2X1 U13986 ( .IN1(n13811), .IN2(n13812), .Q(g33540) );
  OR2X1 U13987 ( .IN1(n13813), .IN2(n13814), .Q(n13812) );
  AND2X1 U13988 ( .IN1(n5731), .IN2(n13815), .Q(n13814) );
  INVX0 U13989 ( .INP(n13816), .ZN(n13813) );
  OR2X1 U13990 ( .IN1(n13817), .IN2(n5731), .Q(n13816) );
  OR2X1 U13991 ( .IN1(n13818), .IN2(n13815), .Q(n13817) );
  AND2X1 U13992 ( .IN1(n10916), .IN2(g925), .Q(n13811) );
  OR2X1 U13993 ( .IN1(n13819), .IN2(n13820), .Q(g33539) );
  OR2X1 U13994 ( .IN1(n13821), .IN2(n13822), .Q(n13820) );
  AND2X1 U13995 ( .IN1(n2980), .IN2(n5332), .Q(n13822) );
  AND2X1 U13996 ( .IN1(n13823), .IN2(g763), .Q(n13821) );
  AND2X1 U13997 ( .IN1(n2404), .IN2(n13824), .Q(n13823) );
  INVX0 U13998 ( .INP(n2980), .ZN(n13824) );
  AND2X1 U13999 ( .IN1(n10916), .IN2(g758), .Q(n13819) );
  OR2X1 U14000 ( .IN1(n13825), .IN2(n13826), .Q(g33538) );
  OR2X1 U14001 ( .IN1(n13827), .IN2(n13828), .Q(n13826) );
  AND2X1 U14002 ( .IN1(n2982), .IN2(n5476), .Q(n13828) );
  AND2X1 U14003 ( .IN1(n13829), .IN2(g595), .Q(n13827) );
  AND2X1 U14004 ( .IN1(n2421), .IN2(n13830), .Q(n13829) );
  INVX0 U14005 ( .INP(n2982), .ZN(n13830) );
  AND2X1 U14006 ( .IN1(n10916), .IN2(g590), .Q(n13825) );
  OR2X1 U14007 ( .IN1(n13831), .IN2(n13832), .Q(g33537) );
  AND2X1 U14008 ( .IN1(n13833), .IN2(n10751), .Q(n13832) );
  AND2X1 U14009 ( .IN1(n2707), .IN2(g142), .Q(n13833) );
  AND2X1 U14010 ( .IN1(n10929), .IN2(g301), .Q(n13831) );
  AND2X1 U14011 ( .IN1(n13834), .IN2(g160), .Q(g33536) );
  OR2X1 U14012 ( .IN1(n2710), .IN2(n10875), .Q(n13834) );
  OR2X1 U14013 ( .IN1(n13835), .IN2(n13836), .Q(g33535) );
  OR2X1 U14014 ( .IN1(n13837), .IN2(n13838), .Q(n13836) );
  AND2X1 U14015 ( .IN1(n3276), .IN2(n5680), .Q(n13838) );
  AND2X1 U14016 ( .IN1(n13839), .IN2(g294), .Q(n13837) );
  AND2X1 U14017 ( .IN1(n10534), .IN2(n13840), .Q(n13839) );
  INVX0 U14018 ( .INP(n3276), .ZN(n13840) );
  AND2X1 U14019 ( .IN1(n10927), .IN2(g291), .Q(n13835) );
  OR2X1 U14020 ( .IN1(n13841), .IN2(n13842), .Q(g33534) );
  OR2X1 U14021 ( .IN1(n13843), .IN2(n13844), .Q(n13842) );
  AND2X1 U14022 ( .IN1(n3277), .IN2(n5677), .Q(n13844) );
  AND2X1 U14023 ( .IN1(n13845), .IN2(g153), .Q(n13843) );
  AND2X1 U14024 ( .IN1(n13055), .IN2(n13846), .Q(n13845) );
  INVX0 U14025 ( .INP(n3277), .ZN(n13846) );
  AND2X1 U14026 ( .IN1(n10927), .IN2(g150), .Q(n13841) );
  INVX0 U14027 ( .INP(n13734), .ZN(g33533) );
  OR2X1 U14028 ( .IN1(n13847), .IN2(n10111), .Q(n13734) );
  AND2X1 U14029 ( .IN1(n13848), .IN2(n5599), .Q(n13847) );
  AND2X1 U14030 ( .IN1(n13598), .IN2(g1171), .Q(n13848) );
  INVX0 U14031 ( .INP(n13849), .ZN(n13598) );
  OR2X1 U14032 ( .IN1(n13850), .IN2(n13851), .Q(n13849) );
  OR2X1 U14033 ( .IN1(g1205), .IN2(n13852), .Q(n13851) );
  OR2X1 U14034 ( .IN1(g1221), .IN2(g1216), .Q(n13852) );
  OR2X1 U14035 ( .IN1(n10499), .IN2(n13853), .Q(n13850) );
  OR2X1 U14036 ( .IN1(test_so76), .IN2(n5320), .Q(n13853) );
  AND2X1 U14037 ( .IN1(n13854), .IN2(n13855), .Q(g33435) );
  OR2X1 U14038 ( .IN1(n5610), .IN2(n12042), .Q(n13855) );
  AND2X1 U14039 ( .IN1(n13856), .IN2(n13857), .Q(n13854) );
  OR2X1 U14040 ( .IN1(g2729), .IN2(n13858), .Q(n13857) );
  OR2X1 U14041 ( .IN1(n13859), .IN2(n13860), .Q(n13858) );
  AND2X1 U14042 ( .IN1(n5544), .IN2(n5301), .Q(n13860) );
  AND2X1 U14043 ( .IN1(n5378), .IN2(g2724), .Q(n13859) );
  OR2X1 U14044 ( .IN1(n5403), .IN2(n12062), .Q(n13856) );
  AND2X1 U14045 ( .IN1(n13861), .IN2(n13862), .Q(g33079) );
  OR2X1 U14046 ( .IN1(n5609), .IN2(n12042), .Q(n13862) );
  AND2X1 U14047 ( .IN1(n13863), .IN2(n13864), .Q(n13861) );
  OR2X1 U14048 ( .IN1(g2729), .IN2(n13865), .Q(n13864) );
  OR2X1 U14049 ( .IN1(n13866), .IN2(n13867), .Q(n13865) );
  AND2X1 U14050 ( .IN1(n5545), .IN2(n5301), .Q(n13867) );
  AND2X1 U14051 ( .IN1(n5379), .IN2(g2724), .Q(n13866) );
  OR2X1 U14052 ( .IN1(n5404), .IN2(n12062), .Q(n13863) );
  OR2X1 U14053 ( .IN1(n10520), .IN2(g2724), .Q(n12062) );
  OR2X1 U14054 ( .IN1(n13868), .IN2(n13869), .Q(g33070) );
  AND2X1 U14055 ( .IN1(n10927), .IN2(g6565), .Q(n13869) );
  AND2X1 U14056 ( .IN1(n13870), .IN2(n13871), .Q(n13868) );
  OR2X1 U14057 ( .IN1(n13872), .IN2(n13873), .Q(n13870) );
  OR2X1 U14058 ( .IN1(n13874), .IN2(n13875), .Q(n13873) );
  AND2X1 U14059 ( .IN1(g25756), .IN2(n5646), .Q(n13875) );
  AND2X1 U14060 ( .IN1(n10818), .IN2(n13876), .Q(n13872) );
  OR2X1 U14061 ( .IN1(n13877), .IN2(n13878), .Q(g33069) );
  AND2X1 U14062 ( .IN1(n13879), .IN2(g6565), .Q(n13878) );
  AND2X1 U14063 ( .IN1(n13880), .IN2(g6561), .Q(n13877) );
  OR2X1 U14064 ( .IN1(n10882), .IN2(n13881), .Q(n13880) );
  AND2X1 U14065 ( .IN1(n5386), .IN2(n13871), .Q(n13881) );
  OR2X1 U14066 ( .IN1(n13882), .IN2(n13883), .Q(g33068) );
  AND2X1 U14067 ( .IN1(n10927), .IN2(g6555), .Q(n13883) );
  AND2X1 U14068 ( .IN1(n13884), .IN2(n5646), .Q(n13882) );
  AND2X1 U14069 ( .IN1(n13871), .IN2(n13885), .Q(n13884) );
  OR2X1 U14070 ( .IN1(n13886), .IN2(n13887), .Q(g33067) );
  AND2X1 U14071 ( .IN1(n10927), .IN2(g6549), .Q(n13887) );
  AND2X1 U14072 ( .IN1(n13888), .IN2(n13871), .Q(n13886) );
  INVX0 U14073 ( .INP(n13889), .ZN(n13888) );
  AND2X1 U14074 ( .IN1(n13890), .IN2(n3407), .Q(n13889) );
  OR2X1 U14075 ( .IN1(n10881), .IN2(n3406), .Q(n13890) );
  OR2X1 U14076 ( .IN1(n13891), .IN2(n13892), .Q(g33065) );
  AND2X1 U14077 ( .IN1(n10927), .IN2(g6219), .Q(n13892) );
  AND2X1 U14078 ( .IN1(n13893), .IN2(n13894), .Q(n13891) );
  OR2X1 U14079 ( .IN1(n13895), .IN2(n13896), .Q(n13893) );
  OR2X1 U14080 ( .IN1(n13897), .IN2(n13898), .Q(n13896) );
  AND2X1 U14081 ( .IN1(g25742), .IN2(n5651), .Q(n13898) );
  AND2X1 U14082 ( .IN1(n10819), .IN2(n13899), .Q(n13895) );
  OR2X1 U14083 ( .IN1(n13900), .IN2(n13901), .Q(g33064) );
  AND2X1 U14084 ( .IN1(n13902), .IN2(g6219), .Q(n13901) );
  AND2X1 U14085 ( .IN1(n13903), .IN2(g6215), .Q(n13900) );
  OR2X1 U14086 ( .IN1(n10881), .IN2(n13904), .Q(n13903) );
  AND2X1 U14087 ( .IN1(n5385), .IN2(n13894), .Q(n13904) );
  OR2X1 U14088 ( .IN1(n13905), .IN2(n13906), .Q(g33063) );
  AND2X1 U14089 ( .IN1(n10927), .IN2(g6209), .Q(n13906) );
  AND2X1 U14090 ( .IN1(n13907), .IN2(n5651), .Q(n13905) );
  AND2X1 U14091 ( .IN1(n13894), .IN2(n13908), .Q(n13907) );
  OR2X1 U14092 ( .IN1(n13909), .IN2(n13910), .Q(g33062) );
  AND2X1 U14093 ( .IN1(n10927), .IN2(g6203), .Q(n13910) );
  AND2X1 U14094 ( .IN1(n13911), .IN2(n13894), .Q(n13909) );
  INVX0 U14095 ( .INP(n13912), .ZN(n13911) );
  AND2X1 U14096 ( .IN1(n13913), .IN2(n3417), .Q(n13912) );
  OR2X1 U14097 ( .IN1(n10880), .IN2(n3416), .Q(n13913) );
  OR2X1 U14098 ( .IN1(n13914), .IN2(n13915), .Q(g33060) );
  AND2X1 U14099 ( .IN1(n10927), .IN2(g5873), .Q(n13915) );
  AND2X1 U14100 ( .IN1(n13916), .IN2(n13917), .Q(n13914) );
  OR2X1 U14101 ( .IN1(n13918), .IN2(n13919), .Q(n13916) );
  OR2X1 U14102 ( .IN1(n13920), .IN2(n13921), .Q(n13919) );
  AND2X1 U14103 ( .IN1(g25728), .IN2(n5649), .Q(n13921) );
  AND2X1 U14104 ( .IN1(n10819), .IN2(n13922), .Q(n13918) );
  OR2X1 U14105 ( .IN1(n13923), .IN2(n13924), .Q(g33059) );
  AND2X1 U14106 ( .IN1(n13925), .IN2(g5873), .Q(n13924) );
  AND2X1 U14107 ( .IN1(n13926), .IN2(g5869), .Q(n13923) );
  OR2X1 U14108 ( .IN1(n10879), .IN2(n13927), .Q(n13926) );
  AND2X1 U14109 ( .IN1(n5388), .IN2(n13917), .Q(n13927) );
  OR2X1 U14110 ( .IN1(n13928), .IN2(n13929), .Q(g33058) );
  AND2X1 U14111 ( .IN1(n10927), .IN2(g5863), .Q(n13929) );
  AND2X1 U14112 ( .IN1(n13930), .IN2(n5649), .Q(n13928) );
  AND2X1 U14113 ( .IN1(n13917), .IN2(n13931), .Q(n13930) );
  OR2X1 U14114 ( .IN1(n13932), .IN2(n13933), .Q(g33057) );
  AND2X1 U14115 ( .IN1(n10927), .IN2(g5857), .Q(n13933) );
  AND2X1 U14116 ( .IN1(n13934), .IN2(n13917), .Q(n13932) );
  INVX0 U14117 ( .INP(n13935), .ZN(n13934) );
  AND2X1 U14118 ( .IN1(n13936), .IN2(n3427), .Q(n13935) );
  OR2X1 U14119 ( .IN1(n10880), .IN2(n3426), .Q(n13936) );
  OR2X1 U14120 ( .IN1(n13937), .IN2(n13938), .Q(g33055) );
  AND2X1 U14121 ( .IN1(n10927), .IN2(g5527), .Q(n13938) );
  AND2X1 U14122 ( .IN1(n13939), .IN2(n13940), .Q(n13937) );
  OR2X1 U14123 ( .IN1(n13941), .IN2(n13942), .Q(n13939) );
  OR2X1 U14124 ( .IN1(n13943), .IN2(n13944), .Q(n13942) );
  AND2X1 U14125 ( .IN1(g25714), .IN2(n5647), .Q(n13944) );
  AND2X1 U14126 ( .IN1(n10819), .IN2(n13945), .Q(n13941) );
  OR2X1 U14127 ( .IN1(n13946), .IN2(n13947), .Q(g33054) );
  AND2X1 U14128 ( .IN1(n13948), .IN2(g5527), .Q(n13947) );
  AND2X1 U14129 ( .IN1(n13949), .IN2(g5523), .Q(n13946) );
  OR2X1 U14130 ( .IN1(n10879), .IN2(n13950), .Q(n13949) );
  AND2X1 U14131 ( .IN1(n5389), .IN2(n13940), .Q(n13950) );
  OR2X1 U14132 ( .IN1(n13951), .IN2(n13952), .Q(g33053) );
  AND2X1 U14133 ( .IN1(n10927), .IN2(g5517), .Q(n13952) );
  AND2X1 U14134 ( .IN1(n13953), .IN2(n5647), .Q(n13951) );
  AND2X1 U14135 ( .IN1(n13940), .IN2(n13954), .Q(n13953) );
  OR2X1 U14136 ( .IN1(n13955), .IN2(n13956), .Q(g33052) );
  AND2X1 U14137 ( .IN1(n10927), .IN2(g5511), .Q(n13956) );
  AND2X1 U14138 ( .IN1(n13957), .IN2(n13940), .Q(n13955) );
  INVX0 U14139 ( .INP(n13958), .ZN(n13957) );
  AND2X1 U14140 ( .IN1(n13959), .IN2(n3437), .Q(n13958) );
  OR2X1 U14141 ( .IN1(n10878), .IN2(n3436), .Q(n13959) );
  OR2X1 U14142 ( .IN1(n13960), .IN2(n13961), .Q(g33050) );
  AND2X1 U14143 ( .IN1(n10927), .IN2(g5180), .Q(n13961) );
  AND2X1 U14144 ( .IN1(n13962), .IN2(n13963), .Q(n13960) );
  OR2X1 U14145 ( .IN1(n13964), .IN2(n13965), .Q(n13962) );
  OR2X1 U14146 ( .IN1(n13966), .IN2(n13967), .Q(n13965) );
  AND2X1 U14147 ( .IN1(g25700), .IN2(n5650), .Q(n13967) );
  AND2X1 U14148 ( .IN1(n10819), .IN2(n13968), .Q(n13964) );
  OR2X1 U14149 ( .IN1(n13969), .IN2(n13970), .Q(g33049) );
  AND2X1 U14150 ( .IN1(n13971), .IN2(g5180), .Q(n13970) );
  AND2X1 U14151 ( .IN1(n13972), .IN2(g5176), .Q(n13969) );
  OR2X1 U14152 ( .IN1(n10878), .IN2(n13973), .Q(n13972) );
  AND2X1 U14153 ( .IN1(n5384), .IN2(n13963), .Q(n13973) );
  OR2X1 U14154 ( .IN1(n13974), .IN2(n13975), .Q(g33048) );
  AND2X1 U14155 ( .IN1(n10927), .IN2(g5170), .Q(n13975) );
  AND2X1 U14156 ( .IN1(n13976), .IN2(n5650), .Q(n13974) );
  AND2X1 U14157 ( .IN1(n13963), .IN2(n13977), .Q(n13976) );
  OR2X1 U14158 ( .IN1(n13978), .IN2(n13979), .Q(g33047) );
  AND2X1 U14159 ( .IN1(n10927), .IN2(g5164), .Q(n13979) );
  AND2X1 U14160 ( .IN1(n13980), .IN2(n13963), .Q(n13978) );
  INVX0 U14161 ( .INP(n13981), .ZN(n13980) );
  AND2X1 U14162 ( .IN1(n13982), .IN2(n3447), .Q(n13981) );
  OR2X1 U14163 ( .IN1(n10878), .IN2(n3446), .Q(n13982) );
  OR2X1 U14164 ( .IN1(n13983), .IN2(n13984), .Q(g33046) );
  OR2X1 U14165 ( .IN1(n13985), .IN2(n13986), .Q(n13984) );
  AND2X1 U14166 ( .IN1(n13987), .IN2(g5057), .Q(n13986) );
  AND2X1 U14167 ( .IN1(n13988), .IN2(n13989), .Q(n13987) );
  INVX0 U14168 ( .INP(n13990), .ZN(n13989) );
  AND2X1 U14169 ( .IN1(n5615), .IN2(n13991), .Q(n13985) );
  OR2X1 U14170 ( .IN1(n13990), .IN2(n13992), .Q(n13991) );
  AND2X1 U14171 ( .IN1(g5052), .IN2(n13993), .Q(n13990) );
  AND2X1 U14172 ( .IN1(n10927), .IN2(g5052), .Q(n13983) );
  OR2X1 U14173 ( .IN1(n13994), .IN2(n13995), .Q(g33045) );
  OR2X1 U14174 ( .IN1(n13996), .IN2(n13997), .Q(n13995) );
  AND2X1 U14175 ( .IN1(n13998), .IN2(g4567), .Q(n13994) );
  OR2X1 U14176 ( .IN1(n13997), .IN2(n13999), .Q(g33044) );
  OR2X1 U14177 ( .IN1(n14000), .IN2(n14001), .Q(n13999) );
  AND2X1 U14178 ( .IN1(test_so93), .IN2(n13998), .Q(n14001) );
  OR2X1 U14179 ( .IN1(n14002), .IN2(n14003), .Q(g33043) );
  OR2X1 U14180 ( .IN1(n14004), .IN2(n14005), .Q(n14003) );
  AND2X1 U14181 ( .IN1(test_so16), .IN2(n13998), .Q(n14002) );
  OR2X1 U14182 ( .IN1(n14006), .IN2(n14007), .Q(g33042) );
  OR2X1 U14183 ( .IN1(n14004), .IN2(n13997), .Q(n14007) );
  AND2X1 U14184 ( .IN1(g4578), .IN2(n14008), .Q(n13997) );
  AND2X1 U14185 ( .IN1(n13998), .IN2(g4540), .Q(n14006) );
  OR2X1 U14186 ( .IN1(n14009), .IN2(n14010), .Q(g33041) );
  OR2X1 U14187 ( .IN1(n13996), .IN2(n14005), .Q(n14010) );
  AND2X1 U14188 ( .IN1(test_so56), .IN2(n13998), .Q(n14009) );
  OR2X1 U14189 ( .IN1(n14011), .IN2(n14012), .Q(g33040) );
  OR2X1 U14190 ( .IN1(n14000), .IN2(n14013), .Q(n14012) );
  AND2X1 U14191 ( .IN1(n13998), .IN2(g4504), .Q(n14013) );
  AND2X1 U14192 ( .IN1(n14008), .IN2(n11594), .Q(n14000) );
  INVX0 U14193 ( .INP(n12429), .ZN(n11594) );
  AND2X1 U14194 ( .IN1(n11628), .IN2(n13030), .Q(n12429) );
  INVX0 U14195 ( .INP(g72), .ZN(n13030) );
  INVX0 U14196 ( .INP(g73), .ZN(n11628) );
  OR2X1 U14197 ( .IN1(n14014), .IN2(n14015), .Q(g33039) );
  OR2X1 U14198 ( .IN1(n13996), .IN2(n14016), .Q(n14015) );
  AND2X1 U14199 ( .IN1(n13998), .IN2(g4501), .Q(n14014) );
  OR2X1 U14200 ( .IN1(n14017), .IN2(n14018), .Q(g33038) );
  OR2X1 U14201 ( .IN1(n13996), .IN2(n14011), .Q(n14018) );
  AND2X1 U14202 ( .IN1(n14019), .IN2(n14008), .Q(n13996) );
  OR2X1 U14203 ( .IN1(n11205), .IN2(g73), .Q(n14019) );
  AND2X1 U14204 ( .IN1(n13998), .IN2(g4498), .Q(n14017) );
  OR2X1 U14205 ( .IN1(n14020), .IN2(n14021), .Q(g33037) );
  OR2X1 U14206 ( .IN1(n14004), .IN2(n14016), .Q(n14021) );
  AND2X1 U14207 ( .IN1(n13998), .IN2(g4495), .Q(n14020) );
  OR2X1 U14208 ( .IN1(n14022), .IN2(n14023), .Q(g33036) );
  OR2X1 U14209 ( .IN1(n14004), .IN2(n14011), .Q(n14023) );
  AND2X1 U14210 ( .IN1(g4572), .IN2(n14008), .Q(n14011) );
  AND2X1 U14211 ( .IN1(n14024), .IN2(n14008), .Q(n14004) );
  OR2X1 U14212 ( .IN1(n13097), .IN2(g72), .Q(n14024) );
  AND2X1 U14213 ( .IN1(n13998), .IN2(g4480), .Q(n14022) );
  INVX0 U14214 ( .INP(n14008), .ZN(n13998) );
  OR2X1 U14215 ( .IN1(n14025), .IN2(n14026), .Q(g33035) );
  OR2X1 U14216 ( .IN1(n10542), .IN2(n14027), .Q(n14026) );
  AND2X1 U14217 ( .IN1(n11208), .IN2(n5715), .Q(n14027) );
  INVX0 U14218 ( .INP(n11202), .ZN(n11208) );
  OR2X1 U14219 ( .IN1(n14028), .IN2(n14029), .Q(n14025) );
  AND2X1 U14220 ( .IN1(n10928), .IN2(g4098), .Q(n14029) );
  AND2X1 U14221 ( .IN1(n14030), .IN2(n10750), .Q(n14028) );
  AND2X1 U14222 ( .IN1(n11202), .IN2(g4108), .Q(n14030) );
  OR2X1 U14223 ( .IN1(n5350), .IN2(n14031), .Q(n11202) );
  OR2X1 U14224 ( .IN1(n14032), .IN2(n14033), .Q(g33034) );
  AND2X1 U14225 ( .IN1(n10928), .IN2(g3873), .Q(n14033) );
  AND2X1 U14226 ( .IN1(n14034), .IN2(n14035), .Q(n14032) );
  OR2X1 U14227 ( .IN1(n14036), .IN2(n14037), .Q(n14034) );
  OR2X1 U14228 ( .IN1(n14038), .IN2(n14039), .Q(n14037) );
  AND2X1 U14229 ( .IN1(g25676), .IN2(n10553), .Q(n14039) );
  AND2X1 U14230 ( .IN1(n10819), .IN2(n14040), .Q(n14036) );
  OR2X1 U14231 ( .IN1(n14041), .IN2(n14042), .Q(g33033) );
  AND2X1 U14232 ( .IN1(n14043), .IN2(g3873), .Q(n14042) );
  AND2X1 U14233 ( .IN1(test_so33), .IN2(n14044), .Q(n14041) );
  OR2X1 U14234 ( .IN1(n10879), .IN2(n14045), .Q(n14044) );
  AND2X1 U14235 ( .IN1(n5387), .IN2(n14035), .Q(n14045) );
  OR2X1 U14236 ( .IN1(n14046), .IN2(n14047), .Q(g33032) );
  AND2X1 U14237 ( .IN1(n10928), .IN2(g3863), .Q(n14047) );
  AND2X1 U14238 ( .IN1(n14048), .IN2(n14035), .Q(n14046) );
  AND2X1 U14239 ( .IN1(n14049), .IN2(n10553), .Q(n14048) );
  INVX0 U14240 ( .INP(n1075), .ZN(n14049) );
  OR2X1 U14241 ( .IN1(n14050), .IN2(n14051), .Q(g33031) );
  AND2X1 U14242 ( .IN1(n10928), .IN2(g3857), .Q(n14051) );
  AND2X1 U14243 ( .IN1(n14052), .IN2(n14035), .Q(n14050) );
  INVX0 U14244 ( .INP(n14053), .ZN(n14052) );
  AND2X1 U14245 ( .IN1(n14054), .IN2(n3482), .Q(n14053) );
  OR2X1 U14246 ( .IN1(n10878), .IN2(n3481), .Q(n14054) );
  OR2X1 U14247 ( .IN1(n14055), .IN2(n14056), .Q(g33029) );
  AND2X1 U14248 ( .IN1(n10928), .IN2(g3522), .Q(n14056) );
  AND2X1 U14249 ( .IN1(n14057), .IN2(n14058), .Q(n14055) );
  OR2X1 U14250 ( .IN1(n14059), .IN2(n14060), .Q(n14057) );
  OR2X1 U14251 ( .IN1(n14061), .IN2(n14062), .Q(n14060) );
  AND2X1 U14252 ( .IN1(g25662), .IN2(n5645), .Q(n14062) );
  AND2X1 U14253 ( .IN1(n10819), .IN2(n14063), .Q(n14059) );
  OR2X1 U14254 ( .IN1(n14064), .IN2(n14065), .Q(g33028) );
  AND2X1 U14255 ( .IN1(n14066), .IN2(g3522), .Q(n14065) );
  AND2X1 U14256 ( .IN1(n14067), .IN2(g3518), .Q(n14064) );
  OR2X1 U14257 ( .IN1(n10879), .IN2(n14068), .Q(n14067) );
  AND2X1 U14258 ( .IN1(n5383), .IN2(n14058), .Q(n14068) );
  OR2X1 U14259 ( .IN1(n14069), .IN2(n14070), .Q(g33027) );
  AND2X1 U14260 ( .IN1(n10928), .IN2(g3512), .Q(n14070) );
  AND2X1 U14261 ( .IN1(n14071), .IN2(n5645), .Q(n14069) );
  AND2X1 U14262 ( .IN1(n14058), .IN2(n14072), .Q(n14071) );
  OR2X1 U14263 ( .IN1(n14073), .IN2(n14074), .Q(g33026) );
  AND2X1 U14264 ( .IN1(n10928), .IN2(g3506), .Q(n14074) );
  AND2X1 U14265 ( .IN1(n14075), .IN2(n14058), .Q(n14073) );
  INVX0 U14266 ( .INP(n14076), .ZN(n14075) );
  AND2X1 U14267 ( .IN1(n14077), .IN2(n3492), .Q(n14076) );
  OR2X1 U14268 ( .IN1(n10877), .IN2(n3491), .Q(n14077) );
  OR2X1 U14269 ( .IN1(n14078), .IN2(n14079), .Q(g33024) );
  OR2X1 U14270 ( .IN1(n14080), .IN2(n14081), .Q(n14079) );
  AND2X1 U14271 ( .IN1(n14082), .IN2(n10750), .Q(n14081) );
  AND2X1 U14272 ( .IN1(n14083), .IN2(n14084), .Q(n14082) );
  OR2X1 U14273 ( .IN1(n14085), .IN2(n14086), .Q(n14083) );
  AND2X1 U14274 ( .IN1(n10928), .IN2(g3171), .Q(n14080) );
  AND2X1 U14275 ( .IN1(g25648), .IN2(n14087), .Q(n14078) );
  OR2X1 U14276 ( .IN1(n14088), .IN2(n14089), .Q(g33023) );
  AND2X1 U14277 ( .IN1(n14090), .IN2(g3167), .Q(n14089) );
  OR2X1 U14278 ( .IN1(n10878), .IN2(n14091), .Q(n14090) );
  AND2X1 U14279 ( .IN1(n5603), .IN2(n14084), .Q(n14091) );
  AND2X1 U14280 ( .IN1(n14092), .IN2(n14087), .Q(n14088) );
  AND2X1 U14281 ( .IN1(n10819), .IN2(g3171), .Q(n14092) );
  OR2X1 U14282 ( .IN1(n14093), .IN2(n14094), .Q(g33022) );
  AND2X1 U14283 ( .IN1(n10928), .IN2(g3161), .Q(n14094) );
  AND2X1 U14284 ( .IN1(n14087), .IN2(n14095), .Q(n14093) );
  OR2X1 U14285 ( .IN1(n14096), .IN2(n14097), .Q(g33021) );
  AND2X1 U14286 ( .IN1(n10928), .IN2(g3155), .Q(n14097) );
  AND2X1 U14287 ( .IN1(n14098), .IN2(n14084), .Q(n14096) );
  INVX0 U14288 ( .INP(n14099), .ZN(n14098) );
  AND2X1 U14289 ( .IN1(n14100), .IN2(n3501), .Q(n14099) );
  OR2X1 U14290 ( .IN1(n10877), .IN2(n3502), .Q(n14100) );
  OR2X1 U14291 ( .IN1(n2787), .IN2(n14101), .Q(g33019) );
  OR2X1 U14292 ( .IN1(n14102), .IN2(n14103), .Q(n14101) );
  AND2X1 U14293 ( .IN1(n14104), .IN2(n10750), .Q(n14103) );
  XOR2X1 U14294 ( .IN1(test_so30), .IN2(n2790), .Q(n14104) );
  AND2X1 U14295 ( .IN1(n10928), .IN2(g2748), .Q(n14102) );
  OR2X1 U14296 ( .IN1(n14105), .IN2(n14106), .Q(g33018) );
  OR2X1 U14297 ( .IN1(n14107), .IN2(n14108), .Q(n14106) );
  AND2X1 U14298 ( .IN1(test_so40), .IN2(n14109), .Q(n14108) );
  OR2X1 U14299 ( .IN1(n14110), .IN2(n14111), .Q(n14109) );
  OR2X1 U14300 ( .IN1(n13293), .IN2(n14112), .Q(n14111) );
  AND2X1 U14301 ( .IN1(n3006), .IN2(n10750), .Q(n14110) );
  INVX0 U14302 ( .INP(n12362), .ZN(n3006) );
  AND2X1 U14303 ( .IN1(n14113), .IN2(n3517), .Q(n14107) );
  AND2X1 U14304 ( .IN1(n3512), .IN2(n11218), .Q(n14113) );
  AND2X1 U14305 ( .IN1(n12362), .IN2(n3524), .Q(n11218) );
  AND2X1 U14306 ( .IN1(n1284), .IN2(n3525), .Q(n12362) );
  OR2X1 U14307 ( .IN1(g2610), .IN2(n14114), .Q(n3512) );
  OR2X1 U14308 ( .IN1(n5508), .IN2(n10531), .Q(n14114) );
  OR2X1 U14309 ( .IN1(n14115), .IN2(n14116), .Q(n14105) );
  AND2X1 U14310 ( .IN1(n14117), .IN2(n10468), .Q(n14116) );
  AND2X1 U14311 ( .IN1(n14118), .IN2(n14119), .Q(n14117) );
  AND2X1 U14312 ( .IN1(n14120), .IN2(g2619), .Q(n14119) );
  AND2X1 U14313 ( .IN1(n3511), .IN2(n12005), .Q(n14118) );
  AND2X1 U14314 ( .IN1(n10928), .IN2(g2610), .Q(n14115) );
  OR2X1 U14315 ( .IN1(n14121), .IN2(n14122), .Q(g33017) );
  OR2X1 U14316 ( .IN1(n14123), .IN2(n14124), .Q(n14122) );
  AND2X1 U14317 ( .IN1(test_so40), .IN2(n10895), .Q(n14124) );
  AND2X1 U14318 ( .IN1(n3517), .IN2(g2610), .Q(n14123) );
  OR2X1 U14319 ( .IN1(n3519), .IN2(n14125), .Q(n14121) );
  AND2X1 U14320 ( .IN1(n14112), .IN2(g2619), .Q(n14125) );
  OR2X1 U14321 ( .IN1(n3519), .IN2(n14126), .Q(g33016) );
  OR2X1 U14322 ( .IN1(n14127), .IN2(n14128), .Q(n14126) );
  AND2X1 U14323 ( .IN1(n14129), .IN2(g2587), .Q(n14128) );
  AND2X1 U14324 ( .IN1(n14112), .IN2(g2610), .Q(n14127) );
  OR2X1 U14325 ( .IN1(n14130), .IN2(n14131), .Q(g33015) );
  OR2X1 U14326 ( .IN1(n14132), .IN2(n14133), .Q(n14131) );
  AND2X1 U14327 ( .IN1(test_so34), .IN2(n10895), .Q(n14133) );
  AND2X1 U14328 ( .IN1(n14112), .IN2(g2587), .Q(n14132) );
  OR2X1 U14329 ( .IN1(n3519), .IN2(n14134), .Q(n14130) );
  AND2X1 U14330 ( .IN1(n14135), .IN2(n3517), .Q(n14134) );
  AND2X1 U14331 ( .IN1(n5508), .IN2(n14136), .Q(n14135) );
  OR2X1 U14332 ( .IN1(n14137), .IN2(n14138), .Q(g33014) );
  OR2X1 U14333 ( .IN1(n14139), .IN2(n14140), .Q(n14138) );
  AND2X1 U14334 ( .IN1(n14141), .IN2(g2491), .Q(n14140) );
  OR2X1 U14335 ( .IN1(n14142), .IN2(n14143), .Q(n14141) );
  OR2X1 U14336 ( .IN1(n13293), .IN2(n14144), .Q(n14143) );
  AND2X1 U14337 ( .IN1(n3007), .IN2(n10750), .Q(n14142) );
  AND2X1 U14338 ( .IN1(n14145), .IN2(n3536), .Q(n14139) );
  AND2X1 U14339 ( .IN1(n3531), .IN2(n11219), .Q(n14145) );
  AND2X1 U14340 ( .IN1(n12360), .IN2(n3524), .Q(n11219) );
  INVX0 U14341 ( .INP(n3007), .ZN(n12360) );
  OR2X1 U14342 ( .IN1(n14146), .IN2(n14147), .Q(n3007) );
  OR2X1 U14343 ( .IN1(n5516), .IN2(g2741), .Q(n14147) );
  OR2X1 U14344 ( .IN1(g2476), .IN2(n14148), .Q(n3531) );
  OR2X1 U14345 ( .IN1(n5509), .IN2(n10531), .Q(n14148) );
  OR2X1 U14346 ( .IN1(n14149), .IN2(n14150), .Q(n14137) );
  AND2X1 U14347 ( .IN1(n14151), .IN2(n10470), .Q(n14150) );
  AND2X1 U14348 ( .IN1(n14152), .IN2(n14153), .Q(n14151) );
  AND2X1 U14349 ( .IN1(n14154), .IN2(g2485), .Q(n14153) );
  AND2X1 U14350 ( .IN1(n3530), .IN2(n12005), .Q(n14152) );
  AND2X1 U14351 ( .IN1(n10928), .IN2(g2476), .Q(n14149) );
  OR2X1 U14352 ( .IN1(n14155), .IN2(n14156), .Q(g33013) );
  OR2X1 U14353 ( .IN1(n14157), .IN2(n14158), .Q(n14156) );
  AND2X1 U14354 ( .IN1(n10928), .IN2(g2491), .Q(n14158) );
  AND2X1 U14355 ( .IN1(n3536), .IN2(g2476), .Q(n14157) );
  OR2X1 U14356 ( .IN1(n3538), .IN2(n14159), .Q(n14155) );
  AND2X1 U14357 ( .IN1(n14144), .IN2(g2485), .Q(n14159) );
  OR2X1 U14358 ( .IN1(n3538), .IN2(n14160), .Q(g33012) );
  OR2X1 U14359 ( .IN1(n14161), .IN2(n14162), .Q(n14160) );
  AND2X1 U14360 ( .IN1(n14163), .IN2(g2453), .Q(n14162) );
  AND2X1 U14361 ( .IN1(n14144), .IN2(g2476), .Q(n14161) );
  OR2X1 U14362 ( .IN1(n14164), .IN2(n14165), .Q(g33011) );
  OR2X1 U14363 ( .IN1(n14166), .IN2(n14167), .Q(n14165) );
  AND2X1 U14364 ( .IN1(n10928), .IN2(g2461), .Q(n14167) );
  AND2X1 U14365 ( .IN1(n14144), .IN2(g2453), .Q(n14166) );
  OR2X1 U14366 ( .IN1(n3538), .IN2(n14168), .Q(n14164) );
  AND2X1 U14367 ( .IN1(n14169), .IN2(n3536), .Q(n14168) );
  AND2X1 U14368 ( .IN1(n5509), .IN2(n14170), .Q(n14169) );
  OR2X1 U14369 ( .IN1(n14171), .IN2(n14172), .Q(g33010) );
  OR2X1 U14370 ( .IN1(n14173), .IN2(n14174), .Q(n14172) );
  AND2X1 U14371 ( .IN1(n14175), .IN2(g2357), .Q(n14174) );
  OR2X1 U14372 ( .IN1(n14176), .IN2(n14177), .Q(n14175) );
  OR2X1 U14373 ( .IN1(n13293), .IN2(n14178), .Q(n14177) );
  AND2X1 U14374 ( .IN1(n3550), .IN2(n10750), .Q(n14176) );
  AND2X1 U14375 ( .IN1(n14179), .IN2(n3555), .Q(n14173) );
  AND2X1 U14376 ( .IN1(n3549), .IN2(n11216), .Q(n14179) );
  AND2X1 U14377 ( .IN1(n12356), .IN2(n3524), .Q(n11216) );
  INVX0 U14378 ( .INP(n3550), .ZN(n12356) );
  OR2X1 U14379 ( .IN1(n14146), .IN2(n14180), .Q(n3550) );
  OR2X1 U14380 ( .IN1(n5349), .IN2(g2748), .Q(n14180) );
  OR2X1 U14381 ( .IN1(n10531), .IN2(n14181), .Q(n3549) );
  OR2X1 U14382 ( .IN1(test_so21), .IN2(n5511), .Q(n14181) );
  OR2X1 U14383 ( .IN1(n14182), .IN2(n14183), .Q(n14171) );
  AND2X1 U14384 ( .IN1(n14184), .IN2(n10555), .Q(n14183) );
  AND2X1 U14385 ( .IN1(n14185), .IN2(n14186), .Q(n14184) );
  AND2X1 U14386 ( .IN1(n14187), .IN2(g2351), .Q(n14186) );
  AND2X1 U14387 ( .IN1(n3548), .IN2(n12005), .Q(n14185) );
  AND2X1 U14388 ( .IN1(test_so21), .IN2(n10894), .Q(n14182) );
  OR2X1 U14389 ( .IN1(n14188), .IN2(n14189), .Q(g33009) );
  OR2X1 U14390 ( .IN1(n14190), .IN2(n14191), .Q(n14189) );
  AND2X1 U14391 ( .IN1(n10928), .IN2(g2357), .Q(n14191) );
  AND2X1 U14392 ( .IN1(n3555), .IN2(test_so21), .Q(n14190) );
  OR2X1 U14393 ( .IN1(n3557), .IN2(n14192), .Q(n14188) );
  AND2X1 U14394 ( .IN1(n14178), .IN2(g2351), .Q(n14192) );
  OR2X1 U14395 ( .IN1(n3557), .IN2(n14193), .Q(g33008) );
  OR2X1 U14396 ( .IN1(n14194), .IN2(n14195), .Q(n14193) );
  AND2X1 U14397 ( .IN1(n14196), .IN2(g2319), .Q(n14195) );
  AND2X1 U14398 ( .IN1(n14178), .IN2(test_so21), .Q(n14194) );
  OR2X1 U14399 ( .IN1(n14197), .IN2(n14198), .Q(g33007) );
  OR2X1 U14400 ( .IN1(n14199), .IN2(n14200), .Q(n14198) );
  AND2X1 U14401 ( .IN1(n10928), .IN2(g2327), .Q(n14200) );
  AND2X1 U14402 ( .IN1(n14178), .IN2(g2319), .Q(n14199) );
  OR2X1 U14403 ( .IN1(n3557), .IN2(n14201), .Q(n14197) );
  AND2X1 U14404 ( .IN1(n14202), .IN2(n3555), .Q(n14201) );
  AND2X1 U14405 ( .IN1(n5511), .IN2(n14203), .Q(n14202) );
  OR2X1 U14406 ( .IN1(n14204), .IN2(n14205), .Q(g33006) );
  OR2X1 U14407 ( .IN1(n14206), .IN2(n14207), .Q(n14205) );
  AND2X1 U14408 ( .IN1(n14208), .IN2(g2223), .Q(n14207) );
  OR2X1 U14409 ( .IN1(n14209), .IN2(n14210), .Q(n14208) );
  OR2X1 U14410 ( .IN1(n13293), .IN2(n14211), .Q(n14210) );
  AND2X1 U14411 ( .IN1(n3569), .IN2(n10750), .Q(n14209) );
  AND2X1 U14412 ( .IN1(n14212), .IN2(n3574), .Q(n14206) );
  AND2X1 U14413 ( .IN1(n3568), .IN2(n11217), .Q(n14212) );
  AND2X1 U14414 ( .IN1(n12354), .IN2(n3524), .Q(n11217) );
  INVX0 U14415 ( .INP(n3569), .ZN(n12354) );
  OR2X1 U14416 ( .IN1(n14146), .IN2(n14213), .Q(n3569) );
  OR2X1 U14417 ( .IN1(g2748), .IN2(g2741), .Q(n14213) );
  INVX0 U14418 ( .INP(n3525), .ZN(n14146) );
  OR2X1 U14419 ( .IN1(g2208), .IN2(n14214), .Q(n3568) );
  OR2X1 U14420 ( .IN1(n5512), .IN2(n10531), .Q(n14214) );
  OR2X1 U14421 ( .IN1(n14215), .IN2(n14216), .Q(n14204) );
  AND2X1 U14422 ( .IN1(n14217), .IN2(n10471), .Q(n14216) );
  AND2X1 U14423 ( .IN1(n14218), .IN2(n14219), .Q(n14217) );
  AND2X1 U14424 ( .IN1(n14220), .IN2(g2217), .Q(n14219) );
  AND2X1 U14425 ( .IN1(n3567), .IN2(n12005), .Q(n14218) );
  AND2X1 U14426 ( .IN1(n10928), .IN2(g2208), .Q(n14215) );
  OR2X1 U14427 ( .IN1(n14221), .IN2(n14222), .Q(g33005) );
  OR2X1 U14428 ( .IN1(n14223), .IN2(n14224), .Q(n14222) );
  AND2X1 U14429 ( .IN1(n10928), .IN2(g2223), .Q(n14224) );
  AND2X1 U14430 ( .IN1(n3574), .IN2(g2208), .Q(n14223) );
  OR2X1 U14431 ( .IN1(n3576), .IN2(n14225), .Q(n14221) );
  AND2X1 U14432 ( .IN1(n14211), .IN2(g2217), .Q(n14225) );
  OR2X1 U14433 ( .IN1(n3576), .IN2(n14226), .Q(g33004) );
  OR2X1 U14434 ( .IN1(n14227), .IN2(n14228), .Q(n14226) );
  AND2X1 U14435 ( .IN1(n14229), .IN2(g2185), .Q(n14228) );
  AND2X1 U14436 ( .IN1(n14211), .IN2(g2208), .Q(n14227) );
  OR2X1 U14437 ( .IN1(n14230), .IN2(n14231), .Q(g33003) );
  OR2X1 U14438 ( .IN1(n14232), .IN2(n14233), .Q(n14231) );
  AND2X1 U14439 ( .IN1(n10929), .IN2(g2193), .Q(n14233) );
  AND2X1 U14440 ( .IN1(n14211), .IN2(g2185), .Q(n14232) );
  OR2X1 U14441 ( .IN1(n3576), .IN2(n14234), .Q(n14230) );
  AND2X1 U14442 ( .IN1(n14235), .IN2(n3574), .Q(n14234) );
  AND2X1 U14443 ( .IN1(n5512), .IN2(n14236), .Q(n14235) );
  OR2X1 U14444 ( .IN1(n14237), .IN2(n14238), .Q(g33002) );
  OR2X1 U14445 ( .IN1(n14239), .IN2(n14240), .Q(n14238) );
  AND2X1 U14446 ( .IN1(n14241), .IN2(g2066), .Q(n14240) );
  OR2X1 U14447 ( .IN1(n14242), .IN2(n14243), .Q(n14241) );
  OR2X1 U14448 ( .IN1(n13293), .IN2(n14244), .Q(n14243) );
  AND2X1 U14449 ( .IN1(n3588), .IN2(n10750), .Q(n14242) );
  AND2X1 U14450 ( .IN1(n14245), .IN2(n3593), .Q(n14239) );
  AND2X1 U14451 ( .IN1(n3587), .IN2(n11077), .Q(n14245) );
  AND2X1 U14452 ( .IN1(n12348), .IN2(n3524), .Q(n11077) );
  INVX0 U14453 ( .INP(n3588), .ZN(n12348) );
  OR2X1 U14454 ( .IN1(n14246), .IN2(n14247), .Q(n3588) );
  OR2X1 U14455 ( .IN1(test_so30), .IN2(n11074), .Q(n14247) );
  INVX0 U14456 ( .INP(n1284), .ZN(n14246) );
  OR2X1 U14457 ( .IN1(g2051), .IN2(n14248), .Q(n3587) );
  OR2X1 U14458 ( .IN1(n5507), .IN2(n10531), .Q(n14248) );
  OR2X1 U14459 ( .IN1(n14249), .IN2(n14250), .Q(n14237) );
  AND2X1 U14460 ( .IN1(n14251), .IN2(n10472), .Q(n14250) );
  AND2X1 U14461 ( .IN1(n14252), .IN2(n14253), .Q(n14251) );
  AND2X1 U14462 ( .IN1(n14254), .IN2(g2060), .Q(n14253) );
  AND2X1 U14463 ( .IN1(n3586), .IN2(n12005), .Q(n14252) );
  AND2X1 U14464 ( .IN1(n10929), .IN2(g2051), .Q(n14249) );
  OR2X1 U14465 ( .IN1(n14255), .IN2(n14256), .Q(g33001) );
  OR2X1 U14466 ( .IN1(n14257), .IN2(n14258), .Q(n14256) );
  AND2X1 U14467 ( .IN1(n10929), .IN2(g2066), .Q(n14258) );
  AND2X1 U14468 ( .IN1(n3593), .IN2(g2051), .Q(n14257) );
  OR2X1 U14469 ( .IN1(n3595), .IN2(n14259), .Q(n14255) );
  AND2X1 U14470 ( .IN1(n14244), .IN2(g2060), .Q(n14259) );
  OR2X1 U14471 ( .IN1(n3595), .IN2(n14260), .Q(g33000) );
  OR2X1 U14472 ( .IN1(n14261), .IN2(n14262), .Q(n14260) );
  AND2X1 U14473 ( .IN1(n14263), .IN2(g2028), .Q(n14262) );
  AND2X1 U14474 ( .IN1(n14244), .IN2(g2051), .Q(n14261) );
  OR2X1 U14475 ( .IN1(n14264), .IN2(n14265), .Q(g32999) );
  OR2X1 U14476 ( .IN1(n14266), .IN2(n14267), .Q(n14265) );
  AND2X1 U14477 ( .IN1(test_so59), .IN2(n10894), .Q(n14267) );
  AND2X1 U14478 ( .IN1(n14244), .IN2(g2028), .Q(n14266) );
  OR2X1 U14479 ( .IN1(n3595), .IN2(n14268), .Q(n14264) );
  AND2X1 U14480 ( .IN1(n14269), .IN2(n3593), .Q(n14268) );
  AND2X1 U14481 ( .IN1(n5507), .IN2(n14270), .Q(n14269) );
  OR2X1 U14482 ( .IN1(n14271), .IN2(n14272), .Q(g32998) );
  OR2X1 U14483 ( .IN1(n14273), .IN2(n14274), .Q(n14272) );
  AND2X1 U14484 ( .IN1(n14275), .IN2(g1932), .Q(n14274) );
  OR2X1 U14485 ( .IN1(n14276), .IN2(n14277), .Q(n14275) );
  OR2X1 U14486 ( .IN1(n13293), .IN2(n14278), .Q(n14277) );
  AND2X1 U14487 ( .IN1(n3606), .IN2(n10749), .Q(n14276) );
  AND2X1 U14488 ( .IN1(n14279), .IN2(n3611), .Q(n14273) );
  AND2X1 U14489 ( .IN1(n3605), .IN2(n11076), .Q(n14279) );
  AND2X1 U14490 ( .IN1(n12346), .IN2(n3524), .Q(n11076) );
  INVX0 U14491 ( .INP(n3606), .ZN(n12346) );
  OR2X1 U14492 ( .IN1(n14280), .IN2(n14281), .Q(n3606) );
  OR2X1 U14493 ( .IN1(g2741), .IN2(n11074), .Q(n14281) );
  OR2X1 U14494 ( .IN1(test_so30), .IN2(n5516), .Q(n14280) );
  OR2X1 U14495 ( .IN1(g1917), .IN2(n14282), .Q(n3605) );
  OR2X1 U14496 ( .IN1(n5510), .IN2(n10531), .Q(n14282) );
  OR2X1 U14497 ( .IN1(n14283), .IN2(n14284), .Q(n14271) );
  AND2X1 U14498 ( .IN1(n14285), .IN2(n10469), .Q(n14284) );
  AND2X1 U14499 ( .IN1(n14286), .IN2(n14287), .Q(n14285) );
  AND2X1 U14500 ( .IN1(n14288), .IN2(g1926), .Q(n14287) );
  AND2X1 U14501 ( .IN1(n3604), .IN2(n12005), .Q(n14286) );
  AND2X1 U14502 ( .IN1(n10929), .IN2(g1917), .Q(n14283) );
  OR2X1 U14503 ( .IN1(n14289), .IN2(n14290), .Q(g32997) );
  OR2X1 U14504 ( .IN1(n14291), .IN2(n14292), .Q(n14290) );
  AND2X1 U14505 ( .IN1(n10929), .IN2(g1932), .Q(n14292) );
  AND2X1 U14506 ( .IN1(n3611), .IN2(g1917), .Q(n14291) );
  OR2X1 U14507 ( .IN1(n3613), .IN2(n14293), .Q(n14289) );
  AND2X1 U14508 ( .IN1(n14278), .IN2(g1926), .Q(n14293) );
  OR2X1 U14509 ( .IN1(n3613), .IN2(n14294), .Q(g32996) );
  OR2X1 U14510 ( .IN1(n14295), .IN2(n14296), .Q(n14294) );
  AND2X1 U14511 ( .IN1(n14297), .IN2(g1894), .Q(n14296) );
  AND2X1 U14512 ( .IN1(n14278), .IN2(g1917), .Q(n14295) );
  OR2X1 U14513 ( .IN1(n14298), .IN2(n14299), .Q(g32995) );
  OR2X1 U14514 ( .IN1(n14300), .IN2(n14301), .Q(n14299) );
  AND2X1 U14515 ( .IN1(n10929), .IN2(g1902), .Q(n14301) );
  AND2X1 U14516 ( .IN1(n14278), .IN2(g1894), .Q(n14300) );
  OR2X1 U14517 ( .IN1(n3613), .IN2(n14302), .Q(n14298) );
  AND2X1 U14518 ( .IN1(n14303), .IN2(n3611), .Q(n14302) );
  AND2X1 U14519 ( .IN1(n5510), .IN2(n14304), .Q(n14303) );
  OR2X1 U14520 ( .IN1(n14305), .IN2(n14306), .Q(g32994) );
  OR2X1 U14521 ( .IN1(n14307), .IN2(n14308), .Q(n14306) );
  AND2X1 U14522 ( .IN1(n14309), .IN2(g1798), .Q(n14308) );
  OR2X1 U14523 ( .IN1(n14310), .IN2(n14311), .Q(n14309) );
  OR2X1 U14524 ( .IN1(n13293), .IN2(n14312), .Q(n14311) );
  AND2X1 U14525 ( .IN1(n10820), .IN2(n1645), .Q(n14310) );
  INVX0 U14526 ( .INP(n3005), .ZN(n1645) );
  AND2X1 U14527 ( .IN1(n14313), .IN2(n3628), .Q(n14307) );
  AND2X1 U14528 ( .IN1(n3623), .IN2(n11215), .Q(n14313) );
  AND2X1 U14529 ( .IN1(n3005), .IN2(n3524), .Q(n11215) );
  OR2X1 U14530 ( .IN1(g1783), .IN2(n14314), .Q(n3623) );
  OR2X1 U14531 ( .IN1(n5359), .IN2(n10531), .Q(n14314) );
  OR2X1 U14532 ( .IN1(n14315), .IN2(n14316), .Q(n14305) );
  AND2X1 U14533 ( .IN1(n14317), .IN2(n5596), .Q(n14316) );
  AND2X1 U14534 ( .IN1(n14318), .IN2(n14319), .Q(n14317) );
  AND2X1 U14535 ( .IN1(n14320), .IN2(g1792), .Q(n14319) );
  AND2X1 U14536 ( .IN1(n3622), .IN2(n12005), .Q(n14318) );
  AND2X1 U14537 ( .IN1(n10929), .IN2(g1783), .Q(n14315) );
  OR2X1 U14538 ( .IN1(n14321), .IN2(n14322), .Q(g32993) );
  OR2X1 U14539 ( .IN1(n14323), .IN2(n14324), .Q(n14322) );
  AND2X1 U14540 ( .IN1(n10929), .IN2(g1798), .Q(n14324) );
  AND2X1 U14541 ( .IN1(n3628), .IN2(g1783), .Q(n14323) );
  OR2X1 U14542 ( .IN1(n3630), .IN2(n14325), .Q(n14321) );
  AND2X1 U14543 ( .IN1(n14312), .IN2(g1792), .Q(n14325) );
  OR2X1 U14544 ( .IN1(n3630), .IN2(n14326), .Q(g32992) );
  OR2X1 U14545 ( .IN1(n14327), .IN2(n14328), .Q(n14326) );
  AND2X1 U14546 ( .IN1(n14329), .IN2(g1760), .Q(n14328) );
  AND2X1 U14547 ( .IN1(n14312), .IN2(g1783), .Q(n14327) );
  OR2X1 U14548 ( .IN1(n14330), .IN2(n14331), .Q(g32991) );
  OR2X1 U14549 ( .IN1(n14332), .IN2(n14333), .Q(n14331) );
  AND2X1 U14550 ( .IN1(n10929), .IN2(g1768), .Q(n14333) );
  AND2X1 U14551 ( .IN1(n14312), .IN2(g1760), .Q(n14332) );
  OR2X1 U14552 ( .IN1(n3630), .IN2(n14334), .Q(n14330) );
  AND2X1 U14553 ( .IN1(n14335), .IN2(n3628), .Q(n14334) );
  AND2X1 U14554 ( .IN1(n5359), .IN2(n14336), .Q(n14335) );
  OR2X1 U14555 ( .IN1(n14337), .IN2(n14338), .Q(g32990) );
  OR2X1 U14556 ( .IN1(n14339), .IN2(n14340), .Q(n14338) );
  AND2X1 U14557 ( .IN1(n14341), .IN2(g1664), .Q(n14340) );
  OR2X1 U14558 ( .IN1(n14342), .IN2(n14343), .Q(n14341) );
  OR2X1 U14559 ( .IN1(n13293), .IN2(n14344), .Q(n14343) );
  AND2X1 U14560 ( .IN1(n1698), .IN2(n10749), .Q(n13293) );
  INVX0 U14561 ( .INP(n2760), .ZN(n1698) );
  AND2X1 U14562 ( .IN1(n3003), .IN2(n10749), .Q(n14342) );
  AND2X1 U14563 ( .IN1(n14345), .IN2(n3646), .Q(n14339) );
  AND2X1 U14564 ( .IN1(n3641), .IN2(n11075), .Q(n14345) );
  AND2X1 U14565 ( .IN1(n12341), .IN2(n3524), .Q(n11075) );
  INVX0 U14566 ( .INP(n3003), .ZN(n12341) );
  OR2X1 U14567 ( .IN1(n11074), .IN2(n14346), .Q(n3003) );
  OR2X1 U14568 ( .IN1(n14347), .IN2(n14348), .Q(n11074) );
  XNOR2X1 U14569 ( .IN1(n10530), .IN2(g72), .Q(n14348) );
  XNOR2X1 U14570 ( .IN1(n10019), .IN2(g73), .Q(n14347) );
  OR2X1 U14571 ( .IN1(n10531), .IN2(n14349), .Q(n3641) );
  OR2X1 U14572 ( .IN1(test_so94), .IN2(n5525), .Q(n14349) );
  OR2X1 U14573 ( .IN1(n14350), .IN2(n14351), .Q(n14337) );
  AND2X1 U14574 ( .IN1(n14352), .IN2(n10556), .Q(n14351) );
  AND2X1 U14575 ( .IN1(n14353), .IN2(n14354), .Q(n14352) );
  AND2X1 U14576 ( .IN1(n14355), .IN2(g1657), .Q(n14354) );
  AND2X1 U14577 ( .IN1(n3640), .IN2(n12005), .Q(n14353) );
  AND2X1 U14578 ( .IN1(test_so94), .IN2(n10895), .Q(n14350) );
  OR2X1 U14579 ( .IN1(n14356), .IN2(n14357), .Q(g32989) );
  OR2X1 U14580 ( .IN1(n14358), .IN2(n14359), .Q(n14357) );
  AND2X1 U14581 ( .IN1(n10929), .IN2(g1664), .Q(n14359) );
  AND2X1 U14582 ( .IN1(n3646), .IN2(test_so94), .Q(n14358) );
  OR2X1 U14583 ( .IN1(n3648), .IN2(n14360), .Q(n14356) );
  AND2X1 U14584 ( .IN1(n14344), .IN2(g1657), .Q(n14360) );
  OR2X1 U14585 ( .IN1(n3648), .IN2(n14361), .Q(g32988) );
  OR2X1 U14586 ( .IN1(n14362), .IN2(n14363), .Q(n14361) );
  INVX0 U14587 ( .INP(n14364), .ZN(n14363) );
  OR2X1 U14588 ( .IN1(n14344), .IN2(n5370), .Q(n14364) );
  AND2X1 U14589 ( .IN1(n14344), .IN2(test_so94), .Q(n14362) );
  OR2X1 U14590 ( .IN1(n14365), .IN2(n14366), .Q(g32987) );
  OR2X1 U14591 ( .IN1(n14367), .IN2(n14368), .Q(n14366) );
  AND2X1 U14592 ( .IN1(n10929), .IN2(g1632), .Q(n14368) );
  AND2X1 U14593 ( .IN1(n14344), .IN2(g1624), .Q(n14367) );
  OR2X1 U14594 ( .IN1(n3648), .IN2(n14369), .Q(n14365) );
  AND2X1 U14595 ( .IN1(n14370), .IN2(n3646), .Q(n14369) );
  AND2X1 U14596 ( .IN1(n5525), .IN2(n14371), .Q(n14370) );
  OR2X1 U14597 ( .IN1(n14372), .IN2(n14373), .Q(g32986) );
  OR2X1 U14598 ( .IN1(n14374), .IN2(n14375), .Q(n14373) );
  AND2X1 U14599 ( .IN1(n10929), .IN2(g1367), .Q(n14375) );
  AND2X1 U14600 ( .IN1(n14376), .IN2(n10749), .Q(n14374) );
  AND2X1 U14601 ( .IN1(n13791), .IN2(g1373), .Q(n14376) );
  AND2X1 U14602 ( .IN1(n14377), .IN2(n14378), .Q(n14372) );
  AND2X1 U14603 ( .IN1(n13786), .IN2(n10462), .Q(n14377) );
  INVX0 U14604 ( .INP(n13791), .ZN(n13786) );
  OR2X1 U14605 ( .IN1(n14379), .IN2(n11214), .Q(n13791) );
  AND2X1 U14606 ( .IN1(n10121), .IN2(n13787), .Q(n14379) );
  AND2X1 U14607 ( .IN1(n14380), .IN2(g1274), .Q(g32985) );
  OR2X1 U14608 ( .IN1(n10892), .IN2(n14381), .Q(n14380) );
  AND2X1 U14609 ( .IN1(n13796), .IN2(n11668), .Q(n14381) );
  AND2X1 U14610 ( .IN1(g1270), .IN2(n3662), .Q(n13796) );
  OR2X1 U14611 ( .IN1(n14382), .IN2(n14383), .Q(g32984) );
  OR2X1 U14612 ( .IN1(n14384), .IN2(n14385), .Q(n14383) );
  AND2X1 U14613 ( .IN1(n5716), .IN2(n3662), .Q(n14385) );
  INVX0 U14614 ( .INP(n14386), .ZN(n14384) );
  OR2X1 U14615 ( .IN1(n14387), .IN2(n5716), .Q(n14386) );
  OR2X1 U14616 ( .IN1(n13799), .IN2(n3662), .Q(n14387) );
  AND2X1 U14617 ( .IN1(n10929), .IN2(g1263), .Q(n14382) );
  OR2X1 U14618 ( .IN1(n14388), .IN2(n14389), .Q(g32983) );
  OR2X1 U14619 ( .IN1(n14390), .IN2(n14391), .Q(n14389) );
  AND2X1 U14620 ( .IN1(n10929), .IN2(g1024), .Q(n14391) );
  AND2X1 U14621 ( .IN1(n14392), .IN2(n10749), .Q(n14390) );
  AND2X1 U14622 ( .IN1(n13810), .IN2(g1030), .Q(n14392) );
  AND2X1 U14623 ( .IN1(n14393), .IN2(n14394), .Q(n14388) );
  AND2X1 U14624 ( .IN1(n13805), .IN2(n10461), .Q(n14393) );
  INVX0 U14625 ( .INP(n13810), .ZN(n13805) );
  OR2X1 U14626 ( .IN1(n14395), .IN2(n11098), .Q(n13810) );
  AND2X1 U14627 ( .IN1(n10122), .IN2(n13806), .Q(n14395) );
  AND2X1 U14628 ( .IN1(n14396), .IN2(g930), .Q(g32982) );
  OR2X1 U14629 ( .IN1(n10892), .IN2(n14397), .Q(n14396) );
  AND2X1 U14630 ( .IN1(n13815), .IN2(n11669), .Q(n14397) );
  AND2X1 U14631 ( .IN1(g925), .IN2(n3671), .Q(n13815) );
  OR2X1 U14632 ( .IN1(n14398), .IN2(n14399), .Q(g32981) );
  OR2X1 U14633 ( .IN1(n14400), .IN2(n14401), .Q(n14399) );
  AND2X1 U14634 ( .IN1(n5725), .IN2(n3671), .Q(n14401) );
  INVX0 U14635 ( .INP(n14402), .ZN(n14400) );
  OR2X1 U14636 ( .IN1(n14403), .IN2(n5725), .Q(n14402) );
  OR2X1 U14637 ( .IN1(n13818), .IN2(n3671), .Q(n14403) );
  AND2X1 U14638 ( .IN1(n10929), .IN2(g918), .Q(n14398) );
  AND2X1 U14639 ( .IN1(n14404), .IN2(n10749), .Q(g32980) );
  AND2X1 U14640 ( .IN1(n14405), .IN2(n14406), .Q(n14404) );
  OR2X1 U14641 ( .IN1(n14407), .IN2(g854), .Q(n14406) );
  INVX0 U14642 ( .INP(n12085), .ZN(n14407) );
  OR2X1 U14643 ( .IN1(n12085), .IN2(n14408), .Q(n14405) );
  INVX0 U14644 ( .INP(n2644), .ZN(n14408) );
  OR2X1 U14645 ( .IN1(n14409), .IN2(n14410), .Q(n12085) );
  OR2X1 U14646 ( .IN1(n10155), .IN2(g385), .Q(n14410) );
  OR2X1 U14647 ( .IN1(n5633), .IN2(n10156), .Q(n14409) );
  OR2X1 U14648 ( .IN1(n14411), .IN2(n14412), .Q(g32979) );
  OR2X1 U14649 ( .IN1(n14413), .IN2(n14414), .Q(n14412) );
  AND2X1 U14650 ( .IN1(n3272), .IN2(n5331), .Q(n14414) );
  AND2X1 U14651 ( .IN1(n14415), .IN2(g758), .Q(n14413) );
  AND2X1 U14652 ( .IN1(n2404), .IN2(n14416), .Q(n14415) );
  INVX0 U14653 ( .INP(n3272), .ZN(n14416) );
  AND2X1 U14654 ( .IN1(test_so2), .IN2(n10894), .Q(n14411) );
  OR2X1 U14655 ( .IN1(n14417), .IN2(n14418), .Q(g32978) );
  OR2X1 U14656 ( .IN1(n14419), .IN2(n14420), .Q(n14418) );
  AND2X1 U14657 ( .IN1(n3274), .IN2(n5472), .Q(n14420) );
  AND2X1 U14658 ( .IN1(n14421), .IN2(g590), .Q(n14419) );
  AND2X1 U14659 ( .IN1(n2421), .IN2(n14422), .Q(n14421) );
  INVX0 U14660 ( .INP(n3274), .ZN(n14422) );
  AND2X1 U14661 ( .IN1(n10929), .IN2(g582), .Q(n14417) );
  OR2X1 U14662 ( .IN1(n14423), .IN2(n14424), .Q(g32977) );
  OR2X1 U14663 ( .IN1(n14425), .IN2(n14426), .Q(n14424) );
  AND2X1 U14664 ( .IN1(n44), .IN2(n5679), .Q(n14426) );
  INVX0 U14665 ( .INP(n14427), .ZN(n44) );
  AND2X1 U14666 ( .IN1(n14428), .IN2(g291), .Q(n14425) );
  AND2X1 U14667 ( .IN1(n10534), .IN2(n14427), .Q(n14428) );
  OR2X1 U14668 ( .IN1(n10558), .IN2(n14429), .Q(n14427) );
  OR2X1 U14669 ( .IN1(n14430), .IN2(n10571), .Q(n14429) );
  AND2X1 U14670 ( .IN1(test_so51), .IN2(n10894), .Q(n14423) );
  OR2X1 U14671 ( .IN1(n14431), .IN2(n14432), .Q(g32976) );
  OR2X1 U14672 ( .IN1(n14433), .IN2(n14434), .Q(n14432) );
  AND2X1 U14673 ( .IN1(n3281), .IN2(n5676), .Q(n14434) );
  AND2X1 U14674 ( .IN1(n14435), .IN2(g150), .Q(n14433) );
  AND2X1 U14675 ( .IN1(n13055), .IN2(n14436), .Q(n14435) );
  INVX0 U14676 ( .INP(n3281), .ZN(n14436) );
  AND2X1 U14677 ( .IN1(n10929), .IN2(g164), .Q(n14431) );
  AND2X1 U14678 ( .IN1(n14437), .IN2(n14438), .Q(g32185) );
  AND2X1 U14679 ( .IN1(n14439), .IN2(n14440), .Q(n14438) );
  AND2X1 U14680 ( .IN1(n14441), .IN2(n14442), .Q(n14440) );
  INVX0 U14681 ( .INP(n14443), .ZN(n14442) );
  AND2X1 U14682 ( .IN1(g2965), .IN2(test_so22), .Q(n14443) );
  OR2X1 U14683 ( .IN1(n10123), .IN2(n10399), .Q(n14441) );
  AND2X1 U14684 ( .IN1(n14444), .IN2(n14445), .Q(n14439) );
  INVX0 U14685 ( .INP(n14446), .ZN(n14445) );
  AND2X1 U14686 ( .IN1(g2902), .IN2(test_so1), .Q(n14446) );
  OR2X1 U14687 ( .IN1(n10124), .IN2(n10398), .Q(n14444) );
  AND2X1 U14688 ( .IN1(n14447), .IN2(n14448), .Q(n14437) );
  OR2X1 U14689 ( .IN1(n10401), .IN2(n10402), .Q(n14448) );
  AND2X1 U14690 ( .IN1(n14449), .IN2(n14450), .Q(n14447) );
  OR2X1 U14691 ( .IN1(n10397), .IN2(n5750), .Q(n14450) );
  OR2X1 U14692 ( .IN1(n10127), .IN2(n10400), .Q(n14449) );
  OR2X1 U14693 ( .IN1(n14451), .IN2(n14452), .Q(g31904) );
  OR2X1 U14694 ( .IN1(n14453), .IN2(n14454), .Q(n14452) );
  AND2X1 U14695 ( .IN1(n10929), .IN2(g5029), .Q(n14454) );
  OR2X1 U14696 ( .IN1(n14455), .IN2(n14456), .Q(n14451) );
  INVX0 U14697 ( .INP(n14457), .ZN(n14456) );
  OR2X1 U14698 ( .IN1(g5033), .IN2(n14458), .Q(n14457) );
  AND2X1 U14699 ( .IN1(n14459), .IN2(g5033), .Q(n14455) );
  AND2X1 U14700 ( .IN1(n14460), .IN2(n13988), .Q(n14459) );
  AND2X1 U14701 ( .IN1(n14461), .IN2(n14458), .Q(n14460) );
  OR2X1 U14702 ( .IN1(n14462), .IN2(n14463), .Q(g31903) );
  OR2X1 U14703 ( .IN1(n13992), .IN2(n14464), .Q(n14463) );
  AND2X1 U14704 ( .IN1(n10930), .IN2(g5046), .Q(n14464) );
  AND2X1 U14705 ( .IN1(n14465), .IN2(n14466), .Q(n13992) );
  AND2X1 U14706 ( .IN1(n10820), .IN2(n5607), .Q(n14466) );
  OR2X1 U14707 ( .IN1(n14467), .IN2(n14468), .Q(n14462) );
  AND2X1 U14708 ( .IN1(n13993), .IN2(n5607), .Q(n14468) );
  AND2X1 U14709 ( .IN1(n14469), .IN2(g5052), .Q(n14467) );
  AND2X1 U14710 ( .IN1(n14470), .IN2(n13988), .Q(n14469) );
  INVX0 U14711 ( .INP(n14471), .ZN(n14470) );
  OR2X1 U14712 ( .IN1(n14465), .IN2(n13993), .Q(n14471) );
  AND2X1 U14713 ( .IN1(g5046), .IN2(n14472), .Q(n13993) );
  OR2X1 U14714 ( .IN1(n14473), .IN2(n14474), .Q(g31902) );
  OR2X1 U14715 ( .IN1(n14475), .IN2(n14476), .Q(n14474) );
  AND2X1 U14716 ( .IN1(n14477), .IN2(g5016), .Q(n14476) );
  OR2X1 U14717 ( .IN1(n10891), .IN2(n14478), .Q(n14477) );
  AND2X1 U14718 ( .IN1(n5601), .IN2(g5062), .Q(n14478) );
  AND2X1 U14719 ( .IN1(n14479), .IN2(n14480), .Q(n14475) );
  AND2X1 U14720 ( .IN1(n14481), .IN2(n14482), .Q(n14480) );
  OR2X1 U14721 ( .IN1(n5369), .IN2(n10508), .Q(n14482) );
  AND2X1 U14722 ( .IN1(n13988), .IN2(g5029), .Q(n14479) );
  AND2X1 U14723 ( .IN1(n14483), .IN2(n10749), .Q(n14473) );
  INVX0 U14724 ( .INP(n14461), .ZN(n14483) );
  OR2X1 U14725 ( .IN1(n14484), .IN2(n14485), .Q(g31901) );
  OR2X1 U14726 ( .IN1(n14486), .IN2(n14487), .Q(n14485) );
  AND2X1 U14727 ( .IN1(n14465), .IN2(n10749), .Q(n14487) );
  AND2X1 U14728 ( .IN1(n5578), .IN2(n14488), .Q(n14465) );
  AND2X1 U14729 ( .IN1(n10930), .IN2(g5041), .Q(n14486) );
  OR2X1 U14730 ( .IN1(n14489), .IN2(n14490), .Q(n14484) );
  AND2X1 U14731 ( .IN1(n14472), .IN2(n5578), .Q(n14490) );
  AND2X1 U14732 ( .IN1(n14491), .IN2(g5046), .Q(n14489) );
  AND2X1 U14733 ( .IN1(n14492), .IN2(n13988), .Q(n14491) );
  AND2X1 U14734 ( .IN1(n14493), .IN2(n14494), .Q(n14492) );
  INVX0 U14735 ( .INP(n14472), .ZN(n14494) );
  AND2X1 U14736 ( .IN1(g5041), .IN2(n14495), .Q(n14472) );
  OR2X1 U14737 ( .IN1(n14496), .IN2(n14497), .Q(g31900) );
  OR2X1 U14738 ( .IN1(n14498), .IN2(n14499), .Q(n14497) );
  AND2X1 U14739 ( .IN1(n14488), .IN2(n10748), .Q(n14499) );
  INVX0 U14740 ( .INP(n14493), .ZN(n14488) );
  OR2X1 U14741 ( .IN1(g5041), .IN2(n14500), .Q(n14493) );
  AND2X1 U14742 ( .IN1(n10930), .IN2(g5037), .Q(n14498) );
  OR2X1 U14743 ( .IN1(n14501), .IN2(n14502), .Q(n14496) );
  AND2X1 U14744 ( .IN1(n14495), .IN2(n5605), .Q(n14502) );
  INVX0 U14745 ( .INP(n14503), .ZN(n14495) );
  AND2X1 U14746 ( .IN1(n14504), .IN2(g5041), .Q(n14501) );
  AND2X1 U14747 ( .IN1(n14505), .IN2(n14506), .Q(n14504) );
  AND2X1 U14748 ( .IN1(n14503), .IN2(n14507), .Q(n14506) );
  OR2X1 U14749 ( .IN1(n5611), .IN2(n14508), .Q(n14503) );
  AND2X1 U14750 ( .IN1(n14509), .IN2(n14500), .Q(n14505) );
  OR2X1 U14751 ( .IN1(n14510), .IN2(g5037), .Q(n14500) );
  OR2X1 U14752 ( .IN1(n14511), .IN2(n14512), .Q(g31899) );
  OR2X1 U14753 ( .IN1(n14513), .IN2(n14514), .Q(n14512) );
  AND2X1 U14754 ( .IN1(n14515), .IN2(g5037), .Q(n14514) );
  AND2X1 U14755 ( .IN1(n14516), .IN2(n13988), .Q(n14515) );
  AND2X1 U14756 ( .IN1(n14510), .IN2(n14508), .Q(n14516) );
  AND2X1 U14757 ( .IN1(n5611), .IN2(n14517), .Q(n14513) );
  OR2X1 U14758 ( .IN1(n14518), .IN2(n14453), .Q(n14517) );
  AND2X1 U14759 ( .IN1(n10821), .IN2(n14519), .Q(n14453) );
  INVX0 U14760 ( .INP(n14510), .ZN(n14519) );
  OR2X1 U14761 ( .IN1(n14461), .IN2(g5033), .Q(n14510) );
  OR2X1 U14762 ( .IN1(g5029), .IN2(n14481), .Q(n14461) );
  OR2X1 U14763 ( .IN1(n10507), .IN2(g5016), .Q(n14481) );
  INVX0 U14764 ( .INP(n14508), .ZN(n14518) );
  OR2X1 U14765 ( .IN1(n10464), .IN2(n14458), .Q(n14508) );
  OR2X1 U14766 ( .IN1(n10508), .IN2(n14520), .Q(n14458) );
  OR2X1 U14767 ( .IN1(n5601), .IN2(n5369), .Q(n14520) );
  AND2X1 U14768 ( .IN1(n10930), .IN2(g5033), .Q(n14511) );
  OR2X1 U14769 ( .IN1(n14521), .IN2(n14522), .Q(g31898) );
  OR2X1 U14770 ( .IN1(n14523), .IN2(n14524), .Q(n14522) );
  AND2X1 U14771 ( .IN1(n10930), .IN2(g5022), .Q(n14524) );
  AND2X1 U14772 ( .IN1(n14525), .IN2(n10748), .Q(n14523) );
  AND2X1 U14773 ( .IN1(n14526), .IN2(g5016), .Q(n14525) );
  INVX0 U14774 ( .INP(n14527), .ZN(n14526) );
  AND2X1 U14775 ( .IN1(n14528), .IN2(n5369), .Q(n14521) );
  AND2X1 U14776 ( .IN1(n13988), .IN2(n14527), .Q(n14528) );
  OR2X1 U14777 ( .IN1(g5022), .IN2(g5062), .Q(n14527) );
  AND2X1 U14778 ( .IN1(n14509), .IN2(n14529), .Q(n13988) );
  OR2X1 U14779 ( .IN1(n14530), .IN2(n14531), .Q(g31897) );
  OR2X1 U14780 ( .IN1(n14005), .IN2(n14532), .Q(n14531) );
  AND2X1 U14781 ( .IN1(n10930), .IN2(g4423), .Q(n14532) );
  AND2X1 U14782 ( .IN1(g4575), .IN2(n14008), .Q(n14005) );
  OR2X1 U14783 ( .IN1(n14530), .IN2(n14533), .Q(g31896) );
  OR2X1 U14784 ( .IN1(n14016), .IN2(n14534), .Q(n14533) );
  INVX0 U14785 ( .INP(n14535), .ZN(n14534) );
  OR2X1 U14786 ( .IN1(n10737), .IN2(n5849), .Q(n14535) );
  AND2X1 U14787 ( .IN1(n14008), .IN2(test_so100), .Q(n14016) );
  OR2X1 U14788 ( .IN1(n14536), .IN2(n14537), .Q(n14530) );
  AND2X1 U14789 ( .IN1(n14008), .IN2(n14538), .Q(n14537) );
  OR2X1 U14790 ( .IN1(n13097), .IN2(n11205), .Q(n14538) );
  INVX0 U14791 ( .INP(g72), .ZN(n11205) );
  INVX0 U14792 ( .INP(g73), .ZN(n13097) );
  AND2X1 U14793 ( .IN1(g4581), .IN2(n10748), .Q(n14008) );
  AND2X1 U14794 ( .IN1(n14539), .IN2(n5670), .Q(n14536) );
  AND2X1 U14795 ( .IN1(n10821), .IN2(g4372), .Q(n14539) );
  OR2X1 U14796 ( .IN1(n14540), .IN2(n12005), .Q(g31895) );
  AND2X1 U14797 ( .IN1(n10821), .IN2(n2760), .Q(n12005) );
  AND2X1 U14798 ( .IN1(n10930), .IN2(g4382), .Q(n14540) );
  OR2X1 U14799 ( .IN1(n10542), .IN2(n14541), .Q(g31894) );
  OR2X1 U14800 ( .IN1(n14542), .IN2(n14543), .Q(n14541) );
  AND2X1 U14801 ( .IN1(n14544), .IN2(n10748), .Q(n14543) );
  XNOR2X1 U14802 ( .IN1(n14031), .IN2(g4098), .Q(n14544) );
  OR2X1 U14803 ( .IN1(n5340), .IN2(n3729), .Q(n14031) );
  OR2X1 U14804 ( .IN1(n5480), .IN2(n14545), .Q(n3729) );
  AND2X1 U14805 ( .IN1(n10930), .IN2(g4093), .Q(n14542) );
  OR2X1 U14806 ( .IN1(n14546), .IN2(n14547), .Q(g31872) );
  AND2X1 U14807 ( .IN1(n10930), .IN2(g2741), .Q(n14547) );
  AND2X1 U14808 ( .IN1(n14548), .IN2(n3730), .Q(n14546) );
  XNOR2X1 U14809 ( .IN1(n14549), .IN2(g2748), .Q(n14548) );
  OR2X1 U14810 ( .IN1(n5349), .IN2(n3506), .Q(n14549) );
  OR2X1 U14811 ( .IN1(n14550), .IN2(n14551), .Q(g31871) );
  OR2X1 U14812 ( .IN1(n14552), .IN2(n14553), .Q(n14551) );
  AND2X1 U14813 ( .IN1(n14554), .IN2(n10749), .Q(n14553) );
  AND2X1 U14814 ( .IN1(n11214), .IN2(g1367), .Q(n14554) );
  OR2X1 U14815 ( .IN1(n14555), .IN2(n11213), .Q(n11214) );
  AND2X1 U14816 ( .IN1(n10459), .IN2(n13787), .Q(n14555) );
  AND2X1 U14817 ( .IN1(n10930), .IN2(g1361), .Q(n14552) );
  AND2X1 U14818 ( .IN1(n3733), .IN2(n14378), .Q(n14550) );
  OR2X1 U14819 ( .IN1(n14556), .IN2(n14557), .Q(g31870) );
  OR2X1 U14820 ( .IN1(n14558), .IN2(n14559), .Q(n14557) );
  AND2X1 U14821 ( .IN1(n3664), .IN2(n5674), .Q(n14559) );
  INVX0 U14822 ( .INP(n14560), .ZN(n14558) );
  OR2X1 U14823 ( .IN1(n14561), .IN2(n5674), .Q(n14560) );
  OR2X1 U14824 ( .IN1(n13799), .IN2(n3664), .Q(n14561) );
  AND2X1 U14825 ( .IN1(n10930), .IN2(g1259), .Q(n14556) );
  OR2X1 U14826 ( .IN1(n14562), .IN2(n14563), .Q(g31869) );
  OR2X1 U14827 ( .IN1(n14564), .IN2(n14565), .Q(n14563) );
  AND2X1 U14828 ( .IN1(n14566), .IN2(n10748), .Q(n14565) );
  AND2X1 U14829 ( .IN1(n11098), .IN2(g1024), .Q(n14566) );
  OR2X1 U14830 ( .IN1(n14567), .IN2(n11097), .Q(n11098) );
  AND2X1 U14831 ( .IN1(n10458), .IN2(n13806), .Q(n14567) );
  AND2X1 U14832 ( .IN1(n10930), .IN2(g1018), .Q(n14564) );
  AND2X1 U14833 ( .IN1(n3738), .IN2(n14394), .Q(n14562) );
  OR2X1 U14834 ( .IN1(n14568), .IN2(n14569), .Q(g31868) );
  OR2X1 U14835 ( .IN1(n14570), .IN2(n14571), .Q(n14569) );
  AND2X1 U14836 ( .IN1(n3673), .IN2(n5673), .Q(n14571) );
  INVX0 U14837 ( .INP(n14572), .ZN(n14570) );
  OR2X1 U14838 ( .IN1(n14573), .IN2(n5673), .Q(n14572) );
  OR2X1 U14839 ( .IN1(n13818), .IN2(n3673), .Q(n14573) );
  AND2X1 U14840 ( .IN1(n10930), .IN2(g914), .Q(n14568) );
  OR2X1 U14841 ( .IN1(n14574), .IN2(n14575), .Q(g31867) );
  OR2X1 U14842 ( .IN1(n14576), .IN2(n14577), .Q(n14575) );
  INVX0 U14843 ( .INP(n14578), .ZN(n14577) );
  OR2X1 U14844 ( .IN1(n14579), .IN2(test_so2), .Q(n14578) );
  AND2X1 U14845 ( .IN1(n14580), .IN2(n14579), .Q(n14576) );
  INVX0 U14846 ( .INP(n3682), .ZN(n14579) );
  AND2X1 U14847 ( .IN1(n2404), .IN2(test_so2), .Q(n14580) );
  AND2X1 U14848 ( .IN1(n10930), .IN2(g744), .Q(n14574) );
  OR2X1 U14849 ( .IN1(n14581), .IN2(n14582), .Q(g31866) );
  OR2X1 U14850 ( .IN1(n14583), .IN2(n14584), .Q(n14582) );
  AND2X1 U14851 ( .IN1(n3684), .IN2(n5552), .Q(n14584) );
  AND2X1 U14852 ( .IN1(n14585), .IN2(g582), .Q(n14583) );
  AND2X1 U14853 ( .IN1(n2421), .IN2(n14586), .Q(n14585) );
  INVX0 U14854 ( .INP(n3684), .ZN(n14586) );
  AND2X1 U14855 ( .IN1(n10930), .IN2(g577), .Q(n14581) );
  OR2X1 U14856 ( .IN1(n14587), .IN2(n14588), .Q(g31865) );
  AND2X1 U14857 ( .IN1(n14589), .IN2(n10558), .Q(n14588) );
  AND2X1 U14858 ( .IN1(n10534), .IN2(test_so51), .Q(n14589) );
  AND2X1 U14859 ( .IN1(test_so55), .IN2(n14590), .Q(n14587) );
  OR2X1 U14860 ( .IN1(n10890), .IN2(n14591), .Q(n14590) );
  AND2X1 U14861 ( .IN1(n14592), .IN2(n10571), .Q(n14591) );
  OR2X1 U14862 ( .IN1(n14593), .IN2(n14594), .Q(g31864) );
  OR2X1 U14863 ( .IN1(n14595), .IN2(n14596), .Q(n14594) );
  AND2X1 U14864 ( .IN1(n3687), .IN2(n5561), .Q(n14596) );
  AND2X1 U14865 ( .IN1(n14597), .IN2(g164), .Q(n14595) );
  AND2X1 U14866 ( .IN1(n13055), .IN2(n14598), .Q(n14597) );
  INVX0 U14867 ( .INP(n3687), .ZN(n14598) );
  AND2X1 U14868 ( .IN1(test_so73), .IN2(n14599), .Q(n3687) );
  AND2X1 U14869 ( .IN1(n14600), .IN2(n14601), .Q(n14599) );
  INVX0 U14870 ( .INP(n14602), .ZN(n14601) );
  AND2X1 U14871 ( .IN1(test_so73), .IN2(n10894), .Q(n14593) );
  AND2X1 U14872 ( .IN1(g1668), .IN2(n5549), .Q(g31862) );
  OR2X1 U14873 ( .IN1(n14603), .IN2(n14604), .Q(g31793) );
  AND2X1 U14874 ( .IN1(n11706), .IN2(n14605), .Q(n14604) );
  AND2X1 U14875 ( .IN1(n14606), .IN2(n10564), .Q(n14605) );
  OR2X1 U14876 ( .IN1(n14607), .IN2(n14608), .Q(n14606) );
  AND2X1 U14877 ( .IN1(n11707), .IN2(n11709), .Q(n14608) );
  AND2X1 U14878 ( .IN1(n14609), .IN2(n10484), .Q(n14607) );
  AND2X1 U14879 ( .IN1(n14610), .IN2(n14611), .Q(n14609) );
  OR2X1 U14880 ( .IN1(n14612), .IN2(n14613), .Q(n14611) );
  OR2X1 U14881 ( .IN1(n11707), .IN2(n11709), .Q(n14610) );
  AND2X1 U14882 ( .IN1(n10456), .IN2(n14614), .Q(n11706) );
  AND2X1 U14883 ( .IN1(n14615), .IN2(n14616), .Q(n14603) );
  AND2X1 U14884 ( .IN1(n14617), .IN2(n11709), .Q(n14616) );
  OR2X1 U14885 ( .IN1(n14618), .IN2(n14614), .Q(n14617) );
  AND2X1 U14886 ( .IN1(n14619), .IN2(n14620), .Q(n14614) );
  AND2X1 U14887 ( .IN1(n14621), .IN2(n10456), .Q(n14618) );
  AND2X1 U14888 ( .IN1(n14622), .IN2(n10564), .Q(n14621) );
  OR2X1 U14889 ( .IN1(n14623), .IN2(n14620), .Q(n14622) );
  AND2X1 U14890 ( .IN1(n14624), .IN2(n14625), .Q(n14620) );
  OR2X1 U14891 ( .IN1(n14626), .IN2(n10875), .Q(n14625) );
  AND2X1 U14892 ( .IN1(n14627), .IN2(n14628), .Q(n14623) );
  OR2X1 U14893 ( .IN1(n10521), .IN2(n10522), .Q(n14628) );
  AND2X1 U14894 ( .IN1(n14629), .IN2(n14619), .Q(n14627) );
  OR2X1 U14895 ( .IN1(n14626), .IN2(n14624), .Q(n14629) );
  AND2X1 U14896 ( .IN1(n10522), .IN2(n10521), .Q(n14626) );
  AND2X1 U14897 ( .IN1(n11707), .IN2(n14630), .Q(n14615) );
  AND2X1 U14898 ( .IN1(n14613), .IN2(n14612), .Q(n11707) );
  OR2X1 U14899 ( .IN1(n10476), .IN2(n13094), .Q(g31665) );
  OR2X1 U14900 ( .IN1(n5488), .IN2(n13094), .Q(g31656) );
  INVX0 U14901 ( .INP(g113), .ZN(n13094) );
  OR2X1 U14902 ( .IN1(n14631), .IN2(n14632), .Q(g30563) );
  OR2X1 U14903 ( .IN1(n14633), .IN2(n14634), .Q(n14632) );
  AND2X1 U14904 ( .IN1(n3765), .IN2(n13075), .Q(n14634) );
  AND2X1 U14905 ( .IN1(n14635), .IN2(g6657), .Q(n14633) );
  AND2X1 U14906 ( .IN1(n10930), .IN2(g6653), .Q(n14631) );
  OR2X1 U14907 ( .IN1(n14636), .IN2(n14637), .Q(g30562) );
  OR2X1 U14908 ( .IN1(n14638), .IN2(n14639), .Q(n14637) );
  AND2X1 U14909 ( .IN1(n10930), .IN2(g6649), .Q(n14639) );
  INVX0 U14910 ( .INP(n14640), .ZN(n14638) );
  OR2X1 U14911 ( .IN1(n14641), .IN2(n10875), .Q(n14640) );
  OR2X1 U14912 ( .IN1(n14642), .IN2(n10368), .Q(n14641) );
  AND2X1 U14913 ( .IN1(n14642), .IN2(n3765), .Q(n14636) );
  AND2X1 U14914 ( .IN1(g6561), .IN2(n13876), .Q(n14642) );
  OR2X1 U14915 ( .IN1(n14643), .IN2(n14644), .Q(g30561) );
  OR2X1 U14916 ( .IN1(n14645), .IN2(n14646), .Q(n14644) );
  AND2X1 U14917 ( .IN1(n10930), .IN2(g6645), .Q(n14646) );
  INVX0 U14918 ( .INP(n14647), .ZN(n14645) );
  OR2X1 U14919 ( .IN1(n14648), .IN2(n10876), .Q(n14647) );
  OR2X1 U14920 ( .IN1(n13874), .IN2(n10343), .Q(n14648) );
  AND2X1 U14921 ( .IN1(n13874), .IN2(n3765), .Q(n14643) );
  AND2X1 U14922 ( .IN1(g6561), .IN2(n14649), .Q(n13874) );
  OR2X1 U14923 ( .IN1(n14650), .IN2(n14651), .Q(g30560) );
  OR2X1 U14924 ( .IN1(n14652), .IN2(n14653), .Q(n14651) );
  AND2X1 U14925 ( .IN1(n10930), .IN2(g6641), .Q(n14653) );
  INVX0 U14926 ( .INP(n14654), .ZN(n14652) );
  OR2X1 U14927 ( .IN1(n14655), .IN2(n10877), .Q(n14654) );
  OR2X1 U14928 ( .IN1(n14656), .IN2(n10313), .Q(n14655) );
  AND2X1 U14929 ( .IN1(n14656), .IN2(n3765), .Q(n14650) );
  AND2X1 U14930 ( .IN1(g6561), .IN2(n14657), .Q(n14656) );
  OR2X1 U14931 ( .IN1(n14658), .IN2(n14659), .Q(g30559) );
  OR2X1 U14932 ( .IN1(n14660), .IN2(n14661), .Q(n14659) );
  AND2X1 U14933 ( .IN1(n14662), .IN2(n10747), .Q(n14661) );
  AND2X1 U14934 ( .IN1(n14663), .IN2(g6653), .Q(n14662) );
  OR2X1 U14935 ( .IN1(n3776), .IN2(n3404), .Q(n14663) );
  AND2X1 U14936 ( .IN1(n10931), .IN2(g6637), .Q(n14660) );
  AND2X1 U14937 ( .IN1(n3774), .IN2(n14664), .Q(n14658) );
  OR2X1 U14938 ( .IN1(n14665), .IN2(n14666), .Q(g30558) );
  OR2X1 U14939 ( .IN1(n14667), .IN2(n14668), .Q(n14666) );
  AND2X1 U14940 ( .IN1(n14669), .IN2(n10747), .Q(n14668) );
  AND2X1 U14941 ( .IN1(n14670), .IN2(g6649), .Q(n14669) );
  OR2X1 U14942 ( .IN1(n3768), .IN2(n3404), .Q(n14670) );
  AND2X1 U14943 ( .IN1(n10931), .IN2(g6633), .Q(n14667) );
  AND2X1 U14944 ( .IN1(n3774), .IN2(n13876), .Q(n14665) );
  OR2X1 U14945 ( .IN1(n14671), .IN2(n14672), .Q(g30557) );
  OR2X1 U14946 ( .IN1(n14673), .IN2(n14674), .Q(n14672) );
  AND2X1 U14947 ( .IN1(n14675), .IN2(n10748), .Q(n14674) );
  AND2X1 U14948 ( .IN1(n14676), .IN2(g6645), .Q(n14675) );
  OR2X1 U14949 ( .IN1(n3770), .IN2(n3404), .Q(n14676) );
  AND2X1 U14950 ( .IN1(n10931), .IN2(g6629), .Q(n14673) );
  AND2X1 U14951 ( .IN1(n3774), .IN2(n14649), .Q(n14671) );
  OR2X1 U14952 ( .IN1(n14677), .IN2(n14678), .Q(g30556) );
  OR2X1 U14953 ( .IN1(n14679), .IN2(n14680), .Q(n14678) );
  AND2X1 U14954 ( .IN1(n14681), .IN2(n10747), .Q(n14680) );
  AND2X1 U14955 ( .IN1(n14682), .IN2(g6641), .Q(n14681) );
  OR2X1 U14956 ( .IN1(n3773), .IN2(n3404), .Q(n14682) );
  INVX0 U14957 ( .INP(n13885), .ZN(n3404) );
  AND2X1 U14958 ( .IN1(g6555), .IN2(g6549), .Q(n13885) );
  AND2X1 U14959 ( .IN1(n10931), .IN2(g6625), .Q(n14679) );
  AND2X1 U14960 ( .IN1(n3774), .IN2(n14657), .Q(n14677) );
  OR2X1 U14961 ( .IN1(n14683), .IN2(n14684), .Q(g30555) );
  OR2X1 U14962 ( .IN1(n14685), .IN2(n14686), .Q(n14684) );
  AND2X1 U14963 ( .IN1(n14687), .IN2(n10748), .Q(n14686) );
  AND2X1 U14964 ( .IN1(n14688), .IN2(g6637), .Q(n14687) );
  OR2X1 U14965 ( .IN1(n3776), .IN2(n3406), .Q(n14688) );
  AND2X1 U14966 ( .IN1(n10931), .IN2(g6621), .Q(n14685) );
  AND2X1 U14967 ( .IN1(n3780), .IN2(n14664), .Q(n14683) );
  OR2X1 U14968 ( .IN1(n14689), .IN2(n14690), .Q(g30554) );
  OR2X1 U14969 ( .IN1(n14691), .IN2(n14692), .Q(n14690) );
  AND2X1 U14970 ( .IN1(n14693), .IN2(n10748), .Q(n14692) );
  AND2X1 U14971 ( .IN1(n14694), .IN2(g6633), .Q(n14693) );
  OR2X1 U14972 ( .IN1(n3768), .IN2(n3406), .Q(n14694) );
  AND2X1 U14973 ( .IN1(n10931), .IN2(g6617), .Q(n14691) );
  AND2X1 U14974 ( .IN1(n3780), .IN2(n13876), .Q(n14689) );
  OR2X1 U14975 ( .IN1(n14695), .IN2(n14696), .Q(g30553) );
  OR2X1 U14976 ( .IN1(n14697), .IN2(n14698), .Q(n14696) );
  AND2X1 U14977 ( .IN1(n14699), .IN2(n10748), .Q(n14698) );
  AND2X1 U14978 ( .IN1(n14700), .IN2(g6629), .Q(n14699) );
  OR2X1 U14979 ( .IN1(n3770), .IN2(n3406), .Q(n14700) );
  AND2X1 U14980 ( .IN1(n10931), .IN2(g6613), .Q(n14697) );
  AND2X1 U14981 ( .IN1(n3780), .IN2(n14649), .Q(n14695) );
  OR2X1 U14982 ( .IN1(n14701), .IN2(n14702), .Q(g30552) );
  OR2X1 U14983 ( .IN1(n14703), .IN2(n14704), .Q(n14702) );
  AND2X1 U14984 ( .IN1(n14705), .IN2(n10747), .Q(n14704) );
  AND2X1 U14985 ( .IN1(n14706), .IN2(g6625), .Q(n14705) );
  OR2X1 U14986 ( .IN1(n3773), .IN2(n3406), .Q(n14706) );
  OR2X1 U14987 ( .IN1(n10431), .IN2(g6549), .Q(n3406) );
  AND2X1 U14988 ( .IN1(n10931), .IN2(g6609), .Q(n14703) );
  AND2X1 U14989 ( .IN1(n3780), .IN2(n14657), .Q(n14701) );
  OR2X1 U14990 ( .IN1(n14707), .IN2(n14708), .Q(g30551) );
  OR2X1 U14991 ( .IN1(n14709), .IN2(n14710), .Q(n14708) );
  AND2X1 U14992 ( .IN1(n14711), .IN2(n10747), .Q(n14710) );
  AND2X1 U14993 ( .IN1(n14712), .IN2(g6621), .Q(n14711) );
  OR2X1 U14994 ( .IN1(n3776), .IN2(n3407), .Q(n14712) );
  INVX0 U14995 ( .INP(n14664), .ZN(n3776) );
  AND2X1 U14996 ( .IN1(n10931), .IN2(g6601), .Q(n14709) );
  AND2X1 U14997 ( .IN1(n3785), .IN2(n14664), .Q(n14707) );
  OR2X1 U14998 ( .IN1(n14713), .IN2(n14714), .Q(g30550) );
  OR2X1 U14999 ( .IN1(n14715), .IN2(n14716), .Q(n14714) );
  AND2X1 U15000 ( .IN1(n14717), .IN2(n10747), .Q(n14716) );
  AND2X1 U15001 ( .IN1(n14718), .IN2(g6617), .Q(n14717) );
  OR2X1 U15002 ( .IN1(n3768), .IN2(n3407), .Q(n14718) );
  INVX0 U15003 ( .INP(n13876), .ZN(n3768) );
  AND2X1 U15004 ( .IN1(n10931), .IN2(g6593), .Q(n14715) );
  AND2X1 U15005 ( .IN1(n3785), .IN2(n13876), .Q(n14713) );
  AND2X1 U15006 ( .IN1(g6573), .IN2(n5386), .Q(n13876) );
  OR2X1 U15007 ( .IN1(n14719), .IN2(n14720), .Q(g30549) );
  OR2X1 U15008 ( .IN1(n14721), .IN2(n14722), .Q(n14720) );
  AND2X1 U15009 ( .IN1(n14723), .IN2(n10747), .Q(n14722) );
  AND2X1 U15010 ( .IN1(n14724), .IN2(g6613), .Q(n14723) );
  OR2X1 U15011 ( .IN1(n3770), .IN2(n3407), .Q(n14724) );
  INVX0 U15012 ( .INP(n14649), .ZN(n3770) );
  AND2X1 U15013 ( .IN1(test_so71), .IN2(n10893), .Q(n14721) );
  AND2X1 U15014 ( .IN1(n3785), .IN2(n14649), .Q(n14719) );
  AND2X1 U15015 ( .IN1(g6565), .IN2(n5563), .Q(n14649) );
  OR2X1 U15016 ( .IN1(n14725), .IN2(n14726), .Q(g30548) );
  OR2X1 U15017 ( .IN1(n14727), .IN2(n14728), .Q(n14726) );
  AND2X1 U15018 ( .IN1(n14729), .IN2(n10740), .Q(n14728) );
  AND2X1 U15019 ( .IN1(n14730), .IN2(g6609), .Q(n14729) );
  OR2X1 U15020 ( .IN1(n3773), .IN2(n3407), .Q(n14730) );
  OR2X1 U15021 ( .IN1(n5571), .IN2(g6555), .Q(n3407) );
  INVX0 U15022 ( .INP(n14657), .ZN(n3773) );
  AND2X1 U15023 ( .IN1(n10931), .IN2(g6581), .Q(n14727) );
  AND2X1 U15024 ( .IN1(n3785), .IN2(n14657), .Q(n14725) );
  AND2X1 U15025 ( .IN1(n5386), .IN2(n5563), .Q(n14657) );
  OR2X1 U15026 ( .IN1(n14731), .IN2(n14732), .Q(g30547) );
  OR2X1 U15027 ( .IN1(n14733), .IN2(n14734), .Q(n14732) );
  AND2X1 U15028 ( .IN1(n3790), .IN2(n3765), .Q(n14734) );
  AND2X1 U15029 ( .IN1(n14735), .IN2(n14736), .Q(n14733) );
  INVX0 U15030 ( .INP(n3790), .ZN(n14736) );
  AND2X1 U15031 ( .IN1(n10823), .IN2(g6601), .Q(n14735) );
  AND2X1 U15032 ( .IN1(n10931), .IN2(g6605), .Q(n14731) );
  OR2X1 U15033 ( .IN1(n14737), .IN2(n14738), .Q(g30546) );
  OR2X1 U15034 ( .IN1(n14739), .IN2(n14740), .Q(n14738) );
  AND2X1 U15035 ( .IN1(n3793), .IN2(n3765), .Q(n14740) );
  AND2X1 U15036 ( .IN1(n14741), .IN2(n14742), .Q(n14739) );
  INVX0 U15037 ( .INP(n3793), .ZN(n14742) );
  AND2X1 U15038 ( .IN1(n10823), .IN2(g6593), .Q(n14741) );
  AND2X1 U15039 ( .IN1(n10931), .IN2(g6597), .Q(n14737) );
  OR2X1 U15040 ( .IN1(n14743), .IN2(n14744), .Q(g30545) );
  OR2X1 U15041 ( .IN1(n14745), .IN2(n14746), .Q(n14744) );
  AND2X1 U15042 ( .IN1(n3795), .IN2(n3765), .Q(n14746) );
  AND2X1 U15043 ( .IN1(n14747), .IN2(n14748), .Q(n14745) );
  INVX0 U15044 ( .INP(n3795), .ZN(n14748) );
  AND2X1 U15045 ( .IN1(test_so71), .IN2(n10754), .Q(n14747) );
  AND2X1 U15046 ( .IN1(n10931), .IN2(g6589), .Q(n14743) );
  OR2X1 U15047 ( .IN1(n14749), .IN2(n14750), .Q(g30544) );
  OR2X1 U15048 ( .IN1(n14751), .IN2(n14752), .Q(n14750) );
  AND2X1 U15049 ( .IN1(n3797), .IN2(n3765), .Q(n14752) );
  AND2X1 U15050 ( .IN1(n14753), .IN2(n14754), .Q(n14751) );
  INVX0 U15051 ( .INP(n3797), .ZN(n14754) );
  AND2X1 U15052 ( .IN1(n10823), .IN2(g6581), .Q(n14753) );
  AND2X1 U15053 ( .IN1(n10931), .IN2(g6573), .Q(n14749) );
  AND2X1 U15054 ( .IN1(n13879), .IN2(n5571), .Q(g30543) );
  AND2X1 U15055 ( .IN1(n5646), .IN2(n14755), .Q(n13879) );
  AND2X1 U15056 ( .IN1(n10824), .IN2(n13871), .Q(n14755) );
  OR2X1 U15057 ( .IN1(n14756), .IN2(n14757), .Q(n13871) );
  OR2X1 U15058 ( .IN1(n14758), .IN2(n14759), .Q(g30542) );
  OR2X1 U15059 ( .IN1(n14760), .IN2(n14761), .Q(n14759) );
  AND2X1 U15060 ( .IN1(n13092), .IN2(n3765), .Q(n14761) );
  AND2X1 U15061 ( .IN1(n14762), .IN2(g6311), .Q(n14760) );
  AND2X1 U15062 ( .IN1(n10931), .IN2(g6307), .Q(n14758) );
  OR2X1 U15063 ( .IN1(n14763), .IN2(n14764), .Q(g30541) );
  OR2X1 U15064 ( .IN1(n14765), .IN2(n14766), .Q(n14764) );
  AND2X1 U15065 ( .IN1(n10931), .IN2(g6303), .Q(n14766) );
  INVX0 U15066 ( .INP(n14767), .ZN(n14765) );
  OR2X1 U15067 ( .IN1(n14768), .IN2(n10877), .Q(n14767) );
  OR2X1 U15068 ( .IN1(n14769), .IN2(n10376), .Q(n14768) );
  AND2X1 U15069 ( .IN1(n14769), .IN2(n3765), .Q(n14763) );
  AND2X1 U15070 ( .IN1(g6215), .IN2(n13899), .Q(n14769) );
  OR2X1 U15071 ( .IN1(n14770), .IN2(n14771), .Q(g30540) );
  OR2X1 U15072 ( .IN1(n14772), .IN2(n14773), .Q(n14771) );
  AND2X1 U15073 ( .IN1(n10931), .IN2(g6299), .Q(n14773) );
  INVX0 U15074 ( .INP(n14774), .ZN(n14772) );
  OR2X1 U15075 ( .IN1(n14775), .IN2(n10877), .Q(n14774) );
  OR2X1 U15076 ( .IN1(n13897), .IN2(n10351), .Q(n14775) );
  AND2X1 U15077 ( .IN1(n13897), .IN2(n3765), .Q(n14770) );
  AND2X1 U15078 ( .IN1(g6215), .IN2(n14776), .Q(n13897) );
  OR2X1 U15079 ( .IN1(n14777), .IN2(n14778), .Q(g30539) );
  OR2X1 U15080 ( .IN1(n14779), .IN2(n14780), .Q(n14778) );
  AND2X1 U15081 ( .IN1(n10931), .IN2(g6295), .Q(n14780) );
  INVX0 U15082 ( .INP(n14781), .ZN(n14779) );
  OR2X1 U15083 ( .IN1(n14782), .IN2(n10877), .Q(n14781) );
  OR2X1 U15084 ( .IN1(n14783), .IN2(n10317), .Q(n14782) );
  AND2X1 U15085 ( .IN1(n14783), .IN2(n3765), .Q(n14777) );
  AND2X1 U15086 ( .IN1(g6215), .IN2(n14784), .Q(n14783) );
  OR2X1 U15087 ( .IN1(n14785), .IN2(n14786), .Q(g30538) );
  OR2X1 U15088 ( .IN1(n14787), .IN2(n14788), .Q(n14786) );
  AND2X1 U15089 ( .IN1(n14789), .IN2(n10754), .Q(n14788) );
  AND2X1 U15090 ( .IN1(n14790), .IN2(g6307), .Q(n14789) );
  OR2X1 U15091 ( .IN1(n3810), .IN2(n3414), .Q(n14790) );
  AND2X1 U15092 ( .IN1(n10932), .IN2(g6291), .Q(n14787) );
  AND2X1 U15093 ( .IN1(n3808), .IN2(n14791), .Q(n14785) );
  OR2X1 U15094 ( .IN1(n14792), .IN2(n14793), .Q(g30537) );
  OR2X1 U15095 ( .IN1(n14794), .IN2(n14795), .Q(n14793) );
  AND2X1 U15096 ( .IN1(n14796), .IN2(n10754), .Q(n14795) );
  AND2X1 U15097 ( .IN1(n14797), .IN2(g6303), .Q(n14796) );
  OR2X1 U15098 ( .IN1(n3802), .IN2(n3414), .Q(n14797) );
  AND2X1 U15099 ( .IN1(n10932), .IN2(g6287), .Q(n14794) );
  AND2X1 U15100 ( .IN1(n3808), .IN2(n13899), .Q(n14792) );
  OR2X1 U15101 ( .IN1(n14798), .IN2(n14799), .Q(g30536) );
  OR2X1 U15102 ( .IN1(n14800), .IN2(n14801), .Q(n14799) );
  AND2X1 U15103 ( .IN1(n14802), .IN2(n10754), .Q(n14801) );
  AND2X1 U15104 ( .IN1(n14803), .IN2(g6299), .Q(n14802) );
  OR2X1 U15105 ( .IN1(n3804), .IN2(n3414), .Q(n14803) );
  AND2X1 U15106 ( .IN1(n10932), .IN2(g6283), .Q(n14800) );
  AND2X1 U15107 ( .IN1(n3808), .IN2(n14776), .Q(n14798) );
  OR2X1 U15108 ( .IN1(n14804), .IN2(n14805), .Q(g30535) );
  OR2X1 U15109 ( .IN1(n14806), .IN2(n14807), .Q(n14805) );
  AND2X1 U15110 ( .IN1(n14808), .IN2(n10755), .Q(n14807) );
  AND2X1 U15111 ( .IN1(n14809), .IN2(g6295), .Q(n14808) );
  OR2X1 U15112 ( .IN1(n3807), .IN2(n3414), .Q(n14809) );
  INVX0 U15113 ( .INP(n13908), .ZN(n3414) );
  AND2X1 U15114 ( .IN1(g6209), .IN2(g6203), .Q(n13908) );
  AND2X1 U15115 ( .IN1(n10932), .IN2(g6279), .Q(n14806) );
  AND2X1 U15116 ( .IN1(n3808), .IN2(n14784), .Q(n14804) );
  OR2X1 U15117 ( .IN1(n14810), .IN2(n14811), .Q(g30534) );
  OR2X1 U15118 ( .IN1(n14812), .IN2(n14813), .Q(n14811) );
  AND2X1 U15119 ( .IN1(n14814), .IN2(n10755), .Q(n14813) );
  AND2X1 U15120 ( .IN1(n14815), .IN2(g6291), .Q(n14814) );
  OR2X1 U15121 ( .IN1(n3810), .IN2(n3416), .Q(n14815) );
  AND2X1 U15122 ( .IN1(n10932), .IN2(g6275), .Q(n14812) );
  AND2X1 U15123 ( .IN1(n3814), .IN2(n14791), .Q(n14810) );
  OR2X1 U15124 ( .IN1(n14816), .IN2(n14817), .Q(g30533) );
  OR2X1 U15125 ( .IN1(n14818), .IN2(n14819), .Q(n14817) );
  AND2X1 U15126 ( .IN1(n14820), .IN2(n10755), .Q(n14819) );
  AND2X1 U15127 ( .IN1(n14821), .IN2(g6287), .Q(n14820) );
  OR2X1 U15128 ( .IN1(n3802), .IN2(n3416), .Q(n14821) );
  AND2X1 U15129 ( .IN1(n10932), .IN2(g6271), .Q(n14818) );
  AND2X1 U15130 ( .IN1(n3814), .IN2(n13899), .Q(n14816) );
  OR2X1 U15131 ( .IN1(n14822), .IN2(n14823), .Q(g30532) );
  OR2X1 U15132 ( .IN1(n14824), .IN2(n14825), .Q(n14823) );
  AND2X1 U15133 ( .IN1(n14826), .IN2(n10755), .Q(n14825) );
  AND2X1 U15134 ( .IN1(n14827), .IN2(g6283), .Q(n14826) );
  OR2X1 U15135 ( .IN1(n3804), .IN2(n3416), .Q(n14827) );
  AND2X1 U15136 ( .IN1(n10932), .IN2(g6267), .Q(n14824) );
  AND2X1 U15137 ( .IN1(n3814), .IN2(n14776), .Q(n14822) );
  OR2X1 U15138 ( .IN1(n14828), .IN2(n14829), .Q(g30531) );
  OR2X1 U15139 ( .IN1(n14830), .IN2(n14831), .Q(n14829) );
  AND2X1 U15140 ( .IN1(n14832), .IN2(n10755), .Q(n14831) );
  AND2X1 U15141 ( .IN1(n14833), .IN2(g6279), .Q(n14832) );
  OR2X1 U15142 ( .IN1(n3807), .IN2(n3416), .Q(n14833) );
  OR2X1 U15143 ( .IN1(n10428), .IN2(g6203), .Q(n3416) );
  AND2X1 U15144 ( .IN1(n10932), .IN2(g6263), .Q(n14830) );
  AND2X1 U15145 ( .IN1(n3814), .IN2(n14784), .Q(n14828) );
  OR2X1 U15146 ( .IN1(n14834), .IN2(n14835), .Q(g30530) );
  OR2X1 U15147 ( .IN1(n14836), .IN2(n14837), .Q(n14835) );
  AND2X1 U15148 ( .IN1(n14838), .IN2(n10755), .Q(n14837) );
  AND2X1 U15149 ( .IN1(n14839), .IN2(g6275), .Q(n14838) );
  OR2X1 U15150 ( .IN1(n3810), .IN2(n3417), .Q(n14839) );
  INVX0 U15151 ( .INP(n14791), .ZN(n3810) );
  AND2X1 U15152 ( .IN1(n10932), .IN2(g6255), .Q(n14836) );
  AND2X1 U15153 ( .IN1(n3819), .IN2(n14791), .Q(n14834) );
  OR2X1 U15154 ( .IN1(n14840), .IN2(n14841), .Q(g30529) );
  OR2X1 U15155 ( .IN1(n14842), .IN2(n14843), .Q(n14841) );
  AND2X1 U15156 ( .IN1(n14844), .IN2(n10755), .Q(n14843) );
  AND2X1 U15157 ( .IN1(n14845), .IN2(g6271), .Q(n14844) );
  OR2X1 U15158 ( .IN1(n3802), .IN2(n3417), .Q(n14845) );
  INVX0 U15159 ( .INP(n13899), .ZN(n3802) );
  AND2X1 U15160 ( .IN1(n10924), .IN2(g6247), .Q(n14842) );
  AND2X1 U15161 ( .IN1(n3819), .IN2(n13899), .Q(n14840) );
  AND2X1 U15162 ( .IN1(g6227), .IN2(n5385), .Q(n13899) );
  OR2X1 U15163 ( .IN1(n14846), .IN2(n14847), .Q(g30528) );
  OR2X1 U15164 ( .IN1(n14848), .IN2(n14849), .Q(n14847) );
  AND2X1 U15165 ( .IN1(n14850), .IN2(n10755), .Q(n14849) );
  AND2X1 U15166 ( .IN1(n14851), .IN2(g6267), .Q(n14850) );
  OR2X1 U15167 ( .IN1(n3804), .IN2(n3417), .Q(n14851) );
  INVX0 U15168 ( .INP(n14776), .ZN(n3804) );
  AND2X1 U15169 ( .IN1(n10921), .IN2(g6239), .Q(n14848) );
  AND2X1 U15170 ( .IN1(n3819), .IN2(n14776), .Q(n14846) );
  AND2X1 U15171 ( .IN1(g6219), .IN2(n5568), .Q(n14776) );
  OR2X1 U15172 ( .IN1(n14852), .IN2(n14853), .Q(g30527) );
  OR2X1 U15173 ( .IN1(n14854), .IN2(n14855), .Q(n14853) );
  AND2X1 U15174 ( .IN1(n14856), .IN2(n10755), .Q(n14855) );
  AND2X1 U15175 ( .IN1(n14857), .IN2(g6263), .Q(n14856) );
  OR2X1 U15176 ( .IN1(n3807), .IN2(n3417), .Q(n14857) );
  OR2X1 U15177 ( .IN1(n5574), .IN2(g6209), .Q(n3417) );
  INVX0 U15178 ( .INP(n14784), .ZN(n3807) );
  AND2X1 U15179 ( .IN1(n10921), .IN2(g6235), .Q(n14854) );
  AND2X1 U15180 ( .IN1(n3819), .IN2(n14784), .Q(n14852) );
  AND2X1 U15181 ( .IN1(n5385), .IN2(n5568), .Q(n14784) );
  OR2X1 U15182 ( .IN1(n14858), .IN2(n14859), .Q(g30526) );
  OR2X1 U15183 ( .IN1(n14860), .IN2(n14861), .Q(n14859) );
  AND2X1 U15184 ( .IN1(n3824), .IN2(n3765), .Q(n14861) );
  AND2X1 U15185 ( .IN1(n14862), .IN2(n14863), .Q(n14860) );
  INVX0 U15186 ( .INP(n3824), .ZN(n14863) );
  AND2X1 U15187 ( .IN1(n10825), .IN2(g6255), .Q(n14862) );
  AND2X1 U15188 ( .IN1(n10921), .IN2(g6259), .Q(n14858) );
  OR2X1 U15189 ( .IN1(n14864), .IN2(n14865), .Q(g30525) );
  OR2X1 U15190 ( .IN1(n14866), .IN2(n14867), .Q(n14865) );
  AND2X1 U15191 ( .IN1(n3827), .IN2(n3765), .Q(n14867) );
  AND2X1 U15192 ( .IN1(n14868), .IN2(n14869), .Q(n14866) );
  INVX0 U15193 ( .INP(n3827), .ZN(n14869) );
  AND2X1 U15194 ( .IN1(n10825), .IN2(g6247), .Q(n14868) );
  AND2X1 U15195 ( .IN1(n10921), .IN2(g6251), .Q(n14864) );
  OR2X1 U15196 ( .IN1(n14870), .IN2(n14871), .Q(g30524) );
  OR2X1 U15197 ( .IN1(n14872), .IN2(n14873), .Q(n14871) );
  AND2X1 U15198 ( .IN1(n3829), .IN2(n3765), .Q(n14873) );
  AND2X1 U15199 ( .IN1(n14874), .IN2(n14875), .Q(n14872) );
  INVX0 U15200 ( .INP(n3829), .ZN(n14875) );
  AND2X1 U15201 ( .IN1(n10825), .IN2(g6239), .Q(n14874) );
  AND2X1 U15202 ( .IN1(n10921), .IN2(g6243), .Q(n14870) );
  OR2X1 U15203 ( .IN1(n14876), .IN2(n14877), .Q(g30523) );
  OR2X1 U15204 ( .IN1(n14878), .IN2(n14879), .Q(n14877) );
  AND2X1 U15205 ( .IN1(n3831), .IN2(n3765), .Q(n14879) );
  AND2X1 U15206 ( .IN1(n14880), .IN2(n14881), .Q(n14878) );
  INVX0 U15207 ( .INP(n3831), .ZN(n14881) );
  AND2X1 U15208 ( .IN1(n10825), .IN2(g6235), .Q(n14880) );
  AND2X1 U15209 ( .IN1(n10921), .IN2(g6227), .Q(n14876) );
  AND2X1 U15210 ( .IN1(n13902), .IN2(n5574), .Q(g30522) );
  AND2X1 U15211 ( .IN1(n5651), .IN2(n14882), .Q(n13902) );
  AND2X1 U15212 ( .IN1(n10826), .IN2(n13894), .Q(n14882) );
  OR2X1 U15213 ( .IN1(n14883), .IN2(n14884), .Q(n13894) );
  OR2X1 U15214 ( .IN1(n14885), .IN2(n14886), .Q(g30521) );
  OR2X1 U15215 ( .IN1(n14887), .IN2(n14888), .Q(n14886) );
  AND2X1 U15216 ( .IN1(n13091), .IN2(n3765), .Q(n14888) );
  AND2X1 U15217 ( .IN1(test_so13), .IN2(n14889), .Q(n14887) );
  AND2X1 U15218 ( .IN1(n10921), .IN2(g5961), .Q(n14885) );
  OR2X1 U15219 ( .IN1(n14890), .IN2(n14891), .Q(g30520) );
  OR2X1 U15220 ( .IN1(n14892), .IN2(n14893), .Q(n14891) );
  AND2X1 U15221 ( .IN1(n10922), .IN2(g5957), .Q(n14893) );
  INVX0 U15222 ( .INP(n14894), .ZN(n14892) );
  OR2X1 U15223 ( .IN1(n14895), .IN2(n10875), .Q(n14894) );
  OR2X1 U15224 ( .IN1(n14896), .IN2(n10356), .Q(n14895) );
  AND2X1 U15225 ( .IN1(n14896), .IN2(n3765), .Q(n14890) );
  AND2X1 U15226 ( .IN1(g5869), .IN2(n13922), .Q(n14896) );
  OR2X1 U15227 ( .IN1(n14897), .IN2(n14898), .Q(g30519) );
  OR2X1 U15228 ( .IN1(n14899), .IN2(n14900), .Q(n14898) );
  AND2X1 U15229 ( .IN1(n10922), .IN2(g5953), .Q(n14900) );
  INVX0 U15230 ( .INP(n14901), .ZN(n14899) );
  OR2X1 U15231 ( .IN1(n14902), .IN2(n10876), .Q(n14901) );
  OR2X1 U15232 ( .IN1(n13920), .IN2(n10332), .Q(n14902) );
  AND2X1 U15233 ( .IN1(n13920), .IN2(n3765), .Q(n14897) );
  AND2X1 U15234 ( .IN1(g5869), .IN2(n14903), .Q(n13920) );
  OR2X1 U15235 ( .IN1(n14904), .IN2(n14905), .Q(g30518) );
  OR2X1 U15236 ( .IN1(n14906), .IN2(n14907), .Q(n14905) );
  AND2X1 U15237 ( .IN1(n10922), .IN2(g5949), .Q(n14907) );
  INVX0 U15238 ( .INP(n14908), .ZN(n14906) );
  OR2X1 U15239 ( .IN1(n14909), .IN2(n10875), .Q(n14908) );
  OR2X1 U15240 ( .IN1(n14910), .IN2(n10308), .Q(n14909) );
  AND2X1 U15241 ( .IN1(n14910), .IN2(n3765), .Q(n14904) );
  AND2X1 U15242 ( .IN1(g5869), .IN2(n14911), .Q(n14910) );
  OR2X1 U15243 ( .IN1(n14912), .IN2(n14913), .Q(g30517) );
  OR2X1 U15244 ( .IN1(n14914), .IN2(n14915), .Q(n14913) );
  AND2X1 U15245 ( .IN1(n14916), .IN2(n10756), .Q(n14915) );
  AND2X1 U15246 ( .IN1(n14917), .IN2(g5961), .Q(n14916) );
  OR2X1 U15247 ( .IN1(n3844), .IN2(n3424), .Q(n14917) );
  AND2X1 U15248 ( .IN1(n10922), .IN2(g5945), .Q(n14914) );
  AND2X1 U15249 ( .IN1(n3842), .IN2(n14918), .Q(n14912) );
  OR2X1 U15250 ( .IN1(n14919), .IN2(n14920), .Q(g30516) );
  OR2X1 U15251 ( .IN1(n14921), .IN2(n14922), .Q(n14920) );
  AND2X1 U15252 ( .IN1(n14923), .IN2(n10756), .Q(n14922) );
  AND2X1 U15253 ( .IN1(n14924), .IN2(g5957), .Q(n14923) );
  OR2X1 U15254 ( .IN1(n3836), .IN2(n3424), .Q(n14924) );
  AND2X1 U15255 ( .IN1(n10922), .IN2(g5941), .Q(n14921) );
  AND2X1 U15256 ( .IN1(n3842), .IN2(n13922), .Q(n14919) );
  OR2X1 U15257 ( .IN1(n14925), .IN2(n14926), .Q(g30515) );
  OR2X1 U15258 ( .IN1(n14927), .IN2(n14928), .Q(n14926) );
  AND2X1 U15259 ( .IN1(n14929), .IN2(n10756), .Q(n14928) );
  AND2X1 U15260 ( .IN1(n14930), .IN2(g5953), .Q(n14929) );
  OR2X1 U15261 ( .IN1(n3838), .IN2(n3424), .Q(n14930) );
  AND2X1 U15262 ( .IN1(n10922), .IN2(g5937), .Q(n14927) );
  AND2X1 U15263 ( .IN1(n3842), .IN2(n14903), .Q(n14925) );
  OR2X1 U15264 ( .IN1(n14931), .IN2(n14932), .Q(g30514) );
  OR2X1 U15265 ( .IN1(n14933), .IN2(n14934), .Q(n14932) );
  AND2X1 U15266 ( .IN1(n14935), .IN2(n10756), .Q(n14934) );
  AND2X1 U15267 ( .IN1(n14936), .IN2(g5949), .Q(n14935) );
  OR2X1 U15268 ( .IN1(n3841), .IN2(n3424), .Q(n14936) );
  INVX0 U15269 ( .INP(n13931), .ZN(n3424) );
  AND2X1 U15270 ( .IN1(g5863), .IN2(g5857), .Q(n13931) );
  AND2X1 U15271 ( .IN1(n10922), .IN2(g5933), .Q(n14933) );
  AND2X1 U15272 ( .IN1(n3842), .IN2(n14911), .Q(n14931) );
  OR2X1 U15273 ( .IN1(n14937), .IN2(n14938), .Q(g30513) );
  OR2X1 U15274 ( .IN1(n14939), .IN2(n14940), .Q(n14938) );
  AND2X1 U15275 ( .IN1(n14941), .IN2(n10756), .Q(n14940) );
  AND2X1 U15276 ( .IN1(n14942), .IN2(g5945), .Q(n14941) );
  OR2X1 U15277 ( .IN1(n3844), .IN2(n3426), .Q(n14942) );
  AND2X1 U15278 ( .IN1(n10922), .IN2(g5929), .Q(n14939) );
  AND2X1 U15279 ( .IN1(n3848), .IN2(n14918), .Q(n14937) );
  OR2X1 U15280 ( .IN1(n14943), .IN2(n14944), .Q(g30512) );
  OR2X1 U15281 ( .IN1(n14945), .IN2(n14946), .Q(n14944) );
  AND2X1 U15282 ( .IN1(n14947), .IN2(n10756), .Q(n14946) );
  AND2X1 U15283 ( .IN1(n14948), .IN2(g5941), .Q(n14947) );
  OR2X1 U15284 ( .IN1(n3836), .IN2(n3426), .Q(n14948) );
  AND2X1 U15285 ( .IN1(n10922), .IN2(g5925), .Q(n14945) );
  AND2X1 U15286 ( .IN1(n3848), .IN2(n13922), .Q(n14943) );
  OR2X1 U15287 ( .IN1(n14949), .IN2(n14950), .Q(g30511) );
  OR2X1 U15288 ( .IN1(n14951), .IN2(n14952), .Q(n14950) );
  AND2X1 U15289 ( .IN1(n14953), .IN2(n10756), .Q(n14952) );
  AND2X1 U15290 ( .IN1(n14954), .IN2(g5937), .Q(n14953) );
  OR2X1 U15291 ( .IN1(n3838), .IN2(n3426), .Q(n14954) );
  AND2X1 U15292 ( .IN1(n10922), .IN2(g5921), .Q(n14951) );
  AND2X1 U15293 ( .IN1(n3848), .IN2(n14903), .Q(n14949) );
  OR2X1 U15294 ( .IN1(n14955), .IN2(n14956), .Q(g30510) );
  OR2X1 U15295 ( .IN1(n14957), .IN2(n14958), .Q(n14956) );
  AND2X1 U15296 ( .IN1(n14959), .IN2(n10756), .Q(n14958) );
  AND2X1 U15297 ( .IN1(n14960), .IN2(g5933), .Q(n14959) );
  OR2X1 U15298 ( .IN1(n3841), .IN2(n3426), .Q(n14960) );
  OR2X1 U15299 ( .IN1(n10430), .IN2(g5857), .Q(n3426) );
  AND2X1 U15300 ( .IN1(test_so28), .IN2(n10895), .Q(n14957) );
  AND2X1 U15301 ( .IN1(n3848), .IN2(n14911), .Q(n14955) );
  OR2X1 U15302 ( .IN1(n14961), .IN2(n14962), .Q(g30509) );
  OR2X1 U15303 ( .IN1(n14963), .IN2(n14964), .Q(n14962) );
  AND2X1 U15304 ( .IN1(n14965), .IN2(n10756), .Q(n14964) );
  AND2X1 U15305 ( .IN1(n14966), .IN2(g5929), .Q(n14965) );
  OR2X1 U15306 ( .IN1(n3844), .IN2(n3427), .Q(n14966) );
  INVX0 U15307 ( .INP(n14918), .ZN(n3844) );
  AND2X1 U15308 ( .IN1(n10922), .IN2(g5909), .Q(n14963) );
  AND2X1 U15309 ( .IN1(n3853), .IN2(n14918), .Q(n14961) );
  OR2X1 U15310 ( .IN1(n14967), .IN2(n14968), .Q(g30508) );
  OR2X1 U15311 ( .IN1(n14969), .IN2(n14970), .Q(n14968) );
  AND2X1 U15312 ( .IN1(n14971), .IN2(n10757), .Q(n14970) );
  AND2X1 U15313 ( .IN1(n14972), .IN2(g5925), .Q(n14971) );
  OR2X1 U15314 ( .IN1(n3836), .IN2(n3427), .Q(n14972) );
  INVX0 U15315 ( .INP(n13922), .ZN(n3836) );
  AND2X1 U15316 ( .IN1(n10922), .IN2(g5901), .Q(n14969) );
  AND2X1 U15317 ( .IN1(n3853), .IN2(n13922), .Q(n14967) );
  AND2X1 U15318 ( .IN1(test_so36), .IN2(n5388), .Q(n13922) );
  OR2X1 U15319 ( .IN1(n14973), .IN2(n14974), .Q(g30507) );
  OR2X1 U15320 ( .IN1(n14975), .IN2(n14976), .Q(n14974) );
  AND2X1 U15321 ( .IN1(n14977), .IN2(n10757), .Q(n14976) );
  AND2X1 U15322 ( .IN1(n14978), .IN2(g5921), .Q(n14977) );
  OR2X1 U15323 ( .IN1(n3838), .IN2(n3427), .Q(n14978) );
  INVX0 U15324 ( .INP(n14903), .ZN(n3838) );
  AND2X1 U15325 ( .IN1(n10922), .IN2(g5893), .Q(n14975) );
  AND2X1 U15326 ( .IN1(n3853), .IN2(n14903), .Q(n14973) );
  AND2X1 U15327 ( .IN1(g5873), .IN2(n10576), .Q(n14903) );
  OR2X1 U15328 ( .IN1(n14979), .IN2(n14980), .Q(g30506) );
  OR2X1 U15329 ( .IN1(n14981), .IN2(n14982), .Q(n14980) );
  AND2X1 U15330 ( .IN1(n14983), .IN2(n10757), .Q(n14982) );
  AND2X1 U15331 ( .IN1(test_so28), .IN2(n14984), .Q(n14983) );
  OR2X1 U15332 ( .IN1(n3841), .IN2(n3427), .Q(n14984) );
  OR2X1 U15333 ( .IN1(n5573), .IN2(g5863), .Q(n3427) );
  INVX0 U15334 ( .INP(n14911), .ZN(n3841) );
  AND2X1 U15335 ( .IN1(n10922), .IN2(g5889), .Q(n14981) );
  AND2X1 U15336 ( .IN1(n3853), .IN2(n14911), .Q(n14979) );
  AND2X1 U15337 ( .IN1(n10576), .IN2(n5388), .Q(n14911) );
  OR2X1 U15338 ( .IN1(n14985), .IN2(n14986), .Q(g30505) );
  OR2X1 U15339 ( .IN1(n14987), .IN2(n14988), .Q(n14986) );
  AND2X1 U15340 ( .IN1(n3858), .IN2(n3765), .Q(n14988) );
  AND2X1 U15341 ( .IN1(n14989), .IN2(n14990), .Q(n14987) );
  INVX0 U15342 ( .INP(n3858), .ZN(n14990) );
  AND2X1 U15343 ( .IN1(n10810), .IN2(g5909), .Q(n14989) );
  AND2X1 U15344 ( .IN1(n10922), .IN2(g5913), .Q(n14985) );
  OR2X1 U15345 ( .IN1(n14991), .IN2(n14992), .Q(g30504) );
  OR2X1 U15346 ( .IN1(n14993), .IN2(n14994), .Q(n14992) );
  AND2X1 U15347 ( .IN1(n3861), .IN2(n3765), .Q(n14994) );
  AND2X1 U15348 ( .IN1(n14995), .IN2(n14996), .Q(n14993) );
  INVX0 U15349 ( .INP(n3861), .ZN(n14996) );
  AND2X1 U15350 ( .IN1(n10808), .IN2(g5901), .Q(n14995) );
  AND2X1 U15351 ( .IN1(n10922), .IN2(g5905), .Q(n14991) );
  OR2X1 U15352 ( .IN1(n14997), .IN2(n14998), .Q(g30503) );
  OR2X1 U15353 ( .IN1(n14999), .IN2(n15000), .Q(n14998) );
  AND2X1 U15354 ( .IN1(n3863), .IN2(n3765), .Q(n15000) );
  AND2X1 U15355 ( .IN1(n15001), .IN2(n15002), .Q(n14999) );
  INVX0 U15356 ( .INP(n3863), .ZN(n15002) );
  AND2X1 U15357 ( .IN1(n10811), .IN2(g5893), .Q(n15001) );
  AND2X1 U15358 ( .IN1(n10922), .IN2(g5897), .Q(n14997) );
  OR2X1 U15359 ( .IN1(n15003), .IN2(n15004), .Q(g30502) );
  OR2X1 U15360 ( .IN1(n15005), .IN2(n15006), .Q(n15004) );
  AND2X1 U15361 ( .IN1(n3865), .IN2(n3765), .Q(n15006) );
  AND2X1 U15362 ( .IN1(n15007), .IN2(n15008), .Q(n15005) );
  INVX0 U15363 ( .INP(n3865), .ZN(n15008) );
  AND2X1 U15364 ( .IN1(n10811), .IN2(g5889), .Q(n15007) );
  AND2X1 U15365 ( .IN1(test_so36), .IN2(n10896), .Q(n15003) );
  AND2X1 U15366 ( .IN1(n13925), .IN2(n5573), .Q(g30501) );
  AND2X1 U15367 ( .IN1(n5649), .IN2(n15009), .Q(n13925) );
  AND2X1 U15368 ( .IN1(n10811), .IN2(n13917), .Q(n15009) );
  OR2X1 U15369 ( .IN1(n14883), .IN2(n15010), .Q(n13917) );
  OR2X1 U15370 ( .IN1(n15011), .IN2(n15012), .Q(g30500) );
  OR2X1 U15371 ( .IN1(n15013), .IN2(n15014), .Q(n15012) );
  AND2X1 U15372 ( .IN1(n3765), .IN2(n13093), .Q(n15014) );
  AND2X1 U15373 ( .IN1(n15015), .IN2(g5619), .Q(n15013) );
  AND2X1 U15374 ( .IN1(n10922), .IN2(g5615), .Q(n15011) );
  OR2X1 U15375 ( .IN1(n15016), .IN2(n15017), .Q(g30499) );
  OR2X1 U15376 ( .IN1(n15018), .IN2(n15019), .Q(n15017) );
  AND2X1 U15377 ( .IN1(n10922), .IN2(g5611), .Q(n15019) );
  INVX0 U15378 ( .INP(n15020), .ZN(n15018) );
  OR2X1 U15379 ( .IN1(n15021), .IN2(n10876), .Q(n15020) );
  OR2X1 U15380 ( .IN1(n15022), .IN2(n10360), .Q(n15021) );
  AND2X1 U15381 ( .IN1(n15022), .IN2(n3765), .Q(n15016) );
  AND2X1 U15382 ( .IN1(g5523), .IN2(n13945), .Q(n15022) );
  OR2X1 U15383 ( .IN1(n15023), .IN2(n15024), .Q(g30498) );
  OR2X1 U15384 ( .IN1(n15025), .IN2(n15026), .Q(n15024) );
  AND2X1 U15385 ( .IN1(n10923), .IN2(g5607), .Q(n15026) );
  AND2X1 U15386 ( .IN1(n15027), .IN2(n10757), .Q(n15025) );
  AND2X1 U15387 ( .IN1(test_so6), .IN2(n15028), .Q(n15027) );
  INVX0 U15388 ( .INP(n13943), .ZN(n15028) );
  AND2X1 U15389 ( .IN1(n13943), .IN2(n3765), .Q(n15023) );
  AND2X1 U15390 ( .IN1(g5523), .IN2(n15029), .Q(n13943) );
  OR2X1 U15391 ( .IN1(n15030), .IN2(n15031), .Q(g30497) );
  OR2X1 U15392 ( .IN1(n15032), .IN2(n15033), .Q(n15031) );
  AND2X1 U15393 ( .IN1(n10923), .IN2(g5603), .Q(n15033) );
  INVX0 U15394 ( .INP(n15034), .ZN(n15032) );
  OR2X1 U15395 ( .IN1(n15035), .IN2(n10876), .Q(n15034) );
  OR2X1 U15396 ( .IN1(n15036), .IN2(n10310), .Q(n15035) );
  AND2X1 U15397 ( .IN1(n15036), .IN2(n3765), .Q(n15030) );
  AND2X1 U15398 ( .IN1(g5523), .IN2(n15037), .Q(n15036) );
  OR2X1 U15399 ( .IN1(n15038), .IN2(n15039), .Q(g30496) );
  OR2X1 U15400 ( .IN1(n15040), .IN2(n15041), .Q(n15039) );
  AND2X1 U15401 ( .IN1(n15042), .IN2(n10757), .Q(n15041) );
  AND2X1 U15402 ( .IN1(n15043), .IN2(g5615), .Q(n15042) );
  OR2X1 U15403 ( .IN1(n3877), .IN2(n3434), .Q(n15043) );
  AND2X1 U15404 ( .IN1(n10923), .IN2(g5599), .Q(n15040) );
  AND2X1 U15405 ( .IN1(n3875), .IN2(n15044), .Q(n15038) );
  OR2X1 U15406 ( .IN1(n15045), .IN2(n15046), .Q(g30495) );
  OR2X1 U15407 ( .IN1(n15047), .IN2(n15048), .Q(n15046) );
  AND2X1 U15408 ( .IN1(n15049), .IN2(n10757), .Q(n15048) );
  AND2X1 U15409 ( .IN1(n15050), .IN2(g5611), .Q(n15049) );
  OR2X1 U15410 ( .IN1(n3869), .IN2(n3434), .Q(n15050) );
  AND2X1 U15411 ( .IN1(n10923), .IN2(g5595), .Q(n15047) );
  AND2X1 U15412 ( .IN1(n3875), .IN2(n13945), .Q(n15045) );
  OR2X1 U15413 ( .IN1(n15051), .IN2(n15052), .Q(g30494) );
  OR2X1 U15414 ( .IN1(n15053), .IN2(n15054), .Q(n15052) );
  AND2X1 U15415 ( .IN1(n15055), .IN2(n10757), .Q(n15054) );
  AND2X1 U15416 ( .IN1(n15056), .IN2(g5607), .Q(n15055) );
  OR2X1 U15417 ( .IN1(n3871), .IN2(n3434), .Q(n15056) );
  AND2X1 U15418 ( .IN1(test_so5), .IN2(n10895), .Q(n15053) );
  AND2X1 U15419 ( .IN1(n3875), .IN2(n15029), .Q(n15051) );
  OR2X1 U15420 ( .IN1(n15057), .IN2(n15058), .Q(g30493) );
  OR2X1 U15421 ( .IN1(n15059), .IN2(n15060), .Q(n15058) );
  AND2X1 U15422 ( .IN1(n15061), .IN2(n10757), .Q(n15060) );
  AND2X1 U15423 ( .IN1(n15062), .IN2(g5603), .Q(n15061) );
  OR2X1 U15424 ( .IN1(n3874), .IN2(n3434), .Q(n15062) );
  INVX0 U15425 ( .INP(n13954), .ZN(n3434) );
  AND2X1 U15426 ( .IN1(g5517), .IN2(g5511), .Q(n13954) );
  AND2X1 U15427 ( .IN1(n10923), .IN2(g5587), .Q(n15059) );
  AND2X1 U15428 ( .IN1(n3875), .IN2(n15037), .Q(n15057) );
  OR2X1 U15429 ( .IN1(n15063), .IN2(n15064), .Q(g30492) );
  OR2X1 U15430 ( .IN1(n15065), .IN2(n15066), .Q(n15064) );
  AND2X1 U15431 ( .IN1(n15067), .IN2(n10757), .Q(n15066) );
  AND2X1 U15432 ( .IN1(n15068), .IN2(g5599), .Q(n15067) );
  OR2X1 U15433 ( .IN1(n3877), .IN2(n3436), .Q(n15068) );
  AND2X1 U15434 ( .IN1(n10923), .IN2(g5583), .Q(n15065) );
  AND2X1 U15435 ( .IN1(n3881), .IN2(n15044), .Q(n15063) );
  OR2X1 U15436 ( .IN1(n15069), .IN2(n15070), .Q(g30491) );
  OR2X1 U15437 ( .IN1(n15071), .IN2(n15072), .Q(n15070) );
  AND2X1 U15438 ( .IN1(n15073), .IN2(n10758), .Q(n15072) );
  AND2X1 U15439 ( .IN1(n15074), .IN2(g5595), .Q(n15073) );
  OR2X1 U15440 ( .IN1(n3869), .IN2(n3436), .Q(n15074) );
  AND2X1 U15441 ( .IN1(n10923), .IN2(g5579), .Q(n15071) );
  AND2X1 U15442 ( .IN1(n3881), .IN2(n13945), .Q(n15069) );
  OR2X1 U15443 ( .IN1(n15075), .IN2(n15076), .Q(g30490) );
  OR2X1 U15444 ( .IN1(n15077), .IN2(n15078), .Q(n15076) );
  AND2X1 U15445 ( .IN1(n15079), .IN2(n10758), .Q(n15078) );
  AND2X1 U15446 ( .IN1(test_so5), .IN2(n15080), .Q(n15079) );
  OR2X1 U15447 ( .IN1(n3871), .IN2(n3436), .Q(n15080) );
  AND2X1 U15448 ( .IN1(n10923), .IN2(g5575), .Q(n15077) );
  AND2X1 U15449 ( .IN1(n3881), .IN2(n15029), .Q(n15075) );
  OR2X1 U15450 ( .IN1(n15081), .IN2(n15082), .Q(g30489) );
  OR2X1 U15451 ( .IN1(n15083), .IN2(n15084), .Q(n15082) );
  AND2X1 U15452 ( .IN1(n15085), .IN2(n10758), .Q(n15084) );
  AND2X1 U15453 ( .IN1(n15086), .IN2(g5587), .Q(n15085) );
  OR2X1 U15454 ( .IN1(n3874), .IN2(n3436), .Q(n15086) );
  OR2X1 U15455 ( .IN1(n10426), .IN2(g5511), .Q(n3436) );
  AND2X1 U15456 ( .IN1(n10923), .IN2(g5571), .Q(n15083) );
  AND2X1 U15457 ( .IN1(n3881), .IN2(n15037), .Q(n15081) );
  OR2X1 U15458 ( .IN1(n15087), .IN2(n15088), .Q(g30488) );
  OR2X1 U15459 ( .IN1(n15089), .IN2(n15090), .Q(n15088) );
  AND2X1 U15460 ( .IN1(n15091), .IN2(n10758), .Q(n15090) );
  AND2X1 U15461 ( .IN1(n15092), .IN2(g5583), .Q(n15091) );
  OR2X1 U15462 ( .IN1(n3877), .IN2(n3437), .Q(n15092) );
  INVX0 U15463 ( .INP(n15044), .ZN(n3877) );
  AND2X1 U15464 ( .IN1(n10923), .IN2(g5563), .Q(n15089) );
  AND2X1 U15465 ( .IN1(n3886), .IN2(n15044), .Q(n15087) );
  OR2X1 U15466 ( .IN1(n15093), .IN2(n15094), .Q(g30487) );
  OR2X1 U15467 ( .IN1(n15095), .IN2(n15096), .Q(n15094) );
  AND2X1 U15468 ( .IN1(n15097), .IN2(n10758), .Q(n15096) );
  AND2X1 U15469 ( .IN1(n15098), .IN2(g5579), .Q(n15097) );
  OR2X1 U15470 ( .IN1(n3869), .IN2(n3437), .Q(n15098) );
  INVX0 U15471 ( .INP(n13945), .ZN(n3869) );
  AND2X1 U15472 ( .IN1(n10923), .IN2(g5555), .Q(n15095) );
  AND2X1 U15473 ( .IN1(n3886), .IN2(n13945), .Q(n15093) );
  AND2X1 U15474 ( .IN1(g5535), .IN2(n5389), .Q(n13945) );
  OR2X1 U15475 ( .IN1(n15099), .IN2(n15100), .Q(g30486) );
  OR2X1 U15476 ( .IN1(n15101), .IN2(n15102), .Q(n15100) );
  AND2X1 U15477 ( .IN1(n15103), .IN2(n10758), .Q(n15102) );
  AND2X1 U15478 ( .IN1(n15104), .IN2(g5575), .Q(n15103) );
  OR2X1 U15479 ( .IN1(n3871), .IN2(n3437), .Q(n15104) );
  INVX0 U15480 ( .INP(n15029), .ZN(n3871) );
  AND2X1 U15481 ( .IN1(n10923), .IN2(g5547), .Q(n15101) );
  AND2X1 U15482 ( .IN1(n3886), .IN2(n15029), .Q(n15099) );
  AND2X1 U15483 ( .IN1(g5527), .IN2(n5566), .Q(n15029) );
  OR2X1 U15484 ( .IN1(n15105), .IN2(n15106), .Q(g30485) );
  OR2X1 U15485 ( .IN1(n15107), .IN2(n15108), .Q(n15106) );
  AND2X1 U15486 ( .IN1(n15109), .IN2(n10758), .Q(n15108) );
  AND2X1 U15487 ( .IN1(n15110), .IN2(g5571), .Q(n15109) );
  OR2X1 U15488 ( .IN1(n3874), .IN2(n3437), .Q(n15110) );
  OR2X1 U15489 ( .IN1(n5575), .IN2(g5517), .Q(n3437) );
  INVX0 U15490 ( .INP(n15037), .ZN(n3874) );
  AND2X1 U15491 ( .IN1(n10923), .IN2(g5543), .Q(n15107) );
  AND2X1 U15492 ( .IN1(n3886), .IN2(n15037), .Q(n15105) );
  AND2X1 U15493 ( .IN1(n5389), .IN2(n5566), .Q(n15037) );
  OR2X1 U15494 ( .IN1(n15111), .IN2(n15112), .Q(g30484) );
  OR2X1 U15495 ( .IN1(n15113), .IN2(n15114), .Q(n15112) );
  AND2X1 U15496 ( .IN1(n3891), .IN2(n3765), .Q(n15114) );
  AND2X1 U15497 ( .IN1(n15115), .IN2(n15116), .Q(n15113) );
  INVX0 U15498 ( .INP(n3891), .ZN(n15116) );
  AND2X1 U15499 ( .IN1(n10811), .IN2(g5563), .Q(n15115) );
  AND2X1 U15500 ( .IN1(n10923), .IN2(g5567), .Q(n15111) );
  OR2X1 U15501 ( .IN1(n15117), .IN2(n15118), .Q(g30483) );
  OR2X1 U15502 ( .IN1(n15119), .IN2(n15120), .Q(n15118) );
  AND2X1 U15503 ( .IN1(n3894), .IN2(n3765), .Q(n15120) );
  AND2X1 U15504 ( .IN1(n15121), .IN2(n15122), .Q(n15119) );
  INVX0 U15505 ( .INP(n3894), .ZN(n15122) );
  AND2X1 U15506 ( .IN1(n10811), .IN2(g5555), .Q(n15121) );
  AND2X1 U15507 ( .IN1(test_so6), .IN2(n10895), .Q(n15117) );
  OR2X1 U15508 ( .IN1(n15123), .IN2(n15124), .Q(g30482) );
  OR2X1 U15509 ( .IN1(n15125), .IN2(n15126), .Q(n15124) );
  AND2X1 U15510 ( .IN1(n3896), .IN2(n3765), .Q(n15126) );
  AND2X1 U15511 ( .IN1(n15127), .IN2(n15128), .Q(n15125) );
  INVX0 U15512 ( .INP(n3896), .ZN(n15128) );
  AND2X1 U15513 ( .IN1(n10812), .IN2(g5547), .Q(n15127) );
  AND2X1 U15514 ( .IN1(n10923), .IN2(g5551), .Q(n15123) );
  OR2X1 U15515 ( .IN1(n15129), .IN2(n15130), .Q(g30481) );
  OR2X1 U15516 ( .IN1(n15131), .IN2(n15132), .Q(n15130) );
  AND2X1 U15517 ( .IN1(n3898), .IN2(n3765), .Q(n15132) );
  AND2X1 U15518 ( .IN1(n15133), .IN2(n15134), .Q(n15131) );
  INVX0 U15519 ( .INP(n3898), .ZN(n15134) );
  AND2X1 U15520 ( .IN1(n10812), .IN2(g5543), .Q(n15133) );
  AND2X1 U15521 ( .IN1(n10923), .IN2(g5535), .Q(n15129) );
  AND2X1 U15522 ( .IN1(n13948), .IN2(n5575), .Q(g30480) );
  AND2X1 U15523 ( .IN1(n5647), .IN2(n15135), .Q(n13948) );
  AND2X1 U15524 ( .IN1(n10812), .IN2(n13940), .Q(n15135) );
  OR2X1 U15525 ( .IN1(n15136), .IN2(n14883), .Q(n13940) );
  OR2X1 U15526 ( .IN1(n15137), .IN2(n15138), .Q(g30479) );
  OR2X1 U15527 ( .IN1(n15139), .IN2(n15140), .Q(n15138) );
  AND2X1 U15528 ( .IN1(n3765), .IN2(g32975), .Q(n15140) );
  AND2X1 U15529 ( .IN1(n15141), .IN2(g5272), .Q(n15139) );
  AND2X1 U15530 ( .IN1(n10923), .IN2(g5268), .Q(n15137) );
  OR2X1 U15531 ( .IN1(n15142), .IN2(n15143), .Q(g30478) );
  OR2X1 U15532 ( .IN1(n15144), .IN2(n15145), .Q(n15143) );
  AND2X1 U15533 ( .IN1(n10923), .IN2(g5264), .Q(n15145) );
  INVX0 U15534 ( .INP(n15146), .ZN(n15144) );
  OR2X1 U15535 ( .IN1(n15147), .IN2(n10874), .Q(n15146) );
  OR2X1 U15536 ( .IN1(n15148), .IN2(n10276), .Q(n15147) );
  AND2X1 U15537 ( .IN1(n15148), .IN2(n3765), .Q(n15142) );
  AND2X1 U15538 ( .IN1(g5176), .IN2(n13968), .Q(n15148) );
  OR2X1 U15539 ( .IN1(n15149), .IN2(n15150), .Q(g30477) );
  OR2X1 U15540 ( .IN1(n15151), .IN2(n15152), .Q(n15150) );
  AND2X1 U15541 ( .IN1(n10923), .IN2(g5260), .Q(n15152) );
  INVX0 U15542 ( .INP(n15153), .ZN(n15151) );
  OR2X1 U15543 ( .IN1(n15154), .IN2(n10874), .Q(n15153) );
  OR2X1 U15544 ( .IN1(n13966), .IN2(n10328), .Q(n15154) );
  AND2X1 U15545 ( .IN1(n13966), .IN2(n3765), .Q(n15149) );
  AND2X1 U15546 ( .IN1(g5176), .IN2(n15155), .Q(n13966) );
  OR2X1 U15547 ( .IN1(n15156), .IN2(n15157), .Q(g30476) );
  OR2X1 U15548 ( .IN1(n15158), .IN2(n15159), .Q(n15157) );
  AND2X1 U15549 ( .IN1(n10924), .IN2(g5256), .Q(n15159) );
  INVX0 U15550 ( .INP(n15160), .ZN(n15158) );
  OR2X1 U15551 ( .IN1(n15161), .IN2(n10875), .Q(n15160) );
  OR2X1 U15552 ( .IN1(n15162), .IN2(n10305), .Q(n15161) );
  AND2X1 U15553 ( .IN1(n15162), .IN2(n3765), .Q(n15156) );
  AND2X1 U15554 ( .IN1(g5176), .IN2(n15163), .Q(n15162) );
  OR2X1 U15555 ( .IN1(n15164), .IN2(n15165), .Q(g30475) );
  OR2X1 U15556 ( .IN1(n15166), .IN2(n15167), .Q(n15165) );
  AND2X1 U15557 ( .IN1(n15168), .IN2(n10758), .Q(n15167) );
  AND2X1 U15558 ( .IN1(n15169), .IN2(g5268), .Q(n15168) );
  OR2X1 U15559 ( .IN1(n3910), .IN2(n3444), .Q(n15169) );
  AND2X1 U15560 ( .IN1(n10924), .IN2(g5252), .Q(n15166) );
  AND2X1 U15561 ( .IN1(n3908), .IN2(n15170), .Q(n15164) );
  OR2X1 U15562 ( .IN1(n15171), .IN2(n15172), .Q(g30474) );
  OR2X1 U15563 ( .IN1(n15173), .IN2(n15174), .Q(n15172) );
  AND2X1 U15564 ( .IN1(n15175), .IN2(n10758), .Q(n15174) );
  AND2X1 U15565 ( .IN1(n15176), .IN2(g5264), .Q(n15175) );
  OR2X1 U15566 ( .IN1(n3902), .IN2(n3444), .Q(n15176) );
  AND2X1 U15567 ( .IN1(n10924), .IN2(g5248), .Q(n15173) );
  AND2X1 U15568 ( .IN1(n3908), .IN2(n13968), .Q(n15171) );
  OR2X1 U15569 ( .IN1(n15177), .IN2(n15178), .Q(g30473) );
  OR2X1 U15570 ( .IN1(n15179), .IN2(n15180), .Q(n15178) );
  AND2X1 U15571 ( .IN1(n15181), .IN2(n10759), .Q(n15180) );
  AND2X1 U15572 ( .IN1(n15182), .IN2(g5260), .Q(n15181) );
  OR2X1 U15573 ( .IN1(n3904), .IN2(n3444), .Q(n15182) );
  AND2X1 U15574 ( .IN1(n10924), .IN2(g5244), .Q(n15179) );
  AND2X1 U15575 ( .IN1(n3908), .IN2(n15155), .Q(n15177) );
  OR2X1 U15576 ( .IN1(n15183), .IN2(n15184), .Q(g30472) );
  OR2X1 U15577 ( .IN1(n15185), .IN2(n15186), .Q(n15184) );
  AND2X1 U15578 ( .IN1(n15187), .IN2(n10759), .Q(n15186) );
  AND2X1 U15579 ( .IN1(n15188), .IN2(g5256), .Q(n15187) );
  OR2X1 U15580 ( .IN1(n3907), .IN2(n3444), .Q(n15188) );
  INVX0 U15581 ( .INP(n13977), .ZN(n3444) );
  AND2X1 U15582 ( .IN1(g5170), .IN2(g5164), .Q(n13977) );
  AND2X1 U15583 ( .IN1(n10924), .IN2(g5240), .Q(n15185) );
  AND2X1 U15584 ( .IN1(n3908), .IN2(n15163), .Q(n15183) );
  OR2X1 U15585 ( .IN1(n15189), .IN2(n15190), .Q(g30471) );
  OR2X1 U15586 ( .IN1(n15191), .IN2(n15192), .Q(n15190) );
  AND2X1 U15587 ( .IN1(n15193), .IN2(n10759), .Q(n15192) );
  AND2X1 U15588 ( .IN1(n15194), .IN2(g5252), .Q(n15193) );
  OR2X1 U15589 ( .IN1(n3910), .IN2(n3446), .Q(n15194) );
  AND2X1 U15590 ( .IN1(n10924), .IN2(g5236), .Q(n15191) );
  AND2X1 U15591 ( .IN1(n3914), .IN2(n15170), .Q(n15189) );
  OR2X1 U15592 ( .IN1(n15195), .IN2(n15196), .Q(g30470) );
  OR2X1 U15593 ( .IN1(n15197), .IN2(n15198), .Q(n15196) );
  AND2X1 U15594 ( .IN1(n15199), .IN2(n10759), .Q(n15198) );
  AND2X1 U15595 ( .IN1(n15200), .IN2(g5248), .Q(n15199) );
  OR2X1 U15596 ( .IN1(n3902), .IN2(n3446), .Q(n15200) );
  AND2X1 U15597 ( .IN1(n10924), .IN2(g5232), .Q(n15197) );
  AND2X1 U15598 ( .IN1(n3914), .IN2(n13968), .Q(n15195) );
  OR2X1 U15599 ( .IN1(n15201), .IN2(n15202), .Q(g30469) );
  OR2X1 U15600 ( .IN1(n15203), .IN2(n15204), .Q(n15202) );
  AND2X1 U15601 ( .IN1(n15205), .IN2(n10759), .Q(n15204) );
  AND2X1 U15602 ( .IN1(n15206), .IN2(g5244), .Q(n15205) );
  OR2X1 U15603 ( .IN1(n3904), .IN2(n3446), .Q(n15206) );
  AND2X1 U15604 ( .IN1(test_so82), .IN2(n10895), .Q(n15203) );
  AND2X1 U15605 ( .IN1(n3914), .IN2(n15155), .Q(n15201) );
  OR2X1 U15606 ( .IN1(n15207), .IN2(n15208), .Q(g30468) );
  OR2X1 U15607 ( .IN1(n15209), .IN2(n15210), .Q(n15208) );
  AND2X1 U15608 ( .IN1(n15211), .IN2(n10759), .Q(n15210) );
  AND2X1 U15609 ( .IN1(n15212), .IN2(g5240), .Q(n15211) );
  OR2X1 U15610 ( .IN1(n3907), .IN2(n3446), .Q(n15212) );
  OR2X1 U15611 ( .IN1(n10429), .IN2(g5164), .Q(n3446) );
  AND2X1 U15612 ( .IN1(n10924), .IN2(g5224), .Q(n15209) );
  AND2X1 U15613 ( .IN1(n3914), .IN2(n15163), .Q(n15207) );
  OR2X1 U15614 ( .IN1(n15213), .IN2(n15214), .Q(g30467) );
  OR2X1 U15615 ( .IN1(n15215), .IN2(n15216), .Q(n15214) );
  AND2X1 U15616 ( .IN1(n15217), .IN2(n10759), .Q(n15216) );
  AND2X1 U15617 ( .IN1(n15218), .IN2(g5236), .Q(n15217) );
  OR2X1 U15618 ( .IN1(n3910), .IN2(n3447), .Q(n15218) );
  INVX0 U15619 ( .INP(n15170), .ZN(n3910) );
  AND2X1 U15620 ( .IN1(n10924), .IN2(g5216), .Q(n15215) );
  AND2X1 U15621 ( .IN1(n3919), .IN2(n15170), .Q(n15213) );
  OR2X1 U15622 ( .IN1(n15219), .IN2(n15220), .Q(g30466) );
  OR2X1 U15623 ( .IN1(n15221), .IN2(n15222), .Q(n15220) );
  AND2X1 U15624 ( .IN1(n15223), .IN2(n10759), .Q(n15222) );
  AND2X1 U15625 ( .IN1(n15224), .IN2(g5232), .Q(n15223) );
  OR2X1 U15626 ( .IN1(n3902), .IN2(n3447), .Q(n15224) );
  INVX0 U15627 ( .INP(n13968), .ZN(n3902) );
  AND2X1 U15628 ( .IN1(n10924), .IN2(g5208), .Q(n15221) );
  AND2X1 U15629 ( .IN1(n3919), .IN2(n13968), .Q(n15219) );
  AND2X1 U15630 ( .IN1(g5188), .IN2(n5384), .Q(n13968) );
  OR2X1 U15631 ( .IN1(n15225), .IN2(n15226), .Q(g30465) );
  OR2X1 U15632 ( .IN1(n15227), .IN2(n15228), .Q(n15226) );
  AND2X1 U15633 ( .IN1(n15229), .IN2(n10759), .Q(n15228) );
  AND2X1 U15634 ( .IN1(test_so82), .IN2(n15230), .Q(n15229) );
  OR2X1 U15635 ( .IN1(n3904), .IN2(n3447), .Q(n15230) );
  INVX0 U15636 ( .INP(n15155), .ZN(n3904) );
  AND2X1 U15637 ( .IN1(n10924), .IN2(g5200), .Q(n15227) );
  AND2X1 U15638 ( .IN1(n3919), .IN2(n15155), .Q(n15225) );
  AND2X1 U15639 ( .IN1(g5180), .IN2(n5567), .Q(n15155) );
  OR2X1 U15640 ( .IN1(n15231), .IN2(n15232), .Q(g30464) );
  OR2X1 U15641 ( .IN1(n15233), .IN2(n15234), .Q(n15232) );
  AND2X1 U15642 ( .IN1(n15235), .IN2(n10760), .Q(n15234) );
  AND2X1 U15643 ( .IN1(n15236), .IN2(g5224), .Q(n15235) );
  OR2X1 U15644 ( .IN1(n3907), .IN2(n3447), .Q(n15236) );
  OR2X1 U15645 ( .IN1(n5570), .IN2(g5170), .Q(n3447) );
  INVX0 U15646 ( .INP(n15163), .ZN(n3907) );
  AND2X1 U15647 ( .IN1(n10924), .IN2(g5196), .Q(n15233) );
  AND2X1 U15648 ( .IN1(n3919), .IN2(n15163), .Q(n15231) );
  AND2X1 U15649 ( .IN1(n5384), .IN2(n5567), .Q(n15163) );
  OR2X1 U15650 ( .IN1(n15237), .IN2(n15238), .Q(g30463) );
  OR2X1 U15651 ( .IN1(n15239), .IN2(n15240), .Q(n15238) );
  AND2X1 U15652 ( .IN1(n3924), .IN2(n3765), .Q(n15240) );
  AND2X1 U15653 ( .IN1(n15241), .IN2(n15242), .Q(n15239) );
  INVX0 U15654 ( .INP(n3924), .ZN(n15242) );
  AND2X1 U15655 ( .IN1(n10812), .IN2(g5216), .Q(n15241) );
  AND2X1 U15656 ( .IN1(n10924), .IN2(g5220), .Q(n15237) );
  OR2X1 U15657 ( .IN1(n15243), .IN2(n15244), .Q(g30462) );
  OR2X1 U15658 ( .IN1(n15245), .IN2(n15246), .Q(n15244) );
  AND2X1 U15659 ( .IN1(n3927), .IN2(n3765), .Q(n15246) );
  AND2X1 U15660 ( .IN1(n15247), .IN2(n15248), .Q(n15245) );
  INVX0 U15661 ( .INP(n3927), .ZN(n15248) );
  AND2X1 U15662 ( .IN1(n10812), .IN2(g5208), .Q(n15247) );
  AND2X1 U15663 ( .IN1(n10924), .IN2(g5212), .Q(n15243) );
  OR2X1 U15664 ( .IN1(n15249), .IN2(n15250), .Q(g30461) );
  OR2X1 U15665 ( .IN1(n15251), .IN2(n15252), .Q(n15250) );
  AND2X1 U15666 ( .IN1(n3929), .IN2(n3765), .Q(n15252) );
  AND2X1 U15667 ( .IN1(n15253), .IN2(n15254), .Q(n15251) );
  INVX0 U15668 ( .INP(n3929), .ZN(n15254) );
  AND2X1 U15669 ( .IN1(n10812), .IN2(g5200), .Q(n15253) );
  AND2X1 U15670 ( .IN1(n10924), .IN2(g5204), .Q(n15249) );
  OR2X1 U15671 ( .IN1(n15255), .IN2(n15256), .Q(g30460) );
  OR2X1 U15672 ( .IN1(n15257), .IN2(n15258), .Q(n15256) );
  AND2X1 U15673 ( .IN1(n3931), .IN2(n3765), .Q(n15258) );
  AND2X1 U15674 ( .IN1(n15259), .IN2(n15260), .Q(n15257) );
  INVX0 U15675 ( .INP(n3931), .ZN(n15260) );
  AND2X1 U15676 ( .IN1(n10812), .IN2(g5196), .Q(n15259) );
  AND2X1 U15677 ( .IN1(n10924), .IN2(g5188), .Q(n15255) );
  AND2X1 U15678 ( .IN1(n13971), .IN2(n5570), .Q(g30459) );
  AND2X1 U15679 ( .IN1(n5650), .IN2(n15261), .Q(n13971) );
  AND2X1 U15680 ( .IN1(n10812), .IN2(n13963), .Q(n15261) );
  OR2X1 U15681 ( .IN1(n14756), .IN2(n14883), .Q(n13963) );
  INVX0 U15682 ( .INP(n3833), .ZN(n14883) );
  OR2X1 U15683 ( .IN1(n10885), .IN2(n15262), .Q(g30458) );
  OR2X1 U15684 ( .IN1(n15263), .IN2(n15264), .Q(n15262) );
  INVX0 U15685 ( .INP(n15265), .ZN(n15264) );
  OR2X1 U15686 ( .IN1(n15266), .IN2(n5846), .Q(n15265) );
  AND2X1 U15687 ( .IN1(n15266), .IN2(g113), .Q(n15263) );
  AND2X1 U15688 ( .IN1(g4473), .IN2(n5765), .Q(n15266) );
  OR2X1 U15689 ( .IN1(n15267), .IN2(n15268), .Q(g30457) );
  AND2X1 U15690 ( .IN1(n15269), .IN2(n10760), .Q(n15268) );
  OR2X1 U15691 ( .IN1(n15270), .IN2(n15271), .Q(n15269) );
  AND2X1 U15692 ( .IN1(n15272), .IN2(n5983), .Q(n15271) );
  XNOR2X1 U15693 ( .IN1(g115), .IN2(n15273), .Q(n15272) );
  AND2X1 U15694 ( .IN1(n15274), .IN2(n5981), .Q(n15270) );
  XNOR2X1 U15695 ( .IN1(g126), .IN2(n15275), .Q(n15274) );
  AND2X1 U15696 ( .IN1(n10924), .IN2(g4122), .Q(n15267) );
  OR2X1 U15697 ( .IN1(n15276), .IN2(n15277), .Q(g30456) );
  OR2X1 U15698 ( .IN1(n15278), .IN2(n15279), .Q(n15277) );
  AND2X1 U15699 ( .IN1(n3941), .IN2(n15280), .Q(n15279) );
  AND2X1 U15700 ( .IN1(n15281), .IN2(n13081), .Q(n15278) );
  INVX0 U15701 ( .INP(n15136), .ZN(n13081) );
  INVX0 U15702 ( .INP(n15282), .ZN(n15281) );
  OR2X1 U15703 ( .IN1(n14545), .IN2(n5729), .Q(n15282) );
  AND2X1 U15704 ( .IN1(n10924), .IN2(g4087), .Q(n15276) );
  OR2X1 U15705 ( .IN1(n15283), .IN2(n15284), .Q(g30455) );
  OR2X1 U15706 ( .IN1(n15285), .IN2(n15286), .Q(n15284) );
  AND2X1 U15707 ( .IN1(n13080), .IN2(n3765), .Q(n15286) );
  AND2X1 U15708 ( .IN1(n15287), .IN2(g3965), .Q(n15285) );
  AND2X1 U15709 ( .IN1(n10925), .IN2(g3961), .Q(n15283) );
  OR2X1 U15710 ( .IN1(n15288), .IN2(n15289), .Q(g30454) );
  OR2X1 U15711 ( .IN1(n15290), .IN2(n15291), .Q(n15289) );
  AND2X1 U15712 ( .IN1(n10925), .IN2(g3957), .Q(n15291) );
  INVX0 U15713 ( .INP(n15292), .ZN(n15290) );
  OR2X1 U15714 ( .IN1(n15293), .IN2(n10874), .Q(n15292) );
  OR2X1 U15715 ( .IN1(n15294), .IN2(n10364), .Q(n15293) );
  AND2X1 U15716 ( .IN1(n15294), .IN2(n3765), .Q(n15288) );
  AND2X1 U15717 ( .IN1(n14040), .IN2(test_so33), .Q(n15294) );
  OR2X1 U15718 ( .IN1(n15295), .IN2(n15296), .Q(g30453) );
  OR2X1 U15719 ( .IN1(n15297), .IN2(n15298), .Q(n15296) );
  AND2X1 U15720 ( .IN1(n10925), .IN2(g3953), .Q(n15298) );
  INVX0 U15721 ( .INP(n15299), .ZN(n15297) );
  OR2X1 U15722 ( .IN1(n15300), .IN2(n10874), .Q(n15299) );
  OR2X1 U15723 ( .IN1(n14038), .IN2(n10339), .Q(n15300) );
  AND2X1 U15724 ( .IN1(n14038), .IN2(n3765), .Q(n15295) );
  AND2X1 U15725 ( .IN1(n15301), .IN2(test_so33), .Q(n14038) );
  OR2X1 U15726 ( .IN1(n15302), .IN2(n15303), .Q(g30452) );
  OR2X1 U15727 ( .IN1(n15304), .IN2(n15305), .Q(n15303) );
  AND2X1 U15728 ( .IN1(test_so65), .IN2(n10896), .Q(n15305) );
  INVX0 U15729 ( .INP(n15306), .ZN(n15304) );
  OR2X1 U15730 ( .IN1(n15307), .IN2(n10874), .Q(n15306) );
  OR2X1 U15731 ( .IN1(n15308), .IN2(n10312), .Q(n15307) );
  AND2X1 U15732 ( .IN1(n15308), .IN2(n3765), .Q(n15302) );
  AND2X1 U15733 ( .IN1(n15309), .IN2(test_so33), .Q(n15308) );
  OR2X1 U15734 ( .IN1(n15310), .IN2(n15311), .Q(g30451) );
  OR2X1 U15735 ( .IN1(n15312), .IN2(n15313), .Q(n15311) );
  AND2X1 U15736 ( .IN1(n15314), .IN2(n10760), .Q(n15313) );
  AND2X1 U15737 ( .IN1(n15315), .IN2(g3961), .Q(n15314) );
  OR2X1 U15738 ( .IN1(n3953), .IN2(n1075), .Q(n15315) );
  AND2X1 U15739 ( .IN1(n10925), .IN2(g3945), .Q(n15312) );
  AND2X1 U15740 ( .IN1(n3951), .IN2(n15316), .Q(n15310) );
  OR2X1 U15741 ( .IN1(n15317), .IN2(n15318), .Q(g30450) );
  OR2X1 U15742 ( .IN1(n15319), .IN2(n15320), .Q(n15318) );
  AND2X1 U15743 ( .IN1(n15321), .IN2(n10760), .Q(n15320) );
  AND2X1 U15744 ( .IN1(n15322), .IN2(g3957), .Q(n15321) );
  OR2X1 U15745 ( .IN1(n3945), .IN2(n1075), .Q(n15322) );
  AND2X1 U15746 ( .IN1(n10925), .IN2(g3941), .Q(n15319) );
  AND2X1 U15747 ( .IN1(n3951), .IN2(n14040), .Q(n15317) );
  OR2X1 U15748 ( .IN1(n15323), .IN2(n15324), .Q(g30449) );
  OR2X1 U15749 ( .IN1(n15325), .IN2(n15326), .Q(n15324) );
  AND2X1 U15750 ( .IN1(n15327), .IN2(n10760), .Q(n15326) );
  AND2X1 U15751 ( .IN1(n15328), .IN2(g3953), .Q(n15327) );
  OR2X1 U15752 ( .IN1(n3947), .IN2(n1075), .Q(n15328) );
  AND2X1 U15753 ( .IN1(n10925), .IN2(g3937), .Q(n15325) );
  AND2X1 U15754 ( .IN1(n3951), .IN2(n15301), .Q(n15323) );
  OR2X1 U15755 ( .IN1(n15329), .IN2(n15330), .Q(g30448) );
  OR2X1 U15756 ( .IN1(n15331), .IN2(n15332), .Q(n15330) );
  AND2X1 U15757 ( .IN1(n15333), .IN2(n10760), .Q(n15332) );
  AND2X1 U15758 ( .IN1(test_so65), .IN2(n15334), .Q(n15333) );
  OR2X1 U15759 ( .IN1(n3950), .IN2(n1075), .Q(n15334) );
  OR2X1 U15760 ( .IN1(n5572), .IN2(n10432), .Q(n1075) );
  AND2X1 U15761 ( .IN1(n10925), .IN2(g3933), .Q(n15331) );
  AND2X1 U15762 ( .IN1(n3951), .IN2(n15309), .Q(n15329) );
  OR2X1 U15763 ( .IN1(n15335), .IN2(n15336), .Q(g30447) );
  OR2X1 U15764 ( .IN1(n15337), .IN2(n15338), .Q(n15336) );
  AND2X1 U15765 ( .IN1(n15339), .IN2(n10760), .Q(n15338) );
  AND2X1 U15766 ( .IN1(n15340), .IN2(g3945), .Q(n15339) );
  OR2X1 U15767 ( .IN1(n3953), .IN2(n3481), .Q(n15340) );
  AND2X1 U15768 ( .IN1(n10925), .IN2(g3929), .Q(n15337) );
  AND2X1 U15769 ( .IN1(n3957), .IN2(n15316), .Q(n15335) );
  OR2X1 U15770 ( .IN1(n15341), .IN2(n15342), .Q(g30446) );
  OR2X1 U15771 ( .IN1(n15343), .IN2(n15344), .Q(n15342) );
  AND2X1 U15772 ( .IN1(n15345), .IN2(n10760), .Q(n15344) );
  AND2X1 U15773 ( .IN1(n15346), .IN2(g3941), .Q(n15345) );
  OR2X1 U15774 ( .IN1(n3945), .IN2(n3481), .Q(n15346) );
  AND2X1 U15775 ( .IN1(n10925), .IN2(g3925), .Q(n15343) );
  AND2X1 U15776 ( .IN1(n3957), .IN2(n14040), .Q(n15341) );
  OR2X1 U15777 ( .IN1(n15347), .IN2(n15348), .Q(g30445) );
  OR2X1 U15778 ( .IN1(n15349), .IN2(n15350), .Q(n15348) );
  AND2X1 U15779 ( .IN1(n15351), .IN2(n10760), .Q(n15350) );
  AND2X1 U15780 ( .IN1(n15352), .IN2(g3937), .Q(n15351) );
  OR2X1 U15781 ( .IN1(n3947), .IN2(n3481), .Q(n15352) );
  AND2X1 U15782 ( .IN1(n10925), .IN2(g3921), .Q(n15349) );
  AND2X1 U15783 ( .IN1(n3957), .IN2(n15301), .Q(n15347) );
  OR2X1 U15784 ( .IN1(n15353), .IN2(n15354), .Q(g30444) );
  OR2X1 U15785 ( .IN1(n15355), .IN2(n15356), .Q(n15354) );
  AND2X1 U15786 ( .IN1(n15357), .IN2(n10761), .Q(n15356) );
  AND2X1 U15787 ( .IN1(n15358), .IN2(g3933), .Q(n15357) );
  OR2X1 U15788 ( .IN1(n3950), .IN2(n3481), .Q(n15358) );
  OR2X1 U15789 ( .IN1(n10432), .IN2(g3857), .Q(n3481) );
  AND2X1 U15790 ( .IN1(n10925), .IN2(g3917), .Q(n15355) );
  AND2X1 U15791 ( .IN1(n3957), .IN2(n15309), .Q(n15353) );
  OR2X1 U15792 ( .IN1(n15359), .IN2(n15360), .Q(g30443) );
  OR2X1 U15793 ( .IN1(n15361), .IN2(n15362), .Q(n15360) );
  AND2X1 U15794 ( .IN1(n15363), .IN2(n10761), .Q(n15362) );
  AND2X1 U15795 ( .IN1(n15364), .IN2(g3929), .Q(n15363) );
  OR2X1 U15796 ( .IN1(n3953), .IN2(n3482), .Q(n15364) );
  INVX0 U15797 ( .INP(n15316), .ZN(n3953) );
  AND2X1 U15798 ( .IN1(n10925), .IN2(g3909), .Q(n15361) );
  AND2X1 U15799 ( .IN1(n3962), .IN2(n15316), .Q(n15359) );
  OR2X1 U15800 ( .IN1(n15365), .IN2(n15366), .Q(g30442) );
  OR2X1 U15801 ( .IN1(n15367), .IN2(n15368), .Q(n15366) );
  AND2X1 U15802 ( .IN1(n15369), .IN2(n10761), .Q(n15368) );
  AND2X1 U15803 ( .IN1(n15370), .IN2(g3925), .Q(n15369) );
  OR2X1 U15804 ( .IN1(n3945), .IN2(n3482), .Q(n15370) );
  INVX0 U15805 ( .INP(n14040), .ZN(n3945) );
  AND2X1 U15806 ( .IN1(n10925), .IN2(g3901), .Q(n15367) );
  AND2X1 U15807 ( .IN1(n3962), .IN2(n14040), .Q(n15365) );
  AND2X1 U15808 ( .IN1(g3881), .IN2(n5387), .Q(n14040) );
  OR2X1 U15809 ( .IN1(n15371), .IN2(n15372), .Q(g30441) );
  OR2X1 U15810 ( .IN1(n15373), .IN2(n15374), .Q(n15372) );
  AND2X1 U15811 ( .IN1(n15375), .IN2(n10761), .Q(n15374) );
  AND2X1 U15812 ( .IN1(n15376), .IN2(g3921), .Q(n15375) );
  OR2X1 U15813 ( .IN1(n3947), .IN2(n3482), .Q(n15376) );
  INVX0 U15814 ( .INP(n15301), .ZN(n3947) );
  AND2X1 U15815 ( .IN1(n10925), .IN2(g3893), .Q(n15373) );
  AND2X1 U15816 ( .IN1(n3962), .IN2(n15301), .Q(n15371) );
  AND2X1 U15817 ( .IN1(g3873), .IN2(n5564), .Q(n15301) );
  OR2X1 U15818 ( .IN1(n15377), .IN2(n15378), .Q(g30440) );
  OR2X1 U15819 ( .IN1(n15379), .IN2(n15380), .Q(n15378) );
  AND2X1 U15820 ( .IN1(n15381), .IN2(n10761), .Q(n15380) );
  AND2X1 U15821 ( .IN1(n15382), .IN2(g3917), .Q(n15381) );
  OR2X1 U15822 ( .IN1(n3950), .IN2(n3482), .Q(n15382) );
  OR2X1 U15823 ( .IN1(n5572), .IN2(g3863), .Q(n3482) );
  INVX0 U15824 ( .INP(n15309), .ZN(n3950) );
  AND2X1 U15825 ( .IN1(test_so24), .IN2(n10896), .Q(n15379) );
  AND2X1 U15826 ( .IN1(n3962), .IN2(n15309), .Q(n15377) );
  AND2X1 U15827 ( .IN1(n5387), .IN2(n5564), .Q(n15309) );
  OR2X1 U15828 ( .IN1(n15383), .IN2(n15384), .Q(g30439) );
  OR2X1 U15829 ( .IN1(n15385), .IN2(n15386), .Q(n15384) );
  AND2X1 U15830 ( .IN1(n3967), .IN2(n3765), .Q(n15386) );
  AND2X1 U15831 ( .IN1(n15387), .IN2(n15388), .Q(n15385) );
  INVX0 U15832 ( .INP(n3967), .ZN(n15388) );
  AND2X1 U15833 ( .IN1(n10814), .IN2(g3909), .Q(n15387) );
  AND2X1 U15834 ( .IN1(n10925), .IN2(g3913), .Q(n15383) );
  OR2X1 U15835 ( .IN1(n15389), .IN2(n15390), .Q(g30438) );
  OR2X1 U15836 ( .IN1(n15391), .IN2(n15392), .Q(n15390) );
  AND2X1 U15837 ( .IN1(n3970), .IN2(n3765), .Q(n15392) );
  AND2X1 U15838 ( .IN1(n15393), .IN2(n15394), .Q(n15391) );
  INVX0 U15839 ( .INP(n3970), .ZN(n15394) );
  AND2X1 U15840 ( .IN1(n10814), .IN2(g3901), .Q(n15393) );
  AND2X1 U15841 ( .IN1(n10925), .IN2(g3905), .Q(n15389) );
  OR2X1 U15842 ( .IN1(n15395), .IN2(n15396), .Q(g30437) );
  OR2X1 U15843 ( .IN1(n15397), .IN2(n15398), .Q(n15396) );
  AND2X1 U15844 ( .IN1(n3972), .IN2(n3765), .Q(n15398) );
  AND2X1 U15845 ( .IN1(n15399), .IN2(n15400), .Q(n15397) );
  INVX0 U15846 ( .INP(n3972), .ZN(n15400) );
  AND2X1 U15847 ( .IN1(n10814), .IN2(g3893), .Q(n15399) );
  AND2X1 U15848 ( .IN1(n10925), .IN2(g3897), .Q(n15395) );
  OR2X1 U15849 ( .IN1(n15401), .IN2(n15402), .Q(g30436) );
  OR2X1 U15850 ( .IN1(n15403), .IN2(n15404), .Q(n15402) );
  AND2X1 U15851 ( .IN1(n3974), .IN2(n3765), .Q(n15404) );
  AND2X1 U15852 ( .IN1(n15405), .IN2(n15406), .Q(n15403) );
  INVX0 U15853 ( .INP(n3974), .ZN(n15406) );
  AND2X1 U15854 ( .IN1(test_so24), .IN2(n10761), .Q(n15405) );
  AND2X1 U15855 ( .IN1(n10925), .IN2(g3881), .Q(n15401) );
  AND2X1 U15856 ( .IN1(n14043), .IN2(n5572), .Q(g30435) );
  AND2X1 U15857 ( .IN1(n14035), .IN2(n15407), .Q(n14043) );
  AND2X1 U15858 ( .IN1(n10553), .IN2(n10761), .Q(n15407) );
  OR2X1 U15859 ( .IN1(n14757), .IN2(n14884), .Q(n14035) );
  OR2X1 U15860 ( .IN1(n5480), .IN2(n5340), .Q(n14884) );
  OR2X1 U15861 ( .IN1(n15408), .IN2(n15409), .Q(g30434) );
  OR2X1 U15862 ( .IN1(n15410), .IN2(n15411), .Q(n15409) );
  AND2X1 U15863 ( .IN1(n13079), .IN2(n3765), .Q(n15411) );
  AND2X1 U15864 ( .IN1(n15412), .IN2(g3614), .Q(n15410) );
  AND2X1 U15865 ( .IN1(n10925), .IN2(g3610), .Q(n15408) );
  OR2X1 U15866 ( .IN1(n15413), .IN2(n15414), .Q(g30433) );
  OR2X1 U15867 ( .IN1(n15415), .IN2(n15416), .Q(n15414) );
  AND2X1 U15868 ( .IN1(n10926), .IN2(g3606), .Q(n15416) );
  INVX0 U15869 ( .INP(n15417), .ZN(n15415) );
  OR2X1 U15870 ( .IN1(n15418), .IN2(n10874), .Q(n15417) );
  OR2X1 U15871 ( .IN1(n15419), .IN2(n10372), .Q(n15418) );
  AND2X1 U15872 ( .IN1(n15419), .IN2(n3765), .Q(n15413) );
  AND2X1 U15873 ( .IN1(g3518), .IN2(n14063), .Q(n15419) );
  OR2X1 U15874 ( .IN1(n15420), .IN2(n15421), .Q(g30432) );
  OR2X1 U15875 ( .IN1(n15422), .IN2(n15423), .Q(n15421) );
  AND2X1 U15876 ( .IN1(test_so43), .IN2(n10897), .Q(n15423) );
  INVX0 U15877 ( .INP(n15424), .ZN(n15422) );
  OR2X1 U15878 ( .IN1(n15425), .IN2(n10874), .Q(n15424) );
  OR2X1 U15879 ( .IN1(n14061), .IN2(n10347), .Q(n15425) );
  AND2X1 U15880 ( .IN1(n14061), .IN2(n3765), .Q(n15420) );
  AND2X1 U15881 ( .IN1(g3518), .IN2(n15426), .Q(n14061) );
  OR2X1 U15882 ( .IN1(n15427), .IN2(n15428), .Q(g30431) );
  OR2X1 U15883 ( .IN1(n15429), .IN2(n15430), .Q(n15428) );
  AND2X1 U15884 ( .IN1(n10926), .IN2(g3598), .Q(n15430) );
  INVX0 U15885 ( .INP(n15431), .ZN(n15429) );
  OR2X1 U15886 ( .IN1(n15432), .IN2(n10874), .Q(n15431) );
  OR2X1 U15887 ( .IN1(n15433), .IN2(n10315), .Q(n15432) );
  AND2X1 U15888 ( .IN1(n15433), .IN2(n3765), .Q(n15427) );
  AND2X1 U15889 ( .IN1(g3518), .IN2(n15434), .Q(n15433) );
  OR2X1 U15890 ( .IN1(n15435), .IN2(n15436), .Q(g30430) );
  OR2X1 U15891 ( .IN1(n15437), .IN2(n15438), .Q(n15436) );
  AND2X1 U15892 ( .IN1(n15439), .IN2(n10761), .Q(n15438) );
  AND2X1 U15893 ( .IN1(n15440), .IN2(g3610), .Q(n15439) );
  OR2X1 U15894 ( .IN1(n3986), .IN2(n3489), .Q(n15440) );
  AND2X1 U15895 ( .IN1(n10926), .IN2(g3594), .Q(n15437) );
  AND2X1 U15896 ( .IN1(n3984), .IN2(n15441), .Q(n15435) );
  OR2X1 U15897 ( .IN1(n15442), .IN2(n15443), .Q(g30429) );
  OR2X1 U15898 ( .IN1(n15444), .IN2(n15445), .Q(n15443) );
  AND2X1 U15899 ( .IN1(n15446), .IN2(n10761), .Q(n15445) );
  AND2X1 U15900 ( .IN1(n15447), .IN2(g3606), .Q(n15446) );
  OR2X1 U15901 ( .IN1(n3978), .IN2(n3489), .Q(n15447) );
  AND2X1 U15902 ( .IN1(n10926), .IN2(g3590), .Q(n15444) );
  AND2X1 U15903 ( .IN1(n3984), .IN2(n14063), .Q(n15442) );
  OR2X1 U15904 ( .IN1(n15448), .IN2(n15449), .Q(g30428) );
  OR2X1 U15905 ( .IN1(n15450), .IN2(n15451), .Q(n15449) );
  AND2X1 U15906 ( .IN1(n15452), .IN2(n10762), .Q(n15451) );
  AND2X1 U15907 ( .IN1(test_so43), .IN2(n15453), .Q(n15452) );
  OR2X1 U15908 ( .IN1(n3980), .IN2(n3489), .Q(n15453) );
  AND2X1 U15909 ( .IN1(n10926), .IN2(g3586), .Q(n15450) );
  AND2X1 U15910 ( .IN1(n3984), .IN2(n15426), .Q(n15448) );
  OR2X1 U15911 ( .IN1(n15454), .IN2(n15455), .Q(g30427) );
  OR2X1 U15912 ( .IN1(n15456), .IN2(n15457), .Q(n15455) );
  AND2X1 U15913 ( .IN1(n15458), .IN2(n10762), .Q(n15457) );
  AND2X1 U15914 ( .IN1(n15459), .IN2(g3598), .Q(n15458) );
  OR2X1 U15915 ( .IN1(n3983), .IN2(n3489), .Q(n15459) );
  INVX0 U15916 ( .INP(n14072), .ZN(n3489) );
  AND2X1 U15917 ( .IN1(g3512), .IN2(g3506), .Q(n14072) );
  AND2X1 U15918 ( .IN1(n10926), .IN2(g3582), .Q(n15456) );
  AND2X1 U15919 ( .IN1(n3984), .IN2(n15434), .Q(n15454) );
  OR2X1 U15920 ( .IN1(n15460), .IN2(n15461), .Q(g30426) );
  OR2X1 U15921 ( .IN1(n15462), .IN2(n15463), .Q(n15461) );
  AND2X1 U15922 ( .IN1(n15464), .IN2(n10762), .Q(n15463) );
  AND2X1 U15923 ( .IN1(n15465), .IN2(g3594), .Q(n15464) );
  OR2X1 U15924 ( .IN1(n3986), .IN2(n3491), .Q(n15465) );
  AND2X1 U15925 ( .IN1(n10926), .IN2(g3578), .Q(n15462) );
  AND2X1 U15926 ( .IN1(n3990), .IN2(n15441), .Q(n15460) );
  OR2X1 U15927 ( .IN1(n15466), .IN2(n15467), .Q(g30425) );
  OR2X1 U15928 ( .IN1(n15468), .IN2(n15469), .Q(n15467) );
  AND2X1 U15929 ( .IN1(n15470), .IN2(n10762), .Q(n15469) );
  AND2X1 U15930 ( .IN1(n15471), .IN2(g3590), .Q(n15470) );
  OR2X1 U15931 ( .IN1(n3978), .IN2(n3491), .Q(n15471) );
  AND2X1 U15932 ( .IN1(n10926), .IN2(g3574), .Q(n15468) );
  AND2X1 U15933 ( .IN1(n3990), .IN2(n14063), .Q(n15466) );
  OR2X1 U15934 ( .IN1(n15472), .IN2(n15473), .Q(g30424) );
  OR2X1 U15935 ( .IN1(n15474), .IN2(n15475), .Q(n15473) );
  AND2X1 U15936 ( .IN1(n15476), .IN2(n10762), .Q(n15475) );
  AND2X1 U15937 ( .IN1(n15477), .IN2(g3586), .Q(n15476) );
  OR2X1 U15938 ( .IN1(n3980), .IN2(n3491), .Q(n15477) );
  AND2X1 U15939 ( .IN1(n10926), .IN2(g3570), .Q(n15474) );
  AND2X1 U15940 ( .IN1(n3990), .IN2(n15426), .Q(n15472) );
  OR2X1 U15941 ( .IN1(n15478), .IN2(n15479), .Q(g30423) );
  OR2X1 U15942 ( .IN1(n15480), .IN2(n15481), .Q(n15479) );
  AND2X1 U15943 ( .IN1(n15482), .IN2(n10762), .Q(n15481) );
  AND2X1 U15944 ( .IN1(n15483), .IN2(g3582), .Q(n15482) );
  OR2X1 U15945 ( .IN1(n3983), .IN2(n3491), .Q(n15483) );
  OR2X1 U15946 ( .IN1(n10427), .IN2(g3506), .Q(n3491) );
  AND2X1 U15947 ( .IN1(n10926), .IN2(g3566), .Q(n15480) );
  AND2X1 U15948 ( .IN1(n3990), .IN2(n15434), .Q(n15478) );
  OR2X1 U15949 ( .IN1(n15484), .IN2(n15485), .Q(g30422) );
  OR2X1 U15950 ( .IN1(n15486), .IN2(n15487), .Q(n15485) );
  AND2X1 U15951 ( .IN1(n15488), .IN2(n10762), .Q(n15487) );
  AND2X1 U15952 ( .IN1(n15489), .IN2(g3578), .Q(n15488) );
  OR2X1 U15953 ( .IN1(n3986), .IN2(n3492), .Q(n15489) );
  INVX0 U15954 ( .INP(n15441), .ZN(n3986) );
  AND2X1 U15955 ( .IN1(n10926), .IN2(g3558), .Q(n15486) );
  AND2X1 U15956 ( .IN1(n3995), .IN2(n15441), .Q(n15484) );
  OR2X1 U15957 ( .IN1(n15490), .IN2(n15491), .Q(g30421) );
  OR2X1 U15958 ( .IN1(n15492), .IN2(n15493), .Q(n15491) );
  AND2X1 U15959 ( .IN1(n15494), .IN2(n10762), .Q(n15493) );
  AND2X1 U15960 ( .IN1(n15495), .IN2(g3574), .Q(n15494) );
  OR2X1 U15961 ( .IN1(n3978), .IN2(n3492), .Q(n15495) );
  INVX0 U15962 ( .INP(n14063), .ZN(n3978) );
  AND2X1 U15963 ( .IN1(n10926), .IN2(g3550), .Q(n15492) );
  AND2X1 U15964 ( .IN1(n3995), .IN2(n14063), .Q(n15490) );
  AND2X1 U15965 ( .IN1(g3530), .IN2(n5383), .Q(n14063) );
  OR2X1 U15966 ( .IN1(n15496), .IN2(n15497), .Q(g30420) );
  OR2X1 U15967 ( .IN1(n15498), .IN2(n15499), .Q(n15497) );
  AND2X1 U15968 ( .IN1(n15500), .IN2(n10762), .Q(n15499) );
  AND2X1 U15969 ( .IN1(n15501), .IN2(g3570), .Q(n15500) );
  OR2X1 U15970 ( .IN1(n3980), .IN2(n3492), .Q(n15501) );
  INVX0 U15971 ( .INP(n15426), .ZN(n3980) );
  AND2X1 U15972 ( .IN1(n10926), .IN2(g3542), .Q(n15498) );
  AND2X1 U15973 ( .IN1(n3995), .IN2(n15426), .Q(n15496) );
  AND2X1 U15974 ( .IN1(g3522), .IN2(n5569), .Q(n15426) );
  OR2X1 U15975 ( .IN1(n15502), .IN2(n15503), .Q(g30419) );
  OR2X1 U15976 ( .IN1(n15504), .IN2(n15505), .Q(n15503) );
  AND2X1 U15977 ( .IN1(n15506), .IN2(n10802), .Q(n15505) );
  AND2X1 U15978 ( .IN1(n15507), .IN2(g3566), .Q(n15506) );
  OR2X1 U15979 ( .IN1(n3983), .IN2(n3492), .Q(n15507) );
  OR2X1 U15980 ( .IN1(n5576), .IN2(g3512), .Q(n3492) );
  INVX0 U15981 ( .INP(n15434), .ZN(n3983) );
  AND2X1 U15982 ( .IN1(n10926), .IN2(g3538), .Q(n15504) );
  AND2X1 U15983 ( .IN1(n3995), .IN2(n15434), .Q(n15502) );
  AND2X1 U15984 ( .IN1(n5383), .IN2(n5569), .Q(n15434) );
  OR2X1 U15985 ( .IN1(n15508), .IN2(n15509), .Q(g30418) );
  OR2X1 U15986 ( .IN1(n15510), .IN2(n15511), .Q(n15509) );
  AND2X1 U15987 ( .IN1(n4000), .IN2(n3765), .Q(n15511) );
  AND2X1 U15988 ( .IN1(n15512), .IN2(n15513), .Q(n15510) );
  INVX0 U15989 ( .INP(n4000), .ZN(n15513) );
  AND2X1 U15990 ( .IN1(n10815), .IN2(g3558), .Q(n15512) );
  AND2X1 U15991 ( .IN1(n10926), .IN2(g3562), .Q(n15508) );
  OR2X1 U15992 ( .IN1(n15514), .IN2(n15515), .Q(g30417) );
  OR2X1 U15993 ( .IN1(n15516), .IN2(n15517), .Q(n15515) );
  AND2X1 U15994 ( .IN1(n4003), .IN2(n3765), .Q(n15517) );
  AND2X1 U15995 ( .IN1(n15518), .IN2(n15519), .Q(n15516) );
  INVX0 U15996 ( .INP(n4003), .ZN(n15519) );
  AND2X1 U15997 ( .IN1(n10815), .IN2(g3550), .Q(n15518) );
  AND2X1 U15998 ( .IN1(n10926), .IN2(g3554), .Q(n15514) );
  OR2X1 U15999 ( .IN1(n15520), .IN2(n15521), .Q(g30416) );
  OR2X1 U16000 ( .IN1(n15522), .IN2(n15523), .Q(n15521) );
  AND2X1 U16001 ( .IN1(n4005), .IN2(n3765), .Q(n15523) );
  AND2X1 U16002 ( .IN1(n15524), .IN2(n15525), .Q(n15522) );
  INVX0 U16003 ( .INP(n4005), .ZN(n15525) );
  AND2X1 U16004 ( .IN1(n10815), .IN2(g3542), .Q(n15524) );
  AND2X1 U16005 ( .IN1(n10926), .IN2(g3546), .Q(n15520) );
  OR2X1 U16006 ( .IN1(n15526), .IN2(n15527), .Q(g30415) );
  OR2X1 U16007 ( .IN1(n15528), .IN2(n15529), .Q(n15527) );
  AND2X1 U16008 ( .IN1(n4007), .IN2(n3765), .Q(n15529) );
  AND2X1 U16009 ( .IN1(n15530), .IN2(n15531), .Q(n15528) );
  INVX0 U16010 ( .INP(n4007), .ZN(n15531) );
  AND2X1 U16011 ( .IN1(n10814), .IN2(g3538), .Q(n15530) );
  AND2X1 U16012 ( .IN1(n10926), .IN2(g3530), .Q(n15526) );
  AND2X1 U16013 ( .IN1(n14066), .IN2(n5576), .Q(g30414) );
  AND2X1 U16014 ( .IN1(n5645), .IN2(n15532), .Q(n14066) );
  AND2X1 U16015 ( .IN1(n10814), .IN2(n14058), .Q(n15532) );
  OR2X1 U16016 ( .IN1(n14757), .IN2(n15010), .Q(n14058) );
  OR2X1 U16017 ( .IN1(n5340), .IN2(g4087), .Q(n15010) );
  OR2X1 U16018 ( .IN1(n15533), .IN2(n15534), .Q(g30413) );
  OR2X1 U16019 ( .IN1(n15535), .IN2(n15536), .Q(n15534) );
  AND2X1 U16020 ( .IN1(n3765), .IN2(n13082), .Q(n15536) );
  AND2X1 U16021 ( .IN1(n15537), .IN2(g3263), .Q(n15535) );
  AND2X1 U16022 ( .IN1(test_so84), .IN2(n10896), .Q(n15533) );
  OR2X1 U16023 ( .IN1(n15538), .IN2(n15539), .Q(g30412) );
  OR2X1 U16024 ( .IN1(n15540), .IN2(n15541), .Q(n15539) );
  AND2X1 U16025 ( .IN1(n10926), .IN2(g3255), .Q(n15541) );
  INVX0 U16026 ( .INP(n15542), .ZN(n15540) );
  OR2X1 U16027 ( .IN1(n15543), .IN2(n10874), .Q(n15542) );
  OR2X1 U16028 ( .IN1(n15544), .IN2(n10352), .Q(n15543) );
  AND2X1 U16029 ( .IN1(n15544), .IN2(n3765), .Q(n15538) );
  AND2X1 U16030 ( .IN1(g3167), .IN2(n14086), .Q(n15544) );
  OR2X1 U16031 ( .IN1(n15545), .IN2(n15546), .Q(g30411) );
  OR2X1 U16032 ( .IN1(n15547), .IN2(n15548), .Q(n15546) );
  AND2X1 U16033 ( .IN1(n10927), .IN2(g3251), .Q(n15548) );
  INVX0 U16034 ( .INP(n15549), .ZN(n15547) );
  OR2X1 U16035 ( .IN1(n15550), .IN2(n10874), .Q(n15549) );
  OR2X1 U16036 ( .IN1(n14085), .IN2(n10324), .Q(n15550) );
  AND2X1 U16037 ( .IN1(n14085), .IN2(n3765), .Q(n15545) );
  AND2X1 U16038 ( .IN1(g3167), .IN2(n15551), .Q(n14085) );
  OR2X1 U16039 ( .IN1(n15552), .IN2(n15553), .Q(g30410) );
  OR2X1 U16040 ( .IN1(n15554), .IN2(n15555), .Q(n15553) );
  AND2X1 U16041 ( .IN1(n10897), .IN2(g3247), .Q(n15555) );
  AND2X1 U16042 ( .IN1(n15556), .IN2(n10807), .Q(n15554) );
  AND2X1 U16043 ( .IN1(test_so88), .IN2(n15557), .Q(n15556) );
  INVX0 U16044 ( .INP(n15558), .ZN(n15557) );
  AND2X1 U16045 ( .IN1(n15558), .IN2(n3765), .Q(n15552) );
  AND2X1 U16046 ( .IN1(g3167), .IN2(n15559), .Q(n15558) );
  OR2X1 U16047 ( .IN1(n15560), .IN2(n15561), .Q(g30409) );
  OR2X1 U16048 ( .IN1(n15562), .IN2(n15563), .Q(n15561) );
  AND2X1 U16049 ( .IN1(n15564), .IN2(n10806), .Q(n15563) );
  AND2X1 U16050 ( .IN1(test_so84), .IN2(n15565), .Q(n15564) );
  OR2X1 U16051 ( .IN1(n4017), .IN2(n3500), .Q(n15565) );
  AND2X1 U16052 ( .IN1(n10897), .IN2(g3243), .Q(n15562) );
  AND2X1 U16053 ( .IN1(n4015), .IN2(n15566), .Q(n15560) );
  OR2X1 U16054 ( .IN1(n15567), .IN2(n15568), .Q(g30408) );
  OR2X1 U16055 ( .IN1(n15569), .IN2(n15570), .Q(n15568) );
  AND2X1 U16056 ( .IN1(n15571), .IN2(n10807), .Q(n15570) );
  AND2X1 U16057 ( .IN1(n15572), .IN2(g3255), .Q(n15571) );
  OR2X1 U16058 ( .IN1(n3500), .IN2(n3495), .Q(n15572) );
  AND2X1 U16059 ( .IN1(n10897), .IN2(g3239), .Q(n15569) );
  AND2X1 U16060 ( .IN1(n4015), .IN2(n14086), .Q(n15567) );
  OR2X1 U16061 ( .IN1(n15573), .IN2(n15574), .Q(g30407) );
  OR2X1 U16062 ( .IN1(n15575), .IN2(n15576), .Q(n15574) );
  AND2X1 U16063 ( .IN1(n15577), .IN2(n10806), .Q(n15576) );
  AND2X1 U16064 ( .IN1(n15578), .IN2(g3251), .Q(n15577) );
  OR2X1 U16065 ( .IN1(n4020), .IN2(n3500), .Q(n15578) );
  AND2X1 U16066 ( .IN1(n10898), .IN2(g3235), .Q(n15575) );
  AND2X1 U16067 ( .IN1(n4015), .IN2(n15551), .Q(n15573) );
  OR2X1 U16068 ( .IN1(n15579), .IN2(n15580), .Q(g30406) );
  OR2X1 U16069 ( .IN1(n15581), .IN2(n15582), .Q(n15580) );
  AND2X1 U16070 ( .IN1(n15583), .IN2(n10807), .Q(n15582) );
  AND2X1 U16071 ( .IN1(n15584), .IN2(g3247), .Q(n15583) );
  OR2X1 U16072 ( .IN1(n4014), .IN2(n3500), .Q(n15584) );
  INVX0 U16073 ( .INP(n14095), .ZN(n3500) );
  AND2X1 U16074 ( .IN1(g3161), .IN2(g3155), .Q(n14095) );
  AND2X1 U16075 ( .IN1(n10897), .IN2(g3231), .Q(n15581) );
  AND2X1 U16076 ( .IN1(n4015), .IN2(n15559), .Q(n15579) );
  OR2X1 U16077 ( .IN1(n15585), .IN2(n15586), .Q(g30405) );
  OR2X1 U16078 ( .IN1(n15587), .IN2(n15588), .Q(n15586) );
  AND2X1 U16079 ( .IN1(n15589), .IN2(n10805), .Q(n15588) );
  AND2X1 U16080 ( .IN1(n15590), .IN2(g3243), .Q(n15589) );
  OR2X1 U16081 ( .IN1(n4017), .IN2(n3502), .Q(n15590) );
  AND2X1 U16082 ( .IN1(n10897), .IN2(g3227), .Q(n15587) );
  AND2X1 U16083 ( .IN1(n4022), .IN2(n15566), .Q(n15585) );
  OR2X1 U16084 ( .IN1(n15591), .IN2(n15592), .Q(g30404) );
  OR2X1 U16085 ( .IN1(n15593), .IN2(n15594), .Q(n15592) );
  AND2X1 U16086 ( .IN1(n15595), .IN2(n10804), .Q(n15594) );
  AND2X1 U16087 ( .IN1(n15596), .IN2(g3239), .Q(n15595) );
  OR2X1 U16088 ( .IN1(n3502), .IN2(n3495), .Q(n15596) );
  AND2X1 U16089 ( .IN1(n10898), .IN2(g3223), .Q(n15593) );
  AND2X1 U16090 ( .IN1(n4022), .IN2(n14086), .Q(n15591) );
  OR2X1 U16091 ( .IN1(n15597), .IN2(n15598), .Q(g30403) );
  OR2X1 U16092 ( .IN1(n15599), .IN2(n15600), .Q(n15598) );
  AND2X1 U16093 ( .IN1(n15601), .IN2(n10806), .Q(n15600) );
  AND2X1 U16094 ( .IN1(n15602), .IN2(g3235), .Q(n15601) );
  OR2X1 U16095 ( .IN1(n4020), .IN2(n3502), .Q(n15602) );
  AND2X1 U16096 ( .IN1(n10897), .IN2(g3219), .Q(n15599) );
  AND2X1 U16097 ( .IN1(n4022), .IN2(n15551), .Q(n15597) );
  OR2X1 U16098 ( .IN1(n15603), .IN2(n15604), .Q(g30402) );
  OR2X1 U16099 ( .IN1(n15605), .IN2(n15606), .Q(n15604) );
  AND2X1 U16100 ( .IN1(n15607), .IN2(n10805), .Q(n15606) );
  AND2X1 U16101 ( .IN1(n15608), .IN2(g3231), .Q(n15607) );
  OR2X1 U16102 ( .IN1(n4014), .IN2(n3502), .Q(n15608) );
  OR2X1 U16103 ( .IN1(n10425), .IN2(g3155), .Q(n3502) );
  AND2X1 U16104 ( .IN1(n10898), .IN2(g3215), .Q(n15605) );
  AND2X1 U16105 ( .IN1(n4022), .IN2(n15559), .Q(n15603) );
  OR2X1 U16106 ( .IN1(n15609), .IN2(n15610), .Q(g30401) );
  OR2X1 U16107 ( .IN1(n15611), .IN2(n15612), .Q(n15610) );
  AND2X1 U16108 ( .IN1(n15613), .IN2(n10805), .Q(n15612) );
  AND2X1 U16109 ( .IN1(n15614), .IN2(g3227), .Q(n15613) );
  OR2X1 U16110 ( .IN1(n4017), .IN2(n3501), .Q(n15614) );
  INVX0 U16111 ( .INP(n15566), .ZN(n4017) );
  AND2X1 U16112 ( .IN1(n10898), .IN2(g3207), .Q(n15611) );
  AND2X1 U16113 ( .IN1(n4027), .IN2(n15566), .Q(n15609) );
  OR2X1 U16114 ( .IN1(n15615), .IN2(n15616), .Q(g30400) );
  OR2X1 U16115 ( .IN1(n15617), .IN2(n15618), .Q(n15616) );
  AND2X1 U16116 ( .IN1(n15619), .IN2(n10804), .Q(n15618) );
  AND2X1 U16117 ( .IN1(n15620), .IN2(g3223), .Q(n15619) );
  OR2X1 U16118 ( .IN1(n3501), .IN2(n3495), .Q(n15620) );
  INVX0 U16119 ( .INP(n14086), .ZN(n3495) );
  AND2X1 U16120 ( .IN1(n10898), .IN2(g3199), .Q(n15617) );
  AND2X1 U16121 ( .IN1(n4027), .IN2(n14086), .Q(n15615) );
  AND2X1 U16122 ( .IN1(g3179), .IN2(n5603), .Q(n14086) );
  OR2X1 U16123 ( .IN1(n15621), .IN2(n15622), .Q(g30399) );
  OR2X1 U16124 ( .IN1(n15623), .IN2(n15624), .Q(n15622) );
  AND2X1 U16125 ( .IN1(n15625), .IN2(n10805), .Q(n15624) );
  AND2X1 U16126 ( .IN1(n15626), .IN2(g3219), .Q(n15625) );
  OR2X1 U16127 ( .IN1(n4020), .IN2(n3501), .Q(n15626) );
  INVX0 U16128 ( .INP(n15551), .ZN(n4020) );
  AND2X1 U16129 ( .IN1(n10899), .IN2(g3191), .Q(n15623) );
  AND2X1 U16130 ( .IN1(n4027), .IN2(n15551), .Q(n15621) );
  AND2X1 U16131 ( .IN1(g3171), .IN2(n5390), .Q(n15551) );
  OR2X1 U16132 ( .IN1(n15627), .IN2(n15628), .Q(g30398) );
  OR2X1 U16133 ( .IN1(n15629), .IN2(n15630), .Q(n15628) );
  AND2X1 U16134 ( .IN1(n15631), .IN2(n10805), .Q(n15630) );
  AND2X1 U16135 ( .IN1(n15632), .IN2(g3215), .Q(n15631) );
  OR2X1 U16136 ( .IN1(n4014), .IN2(n3501), .Q(n15632) );
  OR2X1 U16137 ( .IN1(n5366), .IN2(g3161), .Q(n3501) );
  INVX0 U16138 ( .INP(n15559), .ZN(n4014) );
  AND2X1 U16139 ( .IN1(n10899), .IN2(g3187), .Q(n15629) );
  AND2X1 U16140 ( .IN1(n4027), .IN2(n15559), .Q(n15627) );
  AND2X1 U16141 ( .IN1(n5390), .IN2(n5603), .Q(n15559) );
  OR2X1 U16142 ( .IN1(n15633), .IN2(n15634), .Q(g30397) );
  OR2X1 U16143 ( .IN1(n15635), .IN2(n15636), .Q(n15634) );
  AND2X1 U16144 ( .IN1(n4032), .IN2(n3765), .Q(n15636) );
  AND2X1 U16145 ( .IN1(n15637), .IN2(n15638), .Q(n15635) );
  INVX0 U16146 ( .INP(n4032), .ZN(n15638) );
  AND2X1 U16147 ( .IN1(n10813), .IN2(g3207), .Q(n15637) );
  AND2X1 U16148 ( .IN1(n10899), .IN2(g3211), .Q(n15633) );
  OR2X1 U16149 ( .IN1(n15639), .IN2(n15640), .Q(g30396) );
  OR2X1 U16150 ( .IN1(n15641), .IN2(n15642), .Q(n15640) );
  AND2X1 U16151 ( .IN1(n4035), .IN2(n3765), .Q(n15642) );
  AND2X1 U16152 ( .IN1(n15643), .IN2(n15644), .Q(n15641) );
  INVX0 U16153 ( .INP(n4035), .ZN(n15644) );
  AND2X1 U16154 ( .IN1(n10813), .IN2(g3199), .Q(n15643) );
  AND2X1 U16155 ( .IN1(n10899), .IN2(g3203), .Q(n15639) );
  OR2X1 U16156 ( .IN1(n15645), .IN2(n15646), .Q(g30395) );
  OR2X1 U16157 ( .IN1(n15647), .IN2(n15648), .Q(n15646) );
  AND2X1 U16158 ( .IN1(n4037), .IN2(n3765), .Q(n15648) );
  AND2X1 U16159 ( .IN1(n15649), .IN2(n15650), .Q(n15647) );
  INVX0 U16160 ( .INP(n4037), .ZN(n15650) );
  AND2X1 U16161 ( .IN1(n10813), .IN2(g3191), .Q(n15649) );
  AND2X1 U16162 ( .IN1(test_so88), .IN2(n10896), .Q(n15645) );
  OR2X1 U16163 ( .IN1(n15651), .IN2(n15652), .Q(g30394) );
  OR2X1 U16164 ( .IN1(n15653), .IN2(n15654), .Q(n15652) );
  AND2X1 U16165 ( .IN1(n4039), .IN2(n3765), .Q(n15654) );
  AND2X1 U16166 ( .IN1(n15655), .IN2(n15656), .Q(n15653) );
  INVX0 U16167 ( .INP(n4039), .ZN(n15656) );
  AND2X1 U16168 ( .IN1(n10813), .IN2(g3187), .Q(n15655) );
  AND2X1 U16169 ( .IN1(n10899), .IN2(g3179), .Q(n15651) );
  AND2X1 U16170 ( .IN1(n15657), .IN2(n14087), .Q(g30393) );
  AND2X1 U16171 ( .IN1(n14084), .IN2(n5652), .Q(n14087) );
  OR2X1 U16172 ( .IN1(n15136), .IN2(n14757), .Q(n14084) );
  INVX0 U16173 ( .INP(n3799), .ZN(n14757) );
  AND2X1 U16174 ( .IN1(n5366), .IN2(n10804), .Q(n15657) );
  OR2X1 U16175 ( .IN1(n15658), .IN2(n15659), .Q(g30392) );
  AND2X1 U16176 ( .IN1(n10899), .IN2(g2803), .Q(n15658) );
  OR2X1 U16177 ( .IN1(n15660), .IN2(n15661), .Q(g30391) );
  AND2X1 U16178 ( .IN1(n10900), .IN2(g2771), .Q(n15660) );
  OR2X1 U16179 ( .IN1(n15662), .IN2(n15659), .Q(g30390) );
  AND2X1 U16180 ( .IN1(n10813), .IN2(n15663), .Q(n15659) );
  INVX0 U16181 ( .INP(n15664), .ZN(n15663) );
  OR2X1 U16182 ( .IN1(n15665), .IN2(n15666), .Q(n15664) );
  AND2X1 U16183 ( .IN1(n15667), .IN2(n15668), .Q(n15666) );
  OR2X1 U16184 ( .IN1(n15669), .IN2(n15670), .Q(n15668) );
  OR2X1 U16185 ( .IN1(n15671), .IN2(n15672), .Q(n15670) );
  AND2X1 U16186 ( .IN1(n15673), .IN2(g2807), .Q(n15672) );
  AND2X1 U16187 ( .IN1(n15674), .IN2(g2803), .Q(n15671) );
  OR2X1 U16188 ( .IN1(n15675), .IN2(n15676), .Q(n15669) );
  AND2X1 U16189 ( .IN1(n15677), .IN2(g2819), .Q(n15676) );
  AND2X1 U16190 ( .IN1(n15678), .IN2(g2815), .Q(n15675) );
  AND2X1 U16191 ( .IN1(n15679), .IN2(n15680), .Q(n15665) );
  OR2X1 U16192 ( .IN1(n15681), .IN2(n15682), .Q(n15679) );
  OR2X1 U16193 ( .IN1(n15683), .IN2(n15684), .Q(n15682) );
  AND2X1 U16194 ( .IN1(n10302), .IN2(n15678), .Q(n15684) );
  AND2X1 U16195 ( .IN1(n10195), .IN2(n15673), .Q(n15683) );
  OR2X1 U16196 ( .IN1(n15685), .IN2(n15686), .Q(n15681) );
  AND2X1 U16197 ( .IN1(n10191), .IN2(n15674), .Q(n15686) );
  AND2X1 U16198 ( .IN1(n10201), .IN2(n15677), .Q(n15685) );
  AND2X1 U16199 ( .IN1(g2834), .IN2(n10897), .Q(n15662) );
  OR2X1 U16200 ( .IN1(n15687), .IN2(n15661), .Q(g30389) );
  AND2X1 U16201 ( .IN1(n10812), .IN2(n15688), .Q(n15661) );
  INVX0 U16202 ( .INP(n15689), .ZN(n15688) );
  OR2X1 U16203 ( .IN1(n15690), .IN2(n15691), .Q(n15689) );
  AND2X1 U16204 ( .IN1(n15667), .IN2(n15692), .Q(n15691) );
  OR2X1 U16205 ( .IN1(n15693), .IN2(n15694), .Q(n15692) );
  OR2X1 U16206 ( .IN1(n15695), .IN2(n15696), .Q(n15694) );
  AND2X1 U16207 ( .IN1(n15673), .IN2(g2775), .Q(n15696) );
  AND2X1 U16208 ( .IN1(n15674), .IN2(g2771), .Q(n15695) );
  OR2X1 U16209 ( .IN1(n15697), .IN2(n15698), .Q(n15693) );
  AND2X1 U16210 ( .IN1(n15677), .IN2(g2787), .Q(n15698) );
  AND2X1 U16211 ( .IN1(n15678), .IN2(g2783), .Q(n15697) );
  AND2X1 U16212 ( .IN1(n15699), .IN2(n15680), .Q(n15690) );
  INVX0 U16213 ( .INP(n15667), .ZN(n15680) );
  AND2X1 U16214 ( .IN1(n5600), .IN2(n15700), .Q(n15667) );
  AND2X1 U16215 ( .IN1(n735), .IN2(n12071), .Q(n15700) );
  INVX0 U16216 ( .INP(n14346), .ZN(n735) );
  OR2X1 U16217 ( .IN1(n11197), .IN2(g2741), .Q(n14346) );
  OR2X1 U16218 ( .IN1(n15701), .IN2(n15702), .Q(n15699) );
  OR2X1 U16219 ( .IN1(n15703), .IN2(n15704), .Q(n15702) );
  AND2X1 U16220 ( .IN1(n15678), .IN2(n10572), .Q(n15704) );
  AND2X1 U16221 ( .IN1(n10193), .IN2(n15673), .Q(n15703) );
  OR2X1 U16222 ( .IN1(n15705), .IN2(n15706), .Q(n15701) );
  AND2X1 U16223 ( .IN1(n10197), .IN2(n15674), .Q(n15706) );
  INVX0 U16224 ( .INP(n15707), .ZN(n15674) );
  AND2X1 U16225 ( .IN1(n10198), .IN2(n15677), .Q(n15705) );
  AND2X1 U16226 ( .IN1(g2831), .IN2(n10896), .Q(n15687) );
  OR2X1 U16227 ( .IN1(n15708), .IN2(n15709), .Q(g30388) );
  AND2X1 U16228 ( .IN1(n10900), .IN2(g2735), .Q(n15709) );
  AND2X1 U16229 ( .IN1(n15710), .IN2(n3730), .Q(n15708) );
  XNOR2X1 U16230 ( .IN1(n3506), .IN2(g2741), .Q(n15710) );
  OR2X1 U16231 ( .IN1(n5600), .IN2(n15711), .Q(n3506) );
  OR2X1 U16232 ( .IN1(n15712), .IN2(n15713), .Q(g30387) );
  OR2X1 U16233 ( .IN1(n15714), .IN2(n15715), .Q(n15713) );
  AND2X1 U16234 ( .IN1(n15716), .IN2(n5777), .Q(n15715) );
  AND2X1 U16235 ( .IN1(n15717), .IN2(n5457), .Q(n15716) );
  AND2X1 U16236 ( .IN1(n15718), .IN2(g2681), .Q(n15714) );
  OR2X1 U16237 ( .IN1(n10884), .IN2(n15719), .Q(n15718) );
  AND2X1 U16238 ( .IN1(n15720), .IN2(g2675), .Q(n15719) );
  AND2X1 U16239 ( .IN1(n15721), .IN2(n9262), .Q(n15712) );
  OR2X1 U16240 ( .IN1(n15722), .IN2(n15723), .Q(g30386) );
  AND2X1 U16241 ( .IN1(n15724), .IN2(g2675), .Q(n15723) );
  AND2X1 U16242 ( .IN1(n15721), .IN2(g2681), .Q(n15722) );
  OR2X1 U16243 ( .IN1(n15725), .IN2(n15726), .Q(g30385) );
  OR2X1 U16244 ( .IN1(n15727), .IN2(n15728), .Q(n15726) );
  AND2X1 U16245 ( .IN1(n15717), .IN2(n5418), .Q(n15728) );
  AND2X1 U16246 ( .IN1(n15721), .IN2(g2661), .Q(n15727) );
  INVX0 U16247 ( .INP(n15724), .ZN(n15721) );
  OR2X1 U16248 ( .IN1(n10884), .IN2(n15720), .Q(n15724) );
  AND2X1 U16249 ( .IN1(n10900), .IN2(g2657), .Q(n15725) );
  OR2X1 U16250 ( .IN1(n15729), .IN2(n15730), .Q(g30384) );
  OR2X1 U16251 ( .IN1(n15731), .IN2(n15732), .Q(n15730) );
  AND2X1 U16252 ( .IN1(n15733), .IN2(g2657), .Q(n15732) );
  OR2X1 U16253 ( .IN1(n15734), .IN2(n14112), .Q(n15733) );
  AND2X1 U16254 ( .IN1(n14136), .IN2(n10804), .Q(n15734) );
  INVX0 U16255 ( .INP(n10539), .ZN(n14136) );
  AND2X1 U16256 ( .IN1(n15735), .IN2(n10539), .Q(n15731) );
  AND2X1 U16257 ( .IN1(n3517), .IN2(n15736), .Q(n15735) );
  XNOR2X1 U16258 ( .IN1(g2652), .IN2(n10070), .Q(n15736) );
  AND2X1 U16259 ( .IN1(n10901), .IN2(g2652), .Q(n15729) );
  OR2X1 U16260 ( .IN1(n15737), .IN2(n15738), .Q(g30383) );
  AND2X1 U16261 ( .IN1(n15739), .IN2(n10803), .Q(n15738) );
  OR2X1 U16262 ( .IN1(n15740), .IN2(n15741), .Q(n15739) );
  AND2X1 U16263 ( .IN1(n15742), .IN2(n15743), .Q(n15741) );
  OR2X1 U16264 ( .IN1(n5524), .IN2(g2555), .Q(n15743) );
  AND2X1 U16265 ( .IN1(test_so34), .IN2(n15744), .Q(n15740) );
  AND2X1 U16266 ( .IN1(test_so66), .IN2(n10896), .Q(n15737) );
  OR2X1 U16267 ( .IN1(n15745), .IN2(n15746), .Q(g30382) );
  OR2X1 U16268 ( .IN1(n15747), .IN2(n15748), .Q(n15746) );
  AND2X1 U16269 ( .IN1(n15749), .IN2(n5782), .Q(n15748) );
  AND2X1 U16270 ( .IN1(n15750), .IN2(n5461), .Q(n15749) );
  AND2X1 U16271 ( .IN1(n15751), .IN2(g2547), .Q(n15747) );
  OR2X1 U16272 ( .IN1(n10885), .IN2(n15752), .Q(n15751) );
  AND2X1 U16273 ( .IN1(n15753), .IN2(g2541), .Q(n15752) );
  AND2X1 U16274 ( .IN1(n15754), .IN2(n9295), .Q(n15745) );
  OR2X1 U16275 ( .IN1(n15755), .IN2(n15756), .Q(g30381) );
  AND2X1 U16276 ( .IN1(n15757), .IN2(g2541), .Q(n15756) );
  AND2X1 U16277 ( .IN1(n15754), .IN2(g2547), .Q(n15755) );
  OR2X1 U16278 ( .IN1(n15758), .IN2(n15759), .Q(g30380) );
  OR2X1 U16279 ( .IN1(n15760), .IN2(n15761), .Q(n15759) );
  AND2X1 U16280 ( .IN1(n15750), .IN2(n5420), .Q(n15761) );
  AND2X1 U16281 ( .IN1(n15754), .IN2(g2527), .Q(n15760) );
  INVX0 U16282 ( .INP(n15757), .ZN(n15754) );
  OR2X1 U16283 ( .IN1(n10885), .IN2(n15753), .Q(n15757) );
  AND2X1 U16284 ( .IN1(n10901), .IN2(g2523), .Q(n15758) );
  OR2X1 U16285 ( .IN1(n15762), .IN2(n15763), .Q(g30379) );
  OR2X1 U16286 ( .IN1(n15764), .IN2(n15765), .Q(n15763) );
  AND2X1 U16287 ( .IN1(n15766), .IN2(g2523), .Q(n15765) );
  OR2X1 U16288 ( .IN1(n15767), .IN2(n14144), .Q(n15766) );
  AND2X1 U16289 ( .IN1(n14170), .IN2(n10803), .Q(n15767) );
  INVX0 U16290 ( .INP(n10546), .ZN(n14170) );
  AND2X1 U16291 ( .IN1(n15768), .IN2(n10546), .Q(n15764) );
  AND2X1 U16292 ( .IN1(n3536), .IN2(n15769), .Q(n15768) );
  XNOR2X1 U16293 ( .IN1(g2518), .IN2(n10067), .Q(n15769) );
  AND2X1 U16294 ( .IN1(n10901), .IN2(g2518), .Q(n15762) );
  OR2X1 U16295 ( .IN1(n15770), .IN2(n15771), .Q(g30378) );
  AND2X1 U16296 ( .IN1(n15772), .IN2(n10802), .Q(n15771) );
  OR2X1 U16297 ( .IN1(n15773), .IN2(n15774), .Q(n15772) );
  AND2X1 U16298 ( .IN1(n15775), .IN2(n15776), .Q(n15774) );
  OR2X1 U16299 ( .IN1(n5523), .IN2(test_so79), .Q(n15776) );
  AND2X1 U16300 ( .IN1(n15777), .IN2(g2461), .Q(n15773) );
  AND2X1 U16301 ( .IN1(n10902), .IN2(g2441), .Q(n15770) );
  OR2X1 U16302 ( .IN1(n15778), .IN2(n15779), .Q(g30377) );
  OR2X1 U16303 ( .IN1(n15780), .IN2(n15781), .Q(n15779) );
  AND2X1 U16304 ( .IN1(n15782), .IN2(n10588), .Q(n15781) );
  AND2X1 U16305 ( .IN1(n15783), .IN2(n5459), .Q(n15782) );
  AND2X1 U16306 ( .IN1(test_so89), .IN2(n15784), .Q(n15780) );
  OR2X1 U16307 ( .IN1(n10885), .IN2(n15785), .Q(n15784) );
  AND2X1 U16308 ( .IN1(n15786), .IN2(g2407), .Q(n15785) );
  AND2X1 U16309 ( .IN1(n15787), .IN2(n9324), .Q(n15778) );
  OR2X1 U16310 ( .IN1(n15788), .IN2(n15789), .Q(g30376) );
  AND2X1 U16311 ( .IN1(n15790), .IN2(g2407), .Q(n15789) );
  AND2X1 U16312 ( .IN1(test_so89), .IN2(n15787), .Q(n15788) );
  OR2X1 U16313 ( .IN1(n15791), .IN2(n15792), .Q(g30375) );
  OR2X1 U16314 ( .IN1(n15793), .IN2(n15794), .Q(n15792) );
  AND2X1 U16315 ( .IN1(n15783), .IN2(n5421), .Q(n15794) );
  AND2X1 U16316 ( .IN1(n15787), .IN2(g2393), .Q(n15793) );
  INVX0 U16317 ( .INP(n15790), .ZN(n15787) );
  OR2X1 U16318 ( .IN1(n10885), .IN2(n15786), .Q(n15790) );
  AND2X1 U16319 ( .IN1(n10902), .IN2(g2389), .Q(n15791) );
  OR2X1 U16320 ( .IN1(n15795), .IN2(n15796), .Q(g30374) );
  OR2X1 U16321 ( .IN1(n15797), .IN2(n15798), .Q(n15796) );
  AND2X1 U16322 ( .IN1(n15799), .IN2(g2389), .Q(n15798) );
  OR2X1 U16323 ( .IN1(n15800), .IN2(n14178), .Q(n15799) );
  AND2X1 U16324 ( .IN1(n14203), .IN2(n10802), .Q(n15800) );
  INVX0 U16325 ( .INP(n10541), .ZN(n14203) );
  AND2X1 U16326 ( .IN1(n15801), .IN2(n10541), .Q(n15797) );
  AND2X1 U16327 ( .IN1(n3555), .IN2(n15802), .Q(n15801) );
  XNOR2X1 U16328 ( .IN1(g2384), .IN2(n10066), .Q(n15802) );
  AND2X1 U16329 ( .IN1(n10902), .IN2(g2384), .Q(n15795) );
  OR2X1 U16330 ( .IN1(n15803), .IN2(n15804), .Q(g30373) );
  AND2X1 U16331 ( .IN1(n15805), .IN2(n10802), .Q(n15804) );
  OR2X1 U16332 ( .IN1(n15806), .IN2(n15807), .Q(n15805) );
  AND2X1 U16333 ( .IN1(n15808), .IN2(n15809), .Q(n15807) );
  OR2X1 U16334 ( .IN1(n5513), .IN2(g2287), .Q(n15809) );
  AND2X1 U16335 ( .IN1(n15810), .IN2(g2327), .Q(n15806) );
  AND2X1 U16336 ( .IN1(n10897), .IN2(g2307), .Q(n15803) );
  OR2X1 U16337 ( .IN1(n15811), .IN2(n15812), .Q(g30372) );
  OR2X1 U16338 ( .IN1(n15813), .IN2(n15814), .Q(n15812) );
  AND2X1 U16339 ( .IN1(n15815), .IN2(n5778), .Q(n15814) );
  AND2X1 U16340 ( .IN1(n15816), .IN2(n5458), .Q(n15815) );
  AND2X1 U16341 ( .IN1(n15817), .IN2(g2279), .Q(n15813) );
  OR2X1 U16342 ( .IN1(n10885), .IN2(n15818), .Q(n15817) );
  AND2X1 U16343 ( .IN1(n15819), .IN2(g2273), .Q(n15818) );
  AND2X1 U16344 ( .IN1(n15820), .IN2(n9273), .Q(n15811) );
  OR2X1 U16345 ( .IN1(n15821), .IN2(n15822), .Q(g30371) );
  AND2X1 U16346 ( .IN1(n15823), .IN2(g2273), .Q(n15822) );
  AND2X1 U16347 ( .IN1(n15820), .IN2(g2279), .Q(n15821) );
  OR2X1 U16348 ( .IN1(n15824), .IN2(n15825), .Q(g30370) );
  OR2X1 U16349 ( .IN1(n15826), .IN2(n15827), .Q(n15825) );
  AND2X1 U16350 ( .IN1(n15816), .IN2(n5419), .Q(n15827) );
  AND2X1 U16351 ( .IN1(n15820), .IN2(g2259), .Q(n15826) );
  INVX0 U16352 ( .INP(n15823), .ZN(n15820) );
  OR2X1 U16353 ( .IN1(n10885), .IN2(n15819), .Q(n15823) );
  AND2X1 U16354 ( .IN1(n10902), .IN2(g2255), .Q(n15824) );
  OR2X1 U16355 ( .IN1(n15828), .IN2(n15829), .Q(g30369) );
  OR2X1 U16356 ( .IN1(n15830), .IN2(n15831), .Q(n15829) );
  AND2X1 U16357 ( .IN1(n15832), .IN2(g2255), .Q(n15831) );
  OR2X1 U16358 ( .IN1(n15833), .IN2(n14211), .Q(n15832) );
  AND2X1 U16359 ( .IN1(n14236), .IN2(n10802), .Q(n15833) );
  INVX0 U16360 ( .INP(n10547), .ZN(n14236) );
  AND2X1 U16361 ( .IN1(n15834), .IN2(n10547), .Q(n15830) );
  AND2X1 U16362 ( .IN1(n3574), .IN2(n15835), .Q(n15834) );
  XNOR2X1 U16363 ( .IN1(g2250), .IN2(n10069), .Q(n15835) );
  AND2X1 U16364 ( .IN1(n10902), .IN2(g2250), .Q(n15828) );
  OR2X1 U16365 ( .IN1(n15836), .IN2(n15837), .Q(g30368) );
  AND2X1 U16366 ( .IN1(n15838), .IN2(n10802), .Q(n15837) );
  OR2X1 U16367 ( .IN1(n15839), .IN2(n15840), .Q(n15838) );
  AND2X1 U16368 ( .IN1(n15841), .IN2(n15842), .Q(n15840) );
  OR2X1 U16369 ( .IN1(n5514), .IN2(g2153), .Q(n15842) );
  AND2X1 U16370 ( .IN1(n15843), .IN2(g2193), .Q(n15839) );
  AND2X1 U16371 ( .IN1(n10902), .IN2(g2173), .Q(n15836) );
  OR2X1 U16372 ( .IN1(n15844), .IN2(n15845), .Q(g30367) );
  OR2X1 U16373 ( .IN1(n15846), .IN2(n15847), .Q(n15845) );
  AND2X1 U16374 ( .IN1(n15848), .IN2(n5784), .Q(n15847) );
  AND2X1 U16375 ( .IN1(n15849), .IN2(n5463), .Q(n15848) );
  AND2X1 U16376 ( .IN1(n15850), .IN2(g2122), .Q(n15846) );
  OR2X1 U16377 ( .IN1(n10885), .IN2(n15851), .Q(n15850) );
  AND2X1 U16378 ( .IN1(n15852), .IN2(g2116), .Q(n15851) );
  AND2X1 U16379 ( .IN1(n15853), .IN2(g2126), .Q(n15844) );
  OR2X1 U16380 ( .IN1(n15854), .IN2(n15855), .Q(g30366) );
  AND2X1 U16381 ( .IN1(n15856), .IN2(g2116), .Q(n15855) );
  AND2X1 U16382 ( .IN1(n15853), .IN2(g2122), .Q(n15854) );
  OR2X1 U16383 ( .IN1(n15857), .IN2(n15858), .Q(g30365) );
  OR2X1 U16384 ( .IN1(n15859), .IN2(n15860), .Q(n15858) );
  AND2X1 U16385 ( .IN1(n15849), .IN2(n5666), .Q(n15860) );
  AND2X1 U16386 ( .IN1(n15853), .IN2(g2102), .Q(n15859) );
  INVX0 U16387 ( .INP(n15856), .ZN(n15853) );
  OR2X1 U16388 ( .IN1(n10885), .IN2(n15852), .Q(n15856) );
  AND2X1 U16389 ( .IN1(n10902), .IN2(g2098), .Q(n15857) );
  OR2X1 U16390 ( .IN1(n15861), .IN2(n15862), .Q(g30364) );
  OR2X1 U16391 ( .IN1(n15863), .IN2(n15864), .Q(n15862) );
  AND2X1 U16392 ( .IN1(n15865), .IN2(g2098), .Q(n15864) );
  OR2X1 U16393 ( .IN1(n15866), .IN2(n14244), .Q(n15865) );
  AND2X1 U16394 ( .IN1(n14270), .IN2(n10802), .Q(n15866) );
  AND2X1 U16395 ( .IN1(n15867), .IN2(n15868), .Q(n15863) );
  XNOR2X1 U16396 ( .IN1(n10065), .IN2(test_so78), .Q(n15868) );
  AND2X1 U16397 ( .IN1(n10549), .IN2(n3593), .Q(n15867) );
  AND2X1 U16398 ( .IN1(test_so78), .IN2(n10895), .Q(n15861) );
  OR2X1 U16399 ( .IN1(n15869), .IN2(n15870), .Q(g30363) );
  AND2X1 U16400 ( .IN1(n15871), .IN2(n10801), .Q(n15870) );
  OR2X1 U16401 ( .IN1(n15872), .IN2(n15873), .Q(n15871) );
  AND2X1 U16402 ( .IN1(n15874), .IN2(n15875), .Q(n15873) );
  OR2X1 U16403 ( .IN1(n5505), .IN2(g1996), .Q(n15875) );
  AND2X1 U16404 ( .IN1(test_so59), .IN2(n15876), .Q(n15872) );
  AND2X1 U16405 ( .IN1(n10902), .IN2(g2016), .Q(n15869) );
  OR2X1 U16406 ( .IN1(n15877), .IN2(n15878), .Q(g30362) );
  OR2X1 U16407 ( .IN1(n15879), .IN2(n15880), .Q(n15878) );
  AND2X1 U16408 ( .IN1(n15881), .IN2(n5783), .Q(n15880) );
  AND2X1 U16409 ( .IN1(n15882), .IN2(n5462), .Q(n15881) );
  AND2X1 U16410 ( .IN1(n15883), .IN2(g1988), .Q(n15879) );
  OR2X1 U16411 ( .IN1(n10885), .IN2(n15884), .Q(n15883) );
  AND2X1 U16412 ( .IN1(n15885), .IN2(g1982), .Q(n15884) );
  AND2X1 U16413 ( .IN1(n15886), .IN2(g1992), .Q(n15877) );
  OR2X1 U16414 ( .IN1(n15887), .IN2(n15888), .Q(g30361) );
  AND2X1 U16415 ( .IN1(n15889), .IN2(g1982), .Q(n15888) );
  AND2X1 U16416 ( .IN1(n15886), .IN2(g1988), .Q(n15887) );
  OR2X1 U16417 ( .IN1(n15890), .IN2(n15891), .Q(g30360) );
  OR2X1 U16418 ( .IN1(n15892), .IN2(n15893), .Q(n15891) );
  AND2X1 U16419 ( .IN1(n15882), .IN2(n5664), .Q(n15893) );
  AND2X1 U16420 ( .IN1(n15886), .IN2(g1968), .Q(n15892) );
  INVX0 U16421 ( .INP(n15889), .ZN(n15886) );
  OR2X1 U16422 ( .IN1(n10885), .IN2(n15885), .Q(n15889) );
  AND2X1 U16423 ( .IN1(n10902), .IN2(g1964), .Q(n15890) );
  OR2X1 U16424 ( .IN1(n15894), .IN2(n15895), .Q(g30359) );
  OR2X1 U16425 ( .IN1(n15896), .IN2(n15897), .Q(n15895) );
  AND2X1 U16426 ( .IN1(n15898), .IN2(g1964), .Q(n15897) );
  OR2X1 U16427 ( .IN1(n15899), .IN2(n14278), .Q(n15898) );
  AND2X1 U16428 ( .IN1(n14304), .IN2(n10801), .Q(n15899) );
  INVX0 U16429 ( .INP(n10538), .ZN(n14304) );
  AND2X1 U16430 ( .IN1(n15900), .IN2(n10538), .Q(n15896) );
  AND2X1 U16431 ( .IN1(n3611), .IN2(n15901), .Q(n15900) );
  XNOR2X1 U16432 ( .IN1(g1959), .IN2(n10063), .Q(n15901) );
  AND2X1 U16433 ( .IN1(n10902), .IN2(g1959), .Q(n15894) );
  OR2X1 U16434 ( .IN1(n15902), .IN2(n15903), .Q(g30358) );
  AND2X1 U16435 ( .IN1(n15904), .IN2(n10801), .Q(n15903) );
  OR2X1 U16436 ( .IN1(n15905), .IN2(n15906), .Q(n15904) );
  AND2X1 U16437 ( .IN1(n15907), .IN2(n15908), .Q(n15906) );
  OR2X1 U16438 ( .IN1(n5503), .IN2(test_so8), .Q(n15908) );
  AND2X1 U16439 ( .IN1(n15909), .IN2(g1902), .Q(n15905) );
  AND2X1 U16440 ( .IN1(n10901), .IN2(g1882), .Q(n15902) );
  OR2X1 U16441 ( .IN1(n15910), .IN2(n15911), .Q(g30357) );
  OR2X1 U16442 ( .IN1(n15912), .IN2(n15913), .Q(n15911) );
  AND2X1 U16443 ( .IN1(n15914), .IN2(n5785), .Q(n15913) );
  AND2X1 U16444 ( .IN1(n15915), .IN2(n5464), .Q(n15914) );
  AND2X1 U16445 ( .IN1(n15916), .IN2(g1854), .Q(n15912) );
  OR2X1 U16446 ( .IN1(n10885), .IN2(n15917), .Q(n15916) );
  AND2X1 U16447 ( .IN1(n15918), .IN2(g1848), .Q(n15917) );
  AND2X1 U16448 ( .IN1(n15919), .IN2(g1858), .Q(n15910) );
  OR2X1 U16449 ( .IN1(n15920), .IN2(n15921), .Q(g30356) );
  AND2X1 U16450 ( .IN1(n15922), .IN2(g1848), .Q(n15921) );
  AND2X1 U16451 ( .IN1(n15919), .IN2(g1854), .Q(n15920) );
  OR2X1 U16452 ( .IN1(n15923), .IN2(n15924), .Q(g30355) );
  OR2X1 U16453 ( .IN1(n15925), .IN2(n15926), .Q(n15924) );
  AND2X1 U16454 ( .IN1(n15915), .IN2(n5665), .Q(n15926) );
  AND2X1 U16455 ( .IN1(n15919), .IN2(g1834), .Q(n15925) );
  INVX0 U16456 ( .INP(n15922), .ZN(n15919) );
  OR2X1 U16457 ( .IN1(n10885), .IN2(n15918), .Q(n15922) );
  AND2X1 U16458 ( .IN1(n10901), .IN2(g1830), .Q(n15923) );
  OR2X1 U16459 ( .IN1(n15927), .IN2(n15928), .Q(g30354) );
  OR2X1 U16460 ( .IN1(n15929), .IN2(n15930), .Q(n15928) );
  AND2X1 U16461 ( .IN1(n15931), .IN2(g1830), .Q(n15930) );
  OR2X1 U16462 ( .IN1(n15932), .IN2(n14312), .Q(n15931) );
  AND2X1 U16463 ( .IN1(n14336), .IN2(n10800), .Q(n15932) );
  INVX0 U16464 ( .INP(n10544), .ZN(n14336) );
  AND2X1 U16465 ( .IN1(n15933), .IN2(n10544), .Q(n15929) );
  AND2X1 U16466 ( .IN1(n3628), .IN2(n15934), .Q(n15933) );
  XNOR2X1 U16467 ( .IN1(g1825), .IN2(n10064), .Q(n15934) );
  AND2X1 U16468 ( .IN1(n10901), .IN2(g1825), .Q(n15927) );
  OR2X1 U16469 ( .IN1(n15935), .IN2(n15936), .Q(g30353) );
  AND2X1 U16470 ( .IN1(n15937), .IN2(n10804), .Q(n15936) );
  OR2X1 U16471 ( .IN1(n15938), .IN2(n15939), .Q(n15937) );
  AND2X1 U16472 ( .IN1(n15940), .IN2(n15941), .Q(n15939) );
  OR2X1 U16473 ( .IN1(n5504), .IN2(g1728), .Q(n15941) );
  AND2X1 U16474 ( .IN1(n15942), .IN2(g1768), .Q(n15938) );
  AND2X1 U16475 ( .IN1(n10901), .IN2(g1748), .Q(n15935) );
  OR2X1 U16476 ( .IN1(n15943), .IN2(n15944), .Q(g30352) );
  OR2X1 U16477 ( .IN1(n15945), .IN2(n15946), .Q(n15944) );
  AND2X1 U16478 ( .IN1(n15947), .IN2(n5780), .Q(n15946) );
  AND2X1 U16479 ( .IN1(n15948), .IN2(n15949), .Q(n15947) );
  AND2X1 U16480 ( .IN1(n5460), .IN2(n10800), .Q(n15948) );
  AND2X1 U16481 ( .IN1(n15950), .IN2(g1720), .Q(n15945) );
  OR2X1 U16482 ( .IN1(n10886), .IN2(n15951), .Q(n15950) );
  AND2X1 U16483 ( .IN1(n15949), .IN2(g1714), .Q(n15951) );
  AND2X1 U16484 ( .IN1(n15952), .IN2(n9236), .Q(n15943) );
  OR2X1 U16485 ( .IN1(n15953), .IN2(n15954), .Q(g30351) );
  AND2X1 U16486 ( .IN1(n15955), .IN2(g1714), .Q(n15954) );
  AND2X1 U16487 ( .IN1(n15952), .IN2(g1720), .Q(n15953) );
  OR2X1 U16488 ( .IN1(n15956), .IN2(n15957), .Q(g30350) );
  OR2X1 U16489 ( .IN1(n15958), .IN2(n15959), .Q(n15957) );
  AND2X1 U16490 ( .IN1(n10901), .IN2(g1696), .Q(n15959) );
  AND2X1 U16491 ( .IN1(n15960), .IN2(n10800), .Q(n15958) );
  AND2X1 U16492 ( .IN1(n15949), .IN2(n5417), .Q(n15960) );
  AND2X1 U16493 ( .IN1(n15952), .IN2(g1700), .Q(n15956) );
  INVX0 U16494 ( .INP(n15955), .ZN(n15952) );
  OR2X1 U16495 ( .IN1(n10886), .IN2(n15949), .Q(n15955) );
  OR2X1 U16496 ( .IN1(n15961), .IN2(n15962), .Q(g30349) );
  OR2X1 U16497 ( .IN1(n15963), .IN2(n15964), .Q(n15962) );
  AND2X1 U16498 ( .IN1(n15965), .IN2(g1696), .Q(n15964) );
  OR2X1 U16499 ( .IN1(n15966), .IN2(n14344), .Q(n15965) );
  AND2X1 U16500 ( .IN1(n14371), .IN2(n10800), .Q(n15966) );
  INVX0 U16501 ( .INP(n10548), .ZN(n14371) );
  AND2X1 U16502 ( .IN1(n15967), .IN2(n10548), .Q(n15963) );
  AND2X1 U16503 ( .IN1(n3646), .IN2(n15968), .Q(n15967) );
  XNOR2X1 U16504 ( .IN1(g1691), .IN2(n10068), .Q(n15968) );
  AND2X1 U16505 ( .IN1(n10901), .IN2(g1691), .Q(n15961) );
  OR2X1 U16506 ( .IN1(n15969), .IN2(n15970), .Q(g30348) );
  OR2X1 U16507 ( .IN1(n15971), .IN2(n15972), .Q(n15970) );
  AND2X1 U16508 ( .IN1(n15973), .IN2(g1632), .Q(n15972) );
  OR2X1 U16509 ( .IN1(n15974), .IN2(n14344), .Q(n15973) );
  AND2X1 U16510 ( .IN1(n15975), .IN2(n10800), .Q(n15974) );
  AND2X1 U16511 ( .IN1(n15976), .IN2(n3646), .Q(n15971) );
  AND2X1 U16512 ( .IN1(g25167), .IN2(n15977), .Q(n15976) );
  OR2X1 U16513 ( .IN1(n5549), .IN2(g1592), .Q(n15977) );
  AND2X1 U16514 ( .IN1(n10901), .IN2(g1612), .Q(n15969) );
  OR2X1 U16515 ( .IN1(n15978), .IN2(n15979), .Q(g30347) );
  AND2X1 U16516 ( .IN1(n10901), .IN2(g1542), .Q(n15979) );
  AND2X1 U16517 ( .IN1(n15980), .IN2(n15981), .Q(n15978) );
  AND2X1 U16518 ( .IN1(n15982), .IN2(n15983), .Q(n15980) );
  INVX0 U16519 ( .INP(n15984), .ZN(n15982) );
  AND2X1 U16520 ( .IN1(n15985), .IN2(n15986), .Q(n15984) );
  OR2X1 U16521 ( .IN1(n10886), .IN2(n10528), .Q(n15986) );
  OR2X1 U16522 ( .IN1(n15987), .IN2(n15988), .Q(g30346) );
  AND2X1 U16523 ( .IN1(n15989), .IN2(n10799), .Q(n15988) );
  AND2X1 U16524 ( .IN1(n15990), .IN2(n15981), .Q(n15989) );
  INVX0 U16525 ( .INP(n15991), .ZN(n15981) );
  AND2X1 U16526 ( .IN1(n15992), .IN2(n15985), .Q(n15990) );
  OR2X1 U16527 ( .IN1(n15993), .IN2(g1542), .Q(n15992) );
  AND2X1 U16528 ( .IN1(n10901), .IN2(g1536), .Q(n15987) );
  OR2X1 U16529 ( .IN1(n15994), .IN2(n15995), .Q(g30345) );
  AND2X1 U16530 ( .IN1(n15996), .IN2(g1514), .Q(n15995) );
  OR2X1 U16531 ( .IN1(n10886), .IN2(n15997), .Q(n15996) );
  XNOR2X1 U16532 ( .IN1(test_so49), .IN2(n5302), .Q(n15997) );
  AND2X1 U16533 ( .IN1(n15998), .IN2(n10799), .Q(n15994) );
  OR2X1 U16534 ( .IN1(n13468), .IN2(n15991), .Q(n15998) );
  AND2X1 U16535 ( .IN1(n15999), .IN2(n10799), .Q(g30344) );
  OR2X1 U16536 ( .IN1(n15991), .IN2(n16000), .Q(n15999) );
  XNOR2X1 U16537 ( .IN1(g1514), .IN2(n5302), .Q(n16000) );
  OR2X1 U16538 ( .IN1(n16001), .IN2(n4173), .Q(n15991) );
  AND2X1 U16539 ( .IN1(n4172), .IN2(n13468), .Q(n16001) );
  AND2X1 U16540 ( .IN1(n4895), .IN2(n16002), .Q(n4172) );
  INVX0 U16541 ( .INP(n16003), .ZN(n16002) );
  OR2X1 U16542 ( .IN1(n5302), .IN2(n16004), .Q(n16003) );
  OR2X1 U16543 ( .IN1(n16005), .IN2(n16006), .Q(g30343) );
  OR2X1 U16544 ( .IN1(n16007), .IN2(n16008), .Q(n16006) );
  AND2X1 U16545 ( .IN1(n16009), .IN2(n10799), .Q(n16008) );
  AND2X1 U16546 ( .IN1(n11213), .IN2(g1361), .Q(n16009) );
  OR2X1 U16547 ( .IN1(n16010), .IN2(n16011), .Q(n11213) );
  AND2X1 U16548 ( .IN1(n10511), .IN2(n13787), .Q(n16010) );
  INVX0 U16549 ( .INP(n16012), .ZN(n16007) );
  OR2X1 U16550 ( .IN1(n10738), .IN2(n10511), .Q(n16012) );
  AND2X1 U16551 ( .IN1(n4175), .IN2(n14378), .Q(n16005) );
  OR2X1 U16552 ( .IN1(n16013), .IN2(n16014), .Q(g30342) );
  OR2X1 U16553 ( .IN1(n16015), .IN2(n16016), .Q(n16014) );
  AND2X1 U16554 ( .IN1(n3736), .IN2(n5553), .Q(n16016) );
  INVX0 U16555 ( .INP(n16017), .ZN(n16015) );
  OR2X1 U16556 ( .IN1(n16018), .IN2(n5553), .Q(n16017) );
  OR2X1 U16557 ( .IN1(n13799), .IN2(n3736), .Q(n16018) );
  AND2X1 U16558 ( .IN1(n10902), .IN2(g1256), .Q(n16013) );
  OR2X1 U16559 ( .IN1(n16019), .IN2(n16020), .Q(g30341) );
  AND2X1 U16560 ( .IN1(n10900), .IN2(g1199), .Q(n16020) );
  AND2X1 U16561 ( .IN1(n16021), .IN2(n16022), .Q(n16019) );
  AND2X1 U16562 ( .IN1(n16023), .IN2(n16024), .Q(n16021) );
  INVX0 U16563 ( .INP(n16025), .ZN(n16023) );
  AND2X1 U16564 ( .IN1(n16026), .IN2(n16027), .Q(n16025) );
  OR2X1 U16565 ( .IN1(n10886), .IN2(n10529), .Q(n16027) );
  OR2X1 U16566 ( .IN1(n16028), .IN2(n16029), .Q(g30340) );
  AND2X1 U16567 ( .IN1(n16030), .IN2(n10799), .Q(n16029) );
  AND2X1 U16568 ( .IN1(n16031), .IN2(n16022), .Q(n16030) );
  INVX0 U16569 ( .INP(n16032), .ZN(n16022) );
  AND2X1 U16570 ( .IN1(n16033), .IN2(n16026), .Q(n16031) );
  OR2X1 U16571 ( .IN1(n16034), .IN2(g1199), .Q(n16033) );
  AND2X1 U16572 ( .IN1(n10900), .IN2(g1193), .Q(n16028) );
  OR2X1 U16573 ( .IN1(n16035), .IN2(n16036), .Q(g30339) );
  AND2X1 U16574 ( .IN1(n16037), .IN2(g1171), .Q(n16036) );
  OR2X1 U16575 ( .IN1(n10886), .IN2(n16038), .Q(n16037) );
  XNOR2X1 U16576 ( .IN1(g1183), .IN2(n5304), .Q(n16038) );
  AND2X1 U16577 ( .IN1(n16039), .IN2(n10798), .Q(n16035) );
  OR2X1 U16578 ( .IN1(n13720), .IN2(n16032), .Q(n16039) );
  AND2X1 U16579 ( .IN1(n16040), .IN2(n10798), .Q(g30338) );
  OR2X1 U16580 ( .IN1(n16032), .IN2(n16041), .Q(n16040) );
  XNOR2X1 U16581 ( .IN1(g1171), .IN2(n5304), .Q(n16041) );
  OR2X1 U16582 ( .IN1(n16042), .IN2(n4191), .Q(n16032) );
  AND2X1 U16583 ( .IN1(n4190), .IN2(n13720), .Q(n16042) );
  AND2X1 U16584 ( .IN1(n4920), .IN2(n16043), .Q(n4190) );
  INVX0 U16585 ( .INP(n16044), .ZN(n16043) );
  OR2X1 U16586 ( .IN1(n5304), .IN2(n16045), .Q(n16044) );
  OR2X1 U16587 ( .IN1(n16046), .IN2(n16047), .Q(g30337) );
  OR2X1 U16588 ( .IN1(n16048), .IN2(n16049), .Q(n16047) );
  AND2X1 U16589 ( .IN1(n16050), .IN2(n10798), .Q(n16049) );
  AND2X1 U16590 ( .IN1(n11097), .IN2(g1018), .Q(n16050) );
  OR2X1 U16591 ( .IN1(n16051), .IN2(n16052), .Q(n11097) );
  AND2X1 U16592 ( .IN1(n10510), .IN2(n13806), .Q(n16051) );
  INVX0 U16593 ( .INP(n16053), .ZN(n16048) );
  OR2X1 U16594 ( .IN1(n10738), .IN2(n10510), .Q(n16053) );
  AND2X1 U16595 ( .IN1(n4193), .IN2(n14394), .Q(n16046) );
  OR2X1 U16596 ( .IN1(n16054), .IN2(n16055), .Q(g30336) );
  OR2X1 U16597 ( .IN1(n16056), .IN2(n16057), .Q(n16055) );
  AND2X1 U16598 ( .IN1(n3741), .IN2(n5560), .Q(n16057) );
  INVX0 U16599 ( .INP(n16058), .ZN(n16056) );
  OR2X1 U16600 ( .IN1(n16059), .IN2(n5560), .Q(n16058) );
  OR2X1 U16601 ( .IN1(n13818), .IN2(n3741), .Q(n16059) );
  AND2X1 U16602 ( .IN1(n10900), .IN2(g911), .Q(n16054) );
  OR2X1 U16603 ( .IN1(n16060), .IN2(n16061), .Q(g30335) );
  OR2X1 U16604 ( .IN1(n16062), .IN2(n16063), .Q(n16061) );
  AND2X1 U16605 ( .IN1(n53), .IN2(n5470), .Q(n16063) );
  AND2X1 U16606 ( .IN1(n16064), .IN2(g744), .Q(n16062) );
  AND2X1 U16607 ( .IN1(n2404), .IN2(n16065), .Q(n16064) );
  INVX0 U16608 ( .INP(n53), .ZN(n16065) );
  AND2X1 U16609 ( .IN1(test_so60), .IN2(n16066), .Q(n53) );
  AND2X1 U16610 ( .IN1(n4198), .IN2(n16067), .Q(n16066) );
  OR2X1 U16611 ( .IN1(n5482), .IN2(g736), .Q(n4198) );
  AND2X1 U16612 ( .IN1(test_so60), .IN2(n10895), .Q(n16060) );
  OR2X1 U16613 ( .IN1(n16068), .IN2(n16069), .Q(g30334) );
  OR2X1 U16614 ( .IN1(n16070), .IN2(n16071), .Q(n16069) );
  AND2X1 U16615 ( .IN1(n3745), .IN2(n5294), .Q(n16071) );
  AND2X1 U16616 ( .IN1(n16072), .IN2(g577), .Q(n16070) );
  AND2X1 U16617 ( .IN1(n2421), .IN2(n16073), .Q(n16072) );
  INVX0 U16618 ( .INP(n3745), .ZN(n16073) );
  AND2X1 U16619 ( .IN1(n10900), .IN2(g586), .Q(n16068) );
  OR2X1 U16620 ( .IN1(n16074), .IN2(n16075), .Q(g30333) );
  AND2X1 U16621 ( .IN1(n10900), .IN2(g142), .Q(n16075) );
  AND2X1 U16622 ( .IN1(n13055), .IN2(n16076), .Q(n16074) );
  XOR2X1 U16623 ( .IN1(test_so73), .IN2(n14600), .Q(n16076) );
  INVX0 U16624 ( .INP(n12326), .ZN(n13055) );
  OR2X1 U16625 ( .IN1(n10886), .IN2(n14602), .Q(n12326) );
  OR2X1 U16626 ( .IN1(n16077), .IN2(n16078), .Q(n14602) );
  AND2X1 U16627 ( .IN1(n14600), .IN2(n16079), .Q(n16077) );
  OR2X1 U16628 ( .IN1(test_so72), .IN2(n16080), .Q(n16079) );
  OR2X1 U16629 ( .IN1(n16081), .IN2(n16082), .Q(g29309) );
  OR2X1 U16630 ( .IN1(n16083), .IN2(n16084), .Q(n16082) );
  AND2X1 U16631 ( .IN1(n16085), .IN2(n14635), .Q(n16084) );
  AND2X1 U16632 ( .IN1(n16086), .IN2(g6541), .Q(n16085) );
  AND2X1 U16633 ( .IN1(n3765), .IN2(n16087), .Q(n16081) );
  OR2X1 U16634 ( .IN1(n13075), .IN2(n5739), .Q(n16087) );
  OR2X1 U16635 ( .IN1(n16088), .IN2(n16089), .Q(g29308) );
  OR2X1 U16636 ( .IN1(n16090), .IN2(n16091), .Q(n16089) );
  AND2X1 U16637 ( .IN1(n5659), .IN2(n16092), .Q(n16091) );
  AND2X1 U16638 ( .IN1(n16093), .IN2(g6527), .Q(n16090) );
  AND2X1 U16639 ( .IN1(n10900), .IN2(g6523), .Q(n16088) );
  OR2X1 U16640 ( .IN1(n16094), .IN2(n16095), .Q(g29307) );
  OR2X1 U16641 ( .IN1(n16096), .IN2(n16097), .Q(n16095) );
  AND2X1 U16642 ( .IN1(n16098), .IN2(n5806), .Q(n16097) );
  AND2X1 U16643 ( .IN1(n5426), .IN2(n16092), .Q(n16098) );
  AND2X1 U16644 ( .IN1(n16099), .IN2(g6519), .Q(n16096) );
  OR2X1 U16645 ( .IN1(n10886), .IN2(n16100), .Q(n16099) );
  AND2X1 U16646 ( .IN1(n16101), .IN2(g6513), .Q(n16100) );
  AND2X1 U16647 ( .IN1(n16093), .IN2(g6523), .Q(n16094) );
  OR2X1 U16648 ( .IN1(n16102), .IN2(n16103), .Q(g29306) );
  AND2X1 U16649 ( .IN1(n16104), .IN2(g6513), .Q(n16103) );
  AND2X1 U16650 ( .IN1(n16093), .IN2(g6519), .Q(n16102) );
  INVX0 U16651 ( .INP(n16104), .ZN(n16093) );
  OR2X1 U16652 ( .IN1(n10886), .IN2(n16101), .Q(n16104) );
  OR2X1 U16653 ( .IN1(n16105), .IN2(n16106), .Q(g29305) );
  OR2X1 U16654 ( .IN1(n16107), .IN2(n16108), .Q(n16106) );
  AND2X1 U16655 ( .IN1(n16109), .IN2(n5748), .Q(n16108) );
  AND2X1 U16656 ( .IN1(n16092), .IN2(g6505), .Q(n16109) );
  AND2X1 U16657 ( .IN1(n10810), .IN2(n16101), .Q(n16092) );
  AND2X1 U16658 ( .IN1(n16110), .IN2(g6500), .Q(n16107) );
  OR2X1 U16659 ( .IN1(n10886), .IN2(n16111), .Q(n16110) );
  AND2X1 U16660 ( .IN1(n10101), .IN2(n16101), .Q(n16111) );
  INVX0 U16661 ( .INP(n16112), .ZN(n16105) );
  OR2X1 U16662 ( .IN1(n14630), .IN2(n16101), .Q(n16112) );
  AND2X1 U16663 ( .IN1(n13113), .IN2(n16113), .Q(n16101) );
  OR2X1 U16664 ( .IN1(n10484), .IN2(n10874), .Q(n14630) );
  OR2X1 U16665 ( .IN1(n16114), .IN2(n16115), .Q(g29304) );
  AND2X1 U16666 ( .IN1(n16116), .IN2(n10798), .Q(n16115) );
  OR2X1 U16667 ( .IN1(n16117), .IN2(n16118), .Q(n16116) );
  AND2X1 U16668 ( .IN1(n16119), .IN2(n13113), .Q(n16118) );
  XNOR2X1 U16669 ( .IN1(n16120), .IN2(n16121), .Q(n16119) );
  OR2X1 U16670 ( .IN1(n16113), .IN2(n5748), .Q(n16120) );
  AND2X1 U16671 ( .IN1(n11096), .IN2(n16122), .Q(n16113) );
  AND2X1 U16672 ( .IN1(g6727), .IN2(g17722), .Q(n16122) );
  AND2X1 U16673 ( .IN1(n10540), .IN2(g6500), .Q(n16117) );
  AND2X1 U16674 ( .IN1(n10900), .IN2(g6505), .Q(n16114) );
  OR2X1 U16675 ( .IN1(n16123), .IN2(n16124), .Q(g29303) );
  OR2X1 U16676 ( .IN1(n16083), .IN2(n16125), .Q(n16124) );
  AND2X1 U16677 ( .IN1(n16126), .IN2(n14762), .Q(n16125) );
  AND2X1 U16678 ( .IN1(n16086), .IN2(g6195), .Q(n16126) );
  AND2X1 U16679 ( .IN1(n3765), .IN2(n16127), .Q(n16123) );
  OR2X1 U16680 ( .IN1(n13092), .IN2(n5741), .Q(n16127) );
  OR2X1 U16681 ( .IN1(n16128), .IN2(n16129), .Q(g29302) );
  OR2X1 U16682 ( .IN1(n16130), .IN2(n16131), .Q(n16129) );
  AND2X1 U16683 ( .IN1(n5667), .IN2(n16132), .Q(n16131) );
  AND2X1 U16684 ( .IN1(n16133), .IN2(g6181), .Q(n16130) );
  AND2X1 U16685 ( .IN1(n10899), .IN2(g6177), .Q(n16128) );
  OR2X1 U16686 ( .IN1(n16134), .IN2(n16135), .Q(g29301) );
  OR2X1 U16687 ( .IN1(n16136), .IN2(n16137), .Q(n16135) );
  AND2X1 U16688 ( .IN1(n16138), .IN2(n5810), .Q(n16137) );
  AND2X1 U16689 ( .IN1(n5430), .IN2(n16132), .Q(n16138) );
  AND2X1 U16690 ( .IN1(n16139), .IN2(g6173), .Q(n16136) );
  OR2X1 U16691 ( .IN1(n10886), .IN2(n16140), .Q(n16139) );
  AND2X1 U16692 ( .IN1(n16141), .IN2(g6167), .Q(n16140) );
  AND2X1 U16693 ( .IN1(n16133), .IN2(g6177), .Q(n16134) );
  OR2X1 U16694 ( .IN1(n16142), .IN2(n16143), .Q(g29300) );
  AND2X1 U16695 ( .IN1(n16144), .IN2(g6167), .Q(n16143) );
  AND2X1 U16696 ( .IN1(n16133), .IN2(g6173), .Q(n16142) );
  OR2X1 U16697 ( .IN1(n16145), .IN2(n16146), .Q(g29299) );
  OR2X1 U16698 ( .IN1(n16147), .IN2(n16148), .Q(n16146) );
  AND2X1 U16699 ( .IN1(n16149), .IN2(n5747), .Q(n16148) );
  AND2X1 U16700 ( .IN1(n16132), .IN2(g6159), .Q(n16149) );
  AND2X1 U16701 ( .IN1(n10809), .IN2(n16141), .Q(n16132) );
  AND2X1 U16702 ( .IN1(n16150), .IN2(g6154), .Q(n16147) );
  OR2X1 U16703 ( .IN1(n10887), .IN2(n16151), .Q(n16150) );
  AND2X1 U16704 ( .IN1(n10100), .IN2(n16141), .Q(n16151) );
  AND2X1 U16705 ( .IN1(n16133), .IN2(g6163), .Q(n16145) );
  INVX0 U16706 ( .INP(n16144), .ZN(n16133) );
  OR2X1 U16707 ( .IN1(n10887), .IN2(n16141), .Q(n16144) );
  AND2X1 U16708 ( .IN1(n13133), .IN2(n16152), .Q(n16141) );
  OR2X1 U16709 ( .IN1(n16153), .IN2(n16154), .Q(g29298) );
  AND2X1 U16710 ( .IN1(n16155), .IN2(n10802), .Q(n16154) );
  OR2X1 U16711 ( .IN1(n16156), .IN2(n16157), .Q(n16155) );
  AND2X1 U16712 ( .IN1(n16158), .IN2(n13133), .Q(n16157) );
  XNOR2X1 U16713 ( .IN1(n16159), .IN2(n16160), .Q(n16158) );
  OR2X1 U16714 ( .IN1(n5747), .IN2(n16152), .Q(n16160) );
  AND2X1 U16715 ( .IN1(test_so69), .IN2(n16161), .Q(n16152) );
  AND2X1 U16716 ( .IN1(g17685), .IN2(n12119), .Q(n16161) );
  AND2X1 U16717 ( .IN1(n13137), .IN2(g6154), .Q(n16156) );
  AND2X1 U16718 ( .IN1(n10899), .IN2(g6159), .Q(n16153) );
  OR2X1 U16719 ( .IN1(n16162), .IN2(n16163), .Q(g29297) );
  OR2X1 U16720 ( .IN1(n16083), .IN2(n16164), .Q(n16163) );
  AND2X1 U16721 ( .IN1(n16165), .IN2(n14889), .Q(n16164) );
  AND2X1 U16722 ( .IN1(n16086), .IN2(g5849), .Q(n16165) );
  AND2X1 U16723 ( .IN1(n3765), .IN2(n16166), .Q(n16162) );
  OR2X1 U16724 ( .IN1(n13091), .IN2(n5736), .Q(n16166) );
  OR2X1 U16725 ( .IN1(n16167), .IN2(n16168), .Q(g29296) );
  OR2X1 U16726 ( .IN1(n16169), .IN2(n16170), .Q(n16168) );
  AND2X1 U16727 ( .IN1(n5663), .IN2(n16171), .Q(n16170) );
  AND2X1 U16728 ( .IN1(n16172), .IN2(g5835), .Q(n16169) );
  AND2X1 U16729 ( .IN1(n10899), .IN2(g5831), .Q(n16167) );
  OR2X1 U16730 ( .IN1(n16173), .IN2(n16174), .Q(g29295) );
  OR2X1 U16731 ( .IN1(n16175), .IN2(n16176), .Q(n16174) );
  AND2X1 U16732 ( .IN1(n16177), .IN2(n5809), .Q(n16176) );
  AND2X1 U16733 ( .IN1(n5429), .IN2(n16171), .Q(n16177) );
  AND2X1 U16734 ( .IN1(n16178), .IN2(g5827), .Q(n16175) );
  OR2X1 U16735 ( .IN1(n10887), .IN2(n16179), .Q(n16178) );
  AND2X1 U16736 ( .IN1(n16180), .IN2(g5821), .Q(n16179) );
  AND2X1 U16737 ( .IN1(n16172), .IN2(g5831), .Q(n16173) );
  OR2X1 U16738 ( .IN1(n16181), .IN2(n16182), .Q(g29294) );
  AND2X1 U16739 ( .IN1(n16183), .IN2(g5821), .Q(n16182) );
  AND2X1 U16740 ( .IN1(n16172), .IN2(g5827), .Q(n16181) );
  INVX0 U16741 ( .INP(n16183), .ZN(n16172) );
  OR2X1 U16742 ( .IN1(n10887), .IN2(n16180), .Q(n16183) );
  OR2X1 U16743 ( .IN1(n16184), .IN2(n16185), .Q(g29293) );
  OR2X1 U16744 ( .IN1(n16186), .IN2(n16187), .Q(n16185) );
  AND2X1 U16745 ( .IN1(n16188), .IN2(n5749), .Q(n16187) );
  AND2X1 U16746 ( .IN1(n16171), .IN2(g5813), .Q(n16188) );
  AND2X1 U16747 ( .IN1(n10808), .IN2(n16180), .Q(n16171) );
  AND2X1 U16748 ( .IN1(n16189), .IN2(g5808), .Q(n16186) );
  OR2X1 U16749 ( .IN1(n10887), .IN2(n16190), .Q(n16189) );
  AND2X1 U16750 ( .IN1(n10102), .IN2(n16180), .Q(n16190) );
  INVX0 U16751 ( .INP(n16191), .ZN(n16184) );
  OR2X1 U16752 ( .IN1(n14624), .IN2(n16180), .Q(n16191) );
  AND2X1 U16753 ( .IN1(n13155), .IN2(n16192), .Q(n16180) );
  OR2X1 U16754 ( .IN1(n10523), .IN2(n10876), .Q(n14624) );
  OR2X1 U16755 ( .IN1(n16193), .IN2(n16194), .Q(g29292) );
  AND2X1 U16756 ( .IN1(n16195), .IN2(n10806), .Q(n16194) );
  OR2X1 U16757 ( .IN1(n16196), .IN2(n16197), .Q(n16195) );
  AND2X1 U16758 ( .IN1(n16198), .IN2(n13155), .Q(n16197) );
  XNOR2X1 U16759 ( .IN1(n16199), .IN2(n16200), .Q(n16198) );
  OR2X1 U16760 ( .IN1(n16192), .IN2(n5749), .Q(n16199) );
  AND2X1 U16761 ( .IN1(n12132), .IN2(n16201), .Q(n16192) );
  AND2X1 U16762 ( .IN1(g6035), .IN2(g17646), .Q(n16201) );
  AND2X1 U16763 ( .IN1(n13159), .IN2(g5808), .Q(n16196) );
  AND2X1 U16764 ( .IN1(n10899), .IN2(g5813), .Q(n16193) );
  OR2X1 U16765 ( .IN1(n16202), .IN2(n16203), .Q(g29291) );
  OR2X1 U16766 ( .IN1(n16083), .IN2(n16204), .Q(n16203) );
  AND2X1 U16767 ( .IN1(n16205), .IN2(n15015), .Q(n16204) );
  AND2X1 U16768 ( .IN1(n16086), .IN2(g5503), .Q(n16205) );
  AND2X1 U16769 ( .IN1(n3765), .IN2(n16206), .Q(n16202) );
  OR2X1 U16770 ( .IN1(n13093), .IN2(n5737), .Q(n16206) );
  OR2X1 U16771 ( .IN1(n16207), .IN2(n16208), .Q(g29290) );
  OR2X1 U16772 ( .IN1(n16209), .IN2(n16210), .Q(n16208) );
  AND2X1 U16773 ( .IN1(n5660), .IN2(n16211), .Q(n16210) );
  AND2X1 U16774 ( .IN1(n16212), .IN2(g5489), .Q(n16209) );
  AND2X1 U16775 ( .IN1(n10898), .IN2(g5485), .Q(n16207) );
  OR2X1 U16776 ( .IN1(n16213), .IN2(n16214), .Q(g29289) );
  OR2X1 U16777 ( .IN1(n16215), .IN2(n16216), .Q(n16214) );
  AND2X1 U16778 ( .IN1(n16217), .IN2(n5805), .Q(n16216) );
  AND2X1 U16779 ( .IN1(n5425), .IN2(n16211), .Q(n16217) );
  AND2X1 U16780 ( .IN1(n16218), .IN2(g5481), .Q(n16215) );
  OR2X1 U16781 ( .IN1(n10887), .IN2(n16219), .Q(n16218) );
  AND2X1 U16782 ( .IN1(n16220), .IN2(g5475), .Q(n16219) );
  AND2X1 U16783 ( .IN1(n16212), .IN2(g5485), .Q(n16213) );
  OR2X1 U16784 ( .IN1(n16221), .IN2(n16222), .Q(g29288) );
  AND2X1 U16785 ( .IN1(n16223), .IN2(g5475), .Q(n16222) );
  AND2X1 U16786 ( .IN1(n16212), .IN2(g5481), .Q(n16221) );
  OR2X1 U16787 ( .IN1(n16224), .IN2(n16225), .Q(g29287) );
  OR2X1 U16788 ( .IN1(n16226), .IN2(n16227), .Q(n16225) );
  AND2X1 U16789 ( .IN1(n16228), .IN2(n5744), .Q(n16227) );
  AND2X1 U16790 ( .IN1(n16211), .IN2(g5467), .Q(n16228) );
  AND2X1 U16791 ( .IN1(n10809), .IN2(n16220), .Q(n16211) );
  AND2X1 U16792 ( .IN1(n16229), .IN2(g5462), .Q(n16226) );
  OR2X1 U16793 ( .IN1(n10887), .IN2(n16230), .Q(n16229) );
  AND2X1 U16794 ( .IN1(n10086), .IN2(n16220), .Q(n16230) );
  AND2X1 U16795 ( .IN1(n16212), .IN2(g5471), .Q(n16224) );
  INVX0 U16796 ( .INP(n16223), .ZN(n16212) );
  OR2X1 U16797 ( .IN1(n10887), .IN2(n16220), .Q(n16223) );
  AND2X1 U16798 ( .IN1(n13176), .IN2(n16231), .Q(n16220) );
  OR2X1 U16799 ( .IN1(n16232), .IN2(n16233), .Q(g29286) );
  AND2X1 U16800 ( .IN1(n16234), .IN2(n10798), .Q(n16233) );
  OR2X1 U16801 ( .IN1(n16235), .IN2(n16236), .Q(n16234) );
  AND2X1 U16802 ( .IN1(n16237), .IN2(n13176), .Q(n16236) );
  XNOR2X1 U16803 ( .IN1(n16238), .IN2(n16239), .Q(n16237) );
  OR2X1 U16804 ( .IN1(n16231), .IN2(n5744), .Q(n16238) );
  AND2X1 U16805 ( .IN1(n12124), .IN2(n16240), .Q(n16231) );
  AND2X1 U16806 ( .IN1(g5689), .IN2(g17604), .Q(n16240) );
  AND2X1 U16807 ( .IN1(n13180), .IN2(g5462), .Q(n16235) );
  AND2X1 U16808 ( .IN1(n10898), .IN2(g5467), .Q(n16232) );
  OR2X1 U16809 ( .IN1(n16241), .IN2(n16242), .Q(g29285) );
  OR2X1 U16810 ( .IN1(n16083), .IN2(n16243), .Q(n16242) );
  AND2X1 U16811 ( .IN1(n16244), .IN2(n15141), .Q(n16243) );
  AND2X1 U16812 ( .IN1(n16086), .IN2(g5156), .Q(n16244) );
  AND2X1 U16813 ( .IN1(n3765), .IN2(n16245), .Q(n16241) );
  OR2X1 U16814 ( .IN1(g32975), .IN2(n5734), .Q(n16245) );
  OR2X1 U16815 ( .IN1(n16246), .IN2(n16247), .Q(g29284) );
  OR2X1 U16816 ( .IN1(n16248), .IN2(n16249), .Q(n16247) );
  AND2X1 U16817 ( .IN1(n5658), .IN2(n16250), .Q(n16249) );
  AND2X1 U16818 ( .IN1(n16251), .IN2(g5142), .Q(n16248) );
  AND2X1 U16819 ( .IN1(n10898), .IN2(g5138), .Q(n16246) );
  OR2X1 U16820 ( .IN1(n16252), .IN2(n16253), .Q(g29283) );
  OR2X1 U16821 ( .IN1(n16254), .IN2(n16255), .Q(n16253) );
  AND2X1 U16822 ( .IN1(n16256), .IN2(n5807), .Q(n16255) );
  AND2X1 U16823 ( .IN1(n16250), .IN2(n10577), .Q(n16256) );
  AND2X1 U16824 ( .IN1(n16257), .IN2(g5134), .Q(n16254) );
  OR2X1 U16825 ( .IN1(n10887), .IN2(n16258), .Q(n16257) );
  AND2X1 U16826 ( .IN1(test_so96), .IN2(n16259), .Q(n16258) );
  AND2X1 U16827 ( .IN1(n16251), .IN2(g5138), .Q(n16252) );
  OR2X1 U16828 ( .IN1(n16260), .IN2(n16261), .Q(g29282) );
  AND2X1 U16829 ( .IN1(test_so96), .IN2(n16262), .Q(n16261) );
  AND2X1 U16830 ( .IN1(n16251), .IN2(g5134), .Q(n16260) );
  INVX0 U16831 ( .INP(n16262), .ZN(n16251) );
  OR2X1 U16832 ( .IN1(n10888), .IN2(n16259), .Q(n16262) );
  OR2X1 U16833 ( .IN1(n16263), .IN2(n16264), .Q(g29281) );
  OR2X1 U16834 ( .IN1(n16265), .IN2(n16266), .Q(n16264) );
  AND2X1 U16835 ( .IN1(n16267), .IN2(n5743), .Q(n16266) );
  AND2X1 U16836 ( .IN1(n16250), .IN2(g5120), .Q(n16267) );
  AND2X1 U16837 ( .IN1(n10827), .IN2(n16259), .Q(n16250) );
  AND2X1 U16838 ( .IN1(n16268), .IN2(g5115), .Q(n16265) );
  OR2X1 U16839 ( .IN1(n10888), .IN2(n16269), .Q(n16268) );
  AND2X1 U16840 ( .IN1(n10085), .IN2(n16259), .Q(n16269) );
  INVX0 U16841 ( .INP(n16270), .ZN(n16263) );
  OR2X1 U16842 ( .IN1(n14619), .IN2(n16259), .Q(n16270) );
  AND2X1 U16843 ( .IN1(g33959), .IN2(n16271), .Q(n16259) );
  OR2X1 U16844 ( .IN1(n10525), .IN2(n10877), .Q(n14619) );
  OR2X1 U16845 ( .IN1(n16272), .IN2(n16273), .Q(g29280) );
  AND2X1 U16846 ( .IN1(n16274), .IN2(n10806), .Q(n16273) );
  OR2X1 U16847 ( .IN1(n16275), .IN2(n16276), .Q(n16274) );
  AND2X1 U16848 ( .IN1(n16277), .IN2(g33959), .Q(n16276) );
  XNOR2X1 U16849 ( .IN1(n16278), .IN2(n16279), .Q(n16277) );
  OR2X1 U16850 ( .IN1(n5743), .IN2(n16271), .Q(n16279) );
  AND2X1 U16851 ( .IN1(test_so10), .IN2(n16280), .Q(n16271) );
  AND2X1 U16852 ( .IN1(g17577), .IN2(g31860), .Q(n16280) );
  AND2X1 U16853 ( .IN1(n10535), .IN2(g5115), .Q(n16275) );
  AND2X1 U16854 ( .IN1(n10898), .IN2(g5120), .Q(n16272) );
  OR2X1 U16855 ( .IN1(n16281), .IN2(g29279), .Q(g29278) );
  AND2X1 U16856 ( .IN1(n10898), .IN2(g4572), .Q(n16281) );
  OR2X1 U16857 ( .IN1(n16282), .IN2(g29277), .Q(g29276) );
  AND2X1 U16858 ( .IN1(test_so100), .IN2(n10895), .Q(n16282) );
  OR2X1 U16859 ( .IN1(n16283), .IN2(n16284), .Q(g29275) );
  AND2X1 U16860 ( .IN1(test_so11), .IN2(n10894), .Q(n16284) );
  AND2X1 U16861 ( .IN1(n16285), .IN2(n15280), .Q(n16283) );
  XNOR2X1 U16862 ( .IN1(n14545), .IN2(g4087), .Q(n16285) );
  OR2X1 U16863 ( .IN1(n16286), .IN2(n10554), .Q(n14545) );
  OR2X1 U16864 ( .IN1(n16287), .IN2(n16288), .Q(g29274) );
  OR2X1 U16865 ( .IN1(n16083), .IN2(n16289), .Q(n16288) );
  AND2X1 U16866 ( .IN1(n16290), .IN2(n15287), .Q(n16289) );
  AND2X1 U16867 ( .IN1(n16086), .IN2(g3849), .Q(n16290) );
  AND2X1 U16868 ( .IN1(n3765), .IN2(n16291), .Q(n16287) );
  OR2X1 U16869 ( .IN1(n13080), .IN2(n5735), .Q(n16291) );
  OR2X1 U16870 ( .IN1(n16292), .IN2(n16293), .Q(g29273) );
  OR2X1 U16871 ( .IN1(n16294), .IN2(n16295), .Q(n16293) );
  AND2X1 U16872 ( .IN1(n5662), .IN2(n16296), .Q(n16295) );
  AND2X1 U16873 ( .IN1(n16297), .IN2(g3835), .Q(n16294) );
  AND2X1 U16874 ( .IN1(n10899), .IN2(g3831), .Q(n16292) );
  OR2X1 U16875 ( .IN1(n16298), .IN2(n16299), .Q(g29272) );
  OR2X1 U16876 ( .IN1(n16300), .IN2(n16301), .Q(n16299) );
  AND2X1 U16877 ( .IN1(n16302), .IN2(n5808), .Q(n16301) );
  AND2X1 U16878 ( .IN1(n5428), .IN2(n16296), .Q(n16302) );
  AND2X1 U16879 ( .IN1(n16303), .IN2(g3827), .Q(n16300) );
  OR2X1 U16880 ( .IN1(n10888), .IN2(n16304), .Q(n16303) );
  AND2X1 U16881 ( .IN1(n16305), .IN2(g3821), .Q(n16304) );
  AND2X1 U16882 ( .IN1(n16297), .IN2(g3831), .Q(n16298) );
  OR2X1 U16883 ( .IN1(n16306), .IN2(n16307), .Q(g29271) );
  AND2X1 U16884 ( .IN1(n16308), .IN2(g3821), .Q(n16307) );
  AND2X1 U16885 ( .IN1(n16297), .IN2(g3827), .Q(n16306) );
  INVX0 U16886 ( .INP(n16308), .ZN(n16297) );
  OR2X1 U16887 ( .IN1(n10888), .IN2(n16305), .Q(n16308) );
  OR2X1 U16888 ( .IN1(n16309), .IN2(n16310), .Q(g29270) );
  OR2X1 U16889 ( .IN1(n16311), .IN2(n16312), .Q(n16310) );
  AND2X1 U16890 ( .IN1(n16313), .IN2(n5745), .Q(n16312) );
  AND2X1 U16891 ( .IN1(n16296), .IN2(g3813), .Q(n16313) );
  AND2X1 U16892 ( .IN1(n10825), .IN2(n16305), .Q(n16296) );
  AND2X1 U16893 ( .IN1(n16314), .IN2(g3808), .Q(n16311) );
  OR2X1 U16894 ( .IN1(n10888), .IN2(n16315), .Q(n16314) );
  AND2X1 U16895 ( .IN1(n10087), .IN2(n16305), .Q(n16315) );
  INVX0 U16896 ( .INP(n16316), .ZN(n16309) );
  OR2X1 U16897 ( .IN1(n11709), .IN2(n16305), .Q(n16316) );
  AND2X1 U16898 ( .IN1(n13224), .IN2(n16317), .Q(n16305) );
  OR2X1 U16899 ( .IN1(n10502), .IN2(n10875), .Q(n11709) );
  OR2X1 U16900 ( .IN1(n16318), .IN2(n16319), .Q(g29269) );
  AND2X1 U16901 ( .IN1(n16320), .IN2(n10804), .Q(n16319) );
  OR2X1 U16902 ( .IN1(n16321), .IN2(n16322), .Q(n16320) );
  AND2X1 U16903 ( .IN1(n16323), .IN2(n13224), .Q(n16322) );
  XNOR2X1 U16904 ( .IN1(n16324), .IN2(n16325), .Q(n16323) );
  OR2X1 U16905 ( .IN1(n16317), .IN2(n5745), .Q(n16324) );
  AND2X1 U16906 ( .IN1(n12118), .IN2(n16326), .Q(n16317) );
  AND2X1 U16907 ( .IN1(g4040), .IN2(g16693), .Q(n16326) );
  AND2X1 U16908 ( .IN1(n13228), .IN2(g3808), .Q(n16321) );
  AND2X1 U16909 ( .IN1(n10897), .IN2(g3813), .Q(n16318) );
  OR2X1 U16910 ( .IN1(n16327), .IN2(n16328), .Q(g29268) );
  OR2X1 U16911 ( .IN1(n16083), .IN2(n16329), .Q(n16328) );
  AND2X1 U16912 ( .IN1(n16330), .IN2(n15412), .Q(n16329) );
  AND2X1 U16913 ( .IN1(n16086), .IN2(g3498), .Q(n16330) );
  AND2X1 U16914 ( .IN1(n3765), .IN2(n16331), .Q(n16327) );
  OR2X1 U16915 ( .IN1(n13079), .IN2(n5740), .Q(n16331) );
  OR2X1 U16916 ( .IN1(n16332), .IN2(n16333), .Q(g29267) );
  OR2X1 U16917 ( .IN1(n16334), .IN2(n16335), .Q(n16333) );
  AND2X1 U16918 ( .IN1(n5668), .IN2(n16336), .Q(n16335) );
  AND2X1 U16919 ( .IN1(n16337), .IN2(g3484), .Q(n16334) );
  AND2X1 U16920 ( .IN1(n10898), .IN2(g3480), .Q(n16332) );
  OR2X1 U16921 ( .IN1(n16338), .IN2(n16339), .Q(g29266) );
  OR2X1 U16922 ( .IN1(n16340), .IN2(n16341), .Q(n16339) );
  AND2X1 U16923 ( .IN1(n16342), .IN2(n5786), .Q(n16341) );
  AND2X1 U16924 ( .IN1(n5424), .IN2(n16336), .Q(n16342) );
  AND2X1 U16925 ( .IN1(n16343), .IN2(g3476), .Q(n16340) );
  OR2X1 U16926 ( .IN1(n10888), .IN2(n16344), .Q(n16343) );
  AND2X1 U16927 ( .IN1(n16345), .IN2(g3470), .Q(n16344) );
  AND2X1 U16928 ( .IN1(n16337), .IN2(g3480), .Q(n16338) );
  OR2X1 U16929 ( .IN1(n16346), .IN2(n16347), .Q(g29265) );
  AND2X1 U16930 ( .IN1(n16348), .IN2(g3470), .Q(n16347) );
  AND2X1 U16931 ( .IN1(n16337), .IN2(g3476), .Q(n16346) );
  INVX0 U16932 ( .INP(n16348), .ZN(n16337) );
  OR2X1 U16933 ( .IN1(n10888), .IN2(n16345), .Q(n16348) );
  OR2X1 U16934 ( .IN1(n16349), .IN2(n16350), .Q(g29264) );
  OR2X1 U16935 ( .IN1(n16351), .IN2(n16352), .Q(n16350) );
  AND2X1 U16936 ( .IN1(n16353), .IN2(n10573), .Q(n16352) );
  AND2X1 U16937 ( .IN1(n16336), .IN2(g3462), .Q(n16353) );
  AND2X1 U16938 ( .IN1(n10825), .IN2(n16345), .Q(n16336) );
  AND2X1 U16939 ( .IN1(test_so4), .IN2(n16354), .Q(n16351) );
  OR2X1 U16940 ( .IN1(n10888), .IN2(n16355), .Q(n16354) );
  AND2X1 U16941 ( .IN1(n10088), .IN2(n16345), .Q(n16355) );
  INVX0 U16942 ( .INP(n16356), .ZN(n16349) );
  OR2X1 U16943 ( .IN1(n14613), .IN2(n16345), .Q(n16356) );
  AND2X1 U16944 ( .IN1(n13245), .IN2(n16357), .Q(n16345) );
  OR2X1 U16945 ( .IN1(n10503), .IN2(n10877), .Q(n14613) );
  OR2X1 U16946 ( .IN1(n16358), .IN2(n16359), .Q(g29263) );
  OR2X1 U16947 ( .IN1(n16360), .IN2(n16361), .Q(n16359) );
  AND2X1 U16948 ( .IN1(test_so4), .IN2(n13258), .Q(n16361) );
  AND2X1 U16949 ( .IN1(n13255), .IN2(n16362), .Q(n16360) );
  XNOR2X1 U16950 ( .IN1(n16363), .IN2(n16364), .Q(n16362) );
  OR2X1 U16951 ( .IN1(n16357), .IN2(n10573), .Q(n16363) );
  AND2X1 U16952 ( .IN1(n12131), .IN2(n16365), .Q(n16357) );
  AND2X1 U16953 ( .IN1(g3689), .IN2(g16656), .Q(n16365) );
  AND2X1 U16954 ( .IN1(n10897), .IN2(g3462), .Q(n16358) );
  OR2X1 U16955 ( .IN1(n16366), .IN2(n16367), .Q(g29262) );
  OR2X1 U16956 ( .IN1(n16083), .IN2(n16368), .Q(n16367) );
  AND2X1 U16957 ( .IN1(n16369), .IN2(n15537), .Q(n16368) );
  AND2X1 U16958 ( .IN1(n16086), .IN2(g3147), .Q(n16369) );
  AND2X1 U16959 ( .IN1(n16086), .IN2(n3765), .Q(n16083) );
  INVX0 U16960 ( .INP(n4210), .ZN(n16086) );
  OR2X1 U16961 ( .IN1(n5380), .IN2(g4284), .Q(n4210) );
  AND2X1 U16962 ( .IN1(n3765), .IN2(n16370), .Q(n16366) );
  OR2X1 U16963 ( .IN1(n13082), .IN2(n5738), .Q(n16370) );
  OR2X1 U16964 ( .IN1(n16371), .IN2(n16372), .Q(g29261) );
  OR2X1 U16965 ( .IN1(n16373), .IN2(n16374), .Q(n16372) );
  AND2X1 U16966 ( .IN1(n5661), .IN2(n16375), .Q(n16374) );
  AND2X1 U16967 ( .IN1(n16376), .IN2(g3133), .Q(n16373) );
  AND2X1 U16968 ( .IN1(n10897), .IN2(g3129), .Q(n16371) );
  OR2X1 U16969 ( .IN1(n16377), .IN2(n16378), .Q(g29260) );
  OR2X1 U16970 ( .IN1(n16379), .IN2(n16380), .Q(n16378) );
  AND2X1 U16971 ( .IN1(n16381), .IN2(n5781), .Q(n16380) );
  AND2X1 U16972 ( .IN1(n5423), .IN2(n16375), .Q(n16381) );
  AND2X1 U16973 ( .IN1(n16382), .IN2(g3125), .Q(n16379) );
  OR2X1 U16974 ( .IN1(n10889), .IN2(n16383), .Q(n16382) );
  AND2X1 U16975 ( .IN1(n16384), .IN2(g3119), .Q(n16383) );
  AND2X1 U16976 ( .IN1(n16376), .IN2(g3129), .Q(n16377) );
  OR2X1 U16977 ( .IN1(n16385), .IN2(n16386), .Q(g29259) );
  AND2X1 U16978 ( .IN1(n16387), .IN2(g3119), .Q(n16386) );
  AND2X1 U16979 ( .IN1(n16376), .IN2(g3125), .Q(n16385) );
  INVX0 U16980 ( .INP(n16387), .ZN(n16376) );
  OR2X1 U16981 ( .IN1(n10889), .IN2(n16384), .Q(n16387) );
  OR2X1 U16982 ( .IN1(n16388), .IN2(n16389), .Q(g29258) );
  OR2X1 U16983 ( .IN1(n16390), .IN2(n16391), .Q(n16389) );
  AND2X1 U16984 ( .IN1(n16392), .IN2(n5742), .Q(n16391) );
  AND2X1 U16985 ( .IN1(n16375), .IN2(g3111), .Q(n16392) );
  AND2X1 U16986 ( .IN1(n10825), .IN2(n16384), .Q(n16375) );
  AND2X1 U16987 ( .IN1(n16393), .IN2(g3106), .Q(n16390) );
  OR2X1 U16988 ( .IN1(n10889), .IN2(n16394), .Q(n16393) );
  AND2X1 U16989 ( .IN1(n10084), .IN2(n16384), .Q(n16394) );
  INVX0 U16990 ( .INP(n16395), .ZN(n16388) );
  OR2X1 U16991 ( .IN1(n14612), .IN2(n16384), .Q(n16395) );
  AND2X1 U16992 ( .IN1(n13270), .IN2(n16396), .Q(n16384) );
  OR2X1 U16993 ( .IN1(n10485), .IN2(n10876), .Q(n14612) );
  OR2X1 U16994 ( .IN1(n16397), .IN2(n16398), .Q(g29257) );
  AND2X1 U16995 ( .IN1(n16399), .IN2(n10801), .Q(n16398) );
  OR2X1 U16996 ( .IN1(n16400), .IN2(n16401), .Q(n16399) );
  AND2X1 U16997 ( .IN1(n16402), .IN2(n13270), .Q(n16401) );
  XNOR2X1 U16998 ( .IN1(n16403), .IN2(n16404), .Q(n16402) );
  OR2X1 U16999 ( .IN1(n16396), .IN2(n5742), .Q(n16403) );
  AND2X1 U17000 ( .IN1(n12123), .IN2(n16405), .Q(n16396) );
  AND2X1 U17001 ( .IN1(g3338), .IN2(g16624), .Q(n16405) );
  AND2X1 U17002 ( .IN1(n13268), .IN2(g3106), .Q(n16400) );
  AND2X1 U17003 ( .IN1(n10910), .IN2(g3111), .Q(n16397) );
  OR2X1 U17004 ( .IN1(n16406), .IN2(n16407), .Q(g29256) );
  OR2X1 U17005 ( .IN1(n2787), .IN2(n16408), .Q(n16407) );
  INVX0 U17006 ( .INP(n16409), .ZN(n16408) );
  OR2X1 U17007 ( .IN1(g2735), .IN2(n15711), .Q(n16409) );
  OR2X1 U17008 ( .IN1(n16410), .IN2(n16411), .Q(n16406) );
  AND2X1 U17009 ( .IN1(n10910), .IN2(g2729), .Q(n16411) );
  AND2X1 U17010 ( .IN1(n16412), .IN2(n10801), .Q(n16410) );
  AND2X1 U17011 ( .IN1(n15711), .IN2(g2735), .Q(n16412) );
  OR2X1 U17012 ( .IN1(n16413), .IN2(n12042), .Q(n15711) );
  OR2X1 U17013 ( .IN1(n10520), .IN2(n5301), .Q(n12042) );
  OR2X1 U17014 ( .IN1(n16414), .IN2(n16415), .Q(g29255) );
  AND2X1 U17015 ( .IN1(n16416), .IN2(g2652), .Q(n16415) );
  OR2X1 U17016 ( .IN1(n16417), .IN2(n14112), .Q(n16416) );
  AND2X1 U17017 ( .IN1(n4379), .IN2(n10801), .Q(n16417) );
  AND2X1 U17018 ( .IN1(n16418), .IN2(g2638), .Q(n16414) );
  OR2X1 U17019 ( .IN1(n10889), .IN2(n16419), .Q(n16418) );
  AND2X1 U17020 ( .IN1(n14120), .IN2(n11107), .Q(n16419) );
  OR2X1 U17021 ( .IN1(n10539), .IN2(n10202), .Q(n11107) );
  OR2X1 U17022 ( .IN1(n16420), .IN2(n16421), .Q(g29254) );
  OR2X1 U17023 ( .IN1(n16422), .IN2(n16423), .Q(n16421) );
  OR2X1 U17024 ( .IN1(n16424), .IN2(n16425), .Q(n16423) );
  AND2X1 U17025 ( .IN1(n16426), .IN2(n10801), .Q(n16425) );
  AND2X1 U17026 ( .IN1(n15742), .IN2(g2583), .Q(n16426) );
  INVX0 U17027 ( .INP(n15744), .ZN(n15742) );
  OR2X1 U17028 ( .IN1(g2619), .IN2(n16427), .Q(n15744) );
  OR2X1 U17029 ( .IN1(n10468), .IN2(n16428), .Q(n16427) );
  AND2X1 U17030 ( .IN1(n10910), .IN2(g2619), .Q(n16424) );
  AND2X1 U17031 ( .IN1(n14112), .IN2(g2638), .Q(n16422) );
  INVX0 U17032 ( .INP(n14129), .ZN(n14112) );
  OR2X1 U17033 ( .IN1(n10889), .IN2(n14120), .Q(n14129) );
  OR2X1 U17034 ( .IN1(n16429), .IN2(n16430), .Q(n16420) );
  AND2X1 U17035 ( .IN1(n3517), .IN2(n16431), .Q(n16430) );
  OR2X1 U17036 ( .IN1(n16432), .IN2(n16433), .Q(n16431) );
  OR2X1 U17037 ( .IN1(n16434), .IN2(n16435), .Q(n16433) );
  AND2X1 U17038 ( .IN1(n10468), .IN2(n16436), .Q(n16435) );
  OR2X1 U17039 ( .IN1(n16437), .IN2(n16438), .Q(n16436) );
  AND2X1 U17040 ( .IN1(g2619), .IN2(g2571), .Q(n16438) );
  AND2X1 U17041 ( .IN1(test_so61), .IN2(g2587), .Q(n16437) );
  AND2X1 U17042 ( .IN1(n16439), .IN2(test_so66), .Q(n16434) );
  AND2X1 U17043 ( .IN1(n5508), .IN2(n5372), .Q(n16439) );
  AND2X1 U17044 ( .IN1(n10539), .IN2(g2563), .Q(n16432) );
  AND2X1 U17045 ( .IN1(g2610), .IN2(n5372), .Q(n10539) );
  AND2X1 U17046 ( .IN1(n10824), .IN2(n14120), .Q(n3517) );
  AND2X1 U17047 ( .IN1(n15717), .IN2(g2567), .Q(n16429) );
  AND2X1 U17048 ( .IN1(n10824), .IN2(n15720), .Q(n15717) );
  AND2X1 U17049 ( .IN1(n14120), .IN2(n16440), .Q(n15720) );
  AND2X1 U17050 ( .IN1(g2619), .IN2(g2587), .Q(n16440) );
  INVX0 U17051 ( .INP(n16428), .ZN(n14120) );
  OR2X1 U17052 ( .IN1(n16413), .IN2(n16441), .Q(n16428) );
  OR2X1 U17053 ( .IN1(n16442), .IN2(n16443), .Q(n16441) );
  AND2X1 U17054 ( .IN1(n12071), .IN2(g2819), .Q(n16443) );
  OR2X1 U17055 ( .IN1(n16444), .IN2(n16445), .Q(g29253) );
  AND2X1 U17056 ( .IN1(n16446), .IN2(g2504), .Q(n16445) );
  OR2X1 U17057 ( .IN1(n10889), .IN2(n16447), .Q(n16446) );
  AND2X1 U17058 ( .IN1(n14154), .IN2(n11106), .Q(n16447) );
  OR2X1 U17059 ( .IN1(n10546), .IN2(n10200), .Q(n11106) );
  AND2X1 U17060 ( .IN1(n16448), .IN2(g2518), .Q(n16444) );
  OR2X1 U17061 ( .IN1(n16449), .IN2(n14144), .Q(n16448) );
  AND2X1 U17062 ( .IN1(n4391), .IN2(n10798), .Q(n16449) );
  OR2X1 U17063 ( .IN1(n16450), .IN2(n16451), .Q(g29252) );
  OR2X1 U17064 ( .IN1(n16452), .IN2(n16453), .Q(n16451) );
  OR2X1 U17065 ( .IN1(n16454), .IN2(n16455), .Q(n16453) );
  AND2X1 U17066 ( .IN1(n16456), .IN2(n10798), .Q(n16455) );
  AND2X1 U17067 ( .IN1(n15775), .IN2(g2449), .Q(n16456) );
  INVX0 U17068 ( .INP(n15777), .ZN(n15775) );
  OR2X1 U17069 ( .IN1(g2485), .IN2(n16457), .Q(n15777) );
  OR2X1 U17070 ( .IN1(n10470), .IN2(n16458), .Q(n16457) );
  AND2X1 U17071 ( .IN1(n10910), .IN2(g2485), .Q(n16454) );
  AND2X1 U17072 ( .IN1(n14144), .IN2(g2504), .Q(n16452) );
  INVX0 U17073 ( .INP(n14163), .ZN(n14144) );
  OR2X1 U17074 ( .IN1(n10890), .IN2(n14154), .Q(n14163) );
  OR2X1 U17075 ( .IN1(n16459), .IN2(n16460), .Q(n16450) );
  AND2X1 U17076 ( .IN1(n3536), .IN2(n16461), .Q(n16460) );
  OR2X1 U17077 ( .IN1(n16462), .IN2(n16463), .Q(n16461) );
  OR2X1 U17078 ( .IN1(n16464), .IN2(n16465), .Q(n16463) );
  AND2X1 U17079 ( .IN1(n10470), .IN2(n16466), .Q(n16465) );
  OR2X1 U17080 ( .IN1(n16467), .IN2(n16468), .Q(n16466) );
  AND2X1 U17081 ( .IN1(g2485), .IN2(g2437), .Q(n16468) );
  AND2X1 U17082 ( .IN1(g2453), .IN2(n9274), .Q(n16467) );
  AND2X1 U17083 ( .IN1(n16469), .IN2(n5509), .Q(n16464) );
  AND2X1 U17084 ( .IN1(n5373), .IN2(g2441), .Q(n16469) );
  AND2X1 U17085 ( .IN1(n10546), .IN2(g2429), .Q(n16462) );
  AND2X1 U17086 ( .IN1(g2476), .IN2(n5373), .Q(n10546) );
  AND2X1 U17087 ( .IN1(n10823), .IN2(n14154), .Q(n3536) );
  AND2X1 U17088 ( .IN1(n15750), .IN2(g2433), .Q(n16459) );
  AND2X1 U17089 ( .IN1(n10823), .IN2(n15753), .Q(n15750) );
  AND2X1 U17090 ( .IN1(n14154), .IN2(n16470), .Q(n15753) );
  AND2X1 U17091 ( .IN1(g2485), .IN2(g2453), .Q(n16470) );
  INVX0 U17092 ( .INP(n16458), .ZN(n14154) );
  OR2X1 U17093 ( .IN1(n16471), .IN2(n16472), .Q(n16458) );
  OR2X1 U17094 ( .IN1(n16442), .IN2(n16473), .Q(n16472) );
  AND2X1 U17095 ( .IN1(n12071), .IN2(g2815), .Q(n16473) );
  OR2X1 U17096 ( .IN1(n16474), .IN2(n16475), .Q(g29251) );
  AND2X1 U17097 ( .IN1(n16476), .IN2(g2370), .Q(n16475) );
  OR2X1 U17098 ( .IN1(n10890), .IN2(n16477), .Q(n16476) );
  AND2X1 U17099 ( .IN1(n14187), .IN2(n11105), .Q(n16477) );
  OR2X1 U17100 ( .IN1(n10541), .IN2(n10194), .Q(n11105) );
  AND2X1 U17101 ( .IN1(n16478), .IN2(g2384), .Q(n16474) );
  OR2X1 U17102 ( .IN1(n16479), .IN2(n14178), .Q(n16478) );
  AND2X1 U17103 ( .IN1(n4402), .IN2(n10799), .Q(n16479) );
  OR2X1 U17104 ( .IN1(n16480), .IN2(n16481), .Q(g29250) );
  OR2X1 U17105 ( .IN1(n16482), .IN2(n16483), .Q(n16481) );
  OR2X1 U17106 ( .IN1(n16484), .IN2(n16485), .Q(n16483) );
  AND2X1 U17107 ( .IN1(n16486), .IN2(n10799), .Q(n16485) );
  AND2X1 U17108 ( .IN1(n15808), .IN2(g2315), .Q(n16486) );
  INVX0 U17109 ( .INP(n15810), .ZN(n15808) );
  OR2X1 U17110 ( .IN1(g2351), .IN2(n16487), .Q(n15810) );
  OR2X1 U17111 ( .IN1(n10555), .IN2(n16488), .Q(n16487) );
  AND2X1 U17112 ( .IN1(n10910), .IN2(g2351), .Q(n16484) );
  AND2X1 U17113 ( .IN1(n14178), .IN2(g2370), .Q(n16482) );
  INVX0 U17114 ( .INP(n14196), .ZN(n14178) );
  OR2X1 U17115 ( .IN1(n10890), .IN2(n14187), .Q(n14196) );
  OR2X1 U17116 ( .IN1(n16489), .IN2(n16490), .Q(n16480) );
  AND2X1 U17117 ( .IN1(n3555), .IN2(n16491), .Q(n16490) );
  OR2X1 U17118 ( .IN1(n16492), .IN2(n16493), .Q(n16491) );
  OR2X1 U17119 ( .IN1(n16494), .IN2(n16495), .Q(n16493) );
  AND2X1 U17120 ( .IN1(n16496), .IN2(n10555), .Q(n16495) );
  OR2X1 U17121 ( .IN1(n16497), .IN2(n16498), .Q(n16496) );
  AND2X1 U17122 ( .IN1(g2351), .IN2(g2303), .Q(n16498) );
  AND2X1 U17123 ( .IN1(g2319), .IN2(n9314), .Q(n16497) );
  AND2X1 U17124 ( .IN1(n16499), .IN2(n5511), .Q(n16494) );
  AND2X1 U17125 ( .IN1(n5375), .IN2(g2307), .Q(n16499) );
  AND2X1 U17126 ( .IN1(n10541), .IN2(g2295), .Q(n16492) );
  AND2X1 U17127 ( .IN1(n5375), .IN2(test_so21), .Q(n10541) );
  AND2X1 U17128 ( .IN1(n10822), .IN2(n14187), .Q(n3555) );
  AND2X1 U17129 ( .IN1(n15783), .IN2(g2299), .Q(n16489) );
  AND2X1 U17130 ( .IN1(n10822), .IN2(n15786), .Q(n15783) );
  AND2X1 U17131 ( .IN1(n14187), .IN2(n16500), .Q(n15786) );
  AND2X1 U17132 ( .IN1(g2351), .IN2(g2319), .Q(n16500) );
  INVX0 U17133 ( .INP(n16488), .ZN(n14187) );
  OR2X1 U17134 ( .IN1(n16501), .IN2(n16502), .Q(n16488) );
  AND2X1 U17135 ( .IN1(n12071), .IN2(g2807), .Q(n16501) );
  OR2X1 U17136 ( .IN1(n16503), .IN2(n16504), .Q(g29249) );
  AND2X1 U17137 ( .IN1(n16505), .IN2(g2236), .Q(n16504) );
  OR2X1 U17138 ( .IN1(n10890), .IN2(n16506), .Q(n16505) );
  AND2X1 U17139 ( .IN1(n14220), .IN2(n11104), .Q(n16506) );
  OR2X1 U17140 ( .IN1(n10547), .IN2(n10190), .Q(n11104) );
  AND2X1 U17141 ( .IN1(n16507), .IN2(g2250), .Q(n16503) );
  OR2X1 U17142 ( .IN1(n16508), .IN2(n14211), .Q(n16507) );
  AND2X1 U17143 ( .IN1(n4414), .IN2(n10799), .Q(n16508) );
  OR2X1 U17144 ( .IN1(n16509), .IN2(n16510), .Q(g29248) );
  OR2X1 U17145 ( .IN1(n16511), .IN2(n16512), .Q(n16510) );
  OR2X1 U17146 ( .IN1(n16513), .IN2(n16514), .Q(n16512) );
  AND2X1 U17147 ( .IN1(n16515), .IN2(n10799), .Q(n16514) );
  AND2X1 U17148 ( .IN1(n15841), .IN2(g2181), .Q(n16515) );
  INVX0 U17149 ( .INP(n15843), .ZN(n15841) );
  OR2X1 U17150 ( .IN1(g2217), .IN2(n16516), .Q(n15843) );
  OR2X1 U17151 ( .IN1(n10471), .IN2(n16517), .Q(n16516) );
  AND2X1 U17152 ( .IN1(n10909), .IN2(g2217), .Q(n16513) );
  AND2X1 U17153 ( .IN1(n14211), .IN2(g2236), .Q(n16511) );
  INVX0 U17154 ( .INP(n14229), .ZN(n14211) );
  OR2X1 U17155 ( .IN1(n10891), .IN2(n14220), .Q(n14229) );
  OR2X1 U17156 ( .IN1(n16518), .IN2(n16519), .Q(n16509) );
  AND2X1 U17157 ( .IN1(n3574), .IN2(n16520), .Q(n16519) );
  OR2X1 U17158 ( .IN1(n16521), .IN2(n16522), .Q(n16520) );
  OR2X1 U17159 ( .IN1(n16523), .IN2(n16524), .Q(n16522) );
  AND2X1 U17160 ( .IN1(n10471), .IN2(n16525), .Q(n16524) );
  OR2X1 U17161 ( .IN1(n16526), .IN2(n16527), .Q(n16525) );
  AND2X1 U17162 ( .IN1(g2217), .IN2(g2169), .Q(n16527) );
  AND2X1 U17163 ( .IN1(g2185), .IN2(n9352), .Q(n16526) );
  AND2X1 U17164 ( .IN1(n16528), .IN2(n5512), .Q(n16523) );
  AND2X1 U17165 ( .IN1(n5376), .IN2(g2173), .Q(n16528) );
  AND2X1 U17166 ( .IN1(n10547), .IN2(g2161), .Q(n16521) );
  AND2X1 U17167 ( .IN1(g2208), .IN2(n5376), .Q(n10547) );
  AND2X1 U17168 ( .IN1(n10822), .IN2(n14220), .Q(n3574) );
  AND2X1 U17169 ( .IN1(n15816), .IN2(g2165), .Q(n16518) );
  AND2X1 U17170 ( .IN1(n10822), .IN2(n15819), .Q(n15816) );
  AND2X1 U17171 ( .IN1(n14220), .IN2(n16529), .Q(n15819) );
  AND2X1 U17172 ( .IN1(g2217), .IN2(g2185), .Q(n16529) );
  INVX0 U17173 ( .INP(n16517), .ZN(n14220) );
  OR2X1 U17174 ( .IN1(n15707), .IN2(n16530), .Q(n16517) );
  OR2X1 U17175 ( .IN1(n16442), .IN2(n16531), .Q(n16530) );
  AND2X1 U17176 ( .IN1(n12071), .IN2(g2803), .Q(n16531) );
  OR2X1 U17177 ( .IN1(n16532), .IN2(n16533), .Q(g29247) );
  AND2X1 U17178 ( .IN1(test_so78), .IN2(n16534), .Q(n16533) );
  OR2X1 U17179 ( .IN1(n16535), .IN2(n14244), .Q(n16534) );
  AND2X1 U17180 ( .IN1(n4425), .IN2(n10800), .Q(n16535) );
  AND2X1 U17181 ( .IN1(n16536), .IN2(g2079), .Q(n16532) );
  OR2X1 U17182 ( .IN1(n10890), .IN2(n16537), .Q(n16536) );
  AND2X1 U17183 ( .IN1(n14254), .IN2(n11103), .Q(n16537) );
  INVX0 U17184 ( .INP(n16538), .ZN(n11103) );
  AND2X1 U17185 ( .IN1(n14270), .IN2(test_so78), .Q(n16538) );
  INVX0 U17186 ( .INP(n10549), .ZN(n14270) );
  OR2X1 U17187 ( .IN1(n16539), .IN2(n16540), .Q(g29246) );
  OR2X1 U17188 ( .IN1(n16541), .IN2(n16542), .Q(n16540) );
  OR2X1 U17189 ( .IN1(n16543), .IN2(n16544), .Q(n16542) );
  AND2X1 U17190 ( .IN1(n16545), .IN2(n10800), .Q(n16544) );
  AND2X1 U17191 ( .IN1(n15874), .IN2(g2024), .Q(n16545) );
  INVX0 U17192 ( .INP(n15876), .ZN(n15874) );
  OR2X1 U17193 ( .IN1(g2060), .IN2(n16546), .Q(n15876) );
  OR2X1 U17194 ( .IN1(n10472), .IN2(n16547), .Q(n16546) );
  AND2X1 U17195 ( .IN1(n10909), .IN2(g2060), .Q(n16543) );
  AND2X1 U17196 ( .IN1(n14244), .IN2(g2079), .Q(n16541) );
  INVX0 U17197 ( .INP(n14263), .ZN(n14244) );
  OR2X1 U17198 ( .IN1(n10891), .IN2(n14254), .Q(n14263) );
  OR2X1 U17199 ( .IN1(n16548), .IN2(n16549), .Q(n16539) );
  AND2X1 U17200 ( .IN1(n3593), .IN2(n16550), .Q(n16549) );
  OR2X1 U17201 ( .IN1(n16551), .IN2(n16552), .Q(n16550) );
  OR2X1 U17202 ( .IN1(n16553), .IN2(n16554), .Q(n16552) );
  AND2X1 U17203 ( .IN1(n10472), .IN2(n16555), .Q(n16554) );
  OR2X1 U17204 ( .IN1(n16556), .IN2(n16557), .Q(n16555) );
  AND2X1 U17205 ( .IN1(g2060), .IN2(g2012), .Q(n16557) );
  AND2X1 U17206 ( .IN1(g2028), .IN2(n9312), .Q(n16556) );
  AND2X1 U17207 ( .IN1(n16558), .IN2(n5507), .Q(n16553) );
  AND2X1 U17208 ( .IN1(n5371), .IN2(g2016), .Q(n16558) );
  AND2X1 U17209 ( .IN1(n10549), .IN2(g2004), .Q(n16551) );
  AND2X1 U17210 ( .IN1(g2051), .IN2(n5371), .Q(n10549) );
  AND2X1 U17211 ( .IN1(n10822), .IN2(n14254), .Q(n3593) );
  AND2X1 U17212 ( .IN1(n15849), .IN2(g2008), .Q(n16548) );
  AND2X1 U17213 ( .IN1(n10822), .IN2(n15852), .Q(n15849) );
  AND2X1 U17214 ( .IN1(n14254), .IN2(n16559), .Q(n15852) );
  AND2X1 U17215 ( .IN1(g2060), .IN2(g2028), .Q(n16559) );
  INVX0 U17216 ( .INP(n16547), .ZN(n14254) );
  OR2X1 U17217 ( .IN1(n16413), .IN2(n16560), .Q(n16547) );
  OR2X1 U17218 ( .IN1(n16442), .IN2(n16561), .Q(n16560) );
  AND2X1 U17219 ( .IN1(n12071), .IN2(g2787), .Q(n16561) );
  OR2X1 U17220 ( .IN1(n16562), .IN2(n16563), .Q(g29245) );
  AND2X1 U17221 ( .IN1(test_so53), .IN2(n16564), .Q(n16563) );
  OR2X1 U17222 ( .IN1(n10891), .IN2(n16565), .Q(n16564) );
  AND2X1 U17223 ( .IN1(n14288), .IN2(n11102), .Q(n16565) );
  OR2X1 U17224 ( .IN1(n10538), .IN2(n10199), .Q(n11102) );
  AND2X1 U17225 ( .IN1(n16566), .IN2(g1959), .Q(n16562) );
  OR2X1 U17226 ( .IN1(n16567), .IN2(n14278), .Q(n16566) );
  AND2X1 U17227 ( .IN1(n4436), .IN2(n10800), .Q(n16567) );
  OR2X1 U17228 ( .IN1(n16568), .IN2(n16569), .Q(g29244) );
  OR2X1 U17229 ( .IN1(n16570), .IN2(n16571), .Q(n16569) );
  OR2X1 U17230 ( .IN1(n16572), .IN2(n16573), .Q(n16571) );
  AND2X1 U17231 ( .IN1(n16574), .IN2(n10800), .Q(n16573) );
  AND2X1 U17232 ( .IN1(n15907), .IN2(g1890), .Q(n16574) );
  INVX0 U17233 ( .INP(n15909), .ZN(n15907) );
  OR2X1 U17234 ( .IN1(g1926), .IN2(n16575), .Q(n15909) );
  OR2X1 U17235 ( .IN1(n10469), .IN2(n16576), .Q(n16575) );
  AND2X1 U17236 ( .IN1(n10909), .IN2(g1926), .Q(n16572) );
  AND2X1 U17237 ( .IN1(n14278), .IN2(test_so53), .Q(n16570) );
  INVX0 U17238 ( .INP(n14297), .ZN(n14278) );
  OR2X1 U17239 ( .IN1(n10891), .IN2(n14288), .Q(n14297) );
  OR2X1 U17240 ( .IN1(n16577), .IN2(n16578), .Q(n16568) );
  AND2X1 U17241 ( .IN1(n3611), .IN2(n16579), .Q(n16578) );
  OR2X1 U17242 ( .IN1(n16580), .IN2(n16581), .Q(n16579) );
  OR2X1 U17243 ( .IN1(n16582), .IN2(n16583), .Q(n16581) );
  AND2X1 U17244 ( .IN1(n10469), .IN2(n16584), .Q(n16583) );
  OR2X1 U17245 ( .IN1(n16585), .IN2(n16586), .Q(n16584) );
  AND2X1 U17246 ( .IN1(g1926), .IN2(g1878), .Q(n16586) );
  AND2X1 U17247 ( .IN1(g1894), .IN2(n9280), .Q(n16585) );
  AND2X1 U17248 ( .IN1(n16587), .IN2(n5510), .Q(n16582) );
  AND2X1 U17249 ( .IN1(n5374), .IN2(g1882), .Q(n16587) );
  AND2X1 U17250 ( .IN1(n10538), .IN2(g1870), .Q(n16580) );
  AND2X1 U17251 ( .IN1(g1917), .IN2(n5374), .Q(n10538) );
  AND2X1 U17252 ( .IN1(n10821), .IN2(n14288), .Q(n3611) );
  AND2X1 U17253 ( .IN1(n15882), .IN2(g1874), .Q(n16577) );
  AND2X1 U17254 ( .IN1(n10821), .IN2(n15885), .Q(n15882) );
  AND2X1 U17255 ( .IN1(n14288), .IN2(n16588), .Q(n15885) );
  AND2X1 U17256 ( .IN1(g1926), .IN2(g1894), .Q(n16588) );
  INVX0 U17257 ( .INP(n16576), .ZN(n14288) );
  OR2X1 U17258 ( .IN1(n16471), .IN2(n16589), .Q(n16576) );
  OR2X1 U17259 ( .IN1(n16442), .IN2(n16590), .Q(n16589) );
  AND2X1 U17260 ( .IN1(n12071), .IN2(g2783), .Q(n16590) );
  INVX0 U17261 ( .INP(n15678), .ZN(n16471) );
  OR2X1 U17262 ( .IN1(n16591), .IN2(n16592), .Q(g29243) );
  AND2X1 U17263 ( .IN1(n16593), .IN2(g1811), .Q(n16592) );
  OR2X1 U17264 ( .IN1(n10891), .IN2(n16594), .Q(n16593) );
  AND2X1 U17265 ( .IN1(n14320), .IN2(n11101), .Q(n16594) );
  OR2X1 U17266 ( .IN1(n10544), .IN2(n10192), .Q(n11101) );
  AND2X1 U17267 ( .IN1(n16595), .IN2(g1825), .Q(n16591) );
  OR2X1 U17268 ( .IN1(n16596), .IN2(n14312), .Q(n16595) );
  AND2X1 U17269 ( .IN1(n4447), .IN2(n10801), .Q(n16596) );
  OR2X1 U17270 ( .IN1(n16597), .IN2(n16598), .Q(g29242) );
  OR2X1 U17271 ( .IN1(n16599), .IN2(n16600), .Q(n16598) );
  OR2X1 U17272 ( .IN1(n16601), .IN2(n16602), .Q(n16600) );
  AND2X1 U17273 ( .IN1(n16603), .IN2(n10801), .Q(n16602) );
  AND2X1 U17274 ( .IN1(n15940), .IN2(g1756), .Q(n16603) );
  INVX0 U17275 ( .INP(n15942), .ZN(n15940) );
  OR2X1 U17276 ( .IN1(g1792), .IN2(n16604), .Q(n15942) );
  OR2X1 U17277 ( .IN1(n5596), .IN2(n16605), .Q(n16604) );
  AND2X1 U17278 ( .IN1(n10909), .IN2(g1792), .Q(n16601) );
  AND2X1 U17279 ( .IN1(n14312), .IN2(g1811), .Q(n16599) );
  INVX0 U17280 ( .INP(n14329), .ZN(n14312) );
  OR2X1 U17281 ( .IN1(n10891), .IN2(n14320), .Q(n14329) );
  OR2X1 U17282 ( .IN1(n16606), .IN2(n16607), .Q(n16597) );
  AND2X1 U17283 ( .IN1(n3628), .IN2(n16608), .Q(n16607) );
  OR2X1 U17284 ( .IN1(n16609), .IN2(n16610), .Q(n16608) );
  OR2X1 U17285 ( .IN1(n16611), .IN2(n16612), .Q(n16610) );
  AND2X1 U17286 ( .IN1(n5596), .IN2(n16613), .Q(n16612) );
  OR2X1 U17287 ( .IN1(n16614), .IN2(n16615), .Q(n16613) );
  AND2X1 U17288 ( .IN1(g1760), .IN2(g1752), .Q(n16615) );
  AND2X1 U17289 ( .IN1(g1792), .IN2(g1744), .Q(n16614) );
  AND2X1 U17290 ( .IN1(n16616), .IN2(n5359), .Q(n16611) );
  AND2X1 U17291 ( .IN1(n5602), .IN2(g1748), .Q(n16616) );
  AND2X1 U17292 ( .IN1(n10544), .IN2(g1736), .Q(n16609) );
  AND2X1 U17293 ( .IN1(g1783), .IN2(n5602), .Q(n10544) );
  AND2X1 U17294 ( .IN1(n10820), .IN2(n14320), .Q(n3628) );
  AND2X1 U17295 ( .IN1(n15915), .IN2(g1740), .Q(n16606) );
  AND2X1 U17296 ( .IN1(n10815), .IN2(n15918), .Q(n15915) );
  AND2X1 U17297 ( .IN1(n14320), .IN2(n16617), .Q(n15918) );
  AND2X1 U17298 ( .IN1(g1760), .IN2(g1792), .Q(n16617) );
  INVX0 U17299 ( .INP(n16605), .ZN(n14320) );
  OR2X1 U17300 ( .IN1(n16618), .IN2(n16502), .Q(n16605) );
  OR2X1 U17301 ( .IN1(n4411), .IN2(n16442), .Q(n16502) );
  INVX0 U17302 ( .INP(n15673), .ZN(n4411) );
  AND2X1 U17303 ( .IN1(g2715), .IN2(n5465), .Q(n15673) );
  AND2X1 U17304 ( .IN1(n12071), .IN2(g2775), .Q(n16618) );
  OR2X1 U17305 ( .IN1(n16619), .IN2(n16620), .Q(g29241) );
  AND2X1 U17306 ( .IN1(n16621), .IN2(g1677), .Q(n16620) );
  OR2X1 U17307 ( .IN1(n10891), .IN2(n16622), .Q(n16621) );
  AND2X1 U17308 ( .IN1(n14355), .IN2(n11100), .Q(n16622) );
  OR2X1 U17309 ( .IN1(n10548), .IN2(n10196), .Q(n11100) );
  AND2X1 U17310 ( .IN1(n16623), .IN2(g1691), .Q(n16619) );
  OR2X1 U17311 ( .IN1(n16624), .IN2(n14344), .Q(n16623) );
  AND2X1 U17312 ( .IN1(n4458), .IN2(n10802), .Q(n16624) );
  OR2X1 U17313 ( .IN1(n16625), .IN2(n16626), .Q(g29240) );
  OR2X1 U17314 ( .IN1(n16627), .IN2(n16628), .Q(n16626) );
  AND2X1 U17315 ( .IN1(n10909), .IN2(g1657), .Q(n16628) );
  AND2X1 U17316 ( .IN1(n15949), .IN2(g1604), .Q(n16627) );
  AND2X1 U17317 ( .IN1(n14355), .IN2(n16629), .Q(n15949) );
  AND2X1 U17318 ( .IN1(g1657), .IN2(g1624), .Q(n16629) );
  OR2X1 U17319 ( .IN1(n16630), .IN2(n16631), .Q(n16625) );
  AND2X1 U17320 ( .IN1(n14344), .IN2(g1677), .Q(n16631) );
  AND2X1 U17321 ( .IN1(n10820), .IN2(n16632), .Q(n14344) );
  AND2X1 U17322 ( .IN1(n3646), .IN2(n16633), .Q(n16630) );
  OR2X1 U17323 ( .IN1(n16634), .IN2(n16635), .Q(n16633) );
  OR2X1 U17324 ( .IN1(n16636), .IN2(n16637), .Q(n16635) );
  AND2X1 U17325 ( .IN1(n10548), .IN2(g1600), .Q(n16637) );
  AND2X1 U17326 ( .IN1(n5370), .IN2(test_so94), .Q(n10548) );
  AND2X1 U17327 ( .IN1(g25167), .IN2(g1620), .Q(n16636) );
  OR2X1 U17328 ( .IN1(n16638), .IN2(n16639), .Q(n16634) );
  AND2X1 U17329 ( .IN1(n16640), .IN2(n10556), .Q(n16639) );
  OR2X1 U17330 ( .IN1(n16641), .IN2(n16642), .Q(n16640) );
  AND2X1 U17331 ( .IN1(g1657), .IN2(g1608), .Q(n16642) );
  AND2X1 U17332 ( .IN1(g1624), .IN2(n9303), .Q(n16641) );
  AND2X1 U17333 ( .IN1(n16643), .IN2(n5525), .Q(n16638) );
  AND2X1 U17334 ( .IN1(n5370), .IN2(g1612), .Q(n16643) );
  AND2X1 U17335 ( .IN1(n10820), .IN2(n14355), .Q(n3646) );
  INVX0 U17336 ( .INP(n16632), .ZN(n14355) );
  OR2X1 U17337 ( .IN1(n15707), .IN2(n16644), .Q(n16632) );
  OR2X1 U17338 ( .IN1(n16442), .IN2(n16645), .Q(n16644) );
  AND2X1 U17339 ( .IN1(n12071), .IN2(g2771), .Q(n16645) );
  AND2X1 U17340 ( .IN1(n16646), .IN2(n12071), .Q(n16442) );
  AND2X1 U17341 ( .IN1(n10520), .IN2(n5301), .Q(n12071) );
  INVX0 U17342 ( .INP(n4388), .ZN(n16646) );
  OR2X1 U17343 ( .IN1(g2719), .IN2(g2715), .Q(n15707) );
  OR2X1 U17344 ( .IN1(n16647), .IN2(n16648), .Q(g29239) );
  OR2X1 U17345 ( .IN1(n16649), .IN2(n16650), .Q(n16648) );
  AND2X1 U17346 ( .IN1(n16651), .IN2(n10803), .Q(n16650) );
  AND2X1 U17347 ( .IN1(n16652), .IN2(g1454), .Q(n16651) );
  OR2X1 U17348 ( .IN1(n16653), .IN2(n16654), .Q(n16652) );
  AND2X1 U17349 ( .IN1(n10909), .IN2(g1478), .Q(n16649) );
  AND2X1 U17350 ( .IN1(n16655), .IN2(n16656), .Q(n16647) );
  AND2X1 U17351 ( .IN1(n16653), .IN2(n16657), .Q(n16655) );
  XNOR2X1 U17352 ( .IN1(n16658), .IN2(g1448), .Q(n16653) );
  OR2X1 U17353 ( .IN1(n16659), .IN2(n16660), .Q(g29238) );
  OR2X1 U17354 ( .IN1(n16661), .IN2(n16662), .Q(n16660) );
  AND2X1 U17355 ( .IN1(n16663), .IN2(g1484), .Q(n16662) );
  OR2X1 U17356 ( .IN1(n16664), .IN2(n16665), .Q(n16663) );
  AND2X1 U17357 ( .IN1(n16666), .IN2(n10803), .Q(n16664) );
  AND2X1 U17358 ( .IN1(n16667), .IN2(n16668), .Q(n16661) );
  AND2X1 U17359 ( .IN1(n16666), .IN2(n16656), .Q(n16667) );
  XNOR2X1 U17360 ( .IN1(n16658), .IN2(g1300), .Q(n16666) );
  AND2X1 U17361 ( .IN1(n10909), .IN2(g1472), .Q(n16659) );
  OR2X1 U17362 ( .IN1(n16669), .IN2(n16670), .Q(g29237) );
  OR2X1 U17363 ( .IN1(n16671), .IN2(n16672), .Q(n16670) );
  AND2X1 U17364 ( .IN1(n16673), .IN2(n10803), .Q(n16672) );
  AND2X1 U17365 ( .IN1(n16674), .IN2(g1467), .Q(n16673) );
  OR2X1 U17366 ( .IN1(n16675), .IN2(n16676), .Q(n16674) );
  OR2X1 U17367 ( .IN1(n10474), .IN2(n16677), .Q(n16676) );
  AND2X1 U17368 ( .IN1(n10908), .IN2(g1448), .Q(n16671) );
  AND2X1 U17369 ( .IN1(n16678), .IN2(n16679), .Q(n16669) );
  AND2X1 U17370 ( .IN1(n13407), .IN2(g13272), .Q(n16679) );
  AND2X1 U17371 ( .IN1(n16677), .IN2(n16656), .Q(n16678) );
  XNOR2X1 U17372 ( .IN1(n16658), .IN2(g1472), .Q(n16677) );
  OR2X1 U17373 ( .IN1(n16680), .IN2(n16681), .Q(g29236) );
  OR2X1 U17374 ( .IN1(n16682), .IN2(n16683), .Q(n16681) );
  AND2X1 U17375 ( .IN1(n16684), .IN2(n10803), .Q(n16683) );
  AND2X1 U17376 ( .IN1(n16685), .IN2(g1437), .Q(n16684) );
  OR2X1 U17377 ( .IN1(n16686), .IN2(n16687), .Q(n16685) );
  AND2X1 U17378 ( .IN1(n10908), .IN2(g1442), .Q(n16682) );
  AND2X1 U17379 ( .IN1(n16688), .IN2(n16689), .Q(n16680) );
  INVX0 U17380 ( .INP(n16687), .ZN(n16689) );
  AND2X1 U17381 ( .IN1(n16686), .IN2(n16656), .Q(n16688) );
  AND2X1 U17382 ( .IN1(n5850), .IN2(n16690), .Q(n16656) );
  XNOR2X1 U17383 ( .IN1(n16658), .IN2(g1478), .Q(n16686) );
  OR2X1 U17384 ( .IN1(n11668), .IN2(n9267), .Q(n16658) );
  INVX0 U17385 ( .INP(n13530), .ZN(n11668) );
  OR2X1 U17386 ( .IN1(n16691), .IN2(n16692), .Q(g29235) );
  OR2X1 U17387 ( .IN1(n16693), .IN2(n16694), .Q(n16692) );
  AND2X1 U17388 ( .IN1(n4178), .IN2(n5558), .Q(n16694) );
  INVX0 U17389 ( .INP(n16695), .ZN(n16693) );
  OR2X1 U17390 ( .IN1(n16696), .IN2(n5558), .Q(n16695) );
  OR2X1 U17391 ( .IN1(n13799), .IN2(n4178), .Q(n16696) );
  AND2X1 U17392 ( .IN1(n10908), .IN2(g1252), .Q(n16691) );
  OR2X1 U17393 ( .IN1(n16697), .IN2(n16698), .Q(g29234) );
  OR2X1 U17394 ( .IN1(n16699), .IN2(n16700), .Q(n16698) );
  AND2X1 U17395 ( .IN1(n16701), .IN2(n10803), .Q(n16700) );
  AND2X1 U17396 ( .IN1(test_so90), .IN2(n16702), .Q(n16701) );
  OR2X1 U17397 ( .IN1(n16703), .IN2(n16704), .Q(n16702) );
  INVX0 U17398 ( .INP(n16705), .ZN(n16704) );
  AND2X1 U17399 ( .IN1(n10908), .IN2(g1135), .Q(n16699) );
  AND2X1 U17400 ( .IN1(n16706), .IN2(n16707), .Q(n16697) );
  AND2X1 U17401 ( .IN1(n16703), .IN2(n16705), .Q(n16706) );
  XNOR2X1 U17402 ( .IN1(n16708), .IN2(g1105), .Q(n16703) );
  OR2X1 U17403 ( .IN1(n16709), .IN2(n16710), .Q(g29233) );
  OR2X1 U17404 ( .IN1(n16711), .IN2(n16712), .Q(n16710) );
  AND2X1 U17405 ( .IN1(n16713), .IN2(g1141), .Q(n16712) );
  OR2X1 U17406 ( .IN1(n16714), .IN2(n16715), .Q(n16713) );
  AND2X1 U17407 ( .IN1(n16716), .IN2(n10803), .Q(n16714) );
  AND2X1 U17408 ( .IN1(n16717), .IN2(n16718), .Q(n16711) );
  AND2X1 U17409 ( .IN1(n16716), .IN2(n16707), .Q(n16717) );
  XNOR2X1 U17410 ( .IN1(n16708), .IN2(g956), .Q(n16716) );
  AND2X1 U17411 ( .IN1(n10908), .IN2(g1129), .Q(n16709) );
  OR2X1 U17412 ( .IN1(n16719), .IN2(n16720), .Q(g29232) );
  OR2X1 U17413 ( .IN1(n16721), .IN2(n16722), .Q(n16720) );
  AND2X1 U17414 ( .IN1(n16723), .IN2(n10803), .Q(n16722) );
  AND2X1 U17415 ( .IN1(n16724), .IN2(g1124), .Q(n16723) );
  OR2X1 U17416 ( .IN1(n16725), .IN2(n16726), .Q(n16724) );
  AND2X1 U17417 ( .IN1(n10908), .IN2(g1105), .Q(n16721) );
  AND2X1 U17418 ( .IN1(n16727), .IN2(n16728), .Q(n16719) );
  INVX0 U17419 ( .INP(n16726), .ZN(n16728) );
  AND2X1 U17420 ( .IN1(n16725), .IN2(n16707), .Q(n16727) );
  XNOR2X1 U17421 ( .IN1(n16708), .IN2(g1129), .Q(n16725) );
  OR2X1 U17422 ( .IN1(n16729), .IN2(n16730), .Q(g29231) );
  OR2X1 U17423 ( .IN1(n16731), .IN2(n16732), .Q(n16730) );
  AND2X1 U17424 ( .IN1(n16733), .IN2(n10804), .Q(n16732) );
  AND2X1 U17425 ( .IN1(n16734), .IN2(g1094), .Q(n16733) );
  OR2X1 U17426 ( .IN1(n16735), .IN2(n16736), .Q(n16734) );
  AND2X1 U17427 ( .IN1(test_so7), .IN2(n10894), .Q(n16731) );
  AND2X1 U17428 ( .IN1(n16737), .IN2(n16738), .Q(n16729) );
  INVX0 U17429 ( .INP(n16736), .ZN(n16738) );
  AND2X1 U17430 ( .IN1(n16735), .IN2(n16707), .Q(n16737) );
  AND2X1 U17431 ( .IN1(n5851), .IN2(n16739), .Q(n16707) );
  XNOR2X1 U17432 ( .IN1(n16708), .IN2(g1135), .Q(n16735) );
  OR2X1 U17433 ( .IN1(n11669), .IN2(n9367), .Q(n16708) );
  INVX0 U17434 ( .INP(n13780), .ZN(n11669) );
  OR2X1 U17435 ( .IN1(n16740), .IN2(n16741), .Q(g29230) );
  OR2X1 U17436 ( .IN1(n16742), .IN2(n16743), .Q(n16741) );
  AND2X1 U17437 ( .IN1(n4196), .IN2(n5559), .Q(n16743) );
  INVX0 U17438 ( .INP(n16744), .ZN(n16742) );
  OR2X1 U17439 ( .IN1(n16745), .IN2(n5559), .Q(n16744) );
  OR2X1 U17440 ( .IN1(n13818), .IN2(n4196), .Q(n16745) );
  AND2X1 U17441 ( .IN1(n10908), .IN2(g907), .Q(n16740) );
  OR2X1 U17442 ( .IN1(n16746), .IN2(n16747), .Q(g29229) );
  OR2X1 U17443 ( .IN1(n16748), .IN2(n16749), .Q(n16747) );
  AND2X1 U17444 ( .IN1(n16750), .IN2(n5826), .Q(n16749) );
  AND2X1 U17445 ( .IN1(n4516), .IN2(n16751), .Q(n16750) );
  AND2X1 U17446 ( .IN1(n4517), .IN2(g723), .Q(n16748) );
  AND2X1 U17447 ( .IN1(n10908), .IN2(g827), .Q(n16746) );
  OR2X1 U17448 ( .IN1(n16752), .IN2(n16753), .Q(g29228) );
  AND2X1 U17449 ( .IN1(n10908), .IN2(g736), .Q(n16753) );
  AND2X1 U17450 ( .IN1(n2404), .IN2(n16754), .Q(n16752) );
  XOR2X1 U17451 ( .IN1(test_so60), .IN2(n16067), .Q(n16754) );
  INVX0 U17452 ( .INP(n16755), .ZN(n16067) );
  OR2X1 U17453 ( .IN1(n16756), .IN2(n16757), .Q(n16755) );
  AND2X1 U17454 ( .IN1(n5482), .IN2(g12184), .Q(n16756) );
  OR2X1 U17455 ( .IN1(n16758), .IN2(n16759), .Q(g29227) );
  OR2X1 U17456 ( .IN1(n16760), .IN2(n16761), .Q(n16759) );
  AND2X1 U17457 ( .IN1(n4524), .IN2(test_so70), .Q(n16761) );
  AND2X1 U17458 ( .IN1(n16762), .IN2(n10580), .Q(n16760) );
  AND2X1 U17459 ( .IN1(n4523), .IN2(n16763), .Q(n16762) );
  AND2X1 U17460 ( .IN1(n10908), .IN2(g676), .Q(n16758) );
  OR2X1 U17461 ( .IN1(n16764), .IN2(n16765), .Q(g29226) );
  OR2X1 U17462 ( .IN1(n16766), .IN2(n16767), .Q(n16765) );
  AND2X1 U17463 ( .IN1(n16768), .IN2(n5751), .Q(n16767) );
  AND2X1 U17464 ( .IN1(n4526), .IN2(n16763), .Q(n16768) );
  AND2X1 U17465 ( .IN1(n16769), .IN2(g676), .Q(n16766) );
  AND2X1 U17466 ( .IN1(n4525), .IN2(n16770), .Q(n16769) );
  INVX0 U17467 ( .INP(n4526), .ZN(n16770) );
  INVX0 U17468 ( .INP(n16771), .ZN(n16764) );
  OR2X1 U17469 ( .IN1(n10739), .IN2(n10042), .Q(n16771) );
  OR2X1 U17470 ( .IN1(n16772), .IN2(n16773), .Q(g29225) );
  AND2X1 U17471 ( .IN1(n10908), .IN2(g667), .Q(n16773) );
  AND2X1 U17472 ( .IN1(n16774), .IN2(n4525), .Q(n16772) );
  AND2X1 U17473 ( .IN1(n10820), .IN2(n16763), .Q(n4525) );
  AND2X1 U17474 ( .IN1(g703), .IN2(n16775), .Q(n16763) );
  OR2X1 U17475 ( .IN1(n16776), .IN2(n16777), .Q(n16775) );
  OR2X1 U17476 ( .IN1(n120), .IN2(n10128), .Q(n16777) );
  OR2X1 U17477 ( .IN1(n4535), .IN2(n16778), .Q(n16776) );
  XNOR2X1 U17478 ( .IN1(n10188), .IN2(g655), .Q(n4535) );
  XNOR2X1 U17479 ( .IN1(n16779), .IN2(n10042), .Q(n16774) );
  OR2X1 U17480 ( .IN1(n16780), .IN2(n16781), .Q(g29224) );
  OR2X1 U17481 ( .IN1(n16782), .IN2(n16783), .Q(n16781) );
  AND2X1 U17482 ( .IN1(n4201), .IN2(n5336), .Q(n16783) );
  AND2X1 U17483 ( .IN1(n16784), .IN2(g586), .Q(n16782) );
  AND2X1 U17484 ( .IN1(n2421), .IN2(n16785), .Q(n16784) );
  INVX0 U17485 ( .INP(n4201), .ZN(n16785) );
  AND2X1 U17486 ( .IN1(n10908), .IN2(g572), .Q(n16780) );
  OR2X1 U17487 ( .IN1(n16786), .IN2(n16787), .Q(g29223) );
  OR2X1 U17488 ( .IN1(n16788), .IN2(n16789), .Q(n16787) );
  AND2X1 U17489 ( .IN1(n16790), .IN2(n10804), .Q(n16789) );
  OR2X1 U17490 ( .IN1(n16791), .IN2(n4962), .Q(n16790) );
  AND2X1 U17491 ( .IN1(n16792), .IN2(g490), .Q(n16791) );
  AND2X1 U17492 ( .IN1(n10908), .IN2(g482), .Q(n16788) );
  INVX0 U17493 ( .INP(n16793), .ZN(n16786) );
  OR2X1 U17494 ( .IN1(n16792), .IN2(g490), .Q(n16793) );
  OR2X1 U17495 ( .IN1(n5820), .IN2(n16794), .Q(n16792) );
  OR2X1 U17496 ( .IN1(n16795), .IN2(n16796), .Q(g29222) );
  OR2X1 U17497 ( .IN1(n16797), .IN2(n16798), .Q(n16796) );
  AND2X1 U17498 ( .IN1(n16799), .IN2(n5358), .Q(n16798) );
  AND2X1 U17499 ( .IN1(n16800), .IN2(n3676), .Q(n16799) );
  AND2X1 U17500 ( .IN1(n16801), .IN2(g417), .Q(n16797) );
  OR2X1 U17501 ( .IN1(n10878), .IN2(n16802), .Q(n16801) );
  AND2X1 U17502 ( .IN1(n4948), .IN2(n16803), .Q(n16802) );
  INVX0 U17503 ( .INP(n3676), .ZN(n16803) );
  XNOR2X1 U17504 ( .IN1(n16804), .IN2(g417), .Q(n3676) );
  OR2X1 U17505 ( .IN1(n16805), .IN2(n16806), .Q(n16804) );
  AND2X1 U17506 ( .IN1(n16807), .IN2(n10466), .Q(n16806) );
  OR2X1 U17507 ( .IN1(n16808), .IN2(n16809), .Q(n16807) );
  AND2X1 U17508 ( .IN1(n10465), .IN2(g424), .Q(n16809) );
  AND2X1 U17509 ( .IN1(g437), .IN2(g392), .Q(n16808) );
  AND2X1 U17510 ( .IN1(n16810), .IN2(g405), .Q(n16805) );
  OR2X1 U17511 ( .IN1(n16811), .IN2(n16812), .Q(n16810) );
  AND2X1 U17512 ( .IN1(g401), .IN2(g392), .Q(n16812) );
  AND2X1 U17513 ( .IN1(n10465), .IN2(g437), .Q(n16811) );
  AND2X1 U17514 ( .IN1(n16813), .IN2(g411), .Q(n16795) );
  OR2X1 U17515 ( .IN1(n16814), .IN2(n16815), .Q(g28105) );
  OR2X1 U17516 ( .IN1(n16816), .IN2(n16817), .Q(n16815) );
  AND2X1 U17517 ( .IN1(n16818), .IN2(n10804), .Q(n16817) );
  AND2X1 U17518 ( .IN1(n16121), .IN2(n13113), .Q(n16818) );
  INVX0 U17519 ( .INP(n10540), .ZN(n13113) );
  OR2X1 U17520 ( .IN1(n16819), .IN2(n16820), .Q(n16121) );
  AND2X1 U17521 ( .IN1(n16821), .IN2(g6727), .Q(n16820) );
  OR2X1 U17522 ( .IN1(n16822), .IN2(n16823), .Q(n16821) );
  OR2X1 U17523 ( .IN1(n16824), .IN2(n16825), .Q(n16823) );
  OR2X1 U17524 ( .IN1(n16826), .IN2(n16827), .Q(n16825) );
  AND2X1 U17525 ( .IN1(test_so80), .IN2(n16828), .Q(n16827) );
  OR2X1 U17526 ( .IN1(n16829), .IN2(n16830), .Q(n16828) );
  AND2X1 U17527 ( .IN1(test_so71), .IN2(n11095), .Q(n16829) );
  AND2X1 U17528 ( .IN1(n16831), .IN2(n10557), .Q(n16826) );
  AND2X1 U17529 ( .IN1(n11091), .IN2(n16832), .Q(n16824) );
  OR2X1 U17530 ( .IN1(n16833), .IN2(n16834), .Q(n16832) );
  AND2X1 U17531 ( .IN1(g6581), .IN2(g13099), .Q(n16834) );
  AND2X1 U17532 ( .IN1(g6589), .IN2(g6723), .Q(n16833) );
  OR2X1 U17533 ( .IN1(n16835), .IN2(n16836), .Q(n16822) );
  OR2X1 U17534 ( .IN1(n16837), .IN2(n16838), .Q(n16836) );
  AND2X1 U17535 ( .IN1(n16839), .IN2(n11092), .Q(n16838) );
  AND2X1 U17536 ( .IN1(g6625), .IN2(g14749), .Q(n16839) );
  AND2X1 U17537 ( .IN1(n16840), .IN2(n11095), .Q(n16837) );
  AND2X1 U17538 ( .IN1(g6609), .IN2(g17871), .Q(n16840) );
  AND2X1 U17539 ( .IN1(n11096), .IN2(n16841), .Q(n16835) );
  OR2X1 U17540 ( .IN1(n16842), .IN2(n16843), .Q(n16841) );
  AND2X1 U17541 ( .IN1(g6641), .IN2(g17764), .Q(n16843) );
  AND2X1 U17542 ( .IN1(g6657), .IN2(g17722), .Q(n16842) );
  AND2X1 U17543 ( .IN1(n5531), .IN2(n16844), .Q(n16819) );
  OR2X1 U17544 ( .IN1(n16845), .IN2(n16846), .Q(n16844) );
  OR2X1 U17545 ( .IN1(n16847), .IN2(n16848), .Q(n16846) );
  OR2X1 U17546 ( .IN1(n16849), .IN2(n16850), .Q(n16848) );
  AND2X1 U17547 ( .IN1(test_so80), .IN2(n16851), .Q(n16850) );
  OR2X1 U17548 ( .IN1(n16852), .IN2(n16831), .Q(n16851) );
  OR2X1 U17549 ( .IN1(n16853), .IN2(n16854), .Q(n16831) );
  OR2X1 U17550 ( .IN1(n16855), .IN2(n16856), .Q(n16854) );
  AND2X1 U17551 ( .IN1(n16857), .IN2(n11092), .Q(n16856) );
  AND2X1 U17552 ( .IN1(g6653), .IN2(g17688), .Q(n16857) );
  AND2X1 U17553 ( .IN1(n16858), .IN2(n11095), .Q(n16855) );
  AND2X1 U17554 ( .IN1(g6637), .IN2(g17778), .Q(n16858) );
  AND2X1 U17555 ( .IN1(n16859), .IN2(n11091), .Q(n16853) );
  AND2X1 U17556 ( .IN1(g6621), .IN2(g14828), .Q(n16859) );
  AND2X1 U17557 ( .IN1(n11096), .IN2(g6601), .Q(n16852) );
  AND2X1 U17558 ( .IN1(n16830), .IN2(n10557), .Q(n16849) );
  OR2X1 U17559 ( .IN1(n16860), .IN2(n16861), .Q(n16830) );
  OR2X1 U17560 ( .IN1(n16862), .IN2(n16863), .Q(n16861) );
  AND2X1 U17561 ( .IN1(n16864), .IN2(n11096), .Q(n16863) );
  AND2X1 U17562 ( .IN1(g17778), .IN2(g6629), .Q(n16864) );
  AND2X1 U17563 ( .IN1(n16865), .IN2(n11092), .Q(n16862) );
  AND2X1 U17564 ( .IN1(g6613), .IN2(g14828), .Q(n16865) );
  AND2X1 U17565 ( .IN1(n16866), .IN2(n11091), .Q(n16860) );
  AND2X1 U17566 ( .IN1(g17688), .IN2(g6645), .Q(n16866) );
  AND2X1 U17567 ( .IN1(n11092), .IN2(n16867), .Q(n16847) );
  OR2X1 U17568 ( .IN1(n16868), .IN2(n16869), .Q(n16867) );
  AND2X1 U17569 ( .IN1(g13099), .IN2(g6593), .Q(n16869) );
  AND2X1 U17570 ( .IN1(g6723), .IN2(g6605), .Q(n16868) );
  AND2X1 U17571 ( .IN1(g6682), .IN2(n5398), .Q(n11092) );
  OR2X1 U17572 ( .IN1(n16870), .IN2(n16871), .Q(n16845) );
  OR2X1 U17573 ( .IN1(n16872), .IN2(n16873), .Q(n16871) );
  AND2X1 U17574 ( .IN1(n16874), .IN2(n11091), .Q(n16873) );
  AND2X1 U17575 ( .IN1(n5590), .IN2(n5398), .Q(n11091) );
  AND2X1 U17576 ( .IN1(g6633), .IN2(g14749), .Q(n16874) );
  AND2X1 U17577 ( .IN1(n16875), .IN2(n11096), .Q(n16872) );
  AND2X1 U17578 ( .IN1(g6682), .IN2(g6741), .Q(n11096) );
  AND2X1 U17579 ( .IN1(g17871), .IN2(g6617), .Q(n16875) );
  AND2X1 U17580 ( .IN1(n11095), .IN2(n16876), .Q(n16870) );
  OR2X1 U17581 ( .IN1(n16877), .IN2(n16878), .Q(n16876) );
  AND2X1 U17582 ( .IN1(g17722), .IN2(g6597), .Q(n16878) );
  AND2X1 U17583 ( .IN1(g17764), .IN2(g6649), .Q(n16877) );
  AND2X1 U17584 ( .IN1(g6741), .IN2(n5590), .Q(n11095) );
  AND2X1 U17585 ( .IN1(n10908), .IN2(g6657), .Q(n16816) );
  AND2X1 U17586 ( .IN1(n13125), .IN2(g5011), .Q(n16814) );
  OR2X1 U17587 ( .IN1(n16879), .IN2(n16880), .Q(g28102) );
  OR2X1 U17588 ( .IN1(n16881), .IN2(n16882), .Q(n16880) );
  AND2X1 U17589 ( .IN1(n13147), .IN2(g4826), .Q(n16882) );
  AND2X1 U17590 ( .IN1(n13143), .IN2(n16159), .Q(n16881) );
  OR2X1 U17591 ( .IN1(n16883), .IN2(n16884), .Q(n16159) );
  AND2X1 U17592 ( .IN1(n16885), .IN2(n10563), .Q(n16884) );
  OR2X1 U17593 ( .IN1(n16886), .IN2(n16887), .Q(n16885) );
  OR2X1 U17594 ( .IN1(n16888), .IN2(n16889), .Q(n16887) );
  OR2X1 U17595 ( .IN1(n16890), .IN2(n16891), .Q(n16889) );
  AND2X1 U17596 ( .IN1(n16892), .IN2(g12422), .Q(n16891) );
  OR2X1 U17597 ( .IN1(n16893), .IN2(n16894), .Q(n16892) );
  AND2X1 U17598 ( .IN1(n12119), .IN2(g6255), .Q(n16893) );
  AND2X1 U17599 ( .IN1(n5437), .IN2(n16895), .Q(n16890) );
  AND2X1 U17600 ( .IN1(n13132), .IN2(n16896), .Q(n16888) );
  OR2X1 U17601 ( .IN1(n16897), .IN2(n16898), .Q(n16896) );
  AND2X1 U17602 ( .IN1(g17685), .IN2(g6251), .Q(n16898) );
  AND2X1 U17603 ( .IN1(g17743), .IN2(g6303), .Q(n16897) );
  OR2X1 U17604 ( .IN1(n16899), .IN2(n16900), .Q(n16886) );
  OR2X1 U17605 ( .IN1(n16901), .IN2(n16902), .Q(n16900) );
  AND2X1 U17606 ( .IN1(n16903), .IN2(n16904), .Q(n16902) );
  AND2X1 U17607 ( .IN1(g6287), .IN2(g14705), .Q(n16903) );
  AND2X1 U17608 ( .IN1(n16905), .IN2(n12119), .Q(n16901) );
  AND2X1 U17609 ( .IN1(g17845), .IN2(g6271), .Q(n16905) );
  AND2X1 U17610 ( .IN1(n13136), .IN2(n16906), .Q(n16899) );
  OR2X1 U17611 ( .IN1(n16907), .IN2(n16908), .Q(n16906) );
  AND2X1 U17612 ( .IN1(g13085), .IN2(g6247), .Q(n16908) );
  AND2X1 U17613 ( .IN1(g6377), .IN2(g6259), .Q(n16907) );
  AND2X1 U17614 ( .IN1(test_so69), .IN2(n16909), .Q(n16883) );
  OR2X1 U17615 ( .IN1(n16910), .IN2(n16911), .Q(n16909) );
  OR2X1 U17616 ( .IN1(n16912), .IN2(n16913), .Q(n16911) );
  OR2X1 U17617 ( .IN1(n16914), .IN2(n16915), .Q(n16913) );
  AND2X1 U17618 ( .IN1(n16916), .IN2(g12422), .Q(n16915) );
  OR2X1 U17619 ( .IN1(n16917), .IN2(n16895), .Q(n16916) );
  OR2X1 U17620 ( .IN1(n16918), .IN2(n16919), .Q(n16895) );
  OR2X1 U17621 ( .IN1(n16920), .IN2(n16921), .Q(n16919) );
  AND2X1 U17622 ( .IN1(n16922), .IN2(n13136), .Q(n16921) );
  AND2X1 U17623 ( .IN1(g6267), .IN2(g14779), .Q(n16922) );
  AND2X1 U17624 ( .IN1(n16923), .IN2(n12119), .Q(n16920) );
  AND2X1 U17625 ( .IN1(g17760), .IN2(g6283), .Q(n16923) );
  AND2X1 U17626 ( .IN1(n16924), .IN2(n16904), .Q(n16918) );
  AND2X1 U17627 ( .IN1(g17649), .IN2(g6299), .Q(n16924) );
  AND2X1 U17628 ( .IN1(n13132), .IN2(g6239), .Q(n16917) );
  AND2X1 U17629 ( .IN1(n5437), .IN2(n16894), .Q(n16914) );
  OR2X1 U17630 ( .IN1(n16925), .IN2(n16926), .Q(n16894) );
  OR2X1 U17631 ( .IN1(n16927), .IN2(n16928), .Q(n16926) );
  AND2X1 U17632 ( .IN1(n16929), .IN2(n16904), .Q(n16928) );
  AND2X1 U17633 ( .IN1(g6275), .IN2(g14779), .Q(n16929) );
  AND2X1 U17634 ( .IN1(n16930), .IN2(n13136), .Q(n16927) );
  AND2X1 U17635 ( .IN1(g6307), .IN2(g17649), .Q(n16930) );
  AND2X1 U17636 ( .IN1(n16931), .IN2(n13132), .Q(n16925) );
  AND2X1 U17637 ( .IN1(g6291), .IN2(g17760), .Q(n16931) );
  AND2X1 U17638 ( .IN1(n16904), .IN2(n16932), .Q(n16912) );
  OR2X1 U17639 ( .IN1(n16933), .IN2(n16934), .Q(n16932) );
  AND2X1 U17640 ( .IN1(g6235), .IN2(g13085), .Q(n16934) );
  AND2X1 U17641 ( .IN1(g6243), .IN2(g6377), .Q(n16933) );
  OR2X1 U17642 ( .IN1(n16935), .IN2(n16936), .Q(n16910) );
  OR2X1 U17643 ( .IN1(n16937), .IN2(n16938), .Q(n16936) );
  AND2X1 U17644 ( .IN1(n16939), .IN2(n13132), .Q(n16938) );
  AND2X1 U17645 ( .IN1(g6263), .IN2(g17845), .Q(n16939) );
  AND2X1 U17646 ( .IN1(n16940), .IN2(n13136), .Q(n16937) );
  AND2X1 U17647 ( .IN1(g6279), .IN2(g14705), .Q(n16940) );
  AND2X1 U17648 ( .IN1(n12119), .IN2(n16941), .Q(n16935) );
  OR2X1 U17649 ( .IN1(n16942), .IN2(n16943), .Q(n16941) );
  AND2X1 U17650 ( .IN1(g6295), .IN2(g17743), .Q(n16943) );
  AND2X1 U17651 ( .IN1(g6311), .IN2(g17685), .Q(n16942) );
  AND2X1 U17652 ( .IN1(n10908), .IN2(g6311), .Q(n16879) );
  OR2X1 U17653 ( .IN1(n16944), .IN2(n16945), .Q(g28099) );
  OR2X1 U17654 ( .IN1(n16946), .IN2(n16947), .Q(n16945) );
  AND2X1 U17655 ( .IN1(n13164), .IN2(g4831), .Q(n16947) );
  AND2X1 U17656 ( .IN1(n13166), .IN2(n16200), .Q(n16946) );
  OR2X1 U17657 ( .IN1(n16948), .IN2(n16949), .Q(n16200) );
  AND2X1 U17658 ( .IN1(n16950), .IN2(g6035), .Q(n16949) );
  OR2X1 U17659 ( .IN1(n16951), .IN2(n16952), .Q(n16950) );
  OR2X1 U17660 ( .IN1(n16953), .IN2(n16954), .Q(n16952) );
  OR2X1 U17661 ( .IN1(n16955), .IN2(n16956), .Q(n16954) );
  AND2X1 U17662 ( .IN1(n16957), .IN2(g12350), .Q(n16956) );
  OR2X1 U17663 ( .IN1(n16958), .IN2(n16959), .Q(n16957) );
  AND2X1 U17664 ( .IN1(n13154), .IN2(g5893), .Q(n16958) );
  AND2X1 U17665 ( .IN1(n5432), .IN2(n16960), .Q(n16955) );
  AND2X1 U17666 ( .IN1(n16961), .IN2(n16962), .Q(n16953) );
  OR2X1 U17667 ( .IN1(n16963), .IN2(n16964), .Q(n16962) );
  AND2X1 U17668 ( .IN1(g5889), .IN2(g13068), .Q(n16964) );
  AND2X1 U17669 ( .IN1(g5897), .IN2(g6031), .Q(n16963) );
  OR2X1 U17670 ( .IN1(n16965), .IN2(n16966), .Q(n16951) );
  OR2X1 U17671 ( .IN1(n16967), .IN2(n16968), .Q(n16966) );
  AND2X1 U17672 ( .IN1(n16969), .IN2(test_so28), .Q(n16968) );
  AND2X1 U17673 ( .IN1(n13154), .IN2(g17819), .Q(n16969) );
  AND2X1 U17674 ( .IN1(n16970), .IN2(n13158), .Q(n16967) );
  AND2X1 U17675 ( .IN1(g5933), .IN2(g14673), .Q(n16970) );
  AND2X1 U17676 ( .IN1(n12132), .IN2(n16971), .Q(n16965) );
  OR2X1 U17677 ( .IN1(n16972), .IN2(n16973), .Q(n16971) );
  AND2X1 U17678 ( .IN1(test_so13), .IN2(g17646), .Q(n16973) );
  AND2X1 U17679 ( .IN1(g5949), .IN2(g17715), .Q(n16972) );
  AND2X1 U17680 ( .IN1(n5528), .IN2(n16974), .Q(n16948) );
  OR2X1 U17681 ( .IN1(n16975), .IN2(n16976), .Q(n16974) );
  OR2X1 U17682 ( .IN1(n16977), .IN2(n16978), .Q(n16976) );
  OR2X1 U17683 ( .IN1(n16979), .IN2(n16980), .Q(n16978) );
  AND2X1 U17684 ( .IN1(n16981), .IN2(g12350), .Q(n16980) );
  OR2X1 U17685 ( .IN1(n16982), .IN2(n16960), .Q(n16981) );
  OR2X1 U17686 ( .IN1(n16983), .IN2(n16984), .Q(n16960) );
  OR2X1 U17687 ( .IN1(n16985), .IN2(n16986), .Q(n16984) );
  AND2X1 U17688 ( .IN1(n16987), .IN2(n16961), .Q(n16986) );
  AND2X1 U17689 ( .IN1(g5929), .IN2(g14738), .Q(n16987) );
  AND2X1 U17690 ( .IN1(n16988), .IN2(n13158), .Q(n16985) );
  AND2X1 U17691 ( .IN1(g5961), .IN2(g17607), .Q(n16988) );
  AND2X1 U17692 ( .IN1(n16989), .IN2(n13154), .Q(n16983) );
  AND2X1 U17693 ( .IN1(g5945), .IN2(g17739), .Q(n16989) );
  AND2X1 U17694 ( .IN1(n12132), .IN2(g5909), .Q(n16982) );
  AND2X1 U17695 ( .IN1(n5432), .IN2(n16959), .Q(n16979) );
  OR2X1 U17696 ( .IN1(n16990), .IN2(n16991), .Q(n16959) );
  OR2X1 U17697 ( .IN1(n16992), .IN2(n16993), .Q(n16991) );
  AND2X1 U17698 ( .IN1(n16994), .IN2(n13158), .Q(n16993) );
  AND2X1 U17699 ( .IN1(g5921), .IN2(g14738), .Q(n16994) );
  AND2X1 U17700 ( .IN1(n16995), .IN2(n12132), .Q(n16992) );
  AND2X1 U17701 ( .IN1(g17739), .IN2(g5937), .Q(n16995) );
  AND2X1 U17702 ( .IN1(n16996), .IN2(n16961), .Q(n16990) );
  AND2X1 U17703 ( .IN1(g17607), .IN2(g5953), .Q(n16996) );
  AND2X1 U17704 ( .IN1(n13154), .IN2(n16997), .Q(n16977) );
  OR2X1 U17705 ( .IN1(n16998), .IN2(n16999), .Q(n16997) );
  AND2X1 U17706 ( .IN1(g17646), .IN2(g5905), .Q(n16999) );
  AND2X1 U17707 ( .IN1(g17715), .IN2(g5957), .Q(n16998) );
  OR2X1 U17708 ( .IN1(n17000), .IN2(n17001), .Q(n16975) );
  OR2X1 U17709 ( .IN1(n17002), .IN2(n17003), .Q(n17001) );
  AND2X1 U17710 ( .IN1(n17004), .IN2(n16961), .Q(n17003) );
  AND2X1 U17711 ( .IN1(g5941), .IN2(g14673), .Q(n17004) );
  AND2X1 U17712 ( .IN1(n17005), .IN2(n12132), .Q(n17002) );
  AND2X1 U17713 ( .IN1(g17819), .IN2(g5925), .Q(n17005) );
  AND2X1 U17714 ( .IN1(n13158), .IN2(n17006), .Q(n17000) );
  OR2X1 U17715 ( .IN1(n17007), .IN2(n17008), .Q(n17006) );
  AND2X1 U17716 ( .IN1(g13068), .IN2(g5901), .Q(n17008) );
  AND2X1 U17717 ( .IN1(g6031), .IN2(g5913), .Q(n17007) );
  AND2X1 U17718 ( .IN1(test_so13), .IN2(n10894), .Q(n16944) );
  OR2X1 U17719 ( .IN1(n17009), .IN2(n17010), .Q(g28096) );
  OR2X1 U17720 ( .IN1(n17011), .IN2(n17012), .Q(n17010) );
  AND2X1 U17721 ( .IN1(n17013), .IN2(n10805), .Q(n17012) );
  AND2X1 U17722 ( .IN1(n13176), .IN2(n16239), .Q(n17013) );
  OR2X1 U17723 ( .IN1(n17014), .IN2(n17015), .Q(n16239) );
  AND2X1 U17724 ( .IN1(n17016), .IN2(g5689), .Q(n17015) );
  OR2X1 U17725 ( .IN1(n17017), .IN2(n17018), .Q(n17016) );
  OR2X1 U17726 ( .IN1(n17019), .IN2(n17020), .Q(n17018) );
  OR2X1 U17727 ( .IN1(n17021), .IN2(n17022), .Q(n17020) );
  AND2X1 U17728 ( .IN1(n17023), .IN2(g12300), .Q(n17022) );
  OR2X1 U17729 ( .IN1(n17024), .IN2(n17025), .Q(n17023) );
  AND2X1 U17730 ( .IN1(n13175), .IN2(g5547), .Q(n17024) );
  AND2X1 U17731 ( .IN1(n5439), .IN2(n17026), .Q(n17021) );
  AND2X1 U17732 ( .IN1(n17027), .IN2(n17028), .Q(n17019) );
  OR2X1 U17733 ( .IN1(n17029), .IN2(n17030), .Q(n17028) );
  AND2X1 U17734 ( .IN1(g5543), .IN2(g13049), .Q(n17030) );
  AND2X1 U17735 ( .IN1(g5551), .IN2(g5685), .Q(n17029) );
  OR2X1 U17736 ( .IN1(n17031), .IN2(n17032), .Q(n17017) );
  OR2X1 U17737 ( .IN1(n17033), .IN2(n17034), .Q(n17032) );
  AND2X1 U17738 ( .IN1(n17035), .IN2(n13175), .Q(n17034) );
  AND2X1 U17739 ( .IN1(g5571), .IN2(g17813), .Q(n17035) );
  AND2X1 U17740 ( .IN1(n17036), .IN2(n13179), .Q(n17033) );
  AND2X1 U17741 ( .IN1(g5587), .IN2(g14635), .Q(n17036) );
  AND2X1 U17742 ( .IN1(n12124), .IN2(n17037), .Q(n17031) );
  OR2X1 U17743 ( .IN1(n17038), .IN2(n17039), .Q(n17037) );
  AND2X1 U17744 ( .IN1(g5603), .IN2(g17678), .Q(n17039) );
  AND2X1 U17745 ( .IN1(g5619), .IN2(g17604), .Q(n17038) );
  AND2X1 U17746 ( .IN1(n5529), .IN2(n17040), .Q(n17014) );
  OR2X1 U17747 ( .IN1(n17041), .IN2(n17042), .Q(n17040) );
  OR2X1 U17748 ( .IN1(n17043), .IN2(n17044), .Q(n17042) );
  OR2X1 U17749 ( .IN1(n17045), .IN2(n17046), .Q(n17044) );
  AND2X1 U17750 ( .IN1(n17047), .IN2(g12300), .Q(n17046) );
  OR2X1 U17751 ( .IN1(n17048), .IN2(n17026), .Q(n17047) );
  OR2X1 U17752 ( .IN1(n17049), .IN2(n17050), .Q(n17026) );
  OR2X1 U17753 ( .IN1(n17051), .IN2(n17052), .Q(n17050) );
  AND2X1 U17754 ( .IN1(n17053), .IN2(n17027), .Q(n17052) );
  AND2X1 U17755 ( .IN1(g5583), .IN2(g14694), .Q(n17053) );
  AND2X1 U17756 ( .IN1(n17054), .IN2(n13179), .Q(n17051) );
  AND2X1 U17757 ( .IN1(g5615), .IN2(g17580), .Q(n17054) );
  AND2X1 U17758 ( .IN1(n17055), .IN2(n13175), .Q(n17049) );
  AND2X1 U17759 ( .IN1(g5599), .IN2(g17711), .Q(n17055) );
  AND2X1 U17760 ( .IN1(n12124), .IN2(g5563), .Q(n17048) );
  AND2X1 U17761 ( .IN1(n5439), .IN2(n17025), .Q(n17045) );
  OR2X1 U17762 ( .IN1(n17056), .IN2(n17057), .Q(n17025) );
  OR2X1 U17763 ( .IN1(n17058), .IN2(n17059), .Q(n17057) );
  AND2X1 U17764 ( .IN1(n17060), .IN2(n13179), .Q(n17059) );
  AND2X1 U17765 ( .IN1(g5575), .IN2(g14694), .Q(n17060) );
  AND2X1 U17766 ( .IN1(n17061), .IN2(test_so5), .Q(n17058) );
  AND2X1 U17767 ( .IN1(n12124), .IN2(g17711), .Q(n17061) );
  AND2X1 U17768 ( .IN1(n17062), .IN2(n17027), .Q(n17056) );
  AND2X1 U17769 ( .IN1(g17580), .IN2(g5607), .Q(n17062) );
  AND2X1 U17770 ( .IN1(n13175), .IN2(n17063), .Q(n17043) );
  OR2X1 U17771 ( .IN1(n17064), .IN2(n17065), .Q(n17063) );
  AND2X1 U17772 ( .IN1(test_so6), .IN2(g17604), .Q(n17065) );
  AND2X1 U17773 ( .IN1(g17678), .IN2(g5611), .Q(n17064) );
  OR2X1 U17774 ( .IN1(n17066), .IN2(n17067), .Q(n17041) );
  OR2X1 U17775 ( .IN1(n17068), .IN2(n17069), .Q(n17067) );
  AND2X1 U17776 ( .IN1(n17070), .IN2(n17027), .Q(n17069) );
  AND2X1 U17777 ( .IN1(g5595), .IN2(g14635), .Q(n17070) );
  AND2X1 U17778 ( .IN1(n17071), .IN2(n12124), .Q(n17068) );
  AND2X1 U17779 ( .IN1(g17813), .IN2(g5579), .Q(n17071) );
  AND2X1 U17780 ( .IN1(n13179), .IN2(n17072), .Q(n17066) );
  OR2X1 U17781 ( .IN1(n17073), .IN2(n17074), .Q(n17072) );
  AND2X1 U17782 ( .IN1(g13049), .IN2(g5555), .Q(n17074) );
  AND2X1 U17783 ( .IN1(g5685), .IN2(g5567), .Q(n17073) );
  AND2X1 U17784 ( .IN1(n10908), .IN2(g5619), .Q(n17011) );
  AND2X1 U17785 ( .IN1(n13188), .IN2(g4821), .Q(n17009) );
  OR2X1 U17786 ( .IN1(n17075), .IN2(n17076), .Q(g28093) );
  OR2X1 U17787 ( .IN1(n17077), .IN2(n17078), .Q(n17076) );
  AND2X1 U17788 ( .IN1(n17079), .IN2(n10805), .Q(n17078) );
  AND2X1 U17789 ( .IN1(n16278), .IN2(g33959), .Q(n17079) );
  INVX0 U17790 ( .INP(n10535), .ZN(g33959) );
  OR2X1 U17791 ( .IN1(n17080), .IN2(n17081), .Q(n16278) );
  AND2X1 U17792 ( .IN1(n17082), .IN2(n10562), .Q(n17081) );
  OR2X1 U17793 ( .IN1(n17083), .IN2(n17084), .Q(n17082) );
  OR2X1 U17794 ( .IN1(n17085), .IN2(n17086), .Q(n17084) );
  OR2X1 U17795 ( .IN1(n17087), .IN2(n17088), .Q(n17086) );
  AND2X1 U17796 ( .IN1(n17089), .IN2(g12238), .Q(n17088) );
  OR2X1 U17797 ( .IN1(n17090), .IN2(n17091), .Q(n17089) );
  AND2X1 U17798 ( .IN1(g31860), .IN2(g5216), .Q(n17090) );
  AND2X1 U17799 ( .IN1(n5438), .IN2(n17092), .Q(n17087) );
  AND2X1 U17800 ( .IN1(n11083), .IN2(n17093), .Q(n17085) );
  OR2X1 U17801 ( .IN1(n17094), .IN2(n17095), .Q(n17093) );
  AND2X1 U17802 ( .IN1(g5208), .IN2(g13039), .Q(n17095) );
  AND2X1 U17803 ( .IN1(g5220), .IN2(g5339), .Q(n17094) );
  OR2X1 U17804 ( .IN1(n17096), .IN2(n17097), .Q(n17083) );
  OR2X1 U17805 ( .IN1(n17098), .IN2(n17099), .Q(n17097) );
  AND2X1 U17806 ( .IN1(n17100), .IN2(g31860), .Q(n17099) );
  AND2X1 U17807 ( .IN1(g17787), .IN2(g5232), .Q(n17100) );
  AND2X1 U17808 ( .IN1(n17101), .IN2(n11082), .Q(n17098) );
  AND2X1 U17809 ( .IN1(g5248), .IN2(g14597), .Q(n17101) );
  AND2X1 U17810 ( .IN1(n11086), .IN2(n17102), .Q(n17096) );
  OR2X1 U17811 ( .IN1(n17103), .IN2(n17104), .Q(n17102) );
  AND2X1 U17812 ( .IN1(g17577), .IN2(g5212), .Q(n17104) );
  AND2X1 U17813 ( .IN1(g17639), .IN2(g5264), .Q(n17103) );
  AND2X1 U17814 ( .IN1(test_so10), .IN2(n17105), .Q(n17080) );
  OR2X1 U17815 ( .IN1(n17106), .IN2(n17107), .Q(n17105) );
  OR2X1 U17816 ( .IN1(n17108), .IN2(n17109), .Q(n17107) );
  OR2X1 U17817 ( .IN1(n17110), .IN2(n17111), .Q(n17109) );
  AND2X1 U17818 ( .IN1(n17112), .IN2(g12238), .Q(n17111) );
  OR2X1 U17819 ( .IN1(n17113), .IN2(n17092), .Q(n17112) );
  OR2X1 U17820 ( .IN1(n17114), .IN2(n17115), .Q(n17092) );
  OR2X1 U17821 ( .IN1(n17116), .IN2(n17117), .Q(n17115) );
  AND2X1 U17822 ( .IN1(n17118), .IN2(test_so82), .Q(n17117) );
  AND2X1 U17823 ( .IN1(n11083), .IN2(g14662), .Q(n17118) );
  AND2X1 U17824 ( .IN1(n17119), .IN2(n11082), .Q(n17116) );
  AND2X1 U17825 ( .IN1(g17519), .IN2(g5260), .Q(n17119) );
  AND2X1 U17826 ( .IN1(n17120), .IN2(g31860), .Q(n17114) );
  AND2X1 U17827 ( .IN1(g17674), .IN2(g5244), .Q(n17120) );
  AND2X1 U17828 ( .IN1(n11086), .IN2(g5200), .Q(n17113) );
  AND2X1 U17829 ( .IN1(n5438), .IN2(n17091), .Q(n17110) );
  OR2X1 U17830 ( .IN1(n17121), .IN2(n17122), .Q(n17091) );
  OR2X1 U17831 ( .IN1(n17123), .IN2(n17124), .Q(n17122) );
  AND2X1 U17832 ( .IN1(n17125), .IN2(n11082), .Q(n17124) );
  AND2X1 U17833 ( .IN1(g5236), .IN2(g14662), .Q(n17125) );
  AND2X1 U17834 ( .IN1(n17126), .IN2(n11086), .Q(n17123) );
  AND2X1 U17835 ( .IN1(g5252), .IN2(g17674), .Q(n17126) );
  AND2X1 U17836 ( .IN1(n17127), .IN2(n11083), .Q(n17121) );
  AND2X1 U17837 ( .IN1(g5268), .IN2(g17519), .Q(n17127) );
  AND2X1 U17838 ( .IN1(g31860), .IN2(n17128), .Q(n17108) );
  OR2X1 U17839 ( .IN1(n17129), .IN2(n17130), .Q(n17128) );
  AND2X1 U17840 ( .IN1(g5256), .IN2(g17639), .Q(n17130) );
  AND2X1 U17841 ( .IN1(g5272), .IN2(g17577), .Q(n17129) );
  AND2X1 U17842 ( .IN1(g5297), .IN2(g5357), .Q(g31860) );
  OR2X1 U17843 ( .IN1(n17131), .IN2(n17132), .Q(n17106) );
  OR2X1 U17844 ( .IN1(n17133), .IN2(n17134), .Q(n17132) );
  AND2X1 U17845 ( .IN1(n17135), .IN2(n11083), .Q(n17134) );
  AND2X1 U17846 ( .IN1(g5297), .IN2(n5393), .Q(n11083) );
  AND2X1 U17847 ( .IN1(g5240), .IN2(g14597), .Q(n17135) );
  AND2X1 U17848 ( .IN1(n17136), .IN2(n11086), .Q(n17133) );
  AND2X1 U17849 ( .IN1(g5357), .IN2(n5588), .Q(n11086) );
  AND2X1 U17850 ( .IN1(g5224), .IN2(g17787), .Q(n17136) );
  AND2X1 U17851 ( .IN1(n11082), .IN2(n17137), .Q(n17131) );
  OR2X1 U17852 ( .IN1(n17138), .IN2(n17139), .Q(n17137) );
  AND2X1 U17853 ( .IN1(g13039), .IN2(g5196), .Q(n17139) );
  AND2X1 U17854 ( .IN1(g5339), .IN2(g5204), .Q(n17138) );
  AND2X1 U17855 ( .IN1(n5588), .IN2(n5393), .Q(n11082) );
  AND2X1 U17856 ( .IN1(n10908), .IN2(g5272), .Q(n17077) );
  AND2X1 U17857 ( .IN1(n13206), .IN2(g29220), .Q(n17075) );
  OR2X1 U17858 ( .IN1(n17140), .IN2(n17141), .Q(g28092) );
  AND2X1 U17859 ( .IN1(n14529), .IN2(n10805), .Q(n17141) );
  AND2X1 U17860 ( .IN1(n17142), .IN2(n14507), .Q(n14529) );
  OR2X1 U17861 ( .IN1(g5052), .IN2(n17143), .Q(n14507) );
  OR2X1 U17862 ( .IN1(g84), .IN2(n17144), .Q(n17143) );
  OR2X1 U17863 ( .IN1(g5041), .IN2(n17145), .Q(n17142) );
  OR2X1 U17864 ( .IN1(n17146), .IN2(n17144), .Q(n17145) );
  OR2X1 U17865 ( .IN1(g5046), .IN2(n17147), .Q(n17144) );
  OR2X1 U17866 ( .IN1(n5615), .IN2(n10507), .Q(n17147) );
  AND2X1 U17867 ( .IN1(n10908), .IN2(g5057), .Q(n17140) );
  OR2X1 U17868 ( .IN1(n17148), .IN2(n14509), .Q(g28091) );
  AND2X1 U17869 ( .IN1(n10818), .IN2(n17149), .Q(n14509) );
  INVX0 U17870 ( .INP(n17150), .ZN(n17149) );
  OR2X1 U17871 ( .IN1(n17151), .IN2(n17152), .Q(n17150) );
  AND2X1 U17872 ( .IN1(n17153), .IN2(g84), .Q(n17152) );
  AND2X1 U17873 ( .IN1(n17154), .IN2(g5041), .Q(n17153) );
  AND2X1 U17874 ( .IN1(n17155), .IN2(n17146), .Q(n17151) );
  INVX0 U17875 ( .INP(g84), .ZN(n17146) );
  AND2X1 U17876 ( .IN1(n17154), .IN2(g5052), .Q(n17155) );
  AND2X1 U17877 ( .IN1(n5615), .IN2(n17156), .Q(n17154) );
  AND2X1 U17878 ( .IN1(g5046), .IN2(g5062), .Q(n17156) );
  AND2X1 U17879 ( .IN1(n10907), .IN2(g5069), .Q(n17148) );
  OR2X1 U17880 ( .IN1(n17157), .IN2(n17158), .Q(g28090) );
  AND2X1 U17881 ( .IN1(n17159), .IN2(g4961), .Q(n17158) );
  OR2X1 U17882 ( .IN1(n17160), .IN2(n13237), .Q(n17159) );
  AND2X1 U17883 ( .IN1(n12181), .IN2(n10806), .Q(n17160) );
  AND2X1 U17884 ( .IN1(n17161), .IN2(n12181), .Q(n17157) );
  AND2X1 U17885 ( .IN1(n11165), .IN2(n11154), .Q(n12181) );
  AND2X1 U17886 ( .IN1(n13234), .IN2(n17162), .Q(n17161) );
  OR2X1 U17887 ( .IN1(n17163), .IN2(n17164), .Q(n17162) );
  OR2X1 U17888 ( .IN1(n17165), .IN2(n17166), .Q(n17164) );
  AND2X1 U17889 ( .IN1(n10268), .IN2(n17167), .Q(n17166) );
  AND2X1 U17890 ( .IN1(n13227), .IN2(g4045), .Q(n17165) );
  OR2X1 U17891 ( .IN1(n17168), .IN2(n17169), .Q(n17163) );
  AND2X1 U17892 ( .IN1(n10490), .IN2(n13223), .Q(n17169) );
  AND2X1 U17893 ( .IN1(n12118), .IN2(g4049), .Q(n17168) );
  OR2X1 U17894 ( .IN1(n17170), .IN2(n17171), .Q(g28089) );
  AND2X1 U17895 ( .IN1(n17172), .IN2(g4950), .Q(n17171) );
  OR2X1 U17896 ( .IN1(n17173), .IN2(n13258), .Q(n17172) );
  AND2X1 U17897 ( .IN1(n12192), .IN2(n10806), .Q(n17173) );
  AND2X1 U17898 ( .IN1(n17174), .IN2(n12192), .Q(n17170) );
  AND2X1 U17899 ( .IN1(n11164), .IN2(n11154), .Q(n12192) );
  AND2X1 U17900 ( .IN1(n13255), .IN2(n17175), .Q(n17174) );
  OR2X1 U17901 ( .IN1(n17176), .IN2(n17177), .Q(n17175) );
  OR2X1 U17902 ( .IN1(n17178), .IN2(n17179), .Q(n17177) );
  AND2X1 U17903 ( .IN1(n10266), .IN2(n17180), .Q(n17179) );
  AND2X1 U17904 ( .IN1(n13248), .IN2(g3694), .Q(n17178) );
  OR2X1 U17905 ( .IN1(n17181), .IN2(n17182), .Q(n17176) );
  AND2X1 U17906 ( .IN1(n10498), .IN2(n13244), .Q(n17182) );
  AND2X1 U17907 ( .IN1(n12131), .IN2(g3698), .Q(n17181) );
  OR2X1 U17908 ( .IN1(n17183), .IN2(n17184), .Q(g28088) );
  AND2X1 U17909 ( .IN1(n13279), .IN2(g4939), .Q(n17184) );
  AND2X1 U17910 ( .IN1(n12202), .IN2(n17185), .Q(n17183) );
  AND2X1 U17911 ( .IN1(n17186), .IN2(n10805), .Q(n17185) );
  OR2X1 U17912 ( .IN1(n17187), .IN2(g4939), .Q(n17186) );
  AND2X1 U17913 ( .IN1(n13270), .IN2(n17188), .Q(n17187) );
  OR2X1 U17914 ( .IN1(n17189), .IN2(n17190), .Q(n17188) );
  OR2X1 U17915 ( .IN1(n17191), .IN2(n17192), .Q(n17190) );
  AND2X1 U17916 ( .IN1(n10263), .IN2(n17193), .Q(n17192) );
  AND2X1 U17917 ( .IN1(n13264), .IN2(g3343), .Q(n17191) );
  OR2X1 U17918 ( .IN1(n17194), .IN2(n17195), .Q(n17189) );
  AND2X1 U17919 ( .IN1(n10487), .IN2(n13269), .Q(n17195) );
  AND2X1 U17920 ( .IN1(n12123), .IN2(g3347), .Q(n17194) );
  AND2X1 U17921 ( .IN1(n11154), .IN2(n11169), .Q(n12202) );
  OR2X1 U17922 ( .IN1(n17196), .IN2(n17197), .Q(g28087) );
  AND2X1 U17923 ( .IN1(n13125), .IN2(g4894), .Q(n17197) );
  AND2X1 U17924 ( .IN1(n10816), .IN2(n10540), .Q(n13125) );
  OR2X1 U17925 ( .IN1(n17198), .IN2(n5713), .Q(n10540) );
  AND2X1 U17926 ( .IN1(n13063), .IN2(n17199), .Q(n17198) );
  AND2X1 U17927 ( .IN1(n11169), .IN2(g4888), .Q(n13063) );
  AND2X1 U17928 ( .IN1(n5360), .IN2(n5517), .Q(n11169) );
  AND2X1 U17929 ( .IN1(n17200), .IN2(n11738), .Q(n17196) );
  AND2X1 U17930 ( .IN1(n11168), .IN2(n11154), .Q(n11738) );
  AND2X1 U17931 ( .IN1(g4983), .IN2(n17201), .Q(n11154) );
  AND2X1 U17932 ( .IN1(n10560), .IN2(g4966), .Q(n17201) );
  AND2X1 U17933 ( .IN1(n17202), .IN2(n10806), .Q(n17200) );
  OR2X1 U17934 ( .IN1(n4689), .IN2(g4894), .Q(n17202) );
  OR2X1 U17935 ( .IN1(n17203), .IN2(n17204), .Q(g28086) );
  AND2X1 U17936 ( .IN1(n17205), .IN2(g4771), .Q(n17204) );
  OR2X1 U17937 ( .IN1(n17206), .IN2(n13147), .Q(n17205) );
  AND2X1 U17938 ( .IN1(n10816), .IN2(n13137), .Q(n13147) );
  AND2X1 U17939 ( .IN1(n12229), .IN2(n10806), .Q(n17206) );
  AND2X1 U17940 ( .IN1(n17207), .IN2(n12229), .Q(n17203) );
  AND2X1 U17941 ( .IN1(n11133), .IN2(n11118), .Q(n12229) );
  AND2X1 U17942 ( .IN1(n13143), .IN2(n17208), .Q(n17207) );
  OR2X1 U17943 ( .IN1(n17209), .IN2(n17210), .Q(n17208) );
  OR2X1 U17944 ( .IN1(n17211), .IN2(n17212), .Q(n17210) );
  AND2X1 U17945 ( .IN1(n10264), .IN2(n16904), .Q(n17212) );
  AND2X1 U17946 ( .IN1(n5396), .IN2(n5592), .Q(n16904) );
  AND2X1 U17947 ( .IN1(n13136), .IN2(g6386), .Q(n17211) );
  AND2X1 U17948 ( .IN1(g6336), .IN2(n5396), .Q(n13136) );
  OR2X1 U17949 ( .IN1(n17213), .IN2(n17214), .Q(n17209) );
  AND2X1 U17950 ( .IN1(n10488), .IN2(n13132), .Q(n17214) );
  AND2X1 U17951 ( .IN1(g6395), .IN2(n5592), .Q(n13132) );
  AND2X1 U17952 ( .IN1(n12119), .IN2(g6390), .Q(n17213) );
  AND2X1 U17953 ( .IN1(g6336), .IN2(g6395), .Q(n12119) );
  AND2X1 U17954 ( .IN1(n10815), .IN2(n13133), .Q(n13143) );
  INVX0 U17955 ( .INP(n13137), .ZN(n13133) );
  OR2X1 U17956 ( .IN1(n17215), .IN2(n5656), .Q(n13137) );
  AND2X1 U17957 ( .IN1(n13104), .IN2(n17216), .Q(n17215) );
  AND2X1 U17958 ( .IN1(n11128), .IN2(g4765), .Q(n13104) );
  OR2X1 U17959 ( .IN1(n17217), .IN2(n17218), .Q(g28085) );
  AND2X1 U17960 ( .IN1(n17219), .IN2(g4760), .Q(n17218) );
  OR2X1 U17961 ( .IN1(n17220), .IN2(n13164), .Q(n17219) );
  AND2X1 U17962 ( .IN1(n10815), .IN2(n13159), .Q(n13164) );
  AND2X1 U17963 ( .IN1(n12240), .IN2(n10788), .Q(n17220) );
  AND2X1 U17964 ( .IN1(n17221), .IN2(n12240), .Q(n17217) );
  AND2X1 U17965 ( .IN1(n11132), .IN2(n11118), .Q(n12240) );
  AND2X1 U17966 ( .IN1(n13166), .IN2(n17222), .Q(n17221) );
  OR2X1 U17967 ( .IN1(n17223), .IN2(n17224), .Q(n17222) );
  OR2X1 U17968 ( .IN1(n17225), .IN2(n17226), .Q(n17224) );
  AND2X1 U17969 ( .IN1(n10265), .IN2(n16961), .Q(n17226) );
  AND2X1 U17970 ( .IN1(n10559), .IN2(n5589), .Q(n16961) );
  AND2X1 U17971 ( .IN1(n13158), .IN2(g6040), .Q(n17225) );
  AND2X1 U17972 ( .IN1(n10559), .IN2(g5990), .Q(n13158) );
  OR2X1 U17973 ( .IN1(n17227), .IN2(n17228), .Q(n17223) );
  AND2X1 U17974 ( .IN1(test_so50), .IN2(n12132), .Q(n17228) );
  AND2X1 U17975 ( .IN1(g5990), .IN2(test_so57), .Q(n12132) );
  AND2X1 U17976 ( .IN1(n13154), .IN2(n10579), .Q(n17227) );
  AND2X1 U17977 ( .IN1(test_so57), .IN2(n5589), .Q(n13154) );
  AND2X1 U17978 ( .IN1(n10810), .IN2(n13155), .Q(n13166) );
  INVX0 U17979 ( .INP(n13159), .ZN(n13155) );
  OR2X1 U17980 ( .IN1(n17229), .IN2(n10435), .Q(n13159) );
  AND2X1 U17981 ( .IN1(n13105), .IN2(n17216), .Q(n17229) );
  AND2X1 U17982 ( .IN1(n11133), .IN2(g4754), .Q(n13105) );
  AND2X1 U17983 ( .IN1(g4709), .IN2(n5361), .Q(n11133) );
  OR2X1 U17984 ( .IN1(n17230), .IN2(n17231), .Q(g28084) );
  AND2X1 U17985 ( .IN1(n13188), .IN2(test_so18), .Q(n17231) );
  AND2X1 U17986 ( .IN1(n10821), .IN2(n13180), .Q(n13188) );
  AND2X1 U17987 ( .IN1(n12250), .IN2(n17232), .Q(n17230) );
  AND2X1 U17988 ( .IN1(n17233), .IN2(n10779), .Q(n17232) );
  OR2X1 U17989 ( .IN1(n17234), .IN2(test_so18), .Q(n17233) );
  AND2X1 U17990 ( .IN1(n13176), .IN2(n17235), .Q(n17234) );
  OR2X1 U17991 ( .IN1(n17236), .IN2(n17237), .Q(n17235) );
  OR2X1 U17992 ( .IN1(n17238), .IN2(n17239), .Q(n17237) );
  AND2X1 U17993 ( .IN1(n10267), .IN2(n17027), .Q(n17239) );
  AND2X1 U17994 ( .IN1(n5397), .IN2(n5593), .Q(n17027) );
  AND2X1 U17995 ( .IN1(n13179), .IN2(g5694), .Q(n17238) );
  AND2X1 U17996 ( .IN1(g5644), .IN2(n5397), .Q(n13179) );
  OR2X1 U17997 ( .IN1(n17240), .IN2(n17241), .Q(n17236) );
  AND2X1 U17998 ( .IN1(n10496), .IN2(n13175), .Q(n17241) );
  AND2X1 U17999 ( .IN1(g5703), .IN2(n5593), .Q(n13175) );
  AND2X1 U18000 ( .IN1(n12124), .IN2(g5698), .Q(n17240) );
  AND2X1 U18001 ( .IN1(g5644), .IN2(g5703), .Q(n12124) );
  INVX0 U18002 ( .INP(n13180), .ZN(n13176) );
  OR2X1 U18003 ( .IN1(n17242), .IN2(n5440), .Q(n13180) );
  AND2X1 U18004 ( .IN1(n13106), .IN2(n17216), .Q(n17242) );
  AND2X1 U18005 ( .IN1(n11132), .IN2(g4743), .Q(n13106) );
  AND2X1 U18006 ( .IN1(g4785), .IN2(n5518), .Q(n11132) );
  AND2X1 U18007 ( .IN1(n11118), .IN2(n11129), .Q(n12250) );
  OR2X1 U18008 ( .IN1(n17243), .IN2(n17244), .Q(g28083) );
  AND2X1 U18009 ( .IN1(n13206), .IN2(g4704), .Q(n17244) );
  AND2X1 U18010 ( .IN1(n10815), .IN2(n10535), .Q(n13206) );
  OR2X1 U18011 ( .IN1(n17245), .IN2(n5712), .Q(n10535) );
  AND2X1 U18012 ( .IN1(n13103), .IN2(n17216), .Q(n17245) );
  INVX0 U18013 ( .INP(n17246), .ZN(n17216) );
  OR2X1 U18014 ( .IN1(n17247), .IN2(n17248), .Q(n17246) );
  OR2X1 U18015 ( .IN1(g4793), .IN2(n12426), .Q(n17248) );
  OR2X1 U18016 ( .IN1(n10567), .IN2(n17249), .Q(n12426) );
  OR2X1 U18017 ( .IN1(n10509), .IN2(n10021), .Q(n17249) );
  OR2X1 U18018 ( .IN1(test_so29), .IN2(n5707), .Q(n17247) );
  AND2X1 U18019 ( .IN1(n11129), .IN2(g4698), .Q(n13103) );
  AND2X1 U18020 ( .IN1(n5361), .IN2(n5518), .Q(n11129) );
  AND2X1 U18021 ( .IN1(n17250), .IN2(n11742), .Q(n17243) );
  AND2X1 U18022 ( .IN1(n11128), .IN2(n11118), .Q(n11742) );
  AND2X1 U18023 ( .IN1(g4793), .IN2(n17251), .Q(n11118) );
  AND2X1 U18024 ( .IN1(n10561), .IN2(g4776), .Q(n17251) );
  AND2X1 U18025 ( .IN1(g4709), .IN2(g4785), .Q(n11128) );
  AND2X1 U18026 ( .IN1(n17252), .IN2(n10779), .Q(n17250) );
  OR2X1 U18027 ( .IN1(n4708), .IN2(g4704), .Q(n17252) );
  OR2X1 U18028 ( .IN1(n17253), .IN2(n17254), .Q(g28082) );
  AND2X1 U18029 ( .IN1(n17255), .IN2(n5752), .Q(n17254) );
  AND2X1 U18030 ( .IN1(n11586), .IN2(n10779), .Q(n17255) );
  INVX0 U18031 ( .INP(n17256), .ZN(n11586) );
  AND2X1 U18032 ( .IN1(n17257), .IN2(g4521), .Q(n17253) );
  OR2X1 U18033 ( .IN1(n10878), .IN2(n17258), .Q(n17257) );
  OR2X1 U18034 ( .IN1(n17259), .IN2(n17260), .Q(g28074) );
  OR2X1 U18035 ( .IN1(n17261), .IN2(n17262), .Q(n17260) );
  AND2X1 U18036 ( .IN1(n4714), .IN2(n4721), .Q(n17262) );
  AND2X1 U18037 ( .IN1(n17263), .IN2(n17264), .Q(n17261) );
  INVX0 U18038 ( .INP(n4714), .ZN(n17264) );
  AND2X1 U18039 ( .IN1(n10816), .IN2(g4122), .Q(n17263) );
  AND2X1 U18040 ( .IN1(n10907), .IN2(g4119), .Q(n17259) );
  OR2X1 U18041 ( .IN1(n17265), .IN2(n17266), .Q(g28073) );
  OR2X1 U18042 ( .IN1(n17267), .IN2(n17268), .Q(n17266) );
  AND2X1 U18043 ( .IN1(n10907), .IN2(g4116), .Q(n17268) );
  AND2X1 U18044 ( .IN1(n17269), .IN2(n10779), .Q(n17267) );
  AND2X1 U18045 ( .IN1(n17270), .IN2(g4119), .Q(n17269) );
  AND2X1 U18046 ( .IN1(n17271), .IN2(n4721), .Q(n17265) );
  INVX0 U18047 ( .INP(n17270), .ZN(n17271) );
  OR2X1 U18048 ( .IN1(n5711), .IN2(n17272), .Q(n17270) );
  OR2X1 U18049 ( .IN1(n17273), .IN2(n17274), .Q(g28072) );
  OR2X1 U18050 ( .IN1(n17275), .IN2(n17276), .Q(n17274) );
  AND2X1 U18051 ( .IN1(n10907), .IN2(g4112), .Q(n17276) );
  AND2X1 U18052 ( .IN1(n17277), .IN2(n10779), .Q(n17275) );
  AND2X1 U18053 ( .IN1(n17278), .IN2(g4116), .Q(n17277) );
  AND2X1 U18054 ( .IN1(n17279), .IN2(n4721), .Q(n17273) );
  INVX0 U18055 ( .INP(n17278), .ZN(n17279) );
  OR2X1 U18056 ( .IN1(n11099), .IN2(n17280), .Q(n17278) );
  OR2X1 U18057 ( .IN1(n5416), .IN2(g4057), .Q(n17280) );
  OR2X1 U18058 ( .IN1(n17281), .IN2(n17282), .Q(g28071) );
  INVX0 U18059 ( .INP(n17283), .ZN(n17282) );
  OR2X1 U18060 ( .IN1(n17284), .IN2(n10391), .Q(n17283) );
  AND2X1 U18061 ( .IN1(n17284), .IN2(g4112), .Q(n17281) );
  AND2X1 U18062 ( .IN1(n10816), .IN2(n17285), .Q(n17284) );
  OR2X1 U18063 ( .IN1(n17272), .IN2(g4057), .Q(n17285) );
  OR2X1 U18064 ( .IN1(g4064), .IN2(n11099), .Q(n17272) );
  OR2X1 U18065 ( .IN1(n17286), .IN2(n17287), .Q(n11099) );
  OR2X1 U18066 ( .IN1(g4098), .IN2(g4141), .Q(n17287) );
  OR2X1 U18067 ( .IN1(g4082), .IN2(n17288), .Q(n17286) );
  OR2X1 U18068 ( .IN1(test_so11), .IN2(n14756), .Q(n17288) );
  INVX0 U18069 ( .INP(n12105), .ZN(n14756) );
  AND2X1 U18070 ( .IN1(n5340), .IN2(n5480), .Q(n12105) );
  OR2X1 U18071 ( .IN1(n17289), .IN2(n17290), .Q(g28070) );
  OR2X1 U18072 ( .IN1(n10542), .IN2(n17291), .Q(n17290) );
  AND2X1 U18073 ( .IN1(n17292), .IN2(n10554), .Q(n17291) );
  INVX0 U18074 ( .INP(n16286), .ZN(n17292) );
  OR2X1 U18075 ( .IN1(n17293), .IN2(n17294), .Q(n17289) );
  AND2X1 U18076 ( .IN1(n10907), .IN2(g4082), .Q(n17294) );
  AND2X1 U18077 ( .IN1(n17295), .IN2(n10780), .Q(n17293) );
  AND2X1 U18078 ( .IN1(test_so11), .IN2(n16286), .Q(n17295) );
  OR2X1 U18079 ( .IN1(n10467), .IN2(n17296), .Q(n16286) );
  OR2X1 U18080 ( .IN1(n17297), .IN2(n17298), .Q(g28069) );
  OR2X1 U18081 ( .IN1(n17299), .IN2(n17300), .Q(n17298) );
  AND2X1 U18082 ( .IN1(n13237), .IN2(g4035), .Q(n17300) );
  AND2X1 U18083 ( .IN1(n10816), .IN2(n13228), .Q(n13237) );
  AND2X1 U18084 ( .IN1(n13234), .IN2(n16325), .Q(n17299) );
  OR2X1 U18085 ( .IN1(n17301), .IN2(n17302), .Q(n16325) );
  AND2X1 U18086 ( .IN1(n17303), .IN2(g4040), .Q(n17302) );
  OR2X1 U18087 ( .IN1(n17304), .IN2(n17305), .Q(n17303) );
  OR2X1 U18088 ( .IN1(n17306), .IN2(n17307), .Q(n17305) );
  OR2X1 U18089 ( .IN1(n17308), .IN2(n17309), .Q(n17307) );
  AND2X1 U18090 ( .IN1(n17310), .IN2(g11418), .Q(n17309) );
  OR2X1 U18091 ( .IN1(n17311), .IN2(n17312), .Q(n17310) );
  AND2X1 U18092 ( .IN1(n13223), .IN2(g3893), .Q(n17311) );
  AND2X1 U18093 ( .IN1(n5435), .IN2(n17313), .Q(n17308) );
  AND2X1 U18094 ( .IN1(n17167), .IN2(n17314), .Q(n17306) );
  OR2X1 U18095 ( .IN1(n17315), .IN2(n17316), .Q(n17314) );
  AND2X1 U18096 ( .IN1(test_so24), .IN2(g14518), .Q(n17316) );
  AND2X1 U18097 ( .IN1(g3897), .IN2(g4031), .Q(n17315) );
  OR2X1 U18098 ( .IN1(n17317), .IN2(n17318), .Q(n17304) );
  OR2X1 U18099 ( .IN1(n17319), .IN2(n17320), .Q(n17318) );
  AND2X1 U18100 ( .IN1(n17321), .IN2(n13227), .Q(n17320) );
  AND2X1 U18101 ( .IN1(g3933), .IN2(g13906), .Q(n17321) );
  AND2X1 U18102 ( .IN1(n17322), .IN2(n13223), .Q(n17319) );
  AND2X1 U18103 ( .IN1(g3917), .IN2(g16955), .Q(n17322) );
  AND2X1 U18104 ( .IN1(n12118), .IN2(n17323), .Q(n17317) );
  OR2X1 U18105 ( .IN1(n17324), .IN2(n17325), .Q(n17323) );
  AND2X1 U18106 ( .IN1(test_so65), .IN2(g16748), .Q(n17325) );
  AND2X1 U18107 ( .IN1(g3965), .IN2(g16693), .Q(n17324) );
  AND2X1 U18108 ( .IN1(n5530), .IN2(n17326), .Q(n17301) );
  OR2X1 U18109 ( .IN1(n17327), .IN2(n17328), .Q(n17326) );
  OR2X1 U18110 ( .IN1(n17329), .IN2(n17330), .Q(n17328) );
  OR2X1 U18111 ( .IN1(n17331), .IN2(n17332), .Q(n17330) );
  AND2X1 U18112 ( .IN1(n17333), .IN2(g11418), .Q(n17332) );
  OR2X1 U18113 ( .IN1(n17334), .IN2(n17313), .Q(n17333) );
  OR2X1 U18114 ( .IN1(n17335), .IN2(n17336), .Q(n17313) );
  OR2X1 U18115 ( .IN1(n17337), .IN2(n17338), .Q(n17336) );
  AND2X1 U18116 ( .IN1(n17339), .IN2(n13227), .Q(n17338) );
  AND2X1 U18117 ( .IN1(g3961), .IN2(g16659), .Q(n17339) );
  AND2X1 U18118 ( .IN1(n17340), .IN2(n13223), .Q(n17337) );
  AND2X1 U18119 ( .IN1(g3945), .IN2(g16775), .Q(n17340) );
  AND2X1 U18120 ( .IN1(n17341), .IN2(n17167), .Q(n17335) );
  AND2X1 U18121 ( .IN1(g3929), .IN2(g13966), .Q(n17341) );
  AND2X1 U18122 ( .IN1(n12118), .IN2(g3909), .Q(n17334) );
  AND2X1 U18123 ( .IN1(n5435), .IN2(n17312), .Q(n17331) );
  OR2X1 U18124 ( .IN1(n17342), .IN2(n17343), .Q(n17312) );
  OR2X1 U18125 ( .IN1(n17344), .IN2(n17345), .Q(n17343) );
  AND2X1 U18126 ( .IN1(n17346), .IN2(n12118), .Q(n17345) );
  AND2X1 U18127 ( .IN1(g16775), .IN2(g3937), .Q(n17346) );
  AND2X1 U18128 ( .IN1(n17347), .IN2(n13227), .Q(n17344) );
  AND2X1 U18129 ( .IN1(g3921), .IN2(g13966), .Q(n17347) );
  AND2X1 U18130 ( .IN1(n17348), .IN2(n17167), .Q(n17342) );
  AND2X1 U18131 ( .IN1(g16659), .IN2(g3953), .Q(n17348) );
  AND2X1 U18132 ( .IN1(n13227), .IN2(n17349), .Q(n17329) );
  OR2X1 U18133 ( .IN1(n17350), .IN2(n17351), .Q(n17349) );
  AND2X1 U18134 ( .IN1(g14518), .IN2(g3901), .Q(n17351) );
  AND2X1 U18135 ( .IN1(g4031), .IN2(g3913), .Q(n17350) );
  AND2X1 U18136 ( .IN1(g3990), .IN2(n5395), .Q(n13227) );
  OR2X1 U18137 ( .IN1(n17352), .IN2(n17353), .Q(n17327) );
  OR2X1 U18138 ( .IN1(n17354), .IN2(n17355), .Q(n17353) );
  AND2X1 U18139 ( .IN1(n17356), .IN2(n17167), .Q(n17355) );
  AND2X1 U18140 ( .IN1(n5395), .IN2(n5594), .Q(n17167) );
  AND2X1 U18141 ( .IN1(g3941), .IN2(g13906), .Q(n17356) );
  AND2X1 U18142 ( .IN1(n17357), .IN2(n12118), .Q(n17354) );
  AND2X1 U18143 ( .IN1(g3990), .IN2(g4054), .Q(n12118) );
  AND2X1 U18144 ( .IN1(g16955), .IN2(g3925), .Q(n17357) );
  AND2X1 U18145 ( .IN1(n13223), .IN2(n17358), .Q(n17352) );
  OR2X1 U18146 ( .IN1(n17359), .IN2(n17360), .Q(n17358) );
  AND2X1 U18147 ( .IN1(g16693), .IN2(g3905), .Q(n17360) );
  AND2X1 U18148 ( .IN1(g16748), .IN2(g3957), .Q(n17359) );
  AND2X1 U18149 ( .IN1(g4054), .IN2(n5594), .Q(n13223) );
  AND2X1 U18150 ( .IN1(n10816), .IN2(n13224), .Q(n13234) );
  INVX0 U18151 ( .INP(n13228), .ZN(n13224) );
  OR2X1 U18152 ( .IN1(n17361), .IN2(n5283), .Q(n13228) );
  AND2X1 U18153 ( .IN1(n13064), .IN2(n17199), .Q(n17361) );
  AND2X1 U18154 ( .IN1(n11168), .IN2(g4955), .Q(n13064) );
  AND2X1 U18155 ( .IN1(g4899), .IN2(g4975), .Q(n11168) );
  AND2X1 U18156 ( .IN1(n10907), .IN2(g3965), .Q(n17297) );
  OR2X1 U18157 ( .IN1(n17362), .IN2(n17363), .Q(g28066) );
  OR2X1 U18158 ( .IN1(n17364), .IN2(n17365), .Q(n17363) );
  AND2X1 U18159 ( .IN1(n13258), .IN2(g3684), .Q(n17365) );
  AND2X1 U18160 ( .IN1(n10816), .IN2(n13249), .Q(n13258) );
  AND2X1 U18161 ( .IN1(n13255), .IN2(n16364), .Q(n17364) );
  OR2X1 U18162 ( .IN1(n17366), .IN2(n17367), .Q(n16364) );
  AND2X1 U18163 ( .IN1(n17368), .IN2(g3689), .Q(n17367) );
  OR2X1 U18164 ( .IN1(n17369), .IN2(n17370), .Q(n17368) );
  OR2X1 U18165 ( .IN1(n17371), .IN2(n17372), .Q(n17370) );
  OR2X1 U18166 ( .IN1(n17373), .IN2(n17374), .Q(n17372) );
  AND2X1 U18167 ( .IN1(n17375), .IN2(g11388), .Q(n17374) );
  OR2X1 U18168 ( .IN1(n17376), .IN2(n17377), .Q(n17375) );
  AND2X1 U18169 ( .IN1(n13244), .IN2(g3542), .Q(n17376) );
  AND2X1 U18170 ( .IN1(n5433), .IN2(n17378), .Q(n17373) );
  AND2X1 U18171 ( .IN1(n17180), .IN2(n17379), .Q(n17371) );
  OR2X1 U18172 ( .IN1(n17380), .IN2(n17381), .Q(n17379) );
  AND2X1 U18173 ( .IN1(g3538), .IN2(g14451), .Q(n17381) );
  AND2X1 U18174 ( .IN1(g3546), .IN2(g3680), .Q(n17380) );
  OR2X1 U18175 ( .IN1(n17382), .IN2(n17383), .Q(n17369) );
  OR2X1 U18176 ( .IN1(n17384), .IN2(n17385), .Q(n17383) );
  AND2X1 U18177 ( .IN1(n17386), .IN2(test_so26), .Q(n17385) );
  AND2X1 U18178 ( .IN1(n13248), .IN2(g3582), .Q(n17386) );
  AND2X1 U18179 ( .IN1(n17387), .IN2(n13244), .Q(n17384) );
  AND2X1 U18180 ( .IN1(g3566), .IN2(g16924), .Q(n17387) );
  AND2X1 U18181 ( .IN1(n12131), .IN2(n17388), .Q(n17382) );
  OR2X1 U18182 ( .IN1(n17389), .IN2(n17390), .Q(n17388) );
  AND2X1 U18183 ( .IN1(g3598), .IN2(g16722), .Q(n17390) );
  AND2X1 U18184 ( .IN1(g3614), .IN2(g16656), .Q(n17389) );
  AND2X1 U18185 ( .IN1(n5532), .IN2(n17391), .Q(n17366) );
  OR2X1 U18186 ( .IN1(n17392), .IN2(n17393), .Q(n17391) );
  OR2X1 U18187 ( .IN1(n17394), .IN2(n17395), .Q(n17393) );
  OR2X1 U18188 ( .IN1(n17396), .IN2(n17397), .Q(n17395) );
  AND2X1 U18189 ( .IN1(n17398), .IN2(g11388), .Q(n17397) );
  OR2X1 U18190 ( .IN1(n17399), .IN2(n17378), .Q(n17398) );
  OR2X1 U18191 ( .IN1(n17400), .IN2(n17401), .Q(n17378) );
  OR2X1 U18192 ( .IN1(n17402), .IN2(n17403), .Q(n17401) );
  AND2X1 U18193 ( .IN1(n17404), .IN2(n13248), .Q(n17403) );
  AND2X1 U18194 ( .IN1(g3610), .IN2(g16627), .Q(n17404) );
  AND2X1 U18195 ( .IN1(n17405), .IN2(n13244), .Q(n17402) );
  AND2X1 U18196 ( .IN1(g3594), .IN2(g16744), .Q(n17405) );
  AND2X1 U18197 ( .IN1(n17406), .IN2(n17180), .Q(n17400) );
  AND2X1 U18198 ( .IN1(g3578), .IN2(g13926), .Q(n17406) );
  AND2X1 U18199 ( .IN1(n12131), .IN2(g3558), .Q(n17399) );
  AND2X1 U18200 ( .IN1(n5433), .IN2(n17377), .Q(n17396) );
  OR2X1 U18201 ( .IN1(n17407), .IN2(n17408), .Q(n17377) );
  OR2X1 U18202 ( .IN1(n17409), .IN2(n17410), .Q(n17408) );
  AND2X1 U18203 ( .IN1(n17411), .IN2(n12131), .Q(n17410) );
  AND2X1 U18204 ( .IN1(g16744), .IN2(g3586), .Q(n17411) );
  AND2X1 U18205 ( .IN1(n17412), .IN2(n13248), .Q(n17409) );
  AND2X1 U18206 ( .IN1(g3570), .IN2(g13926), .Q(n17412) );
  AND2X1 U18207 ( .IN1(n17413), .IN2(n17180), .Q(n17407) );
  AND2X1 U18208 ( .IN1(test_so43), .IN2(g16627), .Q(n17413) );
  AND2X1 U18209 ( .IN1(n13248), .IN2(n17414), .Q(n17394) );
  OR2X1 U18210 ( .IN1(n17415), .IN2(n17416), .Q(n17414) );
  AND2X1 U18211 ( .IN1(g14451), .IN2(g3550), .Q(n17416) );
  AND2X1 U18212 ( .IN1(g3680), .IN2(g3562), .Q(n17415) );
  AND2X1 U18213 ( .IN1(g3639), .IN2(n5399), .Q(n13248) );
  OR2X1 U18214 ( .IN1(n17417), .IN2(n17418), .Q(n17392) );
  OR2X1 U18215 ( .IN1(n17419), .IN2(n17420), .Q(n17418) );
  AND2X1 U18216 ( .IN1(n17421), .IN2(n17180), .Q(n17420) );
  AND2X1 U18217 ( .IN1(n5399), .IN2(n5591), .Q(n17180) );
  AND2X1 U18218 ( .IN1(test_so26), .IN2(g3590), .Q(n17421) );
  AND2X1 U18219 ( .IN1(n17422), .IN2(n12131), .Q(n17419) );
  AND2X1 U18220 ( .IN1(g3703), .IN2(g3639), .Q(n12131) );
  AND2X1 U18221 ( .IN1(g16924), .IN2(g3574), .Q(n17422) );
  AND2X1 U18222 ( .IN1(n13244), .IN2(n17423), .Q(n17417) );
  OR2X1 U18223 ( .IN1(n17424), .IN2(n17425), .Q(n17423) );
  AND2X1 U18224 ( .IN1(g16656), .IN2(g3554), .Q(n17425) );
  AND2X1 U18225 ( .IN1(g16722), .IN2(g3606), .Q(n17424) );
  AND2X1 U18226 ( .IN1(g3703), .IN2(n5591), .Q(n13244) );
  AND2X1 U18227 ( .IN1(n10816), .IN2(n13245), .Q(n13255) );
  INVX0 U18228 ( .INP(n13249), .ZN(n13245) );
  OR2X1 U18229 ( .IN1(n17426), .IN2(n5443), .Q(n13249) );
  AND2X1 U18230 ( .IN1(n13061), .IN2(n17199), .Q(n17426) );
  AND2X1 U18231 ( .IN1(n11165), .IN2(g4944), .Q(n13061) );
  AND2X1 U18232 ( .IN1(g4899), .IN2(n5360), .Q(n11165) );
  AND2X1 U18233 ( .IN1(n10907), .IN2(g3614), .Q(n17362) );
  OR2X1 U18234 ( .IN1(n17427), .IN2(n17428), .Q(g28063) );
  OR2X1 U18235 ( .IN1(n17429), .IN2(n17430), .Q(n17428) );
  AND2X1 U18236 ( .IN1(n17431), .IN2(n10780), .Q(n17430) );
  AND2X1 U18237 ( .IN1(n13270), .IN2(n16404), .Q(n17431) );
  OR2X1 U18238 ( .IN1(n17432), .IN2(n17433), .Q(n16404) );
  AND2X1 U18239 ( .IN1(n17434), .IN2(g3338), .Q(n17433) );
  OR2X1 U18240 ( .IN1(n17435), .IN2(n17436), .Q(n17434) );
  OR2X1 U18241 ( .IN1(n17437), .IN2(n17438), .Q(n17436) );
  OR2X1 U18242 ( .IN1(n17439), .IN2(n17440), .Q(n17438) );
  AND2X1 U18243 ( .IN1(n17441), .IN2(g11349), .Q(n17440) );
  OR2X1 U18244 ( .IN1(n17442), .IN2(n17443), .Q(n17441) );
  AND2X1 U18245 ( .IN1(n13269), .IN2(g3191), .Q(n17442) );
  AND2X1 U18246 ( .IN1(n5436), .IN2(n17444), .Q(n17439) );
  AND2X1 U18247 ( .IN1(n17193), .IN2(n17445), .Q(n17437) );
  OR2X1 U18248 ( .IN1(n17446), .IN2(n17447), .Q(n17445) );
  AND2X1 U18249 ( .IN1(test_so91), .IN2(test_so88), .Q(n17447) );
  AND2X1 U18250 ( .IN1(g3187), .IN2(g14421), .Q(n17446) );
  OR2X1 U18251 ( .IN1(n17448), .IN2(n17449), .Q(n17435) );
  OR2X1 U18252 ( .IN1(n17450), .IN2(n17451), .Q(n17449) );
  AND2X1 U18253 ( .IN1(n17452), .IN2(n13264), .Q(n17451) );
  AND2X1 U18254 ( .IN1(g3231), .IN2(g13865), .Q(n17452) );
  AND2X1 U18255 ( .IN1(n17453), .IN2(n13269), .Q(n17450) );
  AND2X1 U18256 ( .IN1(g3215), .IN2(g16874), .Q(n17453) );
  AND2X1 U18257 ( .IN1(n12123), .IN2(n17454), .Q(n17448) );
  OR2X1 U18258 ( .IN1(n17455), .IN2(n17456), .Q(n17454) );
  AND2X1 U18259 ( .IN1(g3247), .IN2(g16686), .Q(n17456) );
  AND2X1 U18260 ( .IN1(g3263), .IN2(g16624), .Q(n17455) );
  AND2X1 U18261 ( .IN1(n5527), .IN2(n17457), .Q(n17432) );
  OR2X1 U18262 ( .IN1(n17458), .IN2(n17459), .Q(n17457) );
  OR2X1 U18263 ( .IN1(n17460), .IN2(n17461), .Q(n17459) );
  OR2X1 U18264 ( .IN1(n17462), .IN2(n17463), .Q(n17461) );
  AND2X1 U18265 ( .IN1(n17464), .IN2(g11349), .Q(n17463) );
  OR2X1 U18266 ( .IN1(n17465), .IN2(n17444), .Q(n17464) );
  OR2X1 U18267 ( .IN1(n17466), .IN2(n17467), .Q(n17444) );
  OR2X1 U18268 ( .IN1(n17468), .IN2(n17469), .Q(n17467) );
  AND2X1 U18269 ( .IN1(n17470), .IN2(n13264), .Q(n17469) );
  AND2X1 U18270 ( .IN1(test_so84), .IN2(g16603), .Q(n17470) );
  AND2X1 U18271 ( .IN1(n17471), .IN2(n13269), .Q(n17468) );
  AND2X1 U18272 ( .IN1(g3243), .IN2(g16718), .Q(n17471) );
  AND2X1 U18273 ( .IN1(n17472), .IN2(n17193), .Q(n17466) );
  AND2X1 U18274 ( .IN1(g3227), .IN2(g13895), .Q(n17472) );
  AND2X1 U18275 ( .IN1(n12123), .IN2(g3207), .Q(n17465) );
  AND2X1 U18276 ( .IN1(n5436), .IN2(n17443), .Q(n17462) );
  OR2X1 U18277 ( .IN1(n17473), .IN2(n17474), .Q(n17443) );
  OR2X1 U18278 ( .IN1(n17475), .IN2(n17476), .Q(n17474) );
  AND2X1 U18279 ( .IN1(n17477), .IN2(n12123), .Q(n17476) );
  AND2X1 U18280 ( .IN1(g16718), .IN2(g3235), .Q(n17477) );
  AND2X1 U18281 ( .IN1(n17478), .IN2(n13264), .Q(n17475) );
  AND2X1 U18282 ( .IN1(g3219), .IN2(g13895), .Q(n17478) );
  AND2X1 U18283 ( .IN1(n17479), .IN2(n17193), .Q(n17473) );
  AND2X1 U18284 ( .IN1(g16603), .IN2(g3251), .Q(n17479) );
  AND2X1 U18285 ( .IN1(n13264), .IN2(n17480), .Q(n17460) );
  OR2X1 U18286 ( .IN1(n17481), .IN2(n17482), .Q(n17480) );
  AND2X1 U18287 ( .IN1(g14421), .IN2(g3199), .Q(n17482) );
  AND2X1 U18288 ( .IN1(test_so91), .IN2(g3211), .Q(n17481) );
  AND2X1 U18289 ( .IN1(g3288), .IN2(n5604), .Q(n13264) );
  OR2X1 U18290 ( .IN1(n17483), .IN2(n17484), .Q(n17458) );
  OR2X1 U18291 ( .IN1(n17485), .IN2(n17486), .Q(n17484) );
  AND2X1 U18292 ( .IN1(n17487), .IN2(n17193), .Q(n17486) );
  AND2X1 U18293 ( .IN1(n5604), .IN2(n5400), .Q(n17193) );
  AND2X1 U18294 ( .IN1(g3239), .IN2(g13865), .Q(n17487) );
  AND2X1 U18295 ( .IN1(n17488), .IN2(n12123), .Q(n17485) );
  AND2X1 U18296 ( .IN1(g3352), .IN2(g3288), .Q(n12123) );
  AND2X1 U18297 ( .IN1(g16874), .IN2(g3223), .Q(n17488) );
  AND2X1 U18298 ( .IN1(n13269), .IN2(n17489), .Q(n17483) );
  OR2X1 U18299 ( .IN1(n17490), .IN2(n17491), .Q(n17489) );
  AND2X1 U18300 ( .IN1(g16624), .IN2(g3203), .Q(n17491) );
  AND2X1 U18301 ( .IN1(g16686), .IN2(g3255), .Q(n17490) );
  AND2X1 U18302 ( .IN1(g3352), .IN2(n5400), .Q(n13269) );
  INVX0 U18303 ( .INP(n13268), .ZN(n13270) );
  AND2X1 U18304 ( .IN1(n10907), .IN2(g3263), .Q(n17429) );
  AND2X1 U18305 ( .IN1(n13279), .IN2(g3333), .Q(n17427) );
  AND2X1 U18306 ( .IN1(n10817), .IN2(n13268), .Q(n13279) );
  OR2X1 U18307 ( .IN1(n17492), .IN2(n5318), .Q(n13268) );
  AND2X1 U18308 ( .IN1(n13062), .IN2(n17199), .Q(n17492) );
  INVX0 U18309 ( .INP(n17493), .ZN(n17199) );
  OR2X1 U18310 ( .IN1(n17494), .IN2(n17495), .Q(n17493) );
  OR2X1 U18311 ( .IN1(g4983), .IN2(n12393), .Q(n17495) );
  OR2X1 U18312 ( .IN1(n10018), .IN2(n17496), .Q(n12393) );
  OR2X1 U18313 ( .IN1(n10506), .IN2(n10478), .Q(n17496) );
  OR2X1 U18314 ( .IN1(test_so58), .IN2(n5706), .Q(n17494) );
  AND2X1 U18315 ( .IN1(n11164), .IN2(g4933), .Q(n13062) );
  AND2X1 U18316 ( .IN1(g4975), .IN2(n5517), .Q(n11164) );
  OR2X1 U18317 ( .IN1(n17497), .IN2(n17498), .Q(g28060) );
  OR2X1 U18318 ( .IN1(n2787), .IN2(n17499), .Q(n17498) );
  INVX0 U18319 ( .INP(n17500), .ZN(n17499) );
  OR2X1 U18320 ( .IN1(n17501), .IN2(g2729), .Q(n17500) );
  OR2X1 U18321 ( .IN1(n17502), .IN2(n17503), .Q(n17497) );
  AND2X1 U18322 ( .IN1(n10907), .IN2(g2724), .Q(n17503) );
  AND2X1 U18323 ( .IN1(n17504), .IN2(n10780), .Q(n17502) );
  AND2X1 U18324 ( .IN1(n17501), .IN2(g2729), .Q(n17504) );
  OR2X1 U18325 ( .IN1(n5301), .IN2(n16413), .Q(n17501) );
  INVX0 U18326 ( .INP(n15677), .ZN(n16413) );
  OR2X1 U18327 ( .IN1(n17505), .IN2(n17506), .Q(g28059) );
  OR2X1 U18328 ( .IN1(n17507), .IN2(n17508), .Q(n17506) );
  AND2X1 U18329 ( .IN1(n4798), .IN2(n16011), .Q(n17508) );
  AND2X1 U18330 ( .IN1(n17509), .IN2(n17510), .Q(n17507) );
  AND2X1 U18331 ( .IN1(n14378), .IN2(n10511), .Q(n17509) );
  AND2X1 U18332 ( .IN1(n10817), .IN2(n13787), .Q(n14378) );
  AND2X1 U18333 ( .IN1(n17511), .IN2(n17512), .Q(n13787) );
  AND2X1 U18334 ( .IN1(n17513), .IN2(n5466), .Q(n17512) );
  INVX0 U18335 ( .INP(n17514), .ZN(n17511) );
  OR2X1 U18336 ( .IN1(n17515), .IN2(n17516), .Q(n17514) );
  AND2X1 U18337 ( .IN1(n17517), .IN2(n17518), .Q(n17516) );
  AND2X1 U18338 ( .IN1(n17519), .IN2(n5322), .Q(n17515) );
  AND2X1 U18339 ( .IN1(n10907), .IN2(g1351), .Q(n17505) );
  OR2X1 U18340 ( .IN1(n17520), .IN2(n17521), .Q(g28058) );
  OR2X1 U18341 ( .IN1(n17522), .IN2(n17523), .Q(n17521) );
  AND2X1 U18342 ( .IN1(n4490), .IN2(n5554), .Q(n17523) );
  INVX0 U18343 ( .INP(n17524), .ZN(n17522) );
  OR2X1 U18344 ( .IN1(n17525), .IN2(n5554), .Q(n17524) );
  OR2X1 U18345 ( .IN1(n13799), .IN2(n4490), .Q(n17525) );
  AND2X1 U18346 ( .IN1(test_so77), .IN2(n10895), .Q(n17520) );
  OR2X1 U18347 ( .IN1(n17526), .IN2(n17527), .Q(g28057) );
  OR2X1 U18348 ( .IN1(n17528), .IN2(n17529), .Q(n17527) );
  AND2X1 U18349 ( .IN1(n4805), .IN2(n16052), .Q(n17529) );
  AND2X1 U18350 ( .IN1(n17530), .IN2(n17531), .Q(n17528) );
  AND2X1 U18351 ( .IN1(n14394), .IN2(n10510), .Q(n17530) );
  AND2X1 U18352 ( .IN1(n10817), .IN2(n13806), .Q(n14394) );
  INVX0 U18353 ( .INP(n17532), .ZN(n13806) );
  OR2X1 U18354 ( .IN1(n17533), .IN2(n17534), .Q(n17532) );
  OR2X1 U18355 ( .IN1(test_so20), .IN2(n17535), .Q(n17534) );
  INVX0 U18356 ( .INP(n17536), .ZN(n17535) );
  OR2X1 U18357 ( .IN1(n17537), .IN2(n17538), .Q(n17533) );
  AND2X1 U18358 ( .IN1(n5321), .IN2(n17539), .Q(n17538) );
  AND2X1 U18359 ( .IN1(n17540), .IN2(n17541), .Q(n17537) );
  AND2X1 U18360 ( .IN1(n10907), .IN2(g1008), .Q(n17526) );
  OR2X1 U18361 ( .IN1(n17542), .IN2(n17543), .Q(g28056) );
  OR2X1 U18362 ( .IN1(n17544), .IN2(n17545), .Q(n17543) );
  AND2X1 U18363 ( .IN1(n4514), .IN2(n5555), .Q(n17545) );
  INVX0 U18364 ( .INP(n17546), .ZN(n17544) );
  OR2X1 U18365 ( .IN1(n17547), .IN2(n5555), .Q(n17546) );
  OR2X1 U18366 ( .IN1(n13818), .IN2(n4514), .Q(n17547) );
  AND2X1 U18367 ( .IN1(n10907), .IN2(g936), .Q(n17542) );
  OR2X1 U18368 ( .IN1(n17548), .IN2(n17549), .Q(g28055) );
  OR2X1 U18369 ( .IN1(n17550), .IN2(n17551), .Q(n17549) );
  AND2X1 U18370 ( .IN1(n17552), .IN2(n5728), .Q(n17551) );
  AND2X1 U18371 ( .IN1(n4519), .IN2(n16751), .Q(n17552) );
  AND2X1 U18372 ( .IN1(n17553), .IN2(g827), .Q(n17550) );
  AND2X1 U18373 ( .IN1(n4518), .IN2(n17554), .Q(n17553) );
  INVX0 U18374 ( .INP(n4519), .ZN(n17554) );
  AND2X1 U18375 ( .IN1(n10906), .IN2(g822), .Q(n17548) );
  OR2X1 U18376 ( .IN1(n17555), .IN2(n17556), .Q(g28054) );
  AND2X1 U18377 ( .IN1(n17557), .IN2(g661), .Q(n17556) );
  AND2X1 U18378 ( .IN1(n17558), .IN2(g728), .Q(n17555) );
  OR2X1 U18379 ( .IN1(n17559), .IN2(n17560), .Q(g28053) );
  OR2X1 U18380 ( .IN1(n17561), .IN2(n17562), .Q(n17560) );
  AND2X1 U18381 ( .IN1(n16813), .IN2(test_so87), .Q(n17562) );
  AND2X1 U18382 ( .IN1(n10906), .IN2(g681), .Q(n17559) );
  OR2X1 U18383 ( .IN1(n17563), .IN2(n17564), .Q(g28052) );
  AND2X1 U18384 ( .IN1(n17557), .IN2(g718), .Q(n17564) );
  AND2X1 U18385 ( .IN1(n17558), .IN2(g661), .Q(n17563) );
  OR2X1 U18386 ( .IN1(n17565), .IN2(n17566), .Q(g28051) );
  AND2X1 U18387 ( .IN1(n17557), .IN2(g655), .Q(n17566) );
  AND2X1 U18388 ( .IN1(n17558), .IN2(g718), .Q(n17565) );
  OR2X1 U18389 ( .IN1(n17567), .IN2(n17568), .Q(g28050) );
  AND2X1 U18390 ( .IN1(n17557), .IN2(g650), .Q(n17568) );
  AND2X1 U18391 ( .IN1(n17558), .IN2(g655), .Q(n17567) );
  OR2X1 U18392 ( .IN1(n17569), .IN2(n17570), .Q(g28049) );
  OR2X1 U18393 ( .IN1(n17571), .IN2(n17572), .Q(n17570) );
  AND2X1 U18394 ( .IN1(n17558), .IN2(g650), .Q(n17572) );
  AND2X1 U18395 ( .IN1(n17561), .IN2(g681), .Q(n17571) );
  AND2X1 U18396 ( .IN1(test_so87), .IN2(n10895), .Q(n17569) );
  OR2X1 U18397 ( .IN1(n17573), .IN2(n17574), .Q(g28048) );
  OR2X1 U18398 ( .IN1(n17575), .IN2(n17576), .Q(n17574) );
  AND2X1 U18399 ( .IN1(n17577), .IN2(n11073), .Q(n17576) );
  AND2X1 U18400 ( .IN1(n17578), .IN2(n17579), .Q(n11073) );
  AND2X1 U18401 ( .IN1(n5520), .IN2(n5112), .Q(n17579) );
  AND2X1 U18402 ( .IN1(g703), .IN2(n17580), .Q(n17578) );
  INVX0 U18403 ( .INP(n16778), .ZN(n17580) );
  OR2X1 U18404 ( .IN1(n17581), .IN2(n17582), .Q(n16778) );
  OR2X1 U18405 ( .IN1(n10582), .IN2(n17583), .Q(n17582) );
  XNOR2X1 U18406 ( .IN1(n10159), .IN2(g661), .Q(n17583) );
  OR2X1 U18407 ( .IN1(g645), .IN2(g650), .Q(n17581) );
  AND2X1 U18408 ( .IN1(n17584), .IN2(g691), .Q(n17575) );
  OR2X1 U18409 ( .IN1(n17585), .IN2(n17586), .Q(n17584) );
  AND2X1 U18410 ( .IN1(n17587), .IN2(n10780), .Q(n17585) );
  AND2X1 U18411 ( .IN1(g703), .IN2(n10580), .Q(n17587) );
  AND2X1 U18412 ( .IN1(n10906), .IN2(g29212), .Q(n17573) );
  OR2X1 U18413 ( .IN1(n17588), .IN2(n17589), .Q(g28047) );
  AND2X1 U18414 ( .IN1(n17557), .IN2(g645), .Q(n17589) );
  INVX0 U18415 ( .INP(n17558), .ZN(n17557) );
  AND2X1 U18416 ( .IN1(n17558), .IN2(g681), .Q(n17588) );
  OR2X1 U18417 ( .IN1(n17590), .IN2(n17591), .Q(g28046) );
  AND2X1 U18418 ( .IN1(n17558), .IN2(g645), .Q(n17591) );
  AND2X1 U18419 ( .IN1(n10817), .IN2(n17592), .Q(n17558) );
  AND2X1 U18420 ( .IN1(n17561), .IN2(g446), .Q(n17590) );
  AND2X1 U18421 ( .IN1(n10817), .IN2(n17593), .Q(n17561) );
  INVX0 U18422 ( .INP(n17592), .ZN(n17593) );
  OR2X1 U18423 ( .IN1(n17594), .IN2(n17595), .Q(n17592) );
  OR2X1 U18424 ( .IN1(n17596), .IN2(n17597), .Q(n17595) );
  AND2X1 U18425 ( .IN1(n5520), .IN2(n17598), .Q(n17597) );
  OR2X1 U18426 ( .IN1(g424), .IN2(n17599), .Q(n17598) );
  OR2X1 U18427 ( .IN1(n5358), .IN2(g411), .Q(n17599) );
  AND2X1 U18428 ( .IN1(n17600), .IN2(g691), .Q(n17596) );
  OR2X1 U18429 ( .IN1(n17601), .IN2(n17602), .Q(g28045) );
  OR2X1 U18430 ( .IN1(n17603), .IN2(n17604), .Q(n17602) );
  AND2X1 U18431 ( .IN1(n4537), .IN2(n5337), .Q(n17604) );
  AND2X1 U18432 ( .IN1(n17605), .IN2(g572), .Q(n17603) );
  AND2X1 U18433 ( .IN1(n2421), .IN2(n17606), .Q(n17605) );
  INVX0 U18434 ( .INP(n4537), .ZN(n17606) );
  AND2X1 U18435 ( .IN1(n10906), .IN2(g568), .Q(n17601) );
  OR2X1 U18436 ( .IN1(n17607), .IN2(n17608), .Q(g28044) );
  AND2X1 U18437 ( .IN1(n17609), .IN2(n10780), .Q(n17608) );
  OR2X1 U18438 ( .IN1(n4962), .IN2(n17610), .Q(n17609) );
  XNOR2X1 U18439 ( .IN1(n16794), .IN2(g482), .Q(n17610) );
  OR2X1 U18440 ( .IN1(n17611), .IN2(n17612), .Q(n16794) );
  AND2X1 U18441 ( .IN1(n5327), .IN2(n17613), .Q(n17611) );
  AND2X1 U18442 ( .IN1(n10906), .IN2(g528), .Q(n17607) );
  OR2X1 U18443 ( .IN1(n17614), .IN2(n17615), .Q(g28043) );
  AND2X1 U18444 ( .IN1(n10906), .IN2(g278), .Q(n17615) );
  AND2X1 U18445 ( .IN1(n10534), .IN2(n10558), .Q(n17614) );
  AND2X1 U18446 ( .IN1(n10817), .IN2(n14592), .Q(n10534) );
  INVX0 U18447 ( .INP(n14430), .ZN(n14592) );
  OR2X1 U18448 ( .IN1(n16078), .IN2(n17616), .Q(n14430) );
  OR2X1 U18449 ( .IN1(n17617), .IN2(n17618), .Q(n17616) );
  AND2X1 U18450 ( .IN1(n17619), .IN2(g278), .Q(n17618) );
  INVX0 U18451 ( .INP(n17620), .ZN(n17617) );
  OR2X1 U18452 ( .IN1(n5520), .IN2(n17621), .Q(n16078) );
  INVX0 U18453 ( .INP(n16757), .ZN(n17621) );
  OR2X1 U18454 ( .IN1(n17622), .IN2(n17623), .Q(n16757) );
  OR2X1 U18455 ( .IN1(n17624), .IN2(n17625), .Q(n17623) );
  AND2X1 U18456 ( .IN1(g554), .IN2(g807), .Q(n17624) );
  OR2X1 U18457 ( .IN1(n17626), .IN2(n17627), .Q(n17622) );
  AND2X1 U18458 ( .IN1(n17628), .IN2(n10189), .Q(n17627) );
  AND2X1 U18459 ( .IN1(n10188), .IN2(n10082), .Q(n17628) );
  AND2X1 U18460 ( .IN1(n17629), .IN2(g655), .Q(n17626) );
  AND2X1 U18461 ( .IN1(g753), .IN2(g718), .Q(n17629) );
  OR2X1 U18462 ( .IN1(g962), .IN2(n17630), .Q(g28042) );
  OR2X1 U18463 ( .IN1(n10880), .IN2(g1306), .Q(n17630) );
  OR2X1 U18464 ( .IN1(n13530), .IN2(n17631), .Q(g28041) );
  OR2X1 U18465 ( .IN1(n10879), .IN2(n13780), .Q(n17631) );
  AND2X1 U18466 ( .IN1(g1193), .IN2(n4837), .Q(n13780) );
  AND2X1 U18467 ( .IN1(n4836), .IN2(g1536), .Q(n13530) );
  OR2X1 U18468 ( .IN1(n17632), .IN2(n17633), .Q(g28030) );
  AND2X1 U18469 ( .IN1(n11696), .IN2(n11699), .Q(n17633) );
  AND2X1 U18470 ( .IN1(n17634), .IN2(n11698), .Q(n17632) );
  OR2X1 U18471 ( .IN1(n10880), .IN2(n17635), .Q(n11698) );
  AND2X1 U18472 ( .IN1(n5883), .IN2(n5871), .Q(n17635) );
  OR2X1 U18473 ( .IN1(n17636), .IN2(n17637), .Q(n17634) );
  AND2X1 U18474 ( .IN1(n11696), .IN2(n17638), .Q(n17637) );
  OR2X1 U18475 ( .IN1(n17639), .IN2(n17640), .Q(n17638) );
  AND2X1 U18476 ( .IN1(n17641), .IN2(n5882), .Q(n17639) );
  AND2X1 U18477 ( .IN1(n5861), .IN2(n17642), .Q(n17641) );
  OR2X1 U18478 ( .IN1(n17643), .IN2(n17644), .Q(n17642) );
  AND2X1 U18479 ( .IN1(n17645), .IN2(n17646), .Q(n11696) );
  OR2X1 U18480 ( .IN1(n17647), .IN2(n10876), .Q(n17645) );
  AND2X1 U18481 ( .IN1(n11699), .IN2(n17648), .Q(n17636) );
  OR2X1 U18482 ( .IN1(n17649), .IN2(n17646), .Q(n17648) );
  AND2X1 U18483 ( .IN1(n17650), .IN2(n17651), .Q(n17646) );
  AND2X1 U18484 ( .IN1(n17647), .IN2(n17652), .Q(n17649) );
  AND2X1 U18485 ( .IN1(n17653), .IN2(n17654), .Q(n17652) );
  OR2X1 U18486 ( .IN1(n17651), .IN2(n17650), .Q(n17654) );
  OR2X1 U18487 ( .IN1(n10880), .IN2(n17655), .Q(n17650) );
  AND2X1 U18488 ( .IN1(n5884), .IN2(n5870), .Q(n17655) );
  AND2X1 U18489 ( .IN1(n17656), .IN2(n17657), .Q(n17651) );
  OR2X1 U18490 ( .IN1(n17657), .IN2(n17656), .Q(n17653) );
  OR2X1 U18491 ( .IN1(n10881), .IN2(n17658), .Q(n17656) );
  AND2X1 U18492 ( .IN1(n5888), .IN2(n5874), .Q(n17658) );
  OR2X1 U18493 ( .IN1(n10881), .IN2(n17659), .Q(n17657) );
  AND2X1 U18494 ( .IN1(n5873), .IN2(n10593), .Q(n17659) );
  AND2X1 U18495 ( .IN1(n5885), .IN2(n5869), .Q(n17647) );
  AND2X1 U18496 ( .IN1(n17640), .IN2(n17660), .Q(n11699) );
  AND2X1 U18497 ( .IN1(n5861), .IN2(n5882), .Q(n17660) );
  AND2X1 U18498 ( .IN1(n17643), .IN2(n17644), .Q(n17640) );
  OR2X1 U18499 ( .IN1(n10882), .IN2(n17661), .Q(n17644) );
  AND2X1 U18500 ( .IN1(n5889), .IN2(n5868), .Q(n17661) );
  OR2X1 U18501 ( .IN1(n10882), .IN2(n17662), .Q(n17643) );
  AND2X1 U18502 ( .IN1(n5886), .IN2(n5872), .Q(n17662) );
  OR2X1 U18503 ( .IN1(n17663), .IN2(n17664), .Q(g26971) );
  AND2X1 U18504 ( .IN1(n17665), .IN2(n10780), .Q(n17664) );
  OR2X1 U18505 ( .IN1(n10486), .IN2(n5670), .Q(n17665) );
  AND2X1 U18506 ( .IN1(n10905), .IN2(g4512), .Q(n17663) );
  OR2X1 U18507 ( .IN1(n17666), .IN2(n17667), .Q(g26970) );
  AND2X1 U18508 ( .IN1(n10905), .IN2(g4459), .Q(n17667) );
  AND2X1 U18509 ( .IN1(n10818), .IN2(g4473), .Q(n17666) );
  OR2X1 U18510 ( .IN1(n17668), .IN2(n17669), .Q(g26969) );
  AND2X1 U18511 ( .IN1(n17670), .IN2(n10780), .Q(n17669) );
  AND2X1 U18512 ( .IN1(n10494), .IN2(n10566), .Q(n17670) );
  AND2X1 U18513 ( .IN1(n10905), .IN2(g4462), .Q(n17668) );
  OR2X1 U18514 ( .IN1(n17671), .IN2(n17672), .Q(g26968) );
  AND2X1 U18515 ( .IN1(n10905), .IN2(g4558), .Q(n17672) );
  OR2X1 U18516 ( .IN1(n17673), .IN2(n17674), .Q(g26967) );
  AND2X1 U18517 ( .IN1(n10905), .IN2(g4561), .Q(n17674) );
  OR2X1 U18518 ( .IN1(n17675), .IN2(n17676), .Q(g26966) );
  AND2X1 U18519 ( .IN1(n10905), .IN2(g4555), .Q(n17676) );
  XOR2X1 U18520 ( .IN1(n9348), .IN2(n17677), .Q(g26965) );
  AND2X1 U18521 ( .IN1(n10818), .IN2(g10306), .Q(n17677) );
  OR2X1 U18522 ( .IN1(n17678), .IN2(n17679), .Q(g26964) );
  AND2X1 U18523 ( .IN1(n17680), .IN2(n10780), .Q(n17679) );
  OR2X1 U18524 ( .IN1(n17681), .IN2(n17682), .Q(n17680) );
  AND2X1 U18525 ( .IN1(n5752), .IN2(n17258), .Q(n17682) );
  XOR2X1 U18526 ( .IN1(n12435), .IN2(g4527), .Q(n17258) );
  AND2X1 U18527 ( .IN1(n17683), .IN2(n17684), .Q(n12435) );
  AND2X1 U18528 ( .IN1(g4483), .IN2(test_so27), .Q(n17684) );
  AND2X1 U18529 ( .IN1(g4492), .IN2(g4489), .Q(n17683) );
  AND2X1 U18530 ( .IN1(g4515), .IN2(g4521), .Q(n17681) );
  AND2X1 U18531 ( .IN1(n10905), .IN2(g4527), .Q(n17678) );
  OR2X1 U18532 ( .IN1(n17673), .IN2(n17685), .Q(g26963) );
  AND2X1 U18533 ( .IN1(n10905), .IN2(g4489), .Q(n17685) );
  AND2X1 U18534 ( .IN1(g6750), .IN2(n10780), .Q(n17673) );
  OR2X1 U18535 ( .IN1(n17686), .IN2(n17671), .Q(g26962) );
  AND2X1 U18536 ( .IN1(g6749), .IN2(n10781), .Q(n17671) );
  AND2X1 U18537 ( .IN1(test_so27), .IN2(n10896), .Q(n17686) );
  OR2X1 U18538 ( .IN1(n17675), .IN2(n17687), .Q(g26961) );
  AND2X1 U18539 ( .IN1(n10905), .IN2(g4483), .Q(n17687) );
  AND2X1 U18540 ( .IN1(g6748), .IN2(n10781), .Q(n17675) );
  OR2X1 U18541 ( .IN1(n17688), .IN2(n17689), .Q(g26958) );
  AND2X1 U18542 ( .IN1(n10904), .IN2(g4455), .Q(n17688) );
  OR2X1 U18543 ( .IN1(n17690), .IN2(n17691), .Q(g26957) );
  AND2X1 U18544 ( .IN1(test_so47), .IN2(n10781), .Q(n17691) );
  AND2X1 U18545 ( .IN1(n17692), .IN2(g4434), .Q(n17690) );
  OR2X1 U18546 ( .IN1(n10883), .IN2(n17693), .Q(n17692) );
  AND2X1 U18547 ( .IN1(n17694), .IN2(g4392), .Q(n17693) );
  OR2X1 U18548 ( .IN1(n17695), .IN2(n9336), .Q(g26956) );
  AND2X1 U18549 ( .IN1(n17696), .IN2(n17697), .Q(n17695) );
  AND2X1 U18550 ( .IN1(n17694), .IN2(g4430), .Q(n17696) );
  OR2X1 U18551 ( .IN1(n17698), .IN2(n17699), .Q(g26955) );
  AND2X1 U18552 ( .IN1(n17700), .IN2(g4438), .Q(n17699) );
  AND2X1 U18553 ( .IN1(n17694), .IN2(n17701), .Q(n17698) );
  OR2X1 U18554 ( .IN1(n17702), .IN2(n17703), .Q(g26954) );
  OR2X1 U18555 ( .IN1(n17704), .IN2(n17705), .Q(n17703) );
  AND2X1 U18556 ( .IN1(n17706), .IN2(g4438), .Q(n17705) );
  AND2X1 U18557 ( .IN1(n17697), .IN2(n17694), .Q(n17704) );
  INVX0 U18558 ( .INP(n17707), .ZN(n17694) );
  OR2X1 U18559 ( .IN1(n17708), .IN2(n17709), .Q(n17707) );
  OR2X1 U18560 ( .IN1(g7260), .IN2(g7245), .Q(n17709) );
  OR2X1 U18561 ( .IN1(n9336), .IN2(n17710), .Q(n17708) );
  OR2X1 U18562 ( .IN1(test_so47), .IN2(g4438), .Q(n17710) );
  AND2X1 U18563 ( .IN1(test_so47), .IN2(n10896), .Q(n17702) );
  OR2X1 U18564 ( .IN1(n17711), .IN2(n17712), .Q(g26952) );
  AND2X1 U18565 ( .IN1(n17713), .IN2(n10781), .Q(n17712) );
  OR2X1 U18566 ( .IN1(n17714), .IN2(n17715), .Q(n17713) );
  XNOR2X1 U18567 ( .IN1(g4434), .IN2(n10080), .Q(n17715) );
  AND2X1 U18568 ( .IN1(n10083), .IN2(g4388), .Q(n17714) );
  AND2X1 U18569 ( .IN1(n17716), .IN2(g4430), .Q(n17711) );
  OR2X1 U18570 ( .IN1(n10482), .IN2(n10875), .Q(n17716) );
  OR2X1 U18571 ( .IN1(n17717), .IN2(g26953), .Q(g26951) );
  AND2X1 U18572 ( .IN1(n10904), .IN2(g4427), .Q(n17717) );
  OR2X1 U18573 ( .IN1(n17718), .IN2(n17689), .Q(g26950) );
  OR2X1 U18574 ( .IN1(n17719), .IN2(n17720), .Q(n17689) );
  AND2X1 U18575 ( .IN1(n17721), .IN2(n10781), .Q(n17720) );
  AND2X1 U18576 ( .IN1(n17701), .IN2(n17722), .Q(n17719) );
  AND2X1 U18577 ( .IN1(n10904), .IN2(g4417), .Q(n17718) );
  OR2X1 U18578 ( .IN1(n17723), .IN2(n17724), .Q(g26949) );
  AND2X1 U18579 ( .IN1(n10818), .IN2(g4411), .Q(n17724) );
  AND2X1 U18580 ( .IN1(n17725), .IN2(g4401), .Q(n17723) );
  OR2X1 U18581 ( .IN1(n10883), .IN2(n17726), .Q(n17725) );
  AND2X1 U18582 ( .IN1(n17727), .IN2(g4392), .Q(n17726) );
  OR2X1 U18583 ( .IN1(n17728), .IN2(g4405), .Q(g26948) );
  AND2X1 U18584 ( .IN1(n17729), .IN2(n17697), .Q(n17728) );
  AND2X1 U18585 ( .IN1(n17727), .IN2(g4388), .Q(n17729) );
  OR2X1 U18586 ( .IN1(n17730), .IN2(n17731), .Q(g26947) );
  OR2X1 U18587 ( .IN1(n17732), .IN2(n17733), .Q(n17731) );
  AND2X1 U18588 ( .IN1(n17734), .IN2(n10781), .Q(n17733) );
  OR2X1 U18589 ( .IN1(n17735), .IN2(n17721), .Q(n17734) );
  AND2X1 U18590 ( .IN1(n5710), .IN2(n17736), .Q(n17721) );
  AND2X1 U18591 ( .IN1(n17727), .IN2(n10007), .Q(n17736) );
  AND2X1 U18592 ( .IN1(n17737), .IN2(n10012), .Q(n17735) );
  AND2X1 U18593 ( .IN1(n17722), .IN2(g4382), .Q(n17737) );
  AND2X1 U18594 ( .IN1(n10904), .IN2(g4388), .Q(n17732) );
  OR2X1 U18595 ( .IN1(n17738), .IN2(n17739), .Q(g26946) );
  AND2X1 U18596 ( .IN1(n17700), .IN2(g4375), .Q(n17739) );
  INVX0 U18597 ( .INP(n17706), .ZN(n17700) );
  AND2X1 U18598 ( .IN1(n17727), .IN2(n17701), .Q(n17738) );
  AND2X1 U18599 ( .IN1(g4392), .IN2(n10781), .Q(n17701) );
  OR2X1 U18600 ( .IN1(n17740), .IN2(n17741), .Q(g26945) );
  OR2X1 U18601 ( .IN1(n17742), .IN2(n17730), .Q(n17741) );
  AND2X1 U18602 ( .IN1(n17706), .IN2(g4375), .Q(n17730) );
  AND2X1 U18603 ( .IN1(n10819), .IN2(n5714), .Q(n17706) );
  AND2X1 U18604 ( .IN1(n17697), .IN2(n17727), .Q(n17742) );
  INVX0 U18605 ( .INP(n17722), .ZN(n17727) );
  OR2X1 U18606 ( .IN1(n17743), .IN2(n17744), .Q(n17722) );
  OR2X1 U18607 ( .IN1(g7257), .IN2(g7243), .Q(n17744) );
  OR2X1 U18608 ( .IN1(g4411), .IN2(n17745), .Q(n17743) );
  OR2X1 U18609 ( .IN1(g4405), .IN2(g4375), .Q(n17745) );
  AND2X1 U18610 ( .IN1(n10819), .IN2(n5710), .Q(n17697) );
  AND2X1 U18611 ( .IN1(n10904), .IN2(g4411), .Q(n17740) );
  AND2X1 U18612 ( .IN1(n17746), .IN2(n10781), .Q(g26944) );
  OR2X1 U18613 ( .IN1(n17747), .IN2(n17748), .Q(n17746) );
  OR2X1 U18614 ( .IN1(n17256), .IN2(n17749), .Q(n17748) );
  OR2X1 U18615 ( .IN1(n12282), .IN2(n10552), .Q(n17749) );
  INVX0 U18616 ( .INP(n11934), .ZN(n12282) );
  OR2X1 U18617 ( .IN1(n17750), .IN2(g135), .Q(n17256) );
  AND2X1 U18618 ( .IN1(n17751), .IN2(n17752), .Q(n17750) );
  OR2X1 U18619 ( .IN1(n17753), .IN2(n17754), .Q(n17752) );
  OR2X1 U18620 ( .IN1(g4616), .IN2(n17755), .Q(n17754) );
  XNOR2X1 U18621 ( .IN1(g4601), .IN2(n5303), .Q(n17755) );
  XNOR2X1 U18622 ( .IN1(g4584), .IN2(n5274), .Q(n17753) );
  AND2X1 U18623 ( .IN1(n17756), .IN2(n17757), .Q(n17751) );
  OR2X1 U18624 ( .IN1(n5539), .IN2(n17758), .Q(n17757) );
  OR2X1 U18625 ( .IN1(g4608), .IN2(n17759), .Q(n17758) );
  OR2X1 U18626 ( .IN1(n5303), .IN2(g4601), .Q(n17759) );
  OR2X1 U18627 ( .IN1(g4584), .IN2(n17760), .Q(n17756) );
  OR2X1 U18628 ( .IN1(n5274), .IN2(g4593), .Q(n17760) );
  OR2X1 U18629 ( .IN1(n5348), .IN2(n17761), .Q(n17747) );
  OR2X1 U18630 ( .IN1(n5844), .IN2(n5653), .Q(n17761) );
  OR2X1 U18631 ( .IN1(n17762), .IN2(n17763), .Q(g26940) );
  AND2X1 U18632 ( .IN1(n15273), .IN2(n10781), .Q(n17763) );
  OR2X1 U18633 ( .IN1(n17764), .IN2(n17765), .Q(n15273) );
  AND2X1 U18634 ( .IN1(g114), .IN2(n5983), .Q(n17765) );
  AND2X1 U18635 ( .IN1(g116), .IN2(g4157), .Q(n17764) );
  AND2X1 U18636 ( .IN1(n10904), .IN2(g4153), .Q(n17762) );
  OR2X1 U18637 ( .IN1(n17766), .IN2(n17767), .Q(g26939) );
  AND2X1 U18638 ( .IN1(n15275), .IN2(n10782), .Q(n17767) );
  OR2X1 U18639 ( .IN1(n17768), .IN2(n17769), .Q(n15275) );
  AND2X1 U18640 ( .IN1(g120), .IN2(n5981), .Q(n17769) );
  AND2X1 U18641 ( .IN1(g124), .IN2(g4146), .Q(n17768) );
  AND2X1 U18642 ( .IN1(n10904), .IN2(g4104), .Q(n17766) );
  OR2X1 U18643 ( .IN1(n10542), .IN2(n17770), .Q(g26938) );
  OR2X1 U18644 ( .IN1(n17771), .IN2(n17772), .Q(n17770) );
  AND2X1 U18645 ( .IN1(n17773), .IN2(n10782), .Q(n17772) );
  XNOR2X1 U18646 ( .IN1(n17296), .IN2(g4082), .Q(n17773) );
  OR2X1 U18647 ( .IN1(n5612), .IN2(n4723), .Q(n17296) );
  INVX0 U18648 ( .INP(n17774), .ZN(n4723) );
  AND2X1 U18649 ( .IN1(n10904), .IN2(g4141), .Q(n17771) );
  OR2X1 U18650 ( .IN1(n17775), .IN2(n17776), .Q(g26934) );
  OR2X1 U18651 ( .IN1(n17777), .IN2(n17778), .Q(n17776) );
  AND2X1 U18652 ( .IN1(test_so37), .IN2(n10896), .Q(n17778) );
  AND2X1 U18653 ( .IN1(n17779), .IN2(n10589), .Q(n17777) );
  AND2X1 U18654 ( .IN1(n4888), .IN2(g2827), .Q(n17775) );
  OR2X1 U18655 ( .IN1(n17780), .IN2(n17781), .Q(g26933) );
  OR2X1 U18656 ( .IN1(n17782), .IN2(n17783), .Q(n17781) );
  AND2X1 U18657 ( .IN1(n10904), .IN2(g2811), .Q(n17783) );
  AND2X1 U18658 ( .IN1(n5840), .IN2(n17779), .Q(n17782) );
  AND2X1 U18659 ( .IN1(test_so37), .IN2(n4888), .Q(n17780) );
  OR2X1 U18660 ( .IN1(n17784), .IN2(n17785), .Q(g26932) );
  OR2X1 U18661 ( .IN1(n17786), .IN2(n17787), .Q(n17785) );
  AND2X1 U18662 ( .IN1(n10903), .IN2(g2799), .Q(n17787) );
  AND2X1 U18663 ( .IN1(n5841), .IN2(n17779), .Q(n17786) );
  AND2X1 U18664 ( .IN1(n4888), .IN2(g2811), .Q(n17784) );
  OR2X1 U18665 ( .IN1(n17788), .IN2(n17789), .Q(g26931) );
  OR2X1 U18666 ( .IN1(n17790), .IN2(n17791), .Q(n17789) );
  AND2X1 U18667 ( .IN1(n10903), .IN2(g29219), .Q(n17791) );
  AND2X1 U18668 ( .IN1(n5839), .IN2(n17779), .Q(n17790) );
  AND2X1 U18669 ( .IN1(n4888), .IN2(g2799), .Q(n17788) );
  OR2X1 U18670 ( .IN1(n17792), .IN2(n17793), .Q(g26930) );
  OR2X1 U18671 ( .IN1(n17794), .IN2(n17795), .Q(n17793) );
  AND2X1 U18672 ( .IN1(n10903), .IN2(g2791), .Q(n17795) );
  AND2X1 U18673 ( .IN1(n17779), .IN2(n10590), .Q(n17794) );
  AND2X1 U18674 ( .IN1(n4888), .IN2(g2795), .Q(n17792) );
  OR2X1 U18675 ( .IN1(n17796), .IN2(n17797), .Q(g26929) );
  OR2X1 U18676 ( .IN1(n17798), .IN2(n17799), .Q(n17797) );
  AND2X1 U18677 ( .IN1(n10903), .IN2(g2779), .Q(n17799) );
  AND2X1 U18678 ( .IN1(n5837), .IN2(n17779), .Q(n17798) );
  AND2X1 U18679 ( .IN1(n4888), .IN2(g2791), .Q(n17796) );
  OR2X1 U18680 ( .IN1(n17800), .IN2(n17801), .Q(g26928) );
  OR2X1 U18681 ( .IN1(n17802), .IN2(n17803), .Q(n17801) );
  AND2X1 U18682 ( .IN1(n10903), .IN2(g2767), .Q(n17803) );
  AND2X1 U18683 ( .IN1(n5834), .IN2(n17779), .Q(n17802) );
  AND2X1 U18684 ( .IN1(n4888), .IN2(g2779), .Q(n17800) );
  OR2X1 U18685 ( .IN1(n17804), .IN2(n17805), .Q(g26927) );
  OR2X1 U18686 ( .IN1(n17806), .IN2(n17807), .Q(n17805) );
  AND2X1 U18687 ( .IN1(n10903), .IN2(g2763), .Q(n17807) );
  AND2X1 U18688 ( .IN1(n5836), .IN2(n17779), .Q(n17806) );
  AND2X1 U18689 ( .IN1(n4888), .IN2(n17808), .Q(n17779) );
  AND2X1 U18690 ( .IN1(n12043), .IN2(n11197), .Q(n17808) );
  OR2X1 U18691 ( .IN1(test_so30), .IN2(g2748), .Q(n11197) );
  INVX0 U18692 ( .INP(n12072), .ZN(n12043) );
  AND2X1 U18693 ( .IN1(test_so30), .IN2(n17809), .Q(n12072) );
  AND2X1 U18694 ( .IN1(g2735), .IN2(n1284), .Q(n17809) );
  AND2X1 U18695 ( .IN1(g2748), .IN2(g2741), .Q(n1284) );
  AND2X1 U18696 ( .IN1(n4888), .IN2(g2767), .Q(n17804) );
  OR2X1 U18697 ( .IN1(n17810), .IN2(n17811), .Q(g26926) );
  AND2X1 U18698 ( .IN1(n10903), .IN2(g2719), .Q(n17811) );
  AND2X1 U18699 ( .IN1(n17812), .IN2(n3730), .Q(n17810) );
  XNOR2X1 U18700 ( .IN1(n15677), .IN2(n5301), .Q(n17812) );
  AND2X1 U18701 ( .IN1(g2715), .IN2(g2719), .Q(n15677) );
  OR2X1 U18702 ( .IN1(n17813), .IN2(n17814), .Q(g26925) );
  AND2X1 U18703 ( .IN1(n17815), .IN2(n10782), .Q(n17814) );
  OR2X1 U18704 ( .IN1(n17816), .IN2(n4173), .Q(n17815) );
  AND2X1 U18705 ( .IN1(n15983), .IN2(g1536), .Q(n17816) );
  OR2X1 U18706 ( .IN1(n10528), .IN2(n15985), .Q(n15983) );
  INVX0 U18707 ( .INP(n17817), .ZN(n15985) );
  AND2X1 U18708 ( .IN1(g1542), .IN2(n15993), .Q(n17817) );
  AND2X1 U18709 ( .IN1(n13468), .IN2(n17818), .Q(n15993) );
  AND2X1 U18710 ( .IN1(g7946), .IN2(n16004), .Q(n17818) );
  OR2X1 U18711 ( .IN1(g1532), .IN2(n17819), .Q(n16004) );
  OR2X1 U18712 ( .IN1(n5577), .IN2(n5381), .Q(n17819) );
  AND2X1 U18713 ( .IN1(n10903), .IN2(g1532), .Q(n17813) );
  OR2X1 U18714 ( .IN1(n17820), .IN2(n17821), .Q(g26924) );
  OR2X1 U18715 ( .IN1(n17822), .IN2(n17823), .Q(n17821) );
  AND2X1 U18716 ( .IN1(n10903), .IN2(g1437), .Q(n17823) );
  AND2X1 U18717 ( .IN1(n17824), .IN2(n10782), .Q(n17822) );
  AND2X1 U18718 ( .IN1(n17825), .IN2(g1478), .Q(n17824) );
  INVX0 U18719 ( .INP(n17826), .ZN(n17820) );
  OR2X1 U18720 ( .IN1(n17825), .IN2(g1478), .Q(n17826) );
  OR2X1 U18721 ( .IN1(n17827), .IN2(n17828), .Q(n17825) );
  OR2X1 U18722 ( .IN1(n5696), .IN2(n16687), .Q(n17828) );
  OR2X1 U18723 ( .IN1(n10474), .IN2(n17829), .Q(n16687) );
  OR2X1 U18724 ( .IN1(test_so49), .IN2(n5364), .Q(n17829) );
  OR2X1 U18725 ( .IN1(n17830), .IN2(n17831), .Q(g26923) );
  OR2X1 U18726 ( .IN1(n17832), .IN2(n17833), .Q(n17831) );
  AND2X1 U18727 ( .IN1(n10903), .IN2(g1467), .Q(n17833) );
  AND2X1 U18728 ( .IN1(n17834), .IN2(n10782), .Q(n17832) );
  AND2X1 U18729 ( .IN1(n17835), .IN2(g1472), .Q(n17834) );
  INVX0 U18730 ( .INP(n17836), .ZN(n17830) );
  OR2X1 U18731 ( .IN1(n17835), .IN2(g1472), .Q(n17836) );
  OR2X1 U18732 ( .IN1(n17837), .IN2(n17838), .Q(n17835) );
  OR2X1 U18733 ( .IN1(n16675), .IN2(n17827), .Q(n17838) );
  OR2X1 U18734 ( .IN1(n5693), .IN2(n10474), .Q(n17837) );
  OR2X1 U18735 ( .IN1(n17839), .IN2(n17840), .Q(g26922) );
  OR2X1 U18736 ( .IN1(n17841), .IN2(n17842), .Q(n17840) );
  AND2X1 U18737 ( .IN1(n10903), .IN2(g1454), .Q(n17842) );
  AND2X1 U18738 ( .IN1(n17843), .IN2(n10782), .Q(n17841) );
  AND2X1 U18739 ( .IN1(n17844), .IN2(g1448), .Q(n17843) );
  INVX0 U18740 ( .INP(n17845), .ZN(n17839) );
  OR2X1 U18741 ( .IN1(n17844), .IN2(g1448), .Q(n17845) );
  OR2X1 U18742 ( .IN1(n17827), .IN2(n17846), .Q(n17844) );
  OR2X1 U18743 ( .IN1(n5866), .IN2(n16654), .Q(n17846) );
  INVX0 U18744 ( .INP(n16657), .ZN(n16654) );
  AND2X1 U18745 ( .IN1(g13272), .IN2(n13468), .Q(n16657) );
  AND2X1 U18746 ( .IN1(test_so49), .IN2(n5364), .Q(n13468) );
  OR2X1 U18747 ( .IN1(n17847), .IN2(n17848), .Q(g26921) );
  AND2X1 U18748 ( .IN1(n17849), .IN2(n10782), .Q(n17848) );
  AND2X1 U18749 ( .IN1(n17850), .IN2(n10550), .Q(n17849) );
  XOR2X1 U18750 ( .IN1(n17851), .IN2(n10500), .Q(n17850) );
  AND2X1 U18751 ( .IN1(n10902), .IN2(g1395), .Q(n17847) );
  OR2X1 U18752 ( .IN1(n17852), .IN2(n17853), .Q(g26920) );
  OR2X1 U18753 ( .IN1(n17854), .IN2(n17855), .Q(n17853) );
  AND2X1 U18754 ( .IN1(n17856), .IN2(n10782), .Q(n17855) );
  INVX0 U18755 ( .INP(n17857), .ZN(n17856) );
  OR2X1 U18756 ( .IN1(n4915), .IN2(n10460), .Q(n17857) );
  AND2X1 U18757 ( .IN1(n17858), .IN2(n17859), .Q(n4915) );
  OR2X1 U18758 ( .IN1(g1384), .IN2(n5322), .Q(n17858) );
  AND2X1 U18759 ( .IN1(n10902), .IN2(g1384), .Q(n17854) );
  AND2X1 U18760 ( .IN1(n4913), .IN2(n17860), .Q(n17852) );
  OR2X1 U18761 ( .IN1(n17861), .IN2(n17862), .Q(g26919) );
  OR2X1 U18762 ( .IN1(n17863), .IN2(n17864), .Q(n17862) );
  INVX0 U18763 ( .INP(n17865), .ZN(n17864) );
  OR2X1 U18764 ( .IN1(n11220), .IN2(test_so77), .Q(n17865) );
  AND2X1 U18765 ( .IN1(n17866), .IN2(n11220), .Q(n17863) );
  OR2X1 U18766 ( .IN1(n10133), .IN2(n17867), .Q(n11220) );
  OR2X1 U18767 ( .IN1(n5655), .IN2(n10512), .Q(n17867) );
  AND2X1 U18768 ( .IN1(test_so77), .IN2(n17868), .Q(n17866) );
  AND2X1 U18769 ( .IN1(n10902), .IN2(g1266), .Q(n17861) );
  OR2X1 U18770 ( .IN1(n17869), .IN2(n17870), .Q(g26918) );
  AND2X1 U18771 ( .IN1(n17871), .IN2(n10782), .Q(n17870) );
  OR2X1 U18772 ( .IN1(n17872), .IN2(n4191), .Q(n17871) );
  AND2X1 U18773 ( .IN1(n16024), .IN2(g1193), .Q(n17872) );
  OR2X1 U18774 ( .IN1(n10529), .IN2(n16026), .Q(n16024) );
  INVX0 U18775 ( .INP(n17873), .ZN(n16026) );
  AND2X1 U18776 ( .IN1(g1199), .IN2(n16034), .Q(n17873) );
  AND2X1 U18777 ( .IN1(n13720), .IN2(n17874), .Q(n16034) );
  AND2X1 U18778 ( .IN1(g7916), .IN2(n16045), .Q(n17874) );
  OR2X1 U18779 ( .IN1(g1189), .IN2(n17875), .Q(n16045) );
  OR2X1 U18780 ( .IN1(n10138), .IN2(n10137), .Q(n17875) );
  AND2X1 U18781 ( .IN1(n10902), .IN2(g1189), .Q(n17869) );
  OR2X1 U18782 ( .IN1(n17876), .IN2(n17877), .Q(g26917) );
  OR2X1 U18783 ( .IN1(n17878), .IN2(n17879), .Q(n17877) );
  AND2X1 U18784 ( .IN1(n10902), .IN2(g1094), .Q(n17879) );
  AND2X1 U18785 ( .IN1(n17880), .IN2(n10783), .Q(n17878) );
  AND2X1 U18786 ( .IN1(n17881), .IN2(g1135), .Q(n17880) );
  INVX0 U18787 ( .INP(n17882), .ZN(n17876) );
  OR2X1 U18788 ( .IN1(n17881), .IN2(g1135), .Q(n17882) );
  OR2X1 U18789 ( .IN1(n17883), .IN2(n17884), .Q(n17881) );
  OR2X1 U18790 ( .IN1(n5697), .IN2(n16736), .Q(n17884) );
  OR2X1 U18791 ( .IN1(g1183), .IN2(n17885), .Q(n16736) );
  OR2X1 U18792 ( .IN1(n5363), .IN2(n10475), .Q(n17885) );
  OR2X1 U18793 ( .IN1(n17886), .IN2(n17887), .Q(g26916) );
  OR2X1 U18794 ( .IN1(n17888), .IN2(n17889), .Q(n17887) );
  AND2X1 U18795 ( .IN1(n10902), .IN2(g1124), .Q(n17889) );
  AND2X1 U18796 ( .IN1(n17890), .IN2(n10783), .Q(n17888) );
  AND2X1 U18797 ( .IN1(n17891), .IN2(g1129), .Q(n17890) );
  INVX0 U18798 ( .INP(n17892), .ZN(n17886) );
  OR2X1 U18799 ( .IN1(n17891), .IN2(g1129), .Q(n17892) );
  OR2X1 U18800 ( .IN1(n17883), .IN2(n17893), .Q(n17891) );
  OR2X1 U18801 ( .IN1(n5692), .IN2(n16726), .Q(n17893) );
  OR2X1 U18802 ( .IN1(n10475), .IN2(n17894), .Q(n16726) );
  OR2X1 U18803 ( .IN1(n17895), .IN2(n17896), .Q(g26915) );
  OR2X1 U18804 ( .IN1(n17897), .IN2(n17898), .Q(n17896) );
  AND2X1 U18805 ( .IN1(test_so90), .IN2(n10896), .Q(n17898) );
  AND2X1 U18806 ( .IN1(n17899), .IN2(n10783), .Q(n17897) );
  AND2X1 U18807 ( .IN1(n17900), .IN2(g1105), .Q(n17899) );
  INVX0 U18808 ( .INP(n17901), .ZN(n17900) );
  AND2X1 U18809 ( .IN1(n17901), .IN2(n5478), .Q(n17895) );
  AND2X1 U18810 ( .IN1(n17902), .IN2(n17903), .Q(n17901) );
  AND2X1 U18811 ( .IN1(n16705), .IN2(test_so90), .Q(n17903) );
  AND2X1 U18812 ( .IN1(g13259), .IN2(n13720), .Q(n16705) );
  AND2X1 U18813 ( .IN1(g1183), .IN2(n5363), .Q(n13720) );
  OR2X1 U18814 ( .IN1(n17904), .IN2(n17905), .Q(g26914) );
  AND2X1 U18815 ( .IN1(n17906), .IN2(n10783), .Q(n17905) );
  AND2X1 U18816 ( .IN1(n5320), .IN2(n17907), .Q(n17906) );
  XOR2X1 U18817 ( .IN1(n17908), .IN2(n10499), .Q(n17907) );
  AND2X1 U18818 ( .IN1(n10902), .IN2(g1052), .Q(n17904) );
  OR2X1 U18819 ( .IN1(n17909), .IN2(n17910), .Q(g26913) );
  OR2X1 U18820 ( .IN1(n17911), .IN2(n17912), .Q(n17910) );
  AND2X1 U18821 ( .IN1(n17913), .IN2(n10783), .Q(n17912) );
  INVX0 U18822 ( .INP(n17914), .ZN(n17913) );
  OR2X1 U18823 ( .IN1(n4940), .IN2(n10452), .Q(n17914) );
  AND2X1 U18824 ( .IN1(n17915), .IN2(n17916), .Q(n4940) );
  OR2X1 U18825 ( .IN1(g1041), .IN2(n5321), .Q(n17915) );
  AND2X1 U18826 ( .IN1(n10906), .IN2(g1041), .Q(n17911) );
  AND2X1 U18827 ( .IN1(n4938), .IN2(n17917), .Q(n17909) );
  OR2X1 U18828 ( .IN1(n17918), .IN2(n17919), .Q(g26912) );
  OR2X1 U18829 ( .IN1(n17920), .IN2(n17921), .Q(n17919) );
  AND2X1 U18830 ( .IN1(n251), .IN2(n5557), .Q(n17921) );
  INVX0 U18831 ( .INP(n17922), .ZN(n251) );
  AND2X1 U18832 ( .IN1(n17923), .IN2(g936), .Q(n17920) );
  AND2X1 U18833 ( .IN1(n17924), .IN2(n17922), .Q(n17923) );
  OR2X1 U18834 ( .IN1(n10132), .IN2(n17925), .Q(n17922) );
  OR2X1 U18835 ( .IN1(n5654), .IN2(n10513), .Q(n17925) );
  AND2X1 U18836 ( .IN1(n10899), .IN2(g921), .Q(n17918) );
  XNOR2X1 U18837 ( .IN1(n5682), .IN2(n17926), .Q(g26910) );
  AND2X1 U18838 ( .IN1(n5305), .IN2(n10783), .Q(n17926) );
  OR2X1 U18839 ( .IN1(n17927), .IN2(n17928), .Q(g26909) );
  AND2X1 U18840 ( .IN1(n17929), .IN2(n10783), .Q(n17928) );
  OR2X1 U18841 ( .IN1(n17930), .IN2(n17931), .Q(n17929) );
  AND2X1 U18842 ( .IN1(n5305), .IN2(g896), .Q(n17931) );
  AND2X1 U18843 ( .IN1(n5431), .IN2(g862), .Q(n17930) );
  AND2X1 U18844 ( .IN1(n10903), .IN2(g890), .Q(n17927) );
  OR2X1 U18845 ( .IN1(n17932), .IN2(n17933), .Q(g26908) );
  OR2X1 U18846 ( .IN1(n17934), .IN2(n17935), .Q(n17933) );
  AND2X1 U18847 ( .IN1(n10903), .IN2(g246), .Q(n17935) );
  AND2X1 U18848 ( .IN1(n17936), .IN2(g872), .Q(n17934) );
  AND2X1 U18849 ( .IN1(n4945), .IN2(g446), .Q(n17932) );
  OR2X1 U18850 ( .IN1(n17937), .IN2(n17938), .Q(g26907) );
  OR2X1 U18851 ( .IN1(n17939), .IN2(n17940), .Q(n17938) );
  AND2X1 U18852 ( .IN1(n10903), .IN2(g269), .Q(n17940) );
  AND2X1 U18853 ( .IN1(n17936), .IN2(g14167), .Q(n17939) );
  AND2X1 U18854 ( .IN1(n4945), .IN2(g246), .Q(n17937) );
  OR2X1 U18855 ( .IN1(n17941), .IN2(n17942), .Q(g26906) );
  OR2X1 U18856 ( .IN1(n17943), .IN2(n17944), .Q(n17942) );
  AND2X1 U18857 ( .IN1(n10903), .IN2(g239), .Q(n17944) );
  AND2X1 U18858 ( .IN1(n17936), .IN2(g14147), .Q(n17943) );
  AND2X1 U18859 ( .IN1(n4945), .IN2(g269), .Q(n17941) );
  OR2X1 U18860 ( .IN1(n17945), .IN2(n17946), .Q(g26905) );
  OR2X1 U18861 ( .IN1(n17947), .IN2(n17948), .Q(n17946) );
  AND2X1 U18862 ( .IN1(n10903), .IN2(g262), .Q(n17948) );
  AND2X1 U18863 ( .IN1(n17936), .IN2(g14125), .Q(n17947) );
  AND2X1 U18864 ( .IN1(n4945), .IN2(g239), .Q(n17945) );
  OR2X1 U18865 ( .IN1(n17949), .IN2(n17950), .Q(g26904) );
  OR2X1 U18866 ( .IN1(n17951), .IN2(n17952), .Q(n17950) );
  AND2X1 U18867 ( .IN1(n10903), .IN2(g232), .Q(n17952) );
  AND2X1 U18868 ( .IN1(n17936), .IN2(g14096), .Q(n17951) );
  AND2X1 U18869 ( .IN1(n4945), .IN2(g262), .Q(n17949) );
  OR2X1 U18870 ( .IN1(n17953), .IN2(n17954), .Q(g26903) );
  OR2X1 U18871 ( .IN1(n17955), .IN2(n17956), .Q(n17954) );
  AND2X1 U18872 ( .IN1(n10903), .IN2(g255), .Q(n17956) );
  AND2X1 U18873 ( .IN1(n17936), .IN2(g14217), .Q(n17955) );
  AND2X1 U18874 ( .IN1(n4945), .IN2(g232), .Q(n17953) );
  OR2X1 U18875 ( .IN1(n17957), .IN2(n17958), .Q(g26902) );
  OR2X1 U18876 ( .IN1(n17959), .IN2(n17960), .Q(n17958) );
  AND2X1 U18877 ( .IN1(n10903), .IN2(g225), .Q(n17960) );
  AND2X1 U18878 ( .IN1(n17936), .IN2(g14201), .Q(n17959) );
  AND2X1 U18879 ( .IN1(n4945), .IN2(g255), .Q(n17957) );
  OR2X1 U18880 ( .IN1(n17961), .IN2(n17962), .Q(g26901) );
  OR2X1 U18881 ( .IN1(n17963), .IN2(n17964), .Q(n17962) );
  AND2X1 U18882 ( .IN1(n10904), .IN2(g872), .Q(n17964) );
  AND2X1 U18883 ( .IN1(n17936), .IN2(g14189), .Q(n17963) );
  AND2X1 U18884 ( .IN1(n17965), .IN2(n10783), .Q(n17936) );
  INVX0 U18885 ( .INP(n4946), .ZN(n17965) );
  OR2X1 U18886 ( .IN1(g862), .IN2(n17966), .Q(n4946) );
  OR2X1 U18887 ( .IN1(n5305), .IN2(g896), .Q(n17966) );
  AND2X1 U18888 ( .IN1(n4945), .IN2(g225), .Q(n17961) );
  OR2X1 U18889 ( .IN1(n17967), .IN2(n17968), .Q(g26899) );
  AND2X1 U18890 ( .IN1(n10904), .IN2(g832), .Q(n17968) );
  AND2X1 U18891 ( .IN1(n17969), .IN2(n4518), .Q(n17967) );
  XNOR2X1 U18892 ( .IN1(n4814), .IN2(n5422), .Q(n17969) );
  AND2X1 U18893 ( .IN1(n4948), .IN2(n17970), .Q(n4814) );
  AND2X1 U18894 ( .IN1(g817), .IN2(g832), .Q(n17970) );
  OR2X1 U18895 ( .IN1(n17971), .IN2(n17972), .Q(g26898) );
  AND2X1 U18896 ( .IN1(n10904), .IN2(g843), .Q(n17972) );
  AND2X1 U18897 ( .IN1(n17973), .IN2(g837), .Q(n17971) );
  AND2X1 U18898 ( .IN1(n17974), .IN2(n17975), .Q(n17973) );
  OR2X1 U18899 ( .IN1(n17976), .IN2(g812), .Q(n17975) );
  AND2X1 U18900 ( .IN1(n17977), .IN2(g843), .Q(n17976) );
  OR2X1 U18901 ( .IN1(n5733), .IN2(n17978), .Q(n17974) );
  OR2X1 U18902 ( .IN1(n16813), .IN2(n17979), .Q(n17978) );
  AND2X1 U18903 ( .IN1(n17980), .IN2(n10783), .Q(n17979) );
  OR2X1 U18904 ( .IN1(n10109), .IN2(n5709), .Q(n17980) );
  OR2X1 U18905 ( .IN1(n17981), .IN2(n17982), .Q(g26897) );
  INVX0 U18906 ( .INP(n17983), .ZN(n17982) );
  OR2X1 U18907 ( .IN1(n17984), .IN2(n5732), .Q(n17983) );
  AND2X1 U18908 ( .IN1(n17984), .IN2(g753), .Q(n17981) );
  AND2X1 U18909 ( .IN1(n10820), .IN2(n17625), .Q(n17984) );
  OR2X1 U18910 ( .IN1(n17985), .IN2(n17986), .Q(g26896) );
  OR2X1 U18911 ( .IN1(n17987), .IN2(n17988), .Q(n17986) );
  AND2X1 U18912 ( .IN1(n17989), .IN2(g728), .Q(n17988) );
  INVX0 U18913 ( .INP(n17990), .ZN(n17987) );
  OR2X1 U18914 ( .IN1(n17989), .IN2(n5657), .Q(n17990) );
  OR2X1 U18915 ( .IN1(n10883), .IN2(n16779), .Q(n17989) );
  AND2X1 U18916 ( .IN1(n4956), .IN2(n16779), .Q(n17985) );
  INVX0 U18917 ( .INP(n120), .ZN(n16779) );
  OR2X1 U18918 ( .IN1(n17991), .IN2(n17992), .Q(n120) );
  OR2X1 U18919 ( .IN1(g504), .IN2(n10581), .Q(n17992) );
  OR2X1 U18920 ( .IN1(n17613), .IN2(n17993), .Q(n17991) );
  OR2X1 U18921 ( .IN1(g528), .IN2(n17994), .Q(n17993) );
  OR2X1 U18922 ( .IN1(n17995), .IN2(n17996), .Q(g26895) );
  OR2X1 U18923 ( .IN1(n17997), .IN2(n17998), .Q(n17996) );
  AND2X1 U18924 ( .IN1(n4826), .IN2(n5335), .Q(n17998) );
  AND2X1 U18925 ( .IN1(n17999), .IN2(g568), .Q(n17997) );
  AND2X1 U18926 ( .IN1(n2421), .IN2(n18000), .Q(n17999) );
  INVX0 U18927 ( .INP(n4826), .ZN(n18000) );
  AND2X1 U18928 ( .IN1(n4959), .IN2(n18001), .Q(n4826) );
  AND2X1 U18929 ( .IN1(g562), .IN2(n18002), .Q(n18001) );
  INVX0 U18930 ( .INP(n18003), .ZN(n18002) );
  AND2X1 U18931 ( .IN1(n10904), .IN2(g562), .Q(n17995) );
  OR2X1 U18932 ( .IN1(n18004), .IN2(n18005), .Q(g26894) );
  AND2X1 U18933 ( .IN1(n18006), .IN2(n10784), .Q(n18005) );
  AND2X1 U18934 ( .IN1(n18007), .IN2(n18008), .Q(n18006) );
  AND2X1 U18935 ( .IN1(n18009), .IN2(n18010), .Q(n18007) );
  OR2X1 U18936 ( .IN1(n5327), .IN2(n17612), .Q(n18010) );
  OR2X1 U18937 ( .IN1(n18011), .IN2(g528), .Q(n18009) );
  AND2X1 U18938 ( .IN1(n18012), .IN2(n17613), .Q(n18011) );
  OR2X1 U18939 ( .IN1(n5708), .IN2(n5820), .Q(n17613) );
  INVX0 U18940 ( .INP(n17612), .ZN(n18012) );
  OR2X1 U18941 ( .IN1(n18013), .IN2(n18014), .Q(n17612) );
  OR2X1 U18942 ( .IN1(n5287), .IN2(g513), .Q(n18014) );
  AND2X1 U18943 ( .IN1(n10904), .IN2(g518), .Q(n18004) );
  OR2X1 U18944 ( .IN1(n18015), .IN2(n18016), .Q(g26893) );
  AND2X1 U18945 ( .IN1(n18017), .IN2(n10784), .Q(n18016) );
  OR2X1 U18946 ( .IN1(n18018), .IN2(n18019), .Q(n18017) );
  AND2X1 U18947 ( .IN1(test_so17), .IN2(n18020), .Q(n18019) );
  AND2X1 U18948 ( .IN1(g29211), .IN2(n10578), .Q(n18018) );
  AND2X1 U18949 ( .IN1(n10904), .IN2(g355), .Q(n18015) );
  OR2X1 U18950 ( .IN1(n18021), .IN2(n18022), .Q(g26892) );
  AND2X1 U18951 ( .IN1(test_so17), .IN2(n10896), .Q(n18022) );
  AND2X1 U18952 ( .IN1(n18023), .IN2(n10578), .Q(n18021) );
  AND2X1 U18953 ( .IN1(n10820), .IN2(n18020), .Q(n18023) );
  OR2X1 U18954 ( .IN1(g333), .IN2(g355), .Q(n18020) );
  OR2X1 U18955 ( .IN1(n18024), .IN2(n18025), .Q(g26891) );
  AND2X1 U18956 ( .IN1(n18026), .IN2(n5860), .Q(n18025) );
  AND2X1 U18957 ( .IN1(n10820), .IN2(g7540), .Q(n18026) );
  INVX0 U18958 ( .INP(n18027), .ZN(n18024) );
  OR2X1 U18959 ( .IN1(n10738), .IN2(n5860), .Q(n18027) );
  OR2X1 U18960 ( .IN1(n18028), .IN2(n18029), .Q(g26890) );
  AND2X1 U18961 ( .IN1(n10904), .IN2(g333), .Q(n18029) );
  AND2X1 U18962 ( .IN1(n5860), .IN2(n10784), .Q(n18028) );
  OR2X1 U18963 ( .IN1(n18030), .IN2(n18031), .Q(g26889) );
  AND2X1 U18964 ( .IN1(n18032), .IN2(n10784), .Q(n18031) );
  AND2X1 U18965 ( .IN1(n18033), .IN2(n18034), .Q(n18032) );
  AND2X1 U18966 ( .IN1(g329), .IN2(DFF_709_n1), .Q(n18033) );
  AND2X1 U18967 ( .IN1(n10904), .IN2(g29211), .Q(n18030) );
  OR2X1 U18968 ( .IN1(n18035), .IN2(n18036), .Q(g26888) );
  AND2X1 U18969 ( .IN1(n10904), .IN2(g29216), .Q(n18036) );
  AND2X1 U18970 ( .IN1(n10821), .IN2(g316), .Q(n18035) );
  OR2X1 U18971 ( .IN1(n18037), .IN2(n18038), .Q(g26887) );
  OR2X1 U18972 ( .IN1(n18039), .IN2(n18040), .Q(n18038) );
  AND2X1 U18973 ( .IN1(n18041), .IN2(n10784), .Q(n18040) );
  AND2X1 U18974 ( .IN1(n5317), .IN2(g324), .Q(n18041) );
  AND2X1 U18975 ( .IN1(n10904), .IN2(g336), .Q(n18039) );
  OR2X1 U18976 ( .IN1(n18042), .IN2(n18043), .Q(g26886) );
  OR2X1 U18977 ( .IN1(n18044), .IN2(n18045), .Q(n18043) );
  AND2X1 U18978 ( .IN1(n10905), .IN2(g311), .Q(n18045) );
  AND2X1 U18979 ( .IN1(n18046), .IN2(n10784), .Q(n18044) );
  AND2X1 U18980 ( .IN1(n18034), .IN2(g336), .Q(n18046) );
  AND2X1 U18981 ( .IN1(n18037), .IN2(n18047), .Q(n18042) );
  OR2X1 U18982 ( .IN1(n18048), .IN2(n18049), .Q(g26884) );
  AND2X1 U18983 ( .IN1(n18050), .IN2(n10784), .Q(n18049) );
  OR2X1 U18984 ( .IN1(n18051), .IN2(n18052), .Q(n18050) );
  AND2X1 U18985 ( .IN1(n18047), .IN2(n18053), .Q(n18052) );
  OR2X1 U18986 ( .IN1(g26885), .IN2(n18054), .Q(n18053) );
  OR2X1 U18987 ( .IN1(n18055), .IN2(n18056), .Q(n18054) );
  AND2X1 U18988 ( .IN1(g305), .IN2(g336), .Q(n18056) );
  AND2X1 U18989 ( .IN1(n5824), .IN2(g311), .Q(n18055) );
  AND2X1 U18990 ( .IN1(n18057), .IN2(n18058), .Q(n18051) );
  AND2X1 U18991 ( .IN1(n5282), .IN2(n5317), .Q(n18058) );
  AND2X1 U18992 ( .IN1(n5766), .IN2(n5456), .Q(n18057) );
  AND2X1 U18993 ( .IN1(n10905), .IN2(g329), .Q(n18048) );
  OR2X1 U18994 ( .IN1(n18059), .IN2(n18060), .Q(g26883) );
  AND2X1 U18995 ( .IN1(n18047), .IN2(n10784), .Q(n18060) );
  INVX0 U18996 ( .INP(n18034), .ZN(n18047) );
  OR2X1 U18997 ( .IN1(n18061), .IN2(n18062), .Q(n18034) );
  AND2X1 U18998 ( .IN1(n5827), .IN2(n5317), .Q(n18062) );
  AND2X1 U18999 ( .IN1(n5282), .IN2(g324), .Q(n18061) );
  AND2X1 U19000 ( .IN1(n10905), .IN2(g324), .Q(n18059) );
  OR2X1 U19001 ( .IN1(n18037), .IN2(n18063), .Q(g26882) );
  OR2X1 U19002 ( .IN1(n18064), .IN2(n18065), .Q(n18063) );
  AND2X1 U19003 ( .IN1(n10905), .IN2(g316), .Q(n18065) );
  AND2X1 U19004 ( .IN1(n10821), .IN2(g311), .Q(n18064) );
  AND2X1 U19005 ( .IN1(g305), .IN2(n10784), .Q(n18037) );
  OR2X1 U19006 ( .IN1(n18066), .IN2(n18067), .Q(g26881) );
  AND2X1 U19007 ( .IN1(n10905), .IN2(g305), .Q(n18067) );
  AND2X1 U19008 ( .IN1(g6744), .IN2(n10785), .Q(n18066) );
  INVX0 U19009 ( .INP(n18068), .ZN(g26877) );
  AND2X1 U19010 ( .IN1(n11690), .IN2(n18069), .Q(n18068) );
  AND2X1 U19011 ( .IN1(n10821), .IN2(n11691), .Q(n18069) );
  OR2X1 U19012 ( .IN1(n18070), .IN2(n18071), .Q(n11691) );
  OR2X1 U19013 ( .IN1(n18072), .IN2(n18073), .Q(n18071) );
  OR2X1 U19014 ( .IN1(g2472), .IN2(g2204), .Q(n18073) );
  OR2X1 U19015 ( .IN1(g2491), .IN2(g2223), .Q(n18072) );
  OR2X1 U19016 ( .IN1(n18074), .IN2(n18075), .Q(n18070) );
  OR2X1 U19017 ( .IN1(g2338), .IN2(g2606), .Q(n18075) );
  OR2X1 U19018 ( .IN1(test_so40), .IN2(g2357), .Q(n18074) );
  OR2X1 U19019 ( .IN1(n18076), .IN2(n18077), .Q(n11690) );
  OR2X1 U19020 ( .IN1(n18078), .IN2(n18079), .Q(n18077) );
  OR2X1 U19021 ( .IN1(g2066), .IN2(g1798), .Q(n18079) );
  OR2X1 U19022 ( .IN1(g1779), .IN2(g2047), .Q(n18078) );
  OR2X1 U19023 ( .IN1(n18080), .IN2(n18081), .Q(n18076) );
  OR2X1 U19024 ( .IN1(g1913), .IN2(g1932), .Q(n18081) );
  OR2X1 U19025 ( .IN1(test_so75), .IN2(g1664), .Q(n18080) );
  INVX0 U19026 ( .INP(n18082), .ZN(g26876) );
  AND2X1 U19027 ( .IN1(n11713), .IN2(n18083), .Q(n18082) );
  AND2X1 U19028 ( .IN1(n10821), .IN2(n11714), .Q(n18083) );
  OR2X1 U19029 ( .IN1(n18084), .IN2(n18085), .Q(n11714) );
  OR2X1 U19030 ( .IN1(n18086), .IN2(n18087), .Q(n18085) );
  OR2X1 U19031 ( .IN1(n9273), .IN2(n9262), .Q(n18087) );
  OR2X1 U19032 ( .IN1(n9324), .IN2(n9295), .Q(n18086) );
  OR2X1 U19033 ( .IN1(n18088), .IN2(n18089), .Q(n18084) );
  OR2X1 U19034 ( .IN1(g2269), .IN2(g2537), .Q(n18089) );
  OR2X1 U19035 ( .IN1(test_so31), .IN2(g2671), .Q(n18088) );
  OR2X1 U19036 ( .IN1(n18090), .IN2(n18091), .Q(n11713) );
  OR2X1 U19037 ( .IN1(n18092), .IN2(n18093), .Q(n18091) );
  OR2X1 U19038 ( .IN1(g1858), .IN2(n9236), .Q(n18093) );
  OR2X1 U19039 ( .IN1(g1992), .IN2(g2126), .Q(n18092) );
  OR2X1 U19040 ( .IN1(n18094), .IN2(n18095), .Q(n18090) );
  OR2X1 U19041 ( .IN1(g1844), .IN2(g2112), .Q(n18095) );
  OR2X1 U19042 ( .IN1(g1710), .IN2(g1978), .Q(n18094) );
  INVX0 U19043 ( .INP(n18096), .ZN(g26875) );
  AND2X1 U19044 ( .IN1(n11718), .IN2(n18097), .Q(n18096) );
  AND2X1 U19045 ( .IN1(n10822), .IN2(n11719), .Q(n18097) );
  OR2X1 U19046 ( .IN1(n18098), .IN2(n18099), .Q(n11719) );
  OR2X1 U19047 ( .IN1(g2255), .IN2(g2389), .Q(n18099) );
  OR2X1 U19048 ( .IN1(g2523), .IN2(g2657), .Q(n18098) );
  OR2X1 U19049 ( .IN1(n18100), .IN2(n18101), .Q(n11718) );
  OR2X1 U19050 ( .IN1(g1830), .IN2(g1696), .Q(n18101) );
  OR2X1 U19051 ( .IN1(g2098), .IN2(g1964), .Q(n18100) );
  OR2X1 U19052 ( .IN1(n18102), .IN2(n18103), .Q(g25764) );
  AND2X1 U19053 ( .IN1(n18104), .IN2(g6541), .Q(n18103) );
  AND2X1 U19054 ( .IN1(n14635), .IN2(g6505), .Q(n18102) );
  OR2X1 U19055 ( .IN1(n18105), .IN2(n18106), .Q(g25763) );
  OR2X1 U19056 ( .IN1(n18107), .IN2(n18108), .Q(n18106) );
  AND2X1 U19057 ( .IN1(n18109), .IN2(n5445), .Q(n18108) );
  AND2X1 U19058 ( .IN1(n18110), .IN2(n5659), .Q(n18109) );
  AND2X1 U19059 ( .IN1(n13075), .IN2(n10785), .Q(n18110) );
  AND2X1 U19060 ( .IN1(n18111), .IN2(g6533), .Q(n18107) );
  OR2X1 U19061 ( .IN1(n10882), .IN2(n18112), .Q(n18111) );
  AND2X1 U19062 ( .IN1(n13075), .IN2(g6527), .Q(n18112) );
  INVX0 U19063 ( .INP(n18113), .ZN(n18105) );
  OR2X1 U19064 ( .IN1(n18104), .IN2(n5884), .Q(n18113) );
  OR2X1 U19065 ( .IN1(n18114), .IN2(n18115), .Q(g25762) );
  AND2X1 U19066 ( .IN1(n18104), .IN2(g6527), .Q(n18115) );
  AND2X1 U19067 ( .IN1(n14635), .IN2(g6533), .Q(n18114) );
  OR2X1 U19068 ( .IN1(n18116), .IN2(n18117), .Q(g25761) );
  OR2X1 U19069 ( .IN1(n18118), .IN2(n18119), .Q(n18117) );
  INVX0 U19070 ( .INP(n18120), .ZN(n18119) );
  OR2X1 U19071 ( .IN1(n10737), .IN2(n10484), .Q(n18120) );
  AND2X1 U19072 ( .IN1(n18121), .IN2(n10785), .Q(n18118) );
  AND2X1 U19073 ( .IN1(n5426), .IN2(n13075), .Q(n18121) );
  AND2X1 U19074 ( .IN1(n14635), .IN2(g6513), .Q(n18116) );
  INVX0 U19075 ( .INP(n18104), .ZN(n14635) );
  OR2X1 U19076 ( .IN1(n10882), .IN2(n13075), .Q(n18104) );
  AND2X1 U19077 ( .IN1(g6561), .IN2(n14664), .Q(n13075) );
  AND2X1 U19078 ( .IN1(g6565), .IN2(g6573), .Q(n14664) );
  OR2X1 U19079 ( .IN1(n18122), .IN2(n18123), .Q(g25758) );
  AND2X1 U19080 ( .IN1(n18124), .IN2(n10785), .Q(n18123) );
  AND2X1 U19081 ( .IN1(n10048), .IN2(n18125), .Q(n18124) );
  OR2X1 U19082 ( .IN1(n18126), .IN2(g6444), .Q(n18125) );
  AND2X1 U19083 ( .IN1(n10049), .IN2(g9743), .Q(n18126) );
  INVX0 U19084 ( .INP(n18127), .ZN(n18122) );
  OR2X1 U19085 ( .IN1(n10737), .IN2(n10049), .Q(n18127) );
  OR2X1 U19086 ( .IN1(n18128), .IN2(n18129), .Q(g25757) );
  AND2X1 U19087 ( .IN1(n10905), .IN2(g6444), .Q(n18129) );
  AND2X1 U19088 ( .IN1(n10822), .IN2(g6727), .Q(n18128) );
  AND2X1 U19089 ( .IN1(g6573), .IN2(n10785), .Q(g25756) );
  OR2X1 U19090 ( .IN1(n18130), .IN2(n18131), .Q(g25750) );
  AND2X1 U19091 ( .IN1(n18132), .IN2(g6195), .Q(n18131) );
  AND2X1 U19092 ( .IN1(n14762), .IN2(g6159), .Q(n18130) );
  OR2X1 U19093 ( .IN1(n18133), .IN2(n18134), .Q(g25749) );
  OR2X1 U19094 ( .IN1(n18135), .IN2(n18136), .Q(n18134) );
  AND2X1 U19095 ( .IN1(n18137), .IN2(n5453), .Q(n18136) );
  AND2X1 U19096 ( .IN1(n18138), .IN2(n5667), .Q(n18137) );
  AND2X1 U19097 ( .IN1(n13092), .IN2(n10785), .Q(n18138) );
  AND2X1 U19098 ( .IN1(n18139), .IN2(g6187), .Q(n18135) );
  OR2X1 U19099 ( .IN1(n10882), .IN2(n18140), .Q(n18139) );
  AND2X1 U19100 ( .IN1(n13092), .IN2(g6181), .Q(n18140) );
  INVX0 U19101 ( .INP(n18141), .ZN(n18133) );
  OR2X1 U19102 ( .IN1(n18132), .IN2(n5888), .Q(n18141) );
  OR2X1 U19103 ( .IN1(n18142), .IN2(n18143), .Q(g25748) );
  AND2X1 U19104 ( .IN1(n18132), .IN2(g6181), .Q(n18143) );
  AND2X1 U19105 ( .IN1(n14762), .IN2(g6187), .Q(n18142) );
  OR2X1 U19106 ( .IN1(n18144), .IN2(n18145), .Q(g25747) );
  OR2X1 U19107 ( .IN1(n18146), .IN2(n18147), .Q(n18145) );
  AND2X1 U19108 ( .IN1(n10905), .IN2(g6163), .Q(n18147) );
  AND2X1 U19109 ( .IN1(n18148), .IN2(n10785), .Q(n18146) );
  AND2X1 U19110 ( .IN1(n5430), .IN2(n13092), .Q(n18148) );
  AND2X1 U19111 ( .IN1(n14762), .IN2(g6167), .Q(n18144) );
  INVX0 U19112 ( .INP(n18132), .ZN(n14762) );
  OR2X1 U19113 ( .IN1(n10882), .IN2(n13092), .Q(n18132) );
  AND2X1 U19114 ( .IN1(g6215), .IN2(n14791), .Q(n13092) );
  AND2X1 U19115 ( .IN1(g6219), .IN2(g6227), .Q(n14791) );
  OR2X1 U19116 ( .IN1(n18149), .IN2(n18150), .Q(g25744) );
  AND2X1 U19117 ( .IN1(n18151), .IN2(n10785), .Q(n18150) );
  AND2X1 U19118 ( .IN1(n10045), .IN2(n18152), .Q(n18151) );
  OR2X1 U19119 ( .IN1(n18153), .IN2(g6098), .Q(n18152) );
  AND2X1 U19120 ( .IN1(test_so92), .IN2(n10046), .Q(n18153) );
  INVX0 U19121 ( .INP(n18154), .ZN(n18149) );
  OR2X1 U19122 ( .IN1(n10737), .IN2(n10046), .Q(n18154) );
  OR2X1 U19123 ( .IN1(n18155), .IN2(n18156), .Q(g25743) );
  AND2X1 U19124 ( .IN1(n10905), .IN2(g6098), .Q(n18156) );
  AND2X1 U19125 ( .IN1(test_so69), .IN2(n10785), .Q(n18155) );
  AND2X1 U19126 ( .IN1(g6227), .IN2(n10786), .Q(g25742) );
  OR2X1 U19127 ( .IN1(n18157), .IN2(n18158), .Q(g25736) );
  AND2X1 U19128 ( .IN1(n18159), .IN2(g5849), .Q(n18158) );
  AND2X1 U19129 ( .IN1(n14889), .IN2(g5813), .Q(n18157) );
  OR2X1 U19130 ( .IN1(n18160), .IN2(n18161), .Q(g25735) );
  OR2X1 U19131 ( .IN1(n18162), .IN2(n18163), .Q(n18161) );
  AND2X1 U19132 ( .IN1(n18164), .IN2(n5449), .Q(n18163) );
  AND2X1 U19133 ( .IN1(n18165), .IN2(n5663), .Q(n18164) );
  AND2X1 U19134 ( .IN1(n13091), .IN2(n10786), .Q(n18165) );
  AND2X1 U19135 ( .IN1(n18166), .IN2(g5841), .Q(n18162) );
  OR2X1 U19136 ( .IN1(n10882), .IN2(n18167), .Q(n18166) );
  AND2X1 U19137 ( .IN1(n13091), .IN2(g5835), .Q(n18167) );
  AND2X1 U19138 ( .IN1(test_so83), .IN2(n14889), .Q(n18160) );
  OR2X1 U19139 ( .IN1(n18168), .IN2(n18169), .Q(g25734) );
  AND2X1 U19140 ( .IN1(n18159), .IN2(g5835), .Q(n18169) );
  AND2X1 U19141 ( .IN1(n14889), .IN2(g5841), .Q(n18168) );
  OR2X1 U19142 ( .IN1(n18170), .IN2(n18171), .Q(g25733) );
  OR2X1 U19143 ( .IN1(n18172), .IN2(n18173), .Q(n18171) );
  AND2X1 U19144 ( .IN1(n10905), .IN2(g5817), .Q(n18173) );
  AND2X1 U19145 ( .IN1(n18174), .IN2(n10786), .Q(n18172) );
  AND2X1 U19146 ( .IN1(n5429), .IN2(n13091), .Q(n18174) );
  AND2X1 U19147 ( .IN1(n14889), .IN2(g5821), .Q(n18170) );
  INVX0 U19148 ( .INP(n18159), .ZN(n14889) );
  OR2X1 U19149 ( .IN1(n10881), .IN2(n13091), .Q(n18159) );
  AND2X1 U19150 ( .IN1(g5869), .IN2(n14918), .Q(n13091) );
  AND2X1 U19151 ( .IN1(g5873), .IN2(test_so36), .Q(n14918) );
  OR2X1 U19152 ( .IN1(n18175), .IN2(n18176), .Q(g25730) );
  AND2X1 U19153 ( .IN1(n18177), .IN2(n10786), .Q(n18176) );
  AND2X1 U19154 ( .IN1(n10057), .IN2(n18178), .Q(n18177) );
  OR2X1 U19155 ( .IN1(n18179), .IN2(g5752), .Q(n18178) );
  AND2X1 U19156 ( .IN1(n10058), .IN2(g9617), .Q(n18179) );
  INVX0 U19157 ( .INP(n18180), .ZN(n18175) );
  OR2X1 U19158 ( .IN1(n10740), .IN2(n10058), .Q(n18180) );
  OR2X1 U19159 ( .IN1(n18181), .IN2(n18182), .Q(g25729) );
  AND2X1 U19160 ( .IN1(n10905), .IN2(g5752), .Q(n18182) );
  AND2X1 U19161 ( .IN1(n10822), .IN2(g6035), .Q(n18181) );
  AND2X1 U19162 ( .IN1(n10823), .IN2(test_so36), .Q(g25728) );
  OR2X1 U19163 ( .IN1(n18183), .IN2(n18184), .Q(g25722) );
  AND2X1 U19164 ( .IN1(n18185), .IN2(g5503), .Q(n18184) );
  AND2X1 U19165 ( .IN1(n15015), .IN2(g5467), .Q(n18183) );
  OR2X1 U19166 ( .IN1(n18186), .IN2(n18187), .Q(g25721) );
  OR2X1 U19167 ( .IN1(n18188), .IN2(n18189), .Q(n18187) );
  AND2X1 U19168 ( .IN1(n18190), .IN2(n5446), .Q(n18189) );
  AND2X1 U19169 ( .IN1(n18191), .IN2(n5660), .Q(n18190) );
  AND2X1 U19170 ( .IN1(n13093), .IN2(n10786), .Q(n18191) );
  AND2X1 U19171 ( .IN1(n18192), .IN2(g5495), .Q(n18188) );
  OR2X1 U19172 ( .IN1(n10881), .IN2(n18193), .Q(n18192) );
  AND2X1 U19173 ( .IN1(n13093), .IN2(g5489), .Q(n18193) );
  INVX0 U19174 ( .INP(n18194), .ZN(n18186) );
  OR2X1 U19175 ( .IN1(n18185), .IN2(n5885), .Q(n18194) );
  OR2X1 U19176 ( .IN1(n18195), .IN2(n18196), .Q(g25720) );
  AND2X1 U19177 ( .IN1(n18185), .IN2(g5489), .Q(n18196) );
  AND2X1 U19178 ( .IN1(n15015), .IN2(g5495), .Q(n18195) );
  OR2X1 U19179 ( .IN1(n18197), .IN2(n18198), .Q(g25719) );
  OR2X1 U19180 ( .IN1(n18199), .IN2(n18200), .Q(n18198) );
  AND2X1 U19181 ( .IN1(n10906), .IN2(g5471), .Q(n18200) );
  AND2X1 U19182 ( .IN1(n18201), .IN2(n10786), .Q(n18199) );
  AND2X1 U19183 ( .IN1(n5425), .IN2(n13093), .Q(n18201) );
  AND2X1 U19184 ( .IN1(n15015), .IN2(g5475), .Q(n18197) );
  INVX0 U19185 ( .INP(n18185), .ZN(n15015) );
  OR2X1 U19186 ( .IN1(n10881), .IN2(n13093), .Q(n18185) );
  AND2X1 U19187 ( .IN1(g5523), .IN2(n15044), .Q(n13093) );
  AND2X1 U19188 ( .IN1(g5527), .IN2(g5535), .Q(n15044) );
  OR2X1 U19189 ( .IN1(n18202), .IN2(n18203), .Q(g25716) );
  AND2X1 U19190 ( .IN1(n18204), .IN2(n10786), .Q(n18203) );
  AND2X1 U19191 ( .IN1(n18205), .IN2(n10051), .Q(n18204) );
  OR2X1 U19192 ( .IN1(n18206), .IN2(g5406), .Q(n18205) );
  AND2X1 U19193 ( .IN1(n10052), .IN2(g9555), .Q(n18206) );
  INVX0 U19194 ( .INP(n18207), .ZN(n18202) );
  OR2X1 U19195 ( .IN1(n10737), .IN2(n10052), .Q(n18207) );
  OR2X1 U19196 ( .IN1(n18208), .IN2(n18209), .Q(g25715) );
  AND2X1 U19197 ( .IN1(n10906), .IN2(g5406), .Q(n18209) );
  AND2X1 U19198 ( .IN1(n10823), .IN2(g5689), .Q(n18208) );
  AND2X1 U19199 ( .IN1(g5535), .IN2(n10786), .Q(g25714) );
  OR2X1 U19200 ( .IN1(n18210), .IN2(n18211), .Q(g25708) );
  AND2X1 U19201 ( .IN1(n18212), .IN2(g5156), .Q(n18211) );
  AND2X1 U19202 ( .IN1(n15141), .IN2(g5120), .Q(n18210) );
  OR2X1 U19203 ( .IN1(n18213), .IN2(n18214), .Q(g25707) );
  OR2X1 U19204 ( .IN1(n18215), .IN2(n18216), .Q(n18214) );
  AND2X1 U19205 ( .IN1(n18217), .IN2(n10591), .Q(n18216) );
  AND2X1 U19206 ( .IN1(n18218), .IN2(n5658), .Q(n18217) );
  AND2X1 U19207 ( .IN1(g32975), .IN2(n10786), .Q(n18218) );
  AND2X1 U19208 ( .IN1(test_so98), .IN2(n18219), .Q(n18215) );
  OR2X1 U19209 ( .IN1(n10881), .IN2(n18220), .Q(n18219) );
  AND2X1 U19210 ( .IN1(g32975), .IN2(g5142), .Q(n18220) );
  INVX0 U19211 ( .INP(n18221), .ZN(n18213) );
  OR2X1 U19212 ( .IN1(n18212), .IN2(n5883), .Q(n18221) );
  OR2X1 U19213 ( .IN1(n18222), .IN2(n18223), .Q(g25706) );
  AND2X1 U19214 ( .IN1(n18212), .IN2(g5142), .Q(n18223) );
  AND2X1 U19215 ( .IN1(test_so98), .IN2(n15141), .Q(n18222) );
  OR2X1 U19216 ( .IN1(n18224), .IN2(n18225), .Q(g25705) );
  OR2X1 U19217 ( .IN1(n18226), .IN2(n18227), .Q(n18225) );
  AND2X1 U19218 ( .IN1(n10906), .IN2(g5124), .Q(n18227) );
  AND2X1 U19219 ( .IN1(n18228), .IN2(n10787), .Q(n18226) );
  AND2X1 U19220 ( .IN1(g32975), .IN2(n10577), .Q(n18228) );
  AND2X1 U19221 ( .IN1(test_so96), .IN2(n15141), .Q(n18224) );
  INVX0 U19222 ( .INP(n18212), .ZN(n15141) );
  OR2X1 U19223 ( .IN1(n10881), .IN2(g32975), .Q(n18212) );
  AND2X1 U19224 ( .IN1(g5176), .IN2(n15170), .Q(g32975) );
  AND2X1 U19225 ( .IN1(g5180), .IN2(g5188), .Q(n15170) );
  AND2X1 U19226 ( .IN1(n18229), .IN2(g5073), .Q(g25704) );
  OR2X1 U19227 ( .IN1(n10880), .IN2(g5069), .Q(n18229) );
  OR2X1 U19228 ( .IN1(n18230), .IN2(n18231), .Q(g25703) );
  AND2X1 U19229 ( .IN1(n18232), .IN2(n10787), .Q(n18231) );
  AND2X1 U19230 ( .IN1(n5689), .IN2(n18233), .Q(n18232) );
  OR2X1 U19231 ( .IN1(n18234), .IN2(g5022), .Q(n18233) );
  AND2X1 U19232 ( .IN1(n10489), .IN2(g9553), .Q(n18234) );
  AND2X1 U19233 ( .IN1(n10906), .IN2(g5112), .Q(n18230) );
  OR2X1 U19234 ( .IN1(n18235), .IN2(n18236), .Q(g25702) );
  AND2X1 U19235 ( .IN1(n18237), .IN2(n10787), .Q(n18236) );
  AND2X1 U19236 ( .IN1(n5690), .IN2(n18238), .Q(n18237) );
  INVX0 U19237 ( .INP(n18239), .ZN(n18238) );
  AND2X1 U19238 ( .IN1(n18240), .IN2(n10508), .Q(n18239) );
  OR2X1 U19239 ( .IN1(n5689), .IN2(test_so32), .Q(n18240) );
  AND2X1 U19240 ( .IN1(test_so32), .IN2(n10895), .Q(n18235) );
  OR2X1 U19241 ( .IN1(n18241), .IN2(n18242), .Q(g25701) );
  AND2X1 U19242 ( .IN1(n10906), .IN2(g5062), .Q(n18242) );
  AND2X1 U19243 ( .IN1(test_so10), .IN2(n10787), .Q(n18241) );
  AND2X1 U19244 ( .IN1(g5188), .IN2(n10787), .Q(g25700) );
  OR2X1 U19245 ( .IN1(n18243), .IN2(n18244), .Q(g25699) );
  OR2X1 U19246 ( .IN1(n18245), .IN2(n18246), .Q(n18244) );
  AND2X1 U19247 ( .IN1(n5014), .IN2(n5669), .Q(n18246) );
  INVX0 U19248 ( .INP(n18247), .ZN(n18245) );
  OR2X1 U19249 ( .IN1(n18248), .IN2(n5669), .Q(n18247) );
  OR2X1 U19250 ( .IN1(n10880), .IN2(n5014), .Q(n18248) );
  AND2X1 U19251 ( .IN1(n10906), .IN2(g5097), .Q(n18243) );
  OR2X1 U19252 ( .IN1(n18249), .IN2(n18250), .Q(g25698) );
  OR2X1 U19253 ( .IN1(n18251), .IN2(n18252), .Q(n18250) );
  AND2X1 U19254 ( .IN1(n5016), .IN2(n5753), .Q(n18252) );
  INVX0 U19255 ( .INP(n18253), .ZN(n18251) );
  OR2X1 U19256 ( .IN1(n18254), .IN2(n5753), .Q(n18253) );
  OR2X1 U19257 ( .IN1(n10880), .IN2(n5016), .Q(n18254) );
  AND2X1 U19258 ( .IN1(n10906), .IN2(g5092), .Q(n18249) );
  XOR2X1 U19259 ( .IN1(g5084), .IN2(n18255), .Q(g25697) );
  AND2X1 U19260 ( .IN1(n10824), .IN2(g5092), .Q(n18255) );
  OR2X1 U19261 ( .IN1(n18256), .IN2(n18257), .Q(g25696) );
  OR2X1 U19262 ( .IN1(n18258), .IN2(n18259), .Q(n18257) );
  AND2X1 U19263 ( .IN1(n18260), .IN2(n5893), .Q(n18259) );
  AND2X1 U19264 ( .IN1(n18261), .IN2(n18262), .Q(n18260) );
  OR2X1 U19265 ( .IN1(n5455), .IN2(g5069), .Q(n18262) );
  INVX0 U19266 ( .INP(n18263), .ZN(n18258) );
  OR2X1 U19267 ( .IN1(n18261), .IN2(n5893), .Q(n18263) );
  AND2X1 U19268 ( .IN1(n10824), .IN2(n5681), .Q(n18261) );
  AND2X1 U19269 ( .IN1(n18264), .IN2(n10481), .Q(n18256) );
  AND2X1 U19270 ( .IN1(n10824), .IN2(g5077), .Q(n18264) );
  AND2X1 U19271 ( .IN1(n18265), .IN2(g5077), .Q(g25695) );
  OR2X1 U19272 ( .IN1(n10879), .IN2(n18266), .Q(n18265) );
  OR2X1 U19273 ( .IN1(n18267), .IN2(n18268), .Q(n18266) );
  AND2X1 U19274 ( .IN1(n10481), .IN2(n5681), .Q(n18268) );
  AND2X1 U19275 ( .IN1(n10091), .IN2(g5084), .Q(n18267) );
  OR2X1 U19276 ( .IN1(n18269), .IN2(n18270), .Q(g25691) );
  INVX0 U19277 ( .INP(n18271), .ZN(n18270) );
  OR2X1 U19278 ( .IN1(n10737), .IN2(n10497), .Q(n18271) );
  AND2X1 U19279 ( .IN1(n10542), .IN2(n18272), .Q(n18269) );
  OR2X1 U19280 ( .IN1(n18273), .IN2(n18274), .Q(n18272) );
  OR2X1 U19281 ( .IN1(g4057), .IN2(n18275), .Q(n18274) );
  OR2X1 U19282 ( .IN1(n15136), .IN2(g4064), .Q(n18275) );
  OR2X1 U19283 ( .IN1(n5480), .IN2(g4093), .Q(n15136) );
  OR2X1 U19284 ( .IN1(n18276), .IN2(n18277), .Q(n18273) );
  OR2X1 U19285 ( .IN1(g4141), .IN2(n10554), .Q(n18277) );
  OR2X1 U19286 ( .IN1(n5350), .IN2(g4082), .Q(n18276) );
  OR2X1 U19287 ( .IN1(n18278), .IN2(n18279), .Q(g25690) );
  AND2X1 U19288 ( .IN1(n18280), .IN2(n10787), .Q(n18279) );
  AND2X1 U19289 ( .IN1(n10497), .IN2(g25689), .Q(n18280) );
  AND2X1 U19290 ( .IN1(n10906), .IN2(g4169), .Q(n18278) );
  OR2X1 U19291 ( .IN1(n18281), .IN2(n18282), .Q(g25687) );
  OR2X1 U19292 ( .IN1(n18283), .IN2(n18284), .Q(n18282) );
  AND2X1 U19293 ( .IN1(n5026), .IN2(n15280), .Q(n18284) );
  AND2X1 U19294 ( .IN1(n18285), .IN2(n5612), .Q(n18283) );
  AND2X1 U19295 ( .IN1(n17774), .IN2(g4169), .Q(n18285) );
  AND2X1 U19296 ( .IN1(g4064), .IN2(g4057), .Q(n17774) );
  AND2X1 U19297 ( .IN1(n10906), .IN2(g4057), .Q(n18281) );
  OR2X1 U19298 ( .IN1(n18286), .IN2(n18287), .Q(g25686) );
  AND2X1 U19299 ( .IN1(n18288), .IN2(n5416), .Q(n18287) );
  AND2X1 U19300 ( .IN1(n15280), .IN2(g4057), .Q(n18288) );
  AND2X1 U19301 ( .IN1(g4169), .IN2(n10787), .Q(n15280) );
  AND2X1 U19302 ( .IN1(n18289), .IN2(g4064), .Q(n18286) );
  OR2X1 U19303 ( .IN1(n10879), .IN2(n18290), .Q(n18289) );
  AND2X1 U19304 ( .IN1(n5711), .IN2(g4169), .Q(n18290) );
  OR2X1 U19305 ( .IN1(n10542), .IN2(n18291), .Q(g25685) );
  OR2X1 U19306 ( .IN1(n18292), .IN2(n18293), .Q(n18291) );
  AND2X1 U19307 ( .IN1(n10906), .IN2(g4072), .Q(n18293) );
  AND2X1 U19308 ( .IN1(n5416), .IN2(n10787), .Q(n18292) );
  AND2X1 U19309 ( .IN1(n10824), .IN2(n5729), .Q(n10542) );
  OR2X1 U19310 ( .IN1(n18294), .IN2(n18295), .Q(g25684) );
  AND2X1 U19311 ( .IN1(n18296), .IN2(g3849), .Q(n18295) );
  AND2X1 U19312 ( .IN1(n15287), .IN2(g3813), .Q(n18294) );
  OR2X1 U19313 ( .IN1(n18297), .IN2(n18298), .Q(g25683) );
  OR2X1 U19314 ( .IN1(n18299), .IN2(n18300), .Q(n18298) );
  AND2X1 U19315 ( .IN1(n18301), .IN2(n10592), .Q(n18300) );
  AND2X1 U19316 ( .IN1(n18302), .IN2(n5662), .Q(n18301) );
  AND2X1 U19317 ( .IN1(n13080), .IN2(n10787), .Q(n18302) );
  AND2X1 U19318 ( .IN1(test_so97), .IN2(n18303), .Q(n18299) );
  OR2X1 U19319 ( .IN1(n10879), .IN2(n18304), .Q(n18303) );
  AND2X1 U19320 ( .IN1(n13080), .IN2(g3835), .Q(n18304) );
  INVX0 U19321 ( .INP(n18305), .ZN(n18297) );
  OR2X1 U19322 ( .IN1(n18296), .IN2(n5886), .Q(n18305) );
  OR2X1 U19323 ( .IN1(n18306), .IN2(n18307), .Q(g25682) );
  AND2X1 U19324 ( .IN1(n18296), .IN2(g3835), .Q(n18307) );
  AND2X1 U19325 ( .IN1(test_so97), .IN2(n15287), .Q(n18306) );
  OR2X1 U19326 ( .IN1(n18308), .IN2(n18309), .Q(g25681) );
  OR2X1 U19327 ( .IN1(n18310), .IN2(n18311), .Q(n18309) );
  AND2X1 U19328 ( .IN1(n10906), .IN2(g3817), .Q(n18311) );
  AND2X1 U19329 ( .IN1(n18312), .IN2(n10788), .Q(n18310) );
  AND2X1 U19330 ( .IN1(n5428), .IN2(n13080), .Q(n18312) );
  AND2X1 U19331 ( .IN1(n15287), .IN2(g3821), .Q(n18308) );
  INVX0 U19332 ( .INP(n18296), .ZN(n15287) );
  OR2X1 U19333 ( .IN1(n10878), .IN2(n13080), .Q(n18296) );
  AND2X1 U19334 ( .IN1(n15316), .IN2(test_so33), .Q(n13080) );
  AND2X1 U19335 ( .IN1(g3873), .IN2(g3881), .Q(n15316) );
  OR2X1 U19336 ( .IN1(n18313), .IN2(n18314), .Q(g25678) );
  AND2X1 U19337 ( .IN1(n18315), .IN2(n10788), .Q(n18314) );
  AND2X1 U19338 ( .IN1(n10053), .IN2(n18316), .Q(n18315) );
  OR2X1 U19339 ( .IN1(n18317), .IN2(g3752), .Q(n18316) );
  AND2X1 U19340 ( .IN1(n10054), .IN2(g8344), .Q(n18317) );
  INVX0 U19341 ( .INP(n18318), .ZN(n18313) );
  OR2X1 U19342 ( .IN1(n10738), .IN2(n10054), .Q(n18318) );
  OR2X1 U19343 ( .IN1(n18319), .IN2(n18320), .Q(g25677) );
  AND2X1 U19344 ( .IN1(n10906), .IN2(g3752), .Q(n18320) );
  AND2X1 U19345 ( .IN1(n10825), .IN2(g4040), .Q(n18319) );
  AND2X1 U19346 ( .IN1(g3881), .IN2(n10788), .Q(g25676) );
  OR2X1 U19347 ( .IN1(n18321), .IN2(n18322), .Q(g25670) );
  AND2X1 U19348 ( .IN1(n18323), .IN2(g3498), .Q(n18322) );
  AND2X1 U19349 ( .IN1(n15412), .IN2(g3462), .Q(n18321) );
  OR2X1 U19350 ( .IN1(n18324), .IN2(n18325), .Q(g25669) );
  OR2X1 U19351 ( .IN1(n18326), .IN2(n18327), .Q(n18325) );
  AND2X1 U19352 ( .IN1(n18328), .IN2(n5454), .Q(n18327) );
  AND2X1 U19353 ( .IN1(n18329), .IN2(n5668), .Q(n18328) );
  AND2X1 U19354 ( .IN1(n13079), .IN2(n10788), .Q(n18329) );
  AND2X1 U19355 ( .IN1(n18330), .IN2(g3490), .Q(n18326) );
  OR2X1 U19356 ( .IN1(n10879), .IN2(n18331), .Q(n18330) );
  AND2X1 U19357 ( .IN1(n13079), .IN2(g3484), .Q(n18331) );
  INVX0 U19358 ( .INP(n18332), .ZN(n18324) );
  OR2X1 U19359 ( .IN1(n18323), .IN2(n5889), .Q(n18332) );
  OR2X1 U19360 ( .IN1(n18333), .IN2(n18334), .Q(g25668) );
  AND2X1 U19361 ( .IN1(n18323), .IN2(g3484), .Q(n18334) );
  AND2X1 U19362 ( .IN1(n15412), .IN2(g3490), .Q(n18333) );
  OR2X1 U19363 ( .IN1(n18335), .IN2(n18336), .Q(g25667) );
  OR2X1 U19364 ( .IN1(n18337), .IN2(n18338), .Q(n18336) );
  AND2X1 U19365 ( .IN1(n10907), .IN2(g3466), .Q(n18338) );
  AND2X1 U19366 ( .IN1(n18339), .IN2(n10788), .Q(n18337) );
  AND2X1 U19367 ( .IN1(n5424), .IN2(n13079), .Q(n18339) );
  AND2X1 U19368 ( .IN1(n15412), .IN2(g3470), .Q(n18335) );
  INVX0 U19369 ( .INP(n18323), .ZN(n15412) );
  OR2X1 U19370 ( .IN1(n10878), .IN2(n13079), .Q(n18323) );
  AND2X1 U19371 ( .IN1(g3518), .IN2(n15441), .Q(n13079) );
  AND2X1 U19372 ( .IN1(g3522), .IN2(g3530), .Q(n15441) );
  OR2X1 U19373 ( .IN1(n18340), .IN2(n18341), .Q(g25664) );
  AND2X1 U19374 ( .IN1(n18342), .IN2(n10788), .Q(n18341) );
  AND2X1 U19375 ( .IN1(n10036), .IN2(n18343), .Q(n18342) );
  OR2X1 U19376 ( .IN1(n18344), .IN2(g3401), .Q(n18343) );
  AND2X1 U19377 ( .IN1(n10037), .IN2(g8279), .Q(n18344) );
  INVX0 U19378 ( .INP(n18345), .ZN(n18340) );
  OR2X1 U19379 ( .IN1(n10738), .IN2(n10037), .Q(n18345) );
  OR2X1 U19380 ( .IN1(n18346), .IN2(n18347), .Q(g25663) );
  AND2X1 U19381 ( .IN1(n10907), .IN2(g3401), .Q(n18347) );
  AND2X1 U19382 ( .IN1(n10825), .IN2(g3689), .Q(n18346) );
  AND2X1 U19383 ( .IN1(g3530), .IN2(n10788), .Q(g25662) );
  OR2X1 U19384 ( .IN1(n18348), .IN2(n18349), .Q(g25656) );
  AND2X1 U19385 ( .IN1(n18350), .IN2(g3147), .Q(n18349) );
  AND2X1 U19386 ( .IN1(n15537), .IN2(g3111), .Q(n18348) );
  OR2X1 U19387 ( .IN1(n18351), .IN2(n18352), .Q(g25655) );
  OR2X1 U19388 ( .IN1(n18353), .IN2(n18354), .Q(n18352) );
  AND2X1 U19389 ( .IN1(n18355), .IN2(n5447), .Q(n18354) );
  AND2X1 U19390 ( .IN1(n18356), .IN2(n5661), .Q(n18355) );
  AND2X1 U19391 ( .IN1(n13082), .IN2(n10788), .Q(n18356) );
  AND2X1 U19392 ( .IN1(n18357), .IN2(g3139), .Q(n18353) );
  OR2X1 U19393 ( .IN1(n10878), .IN2(n18358), .Q(n18357) );
  AND2X1 U19394 ( .IN1(n13082), .IN2(g3133), .Q(n18358) );
  AND2X1 U19395 ( .IN1(n15537), .IN2(g3143), .Q(n18351) );
  OR2X1 U19396 ( .IN1(n18359), .IN2(n18360), .Q(g25654) );
  AND2X1 U19397 ( .IN1(n18350), .IN2(g3133), .Q(n18360) );
  AND2X1 U19398 ( .IN1(n15537), .IN2(g3139), .Q(n18359) );
  OR2X1 U19399 ( .IN1(n18361), .IN2(n18362), .Q(g25653) );
  OR2X1 U19400 ( .IN1(n18363), .IN2(n18364), .Q(n18362) );
  AND2X1 U19401 ( .IN1(n10907), .IN2(g3115), .Q(n18364) );
  AND2X1 U19402 ( .IN1(n18365), .IN2(n10789), .Q(n18363) );
  AND2X1 U19403 ( .IN1(n5423), .IN2(n13082), .Q(n18365) );
  AND2X1 U19404 ( .IN1(n15537), .IN2(g3119), .Q(n18361) );
  INVX0 U19405 ( .INP(n18350), .ZN(n15537) );
  OR2X1 U19406 ( .IN1(n10877), .IN2(n13082), .Q(n18350) );
  AND2X1 U19407 ( .IN1(g3167), .IN2(n15566), .Q(n13082) );
  AND2X1 U19408 ( .IN1(g3179), .IN2(g3171), .Q(n15566) );
  OR2X1 U19409 ( .IN1(n18366), .IN2(n18367), .Q(g25650) );
  AND2X1 U19410 ( .IN1(n18368), .IN2(n10789), .Q(n18367) );
  AND2X1 U19411 ( .IN1(n10059), .IN2(n18369), .Q(n18368) );
  OR2X1 U19412 ( .IN1(n18370), .IN2(g3050), .Q(n18369) );
  AND2X1 U19413 ( .IN1(n10060), .IN2(g8215), .Q(n18370) );
  INVX0 U19414 ( .INP(n18371), .ZN(n18366) );
  OR2X1 U19415 ( .IN1(n10739), .IN2(n10060), .Q(n18371) );
  OR2X1 U19416 ( .IN1(n18372), .IN2(n18373), .Q(g25649) );
  AND2X1 U19417 ( .IN1(n10907), .IN2(g3050), .Q(n18373) );
  AND2X1 U19418 ( .IN1(n10826), .IN2(g3338), .Q(n18372) );
  AND2X1 U19419 ( .IN1(g3179), .IN2(n10789), .Q(g25648) );
  OR2X1 U19420 ( .IN1(n5045), .IN2(n18374), .Q(g25639) );
  OR2X1 U19421 ( .IN1(n18375), .IN2(n18376), .Q(n18374) );
  AND2X1 U19422 ( .IN1(n15678), .IN2(n10789), .Q(n18376) );
  AND2X1 U19423 ( .IN1(g2719), .IN2(n5299), .Q(n15678) );
  AND2X1 U19424 ( .IN1(n10907), .IN2(g2715), .Q(n18375) );
  OR2X1 U19425 ( .IN1(n18377), .IN2(n18378), .Q(g25638) );
  AND2X1 U19426 ( .IN1(n18379), .IN2(n10789), .Q(n18378) );
  OR2X1 U19427 ( .IN1(n18380), .IN2(n18381), .Q(n18379) );
  AND2X1 U19428 ( .IN1(n18382), .IN2(n5441), .Q(n18381) );
  AND2X1 U19429 ( .IN1(n18383), .IN2(g1559), .Q(n18380) );
  AND2X1 U19430 ( .IN1(n10907), .IN2(g1564), .Q(n18377) );
  OR2X1 U19431 ( .IN1(n18384), .IN2(n18385), .Q(g25637) );
  AND2X1 U19432 ( .IN1(n18386), .IN2(g1559), .Q(n18385) );
  OR2X1 U19433 ( .IN1(n10878), .IN2(n18382), .Q(n18386) );
  AND2X1 U19434 ( .IN1(n18387), .IN2(n5768), .Q(n18382) );
  INVX0 U19435 ( .INP(n18383), .ZN(n18387) );
  AND2X1 U19436 ( .IN1(n18388), .IN2(n18383), .Q(n18384) );
  AND2X1 U19437 ( .IN1(n10827), .IN2(g1554), .Q(n18388) );
  OR2X1 U19438 ( .IN1(n18389), .IN2(n18390), .Q(g25636) );
  OR2X1 U19439 ( .IN1(n18391), .IN2(n18392), .Q(n18390) );
  AND2X1 U19440 ( .IN1(n18393), .IN2(n10789), .Q(n18392) );
  AND2X1 U19441 ( .IN1(n18394), .IN2(g1306), .Q(n18393) );
  OR2X1 U19442 ( .IN1(n5302), .IN2(n16675), .Q(n18394) );
  INVX0 U19443 ( .INP(n13407), .ZN(n16675) );
  AND2X1 U19444 ( .IN1(n10907), .IN2(g1521), .Q(n18391) );
  AND2X1 U19445 ( .IN1(n18395), .IN2(n13407), .Q(n18389) );
  AND2X1 U19446 ( .IN1(g1514), .IN2(test_so49), .Q(n13407) );
  OR2X1 U19447 ( .IN1(n18396), .IN2(n18397), .Q(g25635) );
  AND2X1 U19448 ( .IN1(n18398), .IN2(g1300), .Q(n18397) );
  OR2X1 U19449 ( .IN1(n18399), .IN2(n16665), .Q(n18398) );
  AND2X1 U19450 ( .IN1(n18400), .IN2(n10789), .Q(n18399) );
  OR2X1 U19451 ( .IN1(n5865), .IN2(n17827), .Q(n18400) );
  AND2X1 U19452 ( .IN1(n18401), .IN2(g1484), .Q(n18396) );
  OR2X1 U19453 ( .IN1(n10880), .IN2(n18402), .Q(n18401) );
  AND2X1 U19454 ( .IN1(n18403), .IN2(n18404), .Q(n18402) );
  INVX0 U19455 ( .INP(n17827), .ZN(n18404) );
  OR2X1 U19456 ( .IN1(n10433), .IN2(test_so12), .Q(n17827) );
  AND2X1 U19457 ( .IN1(n16668), .IN2(n5483), .Q(n18403) );
  AND2X1 U19458 ( .IN1(n18405), .IN2(n18406), .Q(g25634) );
  OR2X1 U19459 ( .IN1(n18407), .IN2(n18408), .Q(n18406) );
  AND2X1 U19460 ( .IN1(n10809), .IN2(g1395), .Q(n18408) );
  AND2X1 U19461 ( .IN1(n17868), .IN2(n18409), .Q(n18407) );
  INVX0 U19462 ( .INP(n18410), .ZN(n18409) );
  AND2X1 U19463 ( .IN1(n17851), .IN2(n10550), .Q(n18405) );
  OR2X1 U19464 ( .IN1(n18410), .IN2(n18411), .Q(n17851) );
  OR2X1 U19465 ( .IN1(n5655), .IN2(n10319), .Q(n18411) );
  OR2X1 U19466 ( .IN1(n18412), .IN2(n18413), .Q(g25633) );
  OR2X1 U19467 ( .IN1(n18414), .IN2(n18415), .Q(n18413) );
  AND2X1 U19468 ( .IN1(n10908), .IN2(g1379), .Q(n18415) );
  AND2X1 U19469 ( .IN1(n18416), .IN2(n10789), .Q(n18414) );
  AND2X1 U19470 ( .IN1(n18417), .IN2(g1384), .Q(n18416) );
  AND2X1 U19471 ( .IN1(n18418), .IN2(n17860), .Q(n18412) );
  AND2X1 U19472 ( .IN1(n17859), .IN2(n10504), .Q(n18418) );
  OR2X1 U19473 ( .IN1(n18419), .IN2(n18420), .Q(g25632) );
  AND2X1 U19474 ( .IN1(n17860), .IN2(n18421), .Q(n18420) );
  OR2X1 U19475 ( .IN1(n18422), .IN2(n16011), .Q(n18421) );
  AND2X1 U19476 ( .IN1(n18423), .IN2(n17513), .Q(n18422) );
  OR2X1 U19477 ( .IN1(n10459), .IN2(n10462), .Q(n18423) );
  AND2X1 U19478 ( .IN1(g1351), .IN2(n10789), .Q(n17860) );
  AND2X1 U19479 ( .IN1(n18424), .IN2(g1312), .Q(n18419) );
  OR2X1 U19480 ( .IN1(n10892), .IN2(n17859), .Q(n18424) );
  AND2X1 U19481 ( .IN1(n18425), .IN2(n10790), .Q(g25631) );
  OR2X1 U19482 ( .IN1(n18426), .IN2(n18427), .Q(n18425) );
  AND2X1 U19483 ( .IN1(n18417), .IN2(g1312), .Q(n18427) );
  AND2X1 U19484 ( .IN1(n18428), .IN2(n17510), .Q(n18426) );
  OR2X1 U19485 ( .IN1(n18429), .IN2(n18430), .Q(n18428) );
  INVX0 U19486 ( .INP(n18431), .ZN(n18430) );
  OR2X1 U19487 ( .IN1(g1351), .IN2(n4896), .Q(n18431) );
  OR2X1 U19488 ( .IN1(n18432), .IN2(n18433), .Q(n4896) );
  OR2X1 U19489 ( .IN1(n10089), .IN2(n17519), .Q(n18433) );
  OR2X1 U19490 ( .IN1(n10511), .IN2(n10121), .Q(n18432) );
  AND2X1 U19491 ( .IN1(n17517), .IN2(n17513), .Q(n18429) );
  OR2X1 U19492 ( .IN1(n10460), .IN2(n17518), .Q(n17513) );
  INVX0 U19493 ( .INP(n17519), .ZN(n17518) );
  AND2X1 U19494 ( .IN1(g1361), .IN2(n18434), .Q(n17517) );
  AND2X1 U19495 ( .IN1(g1351), .IN2(g1373), .Q(n18434) );
  OR2X1 U19496 ( .IN1(n18435), .IN2(n18436), .Q(g25630) );
  AND2X1 U19497 ( .IN1(g24247), .IN2(g1266), .Q(n18436) );
  INVX0 U19498 ( .INP(n18437), .ZN(n18435) );
  OR2X1 U19499 ( .IN1(n18438), .IN2(n10512), .Q(n18437) );
  AND2X1 U19500 ( .IN1(n10808), .IN2(n18439), .Q(n18438) );
  OR2X1 U19501 ( .IN1(g1266), .IN2(n5655), .Q(n18439) );
  OR2X1 U19502 ( .IN1(n18440), .IN2(n18441), .Q(g25629) );
  AND2X1 U19503 ( .IN1(n18442), .IN2(n10790), .Q(n18441) );
  OR2X1 U19504 ( .IN1(n18443), .IN2(n18444), .Q(n18442) );
  AND2X1 U19505 ( .IN1(n18445), .IN2(n5442), .Q(n18444) );
  AND2X1 U19506 ( .IN1(n18446), .IN2(g1216), .Q(n18443) );
  AND2X1 U19507 ( .IN1(n10909), .IN2(g1221), .Q(n18440) );
  OR2X1 U19508 ( .IN1(n18447), .IN2(n18448), .Q(g25628) );
  AND2X1 U19509 ( .IN1(n18449), .IN2(g1216), .Q(n18448) );
  OR2X1 U19510 ( .IN1(n10892), .IN2(n18445), .Q(n18449) );
  AND2X1 U19511 ( .IN1(n18450), .IN2(n10565), .Q(n18445) );
  AND2X1 U19512 ( .IN1(n18451), .IN2(test_so76), .Q(n18447) );
  AND2X1 U19513 ( .IN1(n18446), .IN2(n10790), .Q(n18451) );
  OR2X1 U19514 ( .IN1(n18452), .IN2(n18453), .Q(g25627) );
  AND2X1 U19515 ( .IN1(n18454), .IN2(n10790), .Q(n18453) );
  OR2X1 U19516 ( .IN1(n18455), .IN2(n18456), .Q(n18454) );
  AND2X1 U19517 ( .IN1(n18457), .IN2(g962), .Q(n18456) );
  INVX0 U19518 ( .INP(n18458), .ZN(n18455) );
  OR2X1 U19519 ( .IN1(n18457), .IN2(n10138), .Q(n18458) );
  OR2X1 U19520 ( .IN1(n5304), .IN2(n17894), .Q(n18457) );
  OR2X1 U19521 ( .IN1(n5599), .IN2(n5363), .Q(n17894) );
  AND2X1 U19522 ( .IN1(n10909), .IN2(g1178), .Q(n18452) );
  OR2X1 U19523 ( .IN1(n18459), .IN2(n18460), .Q(g25626) );
  AND2X1 U19524 ( .IN1(n18461), .IN2(g956), .Q(n18460) );
  OR2X1 U19525 ( .IN1(n18462), .IN2(n16715), .Q(n18461) );
  AND2X1 U19526 ( .IN1(n18463), .IN2(n10790), .Q(n18462) );
  OR2X1 U19527 ( .IN1(n5691), .IN2(n17883), .Q(n18463) );
  INVX0 U19528 ( .INP(n17902), .ZN(n17883) );
  AND2X1 U19529 ( .IN1(n18464), .IN2(g1141), .Q(n18459) );
  OR2X1 U19530 ( .IN1(n10892), .IN2(n18465), .Q(n18464) );
  AND2X1 U19531 ( .IN1(n18466), .IN2(n17902), .Q(n18465) );
  AND2X1 U19532 ( .IN1(test_so7), .IN2(n5618), .Q(n17902) );
  AND2X1 U19533 ( .IN1(n16718), .IN2(n5341), .Q(n18466) );
  AND2X1 U19534 ( .IN1(n18467), .IN2(n5320), .Q(g25625) );
  AND2X1 U19535 ( .IN1(n18468), .IN2(n17908), .Q(n18467) );
  OR2X1 U19536 ( .IN1(n18469), .IN2(n18470), .Q(n17908) );
  OR2X1 U19537 ( .IN1(n5654), .IN2(n10320), .Q(n18470) );
  OR2X1 U19538 ( .IN1(n18471), .IN2(n18472), .Q(n18468) );
  AND2X1 U19539 ( .IN1(n10810), .IN2(g1052), .Q(n18472) );
  AND2X1 U19540 ( .IN1(n17924), .IN2(n18473), .Q(n18471) );
  INVX0 U19541 ( .INP(n18469), .ZN(n18473) );
  OR2X1 U19542 ( .IN1(n18474), .IN2(n18475), .Q(g25624) );
  OR2X1 U19543 ( .IN1(n18476), .IN2(n18477), .Q(n18475) );
  AND2X1 U19544 ( .IN1(n10909), .IN2(g1036), .Q(n18477) );
  AND2X1 U19545 ( .IN1(n18478), .IN2(n10790), .Q(n18476) );
  AND2X1 U19546 ( .IN1(n18479), .IN2(g1041), .Q(n18478) );
  AND2X1 U19547 ( .IN1(n18480), .IN2(n17917), .Q(n18474) );
  AND2X1 U19548 ( .IN1(n17916), .IN2(n10505), .Q(n18480) );
  OR2X1 U19549 ( .IN1(n18481), .IN2(n18482), .Q(g25623) );
  AND2X1 U19550 ( .IN1(n17917), .IN2(n18483), .Q(n18482) );
  OR2X1 U19551 ( .IN1(n18484), .IN2(n16052), .Q(n18483) );
  AND2X1 U19552 ( .IN1(n18485), .IN2(n17536), .Q(n18484) );
  OR2X1 U19553 ( .IN1(n10458), .IN2(n10461), .Q(n18485) );
  AND2X1 U19554 ( .IN1(g1008), .IN2(n10790), .Q(n17917) );
  AND2X1 U19555 ( .IN1(test_so20), .IN2(n18486), .Q(n18481) );
  OR2X1 U19556 ( .IN1(n10891), .IN2(n17916), .Q(n18486) );
  AND2X1 U19557 ( .IN1(n18487), .IN2(n10790), .Q(g25622) );
  OR2X1 U19558 ( .IN1(n18488), .IN2(n18489), .Q(n18487) );
  AND2X1 U19559 ( .IN1(test_so20), .IN2(n18479), .Q(n18489) );
  AND2X1 U19560 ( .IN1(n18490), .IN2(n17531), .Q(n18488) );
  OR2X1 U19561 ( .IN1(n18491), .IN2(n18492), .Q(n18490) );
  INVX0 U19562 ( .INP(n18493), .ZN(n18492) );
  OR2X1 U19563 ( .IN1(g1008), .IN2(n4921), .Q(n18493) );
  OR2X1 U19564 ( .IN1(n18494), .IN2(n18495), .Q(n4921) );
  OR2X1 U19565 ( .IN1(n10090), .IN2(n17539), .Q(n18495) );
  OR2X1 U19566 ( .IN1(n10510), .IN2(n10122), .Q(n18494) );
  AND2X1 U19567 ( .IN1(n17541), .IN2(n17536), .Q(n18491) );
  OR2X1 U19568 ( .IN1(n10452), .IN2(n17540), .Q(n17536) );
  INVX0 U19569 ( .INP(n17539), .ZN(n17540) );
  AND2X1 U19570 ( .IN1(g1018), .IN2(n18496), .Q(n17541) );
  AND2X1 U19571 ( .IN1(g1008), .IN2(g1030), .Q(n18496) );
  OR2X1 U19572 ( .IN1(n18497), .IN2(n18498), .Q(g25621) );
  AND2X1 U19573 ( .IN1(g24231), .IN2(g921), .Q(n18498) );
  INVX0 U19574 ( .INP(n18499), .ZN(n18497) );
  OR2X1 U19575 ( .IN1(n18500), .IN2(n10513), .Q(n18499) );
  AND2X1 U19576 ( .IN1(n10810), .IN2(n18501), .Q(n18500) );
  OR2X1 U19577 ( .IN1(g921), .IN2(n5654), .Q(n18501) );
  AND2X1 U19578 ( .IN1(n18502), .IN2(g837), .Q(g25619) );
  OR2X1 U19579 ( .IN1(n10891), .IN2(n18503), .Q(n18502) );
  XNOR2X1 U19580 ( .IN1(n17977), .IN2(n10109), .Q(n18503) );
  OR2X1 U19581 ( .IN1(n18504), .IN2(n18505), .Q(g25618) );
  AND2X1 U19582 ( .IN1(n18506), .IN2(g817), .Q(n18505) );
  OR2X1 U19583 ( .IN1(n10891), .IN2(n18507), .Q(n18506) );
  AND2X1 U19584 ( .IN1(n18508), .IN2(n10419), .Q(n18507) );
  AND2X1 U19585 ( .IN1(n4948), .IN2(n16751), .Q(n18508) );
  AND2X1 U19586 ( .IN1(n18509), .IN2(g832), .Q(n18504) );
  OR2X1 U19587 ( .IN1(n18510), .IN2(n18511), .Q(n18509) );
  AND2X1 U19588 ( .IN1(n5822), .IN2(n4518), .Q(n18511) );
  AND2X1 U19589 ( .IN1(n10810), .IN2(n16751), .Q(n4518) );
  AND2X1 U19590 ( .IN1(n16813), .IN2(n16751), .Q(n18510) );
  OR2X1 U19591 ( .IN1(n18512), .IN2(n18513), .Q(g25617) );
  AND2X1 U19592 ( .IN1(n10909), .IN2(g812), .Q(n18513) );
  AND2X1 U19593 ( .IN1(n18514), .IN2(n16751), .Q(n18512) );
  OR2X1 U19594 ( .IN1(n18515), .IN2(n5709), .Q(n16751) );
  AND2X1 U19595 ( .IN1(n5733), .IN2(g837), .Q(n18515) );
  AND2X1 U19596 ( .IN1(n18516), .IN2(n18517), .Q(n18514) );
  OR2X1 U19597 ( .IN1(n16800), .IN2(g817), .Q(n18517) );
  OR2X1 U19598 ( .IN1(n5822), .IN2(n16813), .Q(n18516) );
  AND2X1 U19599 ( .IN1(n18518), .IN2(n10790), .Q(g25616) );
  AND2X1 U19600 ( .IN1(n18519), .IN2(n18520), .Q(n18518) );
  OR2X1 U19601 ( .IN1(n18521), .IN2(n18522), .Q(n18520) );
  INVX0 U19602 ( .INP(n18523), .ZN(n18519) );
  AND2X1 U19603 ( .IN1(n18522), .IN2(n18521), .Q(n18523) );
  AND2X1 U19604 ( .IN1(n17625), .IN2(g732), .Q(n18521) );
  OR2X1 U19605 ( .IN1(n18524), .IN2(n18525), .Q(n17625) );
  OR2X1 U19606 ( .IN1(g490), .IN2(g482), .Q(n18525) );
  OR2X1 U19607 ( .IN1(g528), .IN2(n18526), .Q(n18524) );
  OR2X1 U19608 ( .IN1(n17600), .IN2(n17594), .Q(n18526) );
  OR2X1 U19609 ( .IN1(test_so54), .IN2(g518), .Q(n17600) );
  XOR2X1 U19610 ( .IN1(n18527), .IN2(n18528), .Q(n18522) );
  XOR2X1 U19611 ( .IN1(n18529), .IN2(n18530), .Q(n18528) );
  XNOR2X1 U19612 ( .IN1(g239), .IN2(n10270), .Q(n18530) );
  XNOR2X1 U19613 ( .IN1(g246), .IN2(n5597), .Q(n18529) );
  XNOR2X1 U19614 ( .IN1(n10152), .IN2(n18531), .Q(n18527) );
  XNOR2X1 U19615 ( .IN1(g269), .IN2(n10153), .Q(n18531) );
  OR2X1 U19616 ( .IN1(n18532), .IN2(n18533), .Q(g25615) );
  AND2X1 U19617 ( .IN1(n18534), .IN2(g686), .Q(n18533) );
  AND2X1 U19618 ( .IN1(n17586), .IN2(g667), .Q(n18532) );
  OR2X1 U19619 ( .IN1(n18535), .IN2(n18536), .Q(g25614) );
  OR2X1 U19620 ( .IN1(n18537), .IN2(n18538), .Q(n18536) );
  AND2X1 U19621 ( .IN1(n5111), .IN2(n18539), .Q(n18538) );
  AND2X1 U19622 ( .IN1(n17586), .IN2(g686), .Q(n18537) );
  AND2X1 U19623 ( .IN1(n10909), .IN2(g691), .Q(n18535) );
  OR2X1 U19624 ( .IN1(n18540), .IN2(n18541), .Q(g25613) );
  AND2X1 U19625 ( .IN1(n10909), .IN2(g559), .Q(n18541) );
  AND2X1 U19626 ( .IN1(n18542), .IN2(n18543), .Q(n18540) );
  XNOR2X1 U19627 ( .IN1(n18003), .IN2(g562), .Q(n18543) );
  OR2X1 U19628 ( .IN1(n18544), .IN2(n10477), .Q(n18003) );
  AND2X1 U19629 ( .IN1(n10006), .IN2(g12368), .Q(n18544) );
  AND2X1 U19630 ( .IN1(n2421), .IN2(n18545), .Q(n18542) );
  OR2X1 U19631 ( .IN1(n5288), .IN2(n19032), .Q(n18545) );
  OR2X1 U19632 ( .IN1(n18546), .IN2(n18547), .Q(g25612) );
  AND2X1 U19633 ( .IN1(n17586), .IN2(g518), .Q(n18547) );
  AND2X1 U19634 ( .IN1(n18548), .IN2(g513), .Q(n18546) );
  OR2X1 U19635 ( .IN1(n18549), .IN2(n18550), .Q(g25611) );
  AND2X1 U19636 ( .IN1(n17586), .IN2(g513), .Q(n18550) );
  AND2X1 U19637 ( .IN1(n18548), .IN2(g504), .Q(n18549) );
  OR2X1 U19638 ( .IN1(n10891), .IN2(n18551), .Q(n18548) );
  AND2X1 U19639 ( .IN1(n18539), .IN2(n18008), .Q(n18551) );
  INVX0 U19640 ( .INP(n4962), .ZN(n18008) );
  OR2X1 U19641 ( .IN1(n18552), .IN2(n18553), .Q(g25610) );
  OR2X1 U19642 ( .IN1(n18554), .IN2(n18555), .Q(n18553) );
  AND2X1 U19643 ( .IN1(test_so54), .IN2(n18534), .Q(n18555) );
  INVX0 U19644 ( .INP(n17586), .ZN(n18534) );
  AND2X1 U19645 ( .IN1(n17586), .IN2(g504), .Q(n18554) );
  OR2X1 U19646 ( .IN1(n18556), .IN2(n18557), .Q(g25609) );
  OR2X1 U19647 ( .IN1(n18552), .IN2(n18558), .Q(n18557) );
  AND2X1 U19648 ( .IN1(test_so54), .IN2(n18559), .Q(n18558) );
  OR2X1 U19649 ( .IN1(n18560), .IN2(n17586), .Q(n18559) );
  AND2X1 U19650 ( .IN1(n10811), .IN2(n18013), .Q(n17586) );
  AND2X1 U19651 ( .IN1(n5548), .IN2(n10791), .Q(n18560) );
  AND2X1 U19652 ( .IN1(n17577), .IN2(n4962), .Q(n18552) );
  AND2X1 U19653 ( .IN1(n17577), .IN2(n5287), .Q(n18556) );
  AND2X1 U19654 ( .IN1(n10811), .IN2(n18539), .Q(n17577) );
  INVX0 U19655 ( .INP(n18013), .ZN(n18539) );
  OR2X1 U19656 ( .IN1(g376), .IN2(n18561), .Q(n18013) );
  OR2X1 U19657 ( .IN1(n5632), .IN2(n10526), .Q(n18561) );
  OR2X1 U19658 ( .IN1(n18562), .IN2(n18563), .Q(g25605) );
  OR2X1 U19659 ( .IN1(n18564), .IN2(n18565), .Q(n18563) );
  AND2X1 U19660 ( .IN1(n18566), .IN2(n10791), .Q(n18565) );
  AND2X1 U19661 ( .IN1(n18567), .IN2(g246), .Q(n18566) );
  AND2X1 U19662 ( .IN1(n10909), .IN2(g168), .Q(n18564) );
  AND2X1 U19663 ( .IN1(n18568), .IN2(g460), .Q(n18562) );
  OR2X1 U19664 ( .IN1(n18569), .IN2(n18570), .Q(g25604) );
  AND2X1 U19665 ( .IN1(n18571), .IN2(g460), .Q(n18570) );
  AND2X1 U19666 ( .IN1(n18568), .IN2(g452), .Q(n18569) );
  OR2X1 U19667 ( .IN1(n18572), .IN2(n18573), .Q(g25602) );
  OR2X1 U19668 ( .IN1(n18574), .IN2(n18575), .Q(n18573) );
  AND2X1 U19669 ( .IN1(n18576), .IN2(n10791), .Q(n18575) );
  AND2X1 U19670 ( .IN1(n18567), .IN2(g446), .Q(n18576) );
  INVX0 U19671 ( .INP(n17594), .ZN(n18567) );
  AND2X1 U19672 ( .IN1(n10909), .IN2(g405), .Q(n18574) );
  AND2X1 U19673 ( .IN1(n18568), .IN2(test_so72), .Q(n18572) );
  OR2X1 U19674 ( .IN1(n18577), .IN2(n18578), .Q(g25601) );
  AND2X1 U19675 ( .IN1(test_so72), .IN2(n18571), .Q(n18578) );
  AND2X1 U19676 ( .IN1(n18568), .IN2(g174), .Q(n18577) );
  OR2X1 U19677 ( .IN1(n18579), .IN2(n18580), .Q(g25600) );
  AND2X1 U19678 ( .IN1(n18571), .IN2(g174), .Q(n18580) );
  INVX0 U19679 ( .INP(n18568), .ZN(n18571) );
  AND2X1 U19680 ( .IN1(n18568), .IN2(g168), .Q(n18579) );
  AND2X1 U19681 ( .IN1(n10811), .IN2(n17594), .Q(n18568) );
  OR2X1 U19682 ( .IN1(n5121), .IN2(g370), .Q(n17594) );
  OR2X1 U19683 ( .IN1(n18581), .IN2(n18582), .Q(g25599) );
  AND2X1 U19684 ( .IN1(n10909), .IN2(g385), .Q(n18581) );
  OR2X1 U19685 ( .IN1(n18583), .IN2(n18584), .Q(g25598) );
  AND2X1 U19686 ( .IN1(n18585), .IN2(g376), .Q(n18584) );
  OR2X1 U19687 ( .IN1(n10891), .IN2(n18586), .Q(n18585) );
  AND2X1 U19688 ( .IN1(n5121), .IN2(g358), .Q(n18586) );
  AND2X1 U19689 ( .IN1(n18587), .IN2(n5121), .Q(n18583) );
  OR2X1 U19690 ( .IN1(n10526), .IN2(n18588), .Q(n5121) );
  AND2X1 U19691 ( .IN1(n10811), .IN2(g385), .Q(n18587) );
  OR2X1 U19692 ( .IN1(n18589), .IN2(n18590), .Q(g25597) );
  AND2X1 U19693 ( .IN1(n18591), .IN2(n10791), .Q(n18590) );
  XNOR2X1 U19694 ( .IN1(n18582), .IN2(n10156), .Q(n18591) );
  INVX0 U19695 ( .INP(n12083), .ZN(n18582) );
  OR2X1 U19696 ( .IN1(n10155), .IN2(n18588), .Q(n12083) );
  OR2X1 U19697 ( .IN1(n5633), .IN2(n5632), .Q(n18588) );
  AND2X1 U19698 ( .IN1(n10909), .IN2(g358), .Q(n18589) );
  OR2X1 U19699 ( .IN1(n18592), .IN2(n18593), .Q(g25596) );
  AND2X1 U19700 ( .IN1(n18594), .IN2(n10791), .Q(n18593) );
  XNOR2X1 U19701 ( .IN1(g376), .IN2(n10526), .Q(n18594) );
  AND2X1 U19702 ( .IN1(n10909), .IN2(g370), .Q(n18592) );
  AND2X1 U19703 ( .IN1(n18595), .IN2(n10155), .Q(g25595) );
  AND2X1 U19704 ( .IN1(n10526), .IN2(n10791), .Q(n18595) );
  AND2X1 U19705 ( .IN1(n18596), .IN2(n17620), .Q(g25594) );
  OR2X1 U19706 ( .IN1(n18597), .IN2(g278), .Q(n17620) );
  AND2X1 U19707 ( .IN1(n18598), .IN2(n18599), .Q(n18597) );
  AND2X1 U19708 ( .IN1(n18600), .IN2(n18601), .Q(n18599) );
  AND2X1 U19709 ( .IN1(g262), .IN2(g269), .Q(n18601) );
  AND2X1 U19710 ( .IN1(n10270), .IN2(g255), .Q(n18600) );
  AND2X1 U19711 ( .IN1(n18602), .IN2(n6008), .Q(n18598) );
  AND2X1 U19712 ( .IN1(n5597), .IN2(n10271), .Q(n18602) );
  AND2X1 U19713 ( .IN1(n17619), .IN2(n10791), .Q(n18596) );
  OR2X1 U19714 ( .IN1(n18603), .IN2(n18604), .Q(n17619) );
  OR2X1 U19715 ( .IN1(g269), .IN2(n18605), .Q(n18604) );
  OR2X1 U19716 ( .IN1(g255), .IN2(g262), .Q(n18605) );
  OR2X1 U19717 ( .IN1(n18606), .IN2(n18607), .Q(n18603) );
  OR2X1 U19718 ( .IN1(n10271), .IN2(n10270), .Q(n18607) );
  OR2X1 U19719 ( .IN1(n6008), .IN2(n5597), .Q(n18606) );
  OR2X1 U19720 ( .IN1(n18608), .IN2(n18609), .Q(g25593) );
  AND2X1 U19721 ( .IN1(n18610), .IN2(n10791), .Q(n18609) );
  OR2X1 U19722 ( .IN1(n18611), .IN2(n18612), .Q(n18610) );
  AND2X1 U19723 ( .IN1(n18613), .IN2(n18614), .Q(n18612) );
  INVX0 U19724 ( .INP(n18615), .ZN(n18614) );
  AND2X1 U19725 ( .IN1(n18615), .IN2(g209), .Q(n18611) );
  AND2X1 U19726 ( .IN1(n10909), .IN2(g191), .Q(n18608) );
  OR2X1 U19727 ( .IN1(n18616), .IN2(n18617), .Q(g25592) );
  AND2X1 U19728 ( .IN1(n18618), .IN2(n10791), .Q(n18617) );
  XOR2X1 U19729 ( .IN1(n18619), .IN2(n10139), .Q(n18618) );
  OR2X1 U19730 ( .IN1(n18615), .IN2(n18613), .Q(n18619) );
  XOR2X1 U19731 ( .IN1(n10139), .IN2(n10140), .Q(n18613) );
  OR2X1 U19732 ( .IN1(n10422), .IN2(n10421), .Q(n18615) );
  AND2X1 U19733 ( .IN1(n10910), .IN2(g222), .Q(n18616) );
  OR2X1 U19734 ( .IN1(n18620), .IN2(n18621), .Q(g25591) );
  AND2X1 U19735 ( .IN1(n10910), .IN2(g209), .Q(n18621) );
  AND2X1 U19736 ( .IN1(n10422), .IN2(n10792), .Q(n18620) );
  INVX0 U19737 ( .INP(n15975), .ZN(g25167) );
  OR2X1 U19738 ( .IN1(n10556), .IN2(g1657), .Q(n15975) );
  AND2X1 U19739 ( .IN1(n18622), .IN2(g6732), .Q(g24355) );
  OR2X1 U19740 ( .IN1(n10890), .IN2(n18623), .Q(n18622) );
  OR2X1 U19741 ( .IN1(n18624), .IN2(n18625), .Q(g24354) );
  AND2X1 U19742 ( .IN1(n18626), .IN2(n10792), .Q(n18625) );
  AND2X1 U19743 ( .IN1(n10495), .IN2(n18623), .Q(n18626) );
  OR2X1 U19744 ( .IN1(n5531), .IN2(n18627), .Q(n18623) );
  AND2X1 U19745 ( .IN1(n10910), .IN2(g6727), .Q(n18624) );
  OR2X1 U19746 ( .IN1(n18628), .IN2(n18629), .Q(g24353) );
  AND2X1 U19747 ( .IN1(n18630), .IN2(n10792), .Q(n18629) );
  XNOR2X1 U19748 ( .IN1(g6727), .IN2(n18627), .Q(n18630) );
  OR2X1 U19749 ( .IN1(n18631), .IN2(n18632), .Q(n18627) );
  OR2X1 U19750 ( .IN1(n10243), .IN2(n10557), .Q(n18632) );
  OR2X1 U19751 ( .IN1(n5700), .IN2(n10257), .Q(n18631) );
  AND2X1 U19752 ( .IN1(n10910), .IN2(g6723), .Q(n18628) );
  AND2X1 U19753 ( .IN1(n18633), .IN2(n18634), .Q(g24352) );
  AND2X1 U19754 ( .IN1(n18635), .IN2(n10342), .Q(n18634) );
  AND2X1 U19755 ( .IN1(n10243), .IN2(n10792), .Q(n18635) );
  AND2X1 U19756 ( .IN1(n18636), .IN2(n10369), .Q(n18633) );
  AND2X1 U19757 ( .IN1(n18637), .IN2(n18638), .Q(n18636) );
  OR2X1 U19758 ( .IN1(test_so80), .IN2(n5700), .Q(n18638) );
  OR2X1 U19759 ( .IN1(n10257), .IN2(g14828), .Q(n18637) );
  AND2X1 U19760 ( .IN1(n18639), .IN2(g6386), .Q(g24351) );
  OR2X1 U19761 ( .IN1(n10889), .IN2(n18640), .Q(n18639) );
  OR2X1 U19762 ( .IN1(n18641), .IN2(n18642), .Q(g24350) );
  AND2X1 U19763 ( .IN1(n18643), .IN2(n10792), .Q(n18642) );
  AND2X1 U19764 ( .IN1(n10488), .IN2(n18640), .Q(n18643) );
  OR2X1 U19765 ( .IN1(n10563), .IN2(n18644), .Q(n18640) );
  AND2X1 U19766 ( .IN1(test_so69), .IN2(n10894), .Q(n18641) );
  OR2X1 U19767 ( .IN1(n18645), .IN2(n18646), .Q(g24349) );
  AND2X1 U19768 ( .IN1(n18647), .IN2(n10792), .Q(n18646) );
  XNOR2X1 U19769 ( .IN1(test_so69), .IN2(n18644), .Q(n18647) );
  OR2X1 U19770 ( .IN1(n18648), .IN2(n18649), .Q(n18644) );
  OR2X1 U19771 ( .IN1(n10261), .IN2(n10246), .Q(n18649) );
  OR2X1 U19772 ( .IN1(n5703), .IN2(n5437), .Q(n18648) );
  AND2X1 U19773 ( .IN1(n10910), .IN2(g6377), .Q(n18645) );
  AND2X1 U19774 ( .IN1(n18650), .IN2(n18651), .Q(g24348) );
  AND2X1 U19775 ( .IN1(n18652), .IN2(n10350), .Q(n18651) );
  AND2X1 U19776 ( .IN1(n10246), .IN2(n10792), .Q(n18652) );
  AND2X1 U19777 ( .IN1(n18653), .IN2(n10377), .Q(n18650) );
  AND2X1 U19778 ( .IN1(n18654), .IN2(n18655), .Q(n18653) );
  OR2X1 U19779 ( .IN1(n5703), .IN2(g12422), .Q(n18655) );
  OR2X1 U19780 ( .IN1(n10261), .IN2(g14779), .Q(n18654) );
  AND2X1 U19781 ( .IN1(n18656), .IN2(g6040), .Q(g24347) );
  OR2X1 U19782 ( .IN1(n10889), .IN2(n18657), .Q(n18656) );
  OR2X1 U19783 ( .IN1(n18658), .IN2(n18659), .Q(g24346) );
  AND2X1 U19784 ( .IN1(n18660), .IN2(n10792), .Q(n18659) );
  AND2X1 U19785 ( .IN1(n18657), .IN2(n10579), .Q(n18660) );
  OR2X1 U19786 ( .IN1(n5528), .IN2(n18661), .Q(n18657) );
  AND2X1 U19787 ( .IN1(n10910), .IN2(g6035), .Q(n18658) );
  OR2X1 U19788 ( .IN1(n18662), .IN2(n18663), .Q(g24345) );
  AND2X1 U19789 ( .IN1(n18664), .IN2(n10792), .Q(n18663) );
  XNOR2X1 U19790 ( .IN1(n18661), .IN2(g6035), .Q(n18664) );
  OR2X1 U19791 ( .IN1(n18665), .IN2(n18666), .Q(n18661) );
  OR2X1 U19792 ( .IN1(n10252), .IN2(n10237), .Q(n18666) );
  OR2X1 U19793 ( .IN1(n5698), .IN2(n5432), .Q(n18665) );
  AND2X1 U19794 ( .IN1(n10910), .IN2(g6031), .Q(n18662) );
  AND2X1 U19795 ( .IN1(n18667), .IN2(n18668), .Q(g24344) );
  AND2X1 U19796 ( .IN1(n18669), .IN2(n10331), .Q(n18668) );
  AND2X1 U19797 ( .IN1(n10237), .IN2(n10793), .Q(n18669) );
  AND2X1 U19798 ( .IN1(n18670), .IN2(n10357), .Q(n18667) );
  AND2X1 U19799 ( .IN1(n18671), .IN2(n18672), .Q(n18670) );
  OR2X1 U19800 ( .IN1(n5698), .IN2(g12350), .Q(n18672) );
  OR2X1 U19801 ( .IN1(n10252), .IN2(g14738), .Q(n18671) );
  AND2X1 U19802 ( .IN1(n18673), .IN2(g5694), .Q(g24343) );
  OR2X1 U19803 ( .IN1(n10889), .IN2(n18674), .Q(n18673) );
  OR2X1 U19804 ( .IN1(n18675), .IN2(n18676), .Q(g24342) );
  AND2X1 U19805 ( .IN1(n18677), .IN2(n10793), .Q(n18676) );
  AND2X1 U19806 ( .IN1(n10496), .IN2(n18674), .Q(n18677) );
  OR2X1 U19807 ( .IN1(n5529), .IN2(n18678), .Q(n18674) );
  AND2X1 U19808 ( .IN1(n10910), .IN2(g5689), .Q(n18675) );
  OR2X1 U19809 ( .IN1(n18679), .IN2(n18680), .Q(g24341) );
  AND2X1 U19810 ( .IN1(n18681), .IN2(n10798), .Q(n18680) );
  XNOR2X1 U19811 ( .IN1(n18678), .IN2(g5689), .Q(n18681) );
  OR2X1 U19812 ( .IN1(n18682), .IN2(n18683), .Q(n18678) );
  OR2X1 U19813 ( .IN1(n10254), .IN2(n10239), .Q(n18683) );
  OR2X1 U19814 ( .IN1(n5705), .IN2(n5439), .Q(n18682) );
  AND2X1 U19815 ( .IN1(n10899), .IN2(g5685), .Q(n18679) );
  AND2X1 U19816 ( .IN1(n18684), .IN2(n18685), .Q(g24340) );
  AND2X1 U19817 ( .IN1(n18686), .IN2(n10335), .Q(n18685) );
  AND2X1 U19818 ( .IN1(n10239), .IN2(n10793), .Q(n18686) );
  AND2X1 U19819 ( .IN1(n18687), .IN2(n10361), .Q(n18684) );
  AND2X1 U19820 ( .IN1(n18688), .IN2(n18689), .Q(n18687) );
  OR2X1 U19821 ( .IN1(n5705), .IN2(g12300), .Q(n18689) );
  OR2X1 U19822 ( .IN1(n10254), .IN2(g14694), .Q(n18688) );
  AND2X1 U19823 ( .IN1(n18690), .IN2(g5348), .Q(g24339) );
  OR2X1 U19824 ( .IN1(n10889), .IN2(n18691), .Q(n18690) );
  OR2X1 U19825 ( .IN1(n18692), .IN2(n18693), .Q(g24338) );
  AND2X1 U19826 ( .IN1(n18694), .IN2(n10793), .Q(n18693) );
  AND2X1 U19827 ( .IN1(n10514), .IN2(n18691), .Q(n18694) );
  OR2X1 U19828 ( .IN1(n10562), .IN2(n18695), .Q(n18691) );
  AND2X1 U19829 ( .IN1(test_so10), .IN2(n10893), .Q(n18692) );
  OR2X1 U19830 ( .IN1(n18696), .IN2(n18697), .Q(g24337) );
  AND2X1 U19831 ( .IN1(n18698), .IN2(n10793), .Q(n18697) );
  XNOR2X1 U19832 ( .IN1(test_so10), .IN2(n18695), .Q(n18698) );
  OR2X1 U19833 ( .IN1(n18699), .IN2(n18700), .Q(n18695) );
  OR2X1 U19834 ( .IN1(n10250), .IN2(n10235), .Q(n18700) );
  OR2X1 U19835 ( .IN1(n5704), .IN2(n5438), .Q(n18699) );
  AND2X1 U19836 ( .IN1(n10897), .IN2(g5339), .Q(n18696) );
  AND2X1 U19837 ( .IN1(n18701), .IN2(n18702), .Q(g24336) );
  AND2X1 U19838 ( .IN1(n18703), .IN2(n10306), .Q(n18702) );
  AND2X1 U19839 ( .IN1(n10235), .IN2(n10793), .Q(n18703) );
  AND2X1 U19840 ( .IN1(n18704), .IN2(n10327), .Q(n18701) );
  AND2X1 U19841 ( .IN1(n18705), .IN2(n18706), .Q(n18704) );
  OR2X1 U19842 ( .IN1(n5704), .IN2(g12238), .Q(n18706) );
  OR2X1 U19843 ( .IN1(n10250), .IN2(g14662), .Q(n18705) );
  OR2X1 U19844 ( .IN1(n18707), .IN2(n18708), .Q(g24335) );
  AND2X1 U19845 ( .IN1(n10897), .IN2(g18881), .Q(n18708) );
  AND2X1 U19846 ( .IN1(n18709), .IN2(n18710), .Q(n18707) );
  AND2X1 U19847 ( .IN1(n5653), .IN2(g4643), .Q(n18709) );
  OR2X1 U19848 ( .IN1(n18711), .IN2(n18712), .Q(g24334) );
  AND2X1 U19849 ( .IN1(n10897), .IN2(g4358), .Q(n18712) );
  AND2X1 U19850 ( .IN1(n18713), .IN2(n18714), .Q(n18711) );
  AND2X1 U19851 ( .IN1(n18715), .IN2(n18716), .Q(n18714) );
  AND2X1 U19852 ( .IN1(n18717), .IN2(n11934), .Q(n18716) );
  AND2X1 U19853 ( .IN1(n5727), .IN2(test_so3), .Q(n11934) );
  AND2X1 U19854 ( .IN1(g4340), .IN2(g4633), .Q(n18717) );
  AND2X1 U19855 ( .IN1(n5303), .IN2(n5365), .Q(n18715) );
  AND2X1 U19856 ( .IN1(n18718), .IN2(n18719), .Q(n18713) );
  AND2X1 U19857 ( .IN1(n5274), .IN2(n5539), .Q(n18719) );
  AND2X1 U19858 ( .IN1(n18710), .IN2(n5608), .Q(n18718) );
  INVX0 U19859 ( .INP(n18720), .ZN(n18710) );
  OR2X1 U19860 ( .IN1(n18721), .IN2(n18722), .Q(n18720) );
  OR2X1 U19861 ( .IN1(g4358), .IN2(n18723), .Q(n18722) );
  OR2X1 U19862 ( .IN1(g4332), .IN2(g4311), .Q(n18723) );
  OR2X1 U19863 ( .IN1(g4322), .IN2(n18724), .Q(n18721) );
  OR2X1 U19864 ( .IN1(test_so81), .IN2(n10876), .Q(n18724) );
  AND2X1 U19865 ( .IN1(n10897), .IN2(g4392), .Q(g24298) );
  OR2X1 U19866 ( .IN1(n18725), .IN2(n18726), .Q(g24282) );
  AND2X1 U19867 ( .IN1(g24281), .IN2(g9251), .Q(n18726) );
  AND2X1 U19868 ( .IN1(n18727), .IN2(g4308), .Q(n18725) );
  OR2X1 U19869 ( .IN1(n10389), .IN2(n10876), .Q(n18727) );
  AND2X1 U19870 ( .IN1(n10812), .IN2(n10418), .Q(g24281) );
  OR2X1 U19871 ( .IN1(n18728), .IN2(n18729), .Q(g24280) );
  AND2X1 U19872 ( .IN1(n18730), .IN2(g4273), .Q(n18729) );
  OR2X1 U19873 ( .IN1(n18731), .IN2(n18732), .Q(n18730) );
  AND2X1 U19874 ( .IN1(n5763), .IN2(n10793), .Q(n18731) );
  AND2X1 U19875 ( .IN1(n18733), .IN2(g4269), .Q(n18728) );
  OR2X1 U19876 ( .IN1(n10888), .IN2(n18734), .Q(n18733) );
  AND2X1 U19877 ( .IN1(n18735), .IN2(n5764), .Q(n18734) );
  AND2X1 U19878 ( .IN1(g4258), .IN2(g4264), .Q(n18735) );
  OR2X1 U19879 ( .IN1(n18736), .IN2(n18737), .Q(g24279) );
  AND2X1 U19880 ( .IN1(n18738), .IN2(n10793), .Q(n18737) );
  XOR2X1 U19881 ( .IN1(n18739), .IN2(n18740), .Q(n18738) );
  AND2X1 U19882 ( .IN1(n18741), .IN2(n18742), .Q(n18740) );
  OR2X1 U19883 ( .IN1(n5726), .IN2(n10455), .Q(n18742) );
  OR2X1 U19884 ( .IN1(g8870), .IN2(n18743), .Q(n18741) );
  OR2X1 U19885 ( .IN1(n18744), .IN2(g4235), .Q(n18743) );
  AND2X1 U19886 ( .IN1(n18745), .IN2(n18746), .Q(n18744) );
  AND2X1 U19887 ( .IN1(n18747), .IN2(n18748), .Q(n18746) );
  AND2X1 U19888 ( .IN1(n19038), .IN2(n19039), .Q(n18748) );
  AND2X1 U19889 ( .IN1(n19036), .IN2(n19037), .Q(n18747) );
  AND2X1 U19890 ( .IN1(n18749), .IN2(n19033), .Q(n18745) );
  AND2X1 U19891 ( .IN1(n19034), .IN2(n19035), .Q(n18749) );
  AND2X1 U19892 ( .IN1(n10897), .IN2(g4235), .Q(n18736) );
  AND2X1 U19893 ( .IN1(n18750), .IN2(g4045), .Q(g24278) );
  OR2X1 U19894 ( .IN1(n10888), .IN2(n18751), .Q(n18750) );
  OR2X1 U19895 ( .IN1(n18752), .IN2(n18753), .Q(g24277) );
  AND2X1 U19896 ( .IN1(n18754), .IN2(n10794), .Q(n18753) );
  AND2X1 U19897 ( .IN1(n10490), .IN2(n18751), .Q(n18754) );
  OR2X1 U19898 ( .IN1(n5530), .IN2(n18755), .Q(n18751) );
  AND2X1 U19899 ( .IN1(n10898), .IN2(g4040), .Q(n18752) );
  OR2X1 U19900 ( .IN1(n18756), .IN2(n18757), .Q(g24276) );
  AND2X1 U19901 ( .IN1(n18758), .IN2(n10794), .Q(n18757) );
  XNOR2X1 U19902 ( .IN1(n18755), .IN2(g4040), .Q(n18758) );
  OR2X1 U19903 ( .IN1(n18759), .IN2(n18760), .Q(n18755) );
  OR2X1 U19904 ( .IN1(n10255), .IN2(n10241), .Q(n18760) );
  OR2X1 U19905 ( .IN1(n5701), .IN2(n5435), .Q(n18759) );
  AND2X1 U19906 ( .IN1(n10897), .IN2(g4031), .Q(n18756) );
  AND2X1 U19907 ( .IN1(n18761), .IN2(n18762), .Q(g24275) );
  AND2X1 U19908 ( .IN1(n18763), .IN2(n10338), .Q(n18762) );
  AND2X1 U19909 ( .IN1(n10241), .IN2(n10794), .Q(n18763) );
  AND2X1 U19910 ( .IN1(n18764), .IN2(n10365), .Q(n18761) );
  AND2X1 U19911 ( .IN1(n18765), .IN2(n18766), .Q(n18764) );
  OR2X1 U19912 ( .IN1(n5701), .IN2(g11418), .Q(n18766) );
  OR2X1 U19913 ( .IN1(n10255), .IN2(g13966), .Q(n18765) );
  AND2X1 U19914 ( .IN1(n18767), .IN2(g3694), .Q(g24274) );
  OR2X1 U19915 ( .IN1(n10888), .IN2(n18768), .Q(n18767) );
  OR2X1 U19916 ( .IN1(n18769), .IN2(n18770), .Q(g24273) );
  AND2X1 U19917 ( .IN1(n18771), .IN2(n10794), .Q(n18770) );
  AND2X1 U19918 ( .IN1(n10498), .IN2(n18768), .Q(n18771) );
  OR2X1 U19919 ( .IN1(n5532), .IN2(n18772), .Q(n18768) );
  AND2X1 U19920 ( .IN1(n10898), .IN2(g3689), .Q(n18769) );
  OR2X1 U19921 ( .IN1(n18773), .IN2(n18774), .Q(g24272) );
  AND2X1 U19922 ( .IN1(n18775), .IN2(n10794), .Q(n18774) );
  XNOR2X1 U19923 ( .IN1(n18772), .IN2(g3689), .Q(n18775) );
  OR2X1 U19924 ( .IN1(n18776), .IN2(n18777), .Q(n18772) );
  OR2X1 U19925 ( .IN1(n10259), .IN2(n10245), .Q(n18777) );
  OR2X1 U19926 ( .IN1(n5699), .IN2(n5433), .Q(n18776) );
  AND2X1 U19927 ( .IN1(n10898), .IN2(g3680), .Q(n18773) );
  AND2X1 U19928 ( .IN1(n18778), .IN2(n18779), .Q(g24271) );
  AND2X1 U19929 ( .IN1(n18780), .IN2(n10346), .Q(n18779) );
  AND2X1 U19930 ( .IN1(n10245), .IN2(n10794), .Q(n18780) );
  AND2X1 U19931 ( .IN1(n18781), .IN2(n10373), .Q(n18778) );
  AND2X1 U19932 ( .IN1(n18782), .IN2(n18783), .Q(n18781) );
  OR2X1 U19933 ( .IN1(n5699), .IN2(g11388), .Q(n18783) );
  OR2X1 U19934 ( .IN1(n10259), .IN2(g13926), .Q(n18782) );
  AND2X1 U19935 ( .IN1(n18784), .IN2(g3343), .Q(g24270) );
  OR2X1 U19936 ( .IN1(n10888), .IN2(n18785), .Q(n18784) );
  OR2X1 U19937 ( .IN1(n18786), .IN2(n18787), .Q(g24269) );
  AND2X1 U19938 ( .IN1(n18788), .IN2(n10794), .Q(n18787) );
  AND2X1 U19939 ( .IN1(n10487), .IN2(n18785), .Q(n18788) );
  OR2X1 U19940 ( .IN1(n5527), .IN2(n18789), .Q(n18785) );
  AND2X1 U19941 ( .IN1(n10898), .IN2(g3338), .Q(n18786) );
  OR2X1 U19942 ( .IN1(n18790), .IN2(n18791), .Q(g24268) );
  AND2X1 U19943 ( .IN1(n18792), .IN2(n10794), .Q(n18791) );
  XNOR2X1 U19944 ( .IN1(n18789), .IN2(g3338), .Q(n18792) );
  OR2X1 U19945 ( .IN1(n18793), .IN2(n18794), .Q(n18789) );
  OR2X1 U19946 ( .IN1(n10248), .IN2(n10233), .Q(n18794) );
  OR2X1 U19947 ( .IN1(n5702), .IN2(n5436), .Q(n18793) );
  AND2X1 U19948 ( .IN1(test_so91), .IN2(n10894), .Q(n18790) );
  AND2X1 U19949 ( .IN1(n18795), .IN2(n18796), .Q(g24267) );
  AND2X1 U19950 ( .IN1(n18797), .IN2(n10323), .Q(n18796) );
  AND2X1 U19951 ( .IN1(n10233), .IN2(n10794), .Q(n18797) );
  AND2X1 U19952 ( .IN1(n18798), .IN2(n10353), .Q(n18795) );
  AND2X1 U19953 ( .IN1(n18799), .IN2(n18800), .Q(n18798) );
  OR2X1 U19954 ( .IN1(n5702), .IN2(g11349), .Q(n18800) );
  OR2X1 U19955 ( .IN1(n10248), .IN2(g13895), .Q(n18799) );
  OR2X1 U19956 ( .IN1(n18801), .IN2(n18802), .Q(g24266) );
  AND2X1 U19957 ( .IN1(n18803), .IN2(n10795), .Q(n18802) );
  AND2X1 U19958 ( .IN1(test_so9), .IN2(n10493), .Q(n18803) );
  INVX0 U19959 ( .INP(n18804), .ZN(n18801) );
  OR2X1 U19960 ( .IN1(n10740), .IN2(n5963), .Q(n18804) );
  OR2X1 U19961 ( .IN1(n2787), .IN2(n18805), .Q(g24263) );
  OR2X1 U19962 ( .IN1(n18806), .IN2(n18807), .Q(n18805) );
  INVX0 U19963 ( .INP(n18808), .ZN(n18807) );
  OR2X1 U19964 ( .IN1(n10740), .IN2(n10493), .Q(n18808) );
  AND2X1 U19965 ( .IN1(n5299), .IN2(n10795), .Q(n18806) );
  AND2X1 U19966 ( .IN1(n10813), .IN2(n5963), .Q(n2787) );
  OR2X1 U19967 ( .IN1(n18809), .IN2(n18810), .Q(g24262) );
  OR2X1 U19968 ( .IN1(n18811), .IN2(n18812), .Q(n18810) );
  AND2X1 U19969 ( .IN1(n10898), .IN2(g1548), .Q(n18812) );
  AND2X1 U19970 ( .IN1(n18813), .IN2(n10795), .Q(n18811) );
  AND2X1 U19971 ( .IN1(n18814), .IN2(g1564), .Q(n18813) );
  INVX0 U19972 ( .INP(n18815), .ZN(n18809) );
  OR2X1 U19973 ( .IN1(n18814), .IN2(g1564), .Q(n18815) );
  OR2X1 U19974 ( .IN1(n18816), .IN2(n17868), .Q(g24261) );
  AND2X1 U19975 ( .IN1(n10898), .IN2(g1585), .Q(n18816) );
  XNOR2X1 U19976 ( .IN1(n10386), .IN2(n18817), .Q(g24260) );
  AND2X1 U19977 ( .IN1(n10813), .IN2(g1548), .Q(n18817) );
  OR2X1 U19978 ( .IN1(n18818), .IN2(n17868), .Q(g24259) );
  AND2X1 U19979 ( .IN1(n10898), .IN2(g1579), .Q(n18818) );
  OR2X1 U19980 ( .IN1(n18819), .IN2(n18820), .Q(g24258) );
  AND2X1 U19981 ( .IN1(n10898), .IN2(g1554), .Q(n18820) );
  AND2X1 U19982 ( .IN1(n10813), .IN2(g496), .Q(n18819) );
  XOR2X1 U19983 ( .IN1(n5616), .IN2(n18821), .Q(g24257) );
  OR2X1 U19984 ( .IN1(n18822), .IN2(n10877), .Q(n18821) );
  OR2X1 U19985 ( .IN1(n18823), .IN2(n18824), .Q(g24256) );
  AND2X1 U19986 ( .IN1(n18825), .IN2(n10795), .Q(n18824) );
  OR2X1 U19987 ( .IN1(n18826), .IN2(n18827), .Q(n18825) );
  AND2X1 U19988 ( .IN1(n18828), .IN2(n18822), .Q(n18827) );
  INVX0 U19989 ( .INP(n18829), .ZN(n18826) );
  OR2X1 U19990 ( .IN1(n18822), .IN2(n18828), .Q(n18829) );
  AND2X1 U19991 ( .IN1(n18830), .IN2(n10474), .Q(n18828) );
  AND2X1 U19992 ( .IN1(n10061), .IN2(n18410), .Q(n18830) );
  AND2X1 U19993 ( .IN1(n5401), .IN2(n18831), .Q(n18410) );
  AND2X1 U19994 ( .IN1(n5616), .IN2(n5302), .Q(n18831) );
  OR2X1 U19995 ( .IN1(n18832), .IN2(n18833), .Q(n18822) );
  OR2X1 U19996 ( .IN1(n4836), .IN2(n18417), .Q(n18833) );
  INVX0 U19997 ( .INP(n17859), .ZN(n18417) );
  INVX0 U19998 ( .INP(n18834), .ZN(n4836) );
  XNOR2X1 U19999 ( .IN1(n10550), .IN2(n10118), .Q(n18832) );
  AND2X1 U20000 ( .IN1(n10899), .IN2(g1339), .Q(n18823) );
  OR2X1 U20001 ( .IN1(n18835), .IN2(n18836), .Q(g24255) );
  OR2X1 U20002 ( .IN1(n18837), .IN2(n18838), .Q(n18836) );
  AND2X1 U20003 ( .IN1(n10899), .IN2(g1589), .Q(n18838) );
  AND2X1 U20004 ( .IN1(n18839), .IN2(n10795), .Q(n18837) );
  AND2X1 U20005 ( .IN1(n10516), .IN2(g10527), .Q(n18839) );
  INVX0 U20006 ( .INP(n18840), .ZN(n18835) );
  OR2X1 U20007 ( .IN1(n13799), .IN2(n10516), .Q(n18840) );
  AND2X1 U20008 ( .IN1(n18841), .IN2(n18842), .Q(g24254) );
  AND2X1 U20009 ( .IN1(n18843), .IN2(n10516), .Q(n18842) );
  AND2X1 U20010 ( .IN1(n18844), .IN2(n10795), .Q(n18843) );
  OR2X1 U20011 ( .IN1(n18383), .IN2(n18845), .Q(n18844) );
  OR2X1 U20012 ( .IN1(n5768), .IN2(n18846), .Q(n18845) );
  AND2X1 U20013 ( .IN1(n17859), .IN2(n18834), .Q(n18846) );
  AND2X1 U20014 ( .IN1(n5322), .IN2(n5466), .Q(n18834) );
  AND2X1 U20015 ( .IN1(n17510), .IN2(n17519), .Q(n17859) );
  XNOR2X1 U20016 ( .IN1(g1339), .IN2(n10550), .Q(n17519) );
  INVX0 U20017 ( .INP(n16011), .ZN(n17510) );
  AND2X1 U20018 ( .IN1(n10550), .IN2(n5616), .Q(n16011) );
  OR2X1 U20019 ( .IN1(n10385), .IN2(n18814), .Q(n18383) );
  OR2X1 U20020 ( .IN1(n10386), .IN2(n5546), .Q(n18814) );
  AND2X1 U20021 ( .IN1(n10130), .IN2(n10129), .Q(n18841) );
  OR2X1 U20022 ( .IN1(n18847), .IN2(n18848), .Q(g24253) );
  AND2X1 U20023 ( .IN1(n18849), .IN2(n10795), .Q(n18848) );
  OR2X1 U20024 ( .IN1(n18850), .IN2(n18851), .Q(n18849) );
  AND2X1 U20025 ( .IN1(n5302), .IN2(g1532), .Q(n18851) );
  AND2X1 U20026 ( .IN1(g7946), .IN2(g1521), .Q(n18850) );
  AND2X1 U20027 ( .IN1(n10899), .IN2(g1306), .Q(n18847) );
  OR2X1 U20028 ( .IN1(n18395), .IN2(n18852), .Q(g24252) );
  OR2X1 U20029 ( .IN1(n18853), .IN2(n18854), .Q(n18852) );
  AND2X1 U20030 ( .IN1(n18855), .IN2(n10795), .Q(n18854) );
  AND2X1 U20031 ( .IN1(n5302), .IN2(g1521), .Q(n18855) );
  AND2X1 U20032 ( .IN1(test_so49), .IN2(n10894), .Q(n18853) );
  AND2X1 U20033 ( .IN1(n10813), .IN2(n18856), .Q(n18395) );
  AND2X1 U20034 ( .IN1(g1339), .IN2(g7946), .Q(n18856) );
  OR2X1 U20035 ( .IN1(n18857), .IN2(n18858), .Q(g24251) );
  AND2X1 U20036 ( .IN1(test_so12), .IN2(n18859), .Q(n18858) );
  AND2X1 U20037 ( .IN1(n16665), .IN2(g1442), .Q(n18857) );
  OR2X1 U20038 ( .IN1(n18860), .IN2(n18861), .Q(g24250) );
  INVX0 U20039 ( .INP(n18862), .ZN(n18861) );
  OR2X1 U20040 ( .IN1(n16665), .IN2(n5850), .Q(n18862) );
  AND2X1 U20041 ( .IN1(test_so12), .IN2(n16665), .Q(n18860) );
  INVX0 U20042 ( .INP(n18859), .ZN(n16665) );
  OR2X1 U20043 ( .IN1(n18863), .IN2(n18864), .Q(g24249) );
  INVX0 U20044 ( .INP(n18865), .ZN(n18864) );
  OR2X1 U20045 ( .IN1(n18866), .IN2(n5850), .Q(n18865) );
  AND2X1 U20046 ( .IN1(n18867), .IN2(n18859), .Q(n18866) );
  OR2X1 U20047 ( .IN1(n10887), .IN2(n16668), .Q(n18859) );
  OR2X1 U20048 ( .IN1(n10887), .IN2(test_so12), .Q(n18867) );
  AND2X1 U20049 ( .IN1(n16690), .IN2(n16668), .Q(n18863) );
  AND2X1 U20050 ( .IN1(n5364), .IN2(n18868), .Q(n16668) );
  AND2X1 U20051 ( .IN1(n10568), .IN2(g13272), .Q(n18868) );
  AND2X1 U20052 ( .IN1(n10433), .IN2(n10795), .Q(n16690) );
  OR2X1 U20053 ( .IN1(n18869), .IN2(n18870), .Q(g24248) );
  OR2X1 U20054 ( .IN1(n18871), .IN2(n18872), .Q(n18870) );
  AND2X1 U20055 ( .IN1(n5401), .IN2(n10796), .Q(n18872) );
  AND2X1 U20056 ( .IN1(n17868), .IN2(g1395), .Q(n18871) );
  XNOR2X1 U20057 ( .IN1(n10500), .IN2(n18873), .Q(n18869) );
  AND2X1 U20058 ( .IN1(n5655), .IN2(n10796), .Q(n18873) );
  AND2X1 U20059 ( .IN1(n17868), .IN2(n10512), .Q(g24247) );
  INVX0 U20060 ( .INP(n13799), .ZN(n17868) );
  OR2X1 U20061 ( .IN1(n5655), .IN2(n10876), .Q(n13799) );
  OR2X1 U20062 ( .IN1(n18874), .IN2(n18875), .Q(g24246) );
  OR2X1 U20063 ( .IN1(n18876), .IN2(n18877), .Q(n18875) );
  AND2X1 U20064 ( .IN1(n10899), .IN2(g1205), .Q(n18877) );
  AND2X1 U20065 ( .IN1(n18878), .IN2(n10796), .Q(n18876) );
  AND2X1 U20066 ( .IN1(n18879), .IN2(g1221), .Q(n18878) );
  AND2X1 U20067 ( .IN1(n18880), .IN2(n10387), .Q(n18874) );
  OR2X1 U20068 ( .IN1(n18881), .IN2(n17924), .Q(g24245) );
  AND2X1 U20069 ( .IN1(n10899), .IN2(g30332), .Q(n18881) );
  XNOR2X1 U20070 ( .IN1(n10388), .IN2(n18882), .Q(g24244) );
  AND2X1 U20071 ( .IN1(n10813), .IN2(g1205), .Q(n18882) );
  OR2X1 U20072 ( .IN1(n18883), .IN2(n17924), .Q(g24243) );
  AND2X1 U20073 ( .IN1(n10899), .IN2(g1236), .Q(n18883) );
  OR2X1 U20074 ( .IN1(n18884), .IN2(n18885), .Q(g24242) );
  AND2X1 U20075 ( .IN1(test_so76), .IN2(n10895), .Q(n18885) );
  AND2X1 U20076 ( .IN1(n10814), .IN2(g29215), .Q(n18884) );
  XOR2X1 U20077 ( .IN1(n5622), .IN2(n18886), .Q(g24241) );
  OR2X1 U20078 ( .IN1(n18887), .IN2(n10876), .Q(n18886) );
  OR2X1 U20079 ( .IN1(n18888), .IN2(n18889), .Q(g24240) );
  AND2X1 U20080 ( .IN1(n18890), .IN2(n10796), .Q(n18889) );
  OR2X1 U20081 ( .IN1(n18891), .IN2(n18892), .Q(n18890) );
  AND2X1 U20082 ( .IN1(n18893), .IN2(n18887), .Q(n18892) );
  INVX0 U20083 ( .INP(n18894), .ZN(n18891) );
  OR2X1 U20084 ( .IN1(n18887), .IN2(n18893), .Q(n18894) );
  AND2X1 U20085 ( .IN1(n18895), .IN2(n10475), .Q(n18893) );
  AND2X1 U20086 ( .IN1(n10050), .IN2(n18469), .Q(n18895) );
  AND2X1 U20087 ( .IN1(n5392), .IN2(n18896), .Q(n18469) );
  AND2X1 U20088 ( .IN1(n5622), .IN2(n5304), .Q(n18896) );
  OR2X1 U20089 ( .IN1(n18479), .IN2(n18897), .Q(n18887) );
  OR2X1 U20090 ( .IN1(n4837), .IN2(n18898), .Q(n18897) );
  XNOR2X1 U20091 ( .IN1(n10117), .IN2(n5320), .Q(n18898) );
  INVX0 U20092 ( .INP(n17916), .ZN(n18479) );
  AND2X1 U20093 ( .IN1(n10900), .IN2(g996), .Q(n18888) );
  OR2X1 U20094 ( .IN1(n18899), .IN2(n18900), .Q(g24239) );
  OR2X1 U20095 ( .IN1(n18901), .IN2(n18902), .Q(n18900) );
  AND2X1 U20096 ( .IN1(n10900), .IN2(g1246), .Q(n18902) );
  AND2X1 U20097 ( .IN1(n18903), .IN2(n10796), .Q(n18901) );
  AND2X1 U20098 ( .IN1(n10515), .IN2(g10500), .Q(n18903) );
  INVX0 U20099 ( .INP(n18904), .ZN(n18899) );
  OR2X1 U20100 ( .IN1(n13818), .IN2(n10515), .Q(n18904) );
  AND2X1 U20101 ( .IN1(n18905), .IN2(n18906), .Q(g24238) );
  AND2X1 U20102 ( .IN1(n18907), .IN2(n18908), .Q(n18906) );
  OR2X1 U20103 ( .IN1(n10565), .IN2(n18909), .Q(n18908) );
  OR2X1 U20104 ( .IN1(n18910), .IN2(n18446), .Q(n18909) );
  INVX0 U20105 ( .INP(n18450), .ZN(n18446) );
  AND2X1 U20106 ( .IN1(g1221), .IN2(n18880), .Q(n18450) );
  INVX0 U20107 ( .INP(n18879), .ZN(n18880) );
  OR2X1 U20108 ( .IN1(n10388), .IN2(n5547), .Q(n18879) );
  AND2X1 U20109 ( .IN1(n17916), .IN2(n18911), .Q(n18910) );
  INVX0 U20110 ( .INP(n4837), .ZN(n18911) );
  OR2X1 U20111 ( .IN1(test_so20), .IN2(g1008), .Q(n4837) );
  AND2X1 U20112 ( .IN1(n17531), .IN2(n17539), .Q(n17916) );
  XOR2X1 U20113 ( .IN1(n10138), .IN2(n5320), .Q(n17539) );
  INVX0 U20114 ( .INP(n16052), .ZN(n17531) );
  AND2X1 U20115 ( .IN1(n5320), .IN2(n5622), .Q(n16052) );
  AND2X1 U20116 ( .IN1(n10814), .IN2(n10574), .Q(n18907) );
  AND2X1 U20117 ( .IN1(n10111), .IN2(n10515), .Q(n18905) );
  OR2X1 U20118 ( .IN1(n18912), .IN2(n18913), .Q(g24237) );
  AND2X1 U20119 ( .IN1(n18914), .IN2(n10796), .Q(n18913) );
  OR2X1 U20120 ( .IN1(n18915), .IN2(n18916), .Q(n18914) );
  AND2X1 U20121 ( .IN1(g1178), .IN2(g7916), .Q(n18916) );
  AND2X1 U20122 ( .IN1(n5304), .IN2(g1189), .Q(n18915) );
  AND2X1 U20123 ( .IN1(n10900), .IN2(g962), .Q(n18912) );
  OR2X1 U20124 ( .IN1(n18917), .IN2(n18918), .Q(g24236) );
  AND2X1 U20125 ( .IN1(n18919), .IN2(n10796), .Q(n18918) );
  OR2X1 U20126 ( .IN1(n18920), .IN2(n18921), .Q(n18919) );
  AND2X1 U20127 ( .IN1(n5304), .IN2(g1178), .Q(n18921) );
  AND2X1 U20128 ( .IN1(g996), .IN2(g7916), .Q(n18920) );
  AND2X1 U20129 ( .IN1(n10900), .IN2(g1183), .Q(n18917) );
  OR2X1 U20130 ( .IN1(n18922), .IN2(n18923), .Q(g24235) );
  AND2X1 U20131 ( .IN1(n18924), .IN2(g1152), .Q(n18923) );
  AND2X1 U20132 ( .IN1(n16715), .IN2(test_so7), .Q(n18922) );
  OR2X1 U20133 ( .IN1(n18925), .IN2(n18926), .Q(g24234) );
  AND2X1 U20134 ( .IN1(n18924), .IN2(g1146), .Q(n18926) );
  AND2X1 U20135 ( .IN1(n16715), .IN2(g1152), .Q(n18925) );
  OR2X1 U20136 ( .IN1(n18927), .IN2(n18928), .Q(g24233) );
  AND2X1 U20137 ( .IN1(n18929), .IN2(g1146), .Q(n18928) );
  OR2X1 U20138 ( .IN1(n18930), .IN2(n16715), .Q(n18929) );
  INVX0 U20139 ( .INP(n18924), .ZN(n16715) );
  OR2X1 U20140 ( .IN1(n10886), .IN2(n16718), .Q(n18924) );
  AND2X1 U20141 ( .IN1(n5618), .IN2(n10796), .Q(n18930) );
  AND2X1 U20142 ( .IN1(n16739), .IN2(n16718), .Q(n18927) );
  AND2X1 U20143 ( .IN1(n5599), .IN2(n18931), .Q(n16718) );
  AND2X1 U20144 ( .IN1(g13259), .IN2(n5363), .Q(n18931) );
  AND2X1 U20145 ( .IN1(n10814), .IN2(n10583), .Q(n16739) );
  OR2X1 U20146 ( .IN1(n18932), .IN2(n18933), .Q(g24232) );
  OR2X1 U20147 ( .IN1(n18934), .IN2(n18935), .Q(n18933) );
  AND2X1 U20148 ( .IN1(n5392), .IN2(n10796), .Q(n18935) );
  AND2X1 U20149 ( .IN1(n17924), .IN2(g1052), .Q(n18934) );
  XNOR2X1 U20150 ( .IN1(n10499), .IN2(n18936), .Q(n18932) );
  AND2X1 U20151 ( .IN1(n5654), .IN2(n10797), .Q(n18936) );
  AND2X1 U20152 ( .IN1(n17924), .IN2(n10513), .Q(g24231) );
  INVX0 U20153 ( .INP(n13818), .ZN(n17924) );
  OR2X1 U20154 ( .IN1(n5654), .IN2(n10876), .Q(n13818) );
  OR2X1 U20155 ( .IN1(n18937), .IN2(n18938), .Q(g24216) );
  AND2X1 U20156 ( .IN1(n18939), .IN2(g854), .Q(n18938) );
  AND2X1 U20157 ( .IN1(n16813), .IN2(g847), .Q(n18937) );
  OR2X1 U20158 ( .IN1(n18940), .IN2(n18941), .Q(g24215) );
  AND2X1 U20159 ( .IN1(n18942), .IN2(g703), .Q(n18941) );
  OR2X1 U20160 ( .IN1(n10888), .IN2(n18943), .Q(n18942) );
  AND2X1 U20161 ( .IN1(n5562), .IN2(n17977), .Q(n18943) );
  AND2X1 U20162 ( .IN1(g847), .IN2(n4948), .Q(n17977) );
  AND2X1 U20163 ( .IN1(n18944), .IN2(g837), .Q(n18940) );
  OR2X1 U20164 ( .IN1(n18945), .IN2(n16813), .Q(n18944) );
  AND2X1 U20165 ( .IN1(n18946), .IN2(n18947), .Q(n18945) );
  OR2X1 U20166 ( .IN1(n10419), .IN2(n5728), .Q(n18947) );
  AND2X1 U20167 ( .IN1(n18948), .IN2(n10797), .Q(n18946) );
  OR2X1 U20168 ( .IN1(n18949), .IN2(n18950), .Q(g24214) );
  OR2X1 U20169 ( .IN1(n18951), .IN2(n18952), .Q(n18950) );
  AND2X1 U20170 ( .IN1(n18953), .IN2(n5709), .Q(n18952) );
  AND2X1 U20171 ( .IN1(n18954), .IN2(n18955), .Q(n18953) );
  AND2X1 U20172 ( .IN1(g817), .IN2(g723), .Q(n18955) );
  AND2X1 U20173 ( .IN1(n16800), .IN2(g822), .Q(n18954) );
  AND2X1 U20174 ( .IN1(n10900), .IN2(g847), .Q(n18951) );
  AND2X1 U20175 ( .IN1(n18956), .IN2(g703), .Q(n18949) );
  OR2X1 U20176 ( .IN1(n18957), .IN2(n16813), .Q(n18956) );
  AND2X1 U20177 ( .IN1(n18958), .IN2(n10797), .Q(n18957) );
  OR2X1 U20178 ( .IN1(n5562), .IN2(n18948), .Q(n18958) );
  OR2X1 U20179 ( .IN1(n5709), .IN2(n5733), .Q(n18948) );
  OR2X1 U20180 ( .IN1(n18959), .IN2(g24212), .Q(g24213) );
  AND2X1 U20181 ( .IN1(n10900), .IN2(g753), .Q(n18959) );
  OR2X1 U20182 ( .IN1(n18960), .IN2(n18961), .Q(g24211) );
  AND2X1 U20183 ( .IN1(n10900), .IN2(g546), .Q(n18961) );
  AND2X1 U20184 ( .IN1(n2404), .IN2(n18962), .Q(n18960) );
  OR2X1 U20185 ( .IN1(n5520), .IN2(test_so41), .Q(n18962) );
  AND2X1 U20186 ( .IN1(n18963), .IN2(n14600), .Q(g24210) );
  AND2X1 U20187 ( .IN1(n5548), .IN2(n18964), .Q(n14600) );
  INVX0 U20188 ( .INP(n18965), .ZN(n18964) );
  OR2X1 U20189 ( .IN1(n5287), .IN2(n10136), .Q(n18965) );
  AND2X1 U20190 ( .IN1(n18966), .IN2(n10797), .Q(n18963) );
  OR2X1 U20191 ( .IN1(n18967), .IN2(n18968), .Q(n18966) );
  AND2X1 U20192 ( .IN1(g174), .IN2(g168), .Q(n18968) );
  AND2X1 U20193 ( .IN1(test_so72), .IN2(n16080), .Q(n18967) );
  OR2X1 U20194 ( .IN1(g174), .IN2(g168), .Q(n16080) );
  OR2X1 U20195 ( .IN1(n18969), .IN2(n18970), .Q(g24209) );
  AND2X1 U20196 ( .IN1(n16800), .IN2(g446), .Q(n18970) );
  AND2X1 U20197 ( .IN1(n16813), .IN2(g417), .Q(n18969) );
  OR2X1 U20198 ( .IN1(n18971), .IN2(n18972), .Q(g24208) );
  OR2X1 U20199 ( .IN1(n18973), .IN2(n18974), .Q(n18972) );
  AND2X1 U20200 ( .IN1(n16800), .IN2(g246), .Q(n18974) );
  AND2X1 U20201 ( .IN1(n16813), .IN2(g475), .Q(n18973) );
  AND2X1 U20202 ( .IN1(n10900), .IN2(g424), .Q(n18971) );
  OR2X1 U20203 ( .IN1(n18975), .IN2(n18976), .Q(g24207) );
  AND2X1 U20204 ( .IN1(n18939), .IN2(g475), .Q(n18976) );
  AND2X1 U20205 ( .IN1(n16813), .IN2(g441), .Q(n18975) );
  OR2X1 U20206 ( .IN1(n18977), .IN2(n18978), .Q(g24206) );
  AND2X1 U20207 ( .IN1(n18939), .IN2(g441), .Q(n18978) );
  AND2X1 U20208 ( .IN1(n16813), .IN2(g437), .Q(n18977) );
  OR2X1 U20209 ( .IN1(n18979), .IN2(n18980), .Q(g24205) );
  OR2X1 U20210 ( .IN1(n18981), .IN2(n18982), .Q(n18980) );
  AND2X1 U20211 ( .IN1(n16800), .IN2(g269), .Q(n18982) );
  AND2X1 U20212 ( .IN1(test_so23), .IN2(n16813), .Q(n18981) );
  AND2X1 U20213 ( .IN1(n10900), .IN2(g437), .Q(n18979) );
  OR2X1 U20214 ( .IN1(n18983), .IN2(n18984), .Q(g24204) );
  AND2X1 U20215 ( .IN1(test_so23), .IN2(n18939), .Q(n18984) );
  AND2X1 U20216 ( .IN1(n16813), .IN2(g429), .Q(n18983) );
  OR2X1 U20217 ( .IN1(n18985), .IN2(n18986), .Q(g24203) );
  AND2X1 U20218 ( .IN1(n18939), .IN2(g429), .Q(n18986) );
  AND2X1 U20219 ( .IN1(n16813), .IN2(g401), .Q(n18985) );
  OR2X1 U20220 ( .IN1(n18987), .IN2(n18988), .Q(g24202) );
  AND2X1 U20221 ( .IN1(n18939), .IN2(g411), .Q(n18988) );
  AND2X1 U20222 ( .IN1(n16813), .IN2(g424), .Q(n18987) );
  OR2X1 U20223 ( .IN1(n18989), .IN2(n18990), .Q(g24201) );
  AND2X1 U20224 ( .IN1(n18939), .IN2(g392), .Q(n18990) );
  INVX0 U20225 ( .INP(n16813), .ZN(n18939) );
  AND2X1 U20226 ( .IN1(n16813), .IN2(g405), .Q(n18989) );
  OR2X1 U20227 ( .IN1(n18991), .IN2(n18992), .Q(g24200) );
  OR2X1 U20228 ( .IN1(n18993), .IN2(n18994), .Q(n18992) );
  AND2X1 U20229 ( .IN1(n16813), .IN2(g392), .Q(n18994) );
  AND2X1 U20230 ( .IN1(n17994), .IN2(n10797), .Q(n16813) );
  INVX0 U20231 ( .INP(n4948), .ZN(n17994) );
  AND2X1 U20232 ( .IN1(n18995), .IN2(n16800), .Q(n18993) );
  AND2X1 U20233 ( .IN1(n10814), .IN2(n4948), .Q(n16800) );
  AND2X1 U20234 ( .IN1(n5821), .IN2(g854), .Q(n18995) );
  AND2X1 U20235 ( .IN1(n10901), .IN2(g401), .Q(n18991) );
  AND2X1 U20236 ( .IN1(n10527), .IN2(n10473), .Q(g23190) );
  OR2X1 U20237 ( .IN1(n18996), .IN2(n18997), .Q(g21901) );
  AND2X1 U20238 ( .IN1(n18998), .IN2(n10797), .Q(n18997) );
  OR2X1 U20239 ( .IN1(n18999), .IN2(n19000), .Q(n18998) );
  AND2X1 U20240 ( .IN1(n5380), .IN2(n19001), .Q(n19000) );
  OR2X1 U20241 ( .IN1(n19002), .IN2(g8786), .Q(n19001) );
  AND2X1 U20242 ( .IN1(n19003), .IN2(n19004), .Q(n19002) );
  AND2X1 U20243 ( .IN1(n19005), .IN2(n19006), .Q(n19004) );
  AND2X1 U20244 ( .IN1(n10141), .IN2(DFF_1234_n1), .Q(n19006) );
  AND2X1 U20245 ( .IN1(DFF_480_n1), .IN2(DFF_909_n1), .Q(n19005) );
  AND2X1 U20246 ( .IN1(n19007), .IN2(n10144), .Q(n19003) );
  AND2X1 U20247 ( .IN1(n10143), .IN2(n10142), .Q(n19007) );
  AND2X1 U20248 ( .IN1(n5694), .IN2(g4180), .Q(n18999) );
  AND2X1 U20249 ( .IN1(n10901), .IN2(g2946), .Q(n18996) );
  OR2X1 U20250 ( .IN1(n19008), .IN2(n19009), .Q(g21900) );
  AND2X1 U20251 ( .IN1(n19010), .IN2(n10797), .Q(n19009) );
  AND2X1 U20252 ( .IN1(n10492), .IN2(n10491), .Q(n19010) );
  INVX0 U20253 ( .INP(n19011), .ZN(n19008) );
  OR2X1 U20254 ( .IN1(n10738), .IN2(n10104), .Q(n19011) );
  XNOR2X1 U20255 ( .IN1(n10416), .IN2(n19012), .Q(g21899) );
  AND2X1 U20256 ( .IN1(n10814), .IN2(g9019), .Q(n19012) );
  OR2X1 U20257 ( .IN1(n19013), .IN2(n19014), .Q(g21898) );
  AND2X1 U20258 ( .IN1(n10901), .IN2(g4284), .Q(n19014) );
  AND2X1 U20259 ( .IN1(n10416), .IN2(n10797), .Q(n19013) );
  XNOR2X1 U20260 ( .IN1(n10417), .IN2(n19015), .Q(g21897) );
  AND2X1 U20261 ( .IN1(n10815), .IN2(g8839), .Q(n19015) );
  OR2X1 U20262 ( .IN1(n19016), .IN2(n19017), .Q(g21896) );
  AND2X1 U20263 ( .IN1(n10901), .IN2(g4245), .Q(n19017) );
  AND2X1 U20264 ( .IN1(n10417), .IN2(n10797), .Q(n19016) );
  OR2X1 U20265 ( .IN1(n19018), .IN2(n19019), .Q(g21895) );
  AND2X1 U20266 ( .IN1(n18732), .IN2(g4269), .Q(n19019) );
  OR2X1 U20267 ( .IN1(n19020), .IN2(g21893), .Q(n18732) );
  AND2X1 U20268 ( .IN1(n5823), .IN2(n10798), .Q(n19020) );
  AND2X1 U20269 ( .IN1(n19021), .IN2(g4264), .Q(n19018) );
  OR2X1 U20270 ( .IN1(n10886), .IN2(n19022), .Q(n19021) );
  AND2X1 U20271 ( .IN1(n5763), .IN2(g4258), .Q(n19022) );
  OR2X1 U20272 ( .IN1(n19023), .IN2(n19024), .Q(g21894) );
  AND2X1 U20273 ( .IN1(g21893), .IN2(g4264), .Q(n19024) );
  AND2X1 U20274 ( .IN1(n19025), .IN2(g4258), .Q(n19023) );
  OR2X1 U20275 ( .IN1(n5823), .IN2(n10875), .Q(n19025) );
  AND2X1 U20276 ( .IN1(n10815), .IN2(n10501), .Q(g21893) );
  OR2X1 U20277 ( .IN1(n19026), .IN2(n19027), .Q(g21892) );
  AND2X1 U20278 ( .IN1(n10901), .IN2(g4273), .Q(n19027) );
  AND2X1 U20279 ( .IN1(n10104), .IN2(n10793), .Q(n19026) );
  OR2X1 U20280 ( .IN1(n19028), .IN2(n19029), .Q(g21891) );
  AND2X1 U20281 ( .IN1(n18739), .IN2(n10750), .Q(n19029) );
  OR2X1 U20282 ( .IN1(n19030), .IN2(n19031), .Q(n18739) );
  AND2X1 U20283 ( .IN1(n5484), .IN2(n10391), .Q(n19031) );
  AND2X1 U20284 ( .IN1(n10392), .IN2(g4253), .Q(n19030) );
  AND2X1 U20285 ( .IN1(n10901), .IN2(g4180), .Q(n19028) );
  AND2X1 U20286 ( .IN1(n10901), .IN2(n9240), .Q(g21727) );
  AND2X1 U20287 ( .IN1(n10910), .IN2(g2975), .Q(g18597) );
  INVX0 U20288 ( .INP(g5), .ZN(g12833) );
  OR2X1 U5116_U1 ( .IN1(g34783), .IN2(n286), .Q(g34221) );
  OR2X1 U5126_U1 ( .IN1(n4836), .IN2(n4896), .Q(n4895) );
  OR2X1 U5127_U1 ( .IN1(n4837), .IN2(n4921), .Q(n4920) );
  OR2X1 U5128_U1 ( .IN1(n2787), .IN2(n4411), .Q(n5045) );
  OR2X1 U5129_U1 ( .IN1(g559), .IN2(g9048), .Q(n4959) );
  INVX0 U5353_U2 ( .INP(n10540), .ZN(U5353_n1) );
  AND2X1 U5353_U1 ( .IN1(n5960), .IN2(U5353_n1), .Q(n4689) );
  INVX0 U5355_U2 ( .INP(n10535), .ZN(U5355_n1) );
  AND2X1 U5355_U1 ( .IN1(n5961), .IN2(U5355_n1), .Q(n4708) );
  INVX0 U5961_U2 ( .INP(n725), .ZN(U5961_n1) );
  AND2X1 U5961_U1 ( .IN1(n3593), .IN2(U5961_n1), .Q(n3595) );
  INVX0 U5962_U2 ( .INP(n1287), .ZN(U5962_n1) );
  AND2X1 U5962_U1 ( .IN1(n3574), .IN2(U5962_n1), .Q(n3576) );
  INVX0 U5963_U2 ( .INP(n1285), .ZN(U5963_n1) );
  AND2X1 U5963_U1 ( .IN1(n3517), .IN2(U5963_n1), .Q(n3519) );
  INVX0 U5964_U2 ( .INP(n1643), .ZN(U5964_n1) );
  AND2X1 U5964_U1 ( .IN1(n3628), .IN2(U5964_n1), .Q(n3630) );
  INVX0 U5965_U2 ( .INP(n1289), .ZN(U5965_n1) );
  AND2X1 U5965_U1 ( .IN1(n3555), .IN2(U5965_n1), .Q(n3557) );
  INVX0 U5966_U2 ( .INP(n736), .ZN(U5966_n1) );
  AND2X1 U5966_U1 ( .IN1(n3646), .IN2(U5966_n1), .Q(n3648) );
  INVX0 U5967_U2 ( .INP(n1282), .ZN(U5967_n1) );
  AND2X1 U5967_U1 ( .IN1(n3536), .IN2(U5967_n1), .Q(n3538) );
  INVX0 U5968_U2 ( .INP(n727), .ZN(U5968_n1) );
  AND2X1 U5968_U1 ( .IN1(n3611), .IN2(U5968_n1), .Q(n3613) );
  AND2X1 U6100_U2 ( .IN1(n3635), .IN2(U6100_n1), .Q(n4888) );
  INVX0 U6100_U1 ( .INP(n10892), .ZN(U6100_n1) );
  INVX0 U6211_U2 ( .INP(n1645), .ZN(U6211_n1) );
  AND2X1 U6211_U1 ( .IN1(n3623), .IN2(U6211_n1), .Q(n3622) );
  INVX0 U6212_U2 ( .INP(n3588), .ZN(U6212_n1) );
  AND2X1 U6212_U1 ( .IN1(n3587), .IN2(U6212_n1), .Q(n3586) );
  INVX0 U6213_U2 ( .INP(n3606), .ZN(U6213_n1) );
  AND2X1 U6213_U1 ( .IN1(n3605), .IN2(U6213_n1), .Q(n3604) );
  INVX0 U6214_U2 ( .INP(n3569), .ZN(U6214_n1) );
  AND2X1 U6214_U1 ( .IN1(n3568), .IN2(U6214_n1), .Q(n3567) );
  INVX0 U6215_U2 ( .INP(n3550), .ZN(U6215_n1) );
  AND2X1 U6215_U1 ( .IN1(n3549), .IN2(U6215_n1), .Q(n3548) );
  INVX0 U6216_U2 ( .INP(n3006), .ZN(U6216_n1) );
  AND2X1 U6216_U1 ( .IN1(n3512), .IN2(U6216_n1), .Q(n3511) );
  INVX0 U6217_U2 ( .INP(n3007), .ZN(U6217_n1) );
  AND2X1 U6217_U1 ( .IN1(n3531), .IN2(U6217_n1), .Q(n3530) );
  INVX0 U6218_U2 ( .INP(n3003), .ZN(U6218_n1) );
  AND2X1 U6218_U1 ( .IN1(n3641), .IN2(U6218_n1), .Q(n3640) );
  INVX0 U6279_U2 ( .INP(n5337), .ZN(U6279_n1) );
  AND2X1 U6279_U1 ( .IN1(n4537), .IN2(U6279_n1), .Q(n4201) );
  INVX0 U6280_U2 ( .INP(n5336), .ZN(U6280_n1) );
  AND2X1 U6280_U1 ( .IN1(n4201), .IN2(U6280_n1), .Q(n3745) );
  INVX0 U6281_U2 ( .INP(n5294), .ZN(U6281_n1) );
  AND2X1 U6281_U1 ( .IN1(n3745), .IN2(U6281_n1), .Q(n3684) );
  INVX0 U6282_U2 ( .INP(n5552), .ZN(U6282_n1) );
  AND2X1 U6282_U1 ( .IN1(n3684), .IN2(U6282_n1), .Q(n3274) );
  INVX0 U6283_U2 ( .INP(n5472), .ZN(U6283_n1) );
  AND2X1 U6283_U1 ( .IN1(n3274), .IN2(U6283_n1), .Q(n2982) );
  INVX0 U6284_U2 ( .INP(n5476), .ZN(U6284_n1) );
  AND2X1 U6284_U1 ( .IN1(n2982), .IN2(U6284_n1), .Q(n2706) );
  INVX0 U6285_U2 ( .INP(n5550), .ZN(U6285_n1) );
  AND2X1 U6285_U1 ( .IN1(n2706), .IN2(U6285_n1), .Q(n2649) );
  INVX0 U6286_U2 ( .INP(n5473), .ZN(U6286_n1) );
  AND2X1 U6286_U1 ( .IN1(n2649), .IN2(U6286_n1), .Q(n2556) );
  INVX0 U6287_U2 ( .INP(n5475), .ZN(U6287_n1) );
  AND2X1 U6287_U1 ( .IN1(n2556), .IN2(U6287_n1), .Q(n2509) );
  INVX0 U6288_U2 ( .INP(n5474), .ZN(U6288_n1) );
  AND2X1 U6288_U1 ( .IN1(n2509), .IN2(U6288_n1), .Q(n2487) );
  INVX0 U6289_U2 ( .INP(n5339), .ZN(U6289_n1) );
  AND2X1 U6289_U1 ( .IN1(n2487), .IN2(U6289_n1), .Q(n2427) );
  INVX0 U6290_U2 ( .INP(n5672), .ZN(U6290_n1) );
  AND2X1 U6290_U1 ( .IN1(n2427), .IN2(U6290_n1), .Q(n2423) );
  INVX0 U6291_U2 ( .INP(n5335), .ZN(U6291_n1) );
  AND2X1 U6291_U1 ( .IN1(n4826), .IN2(U6291_n1), .Q(n4537) );
  AND2X1 U6292_U2 ( .IN1(n4959), .IN2(U6292_n1), .Q(n2421) );
  INVX0 U6292_U1 ( .INP(n10892), .ZN(U6292_n1) );
  AND2X1 U6338_U2 ( .IN1(n4210), .IN2(U6338_n1), .Q(n3765) );
  INVX0 U6338_U1 ( .INP(n10893), .ZN(U6338_n1) );
  INVX0 U6341_U2 ( .INP(n1075), .ZN(U6341_n1) );
  AND2X1 U6341_U1 ( .IN1(n3765), .IN2(U6341_n1), .Q(n3951) );
  INVX0 U6342_U2 ( .INP(n3404), .ZN(U6342_n1) );
  AND2X1 U6342_U1 ( .IN1(n3765), .IN2(U6342_n1), .Q(n3774) );
  INVX0 U6343_U2 ( .INP(n3424), .ZN(U6343_n1) );
  AND2X1 U6343_U1 ( .IN1(n3765), .IN2(U6343_n1), .Q(n3842) );
  INVX0 U6344_U2 ( .INP(n3414), .ZN(U6344_n1) );
  AND2X1 U6344_U1 ( .IN1(n3765), .IN2(U6344_n1), .Q(n3808) );
  INVX0 U6345_U2 ( .INP(n3444), .ZN(U6345_n1) );
  AND2X1 U6345_U1 ( .IN1(n3765), .IN2(U6345_n1), .Q(n3908) );
  INVX0 U6346_U2 ( .INP(n3489), .ZN(U6346_n1) );
  AND2X1 U6346_U1 ( .IN1(n3765), .IN2(U6346_n1), .Q(n3984) );
  INVX0 U6347_U2 ( .INP(n3434), .ZN(U6347_n1) );
  AND2X1 U6347_U1 ( .IN1(n3765), .IN2(U6347_n1), .Q(n3875) );
  INVX0 U6348_U2 ( .INP(n3500), .ZN(U6348_n1) );
  AND2X1 U6348_U1 ( .IN1(n3765), .IN2(U6348_n1), .Q(n4015) );
  INVX0 U6349_U2 ( .INP(n3446), .ZN(U6349_n1) );
  AND2X1 U6349_U1 ( .IN1(n3765), .IN2(U6349_n1), .Q(n3914) );
  INVX0 U6350_U2 ( .INP(n3406), .ZN(U6350_n1) );
  AND2X1 U6350_U1 ( .IN1(n3765), .IN2(U6350_n1), .Q(n3780) );
  INVX0 U6351_U2 ( .INP(n3481), .ZN(U6351_n1) );
  AND2X1 U6351_U1 ( .IN1(n3765), .IN2(U6351_n1), .Q(n3957) );
  INVX0 U6352_U2 ( .INP(n3426), .ZN(U6352_n1) );
  AND2X1 U6352_U1 ( .IN1(n3765), .IN2(U6352_n1), .Q(n3848) );
  INVX0 U6353_U2 ( .INP(n3491), .ZN(U6353_n1) );
  AND2X1 U6353_U1 ( .IN1(n3765), .IN2(U6353_n1), .Q(n3990) );
  INVX0 U6354_U2 ( .INP(n3416), .ZN(U6354_n1) );
  AND2X1 U6354_U1 ( .IN1(n3765), .IN2(U6354_n1), .Q(n3814) );
  INVX0 U6355_U2 ( .INP(n3436), .ZN(U6355_n1) );
  AND2X1 U6355_U1 ( .IN1(n3765), .IN2(U6355_n1), .Q(n3881) );
  INVX0 U6356_U2 ( .INP(n3502), .ZN(U6356_n1) );
  AND2X1 U6356_U1 ( .IN1(n3765), .IN2(U6356_n1), .Q(n4022) );
  INVX0 U6357_U2 ( .INP(n3501), .ZN(U6357_n1) );
  AND2X1 U6357_U1 ( .IN1(n3765), .IN2(U6357_n1), .Q(n4027) );
  INVX0 U6358_U2 ( .INP(n3407), .ZN(U6358_n1) );
  AND2X1 U6358_U1 ( .IN1(n3765), .IN2(U6358_n1), .Q(n3785) );
  INVX0 U6359_U2 ( .INP(n3482), .ZN(U6359_n1) );
  AND2X1 U6359_U1 ( .IN1(n3765), .IN2(U6359_n1), .Q(n3962) );
  INVX0 U6360_U2 ( .INP(n3427), .ZN(U6360_n1) );
  AND2X1 U6360_U1 ( .IN1(n3765), .IN2(U6360_n1), .Q(n3853) );
  INVX0 U6361_U2 ( .INP(n3437), .ZN(U6361_n1) );
  AND2X1 U6361_U1 ( .IN1(n3765), .IN2(U6361_n1), .Q(n3886) );
  INVX0 U6362_U2 ( .INP(n3417), .ZN(U6362_n1) );
  AND2X1 U6362_U1 ( .IN1(n3765), .IN2(U6362_n1), .Q(n3819) );
  INVX0 U6363_U2 ( .INP(n3492), .ZN(U6363_n1) );
  AND2X1 U6363_U1 ( .IN1(n3765), .IN2(U6363_n1), .Q(n3995) );
  INVX0 U6364_U2 ( .INP(n3447), .ZN(U6364_n1) );
  AND2X1 U6364_U1 ( .IN1(n3765), .IN2(U6364_n1), .Q(n3919) );
  INVX0 U6365_U2 ( .INP(n5471), .ZN(U6365_n1) );
  AND2X1 U6365_U1 ( .IN1(n3682), .IN2(U6365_n1), .Q(n3272) );
  INVX0 U6366_U2 ( .INP(n5331), .ZN(U6366_n1) );
  AND2X1 U6366_U1 ( .IN1(n3272), .IN2(U6366_n1), .Q(n2980) );
  INVX0 U6367_U2 ( .INP(n5332), .ZN(U6367_n1) );
  AND2X1 U6367_U1 ( .IN1(n2980), .IN2(U6367_n1), .Q(n2704) );
  INVX0 U6368_U2 ( .INP(n5333), .ZN(U6368_n1) );
  AND2X1 U6368_U1 ( .IN1(n2704), .IN2(U6368_n1), .Q(n2647) );
  INVX0 U6369_U2 ( .INP(n5334), .ZN(U6369_n1) );
  AND2X1 U6369_U1 ( .IN1(n2647), .IN2(U6369_n1), .Q(n2554) );
  INVX0 U6370_U2 ( .INP(n5330), .ZN(U6370_n1) );
  AND2X1 U6370_U1 ( .IN1(n2554), .IN2(U6370_n1), .Q(n2507) );
  INVX0 U6371_U2 ( .INP(n5551), .ZN(U6371_n1) );
  AND2X1 U6371_U1 ( .IN1(n2507), .IN2(U6371_n1), .Q(n2485) );
  INVX0 U6372_U2 ( .INP(n5293), .ZN(U6372_n1) );
  AND2X1 U6372_U1 ( .IN1(n2485), .IN2(U6372_n1), .Q(n2425) );
  INVX0 U6373_U2 ( .INP(n5292), .ZN(U6373_n1) );
  AND2X1 U6373_U1 ( .IN1(n2425), .IN2(U6373_n1), .Q(n2419) );
  INVX0 U6374_U2 ( .INP(n5470), .ZN(U6374_n1) );
  AND2X1 U6374_U1 ( .IN1(n53), .IN2(U6374_n1), .Q(n3682) );
  INVX0 U6375_U2 ( .INP(n5291), .ZN(U6375_n1) );
  AND2X1 U6375_U1 ( .IN1(n2419), .IN2(U6375_n1), .Q(n2405) );
  AND2X1 U6417_U2 ( .IN1(n4198), .IN2(U6417_n1), .Q(n2404) );
  INVX0 U6417_U1 ( .INP(n10892), .ZN(U6417_n1) );
  INVX0 U6446_U2 ( .INP(n1698), .ZN(U6446_n1) );
  AND2X1 U6446_U1 ( .IN1(g110), .IN2(U6446_n1), .Q(n3524) );
  INVX0 U6465_U2 ( .INP(n5600), .ZN(U6465_n1) );
  AND2X1 U6465_U1 ( .IN1(n735), .IN2(U6465_n1), .Q(n4388) );
  INVX0 U6497_U2 ( .INP(n3635), .ZN(U6497_n1) );
  AND2X1 U6497_U1 ( .IN1(n760), .IN2(U6497_n1), .Q(n3005) );
  AND2X1 U6523_U2 ( .IN1(n4946), .IN2(U6523_n1), .Q(n4945) );
  INVX0 U6523_U1 ( .INP(n10892), .ZN(U6523_n1) );
  INVX0 U6542_U2 ( .INP(n5300), .ZN(U6542_n1) );
  AND2X1 U6542_U1 ( .IN1(n760), .IN2(U6542_n1), .Q(n3525) );
  INVX0 U6552_U2 ( .INP(n5676), .ZN(U6552_n1) );
  AND2X1 U6552_U1 ( .IN1(n3281), .IN2(U6552_n1), .Q(n3277) );
  INVX0 U6553_U2 ( .INP(n5680), .ZN(U6553_n1) );
  AND2X1 U6553_U1 ( .IN1(n3276), .IN2(U6553_n1), .Q(n2989) );
  INVX0 U6554_U2 ( .INP(n5677), .ZN(U6554_n1) );
  AND2X1 U6554_U1 ( .IN1(n3277), .IN2(U6554_n1), .Q(n2991) );
  INVX0 U6555_U2 ( .INP(n5561), .ZN(U6555_n1) );
  AND2X1 U6555_U1 ( .IN1(n3687), .IN2(U6555_n1), .Q(n3281) );
  INVX0 U6556_U2 ( .INP(n5679), .ZN(U6556_n1) );
  AND2X1 U6556_U1 ( .IN1(n44), .IN2(U6556_n1), .Q(n3276) );
  INVX0 U6559_U2 ( .INP(n5678), .ZN(U6559_n1) );
  AND2X1 U6559_U1 ( .IN1(n2991), .IN2(U6559_n1), .Q(n2710) );
  INVX0 U6560_U2 ( .INP(n5675), .ZN(U6560_n1) );
  AND2X1 U6560_U1 ( .IN1(n2989), .IN2(U6560_n1), .Q(n2707) );
  INVX0 U6561_U2 ( .INP(n5327), .ZN(U6561_n1) );
  AND2X1 U6561_U1 ( .IN1(n3174), .IN2(U6561_n1), .Q(n3116) );
  INVX0 U6570_U2 ( .INP(n5477), .ZN(U6570_n1) );
  AND2X1 U6570_U1 ( .IN1(n3362), .IN2(U6570_n1), .Q(n2527) );
  INVX0 U6911_U2 ( .INP(n2726), .ZN(U6911_n1) );
  AND2X1 U6911_U1 ( .IN1(n3115), .IN2(U6911_n1), .Q(n3111) );
  INVX0 U6912_U2 ( .INP(n2727), .ZN(U6912_n1) );
  AND2X1 U6912_U1 ( .IN1(n3115), .IN2(U6912_n1), .Q(n3131) );
  INVX0 U6917_U2 ( .INP(n5350), .ZN(U6917_n1) );
  AND2X1 U6917_U1 ( .IN1(n3933), .IN2(U6917_n1), .Q(n3799) );
  INVX0 U6926_U2 ( .INP(n5674), .ZN(U6926_n1) );
  AND2X1 U6926_U1 ( .IN1(n3664), .IN2(U6926_n1), .Q(n3662) );
  INVX0 U6927_U2 ( .INP(n5673), .ZN(U6927_n1) );
  AND2X1 U6927_U1 ( .IN1(n3673), .IN2(U6927_n1), .Q(n3671) );
  INVX0 U6929_U2 ( .INP(n3506), .ZN(U6929_n1) );
  AND2X1 U6929_U1 ( .IN1(n1284), .IN2(U6929_n1), .Q(n2790) );
  INVX0 U6931_U2 ( .INP(n5554), .ZN(U6931_n1) );
  AND2X1 U6931_U1 ( .IN1(n4490), .IN2(U6931_n1), .Q(n4178) );
  INVX0 U6932_U2 ( .INP(n5555), .ZN(U6932_n1) );
  AND2X1 U6932_U1 ( .IN1(n4514), .IN2(U6932_n1), .Q(n4196) );
  INVX0 U6933_U2 ( .INP(n5558), .ZN(U6933_n1) );
  AND2X1 U6933_U1 ( .IN1(n4178), .IN2(U6933_n1), .Q(n3736) );
  INVX0 U6934_U2 ( .INP(n5559), .ZN(U6934_n1) );
  AND2X1 U6934_U1 ( .IN1(n4196), .IN2(U6934_n1), .Q(n3741) );
  INVX0 U6935_U2 ( .INP(n5553), .ZN(U6935_n1) );
  AND2X1 U6935_U1 ( .IN1(n3736), .IN2(U6935_n1), .Q(n3664) );
  INVX0 U6936_U2 ( .INP(n5560), .ZN(U6936_n1) );
  AND2X1 U6936_U1 ( .IN1(n3741), .IN2(U6936_n1), .Q(n3673) );
  INVX0 U6937_U2 ( .INP(n5303), .ZN(U6937_n1) );
  AND2X1 U6937_U1 ( .IN1(n108), .IN2(U6937_n1), .Q(n2598) );
  INVX0 U6938_U2 ( .INP(n5556), .ZN(U6938_n1) );
  AND2X1 U6938_U1 ( .IN1(n1156), .IN2(U6938_n1), .Q(n4490) );
  INVX0 U6939_U2 ( .INP(n5557), .ZN(U6939_n1) );
  AND2X1 U6939_U1 ( .IN1(n251), .IN2(U6939_n1), .Q(n4514) );
  INVX0 U6940_U2 ( .INP(n5422), .ZN(U6940_n1) );
  AND2X1 U6940_U1 ( .IN1(n4814), .IN2(U6940_n1), .Q(n4519) );
  INVX0 U6941_U2 ( .INP(n5323), .ZN(U6941_n1) );
  AND2X1 U6941_U1 ( .IN1(n2607), .IN2(U6941_n1), .Q(n2594) );
  INVX0 U6944_U2 ( .INP(n5348), .ZN(U6944_n1) );
  AND2X1 U6944_U1 ( .IN1(n3084), .IN2(U6944_n1), .Q(n3033) );
  INVX0 U6950_U2 ( .INP(n5365), .ZN(U6950_n1) );
  AND2X1 U6950_U1 ( .IN1(n2598), .IN2(U6950_n1), .Q(n2590) );
  INVX0 U6954_U2 ( .INP(n2727), .ZN(U6954_n1) );
  AND2X1 U6954_U1 ( .IN1(n662), .IN2(U6954_n1), .Q(n3125) );
  INVX0 U6955_U2 ( .INP(n2726), .ZN(U6955_n1) );
  AND2X1 U6955_U1 ( .IN1(n646), .IN2(U6955_n1), .Q(n3105) );
  INVX0 U6956_U2 ( .INP(n3146), .ZN(U6956_n1) );
  AND2X1 U6956_U1 ( .IN1(n333), .IN2(U6956_n1), .Q(n3145) );
  INVX0 U6957_U2 ( .INP(n3165), .ZN(U6957_n1) );
  AND2X1 U6957_U1 ( .IN1(n658), .IN2(U6957_n1), .Q(n3164) );
  INVX0 U7174_U2 ( .INP(n5288), .ZN(U7174_n1) );
  AND2X1 U7174_U1 ( .IN1(n2423), .IN2(U7174_n1), .Q(n2422) );
  INVX0 U7248_U2 ( .INP(g1536), .ZN(U7248_n1) );
  AND2X1 U7248_U1 ( .IN1(n4172), .IN2(U7248_n1), .Q(n4173) );
  INVX0 U7249_U2 ( .INP(g1193), .ZN(U7249_n1) );
  AND2X1 U7249_U1 ( .IN1(n4190), .IN2(U7249_n1), .Q(n4191) );
  INVX0 U7402_U2 ( .INP(n4020), .ZN(U7402_n1) );
  AND2X1 U7402_U1 ( .IN1(n4034), .IN2(U7402_n1), .Q(n4037) );
  INVX0 U7405_U2 ( .INP(n4014), .ZN(U7405_n1) );
  AND2X1 U7405_U1 ( .IN1(n4034), .IN2(U7405_n1), .Q(n4039) );
  INVX0 U7413_U2 ( .INP(n3947), .ZN(U7413_n1) );
  AND2X1 U7413_U1 ( .IN1(n3969), .IN2(U7413_n1), .Q(n3972) );
  INVX0 U7416_U2 ( .INP(n3904), .ZN(U7416_n1) );
  AND2X1 U7416_U1 ( .IN1(n3926), .IN2(U7416_n1), .Q(n3929) );
  INVX0 U7427_U2 ( .INP(n3838), .ZN(U7427_n1) );
  AND2X1 U7427_U1 ( .IN1(n3860), .IN2(U7427_n1), .Q(n3863) );
  INVX0 U7438_U2 ( .INP(n3978), .ZN(U7438_n1) );
  AND2X1 U7438_U1 ( .IN1(n4002), .IN2(U7438_n1), .Q(n4003) );
  INVX0 U7449_U2 ( .INP(n4017), .ZN(U7449_n1) );
  AND2X1 U7449_U1 ( .IN1(n4034), .IN2(U7449_n1), .Q(n4032) );
  INVX0 U7455_U2 ( .INP(n3495), .ZN(U7455_n1) );
  AND2X1 U7455_U1 ( .IN1(n4034), .IN2(U7455_n1), .Q(n4035) );
  INVX0 U7464_U2 ( .INP(n3773), .ZN(U7464_n1) );
  AND2X1 U7464_U1 ( .IN1(n3792), .IN2(U7464_n1), .Q(n3797) );
  INVX0 U7467_U2 ( .INP(n3776), .ZN(U7467_n1) );
  AND2X1 U7467_U1 ( .IN1(n3792), .IN2(U7467_n1), .Q(n3790) );
  INVX0 U7482_U2 ( .INP(n3770), .ZN(U7482_n1) );
  AND2X1 U7482_U1 ( .IN1(n3792), .IN2(U7482_n1), .Q(n3795) );
  INVX0 U7492_U2 ( .INP(n3877), .ZN(U7492_n1) );
  AND2X1 U7492_U1 ( .IN1(n3893), .IN2(U7492_n1), .Q(n3891) );
  INVX0 U7513_U2 ( .INP(n3802), .ZN(U7513_n1) );
  AND2X1 U7513_U1 ( .IN1(n3826), .IN2(U7513_n1), .Q(n3827) );
  INVX0 U7516_U2 ( .INP(n3871), .ZN(U7516_n1) );
  AND2X1 U7516_U1 ( .IN1(n3893), .IN2(U7516_n1), .Q(n3896) );
  INVX0 U7549_U2 ( .INP(n3983), .ZN(U7549_n1) );
  AND2X1 U7549_U1 ( .IN1(n4002), .IN2(U7549_n1), .Q(n4007) );
  INVX0 U7561_U2 ( .INP(n3907), .ZN(U7561_n1) );
  AND2X1 U7561_U1 ( .IN1(n3926), .IN2(U7561_n1), .Q(n3931) );
  INVX0 U7574_U2 ( .INP(n3768), .ZN(U7574_n1) );
  AND2X1 U7574_U1 ( .IN1(n3792), .IN2(U7574_n1), .Q(n3793) );
  INVX0 U7577_U2 ( .INP(n3910), .ZN(U7577_n1) );
  AND2X1 U7577_U1 ( .IN1(n3926), .IN2(U7577_n1), .Q(n3924) );
  INVX0 U7585_U2 ( .INP(n3807), .ZN(U7585_n1) );
  AND2X1 U7585_U1 ( .IN1(n3826), .IN2(U7585_n1), .Q(n3831) );
  INVX0 U7595_U2 ( .INP(n3804), .ZN(U7595_n1) );
  AND2X1 U7595_U1 ( .IN1(n3826), .IN2(U7595_n1), .Q(n3829) );
  INVX0 U7614_U2 ( .INP(n3902), .ZN(U7614_n1) );
  AND2X1 U7614_U1 ( .IN1(n3926), .IN2(U7614_n1), .Q(n3927) );
  INVX0 U7621_U2 ( .INP(n3950), .ZN(U7621_n1) );
  AND2X1 U7621_U1 ( .IN1(n3969), .IN2(U7621_n1), .Q(n3974) );
  INVX0 U7629_U2 ( .INP(n3874), .ZN(U7629_n1) );
  AND2X1 U7629_U1 ( .IN1(n3893), .IN2(U7629_n1), .Q(n3898) );
  INVX0 U7636_U2 ( .INP(n3945), .ZN(U7636_n1) );
  AND2X1 U7636_U1 ( .IN1(n3969), .IN2(U7636_n1), .Q(n3970) );
  INVX0 U7639_U2 ( .INP(n3986), .ZN(U7639_n1) );
  AND2X1 U7639_U1 ( .IN1(n4002), .IN2(U7639_n1), .Q(n4000) );
  INVX0 U7649_U2 ( .INP(n3841), .ZN(U7649_n1) );
  AND2X1 U7649_U1 ( .IN1(n3860), .IN2(U7649_n1), .Q(n3865) );
  INVX0 U7652_U2 ( .INP(n3836), .ZN(U7652_n1) );
  AND2X1 U7652_U1 ( .IN1(n3860), .IN2(U7652_n1), .Q(n3861) );
  INVX0 U7668_U2 ( .INP(n3810), .ZN(U7668_n1) );
  AND2X1 U7668_U1 ( .IN1(n3826), .IN2(U7668_n1), .Q(n3824) );
  INVX0 U7673_U2 ( .INP(n3869), .ZN(U7673_n1) );
  AND2X1 U7673_U1 ( .IN1(n3893), .IN2(U7673_n1), .Q(n3894) );
  INVX0 U7690_U2 ( .INP(n3953), .ZN(U7690_n1) );
  AND2X1 U7690_U1 ( .IN1(n3969), .IN2(U7690_n1), .Q(n3967) );
  INVX0 U7707_U2 ( .INP(n3844), .ZN(U7707_n1) );
  AND2X1 U7707_U1 ( .IN1(n3860), .IN2(U7707_n1), .Q(n3858) );
  INVX0 U7712_U2 ( .INP(n3980), .ZN(U7712_n1) );
  AND2X1 U7712_U1 ( .IN1(n4002), .IN2(U7712_n1), .Q(n4005) );
  AND2X1 U7792_U2 ( .IN1(g952), .IN2(U7792_n1), .Q(n2505) );
  INVX0 U7792_U1 ( .INP(n10893), .ZN(U7792_n1) );
  AND2X1 U7794_U2 ( .IN1(g1296), .IN2(U7794_n1), .Q(n2499) );
  INVX0 U7794_U1 ( .INP(n10893), .ZN(U7794_n1) );
  INVX0 U7895_U2 ( .INP(g113), .ZN(U7895_n1) );
  AND2X1 U7895_U1 ( .IN1(n2668), .IN2(U7895_n1), .Q(n2760) );
  INVX0 U7897_U2 ( .INP(g31), .ZN(U7897_n1) );
  AND2X1 U7897_U1 ( .IN1(g6), .IN2(U7897_n1), .Q(n3395) );
  AND2X1 U7977_U2 ( .IN1(g661), .IN2(U7977_n1), .Q(n4956) );
  INVX0 U7977_U1 ( .INP(n10892), .ZN(U7977_n1) );
  INVX0 U8034_U2 ( .INP(n5612), .ZN(U8034_n1) );
  AND2X1 U8034_U1 ( .IN1(n4723), .IN2(U8034_n1), .Q(n5026) );
  INVX0 U8036_U2 ( .INP(n5340), .ZN(U8036_n1) );
  AND2X1 U8036_U1 ( .IN1(n3729), .IN2(U8036_n1), .Q(n3941) );
  INVX0 U8050_U2 ( .INP(g1367), .ZN(U8050_n1) );
  AND2X1 U8050_U1 ( .IN1(n173), .IN2(U8050_n1), .Q(n3733) );
  AND2X1 U8055_U2 ( .IN1(g1345), .IN2(U8055_n1), .Q(n4798) );
  INVX0 U8055_U1 ( .INP(n10893), .ZN(U8055_n1) );
  AND2X1 U8060_U2 ( .IN1(g1002), .IN2(U8060_n1), .Q(n4805) );
  INVX0 U8060_U1 ( .INP(n10893), .ZN(U8060_n1) );
  INVX0 U8070_U2 ( .INP(g1361), .ZN(U8070_n1) );
  AND2X1 U8070_U1 ( .IN1(n174), .IN2(U8070_n1), .Q(n4175) );
  INVX0 U8074_U2 ( .INP(g1018), .ZN(U8074_n1) );
  AND2X1 U8074_U1 ( .IN1(n516), .IN2(U8074_n1), .Q(n4193) );
  INVX0 U8088_U2 ( .INP(g1024), .ZN(U8088_n1) );
  AND2X1 U8088_U1 ( .IN1(n515), .IN2(U8088_n1), .Q(n3738) );
  INVX0 U8112_U2 ( .INP(n4523), .ZN(U8112_n1) );
  AND2X1 U8112_U1 ( .IN1(n4525), .IN2(U8112_n1), .Q(n4524) );
  INVX0 U8113_U2 ( .INP(n5751), .ZN(U8113_n1) );
  AND2X1 U8113_U1 ( .IN1(n4526), .IN2(U8113_n1), .Q(n4523) );
  INVX0 U8147_U2 ( .INP(n2573), .ZN(U8147_n1) );
  AND2X1 U8147_U1 ( .IN1(g4659), .IN2(U8147_n1), .Q(n2577) );
  INVX0 U8165_U2 ( .INP(n2563), .ZN(U8165_n1) );
  AND2X1 U8165_U1 ( .IN1(g4849), .IN2(U8165_n1), .Q(n2567) );
  INVX0 U8185_U2 ( .INP(g1046), .ZN(U8185_n1) );
  AND2X1 U8185_U1 ( .IN1(n4940), .IN2(U8185_n1), .Q(n4938) );
  INVX0 U8192_U2 ( .INP(g1389), .ZN(U8192_n1) );
  AND2X1 U8192_U1 ( .IN1(n4915), .IN2(U8192_n1), .Q(n4913) );
  INVX0 U8210_U2 ( .INP(n4723), .ZN(U8210_n1) );
  AND2X1 U8210_U1 ( .IN1(n4722), .IN2(U8210_n1), .Q(n4714) );
  INVX0 U8223_U2 ( .INP(n4516), .ZN(U8223_n1) );
  AND2X1 U8223_U1 ( .IN1(n4518), .IN2(U8223_n1), .Q(n4517) );
  INVX0 U8224_U2 ( .INP(n5728), .ZN(U8224_n1) );
  AND2X1 U8224_U1 ( .IN1(n4519), .IN2(U8224_n1), .Q(n4516) );
  AND2X1 U8281_U2 ( .IN1(n879), .IN2(U8281_n1), .Q(n5111) );
  INVX0 U8281_U1 ( .INP(n10893), .ZN(U8281_n1) );
  AND2X1 U8307_U2 ( .IN1(g29216), .IN2(U8307_n1), .Q(g26900) );
  INVX0 U8307_U1 ( .INP(n10892), .ZN(U8307_n1) );
  INVX0 U8974_U2 ( .INP(test_so25), .ZN(U8974_n1) );
  AND2X1 U8974_U1 ( .IN1(n3362), .IN2(U8974_n1), .Q(n2552) );
  INVX0 U8975_U2 ( .INP(g528), .ZN(U8975_n1) );
  AND2X1 U8975_U1 ( .IN1(n3174), .IN2(U8975_n1), .Q(n3195) );
  AND2X1 U9065_U2 ( .IN1(g4145), .IN2(U9065_n1), .Q(n4721) );
  INVX0 U9065_U1 ( .INP(n10893), .ZN(U9065_n1) );
  AND2X1 U9070_U2 ( .IN1(g2841), .IN2(U9070_n1), .Q(n3730) );
  INVX0 U9070_U1 ( .INP(n10893), .ZN(U9070_n1) );
  INVX0 U9075_U2 ( .INP(g9), .ZN(U9075_n1) );
  AND2X1 U9075_U1 ( .IN1(g19), .IN2(U9075_n1), .Q(n3362) );
  AND2X1 U9076_U2 ( .IN1(g113), .IN2(U9076_n1), .Q(g25694) );
  INVX0 U9076_U1 ( .INP(n10893), .ZN(U9076_n1) );
  AND2X1 U9080_U2 ( .IN1(n4305), .IN2(U9080_n1), .Q(g29277) );
  INVX0 U9080_U1 ( .INP(n10893), .ZN(U9080_n1) );
  AND2X1 U9084_U2 ( .IN1(g4423), .IN2(U9084_n1), .Q(g26953) );
  INVX0 U9084_U1 ( .INP(n10892), .ZN(U9084_n1) );
  AND2X1 U9085_U2 ( .IN1(g64), .IN2(U9085_n1), .Q(g24212) );
  INVX0 U9085_U1 ( .INP(n10893), .ZN(U9085_n1) );
  AND2X1 U9086_U2 ( .IN1(n4283), .IN2(U9086_n1), .Q(g29279) );
  INVX0 U9086_U1 ( .INP(n10892), .ZN(U9086_n1) );
  AND2X1 U9090_U2 ( .IN1(g125), .IN2(U9090_n1), .Q(g25688) );
  INVX0 U9090_U1 ( .INP(n10893), .ZN(U9090_n1) );
  INVX0 U9098_U2 ( .INP(n290), .ZN(U9098_n1) );
  AND2X1 U9098_U1 ( .IN1(g4681), .IN2(U9098_n1), .Q(g34028) );
  INVX0 U9099_U2 ( .INP(n2608), .ZN(U9099_n1) );
  AND2X1 U9099_U1 ( .IN1(n2595), .IN2(U9099_n1), .Q(g34449) );
  AND2X1 U9101_U2 ( .IN1(g6745), .IN2(U9101_n1), .Q(g26880) );
  INVX0 U9101_U1 ( .INP(n10893), .ZN(U9101_n1) );
  INVX0 U9107_U2 ( .INP(n10544), .ZN(U9107_n1) );
  AND2X1 U9107_U1 ( .IN1(n4448), .IN2(U9107_n1), .Q(n4447) );
  INVX0 U9111_U2 ( .INP(n10541), .ZN(U9111_n1) );
  AND2X1 U9111_U1 ( .IN1(n4403), .IN2(U9111_n1), .Q(n4402) );
  INVX0 U9116_U2 ( .INP(n10549), .ZN(U9116_n1) );
  AND2X1 U9116_U1 ( .IN1(n4426), .IN2(U9116_n1), .Q(n4425) );
  INVX0 U9120_U2 ( .INP(n10538), .ZN(U9120_n1) );
  AND2X1 U9120_U1 ( .IN1(n4437), .IN2(U9120_n1), .Q(n4436) );
  INVX0 U9124_U2 ( .INP(n10546), .ZN(U9124_n1) );
  AND2X1 U9124_U1 ( .IN1(n4392), .IN2(U9124_n1), .Q(n4391) );
  INVX0 U9128_U2 ( .INP(n10539), .ZN(U9128_n1) );
  AND2X1 U9128_U1 ( .IN1(n4380), .IN2(U9128_n1), .Q(n4379) );
  INVX0 U9132_U2 ( .INP(n10547), .ZN(U9132_n1) );
  AND2X1 U9132_U1 ( .IN1(n4415), .IN2(U9132_n1), .Q(n4414) );
  INVX0 U9136_U2 ( .INP(n10548), .ZN(U9136_n1) );
  AND2X1 U9136_U1 ( .IN1(n4459), .IN2(U9136_n1), .Q(n4458) );
  INVX0 U9315_U2 ( .INP(n5753), .ZN(U9315_n1) );
  AND2X1 U9315_U1 ( .IN1(n5016), .IN2(U9315_n1), .Q(n5014) );
  INVX0 U9453_U2 ( .INP(n10542), .ZN(U9453_n1) );
  AND2X1 U9453_U1 ( .IN1(n3065), .IN2(U9453_n1), .Q(n3064) );
  INVX0 U9825_U2 ( .INP(n1698), .ZN(U9825_n1) );
  AND2X1 U9825_U1 ( .IN1(g112), .IN2(U9825_n1), .Q(n3115) );
  INVX0 U9886_U2 ( .INP(n5121), .ZN(U9886_n1) );
  AND2X1 U9886_U1 ( .IN1(g370), .IN2(U9886_n1), .Q(n4948) );
  INVX0 U9927_U2 ( .INP(g4098), .ZN(U9927_n1) );
  AND2X1 U9927_U1 ( .IN1(n3933), .IN2(U9927_n1), .Q(n3833) );
  INVX0 U9953_U2 ( .INP(n120), .ZN(U9953_n1) );
  AND2X1 U9953_U1 ( .IN1(g671), .IN2(U9953_n1), .Q(n4526) );
  INVX0 U9957_U2 ( .INP(n5283), .ZN(U9957_n1) );
  AND2X1 U9957_U1 ( .IN1(g4843), .IN2(U9957_n1), .Q(n2563) );
  INVX0 U9958_U2 ( .INP(n5656), .ZN(U9958_n1) );
  AND2X1 U9958_U1 ( .IN1(test_so19), .IN2(U9958_n1), .Q(n2573) );
  INVX0 U9968_U2 ( .INP(g4358), .ZN(U9968_n1) );
  AND2X1 U9968_U1 ( .IN1(n3084), .IN2(U9968_n1), .Q(n3023) );
  INVX0 U9972_U2 ( .INP(n4535), .ZN(U9972_n1) );
  AND2X1 U9972_U1 ( .IN1(g681), .IN2(U9972_n1), .Q(n5112) );
  INVX0 U9992_U2 ( .INP(n3676), .ZN(U9992_n1) );
  AND2X1 U9992_U1 ( .IN1(n3675), .IN2(U9992_n1), .Q(n2644) );
  INVX0 U10314_U2 ( .INP(g686), .ZN(U10314_n1) );
  AND2X1 U10314_U1 ( .IN1(g667), .IN2(U10314_n1), .Q(n4962) );
  INVX0 U10318_U2 ( .INP(n5681), .ZN(U10318_n1) );
  AND2X1 U10318_U1 ( .IN1(g5092), .IN2(U10318_n1), .Q(n5016) );
endmodule

