module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n236_, new_n238_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n186_, new_n365_, new_n339_, new_n197_, new_n401_, new_n389_, new_n456_, new_n246_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n214_, new_n451_, new_n424_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n123_, new_n342_, new_n462_, new_n317_, new_n344_, new_n287_, new_n427_, new_n234_, new_n393_, new_n418_, new_n292_, new_n215_, new_n157_, new_n153_, new_n257_, new_n212_, new_n364_, new_n449_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n124_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n248_, new_n350_, new_n167_, new_n385_, new_n461_, new_n297_, new_n361_, new_n183_, new_n463_, new_n303_, new_n351_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n158_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n423_, new_n205_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n256_, new_n452_, new_n381_, new_n388_, new_n194_, new_n394_, new_n299_, new_n142_, new_n139_, new_n314_, new_n363_, new_n165_, new_n441_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n162_, new_n409_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n371_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n460_, new_n130_, new_n268_, new_n374_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n145_, new_n253_, new_n403_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n182_, new_n407_, new_n151_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n428_, new_n199_, new_n146_, new_n360_, new_n302_, new_n191_, new_n225_, new_n387_, new_n121_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n255_, new_n459_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n340_, new_n285_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n332_, new_n453_, new_n163_, new_n148_, new_n440_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n307_, new_n190_, new_n408_, new_n213_, new_n435_, new_n265_, new_n370_, new_n278_, new_n217_, new_n269_, new_n129_, new_n412_, new_n327_, new_n431_, new_n196_, new_n319_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n467_, new_n404_, new_n193_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n455_, new_n120_, new_n406_, new_n356_, new_n229_, new_n464_, new_n204_, new_n181_, new_n135_, new_n405_;

not g000 ( new_n119_, N29 );
not g001 ( new_n120_, N42 );
not g002 ( new_n121_, N75 );
nor g003 ( N388, new_n119_, new_n120_, new_n121_ );
not g004 ( new_n123_, N36 );
not g005 ( new_n124_, N80 );
nor g006 ( N389, new_n119_, new_n123_, new_n124_ );
nor g007 ( N390, new_n119_, new_n123_, new_n120_ );
and g008 ( N391, N85, N86 );
and g009 ( N418, N1, N8, N13, N17 );
not g010 ( new_n129_, N390 );
and g011 ( new_n130_, N1, N13, N17, N26 );
nand g012 ( N419, new_n129_, new_n130_ );
nand g013 ( N420, N59, N75, N80 );
nand g014 ( N421, N36, N59, N80 );
nand g015 ( N422, N36, N42, N59 );
not g016 ( new_n135_, N90 );
nor g017 ( new_n136_, N87, N88 );
nor g018 ( N423, new_n136_, new_n135_ );
nand g019 ( N446, N390, new_n130_ );
nand g020 ( new_n139_, N1, N26, N51 );
nand g021 ( new_n140_, new_n139_, keyIn_0_0 );
not g022 ( new_n141_, keyIn_0_0 );
nand g023 ( new_n142_, new_n141_, N1, N26, N51 );
nand g024 ( new_n143_, new_n140_, new_n142_ );
not g025 ( N447, new_n143_ );
not g026 ( new_n145_, N68 );
nand g027 ( new_n146_, N1, N8, N13, N55 );
nor g028 ( N448, new_n146_, new_n119_, new_n145_ );
not g029 ( new_n148_, N74 );
nand g030 ( new_n149_, N59, N68 );
nor g031 ( N449, new_n146_, new_n148_, new_n149_ );
not g032 ( new_n151_, N89 );
nor g033 ( N450, new_n136_, new_n151_ );
xnor g034 ( new_n153_, N91, N96 );
xnor g035 ( new_n154_, N101, N106 );
xnor g036 ( new_n155_, new_n153_, new_n154_ );
xnor g037 ( new_n156_, new_n155_, N130 );
xor g038 ( new_n157_, N111, N116 );
xnor g039 ( new_n158_, N121, N126 );
xnor g040 ( new_n159_, new_n157_, new_n158_ );
xnor g041 ( new_n160_, new_n159_, N135 );
xnor g042 ( N767, new_n160_, new_n156_ );
xnor g043 ( new_n162_, N159, N165 );
xnor g044 ( new_n163_, N171, N177 );
xnor g045 ( new_n164_, new_n162_, new_n163_ );
xnor g046 ( new_n165_, new_n164_, N130 );
xor g047 ( new_n166_, N183, N189 );
xnor g048 ( new_n167_, N195, N201 );
xnor g049 ( new_n168_, new_n166_, new_n167_ );
xnor g050 ( new_n169_, new_n168_, N207 );
xnor g051 ( N768, new_n169_, new_n165_ );
not g052 ( new_n171_, keyIn_0_10 );
not g053 ( new_n172_, keyIn_0_9 );
not g054 ( new_n173_, keyIn_0_7 );
not g055 ( new_n174_, keyIn_0_4 );
nand g056 ( new_n175_, new_n143_, new_n174_ );
nand g057 ( new_n176_, new_n140_, keyIn_0_4, new_n142_ );
nand g058 ( new_n177_, new_n175_, new_n176_ );
nand g059 ( new_n178_, new_n177_, new_n173_ );
nand g060 ( new_n179_, new_n175_, keyIn_0_7, new_n176_ );
nand g061 ( new_n180_, new_n178_, new_n179_ );
nand g062 ( new_n181_, N17, N42 );
nand g063 ( new_n182_, new_n181_, keyIn_0_3 );
not g064 ( new_n183_, keyIn_0_3 );
nand g065 ( new_n184_, new_n183_, N17, N42 );
and g066 ( new_n185_, new_n182_, new_n184_ );
not g067 ( new_n186_, N17 );
nand g068 ( new_n187_, new_n186_, new_n120_, keyIn_0_2 );
not g069 ( new_n188_, keyIn_0_2 );
or g070 ( new_n189_, N17, N42 );
nand g071 ( new_n190_, new_n189_, new_n188_ );
nand g072 ( new_n191_, new_n185_, keyIn_0_6, new_n187_, new_n190_ );
and g073 ( new_n192_, N59, N156 );
not g074 ( new_n193_, keyIn_0_6 );
nand g075 ( new_n194_, new_n190_, new_n182_, new_n184_, new_n187_ );
nand g076 ( new_n195_, new_n194_, new_n193_ );
and g077 ( new_n196_, new_n195_, new_n191_, new_n192_ );
nand g078 ( new_n197_, new_n180_, new_n196_ );
nand g079 ( new_n198_, new_n197_, new_n172_ );
nand g080 ( new_n199_, new_n180_, keyIn_0_9, new_n196_ );
nand g081 ( new_n200_, new_n198_, new_n199_ );
nand g082 ( new_n201_, N1, N8, N17, N51 );
xnor g083 ( new_n202_, new_n201_, keyIn_0_1 );
or g084 ( new_n203_, new_n202_, keyIn_0_5 );
nand g085 ( new_n204_, N42, N59, N75 );
nand g086 ( new_n205_, new_n202_, keyIn_0_5 );
nand g087 ( new_n206_, new_n203_, new_n205_, new_n204_ );
xnor g088 ( new_n207_, new_n206_, keyIn_0_8 );
nand g089 ( new_n208_, new_n200_, new_n207_ );
nand g090 ( new_n209_, new_n208_, new_n171_ );
nand g091 ( new_n210_, new_n200_, keyIn_0_10, new_n207_ );
nand g092 ( new_n211_, new_n209_, new_n210_ );
nand g093 ( new_n212_, new_n211_, N126 );
not g094 ( new_n213_, new_n180_ );
nor g095 ( new_n214_, new_n213_, new_n192_ );
nand g096 ( new_n215_, new_n214_, N17 );
nand g097 ( new_n216_, new_n215_, N1 );
nand g098 ( new_n217_, new_n216_, N153 );
not g099 ( new_n218_, N268 );
nor g100 ( new_n219_, new_n213_, new_n119_, new_n121_, new_n124_ );
nand g101 ( new_n220_, new_n219_, N55, new_n218_ );
and g102 ( new_n221_, new_n217_, new_n220_ );
nand g103 ( new_n222_, new_n212_, new_n221_ );
and g104 ( new_n223_, new_n222_, N201 );
not g105 ( new_n224_, N201 );
nand g106 ( new_n225_, new_n212_, new_n224_, new_n221_ );
not g107 ( new_n226_, new_n225_ );
nor g108 ( new_n227_, new_n223_, new_n226_ );
nand g109 ( new_n228_, new_n227_, N261 );
or g110 ( new_n229_, new_n227_, N261 );
nand g111 ( new_n230_, new_n229_, N219, new_n228_ );
nand g112 ( new_n231_, new_n227_, N228 );
and g113 ( new_n232_, new_n223_, N237 );
and g114 ( new_n233_, new_n222_, N246 );
nand g115 ( new_n234_, N42, N72, N73 );
nor g116 ( new_n235_, new_n146_, new_n234_, new_n149_ );
nand g117 ( new_n236_, new_n235_, N201 );
nand g118 ( new_n237_, N255, N267 );
nand g119 ( new_n238_, N121, N210 );
nand g120 ( new_n239_, new_n236_, new_n237_, new_n238_ );
nor g121 ( new_n240_, new_n232_, new_n233_, new_n239_ );
nand g122 ( N850, new_n230_, new_n231_, new_n240_ );
not g123 ( new_n242_, keyIn_0_14 );
nand g124 ( new_n243_, new_n211_, keyIn_0_11, N111 );
nand g125 ( new_n244_, new_n216_, N143 );
not g126 ( new_n245_, keyIn_0_11 );
nand g127 ( new_n246_, new_n211_, N111 );
nand g128 ( new_n247_, new_n246_, new_n245_ );
nand g129 ( new_n248_, new_n247_, keyIn_0_12, new_n243_, new_n244_ );
not g130 ( new_n249_, keyIn_0_12 );
nand g131 ( new_n250_, new_n247_, new_n243_, new_n244_ );
nand g132 ( new_n251_, new_n250_, new_n249_ );
nand g133 ( new_n252_, new_n251_, new_n220_, new_n248_ );
nand g134 ( new_n253_, new_n252_, keyIn_0_13 );
not g135 ( new_n254_, keyIn_0_13 );
nand g136 ( new_n255_, new_n251_, new_n254_, new_n220_, new_n248_ );
nand g137 ( new_n256_, new_n253_, new_n255_ );
nand g138 ( new_n257_, new_n256_, N183 );
nand g139 ( new_n258_, new_n257_, new_n242_ );
nand g140 ( new_n259_, new_n256_, keyIn_0_14, N183 );
nand g141 ( new_n260_, new_n258_, new_n259_ );
not g142 ( new_n261_, new_n260_ );
not g143 ( new_n262_, keyIn_0_15 );
not g144 ( new_n263_, N183 );
nand g145 ( new_n264_, new_n253_, new_n263_, new_n255_ );
nand g146 ( new_n265_, new_n264_, new_n262_ );
or g147 ( new_n266_, new_n264_, new_n262_ );
and g148 ( new_n267_, new_n266_, new_n265_ );
nand g149 ( new_n268_, new_n261_, new_n267_ );
not g150 ( new_n269_, new_n268_ );
not g151 ( new_n270_, keyIn_0_18 );
nand g152 ( new_n271_, new_n211_, N116 );
nand g153 ( new_n272_, new_n216_, N146 );
nand g154 ( new_n273_, new_n271_, new_n220_, new_n272_ );
or g155 ( new_n274_, new_n273_, N189 );
not g156 ( new_n275_, N195 );
nand g157 ( new_n276_, new_n211_, N121 );
nand g158 ( new_n277_, new_n216_, N149 );
and g159 ( new_n278_, new_n277_, new_n220_ );
nand g160 ( new_n279_, new_n276_, new_n275_, new_n278_ );
xnor g161 ( new_n280_, new_n279_, keyIn_0_16 );
and g162 ( new_n281_, new_n225_, N261 );
nand g163 ( new_n282_, new_n280_, new_n274_, new_n281_ );
xnor g164 ( new_n283_, new_n282_, new_n270_ );
nand g165 ( new_n284_, new_n280_, new_n223_, new_n274_ );
nand g166 ( new_n285_, new_n273_, N189 );
nand g167 ( new_n286_, new_n276_, new_n278_ );
and g168 ( new_n287_, new_n286_, N195 );
nand g169 ( new_n288_, new_n274_, new_n287_ );
and g170 ( new_n289_, new_n288_, new_n285_ );
nand g171 ( new_n290_, new_n283_, new_n284_, new_n289_ );
or g172 ( new_n291_, new_n269_, new_n290_ );
nand g173 ( new_n292_, new_n269_, new_n290_ );
nand g174 ( new_n293_, new_n291_, N219, new_n292_ );
nand g175 ( new_n294_, new_n260_, keyIn_0_17 );
not g176 ( new_n295_, keyIn_0_17 );
nand g177 ( new_n296_, new_n258_, new_n295_, new_n259_ );
nand g178 ( new_n297_, new_n294_, new_n296_ );
nand g179 ( new_n298_, new_n297_, N237 );
nand g180 ( new_n299_, new_n269_, N228 );
nand g181 ( new_n300_, new_n256_, N246 );
nand g182 ( new_n301_, N106, N210 );
nand g183 ( new_n302_, new_n235_, N183 );
and g184 ( new_n303_, new_n299_, new_n300_, new_n301_, new_n302_ );
nand g185 ( N863, new_n303_, new_n293_, new_n298_ );
not g186 ( new_n305_, new_n287_ );
nor g187 ( new_n306_, new_n281_, new_n223_ );
not g188 ( new_n307_, new_n306_ );
nand g189 ( new_n308_, new_n307_, new_n280_ );
nand g190 ( new_n309_, new_n308_, new_n305_ );
nand g191 ( new_n310_, new_n274_, new_n285_ );
not g192 ( new_n311_, new_n310_ );
nand g193 ( new_n312_, new_n309_, new_n311_ );
nand g194 ( new_n313_, new_n308_, new_n305_, new_n310_ );
nand g195 ( new_n314_, new_n312_, N219, new_n313_ );
nand g196 ( new_n315_, new_n311_, N228 );
not g197 ( new_n316_, N237 );
nor g198 ( new_n317_, new_n285_, new_n316_ );
and g199 ( new_n318_, new_n273_, N246 );
nand g200 ( new_n319_, new_n235_, N189 );
nand g201 ( new_n320_, N255, N259 );
nand g202 ( new_n321_, N111, N210 );
nand g203 ( new_n322_, new_n319_, new_n320_, new_n321_ );
nor g204 ( new_n323_, new_n317_, new_n318_, new_n322_ );
nand g205 ( N864, new_n314_, new_n315_, new_n323_ );
nand g206 ( new_n325_, new_n280_, new_n305_ );
nand g207 ( new_n326_, new_n325_, new_n306_ );
not g208 ( new_n327_, new_n325_ );
nand g209 ( new_n328_, new_n327_, new_n307_ );
nand g210 ( new_n329_, new_n328_, N219, new_n326_ );
nand g211 ( new_n330_, new_n327_, N228 );
nor g212 ( new_n331_, new_n305_, new_n316_ );
and g213 ( new_n332_, new_n286_, N246 );
nand g214 ( new_n333_, new_n235_, N195 );
nand g215 ( new_n334_, N255, N260 );
nand g216 ( new_n335_, N116, N210 );
nand g217 ( new_n336_, new_n333_, new_n334_, new_n335_ );
nor g218 ( new_n337_, new_n331_, new_n332_, new_n336_ );
nand g219 ( N865, new_n329_, new_n330_, new_n337_ );
nand g220 ( new_n339_, new_n294_, keyIn_0_21, new_n296_ );
not g221 ( new_n340_, keyIn_0_22 );
nand g222 ( new_n341_, new_n290_, new_n265_, new_n266_ );
nand g223 ( new_n342_, new_n341_, new_n340_ );
nand g224 ( new_n343_, new_n290_, keyIn_0_22, new_n266_, new_n265_ );
nand g225 ( new_n344_, new_n342_, new_n343_ );
not g226 ( new_n345_, keyIn_0_21 );
nand g227 ( new_n346_, new_n297_, new_n345_ );
nand g228 ( new_n347_, new_n346_, new_n339_, new_n344_ );
nand g229 ( new_n348_, new_n347_, keyIn_0_23 );
not g230 ( new_n349_, keyIn_0_23 );
nand g231 ( new_n350_, new_n346_, new_n349_, new_n344_, new_n339_ );
nand g232 ( new_n351_, new_n348_, new_n350_ );
nand g233 ( new_n352_, new_n211_, N106 );
and g234 ( new_n353_, new_n214_, N55 );
nand g235 ( new_n354_, new_n353_, N153 );
nand g236 ( new_n355_, N138, N152 );
nand g237 ( new_n356_, new_n219_, N17, new_n218_ );
nand g238 ( new_n357_, new_n352_, new_n354_, new_n355_, new_n356_ );
nor g239 ( new_n358_, new_n357_, N177 );
not g240 ( new_n359_, new_n358_ );
nand g241 ( new_n360_, new_n351_, new_n359_ );
nand g242 ( new_n361_, new_n357_, N177 );
nand g243 ( new_n362_, new_n360_, new_n361_ );
nand g244 ( new_n363_, new_n211_, N101 );
nand g245 ( new_n364_, new_n353_, N149 );
nand g246 ( new_n365_, N17, N138 );
nand g247 ( new_n366_, new_n363_, new_n356_, new_n364_, new_n365_ );
or g248 ( new_n367_, new_n366_, N171 );
nand g249 ( new_n368_, new_n362_, new_n367_ );
nand g250 ( new_n369_, new_n366_, N171 );
nand g251 ( new_n370_, new_n368_, new_n369_ );
nand g252 ( new_n371_, new_n211_, N96 );
nand g253 ( new_n372_, new_n353_, N146 );
nand g254 ( new_n373_, N51, N138 );
nand g255 ( new_n374_, new_n371_, new_n356_, new_n372_, new_n373_ );
or g256 ( new_n375_, new_n374_, N165 );
nand g257 ( new_n376_, new_n370_, new_n375_ );
nand g258 ( new_n377_, new_n374_, N165 );
nand g259 ( new_n378_, new_n376_, new_n377_ );
nand g260 ( new_n379_, new_n211_, N91 );
nand g261 ( new_n380_, new_n353_, N143 );
nand g262 ( new_n381_, N8, N138 );
nand g263 ( new_n382_, new_n379_, new_n356_, new_n380_, new_n381_ );
or g264 ( new_n383_, new_n382_, N159 );
nand g265 ( new_n384_, new_n378_, new_n383_ );
nand g266 ( new_n385_, new_n382_, N159 );
nand g267 ( N866, new_n384_, new_n385_ );
not g268 ( new_n387_, keyIn_0_31 );
not g269 ( new_n388_, keyIn_0_30 );
not g270 ( new_n389_, keyIn_0_27 );
not g271 ( new_n390_, keyIn_0_24 );
nand g272 ( new_n391_, new_n359_, new_n361_ );
nand g273 ( new_n392_, new_n348_, new_n350_, new_n391_ );
nand g274 ( new_n393_, new_n392_, new_n390_ );
not g275 ( new_n394_, new_n391_ );
nand g276 ( new_n395_, new_n351_, new_n394_ );
nand g277 ( new_n396_, new_n395_, keyIn_0_25 );
not g278 ( new_n397_, keyIn_0_25 );
nand g279 ( new_n398_, new_n351_, new_n397_, new_n394_ );
nand g280 ( new_n399_, new_n348_, keyIn_0_24, new_n350_, new_n391_ );
nand g281 ( new_n400_, new_n396_, new_n393_, new_n398_, new_n399_ );
nand g282 ( new_n401_, new_n400_, keyIn_0_26 );
and g283 ( new_n402_, new_n398_, new_n399_ );
not g284 ( new_n403_, keyIn_0_26 );
and g285 ( new_n404_, new_n393_, new_n403_ );
nand g286 ( new_n405_, new_n402_, new_n404_, new_n396_ );
nand g287 ( new_n406_, new_n401_, new_n405_, new_n389_, N219 );
nand g288 ( new_n407_, N101, N210 );
nand g289 ( new_n408_, new_n401_, N219, new_n405_ );
nand g290 ( new_n409_, new_n408_, keyIn_0_27 );
nand g291 ( new_n410_, new_n409_, keyIn_0_28, new_n406_, new_n407_ );
not g292 ( new_n411_, keyIn_0_28 );
nand g293 ( new_n412_, new_n409_, new_n406_, new_n407_ );
nand g294 ( new_n413_, new_n412_, new_n411_ );
and g295 ( new_n414_, new_n394_, N228 );
not g296 ( new_n415_, new_n414_ );
nor g297 ( new_n416_, new_n415_, keyIn_0_20 );
and g298 ( new_n417_, new_n415_, keyIn_0_20 );
nor g299 ( new_n418_, new_n361_, new_n316_ );
nand g300 ( new_n419_, new_n235_, N177 );
nand g301 ( new_n420_, new_n357_, N246 );
nand g302 ( new_n421_, new_n420_, new_n419_ );
nor g303 ( new_n422_, new_n417_, new_n416_, new_n418_, new_n421_ );
nand g304 ( new_n423_, new_n413_, new_n410_, new_n422_ );
nand g305 ( new_n424_, new_n423_, keyIn_0_29 );
not g306 ( new_n425_, keyIn_0_29 );
nand g307 ( new_n426_, new_n413_, new_n425_, new_n410_, new_n422_ );
nand g308 ( new_n427_, new_n424_, new_n426_ );
nand g309 ( new_n428_, new_n427_, new_n388_ );
nand g310 ( new_n429_, new_n424_, keyIn_0_30, new_n426_ );
nand g311 ( new_n430_, new_n428_, new_n429_ );
nand g312 ( new_n431_, new_n430_, new_n387_ );
nand g313 ( new_n432_, new_n428_, keyIn_0_31, new_n429_ );
and g314 ( N874, new_n431_, new_n432_ );
nand g315 ( new_n434_, new_n383_, new_n385_ );
not g316 ( new_n435_, new_n434_ );
nand g317 ( new_n436_, new_n378_, new_n435_ );
nand g318 ( new_n437_, new_n376_, new_n377_, new_n434_ );
nand g319 ( new_n438_, new_n436_, N219, new_n437_ );
nand g320 ( new_n439_, new_n435_, N228 );
nand g321 ( new_n440_, new_n382_, N159, N237 );
nand g322 ( new_n441_, new_n382_, N246 );
nand g323 ( new_n442_, N210, N268 );
nand g324 ( new_n443_, new_n235_, N159 );
and g325 ( new_n444_, new_n440_, new_n441_, new_n442_, new_n443_ );
nand g326 ( N878, new_n438_, new_n439_, new_n444_ );
nand g327 ( new_n446_, new_n375_, new_n377_ );
not g328 ( new_n447_, new_n446_ );
nand g329 ( new_n448_, new_n370_, new_n447_ );
nand g330 ( new_n449_, new_n368_, new_n369_, new_n446_ );
nand g331 ( new_n450_, new_n448_, N219, new_n449_ );
nand g332 ( new_n451_, new_n447_, N228 );
nand g333 ( new_n452_, new_n374_, N165, N237 );
nand g334 ( new_n453_, new_n374_, N246 );
nand g335 ( new_n454_, N91, N210 );
nand g336 ( new_n455_, new_n235_, N165 );
and g337 ( new_n456_, new_n452_, new_n453_, new_n454_, new_n455_ );
nand g338 ( N879, new_n450_, new_n451_, new_n456_ );
and g339 ( new_n458_, new_n367_, new_n369_ );
nand g340 ( new_n459_, new_n362_, new_n458_ );
or g341 ( new_n460_, new_n362_, new_n458_ );
nand g342 ( new_n461_, new_n460_, N219, new_n459_ );
nor g343 ( new_n462_, new_n369_, new_n316_ );
xnor g344 ( new_n463_, new_n462_, keyIn_0_19 );
nand g345 ( new_n464_, new_n458_, N228 );
nand g346 ( new_n465_, new_n366_, N246 );
nand g347 ( new_n466_, N96, N210 );
nand g348 ( new_n467_, new_n235_, N171 );
and g349 ( new_n468_, new_n464_, new_n465_, new_n466_, new_n467_ );
nand g350 ( N880, new_n461_, new_n463_, new_n468_ );
endmodule