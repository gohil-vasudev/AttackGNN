module add_mul_comp_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713;

  OR2_X1 U872 ( .A1(n856), .A2(n857), .ZN(Result_9_) );
  AND2_X1 U873 ( .A1(n858), .A2(n859), .ZN(n857) );
  OR2_X1 U874 ( .A1(n860), .A2(n861), .ZN(n858) );
  INV_X1 U875 ( .A(n862), .ZN(n861) );
  OR2_X1 U876 ( .A1(n863), .A2(n864), .ZN(n862) );
  AND2_X1 U877 ( .A1(n864), .A2(n863), .ZN(n860) );
  AND2_X1 U878 ( .A1(n865), .A2(n866), .ZN(n863) );
  OR2_X1 U879 ( .A1(n867), .A2(n868), .ZN(n866) );
  INV_X1 U880 ( .A(n869), .ZN(n868) );
  OR2_X1 U881 ( .A1(n869), .A2(n870), .ZN(n865) );
  INV_X1 U882 ( .A(n867), .ZN(n870) );
  AND2_X1 U883 ( .A1(n871), .A2(n872), .ZN(n856) );
  OR2_X1 U884 ( .A1(n873), .A2(n874), .ZN(n871) );
  AND2_X1 U885 ( .A1(n875), .A2(n876), .ZN(n874) );
  OR2_X1 U886 ( .A1(n877), .A2(n878), .ZN(n875) );
  AND2_X1 U887 ( .A1(a_1_), .A2(n879), .ZN(n878) );
  AND2_X1 U888 ( .A1(n880), .A2(n881), .ZN(n873) );
  OR2_X1 U889 ( .A1(n882), .A2(n883), .ZN(n881) );
  INV_X1 U890 ( .A(n876), .ZN(n880) );
  OR2_X1 U891 ( .A1(n884), .A2(n885), .ZN(Result_8_) );
  AND2_X1 U892 ( .A1(n886), .A2(n859), .ZN(n885) );
  OR2_X1 U893 ( .A1(n887), .A2(n888), .ZN(n886) );
  AND2_X1 U894 ( .A1(n889), .A2(n890), .ZN(n888) );
  INV_X1 U895 ( .A(n891), .ZN(n887) );
  OR2_X1 U896 ( .A1(n890), .A2(n889), .ZN(n891) );
  OR2_X1 U897 ( .A1(n892), .A2(n893), .ZN(n889) );
  AND2_X1 U898 ( .A1(n894), .A2(n895), .ZN(n893) );
  INV_X1 U899 ( .A(n896), .ZN(n892) );
  OR2_X1 U900 ( .A1(n895), .A2(n894), .ZN(n896) );
  AND2_X1 U901 ( .A1(n897), .A2(n872), .ZN(n884) );
  OR2_X1 U902 ( .A1(n898), .A2(n899), .ZN(n897) );
  INV_X1 U903 ( .A(n900), .ZN(n899) );
  OR2_X1 U904 ( .A1(n901), .A2(n902), .ZN(n900) );
  AND2_X1 U905 ( .A1(n902), .A2(n901), .ZN(n898) );
  OR2_X1 U906 ( .A1(n903), .A2(n883), .ZN(n901) );
  AND2_X1 U907 ( .A1(n904), .A2(n879), .ZN(n883) );
  AND2_X1 U908 ( .A1(n876), .A2(n905), .ZN(n903) );
  OR2_X1 U909 ( .A1(n906), .A2(n907), .ZN(n876) );
  AND2_X1 U910 ( .A1(n908), .A2(n909), .ZN(n906) );
  AND2_X1 U911 ( .A1(n910), .A2(n859), .ZN(Result_7_) );
  AND2_X1 U912 ( .A1(n911), .A2(n912), .ZN(n910) );
  OR2_X1 U913 ( .A1(n913), .A2(n914), .ZN(n911) );
  AND2_X1 U914 ( .A1(n915), .A2(n859), .ZN(Result_6_) );
  AND2_X1 U915 ( .A1(n916), .A2(n917), .ZN(n915) );
  OR2_X1 U916 ( .A1(n918), .A2(n919), .ZN(n916) );
  INV_X1 U917 ( .A(n920), .ZN(n919) );
  AND2_X1 U918 ( .A1(n913), .A2(n914), .ZN(n918) );
  INV_X1 U919 ( .A(n921), .ZN(n914) );
  INV_X1 U920 ( .A(n922), .ZN(n913) );
  AND2_X1 U921 ( .A1(n859), .A2(n923), .ZN(Result_5_) );
  OR2_X1 U922 ( .A1(n924), .A2(n925), .ZN(n923) );
  AND2_X1 U923 ( .A1(n926), .A2(n917), .ZN(n925) );
  INV_X1 U924 ( .A(n927), .ZN(n924) );
  OR2_X1 U925 ( .A1(n917), .A2(n926), .ZN(n927) );
  OR2_X1 U926 ( .A1(n928), .A2(n929), .ZN(n926) );
  AND2_X1 U927 ( .A1(n930), .A2(n931), .ZN(n929) );
  INV_X1 U928 ( .A(n932), .ZN(n930) );
  AND2_X1 U929 ( .A1(n933), .A2(n932), .ZN(n928) );
  AND2_X1 U930 ( .A1(n934), .A2(n859), .ZN(Result_4_) );
  AND2_X1 U931 ( .A1(n935), .A2(n936), .ZN(n934) );
  OR2_X1 U932 ( .A1(n937), .A2(n938), .ZN(n936) );
  OR2_X1 U933 ( .A1(n939), .A2(n940), .ZN(n938) );
  AND2_X1 U934 ( .A1(n941), .A2(n942), .ZN(n940) );
  AND2_X1 U935 ( .A1(n943), .A2(n944), .ZN(n939) );
  OR2_X1 U936 ( .A1(n945), .A2(n943), .ZN(n935) );
  AND2_X1 U937 ( .A1(n946), .A2(n859), .ZN(Result_3_) );
  AND2_X1 U938 ( .A1(n947), .A2(n948), .ZN(n946) );
  INV_X1 U939 ( .A(n949), .ZN(n948) );
  AND2_X1 U940 ( .A1(n950), .A2(n951), .ZN(n949) );
  OR2_X1 U941 ( .A1(n951), .A2(n950), .ZN(n947) );
  INV_X1 U942 ( .A(n952), .ZN(n951) );
  OR2_X1 U943 ( .A1(n953), .A2(n954), .ZN(n952) );
  AND2_X1 U944 ( .A1(n955), .A2(n956), .ZN(n954) );
  OR2_X1 U945 ( .A1(n957), .A2(n958), .ZN(n956) );
  AND2_X1 U946 ( .A1(n959), .A2(n859), .ZN(Result_2_) );
  AND2_X1 U947 ( .A1(n960), .A2(n961), .ZN(n959) );
  OR2_X1 U948 ( .A1(n962), .A2(n963), .ZN(n961) );
  OR2_X1 U949 ( .A1(n964), .A2(n965), .ZN(n960) );
  INV_X1 U950 ( .A(n962), .ZN(n965) );
  OR2_X1 U951 ( .A1(n966), .A2(n967), .ZN(n962) );
  AND2_X1 U952 ( .A1(n968), .A2(n969), .ZN(n967) );
  AND2_X1 U953 ( .A1(n970), .A2(n971), .ZN(n966) );
  INV_X1 U954 ( .A(n969), .ZN(n970) );
  AND2_X1 U955 ( .A1(n972), .A2(n859), .ZN(Result_1_) );
  AND2_X1 U956 ( .A1(n973), .A2(n974), .ZN(n972) );
  OR2_X1 U957 ( .A1(n975), .A2(n976), .ZN(n974) );
  OR2_X1 U958 ( .A1(n977), .A2(n978), .ZN(n976) );
  AND2_X1 U959 ( .A1(n979), .A2(n980), .ZN(n978) );
  AND2_X1 U960 ( .A1(n981), .A2(n982), .ZN(n977) );
  OR2_X1 U961 ( .A1(n980), .A2(n983), .ZN(n973) );
  INV_X1 U962 ( .A(n981), .ZN(n980) );
  OR2_X1 U963 ( .A1(n984), .A2(n985), .ZN(Result_15_) );
  AND2_X1 U964 ( .A1(n986), .A2(n872), .ZN(n985) );
  OR2_X1 U965 ( .A1(n987), .A2(n988), .ZN(n986) );
  INV_X1 U966 ( .A(n989), .ZN(n988) );
  AND2_X1 U967 ( .A1(b_7_), .A2(n990), .ZN(n987) );
  AND2_X1 U968 ( .A1(n991), .A2(n859), .ZN(n984) );
  OR2_X1 U969 ( .A1(n992), .A2(n993), .ZN(Result_14_) );
  AND2_X1 U970 ( .A1(n994), .A2(n859), .ZN(n993) );
  OR2_X1 U971 ( .A1(n995), .A2(n996), .ZN(n994) );
  INV_X1 U972 ( .A(n997), .ZN(n996) );
  OR2_X1 U973 ( .A1(n998), .A2(n999), .ZN(n997) );
  AND2_X1 U974 ( .A1(n999), .A2(n998), .ZN(n995) );
  OR2_X1 U975 ( .A1(n1000), .A2(n1001), .ZN(n998) );
  AND2_X1 U976 ( .A1(n1002), .A2(n872), .ZN(n992) );
  OR2_X1 U977 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
  OR2_X1 U978 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
  AND2_X1 U979 ( .A1(n1007), .A2(b_6_), .ZN(n1006) );
  AND2_X1 U980 ( .A1(n1008), .A2(n1000), .ZN(n1007) );
  AND2_X1 U981 ( .A1(n1009), .A2(n1010), .ZN(n1005) );
  OR2_X1 U982 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
  AND2_X1 U983 ( .A1(n991), .A2(n1000), .ZN(n1012) );
  AND2_X1 U984 ( .A1(a_6_), .A2(n1008), .ZN(n1011) );
  OR2_X1 U985 ( .A1(n1013), .A2(n1014), .ZN(Result_13_) );
  AND2_X1 U986 ( .A1(n1015), .A2(n859), .ZN(n1014) );
  OR2_X1 U987 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
  AND2_X1 U988 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
  INV_X1 U989 ( .A(n1020), .ZN(n1016) );
  OR2_X1 U990 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  OR2_X1 U991 ( .A1(n1021), .A2(n1022), .ZN(n1018) );
  INV_X1 U992 ( .A(n1023), .ZN(n1022) );
  OR2_X1 U993 ( .A1(n1024), .A2(n1003), .ZN(n1023) );
  AND2_X1 U994 ( .A1(n1003), .A2(n1024), .ZN(n1021) );
  INV_X1 U995 ( .A(n1025), .ZN(n1003) );
  AND2_X1 U996 ( .A1(n1026), .A2(n872), .ZN(n1013) );
  OR2_X1 U997 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
  AND2_X1 U998 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
  OR2_X1 U999 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
  AND2_X1 U1000 ( .A1(n1033), .A2(n1034), .ZN(n1027) );
  OR2_X1 U1001 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
  AND2_X1 U1002 ( .A1(a_5_), .A2(n1037), .ZN(n1036) );
  OR2_X1 U1003 ( .A1(n1038), .A2(n1039), .ZN(Result_12_) );
  AND2_X1 U1004 ( .A1(n1040), .A2(n859), .ZN(n1039) );
  OR2_X1 U1005 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
  AND2_X1 U1006 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
  INV_X1 U1007 ( .A(n1045), .ZN(n1041) );
  OR2_X1 U1008 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  OR2_X1 U1009 ( .A1(n1046), .A2(n1047), .ZN(n1043) );
  AND2_X1 U1010 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
  INV_X1 U1011 ( .A(n1050), .ZN(n1046) );
  OR2_X1 U1012 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  INV_X1 U1013 ( .A(n1051), .ZN(n1048) );
  AND2_X1 U1014 ( .A1(n1052), .A2(n872), .ZN(n1038) );
  OR2_X1 U1015 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
  AND2_X1 U1016 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
  INV_X1 U1017 ( .A(n1057), .ZN(n1055) );
  AND2_X1 U1018 ( .A1(n1058), .A2(n1057), .ZN(n1053) );
  OR2_X1 U1019 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
  INV_X1 U1020 ( .A(n1056), .ZN(n1058) );
  OR2_X1 U1021 ( .A1(n1061), .A2(n1062), .ZN(Result_11_) );
  AND2_X1 U1022 ( .A1(n1063), .A2(n859), .ZN(n1062) );
  AND2_X1 U1023 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
  INV_X1 U1024 ( .A(n1066), .ZN(n1065) );
  AND2_X1 U1025 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
  OR2_X1 U1026 ( .A1(n1068), .A2(n1067), .ZN(n1064) );
  AND2_X1 U1027 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
  INV_X1 U1028 ( .A(n1071), .ZN(n1070) );
  AND2_X1 U1029 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
  OR2_X1 U1030 ( .A1(n1073), .A2(n1072), .ZN(n1069) );
  INV_X1 U1031 ( .A(n1074), .ZN(n1072) );
  AND2_X1 U1032 ( .A1(n1075), .A2(n872), .ZN(n1061) );
  OR2_X1 U1033 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
  OR2_X1 U1034 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
  AND2_X1 U1035 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
  AND2_X1 U1036 ( .A1(n1082), .A2(n1083), .ZN(n1078) );
  AND2_X1 U1037 ( .A1(n1084), .A2(n1085), .ZN(n1076) );
  OR2_X1 U1038 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
  AND2_X1 U1039 ( .A1(n1080), .A2(n1088), .ZN(n1087) );
  INV_X1 U1040 ( .A(n1083), .ZN(n1080) );
  AND2_X1 U1041 ( .A1(a_3_), .A2(n1083), .ZN(n1086) );
  OR2_X1 U1042 ( .A1(n1089), .A2(n1090), .ZN(Result_10_) );
  AND2_X1 U1043 ( .A1(n1091), .A2(n859), .ZN(n1090) );
  OR2_X1 U1044 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
  AND2_X1 U1045 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
  INV_X1 U1046 ( .A(n1096), .ZN(n1092) );
  OR2_X1 U1047 ( .A1(n1095), .A2(n1094), .ZN(n1096) );
  OR2_X1 U1048 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
  AND2_X1 U1049 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
  INV_X1 U1050 ( .A(n1101), .ZN(n1097) );
  OR2_X1 U1051 ( .A1(n1100), .A2(n1099), .ZN(n1101) );
  INV_X1 U1052 ( .A(n1102), .ZN(n1099) );
  AND2_X1 U1053 ( .A1(n1103), .A2(n872), .ZN(n1089) );
  OR2_X1 U1054 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
  AND2_X1 U1055 ( .A1(n1106), .A2(n908), .ZN(n1105) );
  INV_X1 U1056 ( .A(n1107), .ZN(n1106) );
  AND2_X1 U1057 ( .A1(n1108), .A2(n1107), .ZN(n1104) );
  OR2_X1 U1058 ( .A1(n907), .A2(n1109), .ZN(n1107) );
  AND2_X1 U1059 ( .A1(n1110), .A2(n1111), .ZN(n907) );
  INV_X1 U1060 ( .A(n908), .ZN(n1108) );
  OR2_X1 U1061 ( .A1(n1112), .A2(n1113), .ZN(n908) );
  AND2_X1 U1062 ( .A1(n1088), .A2(n1085), .ZN(n1113) );
  AND2_X1 U1063 ( .A1(n1083), .A2(n1114), .ZN(n1112) );
  OR2_X1 U1064 ( .A1(n1115), .A2(n1059), .ZN(n1083) );
  AND2_X1 U1065 ( .A1(n1116), .A2(n1117), .ZN(n1059) );
  AND2_X1 U1066 ( .A1(n1056), .A2(n1118), .ZN(n1115) );
  OR2_X1 U1067 ( .A1(n1119), .A2(n1032), .ZN(n1056) );
  AND2_X1 U1068 ( .A1(n1120), .A2(n1037), .ZN(n1032) );
  AND2_X1 U1069 ( .A1(n1033), .A2(n1121), .ZN(n1119) );
  INV_X1 U1070 ( .A(n1030), .ZN(n1033) );
  OR2_X1 U1071 ( .A1(n1122), .A2(n1123), .ZN(n1030) );
  OR2_X1 U1072 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
  AND2_X1 U1073 ( .A1(b_7_), .A2(n999), .ZN(n1125) );
  AND2_X1 U1074 ( .A1(n991), .A2(a_6_), .ZN(n1122) );
  INV_X1 U1075 ( .A(n1008), .ZN(n991) );
  OR2_X1 U1076 ( .A1(n990), .A2(n1001), .ZN(n1008) );
  AND2_X1 U1077 ( .A1(n859), .A2(n1126), .ZN(Result_0_) );
  OR2_X1 U1078 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
  AND2_X1 U1079 ( .A1(n981), .A2(n1129), .ZN(n1128) );
  OR2_X1 U1080 ( .A1(n975), .A2(n979), .ZN(n1129) );
  INV_X1 U1081 ( .A(n983), .ZN(n975) );
  OR2_X1 U1082 ( .A1(n1130), .A2(n969), .ZN(n983) );
  OR2_X1 U1083 ( .A1(n979), .A2(n1131), .ZN(n969) );
  AND2_X1 U1084 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
  INV_X1 U1085 ( .A(n982), .ZN(n979) );
  OR2_X1 U1086 ( .A1(n1132), .A2(n1133), .ZN(n982) );
  AND2_X1 U1087 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
  OR2_X1 U1088 ( .A1(n1111), .A2(n1136), .ZN(n1134) );
  AND2_X1 U1089 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
  INV_X1 U1090 ( .A(n1139), .ZN(n1138) );
  OR2_X1 U1091 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
  AND2_X1 U1092 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
  AND2_X1 U1093 ( .A1(b_0_), .A2(n1144), .ZN(n1140) );
  OR2_X1 U1094 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
  AND2_X1 U1095 ( .A1(a_1_), .A2(n1147), .ZN(n1146) );
  AND2_X1 U1096 ( .A1(n882), .A2(a_2_), .ZN(n1145) );
  AND2_X1 U1097 ( .A1(n968), .A2(n963), .ZN(n1130) );
  INV_X1 U1098 ( .A(n971), .ZN(n968) );
  OR2_X1 U1099 ( .A1(n953), .A2(n1148), .ZN(n971) );
  AND2_X1 U1100 ( .A1(n1149), .A2(n950), .ZN(n1148) );
  OR2_X1 U1101 ( .A1(n1150), .A2(n1151), .ZN(n950) );
  AND2_X1 U1102 ( .A1(n944), .A2(n941), .ZN(n1151) );
  AND2_X1 U1103 ( .A1(n937), .A2(n941), .ZN(n1150) );
  INV_X1 U1104 ( .A(n943), .ZN(n941) );
  AND2_X1 U1105 ( .A1(n1152), .A2(n1153), .ZN(n943) );
  OR2_X1 U1106 ( .A1(n957), .A2(n1154), .ZN(n1153) );
  INV_X1 U1107 ( .A(n1155), .ZN(n957) );
  OR2_X1 U1108 ( .A1(n1155), .A2(n958), .ZN(n1152) );
  INV_X1 U1109 ( .A(n945), .ZN(n937) );
  OR2_X1 U1110 ( .A1(n1156), .A2(n932), .ZN(n945) );
  OR2_X1 U1111 ( .A1(n944), .A2(n1157), .ZN(n932) );
  AND2_X1 U1112 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
  INV_X1 U1113 ( .A(n942), .ZN(n944) );
  OR2_X1 U1114 ( .A1(n1158), .A2(n1159), .ZN(n942) );
  OR2_X1 U1115 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
  AND2_X1 U1116 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
  AND2_X1 U1117 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
  OR2_X1 U1118 ( .A1(n1163), .A2(n1162), .ZN(n1164) );
  AND2_X1 U1119 ( .A1(n1166), .A2(n1167), .ZN(n1158) );
  OR2_X1 U1120 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
  OR2_X1 U1121 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
  INV_X1 U1122 ( .A(n1169), .ZN(n1170) );
  AND2_X1 U1123 ( .A1(n1172), .A2(n1173), .ZN(n1169) );
  OR2_X1 U1124 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
  INV_X1 U1125 ( .A(n1176), .ZN(n1175) );
  OR2_X1 U1126 ( .A1(n1176), .A2(n1177), .ZN(n1172) );
  AND2_X1 U1127 ( .A1(n917), .A2(n931), .ZN(n1156) );
  OR2_X1 U1128 ( .A1(n920), .A2(n912), .ZN(n917) );
  OR2_X1 U1129 ( .A1(n922), .A2(n921), .ZN(n912) );
  OR2_X1 U1130 ( .A1(n1178), .A2(n1179), .ZN(n921) );
  INV_X1 U1131 ( .A(n1180), .ZN(n1179) );
  OR2_X1 U1132 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
  AND2_X1 U1133 ( .A1(n1182), .A2(n1181), .ZN(n1178) );
  AND2_X1 U1134 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
  OR2_X1 U1135 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
  INV_X1 U1136 ( .A(n1187), .ZN(n1186) );
  OR2_X1 U1137 ( .A1(n1187), .A2(n1188), .ZN(n1183) );
  INV_X1 U1138 ( .A(n1185), .ZN(n1188) );
  OR2_X1 U1139 ( .A1(n1189), .A2(n1190), .ZN(n922) );
  AND2_X1 U1140 ( .A1(n1191), .A2(n895), .ZN(n1190) );
  AND2_X1 U1141 ( .A1(n890), .A2(n1192), .ZN(n1189) );
  OR2_X1 U1142 ( .A1(n895), .A2(n1191), .ZN(n1192) );
  INV_X1 U1143 ( .A(n894), .ZN(n1191) );
  AND2_X1 U1144 ( .A1(a_0_), .A2(b_7_), .ZN(n894) );
  OR2_X1 U1145 ( .A1(n1193), .A2(n1194), .ZN(n895) );
  AND2_X1 U1146 ( .A1(n867), .A2(n869), .ZN(n1194) );
  AND2_X1 U1147 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
  OR2_X1 U1148 ( .A1(n869), .A2(n867), .ZN(n1196) );
  OR2_X1 U1149 ( .A1(n904), .A2(n1001), .ZN(n867) );
  OR2_X1 U1150 ( .A1(n1197), .A2(n1198), .ZN(n869) );
  AND2_X1 U1151 ( .A1(n1102), .A2(n1100), .ZN(n1198) );
  AND2_X1 U1152 ( .A1(n1095), .A2(n1199), .ZN(n1197) );
  OR2_X1 U1153 ( .A1(n1102), .A2(n1100), .ZN(n1199) );
  OR2_X1 U1154 ( .A1(n1110), .A2(n1001), .ZN(n1100) );
  OR2_X1 U1155 ( .A1(n1200), .A2(n1201), .ZN(n1102) );
  AND2_X1 U1156 ( .A1(n1074), .A2(n1073), .ZN(n1201) );
  AND2_X1 U1157 ( .A1(n1068), .A2(n1202), .ZN(n1200) );
  OR2_X1 U1158 ( .A1(n1074), .A2(n1073), .ZN(n1202) );
  OR2_X1 U1159 ( .A1(n1088), .A2(n1001), .ZN(n1073) );
  OR2_X1 U1160 ( .A1(n1203), .A2(n1204), .ZN(n1074) );
  AND2_X1 U1161 ( .A1(n1051), .A2(n1049), .ZN(n1204) );
  AND2_X1 U1162 ( .A1(n1044), .A2(n1205), .ZN(n1203) );
  OR2_X1 U1163 ( .A1(n1051), .A2(n1049), .ZN(n1205) );
  OR2_X1 U1164 ( .A1(n1116), .A2(n1001), .ZN(n1049) );
  OR2_X1 U1165 ( .A1(n1206), .A2(n1207), .ZN(n1051) );
  AND2_X1 U1166 ( .A1(n1024), .A2(n1025), .ZN(n1207) );
  AND2_X1 U1167 ( .A1(n1019), .A2(n1208), .ZN(n1206) );
  OR2_X1 U1168 ( .A1(n1024), .A2(n1025), .ZN(n1208) );
  OR2_X1 U1169 ( .A1(n1001), .A2(n1209), .ZN(n1025) );
  OR2_X1 U1170 ( .A1(n1000), .A2(n1210), .ZN(n1209) );
  INV_X1 U1171 ( .A(n999), .ZN(n1210) );
  OR2_X1 U1172 ( .A1(n1120), .A2(n1001), .ZN(n1024) );
  INV_X1 U1173 ( .A(b_7_), .ZN(n1001) );
  AND2_X1 U1174 ( .A1(n1211), .A2(n1212), .ZN(n1019) );
  OR2_X1 U1175 ( .A1(n1213), .A2(n1124), .ZN(n1212) );
  INV_X1 U1176 ( .A(n1214), .ZN(n1211) );
  AND2_X1 U1177 ( .A1(n1124), .A2(n1213), .ZN(n1214) );
  OR2_X1 U1178 ( .A1(n990), .A2(n1037), .ZN(n1213) );
  AND2_X1 U1179 ( .A1(a_6_), .A2(b_6_), .ZN(n1124) );
  AND2_X1 U1180 ( .A1(n1215), .A2(n1216), .ZN(n1044) );
  INV_X1 U1181 ( .A(n1217), .ZN(n1216) );
  AND2_X1 U1182 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
  OR2_X1 U1183 ( .A1(n1219), .A2(n1218), .ZN(n1215) );
  OR2_X1 U1184 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
  INV_X1 U1185 ( .A(n1222), .ZN(n1221) );
  OR2_X1 U1186 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
  AND2_X1 U1187 ( .A1(n1224), .A2(n1223), .ZN(n1220) );
  OR2_X1 U1188 ( .A1(n1225), .A2(n1226), .ZN(n1068) );
  INV_X1 U1189 ( .A(n1227), .ZN(n1226) );
  OR2_X1 U1190 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
  AND2_X1 U1191 ( .A1(n1229), .A2(n1228), .ZN(n1225) );
  AND2_X1 U1192 ( .A1(n1230), .A2(n1231), .ZN(n1228) );
  INV_X1 U1193 ( .A(n1232), .ZN(n1231) );
  AND2_X1 U1194 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
  OR2_X1 U1195 ( .A1(n1234), .A2(n1233), .ZN(n1230) );
  INV_X1 U1196 ( .A(n1235), .ZN(n1233) );
  AND2_X1 U1197 ( .A1(n1236), .A2(n1237), .ZN(n1095) );
  INV_X1 U1198 ( .A(n1238), .ZN(n1237) );
  AND2_X1 U1199 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
  OR2_X1 U1200 ( .A1(n1240), .A2(n1239), .ZN(n1236) );
  OR2_X1 U1201 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
  AND2_X1 U1202 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
  INV_X1 U1203 ( .A(n1245), .ZN(n1241) );
  OR2_X1 U1204 ( .A1(n1244), .A2(n1243), .ZN(n1245) );
  INV_X1 U1205 ( .A(n1246), .ZN(n1243) );
  INV_X1 U1206 ( .A(n864), .ZN(n1195) );
  OR2_X1 U1207 ( .A1(n1247), .A2(n1248), .ZN(n864) );
  AND2_X1 U1208 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
  INV_X1 U1209 ( .A(n1251), .ZN(n1247) );
  OR2_X1 U1210 ( .A1(n1250), .A2(n1249), .ZN(n1251) );
  OR2_X1 U1211 ( .A1(n1252), .A2(n1253), .ZN(n1249) );
  AND2_X1 U1212 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
  INV_X1 U1213 ( .A(n1256), .ZN(n1254) );
  AND2_X1 U1214 ( .A1(n1257), .A2(n1256), .ZN(n1252) );
  INV_X1 U1215 ( .A(n1255), .ZN(n1257) );
  AND2_X1 U1216 ( .A1(n1258), .A2(n1259), .ZN(n890) );
  INV_X1 U1217 ( .A(n1260), .ZN(n1259) );
  AND2_X1 U1218 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
  OR2_X1 U1219 ( .A1(n1262), .A2(n1261), .ZN(n1258) );
  OR2_X1 U1220 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
  AND2_X1 U1221 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
  INV_X1 U1222 ( .A(n1267), .ZN(n1265) );
  AND2_X1 U1223 ( .A1(n1268), .A2(n1267), .ZN(n1263) );
  INV_X1 U1224 ( .A(n1266), .ZN(n1268) );
  OR2_X1 U1225 ( .A1(n933), .A2(n1269), .ZN(n920) );
  AND2_X1 U1226 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
  INV_X1 U1227 ( .A(n931), .ZN(n933) );
  OR2_X1 U1228 ( .A1(n1270), .A2(n1271), .ZN(n931) );
  OR2_X1 U1229 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
  AND2_X1 U1230 ( .A1(n1185), .A2(n1187), .ZN(n1273) );
  AND2_X1 U1231 ( .A1(n1182), .A2(n1274), .ZN(n1272) );
  OR2_X1 U1232 ( .A1(n1187), .A2(n1185), .ZN(n1274) );
  OR2_X1 U1233 ( .A1(n1010), .A2(n1275), .ZN(n1185) );
  OR2_X1 U1234 ( .A1(n1276), .A2(n1277), .ZN(n1187) );
  AND2_X1 U1235 ( .A1(n1267), .A2(n1266), .ZN(n1277) );
  AND2_X1 U1236 ( .A1(n1262), .A2(n1278), .ZN(n1276) );
  OR2_X1 U1237 ( .A1(n1266), .A2(n1267), .ZN(n1278) );
  OR2_X1 U1238 ( .A1(n1010), .A2(n904), .ZN(n1267) );
  OR2_X1 U1239 ( .A1(n1279), .A2(n1280), .ZN(n1266) );
  AND2_X1 U1240 ( .A1(n1256), .A2(n1255), .ZN(n1280) );
  AND2_X1 U1241 ( .A1(n1250), .A2(n1281), .ZN(n1279) );
  OR2_X1 U1242 ( .A1(n1255), .A2(n1256), .ZN(n1281) );
  OR2_X1 U1243 ( .A1(n1010), .A2(n1110), .ZN(n1256) );
  OR2_X1 U1244 ( .A1(n1282), .A2(n1283), .ZN(n1255) );
  AND2_X1 U1245 ( .A1(n1246), .A2(n1244), .ZN(n1283) );
  AND2_X1 U1246 ( .A1(n1240), .A2(n1284), .ZN(n1282) );
  OR2_X1 U1247 ( .A1(n1246), .A2(n1244), .ZN(n1284) );
  OR2_X1 U1248 ( .A1(n1010), .A2(n1088), .ZN(n1244) );
  OR2_X1 U1249 ( .A1(n1285), .A2(n1286), .ZN(n1246) );
  AND2_X1 U1250 ( .A1(n1235), .A2(n1234), .ZN(n1286) );
  AND2_X1 U1251 ( .A1(n1229), .A2(n1287), .ZN(n1285) );
  OR2_X1 U1252 ( .A1(n1235), .A2(n1234), .ZN(n1287) );
  OR2_X1 U1253 ( .A1(n1010), .A2(n1116), .ZN(n1234) );
  OR2_X1 U1254 ( .A1(n1288), .A2(n1289), .ZN(n1235) );
  AND2_X1 U1255 ( .A1(n1223), .A2(n1290), .ZN(n1289) );
  AND2_X1 U1256 ( .A1(n1219), .A2(n1291), .ZN(n1288) );
  OR2_X1 U1257 ( .A1(n1223), .A2(n1290), .ZN(n1291) );
  INV_X1 U1258 ( .A(n1224), .ZN(n1290) );
  AND2_X1 U1259 ( .A1(n1292), .A2(n999), .ZN(n1224) );
  AND2_X1 U1260 ( .A1(a_7_), .A2(b_6_), .ZN(n999) );
  OR2_X1 U1261 ( .A1(n1010), .A2(n1120), .ZN(n1223) );
  INV_X1 U1262 ( .A(b_6_), .ZN(n1010) );
  AND2_X1 U1263 ( .A1(n1293), .A2(n1294), .ZN(n1219) );
  OR2_X1 U1264 ( .A1(n1295), .A2(n1292), .ZN(n1294) );
  INV_X1 U1265 ( .A(n1296), .ZN(n1292) );
  OR2_X1 U1266 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
  OR2_X1 U1267 ( .A1(n1298), .A2(n1299), .ZN(n1229) );
  AND2_X1 U1268 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
  INV_X1 U1269 ( .A(n1302), .ZN(n1298) );
  OR2_X1 U1270 ( .A1(n1300), .A2(n1301), .ZN(n1302) );
  OR2_X1 U1271 ( .A1(n1303), .A2(n1304), .ZN(n1300) );
  AND2_X1 U1272 ( .A1(n1031), .A2(n1305), .ZN(n1304) );
  INV_X1 U1273 ( .A(n1121), .ZN(n1031) );
  AND2_X1 U1274 ( .A1(n1306), .A2(n1121), .ZN(n1303) );
  AND2_X1 U1275 ( .A1(n1307), .A2(n1308), .ZN(n1240) );
  INV_X1 U1276 ( .A(n1309), .ZN(n1308) );
  AND2_X1 U1277 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
  OR2_X1 U1278 ( .A1(n1311), .A2(n1310), .ZN(n1307) );
  OR2_X1 U1279 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
  AND2_X1 U1280 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
  INV_X1 U1281 ( .A(n1316), .ZN(n1312) );
  OR2_X1 U1282 ( .A1(n1315), .A2(n1314), .ZN(n1316) );
  INV_X1 U1283 ( .A(n1317), .ZN(n1314) );
  AND2_X1 U1284 ( .A1(n1318), .A2(n1319), .ZN(n1250) );
  INV_X1 U1285 ( .A(n1320), .ZN(n1319) );
  AND2_X1 U1286 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
  OR2_X1 U1287 ( .A1(n1322), .A2(n1321), .ZN(n1318) );
  OR2_X1 U1288 ( .A1(n1323), .A2(n1324), .ZN(n1321) );
  AND2_X1 U1289 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
  INV_X1 U1290 ( .A(n1327), .ZN(n1325) );
  AND2_X1 U1291 ( .A1(n1328), .A2(n1327), .ZN(n1323) );
  INV_X1 U1292 ( .A(n1326), .ZN(n1328) );
  AND2_X1 U1293 ( .A1(n1329), .A2(n1330), .ZN(n1262) );
  INV_X1 U1294 ( .A(n1331), .ZN(n1330) );
  AND2_X1 U1295 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
  OR2_X1 U1296 ( .A1(n1333), .A2(n1332), .ZN(n1329) );
  OR2_X1 U1297 ( .A1(n1334), .A2(n1335), .ZN(n1332) );
  AND2_X1 U1298 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
  INV_X1 U1299 ( .A(n1338), .ZN(n1336) );
  AND2_X1 U1300 ( .A1(n1339), .A2(n1338), .ZN(n1334) );
  INV_X1 U1301 ( .A(n1337), .ZN(n1339) );
  OR2_X1 U1302 ( .A1(n1340), .A2(n1341), .ZN(n1182) );
  INV_X1 U1303 ( .A(n1342), .ZN(n1341) );
  OR2_X1 U1304 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
  AND2_X1 U1305 ( .A1(n1344), .A2(n1343), .ZN(n1340) );
  AND2_X1 U1306 ( .A1(n1345), .A2(n1346), .ZN(n1343) );
  OR2_X1 U1307 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
  INV_X1 U1308 ( .A(n1349), .ZN(n1348) );
  OR2_X1 U1309 ( .A1(n1349), .A2(n1350), .ZN(n1345) );
  INV_X1 U1310 ( .A(n1347), .ZN(n1350) );
  OR2_X1 U1311 ( .A1(n1351), .A2(n1352), .ZN(n1270) );
  INV_X1 U1312 ( .A(n1353), .ZN(n1352) );
  OR2_X1 U1313 ( .A1(n1354), .A2(n1162), .ZN(n1353) );
  AND2_X1 U1314 ( .A1(n1162), .A2(n1354), .ZN(n1351) );
  AND2_X1 U1315 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
  OR2_X1 U1316 ( .A1(n1163), .A2(n1357), .ZN(n1356) );
  INV_X1 U1317 ( .A(n1165), .ZN(n1357) );
  OR2_X1 U1318 ( .A1(n1165), .A2(n1358), .ZN(n1355) );
  INV_X1 U1319 ( .A(n1163), .ZN(n1358) );
  OR2_X1 U1320 ( .A1(n1037), .A2(n1275), .ZN(n1163) );
  OR2_X1 U1321 ( .A1(n1359), .A2(n1360), .ZN(n1165) );
  AND2_X1 U1322 ( .A1(n1347), .A2(n1349), .ZN(n1360) );
  AND2_X1 U1323 ( .A1(n1344), .A2(n1361), .ZN(n1359) );
  OR2_X1 U1324 ( .A1(n1349), .A2(n1347), .ZN(n1361) );
  OR2_X1 U1325 ( .A1(n1037), .A2(n904), .ZN(n1347) );
  OR2_X1 U1326 ( .A1(n1362), .A2(n1363), .ZN(n1349) );
  AND2_X1 U1327 ( .A1(n1338), .A2(n1337), .ZN(n1363) );
  AND2_X1 U1328 ( .A1(n1333), .A2(n1364), .ZN(n1362) );
  OR2_X1 U1329 ( .A1(n1337), .A2(n1338), .ZN(n1364) );
  OR2_X1 U1330 ( .A1(n1037), .A2(n1110), .ZN(n1338) );
  OR2_X1 U1331 ( .A1(n1365), .A2(n1366), .ZN(n1337) );
  AND2_X1 U1332 ( .A1(n1327), .A2(n1326), .ZN(n1366) );
  AND2_X1 U1333 ( .A1(n1322), .A2(n1367), .ZN(n1365) );
  OR2_X1 U1334 ( .A1(n1326), .A2(n1327), .ZN(n1367) );
  OR2_X1 U1335 ( .A1(n1037), .A2(n1088), .ZN(n1327) );
  OR2_X1 U1336 ( .A1(n1368), .A2(n1369), .ZN(n1326) );
  AND2_X1 U1337 ( .A1(n1317), .A2(n1315), .ZN(n1369) );
  AND2_X1 U1338 ( .A1(n1311), .A2(n1370), .ZN(n1368) );
  OR2_X1 U1339 ( .A1(n1317), .A2(n1315), .ZN(n1370) );
  OR2_X1 U1340 ( .A1(n1037), .A2(n1116), .ZN(n1315) );
  OR2_X1 U1341 ( .A1(n1371), .A2(n1372), .ZN(n1317) );
  AND2_X1 U1342 ( .A1(n1301), .A2(n1121), .ZN(n1372) );
  AND2_X1 U1343 ( .A1(n1306), .A2(n1373), .ZN(n1371) );
  OR2_X1 U1344 ( .A1(n1301), .A2(n1121), .ZN(n1373) );
  OR2_X1 U1345 ( .A1(n1037), .A2(n1120), .ZN(n1121) );
  OR2_X1 U1346 ( .A1(n1295), .A2(n1296), .ZN(n1301) );
  OR2_X1 U1347 ( .A1(n1000), .A2(n1037), .ZN(n1296) );
  INV_X1 U1348 ( .A(b_5_), .ZN(n1037) );
  INV_X1 U1349 ( .A(n1297), .ZN(n1295) );
  INV_X1 U1350 ( .A(n1305), .ZN(n1306) );
  OR2_X1 U1351 ( .A1(n1374), .A2(n1375), .ZN(n1305) );
  AND2_X1 U1352 ( .A1(n1376), .A2(b_3_), .ZN(n1375) );
  AND2_X1 U1353 ( .A1(a_7_), .A2(n1377), .ZN(n1376) );
  OR2_X1 U1354 ( .A1(n1000), .A2(n1117), .ZN(n1377) );
  AND2_X1 U1355 ( .A1(n1378), .A2(b_4_), .ZN(n1374) );
  AND2_X1 U1356 ( .A1(a_6_), .A2(n1379), .ZN(n1378) );
  OR2_X1 U1357 ( .A1(n990), .A2(n1085), .ZN(n1379) );
  AND2_X1 U1358 ( .A1(n1380), .A2(n1381), .ZN(n1311) );
  OR2_X1 U1359 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
  INV_X1 U1360 ( .A(n1384), .ZN(n1382) );
  OR2_X1 U1361 ( .A1(n1385), .A2(n1384), .ZN(n1380) );
  OR2_X1 U1362 ( .A1(n1386), .A2(n1387), .ZN(n1384) );
  AND2_X1 U1363 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
  INV_X1 U1364 ( .A(n1390), .ZN(n1386) );
  OR2_X1 U1365 ( .A1(n1389), .A2(n1388), .ZN(n1390) );
  AND2_X1 U1366 ( .A1(n1391), .A2(n1392), .ZN(n1322) );
  INV_X1 U1367 ( .A(n1393), .ZN(n1392) );
  AND2_X1 U1368 ( .A1(n1394), .A2(n1395), .ZN(n1393) );
  OR2_X1 U1369 ( .A1(n1395), .A2(n1394), .ZN(n1391) );
  OR2_X1 U1370 ( .A1(n1396), .A2(n1397), .ZN(n1394) );
  AND2_X1 U1371 ( .A1(n1398), .A2(n1118), .ZN(n1397) );
  INV_X1 U1372 ( .A(n1399), .ZN(n1398) );
  AND2_X1 U1373 ( .A1(n1060), .A2(n1399), .ZN(n1396) );
  AND2_X1 U1374 ( .A1(n1400), .A2(n1401), .ZN(n1333) );
  INV_X1 U1375 ( .A(n1402), .ZN(n1401) );
  AND2_X1 U1376 ( .A1(n1403), .A2(n1404), .ZN(n1402) );
  OR2_X1 U1377 ( .A1(n1404), .A2(n1403), .ZN(n1400) );
  OR2_X1 U1378 ( .A1(n1405), .A2(n1406), .ZN(n1403) );
  AND2_X1 U1379 ( .A1(n1407), .A2(n1408), .ZN(n1406) );
  INV_X1 U1380 ( .A(n1409), .ZN(n1407) );
  AND2_X1 U1381 ( .A1(n1410), .A2(n1409), .ZN(n1405) );
  INV_X1 U1382 ( .A(n1408), .ZN(n1410) );
  OR2_X1 U1383 ( .A1(n1411), .A2(n1412), .ZN(n1344) );
  INV_X1 U1384 ( .A(n1413), .ZN(n1412) );
  OR2_X1 U1385 ( .A1(n1414), .A2(n1415), .ZN(n1413) );
  AND2_X1 U1386 ( .A1(n1415), .A2(n1414), .ZN(n1411) );
  AND2_X1 U1387 ( .A1(n1416), .A2(n1417), .ZN(n1414) );
  OR2_X1 U1388 ( .A1(n1418), .A2(n1419), .ZN(n1417) );
  INV_X1 U1389 ( .A(n1420), .ZN(n1419) );
  OR2_X1 U1390 ( .A1(n1420), .A2(n1421), .ZN(n1416) );
  INV_X1 U1391 ( .A(n1418), .ZN(n1421) );
  OR2_X1 U1392 ( .A1(n1422), .A2(n1423), .ZN(n1162) );
  INV_X1 U1393 ( .A(n1424), .ZN(n1423) );
  OR2_X1 U1394 ( .A1(n1425), .A2(n1426), .ZN(n1424) );
  AND2_X1 U1395 ( .A1(n1426), .A2(n1425), .ZN(n1422) );
  AND2_X1 U1396 ( .A1(n1427), .A2(n1428), .ZN(n1425) );
  OR2_X1 U1397 ( .A1(n1429), .A2(n1430), .ZN(n1428) );
  INV_X1 U1398 ( .A(n1431), .ZN(n1430) );
  OR2_X1 U1399 ( .A1(n1431), .A2(n1432), .ZN(n1427) );
  INV_X1 U1400 ( .A(n1429), .ZN(n1432) );
  AND2_X1 U1401 ( .A1(n1149), .A2(n1433), .ZN(n953) );
  AND2_X1 U1402 ( .A1(n1155), .A2(n1154), .ZN(n1433) );
  INV_X1 U1403 ( .A(n958), .ZN(n1154) );
  OR2_X1 U1404 ( .A1(n1434), .A2(n1435), .ZN(n958) );
  AND2_X1 U1405 ( .A1(n1174), .A2(n1176), .ZN(n1435) );
  AND2_X1 U1406 ( .A1(n1171), .A2(n1436), .ZN(n1434) );
  OR2_X1 U1407 ( .A1(n1176), .A2(n1174), .ZN(n1436) );
  INV_X1 U1408 ( .A(n1177), .ZN(n1174) );
  AND2_X1 U1409 ( .A1(b_4_), .A2(a_0_), .ZN(n1177) );
  OR2_X1 U1410 ( .A1(n1437), .A2(n1438), .ZN(n1176) );
  AND2_X1 U1411 ( .A1(n1426), .A2(n1429), .ZN(n1438) );
  AND2_X1 U1412 ( .A1(n1439), .A2(n1431), .ZN(n1437) );
  OR2_X1 U1413 ( .A1(n1440), .A2(n1441), .ZN(n1431) );
  AND2_X1 U1414 ( .A1(n1418), .A2(n1420), .ZN(n1441) );
  AND2_X1 U1415 ( .A1(n1415), .A2(n1442), .ZN(n1440) );
  OR2_X1 U1416 ( .A1(n1420), .A2(n1418), .ZN(n1442) );
  OR2_X1 U1417 ( .A1(n1117), .A2(n1110), .ZN(n1418) );
  OR2_X1 U1418 ( .A1(n1443), .A2(n1444), .ZN(n1420) );
  AND2_X1 U1419 ( .A1(n1409), .A2(n1408), .ZN(n1444) );
  AND2_X1 U1420 ( .A1(n1404), .A2(n1445), .ZN(n1443) );
  OR2_X1 U1421 ( .A1(n1408), .A2(n1409), .ZN(n1445) );
  OR2_X1 U1422 ( .A1(n1117), .A2(n1088), .ZN(n1409) );
  OR2_X1 U1423 ( .A1(n1446), .A2(n1447), .ZN(n1408) );
  AND2_X1 U1424 ( .A1(n1399), .A2(n1118), .ZN(n1447) );
  AND2_X1 U1425 ( .A1(n1395), .A2(n1448), .ZN(n1446) );
  OR2_X1 U1426 ( .A1(n1118), .A2(n1399), .ZN(n1448) );
  OR2_X1 U1427 ( .A1(n1449), .A2(n1450), .ZN(n1399) );
  AND2_X1 U1428 ( .A1(n1451), .A2(n1389), .ZN(n1450) );
  AND2_X1 U1429 ( .A1(n1385), .A2(n1452), .ZN(n1449) );
  OR2_X1 U1430 ( .A1(n1451), .A2(n1389), .ZN(n1452) );
  OR2_X1 U1431 ( .A1(n1120), .A2(n1117), .ZN(n1389) );
  INV_X1 U1432 ( .A(n1388), .ZN(n1451) );
  AND2_X1 U1433 ( .A1(n1453), .A2(n1297), .ZN(n1388) );
  AND2_X1 U1434 ( .A1(a_7_), .A2(b_4_), .ZN(n1297) );
  INV_X1 U1435 ( .A(n1383), .ZN(n1385) );
  OR2_X1 U1436 ( .A1(n1454), .A2(n1455), .ZN(n1383) );
  AND2_X1 U1437 ( .A1(n1456), .A2(n1457), .ZN(n1455) );
  AND2_X1 U1438 ( .A1(b_2_), .A2(a_7_), .ZN(n1456) );
  AND2_X1 U1439 ( .A1(n1453), .A2(n1458), .ZN(n1454) );
  INV_X1 U1440 ( .A(n1457), .ZN(n1453) );
  INV_X1 U1441 ( .A(n1060), .ZN(n1118) );
  AND2_X1 U1442 ( .A1(a_4_), .A2(b_4_), .ZN(n1060) );
  AND2_X1 U1443 ( .A1(n1459), .A2(n1460), .ZN(n1395) );
  INV_X1 U1444 ( .A(n1461), .ZN(n1460) );
  AND2_X1 U1445 ( .A1(n1462), .A2(n1463), .ZN(n1461) );
  OR2_X1 U1446 ( .A1(n1463), .A2(n1462), .ZN(n1459) );
  OR2_X1 U1447 ( .A1(n1464), .A2(n1465), .ZN(n1462) );
  AND2_X1 U1448 ( .A1(n1466), .A2(n1467), .ZN(n1465) );
  INV_X1 U1449 ( .A(n1468), .ZN(n1464) );
  OR2_X1 U1450 ( .A1(n1467), .A2(n1466), .ZN(n1468) );
  INV_X1 U1451 ( .A(n1469), .ZN(n1466) );
  AND2_X1 U1452 ( .A1(n1470), .A2(n1471), .ZN(n1404) );
  INV_X1 U1453 ( .A(n1472), .ZN(n1471) );
  AND2_X1 U1454 ( .A1(n1473), .A2(n1474), .ZN(n1472) );
  OR2_X1 U1455 ( .A1(n1474), .A2(n1473), .ZN(n1470) );
  OR2_X1 U1456 ( .A1(n1475), .A2(n1476), .ZN(n1473) );
  AND2_X1 U1457 ( .A1(n1477), .A2(n1478), .ZN(n1476) );
  INV_X1 U1458 ( .A(n1479), .ZN(n1477) );
  AND2_X1 U1459 ( .A1(n1480), .A2(n1479), .ZN(n1475) );
  INV_X1 U1460 ( .A(n1478), .ZN(n1480) );
  OR2_X1 U1461 ( .A1(n1481), .A2(n1482), .ZN(n1415) );
  INV_X1 U1462 ( .A(n1483), .ZN(n1482) );
  OR2_X1 U1463 ( .A1(n1484), .A2(n1485), .ZN(n1483) );
  AND2_X1 U1464 ( .A1(n1485), .A2(n1484), .ZN(n1481) );
  AND2_X1 U1465 ( .A1(n1486), .A2(n1487), .ZN(n1484) );
  OR2_X1 U1466 ( .A1(n1488), .A2(n1081), .ZN(n1487) );
  INV_X1 U1467 ( .A(n1114), .ZN(n1081) );
  OR2_X1 U1468 ( .A1(n1114), .A2(n1489), .ZN(n1486) );
  INV_X1 U1469 ( .A(n1488), .ZN(n1489) );
  OR2_X1 U1470 ( .A1(n1429), .A2(n1426), .ZN(n1439) );
  OR2_X1 U1471 ( .A1(n1490), .A2(n1491), .ZN(n1426) );
  INV_X1 U1472 ( .A(n1492), .ZN(n1491) );
  OR2_X1 U1473 ( .A1(n1493), .A2(n1494), .ZN(n1492) );
  AND2_X1 U1474 ( .A1(n1494), .A2(n1493), .ZN(n1490) );
  AND2_X1 U1475 ( .A1(n1495), .A2(n1496), .ZN(n1493) );
  OR2_X1 U1476 ( .A1(n1497), .A2(n1498), .ZN(n1496) );
  INV_X1 U1477 ( .A(n1499), .ZN(n1498) );
  OR2_X1 U1478 ( .A1(n1499), .A2(n1500), .ZN(n1495) );
  INV_X1 U1479 ( .A(n1497), .ZN(n1500) );
  OR2_X1 U1480 ( .A1(n1117), .A2(n904), .ZN(n1429) );
  INV_X1 U1481 ( .A(b_4_), .ZN(n1117) );
  INV_X1 U1482 ( .A(n1168), .ZN(n1171) );
  OR2_X1 U1483 ( .A1(n1501), .A2(n1502), .ZN(n1168) );
  AND2_X1 U1484 ( .A1(n1503), .A2(n1504), .ZN(n1502) );
  INV_X1 U1485 ( .A(n1505), .ZN(n1501) );
  OR2_X1 U1486 ( .A1(n1504), .A2(n1503), .ZN(n1505) );
  OR2_X1 U1487 ( .A1(n1506), .A2(n1507), .ZN(n1503) );
  AND2_X1 U1488 ( .A1(n1508), .A2(n1509), .ZN(n1507) );
  INV_X1 U1489 ( .A(n1510), .ZN(n1506) );
  OR2_X1 U1490 ( .A1(n1509), .A2(n1508), .ZN(n1510) );
  INV_X1 U1491 ( .A(n1511), .ZN(n1508) );
  OR2_X1 U1492 ( .A1(n1512), .A2(n1513), .ZN(n1155) );
  AND2_X1 U1493 ( .A1(n1514), .A2(n1515), .ZN(n1513) );
  INV_X1 U1494 ( .A(n1516), .ZN(n1512) );
  OR2_X1 U1495 ( .A1(n1515), .A2(n1514), .ZN(n1516) );
  OR2_X1 U1496 ( .A1(n1517), .A2(n1518), .ZN(n1514) );
  AND2_X1 U1497 ( .A1(n1519), .A2(n1520), .ZN(n1518) );
  INV_X1 U1498 ( .A(n1521), .ZN(n1517) );
  OR2_X1 U1499 ( .A1(n1520), .A2(n1519), .ZN(n1521) );
  INV_X1 U1500 ( .A(n1522), .ZN(n1519) );
  INV_X1 U1501 ( .A(n955), .ZN(n1149) );
  OR2_X1 U1502 ( .A1(n1523), .A2(n964), .ZN(n955) );
  INV_X1 U1503 ( .A(n963), .ZN(n964) );
  OR2_X1 U1504 ( .A1(n1524), .A2(n1525), .ZN(n963) );
  AND2_X1 U1505 ( .A1(n1524), .A2(n1525), .ZN(n1523) );
  OR2_X1 U1506 ( .A1(n1526), .A2(n1527), .ZN(n1525) );
  AND2_X1 U1507 ( .A1(n1522), .A2(n1520), .ZN(n1527) );
  AND2_X1 U1508 ( .A1(n1515), .A2(n1528), .ZN(n1526) );
  OR2_X1 U1509 ( .A1(n1520), .A2(n1522), .ZN(n1528) );
  OR2_X1 U1510 ( .A1(n1529), .A2(n1530), .ZN(n1522) );
  AND2_X1 U1511 ( .A1(n1511), .A2(n1509), .ZN(n1530) );
  AND2_X1 U1512 ( .A1(n1504), .A2(n1531), .ZN(n1529) );
  OR2_X1 U1513 ( .A1(n1509), .A2(n1511), .ZN(n1531) );
  OR2_X1 U1514 ( .A1(n1532), .A2(n1533), .ZN(n1511) );
  AND2_X1 U1515 ( .A1(n1497), .A2(n1499), .ZN(n1533) );
  AND2_X1 U1516 ( .A1(n1494), .A2(n1534), .ZN(n1532) );
  OR2_X1 U1517 ( .A1(n1499), .A2(n1497), .ZN(n1534) );
  OR2_X1 U1518 ( .A1(n1085), .A2(n1110), .ZN(n1497) );
  OR2_X1 U1519 ( .A1(n1535), .A2(n1536), .ZN(n1499) );
  AND2_X1 U1520 ( .A1(n1488), .A2(n1114), .ZN(n1536) );
  AND2_X1 U1521 ( .A1(n1485), .A2(n1537), .ZN(n1535) );
  OR2_X1 U1522 ( .A1(n1114), .A2(n1488), .ZN(n1537) );
  OR2_X1 U1523 ( .A1(n1538), .A2(n1539), .ZN(n1488) );
  AND2_X1 U1524 ( .A1(n1479), .A2(n1478), .ZN(n1539) );
  AND2_X1 U1525 ( .A1(n1474), .A2(n1540), .ZN(n1538) );
  OR2_X1 U1526 ( .A1(n1478), .A2(n1479), .ZN(n1540) );
  OR2_X1 U1527 ( .A1(n1116), .A2(n1085), .ZN(n1479) );
  OR2_X1 U1528 ( .A1(n1541), .A2(n1542), .ZN(n1478) );
  AND2_X1 U1529 ( .A1(n1469), .A2(n1467), .ZN(n1542) );
  AND2_X1 U1530 ( .A1(n1463), .A2(n1543), .ZN(n1541) );
  OR2_X1 U1531 ( .A1(n1467), .A2(n1469), .ZN(n1543) );
  OR2_X1 U1532 ( .A1(n1457), .A2(n1458), .ZN(n1469) );
  OR2_X1 U1533 ( .A1(n990), .A2(n1111), .ZN(n1458) );
  OR2_X1 U1534 ( .A1(n1000), .A2(n1085), .ZN(n1457) );
  OR2_X1 U1535 ( .A1(n1120), .A2(n1085), .ZN(n1467) );
  AND2_X1 U1536 ( .A1(n1544), .A2(n1545), .ZN(n1463) );
  OR2_X1 U1537 ( .A1(n1546), .A2(n1547), .ZN(n1545) );
  INV_X1 U1538 ( .A(n1548), .ZN(n1547) );
  OR2_X1 U1539 ( .A1(n1548), .A2(n1549), .ZN(n1544) );
  AND2_X1 U1540 ( .A1(n1550), .A2(n1551), .ZN(n1474) );
  INV_X1 U1541 ( .A(n1552), .ZN(n1551) );
  AND2_X1 U1542 ( .A1(n1553), .A2(n1554), .ZN(n1552) );
  OR2_X1 U1543 ( .A1(n1554), .A2(n1553), .ZN(n1550) );
  OR2_X1 U1544 ( .A1(n1555), .A2(n1556), .ZN(n1553) );
  AND2_X1 U1545 ( .A1(n1557), .A2(n1558), .ZN(n1556) );
  INV_X1 U1546 ( .A(n1559), .ZN(n1555) );
  OR2_X1 U1547 ( .A1(n1558), .A2(n1557), .ZN(n1559) );
  OR2_X1 U1548 ( .A1(n1085), .A2(n1088), .ZN(n1114) );
  OR2_X1 U1549 ( .A1(n1560), .A2(n1561), .ZN(n1485) );
  INV_X1 U1550 ( .A(n1562), .ZN(n1561) );
  OR2_X1 U1551 ( .A1(n1563), .A2(n1564), .ZN(n1562) );
  AND2_X1 U1552 ( .A1(n1564), .A2(n1563), .ZN(n1560) );
  AND2_X1 U1553 ( .A1(n1565), .A2(n1566), .ZN(n1563) );
  OR2_X1 U1554 ( .A1(n1567), .A2(n1568), .ZN(n1566) );
  INV_X1 U1555 ( .A(n1569), .ZN(n1568) );
  OR2_X1 U1556 ( .A1(n1569), .A2(n1570), .ZN(n1565) );
  INV_X1 U1557 ( .A(n1567), .ZN(n1570) );
  OR2_X1 U1558 ( .A1(n1571), .A2(n1572), .ZN(n1494) );
  INV_X1 U1559 ( .A(n1573), .ZN(n1572) );
  OR2_X1 U1560 ( .A1(n1574), .A2(n1575), .ZN(n1573) );
  AND2_X1 U1561 ( .A1(n1575), .A2(n1574), .ZN(n1571) );
  AND2_X1 U1562 ( .A1(n1576), .A2(n1577), .ZN(n1574) );
  OR2_X1 U1563 ( .A1(n1578), .A2(n1579), .ZN(n1577) );
  INV_X1 U1564 ( .A(n1580), .ZN(n1579) );
  OR2_X1 U1565 ( .A1(n1580), .A2(n1581), .ZN(n1576) );
  INV_X1 U1566 ( .A(n1578), .ZN(n1581) );
  OR2_X1 U1567 ( .A1(n1085), .A2(n904), .ZN(n1509) );
  AND2_X1 U1568 ( .A1(n1582), .A2(n1583), .ZN(n1504) );
  INV_X1 U1569 ( .A(n1584), .ZN(n1583) );
  AND2_X1 U1570 ( .A1(n1585), .A2(n1586), .ZN(n1584) );
  OR2_X1 U1571 ( .A1(n1586), .A2(n1585), .ZN(n1582) );
  OR2_X1 U1572 ( .A1(n1587), .A2(n1588), .ZN(n1585) );
  AND2_X1 U1573 ( .A1(n1589), .A2(n909), .ZN(n1588) );
  INV_X1 U1574 ( .A(n1590), .ZN(n1589) );
  AND2_X1 U1575 ( .A1(n1109), .A2(n1590), .ZN(n1587) );
  INV_X1 U1576 ( .A(n909), .ZN(n1109) );
  OR2_X1 U1577 ( .A1(n1085), .A2(n1275), .ZN(n1520) );
  INV_X1 U1578 ( .A(b_3_), .ZN(n1085) );
  AND2_X1 U1579 ( .A1(n1591), .A2(n1592), .ZN(n1515) );
  INV_X1 U1580 ( .A(n1593), .ZN(n1592) );
  AND2_X1 U1581 ( .A1(n1594), .A2(n1595), .ZN(n1593) );
  OR2_X1 U1582 ( .A1(n1595), .A2(n1594), .ZN(n1591) );
  OR2_X1 U1583 ( .A1(n1596), .A2(n1597), .ZN(n1594) );
  AND2_X1 U1584 ( .A1(n1598), .A2(n1599), .ZN(n1597) );
  INV_X1 U1585 ( .A(n1600), .ZN(n1598) );
  AND2_X1 U1586 ( .A1(n1601), .A2(n1600), .ZN(n1596) );
  INV_X1 U1587 ( .A(n1599), .ZN(n1601) );
  AND2_X1 U1588 ( .A1(n1602), .A2(n1603), .ZN(n1524) );
  INV_X1 U1589 ( .A(n1604), .ZN(n1603) );
  AND2_X1 U1590 ( .A1(n1605), .A2(n1136), .ZN(n1604) );
  OR2_X1 U1591 ( .A1(n1136), .A2(n1605), .ZN(n1602) );
  OR2_X1 U1592 ( .A1(n1606), .A2(n1607), .ZN(n1605) );
  AND2_X1 U1593 ( .A1(n1608), .A2(n1135), .ZN(n1607) );
  INV_X1 U1594 ( .A(n1609), .ZN(n1606) );
  OR2_X1 U1595 ( .A1(n1135), .A2(n1608), .ZN(n1609) );
  AND2_X1 U1596 ( .A1(b_2_), .A2(a_0_), .ZN(n1608) );
  OR2_X1 U1597 ( .A1(n1610), .A2(n1611), .ZN(n1135) );
  AND2_X1 U1598 ( .A1(n1600), .A2(n1599), .ZN(n1611) );
  AND2_X1 U1599 ( .A1(n1595), .A2(n1612), .ZN(n1610) );
  OR2_X1 U1600 ( .A1(n1599), .A2(n1600), .ZN(n1612) );
  OR2_X1 U1601 ( .A1(n1111), .A2(n904), .ZN(n1600) );
  OR2_X1 U1602 ( .A1(n1613), .A2(n1614), .ZN(n1599) );
  AND2_X1 U1603 ( .A1(n1590), .A2(n909), .ZN(n1614) );
  AND2_X1 U1604 ( .A1(n1586), .A2(n1615), .ZN(n1613) );
  OR2_X1 U1605 ( .A1(n909), .A2(n1590), .ZN(n1615) );
  OR2_X1 U1606 ( .A1(n1616), .A2(n1617), .ZN(n1590) );
  AND2_X1 U1607 ( .A1(n1578), .A2(n1580), .ZN(n1617) );
  AND2_X1 U1608 ( .A1(n1575), .A2(n1618), .ZN(n1616) );
  OR2_X1 U1609 ( .A1(n1580), .A2(n1578), .ZN(n1618) );
  OR2_X1 U1610 ( .A1(n1088), .A2(n1111), .ZN(n1578) );
  OR2_X1 U1611 ( .A1(n1619), .A2(n1620), .ZN(n1580) );
  AND2_X1 U1612 ( .A1(n1567), .A2(n1569), .ZN(n1620) );
  AND2_X1 U1613 ( .A1(n1564), .A2(n1621), .ZN(n1619) );
  OR2_X1 U1614 ( .A1(n1569), .A2(n1567), .ZN(n1621) );
  OR2_X1 U1615 ( .A1(n1116), .A2(n1111), .ZN(n1567) );
  OR2_X1 U1616 ( .A1(n1622), .A2(n1623), .ZN(n1569) );
  AND2_X1 U1617 ( .A1(n1624), .A2(n1558), .ZN(n1623) );
  AND2_X1 U1618 ( .A1(n1554), .A2(n1625), .ZN(n1622) );
  OR2_X1 U1619 ( .A1(n1558), .A2(n1624), .ZN(n1625) );
  INV_X1 U1620 ( .A(n1557), .ZN(n1624) );
  AND2_X1 U1621 ( .A1(a_5_), .A2(b_2_), .ZN(n1557) );
  OR2_X1 U1622 ( .A1(n1548), .A2(n1546), .ZN(n1558) );
  INV_X1 U1623 ( .A(n1549), .ZN(n1546) );
  AND2_X1 U1624 ( .A1(a_6_), .A2(b_2_), .ZN(n1549) );
  OR2_X1 U1625 ( .A1(n990), .A2(n879), .ZN(n1548) );
  AND2_X1 U1626 ( .A1(n1626), .A2(n1627), .ZN(n1554) );
  OR2_X1 U1627 ( .A1(n1628), .A2(n1629), .ZN(n1627) );
  INV_X1 U1628 ( .A(n1630), .ZN(n1626) );
  AND2_X1 U1629 ( .A1(n1629), .A2(n1628), .ZN(n1630) );
  OR2_X1 U1630 ( .A1(n1631), .A2(n1632), .ZN(n1564) );
  INV_X1 U1631 ( .A(n1633), .ZN(n1632) );
  OR2_X1 U1632 ( .A1(n1634), .A2(n1635), .ZN(n1633) );
  AND2_X1 U1633 ( .A1(n1635), .A2(n1634), .ZN(n1631) );
  OR2_X1 U1634 ( .A1(n1636), .A2(n1637), .ZN(n1634) );
  AND2_X1 U1635 ( .A1(n1638), .A2(b_0_), .ZN(n1637) );
  AND2_X1 U1636 ( .A1(a_6_), .A2(n1639), .ZN(n1638) );
  OR2_X1 U1637 ( .A1(n1120), .A2(n879), .ZN(n1639) );
  AND2_X1 U1638 ( .A1(n1640), .A2(b_1_), .ZN(n1636) );
  AND2_X1 U1639 ( .A1(a_5_), .A2(n1641), .ZN(n1640) );
  OR2_X1 U1640 ( .A1(n1000), .A2(n1143), .ZN(n1641) );
  OR2_X1 U1641 ( .A1(n1642), .A2(n1643), .ZN(n1575) );
  AND2_X1 U1642 ( .A1(n1644), .A2(n1645), .ZN(n1643) );
  INV_X1 U1643 ( .A(n1646), .ZN(n1642) );
  OR2_X1 U1644 ( .A1(n1644), .A2(n1645), .ZN(n1646) );
  OR2_X1 U1645 ( .A1(n1647), .A2(n1648), .ZN(n1644) );
  AND2_X1 U1646 ( .A1(n1649), .A2(n1650), .ZN(n1648) );
  AND2_X1 U1647 ( .A1(n1651), .A2(n1652), .ZN(n1647) );
  OR2_X1 U1648 ( .A1(n1110), .A2(n1111), .ZN(n909) );
  INV_X1 U1649 ( .A(b_2_), .ZN(n1111) );
  AND2_X1 U1650 ( .A1(n1653), .A2(n1654), .ZN(n1586) );
  INV_X1 U1651 ( .A(n1655), .ZN(n1654) );
  AND2_X1 U1652 ( .A1(n1656), .A2(n1657), .ZN(n1655) );
  OR2_X1 U1653 ( .A1(n1656), .A2(n1657), .ZN(n1653) );
  OR2_X1 U1654 ( .A1(n1658), .A2(n1659), .ZN(n1656) );
  INV_X1 U1655 ( .A(n1660), .ZN(n1659) );
  OR2_X1 U1656 ( .A1(n1661), .A2(n1662), .ZN(n1660) );
  AND2_X1 U1657 ( .A1(n1662), .A2(n1661), .ZN(n1658) );
  AND2_X1 U1658 ( .A1(n1663), .A2(n1664), .ZN(n1595) );
  INV_X1 U1659 ( .A(n1665), .ZN(n1664) );
  AND2_X1 U1660 ( .A1(n1666), .A2(n1667), .ZN(n1665) );
  OR2_X1 U1661 ( .A1(n1666), .A2(n1667), .ZN(n1663) );
  OR2_X1 U1662 ( .A1(n1668), .A2(n1669), .ZN(n1666) );
  INV_X1 U1663 ( .A(n1670), .ZN(n1669) );
  OR2_X1 U1664 ( .A1(n1671), .A2(n1672), .ZN(n1670) );
  AND2_X1 U1665 ( .A1(n1672), .A2(n1671), .ZN(n1668) );
  AND2_X1 U1666 ( .A1(n1673), .A2(n1674), .ZN(n1136) );
  INV_X1 U1667 ( .A(n1675), .ZN(n1674) );
  AND2_X1 U1668 ( .A1(n1676), .A2(n1677), .ZN(n1675) );
  OR2_X1 U1669 ( .A1(n1677), .A2(n1676), .ZN(n1673) );
  AND2_X1 U1670 ( .A1(n1137), .A2(n882), .ZN(n1676) );
  INV_X1 U1671 ( .A(n905), .ZN(n882) );
  OR2_X1 U1672 ( .A1(n879), .A2(n904), .ZN(n905) );
  OR2_X1 U1673 ( .A1(n1678), .A2(n1679), .ZN(n1137) );
  AND2_X1 U1674 ( .A1(n1667), .A2(n1671), .ZN(n1679) );
  AND2_X1 U1675 ( .A1(n1680), .A2(n1681), .ZN(n1678) );
  INV_X1 U1676 ( .A(n1672), .ZN(n1681) );
  AND2_X1 U1677 ( .A1(a_3_), .A2(b_0_), .ZN(n1672) );
  OR2_X1 U1678 ( .A1(n1671), .A2(n1667), .ZN(n1680) );
  OR2_X1 U1679 ( .A1(n1110), .A2(n879), .ZN(n1667) );
  OR2_X1 U1680 ( .A1(n1682), .A2(n1683), .ZN(n1671) );
  AND2_X1 U1681 ( .A1(n1657), .A2(n1661), .ZN(n1683) );
  AND2_X1 U1682 ( .A1(n1684), .A2(n1685), .ZN(n1682) );
  INV_X1 U1683 ( .A(n1662), .ZN(n1685) );
  AND2_X1 U1684 ( .A1(a_3_), .A2(b_1_), .ZN(n1662) );
  OR2_X1 U1685 ( .A1(n1661), .A2(n1657), .ZN(n1684) );
  OR2_X1 U1686 ( .A1(n1116), .A2(n1143), .ZN(n1657) );
  OR2_X1 U1687 ( .A1(n1686), .A2(n1687), .ZN(n1661) );
  AND2_X1 U1688 ( .A1(n1645), .A2(n1650), .ZN(n1687) );
  AND2_X1 U1689 ( .A1(n1649), .A2(n1688), .ZN(n1686) );
  OR2_X1 U1690 ( .A1(n1650), .A2(n1645), .ZN(n1688) );
  OR2_X1 U1691 ( .A1(n1116), .A2(n879), .ZN(n1645) );
  INV_X1 U1692 ( .A(b_1_), .ZN(n879) );
  INV_X1 U1693 ( .A(n1652), .ZN(n1649) );
  OR2_X1 U1694 ( .A1(n1689), .A2(n1635), .ZN(n1652) );
  AND2_X1 U1695 ( .A1(n1629), .A2(n1690), .ZN(n1635) );
  INV_X1 U1696 ( .A(n1628), .ZN(n1690) );
  OR2_X1 U1697 ( .A1(n990), .A2(n1143), .ZN(n1628) );
  AND2_X1 U1698 ( .A1(n1651), .A2(n1629), .ZN(n1689) );
  AND2_X1 U1699 ( .A1(a_6_), .A2(b_1_), .ZN(n1629) );
  INV_X1 U1700 ( .A(n1650), .ZN(n1651) );
  OR2_X1 U1701 ( .A1(n1120), .A2(n1143), .ZN(n1650) );
  OR2_X1 U1702 ( .A1(n1110), .A2(n1143), .ZN(n1677) );
  INV_X1 U1703 ( .A(b_0_), .ZN(n1143) );
  AND2_X1 U1704 ( .A1(n1147), .A2(b_0_), .ZN(n981) );
  INV_X1 U1705 ( .A(n1142), .ZN(n1147) );
  AND2_X1 U1706 ( .A1(n1142), .A2(b_0_), .ZN(n1127) );
  AND2_X1 U1707 ( .A1(b_1_), .A2(a_0_), .ZN(n1142) );
  INV_X1 U1708 ( .A(n872), .ZN(n859) );
  OR2_X1 U1709 ( .A1(n1691), .A2(n902), .ZN(n872) );
  AND2_X1 U1710 ( .A1(n1275), .A2(b_0_), .ZN(n902) );
  AND2_X1 U1711 ( .A1(n1692), .A2(n1693), .ZN(n1691) );
  OR2_X1 U1712 ( .A1(b_0_), .A2(n1275), .ZN(n1693) );
  INV_X1 U1713 ( .A(a_0_), .ZN(n1275) );
  AND2_X1 U1714 ( .A1(n1694), .A2(n1695), .ZN(n1692) );
  OR2_X1 U1715 ( .A1(n877), .A2(n1696), .ZN(n1695) );
  OR2_X1 U1716 ( .A1(n1697), .A2(n1698), .ZN(n1696) );
  AND2_X1 U1717 ( .A1(b_2_), .A2(n1110), .ZN(n1698) );
  AND2_X1 U1718 ( .A1(n1699), .A2(n1700), .ZN(n1697) );
  OR2_X1 U1719 ( .A1(b_3_), .A2(n1088), .ZN(n1700) );
  AND2_X1 U1720 ( .A1(n1701), .A2(n1702), .ZN(n1699) );
  OR2_X1 U1721 ( .A1(n1082), .A2(n1703), .ZN(n1702) );
  OR2_X1 U1722 ( .A1(n1704), .A2(n1705), .ZN(n1703) );
  AND2_X1 U1723 ( .A1(b_4_), .A2(n1116), .ZN(n1705) );
  AND2_X1 U1724 ( .A1(n1706), .A2(n1707), .ZN(n1704) );
  OR2_X1 U1725 ( .A1(b_5_), .A2(n1120), .ZN(n1707) );
  AND2_X1 U1726 ( .A1(n1708), .A2(n1709), .ZN(n1706) );
  OR2_X1 U1727 ( .A1(n1710), .A2(n1711), .ZN(n1709) );
  OR2_X1 U1728 ( .A1(n1712), .A2(n1035), .ZN(n1711) );
  AND2_X1 U1729 ( .A1(n1120), .A2(b_5_), .ZN(n1035) );
  INV_X1 U1730 ( .A(a_5_), .ZN(n1120) );
  AND2_X1 U1731 ( .A1(b_6_), .A2(n1713), .ZN(n1712) );
  OR2_X1 U1732 ( .A1(n989), .A2(n1000), .ZN(n1713) );
  AND2_X1 U1733 ( .A1(n1000), .A2(n989), .ZN(n1710) );
  OR2_X1 U1734 ( .A1(b_7_), .A2(n990), .ZN(n989) );
  INV_X1 U1735 ( .A(a_7_), .ZN(n990) );
  INV_X1 U1736 ( .A(a_6_), .ZN(n1000) );
  OR2_X1 U1737 ( .A1(b_4_), .A2(n1116), .ZN(n1708) );
  INV_X1 U1738 ( .A(a_4_), .ZN(n1116) );
  AND2_X1 U1739 ( .A1(n1088), .A2(b_3_), .ZN(n1082) );
  INV_X1 U1740 ( .A(a_3_), .ZN(n1088) );
  OR2_X1 U1741 ( .A1(b_2_), .A2(n1110), .ZN(n1701) );
  INV_X1 U1742 ( .A(a_2_), .ZN(n1110) );
  AND2_X1 U1743 ( .A1(n904), .A2(b_1_), .ZN(n877) );
  OR2_X1 U1744 ( .A1(b_1_), .A2(n904), .ZN(n1694) );
  INV_X1 U1745 ( .A(a_1_), .ZN(n904) );
endmodule

