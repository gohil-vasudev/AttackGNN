module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n552_, new_n342_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n234_, new_n532_, new_n472_, new_n393_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n606_, new_n589_, new_n248_, new_n350_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n397_, new_n399_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n598_, new_n143_, new_n520_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n151_, new_n513_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n417_, new_n591_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n440_, new_n531_, new_n593_, new_n252_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n217_, new_n269_, new_n512_, new_n599_, new_n412_, new_n607_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n567_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n405_;

not g000 ( new_n138_, keyIn_0_41 );
xnor g001 ( new_n139_, N89, N93 );
xnor g002 ( new_n140_, N81, N85 );
xnor g003 ( new_n141_, new_n139_, new_n140_ );
xor g004 ( new_n142_, N65, N69 );
not g005 ( new_n143_, new_n142_ );
not g006 ( new_n144_, keyIn_0_6 );
not g007 ( new_n145_, N73 );
not g008 ( new_n146_, N77 );
nand g009 ( new_n147_, new_n145_, new_n146_ );
nand g010 ( new_n148_, N73, N77 );
nand g011 ( new_n149_, new_n147_, new_n148_ );
nand g012 ( new_n150_, new_n149_, new_n144_ );
nand g013 ( new_n151_, new_n147_, keyIn_0_6, new_n148_ );
nand g014 ( new_n152_, new_n150_, new_n151_ );
xnor g015 ( new_n153_, new_n152_, keyIn_0_5 );
xnor g016 ( new_n154_, new_n153_, new_n143_ );
xnor g017 ( new_n155_, new_n154_, new_n141_ );
nand g018 ( new_n156_, N129, N137 );
xnor g019 ( new_n157_, new_n155_, new_n156_ );
xnor g020 ( new_n158_, N1, N17 );
xnor g021 ( new_n159_, N33, N49 );
xnor g022 ( new_n160_, new_n158_, new_n159_ );
nand g023 ( new_n161_, new_n157_, new_n160_ );
not g024 ( new_n162_, new_n156_ );
xnor g025 ( new_n163_, new_n155_, new_n162_ );
not g026 ( new_n164_, new_n160_ );
nand g027 ( new_n165_, new_n163_, new_n164_ );
nand g028 ( new_n166_, new_n161_, new_n165_ );
not g029 ( new_n167_, keyIn_0_19 );
not g030 ( new_n168_, N121 );
not g031 ( new_n169_, N125 );
nand g032 ( new_n170_, new_n168_, new_n169_ );
nand g033 ( new_n171_, N121, N125 );
nand g034 ( new_n172_, new_n170_, new_n171_ );
nand g035 ( new_n173_, new_n172_, keyIn_0_7 );
not g036 ( new_n174_, keyIn_0_7 );
nand g037 ( new_n175_, new_n170_, new_n174_, new_n171_ );
nand g038 ( new_n176_, new_n173_, new_n175_ );
xor g039 ( new_n177_, N113, N117 );
xnor g040 ( new_n178_, new_n176_, new_n177_ );
xnor g041 ( new_n179_, new_n178_, new_n167_ );
xor g042 ( new_n180_, N97, N101 );
xnor g043 ( new_n181_, N105, N109 );
xnor g044 ( new_n182_, new_n180_, new_n181_ );
xor g045 ( new_n183_, new_n182_, keyIn_0_18 );
nand g046 ( new_n184_, new_n179_, new_n183_ );
xnor g047 ( new_n185_, new_n178_, keyIn_0_19 );
not g048 ( new_n186_, new_n183_ );
nand g049 ( new_n187_, new_n185_, new_n186_ );
nand g050 ( new_n188_, new_n184_, new_n187_ );
nand g051 ( new_n189_, new_n188_, keyIn_0_22 );
not g052 ( new_n190_, keyIn_0_22 );
nand g053 ( new_n191_, new_n184_, new_n187_, new_n190_ );
nand g054 ( new_n192_, new_n189_, new_n191_ );
nand g055 ( new_n193_, new_n192_, keyIn_0_8 );
not g056 ( new_n194_, keyIn_0_8 );
nand g057 ( new_n195_, new_n189_, new_n194_, new_n191_ );
nand g058 ( new_n196_, new_n193_, new_n195_ );
nand g059 ( new_n197_, N130, N137 );
nand g060 ( new_n198_, new_n196_, new_n197_ );
nand g061 ( new_n199_, new_n193_, N130, N137, new_n195_ );
nand g062 ( new_n200_, new_n198_, new_n199_ );
xor g063 ( new_n201_, N5, N21 );
xnor g064 ( new_n202_, new_n201_, keyIn_0_12 );
xor g065 ( new_n203_, N37, N53 );
xnor g066 ( new_n204_, new_n203_, keyIn_0_13 );
xnor g067 ( new_n205_, new_n202_, new_n204_ );
not g068 ( new_n206_, new_n205_ );
xnor g069 ( new_n207_, new_n200_, new_n206_ );
not g070 ( new_n208_, keyIn_0_23 );
xnor g071 ( new_n209_, new_n185_, new_n141_ );
not g072 ( new_n210_, keyIn_0_9 );
nand g073 ( new_n211_, N132, N137 );
nand g074 ( new_n212_, new_n211_, new_n210_ );
nand g075 ( new_n213_, keyIn_0_9, N132, N137 );
nand g076 ( new_n214_, new_n212_, new_n213_ );
xnor g077 ( new_n215_, new_n209_, new_n214_ );
nand g078 ( new_n216_, new_n215_, new_n208_ );
not g079 ( new_n217_, new_n214_ );
xnor g080 ( new_n218_, new_n209_, new_n217_ );
nand g081 ( new_n219_, new_n218_, keyIn_0_23 );
xor g082 ( new_n220_, N45, N61 );
xor g083 ( new_n221_, N13, N29 );
xnor g084 ( new_n222_, new_n221_, keyIn_0_14 );
xnor g085 ( new_n223_, new_n222_, new_n220_ );
not g086 ( new_n224_, new_n223_ );
nand g087 ( new_n225_, new_n216_, new_n219_, new_n224_ );
nand g088 ( new_n226_, new_n216_, new_n219_ );
nand g089 ( new_n227_, new_n226_, new_n223_ );
nand g090 ( new_n228_, new_n227_, new_n225_ );
not g091 ( new_n229_, new_n166_ );
xnor g092 ( new_n230_, new_n153_, new_n142_ );
nand g093 ( new_n231_, new_n230_, new_n183_ );
nand g094 ( new_n232_, new_n154_, new_n186_ );
nand g095 ( new_n233_, new_n231_, new_n232_ );
nand g096 ( new_n234_, N131, N137 );
nand g097 ( new_n235_, new_n233_, new_n234_ );
nand g098 ( new_n236_, new_n231_, new_n232_, N131, N137 );
nand g099 ( new_n237_, new_n235_, new_n236_ );
xnor g100 ( new_n238_, N41, N57 );
xnor g101 ( new_n239_, N9, N25 );
xnor g102 ( new_n240_, new_n238_, new_n239_ );
nand g103 ( new_n241_, new_n237_, new_n240_ );
not g104 ( new_n242_, new_n240_ );
nand g105 ( new_n243_, new_n235_, new_n236_, new_n242_ );
nand g106 ( new_n244_, new_n241_, new_n243_ );
nand g107 ( new_n245_, new_n244_, keyIn_0_24 );
not g108 ( new_n246_, keyIn_0_24 );
nand g109 ( new_n247_, new_n241_, new_n246_, new_n243_ );
nand g110 ( new_n248_, new_n245_, new_n247_ );
nand g111 ( new_n249_, new_n248_, new_n229_ );
not g112 ( new_n250_, new_n249_ );
nand g113 ( new_n251_, new_n207_, new_n228_, new_n250_ );
nand g114 ( new_n252_, new_n248_, keyIn_0_26 );
not g115 ( new_n253_, keyIn_0_26 );
nand g116 ( new_n254_, new_n245_, new_n253_, new_n247_ );
not g117 ( new_n255_, new_n254_ );
nor g118 ( new_n256_, new_n228_, new_n255_ );
nand g119 ( new_n257_, new_n207_, new_n256_, new_n166_, new_n252_ );
nand g120 ( new_n258_, new_n257_, keyIn_0_36 );
not g121 ( new_n259_, new_n228_ );
nand g122 ( new_n260_, new_n198_, new_n199_, new_n206_ );
nand g123 ( new_n261_, new_n200_, new_n205_ );
nand g124 ( new_n262_, new_n261_, new_n260_ );
nand g125 ( new_n263_, new_n262_, new_n250_ );
not g126 ( new_n264_, new_n248_ );
not g127 ( new_n265_, keyIn_0_25 );
nand g128 ( new_n266_, new_n161_, new_n165_, new_n265_ );
nand g129 ( new_n267_, new_n166_, keyIn_0_25 );
nand g130 ( new_n268_, new_n267_, new_n266_ );
nand g131 ( new_n269_, new_n268_, new_n261_, new_n260_, new_n264_ );
nand g132 ( new_n270_, new_n263_, new_n269_ );
nand g133 ( new_n271_, new_n270_, new_n259_ );
not g134 ( new_n272_, keyIn_0_36 );
not g135 ( new_n273_, new_n252_ );
nor g136 ( new_n274_, new_n273_, new_n228_, new_n255_ );
nand g137 ( new_n275_, new_n274_, new_n272_, new_n166_, new_n207_ );
nand g138 ( new_n276_, new_n258_, new_n271_, new_n275_, new_n251_ );
not g139 ( new_n277_, keyIn_0_21 );
not g140 ( new_n278_, keyIn_0_3 );
xnor g141 ( new_n279_, N41, N45 );
nand g142 ( new_n280_, new_n279_, new_n278_ );
not g143 ( new_n281_, N41 );
not g144 ( new_n282_, N45 );
nand g145 ( new_n283_, new_n281_, new_n282_ );
nand g146 ( new_n284_, N41, N45 );
nand g147 ( new_n285_, new_n283_, keyIn_0_3, new_n284_ );
nand g148 ( new_n286_, new_n280_, new_n285_ );
not g149 ( new_n287_, N37 );
not g150 ( new_n288_, N33 );
nand g151 ( new_n289_, new_n288_, keyIn_0_2 );
not g152 ( new_n290_, keyIn_0_2 );
nand g153 ( new_n291_, new_n290_, N33 );
nand g154 ( new_n292_, new_n289_, new_n291_ );
nand g155 ( new_n293_, new_n292_, new_n287_ );
nand g156 ( new_n294_, new_n289_, new_n291_, N37 );
nand g157 ( new_n295_, new_n293_, new_n294_ );
nand g158 ( new_n296_, new_n295_, new_n286_ );
nand g159 ( new_n297_, new_n293_, new_n280_, new_n285_, new_n294_ );
nand g160 ( new_n298_, new_n296_, new_n297_ );
nand g161 ( new_n299_, new_n298_, keyIn_0_17 );
not g162 ( new_n300_, keyIn_0_17 );
nand g163 ( new_n301_, new_n296_, new_n300_, new_n297_ );
nand g164 ( new_n302_, new_n299_, new_n301_ );
xnor g165 ( new_n303_, N9, N13 );
xnor g166 ( new_n304_, N1, N5 );
xnor g167 ( new_n305_, new_n303_, new_n304_ );
xnor g168 ( new_n306_, new_n305_, keyIn_0_16 );
nand g169 ( new_n307_, new_n302_, new_n306_ );
not g170 ( new_n308_, keyIn_0_16 );
xnor g171 ( new_n309_, new_n305_, new_n308_ );
nand g172 ( new_n310_, new_n309_, new_n299_, new_n301_ );
nand g173 ( new_n311_, new_n307_, new_n310_ );
nand g174 ( new_n312_, new_n311_, new_n277_ );
nand g175 ( new_n313_, new_n307_, keyIn_0_21, new_n310_ );
nand g176 ( new_n314_, new_n312_, new_n313_ );
nand g177 ( new_n315_, new_n314_, keyIn_0_10 );
not g178 ( new_n316_, keyIn_0_10 );
nand g179 ( new_n317_, new_n312_, new_n316_, new_n313_ );
nand g180 ( new_n318_, new_n315_, new_n317_ );
nand g181 ( new_n319_, N135, N137 );
nand g182 ( new_n320_, new_n318_, new_n319_ );
nand g183 ( new_n321_, new_n315_, N135, N137, new_n317_ );
nand g184 ( new_n322_, new_n320_, new_n321_ );
xor g185 ( new_n323_, N73, N89 );
xnor g186 ( new_n324_, N105, N121 );
xnor g187 ( new_n325_, new_n323_, new_n324_ );
xor g188 ( new_n326_, new_n325_, keyIn_0_20 );
nand g189 ( new_n327_, new_n322_, new_n326_ );
not g190 ( new_n328_, new_n326_ );
nand g191 ( new_n329_, new_n320_, new_n321_, new_n328_ );
nand g192 ( new_n330_, new_n327_, new_n329_ );
not g193 ( new_n331_, N49 );
not g194 ( new_n332_, N53 );
nand g195 ( new_n333_, new_n331_, new_n332_ );
nand g196 ( new_n334_, N49, N53 );
nand g197 ( new_n335_, new_n333_, new_n334_ );
nand g198 ( new_n336_, new_n335_, keyIn_0_4 );
not g199 ( new_n337_, keyIn_0_4 );
nand g200 ( new_n338_, new_n333_, new_n337_, new_n334_ );
nand g201 ( new_n339_, new_n336_, new_n338_ );
xnor g202 ( new_n340_, N57, N61 );
nand g203 ( new_n341_, new_n339_, new_n340_ );
not g204 ( new_n342_, new_n340_ );
nand g205 ( new_n343_, new_n336_, new_n338_, new_n342_ );
nand g206 ( new_n344_, new_n341_, new_n343_ );
not g207 ( new_n345_, N17 );
not g208 ( new_n346_, N21 );
nand g209 ( new_n347_, new_n345_, new_n346_ );
nand g210 ( new_n348_, N17, N21 );
nand g211 ( new_n349_, new_n347_, new_n348_ );
nand g212 ( new_n350_, new_n349_, keyIn_0_0 );
not g213 ( new_n351_, keyIn_0_0 );
nand g214 ( new_n352_, new_n347_, new_n351_, new_n348_ );
nand g215 ( new_n353_, new_n350_, new_n352_ );
not g216 ( new_n354_, N25 );
not g217 ( new_n355_, N29 );
nand g218 ( new_n356_, new_n354_, new_n355_ );
nand g219 ( new_n357_, N25, N29 );
nand g220 ( new_n358_, new_n356_, new_n357_ );
nand g221 ( new_n359_, new_n358_, keyIn_0_1 );
not g222 ( new_n360_, keyIn_0_1 );
nand g223 ( new_n361_, new_n356_, new_n360_, new_n357_ );
nand g224 ( new_n362_, new_n359_, new_n361_ );
nand g225 ( new_n363_, new_n353_, new_n362_ );
nand g226 ( new_n364_, new_n350_, new_n359_, new_n352_, new_n361_ );
nand g227 ( new_n365_, new_n363_, new_n364_ );
nand g228 ( new_n366_, new_n365_, new_n344_ );
nand g229 ( new_n367_, new_n363_, new_n341_, new_n343_, new_n364_ );
nand g230 ( new_n368_, new_n366_, new_n367_ );
nand g231 ( new_n369_, new_n368_, keyIn_0_11 );
not g232 ( new_n370_, keyIn_0_11 );
nand g233 ( new_n371_, new_n366_, new_n370_, new_n367_ );
nand g234 ( new_n372_, new_n369_, new_n371_ );
nand g235 ( new_n373_, N136, N137 );
nand g236 ( new_n374_, new_n372_, new_n373_ );
nand g237 ( new_n375_, new_n369_, N136, N137, new_n371_ );
nand g238 ( new_n376_, new_n374_, new_n375_ );
xnor g239 ( new_n377_, N109, N125 );
xnor g240 ( new_n378_, N77, N93 );
xnor g241 ( new_n379_, new_n377_, new_n378_ );
not g242 ( new_n380_, new_n379_ );
nand g243 ( new_n381_, new_n376_, new_n380_ );
nand g244 ( new_n382_, new_n374_, new_n375_, new_n379_ );
nand g245 ( new_n383_, new_n381_, new_n382_ );
nand g246 ( new_n384_, new_n302_, new_n344_ );
nand g247 ( new_n385_, new_n299_, new_n301_, new_n341_, new_n343_ );
nand g248 ( new_n386_, new_n384_, new_n385_ );
nand g249 ( new_n387_, N134, N137 );
xnor g250 ( new_n388_, new_n386_, new_n387_ );
xnor g251 ( new_n389_, N101, N117 );
xnor g252 ( new_n390_, N69, N85 );
xnor g253 ( new_n391_, new_n389_, new_n390_ );
xnor g254 ( new_n392_, new_n388_, new_n391_ );
nand g255 ( new_n393_, new_n306_, new_n365_ );
nand g256 ( new_n394_, new_n309_, new_n363_, new_n364_ );
nand g257 ( new_n395_, new_n394_, new_n393_ );
nand g258 ( new_n396_, N133, N137 );
nand g259 ( new_n397_, new_n395_, new_n396_ );
nand g260 ( new_n398_, new_n394_, new_n393_, N133, N137 );
nand g261 ( new_n399_, new_n397_, new_n398_ );
xnor g262 ( new_n400_, N97, N113 );
xnor g263 ( new_n401_, new_n400_, keyIn_0_15 );
xnor g264 ( new_n402_, N65, N81 );
xnor g265 ( new_n403_, new_n401_, new_n402_ );
xnor g266 ( new_n404_, new_n399_, new_n403_ );
not g267 ( new_n405_, new_n404_ );
nor g268 ( new_n406_, new_n392_, new_n405_, new_n383_ );
nand g269 ( new_n407_, new_n276_, new_n330_, new_n406_ );
not g270 ( new_n408_, new_n407_ );
nand g271 ( new_n409_, new_n408_, new_n166_ );
xnor g272 ( new_n410_, new_n409_, new_n138_ );
xnor g273 ( N724, new_n410_, N1 );
nand g274 ( new_n412_, new_n408_, new_n262_ );
xnor g275 ( new_n413_, new_n412_, keyIn_0_42 );
xnor g276 ( N725, new_n413_, N5 );
nand g277 ( new_n415_, new_n408_, new_n264_ );
xnor g278 ( N726, new_n415_, N9 );
nand g279 ( new_n417_, new_n408_, new_n228_ );
xnor g280 ( N727, new_n417_, N13 );
nand g281 ( new_n419_, new_n276_, new_n166_ );
not g282 ( new_n420_, new_n419_ );
not g283 ( new_n421_, new_n330_ );
xor g284 ( new_n422_, new_n388_, new_n391_ );
nand g285 ( new_n423_, new_n421_, new_n383_, new_n422_, new_n404_ );
not g286 ( new_n424_, new_n423_ );
nand g287 ( new_n425_, new_n420_, new_n424_ );
xnor g288 ( new_n426_, new_n425_, N17 );
xnor g289 ( N728, new_n426_, keyIn_0_54 );
nand g290 ( new_n428_, new_n276_, new_n262_ );
not g291 ( new_n429_, new_n428_ );
nand g292 ( new_n430_, new_n429_, new_n424_ );
xnor g293 ( new_n431_, new_n430_, N21 );
xnor g294 ( N729, new_n431_, keyIn_0_55 );
nand g295 ( new_n433_, new_n276_, new_n264_ );
not g296 ( new_n434_, new_n433_ );
nand g297 ( new_n435_, new_n434_, new_n424_ );
xnor g298 ( N730, new_n435_, N25 );
nand g299 ( new_n437_, new_n276_, new_n228_, new_n424_ );
xnor g300 ( new_n438_, new_n437_, keyIn_0_43 );
xnor g301 ( N731, new_n438_, new_n355_ );
nor g302 ( new_n440_, new_n422_, new_n383_, new_n404_ );
nand g303 ( new_n441_, new_n330_, new_n440_ );
not g304 ( new_n442_, new_n441_ );
nand g305 ( new_n443_, new_n420_, new_n442_ );
xnor g306 ( new_n444_, new_n443_, N33 );
xnor g307 ( N732, new_n444_, keyIn_0_56 );
nand g308 ( new_n446_, new_n429_, new_n442_ );
xnor g309 ( new_n447_, new_n446_, new_n287_ );
xnor g310 ( N733, new_n447_, keyIn_0_57 );
nand g311 ( new_n449_, new_n434_, new_n442_ );
xnor g312 ( new_n450_, new_n449_, keyIn_0_44 );
xnor g313 ( N734, new_n450_, new_n281_ );
not g314 ( new_n452_, keyIn_0_45 );
nand g315 ( new_n453_, new_n276_, new_n228_, new_n442_ );
xnor g316 ( new_n454_, new_n453_, new_n452_ );
nand g317 ( new_n455_, new_n454_, N45 );
xnor g318 ( new_n456_, new_n453_, keyIn_0_45 );
nand g319 ( new_n457_, new_n456_, new_n282_ );
nand g320 ( new_n458_, new_n455_, new_n457_ );
nand g321 ( new_n459_, new_n458_, keyIn_0_58 );
not g322 ( new_n460_, keyIn_0_58 );
nand g323 ( new_n461_, new_n455_, new_n457_, new_n460_ );
nand g324 ( N735, new_n459_, new_n461_ );
not g325 ( new_n463_, keyIn_0_39 );
nand g326 ( new_n464_, new_n421_, keyIn_0_27 );
not g327 ( new_n465_, keyIn_0_27 );
nand g328 ( new_n466_, new_n330_, new_n465_ );
nand g329 ( new_n467_, new_n405_, new_n383_ );
not g330 ( new_n468_, new_n467_ );
nand g331 ( new_n469_, new_n464_, new_n392_, new_n466_, new_n468_ );
not g332 ( new_n470_, new_n469_ );
nand g333 ( new_n471_, new_n276_, new_n470_ );
nand g334 ( new_n472_, new_n471_, new_n463_ );
nand g335 ( new_n473_, new_n276_, keyIn_0_39, new_n470_ );
nand g336 ( new_n474_, new_n472_, new_n473_ );
nand g337 ( new_n475_, new_n474_, new_n166_ );
nand g338 ( new_n476_, new_n475_, N49 );
nand g339 ( new_n477_, new_n474_, new_n331_, new_n166_ );
nand g340 ( new_n478_, new_n476_, new_n477_ );
nand g341 ( new_n479_, new_n478_, keyIn_0_59 );
not g342 ( new_n480_, keyIn_0_59 );
nand g343 ( new_n481_, new_n476_, new_n480_, new_n477_ );
nand g344 ( N736, new_n479_, new_n481_ );
nand g345 ( new_n483_, new_n474_, new_n262_ );
nand g346 ( new_n484_, new_n483_, keyIn_0_46 );
not g347 ( new_n485_, keyIn_0_46 );
nand g348 ( new_n486_, new_n474_, new_n485_, new_n262_ );
nand g349 ( new_n487_, new_n484_, new_n486_ );
nand g350 ( new_n488_, new_n487_, N53 );
nand g351 ( new_n489_, new_n484_, new_n332_, new_n486_ );
nand g352 ( N737, new_n488_, new_n489_ );
nand g353 ( new_n491_, new_n474_, new_n264_ );
xnor g354 ( N738, new_n491_, N57 );
nand g355 ( new_n493_, new_n474_, new_n228_ );
xnor g356 ( N739, new_n493_, N61 );
not g357 ( new_n495_, N65 );
not g358 ( new_n496_, keyIn_0_37 );
not g359 ( new_n497_, keyIn_0_31 );
nand g360 ( new_n498_, new_n327_, new_n497_, new_n329_ );
nand g361 ( new_n499_, new_n330_, keyIn_0_31 );
nand g362 ( new_n500_, new_n499_, new_n496_, new_n440_, new_n498_ );
nand g363 ( new_n501_, new_n499_, new_n440_, new_n498_ );
nand g364 ( new_n502_, new_n501_, keyIn_0_37 );
not g365 ( new_n503_, keyIn_0_32 );
nand g366 ( new_n504_, new_n327_, new_n503_, new_n329_ );
nand g367 ( new_n505_, new_n330_, keyIn_0_32 );
nand g368 ( new_n506_, new_n381_, keyIn_0_33, new_n382_ );
not g369 ( new_n507_, keyIn_0_33 );
nand g370 ( new_n508_, new_n383_, new_n507_ );
nand g371 ( new_n509_, new_n422_, new_n508_, new_n404_, new_n506_ );
not g372 ( new_n510_, new_n509_ );
nand g373 ( new_n511_, new_n505_, new_n504_, new_n510_ );
xor g374 ( new_n512_, new_n383_, keyIn_0_30 );
xnor g375 ( new_n513_, new_n404_, keyIn_0_29 );
nor g376 ( new_n514_, new_n513_, new_n392_ );
nand g377 ( new_n515_, new_n330_, new_n514_, new_n512_ );
xnor g378 ( new_n516_, new_n392_, keyIn_0_28 );
nand g379 ( new_n517_, new_n516_, new_n327_, new_n329_, new_n468_ );
nand g380 ( new_n518_, new_n515_, new_n517_ );
not g381 ( new_n519_, new_n518_ );
nand g382 ( new_n520_, new_n502_, new_n519_, new_n500_, new_n511_ );
nand g383 ( new_n521_, new_n520_, keyIn_0_38 );
not g384 ( new_n522_, keyIn_0_38 );
not g385 ( new_n523_, new_n511_ );
nor g386 ( new_n524_, new_n523_, new_n518_ );
nand g387 ( new_n525_, new_n524_, new_n522_, new_n500_, new_n502_ );
nor g388 ( new_n526_, new_n262_, new_n228_, new_n229_, new_n248_ );
nand g389 ( new_n527_, new_n521_, new_n525_, new_n526_ );
nand g390 ( new_n528_, new_n527_, keyIn_0_40 );
not g391 ( new_n529_, keyIn_0_40 );
nand g392 ( new_n530_, new_n521_, new_n525_, new_n529_, new_n526_ );
nand g393 ( new_n531_, new_n528_, new_n530_ );
nand g394 ( new_n532_, new_n531_, new_n404_ );
nand g395 ( new_n533_, new_n532_, keyIn_0_47 );
not g396 ( new_n534_, keyIn_0_47 );
nand g397 ( new_n535_, new_n531_, new_n534_, new_n404_ );
nand g398 ( new_n536_, new_n533_, new_n535_ );
nand g399 ( new_n537_, new_n536_, new_n495_ );
nand g400 ( new_n538_, new_n533_, N65, new_n535_ );
nand g401 ( N740, new_n537_, new_n538_ );
not g402 ( new_n540_, N69 );
nand g403 ( new_n541_, new_n531_, new_n392_ );
nand g404 ( new_n542_, new_n541_, keyIn_0_48 );
not g405 ( new_n543_, keyIn_0_48 );
nand g406 ( new_n544_, new_n531_, new_n543_, new_n392_ );
nand g407 ( new_n545_, new_n542_, new_n544_ );
nand g408 ( new_n546_, new_n545_, new_n540_ );
nand g409 ( new_n547_, new_n542_, N69, new_n544_ );
nand g410 ( N741, new_n546_, new_n547_ );
nand g411 ( new_n549_, new_n531_, new_n330_ );
xnor g412 ( N742, new_n549_, N73 );
nand g413 ( new_n551_, new_n531_, new_n383_ );
nand g414 ( new_n552_, new_n551_, N77 );
nand g415 ( new_n553_, new_n531_, new_n146_, new_n383_ );
nand g416 ( new_n554_, new_n552_, new_n553_ );
nand g417 ( new_n555_, new_n554_, keyIn_0_60 );
not g418 ( new_n556_, keyIn_0_60 );
nand g419 ( new_n557_, new_n552_, new_n556_, new_n553_ );
nand g420 ( N743, new_n555_, new_n557_ );
xnor g421 ( new_n559_, new_n520_, new_n522_ );
nand g422 ( new_n560_, new_n262_, keyIn_0_34 );
not g423 ( new_n561_, new_n560_ );
not g424 ( new_n562_, keyIn_0_34 );
nand g425 ( new_n563_, new_n207_, new_n562_ );
not g426 ( new_n564_, new_n563_ );
nand g427 ( new_n565_, new_n228_, new_n166_, new_n248_ );
nor g428 ( new_n566_, new_n564_, new_n561_, new_n565_ );
nand g429 ( new_n567_, new_n559_, new_n566_ );
not g430 ( new_n568_, new_n567_ );
nand g431 ( new_n569_, new_n568_, new_n404_ );
xnor g432 ( N744, new_n569_, N81 );
nand g433 ( new_n571_, new_n559_, new_n392_, new_n566_ );
xnor g434 ( new_n572_, new_n571_, keyIn_0_49 );
xnor g435 ( N745, new_n572_, N85 );
nand g436 ( new_n574_, new_n559_, new_n330_, new_n566_ );
xnor g437 ( new_n575_, new_n574_, N89 );
xnor g438 ( N746, new_n575_, keyIn_0_61 );
nand g439 ( new_n577_, new_n568_, new_n383_ );
xnor g440 ( N747, new_n577_, N93 );
xnor g441 ( new_n579_, new_n166_, keyIn_0_35 );
nand g442 ( new_n580_, new_n262_, new_n259_, new_n579_, new_n264_ );
not g443 ( new_n581_, new_n580_ );
nand g444 ( new_n582_, new_n559_, new_n581_ );
not g445 ( new_n583_, new_n582_ );
nand g446 ( new_n584_, new_n583_, new_n404_ );
xnor g447 ( N748, new_n584_, N97 );
nand g448 ( new_n586_, new_n559_, new_n392_, new_n581_ );
xnor g449 ( new_n587_, new_n586_, keyIn_0_50 );
xnor g450 ( N749, new_n587_, N101 );
nand g451 ( new_n589_, new_n583_, new_n330_ );
xnor g452 ( N750, new_n589_, N105 );
nand g453 ( new_n591_, new_n583_, new_n383_ );
xnor g454 ( N751, new_n591_, N109 );
nand g455 ( new_n593_, new_n262_, new_n250_, new_n228_ );
not g456 ( new_n594_, new_n593_ );
nand g457 ( new_n595_, new_n559_, new_n404_, new_n594_ );
xnor g458 ( N752, new_n595_, N113 );
not g459 ( new_n597_, N117 );
nand g460 ( new_n598_, new_n559_, new_n392_, new_n594_ );
xnor g461 ( new_n599_, new_n598_, keyIn_0_51 );
xnor g462 ( N753, new_n599_, new_n597_ );
not g463 ( new_n601_, keyIn_0_62 );
nand g464 ( new_n602_, new_n521_, new_n525_, new_n330_, new_n594_ );
xnor g465 ( new_n603_, new_n602_, keyIn_0_52 );
nand g466 ( new_n604_, new_n603_, new_n168_ );
not g467 ( new_n605_, keyIn_0_52 );
xnor g468 ( new_n606_, new_n602_, new_n605_ );
nand g469 ( new_n607_, new_n606_, N121 );
nand g470 ( new_n608_, new_n604_, new_n607_ );
nand g471 ( new_n609_, new_n608_, new_n601_ );
nand g472 ( new_n610_, new_n604_, new_n607_, keyIn_0_62 );
nand g473 ( N754, new_n609_, new_n610_ );
not g474 ( new_n612_, keyIn_0_63 );
nand g475 ( new_n613_, new_n594_, new_n383_ );
not g476 ( new_n614_, new_n613_ );
nand g477 ( new_n615_, new_n521_, new_n525_, new_n614_ );
nand g478 ( new_n616_, new_n615_, keyIn_0_53 );
not g479 ( new_n617_, keyIn_0_53 );
nand g480 ( new_n618_, new_n559_, new_n617_, new_n614_ );
nand g481 ( new_n619_, new_n618_, new_n616_ );
nand g482 ( new_n620_, new_n619_, N125 );
nand g483 ( new_n621_, new_n618_, new_n169_, new_n616_ );
nand g484 ( new_n622_, new_n620_, new_n621_ );
nand g485 ( new_n623_, new_n622_, new_n612_ );
nand g486 ( new_n624_, new_n620_, keyIn_0_63, new_n621_ );
nand g487 ( N755, new_n623_, new_n624_ );
endmodule